// Benchmark "sqrt" written by ABC on Tue Sep  5 18:14:00 2023

module sqrt ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] ,
    \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] , \asqrt[5] ,
    \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] , \asqrt[10] ,
    \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] , \asqrt[15] ,
    \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] , \asqrt[20] ,
    \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] , \asqrt[25] ,
    \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] , \asqrt[30] ,
    \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] , \asqrt[35] ,
    \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] , \asqrt[40] ,
    \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] , \asqrt[45] ,
    \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] , \asqrt[50] ,
    \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] , \asqrt[55] ,
    \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] , \asqrt[60] ,
    \asqrt[61] , \asqrt[62] , \asqrt[63]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] ;
  output \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] ,
    \asqrt[5] , \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] ,
    \asqrt[10] , \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] ,
    \asqrt[15] , \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] ,
    \asqrt[20] , \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] ,
    \asqrt[25] , \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] ,
    \asqrt[30] , \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] ,
    \asqrt[35] , \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] ,
    \asqrt[40] , \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] ,
    \asqrt[45] , \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] ,
    \asqrt[50] , \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] ,
    \asqrt[55] , \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] ,
    \asqrt[60] , \asqrt[61] , \asqrt[62] , \asqrt[63] ;
  wire new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n201_, new_n202_, new_n203_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_,
    new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_,
    new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_,
    new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_,
    new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_,
    new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_,
    new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_,
    new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_,
    new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_,
    new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_,
    new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_,
    new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_,
    new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_,
    new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_,
    new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_,
    new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_,
    new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_,
    new_n3179_, new_n3180_, new_n3181_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_,
    new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_,
    new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_,
    new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_,
    new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_,
    new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_,
    new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_,
    new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_,
    new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_,
    new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_,
    new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_,
    new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_,
    new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_,
    new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_,
    new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_,
    new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_,
    new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_,
    new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_,
    new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_,
    new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_,
    new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_,
    new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_,
    new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_,
    new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_,
    new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_,
    new_n3667_, new_n3668_, new_n3669_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_,
    new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_,
    new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_,
    new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_,
    new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_,
    new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_,
    new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_,
    new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_,
    new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_,
    new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_,
    new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_,
    new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_,
    new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_,
    new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_,
    new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_,
    new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_,
    new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_,
    new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_,
    new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_,
    new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_,
    new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_,
    new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_,
    new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_,
    new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_,
    new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_,
    new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_,
    new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_,
    new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_,
    new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_,
    new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_,
    new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_,
    new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_,
    new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_,
    new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_,
    new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_,
    new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_,
    new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_,
    new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_,
    new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_,
    new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_,
    new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_,
    new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_,
    new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_,
    new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_,
    new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_,
    new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_,
    new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_,
    new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_,
    new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_,
    new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_,
    new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_,
    new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_,
    new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_,
    new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_,
    new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_,
    new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_,
    new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_,
    new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_,
    new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_,
    new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_,
    new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_,
    new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_,
    new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_,
    new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_,
    new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_,
    new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_,
    new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_,
    new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_,
    new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_,
    new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_,
    new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_,
    new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_,
    new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_,
    new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_,
    new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_,
    new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_,
    new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4450_,
    new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_,
    new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_,
    new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_,
    new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_,
    new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_,
    new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_,
    new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_,
    new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_,
    new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_,
    new_n4505_, new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_,
    new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_,
    new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_,
    new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_,
    new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_,
    new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_,
    new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_,
    new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_,
    new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_,
    new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_,
    new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_,
    new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_,
    new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_,
    new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_,
    new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_,
    new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_,
    new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_,
    new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_,
    new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_,
    new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_,
    new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_,
    new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_,
    new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_,
    new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_,
    new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_,
    new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_,
    new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_,
    new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_,
    new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_,
    new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_,
    new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_,
    new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5019_, new_n5020_, new_n5021_, new_n5022_,
    new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_,
    new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_,
    new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_,
    new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_,
    new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_,
    new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_,
    new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_,
    new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_,
    new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_,
    new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_,
    new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_,
    new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_,
    new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_,
    new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_,
    new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_,
    new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_,
    new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_,
    new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_,
    new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_,
    new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_,
    new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_,
    new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_,
    new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_,
    new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_,
    new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_,
    new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_,
    new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_,
    new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_,
    new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_,
    new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_,
    new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5623_, new_n5624_,
    new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_,
    new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_,
    new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_,
    new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_,
    new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_,
    new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_,
    new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_,
    new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_,
    new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_,
    new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_,
    new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_,
    new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_,
    new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_,
    new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_,
    new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_,
    new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_,
    new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_,
    new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_,
    new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_,
    new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_,
    new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_,
    new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_,
    new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_,
    new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_,
    new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_,
    new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_,
    new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_,
    new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_,
    new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_,
    new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_,
    new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_,
    new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_,
    new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_,
    new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_,
    new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_,
    new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_,
    new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_,
    new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_,
    new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_,
    new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_,
    new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_,
    new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_,
    new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_,
    new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_,
    new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_,
    new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_,
    new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5967_,
    new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_,
    new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_,
    new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_,
    new_n6256_, new_n6257_, new_n6258_, new_n6260_, new_n6261_, new_n6262_,
    new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_,
    new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_,
    new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_,
    new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_,
    new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_,
    new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_,
    new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_,
    new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_,
    new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_,
    new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_,
    new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_,
    new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_,
    new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_,
    new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_,
    new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_,
    new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_,
    new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_,
    new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_,
    new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_,
    new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_,
    new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_,
    new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_,
    new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_,
    new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_,
    new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_,
    new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_,
    new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_,
    new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_,
    new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_,
    new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_,
    new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_,
    new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_,
    new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_,
    new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_,
    new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_,
    new_n6599_, new_n6600_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_,
    new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_,
    new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_,
    new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_,
    new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_,
    new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_,
    new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_,
    new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_,
    new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_,
    new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_,
    new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_,
    new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_,
    new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_,
    new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_,
    new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_,
    new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_,
    new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_,
    new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_,
    new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_,
    new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_,
    new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_,
    new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_,
    new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_,
    new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_,
    new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_,
    new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_,
    new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_,
    new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_,
    new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_,
    new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_,
    new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_,
    new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_,
    new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_,
    new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_,
    new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_,
    new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_,
    new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_,
    new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_,
    new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_,
    new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_,
    new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_,
    new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_,
    new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_,
    new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_,
    new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_,
    new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_,
    new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_,
    new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_,
    new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_,
    new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_,
    new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_,
    new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_,
    new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_,
    new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_,
    new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_,
    new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_,
    new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_,
    new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_,
    new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_,
    new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_,
    new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_,
    new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_,
    new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_,
    new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_,
    new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_,
    new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_,
    new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_,
    new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_,
    new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_,
    new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_,
    new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_,
    new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_,
    new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_,
    new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_,
    new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_,
    new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_,
    new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_,
    new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_,
    new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_,
    new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_,
    new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_,
    new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_,
    new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_,
    new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_,
    new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_,
    new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_,
    new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_,
    new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_,
    new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_,
    new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_,
    new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_,
    new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_,
    new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_,
    new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_,
    new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_,
    new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_,
    new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_,
    new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_,
    new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_,
    new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_,
    new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_,
    new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_,
    new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_,
    new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_,
    new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_,
    new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_,
    new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_,
    new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_,
    new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_,
    new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_,
    new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_,
    new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_,
    new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_,
    new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_,
    new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_,
    new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_,
    new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_,
    new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_,
    new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_,
    new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_,
    new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_,
    new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_,
    new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_,
    new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_,
    new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_,
    new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_,
    new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_,
    new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_,
    new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_,
    new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_,
    new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_,
    new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_,
    new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_,
    new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_,
    new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_,
    new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_,
    new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_,
    new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_,
    new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_,
    new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_,
    new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_,
    new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_,
    new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_,
    new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_,
    new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_,
    new_n8380_, new_n8381_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_,
    new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_,
    new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_,
    new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_,
    new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_,
    new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_,
    new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_,
    new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_,
    new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_,
    new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_,
    new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_,
    new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_,
    new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_,
    new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_,
    new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_,
    new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_,
    new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_,
    new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_,
    new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_,
    new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_,
    new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_,
    new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_,
    new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_,
    new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_,
    new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_,
    new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_,
    new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_,
    new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_,
    new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_,
    new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_,
    new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_,
    new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_,
    new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_,
    new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_,
    new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_,
    new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_,
    new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_,
    new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_,
    new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_,
    new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_,
    new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_,
    new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_,
    new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_,
    new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_,
    new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_,
    new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_,
    new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_,
    new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_,
    new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_,
    new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_,
    new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_,
    new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_,
    new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_,
    new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_,
    new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_,
    new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_,
    new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_,
    new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_,
    new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_,
    new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_,
    new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_,
    new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_,
    new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_,
    new_n9156_, new_n9157_, new_n9159_, new_n9160_, new_n9161_, new_n9162_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_,
    new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_,
    new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_,
    new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_,
    new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_,
    new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_,
    new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_,
    new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_,
    new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_,
    new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_,
    new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_,
    new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_,
    new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_,
    new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_,
    new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_,
    new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_,
    new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_,
    new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_,
    new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_,
    new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_,
    new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_,
    new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_,
    new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_,
    new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_,
    new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_,
    new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_,
    new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_,
    new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_,
    new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_,
    new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_,
    new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_,
    new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_,
    new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_,
    new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_,
    new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_,
    new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_,
    new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_,
    new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_,
    new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_,
    new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_,
    new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_,
    new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_,
    new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_,
    new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_,
    new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_,
    new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_,
    new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_,
    new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_,
    new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_,
    new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_,
    new_n9571_, new_n9572_, new_n9574_, new_n9575_, new_n9576_, new_n9577_,
    new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_,
    new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_,
    new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_,
    new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_,
    new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_,
    new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_,
    new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_,
    new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_,
    new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_,
    new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_,
    new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_,
    new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9971_, new_n9972_, new_n9973_, new_n9974_,
    new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_,
    new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_,
    new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_,
    new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_,
    new_n9999_, new_n10000_, new_n10001_, new_n10002_, new_n10003_,
    new_n10004_, new_n10005_, new_n10006_, new_n10007_, new_n10008_,
    new_n10009_, new_n10010_, new_n10011_, new_n10012_, new_n10013_,
    new_n10014_, new_n10015_, new_n10016_, new_n10017_, new_n10018_,
    new_n10019_, new_n10020_, new_n10021_, new_n10022_, new_n10023_,
    new_n10024_, new_n10025_, new_n10026_, new_n10027_, new_n10028_,
    new_n10029_, new_n10030_, new_n10031_, new_n10032_, new_n10033_,
    new_n10034_, new_n10035_, new_n10036_, new_n10037_, new_n10038_,
    new_n10039_, new_n10040_, new_n10041_, new_n10042_, new_n10043_,
    new_n10044_, new_n10045_, new_n10046_, new_n10047_, new_n10048_,
    new_n10049_, new_n10050_, new_n10051_, new_n10052_, new_n10053_,
    new_n10054_, new_n10055_, new_n10056_, new_n10057_, new_n10058_,
    new_n10059_, new_n10060_, new_n10061_, new_n10062_, new_n10063_,
    new_n10064_, new_n10065_, new_n10066_, new_n10067_, new_n10068_,
    new_n10069_, new_n10070_, new_n10071_, new_n10072_, new_n10073_,
    new_n10074_, new_n10075_, new_n10076_, new_n10077_, new_n10078_,
    new_n10079_, new_n10080_, new_n10081_, new_n10082_, new_n10083_,
    new_n10084_, new_n10085_, new_n10086_, new_n10087_, new_n10088_,
    new_n10089_, new_n10090_, new_n10091_, new_n10092_, new_n10093_,
    new_n10094_, new_n10095_, new_n10096_, new_n10097_, new_n10098_,
    new_n10099_, new_n10100_, new_n10101_, new_n10102_, new_n10103_,
    new_n10104_, new_n10105_, new_n10106_, new_n10107_, new_n10108_,
    new_n10109_, new_n10110_, new_n10111_, new_n10112_, new_n10113_,
    new_n10114_, new_n10115_, new_n10116_, new_n10117_, new_n10118_,
    new_n10119_, new_n10120_, new_n10121_, new_n10122_, new_n10123_,
    new_n10124_, new_n10125_, new_n10126_, new_n10127_, new_n10128_,
    new_n10129_, new_n10130_, new_n10131_, new_n10132_, new_n10133_,
    new_n10134_, new_n10135_, new_n10136_, new_n10137_, new_n10138_,
    new_n10139_, new_n10140_, new_n10141_, new_n10142_, new_n10143_,
    new_n10144_, new_n10145_, new_n10146_, new_n10147_, new_n10148_,
    new_n10149_, new_n10150_, new_n10151_, new_n10152_, new_n10153_,
    new_n10154_, new_n10155_, new_n10156_, new_n10157_, new_n10158_,
    new_n10159_, new_n10160_, new_n10161_, new_n10162_, new_n10163_,
    new_n10164_, new_n10165_, new_n10166_, new_n10167_, new_n10168_,
    new_n10169_, new_n10170_, new_n10171_, new_n10172_, new_n10173_,
    new_n10174_, new_n10175_, new_n10176_, new_n10177_, new_n10178_,
    new_n10179_, new_n10180_, new_n10181_, new_n10182_, new_n10183_,
    new_n10184_, new_n10185_, new_n10186_, new_n10187_, new_n10188_,
    new_n10189_, new_n10190_, new_n10191_, new_n10192_, new_n10193_,
    new_n10194_, new_n10195_, new_n10196_, new_n10197_, new_n10198_,
    new_n10199_, new_n10200_, new_n10201_, new_n10202_, new_n10203_,
    new_n10204_, new_n10205_, new_n10206_, new_n10207_, new_n10208_,
    new_n10209_, new_n10210_, new_n10211_, new_n10212_, new_n10213_,
    new_n10214_, new_n10215_, new_n10216_, new_n10217_, new_n10218_,
    new_n10219_, new_n10220_, new_n10221_, new_n10222_, new_n10223_,
    new_n10224_, new_n10225_, new_n10226_, new_n10227_, new_n10228_,
    new_n10229_, new_n10230_, new_n10231_, new_n10232_, new_n10233_,
    new_n10234_, new_n10235_, new_n10236_, new_n10237_, new_n10238_,
    new_n10239_, new_n10240_, new_n10241_, new_n10242_, new_n10243_,
    new_n10244_, new_n10245_, new_n10246_, new_n10247_, new_n10248_,
    new_n10249_, new_n10250_, new_n10251_, new_n10252_, new_n10253_,
    new_n10254_, new_n10255_, new_n10256_, new_n10257_, new_n10258_,
    new_n10259_, new_n10260_, new_n10261_, new_n10262_, new_n10263_,
    new_n10264_, new_n10265_, new_n10266_, new_n10267_, new_n10268_,
    new_n10269_, new_n10270_, new_n10271_, new_n10272_, new_n10273_,
    new_n10274_, new_n10275_, new_n10276_, new_n10277_, new_n10278_,
    new_n10279_, new_n10280_, new_n10281_, new_n10282_, new_n10283_,
    new_n10284_, new_n10285_, new_n10286_, new_n10287_, new_n10288_,
    new_n10289_, new_n10290_, new_n10291_, new_n10292_, new_n10293_,
    new_n10294_, new_n10295_, new_n10296_, new_n10297_, new_n10298_,
    new_n10299_, new_n10300_, new_n10301_, new_n10302_, new_n10303_,
    new_n10304_, new_n10305_, new_n10306_, new_n10307_, new_n10308_,
    new_n10309_, new_n10310_, new_n10311_, new_n10312_, new_n10313_,
    new_n10314_, new_n10315_, new_n10316_, new_n10317_, new_n10318_,
    new_n10319_, new_n10320_, new_n10321_, new_n10322_, new_n10323_,
    new_n10324_, new_n10325_, new_n10326_, new_n10327_, new_n10328_,
    new_n10329_, new_n10330_, new_n10331_, new_n10332_, new_n10333_,
    new_n10334_, new_n10335_, new_n10336_, new_n10337_, new_n10338_,
    new_n10339_, new_n10340_, new_n10341_, new_n10342_, new_n10343_,
    new_n10344_, new_n10345_, new_n10346_, new_n10347_, new_n10348_,
    new_n10349_, new_n10350_, new_n10351_, new_n10352_, new_n10353_,
    new_n10354_, new_n10355_, new_n10356_, new_n10357_, new_n10358_,
    new_n10359_, new_n10360_, new_n10361_, new_n10362_, new_n10363_,
    new_n10364_, new_n10365_, new_n10366_, new_n10367_, new_n10368_,
    new_n10369_, new_n10370_, new_n10371_, new_n10372_, new_n10373_,
    new_n10374_, new_n10375_, new_n10376_, new_n10377_, new_n10378_,
    new_n10379_, new_n10380_, new_n10381_, new_n10382_, new_n10383_,
    new_n10384_, new_n10385_, new_n10386_, new_n10387_, new_n10388_,
    new_n10389_, new_n10390_, new_n10391_, new_n10392_, new_n10393_,
    new_n10394_, new_n10395_, new_n10396_, new_n10397_, new_n10398_,
    new_n10399_, new_n10400_, new_n10401_, new_n10402_, new_n10403_,
    new_n10404_, new_n10405_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10439_,
    new_n10440_, new_n10441_, new_n10442_, new_n10443_, new_n10444_,
    new_n10445_, new_n10446_, new_n10447_, new_n10448_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10453_, new_n10454_,
    new_n10455_, new_n10456_, new_n10457_, new_n10458_, new_n10459_,
    new_n10460_, new_n10461_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11299_, new_n11300_, new_n11301_,
    new_n11302_, new_n11303_, new_n11304_, new_n11305_, new_n11306_,
    new_n11307_, new_n11308_, new_n11309_, new_n11310_, new_n11311_,
    new_n11312_, new_n11313_, new_n11314_, new_n11315_, new_n11316_,
    new_n11317_, new_n11318_, new_n11319_, new_n11320_, new_n11321_,
    new_n11322_, new_n11323_, new_n11324_, new_n11325_, new_n11326_,
    new_n11327_, new_n11328_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11340_, new_n11341_,
    new_n11342_, new_n11343_, new_n11344_, new_n11345_, new_n11346_,
    new_n11347_, new_n11348_, new_n11349_, new_n11350_, new_n11351_,
    new_n11352_, new_n11353_, new_n11354_, new_n11355_, new_n11356_,
    new_n11357_, new_n11358_, new_n11359_, new_n11360_, new_n11361_,
    new_n11362_, new_n11363_, new_n11364_, new_n11365_, new_n11366_,
    new_n11367_, new_n11368_, new_n11369_, new_n11370_, new_n11371_,
    new_n11372_, new_n11373_, new_n11374_, new_n11375_, new_n11376_,
    new_n11377_, new_n11378_, new_n11379_, new_n11380_, new_n11381_,
    new_n11382_, new_n11383_, new_n11384_, new_n11385_, new_n11386_,
    new_n11387_, new_n11388_, new_n11389_, new_n11390_, new_n11391_,
    new_n11392_, new_n11393_, new_n11394_, new_n11395_, new_n11396_,
    new_n11397_, new_n11398_, new_n11399_, new_n11400_, new_n11401_,
    new_n11402_, new_n11403_, new_n11404_, new_n11405_, new_n11406_,
    new_n11407_, new_n11408_, new_n11409_, new_n11410_, new_n11411_,
    new_n11412_, new_n11413_, new_n11414_, new_n11415_, new_n11416_,
    new_n11417_, new_n11418_, new_n11419_, new_n11420_, new_n11421_,
    new_n11422_, new_n11423_, new_n11424_, new_n11425_, new_n11426_,
    new_n11427_, new_n11428_, new_n11429_, new_n11430_, new_n11431_,
    new_n11432_, new_n11433_, new_n11434_, new_n11435_, new_n11436_,
    new_n11437_, new_n11438_, new_n11439_, new_n11440_, new_n11441_,
    new_n11442_, new_n11443_, new_n11444_, new_n11445_, new_n11446_,
    new_n11447_, new_n11448_, new_n11449_, new_n11450_, new_n11451_,
    new_n11452_, new_n11453_, new_n11454_, new_n11455_, new_n11456_,
    new_n11457_, new_n11458_, new_n11459_, new_n11460_, new_n11461_,
    new_n11462_, new_n11463_, new_n11464_, new_n11465_, new_n11466_,
    new_n11467_, new_n11468_, new_n11469_, new_n11470_, new_n11471_,
    new_n11472_, new_n11473_, new_n11474_, new_n11475_, new_n11476_,
    new_n11477_, new_n11478_, new_n11479_, new_n11480_, new_n11481_,
    new_n11482_, new_n11483_, new_n11484_, new_n11485_, new_n11486_,
    new_n11487_, new_n11488_, new_n11489_, new_n11490_, new_n11491_,
    new_n11492_, new_n11493_, new_n11494_, new_n11495_, new_n11496_,
    new_n11497_, new_n11498_, new_n11499_, new_n11500_, new_n11501_,
    new_n11502_, new_n11503_, new_n11504_, new_n11505_, new_n11506_,
    new_n11507_, new_n11508_, new_n11509_, new_n11510_, new_n11511_,
    new_n11512_, new_n11513_, new_n11514_, new_n11515_, new_n11516_,
    new_n11517_, new_n11518_, new_n11519_, new_n11520_, new_n11521_,
    new_n11522_, new_n11523_, new_n11524_, new_n11525_, new_n11526_,
    new_n11527_, new_n11528_, new_n11529_, new_n11530_, new_n11531_,
    new_n11532_, new_n11533_, new_n11534_, new_n11535_, new_n11536_,
    new_n11537_, new_n11538_, new_n11539_, new_n11540_, new_n11541_,
    new_n11542_, new_n11543_, new_n11544_, new_n11545_, new_n11546_,
    new_n11547_, new_n11548_, new_n11549_, new_n11550_, new_n11551_,
    new_n11552_, new_n11553_, new_n11554_, new_n11555_, new_n11556_,
    new_n11557_, new_n11558_, new_n11559_, new_n11560_, new_n11561_,
    new_n11562_, new_n11563_, new_n11564_, new_n11565_, new_n11566_,
    new_n11567_, new_n11568_, new_n11569_, new_n11570_, new_n11571_,
    new_n11572_, new_n11573_, new_n11574_, new_n11575_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11740_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11748_, new_n11749_, new_n11750_, new_n11751_, new_n11752_,
    new_n11753_, new_n11754_, new_n11755_, new_n11756_, new_n11757_,
    new_n11758_, new_n11759_, new_n11760_, new_n11761_, new_n11762_,
    new_n11763_, new_n11764_, new_n11765_, new_n11766_, new_n11767_,
    new_n11768_, new_n11769_, new_n11770_, new_n11771_, new_n11772_,
    new_n11773_, new_n11774_, new_n11775_, new_n11776_, new_n11777_,
    new_n11778_, new_n11779_, new_n11780_, new_n11781_, new_n11782_,
    new_n11783_, new_n11784_, new_n11785_, new_n11786_, new_n11787_,
    new_n11788_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11813_, new_n11814_, new_n11815_, new_n11816_, new_n11817_,
    new_n11818_, new_n11819_, new_n11820_, new_n11821_, new_n11822_,
    new_n11823_, new_n11824_, new_n11825_, new_n11826_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11844_, new_n11845_, new_n11846_, new_n11847_,
    new_n11848_, new_n11849_, new_n11850_, new_n11851_, new_n11852_,
    new_n11853_, new_n11854_, new_n11855_, new_n11856_, new_n11857_,
    new_n11858_, new_n11859_, new_n11860_, new_n11861_, new_n11862_,
    new_n11863_, new_n11864_, new_n11865_, new_n11866_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11873_, new_n11874_, new_n11875_, new_n11876_, new_n11877_,
    new_n11878_, new_n11879_, new_n11880_, new_n11881_, new_n11882_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11925_, new_n11926_, new_n11927_,
    new_n11928_, new_n11929_, new_n11930_, new_n11931_, new_n11932_,
    new_n11933_, new_n11934_, new_n11935_, new_n11936_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11943_, new_n11944_, new_n11945_, new_n11946_, new_n11947_,
    new_n11948_, new_n11949_, new_n11950_, new_n11951_, new_n11952_,
    new_n11953_, new_n11954_, new_n11955_, new_n11956_, new_n11957_,
    new_n11958_, new_n11959_, new_n11960_, new_n11961_, new_n11962_,
    new_n11963_, new_n11964_, new_n11965_, new_n11966_, new_n11967_,
    new_n11968_, new_n11969_, new_n11970_, new_n11971_, new_n11972_,
    new_n11973_, new_n11974_, new_n11975_, new_n11976_, new_n11977_,
    new_n11978_, new_n11979_, new_n11980_, new_n11981_, new_n11982_,
    new_n11983_, new_n11984_, new_n11985_, new_n11986_, new_n11987_,
    new_n11988_, new_n11989_, new_n11990_, new_n11991_, new_n11992_,
    new_n11993_, new_n11994_, new_n11995_, new_n11996_, new_n11997_,
    new_n11998_, new_n11999_, new_n12000_, new_n12001_, new_n12002_,
    new_n12003_, new_n12004_, new_n12005_, new_n12006_, new_n12007_,
    new_n12008_, new_n12009_, new_n12010_, new_n12011_, new_n12012_,
    new_n12013_, new_n12014_, new_n12015_, new_n12016_, new_n12017_,
    new_n12018_, new_n12019_, new_n12020_, new_n12021_, new_n12022_,
    new_n12023_, new_n12024_, new_n12025_, new_n12026_, new_n12027_,
    new_n12028_, new_n12029_, new_n12030_, new_n12031_, new_n12032_,
    new_n12033_, new_n12034_, new_n12035_, new_n12036_, new_n12037_,
    new_n12038_, new_n12039_, new_n12040_, new_n12041_, new_n12042_,
    new_n12043_, new_n12044_, new_n12045_, new_n12046_, new_n12047_,
    new_n12048_, new_n12049_, new_n12050_, new_n12051_, new_n12052_,
    new_n12053_, new_n12054_, new_n12055_, new_n12056_, new_n12057_,
    new_n12058_, new_n12059_, new_n12060_, new_n12061_, new_n12062_,
    new_n12063_, new_n12064_, new_n12065_, new_n12066_, new_n12067_,
    new_n12068_, new_n12069_, new_n12070_, new_n12071_, new_n12072_,
    new_n12073_, new_n12074_, new_n12075_, new_n12076_, new_n12077_,
    new_n12078_, new_n12079_, new_n12080_, new_n12081_, new_n12082_,
    new_n12083_, new_n12084_, new_n12085_, new_n12086_, new_n12087_,
    new_n12088_, new_n12089_, new_n12090_, new_n12091_, new_n12092_,
    new_n12093_, new_n12094_, new_n12095_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12100_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12106_, new_n12107_,
    new_n12108_, new_n12109_, new_n12110_, new_n12111_, new_n12112_,
    new_n12113_, new_n12114_, new_n12115_, new_n12116_, new_n12117_,
    new_n12118_, new_n12119_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12148_, new_n12149_, new_n12150_, new_n12151_, new_n12152_,
    new_n12153_, new_n12154_, new_n12155_, new_n12156_, new_n12157_,
    new_n12158_, new_n12159_, new_n12160_, new_n12161_, new_n12162_,
    new_n12163_, new_n12164_, new_n12165_, new_n12166_, new_n12167_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12173_,
    new_n12174_, new_n12175_, new_n12176_, new_n12177_, new_n12178_,
    new_n12179_, new_n12180_, new_n12181_, new_n12182_, new_n12183_,
    new_n12184_, new_n12185_, new_n12186_, new_n12187_, new_n12188_,
    new_n12189_, new_n12190_, new_n12191_, new_n12192_, new_n12193_,
    new_n12194_, new_n12195_, new_n12196_, new_n12197_, new_n12198_,
    new_n12199_, new_n12200_, new_n12201_, new_n12202_, new_n12203_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12254_, new_n12255_, new_n12256_, new_n12257_, new_n12258_,
    new_n12259_, new_n12260_, new_n12261_, new_n12262_, new_n12263_,
    new_n12264_, new_n12265_, new_n12266_, new_n12267_, new_n12268_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12280_, new_n12281_, new_n12282_, new_n12283_,
    new_n12284_, new_n12285_, new_n12286_, new_n12287_, new_n12288_,
    new_n12289_, new_n12290_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12296_, new_n12297_, new_n12298_,
    new_n12299_, new_n12300_, new_n12301_, new_n12302_, new_n12303_,
    new_n12304_, new_n12305_, new_n12306_, new_n12307_, new_n12308_,
    new_n12309_, new_n12310_, new_n12311_, new_n12312_, new_n12313_,
    new_n12314_, new_n12315_, new_n12316_, new_n12317_, new_n12318_,
    new_n12319_, new_n12320_, new_n12321_, new_n12322_, new_n12323_,
    new_n12324_, new_n12325_, new_n12326_, new_n12327_, new_n12328_,
    new_n12329_, new_n12330_, new_n12331_, new_n12332_, new_n12333_,
    new_n12334_, new_n12335_, new_n12336_, new_n12337_, new_n12338_,
    new_n12339_, new_n12340_, new_n12341_, new_n12342_, new_n12343_,
    new_n12344_, new_n12345_, new_n12346_, new_n12347_, new_n12348_,
    new_n12349_, new_n12350_, new_n12351_, new_n12352_, new_n12353_,
    new_n12354_, new_n12355_, new_n12356_, new_n12357_, new_n12358_,
    new_n12359_, new_n12360_, new_n12361_, new_n12362_, new_n12363_,
    new_n12364_, new_n12365_, new_n12366_, new_n12367_, new_n12368_,
    new_n12369_, new_n12370_, new_n12371_, new_n12372_, new_n12373_,
    new_n12374_, new_n12375_, new_n12376_, new_n12377_, new_n12378_,
    new_n12379_, new_n12380_, new_n12381_, new_n12382_, new_n12383_,
    new_n12384_, new_n12385_, new_n12386_, new_n12387_, new_n12388_,
    new_n12389_, new_n12390_, new_n12391_, new_n12392_, new_n12393_,
    new_n12394_, new_n12395_, new_n12396_, new_n12397_, new_n12398_,
    new_n12399_, new_n12400_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12405_, new_n12406_, new_n12407_, new_n12408_,
    new_n12409_, new_n12410_, new_n12411_, new_n12412_, new_n12413_,
    new_n12414_, new_n12415_, new_n12416_, new_n12417_, new_n12418_,
    new_n12419_, new_n12420_, new_n12421_, new_n12422_, new_n12423_,
    new_n12424_, new_n12425_, new_n12426_, new_n12427_, new_n12428_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12458_,
    new_n12459_, new_n12460_, new_n12461_, new_n12462_, new_n12463_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12470_, new_n12471_, new_n12472_, new_n12473_,
    new_n12474_, new_n12475_, new_n12476_, new_n12477_, new_n12478_,
    new_n12479_, new_n12480_, new_n12481_, new_n12482_, new_n12483_,
    new_n12484_, new_n12485_, new_n12486_, new_n12487_, new_n12488_,
    new_n12489_, new_n12490_, new_n12491_, new_n12492_, new_n12493_,
    new_n12494_, new_n12495_, new_n12496_, new_n12497_, new_n12498_,
    new_n12499_, new_n12500_, new_n12501_, new_n12502_, new_n12503_,
    new_n12504_, new_n12505_, new_n12506_, new_n12507_, new_n12508_,
    new_n12509_, new_n12510_, new_n12511_, new_n12512_, new_n12513_,
    new_n12514_, new_n12515_, new_n12516_, new_n12517_, new_n12518_,
    new_n12519_, new_n12520_, new_n12521_, new_n12522_, new_n12523_,
    new_n12524_, new_n12525_, new_n12526_, new_n12527_, new_n12528_,
    new_n12529_, new_n12530_, new_n12531_, new_n12532_, new_n12533_,
    new_n12534_, new_n12535_, new_n12536_, new_n12537_, new_n12538_,
    new_n12539_, new_n12540_, new_n12541_, new_n12542_, new_n12543_,
    new_n12544_, new_n12545_, new_n12546_, new_n12547_, new_n12548_,
    new_n12549_, new_n12550_, new_n12551_, new_n12552_, new_n12553_,
    new_n12554_, new_n12555_, new_n12556_, new_n12557_, new_n12558_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12566_, new_n12567_, new_n12568_,
    new_n12569_, new_n12570_, new_n12571_, new_n12572_, new_n12573_,
    new_n12574_, new_n12575_, new_n12576_, new_n12577_, new_n12578_,
    new_n12579_, new_n12580_, new_n12581_, new_n12582_, new_n12583_,
    new_n12584_, new_n12585_, new_n12586_, new_n12587_, new_n12588_,
    new_n12589_, new_n12590_, new_n12591_, new_n12592_, new_n12593_,
    new_n12594_, new_n12595_, new_n12596_, new_n12597_, new_n12598_,
    new_n12599_, new_n12600_, new_n12601_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12608_,
    new_n12609_, new_n12611_, new_n12612_, new_n12613_, new_n12614_,
    new_n12615_, new_n12616_, new_n12617_, new_n12618_, new_n12619_,
    new_n12620_, new_n12621_, new_n12622_, new_n12623_, new_n12624_,
    new_n12625_, new_n12626_, new_n12627_, new_n12628_, new_n12629_,
    new_n12630_, new_n12631_, new_n12632_, new_n12633_, new_n12634_,
    new_n12635_, new_n12636_, new_n12637_, new_n12638_, new_n12639_,
    new_n12640_, new_n12641_, new_n12642_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12649_,
    new_n12650_, new_n12651_, new_n12652_, new_n12653_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12663_, new_n12664_,
    new_n12665_, new_n12666_, new_n12667_, new_n12668_, new_n12669_,
    new_n12670_, new_n12671_, new_n12672_, new_n12673_, new_n12674_,
    new_n12675_, new_n12676_, new_n12677_, new_n12678_, new_n12679_,
    new_n12680_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12687_, new_n12688_, new_n12689_,
    new_n12690_, new_n12691_, new_n12692_, new_n12693_, new_n12694_,
    new_n12695_, new_n12696_, new_n12697_, new_n12698_, new_n12699_,
    new_n12700_, new_n12701_, new_n12702_, new_n12703_, new_n12704_,
    new_n12705_, new_n12706_, new_n12707_, new_n12708_, new_n12709_,
    new_n12710_, new_n12711_, new_n12712_, new_n12713_, new_n12714_,
    new_n12715_, new_n12716_, new_n12717_, new_n12718_, new_n12719_,
    new_n12720_, new_n12721_, new_n12722_, new_n12723_, new_n12724_,
    new_n12725_, new_n12726_, new_n12727_, new_n12728_, new_n12729_,
    new_n12730_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13089_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13096_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14069_, new_n14070_, new_n14071_, new_n14072_,
    new_n14073_, new_n14074_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14122_,
    new_n14123_, new_n14124_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14156_, new_n14157_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14170_, new_n14171_, new_n14172_,
    new_n14173_, new_n14174_, new_n14175_, new_n14176_, new_n14177_,
    new_n14178_, new_n14179_, new_n14180_, new_n14181_, new_n14182_,
    new_n14183_, new_n14184_, new_n14185_, new_n14186_, new_n14187_,
    new_n14188_, new_n14189_, new_n14190_, new_n14191_, new_n14192_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14206_, new_n14207_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14217_,
    new_n14218_, new_n14219_, new_n14220_, new_n14221_, new_n14222_,
    new_n14223_, new_n14224_, new_n14225_, new_n14226_, new_n14227_,
    new_n14228_, new_n14229_, new_n14230_, new_n14231_, new_n14232_,
    new_n14233_, new_n14234_, new_n14235_, new_n14236_, new_n14237_,
    new_n14238_, new_n14239_, new_n14240_, new_n14241_, new_n14242_,
    new_n14243_, new_n14244_, new_n14245_, new_n14246_, new_n14247_,
    new_n14248_, new_n14249_, new_n14250_, new_n14251_, new_n14252_,
    new_n14253_, new_n14254_, new_n14255_, new_n14256_, new_n14257_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14302_,
    new_n14303_, new_n14304_, new_n14305_, new_n14306_, new_n14307_,
    new_n14308_, new_n14309_, new_n14310_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14317_,
    new_n14318_, new_n14319_, new_n14320_, new_n14321_, new_n14322_,
    new_n14323_, new_n14324_, new_n14325_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14332_,
    new_n14333_, new_n14334_, new_n14335_, new_n14336_, new_n14337_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14344_, new_n14345_, new_n14346_, new_n14347_,
    new_n14348_, new_n14349_, new_n14350_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14355_, new_n14356_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14362_,
    new_n14363_, new_n14364_, new_n14365_, new_n14366_, new_n14367_,
    new_n14368_, new_n14369_, new_n14370_, new_n14371_, new_n14372_,
    new_n14373_, new_n14374_, new_n14375_, new_n14376_, new_n14377_,
    new_n14378_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14386_, new_n14387_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14393_, new_n14394_, new_n14395_, new_n14396_, new_n14397_,
    new_n14398_, new_n14399_, new_n14400_, new_n14401_, new_n14402_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14409_, new_n14410_, new_n14411_, new_n14412_,
    new_n14413_, new_n14414_, new_n14415_, new_n14416_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14422_,
    new_n14423_, new_n14424_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14544_, new_n14545_, new_n14546_, new_n14547_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14589_, new_n14590_, new_n14591_, new_n14592_, new_n14593_,
    new_n14594_, new_n14595_, new_n14596_, new_n14597_, new_n14598_,
    new_n14599_, new_n14600_, new_n14601_, new_n14602_, new_n14603_,
    new_n14604_, new_n14605_, new_n14606_, new_n14607_, new_n14608_,
    new_n14609_, new_n14610_, new_n14611_, new_n14612_, new_n14613_,
    new_n14614_, new_n14615_, new_n14616_, new_n14617_, new_n14618_,
    new_n14619_, new_n14620_, new_n14621_, new_n14622_, new_n14623_,
    new_n14624_, new_n14625_, new_n14626_, new_n14627_, new_n14628_,
    new_n14629_, new_n14630_, new_n14631_, new_n14632_, new_n14633_,
    new_n14634_, new_n14635_, new_n14636_, new_n14637_, new_n14638_,
    new_n14639_, new_n14640_, new_n14641_, new_n14642_, new_n14643_,
    new_n14644_, new_n14645_, new_n14646_, new_n14647_, new_n14648_,
    new_n14649_, new_n14650_, new_n14651_, new_n14652_, new_n14653_,
    new_n14654_, new_n14655_, new_n14656_, new_n14657_, new_n14658_,
    new_n14659_, new_n14660_, new_n14661_, new_n14662_, new_n14663_,
    new_n14664_, new_n14665_, new_n14666_, new_n14667_, new_n14668_,
    new_n14669_, new_n14670_, new_n14671_, new_n14672_, new_n14673_,
    new_n14674_, new_n14675_, new_n14676_, new_n14677_, new_n14678_,
    new_n14679_, new_n14680_, new_n14681_, new_n14682_, new_n14683_,
    new_n14684_, new_n14685_, new_n14686_, new_n14687_, new_n14688_,
    new_n14689_, new_n14690_, new_n14691_, new_n14692_, new_n14693_,
    new_n14694_, new_n14695_, new_n14696_, new_n14697_, new_n14698_,
    new_n14699_, new_n14700_, new_n14701_, new_n14702_, new_n14703_,
    new_n14704_, new_n14705_, new_n14706_, new_n14707_, new_n14708_,
    new_n14709_, new_n14710_, new_n14711_, new_n14712_, new_n14713_,
    new_n14714_, new_n14715_, new_n14716_, new_n14717_, new_n14718_,
    new_n14719_, new_n14720_, new_n14721_, new_n14722_, new_n14723_,
    new_n14724_, new_n14725_, new_n14726_, new_n14727_, new_n14728_,
    new_n14729_, new_n14730_, new_n14731_, new_n14732_, new_n14733_,
    new_n14734_, new_n14735_, new_n14736_, new_n14737_, new_n14738_,
    new_n14739_, new_n14740_, new_n14741_, new_n14742_, new_n14743_,
    new_n14744_, new_n14745_, new_n14746_, new_n14747_, new_n14748_,
    new_n14749_, new_n14750_, new_n14751_, new_n14752_, new_n14753_,
    new_n14754_, new_n14755_, new_n14756_, new_n14757_, new_n14758_,
    new_n14759_, new_n14760_, new_n14761_, new_n14762_, new_n14763_,
    new_n14764_, new_n14765_, new_n14766_, new_n14767_, new_n14768_,
    new_n14769_, new_n14770_, new_n14771_, new_n14772_, new_n14773_,
    new_n14774_, new_n14775_, new_n14776_, new_n14777_, new_n14778_,
    new_n14779_, new_n14780_, new_n14781_, new_n14782_, new_n14783_,
    new_n14784_, new_n14785_, new_n14786_, new_n14787_, new_n14788_,
    new_n14789_, new_n14790_, new_n14791_, new_n14792_, new_n14793_,
    new_n14794_, new_n14795_, new_n14796_, new_n14797_, new_n14798_,
    new_n14799_, new_n14800_, new_n14801_, new_n14802_, new_n14803_,
    new_n14804_, new_n14805_, new_n14806_, new_n14807_, new_n14808_,
    new_n14809_, new_n14810_, new_n14811_, new_n14812_, new_n14813_,
    new_n14814_, new_n14815_, new_n14816_, new_n14817_, new_n14818_,
    new_n14819_, new_n14820_, new_n14821_, new_n14822_, new_n14823_,
    new_n14824_, new_n14825_, new_n14826_, new_n14827_, new_n14828_,
    new_n14829_, new_n14830_, new_n14831_, new_n14832_, new_n14833_,
    new_n14834_, new_n14835_, new_n14836_, new_n14837_, new_n14838_,
    new_n14839_, new_n14840_, new_n14841_, new_n14842_, new_n14843_,
    new_n14844_, new_n14845_, new_n14846_, new_n14847_, new_n14848_,
    new_n14849_, new_n14850_, new_n14851_, new_n14852_, new_n14853_,
    new_n14854_, new_n14855_, new_n14856_, new_n14857_, new_n14858_,
    new_n14859_, new_n14860_, new_n14861_, new_n14862_, new_n14863_,
    new_n14864_, new_n14865_, new_n14866_, new_n14867_, new_n14868_,
    new_n14869_, new_n14870_, new_n14871_, new_n14872_, new_n14873_,
    new_n14874_, new_n14875_, new_n14876_, new_n14877_, new_n14878_,
    new_n14879_, new_n14880_, new_n14881_, new_n14882_, new_n14883_,
    new_n14884_, new_n14885_, new_n14886_, new_n14887_, new_n14888_,
    new_n14889_, new_n14890_, new_n14891_, new_n14892_, new_n14893_,
    new_n14894_, new_n14895_, new_n14896_, new_n14897_, new_n14898_,
    new_n14899_, new_n14900_, new_n14901_, new_n14902_, new_n14903_,
    new_n14904_, new_n14905_, new_n14906_, new_n14907_, new_n14908_,
    new_n14909_, new_n14910_, new_n14911_, new_n14912_, new_n14913_,
    new_n14914_, new_n14915_, new_n14916_, new_n14917_, new_n14918_,
    new_n14919_, new_n14920_, new_n14921_, new_n14922_, new_n14923_,
    new_n14924_, new_n14925_, new_n14926_, new_n14927_, new_n14928_,
    new_n14929_, new_n14930_, new_n14931_, new_n14932_, new_n14933_,
    new_n14934_, new_n14935_, new_n14936_, new_n14937_, new_n14938_,
    new_n14939_, new_n14940_, new_n14941_, new_n14942_, new_n14943_,
    new_n14944_, new_n14945_, new_n14946_, new_n14947_, new_n14948_,
    new_n14949_, new_n14950_, new_n14951_, new_n14952_, new_n14953_,
    new_n14954_, new_n14955_, new_n14956_, new_n14957_, new_n14958_,
    new_n14959_, new_n14960_, new_n14961_, new_n14962_, new_n14963_,
    new_n14964_, new_n14965_, new_n14966_, new_n14967_, new_n14968_,
    new_n14969_, new_n14970_, new_n14971_, new_n14972_, new_n14973_,
    new_n14974_, new_n14975_, new_n14976_, new_n14977_, new_n14978_,
    new_n14979_, new_n14980_, new_n14981_, new_n14982_, new_n14983_,
    new_n14984_, new_n14985_, new_n14986_, new_n14987_, new_n14988_,
    new_n14989_, new_n14990_, new_n14991_, new_n14992_, new_n14993_,
    new_n14994_, new_n14995_, new_n14996_, new_n14997_, new_n14998_,
    new_n14999_, new_n15000_, new_n15001_, new_n15002_, new_n15003_,
    new_n15004_, new_n15005_, new_n15006_, new_n15007_, new_n15008_,
    new_n15009_, new_n15010_, new_n15011_, new_n15012_, new_n15013_,
    new_n15014_, new_n15015_, new_n15016_, new_n15017_, new_n15018_,
    new_n15019_, new_n15020_, new_n15021_, new_n15022_, new_n15023_,
    new_n15024_, new_n15025_, new_n15026_, new_n15027_, new_n15028_,
    new_n15029_, new_n15030_, new_n15031_, new_n15032_, new_n15033_,
    new_n15034_, new_n15035_, new_n15036_, new_n15037_, new_n15038_,
    new_n15039_, new_n15040_, new_n15041_, new_n15042_, new_n15043_,
    new_n15044_, new_n15045_, new_n15046_, new_n15047_, new_n15048_,
    new_n15049_, new_n15050_, new_n15051_, new_n15052_, new_n15053_,
    new_n15054_, new_n15055_, new_n15056_, new_n15057_, new_n15058_,
    new_n15059_, new_n15060_, new_n15061_, new_n15062_, new_n15063_,
    new_n15064_, new_n15065_, new_n15067_, new_n15068_, new_n15069_,
    new_n15070_, new_n15071_, new_n15072_, new_n15073_, new_n15074_,
    new_n15075_, new_n15076_, new_n15077_, new_n15078_, new_n15079_,
    new_n15080_, new_n15081_, new_n15082_, new_n15083_, new_n15084_,
    new_n15085_, new_n15086_, new_n15087_, new_n15088_, new_n15089_,
    new_n15090_, new_n15091_, new_n15092_, new_n15093_, new_n15094_,
    new_n15095_, new_n15096_, new_n15097_, new_n15098_, new_n15099_,
    new_n15100_, new_n15101_, new_n15102_, new_n15103_, new_n15104_,
    new_n15105_, new_n15106_, new_n15107_, new_n15108_, new_n15109_,
    new_n15110_, new_n15111_, new_n15112_, new_n15113_, new_n15114_,
    new_n15115_, new_n15116_, new_n15117_, new_n15118_, new_n15119_,
    new_n15120_, new_n15121_, new_n15122_, new_n15123_, new_n15124_,
    new_n15125_, new_n15126_, new_n15127_, new_n15128_, new_n15129_,
    new_n15130_, new_n15131_, new_n15132_, new_n15133_, new_n15134_,
    new_n15135_, new_n15136_, new_n15137_, new_n15138_, new_n15139_,
    new_n15140_, new_n15141_, new_n15142_, new_n15143_, new_n15144_,
    new_n15145_, new_n15146_, new_n15147_, new_n15148_, new_n15149_,
    new_n15150_, new_n15151_, new_n15152_, new_n15153_, new_n15154_,
    new_n15155_, new_n15156_, new_n15157_, new_n15158_, new_n15159_,
    new_n15160_, new_n15161_, new_n15162_, new_n15163_, new_n15164_,
    new_n15165_, new_n15166_, new_n15167_, new_n15168_, new_n15169_,
    new_n15170_, new_n15171_, new_n15172_, new_n15173_, new_n15174_,
    new_n15175_, new_n15176_, new_n15177_, new_n15178_, new_n15179_,
    new_n15180_, new_n15181_, new_n15182_, new_n15183_, new_n15184_,
    new_n15185_, new_n15186_, new_n15187_, new_n15188_, new_n15189_,
    new_n15190_, new_n15191_, new_n15192_, new_n15193_, new_n15194_,
    new_n15195_, new_n15196_, new_n15197_, new_n15198_, new_n15199_,
    new_n15200_, new_n15201_, new_n15202_, new_n15203_, new_n15204_,
    new_n15205_, new_n15206_, new_n15207_, new_n15208_, new_n15209_,
    new_n15210_, new_n15211_, new_n15212_, new_n15213_, new_n15214_,
    new_n15215_, new_n15216_, new_n15217_, new_n15218_, new_n15219_,
    new_n15220_, new_n15221_, new_n15222_, new_n15223_, new_n15224_,
    new_n15225_, new_n15226_, new_n15227_, new_n15228_, new_n15229_,
    new_n15230_, new_n15231_, new_n15232_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15369_,
    new_n15370_, new_n15371_, new_n15372_, new_n15373_, new_n15374_,
    new_n15375_, new_n15376_, new_n15377_, new_n15378_, new_n15379_,
    new_n15380_, new_n15381_, new_n15382_, new_n15383_, new_n15384_,
    new_n15385_, new_n15386_, new_n15387_, new_n15388_, new_n15389_,
    new_n15390_, new_n15391_, new_n15392_, new_n15393_, new_n15394_,
    new_n15395_, new_n15396_, new_n15397_, new_n15398_, new_n15399_,
    new_n15400_, new_n15401_, new_n15402_, new_n15403_, new_n15404_,
    new_n15405_, new_n15406_, new_n15407_, new_n15408_, new_n15409_,
    new_n15410_, new_n15411_, new_n15412_, new_n15413_, new_n15414_,
    new_n15415_, new_n15416_, new_n15417_, new_n15418_, new_n15419_,
    new_n15420_, new_n15421_, new_n15422_, new_n15423_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15428_, new_n15429_,
    new_n15430_, new_n15431_, new_n15432_, new_n15433_, new_n15434_,
    new_n15435_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15469_,
    new_n15470_, new_n15471_, new_n15472_, new_n15473_, new_n15474_,
    new_n15475_, new_n15476_, new_n15477_, new_n15478_, new_n15479_,
    new_n15480_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15488_, new_n15489_,
    new_n15490_, new_n15491_, new_n15492_, new_n15493_, new_n15494_,
    new_n15495_, new_n15496_, new_n15497_, new_n15498_, new_n15499_,
    new_n15500_, new_n15501_, new_n15502_, new_n15503_, new_n15504_,
    new_n15505_, new_n15506_, new_n15507_, new_n15508_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16107_, new_n16108_, new_n16109_, new_n16110_, new_n16111_,
    new_n16112_, new_n16113_, new_n16114_, new_n16115_, new_n16116_,
    new_n16117_, new_n16118_, new_n16119_, new_n16120_, new_n16121_,
    new_n16122_, new_n16123_, new_n16124_, new_n16125_, new_n16126_,
    new_n16127_, new_n16128_, new_n16129_, new_n16130_, new_n16131_,
    new_n16132_, new_n16133_, new_n16134_, new_n16135_, new_n16136_,
    new_n16137_, new_n16138_, new_n16139_, new_n16140_, new_n16141_,
    new_n16142_, new_n16143_, new_n16144_, new_n16145_, new_n16146_,
    new_n16147_, new_n16148_, new_n16149_, new_n16150_, new_n16151_,
    new_n16152_, new_n16153_, new_n16154_, new_n16155_, new_n16156_,
    new_n16157_, new_n16158_, new_n16159_, new_n16160_, new_n16161_,
    new_n16162_, new_n16163_, new_n16164_, new_n16165_, new_n16166_,
    new_n16167_, new_n16168_, new_n16169_, new_n16170_, new_n16171_,
    new_n16172_, new_n16173_, new_n16174_, new_n16175_, new_n16176_,
    new_n16177_, new_n16178_, new_n16179_, new_n16180_, new_n16181_,
    new_n16182_, new_n16183_, new_n16184_, new_n16185_, new_n16186_,
    new_n16187_, new_n16188_, new_n16189_, new_n16190_, new_n16191_,
    new_n16192_, new_n16193_, new_n16194_, new_n16195_, new_n16196_,
    new_n16197_, new_n16198_, new_n16199_, new_n16200_, new_n16201_,
    new_n16202_, new_n16203_, new_n16204_, new_n16205_, new_n16206_,
    new_n16207_, new_n16208_, new_n16209_, new_n16210_, new_n16211_,
    new_n16212_, new_n16213_, new_n16214_, new_n16215_, new_n16216_,
    new_n16217_, new_n16218_, new_n16219_, new_n16220_, new_n16221_,
    new_n16222_, new_n16223_, new_n16224_, new_n16225_, new_n16226_,
    new_n16227_, new_n16228_, new_n16229_, new_n16230_, new_n16231_,
    new_n16232_, new_n16233_, new_n16234_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16239_, new_n16240_, new_n16241_,
    new_n16242_, new_n16243_, new_n16244_, new_n16245_, new_n16246_,
    new_n16247_, new_n16248_, new_n16249_, new_n16250_, new_n16251_,
    new_n16252_, new_n16253_, new_n16254_, new_n16255_, new_n16256_,
    new_n16257_, new_n16258_, new_n16259_, new_n16260_, new_n16261_,
    new_n16262_, new_n16263_, new_n16264_, new_n16265_, new_n16266_,
    new_n16267_, new_n16268_, new_n16269_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16274_, new_n16275_, new_n16276_,
    new_n16277_, new_n16278_, new_n16279_, new_n16280_, new_n16281_,
    new_n16282_, new_n16283_, new_n16284_, new_n16285_, new_n16286_,
    new_n16287_, new_n16288_, new_n16289_, new_n16290_, new_n16291_,
    new_n16292_, new_n16293_, new_n16294_, new_n16295_, new_n16296_,
    new_n16297_, new_n16298_, new_n16299_, new_n16300_, new_n16301_,
    new_n16302_, new_n16303_, new_n16304_, new_n16305_, new_n16306_,
    new_n16307_, new_n16308_, new_n16309_, new_n16310_, new_n16311_,
    new_n16312_, new_n16313_, new_n16314_, new_n16315_, new_n16316_,
    new_n16317_, new_n16318_, new_n16319_, new_n16320_, new_n16321_,
    new_n16322_, new_n16323_, new_n16324_, new_n16325_, new_n16326_,
    new_n16327_, new_n16328_, new_n16329_, new_n16330_, new_n16331_,
    new_n16332_, new_n16333_, new_n16334_, new_n16335_, new_n16336_,
    new_n16337_, new_n16338_, new_n16339_, new_n16340_, new_n16341_,
    new_n16342_, new_n16343_, new_n16344_, new_n16345_, new_n16346_,
    new_n16347_, new_n16348_, new_n16349_, new_n16350_, new_n16351_,
    new_n16352_, new_n16353_, new_n16354_, new_n16355_, new_n16356_,
    new_n16357_, new_n16358_, new_n16359_, new_n16360_, new_n16361_,
    new_n16362_, new_n16363_, new_n16364_, new_n16365_, new_n16366_,
    new_n16367_, new_n16368_, new_n16369_, new_n16370_, new_n16371_,
    new_n16372_, new_n16373_, new_n16374_, new_n16375_, new_n16376_,
    new_n16377_, new_n16378_, new_n16379_, new_n16380_, new_n16381_,
    new_n16382_, new_n16383_, new_n16384_, new_n16385_, new_n16386_,
    new_n16387_, new_n16388_, new_n16389_, new_n16390_, new_n16391_,
    new_n16392_, new_n16393_, new_n16394_, new_n16395_, new_n16396_,
    new_n16397_, new_n16398_, new_n16399_, new_n16400_, new_n16401_,
    new_n16402_, new_n16403_, new_n16404_, new_n16405_, new_n16406_,
    new_n16407_, new_n16408_, new_n16409_, new_n16410_, new_n16411_,
    new_n16412_, new_n16413_, new_n16414_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16426_,
    new_n16427_, new_n16428_, new_n16429_, new_n16430_, new_n16431_,
    new_n16432_, new_n16433_, new_n16434_, new_n16435_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16458_, new_n16459_, new_n16460_, new_n16461_,
    new_n16462_, new_n16463_, new_n16464_, new_n16465_, new_n16466_,
    new_n16467_, new_n16468_, new_n16469_, new_n16470_, new_n16471_,
    new_n16472_, new_n16473_, new_n16474_, new_n16475_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16490_, new_n16491_,
    new_n16492_, new_n16493_, new_n16494_, new_n16495_, new_n16496_,
    new_n16497_, new_n16498_, new_n16499_, new_n16500_, new_n16501_,
    new_n16502_, new_n16503_, new_n16504_, new_n16505_, new_n16506_,
    new_n16507_, new_n16508_, new_n16509_, new_n16510_, new_n16511_,
    new_n16512_, new_n16513_, new_n16514_, new_n16515_, new_n16516_,
    new_n16517_, new_n16518_, new_n16519_, new_n16520_, new_n16521_,
    new_n16522_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16530_, new_n16531_,
    new_n16532_, new_n16533_, new_n16534_, new_n16535_, new_n16536_,
    new_n16537_, new_n16538_, new_n16539_, new_n16540_, new_n16541_,
    new_n16542_, new_n16543_, new_n16544_, new_n16545_, new_n16546_,
    new_n16547_, new_n16548_, new_n16549_, new_n16550_, new_n16551_,
    new_n16552_, new_n16553_, new_n16554_, new_n16555_, new_n16556_,
    new_n16557_, new_n16558_, new_n16559_, new_n16560_, new_n16561_,
    new_n16562_, new_n16563_, new_n16564_, new_n16565_, new_n16566_,
    new_n16567_, new_n16568_, new_n16569_, new_n16570_, new_n16571_,
    new_n16572_, new_n16573_, new_n16574_, new_n16575_, new_n16576_,
    new_n16577_, new_n16578_, new_n16579_, new_n16580_, new_n16581_,
    new_n16582_, new_n16583_, new_n16584_, new_n16585_, new_n16586_,
    new_n16587_, new_n16588_, new_n16589_, new_n16590_, new_n16591_,
    new_n16592_, new_n16593_, new_n16594_, new_n16595_, new_n16596_,
    new_n16597_, new_n16598_, new_n16599_, new_n16600_, new_n16601_,
    new_n16602_, new_n16603_, new_n16604_, new_n16605_, new_n16606_,
    new_n16607_, new_n16608_, new_n16609_, new_n16610_, new_n16611_,
    new_n16613_, new_n16614_, new_n16615_, new_n16616_, new_n16617_,
    new_n16618_, new_n16619_, new_n16620_, new_n16621_, new_n16622_,
    new_n16623_, new_n16624_, new_n16625_, new_n16626_, new_n16627_,
    new_n16628_, new_n16629_, new_n16630_, new_n16631_, new_n16632_,
    new_n16633_, new_n16634_, new_n16635_, new_n16636_, new_n16637_,
    new_n16638_, new_n16639_, new_n16640_, new_n16641_, new_n16642_,
    new_n16643_, new_n16644_, new_n16645_, new_n16646_, new_n16647_,
    new_n16648_, new_n16649_, new_n16650_, new_n16651_, new_n16652_,
    new_n16653_, new_n16654_, new_n16655_, new_n16656_, new_n16657_,
    new_n16658_, new_n16659_, new_n16660_, new_n16661_, new_n16662_,
    new_n16663_, new_n16664_, new_n16665_, new_n16666_, new_n16667_,
    new_n16668_, new_n16669_, new_n16670_, new_n16671_, new_n16672_,
    new_n16673_, new_n16674_, new_n16675_, new_n16676_, new_n16677_,
    new_n16678_, new_n16679_, new_n16680_, new_n16681_, new_n16682_,
    new_n16683_, new_n16684_, new_n16685_, new_n16686_, new_n16687_,
    new_n16688_, new_n16689_, new_n16690_, new_n16691_, new_n16692_,
    new_n16693_, new_n16694_, new_n16695_, new_n16696_, new_n16697_,
    new_n16698_, new_n16699_, new_n16700_, new_n16701_, new_n16702_,
    new_n16703_, new_n16704_, new_n16705_, new_n16706_, new_n16707_,
    new_n16708_, new_n16709_, new_n16710_, new_n16711_, new_n16712_,
    new_n16713_, new_n16714_, new_n16715_, new_n16716_, new_n16717_,
    new_n16718_, new_n16719_, new_n16720_, new_n16721_, new_n16722_,
    new_n16723_, new_n16724_, new_n16725_, new_n16726_, new_n16727_,
    new_n16728_, new_n16729_, new_n16730_, new_n16731_, new_n16732_,
    new_n16733_, new_n16734_, new_n16735_, new_n16736_, new_n16737_,
    new_n16738_, new_n16739_, new_n16740_, new_n16741_, new_n16742_,
    new_n16743_, new_n16744_, new_n16745_, new_n16746_, new_n16747_,
    new_n16748_, new_n16749_, new_n16750_, new_n16751_, new_n16752_,
    new_n16753_, new_n16754_, new_n16755_, new_n16756_, new_n16757_,
    new_n16758_, new_n16759_, new_n16760_, new_n16761_, new_n16762_,
    new_n16763_, new_n16764_, new_n16765_, new_n16766_, new_n16767_,
    new_n16768_, new_n16769_, new_n16770_, new_n16771_, new_n16772_,
    new_n16773_, new_n16774_, new_n16775_, new_n16776_, new_n16777_,
    new_n16778_, new_n16779_, new_n16780_, new_n16781_, new_n16782_,
    new_n16783_, new_n16784_, new_n16785_, new_n16786_, new_n16787_,
    new_n16788_, new_n16789_, new_n16790_, new_n16791_, new_n16792_,
    new_n16793_, new_n16794_, new_n16795_, new_n16796_, new_n16797_,
    new_n16798_, new_n16799_, new_n16800_, new_n16801_, new_n16802_,
    new_n16803_, new_n16804_, new_n16805_, new_n16806_, new_n16807_,
    new_n16808_, new_n16809_, new_n16810_, new_n16811_, new_n16812_,
    new_n16813_, new_n16814_, new_n16815_, new_n16816_, new_n16817_,
    new_n16818_, new_n16819_, new_n16820_, new_n16821_, new_n16822_,
    new_n16823_, new_n16824_, new_n16825_, new_n16826_, new_n16827_,
    new_n16828_, new_n16829_, new_n16830_, new_n16831_, new_n16832_,
    new_n16833_, new_n16834_, new_n16835_, new_n16836_, new_n16837_,
    new_n16838_, new_n16839_, new_n16840_, new_n16841_, new_n16842_,
    new_n16843_, new_n16844_, new_n16845_, new_n16846_, new_n16847_,
    new_n16848_, new_n16849_, new_n16850_, new_n16851_, new_n16852_,
    new_n16853_, new_n16854_, new_n16855_, new_n16856_, new_n16857_,
    new_n16858_, new_n16859_, new_n16860_, new_n16861_, new_n16862_,
    new_n16863_, new_n16864_, new_n16865_, new_n16866_, new_n16867_,
    new_n16868_, new_n16869_, new_n16870_, new_n16871_, new_n16872_,
    new_n16873_, new_n16874_, new_n16875_, new_n16876_, new_n16877_,
    new_n16878_, new_n16879_, new_n16880_, new_n16881_, new_n16882_,
    new_n16883_, new_n16884_, new_n16885_, new_n16886_, new_n16887_,
    new_n16888_, new_n16889_, new_n16890_, new_n16891_, new_n16892_,
    new_n16893_, new_n16894_, new_n16895_, new_n16896_, new_n16897_,
    new_n16898_, new_n16899_, new_n16900_, new_n16901_, new_n16902_,
    new_n16903_, new_n16904_, new_n16905_, new_n16906_, new_n16907_,
    new_n16908_, new_n16909_, new_n16910_, new_n16911_, new_n16912_,
    new_n16913_, new_n16914_, new_n16915_, new_n16916_, new_n16917_,
    new_n16918_, new_n16919_, new_n16920_, new_n16921_, new_n16922_,
    new_n16923_, new_n16924_, new_n16925_, new_n16926_, new_n16927_,
    new_n16928_, new_n16929_, new_n16930_, new_n16931_, new_n16932_,
    new_n16933_, new_n16934_, new_n16935_, new_n16936_, new_n16937_,
    new_n16938_, new_n16939_, new_n16940_, new_n16941_, new_n16942_,
    new_n16943_, new_n16944_, new_n16945_, new_n16946_, new_n16947_,
    new_n16948_, new_n16949_, new_n16950_, new_n16951_, new_n16952_,
    new_n16953_, new_n16954_, new_n16955_, new_n16956_, new_n16957_,
    new_n16958_, new_n16959_, new_n16960_, new_n16961_, new_n16962_,
    new_n16963_, new_n16964_, new_n16965_, new_n16966_, new_n16967_,
    new_n16968_, new_n16969_, new_n16970_, new_n16971_, new_n16972_,
    new_n16973_, new_n16974_, new_n16975_, new_n16976_, new_n16977_,
    new_n16978_, new_n16979_, new_n16980_, new_n16981_, new_n16982_,
    new_n16983_, new_n16984_, new_n16985_, new_n16986_, new_n16987_,
    new_n16988_, new_n16989_, new_n16990_, new_n16991_, new_n16992_,
    new_n16993_, new_n16994_, new_n16995_, new_n16996_, new_n16997_,
    new_n16998_, new_n16999_, new_n17000_, new_n17001_, new_n17002_,
    new_n17003_, new_n17004_, new_n17005_, new_n17006_, new_n17007_,
    new_n17008_, new_n17009_, new_n17010_, new_n17011_, new_n17012_,
    new_n17013_, new_n17014_, new_n17015_, new_n17016_, new_n17017_,
    new_n17018_, new_n17019_, new_n17020_, new_n17021_, new_n17022_,
    new_n17023_, new_n17024_, new_n17025_, new_n17026_, new_n17027_,
    new_n17028_, new_n17029_, new_n17030_, new_n17031_, new_n17032_,
    new_n17033_, new_n17034_, new_n17035_, new_n17036_, new_n17037_,
    new_n17038_, new_n17039_, new_n17040_, new_n17041_, new_n17042_,
    new_n17043_, new_n17044_, new_n17045_, new_n17046_, new_n17047_,
    new_n17048_, new_n17049_, new_n17050_, new_n17051_, new_n17052_,
    new_n17053_, new_n17054_, new_n17055_, new_n17056_, new_n17057_,
    new_n17058_, new_n17059_, new_n17060_, new_n17061_, new_n17062_,
    new_n17063_, new_n17064_, new_n17065_, new_n17066_, new_n17067_,
    new_n17068_, new_n17069_, new_n17070_, new_n17071_, new_n17072_,
    new_n17073_, new_n17074_, new_n17075_, new_n17076_, new_n17077_,
    new_n17078_, new_n17079_, new_n17080_, new_n17081_, new_n17082_,
    new_n17083_, new_n17084_, new_n17085_, new_n17086_, new_n17087_,
    new_n17088_, new_n17089_, new_n17090_, new_n17091_, new_n17092_,
    new_n17093_, new_n17094_, new_n17095_, new_n17096_, new_n17097_,
    new_n17098_, new_n17099_, new_n17100_, new_n17101_, new_n17102_,
    new_n17103_, new_n17104_, new_n17105_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17124_, new_n17125_, new_n17126_, new_n17127_,
    new_n17128_, new_n17129_, new_n17130_, new_n17131_, new_n17132_,
    new_n17133_, new_n17134_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17147_,
    new_n17148_, new_n17149_, new_n17150_, new_n17151_, new_n17152_,
    new_n17153_, new_n17154_, new_n17155_, new_n17156_, new_n17157_,
    new_n17158_, new_n17159_, new_n17160_, new_n17161_, new_n17162_,
    new_n17163_, new_n17164_, new_n17165_, new_n17166_, new_n17168_,
    new_n17169_, new_n17170_, new_n17171_, new_n17172_, new_n17173_,
    new_n17174_, new_n17175_, new_n17176_, new_n17177_, new_n17178_,
    new_n17179_, new_n17180_, new_n17181_, new_n17182_, new_n17183_,
    new_n17184_, new_n17185_, new_n17186_, new_n17187_, new_n17188_,
    new_n17189_, new_n17190_, new_n17191_, new_n17192_, new_n17193_,
    new_n17194_, new_n17195_, new_n17196_, new_n17197_, new_n17198_,
    new_n17199_, new_n17200_, new_n17201_, new_n17202_, new_n17203_,
    new_n17204_, new_n17205_, new_n17206_, new_n17207_, new_n17208_,
    new_n17209_, new_n17210_, new_n17211_, new_n17212_, new_n17213_,
    new_n17214_, new_n17215_, new_n17216_, new_n17217_, new_n17218_,
    new_n17219_, new_n17220_, new_n17221_, new_n17222_, new_n17223_,
    new_n17224_, new_n17225_, new_n17226_, new_n17227_, new_n17228_,
    new_n17229_, new_n17230_, new_n17231_, new_n17232_, new_n17233_,
    new_n17234_, new_n17235_, new_n17236_, new_n17237_, new_n17238_,
    new_n17239_, new_n17240_, new_n17241_, new_n17242_, new_n17243_,
    new_n17244_, new_n17245_, new_n17246_, new_n17247_, new_n17248_,
    new_n17249_, new_n17250_, new_n17251_, new_n17252_, new_n17253_,
    new_n17254_, new_n17255_, new_n17256_, new_n17257_, new_n17258_,
    new_n17259_, new_n17260_, new_n17261_, new_n17262_, new_n17263_,
    new_n17264_, new_n17265_, new_n17266_, new_n17267_, new_n17268_,
    new_n17269_, new_n17270_, new_n17271_, new_n17272_, new_n17273_,
    new_n17274_, new_n17275_, new_n17276_, new_n17277_, new_n17278_,
    new_n17279_, new_n17280_, new_n17281_, new_n17282_, new_n17283_,
    new_n17284_, new_n17285_, new_n17286_, new_n17287_, new_n17288_,
    new_n17289_, new_n17290_, new_n17291_, new_n17292_, new_n17293_,
    new_n17294_, new_n17295_, new_n17296_, new_n17297_, new_n17298_,
    new_n17299_, new_n17300_, new_n17301_, new_n17302_, new_n17303_,
    new_n17304_, new_n17305_, new_n17306_, new_n17307_, new_n17308_,
    new_n17309_, new_n17310_, new_n17311_, new_n17312_, new_n17313_,
    new_n17314_, new_n17315_, new_n17316_, new_n17317_, new_n17318_,
    new_n17319_, new_n17320_, new_n17321_, new_n17322_, new_n17323_,
    new_n17324_, new_n17325_, new_n17326_, new_n17327_, new_n17328_,
    new_n17329_, new_n17330_, new_n17331_, new_n17332_, new_n17333_,
    new_n17334_, new_n17335_, new_n17336_, new_n17337_, new_n17338_,
    new_n17339_, new_n17340_, new_n17341_, new_n17342_, new_n17343_,
    new_n17344_, new_n17345_, new_n17346_, new_n17347_, new_n17348_,
    new_n17349_, new_n17350_, new_n17351_, new_n17352_, new_n17353_,
    new_n17354_, new_n17355_, new_n17356_, new_n17357_, new_n17358_,
    new_n17359_, new_n17360_, new_n17361_, new_n17362_, new_n17363_,
    new_n17364_, new_n17365_, new_n17366_, new_n17367_, new_n17368_,
    new_n17369_, new_n17370_, new_n17371_, new_n17372_, new_n17373_,
    new_n17374_, new_n17375_, new_n17376_, new_n17377_, new_n17378_,
    new_n17379_, new_n17380_, new_n17381_, new_n17382_, new_n17383_,
    new_n17384_, new_n17385_, new_n17386_, new_n17387_, new_n17388_,
    new_n17389_, new_n17390_, new_n17391_, new_n17392_, new_n17393_,
    new_n17394_, new_n17395_, new_n17396_, new_n17397_, new_n17398_,
    new_n17399_, new_n17400_, new_n17401_, new_n17402_, new_n17403_,
    new_n17404_, new_n17405_, new_n17406_, new_n17407_, new_n17408_,
    new_n17409_, new_n17410_, new_n17411_, new_n17412_, new_n17413_,
    new_n17414_, new_n17415_, new_n17416_, new_n17417_, new_n17418_,
    new_n17419_, new_n17420_, new_n17421_, new_n17422_, new_n17423_,
    new_n17424_, new_n17425_, new_n17426_, new_n17427_, new_n17428_,
    new_n17429_, new_n17430_, new_n17431_, new_n17432_, new_n17433_,
    new_n17434_, new_n17435_, new_n17436_, new_n17437_, new_n17438_,
    new_n17439_, new_n17440_, new_n17441_, new_n17442_, new_n17443_,
    new_n17444_, new_n17445_, new_n17446_, new_n17447_, new_n17448_,
    new_n17449_, new_n17450_, new_n17451_, new_n17452_, new_n17453_,
    new_n17454_, new_n17455_, new_n17456_, new_n17457_, new_n17458_,
    new_n17459_, new_n17460_, new_n17461_, new_n17462_, new_n17463_,
    new_n17464_, new_n17465_, new_n17466_, new_n17467_, new_n17468_,
    new_n17469_, new_n17470_, new_n17471_, new_n17472_, new_n17473_,
    new_n17474_, new_n17475_, new_n17476_, new_n17477_, new_n17478_,
    new_n17479_, new_n17480_, new_n17481_, new_n17482_, new_n17483_,
    new_n17484_, new_n17485_, new_n17486_, new_n17487_, new_n17488_,
    new_n17489_, new_n17490_, new_n17491_, new_n17492_, new_n17493_,
    new_n17494_, new_n17495_, new_n17496_, new_n17497_, new_n17498_,
    new_n17499_, new_n17500_, new_n17501_, new_n17502_, new_n17503_,
    new_n17504_, new_n17505_, new_n17506_, new_n17507_, new_n17508_,
    new_n17509_, new_n17510_, new_n17511_, new_n17512_, new_n17513_,
    new_n17514_, new_n17515_, new_n17516_, new_n17517_, new_n17518_,
    new_n17519_, new_n17520_, new_n17521_, new_n17522_, new_n17523_,
    new_n17524_, new_n17525_, new_n17526_, new_n17527_, new_n17528_,
    new_n17529_, new_n17530_, new_n17531_, new_n17532_, new_n17533_,
    new_n17534_, new_n17535_, new_n17536_, new_n17537_, new_n17538_,
    new_n17539_, new_n17540_, new_n17541_, new_n17542_, new_n17543_,
    new_n17544_, new_n17545_, new_n17546_, new_n17547_, new_n17548_,
    new_n17549_, new_n17550_, new_n17551_, new_n17552_, new_n17553_,
    new_n17554_, new_n17555_, new_n17556_, new_n17557_, new_n17558_,
    new_n17559_, new_n17560_, new_n17561_, new_n17562_, new_n17563_,
    new_n17564_, new_n17565_, new_n17566_, new_n17567_, new_n17568_,
    new_n17569_, new_n17570_, new_n17571_, new_n17572_, new_n17573_,
    new_n17574_, new_n17575_, new_n17576_, new_n17577_, new_n17578_,
    new_n17579_, new_n17580_, new_n17581_, new_n17582_, new_n17583_,
    new_n17584_, new_n17585_, new_n17586_, new_n17587_, new_n17588_,
    new_n17589_, new_n17590_, new_n17591_, new_n17592_, new_n17593_,
    new_n17594_, new_n17595_, new_n17596_, new_n17597_, new_n17598_,
    new_n17599_, new_n17600_, new_n17601_, new_n17602_, new_n17603_,
    new_n17604_, new_n17605_, new_n17606_, new_n17607_, new_n17608_,
    new_n17609_, new_n17610_, new_n17611_, new_n17612_, new_n17613_,
    new_n17614_, new_n17615_, new_n17616_, new_n17617_, new_n17618_,
    new_n17619_, new_n17620_, new_n17621_, new_n17622_, new_n17623_,
    new_n17624_, new_n17625_, new_n17626_, new_n17627_, new_n17628_,
    new_n17629_, new_n17630_, new_n17631_, new_n17632_, new_n17633_,
    new_n17634_, new_n17635_, new_n17636_, new_n17637_, new_n17638_,
    new_n17639_, new_n17640_, new_n17641_, new_n17642_, new_n17643_,
    new_n17644_, new_n17645_, new_n17646_, new_n17647_, new_n17648_,
    new_n17649_, new_n17650_, new_n17651_, new_n17652_, new_n17653_,
    new_n17654_, new_n17655_, new_n17656_, new_n17657_, new_n17658_,
    new_n17659_, new_n17660_, new_n17661_, new_n17662_, new_n17663_,
    new_n17664_, new_n17665_, new_n17666_, new_n17667_, new_n17668_,
    new_n17669_, new_n17670_, new_n17671_, new_n17672_, new_n17673_,
    new_n17674_, new_n17675_, new_n17676_, new_n17677_, new_n17678_,
    new_n17679_, new_n17680_, new_n17681_, new_n17682_, new_n17683_,
    new_n17684_, new_n17685_, new_n17686_, new_n17687_, new_n17688_,
    new_n17689_, new_n17690_, new_n17692_, new_n17693_, new_n17694_,
    new_n17695_, new_n17696_, new_n17697_, new_n17698_, new_n17699_,
    new_n17700_, new_n17701_, new_n17702_, new_n17703_, new_n17704_,
    new_n17705_, new_n17706_, new_n17707_, new_n17708_, new_n17709_,
    new_n17710_, new_n17711_, new_n17712_, new_n17713_, new_n17714_,
    new_n17715_, new_n17716_, new_n17717_, new_n17718_, new_n17719_,
    new_n17720_, new_n17721_, new_n17722_, new_n17723_, new_n17724_,
    new_n17725_, new_n17726_, new_n17727_, new_n17728_, new_n17729_,
    new_n17730_, new_n17731_, new_n17732_, new_n17733_, new_n17734_,
    new_n17735_, new_n17736_, new_n17737_, new_n17738_, new_n17739_,
    new_n17740_, new_n17741_, new_n17742_, new_n17743_, new_n17744_,
    new_n17745_, new_n17746_, new_n17747_, new_n17748_, new_n17749_,
    new_n17750_, new_n17751_, new_n17752_, new_n17753_, new_n17754_,
    new_n17755_, new_n17756_, new_n17757_, new_n17758_, new_n17759_,
    new_n17760_, new_n17761_, new_n17762_, new_n17763_, new_n17764_,
    new_n17765_, new_n17766_, new_n17767_, new_n17768_, new_n17769_,
    new_n17770_, new_n17771_, new_n17772_, new_n17773_, new_n17774_,
    new_n17775_, new_n17776_, new_n17777_, new_n17778_, new_n17779_,
    new_n17780_, new_n17781_, new_n17782_, new_n17783_, new_n17784_,
    new_n17785_, new_n17786_, new_n17787_, new_n17788_, new_n17789_,
    new_n17790_, new_n17791_, new_n17792_, new_n17793_, new_n17794_,
    new_n17795_, new_n17796_, new_n17797_, new_n17798_, new_n17799_,
    new_n17800_, new_n17801_, new_n17802_, new_n17803_, new_n17804_,
    new_n17805_, new_n17806_, new_n17807_, new_n17808_, new_n17809_,
    new_n17810_, new_n17811_, new_n17812_, new_n17813_, new_n17814_,
    new_n17815_, new_n17816_, new_n17817_, new_n17818_, new_n17819_,
    new_n17820_, new_n17821_, new_n17822_, new_n17823_, new_n17824_,
    new_n17825_, new_n17826_, new_n17827_, new_n17828_, new_n17829_,
    new_n17830_, new_n17831_, new_n17832_, new_n17833_, new_n17834_,
    new_n17835_, new_n17836_, new_n17837_, new_n17838_, new_n17839_,
    new_n17840_, new_n17841_, new_n17842_, new_n17843_, new_n17844_,
    new_n17845_, new_n17846_, new_n17847_, new_n17848_, new_n17849_,
    new_n17850_, new_n17851_, new_n17852_, new_n17853_, new_n17854_,
    new_n17855_, new_n17856_, new_n17857_, new_n17858_, new_n17859_,
    new_n17860_, new_n17861_, new_n17862_, new_n17863_, new_n17864_,
    new_n17865_, new_n17866_, new_n17867_, new_n17868_, new_n17869_,
    new_n17870_, new_n17871_, new_n17872_, new_n17873_, new_n17874_,
    new_n17875_, new_n17876_, new_n17877_, new_n17878_, new_n17879_,
    new_n17880_, new_n17881_, new_n17882_, new_n17883_, new_n17884_,
    new_n17885_, new_n17886_, new_n17887_, new_n17888_, new_n17889_,
    new_n17890_, new_n17891_, new_n17892_, new_n17893_, new_n17894_,
    new_n17895_, new_n17896_, new_n17897_, new_n17898_, new_n17899_,
    new_n17900_, new_n17901_, new_n17902_, new_n17903_, new_n17904_,
    new_n17905_, new_n17906_, new_n17907_, new_n17908_, new_n17909_,
    new_n17910_, new_n17911_, new_n17912_, new_n17913_, new_n17914_,
    new_n17915_, new_n17916_, new_n17917_, new_n17918_, new_n17919_,
    new_n17920_, new_n17921_, new_n17922_, new_n17923_, new_n17924_,
    new_n17925_, new_n17926_, new_n17927_, new_n17928_, new_n17929_,
    new_n17930_, new_n17931_, new_n17932_, new_n17933_, new_n17934_,
    new_n17935_, new_n17936_, new_n17937_, new_n17938_, new_n17939_,
    new_n17940_, new_n17941_, new_n17942_, new_n17943_, new_n17944_,
    new_n17945_, new_n17946_, new_n17947_, new_n17948_, new_n17949_,
    new_n17950_, new_n17951_, new_n17952_, new_n17953_, new_n17954_,
    new_n17955_, new_n17956_, new_n17957_, new_n17958_, new_n17959_,
    new_n17960_, new_n17961_, new_n17962_, new_n17963_, new_n17964_,
    new_n17965_, new_n17966_, new_n17967_, new_n17968_, new_n17969_,
    new_n17970_, new_n17971_, new_n17972_, new_n17973_, new_n17974_,
    new_n17975_, new_n17976_, new_n17977_, new_n17978_, new_n17979_,
    new_n17980_, new_n17981_, new_n17982_, new_n17983_, new_n17984_,
    new_n17985_, new_n17986_, new_n17987_, new_n17988_, new_n17989_,
    new_n17990_, new_n17991_, new_n17992_, new_n17993_, new_n17994_,
    new_n17995_, new_n17996_, new_n17997_, new_n17998_, new_n17999_,
    new_n18000_, new_n18001_, new_n18002_, new_n18003_, new_n18004_,
    new_n18005_, new_n18006_, new_n18007_, new_n18008_, new_n18009_,
    new_n18010_, new_n18011_, new_n18012_, new_n18013_, new_n18014_,
    new_n18015_, new_n18016_, new_n18017_, new_n18018_, new_n18019_,
    new_n18020_, new_n18021_, new_n18022_, new_n18023_, new_n18024_,
    new_n18025_, new_n18026_, new_n18027_, new_n18028_, new_n18029_,
    new_n18030_, new_n18031_, new_n18032_, new_n18033_, new_n18034_,
    new_n18035_, new_n18036_, new_n18037_, new_n18038_, new_n18039_,
    new_n18040_, new_n18041_, new_n18042_, new_n18043_, new_n18044_,
    new_n18045_, new_n18046_, new_n18047_, new_n18048_, new_n18049_,
    new_n18050_, new_n18051_, new_n18052_, new_n18053_, new_n18054_,
    new_n18055_, new_n18056_, new_n18057_, new_n18058_, new_n18059_,
    new_n18060_, new_n18061_, new_n18062_, new_n18063_, new_n18064_,
    new_n18065_, new_n18066_, new_n18067_, new_n18068_, new_n18069_,
    new_n18070_, new_n18071_, new_n18072_, new_n18073_, new_n18074_,
    new_n18075_, new_n18076_, new_n18077_, new_n18078_, new_n18079_,
    new_n18080_, new_n18081_, new_n18082_, new_n18083_, new_n18084_,
    new_n18085_, new_n18086_, new_n18087_, new_n18088_, new_n18089_,
    new_n18090_, new_n18091_, new_n18092_, new_n18093_, new_n18094_,
    new_n18095_, new_n18096_, new_n18097_, new_n18098_, new_n18099_,
    new_n18100_, new_n18101_, new_n18102_, new_n18103_, new_n18104_,
    new_n18105_, new_n18106_, new_n18107_, new_n18108_, new_n18109_,
    new_n18110_, new_n18111_, new_n18112_, new_n18113_, new_n18114_,
    new_n18115_, new_n18116_, new_n18117_, new_n18118_, new_n18119_,
    new_n18120_, new_n18121_, new_n18122_, new_n18123_, new_n18124_,
    new_n18125_, new_n18126_, new_n18127_, new_n18128_, new_n18129_,
    new_n18130_, new_n18131_, new_n18132_, new_n18133_, new_n18134_,
    new_n18135_, new_n18136_, new_n18137_, new_n18138_, new_n18139_,
    new_n18140_, new_n18141_, new_n18142_, new_n18143_, new_n18144_,
    new_n18145_, new_n18146_, new_n18147_, new_n18148_, new_n18149_,
    new_n18150_, new_n18151_, new_n18152_, new_n18153_, new_n18154_,
    new_n18155_, new_n18156_, new_n18157_, new_n18158_, new_n18159_,
    new_n18160_, new_n18161_, new_n18162_, new_n18163_, new_n18164_,
    new_n18165_, new_n18166_, new_n18167_, new_n18168_, new_n18169_,
    new_n18170_, new_n18171_, new_n18172_, new_n18173_, new_n18174_,
    new_n18175_, new_n18176_, new_n18177_, new_n18178_, new_n18179_,
    new_n18180_, new_n18181_, new_n18182_, new_n18183_, new_n18184_,
    new_n18185_, new_n18186_, new_n18187_, new_n18188_, new_n18189_,
    new_n18190_, new_n18191_, new_n18192_, new_n18193_, new_n18194_,
    new_n18195_, new_n18196_, new_n18197_, new_n18198_, new_n18199_,
    new_n18200_, new_n18201_, new_n18202_, new_n18203_, new_n18204_,
    new_n18205_, new_n18206_, new_n18207_, new_n18208_, new_n18209_,
    new_n18210_, new_n18211_, new_n18212_, new_n18213_, new_n18214_,
    new_n18215_, new_n18216_, new_n18217_, new_n18218_, new_n18219_,
    new_n18220_, new_n18221_, new_n18222_, new_n18223_, new_n18224_,
    new_n18225_, new_n18226_, new_n18227_, new_n18228_, new_n18229_,
    new_n18230_, new_n18231_, new_n18232_, new_n18233_, new_n18234_,
    new_n18235_, new_n18236_, new_n18237_, new_n18238_, new_n18239_,
    new_n18240_, new_n18241_, new_n18242_, new_n18243_, new_n18244_,
    new_n18245_, new_n18246_, new_n18247_, new_n18248_, new_n18249_,
    new_n18250_, new_n18251_, new_n18252_, new_n18253_, new_n18254_,
    new_n18255_, new_n18256_, new_n18257_, new_n18258_, new_n18259_,
    new_n18260_, new_n18261_, new_n18262_, new_n18263_, new_n18264_,
    new_n18265_, new_n18266_, new_n18267_, new_n18268_, new_n18269_,
    new_n18270_, new_n18271_, new_n18272_, new_n18273_, new_n18274_,
    new_n18275_, new_n18276_, new_n18277_, new_n18278_, new_n18279_,
    new_n18280_, new_n18281_, new_n18282_, new_n18283_, new_n18284_,
    new_n18285_, new_n18286_, new_n18287_, new_n18288_, new_n18289_,
    new_n18290_, new_n18291_, new_n18292_, new_n18293_, new_n18294_,
    new_n18295_, new_n18296_, new_n18297_, new_n18298_, new_n18299_,
    new_n18300_, new_n18301_, new_n18302_, new_n18303_, new_n18304_,
    new_n18305_, new_n18306_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18338_, new_n18339_, new_n18340_,
    new_n18341_, new_n18342_, new_n18343_, new_n18344_, new_n18345_,
    new_n18346_, new_n18347_, new_n18348_, new_n18349_, new_n18350_,
    new_n18351_, new_n18352_, new_n18353_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18360_,
    new_n18361_, new_n18362_, new_n18363_, new_n18364_, new_n18365_,
    new_n18366_, new_n18367_, new_n18368_, new_n18369_, new_n18370_,
    new_n18371_, new_n18372_, new_n18373_, new_n18374_, new_n18375_,
    new_n18376_, new_n18377_, new_n18378_, new_n18379_, new_n18380_,
    new_n18381_, new_n18382_, new_n18383_, new_n18384_, new_n18385_,
    new_n18386_, new_n18387_, new_n18388_, new_n18389_, new_n18390_,
    new_n18391_, new_n18392_, new_n18393_, new_n18394_, new_n18395_,
    new_n18396_, new_n18397_, new_n18398_, new_n18399_, new_n18400_,
    new_n18401_, new_n18402_, new_n18403_, new_n18404_, new_n18405_,
    new_n18406_, new_n18407_, new_n18408_, new_n18409_, new_n18410_,
    new_n18411_, new_n18412_, new_n18413_, new_n18414_, new_n18415_,
    new_n18416_, new_n18417_, new_n18418_, new_n18419_, new_n18420_,
    new_n18421_, new_n18422_, new_n18423_, new_n18424_, new_n18425_,
    new_n18426_, new_n18427_, new_n18428_, new_n18429_, new_n18430_,
    new_n18431_, new_n18432_, new_n18433_, new_n18434_, new_n18435_,
    new_n18436_, new_n18437_, new_n18438_, new_n18439_, new_n18440_,
    new_n18441_, new_n18442_, new_n18443_, new_n18444_, new_n18445_,
    new_n18446_, new_n18447_, new_n18448_, new_n18449_, new_n18450_,
    new_n18451_, new_n18452_, new_n18453_, new_n18454_, new_n18455_,
    new_n18456_, new_n18457_, new_n18458_, new_n18459_, new_n18460_,
    new_n18461_, new_n18462_, new_n18463_, new_n18464_, new_n18465_,
    new_n18466_, new_n18467_, new_n18468_, new_n18469_, new_n18470_,
    new_n18471_, new_n18472_, new_n18473_, new_n18474_, new_n18475_,
    new_n18476_, new_n18477_, new_n18478_, new_n18479_, new_n18480_,
    new_n18481_, new_n18482_, new_n18483_, new_n18484_, new_n18485_,
    new_n18486_, new_n18487_, new_n18488_, new_n18489_, new_n18490_,
    new_n18491_, new_n18492_, new_n18493_, new_n18494_, new_n18495_,
    new_n18496_, new_n18497_, new_n18498_, new_n18499_, new_n18500_,
    new_n18501_, new_n18502_, new_n18503_, new_n18504_, new_n18505_,
    new_n18506_, new_n18507_, new_n18508_, new_n18509_, new_n18510_,
    new_n18511_, new_n18512_, new_n18513_, new_n18514_, new_n18515_,
    new_n18516_, new_n18517_, new_n18518_, new_n18519_, new_n18520_,
    new_n18521_, new_n18522_, new_n18523_, new_n18524_, new_n18525_,
    new_n18526_, new_n18527_, new_n18528_, new_n18529_, new_n18530_,
    new_n18531_, new_n18532_, new_n18533_, new_n18534_, new_n18535_,
    new_n18536_, new_n18537_, new_n18538_, new_n18539_, new_n18540_,
    new_n18541_, new_n18542_, new_n18543_, new_n18544_, new_n18545_,
    new_n18546_, new_n18547_, new_n18548_, new_n18549_, new_n18550_,
    new_n18551_, new_n18552_, new_n18553_, new_n18554_, new_n18555_,
    new_n18556_, new_n18557_, new_n18558_, new_n18559_, new_n18560_,
    new_n18561_, new_n18562_, new_n18563_, new_n18564_, new_n18565_,
    new_n18566_, new_n18567_, new_n18568_, new_n18569_, new_n18570_,
    new_n18571_, new_n18572_, new_n18573_, new_n18574_, new_n18575_,
    new_n18576_, new_n18577_, new_n18578_, new_n18579_, new_n18580_,
    new_n18581_, new_n18582_, new_n18583_, new_n18584_, new_n18585_,
    new_n18586_, new_n18587_, new_n18588_, new_n18589_, new_n18590_,
    new_n18591_, new_n18592_, new_n18593_, new_n18594_, new_n18595_,
    new_n18596_, new_n18597_, new_n18598_, new_n18599_, new_n18600_,
    new_n18601_, new_n18602_, new_n18603_, new_n18604_, new_n18605_,
    new_n18606_, new_n18607_, new_n18608_, new_n18609_, new_n18610_,
    new_n18611_, new_n18612_, new_n18613_, new_n18614_, new_n18615_,
    new_n18616_, new_n18617_, new_n18618_, new_n18619_, new_n18620_,
    new_n18621_, new_n18622_, new_n18623_, new_n18624_, new_n18625_,
    new_n18626_, new_n18627_, new_n18628_, new_n18629_, new_n18630_,
    new_n18631_, new_n18632_, new_n18633_, new_n18634_, new_n18635_,
    new_n18636_, new_n18637_, new_n18638_, new_n18639_, new_n18640_,
    new_n18641_, new_n18642_, new_n18643_, new_n18644_, new_n18645_,
    new_n18646_, new_n18647_, new_n18648_, new_n18649_, new_n18650_,
    new_n18651_, new_n18652_, new_n18653_, new_n18654_, new_n18655_,
    new_n18656_, new_n18657_, new_n18658_, new_n18659_, new_n18660_,
    new_n18661_, new_n18662_, new_n18663_, new_n18664_, new_n18665_,
    new_n18666_, new_n18667_, new_n18668_, new_n18669_, new_n18670_,
    new_n18671_, new_n18672_, new_n18673_, new_n18674_, new_n18675_,
    new_n18676_, new_n18677_, new_n18678_, new_n18679_, new_n18680_,
    new_n18681_, new_n18682_, new_n18683_, new_n18684_, new_n18685_,
    new_n18686_, new_n18687_, new_n18688_, new_n18689_, new_n18690_,
    new_n18691_, new_n18692_, new_n18693_, new_n18694_, new_n18695_,
    new_n18696_, new_n18697_, new_n18698_, new_n18699_, new_n18700_,
    new_n18701_, new_n18702_, new_n18703_, new_n18704_, new_n18705_,
    new_n18706_, new_n18707_, new_n18708_, new_n18709_, new_n18710_,
    new_n18711_, new_n18712_, new_n18713_, new_n18714_, new_n18715_,
    new_n18716_, new_n18717_, new_n18718_, new_n18719_, new_n18720_,
    new_n18721_, new_n18722_, new_n18723_, new_n18724_, new_n18725_,
    new_n18726_, new_n18727_, new_n18728_, new_n18729_, new_n18730_,
    new_n18731_, new_n18732_, new_n18733_, new_n18734_, new_n18735_,
    new_n18736_, new_n18737_, new_n18738_, new_n18739_, new_n18740_,
    new_n18741_, new_n18742_, new_n18743_, new_n18744_, new_n18745_,
    new_n18746_, new_n18747_, new_n18748_, new_n18749_, new_n18750_,
    new_n18751_, new_n18752_, new_n18753_, new_n18754_, new_n18755_,
    new_n18756_, new_n18757_, new_n18758_, new_n18759_, new_n18760_,
    new_n18761_, new_n18762_, new_n18763_, new_n18764_, new_n18765_,
    new_n18766_, new_n18767_, new_n18768_, new_n18769_, new_n18770_,
    new_n18771_, new_n18772_, new_n18773_, new_n18774_, new_n18775_,
    new_n18776_, new_n18777_, new_n18778_, new_n18779_, new_n18780_,
    new_n18781_, new_n18782_, new_n18783_, new_n18784_, new_n18785_,
    new_n18786_, new_n18787_, new_n18788_, new_n18789_, new_n18790_,
    new_n18791_, new_n18792_, new_n18793_, new_n18794_, new_n18795_,
    new_n18796_, new_n18797_, new_n18798_, new_n18799_, new_n18800_,
    new_n18801_, new_n18802_, new_n18803_, new_n18804_, new_n18805_,
    new_n18806_, new_n18807_, new_n18808_, new_n18809_, new_n18810_,
    new_n18811_, new_n18812_, new_n18813_, new_n18814_, new_n18815_,
    new_n18816_, new_n18817_, new_n18818_, new_n18819_, new_n18820_,
    new_n18821_, new_n18822_, new_n18823_, new_n18824_, new_n18825_,
    new_n18826_, new_n18827_, new_n18828_, new_n18829_, new_n18830_,
    new_n18831_, new_n18832_, new_n18833_, new_n18834_, new_n18835_,
    new_n18836_, new_n18837_, new_n18838_, new_n18839_, new_n18840_,
    new_n18841_, new_n18842_, new_n18843_, new_n18844_, new_n18845_,
    new_n18846_, new_n18847_, new_n18848_, new_n18849_, new_n18850_,
    new_n18851_, new_n18852_, new_n18853_, new_n18854_, new_n18855_,
    new_n18856_, new_n18857_, new_n18858_, new_n18859_, new_n18860_,
    new_n18861_, new_n18862_, new_n18863_, new_n18864_, new_n18865_,
    new_n18866_, new_n18867_, new_n18868_, new_n18869_, new_n18870_,
    new_n18871_, new_n18872_, new_n18873_, new_n18874_, new_n18875_,
    new_n18876_, new_n18877_, new_n18878_, new_n18879_, new_n18880_,
    new_n18881_, new_n18882_, new_n18883_, new_n18884_, new_n18885_,
    new_n18886_, new_n18887_, new_n18888_, new_n18889_, new_n18890_,
    new_n18891_, new_n18892_, new_n18893_, new_n18894_, new_n18895_,
    new_n18896_, new_n18897_, new_n18898_, new_n18899_, new_n18900_,
    new_n18901_, new_n18902_, new_n18903_, new_n18904_, new_n18905_,
    new_n18906_, new_n18907_, new_n18908_, new_n18909_, new_n18910_,
    new_n18911_, new_n18912_, new_n18913_, new_n18914_, new_n18915_,
    new_n18916_, new_n18917_, new_n18918_, new_n18919_, new_n18920_,
    new_n18921_, new_n18922_, new_n18923_, new_n18924_, new_n18925_,
    new_n18926_, new_n18927_, new_n18928_, new_n18929_, new_n18930_,
    new_n18931_, new_n18932_, new_n18933_, new_n18934_, new_n18935_,
    new_n18936_, new_n18937_, new_n18938_, new_n18939_, new_n18940_,
    new_n18941_, new_n18942_, new_n18943_, new_n18944_, new_n18945_,
    new_n18946_, new_n18947_, new_n18948_, new_n18949_, new_n18950_,
    new_n18951_, new_n18952_, new_n18953_, new_n18954_, new_n18955_,
    new_n18956_, new_n18957_, new_n18958_, new_n18959_, new_n18960_,
    new_n18961_, new_n18962_, new_n18963_, new_n18964_, new_n18965_,
    new_n18966_, new_n18967_, new_n18968_, new_n18969_, new_n18970_,
    new_n18971_, new_n18972_, new_n18973_, new_n18974_, new_n18975_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19028_, new_n19029_, new_n19030_, new_n19031_,
    new_n19032_, new_n19033_, new_n19034_, new_n19035_, new_n19036_,
    new_n19037_, new_n19038_, new_n19039_, new_n19040_, new_n19041_,
    new_n19042_, new_n19043_, new_n19044_, new_n19045_, new_n19046_,
    new_n19047_, new_n19048_, new_n19049_, new_n19050_, new_n19051_,
    new_n19052_, new_n19053_, new_n19054_, new_n19055_, new_n19056_,
    new_n19057_, new_n19058_, new_n19059_, new_n19060_, new_n19061_,
    new_n19062_, new_n19063_, new_n19064_, new_n19065_, new_n19066_,
    new_n19067_, new_n19068_, new_n19069_, new_n19070_, new_n19071_,
    new_n19072_, new_n19073_, new_n19074_, new_n19075_, new_n19076_,
    new_n19077_, new_n19078_, new_n19079_, new_n19080_, new_n19081_,
    new_n19082_, new_n19083_, new_n19084_, new_n19085_, new_n19086_,
    new_n19087_, new_n19088_, new_n19089_, new_n19090_, new_n19091_,
    new_n19092_, new_n19093_, new_n19094_, new_n19095_, new_n19096_,
    new_n19097_, new_n19098_, new_n19099_, new_n19100_, new_n19101_,
    new_n19102_, new_n19103_, new_n19104_, new_n19105_, new_n19106_,
    new_n19107_, new_n19108_, new_n19109_, new_n19110_, new_n19111_,
    new_n19112_, new_n19113_, new_n19114_, new_n19115_, new_n19116_,
    new_n19117_, new_n19118_, new_n19119_, new_n19120_, new_n19121_,
    new_n19122_, new_n19123_, new_n19124_, new_n19125_, new_n19126_,
    new_n19127_, new_n19128_, new_n19129_, new_n19130_, new_n19131_,
    new_n19132_, new_n19133_, new_n19134_, new_n19135_, new_n19136_,
    new_n19137_, new_n19138_, new_n19139_, new_n19140_, new_n19141_,
    new_n19142_, new_n19143_, new_n19144_, new_n19145_, new_n19146_,
    new_n19147_, new_n19148_, new_n19149_, new_n19150_, new_n19151_,
    new_n19152_, new_n19153_, new_n19154_, new_n19155_, new_n19156_,
    new_n19157_, new_n19158_, new_n19159_, new_n19160_, new_n19161_,
    new_n19162_, new_n19163_, new_n19164_, new_n19165_, new_n19166_,
    new_n19167_, new_n19168_, new_n19169_, new_n19170_, new_n19171_,
    new_n19172_, new_n19173_, new_n19174_, new_n19175_, new_n19176_,
    new_n19177_, new_n19178_, new_n19179_, new_n19180_, new_n19181_,
    new_n19182_, new_n19183_, new_n19184_, new_n19185_, new_n19186_,
    new_n19187_, new_n19188_, new_n19189_, new_n19190_, new_n19191_,
    new_n19192_, new_n19193_, new_n19194_, new_n19195_, new_n19196_,
    new_n19197_, new_n19198_, new_n19199_, new_n19200_, new_n19201_,
    new_n19202_, new_n19203_, new_n19204_, new_n19205_, new_n19206_,
    new_n19207_, new_n19208_, new_n19209_, new_n19210_, new_n19211_,
    new_n19212_, new_n19213_, new_n19214_, new_n19215_, new_n19216_,
    new_n19217_, new_n19218_, new_n19219_, new_n19220_, new_n19221_,
    new_n19222_, new_n19223_, new_n19224_, new_n19225_, new_n19226_,
    new_n19227_, new_n19228_, new_n19229_, new_n19230_, new_n19231_,
    new_n19232_, new_n19233_, new_n19234_, new_n19235_, new_n19236_,
    new_n19237_, new_n19238_, new_n19239_, new_n19240_, new_n19241_,
    new_n19242_, new_n19243_, new_n19244_, new_n19245_, new_n19246_,
    new_n19247_, new_n19248_, new_n19249_, new_n19250_, new_n19251_,
    new_n19252_, new_n19253_, new_n19254_, new_n19255_, new_n19256_,
    new_n19257_, new_n19258_, new_n19259_, new_n19260_, new_n19261_,
    new_n19262_, new_n19263_, new_n19264_, new_n19265_, new_n19266_,
    new_n19267_, new_n19268_, new_n19269_, new_n19270_, new_n19271_,
    new_n19272_, new_n19273_, new_n19274_, new_n19275_, new_n19276_,
    new_n19277_, new_n19278_, new_n19279_, new_n19280_, new_n19281_,
    new_n19282_, new_n19283_, new_n19284_, new_n19285_, new_n19286_,
    new_n19287_, new_n19288_, new_n19289_, new_n19290_, new_n19291_,
    new_n19292_, new_n19293_, new_n19294_, new_n19295_, new_n19296_,
    new_n19297_, new_n19298_, new_n19299_, new_n19300_, new_n19301_,
    new_n19302_, new_n19303_, new_n19304_, new_n19305_, new_n19306_,
    new_n19307_, new_n19308_, new_n19309_, new_n19310_, new_n19311_,
    new_n19312_, new_n19313_, new_n19314_, new_n19315_, new_n19316_,
    new_n19317_, new_n19318_, new_n19319_, new_n19320_, new_n19321_,
    new_n19322_, new_n19323_, new_n19324_, new_n19325_, new_n19326_,
    new_n19327_, new_n19328_, new_n19329_, new_n19330_, new_n19331_,
    new_n19332_, new_n19333_, new_n19334_, new_n19335_, new_n19336_,
    new_n19337_, new_n19338_, new_n19339_, new_n19340_, new_n19341_,
    new_n19342_, new_n19343_, new_n19344_, new_n19345_, new_n19346_,
    new_n19347_, new_n19348_, new_n19349_, new_n19350_, new_n19351_,
    new_n19352_, new_n19353_, new_n19354_, new_n19355_, new_n19356_,
    new_n19357_, new_n19358_, new_n19359_, new_n19360_, new_n19361_,
    new_n19362_, new_n19363_, new_n19364_, new_n19365_, new_n19366_,
    new_n19367_, new_n19368_, new_n19369_, new_n19370_, new_n19371_,
    new_n19372_, new_n19373_, new_n19374_, new_n19375_, new_n19376_,
    new_n19377_, new_n19378_, new_n19379_, new_n19380_, new_n19381_,
    new_n19382_, new_n19383_, new_n19384_, new_n19385_, new_n19386_,
    new_n19387_, new_n19388_, new_n19389_, new_n19390_, new_n19391_,
    new_n19392_, new_n19393_, new_n19394_, new_n19395_, new_n19396_,
    new_n19397_, new_n19398_, new_n19399_, new_n19400_, new_n19401_,
    new_n19402_, new_n19403_, new_n19404_, new_n19405_, new_n19406_,
    new_n19407_, new_n19408_, new_n19409_, new_n19410_, new_n19411_,
    new_n19412_, new_n19413_, new_n19414_, new_n19415_, new_n19416_,
    new_n19417_, new_n19418_, new_n19419_, new_n19420_, new_n19421_,
    new_n19423_, new_n19424_, new_n19425_, new_n19426_, new_n19427_,
    new_n19428_, new_n19429_, new_n19430_, new_n19431_, new_n19432_,
    new_n19433_, new_n19434_, new_n19435_, new_n19436_, new_n19437_,
    new_n19438_, new_n19439_, new_n19440_, new_n19441_, new_n19442_,
    new_n19443_, new_n19444_, new_n19445_, new_n19446_, new_n19447_,
    new_n19448_, new_n19449_, new_n19450_, new_n19451_, new_n19452_,
    new_n19453_, new_n19454_, new_n19455_, new_n19456_, new_n19457_,
    new_n19458_, new_n19459_, new_n19460_, new_n19461_, new_n19462_,
    new_n19463_, new_n19464_, new_n19465_, new_n19466_, new_n19467_,
    new_n19468_, new_n19469_, new_n19470_, new_n19471_, new_n19472_,
    new_n19473_, new_n19474_, new_n19475_, new_n19476_, new_n19477_,
    new_n19478_, new_n19479_, new_n19480_, new_n19481_, new_n19482_,
    new_n19483_, new_n19484_, new_n19485_, new_n19486_, new_n19487_,
    new_n19488_, new_n19489_, new_n19490_, new_n19491_, new_n19492_,
    new_n19493_, new_n19494_, new_n19495_, new_n19496_, new_n19497_,
    new_n19498_, new_n19499_, new_n19500_, new_n19501_, new_n19502_,
    new_n19503_, new_n19504_, new_n19505_, new_n19506_, new_n19507_,
    new_n19508_, new_n19509_, new_n19510_, new_n19511_, new_n19512_,
    new_n19513_, new_n19514_, new_n19515_, new_n19516_, new_n19517_,
    new_n19518_, new_n19519_, new_n19520_, new_n19521_, new_n19522_,
    new_n19523_, new_n19524_, new_n19525_, new_n19526_, new_n19527_,
    new_n19528_, new_n19529_, new_n19530_, new_n19531_, new_n19532_,
    new_n19533_, new_n19534_, new_n19535_, new_n19536_, new_n19537_,
    new_n19538_, new_n19539_, new_n19540_, new_n19541_, new_n19542_,
    new_n19543_, new_n19544_, new_n19545_, new_n19546_, new_n19547_,
    new_n19548_, new_n19549_, new_n19550_, new_n19551_, new_n19552_,
    new_n19553_, new_n19554_, new_n19555_, new_n19556_, new_n19557_,
    new_n19558_, new_n19559_, new_n19560_, new_n19561_, new_n19562_,
    new_n19563_, new_n19564_, new_n19565_, new_n19566_, new_n19567_,
    new_n19568_, new_n19569_, new_n19570_, new_n19571_, new_n19572_,
    new_n19573_, new_n19574_, new_n19575_, new_n19576_, new_n19577_,
    new_n19578_, new_n19579_, new_n19580_, new_n19581_, new_n19582_,
    new_n19583_, new_n19584_, new_n19585_, new_n19586_, new_n19587_,
    new_n19588_, new_n19589_, new_n19590_, new_n19591_, new_n19592_,
    new_n19593_, new_n19594_, new_n19595_, new_n19596_, new_n19597_,
    new_n19598_, new_n19599_, new_n19600_, new_n19601_, new_n19602_,
    new_n19603_, new_n19604_, new_n19605_, new_n19606_, new_n19607_,
    new_n19608_, new_n19609_, new_n19610_, new_n19611_, new_n19612_,
    new_n19613_, new_n19614_, new_n19615_, new_n19616_, new_n19617_,
    new_n19618_, new_n19619_, new_n19620_, new_n19621_, new_n19622_,
    new_n19623_, new_n19624_, new_n19625_, new_n19626_, new_n19627_,
    new_n19628_, new_n19629_, new_n19630_, new_n19631_, new_n19632_,
    new_n19633_, new_n19634_, new_n19635_, new_n19636_, new_n19637_,
    new_n19638_, new_n19639_, new_n19640_, new_n19641_, new_n19642_,
    new_n19643_, new_n19644_, new_n19645_, new_n19646_, new_n19647_,
    new_n19648_, new_n19649_, new_n19650_, new_n19651_, new_n19652_,
    new_n19653_, new_n19654_, new_n19655_, new_n19656_, new_n19657_,
    new_n19658_, new_n19659_, new_n19660_, new_n19661_, new_n19662_,
    new_n19663_, new_n19664_, new_n19665_, new_n19666_, new_n19667_,
    new_n19668_, new_n19669_, new_n19670_, new_n19671_, new_n19672_,
    new_n19673_, new_n19674_, new_n19675_, new_n19676_, new_n19677_,
    new_n19678_, new_n19679_, new_n19680_, new_n19681_, new_n19682_,
    new_n19683_, new_n19684_, new_n19685_, new_n19686_, new_n19687_,
    new_n19688_, new_n19689_, new_n19690_, new_n19691_, new_n19692_,
    new_n19693_, new_n19694_, new_n19695_, new_n19696_, new_n19697_,
    new_n19698_, new_n19699_, new_n19700_, new_n19701_, new_n19702_,
    new_n19703_, new_n19704_, new_n19705_, new_n19706_, new_n19707_,
    new_n19708_, new_n19709_, new_n19710_, new_n19711_, new_n19712_,
    new_n19713_, new_n19714_, new_n19715_, new_n19716_, new_n19717_,
    new_n19718_, new_n19719_, new_n19720_, new_n19721_, new_n19722_,
    new_n19723_, new_n19724_, new_n19725_, new_n19726_, new_n19727_,
    new_n19728_, new_n19729_, new_n19730_, new_n19731_, new_n19732_,
    new_n19733_, new_n19734_, new_n19735_, new_n19736_, new_n19737_,
    new_n19738_, new_n19739_, new_n19740_, new_n19741_, new_n19742_,
    new_n19743_, new_n19744_, new_n19745_, new_n19746_, new_n19747_,
    new_n19748_, new_n19749_, new_n19750_, new_n19751_, new_n19752_,
    new_n19753_, new_n19754_, new_n19755_, new_n19756_, new_n19757_,
    new_n19758_, new_n19759_, new_n19760_, new_n19761_, new_n19762_,
    new_n19763_, new_n19764_, new_n19765_, new_n19766_, new_n19767_,
    new_n19768_, new_n19769_, new_n19770_, new_n19771_, new_n19772_,
    new_n19773_, new_n19774_, new_n19775_, new_n19776_, new_n19777_,
    new_n19778_, new_n19779_, new_n19780_, new_n19781_, new_n19782_,
    new_n19783_, new_n19784_, new_n19785_, new_n19786_, new_n19787_,
    new_n19788_, new_n19789_, new_n19790_, new_n19791_, new_n19792_,
    new_n19793_, new_n19794_, new_n19795_, new_n19796_, new_n19797_,
    new_n19798_, new_n19799_, new_n19800_, new_n19801_, new_n19802_,
    new_n19803_, new_n19804_, new_n19805_, new_n19806_, new_n19807_,
    new_n19808_, new_n19809_, new_n19810_, new_n19811_, new_n19812_,
    new_n19813_, new_n19814_, new_n19815_, new_n19816_, new_n19817_,
    new_n19818_, new_n19819_, new_n19820_, new_n19821_, new_n19822_,
    new_n19823_, new_n19824_, new_n19825_, new_n19826_, new_n19827_,
    new_n19828_, new_n19829_, new_n19830_, new_n19831_, new_n19832_,
    new_n19833_, new_n19834_, new_n19835_, new_n19836_, new_n19837_,
    new_n19838_, new_n19839_, new_n19840_, new_n19841_, new_n19842_,
    new_n19843_, new_n19844_, new_n19845_, new_n19846_, new_n19847_,
    new_n19848_, new_n19849_, new_n19850_, new_n19851_, new_n19852_,
    new_n19853_, new_n19854_, new_n19855_, new_n19856_, new_n19857_,
    new_n19858_, new_n19859_, new_n19860_, new_n19861_, new_n19862_,
    new_n19863_, new_n19864_, new_n19865_, new_n19866_, new_n19867_,
    new_n19868_, new_n19869_, new_n19870_, new_n19871_, new_n19872_,
    new_n19873_, new_n19874_, new_n19875_, new_n19876_, new_n19877_,
    new_n19878_, new_n19879_, new_n19880_, new_n19881_, new_n19882_,
    new_n19883_, new_n19884_, new_n19885_, new_n19886_, new_n19887_,
    new_n19888_, new_n19889_, new_n19890_, new_n19891_, new_n19892_,
    new_n19893_, new_n19894_, new_n19895_, new_n19896_, new_n19897_,
    new_n19898_, new_n19899_, new_n19900_, new_n19901_, new_n19902_,
    new_n19903_, new_n19904_, new_n19905_, new_n19906_, new_n19907_,
    new_n19908_, new_n19909_, new_n19910_, new_n19911_, new_n19912_,
    new_n19913_, new_n19914_, new_n19915_, new_n19916_, new_n19917_,
    new_n19918_, new_n19919_, new_n19920_, new_n19921_, new_n19922_,
    new_n19923_, new_n19924_, new_n19925_, new_n19926_, new_n19927_,
    new_n19928_, new_n19929_, new_n19930_, new_n19931_, new_n19932_,
    new_n19933_, new_n19934_, new_n19935_, new_n19936_, new_n19937_,
    new_n19938_;
  NOR2_X1    g00000(.A1(\a[126] ), .A2(\a[127] ), .ZN(new_n193_));
  INV_X1     g00001(.I(\a[65] ), .ZN(new_n194_));
  INV_X1     g00002(.I(\a[126] ), .ZN(new_n195_));
  OAI21_X1   g00003(.A1(\a[124] ), .A2(\a[125] ), .B(new_n195_), .ZN(new_n196_));
  INV_X1     g00004(.I(\a[127] ), .ZN(new_n197_));
  NOR2_X1    g00005(.A1(new_n195_), .A2(new_n197_), .ZN(new_n198_));
  INV_X1     g00006(.I(new_n198_), .ZN(new_n199_));
  NAND2_X1   g00007(.A1(new_n199_), .A2(new_n196_), .ZN(\asqrt[62] ));
  INV_X1     g00008(.I(\asqrt[62] ), .ZN(new_n201_));
  INV_X1     g00009(.I(\a[111] ), .ZN(new_n202_));
  INV_X1     g00010(.I(\a[119] ), .ZN(new_n203_));
  INV_X1     g00011(.I(new_n193_), .ZN(\asqrt[63] ));
  NOR2_X1    g00012(.A1(\a[124] ), .A2(\a[126] ), .ZN(new_n205_));
  INV_X1     g00013(.I(\a[124] ), .ZN(new_n206_));
  INV_X1     g00014(.I(\a[125] ), .ZN(new_n207_));
  NAND3_X1   g00015(.A1(new_n206_), .A2(new_n207_), .A3(\a[127] ), .ZN(new_n208_));
  OAI21_X1   g00016(.A1(new_n197_), .A2(\a[124] ), .B(\a[125] ), .ZN(new_n209_));
  AOI21_X1   g00017(.A1(new_n208_), .A2(new_n209_), .B(new_n205_), .ZN(new_n210_));
  NAND3_X1   g00018(.A1(new_n206_), .A2(new_n197_), .A3(\a[126] ), .ZN(new_n211_));
  OR3_X2     g00019(.A1(\a[122] ), .A2(\a[123] ), .A3(\a[124] ), .Z(new_n212_));
  NAND2_X1   g00020(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  AOI21_X1   g00021(.A1(new_n210_), .A2(new_n213_), .B(\asqrt[63] ), .ZN(new_n214_));
  NAND3_X1   g00022(.A1(new_n206_), .A2(new_n207_), .A3(\a[126] ), .ZN(new_n215_));
  AOI21_X1   g00023(.A1(new_n196_), .A2(new_n215_), .B(\a[127] ), .ZN(new_n216_));
  INV_X1     g00024(.I(new_n216_), .ZN(new_n217_));
  INV_X1     g00025(.I(new_n205_), .ZN(new_n218_));
  NOR3_X1    g00026(.A1(new_n197_), .A2(\a[124] ), .A3(\a[125] ), .ZN(new_n219_));
  AOI21_X1   g00027(.A1(new_n206_), .A2(\a[127] ), .B(new_n207_), .ZN(new_n220_));
  OAI21_X1   g00028(.A1(new_n220_), .A2(new_n219_), .B(new_n218_), .ZN(new_n221_));
  NOR2_X1    g00029(.A1(new_n195_), .A2(\a[124] ), .ZN(new_n222_));
  NOR2_X1    g00030(.A1(\a[122] ), .A2(\a[123] ), .ZN(new_n223_));
  AOI22_X1   g00031(.A1(new_n222_), .A2(new_n197_), .B1(new_n206_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1   g00032(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1   g00033(.A1(new_n214_), .A2(new_n225_), .A3(new_n217_), .ZN(\asqrt[61] ));
  INV_X1     g00034(.I(\a[120] ), .ZN(new_n227_));
  NOR2_X1    g00035(.A1(\a[118] ), .A2(\a[119] ), .ZN(new_n228_));
  NAND2_X1   g00036(.A1(new_n210_), .A2(new_n213_), .ZN(new_n229_));
  INV_X1     g00037(.I(new_n229_), .ZN(new_n230_));
  NOR2_X1    g00038(.A1(new_n210_), .A2(new_n213_), .ZN(new_n231_));
  AOI21_X1   g00039(.A1(\asqrt[61] ), .A2(new_n230_), .B(new_n231_), .ZN(new_n232_));
  NAND4_X1   g00040(.A1(new_n214_), .A2(new_n225_), .A3(new_n217_), .A4(\asqrt[62] ), .ZN(new_n233_));
  NAND2_X1   g00041(.A1(\asqrt[61] ), .A2(new_n223_), .ZN(new_n234_));
  AOI21_X1   g00042(.A1(new_n234_), .A2(new_n233_), .B(\a[124] ), .ZN(new_n235_));
  OAI21_X1   g00043(.A1(new_n221_), .A2(new_n224_), .B(new_n193_), .ZN(new_n236_));
  NOR4_X1    g00044(.A1(new_n236_), .A2(new_n201_), .A3(new_n231_), .A4(new_n216_), .ZN(new_n237_));
  INV_X1     g00045(.I(new_n223_), .ZN(new_n238_));
  NOR3_X1    g00046(.A1(new_n236_), .A2(new_n231_), .A3(new_n216_), .ZN(new_n239_));
  NOR2_X1    g00047(.A1(new_n239_), .A2(new_n238_), .ZN(new_n240_));
  NOR3_X1    g00048(.A1(new_n240_), .A2(new_n206_), .A3(new_n237_), .ZN(new_n241_));
  NOR2_X1    g00049(.A1(new_n241_), .A2(new_n235_), .ZN(new_n242_));
  INV_X1     g00050(.I(\a[122] ), .ZN(new_n243_));
  INV_X1     g00051(.I(\a[121] ), .ZN(new_n244_));
  NAND2_X1   g00052(.A1(new_n227_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1   g00053(.A1(new_n199_), .A2(new_n243_), .A3(new_n196_), .A4(new_n245_), .ZN(new_n246_));
  NOR2_X1    g00054(.A1(\asqrt[61] ), .A2(new_n246_), .ZN(new_n247_));
  INV_X1     g00055(.I(\a[123] ), .ZN(new_n248_));
  OAI21_X1   g00056(.A1(new_n239_), .A2(\a[122] ), .B(new_n248_), .ZN(new_n249_));
  NAND3_X1   g00057(.A1(\asqrt[61] ), .A2(new_n243_), .A3(\a[123] ), .ZN(new_n250_));
  AOI21_X1   g00058(.A1(new_n249_), .A2(new_n250_), .B(new_n247_), .ZN(new_n251_));
  NOR2_X1    g00059(.A1(new_n251_), .A2(\asqrt[62] ), .ZN(new_n252_));
  AOI21_X1   g00060(.A1(new_n252_), .A2(new_n242_), .B(new_n232_), .ZN(new_n253_));
  OAI21_X1   g00061(.A1(new_n240_), .A2(new_n237_), .B(new_n206_), .ZN(new_n254_));
  NAND3_X1   g00062(.A1(new_n234_), .A2(\a[124] ), .A3(new_n233_), .ZN(new_n255_));
  OR4_X2     g00063(.A1(new_n236_), .A2(new_n216_), .A3(new_n231_), .A4(new_n246_), .Z(new_n256_));
  AOI21_X1   g00064(.A1(\asqrt[61] ), .A2(new_n243_), .B(\a[123] ), .ZN(new_n257_));
  NOR3_X1    g00065(.A1(new_n239_), .A2(\a[122] ), .A3(new_n248_), .ZN(new_n258_));
  OAI21_X1   g00066(.A1(new_n258_), .A2(new_n257_), .B(new_n256_), .ZN(new_n259_));
  AOI22_X1   g00067(.A1(new_n259_), .A2(new_n201_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n260_));
  NOR2_X1    g00068(.A1(new_n221_), .A2(\asqrt[63] ), .ZN(new_n261_));
  AOI22_X1   g00069(.A1(new_n229_), .A2(new_n225_), .B1(new_n261_), .B2(new_n217_), .ZN(new_n262_));
  NOR4_X1    g00070(.A1(new_n216_), .A2(new_n210_), .A3(new_n224_), .A4(new_n193_), .ZN(new_n263_));
  NOR2_X1    g00071(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1     g00072(.I(new_n264_), .ZN(new_n265_));
  NOR4_X1    g00073(.A1(new_n253_), .A2(\asqrt[63] ), .A3(new_n260_), .A4(new_n265_), .ZN(new_n266_));
  NOR3_X1    g00074(.A1(new_n266_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n267_));
  INV_X1     g00075(.I(new_n228_), .ZN(new_n268_));
  AOI21_X1   g00076(.A1(new_n266_), .A2(\a[120] ), .B(new_n268_), .ZN(new_n269_));
  OAI21_X1   g00077(.A1(new_n267_), .A2(new_n269_), .B(\asqrt[61] ), .ZN(new_n270_));
  INV_X1     g00078(.I(new_n232_), .ZN(new_n271_));
  NAND2_X1   g00079(.A1(new_n254_), .A2(new_n255_), .ZN(new_n272_));
  NAND2_X1   g00080(.A1(new_n259_), .A2(new_n201_), .ZN(new_n273_));
  OAI21_X1   g00081(.A1(new_n273_), .A2(new_n272_), .B(new_n271_), .ZN(new_n274_));
  OAI22_X1   g00082(.A1(new_n251_), .A2(\asqrt[62] ), .B1(new_n241_), .B2(new_n235_), .ZN(new_n275_));
  NAND4_X1   g00083(.A1(new_n274_), .A2(new_n193_), .A3(new_n275_), .A4(new_n264_), .ZN(\asqrt[60] ));
  AOI21_X1   g00084(.A1(\asqrt[60] ), .A2(new_n227_), .B(new_n244_), .ZN(new_n277_));
  NOR3_X1    g00085(.A1(new_n266_), .A2(\a[120] ), .A3(\a[121] ), .ZN(new_n278_));
  NOR3_X1    g00086(.A1(new_n253_), .A2(\asqrt[63] ), .A3(new_n260_), .ZN(new_n279_));
  NAND2_X1   g00087(.A1(new_n228_), .A2(new_n227_), .ZN(new_n280_));
  NAND3_X1   g00088(.A1(new_n225_), .A2(new_n217_), .A3(new_n280_), .ZN(new_n281_));
  OAI21_X1   g00089(.A1(new_n281_), .A2(new_n236_), .B(\a[120] ), .ZN(new_n282_));
  AOI21_X1   g00090(.A1(new_n279_), .A2(new_n264_), .B(new_n282_), .ZN(new_n283_));
  NOR3_X1    g00091(.A1(new_n278_), .A2(new_n277_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1   g00092(.A1(new_n270_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1   g00093(.A1(\asqrt[60] ), .A2(\a[120] ), .A3(new_n268_), .ZN(new_n286_));
  OAI21_X1   g00094(.A1(\asqrt[60] ), .A2(new_n227_), .B(new_n228_), .ZN(new_n287_));
  AOI21_X1   g00095(.A1(new_n287_), .A2(new_n286_), .B(new_n239_), .ZN(new_n288_));
  OAI21_X1   g00096(.A1(new_n266_), .A2(\a[120] ), .B(\a[121] ), .ZN(new_n289_));
  NAND3_X1   g00097(.A1(\asqrt[60] ), .A2(new_n227_), .A3(new_n244_), .ZN(new_n290_));
  INV_X1     g00098(.I(new_n282_), .ZN(new_n291_));
  NAND2_X1   g00099(.A1(\asqrt[60] ), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1   g00100(.A1(new_n289_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  OAI21_X1   g00101(.A1(new_n288_), .A2(new_n293_), .B(new_n201_), .ZN(new_n294_));
  NAND3_X1   g00102(.A1(new_n270_), .A2(new_n284_), .A3(\asqrt[62] ), .ZN(new_n295_));
  NAND2_X1   g00103(.A1(new_n274_), .A2(new_n193_), .ZN(new_n296_));
  NOR4_X1    g00104(.A1(new_n296_), .A2(new_n239_), .A3(new_n260_), .A4(new_n265_), .ZN(new_n297_));
  NOR2_X1    g00105(.A1(new_n266_), .A2(new_n245_), .ZN(new_n298_));
  OAI21_X1   g00106(.A1(new_n298_), .A2(new_n297_), .B(new_n243_), .ZN(new_n299_));
  NAND3_X1   g00107(.A1(new_n279_), .A2(\asqrt[61] ), .A3(new_n264_), .ZN(new_n300_));
  NAND3_X1   g00108(.A1(\asqrt[60] ), .A2(new_n227_), .A3(new_n244_), .ZN(new_n301_));
  NAND3_X1   g00109(.A1(new_n301_), .A2(new_n300_), .A3(\a[122] ), .ZN(new_n302_));
  NAND2_X1   g00110(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  AOI22_X1   g00111(.A1(new_n295_), .A2(new_n294_), .B1(new_n285_), .B2(new_n303_), .ZN(new_n304_));
  NOR2_X1    g00112(.A1(new_n258_), .A2(new_n257_), .ZN(new_n305_));
  INV_X1     g00113(.I(new_n305_), .ZN(new_n306_));
  NOR3_X1    g00114(.A1(new_n266_), .A2(\asqrt[62] ), .A3(new_n247_), .ZN(new_n307_));
  NAND3_X1   g00115(.A1(new_n306_), .A2(new_n201_), .A3(new_n256_), .ZN(new_n308_));
  OAI22_X1   g00116(.A1(new_n307_), .A2(new_n306_), .B1(new_n266_), .B2(new_n308_), .ZN(new_n309_));
  NOR3_X1    g00117(.A1(\asqrt[60] ), .A2(new_n242_), .A3(new_n273_), .ZN(new_n310_));
  NOR2_X1    g00118(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1   g00119(.A1(new_n304_), .A2(new_n311_), .B(new_n193_), .ZN(new_n312_));
  AOI21_X1   g00120(.A1(new_n301_), .A2(new_n300_), .B(\a[122] ), .ZN(new_n313_));
  NOR3_X1    g00121(.A1(new_n298_), .A2(new_n297_), .A3(new_n243_), .ZN(new_n314_));
  NOR2_X1    g00122(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1   g00123(.A1(new_n285_), .A2(\asqrt[62] ), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1   g00124(.A1(new_n285_), .A2(\asqrt[62] ), .ZN(new_n317_));
  NAND3_X1   g00125(.A1(new_n316_), .A2(new_n309_), .A3(new_n317_), .ZN(new_n318_));
  NOR2_X1    g00126(.A1(\asqrt[60] ), .A2(new_n272_), .ZN(new_n319_));
  XOR2_X1    g00127(.A1(new_n252_), .A2(new_n242_), .Z(new_n320_));
  NAND2_X1   g00128(.A1(new_n320_), .A2(\asqrt[63] ), .ZN(new_n321_));
  NOR2_X1    g00129(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1   g00130(.A1(new_n252_), .A2(new_n272_), .A3(new_n264_), .ZN(new_n323_));
  NOR2_X1    g00131(.A1(new_n296_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1    g00132(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1   g00133(.A1(new_n312_), .A2(new_n318_), .A3(new_n325_), .ZN(\asqrt[59] ));
  NOR2_X1    g00134(.A1(new_n288_), .A2(new_n293_), .ZN(new_n327_));
  AOI21_X1   g00135(.A1(new_n270_), .A2(new_n284_), .B(\asqrt[62] ), .ZN(new_n328_));
  NOR3_X1    g00136(.A1(new_n288_), .A2(new_n293_), .A3(new_n201_), .ZN(new_n329_));
  OAI22_X1   g00137(.A1(new_n328_), .A2(new_n329_), .B1(new_n327_), .B2(new_n315_), .ZN(new_n330_));
  INV_X1     g00138(.I(new_n311_), .ZN(new_n331_));
  AOI21_X1   g00139(.A1(new_n330_), .A2(new_n331_), .B(\asqrt[63] ), .ZN(new_n332_));
  AOI21_X1   g00140(.A1(new_n327_), .A2(new_n201_), .B(new_n303_), .ZN(new_n333_));
  OAI21_X1   g00141(.A1(new_n327_), .A2(new_n201_), .B(new_n309_), .ZN(new_n334_));
  NOR2_X1    g00142(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1     g00143(.I(new_n325_), .ZN(new_n336_));
  NOR3_X1    g00144(.A1(new_n332_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NOR2_X1    g00145(.A1(new_n337_), .A2(\a[118] ), .ZN(new_n338_));
  INV_X1     g00146(.I(new_n338_), .ZN(new_n339_));
  NOR2_X1    g00147(.A1(new_n203_), .A2(\a[118] ), .ZN(new_n340_));
  AOI22_X1   g00148(.A1(new_n339_), .A2(new_n203_), .B1(\asqrt[59] ), .B2(new_n340_), .ZN(new_n341_));
  INV_X1     g00149(.I(new_n341_), .ZN(new_n342_));
  NOR2_X1    g00150(.A1(new_n285_), .A2(\asqrt[62] ), .ZN(new_n343_));
  INV_X1     g00151(.I(new_n317_), .ZN(new_n344_));
  OAI21_X1   g00152(.A1(new_n343_), .A2(new_n344_), .B(new_n337_), .ZN(new_n345_));
  NOR2_X1    g00153(.A1(new_n313_), .A2(new_n314_), .ZN(new_n346_));
  AND2_X2    g00154(.A1(new_n345_), .A2(new_n346_), .Z(new_n347_));
  INV_X1     g00155(.I(new_n347_), .ZN(new_n348_));
  INV_X1     g00156(.I(\a[118] ), .ZN(new_n349_));
  NOR2_X1    g00157(.A1(\a[116] ), .A2(\a[117] ), .ZN(new_n350_));
  NOR3_X1    g00158(.A1(new_n337_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1     g00159(.I(new_n350_), .ZN(new_n352_));
  AOI21_X1   g00160(.A1(new_n337_), .A2(\a[118] ), .B(new_n352_), .ZN(new_n353_));
  OAI21_X1   g00161(.A1(new_n351_), .A2(new_n353_), .B(\asqrt[60] ), .ZN(new_n354_));
  AOI21_X1   g00162(.A1(\asqrt[59] ), .A2(new_n349_), .B(new_n203_), .ZN(new_n355_));
  NOR3_X1    g00163(.A1(new_n337_), .A2(\a[118] ), .A3(\a[119] ), .ZN(new_n356_));
  INV_X1     g00164(.I(new_n296_), .ZN(new_n357_));
  NOR2_X1    g00165(.A1(new_n352_), .A2(\a[118] ), .ZN(new_n358_));
  OR3_X2     g00166(.A1(new_n262_), .A2(new_n263_), .A3(new_n358_), .Z(new_n359_));
  NOR2_X1    g00167(.A1(new_n260_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1   g00168(.A1(new_n357_), .A2(new_n360_), .B(new_n349_), .ZN(new_n361_));
  INV_X1     g00169(.I(new_n361_), .ZN(new_n362_));
  NOR2_X1    g00170(.A1(new_n337_), .A2(new_n362_), .ZN(new_n363_));
  NOR3_X1    g00171(.A1(new_n356_), .A2(new_n355_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1   g00172(.A1(new_n354_), .A2(new_n364_), .B(new_n239_), .ZN(new_n365_));
  INV_X1     g00173(.I(new_n322_), .ZN(new_n366_));
  NOR2_X1    g00174(.A1(new_n324_), .A2(new_n266_), .ZN(new_n367_));
  NAND4_X1   g00175(.A1(new_n312_), .A2(new_n318_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  INV_X1     g00176(.I(new_n368_), .ZN(new_n369_));
  NOR2_X1    g00177(.A1(new_n337_), .A2(new_n268_), .ZN(new_n370_));
  OAI21_X1   g00178(.A1(new_n370_), .A2(new_n369_), .B(new_n227_), .ZN(new_n371_));
  NAND2_X1   g00179(.A1(\asqrt[59] ), .A2(new_n228_), .ZN(new_n372_));
  NAND3_X1   g00180(.A1(new_n372_), .A2(new_n368_), .A3(\a[120] ), .ZN(new_n373_));
  NAND2_X1   g00181(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1   g00182(.A1(\asqrt[59] ), .A2(\a[118] ), .A3(new_n352_), .ZN(new_n375_));
  OAI21_X1   g00183(.A1(\asqrt[59] ), .A2(new_n349_), .B(new_n350_), .ZN(new_n376_));
  AOI21_X1   g00184(.A1(new_n376_), .A2(new_n375_), .B(new_n266_), .ZN(new_n377_));
  OAI21_X1   g00185(.A1(new_n337_), .A2(\a[118] ), .B(\a[119] ), .ZN(new_n378_));
  NAND3_X1   g00186(.A1(\asqrt[59] ), .A2(new_n349_), .A3(new_n203_), .ZN(new_n379_));
  NAND2_X1   g00187(.A1(\asqrt[59] ), .A2(new_n361_), .ZN(new_n380_));
  NAND3_X1   g00188(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NOR3_X1    g00189(.A1(new_n377_), .A2(new_n381_), .A3(\asqrt[61] ), .ZN(new_n382_));
  NOR2_X1    g00190(.A1(new_n382_), .A2(new_n374_), .ZN(new_n383_));
  NOR2_X1    g00191(.A1(new_n383_), .A2(new_n365_), .ZN(new_n384_));
  OAI21_X1   g00192(.A1(new_n377_), .A2(new_n381_), .B(\asqrt[61] ), .ZN(new_n385_));
  AOI21_X1   g00193(.A1(new_n372_), .A2(new_n368_), .B(\a[120] ), .ZN(new_n386_));
  NOR3_X1    g00194(.A1(new_n370_), .A2(new_n369_), .A3(new_n227_), .ZN(new_n387_));
  NOR2_X1    g00195(.A1(new_n387_), .A2(new_n386_), .ZN(new_n388_));
  NAND3_X1   g00196(.A1(new_n354_), .A2(new_n364_), .A3(new_n239_), .ZN(new_n389_));
  NAND2_X1   g00197(.A1(new_n389_), .A2(new_n388_), .ZN(new_n390_));
  AOI21_X1   g00198(.A1(new_n390_), .A2(new_n385_), .B(\asqrt[62] ), .ZN(new_n391_));
  NOR3_X1    g00199(.A1(new_n383_), .A2(new_n201_), .A3(new_n365_), .ZN(new_n392_));
  NOR2_X1    g00200(.A1(new_n266_), .A2(\a[120] ), .ZN(new_n393_));
  INV_X1     g00201(.I(new_n393_), .ZN(new_n394_));
  NOR2_X1    g00202(.A1(new_n244_), .A2(\a[120] ), .ZN(new_n395_));
  AOI22_X1   g00203(.A1(new_n394_), .A2(new_n244_), .B1(\asqrt[60] ), .B2(new_n395_), .ZN(new_n396_));
  INV_X1     g00204(.I(new_n396_), .ZN(new_n397_));
  NOR2_X1    g00205(.A1(new_n288_), .A2(new_n283_), .ZN(new_n398_));
  NOR2_X1    g00206(.A1(new_n337_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1    g00207(.A1(new_n399_), .A2(new_n397_), .ZN(new_n400_));
  NOR3_X1    g00208(.A1(new_n337_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n401_));
  NOR2_X1    g00209(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI22_X1   g00210(.A1(new_n391_), .A2(new_n392_), .B1(new_n384_), .B2(new_n402_), .ZN(new_n403_));
  OR2_X2     g00211(.A1(new_n304_), .A2(new_n309_), .Z(new_n404_));
  AOI21_X1   g00212(.A1(new_n337_), .A2(new_n404_), .B(new_n335_), .ZN(new_n405_));
  INV_X1     g00213(.I(new_n405_), .ZN(new_n406_));
  AOI21_X1   g00214(.A1(new_n403_), .A2(new_n348_), .B(new_n406_), .ZN(new_n407_));
  INV_X1     g00215(.I(new_n402_), .ZN(new_n408_));
  AOI21_X1   g00216(.A1(new_n384_), .A2(new_n201_), .B(new_n408_), .ZN(new_n409_));
  NOR2_X1    g00217(.A1(new_n384_), .A2(new_n201_), .ZN(new_n410_));
  NOR3_X1    g00218(.A1(new_n409_), .A2(new_n410_), .A3(new_n348_), .ZN(new_n411_));
  AOI21_X1   g00219(.A1(\asqrt[59] ), .A2(new_n304_), .B(new_n309_), .ZN(new_n412_));
  NOR3_X1    g00220(.A1(new_n412_), .A2(new_n193_), .A3(new_n335_), .ZN(new_n413_));
  NOR2_X1    g00221(.A1(new_n307_), .A2(new_n305_), .ZN(new_n414_));
  INV_X1     g00222(.I(new_n307_), .ZN(new_n415_));
  OAI22_X1   g00223(.A1(new_n415_), .A2(new_n306_), .B1(new_n296_), .B2(new_n323_), .ZN(new_n416_));
  OAI21_X1   g00224(.A1(new_n416_), .A2(new_n414_), .B(new_n366_), .ZN(new_n417_));
  NOR2_X1    g00225(.A1(new_n335_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1   g00226(.A1(new_n418_), .A2(new_n312_), .ZN(new_n419_));
  INV_X1     g00227(.I(new_n419_), .ZN(new_n420_));
  NOR2_X1    g00228(.A1(new_n413_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1     g00229(.I(new_n421_), .ZN(new_n422_));
  NOR4_X1    g00230(.A1(new_n407_), .A2(\asqrt[63] ), .A3(new_n411_), .A4(new_n422_), .ZN(new_n423_));
  NOR2_X1    g00231(.A1(new_n377_), .A2(new_n363_), .ZN(new_n424_));
  NOR2_X1    g00232(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1    g00233(.A1(new_n425_), .A2(new_n342_), .ZN(new_n426_));
  NOR3_X1    g00234(.A1(new_n423_), .A2(new_n341_), .A3(new_n424_), .ZN(new_n427_));
  NOR2_X1    g00235(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1   g00236(.A1(new_n390_), .A2(new_n385_), .ZN(new_n429_));
  OAI21_X1   g00237(.A1(new_n383_), .A2(new_n365_), .B(new_n201_), .ZN(new_n430_));
  NAND3_X1   g00238(.A1(new_n390_), .A2(\asqrt[62] ), .A3(new_n385_), .ZN(new_n431_));
  AOI22_X1   g00239(.A1(new_n430_), .A2(new_n431_), .B1(new_n429_), .B2(new_n408_), .ZN(new_n432_));
  OAI21_X1   g00240(.A1(new_n432_), .A2(new_n347_), .B(new_n405_), .ZN(new_n433_));
  NAND2_X1   g00241(.A1(new_n433_), .A2(new_n193_), .ZN(new_n434_));
  NAND2_X1   g00242(.A1(new_n419_), .A2(\asqrt[59] ), .ZN(new_n435_));
  NOR4_X1    g00243(.A1(new_n434_), .A2(new_n411_), .A3(new_n413_), .A4(new_n435_), .ZN(new_n436_));
  NOR2_X1    g00244(.A1(new_n423_), .A2(new_n352_), .ZN(new_n437_));
  OAI21_X1   g00245(.A1(new_n437_), .A2(new_n436_), .B(new_n349_), .ZN(new_n438_));
  NOR3_X1    g00246(.A1(new_n407_), .A2(\asqrt[63] ), .A3(new_n411_), .ZN(new_n439_));
  NOR2_X1    g00247(.A1(new_n413_), .A2(new_n435_), .ZN(new_n440_));
  NAND2_X1   g00248(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OAI21_X1   g00249(.A1(new_n429_), .A2(\asqrt[62] ), .B(new_n402_), .ZN(new_n442_));
  NAND2_X1   g00250(.A1(new_n429_), .A2(\asqrt[62] ), .ZN(new_n443_));
  NAND3_X1   g00251(.A1(new_n442_), .A2(new_n443_), .A3(new_n347_), .ZN(new_n444_));
  NAND4_X1   g00252(.A1(new_n433_), .A2(new_n193_), .A3(new_n444_), .A4(new_n421_), .ZN(\asqrt[58] ));
  NAND2_X1   g00253(.A1(\asqrt[58] ), .A2(new_n350_), .ZN(new_n446_));
  NAND3_X1   g00254(.A1(new_n446_), .A2(new_n441_), .A3(\a[118] ), .ZN(new_n447_));
  NAND2_X1   g00255(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1    g00256(.A1(\a[114] ), .A2(\a[115] ), .ZN(new_n449_));
  INV_X1     g00257(.I(new_n449_), .ZN(new_n450_));
  NAND3_X1   g00258(.A1(\asqrt[58] ), .A2(\a[116] ), .A3(new_n450_), .ZN(new_n451_));
  INV_X1     g00259(.I(\a[116] ), .ZN(new_n452_));
  OAI21_X1   g00260(.A1(\asqrt[58] ), .A2(new_n452_), .B(new_n449_), .ZN(new_n453_));
  AOI21_X1   g00261(.A1(new_n453_), .A2(new_n451_), .B(new_n337_), .ZN(new_n454_));
  OAI21_X1   g00262(.A1(new_n423_), .A2(\a[116] ), .B(\a[117] ), .ZN(new_n455_));
  INV_X1     g00263(.I(\a[117] ), .ZN(new_n456_));
  NAND3_X1   g00264(.A1(\asqrt[58] ), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_));
  NOR2_X1    g00265(.A1(new_n450_), .A2(\a[116] ), .ZN(new_n458_));
  NOR4_X1    g00266(.A1(new_n335_), .A2(new_n322_), .A3(new_n324_), .A4(new_n458_), .ZN(new_n459_));
  AOI21_X1   g00267(.A1(new_n459_), .A2(new_n312_), .B(new_n452_), .ZN(new_n460_));
  NAND2_X1   g00268(.A1(\asqrt[58] ), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1   g00269(.A1(new_n455_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n462_));
  NOR3_X1    g00270(.A1(new_n454_), .A2(new_n462_), .A3(\asqrt[60] ), .ZN(new_n463_));
  NOR2_X1    g00271(.A1(new_n463_), .A2(new_n448_), .ZN(new_n464_));
  NOR3_X1    g00272(.A1(new_n423_), .A2(new_n452_), .A3(new_n449_), .ZN(new_n465_));
  AOI21_X1   g00273(.A1(new_n423_), .A2(\a[116] ), .B(new_n450_), .ZN(new_n466_));
  OAI21_X1   g00274(.A1(new_n465_), .A2(new_n466_), .B(\asqrt[59] ), .ZN(new_n467_));
  AOI21_X1   g00275(.A1(\asqrt[58] ), .A2(new_n452_), .B(new_n456_), .ZN(new_n468_));
  NOR3_X1    g00276(.A1(new_n423_), .A2(\a[116] ), .A3(\a[117] ), .ZN(new_n469_));
  INV_X1     g00277(.I(new_n460_), .ZN(new_n470_));
  AOI21_X1   g00278(.A1(new_n439_), .A2(new_n421_), .B(new_n470_), .ZN(new_n471_));
  NOR3_X1    g00279(.A1(new_n469_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1   g00280(.A1(new_n467_), .A2(new_n472_), .B(new_n266_), .ZN(new_n473_));
  OAI21_X1   g00281(.A1(new_n464_), .A2(new_n473_), .B(\asqrt[61] ), .ZN(new_n474_));
  AOI21_X1   g00282(.A1(new_n446_), .A2(new_n441_), .B(\a[118] ), .ZN(new_n475_));
  NOR3_X1    g00283(.A1(new_n437_), .A2(new_n436_), .A3(new_n349_), .ZN(new_n476_));
  NOR2_X1    g00284(.A1(new_n476_), .A2(new_n475_), .ZN(new_n477_));
  NAND3_X1   g00285(.A1(new_n467_), .A2(new_n472_), .A3(new_n266_), .ZN(new_n478_));
  NAND2_X1   g00286(.A1(new_n478_), .A2(new_n477_), .ZN(new_n479_));
  OAI21_X1   g00287(.A1(new_n454_), .A2(new_n462_), .B(\asqrt[60] ), .ZN(new_n480_));
  NAND3_X1   g00288(.A1(new_n479_), .A2(new_n239_), .A3(new_n480_), .ZN(new_n481_));
  NOR2_X1    g00289(.A1(new_n429_), .A2(\asqrt[62] ), .ZN(new_n482_));
  NOR2_X1    g00290(.A1(new_n410_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1    g00291(.A1(new_n400_), .A2(new_n401_), .ZN(new_n484_));
  OAI21_X1   g00292(.A1(\asqrt[58] ), .A2(new_n483_), .B(new_n484_), .ZN(new_n485_));
  INV_X1     g00293(.I(new_n485_), .ZN(new_n486_));
  OAI21_X1   g00294(.A1(new_n448_), .A2(new_n463_), .B(new_n480_), .ZN(new_n487_));
  OAI21_X1   g00295(.A1(new_n487_), .A2(\asqrt[61] ), .B(new_n428_), .ZN(new_n488_));
  NAND2_X1   g00296(.A1(new_n488_), .A2(new_n474_), .ZN(new_n489_));
  AOI21_X1   g00297(.A1(new_n479_), .A2(new_n480_), .B(new_n239_), .ZN(new_n490_));
  INV_X1     g00298(.I(new_n428_), .ZN(new_n491_));
  AOI21_X1   g00299(.A1(new_n477_), .A2(new_n478_), .B(new_n473_), .ZN(new_n492_));
  AOI21_X1   g00300(.A1(new_n492_), .A2(new_n239_), .B(new_n491_), .ZN(new_n493_));
  OAI21_X1   g00301(.A1(new_n493_), .A2(new_n490_), .B(new_n201_), .ZN(new_n494_));
  NAND3_X1   g00302(.A1(new_n488_), .A2(\asqrt[62] ), .A3(new_n474_), .ZN(new_n495_));
  AOI21_X1   g00303(.A1(new_n385_), .A2(new_n389_), .B(\asqrt[58] ), .ZN(new_n496_));
  XOR2_X1    g00304(.A1(new_n496_), .A2(new_n388_), .Z(new_n497_));
  INV_X1     g00305(.I(new_n497_), .ZN(new_n498_));
  AOI22_X1   g00306(.A1(new_n494_), .A2(new_n495_), .B1(new_n489_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1    g00307(.A1(new_n432_), .A2(new_n347_), .ZN(new_n500_));
  OAI21_X1   g00308(.A1(\asqrt[58] ), .A2(new_n500_), .B(new_n444_), .ZN(new_n501_));
  INV_X1     g00309(.I(new_n501_), .ZN(new_n502_));
  OAI21_X1   g00310(.A1(new_n499_), .A2(new_n486_), .B(new_n502_), .ZN(new_n503_));
  OAI21_X1   g00311(.A1(new_n489_), .A2(\asqrt[62] ), .B(new_n497_), .ZN(new_n504_));
  NAND2_X1   g00312(.A1(new_n489_), .A2(\asqrt[62] ), .ZN(new_n505_));
  NAND3_X1   g00313(.A1(new_n504_), .A2(new_n505_), .A3(new_n486_), .ZN(new_n506_));
  NAND2_X1   g00314(.A1(new_n423_), .A2(new_n348_), .ZN(new_n507_));
  XOR2_X1    g00315(.A1(new_n432_), .A2(new_n347_), .Z(new_n508_));
  NAND3_X1   g00316(.A1(new_n507_), .A2(\asqrt[63] ), .A3(new_n508_), .ZN(new_n509_));
  INV_X1     g00317(.I(new_n434_), .ZN(new_n510_));
  NOR3_X1    g00318(.A1(new_n411_), .A2(new_n348_), .A3(new_n422_), .ZN(new_n511_));
  NAND2_X1   g00319(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1   g00320(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1     g00321(.I(new_n513_), .ZN(new_n514_));
  NAND4_X1   g00322(.A1(new_n503_), .A2(new_n193_), .A3(new_n506_), .A4(new_n514_), .ZN(\asqrt[57] ));
  AOI21_X1   g00323(.A1(new_n474_), .A2(new_n481_), .B(\asqrt[57] ), .ZN(new_n516_));
  XOR2_X1    g00324(.A1(new_n516_), .A2(new_n428_), .Z(new_n517_));
  NOR2_X1    g00325(.A1(new_n423_), .A2(\a[116] ), .ZN(new_n518_));
  INV_X1     g00326(.I(new_n518_), .ZN(new_n519_));
  NOR2_X1    g00327(.A1(new_n456_), .A2(\a[116] ), .ZN(new_n520_));
  AOI22_X1   g00328(.A1(new_n519_), .A2(new_n456_), .B1(\asqrt[58] ), .B2(new_n520_), .ZN(new_n521_));
  INV_X1     g00329(.I(new_n521_), .ZN(new_n522_));
  AOI21_X1   g00330(.A1(new_n428_), .A2(new_n481_), .B(new_n490_), .ZN(new_n523_));
  AOI21_X1   g00331(.A1(new_n488_), .A2(new_n474_), .B(\asqrt[62] ), .ZN(new_n524_));
  NOR3_X1    g00332(.A1(new_n493_), .A2(new_n201_), .A3(new_n490_), .ZN(new_n525_));
  OAI22_X1   g00333(.A1(new_n525_), .A2(new_n524_), .B1(new_n523_), .B2(new_n497_), .ZN(new_n526_));
  AOI21_X1   g00334(.A1(new_n526_), .A2(new_n485_), .B(new_n501_), .ZN(new_n527_));
  AOI21_X1   g00335(.A1(new_n523_), .A2(new_n201_), .B(new_n498_), .ZN(new_n528_));
  OAI21_X1   g00336(.A1(new_n523_), .A2(new_n201_), .B(new_n486_), .ZN(new_n529_));
  NOR2_X1    g00337(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR4_X1    g00338(.A1(new_n527_), .A2(\asqrt[63] ), .A3(new_n530_), .A4(new_n513_), .ZN(new_n531_));
  NOR2_X1    g00339(.A1(new_n454_), .A2(new_n471_), .ZN(new_n532_));
  NOR2_X1    g00340(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1    g00341(.A1(new_n533_), .A2(new_n522_), .ZN(new_n534_));
  NOR3_X1    g00342(.A1(new_n531_), .A2(new_n521_), .A3(new_n532_), .ZN(new_n535_));
  NOR2_X1    g00343(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1     g00344(.I(new_n536_), .ZN(new_n537_));
  NAND3_X1   g00345(.A1(new_n509_), .A2(\asqrt[58] ), .A3(new_n512_), .ZN(new_n538_));
  OR4_X2     g00346(.A1(\asqrt[63] ), .A2(new_n527_), .A3(new_n530_), .A4(new_n538_), .Z(new_n539_));
  NAND2_X1   g00347(.A1(\asqrt[57] ), .A2(new_n449_), .ZN(new_n540_));
  AOI21_X1   g00348(.A1(new_n540_), .A2(new_n539_), .B(\a[116] ), .ZN(new_n541_));
  NAND2_X1   g00349(.A1(new_n503_), .A2(new_n193_), .ZN(new_n542_));
  NOR3_X1    g00350(.A1(new_n542_), .A2(new_n530_), .A3(new_n538_), .ZN(new_n543_));
  NOR2_X1    g00351(.A1(new_n531_), .A2(new_n450_), .ZN(new_n544_));
  NOR3_X1    g00352(.A1(new_n544_), .A2(new_n543_), .A3(new_n452_), .ZN(new_n545_));
  NOR2_X1    g00353(.A1(new_n545_), .A2(new_n541_), .ZN(new_n546_));
  INV_X1     g00354(.I(\a[114] ), .ZN(new_n547_));
  NOR2_X1    g00355(.A1(\a[112] ), .A2(\a[113] ), .ZN(new_n548_));
  NOR3_X1    g00356(.A1(new_n531_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1     g00357(.I(new_n548_), .ZN(new_n550_));
  AOI21_X1   g00358(.A1(new_n531_), .A2(\a[114] ), .B(new_n550_), .ZN(new_n551_));
  OAI21_X1   g00359(.A1(new_n549_), .A2(new_n551_), .B(\asqrt[58] ), .ZN(new_n552_));
  INV_X1     g00360(.I(\a[115] ), .ZN(new_n553_));
  AOI21_X1   g00361(.A1(\asqrt[57] ), .A2(new_n547_), .B(new_n553_), .ZN(new_n554_));
  NOR3_X1    g00362(.A1(new_n531_), .A2(\a[114] ), .A3(\a[115] ), .ZN(new_n555_));
  NOR2_X1    g00363(.A1(new_n550_), .A2(\a[114] ), .ZN(new_n556_));
  NOR4_X1    g00364(.A1(new_n411_), .A2(new_n413_), .A3(new_n420_), .A4(new_n556_), .ZN(new_n557_));
  AOI21_X1   g00365(.A1(new_n510_), .A2(new_n557_), .B(new_n547_), .ZN(new_n558_));
  INV_X1     g00366(.I(new_n558_), .ZN(new_n559_));
  NOR2_X1    g00367(.A1(new_n531_), .A2(new_n559_), .ZN(new_n560_));
  NOR3_X1    g00368(.A1(new_n555_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1   g00369(.A1(new_n552_), .A2(new_n561_), .A3(new_n337_), .ZN(new_n562_));
  AOI21_X1   g00370(.A1(new_n552_), .A2(new_n561_), .B(new_n337_), .ZN(new_n563_));
  AOI21_X1   g00371(.A1(new_n546_), .A2(new_n562_), .B(new_n563_), .ZN(new_n564_));
  AOI21_X1   g00372(.A1(new_n564_), .A2(new_n266_), .B(new_n537_), .ZN(new_n565_));
  NAND2_X1   g00373(.A1(new_n562_), .A2(new_n546_), .ZN(new_n566_));
  NAND3_X1   g00374(.A1(\asqrt[57] ), .A2(\a[114] ), .A3(new_n550_), .ZN(new_n567_));
  OAI21_X1   g00375(.A1(\asqrt[57] ), .A2(new_n547_), .B(new_n548_), .ZN(new_n568_));
  AOI21_X1   g00376(.A1(new_n568_), .A2(new_n567_), .B(new_n423_), .ZN(new_n569_));
  OAI21_X1   g00377(.A1(new_n531_), .A2(\a[114] ), .B(\a[115] ), .ZN(new_n570_));
  NAND3_X1   g00378(.A1(\asqrt[57] ), .A2(new_n547_), .A3(new_n553_), .ZN(new_n571_));
  NAND2_X1   g00379(.A1(\asqrt[57] ), .A2(new_n558_), .ZN(new_n572_));
  NAND3_X1   g00380(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1   g00381(.A1(new_n569_), .A2(new_n573_), .B(\asqrt[59] ), .ZN(new_n574_));
  AOI21_X1   g00382(.A1(new_n566_), .A2(new_n574_), .B(new_n266_), .ZN(new_n575_));
  OAI21_X1   g00383(.A1(new_n565_), .A2(new_n575_), .B(\asqrt[61] ), .ZN(new_n576_));
  AOI21_X1   g00384(.A1(new_n478_), .A2(new_n480_), .B(\asqrt[57] ), .ZN(new_n577_));
  XOR2_X1    g00385(.A1(new_n577_), .A2(new_n477_), .Z(new_n578_));
  INV_X1     g00386(.I(new_n578_), .ZN(new_n579_));
  NOR3_X1    g00387(.A1(new_n565_), .A2(\asqrt[61] ), .A3(new_n575_), .ZN(new_n580_));
  OAI21_X1   g00388(.A1(new_n579_), .A2(new_n580_), .B(new_n576_), .ZN(new_n581_));
  OAI21_X1   g00389(.A1(new_n581_), .A2(\asqrt[62] ), .B(new_n517_), .ZN(new_n582_));
  OAI21_X1   g00390(.A1(new_n544_), .A2(new_n543_), .B(new_n452_), .ZN(new_n583_));
  NAND3_X1   g00391(.A1(new_n540_), .A2(new_n539_), .A3(\a[116] ), .ZN(new_n584_));
  NAND2_X1   g00392(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NOR3_X1    g00393(.A1(new_n569_), .A2(new_n573_), .A3(\asqrt[59] ), .ZN(new_n586_));
  OAI21_X1   g00394(.A1(new_n585_), .A2(new_n586_), .B(new_n574_), .ZN(new_n587_));
  OAI21_X1   g00395(.A1(new_n587_), .A2(\asqrt[60] ), .B(new_n536_), .ZN(new_n588_));
  NOR2_X1    g00396(.A1(new_n586_), .A2(new_n585_), .ZN(new_n589_));
  OAI21_X1   g00397(.A1(new_n589_), .A2(new_n563_), .B(\asqrt[60] ), .ZN(new_n590_));
  AOI21_X1   g00398(.A1(new_n588_), .A2(new_n590_), .B(new_n239_), .ZN(new_n591_));
  NAND3_X1   g00399(.A1(new_n588_), .A2(new_n239_), .A3(new_n590_), .ZN(new_n592_));
  AOI21_X1   g00400(.A1(new_n578_), .A2(new_n592_), .B(new_n591_), .ZN(new_n593_));
  NOR2_X1    g00401(.A1(new_n489_), .A2(\asqrt[62] ), .ZN(new_n594_));
  INV_X1     g00402(.I(new_n505_), .ZN(new_n595_));
  NOR2_X1    g00403(.A1(new_n595_), .A2(new_n594_), .ZN(new_n596_));
  XOR2_X1    g00404(.A1(new_n496_), .A2(new_n388_), .Z(new_n597_));
  OAI21_X1   g00405(.A1(\asqrt[57] ), .A2(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1     g00406(.I(new_n598_), .ZN(new_n599_));
  OAI21_X1   g00407(.A1(new_n593_), .A2(new_n201_), .B(new_n599_), .ZN(new_n600_));
  INV_X1     g00408(.I(new_n600_), .ZN(new_n601_));
  NAND2_X1   g00409(.A1(new_n601_), .A2(new_n582_), .ZN(new_n602_));
  INV_X1     g00410(.I(new_n517_), .ZN(new_n603_));
  NAND3_X1   g00411(.A1(new_n566_), .A2(new_n266_), .A3(new_n574_), .ZN(new_n604_));
  AOI21_X1   g00412(.A1(new_n536_), .A2(new_n604_), .B(new_n575_), .ZN(new_n605_));
  AOI21_X1   g00413(.A1(new_n605_), .A2(new_n239_), .B(new_n579_), .ZN(new_n606_));
  OAI21_X1   g00414(.A1(new_n606_), .A2(new_n591_), .B(new_n201_), .ZN(new_n607_));
  NAND2_X1   g00415(.A1(new_n592_), .A2(new_n578_), .ZN(new_n608_));
  NAND3_X1   g00416(.A1(new_n608_), .A2(\asqrt[62] ), .A3(new_n576_), .ZN(new_n609_));
  AOI22_X1   g00417(.A1(new_n607_), .A2(new_n609_), .B1(new_n603_), .B2(new_n581_), .ZN(new_n610_));
  NOR2_X1    g00418(.A1(new_n499_), .A2(new_n486_), .ZN(new_n611_));
  OAI21_X1   g00419(.A1(\asqrt[57] ), .A2(new_n611_), .B(new_n506_), .ZN(new_n612_));
  INV_X1     g00420(.I(new_n612_), .ZN(new_n613_));
  OAI21_X1   g00421(.A1(new_n610_), .A2(new_n599_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1   g00422(.A1(new_n531_), .A2(new_n485_), .ZN(new_n615_));
  XOR2_X1    g00423(.A1(new_n526_), .A2(new_n485_), .Z(new_n616_));
  NAND3_X1   g00424(.A1(new_n615_), .A2(\asqrt[63] ), .A3(new_n616_), .ZN(new_n617_));
  INV_X1     g00425(.I(new_n542_), .ZN(new_n618_));
  NOR3_X1    g00426(.A1(new_n530_), .A2(new_n485_), .A3(new_n513_), .ZN(new_n619_));
  NAND2_X1   g00427(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1   g00428(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1     g00429(.I(new_n621_), .ZN(new_n622_));
  NAND4_X1   g00430(.A1(new_n614_), .A2(new_n193_), .A3(new_n602_), .A4(new_n622_), .ZN(\asqrt[56] ));
  NOR2_X1    g00431(.A1(new_n581_), .A2(\asqrt[62] ), .ZN(new_n624_));
  NOR2_X1    g00432(.A1(new_n593_), .A2(new_n201_), .ZN(new_n625_));
  NOR2_X1    g00433(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1    g00434(.A1(\asqrt[56] ), .A2(new_n626_), .ZN(new_n627_));
  INV_X1     g00435(.I(new_n582_), .ZN(new_n628_));
  NOR2_X1    g00436(.A1(new_n628_), .A2(new_n600_), .ZN(new_n629_));
  AOI21_X1   g00437(.A1(new_n608_), .A2(new_n576_), .B(\asqrt[62] ), .ZN(new_n630_));
  NOR3_X1    g00438(.A1(new_n606_), .A2(new_n201_), .A3(new_n591_), .ZN(new_n631_));
  OAI22_X1   g00439(.A1(new_n631_), .A2(new_n630_), .B1(new_n517_), .B2(new_n593_), .ZN(new_n632_));
  AOI21_X1   g00440(.A1(new_n632_), .A2(new_n598_), .B(new_n612_), .ZN(new_n633_));
  NOR4_X1    g00441(.A1(new_n633_), .A2(\asqrt[63] ), .A3(new_n629_), .A4(new_n621_), .ZN(new_n634_));
  XOR2_X1    g00442(.A1(new_n516_), .A2(new_n491_), .Z(new_n635_));
  NOR2_X1    g00443(.A1(new_n627_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1   g00444(.A1(new_n562_), .A2(new_n574_), .B(\asqrt[56] ), .ZN(new_n637_));
  XOR2_X1    g00445(.A1(new_n637_), .A2(new_n546_), .Z(new_n638_));
  INV_X1     g00446(.I(new_n638_), .ZN(new_n639_));
  NOR2_X1    g00447(.A1(new_n531_), .A2(\a[114] ), .ZN(new_n640_));
  INV_X1     g00448(.I(new_n640_), .ZN(new_n641_));
  NOR2_X1    g00449(.A1(new_n553_), .A2(\a[114] ), .ZN(new_n642_));
  AOI22_X1   g00450(.A1(new_n641_), .A2(new_n553_), .B1(\asqrt[57] ), .B2(new_n642_), .ZN(new_n643_));
  INV_X1     g00451(.I(new_n643_), .ZN(new_n644_));
  NOR2_X1    g00452(.A1(new_n569_), .A2(new_n560_), .ZN(new_n645_));
  NOR2_X1    g00453(.A1(new_n634_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1    g00454(.A1(new_n646_), .A2(new_n644_), .ZN(new_n647_));
  NOR3_X1    g00455(.A1(new_n634_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n648_));
  NOR2_X1    g00456(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1   g00457(.A1(new_n617_), .A2(\asqrt[57] ), .A3(new_n620_), .ZN(new_n650_));
  OR4_X2     g00458(.A1(\asqrt[63] ), .A2(new_n633_), .A3(new_n629_), .A4(new_n650_), .Z(new_n651_));
  NAND2_X1   g00459(.A1(\asqrt[56] ), .A2(new_n548_), .ZN(new_n652_));
  AOI21_X1   g00460(.A1(new_n652_), .A2(new_n651_), .B(\a[114] ), .ZN(new_n653_));
  NAND2_X1   g00461(.A1(new_n614_), .A2(new_n193_), .ZN(new_n654_));
  NOR3_X1    g00462(.A1(new_n654_), .A2(new_n629_), .A3(new_n650_), .ZN(new_n655_));
  NOR2_X1    g00463(.A1(new_n634_), .A2(new_n550_), .ZN(new_n656_));
  NOR3_X1    g00464(.A1(new_n656_), .A2(new_n655_), .A3(new_n547_), .ZN(new_n657_));
  NOR2_X1    g00465(.A1(new_n657_), .A2(new_n653_), .ZN(new_n658_));
  INV_X1     g00466(.I(\a[112] ), .ZN(new_n659_));
  NOR2_X1    g00467(.A1(\a[110] ), .A2(\a[111] ), .ZN(new_n660_));
  NOR3_X1    g00468(.A1(new_n634_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1     g00469(.I(new_n660_), .ZN(new_n662_));
  AOI21_X1   g00470(.A1(new_n634_), .A2(\a[112] ), .B(new_n662_), .ZN(new_n663_));
  OAI21_X1   g00471(.A1(new_n661_), .A2(new_n663_), .B(\asqrt[57] ), .ZN(new_n664_));
  INV_X1     g00472(.I(\a[113] ), .ZN(new_n665_));
  AOI21_X1   g00473(.A1(\asqrt[56] ), .A2(new_n659_), .B(new_n665_), .ZN(new_n666_));
  NOR3_X1    g00474(.A1(new_n634_), .A2(\a[112] ), .A3(\a[113] ), .ZN(new_n667_));
  NAND2_X1   g00475(.A1(new_n660_), .A2(new_n659_), .ZN(new_n668_));
  AND4_X2    g00476(.A1(new_n506_), .A2(new_n509_), .A3(new_n512_), .A4(new_n668_), .Z(new_n669_));
  AOI21_X1   g00477(.A1(new_n618_), .A2(new_n669_), .B(new_n659_), .ZN(new_n670_));
  INV_X1     g00478(.I(new_n670_), .ZN(new_n671_));
  NOR2_X1    g00479(.A1(new_n634_), .A2(new_n671_), .ZN(new_n672_));
  NOR3_X1    g00480(.A1(new_n667_), .A2(new_n666_), .A3(new_n672_), .ZN(new_n673_));
  NAND3_X1   g00481(.A1(new_n664_), .A2(new_n673_), .A3(new_n423_), .ZN(new_n674_));
  NAND2_X1   g00482(.A1(new_n674_), .A2(new_n658_), .ZN(new_n675_));
  NAND3_X1   g00483(.A1(\asqrt[56] ), .A2(\a[112] ), .A3(new_n662_), .ZN(new_n676_));
  OAI21_X1   g00484(.A1(\asqrt[56] ), .A2(new_n659_), .B(new_n660_), .ZN(new_n677_));
  AOI21_X1   g00485(.A1(new_n677_), .A2(new_n676_), .B(new_n531_), .ZN(new_n678_));
  OAI21_X1   g00486(.A1(new_n634_), .A2(\a[112] ), .B(\a[113] ), .ZN(new_n679_));
  NAND3_X1   g00487(.A1(\asqrt[56] ), .A2(new_n659_), .A3(new_n665_), .ZN(new_n680_));
  NAND2_X1   g00488(.A1(\asqrt[56] ), .A2(new_n670_), .ZN(new_n681_));
  NAND3_X1   g00489(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1   g00490(.A1(new_n678_), .A2(new_n682_), .B(\asqrt[58] ), .ZN(new_n683_));
  NAND3_X1   g00491(.A1(new_n675_), .A2(new_n337_), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1   g00492(.A1(new_n675_), .A2(new_n683_), .B(new_n337_), .ZN(new_n685_));
  AOI21_X1   g00493(.A1(new_n649_), .A2(new_n684_), .B(new_n685_), .ZN(new_n686_));
  AOI21_X1   g00494(.A1(new_n686_), .A2(new_n266_), .B(new_n639_), .ZN(new_n687_));
  OR2_X2     g00495(.A1(new_n657_), .A2(new_n653_), .Z(new_n688_));
  NOR3_X1    g00496(.A1(new_n678_), .A2(new_n682_), .A3(\asqrt[58] ), .ZN(new_n689_));
  OAI21_X1   g00497(.A1(new_n688_), .A2(new_n689_), .B(new_n683_), .ZN(new_n690_));
  OAI21_X1   g00498(.A1(new_n690_), .A2(\asqrt[59] ), .B(new_n649_), .ZN(new_n691_));
  NAND2_X1   g00499(.A1(new_n690_), .A2(\asqrt[59] ), .ZN(new_n692_));
  AOI21_X1   g00500(.A1(new_n691_), .A2(new_n692_), .B(new_n266_), .ZN(new_n693_));
  OAI21_X1   g00501(.A1(new_n687_), .A2(new_n693_), .B(\asqrt[61] ), .ZN(new_n694_));
  AOI21_X1   g00502(.A1(new_n604_), .A2(new_n590_), .B(\asqrt[56] ), .ZN(new_n695_));
  XOR2_X1    g00503(.A1(new_n695_), .A2(new_n536_), .Z(new_n696_));
  INV_X1     g00504(.I(new_n696_), .ZN(new_n697_));
  NOR3_X1    g00505(.A1(new_n687_), .A2(\asqrt[61] ), .A3(new_n693_), .ZN(new_n698_));
  OAI21_X1   g00506(.A1(new_n697_), .A2(new_n698_), .B(new_n694_), .ZN(new_n699_));
  NAND3_X1   g00507(.A1(new_n691_), .A2(new_n692_), .A3(new_n266_), .ZN(new_n700_));
  NAND2_X1   g00508(.A1(new_n700_), .A2(new_n638_), .ZN(new_n701_));
  INV_X1     g00509(.I(new_n649_), .ZN(new_n702_));
  AOI21_X1   g00510(.A1(new_n664_), .A2(new_n673_), .B(new_n423_), .ZN(new_n703_));
  AOI21_X1   g00511(.A1(new_n658_), .A2(new_n674_), .B(new_n703_), .ZN(new_n704_));
  AOI21_X1   g00512(.A1(new_n704_), .A2(new_n337_), .B(new_n702_), .ZN(new_n705_));
  OAI21_X1   g00513(.A1(new_n705_), .A2(new_n685_), .B(\asqrt[60] ), .ZN(new_n706_));
  AOI21_X1   g00514(.A1(new_n701_), .A2(new_n706_), .B(new_n239_), .ZN(new_n707_));
  AOI21_X1   g00515(.A1(new_n638_), .A2(new_n700_), .B(new_n693_), .ZN(new_n708_));
  AOI21_X1   g00516(.A1(new_n708_), .A2(new_n239_), .B(new_n697_), .ZN(new_n709_));
  OAI21_X1   g00517(.A1(new_n709_), .A2(new_n707_), .B(new_n201_), .ZN(new_n710_));
  NOR3_X1    g00518(.A1(new_n705_), .A2(\asqrt[60] ), .A3(new_n685_), .ZN(new_n711_));
  OAI21_X1   g00519(.A1(new_n639_), .A2(new_n711_), .B(new_n706_), .ZN(new_n712_));
  OAI21_X1   g00520(.A1(new_n712_), .A2(\asqrt[61] ), .B(new_n696_), .ZN(new_n713_));
  NAND3_X1   g00521(.A1(new_n713_), .A2(\asqrt[62] ), .A3(new_n694_), .ZN(new_n714_));
  AOI21_X1   g00522(.A1(new_n576_), .A2(new_n592_), .B(\asqrt[56] ), .ZN(new_n715_));
  XOR2_X1    g00523(.A1(new_n715_), .A2(new_n578_), .Z(new_n716_));
  INV_X1     g00524(.I(new_n716_), .ZN(new_n717_));
  AOI22_X1   g00525(.A1(new_n714_), .A2(new_n710_), .B1(new_n699_), .B2(new_n717_), .ZN(new_n718_));
  NOR2_X1    g00526(.A1(new_n610_), .A2(new_n599_), .ZN(new_n719_));
  OAI21_X1   g00527(.A1(\asqrt[56] ), .A2(new_n719_), .B(new_n602_), .ZN(new_n720_));
  INV_X1     g00528(.I(new_n720_), .ZN(new_n721_));
  OAI21_X1   g00529(.A1(new_n718_), .A2(new_n636_), .B(new_n721_), .ZN(new_n722_));
  OAI21_X1   g00530(.A1(new_n699_), .A2(\asqrt[62] ), .B(new_n716_), .ZN(new_n723_));
  NAND2_X1   g00531(.A1(new_n699_), .A2(\asqrt[62] ), .ZN(new_n724_));
  NAND3_X1   g00532(.A1(new_n723_), .A2(new_n724_), .A3(new_n636_), .ZN(new_n725_));
  NAND2_X1   g00533(.A1(new_n634_), .A2(new_n598_), .ZN(new_n726_));
  XOR2_X1    g00534(.A1(new_n610_), .A2(new_n599_), .Z(new_n727_));
  NAND3_X1   g00535(.A1(new_n726_), .A2(\asqrt[63] ), .A3(new_n727_), .ZN(new_n728_));
  INV_X1     g00536(.I(new_n654_), .ZN(new_n729_));
  NOR3_X1    g00537(.A1(new_n629_), .A2(new_n598_), .A3(new_n621_), .ZN(new_n730_));
  NAND2_X1   g00538(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1   g00539(.A1(new_n728_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1     g00540(.I(new_n732_), .ZN(new_n733_));
  NAND4_X1   g00541(.A1(new_n722_), .A2(new_n193_), .A3(new_n725_), .A4(new_n733_), .ZN(\asqrt[55] ));
  INV_X1     g00542(.I(new_n636_), .ZN(new_n735_));
  NOR2_X1    g00543(.A1(new_n709_), .A2(new_n707_), .ZN(new_n736_));
  AOI21_X1   g00544(.A1(new_n713_), .A2(new_n694_), .B(\asqrt[62] ), .ZN(new_n737_));
  NOR3_X1    g00545(.A1(new_n709_), .A2(new_n201_), .A3(new_n707_), .ZN(new_n738_));
  OAI22_X1   g00546(.A1(new_n737_), .A2(new_n738_), .B1(new_n736_), .B2(new_n716_), .ZN(new_n739_));
  AOI21_X1   g00547(.A1(new_n739_), .A2(new_n735_), .B(new_n720_), .ZN(new_n740_));
  AOI21_X1   g00548(.A1(new_n736_), .A2(new_n201_), .B(new_n717_), .ZN(new_n741_));
  NOR2_X1    g00549(.A1(new_n736_), .A2(new_n201_), .ZN(new_n742_));
  NOR3_X1    g00550(.A1(new_n741_), .A2(new_n742_), .A3(new_n735_), .ZN(new_n743_));
  NOR4_X1    g00551(.A1(new_n740_), .A2(\asqrt[63] ), .A3(new_n743_), .A4(new_n732_), .ZN(new_n744_));
  NOR2_X1    g00552(.A1(new_n744_), .A2(\a[110] ), .ZN(new_n745_));
  INV_X1     g00553(.I(new_n745_), .ZN(new_n746_));
  NOR2_X1    g00554(.A1(new_n202_), .A2(\a[110] ), .ZN(new_n747_));
  AOI22_X1   g00555(.A1(new_n746_), .A2(new_n202_), .B1(\asqrt[55] ), .B2(new_n747_), .ZN(new_n748_));
  INV_X1     g00556(.I(new_n748_), .ZN(new_n749_));
  NOR2_X1    g00557(.A1(new_n699_), .A2(\asqrt[62] ), .ZN(new_n750_));
  NOR2_X1    g00558(.A1(new_n750_), .A2(new_n742_), .ZN(new_n751_));
  NOR2_X1    g00559(.A1(\asqrt[55] ), .A2(new_n751_), .ZN(new_n752_));
  XOR2_X1    g00560(.A1(new_n715_), .A2(new_n579_), .Z(new_n753_));
  NOR2_X1    g00561(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1     g00562(.I(new_n754_), .ZN(new_n755_));
  AOI21_X1   g00563(.A1(new_n684_), .A2(new_n692_), .B(\asqrt[55] ), .ZN(new_n756_));
  XOR2_X1    g00564(.A1(new_n756_), .A2(new_n649_), .Z(new_n757_));
  AOI21_X1   g00565(.A1(new_n674_), .A2(new_n683_), .B(\asqrt[55] ), .ZN(new_n758_));
  XOR2_X1    g00566(.A1(new_n758_), .A2(new_n658_), .Z(new_n759_));
  NOR2_X1    g00567(.A1(new_n634_), .A2(\a[112] ), .ZN(new_n760_));
  INV_X1     g00568(.I(new_n760_), .ZN(new_n761_));
  NOR2_X1    g00569(.A1(new_n665_), .A2(\a[112] ), .ZN(new_n762_));
  AOI22_X1   g00570(.A1(new_n761_), .A2(new_n665_), .B1(\asqrt[56] ), .B2(new_n762_), .ZN(new_n763_));
  INV_X1     g00571(.I(new_n763_), .ZN(new_n764_));
  NOR2_X1    g00572(.A1(new_n678_), .A2(new_n672_), .ZN(new_n765_));
  INV_X1     g00573(.I(new_n765_), .ZN(new_n766_));
  AOI21_X1   g00574(.A1(\asqrt[55] ), .A2(new_n766_), .B(new_n764_), .ZN(new_n767_));
  NOR2_X1    g00575(.A1(new_n765_), .A2(new_n763_), .ZN(new_n768_));
  AOI21_X1   g00576(.A1(\asqrt[55] ), .A2(new_n768_), .B(new_n767_), .ZN(new_n769_));
  NAND2_X1   g00577(.A1(new_n722_), .A2(new_n193_), .ZN(new_n770_));
  NAND3_X1   g00578(.A1(new_n728_), .A2(\asqrt[56] ), .A3(new_n731_), .ZN(new_n771_));
  NOR3_X1    g00579(.A1(new_n770_), .A2(new_n743_), .A3(new_n771_), .ZN(new_n772_));
  NOR2_X1    g00580(.A1(new_n744_), .A2(new_n662_), .ZN(new_n773_));
  OAI21_X1   g00581(.A1(new_n773_), .A2(new_n772_), .B(new_n659_), .ZN(new_n774_));
  OR4_X2     g00582(.A1(\asqrt[63] ), .A2(new_n740_), .A3(new_n743_), .A4(new_n771_), .Z(new_n775_));
  NAND2_X1   g00583(.A1(\asqrt[55] ), .A2(new_n660_), .ZN(new_n776_));
  NAND3_X1   g00584(.A1(new_n776_), .A2(new_n775_), .A3(\a[112] ), .ZN(new_n777_));
  NAND2_X1   g00585(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1    g00586(.A1(\a[108] ), .A2(\a[109] ), .ZN(new_n779_));
  INV_X1     g00587(.I(new_n779_), .ZN(new_n780_));
  NAND3_X1   g00588(.A1(\asqrt[55] ), .A2(\a[110] ), .A3(new_n780_), .ZN(new_n781_));
  INV_X1     g00589(.I(\a[110] ), .ZN(new_n782_));
  OAI21_X1   g00590(.A1(\asqrt[55] ), .A2(new_n782_), .B(new_n779_), .ZN(new_n783_));
  AOI21_X1   g00591(.A1(new_n783_), .A2(new_n781_), .B(new_n634_), .ZN(new_n784_));
  OAI21_X1   g00592(.A1(new_n744_), .A2(\a[110] ), .B(\a[111] ), .ZN(new_n785_));
  NAND3_X1   g00593(.A1(\asqrt[55] ), .A2(new_n782_), .A3(new_n202_), .ZN(new_n786_));
  NAND2_X1   g00594(.A1(new_n779_), .A2(new_n782_), .ZN(new_n787_));
  AND4_X2    g00595(.A1(new_n602_), .A2(new_n617_), .A3(new_n620_), .A4(new_n787_), .Z(new_n788_));
  AOI21_X1   g00596(.A1(new_n729_), .A2(new_n788_), .B(new_n782_), .ZN(new_n789_));
  NAND2_X1   g00597(.A1(\asqrt[55] ), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1   g00598(.A1(new_n785_), .A2(new_n786_), .A3(new_n790_), .ZN(new_n791_));
  NOR3_X1    g00599(.A1(new_n784_), .A2(new_n791_), .A3(\asqrt[57] ), .ZN(new_n792_));
  OAI21_X1   g00600(.A1(new_n784_), .A2(new_n791_), .B(\asqrt[57] ), .ZN(new_n793_));
  OAI21_X1   g00601(.A1(new_n778_), .A2(new_n792_), .B(new_n793_), .ZN(new_n794_));
  OAI21_X1   g00602(.A1(new_n794_), .A2(\asqrt[58] ), .B(new_n769_), .ZN(new_n795_));
  NOR2_X1    g00603(.A1(new_n792_), .A2(new_n778_), .ZN(new_n796_));
  INV_X1     g00604(.I(new_n793_), .ZN(new_n797_));
  OAI21_X1   g00605(.A1(new_n796_), .A2(new_n797_), .B(\asqrt[58] ), .ZN(new_n798_));
  NAND3_X1   g00606(.A1(new_n795_), .A2(new_n337_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1   g00607(.A1(new_n799_), .A2(new_n759_), .ZN(new_n800_));
  INV_X1     g00608(.I(new_n769_), .ZN(new_n801_));
  NOR2_X1    g00609(.A1(new_n796_), .A2(new_n797_), .ZN(new_n802_));
  AOI21_X1   g00610(.A1(new_n802_), .A2(new_n423_), .B(new_n801_), .ZN(new_n803_));
  AOI21_X1   g00611(.A1(new_n776_), .A2(new_n775_), .B(\a[112] ), .ZN(new_n804_));
  NOR3_X1    g00612(.A1(new_n773_), .A2(new_n772_), .A3(new_n659_), .ZN(new_n805_));
  NOR2_X1    g00613(.A1(new_n805_), .A2(new_n804_), .ZN(new_n806_));
  NOR3_X1    g00614(.A1(new_n744_), .A2(new_n782_), .A3(new_n779_), .ZN(new_n807_));
  AOI21_X1   g00615(.A1(new_n744_), .A2(\a[110] ), .B(new_n780_), .ZN(new_n808_));
  OAI21_X1   g00616(.A1(new_n807_), .A2(new_n808_), .B(\asqrt[56] ), .ZN(new_n809_));
  AOI21_X1   g00617(.A1(\asqrt[55] ), .A2(new_n782_), .B(new_n202_), .ZN(new_n810_));
  NOR3_X1    g00618(.A1(new_n744_), .A2(\a[110] ), .A3(\a[111] ), .ZN(new_n811_));
  INV_X1     g00619(.I(new_n789_), .ZN(new_n812_));
  NOR2_X1    g00620(.A1(new_n744_), .A2(new_n812_), .ZN(new_n813_));
  NOR3_X1    g00621(.A1(new_n811_), .A2(new_n810_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1   g00622(.A1(new_n809_), .A2(new_n814_), .A3(new_n531_), .ZN(new_n815_));
  NAND2_X1   g00623(.A1(new_n815_), .A2(new_n806_), .ZN(new_n816_));
  AOI21_X1   g00624(.A1(new_n816_), .A2(new_n793_), .B(new_n423_), .ZN(new_n817_));
  OAI21_X1   g00625(.A1(new_n803_), .A2(new_n817_), .B(\asqrt[59] ), .ZN(new_n818_));
  NAND3_X1   g00626(.A1(new_n800_), .A2(new_n266_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1   g00627(.A1(new_n819_), .A2(new_n757_), .ZN(new_n820_));
  INV_X1     g00628(.I(new_n759_), .ZN(new_n821_));
  NAND3_X1   g00629(.A1(new_n816_), .A2(new_n423_), .A3(new_n793_), .ZN(new_n822_));
  AOI21_X1   g00630(.A1(new_n769_), .A2(new_n822_), .B(new_n817_), .ZN(new_n823_));
  AOI21_X1   g00631(.A1(new_n823_), .A2(new_n337_), .B(new_n821_), .ZN(new_n824_));
  NOR2_X1    g00632(.A1(new_n823_), .A2(new_n337_), .ZN(new_n825_));
  OAI21_X1   g00633(.A1(new_n824_), .A2(new_n825_), .B(\asqrt[60] ), .ZN(new_n826_));
  AOI21_X1   g00634(.A1(new_n820_), .A2(new_n826_), .B(new_n239_), .ZN(new_n827_));
  AOI21_X1   g00635(.A1(new_n800_), .A2(new_n818_), .B(new_n266_), .ZN(new_n828_));
  AOI21_X1   g00636(.A1(new_n757_), .A2(new_n819_), .B(new_n828_), .ZN(new_n829_));
  AOI21_X1   g00637(.A1(new_n700_), .A2(new_n706_), .B(\asqrt[55] ), .ZN(new_n830_));
  XOR2_X1    g00638(.A1(new_n830_), .A2(new_n638_), .Z(new_n831_));
  INV_X1     g00639(.I(new_n831_), .ZN(new_n832_));
  AOI21_X1   g00640(.A1(new_n829_), .A2(new_n239_), .B(new_n832_), .ZN(new_n833_));
  NOR2_X1    g00641(.A1(new_n833_), .A2(new_n827_), .ZN(new_n834_));
  INV_X1     g00642(.I(new_n757_), .ZN(new_n835_));
  NOR3_X1    g00643(.A1(new_n824_), .A2(new_n825_), .A3(\asqrt[60] ), .ZN(new_n836_));
  OAI21_X1   g00644(.A1(new_n835_), .A2(new_n836_), .B(new_n826_), .ZN(new_n837_));
  NAND2_X1   g00645(.A1(new_n837_), .A2(\asqrt[61] ), .ZN(new_n838_));
  OAI21_X1   g00646(.A1(new_n837_), .A2(\asqrt[61] ), .B(new_n831_), .ZN(new_n839_));
  AOI21_X1   g00647(.A1(new_n839_), .A2(new_n838_), .B(\asqrt[62] ), .ZN(new_n840_));
  NOR3_X1    g00648(.A1(new_n833_), .A2(new_n201_), .A3(new_n827_), .ZN(new_n841_));
  NOR2_X1    g00649(.A1(new_n698_), .A2(new_n707_), .ZN(new_n842_));
  NOR2_X1    g00650(.A1(\asqrt[55] ), .A2(new_n842_), .ZN(new_n843_));
  XOR2_X1    g00651(.A1(new_n843_), .A2(new_n696_), .Z(new_n844_));
  OAI22_X1   g00652(.A1(new_n840_), .A2(new_n841_), .B1(new_n834_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1    g00653(.A1(new_n718_), .A2(new_n636_), .ZN(new_n846_));
  OAI21_X1   g00654(.A1(\asqrt[55] ), .A2(new_n846_), .B(new_n725_), .ZN(new_n847_));
  AOI21_X1   g00655(.A1(new_n845_), .A2(new_n755_), .B(new_n847_), .ZN(new_n848_));
  INV_X1     g00656(.I(new_n844_), .ZN(new_n849_));
  AOI21_X1   g00657(.A1(new_n834_), .A2(new_n201_), .B(new_n849_), .ZN(new_n850_));
  NOR2_X1    g00658(.A1(new_n834_), .A2(new_n201_), .ZN(new_n851_));
  NOR3_X1    g00659(.A1(new_n850_), .A2(new_n851_), .A3(new_n755_), .ZN(new_n852_));
  NAND2_X1   g00660(.A1(new_n744_), .A2(new_n735_), .ZN(new_n853_));
  XOR2_X1    g00661(.A1(new_n739_), .A2(new_n735_), .Z(new_n854_));
  NAND3_X1   g00662(.A1(new_n853_), .A2(\asqrt[63] ), .A3(new_n854_), .ZN(new_n855_));
  INV_X1     g00663(.I(new_n770_), .ZN(new_n856_));
  NOR3_X1    g00664(.A1(new_n743_), .A2(new_n735_), .A3(new_n732_), .ZN(new_n857_));
  NAND2_X1   g00665(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1   g00666(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  NOR4_X1    g00667(.A1(new_n848_), .A2(\asqrt[63] ), .A3(new_n852_), .A4(new_n859_), .ZN(new_n860_));
  NOR2_X1    g00668(.A1(new_n784_), .A2(new_n813_), .ZN(new_n861_));
  NOR2_X1    g00669(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1    g00670(.A1(new_n862_), .A2(new_n749_), .ZN(new_n863_));
  NOR3_X1    g00671(.A1(new_n860_), .A2(new_n748_), .A3(new_n861_), .ZN(new_n864_));
  NOR2_X1    g00672(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1   g00673(.A1(new_n839_), .A2(new_n838_), .ZN(new_n866_));
  OAI21_X1   g00674(.A1(new_n833_), .A2(new_n827_), .B(new_n201_), .ZN(new_n867_));
  NAND3_X1   g00675(.A1(new_n839_), .A2(new_n838_), .A3(\asqrt[62] ), .ZN(new_n868_));
  AOI22_X1   g00676(.A1(new_n868_), .A2(new_n867_), .B1(new_n866_), .B2(new_n849_), .ZN(new_n869_));
  INV_X1     g00677(.I(new_n847_), .ZN(new_n870_));
  OAI21_X1   g00678(.A1(new_n869_), .A2(new_n754_), .B(new_n870_), .ZN(new_n871_));
  NAND2_X1   g00679(.A1(new_n871_), .A2(new_n193_), .ZN(new_n872_));
  INV_X1     g00680(.I(new_n858_), .ZN(new_n873_));
  NOR2_X1    g00681(.A1(new_n873_), .A2(new_n744_), .ZN(new_n874_));
  NAND2_X1   g00682(.A1(new_n874_), .A2(new_n855_), .ZN(new_n875_));
  NOR3_X1    g00683(.A1(new_n872_), .A2(new_n852_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1     g00684(.I(new_n876_), .ZN(new_n877_));
  OAI21_X1   g00685(.A1(new_n866_), .A2(\asqrt[62] ), .B(new_n844_), .ZN(new_n878_));
  NAND2_X1   g00686(.A1(new_n866_), .A2(\asqrt[62] ), .ZN(new_n879_));
  NAND3_X1   g00687(.A1(new_n878_), .A2(new_n879_), .A3(new_n754_), .ZN(new_n880_));
  INV_X1     g00688(.I(new_n859_), .ZN(new_n881_));
  NAND4_X1   g00689(.A1(new_n871_), .A2(new_n193_), .A3(new_n880_), .A4(new_n881_), .ZN(\asqrt[54] ));
  NAND2_X1   g00690(.A1(\asqrt[54] ), .A2(new_n779_), .ZN(new_n883_));
  AOI21_X1   g00691(.A1(new_n877_), .A2(new_n883_), .B(\a[110] ), .ZN(new_n884_));
  NOR2_X1    g00692(.A1(new_n860_), .A2(new_n780_), .ZN(new_n885_));
  NOR3_X1    g00693(.A1(new_n885_), .A2(new_n876_), .A3(new_n782_), .ZN(new_n886_));
  NOR2_X1    g00694(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1     g00695(.I(\a[108] ), .ZN(new_n888_));
  NOR2_X1    g00696(.A1(\a[106] ), .A2(\a[107] ), .ZN(new_n889_));
  NOR3_X1    g00697(.A1(new_n860_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1     g00698(.I(new_n889_), .ZN(new_n891_));
  AOI21_X1   g00699(.A1(new_n860_), .A2(\a[108] ), .B(new_n891_), .ZN(new_n892_));
  OAI21_X1   g00700(.A1(new_n890_), .A2(new_n892_), .B(\asqrt[55] ), .ZN(new_n893_));
  INV_X1     g00701(.I(\a[109] ), .ZN(new_n894_));
  AOI21_X1   g00702(.A1(\asqrt[54] ), .A2(new_n888_), .B(new_n894_), .ZN(new_n895_));
  NOR3_X1    g00703(.A1(new_n860_), .A2(\a[108] ), .A3(\a[109] ), .ZN(new_n896_));
  NOR3_X1    g00704(.A1(new_n848_), .A2(\asqrt[63] ), .A3(new_n852_), .ZN(new_n897_));
  NAND2_X1   g00705(.A1(new_n889_), .A2(new_n888_), .ZN(new_n898_));
  AND4_X2    g00706(.A1(new_n725_), .A2(new_n728_), .A3(new_n731_), .A4(new_n898_), .Z(new_n899_));
  AOI21_X1   g00707(.A1(new_n856_), .A2(new_n899_), .B(new_n888_), .ZN(new_n900_));
  INV_X1     g00708(.I(new_n900_), .ZN(new_n901_));
  AOI21_X1   g00709(.A1(new_n897_), .A2(new_n881_), .B(new_n901_), .ZN(new_n902_));
  NOR3_X1    g00710(.A1(new_n896_), .A2(new_n895_), .A3(new_n902_), .ZN(new_n903_));
  NAND3_X1   g00711(.A1(new_n893_), .A2(new_n903_), .A3(new_n634_), .ZN(new_n904_));
  AOI21_X1   g00712(.A1(new_n893_), .A2(new_n903_), .B(new_n634_), .ZN(new_n905_));
  AOI21_X1   g00713(.A1(new_n887_), .A2(new_n904_), .B(new_n905_), .ZN(new_n906_));
  NAND2_X1   g00714(.A1(new_n906_), .A2(new_n531_), .ZN(new_n907_));
  OAI21_X1   g00715(.A1(new_n885_), .A2(new_n876_), .B(new_n782_), .ZN(new_n908_));
  INV_X1     g00716(.I(new_n886_), .ZN(new_n909_));
  NAND2_X1   g00717(.A1(new_n909_), .A2(new_n908_), .ZN(new_n910_));
  NAND3_X1   g00718(.A1(\asqrt[54] ), .A2(\a[108] ), .A3(new_n891_), .ZN(new_n911_));
  OAI21_X1   g00719(.A1(\asqrt[54] ), .A2(new_n888_), .B(new_n889_), .ZN(new_n912_));
  AOI21_X1   g00720(.A1(new_n912_), .A2(new_n911_), .B(new_n744_), .ZN(new_n913_));
  OAI21_X1   g00721(.A1(new_n860_), .A2(\a[108] ), .B(\a[109] ), .ZN(new_n914_));
  NAND3_X1   g00722(.A1(\asqrt[54] ), .A2(new_n888_), .A3(new_n894_), .ZN(new_n915_));
  NAND2_X1   g00723(.A1(\asqrt[54] ), .A2(new_n900_), .ZN(new_n916_));
  NAND3_X1   g00724(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  NOR3_X1    g00725(.A1(new_n913_), .A2(new_n917_), .A3(\asqrt[56] ), .ZN(new_n918_));
  OAI21_X1   g00726(.A1(new_n913_), .A2(new_n917_), .B(\asqrt[56] ), .ZN(new_n919_));
  OAI21_X1   g00727(.A1(new_n910_), .A2(new_n918_), .B(new_n919_), .ZN(new_n920_));
  NAND2_X1   g00728(.A1(new_n920_), .A2(\asqrt[57] ), .ZN(new_n921_));
  NOR2_X1    g00729(.A1(new_n866_), .A2(\asqrt[62] ), .ZN(new_n922_));
  NOR2_X1    g00730(.A1(new_n922_), .A2(new_n851_), .ZN(new_n923_));
  XOR2_X1    g00731(.A1(new_n843_), .A2(new_n696_), .Z(new_n924_));
  OAI21_X1   g00732(.A1(\asqrt[54] ), .A2(new_n923_), .B(new_n924_), .ZN(new_n925_));
  INV_X1     g00733(.I(new_n925_), .ZN(new_n926_));
  AOI21_X1   g00734(.A1(new_n799_), .A2(new_n818_), .B(\asqrt[54] ), .ZN(new_n927_));
  XOR2_X1    g00735(.A1(new_n927_), .A2(new_n759_), .Z(new_n928_));
  INV_X1     g00736(.I(new_n928_), .ZN(new_n929_));
  AOI21_X1   g00737(.A1(new_n822_), .A2(new_n798_), .B(\asqrt[54] ), .ZN(new_n930_));
  XOR2_X1    g00738(.A1(new_n930_), .A2(new_n769_), .Z(new_n931_));
  INV_X1     g00739(.I(new_n931_), .ZN(new_n932_));
  AOI21_X1   g00740(.A1(new_n815_), .A2(new_n793_), .B(\asqrt[54] ), .ZN(new_n933_));
  XOR2_X1    g00741(.A1(new_n933_), .A2(new_n806_), .Z(new_n934_));
  OAI21_X1   g00742(.A1(new_n920_), .A2(\asqrt[57] ), .B(new_n865_), .ZN(new_n935_));
  NAND3_X1   g00743(.A1(new_n935_), .A2(new_n921_), .A3(new_n423_), .ZN(new_n936_));
  AOI21_X1   g00744(.A1(new_n935_), .A2(new_n921_), .B(new_n423_), .ZN(new_n937_));
  AOI21_X1   g00745(.A1(new_n934_), .A2(new_n936_), .B(new_n937_), .ZN(new_n938_));
  AOI21_X1   g00746(.A1(new_n938_), .A2(new_n337_), .B(new_n932_), .ZN(new_n939_));
  NAND2_X1   g00747(.A1(new_n936_), .A2(new_n934_), .ZN(new_n940_));
  INV_X1     g00748(.I(new_n865_), .ZN(new_n941_));
  AOI21_X1   g00749(.A1(new_n906_), .A2(new_n531_), .B(new_n941_), .ZN(new_n942_));
  NAND2_X1   g00750(.A1(new_n904_), .A2(new_n887_), .ZN(new_n943_));
  AOI21_X1   g00751(.A1(new_n943_), .A2(new_n919_), .B(new_n531_), .ZN(new_n944_));
  OAI21_X1   g00752(.A1(new_n942_), .A2(new_n944_), .B(\asqrt[58] ), .ZN(new_n945_));
  AOI21_X1   g00753(.A1(new_n940_), .A2(new_n945_), .B(new_n337_), .ZN(new_n946_));
  NOR3_X1    g00754(.A1(new_n939_), .A2(\asqrt[60] ), .A3(new_n946_), .ZN(new_n947_));
  NOR2_X1    g00755(.A1(new_n947_), .A2(new_n929_), .ZN(new_n948_));
  INV_X1     g00756(.I(new_n934_), .ZN(new_n949_));
  NOR3_X1    g00757(.A1(new_n942_), .A2(\asqrt[58] ), .A3(new_n944_), .ZN(new_n950_));
  OAI21_X1   g00758(.A1(new_n949_), .A2(new_n950_), .B(new_n945_), .ZN(new_n951_));
  OAI21_X1   g00759(.A1(new_n951_), .A2(\asqrt[59] ), .B(new_n931_), .ZN(new_n952_));
  NOR2_X1    g00760(.A1(new_n950_), .A2(new_n949_), .ZN(new_n953_));
  OAI21_X1   g00761(.A1(new_n953_), .A2(new_n937_), .B(\asqrt[59] ), .ZN(new_n954_));
  AOI21_X1   g00762(.A1(new_n952_), .A2(new_n954_), .B(new_n266_), .ZN(new_n955_));
  OAI21_X1   g00763(.A1(new_n948_), .A2(new_n955_), .B(\asqrt[61] ), .ZN(new_n956_));
  OAI21_X1   g00764(.A1(new_n939_), .A2(new_n946_), .B(\asqrt[60] ), .ZN(new_n957_));
  OAI21_X1   g00765(.A1(new_n929_), .A2(new_n947_), .B(new_n957_), .ZN(new_n958_));
  AOI21_X1   g00766(.A1(new_n819_), .A2(new_n826_), .B(\asqrt[54] ), .ZN(new_n959_));
  XOR2_X1    g00767(.A1(new_n959_), .A2(new_n757_), .Z(new_n960_));
  OAI21_X1   g00768(.A1(new_n958_), .A2(\asqrt[61] ), .B(new_n960_), .ZN(new_n961_));
  NAND2_X1   g00769(.A1(new_n961_), .A2(new_n956_), .ZN(new_n962_));
  NAND3_X1   g00770(.A1(new_n952_), .A2(new_n266_), .A3(new_n954_), .ZN(new_n963_));
  NAND2_X1   g00771(.A1(new_n963_), .A2(new_n928_), .ZN(new_n964_));
  AOI21_X1   g00772(.A1(new_n964_), .A2(new_n957_), .B(new_n239_), .ZN(new_n965_));
  AOI21_X1   g00773(.A1(new_n928_), .A2(new_n963_), .B(new_n955_), .ZN(new_n966_));
  INV_X1     g00774(.I(new_n960_), .ZN(new_n967_));
  AOI21_X1   g00775(.A1(new_n966_), .A2(new_n239_), .B(new_n967_), .ZN(new_n968_));
  OAI21_X1   g00776(.A1(new_n968_), .A2(new_n965_), .B(new_n201_), .ZN(new_n969_));
  NAND3_X1   g00777(.A1(new_n961_), .A2(\asqrt[62] ), .A3(new_n956_), .ZN(new_n970_));
  NAND2_X1   g00778(.A1(new_n829_), .A2(new_n239_), .ZN(new_n971_));
  AOI21_X1   g00779(.A1(new_n838_), .A2(new_n971_), .B(\asqrt[54] ), .ZN(new_n972_));
  XOR2_X1    g00780(.A1(new_n972_), .A2(new_n831_), .Z(new_n973_));
  INV_X1     g00781(.I(new_n973_), .ZN(new_n974_));
  AOI22_X1   g00782(.A1(new_n969_), .A2(new_n970_), .B1(new_n962_), .B2(new_n974_), .ZN(new_n975_));
  NOR2_X1    g00783(.A1(new_n869_), .A2(new_n754_), .ZN(new_n976_));
  OAI21_X1   g00784(.A1(\asqrt[54] ), .A2(new_n976_), .B(new_n880_), .ZN(new_n977_));
  INV_X1     g00785(.I(new_n977_), .ZN(new_n978_));
  OAI21_X1   g00786(.A1(new_n975_), .A2(new_n926_), .B(new_n978_), .ZN(new_n979_));
  OAI21_X1   g00787(.A1(new_n962_), .A2(\asqrt[62] ), .B(new_n973_), .ZN(new_n980_));
  NAND2_X1   g00788(.A1(new_n962_), .A2(\asqrt[62] ), .ZN(new_n981_));
  NAND3_X1   g00789(.A1(new_n980_), .A2(new_n981_), .A3(new_n926_), .ZN(new_n982_));
  NAND2_X1   g00790(.A1(new_n860_), .A2(new_n755_), .ZN(new_n983_));
  XOR2_X1    g00791(.A1(new_n845_), .A2(new_n755_), .Z(new_n984_));
  NAND3_X1   g00792(.A1(new_n983_), .A2(\asqrt[63] ), .A3(new_n984_), .ZN(new_n985_));
  INV_X1     g00793(.I(new_n872_), .ZN(new_n986_));
  NOR3_X1    g00794(.A1(new_n852_), .A2(new_n755_), .A3(new_n859_), .ZN(new_n987_));
  NAND2_X1   g00795(.A1(new_n986_), .A2(new_n987_), .ZN(new_n988_));
  NAND2_X1   g00796(.A1(new_n985_), .A2(new_n988_), .ZN(new_n989_));
  INV_X1     g00797(.I(new_n989_), .ZN(new_n990_));
  NAND4_X1   g00798(.A1(new_n979_), .A2(new_n193_), .A3(new_n982_), .A4(new_n990_), .ZN(\asqrt[53] ));
  AOI21_X1   g00799(.A1(new_n907_), .A2(new_n921_), .B(\asqrt[53] ), .ZN(new_n992_));
  XOR2_X1    g00800(.A1(new_n992_), .A2(new_n865_), .Z(new_n993_));
  NOR2_X1    g00801(.A1(new_n962_), .A2(\asqrt[62] ), .ZN(new_n994_));
  INV_X1     g00802(.I(new_n981_), .ZN(new_n995_));
  NOR2_X1    g00803(.A1(new_n995_), .A2(new_n994_), .ZN(new_n996_));
  NAND3_X1   g00804(.A1(new_n964_), .A2(new_n239_), .A3(new_n957_), .ZN(new_n997_));
  AOI21_X1   g00805(.A1(new_n960_), .A2(new_n997_), .B(new_n965_), .ZN(new_n998_));
  AOI21_X1   g00806(.A1(new_n961_), .A2(new_n956_), .B(\asqrt[62] ), .ZN(new_n999_));
  NOR3_X1    g00807(.A1(new_n968_), .A2(new_n201_), .A3(new_n965_), .ZN(new_n1000_));
  OAI22_X1   g00808(.A1(new_n1000_), .A2(new_n999_), .B1(new_n998_), .B2(new_n973_), .ZN(new_n1001_));
  AOI21_X1   g00809(.A1(new_n1001_), .A2(new_n925_), .B(new_n977_), .ZN(new_n1002_));
  AOI21_X1   g00810(.A1(new_n998_), .A2(new_n201_), .B(new_n974_), .ZN(new_n1003_));
  OAI21_X1   g00811(.A1(new_n998_), .A2(new_n201_), .B(new_n926_), .ZN(new_n1004_));
  NOR2_X1    g00812(.A1(new_n1003_), .A2(new_n1004_), .ZN(new_n1005_));
  NOR4_X1    g00813(.A1(new_n1002_), .A2(\asqrt[63] ), .A3(new_n1005_), .A4(new_n989_), .ZN(new_n1006_));
  XOR2_X1    g00814(.A1(new_n972_), .A2(new_n831_), .Z(new_n1007_));
  OAI21_X1   g00815(.A1(\asqrt[53] ), .A2(new_n996_), .B(new_n1007_), .ZN(new_n1008_));
  INV_X1     g00816(.I(new_n1008_), .ZN(new_n1009_));
  NAND2_X1   g00817(.A1(new_n938_), .A2(new_n337_), .ZN(new_n1010_));
  AOI21_X1   g00818(.A1(new_n1010_), .A2(new_n954_), .B(\asqrt[53] ), .ZN(new_n1011_));
  XOR2_X1    g00819(.A1(new_n1011_), .A2(new_n931_), .Z(new_n1012_));
  INV_X1     g00820(.I(new_n1012_), .ZN(new_n1013_));
  AOI21_X1   g00821(.A1(new_n936_), .A2(new_n945_), .B(\asqrt[53] ), .ZN(new_n1014_));
  XOR2_X1    g00822(.A1(new_n1014_), .A2(new_n934_), .Z(new_n1015_));
  INV_X1     g00823(.I(new_n1015_), .ZN(new_n1016_));
  INV_X1     g00824(.I(new_n993_), .ZN(new_n1017_));
  AOI21_X1   g00825(.A1(new_n904_), .A2(new_n919_), .B(\asqrt[53] ), .ZN(new_n1018_));
  XOR2_X1    g00826(.A1(new_n1018_), .A2(new_n887_), .Z(new_n1019_));
  NOR2_X1    g00827(.A1(new_n860_), .A2(\a[108] ), .ZN(new_n1020_));
  INV_X1     g00828(.I(new_n1020_), .ZN(new_n1021_));
  NOR2_X1    g00829(.A1(new_n894_), .A2(\a[108] ), .ZN(new_n1022_));
  AOI22_X1   g00830(.A1(new_n1021_), .A2(new_n894_), .B1(\asqrt[54] ), .B2(new_n1022_), .ZN(new_n1023_));
  INV_X1     g00831(.I(new_n1023_), .ZN(new_n1024_));
  NOR2_X1    g00832(.A1(new_n913_), .A2(new_n902_), .ZN(new_n1025_));
  INV_X1     g00833(.I(new_n1025_), .ZN(new_n1026_));
  AOI21_X1   g00834(.A1(\asqrt[53] ), .A2(new_n1026_), .B(new_n1024_), .ZN(new_n1027_));
  NOR2_X1    g00835(.A1(new_n1025_), .A2(new_n1023_), .ZN(new_n1028_));
  AOI21_X1   g00836(.A1(\asqrt[53] ), .A2(new_n1028_), .B(new_n1027_), .ZN(new_n1029_));
  NAND3_X1   g00837(.A1(new_n985_), .A2(\asqrt[54] ), .A3(new_n988_), .ZN(new_n1030_));
  OR4_X2     g00838(.A1(\asqrt[63] ), .A2(new_n1002_), .A3(new_n1005_), .A4(new_n1030_), .Z(new_n1031_));
  NAND2_X1   g00839(.A1(\asqrt[53] ), .A2(new_n889_), .ZN(new_n1032_));
  AOI21_X1   g00840(.A1(new_n1032_), .A2(new_n1031_), .B(\a[108] ), .ZN(new_n1033_));
  NAND2_X1   g00841(.A1(new_n979_), .A2(new_n193_), .ZN(new_n1034_));
  NOR3_X1    g00842(.A1(new_n1034_), .A2(new_n1005_), .A3(new_n1030_), .ZN(new_n1035_));
  NOR2_X1    g00843(.A1(new_n1006_), .A2(new_n891_), .ZN(new_n1036_));
  NOR3_X1    g00844(.A1(new_n1036_), .A2(new_n1035_), .A3(new_n888_), .ZN(new_n1037_));
  OR2_X2     g00845(.A1(new_n1037_), .A2(new_n1033_), .Z(new_n1038_));
  NOR2_X1    g00846(.A1(\a[104] ), .A2(\a[105] ), .ZN(new_n1039_));
  INV_X1     g00847(.I(new_n1039_), .ZN(new_n1040_));
  NAND3_X1   g00848(.A1(\asqrt[53] ), .A2(\a[106] ), .A3(new_n1040_), .ZN(new_n1041_));
  INV_X1     g00849(.I(\a[106] ), .ZN(new_n1042_));
  OAI21_X1   g00850(.A1(\asqrt[53] ), .A2(new_n1042_), .B(new_n1039_), .ZN(new_n1043_));
  AOI21_X1   g00851(.A1(new_n1043_), .A2(new_n1041_), .B(new_n860_), .ZN(new_n1044_));
  OAI21_X1   g00852(.A1(new_n1006_), .A2(\a[106] ), .B(\a[107] ), .ZN(new_n1045_));
  INV_X1     g00853(.I(\a[107] ), .ZN(new_n1046_));
  NAND3_X1   g00854(.A1(\asqrt[53] ), .A2(new_n1042_), .A3(new_n1046_), .ZN(new_n1047_));
  AOI21_X1   g00855(.A1(new_n1042_), .A2(new_n1039_), .B(new_n873_), .ZN(new_n1048_));
  AND3_X2    g00856(.A1(new_n880_), .A2(new_n855_), .A3(new_n1048_), .Z(new_n1049_));
  AOI21_X1   g00857(.A1(new_n986_), .A2(new_n1049_), .B(new_n1042_), .ZN(new_n1050_));
  NAND2_X1   g00858(.A1(\asqrt[53] ), .A2(new_n1050_), .ZN(new_n1051_));
  NAND3_X1   g00859(.A1(new_n1045_), .A2(new_n1047_), .A3(new_n1051_), .ZN(new_n1052_));
  NOR3_X1    g00860(.A1(new_n1044_), .A2(new_n1052_), .A3(\asqrt[55] ), .ZN(new_n1053_));
  OAI21_X1   g00861(.A1(new_n1044_), .A2(new_n1052_), .B(\asqrt[55] ), .ZN(new_n1054_));
  OAI21_X1   g00862(.A1(new_n1038_), .A2(new_n1053_), .B(new_n1054_), .ZN(new_n1055_));
  OAI21_X1   g00863(.A1(new_n1055_), .A2(\asqrt[56] ), .B(new_n1029_), .ZN(new_n1056_));
  NAND2_X1   g00864(.A1(new_n1055_), .A2(\asqrt[56] ), .ZN(new_n1057_));
  NAND3_X1   g00865(.A1(new_n1056_), .A2(new_n1057_), .A3(new_n531_), .ZN(new_n1058_));
  AOI21_X1   g00866(.A1(new_n1056_), .A2(new_n1057_), .B(new_n531_), .ZN(new_n1059_));
  AOI21_X1   g00867(.A1(new_n1019_), .A2(new_n1058_), .B(new_n1059_), .ZN(new_n1060_));
  AOI21_X1   g00868(.A1(new_n1060_), .A2(new_n423_), .B(new_n1017_), .ZN(new_n1061_));
  NAND2_X1   g00869(.A1(new_n1058_), .A2(new_n1019_), .ZN(new_n1062_));
  INV_X1     g00870(.I(new_n1059_), .ZN(new_n1063_));
  AOI21_X1   g00871(.A1(new_n1062_), .A2(new_n1063_), .B(new_n423_), .ZN(new_n1064_));
  NOR3_X1    g00872(.A1(new_n1061_), .A2(\asqrt[59] ), .A3(new_n1064_), .ZN(new_n1065_));
  NOR2_X1    g00873(.A1(new_n1065_), .A2(new_n1016_), .ZN(new_n1066_));
  OAI21_X1   g00874(.A1(new_n1061_), .A2(new_n1064_), .B(\asqrt[59] ), .ZN(new_n1067_));
  INV_X1     g00875(.I(new_n1067_), .ZN(new_n1068_));
  NOR2_X1    g00876(.A1(new_n1066_), .A2(new_n1068_), .ZN(new_n1069_));
  AOI21_X1   g00877(.A1(new_n1069_), .A2(new_n266_), .B(new_n1013_), .ZN(new_n1070_));
  INV_X1     g00878(.I(new_n1019_), .ZN(new_n1071_));
  NOR2_X1    g00879(.A1(new_n1037_), .A2(new_n1033_), .ZN(new_n1072_));
  NOR3_X1    g00880(.A1(new_n1006_), .A2(new_n1042_), .A3(new_n1039_), .ZN(new_n1073_));
  AOI21_X1   g00881(.A1(new_n1006_), .A2(\a[106] ), .B(new_n1040_), .ZN(new_n1074_));
  OAI21_X1   g00882(.A1(new_n1073_), .A2(new_n1074_), .B(\asqrt[54] ), .ZN(new_n1075_));
  AOI21_X1   g00883(.A1(\asqrt[53] ), .A2(new_n1042_), .B(new_n1046_), .ZN(new_n1076_));
  NOR3_X1    g00884(.A1(new_n1006_), .A2(\a[106] ), .A3(\a[107] ), .ZN(new_n1077_));
  INV_X1     g00885(.I(new_n1050_), .ZN(new_n1078_));
  NOR2_X1    g00886(.A1(new_n1006_), .A2(new_n1078_), .ZN(new_n1079_));
  NOR3_X1    g00887(.A1(new_n1077_), .A2(new_n1076_), .A3(new_n1079_), .ZN(new_n1080_));
  NAND3_X1   g00888(.A1(new_n1075_), .A2(new_n1080_), .A3(new_n744_), .ZN(new_n1081_));
  NAND2_X1   g00889(.A1(new_n1081_), .A2(new_n1072_), .ZN(new_n1082_));
  NAND3_X1   g00890(.A1(new_n1082_), .A2(new_n634_), .A3(new_n1054_), .ZN(new_n1083_));
  AOI21_X1   g00891(.A1(new_n1082_), .A2(new_n1054_), .B(new_n634_), .ZN(new_n1084_));
  AOI21_X1   g00892(.A1(new_n1029_), .A2(new_n1083_), .B(new_n1084_), .ZN(new_n1085_));
  AOI21_X1   g00893(.A1(new_n1085_), .A2(new_n531_), .B(new_n1071_), .ZN(new_n1086_));
  NOR3_X1    g00894(.A1(new_n1086_), .A2(\asqrt[58] ), .A3(new_n1059_), .ZN(new_n1087_));
  OAI21_X1   g00895(.A1(new_n1086_), .A2(new_n1059_), .B(\asqrt[58] ), .ZN(new_n1088_));
  OAI21_X1   g00896(.A1(new_n1017_), .A2(new_n1087_), .B(new_n1088_), .ZN(new_n1089_));
  OAI21_X1   g00897(.A1(new_n1089_), .A2(\asqrt[59] ), .B(new_n1015_), .ZN(new_n1090_));
  AOI21_X1   g00898(.A1(new_n1090_), .A2(new_n1067_), .B(new_n266_), .ZN(new_n1091_));
  OAI21_X1   g00899(.A1(new_n1070_), .A2(new_n1091_), .B(\asqrt[61] ), .ZN(new_n1092_));
  AOI21_X1   g00900(.A1(new_n963_), .A2(new_n957_), .B(\asqrt[53] ), .ZN(new_n1093_));
  XOR2_X1    g00901(.A1(new_n1093_), .A2(new_n928_), .Z(new_n1094_));
  OAI21_X1   g00902(.A1(new_n1016_), .A2(new_n1065_), .B(new_n1067_), .ZN(new_n1095_));
  OAI21_X1   g00903(.A1(new_n1095_), .A2(\asqrt[60] ), .B(new_n1012_), .ZN(new_n1096_));
  OAI21_X1   g00904(.A1(new_n1066_), .A2(new_n1068_), .B(\asqrt[60] ), .ZN(new_n1097_));
  NAND3_X1   g00905(.A1(new_n1096_), .A2(new_n239_), .A3(new_n1097_), .ZN(new_n1098_));
  NAND2_X1   g00906(.A1(new_n1098_), .A2(new_n1094_), .ZN(new_n1099_));
  NAND2_X1   g00907(.A1(new_n1099_), .A2(new_n1092_), .ZN(new_n1100_));
  AOI21_X1   g00908(.A1(new_n1096_), .A2(new_n1097_), .B(new_n239_), .ZN(new_n1101_));
  NAND3_X1   g00909(.A1(new_n1090_), .A2(new_n266_), .A3(new_n1067_), .ZN(new_n1102_));
  AOI21_X1   g00910(.A1(new_n1012_), .A2(new_n1102_), .B(new_n1091_), .ZN(new_n1103_));
  INV_X1     g00911(.I(new_n1094_), .ZN(new_n1104_));
  AOI21_X1   g00912(.A1(new_n1103_), .A2(new_n239_), .B(new_n1104_), .ZN(new_n1105_));
  OAI21_X1   g00913(.A1(new_n1105_), .A2(new_n1101_), .B(new_n201_), .ZN(new_n1106_));
  NAND3_X1   g00914(.A1(new_n1099_), .A2(\asqrt[62] ), .A3(new_n1092_), .ZN(new_n1107_));
  AOI21_X1   g00915(.A1(new_n956_), .A2(new_n997_), .B(\asqrt[53] ), .ZN(new_n1108_));
  XOR2_X1    g00916(.A1(new_n1108_), .A2(new_n960_), .Z(new_n1109_));
  INV_X1     g00917(.I(new_n1109_), .ZN(new_n1110_));
  AOI22_X1   g00918(.A1(new_n1106_), .A2(new_n1107_), .B1(new_n1100_), .B2(new_n1110_), .ZN(new_n1111_));
  NOR2_X1    g00919(.A1(new_n975_), .A2(new_n926_), .ZN(new_n1112_));
  OAI21_X1   g00920(.A1(\asqrt[53] ), .A2(new_n1112_), .B(new_n982_), .ZN(new_n1113_));
  INV_X1     g00921(.I(new_n1113_), .ZN(new_n1114_));
  OAI21_X1   g00922(.A1(new_n1111_), .A2(new_n1009_), .B(new_n1114_), .ZN(new_n1115_));
  AOI21_X1   g00923(.A1(new_n1094_), .A2(new_n1098_), .B(new_n1101_), .ZN(new_n1116_));
  AOI21_X1   g00924(.A1(new_n1116_), .A2(new_n201_), .B(new_n1110_), .ZN(new_n1117_));
  OAI21_X1   g00925(.A1(new_n1116_), .A2(new_n201_), .B(new_n1009_), .ZN(new_n1118_));
  OR2_X2     g00926(.A1(new_n1117_), .A2(new_n1118_), .Z(new_n1119_));
  NAND2_X1   g00927(.A1(new_n975_), .A2(new_n925_), .ZN(new_n1120_));
  NAND2_X1   g00928(.A1(new_n1001_), .A2(new_n926_), .ZN(new_n1121_));
  AOI21_X1   g00929(.A1(new_n1121_), .A2(new_n1120_), .B(new_n193_), .ZN(new_n1122_));
  OAI21_X1   g00930(.A1(\asqrt[53] ), .A2(new_n926_), .B(new_n1122_), .ZN(new_n1123_));
  INV_X1     g00931(.I(new_n1034_), .ZN(new_n1124_));
  NOR3_X1    g00932(.A1(new_n1005_), .A2(new_n925_), .A3(new_n989_), .ZN(new_n1125_));
  NAND2_X1   g00933(.A1(new_n1124_), .A2(new_n1125_), .ZN(new_n1126_));
  NAND2_X1   g00934(.A1(new_n1126_), .A2(new_n1123_), .ZN(new_n1127_));
  INV_X1     g00935(.I(new_n1127_), .ZN(new_n1128_));
  NAND4_X1   g00936(.A1(new_n1115_), .A2(new_n193_), .A3(new_n1119_), .A4(new_n1128_), .ZN(\asqrt[52] ));
  NOR2_X1    g00937(.A1(new_n1087_), .A2(new_n1064_), .ZN(new_n1130_));
  NOR2_X1    g00938(.A1(\asqrt[52] ), .A2(new_n1130_), .ZN(new_n1131_));
  XOR2_X1    g00939(.A1(new_n1131_), .A2(new_n993_), .Z(new_n1132_));
  AOI21_X1   g00940(.A1(new_n1058_), .A2(new_n1063_), .B(\asqrt[52] ), .ZN(new_n1133_));
  XOR2_X1    g00941(.A1(new_n1133_), .A2(new_n1019_), .Z(new_n1134_));
  AOI21_X1   g00942(.A1(new_n1083_), .A2(new_n1057_), .B(\asqrt[52] ), .ZN(new_n1135_));
  XOR2_X1    g00943(.A1(new_n1135_), .A2(new_n1029_), .Z(new_n1136_));
  AOI21_X1   g00944(.A1(new_n1081_), .A2(new_n1054_), .B(\asqrt[52] ), .ZN(new_n1137_));
  XOR2_X1    g00945(.A1(new_n1137_), .A2(new_n1072_), .Z(new_n1138_));
  INV_X1     g00946(.I(new_n1138_), .ZN(new_n1139_));
  NOR2_X1    g00947(.A1(new_n1006_), .A2(\a[106] ), .ZN(new_n1140_));
  INV_X1     g00948(.I(new_n1140_), .ZN(new_n1141_));
  NOR2_X1    g00949(.A1(new_n1046_), .A2(\a[106] ), .ZN(new_n1142_));
  AOI22_X1   g00950(.A1(new_n1141_), .A2(new_n1046_), .B1(\asqrt[53] ), .B2(new_n1142_), .ZN(new_n1143_));
  INV_X1     g00951(.I(new_n1143_), .ZN(new_n1144_));
  AOI21_X1   g00952(.A1(new_n1099_), .A2(new_n1092_), .B(\asqrt[62] ), .ZN(new_n1145_));
  NOR3_X1    g00953(.A1(new_n1105_), .A2(new_n201_), .A3(new_n1101_), .ZN(new_n1146_));
  OAI22_X1   g00954(.A1(new_n1146_), .A2(new_n1145_), .B1(new_n1116_), .B2(new_n1109_), .ZN(new_n1147_));
  AOI21_X1   g00955(.A1(new_n1147_), .A2(new_n1008_), .B(new_n1113_), .ZN(new_n1148_));
  NOR2_X1    g00956(.A1(new_n1117_), .A2(new_n1118_), .ZN(new_n1149_));
  NOR4_X1    g00957(.A1(new_n1148_), .A2(\asqrt[63] ), .A3(new_n1149_), .A4(new_n1127_), .ZN(new_n1150_));
  NOR2_X1    g00958(.A1(new_n1044_), .A2(new_n1079_), .ZN(new_n1151_));
  NOR2_X1    g00959(.A1(new_n1150_), .A2(new_n1151_), .ZN(new_n1152_));
  NOR2_X1    g00960(.A1(new_n1152_), .A2(new_n1144_), .ZN(new_n1153_));
  NOR3_X1    g00961(.A1(new_n1150_), .A2(new_n1143_), .A3(new_n1151_), .ZN(new_n1154_));
  NOR2_X1    g00962(.A1(new_n1153_), .A2(new_n1154_), .ZN(new_n1155_));
  INV_X1     g00963(.I(new_n1155_), .ZN(new_n1156_));
  NAND2_X1   g00964(.A1(new_n1115_), .A2(new_n193_), .ZN(new_n1157_));
  NAND3_X1   g00965(.A1(new_n1126_), .A2(new_n1123_), .A3(\asqrt[53] ), .ZN(new_n1158_));
  NOR3_X1    g00966(.A1(new_n1157_), .A2(new_n1149_), .A3(new_n1158_), .ZN(new_n1159_));
  NOR2_X1    g00967(.A1(new_n1150_), .A2(new_n1040_), .ZN(new_n1160_));
  OAI21_X1   g00968(.A1(new_n1160_), .A2(new_n1159_), .B(new_n1042_), .ZN(new_n1161_));
  INV_X1     g00969(.I(new_n1161_), .ZN(new_n1162_));
  NOR3_X1    g00970(.A1(new_n1160_), .A2(new_n1159_), .A3(new_n1042_), .ZN(new_n1163_));
  NOR2_X1    g00971(.A1(new_n1162_), .A2(new_n1163_), .ZN(new_n1164_));
  INV_X1     g00972(.I(\a[104] ), .ZN(new_n1165_));
  NOR2_X1    g00973(.A1(\a[102] ), .A2(\a[103] ), .ZN(new_n1166_));
  NOR3_X1    g00974(.A1(new_n1150_), .A2(new_n1165_), .A3(new_n1166_), .ZN(new_n1167_));
  INV_X1     g00975(.I(new_n1166_), .ZN(new_n1168_));
  AOI21_X1   g00976(.A1(new_n1150_), .A2(\a[104] ), .B(new_n1168_), .ZN(new_n1169_));
  OAI21_X1   g00977(.A1(new_n1167_), .A2(new_n1169_), .B(\asqrt[53] ), .ZN(new_n1170_));
  INV_X1     g00978(.I(\a[105] ), .ZN(new_n1171_));
  AOI21_X1   g00979(.A1(\asqrt[52] ), .A2(new_n1165_), .B(new_n1171_), .ZN(new_n1172_));
  NOR3_X1    g00980(.A1(new_n1150_), .A2(\a[104] ), .A3(\a[105] ), .ZN(new_n1173_));
  NAND2_X1   g00981(.A1(new_n1166_), .A2(new_n1165_), .ZN(new_n1174_));
  AND4_X2    g00982(.A1(new_n982_), .A2(new_n985_), .A3(new_n988_), .A4(new_n1174_), .Z(new_n1175_));
  AOI21_X1   g00983(.A1(new_n1124_), .A2(new_n1175_), .B(new_n1165_), .ZN(new_n1176_));
  INV_X1     g00984(.I(new_n1176_), .ZN(new_n1177_));
  NOR2_X1    g00985(.A1(new_n1150_), .A2(new_n1177_), .ZN(new_n1178_));
  NOR3_X1    g00986(.A1(new_n1173_), .A2(new_n1172_), .A3(new_n1178_), .ZN(new_n1179_));
  NAND3_X1   g00987(.A1(new_n1170_), .A2(new_n1179_), .A3(new_n860_), .ZN(new_n1180_));
  AOI21_X1   g00988(.A1(new_n1170_), .A2(new_n1179_), .B(new_n860_), .ZN(new_n1181_));
  AOI21_X1   g00989(.A1(new_n1164_), .A2(new_n1180_), .B(new_n1181_), .ZN(new_n1182_));
  AOI21_X1   g00990(.A1(new_n1182_), .A2(new_n744_), .B(new_n1156_), .ZN(new_n1183_));
  NOR2_X1    g00991(.A1(new_n1182_), .A2(new_n744_), .ZN(new_n1184_));
  NOR3_X1    g00992(.A1(new_n1183_), .A2(new_n1184_), .A3(\asqrt[56] ), .ZN(new_n1185_));
  OAI21_X1   g00993(.A1(new_n1183_), .A2(new_n1184_), .B(\asqrt[56] ), .ZN(new_n1186_));
  OAI21_X1   g00994(.A1(new_n1139_), .A2(new_n1185_), .B(new_n1186_), .ZN(new_n1187_));
  OAI21_X1   g00995(.A1(new_n1187_), .A2(\asqrt[57] ), .B(new_n1136_), .ZN(new_n1188_));
  NOR2_X1    g00996(.A1(new_n1185_), .A2(new_n1139_), .ZN(new_n1189_));
  INV_X1     g00997(.I(new_n1163_), .ZN(new_n1190_));
  NAND2_X1   g00998(.A1(new_n1190_), .A2(new_n1161_), .ZN(new_n1191_));
  NAND3_X1   g00999(.A1(\asqrt[52] ), .A2(\a[104] ), .A3(new_n1168_), .ZN(new_n1192_));
  OAI21_X1   g01000(.A1(\asqrt[52] ), .A2(new_n1165_), .B(new_n1166_), .ZN(new_n1193_));
  AOI21_X1   g01001(.A1(new_n1193_), .A2(new_n1192_), .B(new_n1006_), .ZN(new_n1194_));
  OAI21_X1   g01002(.A1(new_n1150_), .A2(\a[104] ), .B(\a[105] ), .ZN(new_n1195_));
  NAND3_X1   g01003(.A1(\asqrt[52] ), .A2(new_n1165_), .A3(new_n1171_), .ZN(new_n1196_));
  NAND2_X1   g01004(.A1(\asqrt[52] ), .A2(new_n1176_), .ZN(new_n1197_));
  NAND3_X1   g01005(.A1(new_n1195_), .A2(new_n1196_), .A3(new_n1197_), .ZN(new_n1198_));
  NOR3_X1    g01006(.A1(new_n1194_), .A2(new_n1198_), .A3(\asqrt[54] ), .ZN(new_n1199_));
  OAI21_X1   g01007(.A1(new_n1194_), .A2(new_n1198_), .B(\asqrt[54] ), .ZN(new_n1200_));
  OAI21_X1   g01008(.A1(new_n1191_), .A2(new_n1199_), .B(new_n1200_), .ZN(new_n1201_));
  OAI21_X1   g01009(.A1(new_n1201_), .A2(\asqrt[55] ), .B(new_n1155_), .ZN(new_n1202_));
  NAND2_X1   g01010(.A1(new_n1201_), .A2(\asqrt[55] ), .ZN(new_n1203_));
  AOI21_X1   g01011(.A1(new_n1202_), .A2(new_n1203_), .B(new_n634_), .ZN(new_n1204_));
  OAI21_X1   g01012(.A1(new_n1189_), .A2(new_n1204_), .B(\asqrt[57] ), .ZN(new_n1205_));
  NAND3_X1   g01013(.A1(new_n1188_), .A2(new_n423_), .A3(new_n1205_), .ZN(new_n1206_));
  NAND2_X1   g01014(.A1(new_n1206_), .A2(new_n1134_), .ZN(new_n1207_));
  INV_X1     g01015(.I(new_n1136_), .ZN(new_n1208_));
  NAND3_X1   g01016(.A1(new_n1202_), .A2(new_n1203_), .A3(new_n634_), .ZN(new_n1209_));
  AOI21_X1   g01017(.A1(new_n1138_), .A2(new_n1209_), .B(new_n1204_), .ZN(new_n1210_));
  AOI21_X1   g01018(.A1(new_n1210_), .A2(new_n531_), .B(new_n1208_), .ZN(new_n1211_));
  NAND2_X1   g01019(.A1(new_n1209_), .A2(new_n1138_), .ZN(new_n1212_));
  AOI21_X1   g01020(.A1(new_n1212_), .A2(new_n1186_), .B(new_n531_), .ZN(new_n1213_));
  OAI21_X1   g01021(.A1(new_n1211_), .A2(new_n1213_), .B(\asqrt[58] ), .ZN(new_n1214_));
  NAND3_X1   g01022(.A1(new_n1207_), .A2(new_n337_), .A3(new_n1214_), .ZN(new_n1215_));
  INV_X1     g01023(.I(new_n1134_), .ZN(new_n1216_));
  NOR3_X1    g01024(.A1(new_n1211_), .A2(\asqrt[58] ), .A3(new_n1213_), .ZN(new_n1217_));
  OAI21_X1   g01025(.A1(new_n1216_), .A2(new_n1217_), .B(new_n1214_), .ZN(new_n1218_));
  NAND2_X1   g01026(.A1(new_n1218_), .A2(\asqrt[59] ), .ZN(new_n1219_));
  NOR2_X1    g01027(.A1(new_n1100_), .A2(\asqrt[62] ), .ZN(new_n1220_));
  NAND2_X1   g01028(.A1(new_n1100_), .A2(\asqrt[62] ), .ZN(new_n1221_));
  INV_X1     g01029(.I(new_n1221_), .ZN(new_n1222_));
  NOR2_X1    g01030(.A1(new_n1222_), .A2(new_n1220_), .ZN(new_n1223_));
  XOR2_X1    g01031(.A1(new_n1108_), .A2(new_n960_), .Z(new_n1224_));
  OAI21_X1   g01032(.A1(\asqrt[52] ), .A2(new_n1223_), .B(new_n1224_), .ZN(new_n1225_));
  INV_X1     g01033(.I(new_n1225_), .ZN(new_n1226_));
  NOR2_X1    g01034(.A1(new_n1068_), .A2(new_n1065_), .ZN(new_n1227_));
  NOR2_X1    g01035(.A1(\asqrt[52] ), .A2(new_n1227_), .ZN(new_n1228_));
  XOR2_X1    g01036(.A1(new_n1228_), .A2(new_n1015_), .Z(new_n1229_));
  INV_X1     g01037(.I(new_n1229_), .ZN(new_n1230_));
  AOI21_X1   g01038(.A1(new_n1207_), .A2(new_n1214_), .B(new_n337_), .ZN(new_n1231_));
  AOI21_X1   g01039(.A1(new_n1132_), .A2(new_n1215_), .B(new_n1231_), .ZN(new_n1232_));
  AOI21_X1   g01040(.A1(new_n1232_), .A2(new_n266_), .B(new_n1230_), .ZN(new_n1233_));
  OAI21_X1   g01041(.A1(new_n1218_), .A2(\asqrt[59] ), .B(new_n1132_), .ZN(new_n1234_));
  AOI21_X1   g01042(.A1(new_n1234_), .A2(new_n1219_), .B(new_n266_), .ZN(new_n1235_));
  OAI21_X1   g01043(.A1(new_n1233_), .A2(new_n1235_), .B(\asqrt[61] ), .ZN(new_n1236_));
  AOI21_X1   g01044(.A1(new_n1102_), .A2(new_n1097_), .B(\asqrt[52] ), .ZN(new_n1237_));
  XOR2_X1    g01045(.A1(new_n1237_), .A2(new_n1012_), .Z(new_n1238_));
  INV_X1     g01046(.I(new_n1238_), .ZN(new_n1239_));
  NOR3_X1    g01047(.A1(new_n1233_), .A2(\asqrt[61] ), .A3(new_n1235_), .ZN(new_n1240_));
  OAI21_X1   g01048(.A1(new_n1239_), .A2(new_n1240_), .B(new_n1236_), .ZN(new_n1241_));
  NAND3_X1   g01049(.A1(new_n1234_), .A2(new_n1219_), .A3(new_n266_), .ZN(new_n1242_));
  NAND2_X1   g01050(.A1(new_n1242_), .A2(new_n1229_), .ZN(new_n1243_));
  INV_X1     g01051(.I(new_n1132_), .ZN(new_n1244_));
  AOI21_X1   g01052(.A1(new_n1188_), .A2(new_n1205_), .B(new_n423_), .ZN(new_n1245_));
  AOI21_X1   g01053(.A1(new_n1134_), .A2(new_n1206_), .B(new_n1245_), .ZN(new_n1246_));
  AOI21_X1   g01054(.A1(new_n1246_), .A2(new_n337_), .B(new_n1244_), .ZN(new_n1247_));
  OAI21_X1   g01055(.A1(new_n1247_), .A2(new_n1231_), .B(\asqrt[60] ), .ZN(new_n1248_));
  AOI21_X1   g01056(.A1(new_n1243_), .A2(new_n1248_), .B(new_n239_), .ZN(new_n1249_));
  AOI21_X1   g01057(.A1(new_n1229_), .A2(new_n1242_), .B(new_n1235_), .ZN(new_n1250_));
  AOI21_X1   g01058(.A1(new_n1250_), .A2(new_n239_), .B(new_n1239_), .ZN(new_n1251_));
  OAI21_X1   g01059(.A1(new_n1251_), .A2(new_n1249_), .B(new_n201_), .ZN(new_n1252_));
  NOR3_X1    g01060(.A1(new_n1247_), .A2(\asqrt[60] ), .A3(new_n1231_), .ZN(new_n1253_));
  OAI21_X1   g01061(.A1(new_n1230_), .A2(new_n1253_), .B(new_n1248_), .ZN(new_n1254_));
  OAI21_X1   g01062(.A1(new_n1254_), .A2(\asqrt[61] ), .B(new_n1238_), .ZN(new_n1255_));
  NAND3_X1   g01063(.A1(new_n1255_), .A2(\asqrt[62] ), .A3(new_n1236_), .ZN(new_n1256_));
  AOI21_X1   g01064(.A1(new_n1092_), .A2(new_n1098_), .B(\asqrt[52] ), .ZN(new_n1257_));
  XOR2_X1    g01065(.A1(new_n1257_), .A2(new_n1094_), .Z(new_n1258_));
  INV_X1     g01066(.I(new_n1258_), .ZN(new_n1259_));
  AOI22_X1   g01067(.A1(new_n1256_), .A2(new_n1252_), .B1(new_n1241_), .B2(new_n1259_), .ZN(new_n1260_));
  NOR2_X1    g01068(.A1(new_n1111_), .A2(new_n1009_), .ZN(new_n1261_));
  OAI21_X1   g01069(.A1(\asqrt[52] ), .A2(new_n1261_), .B(new_n1119_), .ZN(new_n1262_));
  INV_X1     g01070(.I(new_n1262_), .ZN(new_n1263_));
  OAI21_X1   g01071(.A1(new_n1260_), .A2(new_n1226_), .B(new_n1263_), .ZN(new_n1264_));
  OAI21_X1   g01072(.A1(new_n1241_), .A2(\asqrt[62] ), .B(new_n1258_), .ZN(new_n1265_));
  NAND2_X1   g01073(.A1(new_n1241_), .A2(\asqrt[62] ), .ZN(new_n1266_));
  NAND3_X1   g01074(.A1(new_n1265_), .A2(new_n1266_), .A3(new_n1226_), .ZN(new_n1267_));
  NAND2_X1   g01075(.A1(new_n1150_), .A2(new_n1008_), .ZN(new_n1268_));
  XOR2_X1    g01076(.A1(new_n1111_), .A2(new_n1009_), .Z(new_n1269_));
  NAND3_X1   g01077(.A1(new_n1268_), .A2(\asqrt[63] ), .A3(new_n1269_), .ZN(new_n1270_));
  INV_X1     g01078(.I(new_n1157_), .ZN(new_n1271_));
  NAND4_X1   g01079(.A1(new_n1271_), .A2(new_n1009_), .A3(new_n1119_), .A4(new_n1128_), .ZN(new_n1272_));
  NAND2_X1   g01080(.A1(new_n1270_), .A2(new_n1272_), .ZN(new_n1273_));
  INV_X1     g01081(.I(new_n1273_), .ZN(new_n1274_));
  NAND4_X1   g01082(.A1(new_n1264_), .A2(new_n193_), .A3(new_n1267_), .A4(new_n1274_), .ZN(\asqrt[51] ));
  AOI21_X1   g01083(.A1(new_n1215_), .A2(new_n1219_), .B(\asqrt[51] ), .ZN(new_n1276_));
  XOR2_X1    g01084(.A1(new_n1276_), .A2(new_n1132_), .Z(new_n1277_));
  AOI21_X1   g01085(.A1(new_n1206_), .A2(new_n1214_), .B(\asqrt[51] ), .ZN(new_n1278_));
  XOR2_X1    g01086(.A1(new_n1278_), .A2(new_n1134_), .Z(new_n1279_));
  NAND2_X1   g01087(.A1(new_n1210_), .A2(new_n531_), .ZN(new_n1280_));
  AOI21_X1   g01088(.A1(new_n1280_), .A2(new_n1205_), .B(\asqrt[51] ), .ZN(new_n1281_));
  XOR2_X1    g01089(.A1(new_n1281_), .A2(new_n1136_), .Z(new_n1282_));
  AOI21_X1   g01090(.A1(new_n1209_), .A2(new_n1186_), .B(\asqrt[51] ), .ZN(new_n1283_));
  XOR2_X1    g01091(.A1(new_n1283_), .A2(new_n1138_), .Z(new_n1284_));
  INV_X1     g01092(.I(new_n1284_), .ZN(new_n1285_));
  NAND2_X1   g01093(.A1(new_n1182_), .A2(new_n744_), .ZN(new_n1286_));
  AOI21_X1   g01094(.A1(new_n1286_), .A2(new_n1203_), .B(\asqrt[51] ), .ZN(new_n1287_));
  XOR2_X1    g01095(.A1(new_n1287_), .A2(new_n1155_), .Z(new_n1288_));
  INV_X1     g01096(.I(new_n1288_), .ZN(new_n1289_));
  AOI21_X1   g01097(.A1(new_n1180_), .A2(new_n1200_), .B(\asqrt[51] ), .ZN(new_n1290_));
  XOR2_X1    g01098(.A1(new_n1290_), .A2(new_n1164_), .Z(new_n1291_));
  NOR2_X1    g01099(.A1(new_n1150_), .A2(\a[104] ), .ZN(new_n1292_));
  INV_X1     g01100(.I(new_n1292_), .ZN(new_n1293_));
  NOR2_X1    g01101(.A1(new_n1171_), .A2(\a[104] ), .ZN(new_n1294_));
  AOI22_X1   g01102(.A1(new_n1293_), .A2(new_n1171_), .B1(\asqrt[52] ), .B2(new_n1294_), .ZN(new_n1295_));
  INV_X1     g01103(.I(new_n1295_), .ZN(new_n1296_));
  NOR2_X1    g01104(.A1(new_n1251_), .A2(new_n1249_), .ZN(new_n1297_));
  AOI21_X1   g01105(.A1(new_n1255_), .A2(new_n1236_), .B(\asqrt[62] ), .ZN(new_n1298_));
  NOR3_X1    g01106(.A1(new_n1251_), .A2(new_n201_), .A3(new_n1249_), .ZN(new_n1299_));
  OAI22_X1   g01107(.A1(new_n1298_), .A2(new_n1299_), .B1(new_n1297_), .B2(new_n1258_), .ZN(new_n1300_));
  AOI21_X1   g01108(.A1(new_n1300_), .A2(new_n1225_), .B(new_n1262_), .ZN(new_n1301_));
  AOI21_X1   g01109(.A1(new_n1297_), .A2(new_n201_), .B(new_n1259_), .ZN(new_n1302_));
  NOR2_X1    g01110(.A1(new_n1297_), .A2(new_n201_), .ZN(new_n1303_));
  NOR3_X1    g01111(.A1(new_n1302_), .A2(new_n1303_), .A3(new_n1225_), .ZN(new_n1304_));
  NOR4_X1    g01112(.A1(new_n1301_), .A2(\asqrt[63] ), .A3(new_n1304_), .A4(new_n1273_), .ZN(new_n1305_));
  NOR2_X1    g01113(.A1(new_n1194_), .A2(new_n1178_), .ZN(new_n1306_));
  NOR2_X1    g01114(.A1(new_n1305_), .A2(new_n1306_), .ZN(new_n1307_));
  NOR2_X1    g01115(.A1(new_n1307_), .A2(new_n1296_), .ZN(new_n1308_));
  NOR2_X1    g01116(.A1(new_n1306_), .A2(new_n1295_), .ZN(new_n1309_));
  AOI21_X1   g01117(.A1(\asqrt[51] ), .A2(new_n1309_), .B(new_n1308_), .ZN(new_n1310_));
  NAND3_X1   g01118(.A1(new_n1270_), .A2(\asqrt[52] ), .A3(new_n1272_), .ZN(new_n1311_));
  NOR4_X1    g01119(.A1(new_n1301_), .A2(\asqrt[63] ), .A3(new_n1304_), .A4(new_n1311_), .ZN(new_n1312_));
  INV_X1     g01120(.I(new_n1312_), .ZN(new_n1313_));
  NAND2_X1   g01121(.A1(\asqrt[51] ), .A2(new_n1166_), .ZN(new_n1314_));
  AOI21_X1   g01122(.A1(new_n1314_), .A2(new_n1313_), .B(\a[104] ), .ZN(new_n1315_));
  NOR2_X1    g01123(.A1(new_n1305_), .A2(new_n1168_), .ZN(new_n1316_));
  NOR3_X1    g01124(.A1(new_n1316_), .A2(new_n1165_), .A3(new_n1312_), .ZN(new_n1317_));
  OR2_X2     g01125(.A1(new_n1317_), .A2(new_n1315_), .Z(new_n1318_));
  NOR2_X1    g01126(.A1(\a[100] ), .A2(\a[101] ), .ZN(new_n1319_));
  INV_X1     g01127(.I(new_n1319_), .ZN(new_n1320_));
  NAND3_X1   g01128(.A1(\asqrt[51] ), .A2(\a[102] ), .A3(new_n1320_), .ZN(new_n1321_));
  INV_X1     g01129(.I(\a[102] ), .ZN(new_n1322_));
  OAI21_X1   g01130(.A1(\asqrt[51] ), .A2(new_n1322_), .B(new_n1319_), .ZN(new_n1323_));
  AOI21_X1   g01131(.A1(new_n1323_), .A2(new_n1321_), .B(new_n1150_), .ZN(new_n1324_));
  OAI21_X1   g01132(.A1(new_n1305_), .A2(\a[102] ), .B(\a[103] ), .ZN(new_n1325_));
  INV_X1     g01133(.I(\a[103] ), .ZN(new_n1326_));
  NAND3_X1   g01134(.A1(\asqrt[51] ), .A2(new_n1322_), .A3(new_n1326_), .ZN(new_n1327_));
  NAND2_X1   g01135(.A1(new_n1319_), .A2(new_n1322_), .ZN(new_n1328_));
  AND4_X2    g01136(.A1(new_n1119_), .A2(new_n1123_), .A3(new_n1126_), .A4(new_n1328_), .Z(new_n1329_));
  AOI21_X1   g01137(.A1(new_n1271_), .A2(new_n1329_), .B(new_n1322_), .ZN(new_n1330_));
  NAND2_X1   g01138(.A1(\asqrt[51] ), .A2(new_n1330_), .ZN(new_n1331_));
  NAND3_X1   g01139(.A1(new_n1325_), .A2(new_n1327_), .A3(new_n1331_), .ZN(new_n1332_));
  NOR3_X1    g01140(.A1(new_n1324_), .A2(new_n1332_), .A3(\asqrt[53] ), .ZN(new_n1333_));
  OAI21_X1   g01141(.A1(new_n1324_), .A2(new_n1332_), .B(\asqrt[53] ), .ZN(new_n1334_));
  OAI21_X1   g01142(.A1(new_n1318_), .A2(new_n1333_), .B(new_n1334_), .ZN(new_n1335_));
  OAI21_X1   g01143(.A1(new_n1335_), .A2(\asqrt[54] ), .B(new_n1310_), .ZN(new_n1336_));
  NAND2_X1   g01144(.A1(new_n1335_), .A2(\asqrt[54] ), .ZN(new_n1337_));
  NAND3_X1   g01145(.A1(new_n1336_), .A2(new_n1337_), .A3(new_n744_), .ZN(new_n1338_));
  AOI21_X1   g01146(.A1(new_n1336_), .A2(new_n1337_), .B(new_n744_), .ZN(new_n1339_));
  AOI21_X1   g01147(.A1(new_n1291_), .A2(new_n1338_), .B(new_n1339_), .ZN(new_n1340_));
  AOI21_X1   g01148(.A1(new_n1340_), .A2(new_n634_), .B(new_n1289_), .ZN(new_n1341_));
  NAND2_X1   g01149(.A1(new_n1338_), .A2(new_n1291_), .ZN(new_n1342_));
  INV_X1     g01150(.I(new_n1339_), .ZN(new_n1343_));
  AOI21_X1   g01151(.A1(new_n1342_), .A2(new_n1343_), .B(new_n634_), .ZN(new_n1344_));
  NOR3_X1    g01152(.A1(new_n1341_), .A2(\asqrt[57] ), .A3(new_n1344_), .ZN(new_n1345_));
  OAI21_X1   g01153(.A1(new_n1341_), .A2(new_n1344_), .B(\asqrt[57] ), .ZN(new_n1346_));
  OAI21_X1   g01154(.A1(new_n1285_), .A2(new_n1345_), .B(new_n1346_), .ZN(new_n1347_));
  OAI21_X1   g01155(.A1(new_n1347_), .A2(\asqrt[58] ), .B(new_n1282_), .ZN(new_n1348_));
  NOR2_X1    g01156(.A1(new_n1345_), .A2(new_n1285_), .ZN(new_n1349_));
  INV_X1     g01157(.I(new_n1346_), .ZN(new_n1350_));
  OAI21_X1   g01158(.A1(new_n1349_), .A2(new_n1350_), .B(\asqrt[58] ), .ZN(new_n1351_));
  NAND3_X1   g01159(.A1(new_n1348_), .A2(new_n337_), .A3(new_n1351_), .ZN(new_n1352_));
  NAND2_X1   g01160(.A1(new_n1352_), .A2(new_n1279_), .ZN(new_n1353_));
  INV_X1     g01161(.I(new_n1282_), .ZN(new_n1354_));
  NOR2_X1    g01162(.A1(new_n1349_), .A2(new_n1350_), .ZN(new_n1355_));
  AOI21_X1   g01163(.A1(new_n1355_), .A2(new_n423_), .B(new_n1354_), .ZN(new_n1356_));
  INV_X1     g01164(.I(new_n1291_), .ZN(new_n1357_));
  NOR2_X1    g01165(.A1(new_n1317_), .A2(new_n1315_), .ZN(new_n1358_));
  NOR3_X1    g01166(.A1(new_n1305_), .A2(new_n1322_), .A3(new_n1319_), .ZN(new_n1359_));
  AOI21_X1   g01167(.A1(new_n1305_), .A2(\a[102] ), .B(new_n1320_), .ZN(new_n1360_));
  OAI21_X1   g01168(.A1(new_n1359_), .A2(new_n1360_), .B(\asqrt[52] ), .ZN(new_n1361_));
  AOI21_X1   g01169(.A1(\asqrt[51] ), .A2(new_n1322_), .B(new_n1326_), .ZN(new_n1362_));
  NOR3_X1    g01170(.A1(new_n1305_), .A2(\a[102] ), .A3(\a[103] ), .ZN(new_n1363_));
  INV_X1     g01171(.I(new_n1330_), .ZN(new_n1364_));
  NOR2_X1    g01172(.A1(new_n1305_), .A2(new_n1364_), .ZN(new_n1365_));
  NOR3_X1    g01173(.A1(new_n1363_), .A2(new_n1362_), .A3(new_n1365_), .ZN(new_n1366_));
  NAND3_X1   g01174(.A1(new_n1361_), .A2(new_n1366_), .A3(new_n1006_), .ZN(new_n1367_));
  NAND2_X1   g01175(.A1(new_n1367_), .A2(new_n1358_), .ZN(new_n1368_));
  NAND3_X1   g01176(.A1(new_n1368_), .A2(new_n860_), .A3(new_n1334_), .ZN(new_n1369_));
  AOI21_X1   g01177(.A1(new_n1368_), .A2(new_n1334_), .B(new_n860_), .ZN(new_n1370_));
  AOI21_X1   g01178(.A1(new_n1310_), .A2(new_n1369_), .B(new_n1370_), .ZN(new_n1371_));
  AOI21_X1   g01179(.A1(new_n1371_), .A2(new_n744_), .B(new_n1357_), .ZN(new_n1372_));
  NOR3_X1    g01180(.A1(new_n1372_), .A2(\asqrt[56] ), .A3(new_n1339_), .ZN(new_n1373_));
  OAI21_X1   g01181(.A1(new_n1372_), .A2(new_n1339_), .B(\asqrt[56] ), .ZN(new_n1374_));
  OAI21_X1   g01182(.A1(new_n1289_), .A2(new_n1373_), .B(new_n1374_), .ZN(new_n1375_));
  OAI21_X1   g01183(.A1(new_n1375_), .A2(\asqrt[57] ), .B(new_n1284_), .ZN(new_n1376_));
  AOI21_X1   g01184(.A1(new_n1376_), .A2(new_n1346_), .B(new_n423_), .ZN(new_n1377_));
  OAI21_X1   g01185(.A1(new_n1356_), .A2(new_n1377_), .B(\asqrt[59] ), .ZN(new_n1378_));
  NAND3_X1   g01186(.A1(new_n1353_), .A2(new_n266_), .A3(new_n1378_), .ZN(new_n1379_));
  INV_X1     g01187(.I(new_n1279_), .ZN(new_n1380_));
  NAND3_X1   g01188(.A1(new_n1376_), .A2(new_n423_), .A3(new_n1346_), .ZN(new_n1381_));
  AOI21_X1   g01189(.A1(new_n1282_), .A2(new_n1381_), .B(new_n1377_), .ZN(new_n1382_));
  AOI21_X1   g01190(.A1(new_n1382_), .A2(new_n337_), .B(new_n1380_), .ZN(new_n1383_));
  NOR2_X1    g01191(.A1(new_n1382_), .A2(new_n337_), .ZN(new_n1384_));
  OAI21_X1   g01192(.A1(new_n1383_), .A2(new_n1384_), .B(\asqrt[60] ), .ZN(new_n1385_));
  NOR2_X1    g01193(.A1(new_n1241_), .A2(\asqrt[62] ), .ZN(new_n1386_));
  NOR2_X1    g01194(.A1(new_n1386_), .A2(new_n1303_), .ZN(new_n1387_));
  NOR2_X1    g01195(.A1(\asqrt[51] ), .A2(new_n1387_), .ZN(new_n1388_));
  XOR2_X1    g01196(.A1(new_n1257_), .A2(new_n1104_), .Z(new_n1389_));
  NOR2_X1    g01197(.A1(new_n1388_), .A2(new_n1389_), .ZN(new_n1390_));
  INV_X1     g01198(.I(new_n1277_), .ZN(new_n1391_));
  NOR3_X1    g01199(.A1(new_n1383_), .A2(new_n1384_), .A3(\asqrt[60] ), .ZN(new_n1392_));
  OAI21_X1   g01200(.A1(new_n1391_), .A2(new_n1392_), .B(new_n1385_), .ZN(new_n1393_));
  NAND2_X1   g01201(.A1(new_n1393_), .A2(\asqrt[61] ), .ZN(new_n1394_));
  AOI21_X1   g01202(.A1(new_n1242_), .A2(new_n1248_), .B(\asqrt[51] ), .ZN(new_n1395_));
  XOR2_X1    g01203(.A1(new_n1395_), .A2(new_n1229_), .Z(new_n1396_));
  OAI21_X1   g01204(.A1(new_n1393_), .A2(\asqrt[61] ), .B(new_n1396_), .ZN(new_n1397_));
  NAND2_X1   g01205(.A1(new_n1397_), .A2(new_n1394_), .ZN(new_n1398_));
  NAND2_X1   g01206(.A1(new_n1379_), .A2(new_n1277_), .ZN(new_n1399_));
  AOI21_X1   g01207(.A1(new_n1399_), .A2(new_n1385_), .B(new_n239_), .ZN(new_n1400_));
  AOI21_X1   g01208(.A1(new_n1353_), .A2(new_n1378_), .B(new_n266_), .ZN(new_n1401_));
  AOI21_X1   g01209(.A1(new_n1277_), .A2(new_n1379_), .B(new_n1401_), .ZN(new_n1402_));
  INV_X1     g01210(.I(new_n1396_), .ZN(new_n1403_));
  AOI21_X1   g01211(.A1(new_n1402_), .A2(new_n239_), .B(new_n1403_), .ZN(new_n1404_));
  OAI21_X1   g01212(.A1(new_n1404_), .A2(new_n1400_), .B(new_n201_), .ZN(new_n1405_));
  NAND3_X1   g01213(.A1(new_n1397_), .A2(new_n1394_), .A3(\asqrt[62] ), .ZN(new_n1406_));
  NOR2_X1    g01214(.A1(new_n1240_), .A2(new_n1249_), .ZN(new_n1407_));
  NOR2_X1    g01215(.A1(\asqrt[51] ), .A2(new_n1407_), .ZN(new_n1408_));
  XOR2_X1    g01216(.A1(new_n1408_), .A2(new_n1238_), .Z(new_n1409_));
  INV_X1     g01217(.I(new_n1409_), .ZN(new_n1410_));
  AOI22_X1   g01218(.A1(new_n1406_), .A2(new_n1405_), .B1(new_n1398_), .B2(new_n1410_), .ZN(new_n1411_));
  NOR2_X1    g01219(.A1(new_n1260_), .A2(new_n1226_), .ZN(new_n1412_));
  OAI21_X1   g01220(.A1(\asqrt[51] ), .A2(new_n1412_), .B(new_n1267_), .ZN(new_n1413_));
  INV_X1     g01221(.I(new_n1413_), .ZN(new_n1414_));
  OAI21_X1   g01222(.A1(new_n1411_), .A2(new_n1390_), .B(new_n1414_), .ZN(new_n1415_));
  OAI21_X1   g01223(.A1(new_n1398_), .A2(\asqrt[62] ), .B(new_n1409_), .ZN(new_n1416_));
  NAND2_X1   g01224(.A1(new_n1398_), .A2(\asqrt[62] ), .ZN(new_n1417_));
  NAND3_X1   g01225(.A1(new_n1416_), .A2(new_n1417_), .A3(new_n1390_), .ZN(new_n1418_));
  NAND2_X1   g01226(.A1(new_n1305_), .A2(new_n1225_), .ZN(new_n1419_));
  XOR2_X1    g01227(.A1(new_n1300_), .A2(new_n1225_), .Z(new_n1420_));
  NAND3_X1   g01228(.A1(new_n1419_), .A2(\asqrt[63] ), .A3(new_n1420_), .ZN(new_n1421_));
  NOR2_X1    g01229(.A1(new_n1273_), .A2(new_n1225_), .ZN(new_n1422_));
  NAND4_X1   g01230(.A1(new_n1264_), .A2(new_n193_), .A3(new_n1267_), .A4(new_n1422_), .ZN(new_n1423_));
  NAND2_X1   g01231(.A1(new_n1421_), .A2(new_n1423_), .ZN(new_n1424_));
  INV_X1     g01232(.I(new_n1424_), .ZN(new_n1425_));
  NAND4_X1   g01233(.A1(new_n1415_), .A2(new_n193_), .A3(new_n1418_), .A4(new_n1425_), .ZN(\asqrt[50] ));
  AOI21_X1   g01234(.A1(new_n1379_), .A2(new_n1385_), .B(\asqrt[50] ), .ZN(new_n1427_));
  XOR2_X1    g01235(.A1(new_n1427_), .A2(new_n1277_), .Z(new_n1428_));
  AOI21_X1   g01236(.A1(new_n1352_), .A2(new_n1378_), .B(\asqrt[50] ), .ZN(new_n1429_));
  XOR2_X1    g01237(.A1(new_n1429_), .A2(new_n1279_), .Z(new_n1430_));
  INV_X1     g01238(.I(new_n1430_), .ZN(new_n1431_));
  AOI21_X1   g01239(.A1(new_n1381_), .A2(new_n1351_), .B(\asqrt[50] ), .ZN(new_n1432_));
  XOR2_X1    g01240(.A1(new_n1432_), .A2(new_n1282_), .Z(new_n1433_));
  INV_X1     g01241(.I(new_n1433_), .ZN(new_n1434_));
  NOR2_X1    g01242(.A1(new_n1350_), .A2(new_n1345_), .ZN(new_n1435_));
  NOR2_X1    g01243(.A1(\asqrt[50] ), .A2(new_n1435_), .ZN(new_n1436_));
  XOR2_X1    g01244(.A1(new_n1436_), .A2(new_n1284_), .Z(new_n1437_));
  NOR2_X1    g01245(.A1(new_n1373_), .A2(new_n1344_), .ZN(new_n1438_));
  NOR2_X1    g01246(.A1(\asqrt[50] ), .A2(new_n1438_), .ZN(new_n1439_));
  XOR2_X1    g01247(.A1(new_n1439_), .A2(new_n1288_), .Z(new_n1440_));
  AOI21_X1   g01248(.A1(new_n1338_), .A2(new_n1343_), .B(\asqrt[50] ), .ZN(new_n1441_));
  XOR2_X1    g01249(.A1(new_n1441_), .A2(new_n1291_), .Z(new_n1442_));
  INV_X1     g01250(.I(new_n1442_), .ZN(new_n1443_));
  AOI21_X1   g01251(.A1(new_n1369_), .A2(new_n1337_), .B(\asqrt[50] ), .ZN(new_n1444_));
  XOR2_X1    g01252(.A1(new_n1444_), .A2(new_n1310_), .Z(new_n1445_));
  INV_X1     g01253(.I(new_n1445_), .ZN(new_n1446_));
  AOI21_X1   g01254(.A1(new_n1367_), .A2(new_n1334_), .B(\asqrt[50] ), .ZN(new_n1447_));
  XOR2_X1    g01255(.A1(new_n1447_), .A2(new_n1358_), .Z(new_n1448_));
  NOR2_X1    g01256(.A1(new_n1305_), .A2(\a[102] ), .ZN(new_n1449_));
  INV_X1     g01257(.I(new_n1449_), .ZN(new_n1450_));
  NOR2_X1    g01258(.A1(new_n1326_), .A2(\a[102] ), .ZN(new_n1451_));
  AOI22_X1   g01259(.A1(new_n1450_), .A2(new_n1326_), .B1(\asqrt[51] ), .B2(new_n1451_), .ZN(new_n1452_));
  INV_X1     g01260(.I(new_n1452_), .ZN(new_n1453_));
  INV_X1     g01261(.I(new_n1390_), .ZN(new_n1454_));
  NOR2_X1    g01262(.A1(new_n1404_), .A2(new_n1400_), .ZN(new_n1455_));
  AOI21_X1   g01263(.A1(new_n1397_), .A2(new_n1394_), .B(\asqrt[62] ), .ZN(new_n1456_));
  NOR3_X1    g01264(.A1(new_n1404_), .A2(new_n201_), .A3(new_n1400_), .ZN(new_n1457_));
  OAI22_X1   g01265(.A1(new_n1456_), .A2(new_n1457_), .B1(new_n1455_), .B2(new_n1409_), .ZN(new_n1458_));
  AOI21_X1   g01266(.A1(new_n1458_), .A2(new_n1454_), .B(new_n1413_), .ZN(new_n1459_));
  AOI21_X1   g01267(.A1(new_n1455_), .A2(new_n201_), .B(new_n1410_), .ZN(new_n1460_));
  NOR2_X1    g01268(.A1(new_n1455_), .A2(new_n201_), .ZN(new_n1461_));
  NOR3_X1    g01269(.A1(new_n1460_), .A2(new_n1461_), .A3(new_n1454_), .ZN(new_n1462_));
  NOR4_X1    g01270(.A1(new_n1459_), .A2(\asqrt[63] ), .A3(new_n1462_), .A4(new_n1424_), .ZN(new_n1463_));
  NOR2_X1    g01271(.A1(new_n1324_), .A2(new_n1365_), .ZN(new_n1464_));
  NOR2_X1    g01272(.A1(new_n1463_), .A2(new_n1464_), .ZN(new_n1465_));
  NOR2_X1    g01273(.A1(new_n1465_), .A2(new_n1453_), .ZN(new_n1466_));
  NOR3_X1    g01274(.A1(new_n1463_), .A2(new_n1452_), .A3(new_n1464_), .ZN(new_n1467_));
  NOR2_X1    g01275(.A1(new_n1466_), .A2(new_n1467_), .ZN(new_n1468_));
  NOR3_X1    g01276(.A1(new_n1459_), .A2(\asqrt[63] ), .A3(new_n1462_), .ZN(new_n1469_));
  NAND4_X1   g01277(.A1(new_n1469_), .A2(\asqrt[51] ), .A3(new_n1421_), .A4(new_n1423_), .ZN(new_n1470_));
  NAND2_X1   g01278(.A1(\asqrt[50] ), .A2(new_n1319_), .ZN(new_n1471_));
  AOI21_X1   g01279(.A1(new_n1470_), .A2(new_n1471_), .B(\a[102] ), .ZN(new_n1472_));
  NAND2_X1   g01280(.A1(new_n1415_), .A2(new_n193_), .ZN(new_n1473_));
  NAND3_X1   g01281(.A1(new_n1421_), .A2(\asqrt[51] ), .A3(new_n1423_), .ZN(new_n1474_));
  NOR3_X1    g01282(.A1(new_n1473_), .A2(new_n1462_), .A3(new_n1474_), .ZN(new_n1475_));
  NOR2_X1    g01283(.A1(new_n1463_), .A2(new_n1320_), .ZN(new_n1476_));
  NOR3_X1    g01284(.A1(new_n1476_), .A2(new_n1475_), .A3(new_n1322_), .ZN(new_n1477_));
  OR2_X2     g01285(.A1(new_n1472_), .A2(new_n1477_), .Z(new_n1478_));
  NOR2_X1    g01286(.A1(\a[98] ), .A2(\a[99] ), .ZN(new_n1479_));
  INV_X1     g01287(.I(new_n1479_), .ZN(new_n1480_));
  NAND3_X1   g01288(.A1(\asqrt[50] ), .A2(\a[100] ), .A3(new_n1480_), .ZN(new_n1481_));
  INV_X1     g01289(.I(\a[100] ), .ZN(new_n1482_));
  OAI21_X1   g01290(.A1(\asqrt[50] ), .A2(new_n1482_), .B(new_n1479_), .ZN(new_n1483_));
  AOI21_X1   g01291(.A1(new_n1483_), .A2(new_n1481_), .B(new_n1305_), .ZN(new_n1484_));
  NOR3_X1    g01292(.A1(new_n1301_), .A2(\asqrt[63] ), .A3(new_n1304_), .ZN(new_n1485_));
  NAND2_X1   g01293(.A1(new_n1479_), .A2(new_n1482_), .ZN(new_n1486_));
  NAND3_X1   g01294(.A1(new_n1270_), .A2(new_n1272_), .A3(new_n1486_), .ZN(new_n1487_));
  NAND2_X1   g01295(.A1(new_n1485_), .A2(new_n1487_), .ZN(new_n1488_));
  NAND3_X1   g01296(.A1(\asqrt[50] ), .A2(\a[100] ), .A3(new_n1488_), .ZN(new_n1489_));
  INV_X1     g01297(.I(\a[101] ), .ZN(new_n1490_));
  NAND3_X1   g01298(.A1(\asqrt[50] ), .A2(new_n1482_), .A3(new_n1490_), .ZN(new_n1491_));
  OAI21_X1   g01299(.A1(new_n1463_), .A2(\a[100] ), .B(\a[101] ), .ZN(new_n1492_));
  NAND3_X1   g01300(.A1(new_n1489_), .A2(new_n1492_), .A3(new_n1491_), .ZN(new_n1493_));
  NOR3_X1    g01301(.A1(new_n1493_), .A2(new_n1484_), .A3(\asqrt[52] ), .ZN(new_n1494_));
  OAI21_X1   g01302(.A1(new_n1493_), .A2(new_n1484_), .B(\asqrt[52] ), .ZN(new_n1495_));
  OAI21_X1   g01303(.A1(new_n1478_), .A2(new_n1494_), .B(new_n1495_), .ZN(new_n1496_));
  OAI21_X1   g01304(.A1(new_n1496_), .A2(\asqrt[53] ), .B(new_n1468_), .ZN(new_n1497_));
  NAND2_X1   g01305(.A1(new_n1496_), .A2(\asqrt[53] ), .ZN(new_n1498_));
  NAND3_X1   g01306(.A1(new_n1497_), .A2(new_n1498_), .A3(new_n860_), .ZN(new_n1499_));
  AOI21_X1   g01307(.A1(new_n1497_), .A2(new_n1498_), .B(new_n860_), .ZN(new_n1500_));
  AOI21_X1   g01308(.A1(new_n1448_), .A2(new_n1499_), .B(new_n1500_), .ZN(new_n1501_));
  AOI21_X1   g01309(.A1(new_n1501_), .A2(new_n744_), .B(new_n1446_), .ZN(new_n1502_));
  NAND2_X1   g01310(.A1(new_n1499_), .A2(new_n1448_), .ZN(new_n1503_));
  INV_X1     g01311(.I(new_n1468_), .ZN(new_n1504_));
  NOR2_X1    g01312(.A1(new_n1472_), .A2(new_n1477_), .ZN(new_n1505_));
  NOR3_X1    g01313(.A1(new_n1463_), .A2(new_n1482_), .A3(new_n1479_), .ZN(new_n1506_));
  AOI21_X1   g01314(.A1(new_n1463_), .A2(\a[100] ), .B(new_n1480_), .ZN(new_n1507_));
  OAI21_X1   g01315(.A1(new_n1506_), .A2(new_n1507_), .B(\asqrt[51] ), .ZN(new_n1508_));
  INV_X1     g01316(.I(new_n1488_), .ZN(new_n1509_));
  NOR3_X1    g01317(.A1(new_n1463_), .A2(new_n1482_), .A3(new_n1509_), .ZN(new_n1510_));
  NOR3_X1    g01318(.A1(new_n1463_), .A2(\a[100] ), .A3(\a[101] ), .ZN(new_n1511_));
  AOI21_X1   g01319(.A1(\asqrt[50] ), .A2(new_n1482_), .B(new_n1490_), .ZN(new_n1512_));
  NOR3_X1    g01320(.A1(new_n1510_), .A2(new_n1511_), .A3(new_n1512_), .ZN(new_n1513_));
  NAND3_X1   g01321(.A1(new_n1513_), .A2(new_n1508_), .A3(new_n1150_), .ZN(new_n1514_));
  AOI21_X1   g01322(.A1(new_n1513_), .A2(new_n1508_), .B(new_n1150_), .ZN(new_n1515_));
  AOI21_X1   g01323(.A1(new_n1505_), .A2(new_n1514_), .B(new_n1515_), .ZN(new_n1516_));
  AOI21_X1   g01324(.A1(new_n1516_), .A2(new_n1006_), .B(new_n1504_), .ZN(new_n1517_));
  NAND2_X1   g01325(.A1(new_n1514_), .A2(new_n1505_), .ZN(new_n1518_));
  AOI21_X1   g01326(.A1(new_n1518_), .A2(new_n1495_), .B(new_n1006_), .ZN(new_n1519_));
  OAI21_X1   g01327(.A1(new_n1517_), .A2(new_n1519_), .B(\asqrt[54] ), .ZN(new_n1520_));
  AOI21_X1   g01328(.A1(new_n1503_), .A2(new_n1520_), .B(new_n744_), .ZN(new_n1521_));
  NOR3_X1    g01329(.A1(new_n1502_), .A2(\asqrt[56] ), .A3(new_n1521_), .ZN(new_n1522_));
  OAI21_X1   g01330(.A1(new_n1502_), .A2(new_n1521_), .B(\asqrt[56] ), .ZN(new_n1523_));
  OAI21_X1   g01331(.A1(new_n1443_), .A2(new_n1522_), .B(new_n1523_), .ZN(new_n1524_));
  OAI21_X1   g01332(.A1(new_n1524_), .A2(\asqrt[57] ), .B(new_n1440_), .ZN(new_n1525_));
  NAND2_X1   g01333(.A1(new_n1524_), .A2(\asqrt[57] ), .ZN(new_n1526_));
  NAND3_X1   g01334(.A1(new_n1525_), .A2(new_n1526_), .A3(new_n423_), .ZN(new_n1527_));
  AOI21_X1   g01335(.A1(new_n1525_), .A2(new_n1526_), .B(new_n423_), .ZN(new_n1528_));
  AOI21_X1   g01336(.A1(new_n1437_), .A2(new_n1527_), .B(new_n1528_), .ZN(new_n1529_));
  AOI21_X1   g01337(.A1(new_n1529_), .A2(new_n337_), .B(new_n1434_), .ZN(new_n1530_));
  NAND2_X1   g01338(.A1(new_n1527_), .A2(new_n1437_), .ZN(new_n1531_));
  INV_X1     g01339(.I(new_n1440_), .ZN(new_n1532_));
  INV_X1     g01340(.I(new_n1448_), .ZN(new_n1533_));
  NOR3_X1    g01341(.A1(new_n1517_), .A2(\asqrt[54] ), .A3(new_n1519_), .ZN(new_n1534_));
  OAI21_X1   g01342(.A1(new_n1533_), .A2(new_n1534_), .B(new_n1520_), .ZN(new_n1535_));
  OAI21_X1   g01343(.A1(new_n1535_), .A2(\asqrt[55] ), .B(new_n1445_), .ZN(new_n1536_));
  NAND2_X1   g01344(.A1(new_n1535_), .A2(\asqrt[55] ), .ZN(new_n1537_));
  NAND3_X1   g01345(.A1(new_n1536_), .A2(new_n1537_), .A3(new_n634_), .ZN(new_n1538_));
  AOI21_X1   g01346(.A1(new_n1536_), .A2(new_n1537_), .B(new_n634_), .ZN(new_n1539_));
  AOI21_X1   g01347(.A1(new_n1442_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n1540_));
  AOI21_X1   g01348(.A1(new_n1540_), .A2(new_n531_), .B(new_n1532_), .ZN(new_n1541_));
  NAND2_X1   g01349(.A1(new_n1538_), .A2(new_n1442_), .ZN(new_n1542_));
  AOI21_X1   g01350(.A1(new_n1542_), .A2(new_n1523_), .B(new_n531_), .ZN(new_n1543_));
  OAI21_X1   g01351(.A1(new_n1541_), .A2(new_n1543_), .B(\asqrt[58] ), .ZN(new_n1544_));
  AOI21_X1   g01352(.A1(new_n1531_), .A2(new_n1544_), .B(new_n337_), .ZN(new_n1545_));
  NOR3_X1    g01353(.A1(new_n1530_), .A2(\asqrt[60] ), .A3(new_n1545_), .ZN(new_n1546_));
  NOR2_X1    g01354(.A1(new_n1546_), .A2(new_n1431_), .ZN(new_n1547_));
  INV_X1     g01355(.I(new_n1437_), .ZN(new_n1548_));
  NOR3_X1    g01356(.A1(new_n1541_), .A2(\asqrt[58] ), .A3(new_n1543_), .ZN(new_n1549_));
  OAI21_X1   g01357(.A1(new_n1548_), .A2(new_n1549_), .B(new_n1544_), .ZN(new_n1550_));
  OAI21_X1   g01358(.A1(new_n1550_), .A2(\asqrt[59] ), .B(new_n1433_), .ZN(new_n1551_));
  NOR2_X1    g01359(.A1(new_n1549_), .A2(new_n1548_), .ZN(new_n1552_));
  OAI21_X1   g01360(.A1(new_n1552_), .A2(new_n1528_), .B(\asqrt[59] ), .ZN(new_n1553_));
  AOI21_X1   g01361(.A1(new_n1551_), .A2(new_n1553_), .B(new_n266_), .ZN(new_n1554_));
  OAI21_X1   g01362(.A1(new_n1547_), .A2(new_n1554_), .B(\asqrt[61] ), .ZN(new_n1555_));
  NAND3_X1   g01363(.A1(new_n1551_), .A2(new_n266_), .A3(new_n1553_), .ZN(new_n1556_));
  NAND2_X1   g01364(.A1(new_n1556_), .A2(new_n1430_), .ZN(new_n1557_));
  OAI21_X1   g01365(.A1(new_n1530_), .A2(new_n1545_), .B(\asqrt[60] ), .ZN(new_n1558_));
  NAND3_X1   g01366(.A1(new_n1557_), .A2(new_n239_), .A3(new_n1558_), .ZN(new_n1559_));
  NOR2_X1    g01367(.A1(new_n1398_), .A2(\asqrt[62] ), .ZN(new_n1560_));
  NOR2_X1    g01368(.A1(new_n1560_), .A2(new_n1461_), .ZN(new_n1561_));
  XOR2_X1    g01369(.A1(new_n1408_), .A2(new_n1238_), .Z(new_n1562_));
  OAI21_X1   g01370(.A1(\asqrt[50] ), .A2(new_n1561_), .B(new_n1562_), .ZN(new_n1563_));
  INV_X1     g01371(.I(new_n1563_), .ZN(new_n1564_));
  OAI21_X1   g01372(.A1(new_n1431_), .A2(new_n1546_), .B(new_n1558_), .ZN(new_n1565_));
  OAI21_X1   g01373(.A1(new_n1565_), .A2(\asqrt[61] ), .B(new_n1428_), .ZN(new_n1566_));
  NAND2_X1   g01374(.A1(new_n1566_), .A2(new_n1555_), .ZN(new_n1567_));
  AOI21_X1   g01375(.A1(new_n1557_), .A2(new_n1558_), .B(new_n239_), .ZN(new_n1568_));
  INV_X1     g01376(.I(new_n1428_), .ZN(new_n1569_));
  AOI21_X1   g01377(.A1(new_n1430_), .A2(new_n1556_), .B(new_n1554_), .ZN(new_n1570_));
  AOI21_X1   g01378(.A1(new_n1570_), .A2(new_n239_), .B(new_n1569_), .ZN(new_n1571_));
  OAI21_X1   g01379(.A1(new_n1571_), .A2(new_n1568_), .B(new_n201_), .ZN(new_n1572_));
  NAND3_X1   g01380(.A1(new_n1566_), .A2(\asqrt[62] ), .A3(new_n1555_), .ZN(new_n1573_));
  NAND2_X1   g01381(.A1(new_n1402_), .A2(new_n239_), .ZN(new_n1574_));
  AOI21_X1   g01382(.A1(new_n1394_), .A2(new_n1574_), .B(\asqrt[50] ), .ZN(new_n1575_));
  XOR2_X1    g01383(.A1(new_n1575_), .A2(new_n1396_), .Z(new_n1576_));
  INV_X1     g01384(.I(new_n1576_), .ZN(new_n1577_));
  AOI22_X1   g01385(.A1(new_n1572_), .A2(new_n1573_), .B1(new_n1567_), .B2(new_n1577_), .ZN(new_n1578_));
  NOR2_X1    g01386(.A1(new_n1411_), .A2(new_n1390_), .ZN(new_n1579_));
  OAI21_X1   g01387(.A1(\asqrt[50] ), .A2(new_n1579_), .B(new_n1418_), .ZN(new_n1580_));
  INV_X1     g01388(.I(new_n1580_), .ZN(new_n1581_));
  OAI21_X1   g01389(.A1(new_n1578_), .A2(new_n1564_), .B(new_n1581_), .ZN(new_n1582_));
  OAI21_X1   g01390(.A1(new_n1567_), .A2(\asqrt[62] ), .B(new_n1576_), .ZN(new_n1583_));
  NAND2_X1   g01391(.A1(new_n1567_), .A2(\asqrt[62] ), .ZN(new_n1584_));
  NAND3_X1   g01392(.A1(new_n1583_), .A2(new_n1584_), .A3(new_n1564_), .ZN(new_n1585_));
  NAND2_X1   g01393(.A1(new_n1463_), .A2(new_n1454_), .ZN(new_n1586_));
  XOR2_X1    g01394(.A1(new_n1458_), .A2(new_n1454_), .Z(new_n1587_));
  NAND3_X1   g01395(.A1(new_n1586_), .A2(\asqrt[63] ), .A3(new_n1587_), .ZN(new_n1588_));
  INV_X1     g01396(.I(new_n1473_), .ZN(new_n1589_));
  NAND4_X1   g01397(.A1(new_n1589_), .A2(new_n1390_), .A3(new_n1418_), .A4(new_n1425_), .ZN(new_n1590_));
  NAND2_X1   g01398(.A1(new_n1588_), .A2(new_n1590_), .ZN(new_n1591_));
  INV_X1     g01399(.I(new_n1591_), .ZN(new_n1592_));
  NAND4_X1   g01400(.A1(new_n1582_), .A2(new_n193_), .A3(new_n1585_), .A4(new_n1592_), .ZN(\asqrt[49] ));
  AOI21_X1   g01401(.A1(new_n1555_), .A2(new_n1559_), .B(\asqrt[49] ), .ZN(new_n1594_));
  XOR2_X1    g01402(.A1(new_n1594_), .A2(new_n1428_), .Z(new_n1595_));
  INV_X1     g01403(.I(new_n1595_), .ZN(new_n1596_));
  NAND2_X1   g01404(.A1(new_n1529_), .A2(new_n337_), .ZN(new_n1597_));
  AOI21_X1   g01405(.A1(new_n1597_), .A2(new_n1553_), .B(\asqrt[49] ), .ZN(new_n1598_));
  XOR2_X1    g01406(.A1(new_n1598_), .A2(new_n1433_), .Z(new_n1599_));
  AOI21_X1   g01407(.A1(new_n1527_), .A2(new_n1544_), .B(\asqrt[49] ), .ZN(new_n1600_));
  XOR2_X1    g01408(.A1(new_n1600_), .A2(new_n1437_), .Z(new_n1601_));
  INV_X1     g01409(.I(new_n1601_), .ZN(new_n1602_));
  NAND2_X1   g01410(.A1(new_n1540_), .A2(new_n531_), .ZN(new_n1603_));
  AOI21_X1   g01411(.A1(new_n1603_), .A2(new_n1526_), .B(\asqrt[49] ), .ZN(new_n1604_));
  XOR2_X1    g01412(.A1(new_n1604_), .A2(new_n1440_), .Z(new_n1605_));
  INV_X1     g01413(.I(new_n1605_), .ZN(new_n1606_));
  AOI21_X1   g01414(.A1(new_n1538_), .A2(new_n1523_), .B(\asqrt[49] ), .ZN(new_n1607_));
  XOR2_X1    g01415(.A1(new_n1607_), .A2(new_n1442_), .Z(new_n1608_));
  NAND2_X1   g01416(.A1(new_n1501_), .A2(new_n744_), .ZN(new_n1609_));
  AOI21_X1   g01417(.A1(new_n1609_), .A2(new_n1537_), .B(\asqrt[49] ), .ZN(new_n1610_));
  XOR2_X1    g01418(.A1(new_n1610_), .A2(new_n1445_), .Z(new_n1611_));
  AOI21_X1   g01419(.A1(new_n1499_), .A2(new_n1520_), .B(\asqrt[49] ), .ZN(new_n1612_));
  XOR2_X1    g01420(.A1(new_n1612_), .A2(new_n1448_), .Z(new_n1613_));
  INV_X1     g01421(.I(new_n1613_), .ZN(new_n1614_));
  NAND2_X1   g01422(.A1(new_n1516_), .A2(new_n1006_), .ZN(new_n1615_));
  AOI21_X1   g01423(.A1(new_n1615_), .A2(new_n1498_), .B(\asqrt[49] ), .ZN(new_n1616_));
  XOR2_X1    g01424(.A1(new_n1616_), .A2(new_n1468_), .Z(new_n1617_));
  INV_X1     g01425(.I(new_n1617_), .ZN(new_n1618_));
  AOI21_X1   g01426(.A1(new_n1514_), .A2(new_n1495_), .B(\asqrt[49] ), .ZN(new_n1619_));
  XOR2_X1    g01427(.A1(new_n1619_), .A2(new_n1505_), .Z(new_n1620_));
  NAND2_X1   g01428(.A1(\asqrt[50] ), .A2(new_n1482_), .ZN(new_n1621_));
  NOR2_X1    g01429(.A1(new_n1490_), .A2(\a[100] ), .ZN(new_n1622_));
  AOI22_X1   g01430(.A1(new_n1621_), .A2(new_n1490_), .B1(\asqrt[50] ), .B2(new_n1622_), .ZN(new_n1623_));
  AOI21_X1   g01431(.A1(new_n1428_), .A2(new_n1559_), .B(new_n1568_), .ZN(new_n1624_));
  AOI21_X1   g01432(.A1(new_n1566_), .A2(new_n1555_), .B(\asqrt[62] ), .ZN(new_n1625_));
  NOR3_X1    g01433(.A1(new_n1571_), .A2(new_n201_), .A3(new_n1568_), .ZN(new_n1626_));
  OAI22_X1   g01434(.A1(new_n1626_), .A2(new_n1625_), .B1(new_n1624_), .B2(new_n1576_), .ZN(new_n1627_));
  AOI21_X1   g01435(.A1(new_n1627_), .A2(new_n1563_), .B(new_n1580_), .ZN(new_n1628_));
  AOI21_X1   g01436(.A1(new_n1624_), .A2(new_n201_), .B(new_n1577_), .ZN(new_n1629_));
  OAI21_X1   g01437(.A1(new_n1624_), .A2(new_n201_), .B(new_n1564_), .ZN(new_n1630_));
  NOR2_X1    g01438(.A1(new_n1629_), .A2(new_n1630_), .ZN(new_n1631_));
  NOR4_X1    g01439(.A1(new_n1628_), .A2(\asqrt[63] ), .A3(new_n1631_), .A4(new_n1591_), .ZN(new_n1632_));
  AOI21_X1   g01440(.A1(\asqrt[50] ), .A2(\a[100] ), .B(new_n1488_), .ZN(new_n1633_));
  OAI21_X1   g01441(.A1(new_n1484_), .A2(new_n1633_), .B(new_n1632_), .ZN(new_n1634_));
  XNOR2_X1   g01442(.A1(new_n1634_), .A2(new_n1623_), .ZN(new_n1635_));
  NOR3_X1    g01443(.A1(new_n1628_), .A2(\asqrt[63] ), .A3(new_n1631_), .ZN(new_n1636_));
  NAND3_X1   g01444(.A1(new_n1588_), .A2(\asqrt[50] ), .A3(new_n1590_), .ZN(new_n1637_));
  INV_X1     g01445(.I(new_n1637_), .ZN(new_n1638_));
  NAND2_X1   g01446(.A1(new_n1636_), .A2(new_n1638_), .ZN(new_n1639_));
  NAND2_X1   g01447(.A1(\asqrt[49] ), .A2(new_n1479_), .ZN(new_n1640_));
  AOI21_X1   g01448(.A1(new_n1640_), .A2(new_n1639_), .B(\a[100] ), .ZN(new_n1641_));
  NAND2_X1   g01449(.A1(new_n1582_), .A2(new_n193_), .ZN(new_n1642_));
  NOR3_X1    g01450(.A1(new_n1642_), .A2(new_n1631_), .A3(new_n1637_), .ZN(new_n1643_));
  NOR2_X1    g01451(.A1(new_n1632_), .A2(new_n1480_), .ZN(new_n1644_));
  NOR3_X1    g01452(.A1(new_n1644_), .A2(new_n1643_), .A3(new_n1482_), .ZN(new_n1645_));
  OR2_X2     g01453(.A1(new_n1645_), .A2(new_n1641_), .Z(new_n1646_));
  NOR2_X1    g01454(.A1(\a[96] ), .A2(\a[97] ), .ZN(new_n1647_));
  INV_X1     g01455(.I(new_n1647_), .ZN(new_n1648_));
  NAND3_X1   g01456(.A1(\asqrt[49] ), .A2(\a[98] ), .A3(new_n1648_), .ZN(new_n1649_));
  INV_X1     g01457(.I(\a[98] ), .ZN(new_n1650_));
  OAI21_X1   g01458(.A1(\asqrt[49] ), .A2(new_n1650_), .B(new_n1647_), .ZN(new_n1651_));
  AOI21_X1   g01459(.A1(new_n1651_), .A2(new_n1649_), .B(new_n1463_), .ZN(new_n1652_));
  NAND2_X1   g01460(.A1(new_n1647_), .A2(new_n1650_), .ZN(new_n1653_));
  NAND3_X1   g01461(.A1(new_n1421_), .A2(new_n1423_), .A3(new_n1653_), .ZN(new_n1654_));
  NAND2_X1   g01462(.A1(new_n1469_), .A2(new_n1654_), .ZN(new_n1655_));
  NAND3_X1   g01463(.A1(\asqrt[49] ), .A2(\a[98] ), .A3(new_n1655_), .ZN(new_n1656_));
  INV_X1     g01464(.I(\a[99] ), .ZN(new_n1657_));
  NAND3_X1   g01465(.A1(\asqrt[49] ), .A2(new_n1650_), .A3(new_n1657_), .ZN(new_n1658_));
  OAI21_X1   g01466(.A1(new_n1632_), .A2(\a[98] ), .B(\a[99] ), .ZN(new_n1659_));
  NAND3_X1   g01467(.A1(new_n1656_), .A2(new_n1659_), .A3(new_n1658_), .ZN(new_n1660_));
  NOR3_X1    g01468(.A1(new_n1660_), .A2(new_n1652_), .A3(\asqrt[51] ), .ZN(new_n1661_));
  OAI21_X1   g01469(.A1(new_n1660_), .A2(new_n1652_), .B(\asqrt[51] ), .ZN(new_n1662_));
  OAI21_X1   g01470(.A1(new_n1646_), .A2(new_n1661_), .B(new_n1662_), .ZN(new_n1663_));
  OAI21_X1   g01471(.A1(new_n1663_), .A2(\asqrt[52] ), .B(new_n1635_), .ZN(new_n1664_));
  NAND2_X1   g01472(.A1(new_n1663_), .A2(\asqrt[52] ), .ZN(new_n1665_));
  NAND3_X1   g01473(.A1(new_n1664_), .A2(new_n1665_), .A3(new_n1006_), .ZN(new_n1666_));
  AOI21_X1   g01474(.A1(new_n1664_), .A2(new_n1665_), .B(new_n1006_), .ZN(new_n1667_));
  AOI21_X1   g01475(.A1(new_n1620_), .A2(new_n1666_), .B(new_n1667_), .ZN(new_n1668_));
  AOI21_X1   g01476(.A1(new_n1668_), .A2(new_n860_), .B(new_n1618_), .ZN(new_n1669_));
  NAND2_X1   g01477(.A1(new_n1666_), .A2(new_n1620_), .ZN(new_n1670_));
  INV_X1     g01478(.I(new_n1667_), .ZN(new_n1671_));
  AOI21_X1   g01479(.A1(new_n1670_), .A2(new_n1671_), .B(new_n860_), .ZN(new_n1672_));
  NOR3_X1    g01480(.A1(new_n1669_), .A2(\asqrt[55] ), .A3(new_n1672_), .ZN(new_n1673_));
  OAI21_X1   g01481(.A1(new_n1669_), .A2(new_n1672_), .B(\asqrt[55] ), .ZN(new_n1674_));
  OAI21_X1   g01482(.A1(new_n1614_), .A2(new_n1673_), .B(new_n1674_), .ZN(new_n1675_));
  OAI21_X1   g01483(.A1(new_n1675_), .A2(\asqrt[56] ), .B(new_n1611_), .ZN(new_n1676_));
  NAND2_X1   g01484(.A1(new_n1675_), .A2(\asqrt[56] ), .ZN(new_n1677_));
  NAND3_X1   g01485(.A1(new_n1676_), .A2(new_n1677_), .A3(new_n531_), .ZN(new_n1678_));
  AOI21_X1   g01486(.A1(new_n1676_), .A2(new_n1677_), .B(new_n531_), .ZN(new_n1679_));
  AOI21_X1   g01487(.A1(new_n1608_), .A2(new_n1678_), .B(new_n1679_), .ZN(new_n1680_));
  AOI21_X1   g01488(.A1(new_n1680_), .A2(new_n423_), .B(new_n1606_), .ZN(new_n1681_));
  NAND2_X1   g01489(.A1(new_n1678_), .A2(new_n1608_), .ZN(new_n1682_));
  INV_X1     g01490(.I(new_n1611_), .ZN(new_n1683_));
  NOR2_X1    g01491(.A1(new_n1673_), .A2(new_n1614_), .ZN(new_n1684_));
  INV_X1     g01492(.I(new_n1674_), .ZN(new_n1685_));
  NOR2_X1    g01493(.A1(new_n1684_), .A2(new_n1685_), .ZN(new_n1686_));
  AOI21_X1   g01494(.A1(new_n1686_), .A2(new_n634_), .B(new_n1683_), .ZN(new_n1687_));
  INV_X1     g01495(.I(new_n1620_), .ZN(new_n1688_));
  NOR2_X1    g01496(.A1(new_n1645_), .A2(new_n1641_), .ZN(new_n1689_));
  NOR3_X1    g01497(.A1(new_n1632_), .A2(new_n1650_), .A3(new_n1647_), .ZN(new_n1690_));
  AOI21_X1   g01498(.A1(new_n1632_), .A2(\a[98] ), .B(new_n1648_), .ZN(new_n1691_));
  OAI21_X1   g01499(.A1(new_n1690_), .A2(new_n1691_), .B(\asqrt[50] ), .ZN(new_n1692_));
  INV_X1     g01500(.I(new_n1655_), .ZN(new_n1693_));
  NOR3_X1    g01501(.A1(new_n1632_), .A2(new_n1650_), .A3(new_n1693_), .ZN(new_n1694_));
  NOR3_X1    g01502(.A1(new_n1632_), .A2(\a[98] ), .A3(\a[99] ), .ZN(new_n1695_));
  AOI21_X1   g01503(.A1(\asqrt[49] ), .A2(new_n1650_), .B(new_n1657_), .ZN(new_n1696_));
  NOR3_X1    g01504(.A1(new_n1694_), .A2(new_n1695_), .A3(new_n1696_), .ZN(new_n1697_));
  NAND3_X1   g01505(.A1(new_n1697_), .A2(new_n1692_), .A3(new_n1305_), .ZN(new_n1698_));
  NAND2_X1   g01506(.A1(new_n1698_), .A2(new_n1689_), .ZN(new_n1699_));
  NAND3_X1   g01507(.A1(new_n1699_), .A2(new_n1150_), .A3(new_n1662_), .ZN(new_n1700_));
  AOI21_X1   g01508(.A1(new_n1699_), .A2(new_n1662_), .B(new_n1150_), .ZN(new_n1701_));
  AOI21_X1   g01509(.A1(new_n1635_), .A2(new_n1700_), .B(new_n1701_), .ZN(new_n1702_));
  AOI21_X1   g01510(.A1(new_n1702_), .A2(new_n1006_), .B(new_n1688_), .ZN(new_n1703_));
  NOR3_X1    g01511(.A1(new_n1703_), .A2(\asqrt[54] ), .A3(new_n1667_), .ZN(new_n1704_));
  OAI21_X1   g01512(.A1(new_n1703_), .A2(new_n1667_), .B(\asqrt[54] ), .ZN(new_n1705_));
  OAI21_X1   g01513(.A1(new_n1618_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n1706_));
  OAI21_X1   g01514(.A1(new_n1706_), .A2(\asqrt[55] ), .B(new_n1613_), .ZN(new_n1707_));
  AOI21_X1   g01515(.A1(new_n1707_), .A2(new_n1674_), .B(new_n634_), .ZN(new_n1708_));
  OAI21_X1   g01516(.A1(new_n1687_), .A2(new_n1708_), .B(\asqrt[57] ), .ZN(new_n1709_));
  AOI21_X1   g01517(.A1(new_n1682_), .A2(new_n1709_), .B(new_n423_), .ZN(new_n1710_));
  NOR3_X1    g01518(.A1(new_n1681_), .A2(\asqrt[59] ), .A3(new_n1710_), .ZN(new_n1711_));
  OAI21_X1   g01519(.A1(new_n1681_), .A2(new_n1710_), .B(\asqrt[59] ), .ZN(new_n1712_));
  OAI21_X1   g01520(.A1(new_n1602_), .A2(new_n1711_), .B(new_n1712_), .ZN(new_n1713_));
  OAI21_X1   g01521(.A1(new_n1713_), .A2(\asqrt[60] ), .B(new_n1599_), .ZN(new_n1714_));
  NOR2_X1    g01522(.A1(new_n1711_), .A2(new_n1602_), .ZN(new_n1715_));
  NAND3_X1   g01523(.A1(new_n1682_), .A2(new_n423_), .A3(new_n1709_), .ZN(new_n1716_));
  NAND2_X1   g01524(.A1(new_n1716_), .A2(new_n1605_), .ZN(new_n1717_));
  INV_X1     g01525(.I(new_n1608_), .ZN(new_n1718_));
  NAND3_X1   g01526(.A1(new_n1707_), .A2(new_n634_), .A3(new_n1674_), .ZN(new_n1719_));
  AOI21_X1   g01527(.A1(new_n1611_), .A2(new_n1719_), .B(new_n1708_), .ZN(new_n1720_));
  AOI21_X1   g01528(.A1(new_n1720_), .A2(new_n531_), .B(new_n1718_), .ZN(new_n1721_));
  OAI21_X1   g01529(.A1(new_n1721_), .A2(new_n1679_), .B(\asqrt[58] ), .ZN(new_n1722_));
  AOI21_X1   g01530(.A1(new_n1717_), .A2(new_n1722_), .B(new_n337_), .ZN(new_n1723_));
  OAI21_X1   g01531(.A1(new_n1715_), .A2(new_n1723_), .B(\asqrt[60] ), .ZN(new_n1724_));
  AOI21_X1   g01532(.A1(new_n1714_), .A2(new_n1724_), .B(new_n239_), .ZN(new_n1725_));
  AOI21_X1   g01533(.A1(new_n1556_), .A2(new_n1558_), .B(\asqrt[49] ), .ZN(new_n1726_));
  XOR2_X1    g01534(.A1(new_n1726_), .A2(new_n1430_), .Z(new_n1727_));
  NAND3_X1   g01535(.A1(new_n1714_), .A2(new_n239_), .A3(new_n1724_), .ZN(new_n1728_));
  AOI21_X1   g01536(.A1(new_n1727_), .A2(new_n1728_), .B(new_n1725_), .ZN(new_n1729_));
  AOI21_X1   g01537(.A1(new_n1729_), .A2(new_n201_), .B(new_n1596_), .ZN(new_n1730_));
  NOR2_X1    g01538(.A1(new_n1567_), .A2(\asqrt[62] ), .ZN(new_n1731_));
  INV_X1     g01539(.I(new_n1584_), .ZN(new_n1732_));
  NOR2_X1    g01540(.A1(new_n1732_), .A2(new_n1731_), .ZN(new_n1733_));
  XOR2_X1    g01541(.A1(new_n1575_), .A2(new_n1396_), .Z(new_n1734_));
  OAI21_X1   g01542(.A1(\asqrt[49] ), .A2(new_n1733_), .B(new_n1734_), .ZN(new_n1735_));
  NOR2_X1    g01543(.A1(new_n1729_), .A2(new_n201_), .ZN(new_n1736_));
  OR3_X2     g01544(.A1(new_n1730_), .A2(new_n1735_), .A3(new_n1736_), .Z(new_n1737_));
  INV_X1     g01545(.I(new_n1735_), .ZN(new_n1738_));
  INV_X1     g01546(.I(new_n1599_), .ZN(new_n1739_));
  NAND3_X1   g01547(.A1(new_n1717_), .A2(new_n337_), .A3(new_n1722_), .ZN(new_n1740_));
  AOI21_X1   g01548(.A1(new_n1601_), .A2(new_n1740_), .B(new_n1723_), .ZN(new_n1741_));
  AOI21_X1   g01549(.A1(new_n1741_), .A2(new_n266_), .B(new_n1739_), .ZN(new_n1742_));
  NOR3_X1    g01550(.A1(new_n1721_), .A2(\asqrt[58] ), .A3(new_n1679_), .ZN(new_n1743_));
  OAI21_X1   g01551(.A1(new_n1606_), .A2(new_n1743_), .B(new_n1722_), .ZN(new_n1744_));
  OAI21_X1   g01552(.A1(new_n1744_), .A2(\asqrt[59] ), .B(new_n1601_), .ZN(new_n1745_));
  AOI21_X1   g01553(.A1(new_n1745_), .A2(new_n1712_), .B(new_n266_), .ZN(new_n1746_));
  OAI21_X1   g01554(.A1(new_n1742_), .A2(new_n1746_), .B(\asqrt[61] ), .ZN(new_n1747_));
  INV_X1     g01555(.I(new_n1727_), .ZN(new_n1748_));
  NOR3_X1    g01556(.A1(new_n1742_), .A2(\asqrt[61] ), .A3(new_n1746_), .ZN(new_n1749_));
  OAI21_X1   g01557(.A1(new_n1748_), .A2(new_n1749_), .B(new_n1747_), .ZN(new_n1750_));
  NAND3_X1   g01558(.A1(new_n1745_), .A2(new_n266_), .A3(new_n1712_), .ZN(new_n1751_));
  AOI21_X1   g01559(.A1(new_n1599_), .A2(new_n1751_), .B(new_n1746_), .ZN(new_n1752_));
  AOI21_X1   g01560(.A1(new_n1752_), .A2(new_n239_), .B(new_n1748_), .ZN(new_n1753_));
  OAI21_X1   g01561(.A1(new_n1753_), .A2(new_n1725_), .B(new_n201_), .ZN(new_n1754_));
  NAND2_X1   g01562(.A1(new_n1728_), .A2(new_n1727_), .ZN(new_n1755_));
  NAND3_X1   g01563(.A1(new_n1755_), .A2(\asqrt[62] ), .A3(new_n1747_), .ZN(new_n1756_));
  AOI22_X1   g01564(.A1(new_n1754_), .A2(new_n1756_), .B1(new_n1596_), .B2(new_n1750_), .ZN(new_n1757_));
  NOR2_X1    g01565(.A1(new_n1578_), .A2(new_n1564_), .ZN(new_n1758_));
  OAI21_X1   g01566(.A1(\asqrt[49] ), .A2(new_n1758_), .B(new_n1585_), .ZN(new_n1759_));
  INV_X1     g01567(.I(new_n1759_), .ZN(new_n1760_));
  OAI21_X1   g01568(.A1(new_n1757_), .A2(new_n1738_), .B(new_n1760_), .ZN(new_n1761_));
  NAND2_X1   g01569(.A1(new_n1632_), .A2(new_n1563_), .ZN(new_n1762_));
  XOR2_X1    g01570(.A1(new_n1578_), .A2(new_n1564_), .Z(new_n1763_));
  NAND3_X1   g01571(.A1(new_n1762_), .A2(\asqrt[63] ), .A3(new_n1763_), .ZN(new_n1764_));
  INV_X1     g01572(.I(new_n1642_), .ZN(new_n1765_));
  NAND4_X1   g01573(.A1(new_n1765_), .A2(new_n1564_), .A3(new_n1585_), .A4(new_n1592_), .ZN(new_n1766_));
  NAND2_X1   g01574(.A1(new_n1764_), .A2(new_n1766_), .ZN(new_n1767_));
  INV_X1     g01575(.I(new_n1767_), .ZN(new_n1768_));
  NAND4_X1   g01576(.A1(new_n1761_), .A2(new_n193_), .A3(new_n1737_), .A4(new_n1768_), .ZN(\asqrt[48] ));
  NAND2_X1   g01577(.A1(new_n1729_), .A2(new_n201_), .ZN(new_n1770_));
  INV_X1     g01578(.I(new_n1770_), .ZN(new_n1771_));
  NOR2_X1    g01579(.A1(new_n1771_), .A2(new_n1736_), .ZN(new_n1772_));
  NOR3_X1    g01580(.A1(new_n1730_), .A2(new_n1736_), .A3(new_n1735_), .ZN(new_n1773_));
  AOI21_X1   g01581(.A1(new_n1755_), .A2(new_n1747_), .B(\asqrt[62] ), .ZN(new_n1774_));
  NOR3_X1    g01582(.A1(new_n1753_), .A2(new_n201_), .A3(new_n1725_), .ZN(new_n1775_));
  OAI22_X1   g01583(.A1(new_n1775_), .A2(new_n1774_), .B1(new_n1595_), .B2(new_n1729_), .ZN(new_n1776_));
  AOI21_X1   g01584(.A1(new_n1776_), .A2(new_n1735_), .B(new_n1759_), .ZN(new_n1777_));
  NOR4_X1    g01585(.A1(new_n1777_), .A2(\asqrt[63] ), .A3(new_n1773_), .A4(new_n1767_), .ZN(new_n1778_));
  XOR2_X1    g01586(.A1(new_n1594_), .A2(new_n1428_), .Z(new_n1779_));
  OAI21_X1   g01587(.A1(\asqrt[48] ), .A2(new_n1772_), .B(new_n1779_), .ZN(new_n1780_));
  INV_X1     g01588(.I(new_n1780_), .ZN(new_n1781_));
  AOI21_X1   g01589(.A1(new_n1740_), .A2(new_n1712_), .B(\asqrt[48] ), .ZN(new_n1782_));
  XOR2_X1    g01590(.A1(new_n1782_), .A2(new_n1601_), .Z(new_n1783_));
  INV_X1     g01591(.I(new_n1783_), .ZN(new_n1784_));
  AOI21_X1   g01592(.A1(new_n1716_), .A2(new_n1722_), .B(\asqrt[48] ), .ZN(new_n1785_));
  XOR2_X1    g01593(.A1(new_n1785_), .A2(new_n1605_), .Z(new_n1786_));
  INV_X1     g01594(.I(new_n1786_), .ZN(new_n1787_));
  AOI21_X1   g01595(.A1(new_n1678_), .A2(new_n1709_), .B(\asqrt[48] ), .ZN(new_n1788_));
  XOR2_X1    g01596(.A1(new_n1788_), .A2(new_n1608_), .Z(new_n1789_));
  AOI21_X1   g01597(.A1(new_n1719_), .A2(new_n1677_), .B(\asqrt[48] ), .ZN(new_n1790_));
  XOR2_X1    g01598(.A1(new_n1790_), .A2(new_n1611_), .Z(new_n1791_));
  NOR2_X1    g01599(.A1(new_n1685_), .A2(new_n1673_), .ZN(new_n1792_));
  NOR2_X1    g01600(.A1(\asqrt[48] ), .A2(new_n1792_), .ZN(new_n1793_));
  XOR2_X1    g01601(.A1(new_n1793_), .A2(new_n1613_), .Z(new_n1794_));
  INV_X1     g01602(.I(new_n1794_), .ZN(new_n1795_));
  NOR2_X1    g01603(.A1(new_n1704_), .A2(new_n1672_), .ZN(new_n1796_));
  NOR2_X1    g01604(.A1(\asqrt[48] ), .A2(new_n1796_), .ZN(new_n1797_));
  XOR2_X1    g01605(.A1(new_n1797_), .A2(new_n1617_), .Z(new_n1798_));
  INV_X1     g01606(.I(new_n1798_), .ZN(new_n1799_));
  AOI21_X1   g01607(.A1(new_n1666_), .A2(new_n1671_), .B(\asqrt[48] ), .ZN(new_n1800_));
  XOR2_X1    g01608(.A1(new_n1800_), .A2(new_n1620_), .Z(new_n1801_));
  AOI21_X1   g01609(.A1(new_n1700_), .A2(new_n1665_), .B(\asqrt[48] ), .ZN(new_n1802_));
  XOR2_X1    g01610(.A1(new_n1802_), .A2(new_n1635_), .Z(new_n1803_));
  AOI21_X1   g01611(.A1(new_n1698_), .A2(new_n1662_), .B(\asqrt[48] ), .ZN(new_n1804_));
  XOR2_X1    g01612(.A1(new_n1804_), .A2(new_n1689_), .Z(new_n1805_));
  INV_X1     g01613(.I(new_n1805_), .ZN(new_n1806_));
  NAND2_X1   g01614(.A1(\asqrt[49] ), .A2(new_n1650_), .ZN(new_n1807_));
  NOR2_X1    g01615(.A1(new_n1657_), .A2(\a[98] ), .ZN(new_n1808_));
  AOI22_X1   g01616(.A1(new_n1807_), .A2(new_n1657_), .B1(\asqrt[49] ), .B2(new_n1808_), .ZN(new_n1809_));
  AOI21_X1   g01617(.A1(\asqrt[49] ), .A2(\a[98] ), .B(new_n1655_), .ZN(new_n1810_));
  OAI21_X1   g01618(.A1(new_n1652_), .A2(new_n1810_), .B(new_n1778_), .ZN(new_n1811_));
  XNOR2_X1   g01619(.A1(new_n1811_), .A2(new_n1809_), .ZN(new_n1812_));
  INV_X1     g01620(.I(new_n1812_), .ZN(new_n1813_));
  NAND2_X1   g01621(.A1(new_n1761_), .A2(new_n193_), .ZN(new_n1814_));
  NAND3_X1   g01622(.A1(new_n1764_), .A2(\asqrt[49] ), .A3(new_n1766_), .ZN(new_n1815_));
  NOR3_X1    g01623(.A1(new_n1814_), .A2(new_n1773_), .A3(new_n1815_), .ZN(new_n1816_));
  NOR2_X1    g01624(.A1(new_n1778_), .A2(new_n1648_), .ZN(new_n1817_));
  OAI21_X1   g01625(.A1(new_n1817_), .A2(new_n1816_), .B(new_n1650_), .ZN(new_n1818_));
  NOR3_X1    g01626(.A1(new_n1777_), .A2(\asqrt[63] ), .A3(new_n1773_), .ZN(new_n1819_));
  NAND4_X1   g01627(.A1(new_n1819_), .A2(\asqrt[49] ), .A3(new_n1764_), .A4(new_n1766_), .ZN(new_n1820_));
  NAND2_X1   g01628(.A1(\asqrt[48] ), .A2(new_n1647_), .ZN(new_n1821_));
  NAND3_X1   g01629(.A1(new_n1820_), .A2(new_n1821_), .A3(\a[98] ), .ZN(new_n1822_));
  NAND2_X1   g01630(.A1(new_n1822_), .A2(new_n1818_), .ZN(new_n1823_));
  INV_X1     g01631(.I(new_n1823_), .ZN(new_n1824_));
  INV_X1     g01632(.I(\a[96] ), .ZN(new_n1825_));
  NOR2_X1    g01633(.A1(\a[94] ), .A2(\a[95] ), .ZN(new_n1826_));
  NOR3_X1    g01634(.A1(new_n1778_), .A2(new_n1825_), .A3(new_n1826_), .ZN(new_n1827_));
  INV_X1     g01635(.I(new_n1826_), .ZN(new_n1828_));
  AOI21_X1   g01636(.A1(new_n1778_), .A2(\a[96] ), .B(new_n1828_), .ZN(new_n1829_));
  OAI21_X1   g01637(.A1(new_n1827_), .A2(new_n1829_), .B(\asqrt[49] ), .ZN(new_n1830_));
  NAND2_X1   g01638(.A1(new_n1826_), .A2(new_n1825_), .ZN(new_n1831_));
  NAND3_X1   g01639(.A1(new_n1588_), .A2(new_n1590_), .A3(new_n1831_), .ZN(new_n1832_));
  NAND2_X1   g01640(.A1(new_n1636_), .A2(new_n1832_), .ZN(new_n1833_));
  INV_X1     g01641(.I(new_n1833_), .ZN(new_n1834_));
  NOR3_X1    g01642(.A1(new_n1778_), .A2(new_n1825_), .A3(new_n1834_), .ZN(new_n1835_));
  NOR3_X1    g01643(.A1(new_n1778_), .A2(\a[96] ), .A3(\a[97] ), .ZN(new_n1836_));
  INV_X1     g01644(.I(\a[97] ), .ZN(new_n1837_));
  AOI21_X1   g01645(.A1(\asqrt[48] ), .A2(new_n1825_), .B(new_n1837_), .ZN(new_n1838_));
  NOR3_X1    g01646(.A1(new_n1835_), .A2(new_n1836_), .A3(new_n1838_), .ZN(new_n1839_));
  NAND3_X1   g01647(.A1(new_n1839_), .A2(new_n1830_), .A3(new_n1463_), .ZN(new_n1840_));
  AOI21_X1   g01648(.A1(new_n1839_), .A2(new_n1830_), .B(new_n1463_), .ZN(new_n1841_));
  AOI21_X1   g01649(.A1(new_n1824_), .A2(new_n1840_), .B(new_n1841_), .ZN(new_n1842_));
  AOI21_X1   g01650(.A1(new_n1842_), .A2(new_n1305_), .B(new_n1813_), .ZN(new_n1843_));
  NAND2_X1   g01651(.A1(new_n1824_), .A2(new_n1840_), .ZN(new_n1844_));
  NAND3_X1   g01652(.A1(\asqrt[48] ), .A2(\a[96] ), .A3(new_n1828_), .ZN(new_n1845_));
  OAI21_X1   g01653(.A1(\asqrt[48] ), .A2(new_n1825_), .B(new_n1826_), .ZN(new_n1846_));
  AOI21_X1   g01654(.A1(new_n1846_), .A2(new_n1845_), .B(new_n1632_), .ZN(new_n1847_));
  NAND3_X1   g01655(.A1(\asqrt[48] ), .A2(\a[96] ), .A3(new_n1833_), .ZN(new_n1848_));
  NAND3_X1   g01656(.A1(\asqrt[48] ), .A2(new_n1825_), .A3(new_n1837_), .ZN(new_n1849_));
  OAI21_X1   g01657(.A1(new_n1778_), .A2(\a[96] ), .B(\a[97] ), .ZN(new_n1850_));
  NAND3_X1   g01658(.A1(new_n1848_), .A2(new_n1850_), .A3(new_n1849_), .ZN(new_n1851_));
  OAI21_X1   g01659(.A1(new_n1851_), .A2(new_n1847_), .B(\asqrt[50] ), .ZN(new_n1852_));
  AOI21_X1   g01660(.A1(new_n1844_), .A2(new_n1852_), .B(new_n1305_), .ZN(new_n1853_));
  NOR3_X1    g01661(.A1(new_n1843_), .A2(\asqrt[52] ), .A3(new_n1853_), .ZN(new_n1854_));
  OAI21_X1   g01662(.A1(new_n1843_), .A2(new_n1853_), .B(\asqrt[52] ), .ZN(new_n1855_));
  OAI21_X1   g01663(.A1(new_n1806_), .A2(new_n1854_), .B(new_n1855_), .ZN(new_n1856_));
  OAI21_X1   g01664(.A1(new_n1856_), .A2(\asqrt[53] ), .B(new_n1803_), .ZN(new_n1857_));
  NAND2_X1   g01665(.A1(new_n1856_), .A2(\asqrt[53] ), .ZN(new_n1858_));
  NAND3_X1   g01666(.A1(new_n1857_), .A2(new_n1858_), .A3(new_n860_), .ZN(new_n1859_));
  AOI21_X1   g01667(.A1(new_n1857_), .A2(new_n1858_), .B(new_n860_), .ZN(new_n1860_));
  AOI21_X1   g01668(.A1(new_n1801_), .A2(new_n1859_), .B(new_n1860_), .ZN(new_n1861_));
  AOI21_X1   g01669(.A1(new_n1861_), .A2(new_n744_), .B(new_n1799_), .ZN(new_n1862_));
  NAND2_X1   g01670(.A1(new_n1859_), .A2(new_n1801_), .ZN(new_n1863_));
  INV_X1     g01671(.I(new_n1803_), .ZN(new_n1864_));
  NOR3_X1    g01672(.A1(new_n1851_), .A2(new_n1847_), .A3(\asqrt[50] ), .ZN(new_n1865_));
  OAI21_X1   g01673(.A1(new_n1823_), .A2(new_n1865_), .B(new_n1852_), .ZN(new_n1866_));
  OAI21_X1   g01674(.A1(new_n1866_), .A2(\asqrt[51] ), .B(new_n1812_), .ZN(new_n1867_));
  NAND2_X1   g01675(.A1(new_n1866_), .A2(\asqrt[51] ), .ZN(new_n1868_));
  NAND3_X1   g01676(.A1(new_n1867_), .A2(new_n1868_), .A3(new_n1150_), .ZN(new_n1869_));
  AOI21_X1   g01677(.A1(new_n1867_), .A2(new_n1868_), .B(new_n1150_), .ZN(new_n1870_));
  AOI21_X1   g01678(.A1(new_n1805_), .A2(new_n1869_), .B(new_n1870_), .ZN(new_n1871_));
  AOI21_X1   g01679(.A1(new_n1871_), .A2(new_n1006_), .B(new_n1864_), .ZN(new_n1872_));
  NAND2_X1   g01680(.A1(new_n1869_), .A2(new_n1805_), .ZN(new_n1873_));
  AOI21_X1   g01681(.A1(new_n1873_), .A2(new_n1855_), .B(new_n1006_), .ZN(new_n1874_));
  OAI21_X1   g01682(.A1(new_n1872_), .A2(new_n1874_), .B(\asqrt[54] ), .ZN(new_n1875_));
  AOI21_X1   g01683(.A1(new_n1863_), .A2(new_n1875_), .B(new_n744_), .ZN(new_n1876_));
  NOR3_X1    g01684(.A1(new_n1862_), .A2(\asqrt[56] ), .A3(new_n1876_), .ZN(new_n1877_));
  OAI21_X1   g01685(.A1(new_n1862_), .A2(new_n1876_), .B(\asqrt[56] ), .ZN(new_n1878_));
  OAI21_X1   g01686(.A1(new_n1795_), .A2(new_n1877_), .B(new_n1878_), .ZN(new_n1879_));
  OAI21_X1   g01687(.A1(new_n1879_), .A2(\asqrt[57] ), .B(new_n1791_), .ZN(new_n1880_));
  NAND2_X1   g01688(.A1(new_n1879_), .A2(\asqrt[57] ), .ZN(new_n1881_));
  NAND3_X1   g01689(.A1(new_n1880_), .A2(new_n1881_), .A3(new_n423_), .ZN(new_n1882_));
  AOI21_X1   g01690(.A1(new_n1880_), .A2(new_n1881_), .B(new_n423_), .ZN(new_n1883_));
  AOI21_X1   g01691(.A1(new_n1789_), .A2(new_n1882_), .B(new_n1883_), .ZN(new_n1884_));
  AOI21_X1   g01692(.A1(new_n1884_), .A2(new_n337_), .B(new_n1787_), .ZN(new_n1885_));
  NAND2_X1   g01693(.A1(new_n1882_), .A2(new_n1789_), .ZN(new_n1886_));
  INV_X1     g01694(.I(new_n1791_), .ZN(new_n1887_));
  INV_X1     g01695(.I(new_n1801_), .ZN(new_n1888_));
  NOR3_X1    g01696(.A1(new_n1872_), .A2(\asqrt[54] ), .A3(new_n1874_), .ZN(new_n1889_));
  OAI21_X1   g01697(.A1(new_n1888_), .A2(new_n1889_), .B(new_n1875_), .ZN(new_n1890_));
  OAI21_X1   g01698(.A1(new_n1890_), .A2(\asqrt[55] ), .B(new_n1798_), .ZN(new_n1891_));
  NAND2_X1   g01699(.A1(new_n1890_), .A2(\asqrt[55] ), .ZN(new_n1892_));
  NAND3_X1   g01700(.A1(new_n1891_), .A2(new_n1892_), .A3(new_n634_), .ZN(new_n1893_));
  AOI21_X1   g01701(.A1(new_n1891_), .A2(new_n1892_), .B(new_n634_), .ZN(new_n1894_));
  AOI21_X1   g01702(.A1(new_n1794_), .A2(new_n1893_), .B(new_n1894_), .ZN(new_n1895_));
  AOI21_X1   g01703(.A1(new_n1895_), .A2(new_n531_), .B(new_n1887_), .ZN(new_n1896_));
  NAND2_X1   g01704(.A1(new_n1893_), .A2(new_n1794_), .ZN(new_n1897_));
  AOI21_X1   g01705(.A1(new_n1897_), .A2(new_n1878_), .B(new_n531_), .ZN(new_n1898_));
  OAI21_X1   g01706(.A1(new_n1896_), .A2(new_n1898_), .B(\asqrt[58] ), .ZN(new_n1899_));
  AOI21_X1   g01707(.A1(new_n1886_), .A2(new_n1899_), .B(new_n337_), .ZN(new_n1900_));
  NOR3_X1    g01708(.A1(new_n1885_), .A2(\asqrt[60] ), .A3(new_n1900_), .ZN(new_n1901_));
  NOR2_X1    g01709(.A1(new_n1901_), .A2(new_n1784_), .ZN(new_n1902_));
  INV_X1     g01710(.I(new_n1789_), .ZN(new_n1903_));
  NOR3_X1    g01711(.A1(new_n1896_), .A2(\asqrt[58] ), .A3(new_n1898_), .ZN(new_n1904_));
  OAI21_X1   g01712(.A1(new_n1903_), .A2(new_n1904_), .B(new_n1899_), .ZN(new_n1905_));
  OAI21_X1   g01713(.A1(new_n1905_), .A2(\asqrt[59] ), .B(new_n1786_), .ZN(new_n1906_));
  NAND2_X1   g01714(.A1(new_n1905_), .A2(\asqrt[59] ), .ZN(new_n1907_));
  AOI21_X1   g01715(.A1(new_n1906_), .A2(new_n1907_), .B(new_n266_), .ZN(new_n1908_));
  OAI21_X1   g01716(.A1(new_n1902_), .A2(new_n1908_), .B(\asqrt[61] ), .ZN(new_n1909_));
  OAI21_X1   g01717(.A1(new_n1885_), .A2(new_n1900_), .B(\asqrt[60] ), .ZN(new_n1910_));
  OAI21_X1   g01718(.A1(new_n1784_), .A2(new_n1901_), .B(new_n1910_), .ZN(new_n1911_));
  AOI21_X1   g01719(.A1(new_n1751_), .A2(new_n1724_), .B(\asqrt[48] ), .ZN(new_n1912_));
  XOR2_X1    g01720(.A1(new_n1912_), .A2(new_n1599_), .Z(new_n1913_));
  OAI21_X1   g01721(.A1(new_n1911_), .A2(\asqrt[61] ), .B(new_n1913_), .ZN(new_n1914_));
  NAND2_X1   g01722(.A1(new_n1914_), .A2(new_n1909_), .ZN(new_n1915_));
  NAND3_X1   g01723(.A1(new_n1906_), .A2(new_n1907_), .A3(new_n266_), .ZN(new_n1916_));
  NAND2_X1   g01724(.A1(new_n1916_), .A2(new_n1783_), .ZN(new_n1917_));
  AOI21_X1   g01725(.A1(new_n1917_), .A2(new_n1910_), .B(new_n239_), .ZN(new_n1918_));
  AOI21_X1   g01726(.A1(new_n1783_), .A2(new_n1916_), .B(new_n1908_), .ZN(new_n1919_));
  INV_X1     g01727(.I(new_n1913_), .ZN(new_n1920_));
  AOI21_X1   g01728(.A1(new_n1919_), .A2(new_n239_), .B(new_n1920_), .ZN(new_n1921_));
  OAI21_X1   g01729(.A1(new_n1921_), .A2(new_n1918_), .B(new_n201_), .ZN(new_n1922_));
  NAND3_X1   g01730(.A1(new_n1914_), .A2(\asqrt[62] ), .A3(new_n1909_), .ZN(new_n1923_));
  AOI21_X1   g01731(.A1(new_n1747_), .A2(new_n1728_), .B(\asqrt[48] ), .ZN(new_n1924_));
  XOR2_X1    g01732(.A1(new_n1924_), .A2(new_n1727_), .Z(new_n1925_));
  INV_X1     g01733(.I(new_n1925_), .ZN(new_n1926_));
  AOI22_X1   g01734(.A1(new_n1923_), .A2(new_n1922_), .B1(new_n1915_), .B2(new_n1926_), .ZN(new_n1927_));
  NOR2_X1    g01735(.A1(new_n1757_), .A2(new_n1738_), .ZN(new_n1928_));
  OAI21_X1   g01736(.A1(\asqrt[48] ), .A2(new_n1928_), .B(new_n1737_), .ZN(new_n1929_));
  INV_X1     g01737(.I(new_n1929_), .ZN(new_n1930_));
  OAI21_X1   g01738(.A1(new_n1927_), .A2(new_n1781_), .B(new_n1930_), .ZN(new_n1931_));
  OAI21_X1   g01739(.A1(new_n1915_), .A2(\asqrt[62] ), .B(new_n1925_), .ZN(new_n1932_));
  NAND2_X1   g01740(.A1(new_n1915_), .A2(\asqrt[62] ), .ZN(new_n1933_));
  NAND3_X1   g01741(.A1(new_n1932_), .A2(new_n1933_), .A3(new_n1781_), .ZN(new_n1934_));
  NAND2_X1   g01742(.A1(new_n1778_), .A2(new_n1735_), .ZN(new_n1935_));
  XOR2_X1    g01743(.A1(new_n1757_), .A2(new_n1738_), .Z(new_n1936_));
  NAND3_X1   g01744(.A1(new_n1935_), .A2(\asqrt[63] ), .A3(new_n1936_), .ZN(new_n1937_));
  INV_X1     g01745(.I(new_n1814_), .ZN(new_n1938_));
  NAND4_X1   g01746(.A1(new_n1938_), .A2(new_n1738_), .A3(new_n1737_), .A4(new_n1768_), .ZN(new_n1939_));
  NAND2_X1   g01747(.A1(new_n1937_), .A2(new_n1939_), .ZN(new_n1940_));
  INV_X1     g01748(.I(new_n1940_), .ZN(new_n1941_));
  NAND4_X1   g01749(.A1(new_n1931_), .A2(new_n193_), .A3(new_n1934_), .A4(new_n1941_), .ZN(\asqrt[47] ));
  NOR2_X1    g01750(.A1(new_n1915_), .A2(\asqrt[62] ), .ZN(new_n1943_));
  NOR2_X1    g01751(.A1(new_n1921_), .A2(new_n1918_), .ZN(new_n1944_));
  NOR2_X1    g01752(.A1(new_n1944_), .A2(new_n201_), .ZN(new_n1945_));
  NOR2_X1    g01753(.A1(new_n1943_), .A2(new_n1945_), .ZN(new_n1946_));
  AOI21_X1   g01754(.A1(new_n1914_), .A2(new_n1909_), .B(\asqrt[62] ), .ZN(new_n1947_));
  NOR3_X1    g01755(.A1(new_n1921_), .A2(new_n201_), .A3(new_n1918_), .ZN(new_n1948_));
  OAI22_X1   g01756(.A1(new_n1947_), .A2(new_n1948_), .B1(new_n1944_), .B2(new_n1925_), .ZN(new_n1949_));
  AOI21_X1   g01757(.A1(new_n1949_), .A2(new_n1780_), .B(new_n1929_), .ZN(new_n1950_));
  AOI21_X1   g01758(.A1(new_n1944_), .A2(new_n201_), .B(new_n1926_), .ZN(new_n1951_));
  NOR3_X1    g01759(.A1(new_n1951_), .A2(new_n1945_), .A3(new_n1780_), .ZN(new_n1952_));
  NOR4_X1    g01760(.A1(new_n1950_), .A2(\asqrt[63] ), .A3(new_n1952_), .A4(new_n1940_), .ZN(new_n1953_));
  XOR2_X1    g01761(.A1(new_n1924_), .A2(new_n1727_), .Z(new_n1954_));
  OAI21_X1   g01762(.A1(\asqrt[47] ), .A2(new_n1946_), .B(new_n1954_), .ZN(new_n1955_));
  INV_X1     g01763(.I(new_n1955_), .ZN(new_n1956_));
  NAND2_X1   g01764(.A1(new_n1884_), .A2(new_n337_), .ZN(new_n1957_));
  AOI21_X1   g01765(.A1(new_n1957_), .A2(new_n1907_), .B(\asqrt[47] ), .ZN(new_n1958_));
  XOR2_X1    g01766(.A1(new_n1958_), .A2(new_n1786_), .Z(new_n1959_));
  INV_X1     g01767(.I(new_n1959_), .ZN(new_n1960_));
  AOI21_X1   g01768(.A1(new_n1882_), .A2(new_n1899_), .B(\asqrt[47] ), .ZN(new_n1961_));
  XOR2_X1    g01769(.A1(new_n1961_), .A2(new_n1789_), .Z(new_n1962_));
  INV_X1     g01770(.I(new_n1962_), .ZN(new_n1963_));
  NAND2_X1   g01771(.A1(new_n1895_), .A2(new_n531_), .ZN(new_n1964_));
  AOI21_X1   g01772(.A1(new_n1964_), .A2(new_n1881_), .B(\asqrt[47] ), .ZN(new_n1965_));
  XOR2_X1    g01773(.A1(new_n1965_), .A2(new_n1791_), .Z(new_n1966_));
  AOI21_X1   g01774(.A1(new_n1893_), .A2(new_n1878_), .B(\asqrt[47] ), .ZN(new_n1967_));
  XOR2_X1    g01775(.A1(new_n1967_), .A2(new_n1794_), .Z(new_n1968_));
  NAND2_X1   g01776(.A1(new_n1861_), .A2(new_n744_), .ZN(new_n1969_));
  AOI21_X1   g01777(.A1(new_n1969_), .A2(new_n1892_), .B(\asqrt[47] ), .ZN(new_n1970_));
  XOR2_X1    g01778(.A1(new_n1970_), .A2(new_n1798_), .Z(new_n1971_));
  INV_X1     g01779(.I(new_n1971_), .ZN(new_n1972_));
  AOI21_X1   g01780(.A1(new_n1859_), .A2(new_n1875_), .B(\asqrt[47] ), .ZN(new_n1973_));
  XOR2_X1    g01781(.A1(new_n1973_), .A2(new_n1801_), .Z(new_n1974_));
  INV_X1     g01782(.I(new_n1974_), .ZN(new_n1975_));
  NAND2_X1   g01783(.A1(new_n1871_), .A2(new_n1006_), .ZN(new_n1976_));
  AOI21_X1   g01784(.A1(new_n1976_), .A2(new_n1858_), .B(\asqrt[47] ), .ZN(new_n1977_));
  XOR2_X1    g01785(.A1(new_n1977_), .A2(new_n1803_), .Z(new_n1978_));
  AOI21_X1   g01786(.A1(new_n1869_), .A2(new_n1855_), .B(\asqrt[47] ), .ZN(new_n1979_));
  XOR2_X1    g01787(.A1(new_n1979_), .A2(new_n1805_), .Z(new_n1980_));
  NAND2_X1   g01788(.A1(new_n1842_), .A2(new_n1305_), .ZN(new_n1981_));
  AOI21_X1   g01789(.A1(new_n1981_), .A2(new_n1868_), .B(\asqrt[47] ), .ZN(new_n1982_));
  XOR2_X1    g01790(.A1(new_n1982_), .A2(new_n1812_), .Z(new_n1983_));
  INV_X1     g01791(.I(new_n1983_), .ZN(new_n1984_));
  AOI21_X1   g01792(.A1(new_n1840_), .A2(new_n1852_), .B(\asqrt[47] ), .ZN(new_n1985_));
  XOR2_X1    g01793(.A1(new_n1985_), .A2(new_n1824_), .Z(new_n1986_));
  INV_X1     g01794(.I(new_n1986_), .ZN(new_n1987_));
  NAND2_X1   g01795(.A1(\asqrt[48] ), .A2(new_n1825_), .ZN(new_n1988_));
  NOR2_X1    g01796(.A1(new_n1837_), .A2(\a[96] ), .ZN(new_n1989_));
  AOI22_X1   g01797(.A1(new_n1988_), .A2(new_n1837_), .B1(\asqrt[48] ), .B2(new_n1989_), .ZN(new_n1990_));
  AOI21_X1   g01798(.A1(\asqrt[48] ), .A2(\a[96] ), .B(new_n1833_), .ZN(new_n1991_));
  OAI21_X1   g01799(.A1(new_n1847_), .A2(new_n1991_), .B(new_n1953_), .ZN(new_n1992_));
  XNOR2_X1   g01800(.A1(new_n1992_), .A2(new_n1990_), .ZN(new_n1993_));
  NOR3_X1    g01801(.A1(new_n1950_), .A2(\asqrt[63] ), .A3(new_n1952_), .ZN(new_n1994_));
  NAND4_X1   g01802(.A1(new_n1994_), .A2(\asqrt[48] ), .A3(new_n1937_), .A4(new_n1939_), .ZN(new_n1995_));
  NAND2_X1   g01803(.A1(\asqrt[47] ), .A2(new_n1826_), .ZN(new_n1996_));
  AOI21_X1   g01804(.A1(new_n1995_), .A2(new_n1996_), .B(\a[96] ), .ZN(new_n1997_));
  NAND2_X1   g01805(.A1(new_n1931_), .A2(new_n193_), .ZN(new_n1998_));
  NAND3_X1   g01806(.A1(new_n1937_), .A2(\asqrt[48] ), .A3(new_n1939_), .ZN(new_n1999_));
  NOR3_X1    g01807(.A1(new_n1998_), .A2(new_n1952_), .A3(new_n1999_), .ZN(new_n2000_));
  NOR2_X1    g01808(.A1(new_n1953_), .A2(new_n1828_), .ZN(new_n2001_));
  NOR3_X1    g01809(.A1(new_n2001_), .A2(new_n2000_), .A3(new_n1825_), .ZN(new_n2002_));
  NOR2_X1    g01810(.A1(new_n1997_), .A2(new_n2002_), .ZN(new_n2003_));
  INV_X1     g01811(.I(\a[94] ), .ZN(new_n2004_));
  NOR2_X1    g01812(.A1(\a[92] ), .A2(\a[93] ), .ZN(new_n2005_));
  NOR3_X1    g01813(.A1(new_n1953_), .A2(new_n2004_), .A3(new_n2005_), .ZN(new_n2006_));
  INV_X1     g01814(.I(new_n2005_), .ZN(new_n2007_));
  AOI21_X1   g01815(.A1(new_n1953_), .A2(\a[94] ), .B(new_n2007_), .ZN(new_n2008_));
  OAI21_X1   g01816(.A1(new_n2006_), .A2(new_n2008_), .B(\asqrt[48] ), .ZN(new_n2009_));
  NAND2_X1   g01817(.A1(new_n2005_), .A2(new_n2004_), .ZN(new_n2010_));
  NAND3_X1   g01818(.A1(new_n1764_), .A2(new_n1766_), .A3(new_n2010_), .ZN(new_n2011_));
  NAND2_X1   g01819(.A1(new_n1819_), .A2(new_n2011_), .ZN(new_n2012_));
  NAND3_X1   g01820(.A1(\asqrt[47] ), .A2(\a[94] ), .A3(new_n2012_), .ZN(new_n2013_));
  NOR3_X1    g01821(.A1(new_n1953_), .A2(\a[94] ), .A3(\a[95] ), .ZN(new_n2014_));
  INV_X1     g01822(.I(\a[95] ), .ZN(new_n2015_));
  AOI21_X1   g01823(.A1(\asqrt[47] ), .A2(new_n2004_), .B(new_n2015_), .ZN(new_n2016_));
  NOR2_X1    g01824(.A1(new_n2014_), .A2(new_n2016_), .ZN(new_n2017_));
  NAND4_X1   g01825(.A1(new_n2009_), .A2(new_n2017_), .A3(new_n1632_), .A4(new_n2013_), .ZN(new_n2018_));
  NAND2_X1   g01826(.A1(new_n2018_), .A2(new_n2003_), .ZN(new_n2019_));
  NAND3_X1   g01827(.A1(\asqrt[47] ), .A2(\a[94] ), .A3(new_n2007_), .ZN(new_n2020_));
  OAI21_X1   g01828(.A1(\asqrt[47] ), .A2(new_n2004_), .B(new_n2005_), .ZN(new_n2021_));
  AOI21_X1   g01829(.A1(new_n2021_), .A2(new_n2020_), .B(new_n1778_), .ZN(new_n2022_));
  NAND3_X1   g01830(.A1(\asqrt[47] ), .A2(new_n2004_), .A3(new_n2015_), .ZN(new_n2023_));
  OAI21_X1   g01831(.A1(new_n1953_), .A2(\a[94] ), .B(\a[95] ), .ZN(new_n2024_));
  NAND3_X1   g01832(.A1(new_n2013_), .A2(new_n2024_), .A3(new_n2023_), .ZN(new_n2025_));
  OAI21_X1   g01833(.A1(new_n2025_), .A2(new_n2022_), .B(\asqrt[49] ), .ZN(new_n2026_));
  NAND3_X1   g01834(.A1(new_n2019_), .A2(new_n1463_), .A3(new_n2026_), .ZN(new_n2027_));
  AOI21_X1   g01835(.A1(new_n2019_), .A2(new_n2026_), .B(new_n1463_), .ZN(new_n2028_));
  AOI21_X1   g01836(.A1(new_n1993_), .A2(new_n2027_), .B(new_n2028_), .ZN(new_n2029_));
  AOI21_X1   g01837(.A1(new_n2029_), .A2(new_n1305_), .B(new_n1987_), .ZN(new_n2030_));
  OR2_X2     g01838(.A1(new_n1997_), .A2(new_n2002_), .Z(new_n2031_));
  NOR3_X1    g01839(.A1(new_n2025_), .A2(new_n2022_), .A3(\asqrt[49] ), .ZN(new_n2032_));
  OAI21_X1   g01840(.A1(new_n2031_), .A2(new_n2032_), .B(new_n2026_), .ZN(new_n2033_));
  OAI21_X1   g01841(.A1(new_n2033_), .A2(\asqrt[50] ), .B(new_n1993_), .ZN(new_n2034_));
  NAND2_X1   g01842(.A1(new_n2033_), .A2(\asqrt[50] ), .ZN(new_n2035_));
  AOI21_X1   g01843(.A1(new_n2034_), .A2(new_n2035_), .B(new_n1305_), .ZN(new_n2036_));
  NOR3_X1    g01844(.A1(new_n2030_), .A2(\asqrt[52] ), .A3(new_n2036_), .ZN(new_n2037_));
  OAI21_X1   g01845(.A1(new_n2030_), .A2(new_n2036_), .B(\asqrt[52] ), .ZN(new_n2038_));
  OAI21_X1   g01846(.A1(new_n1984_), .A2(new_n2037_), .B(new_n2038_), .ZN(new_n2039_));
  OAI21_X1   g01847(.A1(new_n2039_), .A2(\asqrt[53] ), .B(new_n1980_), .ZN(new_n2040_));
  NAND3_X1   g01848(.A1(new_n2034_), .A2(new_n2035_), .A3(new_n1305_), .ZN(new_n2041_));
  AOI21_X1   g01849(.A1(new_n1986_), .A2(new_n2041_), .B(new_n2036_), .ZN(new_n2042_));
  AOI21_X1   g01850(.A1(new_n2042_), .A2(new_n1150_), .B(new_n1984_), .ZN(new_n2043_));
  NAND2_X1   g01851(.A1(new_n2041_), .A2(new_n1986_), .ZN(new_n2044_));
  INV_X1     g01852(.I(new_n2036_), .ZN(new_n2045_));
  AOI21_X1   g01853(.A1(new_n2044_), .A2(new_n2045_), .B(new_n1150_), .ZN(new_n2046_));
  OAI21_X1   g01854(.A1(new_n2043_), .A2(new_n2046_), .B(\asqrt[53] ), .ZN(new_n2047_));
  NAND3_X1   g01855(.A1(new_n2040_), .A2(new_n860_), .A3(new_n2047_), .ZN(new_n2048_));
  AOI21_X1   g01856(.A1(new_n2040_), .A2(new_n2047_), .B(new_n860_), .ZN(new_n2049_));
  AOI21_X1   g01857(.A1(new_n1978_), .A2(new_n2048_), .B(new_n2049_), .ZN(new_n2050_));
  AOI21_X1   g01858(.A1(new_n2050_), .A2(new_n744_), .B(new_n1975_), .ZN(new_n2051_));
  INV_X1     g01859(.I(new_n1980_), .ZN(new_n2052_));
  NOR3_X1    g01860(.A1(new_n2043_), .A2(\asqrt[53] ), .A3(new_n2046_), .ZN(new_n2053_));
  OAI21_X1   g01861(.A1(new_n2052_), .A2(new_n2053_), .B(new_n2047_), .ZN(new_n2054_));
  OAI21_X1   g01862(.A1(new_n2054_), .A2(\asqrt[54] ), .B(new_n1978_), .ZN(new_n2055_));
  NAND2_X1   g01863(.A1(new_n2054_), .A2(\asqrt[54] ), .ZN(new_n2056_));
  AOI21_X1   g01864(.A1(new_n2055_), .A2(new_n2056_), .B(new_n744_), .ZN(new_n2057_));
  NOR3_X1    g01865(.A1(new_n2051_), .A2(\asqrt[56] ), .A3(new_n2057_), .ZN(new_n2058_));
  OAI21_X1   g01866(.A1(new_n2051_), .A2(new_n2057_), .B(\asqrt[56] ), .ZN(new_n2059_));
  OAI21_X1   g01867(.A1(new_n1972_), .A2(new_n2058_), .B(new_n2059_), .ZN(new_n2060_));
  OAI21_X1   g01868(.A1(new_n2060_), .A2(\asqrt[57] ), .B(new_n1968_), .ZN(new_n2061_));
  NAND3_X1   g01869(.A1(new_n2055_), .A2(new_n2056_), .A3(new_n744_), .ZN(new_n2062_));
  AOI21_X1   g01870(.A1(new_n1974_), .A2(new_n2062_), .B(new_n2057_), .ZN(new_n2063_));
  AOI21_X1   g01871(.A1(new_n2063_), .A2(new_n634_), .B(new_n1972_), .ZN(new_n2064_));
  NAND2_X1   g01872(.A1(new_n2062_), .A2(new_n1974_), .ZN(new_n2065_));
  INV_X1     g01873(.I(new_n2057_), .ZN(new_n2066_));
  AOI21_X1   g01874(.A1(new_n2065_), .A2(new_n2066_), .B(new_n634_), .ZN(new_n2067_));
  OAI21_X1   g01875(.A1(new_n2064_), .A2(new_n2067_), .B(\asqrt[57] ), .ZN(new_n2068_));
  NAND3_X1   g01876(.A1(new_n2061_), .A2(new_n423_), .A3(new_n2068_), .ZN(new_n2069_));
  AOI21_X1   g01877(.A1(new_n2061_), .A2(new_n2068_), .B(new_n423_), .ZN(new_n2070_));
  AOI21_X1   g01878(.A1(new_n1966_), .A2(new_n2069_), .B(new_n2070_), .ZN(new_n2071_));
  AOI21_X1   g01879(.A1(new_n2071_), .A2(new_n337_), .B(new_n1963_), .ZN(new_n2072_));
  NOR2_X1    g01880(.A1(new_n2071_), .A2(new_n337_), .ZN(new_n2073_));
  NOR3_X1    g01881(.A1(new_n2072_), .A2(new_n2073_), .A3(\asqrt[60] ), .ZN(new_n2074_));
  OAI21_X1   g01882(.A1(new_n2072_), .A2(new_n2073_), .B(\asqrt[60] ), .ZN(new_n2075_));
  OAI21_X1   g01883(.A1(new_n1960_), .A2(new_n2074_), .B(new_n2075_), .ZN(new_n2076_));
  NAND2_X1   g01884(.A1(new_n2076_), .A2(\asqrt[61] ), .ZN(new_n2077_));
  AOI21_X1   g01885(.A1(new_n1916_), .A2(new_n1910_), .B(\asqrt[47] ), .ZN(new_n2078_));
  XOR2_X1    g01886(.A1(new_n2078_), .A2(new_n1783_), .Z(new_n2079_));
  OAI21_X1   g01887(.A1(new_n2076_), .A2(\asqrt[61] ), .B(new_n2079_), .ZN(new_n2080_));
  NAND2_X1   g01888(.A1(new_n2080_), .A2(new_n2077_), .ZN(new_n2081_));
  INV_X1     g01889(.I(new_n1968_), .ZN(new_n2082_));
  NOR3_X1    g01890(.A1(new_n2064_), .A2(\asqrt[57] ), .A3(new_n2067_), .ZN(new_n2083_));
  OAI21_X1   g01891(.A1(new_n2082_), .A2(new_n2083_), .B(new_n2068_), .ZN(new_n2084_));
  OAI21_X1   g01892(.A1(new_n2084_), .A2(\asqrt[58] ), .B(new_n1966_), .ZN(new_n2085_));
  NOR2_X1    g01893(.A1(new_n2083_), .A2(new_n2082_), .ZN(new_n2086_));
  INV_X1     g01894(.I(new_n2068_), .ZN(new_n2087_));
  OAI21_X1   g01895(.A1(new_n2086_), .A2(new_n2087_), .B(\asqrt[58] ), .ZN(new_n2088_));
  NAND3_X1   g01896(.A1(new_n2085_), .A2(new_n337_), .A3(new_n2088_), .ZN(new_n2089_));
  NAND2_X1   g01897(.A1(new_n2089_), .A2(new_n1962_), .ZN(new_n2090_));
  INV_X1     g01898(.I(new_n1966_), .ZN(new_n2091_));
  NOR2_X1    g01899(.A1(new_n2086_), .A2(new_n2087_), .ZN(new_n2092_));
  AOI21_X1   g01900(.A1(new_n2092_), .A2(new_n423_), .B(new_n2091_), .ZN(new_n2093_));
  OAI21_X1   g01901(.A1(new_n2093_), .A2(new_n2070_), .B(\asqrt[59] ), .ZN(new_n2094_));
  NAND3_X1   g01902(.A1(new_n2090_), .A2(new_n266_), .A3(new_n2094_), .ZN(new_n2095_));
  NAND2_X1   g01903(.A1(new_n2095_), .A2(new_n1959_), .ZN(new_n2096_));
  AOI21_X1   g01904(.A1(new_n2096_), .A2(new_n2075_), .B(new_n239_), .ZN(new_n2097_));
  AOI21_X1   g01905(.A1(new_n2090_), .A2(new_n2094_), .B(new_n266_), .ZN(new_n2098_));
  AOI21_X1   g01906(.A1(new_n1959_), .A2(new_n2095_), .B(new_n2098_), .ZN(new_n2099_));
  INV_X1     g01907(.I(new_n2079_), .ZN(new_n2100_));
  AOI21_X1   g01908(.A1(new_n2099_), .A2(new_n239_), .B(new_n2100_), .ZN(new_n2101_));
  OAI21_X1   g01909(.A1(new_n2101_), .A2(new_n2097_), .B(new_n201_), .ZN(new_n2102_));
  NAND3_X1   g01910(.A1(new_n2080_), .A2(new_n2077_), .A3(\asqrt[62] ), .ZN(new_n2103_));
  NAND2_X1   g01911(.A1(new_n1919_), .A2(new_n239_), .ZN(new_n2104_));
  AOI21_X1   g01912(.A1(new_n1909_), .A2(new_n2104_), .B(\asqrt[47] ), .ZN(new_n2105_));
  XOR2_X1    g01913(.A1(new_n2105_), .A2(new_n1913_), .Z(new_n2106_));
  INV_X1     g01914(.I(new_n2106_), .ZN(new_n2107_));
  AOI22_X1   g01915(.A1(new_n2103_), .A2(new_n2102_), .B1(new_n2081_), .B2(new_n2107_), .ZN(new_n2108_));
  NOR2_X1    g01916(.A1(new_n1927_), .A2(new_n1781_), .ZN(new_n2109_));
  OAI21_X1   g01917(.A1(\asqrt[47] ), .A2(new_n2109_), .B(new_n1934_), .ZN(new_n2110_));
  INV_X1     g01918(.I(new_n2110_), .ZN(new_n2111_));
  OAI21_X1   g01919(.A1(new_n2108_), .A2(new_n1956_), .B(new_n2111_), .ZN(new_n2112_));
  OAI21_X1   g01920(.A1(new_n2081_), .A2(\asqrt[62] ), .B(new_n2106_), .ZN(new_n2113_));
  NAND2_X1   g01921(.A1(new_n2081_), .A2(\asqrt[62] ), .ZN(new_n2114_));
  NAND3_X1   g01922(.A1(new_n2113_), .A2(new_n2114_), .A3(new_n1956_), .ZN(new_n2115_));
  NAND2_X1   g01923(.A1(new_n1953_), .A2(new_n1780_), .ZN(new_n2116_));
  XOR2_X1    g01924(.A1(new_n1949_), .A2(new_n1780_), .Z(new_n2117_));
  NAND3_X1   g01925(.A1(new_n2116_), .A2(\asqrt[63] ), .A3(new_n2117_), .ZN(new_n2118_));
  INV_X1     g01926(.I(new_n1998_), .ZN(new_n2119_));
  NAND4_X1   g01927(.A1(new_n2119_), .A2(new_n1781_), .A3(new_n1934_), .A4(new_n1941_), .ZN(new_n2120_));
  NAND2_X1   g01928(.A1(new_n2118_), .A2(new_n2120_), .ZN(new_n2121_));
  INV_X1     g01929(.I(new_n2121_), .ZN(new_n2122_));
  NAND4_X1   g01930(.A1(new_n2112_), .A2(new_n193_), .A3(new_n2115_), .A4(new_n2122_), .ZN(\asqrt[46] ));
  NOR2_X1    g01931(.A1(new_n2081_), .A2(\asqrt[62] ), .ZN(new_n2124_));
  NOR2_X1    g01932(.A1(new_n2101_), .A2(new_n2097_), .ZN(new_n2125_));
  NOR2_X1    g01933(.A1(new_n2125_), .A2(new_n201_), .ZN(new_n2126_));
  NOR2_X1    g01934(.A1(new_n2124_), .A2(new_n2126_), .ZN(new_n2127_));
  AOI21_X1   g01935(.A1(new_n2080_), .A2(new_n2077_), .B(\asqrt[62] ), .ZN(new_n2128_));
  NOR3_X1    g01936(.A1(new_n2101_), .A2(new_n201_), .A3(new_n2097_), .ZN(new_n2129_));
  OAI22_X1   g01937(.A1(new_n2128_), .A2(new_n2129_), .B1(new_n2125_), .B2(new_n2106_), .ZN(new_n2130_));
  AOI21_X1   g01938(.A1(new_n2130_), .A2(new_n1955_), .B(new_n2110_), .ZN(new_n2131_));
  AOI21_X1   g01939(.A1(new_n2125_), .A2(new_n201_), .B(new_n2107_), .ZN(new_n2132_));
  NOR3_X1    g01940(.A1(new_n2132_), .A2(new_n2126_), .A3(new_n1955_), .ZN(new_n2133_));
  NOR4_X1    g01941(.A1(new_n2131_), .A2(\asqrt[63] ), .A3(new_n2133_), .A4(new_n2121_), .ZN(new_n2134_));
  XOR2_X1    g01942(.A1(new_n2105_), .A2(new_n1913_), .Z(new_n2135_));
  OAI21_X1   g01943(.A1(\asqrt[46] ), .A2(new_n2127_), .B(new_n2135_), .ZN(new_n2136_));
  INV_X1     g01944(.I(new_n2136_), .ZN(new_n2137_));
  AOI21_X1   g01945(.A1(new_n2089_), .A2(new_n2094_), .B(\asqrt[46] ), .ZN(new_n2138_));
  XOR2_X1    g01946(.A1(new_n2138_), .A2(new_n1962_), .Z(new_n2139_));
  INV_X1     g01947(.I(new_n2139_), .ZN(new_n2140_));
  AOI21_X1   g01948(.A1(new_n2069_), .A2(new_n2088_), .B(\asqrt[46] ), .ZN(new_n2141_));
  XOR2_X1    g01949(.A1(new_n2141_), .A2(new_n1966_), .Z(new_n2142_));
  INV_X1     g01950(.I(new_n2142_), .ZN(new_n2143_));
  NOR2_X1    g01951(.A1(new_n2087_), .A2(new_n2083_), .ZN(new_n2144_));
  NOR2_X1    g01952(.A1(\asqrt[46] ), .A2(new_n2144_), .ZN(new_n2145_));
  XOR2_X1    g01953(.A1(new_n2145_), .A2(new_n1968_), .Z(new_n2146_));
  NOR2_X1    g01954(.A1(new_n2058_), .A2(new_n2067_), .ZN(new_n2147_));
  NOR2_X1    g01955(.A1(\asqrt[46] ), .A2(new_n2147_), .ZN(new_n2148_));
  XOR2_X1    g01956(.A1(new_n2148_), .A2(new_n1971_), .Z(new_n2149_));
  AOI21_X1   g01957(.A1(new_n2062_), .A2(new_n2066_), .B(\asqrt[46] ), .ZN(new_n2150_));
  XOR2_X1    g01958(.A1(new_n2150_), .A2(new_n1974_), .Z(new_n2151_));
  INV_X1     g01959(.I(new_n2151_), .ZN(new_n2152_));
  AOI21_X1   g01960(.A1(new_n2048_), .A2(new_n2056_), .B(\asqrt[46] ), .ZN(new_n2153_));
  XOR2_X1    g01961(.A1(new_n2153_), .A2(new_n1978_), .Z(new_n2154_));
  INV_X1     g01962(.I(new_n2154_), .ZN(new_n2155_));
  XOR2_X1    g01963(.A1(new_n2039_), .A2(\asqrt[53] ), .Z(new_n2156_));
  NOR2_X1    g01964(.A1(\asqrt[46] ), .A2(new_n2156_), .ZN(new_n2157_));
  XOR2_X1    g01965(.A1(new_n2157_), .A2(new_n1980_), .Z(new_n2158_));
  NOR2_X1    g01966(.A1(new_n2037_), .A2(new_n2046_), .ZN(new_n2159_));
  NOR2_X1    g01967(.A1(\asqrt[46] ), .A2(new_n2159_), .ZN(new_n2160_));
  XOR2_X1    g01968(.A1(new_n2160_), .A2(new_n1983_), .Z(new_n2161_));
  AOI21_X1   g01969(.A1(new_n2041_), .A2(new_n2045_), .B(\asqrt[46] ), .ZN(new_n2162_));
  XOR2_X1    g01970(.A1(new_n2162_), .A2(new_n1986_), .Z(new_n2163_));
  INV_X1     g01971(.I(new_n2163_), .ZN(new_n2164_));
  AOI21_X1   g01972(.A1(new_n2027_), .A2(new_n2035_), .B(\asqrt[46] ), .ZN(new_n2165_));
  XOR2_X1    g01973(.A1(new_n2165_), .A2(new_n1993_), .Z(new_n2166_));
  INV_X1     g01974(.I(new_n2166_), .ZN(new_n2167_));
  AOI21_X1   g01975(.A1(new_n2018_), .A2(new_n2026_), .B(\asqrt[46] ), .ZN(new_n2168_));
  XOR2_X1    g01976(.A1(new_n2168_), .A2(new_n2003_), .Z(new_n2169_));
  NAND2_X1   g01977(.A1(\asqrt[47] ), .A2(new_n2004_), .ZN(new_n2170_));
  NOR2_X1    g01978(.A1(new_n2015_), .A2(\a[94] ), .ZN(new_n2171_));
  AOI22_X1   g01979(.A1(new_n2170_), .A2(new_n2015_), .B1(\asqrt[47] ), .B2(new_n2171_), .ZN(new_n2172_));
  AOI21_X1   g01980(.A1(\asqrt[47] ), .A2(\a[94] ), .B(new_n2012_), .ZN(new_n2173_));
  OAI21_X1   g01981(.A1(new_n2022_), .A2(new_n2173_), .B(new_n2134_), .ZN(new_n2174_));
  XNOR2_X1   g01982(.A1(new_n2174_), .A2(new_n2172_), .ZN(new_n2175_));
  NOR3_X1    g01983(.A1(new_n2131_), .A2(\asqrt[63] ), .A3(new_n2133_), .ZN(new_n2176_));
  NAND4_X1   g01984(.A1(new_n2176_), .A2(\asqrt[47] ), .A3(new_n2118_), .A4(new_n2120_), .ZN(new_n2177_));
  NAND2_X1   g01985(.A1(\asqrt[46] ), .A2(new_n2005_), .ZN(new_n2178_));
  AOI21_X1   g01986(.A1(new_n2177_), .A2(new_n2178_), .B(\a[94] ), .ZN(new_n2179_));
  NAND2_X1   g01987(.A1(new_n2112_), .A2(new_n193_), .ZN(new_n2180_));
  NAND3_X1   g01988(.A1(new_n2118_), .A2(\asqrt[47] ), .A3(new_n2120_), .ZN(new_n2181_));
  NOR3_X1    g01989(.A1(new_n2180_), .A2(new_n2133_), .A3(new_n2181_), .ZN(new_n2182_));
  NOR2_X1    g01990(.A1(new_n2134_), .A2(new_n2007_), .ZN(new_n2183_));
  NOR3_X1    g01991(.A1(new_n2183_), .A2(new_n2182_), .A3(new_n2004_), .ZN(new_n2184_));
  OR2_X2     g01992(.A1(new_n2179_), .A2(new_n2184_), .Z(new_n2185_));
  NOR2_X1    g01993(.A1(\a[90] ), .A2(\a[91] ), .ZN(new_n2186_));
  INV_X1     g01994(.I(new_n2186_), .ZN(new_n2187_));
  NAND3_X1   g01995(.A1(\asqrt[46] ), .A2(\a[92] ), .A3(new_n2187_), .ZN(new_n2188_));
  INV_X1     g01996(.I(\a[92] ), .ZN(new_n2189_));
  OAI21_X1   g01997(.A1(\asqrt[46] ), .A2(new_n2189_), .B(new_n2186_), .ZN(new_n2190_));
  AOI21_X1   g01998(.A1(new_n2190_), .A2(new_n2188_), .B(new_n1953_), .ZN(new_n2191_));
  NAND2_X1   g01999(.A1(new_n2186_), .A2(new_n2189_), .ZN(new_n2192_));
  NAND3_X1   g02000(.A1(new_n1937_), .A2(new_n1939_), .A3(new_n2192_), .ZN(new_n2193_));
  NAND2_X1   g02001(.A1(new_n1994_), .A2(new_n2193_), .ZN(new_n2194_));
  NAND3_X1   g02002(.A1(\asqrt[46] ), .A2(\a[92] ), .A3(new_n2194_), .ZN(new_n2195_));
  INV_X1     g02003(.I(\a[93] ), .ZN(new_n2196_));
  NAND3_X1   g02004(.A1(\asqrt[46] ), .A2(new_n2189_), .A3(new_n2196_), .ZN(new_n2197_));
  OAI21_X1   g02005(.A1(new_n2134_), .A2(\a[92] ), .B(\a[93] ), .ZN(new_n2198_));
  NAND3_X1   g02006(.A1(new_n2195_), .A2(new_n2198_), .A3(new_n2197_), .ZN(new_n2199_));
  NOR3_X1    g02007(.A1(new_n2199_), .A2(new_n2191_), .A3(\asqrt[48] ), .ZN(new_n2200_));
  OAI21_X1   g02008(.A1(new_n2199_), .A2(new_n2191_), .B(\asqrt[48] ), .ZN(new_n2201_));
  OAI21_X1   g02009(.A1(new_n2185_), .A2(new_n2200_), .B(new_n2201_), .ZN(new_n2202_));
  OAI21_X1   g02010(.A1(new_n2202_), .A2(\asqrt[49] ), .B(new_n2175_), .ZN(new_n2203_));
  NAND2_X1   g02011(.A1(new_n2202_), .A2(\asqrt[49] ), .ZN(new_n2204_));
  NAND3_X1   g02012(.A1(new_n2203_), .A2(new_n2204_), .A3(new_n1463_), .ZN(new_n2205_));
  AOI21_X1   g02013(.A1(new_n2203_), .A2(new_n2204_), .B(new_n1463_), .ZN(new_n2206_));
  AOI21_X1   g02014(.A1(new_n2169_), .A2(new_n2205_), .B(new_n2206_), .ZN(new_n2207_));
  AOI21_X1   g02015(.A1(new_n2207_), .A2(new_n1305_), .B(new_n2167_), .ZN(new_n2208_));
  NAND2_X1   g02016(.A1(new_n2205_), .A2(new_n2169_), .ZN(new_n2209_));
  INV_X1     g02017(.I(new_n2175_), .ZN(new_n2210_));
  NOR2_X1    g02018(.A1(new_n2179_), .A2(new_n2184_), .ZN(new_n2211_));
  NOR3_X1    g02019(.A1(new_n2134_), .A2(new_n2189_), .A3(new_n2186_), .ZN(new_n2212_));
  AOI21_X1   g02020(.A1(new_n2134_), .A2(\a[92] ), .B(new_n2187_), .ZN(new_n2213_));
  OAI21_X1   g02021(.A1(new_n2212_), .A2(new_n2213_), .B(\asqrt[47] ), .ZN(new_n2214_));
  INV_X1     g02022(.I(new_n2194_), .ZN(new_n2215_));
  NOR3_X1    g02023(.A1(new_n2134_), .A2(new_n2189_), .A3(new_n2215_), .ZN(new_n2216_));
  NOR3_X1    g02024(.A1(new_n2134_), .A2(\a[92] ), .A3(\a[93] ), .ZN(new_n2217_));
  AOI21_X1   g02025(.A1(\asqrt[46] ), .A2(new_n2189_), .B(new_n2196_), .ZN(new_n2218_));
  NOR3_X1    g02026(.A1(new_n2216_), .A2(new_n2217_), .A3(new_n2218_), .ZN(new_n2219_));
  NAND3_X1   g02027(.A1(new_n2219_), .A2(new_n2214_), .A3(new_n1778_), .ZN(new_n2220_));
  AOI21_X1   g02028(.A1(new_n2219_), .A2(new_n2214_), .B(new_n1778_), .ZN(new_n2221_));
  AOI21_X1   g02029(.A1(new_n2211_), .A2(new_n2220_), .B(new_n2221_), .ZN(new_n2222_));
  AOI21_X1   g02030(.A1(new_n2222_), .A2(new_n1632_), .B(new_n2210_), .ZN(new_n2223_));
  NAND2_X1   g02031(.A1(new_n2220_), .A2(new_n2211_), .ZN(new_n2224_));
  AOI21_X1   g02032(.A1(new_n2224_), .A2(new_n2201_), .B(new_n1632_), .ZN(new_n2225_));
  OAI21_X1   g02033(.A1(new_n2223_), .A2(new_n2225_), .B(\asqrt[50] ), .ZN(new_n2226_));
  AOI21_X1   g02034(.A1(new_n2209_), .A2(new_n2226_), .B(new_n1305_), .ZN(new_n2227_));
  NOR3_X1    g02035(.A1(new_n2208_), .A2(\asqrt[52] ), .A3(new_n2227_), .ZN(new_n2228_));
  OAI21_X1   g02036(.A1(new_n2208_), .A2(new_n2227_), .B(\asqrt[52] ), .ZN(new_n2229_));
  OAI21_X1   g02037(.A1(new_n2164_), .A2(new_n2228_), .B(new_n2229_), .ZN(new_n2230_));
  OAI21_X1   g02038(.A1(new_n2230_), .A2(\asqrt[53] ), .B(new_n2161_), .ZN(new_n2231_));
  NAND2_X1   g02039(.A1(new_n2230_), .A2(\asqrt[53] ), .ZN(new_n2232_));
  NAND3_X1   g02040(.A1(new_n2231_), .A2(new_n2232_), .A3(new_n860_), .ZN(new_n2233_));
  AOI21_X1   g02041(.A1(new_n2231_), .A2(new_n2232_), .B(new_n860_), .ZN(new_n2234_));
  AOI21_X1   g02042(.A1(new_n2158_), .A2(new_n2233_), .B(new_n2234_), .ZN(new_n2235_));
  AOI21_X1   g02043(.A1(new_n2235_), .A2(new_n744_), .B(new_n2155_), .ZN(new_n2236_));
  NAND2_X1   g02044(.A1(new_n2233_), .A2(new_n2158_), .ZN(new_n2237_));
  INV_X1     g02045(.I(new_n2161_), .ZN(new_n2238_));
  INV_X1     g02046(.I(new_n2169_), .ZN(new_n2239_));
  NOR3_X1    g02047(.A1(new_n2223_), .A2(\asqrt[50] ), .A3(new_n2225_), .ZN(new_n2240_));
  OAI21_X1   g02048(.A1(new_n2239_), .A2(new_n2240_), .B(new_n2226_), .ZN(new_n2241_));
  OAI21_X1   g02049(.A1(new_n2241_), .A2(\asqrt[51] ), .B(new_n2166_), .ZN(new_n2242_));
  NAND2_X1   g02050(.A1(new_n2241_), .A2(\asqrt[51] ), .ZN(new_n2243_));
  NAND3_X1   g02051(.A1(new_n2242_), .A2(new_n2243_), .A3(new_n1150_), .ZN(new_n2244_));
  AOI21_X1   g02052(.A1(new_n2242_), .A2(new_n2243_), .B(new_n1150_), .ZN(new_n2245_));
  AOI21_X1   g02053(.A1(new_n2163_), .A2(new_n2244_), .B(new_n2245_), .ZN(new_n2246_));
  AOI21_X1   g02054(.A1(new_n2246_), .A2(new_n1006_), .B(new_n2238_), .ZN(new_n2247_));
  NAND2_X1   g02055(.A1(new_n2244_), .A2(new_n2163_), .ZN(new_n2248_));
  AOI21_X1   g02056(.A1(new_n2248_), .A2(new_n2229_), .B(new_n1006_), .ZN(new_n2249_));
  OAI21_X1   g02057(.A1(new_n2247_), .A2(new_n2249_), .B(\asqrt[54] ), .ZN(new_n2250_));
  AOI21_X1   g02058(.A1(new_n2237_), .A2(new_n2250_), .B(new_n744_), .ZN(new_n2251_));
  NOR3_X1    g02059(.A1(new_n2236_), .A2(\asqrt[56] ), .A3(new_n2251_), .ZN(new_n2252_));
  OAI21_X1   g02060(.A1(new_n2236_), .A2(new_n2251_), .B(\asqrt[56] ), .ZN(new_n2253_));
  OAI21_X1   g02061(.A1(new_n2152_), .A2(new_n2252_), .B(new_n2253_), .ZN(new_n2254_));
  OAI21_X1   g02062(.A1(new_n2254_), .A2(\asqrt[57] ), .B(new_n2149_), .ZN(new_n2255_));
  NAND2_X1   g02063(.A1(new_n2254_), .A2(\asqrt[57] ), .ZN(new_n2256_));
  NAND3_X1   g02064(.A1(new_n2255_), .A2(new_n2256_), .A3(new_n423_), .ZN(new_n2257_));
  AOI21_X1   g02065(.A1(new_n2255_), .A2(new_n2256_), .B(new_n423_), .ZN(new_n2258_));
  AOI21_X1   g02066(.A1(new_n2146_), .A2(new_n2257_), .B(new_n2258_), .ZN(new_n2259_));
  AOI21_X1   g02067(.A1(new_n2259_), .A2(new_n337_), .B(new_n2143_), .ZN(new_n2260_));
  NAND2_X1   g02068(.A1(new_n2257_), .A2(new_n2146_), .ZN(new_n2261_));
  INV_X1     g02069(.I(new_n2149_), .ZN(new_n2262_));
  INV_X1     g02070(.I(new_n2158_), .ZN(new_n2263_));
  NOR3_X1    g02071(.A1(new_n2247_), .A2(\asqrt[54] ), .A3(new_n2249_), .ZN(new_n2264_));
  OAI21_X1   g02072(.A1(new_n2263_), .A2(new_n2264_), .B(new_n2250_), .ZN(new_n2265_));
  OAI21_X1   g02073(.A1(new_n2265_), .A2(\asqrt[55] ), .B(new_n2154_), .ZN(new_n2266_));
  NAND2_X1   g02074(.A1(new_n2265_), .A2(\asqrt[55] ), .ZN(new_n2267_));
  NAND3_X1   g02075(.A1(new_n2266_), .A2(new_n2267_), .A3(new_n634_), .ZN(new_n2268_));
  AOI21_X1   g02076(.A1(new_n2266_), .A2(new_n2267_), .B(new_n634_), .ZN(new_n2269_));
  AOI21_X1   g02077(.A1(new_n2151_), .A2(new_n2268_), .B(new_n2269_), .ZN(new_n2270_));
  AOI21_X1   g02078(.A1(new_n2270_), .A2(new_n531_), .B(new_n2262_), .ZN(new_n2271_));
  NAND2_X1   g02079(.A1(new_n2268_), .A2(new_n2151_), .ZN(new_n2272_));
  AOI21_X1   g02080(.A1(new_n2272_), .A2(new_n2253_), .B(new_n531_), .ZN(new_n2273_));
  OAI21_X1   g02081(.A1(new_n2271_), .A2(new_n2273_), .B(\asqrt[58] ), .ZN(new_n2274_));
  AOI21_X1   g02082(.A1(new_n2261_), .A2(new_n2274_), .B(new_n337_), .ZN(new_n2275_));
  NOR3_X1    g02083(.A1(new_n2260_), .A2(\asqrt[60] ), .A3(new_n2275_), .ZN(new_n2276_));
  NOR2_X1    g02084(.A1(new_n2276_), .A2(new_n2140_), .ZN(new_n2277_));
  INV_X1     g02085(.I(new_n2146_), .ZN(new_n2278_));
  NOR3_X1    g02086(.A1(new_n2271_), .A2(\asqrt[58] ), .A3(new_n2273_), .ZN(new_n2279_));
  OAI21_X1   g02087(.A1(new_n2278_), .A2(new_n2279_), .B(new_n2274_), .ZN(new_n2280_));
  OAI21_X1   g02088(.A1(new_n2280_), .A2(\asqrt[59] ), .B(new_n2142_), .ZN(new_n2281_));
  NOR2_X1    g02089(.A1(new_n2279_), .A2(new_n2278_), .ZN(new_n2282_));
  OAI21_X1   g02090(.A1(new_n2282_), .A2(new_n2258_), .B(\asqrt[59] ), .ZN(new_n2283_));
  AOI21_X1   g02091(.A1(new_n2281_), .A2(new_n2283_), .B(new_n266_), .ZN(new_n2284_));
  OAI21_X1   g02092(.A1(new_n2277_), .A2(new_n2284_), .B(\asqrt[61] ), .ZN(new_n2285_));
  OAI21_X1   g02093(.A1(new_n2260_), .A2(new_n2275_), .B(\asqrt[60] ), .ZN(new_n2286_));
  OAI21_X1   g02094(.A1(new_n2140_), .A2(new_n2276_), .B(new_n2286_), .ZN(new_n2287_));
  AOI21_X1   g02095(.A1(new_n2095_), .A2(new_n2075_), .B(\asqrt[46] ), .ZN(new_n2288_));
  XOR2_X1    g02096(.A1(new_n2288_), .A2(new_n1959_), .Z(new_n2289_));
  OAI21_X1   g02097(.A1(new_n2287_), .A2(\asqrt[61] ), .B(new_n2289_), .ZN(new_n2290_));
  NAND2_X1   g02098(.A1(new_n2290_), .A2(new_n2285_), .ZN(new_n2291_));
  NAND3_X1   g02099(.A1(new_n2281_), .A2(new_n266_), .A3(new_n2283_), .ZN(new_n2292_));
  NAND2_X1   g02100(.A1(new_n2292_), .A2(new_n2139_), .ZN(new_n2293_));
  AOI21_X1   g02101(.A1(new_n2293_), .A2(new_n2286_), .B(new_n239_), .ZN(new_n2294_));
  AOI21_X1   g02102(.A1(new_n2139_), .A2(new_n2292_), .B(new_n2284_), .ZN(new_n2295_));
  INV_X1     g02103(.I(new_n2289_), .ZN(new_n2296_));
  AOI21_X1   g02104(.A1(new_n2295_), .A2(new_n239_), .B(new_n2296_), .ZN(new_n2297_));
  OAI21_X1   g02105(.A1(new_n2297_), .A2(new_n2294_), .B(new_n201_), .ZN(new_n2298_));
  NAND3_X1   g02106(.A1(new_n2290_), .A2(\asqrt[62] ), .A3(new_n2285_), .ZN(new_n2299_));
  NAND2_X1   g02107(.A1(new_n2099_), .A2(new_n239_), .ZN(new_n2300_));
  AOI21_X1   g02108(.A1(new_n2077_), .A2(new_n2300_), .B(\asqrt[46] ), .ZN(new_n2301_));
  XOR2_X1    g02109(.A1(new_n2301_), .A2(new_n2079_), .Z(new_n2302_));
  INV_X1     g02110(.I(new_n2302_), .ZN(new_n2303_));
  AOI22_X1   g02111(.A1(new_n2298_), .A2(new_n2299_), .B1(new_n2291_), .B2(new_n2303_), .ZN(new_n2304_));
  NOR2_X1    g02112(.A1(new_n2108_), .A2(new_n1956_), .ZN(new_n2305_));
  OAI21_X1   g02113(.A1(\asqrt[46] ), .A2(new_n2305_), .B(new_n2115_), .ZN(new_n2306_));
  INV_X1     g02114(.I(new_n2306_), .ZN(new_n2307_));
  OAI21_X1   g02115(.A1(new_n2304_), .A2(new_n2137_), .B(new_n2307_), .ZN(new_n2308_));
  OAI21_X1   g02116(.A1(new_n2291_), .A2(\asqrt[62] ), .B(new_n2302_), .ZN(new_n2309_));
  NAND2_X1   g02117(.A1(new_n2291_), .A2(\asqrt[62] ), .ZN(new_n2310_));
  NAND3_X1   g02118(.A1(new_n2309_), .A2(new_n2310_), .A3(new_n2137_), .ZN(new_n2311_));
  NAND2_X1   g02119(.A1(new_n2134_), .A2(new_n1955_), .ZN(new_n2312_));
  XOR2_X1    g02120(.A1(new_n2130_), .A2(new_n1955_), .Z(new_n2313_));
  NAND3_X1   g02121(.A1(new_n2312_), .A2(\asqrt[63] ), .A3(new_n2313_), .ZN(new_n2314_));
  INV_X1     g02122(.I(new_n2180_), .ZN(new_n2315_));
  NAND4_X1   g02123(.A1(new_n2315_), .A2(new_n1956_), .A3(new_n2115_), .A4(new_n2122_), .ZN(new_n2316_));
  NAND2_X1   g02124(.A1(new_n2314_), .A2(new_n2316_), .ZN(new_n2317_));
  INV_X1     g02125(.I(new_n2317_), .ZN(new_n2318_));
  NAND4_X1   g02126(.A1(new_n2308_), .A2(new_n193_), .A3(new_n2311_), .A4(new_n2318_), .ZN(\asqrt[45] ));
  NOR2_X1    g02127(.A1(new_n2291_), .A2(\asqrt[62] ), .ZN(new_n2320_));
  INV_X1     g02128(.I(new_n2310_), .ZN(new_n2321_));
  NOR2_X1    g02129(.A1(new_n2321_), .A2(new_n2320_), .ZN(new_n2322_));
  NAND3_X1   g02130(.A1(new_n2293_), .A2(new_n239_), .A3(new_n2286_), .ZN(new_n2323_));
  AOI21_X1   g02131(.A1(new_n2289_), .A2(new_n2323_), .B(new_n2294_), .ZN(new_n2324_));
  AOI21_X1   g02132(.A1(new_n2290_), .A2(new_n2285_), .B(\asqrt[62] ), .ZN(new_n2325_));
  NOR3_X1    g02133(.A1(new_n2297_), .A2(new_n201_), .A3(new_n2294_), .ZN(new_n2326_));
  OAI22_X1   g02134(.A1(new_n2326_), .A2(new_n2325_), .B1(new_n2324_), .B2(new_n2302_), .ZN(new_n2327_));
  AOI21_X1   g02135(.A1(new_n2327_), .A2(new_n2136_), .B(new_n2306_), .ZN(new_n2328_));
  AOI21_X1   g02136(.A1(new_n2324_), .A2(new_n201_), .B(new_n2303_), .ZN(new_n2329_));
  OAI21_X1   g02137(.A1(new_n2324_), .A2(new_n201_), .B(new_n2137_), .ZN(new_n2330_));
  NOR2_X1    g02138(.A1(new_n2329_), .A2(new_n2330_), .ZN(new_n2331_));
  NOR4_X1    g02139(.A1(new_n2328_), .A2(\asqrt[63] ), .A3(new_n2331_), .A4(new_n2317_), .ZN(new_n2332_));
  XOR2_X1    g02140(.A1(new_n2301_), .A2(new_n2079_), .Z(new_n2333_));
  OAI21_X1   g02141(.A1(\asqrt[45] ), .A2(new_n2322_), .B(new_n2333_), .ZN(new_n2334_));
  INV_X1     g02142(.I(new_n2334_), .ZN(new_n2335_));
  NAND2_X1   g02143(.A1(new_n2259_), .A2(new_n337_), .ZN(new_n2336_));
  AOI21_X1   g02144(.A1(new_n2336_), .A2(new_n2283_), .B(\asqrt[45] ), .ZN(new_n2337_));
  XOR2_X1    g02145(.A1(new_n2337_), .A2(new_n2142_), .Z(new_n2338_));
  INV_X1     g02146(.I(new_n2338_), .ZN(new_n2339_));
  AOI21_X1   g02147(.A1(new_n2257_), .A2(new_n2274_), .B(\asqrt[45] ), .ZN(new_n2340_));
  XOR2_X1    g02148(.A1(new_n2340_), .A2(new_n2146_), .Z(new_n2341_));
  INV_X1     g02149(.I(new_n2341_), .ZN(new_n2342_));
  NAND2_X1   g02150(.A1(new_n2270_), .A2(new_n531_), .ZN(new_n2343_));
  AOI21_X1   g02151(.A1(new_n2343_), .A2(new_n2256_), .B(\asqrt[45] ), .ZN(new_n2344_));
  XOR2_X1    g02152(.A1(new_n2344_), .A2(new_n2149_), .Z(new_n2345_));
  INV_X1     g02153(.I(new_n2345_), .ZN(new_n2346_));
  AOI21_X1   g02154(.A1(new_n2268_), .A2(new_n2253_), .B(\asqrt[45] ), .ZN(new_n2347_));
  XOR2_X1    g02155(.A1(new_n2347_), .A2(new_n2151_), .Z(new_n2348_));
  NAND2_X1   g02156(.A1(new_n2235_), .A2(new_n744_), .ZN(new_n2349_));
  AOI21_X1   g02157(.A1(new_n2349_), .A2(new_n2267_), .B(\asqrt[45] ), .ZN(new_n2350_));
  XOR2_X1    g02158(.A1(new_n2350_), .A2(new_n2154_), .Z(new_n2351_));
  AOI21_X1   g02159(.A1(new_n2233_), .A2(new_n2250_), .B(\asqrt[45] ), .ZN(new_n2352_));
  XOR2_X1    g02160(.A1(new_n2352_), .A2(new_n2158_), .Z(new_n2353_));
  INV_X1     g02161(.I(new_n2353_), .ZN(new_n2354_));
  NAND2_X1   g02162(.A1(new_n2246_), .A2(new_n1006_), .ZN(new_n2355_));
  AOI21_X1   g02163(.A1(new_n2355_), .A2(new_n2232_), .B(\asqrt[45] ), .ZN(new_n2356_));
  XOR2_X1    g02164(.A1(new_n2356_), .A2(new_n2161_), .Z(new_n2357_));
  INV_X1     g02165(.I(new_n2357_), .ZN(new_n2358_));
  AOI21_X1   g02166(.A1(new_n2244_), .A2(new_n2229_), .B(\asqrt[45] ), .ZN(new_n2359_));
  XOR2_X1    g02167(.A1(new_n2359_), .A2(new_n2163_), .Z(new_n2360_));
  NAND2_X1   g02168(.A1(new_n2207_), .A2(new_n1305_), .ZN(new_n2361_));
  AOI21_X1   g02169(.A1(new_n2361_), .A2(new_n2243_), .B(\asqrt[45] ), .ZN(new_n2362_));
  XOR2_X1    g02170(.A1(new_n2362_), .A2(new_n2166_), .Z(new_n2363_));
  AOI21_X1   g02171(.A1(new_n2205_), .A2(new_n2226_), .B(\asqrt[45] ), .ZN(new_n2364_));
  XOR2_X1    g02172(.A1(new_n2364_), .A2(new_n2169_), .Z(new_n2365_));
  INV_X1     g02173(.I(new_n2365_), .ZN(new_n2366_));
  NAND2_X1   g02174(.A1(new_n2222_), .A2(new_n1632_), .ZN(new_n2367_));
  AOI21_X1   g02175(.A1(new_n2367_), .A2(new_n2204_), .B(\asqrt[45] ), .ZN(new_n2368_));
  XOR2_X1    g02176(.A1(new_n2368_), .A2(new_n2175_), .Z(new_n2369_));
  INV_X1     g02177(.I(new_n2369_), .ZN(new_n2370_));
  AOI21_X1   g02178(.A1(new_n2220_), .A2(new_n2201_), .B(\asqrt[45] ), .ZN(new_n2371_));
  XOR2_X1    g02179(.A1(new_n2371_), .A2(new_n2211_), .Z(new_n2372_));
  NAND2_X1   g02180(.A1(\asqrt[46] ), .A2(new_n2189_), .ZN(new_n2373_));
  NOR2_X1    g02181(.A1(new_n2196_), .A2(\a[92] ), .ZN(new_n2374_));
  AOI22_X1   g02182(.A1(new_n2373_), .A2(new_n2196_), .B1(\asqrt[46] ), .B2(new_n2374_), .ZN(new_n2375_));
  AOI21_X1   g02183(.A1(\asqrt[46] ), .A2(\a[92] ), .B(new_n2194_), .ZN(new_n2376_));
  OAI21_X1   g02184(.A1(new_n2191_), .A2(new_n2376_), .B(new_n2332_), .ZN(new_n2377_));
  XNOR2_X1   g02185(.A1(new_n2377_), .A2(new_n2375_), .ZN(new_n2378_));
  NOR3_X1    g02186(.A1(new_n2328_), .A2(\asqrt[63] ), .A3(new_n2331_), .ZN(new_n2379_));
  NAND3_X1   g02187(.A1(new_n2314_), .A2(\asqrt[46] ), .A3(new_n2316_), .ZN(new_n2380_));
  INV_X1     g02188(.I(new_n2380_), .ZN(new_n2381_));
  NAND2_X1   g02189(.A1(new_n2379_), .A2(new_n2381_), .ZN(new_n2382_));
  NAND2_X1   g02190(.A1(\asqrt[45] ), .A2(new_n2186_), .ZN(new_n2383_));
  AOI21_X1   g02191(.A1(new_n2383_), .A2(new_n2382_), .B(\a[92] ), .ZN(new_n2384_));
  NAND2_X1   g02192(.A1(new_n2308_), .A2(new_n193_), .ZN(new_n2385_));
  NOR3_X1    g02193(.A1(new_n2385_), .A2(new_n2331_), .A3(new_n2380_), .ZN(new_n2386_));
  NOR2_X1    g02194(.A1(new_n2332_), .A2(new_n2187_), .ZN(new_n2387_));
  NOR3_X1    g02195(.A1(new_n2387_), .A2(new_n2386_), .A3(new_n2189_), .ZN(new_n2388_));
  OR2_X2     g02196(.A1(new_n2388_), .A2(new_n2384_), .Z(new_n2389_));
  NOR2_X1    g02197(.A1(\a[88] ), .A2(\a[89] ), .ZN(new_n2390_));
  INV_X1     g02198(.I(new_n2390_), .ZN(new_n2391_));
  NAND3_X1   g02199(.A1(\asqrt[45] ), .A2(\a[90] ), .A3(new_n2391_), .ZN(new_n2392_));
  INV_X1     g02200(.I(\a[90] ), .ZN(new_n2393_));
  OAI21_X1   g02201(.A1(\asqrt[45] ), .A2(new_n2393_), .B(new_n2390_), .ZN(new_n2394_));
  AOI21_X1   g02202(.A1(new_n2394_), .A2(new_n2392_), .B(new_n2134_), .ZN(new_n2395_));
  NAND2_X1   g02203(.A1(new_n2390_), .A2(new_n2393_), .ZN(new_n2396_));
  NAND3_X1   g02204(.A1(new_n2118_), .A2(new_n2120_), .A3(new_n2396_), .ZN(new_n2397_));
  NAND2_X1   g02205(.A1(new_n2176_), .A2(new_n2397_), .ZN(new_n2398_));
  NAND3_X1   g02206(.A1(\asqrt[45] ), .A2(\a[90] ), .A3(new_n2398_), .ZN(new_n2399_));
  INV_X1     g02207(.I(\a[91] ), .ZN(new_n2400_));
  NAND3_X1   g02208(.A1(\asqrt[45] ), .A2(new_n2393_), .A3(new_n2400_), .ZN(new_n2401_));
  OAI21_X1   g02209(.A1(new_n2332_), .A2(\a[90] ), .B(\a[91] ), .ZN(new_n2402_));
  NAND3_X1   g02210(.A1(new_n2399_), .A2(new_n2402_), .A3(new_n2401_), .ZN(new_n2403_));
  NOR3_X1    g02211(.A1(new_n2403_), .A2(new_n2395_), .A3(\asqrt[47] ), .ZN(new_n2404_));
  OAI21_X1   g02212(.A1(new_n2403_), .A2(new_n2395_), .B(\asqrt[47] ), .ZN(new_n2405_));
  OAI21_X1   g02213(.A1(new_n2389_), .A2(new_n2404_), .B(new_n2405_), .ZN(new_n2406_));
  OAI21_X1   g02214(.A1(new_n2406_), .A2(\asqrt[48] ), .B(new_n2378_), .ZN(new_n2407_));
  NAND2_X1   g02215(.A1(new_n2406_), .A2(\asqrt[48] ), .ZN(new_n2408_));
  NAND3_X1   g02216(.A1(new_n2407_), .A2(new_n2408_), .A3(new_n1632_), .ZN(new_n2409_));
  AOI21_X1   g02217(.A1(new_n2407_), .A2(new_n2408_), .B(new_n1632_), .ZN(new_n2410_));
  AOI21_X1   g02218(.A1(new_n2372_), .A2(new_n2409_), .B(new_n2410_), .ZN(new_n2411_));
  AOI21_X1   g02219(.A1(new_n2411_), .A2(new_n1463_), .B(new_n2370_), .ZN(new_n2412_));
  NAND2_X1   g02220(.A1(new_n2409_), .A2(new_n2372_), .ZN(new_n2413_));
  INV_X1     g02221(.I(new_n2410_), .ZN(new_n2414_));
  AOI21_X1   g02222(.A1(new_n2413_), .A2(new_n2414_), .B(new_n1463_), .ZN(new_n2415_));
  NOR3_X1    g02223(.A1(new_n2412_), .A2(\asqrt[51] ), .A3(new_n2415_), .ZN(new_n2416_));
  OAI21_X1   g02224(.A1(new_n2412_), .A2(new_n2415_), .B(\asqrt[51] ), .ZN(new_n2417_));
  OAI21_X1   g02225(.A1(new_n2366_), .A2(new_n2416_), .B(new_n2417_), .ZN(new_n2418_));
  OAI21_X1   g02226(.A1(new_n2418_), .A2(\asqrt[52] ), .B(new_n2363_), .ZN(new_n2419_));
  NAND2_X1   g02227(.A1(new_n2418_), .A2(\asqrt[52] ), .ZN(new_n2420_));
  NAND3_X1   g02228(.A1(new_n2419_), .A2(new_n2420_), .A3(new_n1006_), .ZN(new_n2421_));
  AOI21_X1   g02229(.A1(new_n2419_), .A2(new_n2420_), .B(new_n1006_), .ZN(new_n2422_));
  AOI21_X1   g02230(.A1(new_n2360_), .A2(new_n2421_), .B(new_n2422_), .ZN(new_n2423_));
  AOI21_X1   g02231(.A1(new_n2423_), .A2(new_n860_), .B(new_n2358_), .ZN(new_n2424_));
  NAND2_X1   g02232(.A1(new_n2421_), .A2(new_n2360_), .ZN(new_n2425_));
  INV_X1     g02233(.I(new_n2422_), .ZN(new_n2426_));
  AOI21_X1   g02234(.A1(new_n2425_), .A2(new_n2426_), .B(new_n860_), .ZN(new_n2427_));
  NOR3_X1    g02235(.A1(new_n2424_), .A2(\asqrt[55] ), .A3(new_n2427_), .ZN(new_n2428_));
  OAI21_X1   g02236(.A1(new_n2424_), .A2(new_n2427_), .B(\asqrt[55] ), .ZN(new_n2429_));
  OAI21_X1   g02237(.A1(new_n2354_), .A2(new_n2428_), .B(new_n2429_), .ZN(new_n2430_));
  OAI21_X1   g02238(.A1(new_n2430_), .A2(\asqrt[56] ), .B(new_n2351_), .ZN(new_n2431_));
  NAND2_X1   g02239(.A1(new_n2430_), .A2(\asqrt[56] ), .ZN(new_n2432_));
  NAND3_X1   g02240(.A1(new_n2431_), .A2(new_n2432_), .A3(new_n531_), .ZN(new_n2433_));
  AOI21_X1   g02241(.A1(new_n2431_), .A2(new_n2432_), .B(new_n531_), .ZN(new_n2434_));
  AOI21_X1   g02242(.A1(new_n2348_), .A2(new_n2433_), .B(new_n2434_), .ZN(new_n2435_));
  AOI21_X1   g02243(.A1(new_n2435_), .A2(new_n423_), .B(new_n2346_), .ZN(new_n2436_));
  NAND2_X1   g02244(.A1(new_n2433_), .A2(new_n2348_), .ZN(new_n2437_));
  INV_X1     g02245(.I(new_n2434_), .ZN(new_n2438_));
  AOI21_X1   g02246(.A1(new_n2437_), .A2(new_n2438_), .B(new_n423_), .ZN(new_n2439_));
  NOR3_X1    g02247(.A1(new_n2436_), .A2(\asqrt[59] ), .A3(new_n2439_), .ZN(new_n2440_));
  NOR2_X1    g02248(.A1(new_n2440_), .A2(new_n2342_), .ZN(new_n2441_));
  OAI21_X1   g02249(.A1(new_n2436_), .A2(new_n2439_), .B(\asqrt[59] ), .ZN(new_n2442_));
  INV_X1     g02250(.I(new_n2442_), .ZN(new_n2443_));
  NOR2_X1    g02251(.A1(new_n2441_), .A2(new_n2443_), .ZN(new_n2444_));
  AOI21_X1   g02252(.A1(new_n2444_), .A2(new_n266_), .B(new_n2339_), .ZN(new_n2445_));
  INV_X1     g02253(.I(new_n2348_), .ZN(new_n2446_));
  INV_X1     g02254(.I(new_n2360_), .ZN(new_n2447_));
  INV_X1     g02255(.I(new_n2372_), .ZN(new_n2448_));
  NOR2_X1    g02256(.A1(new_n2388_), .A2(new_n2384_), .ZN(new_n2449_));
  NOR3_X1    g02257(.A1(new_n2332_), .A2(new_n2393_), .A3(new_n2390_), .ZN(new_n2450_));
  AOI21_X1   g02258(.A1(new_n2332_), .A2(\a[90] ), .B(new_n2391_), .ZN(new_n2451_));
  OAI21_X1   g02259(.A1(new_n2450_), .A2(new_n2451_), .B(\asqrt[46] ), .ZN(new_n2452_));
  INV_X1     g02260(.I(new_n2398_), .ZN(new_n2453_));
  NOR3_X1    g02261(.A1(new_n2332_), .A2(new_n2393_), .A3(new_n2453_), .ZN(new_n2454_));
  NOR3_X1    g02262(.A1(new_n2332_), .A2(\a[90] ), .A3(\a[91] ), .ZN(new_n2455_));
  AOI21_X1   g02263(.A1(\asqrt[45] ), .A2(new_n2393_), .B(new_n2400_), .ZN(new_n2456_));
  NOR3_X1    g02264(.A1(new_n2454_), .A2(new_n2455_), .A3(new_n2456_), .ZN(new_n2457_));
  NAND3_X1   g02265(.A1(new_n2457_), .A2(new_n2452_), .A3(new_n1953_), .ZN(new_n2458_));
  NAND2_X1   g02266(.A1(new_n2458_), .A2(new_n2449_), .ZN(new_n2459_));
  NAND3_X1   g02267(.A1(new_n2459_), .A2(new_n1778_), .A3(new_n2405_), .ZN(new_n2460_));
  AOI21_X1   g02268(.A1(new_n2459_), .A2(new_n2405_), .B(new_n1778_), .ZN(new_n2461_));
  AOI21_X1   g02269(.A1(new_n2378_), .A2(new_n2460_), .B(new_n2461_), .ZN(new_n2462_));
  AOI21_X1   g02270(.A1(new_n2462_), .A2(new_n1632_), .B(new_n2448_), .ZN(new_n2463_));
  NOR3_X1    g02271(.A1(new_n2463_), .A2(\asqrt[50] ), .A3(new_n2410_), .ZN(new_n2464_));
  OAI21_X1   g02272(.A1(new_n2463_), .A2(new_n2410_), .B(\asqrt[50] ), .ZN(new_n2465_));
  OAI21_X1   g02273(.A1(new_n2370_), .A2(new_n2464_), .B(new_n2465_), .ZN(new_n2466_));
  OAI21_X1   g02274(.A1(new_n2466_), .A2(\asqrt[51] ), .B(new_n2365_), .ZN(new_n2467_));
  NAND3_X1   g02275(.A1(new_n2467_), .A2(new_n1150_), .A3(new_n2417_), .ZN(new_n2468_));
  AOI21_X1   g02276(.A1(new_n2467_), .A2(new_n2417_), .B(new_n1150_), .ZN(new_n2469_));
  AOI21_X1   g02277(.A1(new_n2363_), .A2(new_n2468_), .B(new_n2469_), .ZN(new_n2470_));
  AOI21_X1   g02278(.A1(new_n2470_), .A2(new_n1006_), .B(new_n2447_), .ZN(new_n2471_));
  NOR3_X1    g02279(.A1(new_n2471_), .A2(\asqrt[54] ), .A3(new_n2422_), .ZN(new_n2472_));
  OAI21_X1   g02280(.A1(new_n2471_), .A2(new_n2422_), .B(\asqrt[54] ), .ZN(new_n2473_));
  OAI21_X1   g02281(.A1(new_n2358_), .A2(new_n2472_), .B(new_n2473_), .ZN(new_n2474_));
  OAI21_X1   g02282(.A1(new_n2474_), .A2(\asqrt[55] ), .B(new_n2353_), .ZN(new_n2475_));
  NAND3_X1   g02283(.A1(new_n2475_), .A2(new_n634_), .A3(new_n2429_), .ZN(new_n2476_));
  AOI21_X1   g02284(.A1(new_n2475_), .A2(new_n2429_), .B(new_n634_), .ZN(new_n2477_));
  AOI21_X1   g02285(.A1(new_n2351_), .A2(new_n2476_), .B(new_n2477_), .ZN(new_n2478_));
  AOI21_X1   g02286(.A1(new_n2478_), .A2(new_n531_), .B(new_n2446_), .ZN(new_n2479_));
  NOR3_X1    g02287(.A1(new_n2479_), .A2(\asqrt[58] ), .A3(new_n2434_), .ZN(new_n2480_));
  OAI21_X1   g02288(.A1(new_n2479_), .A2(new_n2434_), .B(\asqrt[58] ), .ZN(new_n2481_));
  OAI21_X1   g02289(.A1(new_n2346_), .A2(new_n2480_), .B(new_n2481_), .ZN(new_n2482_));
  OAI21_X1   g02290(.A1(new_n2482_), .A2(\asqrt[59] ), .B(new_n2341_), .ZN(new_n2483_));
  AOI21_X1   g02291(.A1(new_n2483_), .A2(new_n2442_), .B(new_n266_), .ZN(new_n2484_));
  OAI21_X1   g02292(.A1(new_n2445_), .A2(new_n2484_), .B(\asqrt[61] ), .ZN(new_n2485_));
  AOI21_X1   g02293(.A1(new_n2292_), .A2(new_n2286_), .B(\asqrt[45] ), .ZN(new_n2486_));
  XOR2_X1    g02294(.A1(new_n2486_), .A2(new_n2139_), .Z(new_n2487_));
  OAI21_X1   g02295(.A1(new_n2342_), .A2(new_n2440_), .B(new_n2442_), .ZN(new_n2488_));
  OAI21_X1   g02296(.A1(new_n2488_), .A2(\asqrt[60] ), .B(new_n2338_), .ZN(new_n2489_));
  OAI21_X1   g02297(.A1(new_n2441_), .A2(new_n2443_), .B(\asqrt[60] ), .ZN(new_n2490_));
  NAND3_X1   g02298(.A1(new_n2489_), .A2(new_n239_), .A3(new_n2490_), .ZN(new_n2491_));
  NAND2_X1   g02299(.A1(new_n2491_), .A2(new_n2487_), .ZN(new_n2492_));
  NAND2_X1   g02300(.A1(new_n2492_), .A2(new_n2485_), .ZN(new_n2493_));
  AOI21_X1   g02301(.A1(new_n2489_), .A2(new_n2490_), .B(new_n239_), .ZN(new_n2494_));
  NAND3_X1   g02302(.A1(new_n2483_), .A2(new_n266_), .A3(new_n2442_), .ZN(new_n2495_));
  AOI21_X1   g02303(.A1(new_n2338_), .A2(new_n2495_), .B(new_n2484_), .ZN(new_n2496_));
  INV_X1     g02304(.I(new_n2487_), .ZN(new_n2497_));
  AOI21_X1   g02305(.A1(new_n2496_), .A2(new_n239_), .B(new_n2497_), .ZN(new_n2498_));
  OAI21_X1   g02306(.A1(new_n2498_), .A2(new_n2494_), .B(new_n201_), .ZN(new_n2499_));
  NAND3_X1   g02307(.A1(new_n2492_), .A2(\asqrt[62] ), .A3(new_n2485_), .ZN(new_n2500_));
  AOI21_X1   g02308(.A1(new_n2285_), .A2(new_n2323_), .B(\asqrt[45] ), .ZN(new_n2501_));
  XOR2_X1    g02309(.A1(new_n2501_), .A2(new_n2289_), .Z(new_n2502_));
  INV_X1     g02310(.I(new_n2502_), .ZN(new_n2503_));
  AOI22_X1   g02311(.A1(new_n2499_), .A2(new_n2500_), .B1(new_n2493_), .B2(new_n2503_), .ZN(new_n2504_));
  NOR2_X1    g02312(.A1(new_n2304_), .A2(new_n2137_), .ZN(new_n2505_));
  OAI21_X1   g02313(.A1(\asqrt[45] ), .A2(new_n2505_), .B(new_n2311_), .ZN(new_n2506_));
  INV_X1     g02314(.I(new_n2506_), .ZN(new_n2507_));
  OAI21_X1   g02315(.A1(new_n2504_), .A2(new_n2335_), .B(new_n2507_), .ZN(new_n2508_));
  OAI21_X1   g02316(.A1(new_n2493_), .A2(\asqrt[62] ), .B(new_n2502_), .ZN(new_n2509_));
  NAND2_X1   g02317(.A1(new_n2493_), .A2(\asqrt[62] ), .ZN(new_n2510_));
  NAND3_X1   g02318(.A1(new_n2509_), .A2(new_n2510_), .A3(new_n2335_), .ZN(new_n2511_));
  NAND2_X1   g02319(.A1(new_n2332_), .A2(new_n2136_), .ZN(new_n2512_));
  XOR2_X1    g02320(.A1(new_n2304_), .A2(new_n2137_), .Z(new_n2513_));
  NAND3_X1   g02321(.A1(new_n2512_), .A2(\asqrt[63] ), .A3(new_n2513_), .ZN(new_n2514_));
  INV_X1     g02322(.I(new_n2385_), .ZN(new_n2515_));
  NAND4_X1   g02323(.A1(new_n2515_), .A2(new_n2137_), .A3(new_n2311_), .A4(new_n2318_), .ZN(new_n2516_));
  NAND2_X1   g02324(.A1(new_n2514_), .A2(new_n2516_), .ZN(new_n2517_));
  INV_X1     g02325(.I(new_n2517_), .ZN(new_n2518_));
  NAND4_X1   g02326(.A1(new_n2508_), .A2(new_n193_), .A3(new_n2511_), .A4(new_n2518_), .ZN(\asqrt[44] ));
  NOR2_X1    g02327(.A1(new_n2493_), .A2(\asqrt[62] ), .ZN(new_n2520_));
  INV_X1     g02328(.I(new_n2510_), .ZN(new_n2521_));
  NOR2_X1    g02329(.A1(new_n2521_), .A2(new_n2520_), .ZN(new_n2522_));
  NOR2_X1    g02330(.A1(new_n2498_), .A2(new_n2494_), .ZN(new_n2523_));
  AOI21_X1   g02331(.A1(new_n2492_), .A2(new_n2485_), .B(\asqrt[62] ), .ZN(new_n2524_));
  NOR3_X1    g02332(.A1(new_n2498_), .A2(new_n201_), .A3(new_n2494_), .ZN(new_n2525_));
  OAI22_X1   g02333(.A1(new_n2525_), .A2(new_n2524_), .B1(new_n2523_), .B2(new_n2502_), .ZN(new_n2526_));
  AOI21_X1   g02334(.A1(new_n2526_), .A2(new_n2334_), .B(new_n2506_), .ZN(new_n2527_));
  AOI21_X1   g02335(.A1(new_n2523_), .A2(new_n201_), .B(new_n2503_), .ZN(new_n2528_));
  OAI21_X1   g02336(.A1(new_n2523_), .A2(new_n201_), .B(new_n2335_), .ZN(new_n2529_));
  NOR2_X1    g02337(.A1(new_n2528_), .A2(new_n2529_), .ZN(new_n2530_));
  NOR4_X1    g02338(.A1(new_n2527_), .A2(\asqrt[63] ), .A3(new_n2530_), .A4(new_n2517_), .ZN(new_n2531_));
  XOR2_X1    g02339(.A1(new_n2501_), .A2(new_n2289_), .Z(new_n2532_));
  OAI21_X1   g02340(.A1(\asqrt[44] ), .A2(new_n2522_), .B(new_n2532_), .ZN(new_n2533_));
  INV_X1     g02341(.I(new_n2533_), .ZN(new_n2534_));
  NOR2_X1    g02342(.A1(new_n2443_), .A2(new_n2440_), .ZN(new_n2535_));
  NOR2_X1    g02343(.A1(\asqrt[44] ), .A2(new_n2535_), .ZN(new_n2536_));
  XOR2_X1    g02344(.A1(new_n2536_), .A2(new_n2341_), .Z(new_n2537_));
  INV_X1     g02345(.I(new_n2537_), .ZN(new_n2538_));
  NOR2_X1    g02346(.A1(new_n2480_), .A2(new_n2439_), .ZN(new_n2539_));
  NOR2_X1    g02347(.A1(\asqrt[44] ), .A2(new_n2539_), .ZN(new_n2540_));
  XOR2_X1    g02348(.A1(new_n2540_), .A2(new_n2345_), .Z(new_n2541_));
  AOI21_X1   g02349(.A1(new_n2433_), .A2(new_n2438_), .B(\asqrt[44] ), .ZN(new_n2542_));
  XOR2_X1    g02350(.A1(new_n2542_), .A2(new_n2348_), .Z(new_n2543_));
  AOI21_X1   g02351(.A1(new_n2476_), .A2(new_n2432_), .B(\asqrt[44] ), .ZN(new_n2544_));
  XOR2_X1    g02352(.A1(new_n2544_), .A2(new_n2351_), .Z(new_n2545_));
  INV_X1     g02353(.I(new_n2429_), .ZN(new_n2546_));
  NOR2_X1    g02354(.A1(new_n2546_), .A2(new_n2428_), .ZN(new_n2547_));
  NOR2_X1    g02355(.A1(\asqrt[44] ), .A2(new_n2547_), .ZN(new_n2548_));
  XOR2_X1    g02356(.A1(new_n2548_), .A2(new_n2353_), .Z(new_n2549_));
  INV_X1     g02357(.I(new_n2549_), .ZN(new_n2550_));
  NOR2_X1    g02358(.A1(new_n2472_), .A2(new_n2427_), .ZN(new_n2551_));
  NOR2_X1    g02359(.A1(\asqrt[44] ), .A2(new_n2551_), .ZN(new_n2552_));
  XOR2_X1    g02360(.A1(new_n2552_), .A2(new_n2357_), .Z(new_n2553_));
  INV_X1     g02361(.I(new_n2553_), .ZN(new_n2554_));
  AOI21_X1   g02362(.A1(new_n2421_), .A2(new_n2426_), .B(\asqrt[44] ), .ZN(new_n2555_));
  XOR2_X1    g02363(.A1(new_n2555_), .A2(new_n2360_), .Z(new_n2556_));
  AOI21_X1   g02364(.A1(new_n2468_), .A2(new_n2420_), .B(\asqrt[44] ), .ZN(new_n2557_));
  XOR2_X1    g02365(.A1(new_n2557_), .A2(new_n2363_), .Z(new_n2558_));
  XOR2_X1    g02366(.A1(new_n2466_), .A2(\asqrt[51] ), .Z(new_n2559_));
  NOR2_X1    g02367(.A1(\asqrt[44] ), .A2(new_n2559_), .ZN(new_n2560_));
  XOR2_X1    g02368(.A1(new_n2560_), .A2(new_n2365_), .Z(new_n2561_));
  INV_X1     g02369(.I(new_n2561_), .ZN(new_n2562_));
  NOR2_X1    g02370(.A1(new_n2464_), .A2(new_n2415_), .ZN(new_n2563_));
  NOR2_X1    g02371(.A1(\asqrt[44] ), .A2(new_n2563_), .ZN(new_n2564_));
  XOR2_X1    g02372(.A1(new_n2564_), .A2(new_n2369_), .Z(new_n2565_));
  INV_X1     g02373(.I(new_n2565_), .ZN(new_n2566_));
  AOI21_X1   g02374(.A1(new_n2409_), .A2(new_n2414_), .B(\asqrt[44] ), .ZN(new_n2567_));
  XOR2_X1    g02375(.A1(new_n2567_), .A2(new_n2372_), .Z(new_n2568_));
  AOI21_X1   g02376(.A1(new_n2460_), .A2(new_n2408_), .B(\asqrt[44] ), .ZN(new_n2569_));
  XOR2_X1    g02377(.A1(new_n2569_), .A2(new_n2378_), .Z(new_n2570_));
  AOI21_X1   g02378(.A1(new_n2458_), .A2(new_n2405_), .B(\asqrt[44] ), .ZN(new_n2571_));
  XOR2_X1    g02379(.A1(new_n2571_), .A2(new_n2449_), .Z(new_n2572_));
  INV_X1     g02380(.I(new_n2572_), .ZN(new_n2573_));
  NAND2_X1   g02381(.A1(\asqrt[45] ), .A2(new_n2393_), .ZN(new_n2574_));
  NOR2_X1    g02382(.A1(new_n2400_), .A2(\a[90] ), .ZN(new_n2575_));
  AOI22_X1   g02383(.A1(new_n2574_), .A2(new_n2400_), .B1(\asqrt[45] ), .B2(new_n2575_), .ZN(new_n2576_));
  AOI21_X1   g02384(.A1(\asqrt[45] ), .A2(\a[90] ), .B(new_n2398_), .ZN(new_n2577_));
  OAI21_X1   g02385(.A1(new_n2395_), .A2(new_n2577_), .B(new_n2531_), .ZN(new_n2578_));
  XNOR2_X1   g02386(.A1(new_n2578_), .A2(new_n2576_), .ZN(new_n2579_));
  INV_X1     g02387(.I(new_n2579_), .ZN(new_n2580_));
  NAND2_X1   g02388(.A1(new_n2508_), .A2(new_n193_), .ZN(new_n2581_));
  NAND3_X1   g02389(.A1(new_n2514_), .A2(\asqrt[45] ), .A3(new_n2516_), .ZN(new_n2582_));
  NOR3_X1    g02390(.A1(new_n2581_), .A2(new_n2530_), .A3(new_n2582_), .ZN(new_n2583_));
  NOR2_X1    g02391(.A1(new_n2531_), .A2(new_n2391_), .ZN(new_n2584_));
  OAI21_X1   g02392(.A1(new_n2584_), .A2(new_n2583_), .B(new_n2393_), .ZN(new_n2585_));
  NOR3_X1    g02393(.A1(new_n2527_), .A2(\asqrt[63] ), .A3(new_n2530_), .ZN(new_n2586_));
  NAND4_X1   g02394(.A1(new_n2586_), .A2(\asqrt[45] ), .A3(new_n2514_), .A4(new_n2516_), .ZN(new_n2587_));
  NAND2_X1   g02395(.A1(\asqrt[44] ), .A2(new_n2390_), .ZN(new_n2588_));
  NAND3_X1   g02396(.A1(new_n2587_), .A2(new_n2588_), .A3(\a[90] ), .ZN(new_n2589_));
  NAND2_X1   g02397(.A1(new_n2589_), .A2(new_n2585_), .ZN(new_n2590_));
  INV_X1     g02398(.I(new_n2590_), .ZN(new_n2591_));
  INV_X1     g02399(.I(\a[88] ), .ZN(new_n2592_));
  NOR2_X1    g02400(.A1(\a[86] ), .A2(\a[87] ), .ZN(new_n2593_));
  NOR3_X1    g02401(.A1(new_n2531_), .A2(new_n2592_), .A3(new_n2593_), .ZN(new_n2594_));
  INV_X1     g02402(.I(new_n2593_), .ZN(new_n2595_));
  AOI21_X1   g02403(.A1(new_n2531_), .A2(\a[88] ), .B(new_n2595_), .ZN(new_n2596_));
  OAI21_X1   g02404(.A1(new_n2594_), .A2(new_n2596_), .B(\asqrt[45] ), .ZN(new_n2597_));
  NAND2_X1   g02405(.A1(new_n2593_), .A2(new_n2592_), .ZN(new_n2598_));
  NAND3_X1   g02406(.A1(new_n2314_), .A2(new_n2316_), .A3(new_n2598_), .ZN(new_n2599_));
  NAND2_X1   g02407(.A1(new_n2379_), .A2(new_n2599_), .ZN(new_n2600_));
  INV_X1     g02408(.I(new_n2600_), .ZN(new_n2601_));
  NOR3_X1    g02409(.A1(new_n2531_), .A2(new_n2592_), .A3(new_n2601_), .ZN(new_n2602_));
  NOR3_X1    g02410(.A1(new_n2531_), .A2(\a[88] ), .A3(\a[89] ), .ZN(new_n2603_));
  INV_X1     g02411(.I(\a[89] ), .ZN(new_n2604_));
  AOI21_X1   g02412(.A1(\asqrt[44] ), .A2(new_n2592_), .B(new_n2604_), .ZN(new_n2605_));
  NOR3_X1    g02413(.A1(new_n2602_), .A2(new_n2603_), .A3(new_n2605_), .ZN(new_n2606_));
  NAND3_X1   g02414(.A1(new_n2597_), .A2(new_n2606_), .A3(new_n2134_), .ZN(new_n2607_));
  AOI21_X1   g02415(.A1(new_n2597_), .A2(new_n2606_), .B(new_n2134_), .ZN(new_n2608_));
  AOI21_X1   g02416(.A1(new_n2591_), .A2(new_n2607_), .B(new_n2608_), .ZN(new_n2609_));
  AOI21_X1   g02417(.A1(new_n2609_), .A2(new_n1953_), .B(new_n2580_), .ZN(new_n2610_));
  NAND2_X1   g02418(.A1(new_n2591_), .A2(new_n2607_), .ZN(new_n2611_));
  NAND3_X1   g02419(.A1(\asqrt[44] ), .A2(\a[88] ), .A3(new_n2595_), .ZN(new_n2612_));
  OAI21_X1   g02420(.A1(\asqrt[44] ), .A2(new_n2592_), .B(new_n2593_), .ZN(new_n2613_));
  AOI21_X1   g02421(.A1(new_n2613_), .A2(new_n2612_), .B(new_n2332_), .ZN(new_n2614_));
  NAND3_X1   g02422(.A1(\asqrt[44] ), .A2(\a[88] ), .A3(new_n2600_), .ZN(new_n2615_));
  NAND3_X1   g02423(.A1(\asqrt[44] ), .A2(new_n2592_), .A3(new_n2604_), .ZN(new_n2616_));
  OAI21_X1   g02424(.A1(new_n2531_), .A2(\a[88] ), .B(\a[89] ), .ZN(new_n2617_));
  NAND3_X1   g02425(.A1(new_n2617_), .A2(new_n2615_), .A3(new_n2616_), .ZN(new_n2618_));
  OAI21_X1   g02426(.A1(new_n2618_), .A2(new_n2614_), .B(\asqrt[46] ), .ZN(new_n2619_));
  AOI21_X1   g02427(.A1(new_n2611_), .A2(new_n2619_), .B(new_n1953_), .ZN(new_n2620_));
  NOR3_X1    g02428(.A1(new_n2610_), .A2(\asqrt[48] ), .A3(new_n2620_), .ZN(new_n2621_));
  OAI21_X1   g02429(.A1(new_n2610_), .A2(new_n2620_), .B(\asqrt[48] ), .ZN(new_n2622_));
  OAI21_X1   g02430(.A1(new_n2573_), .A2(new_n2621_), .B(new_n2622_), .ZN(new_n2623_));
  OAI21_X1   g02431(.A1(new_n2623_), .A2(\asqrt[49] ), .B(new_n2570_), .ZN(new_n2624_));
  NAND2_X1   g02432(.A1(new_n2623_), .A2(\asqrt[49] ), .ZN(new_n2625_));
  NAND3_X1   g02433(.A1(new_n2624_), .A2(new_n2625_), .A3(new_n1463_), .ZN(new_n2626_));
  AOI21_X1   g02434(.A1(new_n2624_), .A2(new_n2625_), .B(new_n1463_), .ZN(new_n2627_));
  AOI21_X1   g02435(.A1(new_n2568_), .A2(new_n2626_), .B(new_n2627_), .ZN(new_n2628_));
  AOI21_X1   g02436(.A1(new_n2628_), .A2(new_n1305_), .B(new_n2566_), .ZN(new_n2629_));
  NAND2_X1   g02437(.A1(new_n2626_), .A2(new_n2568_), .ZN(new_n2630_));
  INV_X1     g02438(.I(new_n2570_), .ZN(new_n2631_));
  NOR3_X1    g02439(.A1(new_n2618_), .A2(new_n2614_), .A3(\asqrt[46] ), .ZN(new_n2632_));
  OAI21_X1   g02440(.A1(new_n2590_), .A2(new_n2632_), .B(new_n2619_), .ZN(new_n2633_));
  OAI21_X1   g02441(.A1(new_n2633_), .A2(\asqrt[47] ), .B(new_n2579_), .ZN(new_n2634_));
  NAND2_X1   g02442(.A1(new_n2633_), .A2(\asqrt[47] ), .ZN(new_n2635_));
  NAND3_X1   g02443(.A1(new_n2634_), .A2(new_n2635_), .A3(new_n1778_), .ZN(new_n2636_));
  AOI21_X1   g02444(.A1(new_n2634_), .A2(new_n2635_), .B(new_n1778_), .ZN(new_n2637_));
  AOI21_X1   g02445(.A1(new_n2572_), .A2(new_n2636_), .B(new_n2637_), .ZN(new_n2638_));
  AOI21_X1   g02446(.A1(new_n2638_), .A2(new_n1632_), .B(new_n2631_), .ZN(new_n2639_));
  NAND2_X1   g02447(.A1(new_n2636_), .A2(new_n2572_), .ZN(new_n2640_));
  AOI21_X1   g02448(.A1(new_n2640_), .A2(new_n2622_), .B(new_n1632_), .ZN(new_n2641_));
  OAI21_X1   g02449(.A1(new_n2639_), .A2(new_n2641_), .B(\asqrt[50] ), .ZN(new_n2642_));
  AOI21_X1   g02450(.A1(new_n2630_), .A2(new_n2642_), .B(new_n1305_), .ZN(new_n2643_));
  NOR3_X1    g02451(.A1(new_n2629_), .A2(\asqrt[52] ), .A3(new_n2643_), .ZN(new_n2644_));
  OAI21_X1   g02452(.A1(new_n2629_), .A2(new_n2643_), .B(\asqrt[52] ), .ZN(new_n2645_));
  OAI21_X1   g02453(.A1(new_n2562_), .A2(new_n2644_), .B(new_n2645_), .ZN(new_n2646_));
  OAI21_X1   g02454(.A1(new_n2646_), .A2(\asqrt[53] ), .B(new_n2558_), .ZN(new_n2647_));
  NAND2_X1   g02455(.A1(new_n2646_), .A2(\asqrt[53] ), .ZN(new_n2648_));
  NAND3_X1   g02456(.A1(new_n2647_), .A2(new_n2648_), .A3(new_n860_), .ZN(new_n2649_));
  AOI21_X1   g02457(.A1(new_n2647_), .A2(new_n2648_), .B(new_n860_), .ZN(new_n2650_));
  AOI21_X1   g02458(.A1(new_n2556_), .A2(new_n2649_), .B(new_n2650_), .ZN(new_n2651_));
  AOI21_X1   g02459(.A1(new_n2651_), .A2(new_n744_), .B(new_n2554_), .ZN(new_n2652_));
  NAND2_X1   g02460(.A1(new_n2649_), .A2(new_n2556_), .ZN(new_n2653_));
  INV_X1     g02461(.I(new_n2558_), .ZN(new_n2654_));
  INV_X1     g02462(.I(new_n2568_), .ZN(new_n2655_));
  NOR3_X1    g02463(.A1(new_n2639_), .A2(\asqrt[50] ), .A3(new_n2641_), .ZN(new_n2656_));
  OAI21_X1   g02464(.A1(new_n2655_), .A2(new_n2656_), .B(new_n2642_), .ZN(new_n2657_));
  OAI21_X1   g02465(.A1(new_n2657_), .A2(\asqrt[51] ), .B(new_n2565_), .ZN(new_n2658_));
  NAND2_X1   g02466(.A1(new_n2657_), .A2(\asqrt[51] ), .ZN(new_n2659_));
  NAND3_X1   g02467(.A1(new_n2658_), .A2(new_n2659_), .A3(new_n1150_), .ZN(new_n2660_));
  AOI21_X1   g02468(.A1(new_n2658_), .A2(new_n2659_), .B(new_n1150_), .ZN(new_n2661_));
  AOI21_X1   g02469(.A1(new_n2561_), .A2(new_n2660_), .B(new_n2661_), .ZN(new_n2662_));
  AOI21_X1   g02470(.A1(new_n2662_), .A2(new_n1006_), .B(new_n2654_), .ZN(new_n2663_));
  NAND2_X1   g02471(.A1(new_n2660_), .A2(new_n2561_), .ZN(new_n2664_));
  AOI21_X1   g02472(.A1(new_n2664_), .A2(new_n2645_), .B(new_n1006_), .ZN(new_n2665_));
  OAI21_X1   g02473(.A1(new_n2663_), .A2(new_n2665_), .B(\asqrt[54] ), .ZN(new_n2666_));
  AOI21_X1   g02474(.A1(new_n2653_), .A2(new_n2666_), .B(new_n744_), .ZN(new_n2667_));
  NOR3_X1    g02475(.A1(new_n2652_), .A2(\asqrt[56] ), .A3(new_n2667_), .ZN(new_n2668_));
  OAI21_X1   g02476(.A1(new_n2652_), .A2(new_n2667_), .B(\asqrt[56] ), .ZN(new_n2669_));
  OAI21_X1   g02477(.A1(new_n2550_), .A2(new_n2668_), .B(new_n2669_), .ZN(new_n2670_));
  OAI21_X1   g02478(.A1(new_n2670_), .A2(\asqrt[57] ), .B(new_n2545_), .ZN(new_n2671_));
  NOR2_X1    g02479(.A1(new_n2668_), .A2(new_n2550_), .ZN(new_n2672_));
  INV_X1     g02480(.I(new_n2556_), .ZN(new_n2673_));
  NOR3_X1    g02481(.A1(new_n2663_), .A2(\asqrt[54] ), .A3(new_n2665_), .ZN(new_n2674_));
  OAI21_X1   g02482(.A1(new_n2673_), .A2(new_n2674_), .B(new_n2666_), .ZN(new_n2675_));
  OAI21_X1   g02483(.A1(new_n2675_), .A2(\asqrt[55] ), .B(new_n2553_), .ZN(new_n2676_));
  NAND2_X1   g02484(.A1(new_n2675_), .A2(\asqrt[55] ), .ZN(new_n2677_));
  AOI21_X1   g02485(.A1(new_n2676_), .A2(new_n2677_), .B(new_n634_), .ZN(new_n2678_));
  OAI21_X1   g02486(.A1(new_n2672_), .A2(new_n2678_), .B(\asqrt[57] ), .ZN(new_n2679_));
  NAND3_X1   g02487(.A1(new_n2671_), .A2(new_n423_), .A3(new_n2679_), .ZN(new_n2680_));
  NAND2_X1   g02488(.A1(new_n2680_), .A2(new_n2543_), .ZN(new_n2681_));
  INV_X1     g02489(.I(new_n2545_), .ZN(new_n2682_));
  NAND3_X1   g02490(.A1(new_n2676_), .A2(new_n2677_), .A3(new_n634_), .ZN(new_n2683_));
  AOI21_X1   g02491(.A1(new_n2549_), .A2(new_n2683_), .B(new_n2678_), .ZN(new_n2684_));
  AOI21_X1   g02492(.A1(new_n2684_), .A2(new_n531_), .B(new_n2682_), .ZN(new_n2685_));
  NAND2_X1   g02493(.A1(new_n2683_), .A2(new_n2549_), .ZN(new_n2686_));
  AOI21_X1   g02494(.A1(new_n2686_), .A2(new_n2669_), .B(new_n531_), .ZN(new_n2687_));
  OAI21_X1   g02495(.A1(new_n2685_), .A2(new_n2687_), .B(\asqrt[58] ), .ZN(new_n2688_));
  NAND3_X1   g02496(.A1(new_n2681_), .A2(new_n337_), .A3(new_n2688_), .ZN(new_n2689_));
  AOI21_X1   g02497(.A1(new_n2681_), .A2(new_n2688_), .B(new_n337_), .ZN(new_n2690_));
  AOI21_X1   g02498(.A1(new_n2541_), .A2(new_n2689_), .B(new_n2690_), .ZN(new_n2691_));
  AOI21_X1   g02499(.A1(new_n2691_), .A2(new_n266_), .B(new_n2538_), .ZN(new_n2692_));
  INV_X1     g02500(.I(new_n2543_), .ZN(new_n2693_));
  NOR3_X1    g02501(.A1(new_n2685_), .A2(\asqrt[58] ), .A3(new_n2687_), .ZN(new_n2694_));
  OAI21_X1   g02502(.A1(new_n2693_), .A2(new_n2694_), .B(new_n2688_), .ZN(new_n2695_));
  OAI21_X1   g02503(.A1(new_n2695_), .A2(\asqrt[59] ), .B(new_n2541_), .ZN(new_n2696_));
  NAND2_X1   g02504(.A1(new_n2695_), .A2(\asqrt[59] ), .ZN(new_n2697_));
  AOI21_X1   g02505(.A1(new_n2696_), .A2(new_n2697_), .B(new_n266_), .ZN(new_n2698_));
  OAI21_X1   g02506(.A1(new_n2692_), .A2(new_n2698_), .B(\asqrt[61] ), .ZN(new_n2699_));
  AOI21_X1   g02507(.A1(new_n2495_), .A2(new_n2490_), .B(\asqrt[44] ), .ZN(new_n2700_));
  XOR2_X1    g02508(.A1(new_n2700_), .A2(new_n2338_), .Z(new_n2701_));
  INV_X1     g02509(.I(new_n2701_), .ZN(new_n2702_));
  NOR3_X1    g02510(.A1(new_n2692_), .A2(\asqrt[61] ), .A3(new_n2698_), .ZN(new_n2703_));
  OAI21_X1   g02511(.A1(new_n2702_), .A2(new_n2703_), .B(new_n2699_), .ZN(new_n2704_));
  NAND3_X1   g02512(.A1(new_n2696_), .A2(new_n2697_), .A3(new_n266_), .ZN(new_n2705_));
  NAND2_X1   g02513(.A1(new_n2705_), .A2(new_n2537_), .ZN(new_n2706_));
  INV_X1     g02514(.I(new_n2541_), .ZN(new_n2707_));
  AOI21_X1   g02515(.A1(new_n2671_), .A2(new_n2679_), .B(new_n423_), .ZN(new_n2708_));
  AOI21_X1   g02516(.A1(new_n2543_), .A2(new_n2680_), .B(new_n2708_), .ZN(new_n2709_));
  AOI21_X1   g02517(.A1(new_n2709_), .A2(new_n337_), .B(new_n2707_), .ZN(new_n2710_));
  OAI21_X1   g02518(.A1(new_n2710_), .A2(new_n2690_), .B(\asqrt[60] ), .ZN(new_n2711_));
  AOI21_X1   g02519(.A1(new_n2706_), .A2(new_n2711_), .B(new_n239_), .ZN(new_n2712_));
  AOI21_X1   g02520(.A1(new_n2537_), .A2(new_n2705_), .B(new_n2698_), .ZN(new_n2713_));
  AOI21_X1   g02521(.A1(new_n2713_), .A2(new_n239_), .B(new_n2702_), .ZN(new_n2714_));
  OAI21_X1   g02522(.A1(new_n2714_), .A2(new_n2712_), .B(new_n201_), .ZN(new_n2715_));
  NOR3_X1    g02523(.A1(new_n2710_), .A2(\asqrt[60] ), .A3(new_n2690_), .ZN(new_n2716_));
  OAI21_X1   g02524(.A1(new_n2538_), .A2(new_n2716_), .B(new_n2711_), .ZN(new_n2717_));
  OAI21_X1   g02525(.A1(new_n2717_), .A2(\asqrt[61] ), .B(new_n2701_), .ZN(new_n2718_));
  NAND3_X1   g02526(.A1(new_n2718_), .A2(\asqrt[62] ), .A3(new_n2699_), .ZN(new_n2719_));
  AOI21_X1   g02527(.A1(new_n2485_), .A2(new_n2491_), .B(\asqrt[44] ), .ZN(new_n2720_));
  XOR2_X1    g02528(.A1(new_n2720_), .A2(new_n2487_), .Z(new_n2721_));
  INV_X1     g02529(.I(new_n2721_), .ZN(new_n2722_));
  AOI22_X1   g02530(.A1(new_n2719_), .A2(new_n2715_), .B1(new_n2704_), .B2(new_n2722_), .ZN(new_n2723_));
  NOR2_X1    g02531(.A1(new_n2504_), .A2(new_n2335_), .ZN(new_n2724_));
  OAI21_X1   g02532(.A1(\asqrt[44] ), .A2(new_n2724_), .B(new_n2511_), .ZN(new_n2725_));
  INV_X1     g02533(.I(new_n2725_), .ZN(new_n2726_));
  OAI21_X1   g02534(.A1(new_n2723_), .A2(new_n2534_), .B(new_n2726_), .ZN(new_n2727_));
  OAI21_X1   g02535(.A1(new_n2704_), .A2(\asqrt[62] ), .B(new_n2721_), .ZN(new_n2728_));
  NAND2_X1   g02536(.A1(new_n2704_), .A2(\asqrt[62] ), .ZN(new_n2729_));
  NAND3_X1   g02537(.A1(new_n2728_), .A2(new_n2729_), .A3(new_n2534_), .ZN(new_n2730_));
  NAND2_X1   g02538(.A1(new_n2531_), .A2(new_n2334_), .ZN(new_n2731_));
  XOR2_X1    g02539(.A1(new_n2504_), .A2(new_n2335_), .Z(new_n2732_));
  NAND3_X1   g02540(.A1(new_n2731_), .A2(\asqrt[63] ), .A3(new_n2732_), .ZN(new_n2733_));
  INV_X1     g02541(.I(new_n2581_), .ZN(new_n2734_));
  NAND4_X1   g02542(.A1(new_n2734_), .A2(new_n2335_), .A3(new_n2511_), .A4(new_n2518_), .ZN(new_n2735_));
  NAND2_X1   g02543(.A1(new_n2733_), .A2(new_n2735_), .ZN(new_n2736_));
  INV_X1     g02544(.I(new_n2736_), .ZN(new_n2737_));
  NAND4_X1   g02545(.A1(new_n2727_), .A2(new_n193_), .A3(new_n2730_), .A4(new_n2737_), .ZN(\asqrt[43] ));
  NOR2_X1    g02546(.A1(new_n2704_), .A2(\asqrt[62] ), .ZN(new_n2739_));
  NOR2_X1    g02547(.A1(new_n2714_), .A2(new_n2712_), .ZN(new_n2740_));
  NOR2_X1    g02548(.A1(new_n2740_), .A2(new_n201_), .ZN(new_n2741_));
  NOR2_X1    g02549(.A1(new_n2739_), .A2(new_n2741_), .ZN(new_n2742_));
  AOI21_X1   g02550(.A1(new_n2718_), .A2(new_n2699_), .B(\asqrt[62] ), .ZN(new_n2743_));
  NOR3_X1    g02551(.A1(new_n2714_), .A2(new_n201_), .A3(new_n2712_), .ZN(new_n2744_));
  OAI22_X1   g02552(.A1(new_n2743_), .A2(new_n2744_), .B1(new_n2740_), .B2(new_n2721_), .ZN(new_n2745_));
  AOI21_X1   g02553(.A1(new_n2745_), .A2(new_n2533_), .B(new_n2725_), .ZN(new_n2746_));
  AOI21_X1   g02554(.A1(new_n2740_), .A2(new_n201_), .B(new_n2722_), .ZN(new_n2747_));
  NOR3_X1    g02555(.A1(new_n2747_), .A2(new_n2741_), .A3(new_n2533_), .ZN(new_n2748_));
  NOR4_X1    g02556(.A1(new_n2746_), .A2(\asqrt[63] ), .A3(new_n2748_), .A4(new_n2736_), .ZN(new_n2749_));
  XOR2_X1    g02557(.A1(new_n2720_), .A2(new_n2487_), .Z(new_n2750_));
  OAI21_X1   g02558(.A1(\asqrt[43] ), .A2(new_n2742_), .B(new_n2750_), .ZN(new_n2751_));
  INV_X1     g02559(.I(new_n2751_), .ZN(new_n2752_));
  AOI21_X1   g02560(.A1(new_n2689_), .A2(new_n2697_), .B(\asqrt[43] ), .ZN(new_n2753_));
  XOR2_X1    g02561(.A1(new_n2753_), .A2(new_n2541_), .Z(new_n2754_));
  INV_X1     g02562(.I(new_n2754_), .ZN(new_n2755_));
  AOI21_X1   g02563(.A1(new_n2680_), .A2(new_n2688_), .B(\asqrt[43] ), .ZN(new_n2756_));
  XOR2_X1    g02564(.A1(new_n2756_), .A2(new_n2543_), .Z(new_n2757_));
  INV_X1     g02565(.I(new_n2757_), .ZN(new_n2758_));
  NAND2_X1   g02566(.A1(new_n2684_), .A2(new_n531_), .ZN(new_n2759_));
  AOI21_X1   g02567(.A1(new_n2759_), .A2(new_n2679_), .B(\asqrt[43] ), .ZN(new_n2760_));
  XOR2_X1    g02568(.A1(new_n2760_), .A2(new_n2545_), .Z(new_n2761_));
  AOI21_X1   g02569(.A1(new_n2683_), .A2(new_n2669_), .B(\asqrt[43] ), .ZN(new_n2762_));
  XOR2_X1    g02570(.A1(new_n2762_), .A2(new_n2549_), .Z(new_n2763_));
  NAND2_X1   g02571(.A1(new_n2651_), .A2(new_n744_), .ZN(new_n2764_));
  AOI21_X1   g02572(.A1(new_n2764_), .A2(new_n2677_), .B(\asqrt[43] ), .ZN(new_n2765_));
  XOR2_X1    g02573(.A1(new_n2765_), .A2(new_n2553_), .Z(new_n2766_));
  INV_X1     g02574(.I(new_n2766_), .ZN(new_n2767_));
  AOI21_X1   g02575(.A1(new_n2649_), .A2(new_n2666_), .B(\asqrt[43] ), .ZN(new_n2768_));
  XOR2_X1    g02576(.A1(new_n2768_), .A2(new_n2556_), .Z(new_n2769_));
  INV_X1     g02577(.I(new_n2769_), .ZN(new_n2770_));
  NAND2_X1   g02578(.A1(new_n2662_), .A2(new_n1006_), .ZN(new_n2771_));
  AOI21_X1   g02579(.A1(new_n2771_), .A2(new_n2648_), .B(\asqrt[43] ), .ZN(new_n2772_));
  XOR2_X1    g02580(.A1(new_n2772_), .A2(new_n2558_), .Z(new_n2773_));
  AOI21_X1   g02581(.A1(new_n2660_), .A2(new_n2645_), .B(\asqrt[43] ), .ZN(new_n2774_));
  XOR2_X1    g02582(.A1(new_n2774_), .A2(new_n2561_), .Z(new_n2775_));
  NAND2_X1   g02583(.A1(new_n2628_), .A2(new_n1305_), .ZN(new_n2776_));
  AOI21_X1   g02584(.A1(new_n2776_), .A2(new_n2659_), .B(\asqrt[43] ), .ZN(new_n2777_));
  XOR2_X1    g02585(.A1(new_n2777_), .A2(new_n2565_), .Z(new_n2778_));
  INV_X1     g02586(.I(new_n2778_), .ZN(new_n2779_));
  AOI21_X1   g02587(.A1(new_n2626_), .A2(new_n2642_), .B(\asqrt[43] ), .ZN(new_n2780_));
  XOR2_X1    g02588(.A1(new_n2780_), .A2(new_n2568_), .Z(new_n2781_));
  INV_X1     g02589(.I(new_n2781_), .ZN(new_n2782_));
  NAND2_X1   g02590(.A1(new_n2638_), .A2(new_n1632_), .ZN(new_n2783_));
  AOI21_X1   g02591(.A1(new_n2783_), .A2(new_n2625_), .B(\asqrt[43] ), .ZN(new_n2784_));
  XOR2_X1    g02592(.A1(new_n2784_), .A2(new_n2570_), .Z(new_n2785_));
  AOI21_X1   g02593(.A1(new_n2636_), .A2(new_n2622_), .B(\asqrt[43] ), .ZN(new_n2786_));
  XOR2_X1    g02594(.A1(new_n2786_), .A2(new_n2572_), .Z(new_n2787_));
  NAND2_X1   g02595(.A1(new_n2609_), .A2(new_n1953_), .ZN(new_n2788_));
  AOI21_X1   g02596(.A1(new_n2788_), .A2(new_n2635_), .B(\asqrt[43] ), .ZN(new_n2789_));
  XOR2_X1    g02597(.A1(new_n2789_), .A2(new_n2579_), .Z(new_n2790_));
  INV_X1     g02598(.I(new_n2790_), .ZN(new_n2791_));
  AOI21_X1   g02599(.A1(new_n2607_), .A2(new_n2619_), .B(\asqrt[43] ), .ZN(new_n2792_));
  XOR2_X1    g02600(.A1(new_n2792_), .A2(new_n2591_), .Z(new_n2793_));
  INV_X1     g02601(.I(new_n2793_), .ZN(new_n2794_));
  NAND2_X1   g02602(.A1(\asqrt[44] ), .A2(new_n2592_), .ZN(new_n2795_));
  NOR2_X1    g02603(.A1(new_n2604_), .A2(\a[88] ), .ZN(new_n2796_));
  AOI22_X1   g02604(.A1(new_n2795_), .A2(new_n2604_), .B1(\asqrt[44] ), .B2(new_n2796_), .ZN(new_n2797_));
  AOI21_X1   g02605(.A1(\asqrt[44] ), .A2(\a[88] ), .B(new_n2600_), .ZN(new_n2798_));
  OAI21_X1   g02606(.A1(new_n2614_), .A2(new_n2798_), .B(new_n2749_), .ZN(new_n2799_));
  XNOR2_X1   g02607(.A1(new_n2799_), .A2(new_n2797_), .ZN(new_n2800_));
  NAND3_X1   g02608(.A1(new_n2733_), .A2(\asqrt[44] ), .A3(new_n2735_), .ZN(new_n2801_));
  NOR4_X1    g02609(.A1(new_n2746_), .A2(\asqrt[63] ), .A3(new_n2748_), .A4(new_n2801_), .ZN(new_n2802_));
  INV_X1     g02610(.I(new_n2802_), .ZN(new_n2803_));
  NAND2_X1   g02611(.A1(\asqrt[43] ), .A2(new_n2593_), .ZN(new_n2804_));
  AOI21_X1   g02612(.A1(new_n2804_), .A2(new_n2803_), .B(\a[88] ), .ZN(new_n2805_));
  NOR2_X1    g02613(.A1(new_n2749_), .A2(new_n2595_), .ZN(new_n2806_));
  NOR3_X1    g02614(.A1(new_n2806_), .A2(new_n2592_), .A3(new_n2802_), .ZN(new_n2807_));
  NOR2_X1    g02615(.A1(new_n2807_), .A2(new_n2805_), .ZN(new_n2808_));
  INV_X1     g02616(.I(\a[86] ), .ZN(new_n2809_));
  NOR2_X1    g02617(.A1(\a[84] ), .A2(\a[85] ), .ZN(new_n2810_));
  NOR3_X1    g02618(.A1(new_n2749_), .A2(new_n2809_), .A3(new_n2810_), .ZN(new_n2811_));
  INV_X1     g02619(.I(new_n2810_), .ZN(new_n2812_));
  AOI21_X1   g02620(.A1(new_n2749_), .A2(\a[86] ), .B(new_n2812_), .ZN(new_n2813_));
  OAI21_X1   g02621(.A1(new_n2811_), .A2(new_n2813_), .B(\asqrt[44] ), .ZN(new_n2814_));
  NAND2_X1   g02622(.A1(new_n2810_), .A2(new_n2809_), .ZN(new_n2815_));
  NAND3_X1   g02623(.A1(new_n2514_), .A2(new_n2516_), .A3(new_n2815_), .ZN(new_n2816_));
  NAND2_X1   g02624(.A1(new_n2586_), .A2(new_n2816_), .ZN(new_n2817_));
  NAND3_X1   g02625(.A1(\asqrt[43] ), .A2(\a[86] ), .A3(new_n2817_), .ZN(new_n2818_));
  NOR3_X1    g02626(.A1(new_n2749_), .A2(\a[86] ), .A3(\a[87] ), .ZN(new_n2819_));
  INV_X1     g02627(.I(\a[87] ), .ZN(new_n2820_));
  AOI21_X1   g02628(.A1(\asqrt[43] ), .A2(new_n2809_), .B(new_n2820_), .ZN(new_n2821_));
  NOR2_X1    g02629(.A1(new_n2819_), .A2(new_n2821_), .ZN(new_n2822_));
  NAND4_X1   g02630(.A1(new_n2814_), .A2(new_n2822_), .A3(new_n2332_), .A4(new_n2818_), .ZN(new_n2823_));
  NAND2_X1   g02631(.A1(new_n2823_), .A2(new_n2808_), .ZN(new_n2824_));
  NAND3_X1   g02632(.A1(\asqrt[43] ), .A2(\a[86] ), .A3(new_n2812_), .ZN(new_n2825_));
  OAI21_X1   g02633(.A1(\asqrt[43] ), .A2(new_n2809_), .B(new_n2810_), .ZN(new_n2826_));
  AOI21_X1   g02634(.A1(new_n2826_), .A2(new_n2825_), .B(new_n2531_), .ZN(new_n2827_));
  NAND3_X1   g02635(.A1(\asqrt[43] ), .A2(new_n2809_), .A3(new_n2820_), .ZN(new_n2828_));
  OAI21_X1   g02636(.A1(new_n2749_), .A2(\a[86] ), .B(\a[87] ), .ZN(new_n2829_));
  NAND3_X1   g02637(.A1(new_n2818_), .A2(new_n2829_), .A3(new_n2828_), .ZN(new_n2830_));
  OAI21_X1   g02638(.A1(new_n2830_), .A2(new_n2827_), .B(\asqrt[45] ), .ZN(new_n2831_));
  NAND3_X1   g02639(.A1(new_n2824_), .A2(new_n2134_), .A3(new_n2831_), .ZN(new_n2832_));
  AOI21_X1   g02640(.A1(new_n2824_), .A2(new_n2831_), .B(new_n2134_), .ZN(new_n2833_));
  AOI21_X1   g02641(.A1(new_n2800_), .A2(new_n2832_), .B(new_n2833_), .ZN(new_n2834_));
  AOI21_X1   g02642(.A1(new_n2834_), .A2(new_n1953_), .B(new_n2794_), .ZN(new_n2835_));
  OR2_X2     g02643(.A1(new_n2807_), .A2(new_n2805_), .Z(new_n2836_));
  NOR3_X1    g02644(.A1(new_n2830_), .A2(new_n2827_), .A3(\asqrt[45] ), .ZN(new_n2837_));
  OAI21_X1   g02645(.A1(new_n2836_), .A2(new_n2837_), .B(new_n2831_), .ZN(new_n2838_));
  OAI21_X1   g02646(.A1(new_n2838_), .A2(\asqrt[46] ), .B(new_n2800_), .ZN(new_n2839_));
  NAND2_X1   g02647(.A1(new_n2838_), .A2(\asqrt[46] ), .ZN(new_n2840_));
  AOI21_X1   g02648(.A1(new_n2839_), .A2(new_n2840_), .B(new_n1953_), .ZN(new_n2841_));
  NOR3_X1    g02649(.A1(new_n2835_), .A2(\asqrt[48] ), .A3(new_n2841_), .ZN(new_n2842_));
  OAI21_X1   g02650(.A1(new_n2835_), .A2(new_n2841_), .B(\asqrt[48] ), .ZN(new_n2843_));
  OAI21_X1   g02651(.A1(new_n2791_), .A2(new_n2842_), .B(new_n2843_), .ZN(new_n2844_));
  OAI21_X1   g02652(.A1(new_n2844_), .A2(\asqrt[49] ), .B(new_n2787_), .ZN(new_n2845_));
  NAND3_X1   g02653(.A1(new_n2839_), .A2(new_n2840_), .A3(new_n1953_), .ZN(new_n2846_));
  AOI21_X1   g02654(.A1(new_n2793_), .A2(new_n2846_), .B(new_n2841_), .ZN(new_n2847_));
  AOI21_X1   g02655(.A1(new_n2847_), .A2(new_n1778_), .B(new_n2791_), .ZN(new_n2848_));
  NAND2_X1   g02656(.A1(new_n2846_), .A2(new_n2793_), .ZN(new_n2849_));
  INV_X1     g02657(.I(new_n2841_), .ZN(new_n2850_));
  AOI21_X1   g02658(.A1(new_n2849_), .A2(new_n2850_), .B(new_n1778_), .ZN(new_n2851_));
  OAI21_X1   g02659(.A1(new_n2848_), .A2(new_n2851_), .B(\asqrt[49] ), .ZN(new_n2852_));
  NAND3_X1   g02660(.A1(new_n2845_), .A2(new_n1463_), .A3(new_n2852_), .ZN(new_n2853_));
  AOI21_X1   g02661(.A1(new_n2845_), .A2(new_n2852_), .B(new_n1463_), .ZN(new_n2854_));
  AOI21_X1   g02662(.A1(new_n2785_), .A2(new_n2853_), .B(new_n2854_), .ZN(new_n2855_));
  AOI21_X1   g02663(.A1(new_n2855_), .A2(new_n1305_), .B(new_n2782_), .ZN(new_n2856_));
  INV_X1     g02664(.I(new_n2787_), .ZN(new_n2857_));
  NOR3_X1    g02665(.A1(new_n2848_), .A2(\asqrt[49] ), .A3(new_n2851_), .ZN(new_n2858_));
  OAI21_X1   g02666(.A1(new_n2857_), .A2(new_n2858_), .B(new_n2852_), .ZN(new_n2859_));
  OAI21_X1   g02667(.A1(new_n2859_), .A2(\asqrt[50] ), .B(new_n2785_), .ZN(new_n2860_));
  NAND2_X1   g02668(.A1(new_n2859_), .A2(\asqrt[50] ), .ZN(new_n2861_));
  AOI21_X1   g02669(.A1(new_n2860_), .A2(new_n2861_), .B(new_n1305_), .ZN(new_n2862_));
  NOR3_X1    g02670(.A1(new_n2856_), .A2(\asqrt[52] ), .A3(new_n2862_), .ZN(new_n2863_));
  OAI21_X1   g02671(.A1(new_n2856_), .A2(new_n2862_), .B(\asqrt[52] ), .ZN(new_n2864_));
  OAI21_X1   g02672(.A1(new_n2779_), .A2(new_n2863_), .B(new_n2864_), .ZN(new_n2865_));
  OAI21_X1   g02673(.A1(new_n2865_), .A2(\asqrt[53] ), .B(new_n2775_), .ZN(new_n2866_));
  NAND3_X1   g02674(.A1(new_n2860_), .A2(new_n2861_), .A3(new_n1305_), .ZN(new_n2867_));
  AOI21_X1   g02675(.A1(new_n2781_), .A2(new_n2867_), .B(new_n2862_), .ZN(new_n2868_));
  AOI21_X1   g02676(.A1(new_n2868_), .A2(new_n1150_), .B(new_n2779_), .ZN(new_n2869_));
  NAND2_X1   g02677(.A1(new_n2867_), .A2(new_n2781_), .ZN(new_n2870_));
  INV_X1     g02678(.I(new_n2862_), .ZN(new_n2871_));
  AOI21_X1   g02679(.A1(new_n2870_), .A2(new_n2871_), .B(new_n1150_), .ZN(new_n2872_));
  OAI21_X1   g02680(.A1(new_n2869_), .A2(new_n2872_), .B(\asqrt[53] ), .ZN(new_n2873_));
  NAND3_X1   g02681(.A1(new_n2866_), .A2(new_n860_), .A3(new_n2873_), .ZN(new_n2874_));
  AOI21_X1   g02682(.A1(new_n2866_), .A2(new_n2873_), .B(new_n860_), .ZN(new_n2875_));
  AOI21_X1   g02683(.A1(new_n2773_), .A2(new_n2874_), .B(new_n2875_), .ZN(new_n2876_));
  AOI21_X1   g02684(.A1(new_n2876_), .A2(new_n744_), .B(new_n2770_), .ZN(new_n2877_));
  INV_X1     g02685(.I(new_n2775_), .ZN(new_n2878_));
  NOR3_X1    g02686(.A1(new_n2869_), .A2(\asqrt[53] ), .A3(new_n2872_), .ZN(new_n2879_));
  OAI21_X1   g02687(.A1(new_n2878_), .A2(new_n2879_), .B(new_n2873_), .ZN(new_n2880_));
  OAI21_X1   g02688(.A1(new_n2880_), .A2(\asqrt[54] ), .B(new_n2773_), .ZN(new_n2881_));
  NAND2_X1   g02689(.A1(new_n2880_), .A2(\asqrt[54] ), .ZN(new_n2882_));
  AOI21_X1   g02690(.A1(new_n2881_), .A2(new_n2882_), .B(new_n744_), .ZN(new_n2883_));
  NOR3_X1    g02691(.A1(new_n2877_), .A2(\asqrt[56] ), .A3(new_n2883_), .ZN(new_n2884_));
  OAI21_X1   g02692(.A1(new_n2877_), .A2(new_n2883_), .B(\asqrt[56] ), .ZN(new_n2885_));
  OAI21_X1   g02693(.A1(new_n2767_), .A2(new_n2884_), .B(new_n2885_), .ZN(new_n2886_));
  OAI21_X1   g02694(.A1(new_n2886_), .A2(\asqrt[57] ), .B(new_n2763_), .ZN(new_n2887_));
  NAND3_X1   g02695(.A1(new_n2881_), .A2(new_n2882_), .A3(new_n744_), .ZN(new_n2888_));
  AOI21_X1   g02696(.A1(new_n2769_), .A2(new_n2888_), .B(new_n2883_), .ZN(new_n2889_));
  AOI21_X1   g02697(.A1(new_n2889_), .A2(new_n634_), .B(new_n2767_), .ZN(new_n2890_));
  NAND2_X1   g02698(.A1(new_n2888_), .A2(new_n2769_), .ZN(new_n2891_));
  INV_X1     g02699(.I(new_n2883_), .ZN(new_n2892_));
  AOI21_X1   g02700(.A1(new_n2891_), .A2(new_n2892_), .B(new_n634_), .ZN(new_n2893_));
  OAI21_X1   g02701(.A1(new_n2890_), .A2(new_n2893_), .B(\asqrt[57] ), .ZN(new_n2894_));
  NAND3_X1   g02702(.A1(new_n2887_), .A2(new_n423_), .A3(new_n2894_), .ZN(new_n2895_));
  AOI21_X1   g02703(.A1(new_n2887_), .A2(new_n2894_), .B(new_n423_), .ZN(new_n2896_));
  AOI21_X1   g02704(.A1(new_n2761_), .A2(new_n2895_), .B(new_n2896_), .ZN(new_n2897_));
  AOI21_X1   g02705(.A1(new_n2897_), .A2(new_n337_), .B(new_n2758_), .ZN(new_n2898_));
  NOR2_X1    g02706(.A1(new_n2897_), .A2(new_n337_), .ZN(new_n2899_));
  NOR3_X1    g02707(.A1(new_n2898_), .A2(new_n2899_), .A3(\asqrt[60] ), .ZN(new_n2900_));
  OAI21_X1   g02708(.A1(new_n2898_), .A2(new_n2899_), .B(\asqrt[60] ), .ZN(new_n2901_));
  OAI21_X1   g02709(.A1(new_n2755_), .A2(new_n2900_), .B(new_n2901_), .ZN(new_n2902_));
  NAND2_X1   g02710(.A1(new_n2902_), .A2(\asqrt[61] ), .ZN(new_n2903_));
  AOI21_X1   g02711(.A1(new_n2705_), .A2(new_n2711_), .B(\asqrt[43] ), .ZN(new_n2904_));
  XOR2_X1    g02712(.A1(new_n2904_), .A2(new_n2537_), .Z(new_n2905_));
  OAI21_X1   g02713(.A1(new_n2902_), .A2(\asqrt[61] ), .B(new_n2905_), .ZN(new_n2906_));
  NAND2_X1   g02714(.A1(new_n2906_), .A2(new_n2903_), .ZN(new_n2907_));
  INV_X1     g02715(.I(new_n2763_), .ZN(new_n2908_));
  NOR3_X1    g02716(.A1(new_n2890_), .A2(\asqrt[57] ), .A3(new_n2893_), .ZN(new_n2909_));
  OAI21_X1   g02717(.A1(new_n2908_), .A2(new_n2909_), .B(new_n2894_), .ZN(new_n2910_));
  OAI21_X1   g02718(.A1(new_n2910_), .A2(\asqrt[58] ), .B(new_n2761_), .ZN(new_n2911_));
  NOR2_X1    g02719(.A1(new_n2909_), .A2(new_n2908_), .ZN(new_n2912_));
  INV_X1     g02720(.I(new_n2894_), .ZN(new_n2913_));
  OAI21_X1   g02721(.A1(new_n2912_), .A2(new_n2913_), .B(\asqrt[58] ), .ZN(new_n2914_));
  NAND3_X1   g02722(.A1(new_n2911_), .A2(new_n337_), .A3(new_n2914_), .ZN(new_n2915_));
  NAND2_X1   g02723(.A1(new_n2915_), .A2(new_n2757_), .ZN(new_n2916_));
  INV_X1     g02724(.I(new_n2761_), .ZN(new_n2917_));
  NOR2_X1    g02725(.A1(new_n2912_), .A2(new_n2913_), .ZN(new_n2918_));
  AOI21_X1   g02726(.A1(new_n2918_), .A2(new_n423_), .B(new_n2917_), .ZN(new_n2919_));
  OAI21_X1   g02727(.A1(new_n2919_), .A2(new_n2896_), .B(\asqrt[59] ), .ZN(new_n2920_));
  NAND3_X1   g02728(.A1(new_n2916_), .A2(new_n266_), .A3(new_n2920_), .ZN(new_n2921_));
  NAND2_X1   g02729(.A1(new_n2921_), .A2(new_n2754_), .ZN(new_n2922_));
  AOI21_X1   g02730(.A1(new_n2922_), .A2(new_n2901_), .B(new_n239_), .ZN(new_n2923_));
  AOI21_X1   g02731(.A1(new_n2916_), .A2(new_n2920_), .B(new_n266_), .ZN(new_n2924_));
  AOI21_X1   g02732(.A1(new_n2754_), .A2(new_n2921_), .B(new_n2924_), .ZN(new_n2925_));
  INV_X1     g02733(.I(new_n2905_), .ZN(new_n2926_));
  AOI21_X1   g02734(.A1(new_n2925_), .A2(new_n239_), .B(new_n2926_), .ZN(new_n2927_));
  OAI21_X1   g02735(.A1(new_n2927_), .A2(new_n2923_), .B(new_n201_), .ZN(new_n2928_));
  NAND3_X1   g02736(.A1(new_n2906_), .A2(new_n2903_), .A3(\asqrt[62] ), .ZN(new_n2929_));
  NOR2_X1    g02737(.A1(new_n2703_), .A2(new_n2712_), .ZN(new_n2930_));
  NOR2_X1    g02738(.A1(\asqrt[43] ), .A2(new_n2930_), .ZN(new_n2931_));
  XOR2_X1    g02739(.A1(new_n2931_), .A2(new_n2701_), .Z(new_n2932_));
  INV_X1     g02740(.I(new_n2932_), .ZN(new_n2933_));
  AOI22_X1   g02741(.A1(new_n2929_), .A2(new_n2928_), .B1(new_n2907_), .B2(new_n2933_), .ZN(new_n2934_));
  NOR2_X1    g02742(.A1(new_n2723_), .A2(new_n2534_), .ZN(new_n2935_));
  OAI21_X1   g02743(.A1(\asqrt[43] ), .A2(new_n2935_), .B(new_n2730_), .ZN(new_n2936_));
  INV_X1     g02744(.I(new_n2936_), .ZN(new_n2937_));
  OAI21_X1   g02745(.A1(new_n2934_), .A2(new_n2752_), .B(new_n2937_), .ZN(new_n2938_));
  OAI21_X1   g02746(.A1(new_n2907_), .A2(\asqrt[62] ), .B(new_n2932_), .ZN(new_n2939_));
  NAND2_X1   g02747(.A1(new_n2907_), .A2(\asqrt[62] ), .ZN(new_n2940_));
  NAND3_X1   g02748(.A1(new_n2939_), .A2(new_n2940_), .A3(new_n2752_), .ZN(new_n2941_));
  NAND2_X1   g02749(.A1(new_n2749_), .A2(new_n2533_), .ZN(new_n2942_));
  XOR2_X1    g02750(.A1(new_n2745_), .A2(new_n2533_), .Z(new_n2943_));
  NAND3_X1   g02751(.A1(new_n2942_), .A2(\asqrt[63] ), .A3(new_n2943_), .ZN(new_n2944_));
  NOR2_X1    g02752(.A1(new_n2736_), .A2(new_n2533_), .ZN(new_n2945_));
  NAND4_X1   g02753(.A1(new_n2727_), .A2(new_n193_), .A3(new_n2730_), .A4(new_n2945_), .ZN(new_n2946_));
  NAND2_X1   g02754(.A1(new_n2944_), .A2(new_n2946_), .ZN(new_n2947_));
  INV_X1     g02755(.I(new_n2947_), .ZN(new_n2948_));
  NAND4_X1   g02756(.A1(new_n2938_), .A2(new_n193_), .A3(new_n2941_), .A4(new_n2948_), .ZN(\asqrt[42] ));
  NOR2_X1    g02757(.A1(new_n2907_), .A2(\asqrt[62] ), .ZN(new_n2950_));
  NOR2_X1    g02758(.A1(new_n2927_), .A2(new_n2923_), .ZN(new_n2951_));
  NOR2_X1    g02759(.A1(new_n2951_), .A2(new_n201_), .ZN(new_n2952_));
  NOR2_X1    g02760(.A1(new_n2950_), .A2(new_n2952_), .ZN(new_n2953_));
  AOI21_X1   g02761(.A1(new_n2906_), .A2(new_n2903_), .B(\asqrt[62] ), .ZN(new_n2954_));
  NOR3_X1    g02762(.A1(new_n2927_), .A2(new_n201_), .A3(new_n2923_), .ZN(new_n2955_));
  OAI22_X1   g02763(.A1(new_n2954_), .A2(new_n2955_), .B1(new_n2951_), .B2(new_n2932_), .ZN(new_n2956_));
  AOI21_X1   g02764(.A1(new_n2956_), .A2(new_n2751_), .B(new_n2936_), .ZN(new_n2957_));
  AOI21_X1   g02765(.A1(new_n2951_), .A2(new_n201_), .B(new_n2933_), .ZN(new_n2958_));
  NOR3_X1    g02766(.A1(new_n2958_), .A2(new_n2952_), .A3(new_n2751_), .ZN(new_n2959_));
  NOR4_X1    g02767(.A1(new_n2957_), .A2(\asqrt[63] ), .A3(new_n2959_), .A4(new_n2947_), .ZN(new_n2960_));
  XOR2_X1    g02768(.A1(new_n2931_), .A2(new_n2701_), .Z(new_n2961_));
  OAI21_X1   g02769(.A1(\asqrt[42] ), .A2(new_n2953_), .B(new_n2961_), .ZN(new_n2962_));
  INV_X1     g02770(.I(new_n2962_), .ZN(new_n2963_));
  AOI21_X1   g02771(.A1(new_n2915_), .A2(new_n2920_), .B(\asqrt[42] ), .ZN(new_n2964_));
  XOR2_X1    g02772(.A1(new_n2964_), .A2(new_n2757_), .Z(new_n2965_));
  INV_X1     g02773(.I(new_n2965_), .ZN(new_n2966_));
  AOI21_X1   g02774(.A1(new_n2895_), .A2(new_n2914_), .B(\asqrt[42] ), .ZN(new_n2967_));
  XOR2_X1    g02775(.A1(new_n2967_), .A2(new_n2761_), .Z(new_n2968_));
  INV_X1     g02776(.I(new_n2968_), .ZN(new_n2969_));
  NOR2_X1    g02777(.A1(new_n2913_), .A2(new_n2909_), .ZN(new_n2970_));
  NOR2_X1    g02778(.A1(\asqrt[42] ), .A2(new_n2970_), .ZN(new_n2971_));
  XOR2_X1    g02779(.A1(new_n2971_), .A2(new_n2763_), .Z(new_n2972_));
  NOR2_X1    g02780(.A1(new_n2884_), .A2(new_n2893_), .ZN(new_n2973_));
  NOR2_X1    g02781(.A1(\asqrt[42] ), .A2(new_n2973_), .ZN(new_n2974_));
  XOR2_X1    g02782(.A1(new_n2974_), .A2(new_n2766_), .Z(new_n2975_));
  AOI21_X1   g02783(.A1(new_n2888_), .A2(new_n2892_), .B(\asqrt[42] ), .ZN(new_n2976_));
  XOR2_X1    g02784(.A1(new_n2976_), .A2(new_n2769_), .Z(new_n2977_));
  INV_X1     g02785(.I(new_n2977_), .ZN(new_n2978_));
  AOI21_X1   g02786(.A1(new_n2874_), .A2(new_n2882_), .B(\asqrt[42] ), .ZN(new_n2979_));
  XOR2_X1    g02787(.A1(new_n2979_), .A2(new_n2773_), .Z(new_n2980_));
  INV_X1     g02788(.I(new_n2980_), .ZN(new_n2981_));
  XOR2_X1    g02789(.A1(new_n2865_), .A2(\asqrt[53] ), .Z(new_n2982_));
  NOR2_X1    g02790(.A1(\asqrt[42] ), .A2(new_n2982_), .ZN(new_n2983_));
  XOR2_X1    g02791(.A1(new_n2983_), .A2(new_n2775_), .Z(new_n2984_));
  NOR2_X1    g02792(.A1(new_n2863_), .A2(new_n2872_), .ZN(new_n2985_));
  NOR2_X1    g02793(.A1(\asqrt[42] ), .A2(new_n2985_), .ZN(new_n2986_));
  XOR2_X1    g02794(.A1(new_n2986_), .A2(new_n2778_), .Z(new_n2987_));
  AOI21_X1   g02795(.A1(new_n2867_), .A2(new_n2871_), .B(\asqrt[42] ), .ZN(new_n2988_));
  XOR2_X1    g02796(.A1(new_n2988_), .A2(new_n2781_), .Z(new_n2989_));
  INV_X1     g02797(.I(new_n2989_), .ZN(new_n2990_));
  AOI21_X1   g02798(.A1(new_n2853_), .A2(new_n2861_), .B(\asqrt[42] ), .ZN(new_n2991_));
  XOR2_X1    g02799(.A1(new_n2991_), .A2(new_n2785_), .Z(new_n2992_));
  INV_X1     g02800(.I(new_n2992_), .ZN(new_n2993_));
  XOR2_X1    g02801(.A1(new_n2844_), .A2(\asqrt[49] ), .Z(new_n2994_));
  NOR2_X1    g02802(.A1(\asqrt[42] ), .A2(new_n2994_), .ZN(new_n2995_));
  XOR2_X1    g02803(.A1(new_n2995_), .A2(new_n2787_), .Z(new_n2996_));
  NOR2_X1    g02804(.A1(new_n2842_), .A2(new_n2851_), .ZN(new_n2997_));
  NOR2_X1    g02805(.A1(\asqrt[42] ), .A2(new_n2997_), .ZN(new_n2998_));
  XOR2_X1    g02806(.A1(new_n2998_), .A2(new_n2790_), .Z(new_n2999_));
  AOI21_X1   g02807(.A1(new_n2846_), .A2(new_n2850_), .B(\asqrt[42] ), .ZN(new_n3000_));
  XOR2_X1    g02808(.A1(new_n3000_), .A2(new_n2793_), .Z(new_n3001_));
  INV_X1     g02809(.I(new_n3001_), .ZN(new_n3002_));
  AOI21_X1   g02810(.A1(new_n2832_), .A2(new_n2840_), .B(\asqrt[42] ), .ZN(new_n3003_));
  XOR2_X1    g02811(.A1(new_n3003_), .A2(new_n2800_), .Z(new_n3004_));
  INV_X1     g02812(.I(new_n3004_), .ZN(new_n3005_));
  AOI21_X1   g02813(.A1(new_n2823_), .A2(new_n2831_), .B(\asqrt[42] ), .ZN(new_n3006_));
  XOR2_X1    g02814(.A1(new_n3006_), .A2(new_n2808_), .Z(new_n3007_));
  NAND2_X1   g02815(.A1(\asqrt[43] ), .A2(new_n2809_), .ZN(new_n3008_));
  NOR2_X1    g02816(.A1(new_n2820_), .A2(\a[86] ), .ZN(new_n3009_));
  AOI22_X1   g02817(.A1(new_n3008_), .A2(new_n2820_), .B1(\asqrt[43] ), .B2(new_n3009_), .ZN(new_n3010_));
  AOI21_X1   g02818(.A1(\asqrt[43] ), .A2(\a[86] ), .B(new_n2817_), .ZN(new_n3011_));
  OAI21_X1   g02819(.A1(new_n2827_), .A2(new_n3011_), .B(new_n2960_), .ZN(new_n3012_));
  XNOR2_X1   g02820(.A1(new_n3012_), .A2(new_n3010_), .ZN(new_n3013_));
  NOR3_X1    g02821(.A1(new_n2957_), .A2(\asqrt[63] ), .A3(new_n2959_), .ZN(new_n3014_));
  NAND4_X1   g02822(.A1(new_n3014_), .A2(\asqrt[43] ), .A3(new_n2944_), .A4(new_n2946_), .ZN(new_n3015_));
  NAND2_X1   g02823(.A1(\asqrt[42] ), .A2(new_n2810_), .ZN(new_n3016_));
  AOI21_X1   g02824(.A1(new_n3015_), .A2(new_n3016_), .B(\a[86] ), .ZN(new_n3017_));
  NAND2_X1   g02825(.A1(new_n2938_), .A2(new_n193_), .ZN(new_n3018_));
  NAND3_X1   g02826(.A1(new_n2944_), .A2(\asqrt[43] ), .A3(new_n2946_), .ZN(new_n3019_));
  NOR3_X1    g02827(.A1(new_n3018_), .A2(new_n2959_), .A3(new_n3019_), .ZN(new_n3020_));
  NOR2_X1    g02828(.A1(new_n2960_), .A2(new_n2812_), .ZN(new_n3021_));
  NOR3_X1    g02829(.A1(new_n3021_), .A2(new_n3020_), .A3(new_n2809_), .ZN(new_n3022_));
  OR2_X2     g02830(.A1(new_n3017_), .A2(new_n3022_), .Z(new_n3023_));
  NOR2_X1    g02831(.A1(\a[82] ), .A2(\a[83] ), .ZN(new_n3024_));
  INV_X1     g02832(.I(new_n3024_), .ZN(new_n3025_));
  NAND3_X1   g02833(.A1(\asqrt[42] ), .A2(\a[84] ), .A3(new_n3025_), .ZN(new_n3026_));
  INV_X1     g02834(.I(\a[84] ), .ZN(new_n3027_));
  OAI21_X1   g02835(.A1(\asqrt[42] ), .A2(new_n3027_), .B(new_n3024_), .ZN(new_n3028_));
  AOI21_X1   g02836(.A1(new_n3028_), .A2(new_n3026_), .B(new_n2749_), .ZN(new_n3029_));
  NOR3_X1    g02837(.A1(new_n2746_), .A2(\asqrt[63] ), .A3(new_n2748_), .ZN(new_n3030_));
  NAND2_X1   g02838(.A1(new_n3024_), .A2(new_n3027_), .ZN(new_n3031_));
  NAND3_X1   g02839(.A1(new_n2733_), .A2(new_n2735_), .A3(new_n3031_), .ZN(new_n3032_));
  NAND2_X1   g02840(.A1(new_n3030_), .A2(new_n3032_), .ZN(new_n3033_));
  NAND3_X1   g02841(.A1(\asqrt[42] ), .A2(\a[84] ), .A3(new_n3033_), .ZN(new_n3034_));
  INV_X1     g02842(.I(\a[85] ), .ZN(new_n3035_));
  NAND3_X1   g02843(.A1(\asqrt[42] ), .A2(new_n3027_), .A3(new_n3035_), .ZN(new_n3036_));
  OAI21_X1   g02844(.A1(new_n2960_), .A2(\a[84] ), .B(\a[85] ), .ZN(new_n3037_));
  NAND3_X1   g02845(.A1(new_n3034_), .A2(new_n3037_), .A3(new_n3036_), .ZN(new_n3038_));
  NOR3_X1    g02846(.A1(new_n3038_), .A2(new_n3029_), .A3(\asqrt[44] ), .ZN(new_n3039_));
  OAI21_X1   g02847(.A1(new_n3038_), .A2(new_n3029_), .B(\asqrt[44] ), .ZN(new_n3040_));
  OAI21_X1   g02848(.A1(new_n3023_), .A2(new_n3039_), .B(new_n3040_), .ZN(new_n3041_));
  OAI21_X1   g02849(.A1(new_n3041_), .A2(\asqrt[45] ), .B(new_n3013_), .ZN(new_n3042_));
  NAND2_X1   g02850(.A1(new_n3041_), .A2(\asqrt[45] ), .ZN(new_n3043_));
  NAND3_X1   g02851(.A1(new_n3042_), .A2(new_n3043_), .A3(new_n2134_), .ZN(new_n3044_));
  AOI21_X1   g02852(.A1(new_n3042_), .A2(new_n3043_), .B(new_n2134_), .ZN(new_n3045_));
  AOI21_X1   g02853(.A1(new_n3007_), .A2(new_n3044_), .B(new_n3045_), .ZN(new_n3046_));
  AOI21_X1   g02854(.A1(new_n3046_), .A2(new_n1953_), .B(new_n3005_), .ZN(new_n3047_));
  NAND2_X1   g02855(.A1(new_n3044_), .A2(new_n3007_), .ZN(new_n3048_));
  INV_X1     g02856(.I(new_n3013_), .ZN(new_n3049_));
  NOR2_X1    g02857(.A1(new_n3017_), .A2(new_n3022_), .ZN(new_n3050_));
  NOR3_X1    g02858(.A1(new_n2960_), .A2(new_n3027_), .A3(new_n3024_), .ZN(new_n3051_));
  AOI21_X1   g02859(.A1(new_n2960_), .A2(\a[84] ), .B(new_n3025_), .ZN(new_n3052_));
  OAI21_X1   g02860(.A1(new_n3051_), .A2(new_n3052_), .B(\asqrt[43] ), .ZN(new_n3053_));
  INV_X1     g02861(.I(new_n3033_), .ZN(new_n3054_));
  NOR3_X1    g02862(.A1(new_n2960_), .A2(new_n3027_), .A3(new_n3054_), .ZN(new_n3055_));
  NOR3_X1    g02863(.A1(new_n2960_), .A2(\a[84] ), .A3(\a[85] ), .ZN(new_n3056_));
  AOI21_X1   g02864(.A1(\asqrt[42] ), .A2(new_n3027_), .B(new_n3035_), .ZN(new_n3057_));
  NOR3_X1    g02865(.A1(new_n3055_), .A2(new_n3056_), .A3(new_n3057_), .ZN(new_n3058_));
  NAND3_X1   g02866(.A1(new_n3058_), .A2(new_n3053_), .A3(new_n2531_), .ZN(new_n3059_));
  AOI21_X1   g02867(.A1(new_n3058_), .A2(new_n3053_), .B(new_n2531_), .ZN(new_n3060_));
  AOI21_X1   g02868(.A1(new_n3050_), .A2(new_n3059_), .B(new_n3060_), .ZN(new_n3061_));
  AOI21_X1   g02869(.A1(new_n3061_), .A2(new_n2332_), .B(new_n3049_), .ZN(new_n3062_));
  NAND2_X1   g02870(.A1(new_n3059_), .A2(new_n3050_), .ZN(new_n3063_));
  AOI21_X1   g02871(.A1(new_n3063_), .A2(new_n3040_), .B(new_n2332_), .ZN(new_n3064_));
  OAI21_X1   g02872(.A1(new_n3062_), .A2(new_n3064_), .B(\asqrt[46] ), .ZN(new_n3065_));
  AOI21_X1   g02873(.A1(new_n3048_), .A2(new_n3065_), .B(new_n1953_), .ZN(new_n3066_));
  NOR3_X1    g02874(.A1(new_n3047_), .A2(\asqrt[48] ), .A3(new_n3066_), .ZN(new_n3067_));
  OAI21_X1   g02875(.A1(new_n3047_), .A2(new_n3066_), .B(\asqrt[48] ), .ZN(new_n3068_));
  OAI21_X1   g02876(.A1(new_n3002_), .A2(new_n3067_), .B(new_n3068_), .ZN(new_n3069_));
  OAI21_X1   g02877(.A1(new_n3069_), .A2(\asqrt[49] ), .B(new_n2999_), .ZN(new_n3070_));
  NAND2_X1   g02878(.A1(new_n3069_), .A2(\asqrt[49] ), .ZN(new_n3071_));
  NAND3_X1   g02879(.A1(new_n3070_), .A2(new_n3071_), .A3(new_n1463_), .ZN(new_n3072_));
  AOI21_X1   g02880(.A1(new_n3070_), .A2(new_n3071_), .B(new_n1463_), .ZN(new_n3073_));
  AOI21_X1   g02881(.A1(new_n2996_), .A2(new_n3072_), .B(new_n3073_), .ZN(new_n3074_));
  AOI21_X1   g02882(.A1(new_n3074_), .A2(new_n1305_), .B(new_n2993_), .ZN(new_n3075_));
  NAND2_X1   g02883(.A1(new_n3072_), .A2(new_n2996_), .ZN(new_n3076_));
  INV_X1     g02884(.I(new_n2999_), .ZN(new_n3077_));
  INV_X1     g02885(.I(new_n3007_), .ZN(new_n3078_));
  NOR3_X1    g02886(.A1(new_n3062_), .A2(\asqrt[46] ), .A3(new_n3064_), .ZN(new_n3079_));
  OAI21_X1   g02887(.A1(new_n3078_), .A2(new_n3079_), .B(new_n3065_), .ZN(new_n3080_));
  OAI21_X1   g02888(.A1(new_n3080_), .A2(\asqrt[47] ), .B(new_n3004_), .ZN(new_n3081_));
  NAND2_X1   g02889(.A1(new_n3080_), .A2(\asqrt[47] ), .ZN(new_n3082_));
  NAND3_X1   g02890(.A1(new_n3081_), .A2(new_n3082_), .A3(new_n1778_), .ZN(new_n3083_));
  AOI21_X1   g02891(.A1(new_n3081_), .A2(new_n3082_), .B(new_n1778_), .ZN(new_n3084_));
  AOI21_X1   g02892(.A1(new_n3001_), .A2(new_n3083_), .B(new_n3084_), .ZN(new_n3085_));
  AOI21_X1   g02893(.A1(new_n3085_), .A2(new_n1632_), .B(new_n3077_), .ZN(new_n3086_));
  NAND2_X1   g02894(.A1(new_n3083_), .A2(new_n3001_), .ZN(new_n3087_));
  AOI21_X1   g02895(.A1(new_n3087_), .A2(new_n3068_), .B(new_n1632_), .ZN(new_n3088_));
  OAI21_X1   g02896(.A1(new_n3086_), .A2(new_n3088_), .B(\asqrt[50] ), .ZN(new_n3089_));
  AOI21_X1   g02897(.A1(new_n3076_), .A2(new_n3089_), .B(new_n1305_), .ZN(new_n3090_));
  NOR3_X1    g02898(.A1(new_n3075_), .A2(\asqrt[52] ), .A3(new_n3090_), .ZN(new_n3091_));
  OAI21_X1   g02899(.A1(new_n3075_), .A2(new_n3090_), .B(\asqrt[52] ), .ZN(new_n3092_));
  OAI21_X1   g02900(.A1(new_n2990_), .A2(new_n3091_), .B(new_n3092_), .ZN(new_n3093_));
  OAI21_X1   g02901(.A1(new_n3093_), .A2(\asqrt[53] ), .B(new_n2987_), .ZN(new_n3094_));
  NAND2_X1   g02902(.A1(new_n3093_), .A2(\asqrt[53] ), .ZN(new_n3095_));
  NAND3_X1   g02903(.A1(new_n3094_), .A2(new_n3095_), .A3(new_n860_), .ZN(new_n3096_));
  AOI21_X1   g02904(.A1(new_n3094_), .A2(new_n3095_), .B(new_n860_), .ZN(new_n3097_));
  AOI21_X1   g02905(.A1(new_n2984_), .A2(new_n3096_), .B(new_n3097_), .ZN(new_n3098_));
  AOI21_X1   g02906(.A1(new_n3098_), .A2(new_n744_), .B(new_n2981_), .ZN(new_n3099_));
  NAND2_X1   g02907(.A1(new_n3096_), .A2(new_n2984_), .ZN(new_n3100_));
  INV_X1     g02908(.I(new_n2987_), .ZN(new_n3101_));
  INV_X1     g02909(.I(new_n2996_), .ZN(new_n3102_));
  NOR3_X1    g02910(.A1(new_n3086_), .A2(\asqrt[50] ), .A3(new_n3088_), .ZN(new_n3103_));
  OAI21_X1   g02911(.A1(new_n3102_), .A2(new_n3103_), .B(new_n3089_), .ZN(new_n3104_));
  OAI21_X1   g02912(.A1(new_n3104_), .A2(\asqrt[51] ), .B(new_n2992_), .ZN(new_n3105_));
  NAND2_X1   g02913(.A1(new_n3104_), .A2(\asqrt[51] ), .ZN(new_n3106_));
  NAND3_X1   g02914(.A1(new_n3105_), .A2(new_n3106_), .A3(new_n1150_), .ZN(new_n3107_));
  AOI21_X1   g02915(.A1(new_n3105_), .A2(new_n3106_), .B(new_n1150_), .ZN(new_n3108_));
  AOI21_X1   g02916(.A1(new_n2989_), .A2(new_n3107_), .B(new_n3108_), .ZN(new_n3109_));
  AOI21_X1   g02917(.A1(new_n3109_), .A2(new_n1006_), .B(new_n3101_), .ZN(new_n3110_));
  NAND2_X1   g02918(.A1(new_n3107_), .A2(new_n2989_), .ZN(new_n3111_));
  AOI21_X1   g02919(.A1(new_n3111_), .A2(new_n3092_), .B(new_n1006_), .ZN(new_n3112_));
  OAI21_X1   g02920(.A1(new_n3110_), .A2(new_n3112_), .B(\asqrt[54] ), .ZN(new_n3113_));
  AOI21_X1   g02921(.A1(new_n3100_), .A2(new_n3113_), .B(new_n744_), .ZN(new_n3114_));
  NOR3_X1    g02922(.A1(new_n3099_), .A2(\asqrt[56] ), .A3(new_n3114_), .ZN(new_n3115_));
  OAI21_X1   g02923(.A1(new_n3099_), .A2(new_n3114_), .B(\asqrt[56] ), .ZN(new_n3116_));
  OAI21_X1   g02924(.A1(new_n2978_), .A2(new_n3115_), .B(new_n3116_), .ZN(new_n3117_));
  OAI21_X1   g02925(.A1(new_n3117_), .A2(\asqrt[57] ), .B(new_n2975_), .ZN(new_n3118_));
  NAND2_X1   g02926(.A1(new_n3117_), .A2(\asqrt[57] ), .ZN(new_n3119_));
  NAND3_X1   g02927(.A1(new_n3118_), .A2(new_n3119_), .A3(new_n423_), .ZN(new_n3120_));
  AOI21_X1   g02928(.A1(new_n3118_), .A2(new_n3119_), .B(new_n423_), .ZN(new_n3121_));
  AOI21_X1   g02929(.A1(new_n2972_), .A2(new_n3120_), .B(new_n3121_), .ZN(new_n3122_));
  AOI21_X1   g02930(.A1(new_n3122_), .A2(new_n337_), .B(new_n2969_), .ZN(new_n3123_));
  NAND2_X1   g02931(.A1(new_n3120_), .A2(new_n2972_), .ZN(new_n3124_));
  INV_X1     g02932(.I(new_n2975_), .ZN(new_n3125_));
  INV_X1     g02933(.I(new_n2984_), .ZN(new_n3126_));
  NOR3_X1    g02934(.A1(new_n3110_), .A2(\asqrt[54] ), .A3(new_n3112_), .ZN(new_n3127_));
  OAI21_X1   g02935(.A1(new_n3126_), .A2(new_n3127_), .B(new_n3113_), .ZN(new_n3128_));
  OAI21_X1   g02936(.A1(new_n3128_), .A2(\asqrt[55] ), .B(new_n2980_), .ZN(new_n3129_));
  NAND2_X1   g02937(.A1(new_n3128_), .A2(\asqrt[55] ), .ZN(new_n3130_));
  NAND3_X1   g02938(.A1(new_n3129_), .A2(new_n3130_), .A3(new_n634_), .ZN(new_n3131_));
  AOI21_X1   g02939(.A1(new_n3129_), .A2(new_n3130_), .B(new_n634_), .ZN(new_n3132_));
  AOI21_X1   g02940(.A1(new_n2977_), .A2(new_n3131_), .B(new_n3132_), .ZN(new_n3133_));
  AOI21_X1   g02941(.A1(new_n3133_), .A2(new_n531_), .B(new_n3125_), .ZN(new_n3134_));
  NAND2_X1   g02942(.A1(new_n3131_), .A2(new_n2977_), .ZN(new_n3135_));
  AOI21_X1   g02943(.A1(new_n3135_), .A2(new_n3116_), .B(new_n531_), .ZN(new_n3136_));
  OAI21_X1   g02944(.A1(new_n3134_), .A2(new_n3136_), .B(\asqrt[58] ), .ZN(new_n3137_));
  AOI21_X1   g02945(.A1(new_n3124_), .A2(new_n3137_), .B(new_n337_), .ZN(new_n3138_));
  NOR3_X1    g02946(.A1(new_n3123_), .A2(\asqrt[60] ), .A3(new_n3138_), .ZN(new_n3139_));
  NOR2_X1    g02947(.A1(new_n3139_), .A2(new_n2966_), .ZN(new_n3140_));
  INV_X1     g02948(.I(new_n2972_), .ZN(new_n3141_));
  NOR3_X1    g02949(.A1(new_n3134_), .A2(\asqrt[58] ), .A3(new_n3136_), .ZN(new_n3142_));
  OAI21_X1   g02950(.A1(new_n3141_), .A2(new_n3142_), .B(new_n3137_), .ZN(new_n3143_));
  OAI21_X1   g02951(.A1(new_n3143_), .A2(\asqrt[59] ), .B(new_n2968_), .ZN(new_n3144_));
  NOR2_X1    g02952(.A1(new_n3142_), .A2(new_n3141_), .ZN(new_n3145_));
  OAI21_X1   g02953(.A1(new_n3145_), .A2(new_n3121_), .B(\asqrt[59] ), .ZN(new_n3146_));
  AOI21_X1   g02954(.A1(new_n3144_), .A2(new_n3146_), .B(new_n266_), .ZN(new_n3147_));
  OAI21_X1   g02955(.A1(new_n3140_), .A2(new_n3147_), .B(\asqrt[61] ), .ZN(new_n3148_));
  OAI21_X1   g02956(.A1(new_n3123_), .A2(new_n3138_), .B(\asqrt[60] ), .ZN(new_n3149_));
  OAI21_X1   g02957(.A1(new_n2966_), .A2(new_n3139_), .B(new_n3149_), .ZN(new_n3150_));
  AOI21_X1   g02958(.A1(new_n2921_), .A2(new_n2901_), .B(\asqrt[42] ), .ZN(new_n3151_));
  XOR2_X1    g02959(.A1(new_n3151_), .A2(new_n2754_), .Z(new_n3152_));
  OAI21_X1   g02960(.A1(new_n3150_), .A2(\asqrt[61] ), .B(new_n3152_), .ZN(new_n3153_));
  NAND2_X1   g02961(.A1(new_n3153_), .A2(new_n3148_), .ZN(new_n3154_));
  NAND3_X1   g02962(.A1(new_n3144_), .A2(new_n266_), .A3(new_n3146_), .ZN(new_n3155_));
  NAND2_X1   g02963(.A1(new_n3155_), .A2(new_n2965_), .ZN(new_n3156_));
  AOI21_X1   g02964(.A1(new_n3156_), .A2(new_n3149_), .B(new_n239_), .ZN(new_n3157_));
  AOI21_X1   g02965(.A1(new_n2965_), .A2(new_n3155_), .B(new_n3147_), .ZN(new_n3158_));
  INV_X1     g02966(.I(new_n3152_), .ZN(new_n3159_));
  AOI21_X1   g02967(.A1(new_n3158_), .A2(new_n239_), .B(new_n3159_), .ZN(new_n3160_));
  OAI21_X1   g02968(.A1(new_n3160_), .A2(new_n3157_), .B(new_n201_), .ZN(new_n3161_));
  NAND3_X1   g02969(.A1(new_n3153_), .A2(\asqrt[62] ), .A3(new_n3148_), .ZN(new_n3162_));
  NAND2_X1   g02970(.A1(new_n2925_), .A2(new_n239_), .ZN(new_n3163_));
  AOI21_X1   g02971(.A1(new_n2903_), .A2(new_n3163_), .B(\asqrt[42] ), .ZN(new_n3164_));
  XOR2_X1    g02972(.A1(new_n3164_), .A2(new_n2905_), .Z(new_n3165_));
  INV_X1     g02973(.I(new_n3165_), .ZN(new_n3166_));
  AOI22_X1   g02974(.A1(new_n3161_), .A2(new_n3162_), .B1(new_n3154_), .B2(new_n3166_), .ZN(new_n3167_));
  NOR2_X1    g02975(.A1(new_n2934_), .A2(new_n2752_), .ZN(new_n3168_));
  OAI21_X1   g02976(.A1(\asqrt[42] ), .A2(new_n3168_), .B(new_n2941_), .ZN(new_n3169_));
  INV_X1     g02977(.I(new_n3169_), .ZN(new_n3170_));
  OAI21_X1   g02978(.A1(new_n3167_), .A2(new_n2963_), .B(new_n3170_), .ZN(new_n3171_));
  OAI21_X1   g02979(.A1(new_n3154_), .A2(\asqrt[62] ), .B(new_n3165_), .ZN(new_n3172_));
  NAND2_X1   g02980(.A1(new_n3154_), .A2(\asqrt[62] ), .ZN(new_n3173_));
  NAND3_X1   g02981(.A1(new_n3172_), .A2(new_n3173_), .A3(new_n2963_), .ZN(new_n3174_));
  NAND2_X1   g02982(.A1(new_n2960_), .A2(new_n2751_), .ZN(new_n3175_));
  XOR2_X1    g02983(.A1(new_n2956_), .A2(new_n2751_), .Z(new_n3176_));
  NAND3_X1   g02984(.A1(new_n3175_), .A2(\asqrt[63] ), .A3(new_n3176_), .ZN(new_n3177_));
  INV_X1     g02985(.I(new_n3018_), .ZN(new_n3178_));
  NAND4_X1   g02986(.A1(new_n3178_), .A2(new_n2752_), .A3(new_n2941_), .A4(new_n2948_), .ZN(new_n3179_));
  NAND2_X1   g02987(.A1(new_n3177_), .A2(new_n3179_), .ZN(new_n3180_));
  INV_X1     g02988(.I(new_n3180_), .ZN(new_n3181_));
  NAND4_X1   g02989(.A1(new_n3171_), .A2(new_n193_), .A3(new_n3174_), .A4(new_n3181_), .ZN(\asqrt[41] ));
  NOR2_X1    g02990(.A1(new_n3154_), .A2(\asqrt[62] ), .ZN(new_n3183_));
  INV_X1     g02991(.I(new_n3173_), .ZN(new_n3184_));
  NOR2_X1    g02992(.A1(new_n3184_), .A2(new_n3183_), .ZN(new_n3185_));
  NAND3_X1   g02993(.A1(new_n3156_), .A2(new_n239_), .A3(new_n3149_), .ZN(new_n3186_));
  AOI21_X1   g02994(.A1(new_n3152_), .A2(new_n3186_), .B(new_n3157_), .ZN(new_n3187_));
  AOI21_X1   g02995(.A1(new_n3153_), .A2(new_n3148_), .B(\asqrt[62] ), .ZN(new_n3188_));
  NOR3_X1    g02996(.A1(new_n3160_), .A2(new_n201_), .A3(new_n3157_), .ZN(new_n3189_));
  OAI22_X1   g02997(.A1(new_n3189_), .A2(new_n3188_), .B1(new_n3187_), .B2(new_n3165_), .ZN(new_n3190_));
  AOI21_X1   g02998(.A1(new_n3190_), .A2(new_n2962_), .B(new_n3169_), .ZN(new_n3191_));
  AOI21_X1   g02999(.A1(new_n3187_), .A2(new_n201_), .B(new_n3166_), .ZN(new_n3192_));
  OAI21_X1   g03000(.A1(new_n3187_), .A2(new_n201_), .B(new_n2963_), .ZN(new_n3193_));
  NOR2_X1    g03001(.A1(new_n3192_), .A2(new_n3193_), .ZN(new_n3194_));
  NOR4_X1    g03002(.A1(new_n3191_), .A2(\asqrt[63] ), .A3(new_n3194_), .A4(new_n3180_), .ZN(new_n3195_));
  XOR2_X1    g03003(.A1(new_n3164_), .A2(new_n2905_), .Z(new_n3196_));
  OAI21_X1   g03004(.A1(\asqrt[41] ), .A2(new_n3185_), .B(new_n3196_), .ZN(new_n3197_));
  INV_X1     g03005(.I(new_n3197_), .ZN(new_n3198_));
  NAND2_X1   g03006(.A1(new_n3122_), .A2(new_n337_), .ZN(new_n3199_));
  AOI21_X1   g03007(.A1(new_n3199_), .A2(new_n3146_), .B(\asqrt[41] ), .ZN(new_n3200_));
  XOR2_X1    g03008(.A1(new_n3200_), .A2(new_n2968_), .Z(new_n3201_));
  INV_X1     g03009(.I(new_n3201_), .ZN(new_n3202_));
  AOI21_X1   g03010(.A1(new_n3120_), .A2(new_n3137_), .B(\asqrt[41] ), .ZN(new_n3203_));
  XOR2_X1    g03011(.A1(new_n3203_), .A2(new_n2972_), .Z(new_n3204_));
  INV_X1     g03012(.I(new_n3204_), .ZN(new_n3205_));
  NAND2_X1   g03013(.A1(new_n3133_), .A2(new_n531_), .ZN(new_n3206_));
  AOI21_X1   g03014(.A1(new_n3206_), .A2(new_n3119_), .B(\asqrt[41] ), .ZN(new_n3207_));
  XOR2_X1    g03015(.A1(new_n3207_), .A2(new_n2975_), .Z(new_n3208_));
  INV_X1     g03016(.I(new_n3208_), .ZN(new_n3209_));
  AOI21_X1   g03017(.A1(new_n3131_), .A2(new_n3116_), .B(\asqrt[41] ), .ZN(new_n3210_));
  XOR2_X1    g03018(.A1(new_n3210_), .A2(new_n2977_), .Z(new_n3211_));
  NAND2_X1   g03019(.A1(new_n3098_), .A2(new_n744_), .ZN(new_n3212_));
  AOI21_X1   g03020(.A1(new_n3212_), .A2(new_n3130_), .B(\asqrt[41] ), .ZN(new_n3213_));
  XOR2_X1    g03021(.A1(new_n3213_), .A2(new_n2980_), .Z(new_n3214_));
  AOI21_X1   g03022(.A1(new_n3096_), .A2(new_n3113_), .B(\asqrt[41] ), .ZN(new_n3215_));
  XOR2_X1    g03023(.A1(new_n3215_), .A2(new_n2984_), .Z(new_n3216_));
  INV_X1     g03024(.I(new_n3216_), .ZN(new_n3217_));
  NAND2_X1   g03025(.A1(new_n3109_), .A2(new_n1006_), .ZN(new_n3218_));
  AOI21_X1   g03026(.A1(new_n3218_), .A2(new_n3095_), .B(\asqrt[41] ), .ZN(new_n3219_));
  XOR2_X1    g03027(.A1(new_n3219_), .A2(new_n2987_), .Z(new_n3220_));
  INV_X1     g03028(.I(new_n3220_), .ZN(new_n3221_));
  AOI21_X1   g03029(.A1(new_n3107_), .A2(new_n3092_), .B(\asqrt[41] ), .ZN(new_n3222_));
  XOR2_X1    g03030(.A1(new_n3222_), .A2(new_n2989_), .Z(new_n3223_));
  NAND2_X1   g03031(.A1(new_n3074_), .A2(new_n1305_), .ZN(new_n3224_));
  AOI21_X1   g03032(.A1(new_n3224_), .A2(new_n3106_), .B(\asqrt[41] ), .ZN(new_n3225_));
  XOR2_X1    g03033(.A1(new_n3225_), .A2(new_n2992_), .Z(new_n3226_));
  AOI21_X1   g03034(.A1(new_n3072_), .A2(new_n3089_), .B(\asqrt[41] ), .ZN(new_n3227_));
  XOR2_X1    g03035(.A1(new_n3227_), .A2(new_n2996_), .Z(new_n3228_));
  INV_X1     g03036(.I(new_n3228_), .ZN(new_n3229_));
  NAND2_X1   g03037(.A1(new_n3085_), .A2(new_n1632_), .ZN(new_n3230_));
  AOI21_X1   g03038(.A1(new_n3230_), .A2(new_n3071_), .B(\asqrt[41] ), .ZN(new_n3231_));
  XOR2_X1    g03039(.A1(new_n3231_), .A2(new_n2999_), .Z(new_n3232_));
  INV_X1     g03040(.I(new_n3232_), .ZN(new_n3233_));
  AOI21_X1   g03041(.A1(new_n3083_), .A2(new_n3068_), .B(\asqrt[41] ), .ZN(new_n3234_));
  XOR2_X1    g03042(.A1(new_n3234_), .A2(new_n3001_), .Z(new_n3235_));
  NAND2_X1   g03043(.A1(new_n3046_), .A2(new_n1953_), .ZN(new_n3236_));
  AOI21_X1   g03044(.A1(new_n3236_), .A2(new_n3082_), .B(\asqrt[41] ), .ZN(new_n3237_));
  XOR2_X1    g03045(.A1(new_n3237_), .A2(new_n3004_), .Z(new_n3238_));
  AOI21_X1   g03046(.A1(new_n3044_), .A2(new_n3065_), .B(\asqrt[41] ), .ZN(new_n3239_));
  XOR2_X1    g03047(.A1(new_n3239_), .A2(new_n3007_), .Z(new_n3240_));
  INV_X1     g03048(.I(new_n3240_), .ZN(new_n3241_));
  NAND2_X1   g03049(.A1(new_n3061_), .A2(new_n2332_), .ZN(new_n3242_));
  AOI21_X1   g03050(.A1(new_n3242_), .A2(new_n3043_), .B(\asqrt[41] ), .ZN(new_n3243_));
  XOR2_X1    g03051(.A1(new_n3243_), .A2(new_n3013_), .Z(new_n3244_));
  INV_X1     g03052(.I(new_n3244_), .ZN(new_n3245_));
  AOI21_X1   g03053(.A1(new_n3059_), .A2(new_n3040_), .B(\asqrt[41] ), .ZN(new_n3246_));
  XOR2_X1    g03054(.A1(new_n3246_), .A2(new_n3050_), .Z(new_n3247_));
  NAND2_X1   g03055(.A1(\asqrt[42] ), .A2(new_n3027_), .ZN(new_n3248_));
  NOR2_X1    g03056(.A1(new_n3035_), .A2(\a[84] ), .ZN(new_n3249_));
  AOI22_X1   g03057(.A1(new_n3248_), .A2(new_n3035_), .B1(\asqrt[42] ), .B2(new_n3249_), .ZN(new_n3250_));
  AOI21_X1   g03058(.A1(\asqrt[42] ), .A2(\a[84] ), .B(new_n3033_), .ZN(new_n3251_));
  OAI21_X1   g03059(.A1(new_n3029_), .A2(new_n3251_), .B(new_n3195_), .ZN(new_n3252_));
  XNOR2_X1   g03060(.A1(new_n3252_), .A2(new_n3250_), .ZN(new_n3253_));
  NOR3_X1    g03061(.A1(new_n3191_), .A2(\asqrt[63] ), .A3(new_n3194_), .ZN(new_n3254_));
  NAND3_X1   g03062(.A1(new_n3177_), .A2(\asqrt[42] ), .A3(new_n3179_), .ZN(new_n3255_));
  INV_X1     g03063(.I(new_n3255_), .ZN(new_n3256_));
  NAND2_X1   g03064(.A1(new_n3254_), .A2(new_n3256_), .ZN(new_n3257_));
  NAND2_X1   g03065(.A1(\asqrt[41] ), .A2(new_n3024_), .ZN(new_n3258_));
  AOI21_X1   g03066(.A1(new_n3258_), .A2(new_n3257_), .B(\a[84] ), .ZN(new_n3259_));
  NAND2_X1   g03067(.A1(new_n3171_), .A2(new_n193_), .ZN(new_n3260_));
  NOR3_X1    g03068(.A1(new_n3260_), .A2(new_n3194_), .A3(new_n3255_), .ZN(new_n3261_));
  NOR2_X1    g03069(.A1(new_n3195_), .A2(new_n3025_), .ZN(new_n3262_));
  NOR3_X1    g03070(.A1(new_n3262_), .A2(new_n3261_), .A3(new_n3027_), .ZN(new_n3263_));
  OR2_X2     g03071(.A1(new_n3263_), .A2(new_n3259_), .Z(new_n3264_));
  NOR2_X1    g03072(.A1(\a[80] ), .A2(\a[81] ), .ZN(new_n3265_));
  INV_X1     g03073(.I(new_n3265_), .ZN(new_n3266_));
  NAND3_X1   g03074(.A1(\asqrt[41] ), .A2(\a[82] ), .A3(new_n3266_), .ZN(new_n3267_));
  INV_X1     g03075(.I(\a[82] ), .ZN(new_n3268_));
  OAI21_X1   g03076(.A1(\asqrt[41] ), .A2(new_n3268_), .B(new_n3265_), .ZN(new_n3269_));
  AOI21_X1   g03077(.A1(new_n3269_), .A2(new_n3267_), .B(new_n2960_), .ZN(new_n3270_));
  NAND2_X1   g03078(.A1(new_n3265_), .A2(new_n3268_), .ZN(new_n3271_));
  NAND3_X1   g03079(.A1(new_n2944_), .A2(new_n2946_), .A3(new_n3271_), .ZN(new_n3272_));
  NAND2_X1   g03080(.A1(new_n3014_), .A2(new_n3272_), .ZN(new_n3273_));
  NAND3_X1   g03081(.A1(\asqrt[41] ), .A2(\a[82] ), .A3(new_n3273_), .ZN(new_n3274_));
  INV_X1     g03082(.I(\a[83] ), .ZN(new_n3275_));
  NAND3_X1   g03083(.A1(\asqrt[41] ), .A2(new_n3268_), .A3(new_n3275_), .ZN(new_n3276_));
  OAI21_X1   g03084(.A1(new_n3195_), .A2(\a[82] ), .B(\a[83] ), .ZN(new_n3277_));
  NAND3_X1   g03085(.A1(new_n3274_), .A2(new_n3277_), .A3(new_n3276_), .ZN(new_n3278_));
  NOR3_X1    g03086(.A1(new_n3278_), .A2(new_n3270_), .A3(\asqrt[43] ), .ZN(new_n3279_));
  OAI21_X1   g03087(.A1(new_n3278_), .A2(new_n3270_), .B(\asqrt[43] ), .ZN(new_n3280_));
  OAI21_X1   g03088(.A1(new_n3264_), .A2(new_n3279_), .B(new_n3280_), .ZN(new_n3281_));
  OAI21_X1   g03089(.A1(new_n3281_), .A2(\asqrt[44] ), .B(new_n3253_), .ZN(new_n3282_));
  NAND2_X1   g03090(.A1(new_n3281_), .A2(\asqrt[44] ), .ZN(new_n3283_));
  NAND3_X1   g03091(.A1(new_n3282_), .A2(new_n3283_), .A3(new_n2332_), .ZN(new_n3284_));
  AOI21_X1   g03092(.A1(new_n3282_), .A2(new_n3283_), .B(new_n2332_), .ZN(new_n3285_));
  AOI21_X1   g03093(.A1(new_n3247_), .A2(new_n3284_), .B(new_n3285_), .ZN(new_n3286_));
  AOI21_X1   g03094(.A1(new_n3286_), .A2(new_n2134_), .B(new_n3245_), .ZN(new_n3287_));
  NAND2_X1   g03095(.A1(new_n3284_), .A2(new_n3247_), .ZN(new_n3288_));
  INV_X1     g03096(.I(new_n3285_), .ZN(new_n3289_));
  AOI21_X1   g03097(.A1(new_n3288_), .A2(new_n3289_), .B(new_n2134_), .ZN(new_n3290_));
  NOR3_X1    g03098(.A1(new_n3287_), .A2(\asqrt[47] ), .A3(new_n3290_), .ZN(new_n3291_));
  OAI21_X1   g03099(.A1(new_n3287_), .A2(new_n3290_), .B(\asqrt[47] ), .ZN(new_n3292_));
  OAI21_X1   g03100(.A1(new_n3241_), .A2(new_n3291_), .B(new_n3292_), .ZN(new_n3293_));
  OAI21_X1   g03101(.A1(new_n3293_), .A2(\asqrt[48] ), .B(new_n3238_), .ZN(new_n3294_));
  NAND2_X1   g03102(.A1(new_n3293_), .A2(\asqrt[48] ), .ZN(new_n3295_));
  NAND3_X1   g03103(.A1(new_n3294_), .A2(new_n3295_), .A3(new_n1632_), .ZN(new_n3296_));
  AOI21_X1   g03104(.A1(new_n3294_), .A2(new_n3295_), .B(new_n1632_), .ZN(new_n3297_));
  AOI21_X1   g03105(.A1(new_n3235_), .A2(new_n3296_), .B(new_n3297_), .ZN(new_n3298_));
  AOI21_X1   g03106(.A1(new_n3298_), .A2(new_n1463_), .B(new_n3233_), .ZN(new_n3299_));
  NAND2_X1   g03107(.A1(new_n3296_), .A2(new_n3235_), .ZN(new_n3300_));
  INV_X1     g03108(.I(new_n3297_), .ZN(new_n3301_));
  AOI21_X1   g03109(.A1(new_n3300_), .A2(new_n3301_), .B(new_n1463_), .ZN(new_n3302_));
  NOR3_X1    g03110(.A1(new_n3299_), .A2(\asqrt[51] ), .A3(new_n3302_), .ZN(new_n3303_));
  OAI21_X1   g03111(.A1(new_n3299_), .A2(new_n3302_), .B(\asqrt[51] ), .ZN(new_n3304_));
  OAI21_X1   g03112(.A1(new_n3229_), .A2(new_n3303_), .B(new_n3304_), .ZN(new_n3305_));
  OAI21_X1   g03113(.A1(new_n3305_), .A2(\asqrt[52] ), .B(new_n3226_), .ZN(new_n3306_));
  NAND2_X1   g03114(.A1(new_n3305_), .A2(\asqrt[52] ), .ZN(new_n3307_));
  NAND3_X1   g03115(.A1(new_n3306_), .A2(new_n3307_), .A3(new_n1006_), .ZN(new_n3308_));
  AOI21_X1   g03116(.A1(new_n3306_), .A2(new_n3307_), .B(new_n1006_), .ZN(new_n3309_));
  AOI21_X1   g03117(.A1(new_n3223_), .A2(new_n3308_), .B(new_n3309_), .ZN(new_n3310_));
  AOI21_X1   g03118(.A1(new_n3310_), .A2(new_n860_), .B(new_n3221_), .ZN(new_n3311_));
  NAND2_X1   g03119(.A1(new_n3308_), .A2(new_n3223_), .ZN(new_n3312_));
  INV_X1     g03120(.I(new_n3309_), .ZN(new_n3313_));
  AOI21_X1   g03121(.A1(new_n3312_), .A2(new_n3313_), .B(new_n860_), .ZN(new_n3314_));
  NOR3_X1    g03122(.A1(new_n3311_), .A2(\asqrt[55] ), .A3(new_n3314_), .ZN(new_n3315_));
  OAI21_X1   g03123(.A1(new_n3311_), .A2(new_n3314_), .B(\asqrt[55] ), .ZN(new_n3316_));
  OAI21_X1   g03124(.A1(new_n3217_), .A2(new_n3315_), .B(new_n3316_), .ZN(new_n3317_));
  OAI21_X1   g03125(.A1(new_n3317_), .A2(\asqrt[56] ), .B(new_n3214_), .ZN(new_n3318_));
  NAND2_X1   g03126(.A1(new_n3317_), .A2(\asqrt[56] ), .ZN(new_n3319_));
  NAND3_X1   g03127(.A1(new_n3318_), .A2(new_n3319_), .A3(new_n531_), .ZN(new_n3320_));
  AOI21_X1   g03128(.A1(new_n3318_), .A2(new_n3319_), .B(new_n531_), .ZN(new_n3321_));
  AOI21_X1   g03129(.A1(new_n3211_), .A2(new_n3320_), .B(new_n3321_), .ZN(new_n3322_));
  AOI21_X1   g03130(.A1(new_n3322_), .A2(new_n423_), .B(new_n3209_), .ZN(new_n3323_));
  NAND2_X1   g03131(.A1(new_n3320_), .A2(new_n3211_), .ZN(new_n3324_));
  INV_X1     g03132(.I(new_n3321_), .ZN(new_n3325_));
  AOI21_X1   g03133(.A1(new_n3324_), .A2(new_n3325_), .B(new_n423_), .ZN(new_n3326_));
  NOR3_X1    g03134(.A1(new_n3323_), .A2(\asqrt[59] ), .A3(new_n3326_), .ZN(new_n3327_));
  NOR2_X1    g03135(.A1(new_n3327_), .A2(new_n3205_), .ZN(new_n3328_));
  OAI21_X1   g03136(.A1(new_n3323_), .A2(new_n3326_), .B(\asqrt[59] ), .ZN(new_n3329_));
  INV_X1     g03137(.I(new_n3329_), .ZN(new_n3330_));
  NOR2_X1    g03138(.A1(new_n3328_), .A2(new_n3330_), .ZN(new_n3331_));
  AOI21_X1   g03139(.A1(new_n3331_), .A2(new_n266_), .B(new_n3202_), .ZN(new_n3332_));
  INV_X1     g03140(.I(new_n3211_), .ZN(new_n3333_));
  INV_X1     g03141(.I(new_n3223_), .ZN(new_n3334_));
  INV_X1     g03142(.I(new_n3235_), .ZN(new_n3335_));
  INV_X1     g03143(.I(new_n3247_), .ZN(new_n3336_));
  NOR2_X1    g03144(.A1(new_n3263_), .A2(new_n3259_), .ZN(new_n3337_));
  NOR3_X1    g03145(.A1(new_n3195_), .A2(new_n3268_), .A3(new_n3265_), .ZN(new_n3338_));
  AOI21_X1   g03146(.A1(new_n3195_), .A2(\a[82] ), .B(new_n3266_), .ZN(new_n3339_));
  OAI21_X1   g03147(.A1(new_n3338_), .A2(new_n3339_), .B(\asqrt[42] ), .ZN(new_n3340_));
  INV_X1     g03148(.I(new_n3273_), .ZN(new_n3341_));
  NOR3_X1    g03149(.A1(new_n3195_), .A2(new_n3268_), .A3(new_n3341_), .ZN(new_n3342_));
  NOR3_X1    g03150(.A1(new_n3195_), .A2(\a[82] ), .A3(\a[83] ), .ZN(new_n3343_));
  AOI21_X1   g03151(.A1(\asqrt[41] ), .A2(new_n3268_), .B(new_n3275_), .ZN(new_n3344_));
  NOR3_X1    g03152(.A1(new_n3342_), .A2(new_n3343_), .A3(new_n3344_), .ZN(new_n3345_));
  NAND3_X1   g03153(.A1(new_n3345_), .A2(new_n3340_), .A3(new_n2749_), .ZN(new_n3346_));
  NAND2_X1   g03154(.A1(new_n3346_), .A2(new_n3337_), .ZN(new_n3347_));
  NAND3_X1   g03155(.A1(new_n3347_), .A2(new_n2531_), .A3(new_n3280_), .ZN(new_n3348_));
  AOI21_X1   g03156(.A1(new_n3347_), .A2(new_n3280_), .B(new_n2531_), .ZN(new_n3349_));
  AOI21_X1   g03157(.A1(new_n3253_), .A2(new_n3348_), .B(new_n3349_), .ZN(new_n3350_));
  AOI21_X1   g03158(.A1(new_n3350_), .A2(new_n2332_), .B(new_n3336_), .ZN(new_n3351_));
  NOR3_X1    g03159(.A1(new_n3351_), .A2(\asqrt[46] ), .A3(new_n3285_), .ZN(new_n3352_));
  OAI21_X1   g03160(.A1(new_n3351_), .A2(new_n3285_), .B(\asqrt[46] ), .ZN(new_n3353_));
  OAI21_X1   g03161(.A1(new_n3245_), .A2(new_n3352_), .B(new_n3353_), .ZN(new_n3354_));
  OAI21_X1   g03162(.A1(new_n3354_), .A2(\asqrt[47] ), .B(new_n3240_), .ZN(new_n3355_));
  NAND3_X1   g03163(.A1(new_n3355_), .A2(new_n1778_), .A3(new_n3292_), .ZN(new_n3356_));
  AOI21_X1   g03164(.A1(new_n3355_), .A2(new_n3292_), .B(new_n1778_), .ZN(new_n3357_));
  AOI21_X1   g03165(.A1(new_n3238_), .A2(new_n3356_), .B(new_n3357_), .ZN(new_n3358_));
  AOI21_X1   g03166(.A1(new_n3358_), .A2(new_n1632_), .B(new_n3335_), .ZN(new_n3359_));
  NOR3_X1    g03167(.A1(new_n3359_), .A2(\asqrt[50] ), .A3(new_n3297_), .ZN(new_n3360_));
  OAI21_X1   g03168(.A1(new_n3359_), .A2(new_n3297_), .B(\asqrt[50] ), .ZN(new_n3361_));
  OAI21_X1   g03169(.A1(new_n3233_), .A2(new_n3360_), .B(new_n3361_), .ZN(new_n3362_));
  OAI21_X1   g03170(.A1(new_n3362_), .A2(\asqrt[51] ), .B(new_n3228_), .ZN(new_n3363_));
  NAND3_X1   g03171(.A1(new_n3363_), .A2(new_n1150_), .A3(new_n3304_), .ZN(new_n3364_));
  AOI21_X1   g03172(.A1(new_n3363_), .A2(new_n3304_), .B(new_n1150_), .ZN(new_n3365_));
  AOI21_X1   g03173(.A1(new_n3226_), .A2(new_n3364_), .B(new_n3365_), .ZN(new_n3366_));
  AOI21_X1   g03174(.A1(new_n3366_), .A2(new_n1006_), .B(new_n3334_), .ZN(new_n3367_));
  NOR3_X1    g03175(.A1(new_n3367_), .A2(\asqrt[54] ), .A3(new_n3309_), .ZN(new_n3368_));
  OAI21_X1   g03176(.A1(new_n3367_), .A2(new_n3309_), .B(\asqrt[54] ), .ZN(new_n3369_));
  OAI21_X1   g03177(.A1(new_n3221_), .A2(new_n3368_), .B(new_n3369_), .ZN(new_n3370_));
  OAI21_X1   g03178(.A1(new_n3370_), .A2(\asqrt[55] ), .B(new_n3216_), .ZN(new_n3371_));
  NAND3_X1   g03179(.A1(new_n3371_), .A2(new_n634_), .A3(new_n3316_), .ZN(new_n3372_));
  AOI21_X1   g03180(.A1(new_n3371_), .A2(new_n3316_), .B(new_n634_), .ZN(new_n3373_));
  AOI21_X1   g03181(.A1(new_n3214_), .A2(new_n3372_), .B(new_n3373_), .ZN(new_n3374_));
  AOI21_X1   g03182(.A1(new_n3374_), .A2(new_n531_), .B(new_n3333_), .ZN(new_n3375_));
  NOR3_X1    g03183(.A1(new_n3375_), .A2(\asqrt[58] ), .A3(new_n3321_), .ZN(new_n3376_));
  OAI21_X1   g03184(.A1(new_n3375_), .A2(new_n3321_), .B(\asqrt[58] ), .ZN(new_n3377_));
  OAI21_X1   g03185(.A1(new_n3209_), .A2(new_n3376_), .B(new_n3377_), .ZN(new_n3378_));
  OAI21_X1   g03186(.A1(new_n3378_), .A2(\asqrt[59] ), .B(new_n3204_), .ZN(new_n3379_));
  AOI21_X1   g03187(.A1(new_n3379_), .A2(new_n3329_), .B(new_n266_), .ZN(new_n3380_));
  OAI21_X1   g03188(.A1(new_n3332_), .A2(new_n3380_), .B(\asqrt[61] ), .ZN(new_n3381_));
  AOI21_X1   g03189(.A1(new_n3155_), .A2(new_n3149_), .B(\asqrt[41] ), .ZN(new_n3382_));
  XOR2_X1    g03190(.A1(new_n3382_), .A2(new_n2965_), .Z(new_n3383_));
  OAI21_X1   g03191(.A1(new_n3205_), .A2(new_n3327_), .B(new_n3329_), .ZN(new_n3384_));
  OAI21_X1   g03192(.A1(new_n3384_), .A2(\asqrt[60] ), .B(new_n3201_), .ZN(new_n3385_));
  OAI21_X1   g03193(.A1(new_n3328_), .A2(new_n3330_), .B(\asqrt[60] ), .ZN(new_n3386_));
  NAND3_X1   g03194(.A1(new_n3385_), .A2(new_n239_), .A3(new_n3386_), .ZN(new_n3387_));
  NAND2_X1   g03195(.A1(new_n3387_), .A2(new_n3383_), .ZN(new_n3388_));
  NAND2_X1   g03196(.A1(new_n3388_), .A2(new_n3381_), .ZN(new_n3389_));
  AOI21_X1   g03197(.A1(new_n3385_), .A2(new_n3386_), .B(new_n239_), .ZN(new_n3390_));
  NAND3_X1   g03198(.A1(new_n3379_), .A2(new_n266_), .A3(new_n3329_), .ZN(new_n3391_));
  AOI21_X1   g03199(.A1(new_n3201_), .A2(new_n3391_), .B(new_n3380_), .ZN(new_n3392_));
  INV_X1     g03200(.I(new_n3383_), .ZN(new_n3393_));
  AOI21_X1   g03201(.A1(new_n3392_), .A2(new_n239_), .B(new_n3393_), .ZN(new_n3394_));
  OAI21_X1   g03202(.A1(new_n3394_), .A2(new_n3390_), .B(new_n201_), .ZN(new_n3395_));
  NAND3_X1   g03203(.A1(new_n3388_), .A2(\asqrt[62] ), .A3(new_n3381_), .ZN(new_n3396_));
  AOI21_X1   g03204(.A1(new_n3148_), .A2(new_n3186_), .B(\asqrt[41] ), .ZN(new_n3397_));
  XOR2_X1    g03205(.A1(new_n3397_), .A2(new_n3152_), .Z(new_n3398_));
  INV_X1     g03206(.I(new_n3398_), .ZN(new_n3399_));
  AOI22_X1   g03207(.A1(new_n3395_), .A2(new_n3396_), .B1(new_n3389_), .B2(new_n3399_), .ZN(new_n3400_));
  NOR2_X1    g03208(.A1(new_n3167_), .A2(new_n2963_), .ZN(new_n3401_));
  OAI21_X1   g03209(.A1(\asqrt[41] ), .A2(new_n3401_), .B(new_n3174_), .ZN(new_n3402_));
  INV_X1     g03210(.I(new_n3402_), .ZN(new_n3403_));
  OAI21_X1   g03211(.A1(new_n3400_), .A2(new_n3198_), .B(new_n3403_), .ZN(new_n3404_));
  OAI21_X1   g03212(.A1(new_n3389_), .A2(\asqrt[62] ), .B(new_n3398_), .ZN(new_n3405_));
  NAND2_X1   g03213(.A1(new_n3389_), .A2(\asqrt[62] ), .ZN(new_n3406_));
  NAND3_X1   g03214(.A1(new_n3405_), .A2(new_n3406_), .A3(new_n3198_), .ZN(new_n3407_));
  NAND2_X1   g03215(.A1(new_n3195_), .A2(new_n2962_), .ZN(new_n3408_));
  XOR2_X1    g03216(.A1(new_n3167_), .A2(new_n2963_), .Z(new_n3409_));
  NAND3_X1   g03217(.A1(new_n3408_), .A2(\asqrt[63] ), .A3(new_n3409_), .ZN(new_n3410_));
  INV_X1     g03218(.I(new_n3260_), .ZN(new_n3411_));
  NAND4_X1   g03219(.A1(new_n3411_), .A2(new_n2963_), .A3(new_n3174_), .A4(new_n3181_), .ZN(new_n3412_));
  NAND2_X1   g03220(.A1(new_n3410_), .A2(new_n3412_), .ZN(new_n3413_));
  INV_X1     g03221(.I(new_n3413_), .ZN(new_n3414_));
  NAND4_X1   g03222(.A1(new_n3404_), .A2(new_n193_), .A3(new_n3407_), .A4(new_n3414_), .ZN(\asqrt[40] ));
  NOR2_X1    g03223(.A1(new_n3389_), .A2(\asqrt[62] ), .ZN(new_n3416_));
  INV_X1     g03224(.I(new_n3406_), .ZN(new_n3417_));
  NOR2_X1    g03225(.A1(new_n3417_), .A2(new_n3416_), .ZN(new_n3418_));
  NOR2_X1    g03226(.A1(new_n3394_), .A2(new_n3390_), .ZN(new_n3419_));
  AOI21_X1   g03227(.A1(new_n3388_), .A2(new_n3381_), .B(\asqrt[62] ), .ZN(new_n3420_));
  NOR3_X1    g03228(.A1(new_n3394_), .A2(new_n201_), .A3(new_n3390_), .ZN(new_n3421_));
  OAI22_X1   g03229(.A1(new_n3421_), .A2(new_n3420_), .B1(new_n3419_), .B2(new_n3398_), .ZN(new_n3422_));
  AOI21_X1   g03230(.A1(new_n3422_), .A2(new_n3197_), .B(new_n3402_), .ZN(new_n3423_));
  AOI21_X1   g03231(.A1(new_n3419_), .A2(new_n201_), .B(new_n3399_), .ZN(new_n3424_));
  OAI21_X1   g03232(.A1(new_n3419_), .A2(new_n201_), .B(new_n3198_), .ZN(new_n3425_));
  NOR2_X1    g03233(.A1(new_n3424_), .A2(new_n3425_), .ZN(new_n3426_));
  NOR4_X1    g03234(.A1(new_n3423_), .A2(\asqrt[63] ), .A3(new_n3426_), .A4(new_n3413_), .ZN(new_n3427_));
  XOR2_X1    g03235(.A1(new_n3397_), .A2(new_n3152_), .Z(new_n3428_));
  OAI21_X1   g03236(.A1(\asqrt[40] ), .A2(new_n3418_), .B(new_n3428_), .ZN(new_n3429_));
  INV_X1     g03237(.I(new_n3429_), .ZN(new_n3430_));
  NOR2_X1    g03238(.A1(new_n3330_), .A2(new_n3327_), .ZN(new_n3431_));
  NOR2_X1    g03239(.A1(\asqrt[40] ), .A2(new_n3431_), .ZN(new_n3432_));
  XOR2_X1    g03240(.A1(new_n3432_), .A2(new_n3204_), .Z(new_n3433_));
  INV_X1     g03241(.I(new_n3433_), .ZN(new_n3434_));
  NOR2_X1    g03242(.A1(new_n3376_), .A2(new_n3326_), .ZN(new_n3435_));
  NOR2_X1    g03243(.A1(\asqrt[40] ), .A2(new_n3435_), .ZN(new_n3436_));
  XOR2_X1    g03244(.A1(new_n3436_), .A2(new_n3208_), .Z(new_n3437_));
  AOI21_X1   g03245(.A1(new_n3320_), .A2(new_n3325_), .B(\asqrt[40] ), .ZN(new_n3438_));
  XOR2_X1    g03246(.A1(new_n3438_), .A2(new_n3211_), .Z(new_n3439_));
  AOI21_X1   g03247(.A1(new_n3372_), .A2(new_n3319_), .B(\asqrt[40] ), .ZN(new_n3440_));
  XOR2_X1    g03248(.A1(new_n3440_), .A2(new_n3214_), .Z(new_n3441_));
  INV_X1     g03249(.I(new_n3316_), .ZN(new_n3442_));
  NOR2_X1    g03250(.A1(new_n3442_), .A2(new_n3315_), .ZN(new_n3443_));
  NOR2_X1    g03251(.A1(\asqrt[40] ), .A2(new_n3443_), .ZN(new_n3444_));
  XOR2_X1    g03252(.A1(new_n3444_), .A2(new_n3216_), .Z(new_n3445_));
  INV_X1     g03253(.I(new_n3445_), .ZN(new_n3446_));
  NOR2_X1    g03254(.A1(new_n3368_), .A2(new_n3314_), .ZN(new_n3447_));
  NOR2_X1    g03255(.A1(\asqrt[40] ), .A2(new_n3447_), .ZN(new_n3448_));
  XOR2_X1    g03256(.A1(new_n3448_), .A2(new_n3220_), .Z(new_n3449_));
  INV_X1     g03257(.I(new_n3449_), .ZN(new_n3450_));
  AOI21_X1   g03258(.A1(new_n3308_), .A2(new_n3313_), .B(\asqrt[40] ), .ZN(new_n3451_));
  XOR2_X1    g03259(.A1(new_n3451_), .A2(new_n3223_), .Z(new_n3452_));
  AOI21_X1   g03260(.A1(new_n3364_), .A2(new_n3307_), .B(\asqrt[40] ), .ZN(new_n3453_));
  XOR2_X1    g03261(.A1(new_n3453_), .A2(new_n3226_), .Z(new_n3454_));
  XOR2_X1    g03262(.A1(new_n3362_), .A2(\asqrt[51] ), .Z(new_n3455_));
  NOR2_X1    g03263(.A1(\asqrt[40] ), .A2(new_n3455_), .ZN(new_n3456_));
  XOR2_X1    g03264(.A1(new_n3456_), .A2(new_n3228_), .Z(new_n3457_));
  INV_X1     g03265(.I(new_n3457_), .ZN(new_n3458_));
  NOR2_X1    g03266(.A1(new_n3360_), .A2(new_n3302_), .ZN(new_n3459_));
  NOR2_X1    g03267(.A1(\asqrt[40] ), .A2(new_n3459_), .ZN(new_n3460_));
  XOR2_X1    g03268(.A1(new_n3460_), .A2(new_n3232_), .Z(new_n3461_));
  INV_X1     g03269(.I(new_n3461_), .ZN(new_n3462_));
  AOI21_X1   g03270(.A1(new_n3296_), .A2(new_n3301_), .B(\asqrt[40] ), .ZN(new_n3463_));
  XOR2_X1    g03271(.A1(new_n3463_), .A2(new_n3235_), .Z(new_n3464_));
  AOI21_X1   g03272(.A1(new_n3356_), .A2(new_n3295_), .B(\asqrt[40] ), .ZN(new_n3465_));
  XOR2_X1    g03273(.A1(new_n3465_), .A2(new_n3238_), .Z(new_n3466_));
  XOR2_X1    g03274(.A1(new_n3354_), .A2(\asqrt[47] ), .Z(new_n3467_));
  NOR2_X1    g03275(.A1(\asqrt[40] ), .A2(new_n3467_), .ZN(new_n3468_));
  XOR2_X1    g03276(.A1(new_n3468_), .A2(new_n3240_), .Z(new_n3469_));
  INV_X1     g03277(.I(new_n3469_), .ZN(new_n3470_));
  NOR2_X1    g03278(.A1(new_n3352_), .A2(new_n3290_), .ZN(new_n3471_));
  NOR2_X1    g03279(.A1(\asqrt[40] ), .A2(new_n3471_), .ZN(new_n3472_));
  XOR2_X1    g03280(.A1(new_n3472_), .A2(new_n3244_), .Z(new_n3473_));
  INV_X1     g03281(.I(new_n3473_), .ZN(new_n3474_));
  AOI21_X1   g03282(.A1(new_n3284_), .A2(new_n3289_), .B(\asqrt[40] ), .ZN(new_n3475_));
  XOR2_X1    g03283(.A1(new_n3475_), .A2(new_n3247_), .Z(new_n3476_));
  AOI21_X1   g03284(.A1(new_n3348_), .A2(new_n3283_), .B(\asqrt[40] ), .ZN(new_n3477_));
  XOR2_X1    g03285(.A1(new_n3477_), .A2(new_n3253_), .Z(new_n3478_));
  AOI21_X1   g03286(.A1(new_n3346_), .A2(new_n3280_), .B(\asqrt[40] ), .ZN(new_n3479_));
  XOR2_X1    g03287(.A1(new_n3479_), .A2(new_n3337_), .Z(new_n3480_));
  INV_X1     g03288(.I(new_n3480_), .ZN(new_n3481_));
  NAND2_X1   g03289(.A1(\asqrt[41] ), .A2(new_n3268_), .ZN(new_n3482_));
  NOR2_X1    g03290(.A1(new_n3275_), .A2(\a[82] ), .ZN(new_n3483_));
  AOI22_X1   g03291(.A1(new_n3482_), .A2(new_n3275_), .B1(\asqrt[41] ), .B2(new_n3483_), .ZN(new_n3484_));
  AOI21_X1   g03292(.A1(\asqrt[41] ), .A2(\a[82] ), .B(new_n3273_), .ZN(new_n3485_));
  OAI21_X1   g03293(.A1(new_n3270_), .A2(new_n3485_), .B(new_n3427_), .ZN(new_n3486_));
  XNOR2_X1   g03294(.A1(new_n3486_), .A2(new_n3484_), .ZN(new_n3487_));
  INV_X1     g03295(.I(new_n3487_), .ZN(new_n3488_));
  NAND2_X1   g03296(.A1(new_n3404_), .A2(new_n193_), .ZN(new_n3489_));
  NAND3_X1   g03297(.A1(new_n3410_), .A2(\asqrt[41] ), .A3(new_n3412_), .ZN(new_n3490_));
  NOR3_X1    g03298(.A1(new_n3489_), .A2(new_n3426_), .A3(new_n3490_), .ZN(new_n3491_));
  NOR2_X1    g03299(.A1(new_n3427_), .A2(new_n3266_), .ZN(new_n3492_));
  OAI21_X1   g03300(.A1(new_n3492_), .A2(new_n3491_), .B(new_n3268_), .ZN(new_n3493_));
  NOR3_X1    g03301(.A1(new_n3423_), .A2(\asqrt[63] ), .A3(new_n3426_), .ZN(new_n3494_));
  NAND4_X1   g03302(.A1(new_n3494_), .A2(\asqrt[41] ), .A3(new_n3410_), .A4(new_n3412_), .ZN(new_n3495_));
  NAND2_X1   g03303(.A1(\asqrt[40] ), .A2(new_n3265_), .ZN(new_n3496_));
  NAND3_X1   g03304(.A1(new_n3495_), .A2(new_n3496_), .A3(\a[82] ), .ZN(new_n3497_));
  NAND2_X1   g03305(.A1(new_n3497_), .A2(new_n3493_), .ZN(new_n3498_));
  INV_X1     g03306(.I(new_n3498_), .ZN(new_n3499_));
  INV_X1     g03307(.I(\a[80] ), .ZN(new_n3500_));
  NOR2_X1    g03308(.A1(\a[78] ), .A2(\a[79] ), .ZN(new_n3501_));
  NOR3_X1    g03309(.A1(new_n3427_), .A2(new_n3500_), .A3(new_n3501_), .ZN(new_n3502_));
  INV_X1     g03310(.I(new_n3501_), .ZN(new_n3503_));
  AOI21_X1   g03311(.A1(new_n3427_), .A2(\a[80] ), .B(new_n3503_), .ZN(new_n3504_));
  OAI21_X1   g03312(.A1(new_n3502_), .A2(new_n3504_), .B(\asqrt[41] ), .ZN(new_n3505_));
  NAND2_X1   g03313(.A1(new_n3501_), .A2(new_n3500_), .ZN(new_n3506_));
  NAND3_X1   g03314(.A1(new_n3177_), .A2(new_n3179_), .A3(new_n3506_), .ZN(new_n3507_));
  NAND2_X1   g03315(.A1(new_n3254_), .A2(new_n3507_), .ZN(new_n3508_));
  INV_X1     g03316(.I(new_n3508_), .ZN(new_n3509_));
  NOR3_X1    g03317(.A1(new_n3427_), .A2(new_n3500_), .A3(new_n3509_), .ZN(new_n3510_));
  NOR3_X1    g03318(.A1(new_n3427_), .A2(\a[80] ), .A3(\a[81] ), .ZN(new_n3511_));
  INV_X1     g03319(.I(\a[81] ), .ZN(new_n3512_));
  AOI21_X1   g03320(.A1(\asqrt[40] ), .A2(new_n3500_), .B(new_n3512_), .ZN(new_n3513_));
  NOR3_X1    g03321(.A1(new_n3510_), .A2(new_n3511_), .A3(new_n3513_), .ZN(new_n3514_));
  NAND3_X1   g03322(.A1(new_n3505_), .A2(new_n3514_), .A3(new_n2960_), .ZN(new_n3515_));
  AOI21_X1   g03323(.A1(new_n3505_), .A2(new_n3514_), .B(new_n2960_), .ZN(new_n3516_));
  AOI21_X1   g03324(.A1(new_n3499_), .A2(new_n3515_), .B(new_n3516_), .ZN(new_n3517_));
  AOI21_X1   g03325(.A1(new_n3517_), .A2(new_n2749_), .B(new_n3488_), .ZN(new_n3518_));
  NAND2_X1   g03326(.A1(new_n3499_), .A2(new_n3515_), .ZN(new_n3519_));
  NAND3_X1   g03327(.A1(\asqrt[40] ), .A2(\a[80] ), .A3(new_n3503_), .ZN(new_n3520_));
  OAI21_X1   g03328(.A1(\asqrt[40] ), .A2(new_n3500_), .B(new_n3501_), .ZN(new_n3521_));
  AOI21_X1   g03329(.A1(new_n3521_), .A2(new_n3520_), .B(new_n3195_), .ZN(new_n3522_));
  NAND3_X1   g03330(.A1(\asqrt[40] ), .A2(\a[80] ), .A3(new_n3508_), .ZN(new_n3523_));
  NAND3_X1   g03331(.A1(\asqrt[40] ), .A2(new_n3500_), .A3(new_n3512_), .ZN(new_n3524_));
  OAI21_X1   g03332(.A1(new_n3427_), .A2(\a[80] ), .B(\a[81] ), .ZN(new_n3525_));
  NAND3_X1   g03333(.A1(new_n3525_), .A2(new_n3523_), .A3(new_n3524_), .ZN(new_n3526_));
  OAI21_X1   g03334(.A1(new_n3526_), .A2(new_n3522_), .B(\asqrt[42] ), .ZN(new_n3527_));
  AOI21_X1   g03335(.A1(new_n3519_), .A2(new_n3527_), .B(new_n2749_), .ZN(new_n3528_));
  NOR3_X1    g03336(.A1(new_n3518_), .A2(\asqrt[44] ), .A3(new_n3528_), .ZN(new_n3529_));
  OAI21_X1   g03337(.A1(new_n3518_), .A2(new_n3528_), .B(\asqrt[44] ), .ZN(new_n3530_));
  OAI21_X1   g03338(.A1(new_n3481_), .A2(new_n3529_), .B(new_n3530_), .ZN(new_n3531_));
  OAI21_X1   g03339(.A1(new_n3531_), .A2(\asqrt[45] ), .B(new_n3478_), .ZN(new_n3532_));
  NAND2_X1   g03340(.A1(new_n3531_), .A2(\asqrt[45] ), .ZN(new_n3533_));
  NAND3_X1   g03341(.A1(new_n3532_), .A2(new_n3533_), .A3(new_n2134_), .ZN(new_n3534_));
  AOI21_X1   g03342(.A1(new_n3532_), .A2(new_n3533_), .B(new_n2134_), .ZN(new_n3535_));
  AOI21_X1   g03343(.A1(new_n3476_), .A2(new_n3534_), .B(new_n3535_), .ZN(new_n3536_));
  AOI21_X1   g03344(.A1(new_n3536_), .A2(new_n1953_), .B(new_n3474_), .ZN(new_n3537_));
  NAND2_X1   g03345(.A1(new_n3534_), .A2(new_n3476_), .ZN(new_n3538_));
  INV_X1     g03346(.I(new_n3478_), .ZN(new_n3539_));
  NOR3_X1    g03347(.A1(new_n3526_), .A2(new_n3522_), .A3(\asqrt[42] ), .ZN(new_n3540_));
  OAI21_X1   g03348(.A1(new_n3498_), .A2(new_n3540_), .B(new_n3527_), .ZN(new_n3541_));
  OAI21_X1   g03349(.A1(new_n3541_), .A2(\asqrt[43] ), .B(new_n3487_), .ZN(new_n3542_));
  NAND2_X1   g03350(.A1(new_n3541_), .A2(\asqrt[43] ), .ZN(new_n3543_));
  NAND3_X1   g03351(.A1(new_n3542_), .A2(new_n3543_), .A3(new_n2531_), .ZN(new_n3544_));
  AOI21_X1   g03352(.A1(new_n3542_), .A2(new_n3543_), .B(new_n2531_), .ZN(new_n3545_));
  AOI21_X1   g03353(.A1(new_n3480_), .A2(new_n3544_), .B(new_n3545_), .ZN(new_n3546_));
  AOI21_X1   g03354(.A1(new_n3546_), .A2(new_n2332_), .B(new_n3539_), .ZN(new_n3547_));
  NAND2_X1   g03355(.A1(new_n3544_), .A2(new_n3480_), .ZN(new_n3548_));
  AOI21_X1   g03356(.A1(new_n3548_), .A2(new_n3530_), .B(new_n2332_), .ZN(new_n3549_));
  OAI21_X1   g03357(.A1(new_n3547_), .A2(new_n3549_), .B(\asqrt[46] ), .ZN(new_n3550_));
  AOI21_X1   g03358(.A1(new_n3538_), .A2(new_n3550_), .B(new_n1953_), .ZN(new_n3551_));
  NOR3_X1    g03359(.A1(new_n3537_), .A2(\asqrt[48] ), .A3(new_n3551_), .ZN(new_n3552_));
  OAI21_X1   g03360(.A1(new_n3537_), .A2(new_n3551_), .B(\asqrt[48] ), .ZN(new_n3553_));
  OAI21_X1   g03361(.A1(new_n3470_), .A2(new_n3552_), .B(new_n3553_), .ZN(new_n3554_));
  OAI21_X1   g03362(.A1(new_n3554_), .A2(\asqrt[49] ), .B(new_n3466_), .ZN(new_n3555_));
  NAND2_X1   g03363(.A1(new_n3554_), .A2(\asqrt[49] ), .ZN(new_n3556_));
  NAND3_X1   g03364(.A1(new_n3555_), .A2(new_n3556_), .A3(new_n1463_), .ZN(new_n3557_));
  AOI21_X1   g03365(.A1(new_n3555_), .A2(new_n3556_), .B(new_n1463_), .ZN(new_n3558_));
  AOI21_X1   g03366(.A1(new_n3464_), .A2(new_n3557_), .B(new_n3558_), .ZN(new_n3559_));
  AOI21_X1   g03367(.A1(new_n3559_), .A2(new_n1305_), .B(new_n3462_), .ZN(new_n3560_));
  NAND2_X1   g03368(.A1(new_n3557_), .A2(new_n3464_), .ZN(new_n3561_));
  INV_X1     g03369(.I(new_n3466_), .ZN(new_n3562_));
  INV_X1     g03370(.I(new_n3476_), .ZN(new_n3563_));
  NOR3_X1    g03371(.A1(new_n3547_), .A2(\asqrt[46] ), .A3(new_n3549_), .ZN(new_n3564_));
  OAI21_X1   g03372(.A1(new_n3563_), .A2(new_n3564_), .B(new_n3550_), .ZN(new_n3565_));
  OAI21_X1   g03373(.A1(new_n3565_), .A2(\asqrt[47] ), .B(new_n3473_), .ZN(new_n3566_));
  NAND2_X1   g03374(.A1(new_n3565_), .A2(\asqrt[47] ), .ZN(new_n3567_));
  NAND3_X1   g03375(.A1(new_n3566_), .A2(new_n3567_), .A3(new_n1778_), .ZN(new_n3568_));
  AOI21_X1   g03376(.A1(new_n3566_), .A2(new_n3567_), .B(new_n1778_), .ZN(new_n3569_));
  AOI21_X1   g03377(.A1(new_n3469_), .A2(new_n3568_), .B(new_n3569_), .ZN(new_n3570_));
  AOI21_X1   g03378(.A1(new_n3570_), .A2(new_n1632_), .B(new_n3562_), .ZN(new_n3571_));
  NAND2_X1   g03379(.A1(new_n3568_), .A2(new_n3469_), .ZN(new_n3572_));
  AOI21_X1   g03380(.A1(new_n3572_), .A2(new_n3553_), .B(new_n1632_), .ZN(new_n3573_));
  OAI21_X1   g03381(.A1(new_n3571_), .A2(new_n3573_), .B(\asqrt[50] ), .ZN(new_n3574_));
  AOI21_X1   g03382(.A1(new_n3561_), .A2(new_n3574_), .B(new_n1305_), .ZN(new_n3575_));
  NOR3_X1    g03383(.A1(new_n3560_), .A2(\asqrt[52] ), .A3(new_n3575_), .ZN(new_n3576_));
  OAI21_X1   g03384(.A1(new_n3560_), .A2(new_n3575_), .B(\asqrt[52] ), .ZN(new_n3577_));
  OAI21_X1   g03385(.A1(new_n3458_), .A2(new_n3576_), .B(new_n3577_), .ZN(new_n3578_));
  OAI21_X1   g03386(.A1(new_n3578_), .A2(\asqrt[53] ), .B(new_n3454_), .ZN(new_n3579_));
  NAND2_X1   g03387(.A1(new_n3578_), .A2(\asqrt[53] ), .ZN(new_n3580_));
  NAND3_X1   g03388(.A1(new_n3579_), .A2(new_n3580_), .A3(new_n860_), .ZN(new_n3581_));
  AOI21_X1   g03389(.A1(new_n3579_), .A2(new_n3580_), .B(new_n860_), .ZN(new_n3582_));
  AOI21_X1   g03390(.A1(new_n3452_), .A2(new_n3581_), .B(new_n3582_), .ZN(new_n3583_));
  AOI21_X1   g03391(.A1(new_n3583_), .A2(new_n744_), .B(new_n3450_), .ZN(new_n3584_));
  NAND2_X1   g03392(.A1(new_n3581_), .A2(new_n3452_), .ZN(new_n3585_));
  INV_X1     g03393(.I(new_n3454_), .ZN(new_n3586_));
  INV_X1     g03394(.I(new_n3464_), .ZN(new_n3587_));
  NOR3_X1    g03395(.A1(new_n3571_), .A2(\asqrt[50] ), .A3(new_n3573_), .ZN(new_n3588_));
  OAI21_X1   g03396(.A1(new_n3587_), .A2(new_n3588_), .B(new_n3574_), .ZN(new_n3589_));
  OAI21_X1   g03397(.A1(new_n3589_), .A2(\asqrt[51] ), .B(new_n3461_), .ZN(new_n3590_));
  NAND2_X1   g03398(.A1(new_n3589_), .A2(\asqrt[51] ), .ZN(new_n3591_));
  NAND3_X1   g03399(.A1(new_n3590_), .A2(new_n3591_), .A3(new_n1150_), .ZN(new_n3592_));
  AOI21_X1   g03400(.A1(new_n3590_), .A2(new_n3591_), .B(new_n1150_), .ZN(new_n3593_));
  AOI21_X1   g03401(.A1(new_n3457_), .A2(new_n3592_), .B(new_n3593_), .ZN(new_n3594_));
  AOI21_X1   g03402(.A1(new_n3594_), .A2(new_n1006_), .B(new_n3586_), .ZN(new_n3595_));
  NAND2_X1   g03403(.A1(new_n3592_), .A2(new_n3457_), .ZN(new_n3596_));
  AOI21_X1   g03404(.A1(new_n3596_), .A2(new_n3577_), .B(new_n1006_), .ZN(new_n3597_));
  OAI21_X1   g03405(.A1(new_n3595_), .A2(new_n3597_), .B(\asqrt[54] ), .ZN(new_n3598_));
  AOI21_X1   g03406(.A1(new_n3585_), .A2(new_n3598_), .B(new_n744_), .ZN(new_n3599_));
  NOR3_X1    g03407(.A1(new_n3584_), .A2(\asqrt[56] ), .A3(new_n3599_), .ZN(new_n3600_));
  OAI21_X1   g03408(.A1(new_n3584_), .A2(new_n3599_), .B(\asqrt[56] ), .ZN(new_n3601_));
  OAI21_X1   g03409(.A1(new_n3446_), .A2(new_n3600_), .B(new_n3601_), .ZN(new_n3602_));
  OAI21_X1   g03410(.A1(new_n3602_), .A2(\asqrt[57] ), .B(new_n3441_), .ZN(new_n3603_));
  NOR2_X1    g03411(.A1(new_n3600_), .A2(new_n3446_), .ZN(new_n3604_));
  INV_X1     g03412(.I(new_n3452_), .ZN(new_n3605_));
  NOR3_X1    g03413(.A1(new_n3595_), .A2(\asqrt[54] ), .A3(new_n3597_), .ZN(new_n3606_));
  OAI21_X1   g03414(.A1(new_n3605_), .A2(new_n3606_), .B(new_n3598_), .ZN(new_n3607_));
  OAI21_X1   g03415(.A1(new_n3607_), .A2(\asqrt[55] ), .B(new_n3449_), .ZN(new_n3608_));
  NAND2_X1   g03416(.A1(new_n3607_), .A2(\asqrt[55] ), .ZN(new_n3609_));
  AOI21_X1   g03417(.A1(new_n3608_), .A2(new_n3609_), .B(new_n634_), .ZN(new_n3610_));
  OAI21_X1   g03418(.A1(new_n3604_), .A2(new_n3610_), .B(\asqrt[57] ), .ZN(new_n3611_));
  NAND3_X1   g03419(.A1(new_n3603_), .A2(new_n423_), .A3(new_n3611_), .ZN(new_n3612_));
  NAND2_X1   g03420(.A1(new_n3612_), .A2(new_n3439_), .ZN(new_n3613_));
  INV_X1     g03421(.I(new_n3441_), .ZN(new_n3614_));
  NAND3_X1   g03422(.A1(new_n3608_), .A2(new_n3609_), .A3(new_n634_), .ZN(new_n3615_));
  AOI21_X1   g03423(.A1(new_n3445_), .A2(new_n3615_), .B(new_n3610_), .ZN(new_n3616_));
  AOI21_X1   g03424(.A1(new_n3616_), .A2(new_n531_), .B(new_n3614_), .ZN(new_n3617_));
  NAND2_X1   g03425(.A1(new_n3615_), .A2(new_n3445_), .ZN(new_n3618_));
  AOI21_X1   g03426(.A1(new_n3618_), .A2(new_n3601_), .B(new_n531_), .ZN(new_n3619_));
  OAI21_X1   g03427(.A1(new_n3617_), .A2(new_n3619_), .B(\asqrt[58] ), .ZN(new_n3620_));
  NAND3_X1   g03428(.A1(new_n3613_), .A2(new_n337_), .A3(new_n3620_), .ZN(new_n3621_));
  AOI21_X1   g03429(.A1(new_n3613_), .A2(new_n3620_), .B(new_n337_), .ZN(new_n3622_));
  AOI21_X1   g03430(.A1(new_n3437_), .A2(new_n3621_), .B(new_n3622_), .ZN(new_n3623_));
  AOI21_X1   g03431(.A1(new_n3623_), .A2(new_n266_), .B(new_n3434_), .ZN(new_n3624_));
  INV_X1     g03432(.I(new_n3439_), .ZN(new_n3625_));
  NOR3_X1    g03433(.A1(new_n3617_), .A2(\asqrt[58] ), .A3(new_n3619_), .ZN(new_n3626_));
  OAI21_X1   g03434(.A1(new_n3625_), .A2(new_n3626_), .B(new_n3620_), .ZN(new_n3627_));
  OAI21_X1   g03435(.A1(new_n3627_), .A2(\asqrt[59] ), .B(new_n3437_), .ZN(new_n3628_));
  NAND2_X1   g03436(.A1(new_n3627_), .A2(\asqrt[59] ), .ZN(new_n3629_));
  AOI21_X1   g03437(.A1(new_n3628_), .A2(new_n3629_), .B(new_n266_), .ZN(new_n3630_));
  OAI21_X1   g03438(.A1(new_n3624_), .A2(new_n3630_), .B(\asqrt[61] ), .ZN(new_n3631_));
  AOI21_X1   g03439(.A1(new_n3391_), .A2(new_n3386_), .B(\asqrt[40] ), .ZN(new_n3632_));
  XOR2_X1    g03440(.A1(new_n3632_), .A2(new_n3201_), .Z(new_n3633_));
  INV_X1     g03441(.I(new_n3633_), .ZN(new_n3634_));
  NOR3_X1    g03442(.A1(new_n3624_), .A2(\asqrt[61] ), .A3(new_n3630_), .ZN(new_n3635_));
  OAI21_X1   g03443(.A1(new_n3634_), .A2(new_n3635_), .B(new_n3631_), .ZN(new_n3636_));
  NAND3_X1   g03444(.A1(new_n3628_), .A2(new_n3629_), .A3(new_n266_), .ZN(new_n3637_));
  NAND2_X1   g03445(.A1(new_n3637_), .A2(new_n3433_), .ZN(new_n3638_));
  INV_X1     g03446(.I(new_n3437_), .ZN(new_n3639_));
  AOI21_X1   g03447(.A1(new_n3603_), .A2(new_n3611_), .B(new_n423_), .ZN(new_n3640_));
  AOI21_X1   g03448(.A1(new_n3439_), .A2(new_n3612_), .B(new_n3640_), .ZN(new_n3641_));
  AOI21_X1   g03449(.A1(new_n3641_), .A2(new_n337_), .B(new_n3639_), .ZN(new_n3642_));
  OAI21_X1   g03450(.A1(new_n3642_), .A2(new_n3622_), .B(\asqrt[60] ), .ZN(new_n3643_));
  AOI21_X1   g03451(.A1(new_n3638_), .A2(new_n3643_), .B(new_n239_), .ZN(new_n3644_));
  AOI21_X1   g03452(.A1(new_n3433_), .A2(new_n3637_), .B(new_n3630_), .ZN(new_n3645_));
  AOI21_X1   g03453(.A1(new_n3645_), .A2(new_n239_), .B(new_n3634_), .ZN(new_n3646_));
  OAI21_X1   g03454(.A1(new_n3646_), .A2(new_n3644_), .B(new_n201_), .ZN(new_n3647_));
  NOR3_X1    g03455(.A1(new_n3642_), .A2(\asqrt[60] ), .A3(new_n3622_), .ZN(new_n3648_));
  OAI21_X1   g03456(.A1(new_n3434_), .A2(new_n3648_), .B(new_n3643_), .ZN(new_n3649_));
  OAI21_X1   g03457(.A1(new_n3649_), .A2(\asqrt[61] ), .B(new_n3633_), .ZN(new_n3650_));
  NAND3_X1   g03458(.A1(new_n3650_), .A2(\asqrt[62] ), .A3(new_n3631_), .ZN(new_n3651_));
  AOI21_X1   g03459(.A1(new_n3381_), .A2(new_n3387_), .B(\asqrt[40] ), .ZN(new_n3652_));
  XOR2_X1    g03460(.A1(new_n3652_), .A2(new_n3383_), .Z(new_n3653_));
  INV_X1     g03461(.I(new_n3653_), .ZN(new_n3654_));
  AOI22_X1   g03462(.A1(new_n3651_), .A2(new_n3647_), .B1(new_n3636_), .B2(new_n3654_), .ZN(new_n3655_));
  NOR2_X1    g03463(.A1(new_n3400_), .A2(new_n3198_), .ZN(new_n3656_));
  OAI21_X1   g03464(.A1(\asqrt[40] ), .A2(new_n3656_), .B(new_n3407_), .ZN(new_n3657_));
  INV_X1     g03465(.I(new_n3657_), .ZN(new_n3658_));
  OAI21_X1   g03466(.A1(new_n3655_), .A2(new_n3430_), .B(new_n3658_), .ZN(new_n3659_));
  OAI21_X1   g03467(.A1(new_n3636_), .A2(\asqrt[62] ), .B(new_n3653_), .ZN(new_n3660_));
  NAND2_X1   g03468(.A1(new_n3636_), .A2(\asqrt[62] ), .ZN(new_n3661_));
  NAND3_X1   g03469(.A1(new_n3660_), .A2(new_n3661_), .A3(new_n3430_), .ZN(new_n3662_));
  NAND2_X1   g03470(.A1(new_n3427_), .A2(new_n3197_), .ZN(new_n3663_));
  XOR2_X1    g03471(.A1(new_n3400_), .A2(new_n3198_), .Z(new_n3664_));
  NAND3_X1   g03472(.A1(new_n3663_), .A2(\asqrt[63] ), .A3(new_n3664_), .ZN(new_n3665_));
  INV_X1     g03473(.I(new_n3489_), .ZN(new_n3666_));
  NAND4_X1   g03474(.A1(new_n3666_), .A2(new_n3198_), .A3(new_n3407_), .A4(new_n3414_), .ZN(new_n3667_));
  NAND2_X1   g03475(.A1(new_n3665_), .A2(new_n3667_), .ZN(new_n3668_));
  INV_X1     g03476(.I(new_n3668_), .ZN(new_n3669_));
  NAND4_X1   g03477(.A1(new_n3659_), .A2(new_n193_), .A3(new_n3662_), .A4(new_n3669_), .ZN(\asqrt[39] ));
  NOR2_X1    g03478(.A1(new_n3636_), .A2(\asqrt[62] ), .ZN(new_n3671_));
  NOR2_X1    g03479(.A1(new_n3646_), .A2(new_n3644_), .ZN(new_n3672_));
  NOR2_X1    g03480(.A1(new_n3672_), .A2(new_n201_), .ZN(new_n3673_));
  NOR2_X1    g03481(.A1(new_n3671_), .A2(new_n3673_), .ZN(new_n3674_));
  AOI21_X1   g03482(.A1(new_n3650_), .A2(new_n3631_), .B(\asqrt[62] ), .ZN(new_n3675_));
  NOR3_X1    g03483(.A1(new_n3646_), .A2(new_n201_), .A3(new_n3644_), .ZN(new_n3676_));
  OAI22_X1   g03484(.A1(new_n3675_), .A2(new_n3676_), .B1(new_n3672_), .B2(new_n3653_), .ZN(new_n3677_));
  AOI21_X1   g03485(.A1(new_n3677_), .A2(new_n3429_), .B(new_n3657_), .ZN(new_n3678_));
  AOI21_X1   g03486(.A1(new_n3672_), .A2(new_n201_), .B(new_n3654_), .ZN(new_n3679_));
  NOR3_X1    g03487(.A1(new_n3679_), .A2(new_n3673_), .A3(new_n3429_), .ZN(new_n3680_));
  NOR4_X1    g03488(.A1(new_n3678_), .A2(\asqrt[63] ), .A3(new_n3680_), .A4(new_n3668_), .ZN(new_n3681_));
  XOR2_X1    g03489(.A1(new_n3652_), .A2(new_n3383_), .Z(new_n3682_));
  OAI21_X1   g03490(.A1(\asqrt[39] ), .A2(new_n3674_), .B(new_n3682_), .ZN(new_n3683_));
  INV_X1     g03491(.I(new_n3683_), .ZN(new_n3684_));
  AOI21_X1   g03492(.A1(new_n3621_), .A2(new_n3629_), .B(\asqrt[39] ), .ZN(new_n3685_));
  XOR2_X1    g03493(.A1(new_n3685_), .A2(new_n3437_), .Z(new_n3686_));
  INV_X1     g03494(.I(new_n3686_), .ZN(new_n3687_));
  AOI21_X1   g03495(.A1(new_n3612_), .A2(new_n3620_), .B(\asqrt[39] ), .ZN(new_n3688_));
  XOR2_X1    g03496(.A1(new_n3688_), .A2(new_n3439_), .Z(new_n3689_));
  INV_X1     g03497(.I(new_n3689_), .ZN(new_n3690_));
  NAND2_X1   g03498(.A1(new_n3616_), .A2(new_n531_), .ZN(new_n3691_));
  AOI21_X1   g03499(.A1(new_n3691_), .A2(new_n3611_), .B(\asqrt[39] ), .ZN(new_n3692_));
  XOR2_X1    g03500(.A1(new_n3692_), .A2(new_n3441_), .Z(new_n3693_));
  AOI21_X1   g03501(.A1(new_n3615_), .A2(new_n3601_), .B(\asqrt[39] ), .ZN(new_n3694_));
  XOR2_X1    g03502(.A1(new_n3694_), .A2(new_n3445_), .Z(new_n3695_));
  NAND2_X1   g03503(.A1(new_n3583_), .A2(new_n744_), .ZN(new_n3696_));
  AOI21_X1   g03504(.A1(new_n3696_), .A2(new_n3609_), .B(\asqrt[39] ), .ZN(new_n3697_));
  XOR2_X1    g03505(.A1(new_n3697_), .A2(new_n3449_), .Z(new_n3698_));
  INV_X1     g03506(.I(new_n3698_), .ZN(new_n3699_));
  AOI21_X1   g03507(.A1(new_n3581_), .A2(new_n3598_), .B(\asqrt[39] ), .ZN(new_n3700_));
  XOR2_X1    g03508(.A1(new_n3700_), .A2(new_n3452_), .Z(new_n3701_));
  INV_X1     g03509(.I(new_n3701_), .ZN(new_n3702_));
  NAND2_X1   g03510(.A1(new_n3594_), .A2(new_n1006_), .ZN(new_n3703_));
  AOI21_X1   g03511(.A1(new_n3703_), .A2(new_n3580_), .B(\asqrt[39] ), .ZN(new_n3704_));
  XOR2_X1    g03512(.A1(new_n3704_), .A2(new_n3454_), .Z(new_n3705_));
  AOI21_X1   g03513(.A1(new_n3592_), .A2(new_n3577_), .B(\asqrt[39] ), .ZN(new_n3706_));
  XOR2_X1    g03514(.A1(new_n3706_), .A2(new_n3457_), .Z(new_n3707_));
  NAND2_X1   g03515(.A1(new_n3559_), .A2(new_n1305_), .ZN(new_n3708_));
  AOI21_X1   g03516(.A1(new_n3708_), .A2(new_n3591_), .B(\asqrt[39] ), .ZN(new_n3709_));
  XOR2_X1    g03517(.A1(new_n3709_), .A2(new_n3461_), .Z(new_n3710_));
  INV_X1     g03518(.I(new_n3710_), .ZN(new_n3711_));
  AOI21_X1   g03519(.A1(new_n3557_), .A2(new_n3574_), .B(\asqrt[39] ), .ZN(new_n3712_));
  XOR2_X1    g03520(.A1(new_n3712_), .A2(new_n3464_), .Z(new_n3713_));
  INV_X1     g03521(.I(new_n3713_), .ZN(new_n3714_));
  NAND2_X1   g03522(.A1(new_n3570_), .A2(new_n1632_), .ZN(new_n3715_));
  AOI21_X1   g03523(.A1(new_n3715_), .A2(new_n3556_), .B(\asqrt[39] ), .ZN(new_n3716_));
  XOR2_X1    g03524(.A1(new_n3716_), .A2(new_n3466_), .Z(new_n3717_));
  AOI21_X1   g03525(.A1(new_n3568_), .A2(new_n3553_), .B(\asqrt[39] ), .ZN(new_n3718_));
  XOR2_X1    g03526(.A1(new_n3718_), .A2(new_n3469_), .Z(new_n3719_));
  NAND2_X1   g03527(.A1(new_n3536_), .A2(new_n1953_), .ZN(new_n3720_));
  AOI21_X1   g03528(.A1(new_n3720_), .A2(new_n3567_), .B(\asqrt[39] ), .ZN(new_n3721_));
  XOR2_X1    g03529(.A1(new_n3721_), .A2(new_n3473_), .Z(new_n3722_));
  INV_X1     g03530(.I(new_n3722_), .ZN(new_n3723_));
  AOI21_X1   g03531(.A1(new_n3534_), .A2(new_n3550_), .B(\asqrt[39] ), .ZN(new_n3724_));
  XOR2_X1    g03532(.A1(new_n3724_), .A2(new_n3476_), .Z(new_n3725_));
  INV_X1     g03533(.I(new_n3725_), .ZN(new_n3726_));
  NAND2_X1   g03534(.A1(new_n3546_), .A2(new_n2332_), .ZN(new_n3727_));
  AOI21_X1   g03535(.A1(new_n3727_), .A2(new_n3533_), .B(\asqrt[39] ), .ZN(new_n3728_));
  XOR2_X1    g03536(.A1(new_n3728_), .A2(new_n3478_), .Z(new_n3729_));
  AOI21_X1   g03537(.A1(new_n3544_), .A2(new_n3530_), .B(\asqrt[39] ), .ZN(new_n3730_));
  XOR2_X1    g03538(.A1(new_n3730_), .A2(new_n3480_), .Z(new_n3731_));
  NAND2_X1   g03539(.A1(new_n3517_), .A2(new_n2749_), .ZN(new_n3732_));
  AOI21_X1   g03540(.A1(new_n3732_), .A2(new_n3543_), .B(\asqrt[39] ), .ZN(new_n3733_));
  XOR2_X1    g03541(.A1(new_n3733_), .A2(new_n3487_), .Z(new_n3734_));
  INV_X1     g03542(.I(new_n3734_), .ZN(new_n3735_));
  AOI21_X1   g03543(.A1(new_n3515_), .A2(new_n3527_), .B(\asqrt[39] ), .ZN(new_n3736_));
  XOR2_X1    g03544(.A1(new_n3736_), .A2(new_n3499_), .Z(new_n3737_));
  INV_X1     g03545(.I(new_n3737_), .ZN(new_n3738_));
  NAND2_X1   g03546(.A1(\asqrt[40] ), .A2(new_n3500_), .ZN(new_n3739_));
  NOR2_X1    g03547(.A1(new_n3512_), .A2(\a[80] ), .ZN(new_n3740_));
  AOI22_X1   g03548(.A1(new_n3739_), .A2(new_n3512_), .B1(\asqrt[40] ), .B2(new_n3740_), .ZN(new_n3741_));
  AOI21_X1   g03549(.A1(\asqrt[40] ), .A2(\a[80] ), .B(new_n3508_), .ZN(new_n3742_));
  OAI21_X1   g03550(.A1(new_n3522_), .A2(new_n3742_), .B(new_n3681_), .ZN(new_n3743_));
  XNOR2_X1   g03551(.A1(new_n3743_), .A2(new_n3741_), .ZN(new_n3744_));
  NAND3_X1   g03552(.A1(new_n3665_), .A2(\asqrt[40] ), .A3(new_n3667_), .ZN(new_n3745_));
  NOR4_X1    g03553(.A1(new_n3678_), .A2(\asqrt[63] ), .A3(new_n3680_), .A4(new_n3745_), .ZN(new_n3746_));
  INV_X1     g03554(.I(new_n3746_), .ZN(new_n3747_));
  NAND2_X1   g03555(.A1(\asqrt[39] ), .A2(new_n3501_), .ZN(new_n3748_));
  AOI21_X1   g03556(.A1(new_n3748_), .A2(new_n3747_), .B(\a[80] ), .ZN(new_n3749_));
  NOR2_X1    g03557(.A1(new_n3681_), .A2(new_n3503_), .ZN(new_n3750_));
  NOR3_X1    g03558(.A1(new_n3750_), .A2(new_n3500_), .A3(new_n3746_), .ZN(new_n3751_));
  NOR2_X1    g03559(.A1(new_n3751_), .A2(new_n3749_), .ZN(new_n3752_));
  INV_X1     g03560(.I(\a[78] ), .ZN(new_n3753_));
  NOR2_X1    g03561(.A1(\a[76] ), .A2(\a[77] ), .ZN(new_n3754_));
  NOR3_X1    g03562(.A1(new_n3681_), .A2(new_n3753_), .A3(new_n3754_), .ZN(new_n3755_));
  INV_X1     g03563(.I(new_n3754_), .ZN(new_n3756_));
  AOI21_X1   g03564(.A1(new_n3681_), .A2(\a[78] ), .B(new_n3756_), .ZN(new_n3757_));
  OAI21_X1   g03565(.A1(new_n3755_), .A2(new_n3757_), .B(\asqrt[40] ), .ZN(new_n3758_));
  NAND2_X1   g03566(.A1(new_n3754_), .A2(new_n3753_), .ZN(new_n3759_));
  NAND3_X1   g03567(.A1(new_n3410_), .A2(new_n3412_), .A3(new_n3759_), .ZN(new_n3760_));
  NAND2_X1   g03568(.A1(new_n3494_), .A2(new_n3760_), .ZN(new_n3761_));
  NAND3_X1   g03569(.A1(\asqrt[39] ), .A2(\a[78] ), .A3(new_n3761_), .ZN(new_n3762_));
  NOR3_X1    g03570(.A1(new_n3681_), .A2(\a[78] ), .A3(\a[79] ), .ZN(new_n3763_));
  INV_X1     g03571(.I(\a[79] ), .ZN(new_n3764_));
  AOI21_X1   g03572(.A1(\asqrt[39] ), .A2(new_n3753_), .B(new_n3764_), .ZN(new_n3765_));
  NOR2_X1    g03573(.A1(new_n3763_), .A2(new_n3765_), .ZN(new_n3766_));
  NAND4_X1   g03574(.A1(new_n3758_), .A2(new_n3766_), .A3(new_n3195_), .A4(new_n3762_), .ZN(new_n3767_));
  NAND2_X1   g03575(.A1(new_n3767_), .A2(new_n3752_), .ZN(new_n3768_));
  NAND3_X1   g03576(.A1(\asqrt[39] ), .A2(\a[78] ), .A3(new_n3756_), .ZN(new_n3769_));
  OAI21_X1   g03577(.A1(\asqrt[39] ), .A2(new_n3753_), .B(new_n3754_), .ZN(new_n3770_));
  AOI21_X1   g03578(.A1(new_n3770_), .A2(new_n3769_), .B(new_n3427_), .ZN(new_n3771_));
  NAND3_X1   g03579(.A1(\asqrt[39] ), .A2(new_n3753_), .A3(new_n3764_), .ZN(new_n3772_));
  OAI21_X1   g03580(.A1(new_n3681_), .A2(\a[78] ), .B(\a[79] ), .ZN(new_n3773_));
  NAND3_X1   g03581(.A1(new_n3762_), .A2(new_n3773_), .A3(new_n3772_), .ZN(new_n3774_));
  OAI21_X1   g03582(.A1(new_n3774_), .A2(new_n3771_), .B(\asqrt[41] ), .ZN(new_n3775_));
  NAND3_X1   g03583(.A1(new_n3768_), .A2(new_n2960_), .A3(new_n3775_), .ZN(new_n3776_));
  AOI21_X1   g03584(.A1(new_n3768_), .A2(new_n3775_), .B(new_n2960_), .ZN(new_n3777_));
  AOI21_X1   g03585(.A1(new_n3744_), .A2(new_n3776_), .B(new_n3777_), .ZN(new_n3778_));
  AOI21_X1   g03586(.A1(new_n3778_), .A2(new_n2749_), .B(new_n3738_), .ZN(new_n3779_));
  OR2_X2     g03587(.A1(new_n3751_), .A2(new_n3749_), .Z(new_n3780_));
  NOR3_X1    g03588(.A1(new_n3774_), .A2(new_n3771_), .A3(\asqrt[41] ), .ZN(new_n3781_));
  OAI21_X1   g03589(.A1(new_n3780_), .A2(new_n3781_), .B(new_n3775_), .ZN(new_n3782_));
  OAI21_X1   g03590(.A1(new_n3782_), .A2(\asqrt[42] ), .B(new_n3744_), .ZN(new_n3783_));
  NAND2_X1   g03591(.A1(new_n3782_), .A2(\asqrt[42] ), .ZN(new_n3784_));
  AOI21_X1   g03592(.A1(new_n3783_), .A2(new_n3784_), .B(new_n2749_), .ZN(new_n3785_));
  NOR3_X1    g03593(.A1(new_n3779_), .A2(\asqrt[44] ), .A3(new_n3785_), .ZN(new_n3786_));
  OAI21_X1   g03594(.A1(new_n3779_), .A2(new_n3785_), .B(\asqrt[44] ), .ZN(new_n3787_));
  OAI21_X1   g03595(.A1(new_n3735_), .A2(new_n3786_), .B(new_n3787_), .ZN(new_n3788_));
  OAI21_X1   g03596(.A1(new_n3788_), .A2(\asqrt[45] ), .B(new_n3731_), .ZN(new_n3789_));
  NAND3_X1   g03597(.A1(new_n3783_), .A2(new_n3784_), .A3(new_n2749_), .ZN(new_n3790_));
  AOI21_X1   g03598(.A1(new_n3737_), .A2(new_n3790_), .B(new_n3785_), .ZN(new_n3791_));
  AOI21_X1   g03599(.A1(new_n3791_), .A2(new_n2531_), .B(new_n3735_), .ZN(new_n3792_));
  NAND2_X1   g03600(.A1(new_n3790_), .A2(new_n3737_), .ZN(new_n3793_));
  INV_X1     g03601(.I(new_n3785_), .ZN(new_n3794_));
  AOI21_X1   g03602(.A1(new_n3793_), .A2(new_n3794_), .B(new_n2531_), .ZN(new_n3795_));
  OAI21_X1   g03603(.A1(new_n3792_), .A2(new_n3795_), .B(\asqrt[45] ), .ZN(new_n3796_));
  NAND3_X1   g03604(.A1(new_n3789_), .A2(new_n2134_), .A3(new_n3796_), .ZN(new_n3797_));
  AOI21_X1   g03605(.A1(new_n3789_), .A2(new_n3796_), .B(new_n2134_), .ZN(new_n3798_));
  AOI21_X1   g03606(.A1(new_n3729_), .A2(new_n3797_), .B(new_n3798_), .ZN(new_n3799_));
  AOI21_X1   g03607(.A1(new_n3799_), .A2(new_n1953_), .B(new_n3726_), .ZN(new_n3800_));
  INV_X1     g03608(.I(new_n3731_), .ZN(new_n3801_));
  NOR3_X1    g03609(.A1(new_n3792_), .A2(\asqrt[45] ), .A3(new_n3795_), .ZN(new_n3802_));
  OAI21_X1   g03610(.A1(new_n3801_), .A2(new_n3802_), .B(new_n3796_), .ZN(new_n3803_));
  OAI21_X1   g03611(.A1(new_n3803_), .A2(\asqrt[46] ), .B(new_n3729_), .ZN(new_n3804_));
  NAND2_X1   g03612(.A1(new_n3803_), .A2(\asqrt[46] ), .ZN(new_n3805_));
  AOI21_X1   g03613(.A1(new_n3804_), .A2(new_n3805_), .B(new_n1953_), .ZN(new_n3806_));
  NOR3_X1    g03614(.A1(new_n3800_), .A2(\asqrt[48] ), .A3(new_n3806_), .ZN(new_n3807_));
  OAI21_X1   g03615(.A1(new_n3800_), .A2(new_n3806_), .B(\asqrt[48] ), .ZN(new_n3808_));
  OAI21_X1   g03616(.A1(new_n3723_), .A2(new_n3807_), .B(new_n3808_), .ZN(new_n3809_));
  OAI21_X1   g03617(.A1(new_n3809_), .A2(\asqrt[49] ), .B(new_n3719_), .ZN(new_n3810_));
  NAND3_X1   g03618(.A1(new_n3804_), .A2(new_n3805_), .A3(new_n1953_), .ZN(new_n3811_));
  AOI21_X1   g03619(.A1(new_n3725_), .A2(new_n3811_), .B(new_n3806_), .ZN(new_n3812_));
  AOI21_X1   g03620(.A1(new_n3812_), .A2(new_n1778_), .B(new_n3723_), .ZN(new_n3813_));
  NAND2_X1   g03621(.A1(new_n3811_), .A2(new_n3725_), .ZN(new_n3814_));
  INV_X1     g03622(.I(new_n3806_), .ZN(new_n3815_));
  AOI21_X1   g03623(.A1(new_n3814_), .A2(new_n3815_), .B(new_n1778_), .ZN(new_n3816_));
  OAI21_X1   g03624(.A1(new_n3813_), .A2(new_n3816_), .B(\asqrt[49] ), .ZN(new_n3817_));
  NAND3_X1   g03625(.A1(new_n3810_), .A2(new_n1463_), .A3(new_n3817_), .ZN(new_n3818_));
  AOI21_X1   g03626(.A1(new_n3810_), .A2(new_n3817_), .B(new_n1463_), .ZN(new_n3819_));
  AOI21_X1   g03627(.A1(new_n3717_), .A2(new_n3818_), .B(new_n3819_), .ZN(new_n3820_));
  AOI21_X1   g03628(.A1(new_n3820_), .A2(new_n1305_), .B(new_n3714_), .ZN(new_n3821_));
  INV_X1     g03629(.I(new_n3719_), .ZN(new_n3822_));
  NOR3_X1    g03630(.A1(new_n3813_), .A2(\asqrt[49] ), .A3(new_n3816_), .ZN(new_n3823_));
  OAI21_X1   g03631(.A1(new_n3822_), .A2(new_n3823_), .B(new_n3817_), .ZN(new_n3824_));
  OAI21_X1   g03632(.A1(new_n3824_), .A2(\asqrt[50] ), .B(new_n3717_), .ZN(new_n3825_));
  NAND2_X1   g03633(.A1(new_n3824_), .A2(\asqrt[50] ), .ZN(new_n3826_));
  AOI21_X1   g03634(.A1(new_n3825_), .A2(new_n3826_), .B(new_n1305_), .ZN(new_n3827_));
  NOR3_X1    g03635(.A1(new_n3821_), .A2(\asqrt[52] ), .A3(new_n3827_), .ZN(new_n3828_));
  OAI21_X1   g03636(.A1(new_n3821_), .A2(new_n3827_), .B(\asqrt[52] ), .ZN(new_n3829_));
  OAI21_X1   g03637(.A1(new_n3711_), .A2(new_n3828_), .B(new_n3829_), .ZN(new_n3830_));
  OAI21_X1   g03638(.A1(new_n3830_), .A2(\asqrt[53] ), .B(new_n3707_), .ZN(new_n3831_));
  NAND3_X1   g03639(.A1(new_n3825_), .A2(new_n3826_), .A3(new_n1305_), .ZN(new_n3832_));
  AOI21_X1   g03640(.A1(new_n3713_), .A2(new_n3832_), .B(new_n3827_), .ZN(new_n3833_));
  AOI21_X1   g03641(.A1(new_n3833_), .A2(new_n1150_), .B(new_n3711_), .ZN(new_n3834_));
  NAND2_X1   g03642(.A1(new_n3832_), .A2(new_n3713_), .ZN(new_n3835_));
  INV_X1     g03643(.I(new_n3827_), .ZN(new_n3836_));
  AOI21_X1   g03644(.A1(new_n3835_), .A2(new_n3836_), .B(new_n1150_), .ZN(new_n3837_));
  OAI21_X1   g03645(.A1(new_n3834_), .A2(new_n3837_), .B(\asqrt[53] ), .ZN(new_n3838_));
  NAND3_X1   g03646(.A1(new_n3831_), .A2(new_n860_), .A3(new_n3838_), .ZN(new_n3839_));
  AOI21_X1   g03647(.A1(new_n3831_), .A2(new_n3838_), .B(new_n860_), .ZN(new_n3840_));
  AOI21_X1   g03648(.A1(new_n3705_), .A2(new_n3839_), .B(new_n3840_), .ZN(new_n3841_));
  AOI21_X1   g03649(.A1(new_n3841_), .A2(new_n744_), .B(new_n3702_), .ZN(new_n3842_));
  INV_X1     g03650(.I(new_n3707_), .ZN(new_n3843_));
  NOR3_X1    g03651(.A1(new_n3834_), .A2(\asqrt[53] ), .A3(new_n3837_), .ZN(new_n3844_));
  OAI21_X1   g03652(.A1(new_n3843_), .A2(new_n3844_), .B(new_n3838_), .ZN(new_n3845_));
  OAI21_X1   g03653(.A1(new_n3845_), .A2(\asqrt[54] ), .B(new_n3705_), .ZN(new_n3846_));
  NAND2_X1   g03654(.A1(new_n3845_), .A2(\asqrt[54] ), .ZN(new_n3847_));
  AOI21_X1   g03655(.A1(new_n3846_), .A2(new_n3847_), .B(new_n744_), .ZN(new_n3848_));
  NOR3_X1    g03656(.A1(new_n3842_), .A2(\asqrt[56] ), .A3(new_n3848_), .ZN(new_n3849_));
  OAI21_X1   g03657(.A1(new_n3842_), .A2(new_n3848_), .B(\asqrt[56] ), .ZN(new_n3850_));
  OAI21_X1   g03658(.A1(new_n3699_), .A2(new_n3849_), .B(new_n3850_), .ZN(new_n3851_));
  OAI21_X1   g03659(.A1(new_n3851_), .A2(\asqrt[57] ), .B(new_n3695_), .ZN(new_n3852_));
  NAND3_X1   g03660(.A1(new_n3846_), .A2(new_n3847_), .A3(new_n744_), .ZN(new_n3853_));
  AOI21_X1   g03661(.A1(new_n3701_), .A2(new_n3853_), .B(new_n3848_), .ZN(new_n3854_));
  AOI21_X1   g03662(.A1(new_n3854_), .A2(new_n634_), .B(new_n3699_), .ZN(new_n3855_));
  NAND2_X1   g03663(.A1(new_n3853_), .A2(new_n3701_), .ZN(new_n3856_));
  INV_X1     g03664(.I(new_n3848_), .ZN(new_n3857_));
  AOI21_X1   g03665(.A1(new_n3856_), .A2(new_n3857_), .B(new_n634_), .ZN(new_n3858_));
  OAI21_X1   g03666(.A1(new_n3855_), .A2(new_n3858_), .B(\asqrt[57] ), .ZN(new_n3859_));
  NAND3_X1   g03667(.A1(new_n3852_), .A2(new_n423_), .A3(new_n3859_), .ZN(new_n3860_));
  AOI21_X1   g03668(.A1(new_n3852_), .A2(new_n3859_), .B(new_n423_), .ZN(new_n3861_));
  AOI21_X1   g03669(.A1(new_n3693_), .A2(new_n3860_), .B(new_n3861_), .ZN(new_n3862_));
  AOI21_X1   g03670(.A1(new_n3862_), .A2(new_n337_), .B(new_n3690_), .ZN(new_n3863_));
  NOR2_X1    g03671(.A1(new_n3862_), .A2(new_n337_), .ZN(new_n3864_));
  NOR3_X1    g03672(.A1(new_n3863_), .A2(new_n3864_), .A3(\asqrt[60] ), .ZN(new_n3865_));
  OAI21_X1   g03673(.A1(new_n3863_), .A2(new_n3864_), .B(\asqrt[60] ), .ZN(new_n3866_));
  OAI21_X1   g03674(.A1(new_n3687_), .A2(new_n3865_), .B(new_n3866_), .ZN(new_n3867_));
  NAND2_X1   g03675(.A1(new_n3867_), .A2(\asqrt[61] ), .ZN(new_n3868_));
  AOI21_X1   g03676(.A1(new_n3637_), .A2(new_n3643_), .B(\asqrt[39] ), .ZN(new_n3869_));
  XOR2_X1    g03677(.A1(new_n3869_), .A2(new_n3433_), .Z(new_n3870_));
  OAI21_X1   g03678(.A1(new_n3867_), .A2(\asqrt[61] ), .B(new_n3870_), .ZN(new_n3871_));
  NAND2_X1   g03679(.A1(new_n3871_), .A2(new_n3868_), .ZN(new_n3872_));
  INV_X1     g03680(.I(new_n3695_), .ZN(new_n3873_));
  NOR3_X1    g03681(.A1(new_n3855_), .A2(\asqrt[57] ), .A3(new_n3858_), .ZN(new_n3874_));
  OAI21_X1   g03682(.A1(new_n3873_), .A2(new_n3874_), .B(new_n3859_), .ZN(new_n3875_));
  OAI21_X1   g03683(.A1(new_n3875_), .A2(\asqrt[58] ), .B(new_n3693_), .ZN(new_n3876_));
  NOR2_X1    g03684(.A1(new_n3874_), .A2(new_n3873_), .ZN(new_n3877_));
  INV_X1     g03685(.I(new_n3859_), .ZN(new_n3878_));
  OAI21_X1   g03686(.A1(new_n3877_), .A2(new_n3878_), .B(\asqrt[58] ), .ZN(new_n3879_));
  NAND3_X1   g03687(.A1(new_n3876_), .A2(new_n337_), .A3(new_n3879_), .ZN(new_n3880_));
  NAND2_X1   g03688(.A1(new_n3880_), .A2(new_n3689_), .ZN(new_n3881_));
  INV_X1     g03689(.I(new_n3693_), .ZN(new_n3882_));
  NOR2_X1    g03690(.A1(new_n3877_), .A2(new_n3878_), .ZN(new_n3883_));
  AOI21_X1   g03691(.A1(new_n3883_), .A2(new_n423_), .B(new_n3882_), .ZN(new_n3884_));
  OAI21_X1   g03692(.A1(new_n3884_), .A2(new_n3861_), .B(\asqrt[59] ), .ZN(new_n3885_));
  NAND3_X1   g03693(.A1(new_n3881_), .A2(new_n266_), .A3(new_n3885_), .ZN(new_n3886_));
  NAND2_X1   g03694(.A1(new_n3886_), .A2(new_n3686_), .ZN(new_n3887_));
  AOI21_X1   g03695(.A1(new_n3887_), .A2(new_n3866_), .B(new_n239_), .ZN(new_n3888_));
  AOI21_X1   g03696(.A1(new_n3881_), .A2(new_n3885_), .B(new_n266_), .ZN(new_n3889_));
  AOI21_X1   g03697(.A1(new_n3686_), .A2(new_n3886_), .B(new_n3889_), .ZN(new_n3890_));
  INV_X1     g03698(.I(new_n3870_), .ZN(new_n3891_));
  AOI21_X1   g03699(.A1(new_n3890_), .A2(new_n239_), .B(new_n3891_), .ZN(new_n3892_));
  OAI21_X1   g03700(.A1(new_n3892_), .A2(new_n3888_), .B(new_n201_), .ZN(new_n3893_));
  NAND3_X1   g03701(.A1(new_n3871_), .A2(new_n3868_), .A3(\asqrt[62] ), .ZN(new_n3894_));
  NOR2_X1    g03702(.A1(new_n3635_), .A2(new_n3644_), .ZN(new_n3895_));
  NOR2_X1    g03703(.A1(\asqrt[39] ), .A2(new_n3895_), .ZN(new_n3896_));
  XOR2_X1    g03704(.A1(new_n3896_), .A2(new_n3633_), .Z(new_n3897_));
  INV_X1     g03705(.I(new_n3897_), .ZN(new_n3898_));
  AOI22_X1   g03706(.A1(new_n3894_), .A2(new_n3893_), .B1(new_n3872_), .B2(new_n3898_), .ZN(new_n3899_));
  NOR2_X1    g03707(.A1(new_n3655_), .A2(new_n3430_), .ZN(new_n3900_));
  OAI21_X1   g03708(.A1(\asqrt[39] ), .A2(new_n3900_), .B(new_n3662_), .ZN(new_n3901_));
  INV_X1     g03709(.I(new_n3901_), .ZN(new_n3902_));
  OAI21_X1   g03710(.A1(new_n3899_), .A2(new_n3684_), .B(new_n3902_), .ZN(new_n3903_));
  OAI21_X1   g03711(.A1(new_n3872_), .A2(\asqrt[62] ), .B(new_n3897_), .ZN(new_n3904_));
  NAND2_X1   g03712(.A1(new_n3872_), .A2(\asqrt[62] ), .ZN(new_n3905_));
  NAND3_X1   g03713(.A1(new_n3904_), .A2(new_n3905_), .A3(new_n3684_), .ZN(new_n3906_));
  NAND2_X1   g03714(.A1(new_n3681_), .A2(new_n3429_), .ZN(new_n3907_));
  XOR2_X1    g03715(.A1(new_n3677_), .A2(new_n3429_), .Z(new_n3908_));
  NAND3_X1   g03716(.A1(new_n3907_), .A2(\asqrt[63] ), .A3(new_n3908_), .ZN(new_n3909_));
  NOR2_X1    g03717(.A1(new_n3668_), .A2(new_n3429_), .ZN(new_n3910_));
  NAND4_X1   g03718(.A1(new_n3659_), .A2(new_n193_), .A3(new_n3662_), .A4(new_n3910_), .ZN(new_n3911_));
  NAND2_X1   g03719(.A1(new_n3909_), .A2(new_n3911_), .ZN(new_n3912_));
  INV_X1     g03720(.I(new_n3912_), .ZN(new_n3913_));
  NAND4_X1   g03721(.A1(new_n3903_), .A2(new_n193_), .A3(new_n3906_), .A4(new_n3913_), .ZN(\asqrt[38] ));
  NOR2_X1    g03722(.A1(new_n3872_), .A2(\asqrt[62] ), .ZN(new_n3915_));
  NOR2_X1    g03723(.A1(new_n3892_), .A2(new_n3888_), .ZN(new_n3916_));
  NOR2_X1    g03724(.A1(new_n3916_), .A2(new_n201_), .ZN(new_n3917_));
  NOR2_X1    g03725(.A1(new_n3915_), .A2(new_n3917_), .ZN(new_n3918_));
  AOI21_X1   g03726(.A1(new_n3871_), .A2(new_n3868_), .B(\asqrt[62] ), .ZN(new_n3919_));
  NOR3_X1    g03727(.A1(new_n3892_), .A2(new_n201_), .A3(new_n3888_), .ZN(new_n3920_));
  OAI22_X1   g03728(.A1(new_n3919_), .A2(new_n3920_), .B1(new_n3916_), .B2(new_n3897_), .ZN(new_n3921_));
  AOI21_X1   g03729(.A1(new_n3921_), .A2(new_n3683_), .B(new_n3901_), .ZN(new_n3922_));
  AOI21_X1   g03730(.A1(new_n3916_), .A2(new_n201_), .B(new_n3898_), .ZN(new_n3923_));
  NOR3_X1    g03731(.A1(new_n3923_), .A2(new_n3917_), .A3(new_n3683_), .ZN(new_n3924_));
  NOR4_X1    g03732(.A1(new_n3922_), .A2(\asqrt[63] ), .A3(new_n3924_), .A4(new_n3912_), .ZN(new_n3925_));
  XOR2_X1    g03733(.A1(new_n3896_), .A2(new_n3633_), .Z(new_n3926_));
  OAI21_X1   g03734(.A1(\asqrt[38] ), .A2(new_n3918_), .B(new_n3926_), .ZN(new_n3927_));
  INV_X1     g03735(.I(new_n3927_), .ZN(new_n3928_));
  AOI21_X1   g03736(.A1(new_n3880_), .A2(new_n3885_), .B(\asqrt[38] ), .ZN(new_n3929_));
  XOR2_X1    g03737(.A1(new_n3929_), .A2(new_n3689_), .Z(new_n3930_));
  INV_X1     g03738(.I(new_n3930_), .ZN(new_n3931_));
  AOI21_X1   g03739(.A1(new_n3860_), .A2(new_n3879_), .B(\asqrt[38] ), .ZN(new_n3932_));
  XOR2_X1    g03740(.A1(new_n3932_), .A2(new_n3693_), .Z(new_n3933_));
  INV_X1     g03741(.I(new_n3933_), .ZN(new_n3934_));
  NOR2_X1    g03742(.A1(new_n3878_), .A2(new_n3874_), .ZN(new_n3935_));
  NOR2_X1    g03743(.A1(\asqrt[38] ), .A2(new_n3935_), .ZN(new_n3936_));
  XOR2_X1    g03744(.A1(new_n3936_), .A2(new_n3695_), .Z(new_n3937_));
  NOR2_X1    g03745(.A1(new_n3849_), .A2(new_n3858_), .ZN(new_n3938_));
  NOR2_X1    g03746(.A1(\asqrt[38] ), .A2(new_n3938_), .ZN(new_n3939_));
  XOR2_X1    g03747(.A1(new_n3939_), .A2(new_n3698_), .Z(new_n3940_));
  AOI21_X1   g03748(.A1(new_n3853_), .A2(new_n3857_), .B(\asqrt[38] ), .ZN(new_n3941_));
  XOR2_X1    g03749(.A1(new_n3941_), .A2(new_n3701_), .Z(new_n3942_));
  INV_X1     g03750(.I(new_n3942_), .ZN(new_n3943_));
  AOI21_X1   g03751(.A1(new_n3839_), .A2(new_n3847_), .B(\asqrt[38] ), .ZN(new_n3944_));
  XOR2_X1    g03752(.A1(new_n3944_), .A2(new_n3705_), .Z(new_n3945_));
  INV_X1     g03753(.I(new_n3945_), .ZN(new_n3946_));
  XOR2_X1    g03754(.A1(new_n3830_), .A2(\asqrt[53] ), .Z(new_n3947_));
  NOR2_X1    g03755(.A1(\asqrt[38] ), .A2(new_n3947_), .ZN(new_n3948_));
  XOR2_X1    g03756(.A1(new_n3948_), .A2(new_n3707_), .Z(new_n3949_));
  NOR2_X1    g03757(.A1(new_n3828_), .A2(new_n3837_), .ZN(new_n3950_));
  NOR2_X1    g03758(.A1(\asqrt[38] ), .A2(new_n3950_), .ZN(new_n3951_));
  XOR2_X1    g03759(.A1(new_n3951_), .A2(new_n3710_), .Z(new_n3952_));
  AOI21_X1   g03760(.A1(new_n3832_), .A2(new_n3836_), .B(\asqrt[38] ), .ZN(new_n3953_));
  XOR2_X1    g03761(.A1(new_n3953_), .A2(new_n3713_), .Z(new_n3954_));
  INV_X1     g03762(.I(new_n3954_), .ZN(new_n3955_));
  AOI21_X1   g03763(.A1(new_n3818_), .A2(new_n3826_), .B(\asqrt[38] ), .ZN(new_n3956_));
  XOR2_X1    g03764(.A1(new_n3956_), .A2(new_n3717_), .Z(new_n3957_));
  INV_X1     g03765(.I(new_n3957_), .ZN(new_n3958_));
  XOR2_X1    g03766(.A1(new_n3809_), .A2(\asqrt[49] ), .Z(new_n3959_));
  NOR2_X1    g03767(.A1(\asqrt[38] ), .A2(new_n3959_), .ZN(new_n3960_));
  XOR2_X1    g03768(.A1(new_n3960_), .A2(new_n3719_), .Z(new_n3961_));
  NOR2_X1    g03769(.A1(new_n3807_), .A2(new_n3816_), .ZN(new_n3962_));
  NOR2_X1    g03770(.A1(\asqrt[38] ), .A2(new_n3962_), .ZN(new_n3963_));
  XOR2_X1    g03771(.A1(new_n3963_), .A2(new_n3722_), .Z(new_n3964_));
  AOI21_X1   g03772(.A1(new_n3811_), .A2(new_n3815_), .B(\asqrt[38] ), .ZN(new_n3965_));
  XOR2_X1    g03773(.A1(new_n3965_), .A2(new_n3725_), .Z(new_n3966_));
  INV_X1     g03774(.I(new_n3966_), .ZN(new_n3967_));
  AOI21_X1   g03775(.A1(new_n3797_), .A2(new_n3805_), .B(\asqrt[38] ), .ZN(new_n3968_));
  XOR2_X1    g03776(.A1(new_n3968_), .A2(new_n3729_), .Z(new_n3969_));
  INV_X1     g03777(.I(new_n3969_), .ZN(new_n3970_));
  XOR2_X1    g03778(.A1(new_n3788_), .A2(\asqrt[45] ), .Z(new_n3971_));
  NOR2_X1    g03779(.A1(\asqrt[38] ), .A2(new_n3971_), .ZN(new_n3972_));
  XOR2_X1    g03780(.A1(new_n3972_), .A2(new_n3731_), .Z(new_n3973_));
  NOR2_X1    g03781(.A1(new_n3786_), .A2(new_n3795_), .ZN(new_n3974_));
  NOR2_X1    g03782(.A1(\asqrt[38] ), .A2(new_n3974_), .ZN(new_n3975_));
  XOR2_X1    g03783(.A1(new_n3975_), .A2(new_n3734_), .Z(new_n3976_));
  AOI21_X1   g03784(.A1(new_n3790_), .A2(new_n3794_), .B(\asqrt[38] ), .ZN(new_n3977_));
  XOR2_X1    g03785(.A1(new_n3977_), .A2(new_n3737_), .Z(new_n3978_));
  INV_X1     g03786(.I(new_n3978_), .ZN(new_n3979_));
  AOI21_X1   g03787(.A1(new_n3776_), .A2(new_n3784_), .B(\asqrt[38] ), .ZN(new_n3980_));
  XOR2_X1    g03788(.A1(new_n3980_), .A2(new_n3744_), .Z(new_n3981_));
  INV_X1     g03789(.I(new_n3981_), .ZN(new_n3982_));
  AOI21_X1   g03790(.A1(new_n3767_), .A2(new_n3775_), .B(\asqrt[38] ), .ZN(new_n3983_));
  XOR2_X1    g03791(.A1(new_n3983_), .A2(new_n3752_), .Z(new_n3984_));
  NAND2_X1   g03792(.A1(\asqrt[39] ), .A2(new_n3753_), .ZN(new_n3985_));
  NOR2_X1    g03793(.A1(new_n3764_), .A2(\a[78] ), .ZN(new_n3986_));
  AOI22_X1   g03794(.A1(new_n3985_), .A2(new_n3764_), .B1(\asqrt[39] ), .B2(new_n3986_), .ZN(new_n3987_));
  AOI21_X1   g03795(.A1(\asqrt[39] ), .A2(\a[78] ), .B(new_n3761_), .ZN(new_n3988_));
  OAI21_X1   g03796(.A1(new_n3771_), .A2(new_n3988_), .B(new_n3925_), .ZN(new_n3989_));
  XNOR2_X1   g03797(.A1(new_n3989_), .A2(new_n3987_), .ZN(new_n3990_));
  NOR3_X1    g03798(.A1(new_n3922_), .A2(\asqrt[63] ), .A3(new_n3924_), .ZN(new_n3991_));
  NAND4_X1   g03799(.A1(new_n3991_), .A2(\asqrt[39] ), .A3(new_n3909_), .A4(new_n3911_), .ZN(new_n3992_));
  NAND2_X1   g03800(.A1(\asqrt[38] ), .A2(new_n3754_), .ZN(new_n3993_));
  AOI21_X1   g03801(.A1(new_n3992_), .A2(new_n3993_), .B(\a[78] ), .ZN(new_n3994_));
  NAND2_X1   g03802(.A1(new_n3903_), .A2(new_n193_), .ZN(new_n3995_));
  NAND3_X1   g03803(.A1(new_n3909_), .A2(\asqrt[39] ), .A3(new_n3911_), .ZN(new_n3996_));
  NOR3_X1    g03804(.A1(new_n3995_), .A2(new_n3924_), .A3(new_n3996_), .ZN(new_n3997_));
  NOR2_X1    g03805(.A1(new_n3925_), .A2(new_n3756_), .ZN(new_n3998_));
  NOR3_X1    g03806(.A1(new_n3998_), .A2(new_n3997_), .A3(new_n3753_), .ZN(new_n3999_));
  OR2_X2     g03807(.A1(new_n3994_), .A2(new_n3999_), .Z(new_n4000_));
  NOR2_X1    g03808(.A1(\a[74] ), .A2(\a[75] ), .ZN(new_n4001_));
  INV_X1     g03809(.I(new_n4001_), .ZN(new_n4002_));
  NAND3_X1   g03810(.A1(\asqrt[38] ), .A2(\a[76] ), .A3(new_n4002_), .ZN(new_n4003_));
  INV_X1     g03811(.I(\a[76] ), .ZN(new_n4004_));
  OAI21_X1   g03812(.A1(\asqrt[38] ), .A2(new_n4004_), .B(new_n4001_), .ZN(new_n4005_));
  AOI21_X1   g03813(.A1(new_n4005_), .A2(new_n4003_), .B(new_n3681_), .ZN(new_n4006_));
  NOR3_X1    g03814(.A1(new_n3678_), .A2(\asqrt[63] ), .A3(new_n3680_), .ZN(new_n4007_));
  NAND2_X1   g03815(.A1(new_n4001_), .A2(new_n4004_), .ZN(new_n4008_));
  NAND3_X1   g03816(.A1(new_n3665_), .A2(new_n3667_), .A3(new_n4008_), .ZN(new_n4009_));
  NAND2_X1   g03817(.A1(new_n4007_), .A2(new_n4009_), .ZN(new_n4010_));
  NAND3_X1   g03818(.A1(\asqrt[38] ), .A2(\a[76] ), .A3(new_n4010_), .ZN(new_n4011_));
  INV_X1     g03819(.I(\a[77] ), .ZN(new_n4012_));
  NAND3_X1   g03820(.A1(\asqrt[38] ), .A2(new_n4004_), .A3(new_n4012_), .ZN(new_n4013_));
  OAI21_X1   g03821(.A1(new_n3925_), .A2(\a[76] ), .B(\a[77] ), .ZN(new_n4014_));
  NAND3_X1   g03822(.A1(new_n4011_), .A2(new_n4014_), .A3(new_n4013_), .ZN(new_n4015_));
  NOR3_X1    g03823(.A1(new_n4015_), .A2(new_n4006_), .A3(\asqrt[40] ), .ZN(new_n4016_));
  OAI21_X1   g03824(.A1(new_n4015_), .A2(new_n4006_), .B(\asqrt[40] ), .ZN(new_n4017_));
  OAI21_X1   g03825(.A1(new_n4000_), .A2(new_n4016_), .B(new_n4017_), .ZN(new_n4018_));
  OAI21_X1   g03826(.A1(new_n4018_), .A2(\asqrt[41] ), .B(new_n3990_), .ZN(new_n4019_));
  NAND2_X1   g03827(.A1(new_n4018_), .A2(\asqrt[41] ), .ZN(new_n4020_));
  NAND3_X1   g03828(.A1(new_n4019_), .A2(new_n4020_), .A3(new_n2960_), .ZN(new_n4021_));
  AOI21_X1   g03829(.A1(new_n4019_), .A2(new_n4020_), .B(new_n2960_), .ZN(new_n4022_));
  AOI21_X1   g03830(.A1(new_n3984_), .A2(new_n4021_), .B(new_n4022_), .ZN(new_n4023_));
  AOI21_X1   g03831(.A1(new_n4023_), .A2(new_n2749_), .B(new_n3982_), .ZN(new_n4024_));
  NAND2_X1   g03832(.A1(new_n4021_), .A2(new_n3984_), .ZN(new_n4025_));
  INV_X1     g03833(.I(new_n3990_), .ZN(new_n4026_));
  NOR2_X1    g03834(.A1(new_n3994_), .A2(new_n3999_), .ZN(new_n4027_));
  NOR3_X1    g03835(.A1(new_n3925_), .A2(new_n4004_), .A3(new_n4001_), .ZN(new_n4028_));
  AOI21_X1   g03836(.A1(new_n3925_), .A2(\a[76] ), .B(new_n4002_), .ZN(new_n4029_));
  OAI21_X1   g03837(.A1(new_n4028_), .A2(new_n4029_), .B(\asqrt[39] ), .ZN(new_n4030_));
  INV_X1     g03838(.I(new_n4010_), .ZN(new_n4031_));
  NOR3_X1    g03839(.A1(new_n3925_), .A2(new_n4004_), .A3(new_n4031_), .ZN(new_n4032_));
  NOR3_X1    g03840(.A1(new_n3925_), .A2(\a[76] ), .A3(\a[77] ), .ZN(new_n4033_));
  AOI21_X1   g03841(.A1(\asqrt[38] ), .A2(new_n4004_), .B(new_n4012_), .ZN(new_n4034_));
  NOR3_X1    g03842(.A1(new_n4032_), .A2(new_n4033_), .A3(new_n4034_), .ZN(new_n4035_));
  NAND3_X1   g03843(.A1(new_n4035_), .A2(new_n4030_), .A3(new_n3427_), .ZN(new_n4036_));
  AOI21_X1   g03844(.A1(new_n4035_), .A2(new_n4030_), .B(new_n3427_), .ZN(new_n4037_));
  AOI21_X1   g03845(.A1(new_n4027_), .A2(new_n4036_), .B(new_n4037_), .ZN(new_n4038_));
  AOI21_X1   g03846(.A1(new_n4038_), .A2(new_n3195_), .B(new_n4026_), .ZN(new_n4039_));
  NAND2_X1   g03847(.A1(new_n4036_), .A2(new_n4027_), .ZN(new_n4040_));
  AOI21_X1   g03848(.A1(new_n4040_), .A2(new_n4017_), .B(new_n3195_), .ZN(new_n4041_));
  OAI21_X1   g03849(.A1(new_n4039_), .A2(new_n4041_), .B(\asqrt[42] ), .ZN(new_n4042_));
  AOI21_X1   g03850(.A1(new_n4025_), .A2(new_n4042_), .B(new_n2749_), .ZN(new_n4043_));
  NOR3_X1    g03851(.A1(new_n4024_), .A2(\asqrt[44] ), .A3(new_n4043_), .ZN(new_n4044_));
  OAI21_X1   g03852(.A1(new_n4024_), .A2(new_n4043_), .B(\asqrt[44] ), .ZN(new_n4045_));
  OAI21_X1   g03853(.A1(new_n3979_), .A2(new_n4044_), .B(new_n4045_), .ZN(new_n4046_));
  OAI21_X1   g03854(.A1(new_n4046_), .A2(\asqrt[45] ), .B(new_n3976_), .ZN(new_n4047_));
  NAND2_X1   g03855(.A1(new_n4046_), .A2(\asqrt[45] ), .ZN(new_n4048_));
  NAND3_X1   g03856(.A1(new_n4047_), .A2(new_n4048_), .A3(new_n2134_), .ZN(new_n4049_));
  AOI21_X1   g03857(.A1(new_n4047_), .A2(new_n4048_), .B(new_n2134_), .ZN(new_n4050_));
  AOI21_X1   g03858(.A1(new_n3973_), .A2(new_n4049_), .B(new_n4050_), .ZN(new_n4051_));
  AOI21_X1   g03859(.A1(new_n4051_), .A2(new_n1953_), .B(new_n3970_), .ZN(new_n4052_));
  NAND2_X1   g03860(.A1(new_n4049_), .A2(new_n3973_), .ZN(new_n4053_));
  INV_X1     g03861(.I(new_n3976_), .ZN(new_n4054_));
  INV_X1     g03862(.I(new_n3984_), .ZN(new_n4055_));
  NOR3_X1    g03863(.A1(new_n4039_), .A2(\asqrt[42] ), .A3(new_n4041_), .ZN(new_n4056_));
  OAI21_X1   g03864(.A1(new_n4055_), .A2(new_n4056_), .B(new_n4042_), .ZN(new_n4057_));
  OAI21_X1   g03865(.A1(new_n4057_), .A2(\asqrt[43] ), .B(new_n3981_), .ZN(new_n4058_));
  NAND2_X1   g03866(.A1(new_n4057_), .A2(\asqrt[43] ), .ZN(new_n4059_));
  NAND3_X1   g03867(.A1(new_n4058_), .A2(new_n4059_), .A3(new_n2531_), .ZN(new_n4060_));
  AOI21_X1   g03868(.A1(new_n4058_), .A2(new_n4059_), .B(new_n2531_), .ZN(new_n4061_));
  AOI21_X1   g03869(.A1(new_n3978_), .A2(new_n4060_), .B(new_n4061_), .ZN(new_n4062_));
  AOI21_X1   g03870(.A1(new_n4062_), .A2(new_n2332_), .B(new_n4054_), .ZN(new_n4063_));
  NAND2_X1   g03871(.A1(new_n4060_), .A2(new_n3978_), .ZN(new_n4064_));
  AOI21_X1   g03872(.A1(new_n4064_), .A2(new_n4045_), .B(new_n2332_), .ZN(new_n4065_));
  OAI21_X1   g03873(.A1(new_n4063_), .A2(new_n4065_), .B(\asqrt[46] ), .ZN(new_n4066_));
  AOI21_X1   g03874(.A1(new_n4053_), .A2(new_n4066_), .B(new_n1953_), .ZN(new_n4067_));
  NOR3_X1    g03875(.A1(new_n4052_), .A2(\asqrt[48] ), .A3(new_n4067_), .ZN(new_n4068_));
  OAI21_X1   g03876(.A1(new_n4052_), .A2(new_n4067_), .B(\asqrt[48] ), .ZN(new_n4069_));
  OAI21_X1   g03877(.A1(new_n3967_), .A2(new_n4068_), .B(new_n4069_), .ZN(new_n4070_));
  OAI21_X1   g03878(.A1(new_n4070_), .A2(\asqrt[49] ), .B(new_n3964_), .ZN(new_n4071_));
  NAND2_X1   g03879(.A1(new_n4070_), .A2(\asqrt[49] ), .ZN(new_n4072_));
  NAND3_X1   g03880(.A1(new_n4071_), .A2(new_n4072_), .A3(new_n1463_), .ZN(new_n4073_));
  AOI21_X1   g03881(.A1(new_n4071_), .A2(new_n4072_), .B(new_n1463_), .ZN(new_n4074_));
  AOI21_X1   g03882(.A1(new_n3961_), .A2(new_n4073_), .B(new_n4074_), .ZN(new_n4075_));
  AOI21_X1   g03883(.A1(new_n4075_), .A2(new_n1305_), .B(new_n3958_), .ZN(new_n4076_));
  NAND2_X1   g03884(.A1(new_n4073_), .A2(new_n3961_), .ZN(new_n4077_));
  INV_X1     g03885(.I(new_n3964_), .ZN(new_n4078_));
  INV_X1     g03886(.I(new_n3973_), .ZN(new_n4079_));
  NOR3_X1    g03887(.A1(new_n4063_), .A2(\asqrt[46] ), .A3(new_n4065_), .ZN(new_n4080_));
  OAI21_X1   g03888(.A1(new_n4079_), .A2(new_n4080_), .B(new_n4066_), .ZN(new_n4081_));
  OAI21_X1   g03889(.A1(new_n4081_), .A2(\asqrt[47] ), .B(new_n3969_), .ZN(new_n4082_));
  NAND2_X1   g03890(.A1(new_n4081_), .A2(\asqrt[47] ), .ZN(new_n4083_));
  NAND3_X1   g03891(.A1(new_n4082_), .A2(new_n4083_), .A3(new_n1778_), .ZN(new_n4084_));
  AOI21_X1   g03892(.A1(new_n4082_), .A2(new_n4083_), .B(new_n1778_), .ZN(new_n4085_));
  AOI21_X1   g03893(.A1(new_n3966_), .A2(new_n4084_), .B(new_n4085_), .ZN(new_n4086_));
  AOI21_X1   g03894(.A1(new_n4086_), .A2(new_n1632_), .B(new_n4078_), .ZN(new_n4087_));
  NAND2_X1   g03895(.A1(new_n4084_), .A2(new_n3966_), .ZN(new_n4088_));
  AOI21_X1   g03896(.A1(new_n4088_), .A2(new_n4069_), .B(new_n1632_), .ZN(new_n4089_));
  OAI21_X1   g03897(.A1(new_n4087_), .A2(new_n4089_), .B(\asqrt[50] ), .ZN(new_n4090_));
  AOI21_X1   g03898(.A1(new_n4077_), .A2(new_n4090_), .B(new_n1305_), .ZN(new_n4091_));
  NOR3_X1    g03899(.A1(new_n4076_), .A2(\asqrt[52] ), .A3(new_n4091_), .ZN(new_n4092_));
  OAI21_X1   g03900(.A1(new_n4076_), .A2(new_n4091_), .B(\asqrt[52] ), .ZN(new_n4093_));
  OAI21_X1   g03901(.A1(new_n3955_), .A2(new_n4092_), .B(new_n4093_), .ZN(new_n4094_));
  OAI21_X1   g03902(.A1(new_n4094_), .A2(\asqrt[53] ), .B(new_n3952_), .ZN(new_n4095_));
  NAND2_X1   g03903(.A1(new_n4094_), .A2(\asqrt[53] ), .ZN(new_n4096_));
  NAND3_X1   g03904(.A1(new_n4095_), .A2(new_n4096_), .A3(new_n860_), .ZN(new_n4097_));
  AOI21_X1   g03905(.A1(new_n4095_), .A2(new_n4096_), .B(new_n860_), .ZN(new_n4098_));
  AOI21_X1   g03906(.A1(new_n3949_), .A2(new_n4097_), .B(new_n4098_), .ZN(new_n4099_));
  AOI21_X1   g03907(.A1(new_n4099_), .A2(new_n744_), .B(new_n3946_), .ZN(new_n4100_));
  NAND2_X1   g03908(.A1(new_n4097_), .A2(new_n3949_), .ZN(new_n4101_));
  INV_X1     g03909(.I(new_n3952_), .ZN(new_n4102_));
  INV_X1     g03910(.I(new_n3961_), .ZN(new_n4103_));
  NOR3_X1    g03911(.A1(new_n4087_), .A2(\asqrt[50] ), .A3(new_n4089_), .ZN(new_n4104_));
  OAI21_X1   g03912(.A1(new_n4103_), .A2(new_n4104_), .B(new_n4090_), .ZN(new_n4105_));
  OAI21_X1   g03913(.A1(new_n4105_), .A2(\asqrt[51] ), .B(new_n3957_), .ZN(new_n4106_));
  NAND2_X1   g03914(.A1(new_n4105_), .A2(\asqrt[51] ), .ZN(new_n4107_));
  NAND3_X1   g03915(.A1(new_n4106_), .A2(new_n4107_), .A3(new_n1150_), .ZN(new_n4108_));
  AOI21_X1   g03916(.A1(new_n4106_), .A2(new_n4107_), .B(new_n1150_), .ZN(new_n4109_));
  AOI21_X1   g03917(.A1(new_n3954_), .A2(new_n4108_), .B(new_n4109_), .ZN(new_n4110_));
  AOI21_X1   g03918(.A1(new_n4110_), .A2(new_n1006_), .B(new_n4102_), .ZN(new_n4111_));
  NAND2_X1   g03919(.A1(new_n4108_), .A2(new_n3954_), .ZN(new_n4112_));
  AOI21_X1   g03920(.A1(new_n4112_), .A2(new_n4093_), .B(new_n1006_), .ZN(new_n4113_));
  OAI21_X1   g03921(.A1(new_n4111_), .A2(new_n4113_), .B(\asqrt[54] ), .ZN(new_n4114_));
  AOI21_X1   g03922(.A1(new_n4101_), .A2(new_n4114_), .B(new_n744_), .ZN(new_n4115_));
  NOR3_X1    g03923(.A1(new_n4100_), .A2(\asqrt[56] ), .A3(new_n4115_), .ZN(new_n4116_));
  OAI21_X1   g03924(.A1(new_n4100_), .A2(new_n4115_), .B(\asqrt[56] ), .ZN(new_n4117_));
  OAI21_X1   g03925(.A1(new_n3943_), .A2(new_n4116_), .B(new_n4117_), .ZN(new_n4118_));
  OAI21_X1   g03926(.A1(new_n4118_), .A2(\asqrt[57] ), .B(new_n3940_), .ZN(new_n4119_));
  NAND2_X1   g03927(.A1(new_n4118_), .A2(\asqrt[57] ), .ZN(new_n4120_));
  NAND3_X1   g03928(.A1(new_n4119_), .A2(new_n4120_), .A3(new_n423_), .ZN(new_n4121_));
  AOI21_X1   g03929(.A1(new_n4119_), .A2(new_n4120_), .B(new_n423_), .ZN(new_n4122_));
  AOI21_X1   g03930(.A1(new_n3937_), .A2(new_n4121_), .B(new_n4122_), .ZN(new_n4123_));
  AOI21_X1   g03931(.A1(new_n4123_), .A2(new_n337_), .B(new_n3934_), .ZN(new_n4124_));
  NAND2_X1   g03932(.A1(new_n4121_), .A2(new_n3937_), .ZN(new_n4125_));
  INV_X1     g03933(.I(new_n3940_), .ZN(new_n4126_));
  INV_X1     g03934(.I(new_n3949_), .ZN(new_n4127_));
  NOR3_X1    g03935(.A1(new_n4111_), .A2(\asqrt[54] ), .A3(new_n4113_), .ZN(new_n4128_));
  OAI21_X1   g03936(.A1(new_n4127_), .A2(new_n4128_), .B(new_n4114_), .ZN(new_n4129_));
  OAI21_X1   g03937(.A1(new_n4129_), .A2(\asqrt[55] ), .B(new_n3945_), .ZN(new_n4130_));
  NAND2_X1   g03938(.A1(new_n4129_), .A2(\asqrt[55] ), .ZN(new_n4131_));
  NAND3_X1   g03939(.A1(new_n4130_), .A2(new_n4131_), .A3(new_n634_), .ZN(new_n4132_));
  AOI21_X1   g03940(.A1(new_n4130_), .A2(new_n4131_), .B(new_n634_), .ZN(new_n4133_));
  AOI21_X1   g03941(.A1(new_n3942_), .A2(new_n4132_), .B(new_n4133_), .ZN(new_n4134_));
  AOI21_X1   g03942(.A1(new_n4134_), .A2(new_n531_), .B(new_n4126_), .ZN(new_n4135_));
  NAND2_X1   g03943(.A1(new_n4132_), .A2(new_n3942_), .ZN(new_n4136_));
  AOI21_X1   g03944(.A1(new_n4136_), .A2(new_n4117_), .B(new_n531_), .ZN(new_n4137_));
  OAI21_X1   g03945(.A1(new_n4135_), .A2(new_n4137_), .B(\asqrt[58] ), .ZN(new_n4138_));
  AOI21_X1   g03946(.A1(new_n4125_), .A2(new_n4138_), .B(new_n337_), .ZN(new_n4139_));
  NOR3_X1    g03947(.A1(new_n4124_), .A2(\asqrt[60] ), .A3(new_n4139_), .ZN(new_n4140_));
  NOR2_X1    g03948(.A1(new_n4140_), .A2(new_n3931_), .ZN(new_n4141_));
  INV_X1     g03949(.I(new_n3937_), .ZN(new_n4142_));
  NOR3_X1    g03950(.A1(new_n4135_), .A2(\asqrt[58] ), .A3(new_n4137_), .ZN(new_n4143_));
  OAI21_X1   g03951(.A1(new_n4142_), .A2(new_n4143_), .B(new_n4138_), .ZN(new_n4144_));
  OAI21_X1   g03952(.A1(new_n4144_), .A2(\asqrt[59] ), .B(new_n3933_), .ZN(new_n4145_));
  NOR2_X1    g03953(.A1(new_n4143_), .A2(new_n4142_), .ZN(new_n4146_));
  OAI21_X1   g03954(.A1(new_n4146_), .A2(new_n4122_), .B(\asqrt[59] ), .ZN(new_n4147_));
  AOI21_X1   g03955(.A1(new_n4145_), .A2(new_n4147_), .B(new_n266_), .ZN(new_n4148_));
  OAI21_X1   g03956(.A1(new_n4141_), .A2(new_n4148_), .B(\asqrt[61] ), .ZN(new_n4149_));
  OAI21_X1   g03957(.A1(new_n4124_), .A2(new_n4139_), .B(\asqrt[60] ), .ZN(new_n4150_));
  OAI21_X1   g03958(.A1(new_n3931_), .A2(new_n4140_), .B(new_n4150_), .ZN(new_n4151_));
  AOI21_X1   g03959(.A1(new_n3886_), .A2(new_n3866_), .B(\asqrt[38] ), .ZN(new_n4152_));
  XOR2_X1    g03960(.A1(new_n4152_), .A2(new_n3686_), .Z(new_n4153_));
  OAI21_X1   g03961(.A1(new_n4151_), .A2(\asqrt[61] ), .B(new_n4153_), .ZN(new_n4154_));
  NAND2_X1   g03962(.A1(new_n4154_), .A2(new_n4149_), .ZN(new_n4155_));
  NAND3_X1   g03963(.A1(new_n4145_), .A2(new_n266_), .A3(new_n4147_), .ZN(new_n4156_));
  NAND2_X1   g03964(.A1(new_n4156_), .A2(new_n3930_), .ZN(new_n4157_));
  AOI21_X1   g03965(.A1(new_n4157_), .A2(new_n4150_), .B(new_n239_), .ZN(new_n4158_));
  AOI21_X1   g03966(.A1(new_n3930_), .A2(new_n4156_), .B(new_n4148_), .ZN(new_n4159_));
  INV_X1     g03967(.I(new_n4153_), .ZN(new_n4160_));
  AOI21_X1   g03968(.A1(new_n4159_), .A2(new_n239_), .B(new_n4160_), .ZN(new_n4161_));
  OAI21_X1   g03969(.A1(new_n4161_), .A2(new_n4158_), .B(new_n201_), .ZN(new_n4162_));
  NAND3_X1   g03970(.A1(new_n4154_), .A2(\asqrt[62] ), .A3(new_n4149_), .ZN(new_n4163_));
  NAND2_X1   g03971(.A1(new_n3890_), .A2(new_n239_), .ZN(new_n4164_));
  AOI21_X1   g03972(.A1(new_n3868_), .A2(new_n4164_), .B(\asqrt[38] ), .ZN(new_n4165_));
  XOR2_X1    g03973(.A1(new_n4165_), .A2(new_n3870_), .Z(new_n4166_));
  INV_X1     g03974(.I(new_n4166_), .ZN(new_n4167_));
  AOI22_X1   g03975(.A1(new_n4162_), .A2(new_n4163_), .B1(new_n4155_), .B2(new_n4167_), .ZN(new_n4168_));
  NOR2_X1    g03976(.A1(new_n3899_), .A2(new_n3684_), .ZN(new_n4169_));
  OAI21_X1   g03977(.A1(\asqrt[38] ), .A2(new_n4169_), .B(new_n3906_), .ZN(new_n4170_));
  INV_X1     g03978(.I(new_n4170_), .ZN(new_n4171_));
  OAI21_X1   g03979(.A1(new_n4168_), .A2(new_n3928_), .B(new_n4171_), .ZN(new_n4172_));
  OAI21_X1   g03980(.A1(new_n4155_), .A2(\asqrt[62] ), .B(new_n4166_), .ZN(new_n4173_));
  NAND2_X1   g03981(.A1(new_n4155_), .A2(\asqrt[62] ), .ZN(new_n4174_));
  NAND3_X1   g03982(.A1(new_n4173_), .A2(new_n4174_), .A3(new_n3928_), .ZN(new_n4175_));
  NAND2_X1   g03983(.A1(new_n3925_), .A2(new_n3683_), .ZN(new_n4176_));
  XOR2_X1    g03984(.A1(new_n3921_), .A2(new_n3683_), .Z(new_n4177_));
  NAND3_X1   g03985(.A1(new_n4176_), .A2(\asqrt[63] ), .A3(new_n4177_), .ZN(new_n4178_));
  INV_X1     g03986(.I(new_n3995_), .ZN(new_n4179_));
  NAND4_X1   g03987(.A1(new_n4179_), .A2(new_n3684_), .A3(new_n3906_), .A4(new_n3913_), .ZN(new_n4180_));
  NAND2_X1   g03988(.A1(new_n4178_), .A2(new_n4180_), .ZN(new_n4181_));
  INV_X1     g03989(.I(new_n4181_), .ZN(new_n4182_));
  NAND4_X1   g03990(.A1(new_n4172_), .A2(new_n193_), .A3(new_n4175_), .A4(new_n4182_), .ZN(\asqrt[37] ));
  NOR2_X1    g03991(.A1(new_n4155_), .A2(\asqrt[62] ), .ZN(new_n4184_));
  INV_X1     g03992(.I(new_n4174_), .ZN(new_n4185_));
  NOR2_X1    g03993(.A1(new_n4185_), .A2(new_n4184_), .ZN(new_n4186_));
  NAND3_X1   g03994(.A1(new_n4157_), .A2(new_n239_), .A3(new_n4150_), .ZN(new_n4187_));
  AOI21_X1   g03995(.A1(new_n4153_), .A2(new_n4187_), .B(new_n4158_), .ZN(new_n4188_));
  AOI21_X1   g03996(.A1(new_n4154_), .A2(new_n4149_), .B(\asqrt[62] ), .ZN(new_n4189_));
  NOR3_X1    g03997(.A1(new_n4161_), .A2(new_n201_), .A3(new_n4158_), .ZN(new_n4190_));
  OAI22_X1   g03998(.A1(new_n4190_), .A2(new_n4189_), .B1(new_n4188_), .B2(new_n4166_), .ZN(new_n4191_));
  AOI21_X1   g03999(.A1(new_n4191_), .A2(new_n3927_), .B(new_n4170_), .ZN(new_n4192_));
  AOI21_X1   g04000(.A1(new_n4188_), .A2(new_n201_), .B(new_n4167_), .ZN(new_n4193_));
  OAI21_X1   g04001(.A1(new_n4188_), .A2(new_n201_), .B(new_n3928_), .ZN(new_n4194_));
  NOR2_X1    g04002(.A1(new_n4193_), .A2(new_n4194_), .ZN(new_n4195_));
  NOR4_X1    g04003(.A1(new_n4192_), .A2(\asqrt[63] ), .A3(new_n4195_), .A4(new_n4181_), .ZN(new_n4196_));
  XOR2_X1    g04004(.A1(new_n4165_), .A2(new_n3870_), .Z(new_n4197_));
  OAI21_X1   g04005(.A1(\asqrt[37] ), .A2(new_n4186_), .B(new_n4197_), .ZN(new_n4198_));
  INV_X1     g04006(.I(new_n4198_), .ZN(new_n4199_));
  NAND2_X1   g04007(.A1(new_n4123_), .A2(new_n337_), .ZN(new_n4200_));
  AOI21_X1   g04008(.A1(new_n4200_), .A2(new_n4147_), .B(\asqrt[37] ), .ZN(new_n4201_));
  XOR2_X1    g04009(.A1(new_n4201_), .A2(new_n3933_), .Z(new_n4202_));
  INV_X1     g04010(.I(new_n4202_), .ZN(new_n4203_));
  AOI21_X1   g04011(.A1(new_n4121_), .A2(new_n4138_), .B(\asqrt[37] ), .ZN(new_n4204_));
  XOR2_X1    g04012(.A1(new_n4204_), .A2(new_n3937_), .Z(new_n4205_));
  INV_X1     g04013(.I(new_n4205_), .ZN(new_n4206_));
  NAND2_X1   g04014(.A1(new_n4134_), .A2(new_n531_), .ZN(new_n4207_));
  AOI21_X1   g04015(.A1(new_n4207_), .A2(new_n4120_), .B(\asqrt[37] ), .ZN(new_n4208_));
  XOR2_X1    g04016(.A1(new_n4208_), .A2(new_n3940_), .Z(new_n4209_));
  INV_X1     g04017(.I(new_n4209_), .ZN(new_n4210_));
  AOI21_X1   g04018(.A1(new_n4132_), .A2(new_n4117_), .B(\asqrt[37] ), .ZN(new_n4211_));
  XOR2_X1    g04019(.A1(new_n4211_), .A2(new_n3942_), .Z(new_n4212_));
  NAND2_X1   g04020(.A1(new_n4099_), .A2(new_n744_), .ZN(new_n4213_));
  AOI21_X1   g04021(.A1(new_n4213_), .A2(new_n4131_), .B(\asqrt[37] ), .ZN(new_n4214_));
  XOR2_X1    g04022(.A1(new_n4214_), .A2(new_n3945_), .Z(new_n4215_));
  AOI21_X1   g04023(.A1(new_n4097_), .A2(new_n4114_), .B(\asqrt[37] ), .ZN(new_n4216_));
  XOR2_X1    g04024(.A1(new_n4216_), .A2(new_n3949_), .Z(new_n4217_));
  INV_X1     g04025(.I(new_n4217_), .ZN(new_n4218_));
  NAND2_X1   g04026(.A1(new_n4110_), .A2(new_n1006_), .ZN(new_n4219_));
  AOI21_X1   g04027(.A1(new_n4219_), .A2(new_n4096_), .B(\asqrt[37] ), .ZN(new_n4220_));
  XOR2_X1    g04028(.A1(new_n4220_), .A2(new_n3952_), .Z(new_n4221_));
  INV_X1     g04029(.I(new_n4221_), .ZN(new_n4222_));
  AOI21_X1   g04030(.A1(new_n4108_), .A2(new_n4093_), .B(\asqrt[37] ), .ZN(new_n4223_));
  XOR2_X1    g04031(.A1(new_n4223_), .A2(new_n3954_), .Z(new_n4224_));
  NAND2_X1   g04032(.A1(new_n4075_), .A2(new_n1305_), .ZN(new_n4225_));
  AOI21_X1   g04033(.A1(new_n4225_), .A2(new_n4107_), .B(\asqrt[37] ), .ZN(new_n4226_));
  XOR2_X1    g04034(.A1(new_n4226_), .A2(new_n3957_), .Z(new_n4227_));
  AOI21_X1   g04035(.A1(new_n4073_), .A2(new_n4090_), .B(\asqrt[37] ), .ZN(new_n4228_));
  XOR2_X1    g04036(.A1(new_n4228_), .A2(new_n3961_), .Z(new_n4229_));
  INV_X1     g04037(.I(new_n4229_), .ZN(new_n4230_));
  NAND2_X1   g04038(.A1(new_n4086_), .A2(new_n1632_), .ZN(new_n4231_));
  AOI21_X1   g04039(.A1(new_n4231_), .A2(new_n4072_), .B(\asqrt[37] ), .ZN(new_n4232_));
  XOR2_X1    g04040(.A1(new_n4232_), .A2(new_n3964_), .Z(new_n4233_));
  INV_X1     g04041(.I(new_n4233_), .ZN(new_n4234_));
  AOI21_X1   g04042(.A1(new_n4084_), .A2(new_n4069_), .B(\asqrt[37] ), .ZN(new_n4235_));
  XOR2_X1    g04043(.A1(new_n4235_), .A2(new_n3966_), .Z(new_n4236_));
  NAND2_X1   g04044(.A1(new_n4051_), .A2(new_n1953_), .ZN(new_n4237_));
  AOI21_X1   g04045(.A1(new_n4237_), .A2(new_n4083_), .B(\asqrt[37] ), .ZN(new_n4238_));
  XOR2_X1    g04046(.A1(new_n4238_), .A2(new_n3969_), .Z(new_n4239_));
  AOI21_X1   g04047(.A1(new_n4049_), .A2(new_n4066_), .B(\asqrt[37] ), .ZN(new_n4240_));
  XOR2_X1    g04048(.A1(new_n4240_), .A2(new_n3973_), .Z(new_n4241_));
  INV_X1     g04049(.I(new_n4241_), .ZN(new_n4242_));
  NAND2_X1   g04050(.A1(new_n4062_), .A2(new_n2332_), .ZN(new_n4243_));
  AOI21_X1   g04051(.A1(new_n4243_), .A2(new_n4048_), .B(\asqrt[37] ), .ZN(new_n4244_));
  XOR2_X1    g04052(.A1(new_n4244_), .A2(new_n3976_), .Z(new_n4245_));
  INV_X1     g04053(.I(new_n4245_), .ZN(new_n4246_));
  AOI21_X1   g04054(.A1(new_n4060_), .A2(new_n4045_), .B(\asqrt[37] ), .ZN(new_n4247_));
  XOR2_X1    g04055(.A1(new_n4247_), .A2(new_n3978_), .Z(new_n4248_));
  NAND2_X1   g04056(.A1(new_n4023_), .A2(new_n2749_), .ZN(new_n4249_));
  AOI21_X1   g04057(.A1(new_n4249_), .A2(new_n4059_), .B(\asqrt[37] ), .ZN(new_n4250_));
  XOR2_X1    g04058(.A1(new_n4250_), .A2(new_n3981_), .Z(new_n4251_));
  AOI21_X1   g04059(.A1(new_n4021_), .A2(new_n4042_), .B(\asqrt[37] ), .ZN(new_n4252_));
  XOR2_X1    g04060(.A1(new_n4252_), .A2(new_n3984_), .Z(new_n4253_));
  INV_X1     g04061(.I(new_n4253_), .ZN(new_n4254_));
  NAND2_X1   g04062(.A1(new_n4038_), .A2(new_n3195_), .ZN(new_n4255_));
  AOI21_X1   g04063(.A1(new_n4255_), .A2(new_n4020_), .B(\asqrt[37] ), .ZN(new_n4256_));
  XOR2_X1    g04064(.A1(new_n4256_), .A2(new_n3990_), .Z(new_n4257_));
  INV_X1     g04065(.I(new_n4257_), .ZN(new_n4258_));
  AOI21_X1   g04066(.A1(new_n4036_), .A2(new_n4017_), .B(\asqrt[37] ), .ZN(new_n4259_));
  XOR2_X1    g04067(.A1(new_n4259_), .A2(new_n4027_), .Z(new_n4260_));
  NAND2_X1   g04068(.A1(\asqrt[38] ), .A2(new_n4004_), .ZN(new_n4261_));
  NOR2_X1    g04069(.A1(new_n4012_), .A2(\a[76] ), .ZN(new_n4262_));
  AOI22_X1   g04070(.A1(new_n4261_), .A2(new_n4012_), .B1(\asqrt[38] ), .B2(new_n4262_), .ZN(new_n4263_));
  AOI21_X1   g04071(.A1(\asqrt[38] ), .A2(\a[76] ), .B(new_n4010_), .ZN(new_n4264_));
  OAI21_X1   g04072(.A1(new_n4006_), .A2(new_n4264_), .B(new_n4196_), .ZN(new_n4265_));
  XNOR2_X1   g04073(.A1(new_n4265_), .A2(new_n4263_), .ZN(new_n4266_));
  NOR3_X1    g04074(.A1(new_n4192_), .A2(\asqrt[63] ), .A3(new_n4195_), .ZN(new_n4267_));
  NAND3_X1   g04075(.A1(new_n4178_), .A2(\asqrt[38] ), .A3(new_n4180_), .ZN(new_n4268_));
  INV_X1     g04076(.I(new_n4268_), .ZN(new_n4269_));
  NAND2_X1   g04077(.A1(new_n4267_), .A2(new_n4269_), .ZN(new_n4270_));
  NAND2_X1   g04078(.A1(\asqrt[37] ), .A2(new_n4001_), .ZN(new_n4271_));
  AOI21_X1   g04079(.A1(new_n4271_), .A2(new_n4270_), .B(\a[76] ), .ZN(new_n4272_));
  NAND2_X1   g04080(.A1(new_n4172_), .A2(new_n193_), .ZN(new_n4273_));
  NOR3_X1    g04081(.A1(new_n4273_), .A2(new_n4195_), .A3(new_n4268_), .ZN(new_n4274_));
  NOR2_X1    g04082(.A1(new_n4196_), .A2(new_n4002_), .ZN(new_n4275_));
  NOR3_X1    g04083(.A1(new_n4275_), .A2(new_n4274_), .A3(new_n4004_), .ZN(new_n4276_));
  OR2_X2     g04084(.A1(new_n4276_), .A2(new_n4272_), .Z(new_n4277_));
  NOR2_X1    g04085(.A1(\a[72] ), .A2(\a[73] ), .ZN(new_n4278_));
  INV_X1     g04086(.I(new_n4278_), .ZN(new_n4279_));
  NAND3_X1   g04087(.A1(\asqrt[37] ), .A2(\a[74] ), .A3(new_n4279_), .ZN(new_n4280_));
  INV_X1     g04088(.I(\a[74] ), .ZN(new_n4281_));
  OAI21_X1   g04089(.A1(\asqrt[37] ), .A2(new_n4281_), .B(new_n4278_), .ZN(new_n4282_));
  AOI21_X1   g04090(.A1(new_n4282_), .A2(new_n4280_), .B(new_n3925_), .ZN(new_n4283_));
  NAND2_X1   g04091(.A1(new_n4278_), .A2(new_n4281_), .ZN(new_n4284_));
  NAND3_X1   g04092(.A1(new_n3909_), .A2(new_n3911_), .A3(new_n4284_), .ZN(new_n4285_));
  NAND2_X1   g04093(.A1(new_n3991_), .A2(new_n4285_), .ZN(new_n4286_));
  NAND3_X1   g04094(.A1(\asqrt[37] ), .A2(\a[74] ), .A3(new_n4286_), .ZN(new_n4287_));
  INV_X1     g04095(.I(\a[75] ), .ZN(new_n4288_));
  NAND3_X1   g04096(.A1(\asqrt[37] ), .A2(new_n4281_), .A3(new_n4288_), .ZN(new_n4289_));
  OAI21_X1   g04097(.A1(new_n4196_), .A2(\a[74] ), .B(\a[75] ), .ZN(new_n4290_));
  NAND3_X1   g04098(.A1(new_n4287_), .A2(new_n4290_), .A3(new_n4289_), .ZN(new_n4291_));
  NOR3_X1    g04099(.A1(new_n4291_), .A2(new_n4283_), .A3(\asqrt[39] ), .ZN(new_n4292_));
  OAI21_X1   g04100(.A1(new_n4291_), .A2(new_n4283_), .B(\asqrt[39] ), .ZN(new_n4293_));
  OAI21_X1   g04101(.A1(new_n4277_), .A2(new_n4292_), .B(new_n4293_), .ZN(new_n4294_));
  OAI21_X1   g04102(.A1(new_n4294_), .A2(\asqrt[40] ), .B(new_n4266_), .ZN(new_n4295_));
  NAND2_X1   g04103(.A1(new_n4294_), .A2(\asqrt[40] ), .ZN(new_n4296_));
  NAND3_X1   g04104(.A1(new_n4295_), .A2(new_n4296_), .A3(new_n3195_), .ZN(new_n4297_));
  AOI21_X1   g04105(.A1(new_n4295_), .A2(new_n4296_), .B(new_n3195_), .ZN(new_n4298_));
  AOI21_X1   g04106(.A1(new_n4260_), .A2(new_n4297_), .B(new_n4298_), .ZN(new_n4299_));
  AOI21_X1   g04107(.A1(new_n4299_), .A2(new_n2960_), .B(new_n4258_), .ZN(new_n4300_));
  NAND2_X1   g04108(.A1(new_n4297_), .A2(new_n4260_), .ZN(new_n4301_));
  INV_X1     g04109(.I(new_n4298_), .ZN(new_n4302_));
  AOI21_X1   g04110(.A1(new_n4301_), .A2(new_n4302_), .B(new_n2960_), .ZN(new_n4303_));
  NOR3_X1    g04111(.A1(new_n4300_), .A2(\asqrt[43] ), .A3(new_n4303_), .ZN(new_n4304_));
  OAI21_X1   g04112(.A1(new_n4300_), .A2(new_n4303_), .B(\asqrt[43] ), .ZN(new_n4305_));
  OAI21_X1   g04113(.A1(new_n4254_), .A2(new_n4304_), .B(new_n4305_), .ZN(new_n4306_));
  OAI21_X1   g04114(.A1(new_n4306_), .A2(\asqrt[44] ), .B(new_n4251_), .ZN(new_n4307_));
  NAND2_X1   g04115(.A1(new_n4306_), .A2(\asqrt[44] ), .ZN(new_n4308_));
  NAND3_X1   g04116(.A1(new_n4307_), .A2(new_n4308_), .A3(new_n2332_), .ZN(new_n4309_));
  AOI21_X1   g04117(.A1(new_n4307_), .A2(new_n4308_), .B(new_n2332_), .ZN(new_n4310_));
  AOI21_X1   g04118(.A1(new_n4248_), .A2(new_n4309_), .B(new_n4310_), .ZN(new_n4311_));
  AOI21_X1   g04119(.A1(new_n4311_), .A2(new_n2134_), .B(new_n4246_), .ZN(new_n4312_));
  NAND2_X1   g04120(.A1(new_n4309_), .A2(new_n4248_), .ZN(new_n4313_));
  INV_X1     g04121(.I(new_n4310_), .ZN(new_n4314_));
  AOI21_X1   g04122(.A1(new_n4313_), .A2(new_n4314_), .B(new_n2134_), .ZN(new_n4315_));
  NOR3_X1    g04123(.A1(new_n4312_), .A2(\asqrt[47] ), .A3(new_n4315_), .ZN(new_n4316_));
  OAI21_X1   g04124(.A1(new_n4312_), .A2(new_n4315_), .B(\asqrt[47] ), .ZN(new_n4317_));
  OAI21_X1   g04125(.A1(new_n4242_), .A2(new_n4316_), .B(new_n4317_), .ZN(new_n4318_));
  OAI21_X1   g04126(.A1(new_n4318_), .A2(\asqrt[48] ), .B(new_n4239_), .ZN(new_n4319_));
  NAND2_X1   g04127(.A1(new_n4318_), .A2(\asqrt[48] ), .ZN(new_n4320_));
  NAND3_X1   g04128(.A1(new_n4319_), .A2(new_n4320_), .A3(new_n1632_), .ZN(new_n4321_));
  AOI21_X1   g04129(.A1(new_n4319_), .A2(new_n4320_), .B(new_n1632_), .ZN(new_n4322_));
  AOI21_X1   g04130(.A1(new_n4236_), .A2(new_n4321_), .B(new_n4322_), .ZN(new_n4323_));
  AOI21_X1   g04131(.A1(new_n4323_), .A2(new_n1463_), .B(new_n4234_), .ZN(new_n4324_));
  NAND2_X1   g04132(.A1(new_n4321_), .A2(new_n4236_), .ZN(new_n4325_));
  INV_X1     g04133(.I(new_n4322_), .ZN(new_n4326_));
  AOI21_X1   g04134(.A1(new_n4325_), .A2(new_n4326_), .B(new_n1463_), .ZN(new_n4327_));
  NOR3_X1    g04135(.A1(new_n4324_), .A2(\asqrt[51] ), .A3(new_n4327_), .ZN(new_n4328_));
  OAI21_X1   g04136(.A1(new_n4324_), .A2(new_n4327_), .B(\asqrt[51] ), .ZN(new_n4329_));
  OAI21_X1   g04137(.A1(new_n4230_), .A2(new_n4328_), .B(new_n4329_), .ZN(new_n4330_));
  OAI21_X1   g04138(.A1(new_n4330_), .A2(\asqrt[52] ), .B(new_n4227_), .ZN(new_n4331_));
  NAND2_X1   g04139(.A1(new_n4330_), .A2(\asqrt[52] ), .ZN(new_n4332_));
  NAND3_X1   g04140(.A1(new_n4331_), .A2(new_n4332_), .A3(new_n1006_), .ZN(new_n4333_));
  AOI21_X1   g04141(.A1(new_n4331_), .A2(new_n4332_), .B(new_n1006_), .ZN(new_n4334_));
  AOI21_X1   g04142(.A1(new_n4224_), .A2(new_n4333_), .B(new_n4334_), .ZN(new_n4335_));
  AOI21_X1   g04143(.A1(new_n4335_), .A2(new_n860_), .B(new_n4222_), .ZN(new_n4336_));
  NAND2_X1   g04144(.A1(new_n4333_), .A2(new_n4224_), .ZN(new_n4337_));
  INV_X1     g04145(.I(new_n4334_), .ZN(new_n4338_));
  AOI21_X1   g04146(.A1(new_n4337_), .A2(new_n4338_), .B(new_n860_), .ZN(new_n4339_));
  NOR3_X1    g04147(.A1(new_n4336_), .A2(\asqrt[55] ), .A3(new_n4339_), .ZN(new_n4340_));
  OAI21_X1   g04148(.A1(new_n4336_), .A2(new_n4339_), .B(\asqrt[55] ), .ZN(new_n4341_));
  OAI21_X1   g04149(.A1(new_n4218_), .A2(new_n4340_), .B(new_n4341_), .ZN(new_n4342_));
  OAI21_X1   g04150(.A1(new_n4342_), .A2(\asqrt[56] ), .B(new_n4215_), .ZN(new_n4343_));
  NAND2_X1   g04151(.A1(new_n4342_), .A2(\asqrt[56] ), .ZN(new_n4344_));
  NAND3_X1   g04152(.A1(new_n4343_), .A2(new_n4344_), .A3(new_n531_), .ZN(new_n4345_));
  AOI21_X1   g04153(.A1(new_n4343_), .A2(new_n4344_), .B(new_n531_), .ZN(new_n4346_));
  AOI21_X1   g04154(.A1(new_n4212_), .A2(new_n4345_), .B(new_n4346_), .ZN(new_n4347_));
  AOI21_X1   g04155(.A1(new_n4347_), .A2(new_n423_), .B(new_n4210_), .ZN(new_n4348_));
  NAND2_X1   g04156(.A1(new_n4345_), .A2(new_n4212_), .ZN(new_n4349_));
  INV_X1     g04157(.I(new_n4346_), .ZN(new_n4350_));
  AOI21_X1   g04158(.A1(new_n4349_), .A2(new_n4350_), .B(new_n423_), .ZN(new_n4351_));
  NOR3_X1    g04159(.A1(new_n4348_), .A2(\asqrt[59] ), .A3(new_n4351_), .ZN(new_n4352_));
  NOR2_X1    g04160(.A1(new_n4352_), .A2(new_n4206_), .ZN(new_n4353_));
  OAI21_X1   g04161(.A1(new_n4348_), .A2(new_n4351_), .B(\asqrt[59] ), .ZN(new_n4354_));
  INV_X1     g04162(.I(new_n4354_), .ZN(new_n4355_));
  NOR2_X1    g04163(.A1(new_n4353_), .A2(new_n4355_), .ZN(new_n4356_));
  AOI21_X1   g04164(.A1(new_n4356_), .A2(new_n266_), .B(new_n4203_), .ZN(new_n4357_));
  INV_X1     g04165(.I(new_n4212_), .ZN(new_n4358_));
  INV_X1     g04166(.I(new_n4224_), .ZN(new_n4359_));
  INV_X1     g04167(.I(new_n4236_), .ZN(new_n4360_));
  INV_X1     g04168(.I(new_n4248_), .ZN(new_n4361_));
  INV_X1     g04169(.I(new_n4260_), .ZN(new_n4362_));
  NOR2_X1    g04170(.A1(new_n4276_), .A2(new_n4272_), .ZN(new_n4363_));
  NOR3_X1    g04171(.A1(new_n4196_), .A2(new_n4281_), .A3(new_n4278_), .ZN(new_n4364_));
  AOI21_X1   g04172(.A1(new_n4196_), .A2(\a[74] ), .B(new_n4279_), .ZN(new_n4365_));
  OAI21_X1   g04173(.A1(new_n4364_), .A2(new_n4365_), .B(\asqrt[38] ), .ZN(new_n4366_));
  INV_X1     g04174(.I(new_n4286_), .ZN(new_n4367_));
  NOR3_X1    g04175(.A1(new_n4196_), .A2(new_n4281_), .A3(new_n4367_), .ZN(new_n4368_));
  NOR3_X1    g04176(.A1(new_n4196_), .A2(\a[74] ), .A3(\a[75] ), .ZN(new_n4369_));
  AOI21_X1   g04177(.A1(\asqrt[37] ), .A2(new_n4281_), .B(new_n4288_), .ZN(new_n4370_));
  NOR3_X1    g04178(.A1(new_n4368_), .A2(new_n4369_), .A3(new_n4370_), .ZN(new_n4371_));
  NAND3_X1   g04179(.A1(new_n4371_), .A2(new_n4366_), .A3(new_n3681_), .ZN(new_n4372_));
  NAND2_X1   g04180(.A1(new_n4372_), .A2(new_n4363_), .ZN(new_n4373_));
  NAND3_X1   g04181(.A1(new_n4373_), .A2(new_n3427_), .A3(new_n4293_), .ZN(new_n4374_));
  AOI21_X1   g04182(.A1(new_n4373_), .A2(new_n4293_), .B(new_n3427_), .ZN(new_n4375_));
  AOI21_X1   g04183(.A1(new_n4266_), .A2(new_n4374_), .B(new_n4375_), .ZN(new_n4376_));
  AOI21_X1   g04184(.A1(new_n4376_), .A2(new_n3195_), .B(new_n4362_), .ZN(new_n4377_));
  NOR3_X1    g04185(.A1(new_n4377_), .A2(\asqrt[42] ), .A3(new_n4298_), .ZN(new_n4378_));
  OAI21_X1   g04186(.A1(new_n4377_), .A2(new_n4298_), .B(\asqrt[42] ), .ZN(new_n4379_));
  OAI21_X1   g04187(.A1(new_n4258_), .A2(new_n4378_), .B(new_n4379_), .ZN(new_n4380_));
  OAI21_X1   g04188(.A1(new_n4380_), .A2(\asqrt[43] ), .B(new_n4253_), .ZN(new_n4381_));
  NAND3_X1   g04189(.A1(new_n4381_), .A2(new_n2531_), .A3(new_n4305_), .ZN(new_n4382_));
  AOI21_X1   g04190(.A1(new_n4381_), .A2(new_n4305_), .B(new_n2531_), .ZN(new_n4383_));
  AOI21_X1   g04191(.A1(new_n4251_), .A2(new_n4382_), .B(new_n4383_), .ZN(new_n4384_));
  AOI21_X1   g04192(.A1(new_n4384_), .A2(new_n2332_), .B(new_n4361_), .ZN(new_n4385_));
  NOR3_X1    g04193(.A1(new_n4385_), .A2(\asqrt[46] ), .A3(new_n4310_), .ZN(new_n4386_));
  OAI21_X1   g04194(.A1(new_n4385_), .A2(new_n4310_), .B(\asqrt[46] ), .ZN(new_n4387_));
  OAI21_X1   g04195(.A1(new_n4246_), .A2(new_n4386_), .B(new_n4387_), .ZN(new_n4388_));
  OAI21_X1   g04196(.A1(new_n4388_), .A2(\asqrt[47] ), .B(new_n4241_), .ZN(new_n4389_));
  NAND3_X1   g04197(.A1(new_n4389_), .A2(new_n1778_), .A3(new_n4317_), .ZN(new_n4390_));
  AOI21_X1   g04198(.A1(new_n4389_), .A2(new_n4317_), .B(new_n1778_), .ZN(new_n4391_));
  AOI21_X1   g04199(.A1(new_n4239_), .A2(new_n4390_), .B(new_n4391_), .ZN(new_n4392_));
  AOI21_X1   g04200(.A1(new_n4392_), .A2(new_n1632_), .B(new_n4360_), .ZN(new_n4393_));
  NOR3_X1    g04201(.A1(new_n4393_), .A2(\asqrt[50] ), .A3(new_n4322_), .ZN(new_n4394_));
  OAI21_X1   g04202(.A1(new_n4393_), .A2(new_n4322_), .B(\asqrt[50] ), .ZN(new_n4395_));
  OAI21_X1   g04203(.A1(new_n4234_), .A2(new_n4394_), .B(new_n4395_), .ZN(new_n4396_));
  OAI21_X1   g04204(.A1(new_n4396_), .A2(\asqrt[51] ), .B(new_n4229_), .ZN(new_n4397_));
  NAND3_X1   g04205(.A1(new_n4397_), .A2(new_n1150_), .A3(new_n4329_), .ZN(new_n4398_));
  AOI21_X1   g04206(.A1(new_n4397_), .A2(new_n4329_), .B(new_n1150_), .ZN(new_n4399_));
  AOI21_X1   g04207(.A1(new_n4227_), .A2(new_n4398_), .B(new_n4399_), .ZN(new_n4400_));
  AOI21_X1   g04208(.A1(new_n4400_), .A2(new_n1006_), .B(new_n4359_), .ZN(new_n4401_));
  NOR3_X1    g04209(.A1(new_n4401_), .A2(\asqrt[54] ), .A3(new_n4334_), .ZN(new_n4402_));
  OAI21_X1   g04210(.A1(new_n4401_), .A2(new_n4334_), .B(\asqrt[54] ), .ZN(new_n4403_));
  OAI21_X1   g04211(.A1(new_n4222_), .A2(new_n4402_), .B(new_n4403_), .ZN(new_n4404_));
  OAI21_X1   g04212(.A1(new_n4404_), .A2(\asqrt[55] ), .B(new_n4217_), .ZN(new_n4405_));
  NAND3_X1   g04213(.A1(new_n4405_), .A2(new_n634_), .A3(new_n4341_), .ZN(new_n4406_));
  AOI21_X1   g04214(.A1(new_n4405_), .A2(new_n4341_), .B(new_n634_), .ZN(new_n4407_));
  AOI21_X1   g04215(.A1(new_n4215_), .A2(new_n4406_), .B(new_n4407_), .ZN(new_n4408_));
  AOI21_X1   g04216(.A1(new_n4408_), .A2(new_n531_), .B(new_n4358_), .ZN(new_n4409_));
  NOR3_X1    g04217(.A1(new_n4409_), .A2(\asqrt[58] ), .A3(new_n4346_), .ZN(new_n4410_));
  OAI21_X1   g04218(.A1(new_n4409_), .A2(new_n4346_), .B(\asqrt[58] ), .ZN(new_n4411_));
  OAI21_X1   g04219(.A1(new_n4210_), .A2(new_n4410_), .B(new_n4411_), .ZN(new_n4412_));
  OAI21_X1   g04220(.A1(new_n4412_), .A2(\asqrt[59] ), .B(new_n4205_), .ZN(new_n4413_));
  AOI21_X1   g04221(.A1(new_n4413_), .A2(new_n4354_), .B(new_n266_), .ZN(new_n4414_));
  OAI21_X1   g04222(.A1(new_n4357_), .A2(new_n4414_), .B(\asqrt[61] ), .ZN(new_n4415_));
  AOI21_X1   g04223(.A1(new_n4156_), .A2(new_n4150_), .B(\asqrt[37] ), .ZN(new_n4416_));
  XOR2_X1    g04224(.A1(new_n4416_), .A2(new_n3930_), .Z(new_n4417_));
  OAI21_X1   g04225(.A1(new_n4206_), .A2(new_n4352_), .B(new_n4354_), .ZN(new_n4418_));
  OAI21_X1   g04226(.A1(new_n4418_), .A2(\asqrt[60] ), .B(new_n4202_), .ZN(new_n4419_));
  OAI21_X1   g04227(.A1(new_n4353_), .A2(new_n4355_), .B(\asqrt[60] ), .ZN(new_n4420_));
  NAND3_X1   g04228(.A1(new_n4419_), .A2(new_n239_), .A3(new_n4420_), .ZN(new_n4421_));
  NAND2_X1   g04229(.A1(new_n4421_), .A2(new_n4417_), .ZN(new_n4422_));
  NAND2_X1   g04230(.A1(new_n4422_), .A2(new_n4415_), .ZN(new_n4423_));
  AOI21_X1   g04231(.A1(new_n4419_), .A2(new_n4420_), .B(new_n239_), .ZN(new_n4424_));
  NAND3_X1   g04232(.A1(new_n4413_), .A2(new_n266_), .A3(new_n4354_), .ZN(new_n4425_));
  AOI21_X1   g04233(.A1(new_n4202_), .A2(new_n4425_), .B(new_n4414_), .ZN(new_n4426_));
  INV_X1     g04234(.I(new_n4417_), .ZN(new_n4427_));
  AOI21_X1   g04235(.A1(new_n4426_), .A2(new_n239_), .B(new_n4427_), .ZN(new_n4428_));
  OAI21_X1   g04236(.A1(new_n4428_), .A2(new_n4424_), .B(new_n201_), .ZN(new_n4429_));
  NAND3_X1   g04237(.A1(new_n4422_), .A2(\asqrt[62] ), .A3(new_n4415_), .ZN(new_n4430_));
  AOI21_X1   g04238(.A1(new_n4149_), .A2(new_n4187_), .B(\asqrt[37] ), .ZN(new_n4431_));
  XOR2_X1    g04239(.A1(new_n4431_), .A2(new_n4153_), .Z(new_n4432_));
  INV_X1     g04240(.I(new_n4432_), .ZN(new_n4433_));
  AOI22_X1   g04241(.A1(new_n4429_), .A2(new_n4430_), .B1(new_n4423_), .B2(new_n4433_), .ZN(new_n4434_));
  NOR2_X1    g04242(.A1(new_n4168_), .A2(new_n3928_), .ZN(new_n4435_));
  OAI21_X1   g04243(.A1(\asqrt[37] ), .A2(new_n4435_), .B(new_n4175_), .ZN(new_n4436_));
  INV_X1     g04244(.I(new_n4436_), .ZN(new_n4437_));
  OAI21_X1   g04245(.A1(new_n4434_), .A2(new_n4199_), .B(new_n4437_), .ZN(new_n4438_));
  OAI21_X1   g04246(.A1(new_n4423_), .A2(\asqrt[62] ), .B(new_n4432_), .ZN(new_n4439_));
  NAND2_X1   g04247(.A1(new_n4423_), .A2(\asqrt[62] ), .ZN(new_n4440_));
  NAND3_X1   g04248(.A1(new_n4439_), .A2(new_n4440_), .A3(new_n4199_), .ZN(new_n4441_));
  NAND2_X1   g04249(.A1(new_n4196_), .A2(new_n3927_), .ZN(new_n4442_));
  XOR2_X1    g04250(.A1(new_n4168_), .A2(new_n3928_), .Z(new_n4443_));
  NAND3_X1   g04251(.A1(new_n4442_), .A2(\asqrt[63] ), .A3(new_n4443_), .ZN(new_n4444_));
  INV_X1     g04252(.I(new_n4273_), .ZN(new_n4445_));
  NAND4_X1   g04253(.A1(new_n4445_), .A2(new_n3928_), .A3(new_n4175_), .A4(new_n4182_), .ZN(new_n4446_));
  NAND2_X1   g04254(.A1(new_n4444_), .A2(new_n4446_), .ZN(new_n4447_));
  INV_X1     g04255(.I(new_n4447_), .ZN(new_n4448_));
  NAND4_X1   g04256(.A1(new_n4438_), .A2(new_n193_), .A3(new_n4441_), .A4(new_n4448_), .ZN(\asqrt[36] ));
  NOR2_X1    g04257(.A1(new_n4423_), .A2(\asqrt[62] ), .ZN(new_n4450_));
  INV_X1     g04258(.I(new_n4440_), .ZN(new_n4451_));
  NOR2_X1    g04259(.A1(new_n4451_), .A2(new_n4450_), .ZN(new_n4452_));
  NOR2_X1    g04260(.A1(new_n4428_), .A2(new_n4424_), .ZN(new_n4453_));
  AOI21_X1   g04261(.A1(new_n4422_), .A2(new_n4415_), .B(\asqrt[62] ), .ZN(new_n4454_));
  NOR3_X1    g04262(.A1(new_n4428_), .A2(new_n201_), .A3(new_n4424_), .ZN(new_n4455_));
  OAI22_X1   g04263(.A1(new_n4455_), .A2(new_n4454_), .B1(new_n4453_), .B2(new_n4432_), .ZN(new_n4456_));
  AOI21_X1   g04264(.A1(new_n4456_), .A2(new_n4198_), .B(new_n4436_), .ZN(new_n4457_));
  AOI21_X1   g04265(.A1(new_n4453_), .A2(new_n201_), .B(new_n4433_), .ZN(new_n4458_));
  OAI21_X1   g04266(.A1(new_n4453_), .A2(new_n201_), .B(new_n4199_), .ZN(new_n4459_));
  NOR2_X1    g04267(.A1(new_n4458_), .A2(new_n4459_), .ZN(new_n4460_));
  NOR4_X1    g04268(.A1(new_n4457_), .A2(\asqrt[63] ), .A3(new_n4460_), .A4(new_n4447_), .ZN(new_n4461_));
  XOR2_X1    g04269(.A1(new_n4431_), .A2(new_n4153_), .Z(new_n4462_));
  OAI21_X1   g04270(.A1(\asqrt[36] ), .A2(new_n4452_), .B(new_n4462_), .ZN(new_n4463_));
  INV_X1     g04271(.I(new_n4463_), .ZN(new_n4464_));
  NOR2_X1    g04272(.A1(new_n4355_), .A2(new_n4352_), .ZN(new_n4465_));
  NOR2_X1    g04273(.A1(\asqrt[36] ), .A2(new_n4465_), .ZN(new_n4466_));
  XOR2_X1    g04274(.A1(new_n4466_), .A2(new_n4205_), .Z(new_n4467_));
  INV_X1     g04275(.I(new_n4467_), .ZN(new_n4468_));
  NOR2_X1    g04276(.A1(new_n4410_), .A2(new_n4351_), .ZN(new_n4469_));
  NOR2_X1    g04277(.A1(\asqrt[36] ), .A2(new_n4469_), .ZN(new_n4470_));
  XOR2_X1    g04278(.A1(new_n4470_), .A2(new_n4209_), .Z(new_n4471_));
  AOI21_X1   g04279(.A1(new_n4345_), .A2(new_n4350_), .B(\asqrt[36] ), .ZN(new_n4472_));
  XOR2_X1    g04280(.A1(new_n4472_), .A2(new_n4212_), .Z(new_n4473_));
  AOI21_X1   g04281(.A1(new_n4406_), .A2(new_n4344_), .B(\asqrt[36] ), .ZN(new_n4474_));
  XOR2_X1    g04282(.A1(new_n4474_), .A2(new_n4215_), .Z(new_n4475_));
  INV_X1     g04283(.I(new_n4341_), .ZN(new_n4476_));
  NOR2_X1    g04284(.A1(new_n4476_), .A2(new_n4340_), .ZN(new_n4477_));
  NOR2_X1    g04285(.A1(\asqrt[36] ), .A2(new_n4477_), .ZN(new_n4478_));
  XOR2_X1    g04286(.A1(new_n4478_), .A2(new_n4217_), .Z(new_n4479_));
  INV_X1     g04287(.I(new_n4479_), .ZN(new_n4480_));
  NOR2_X1    g04288(.A1(new_n4402_), .A2(new_n4339_), .ZN(new_n4481_));
  NOR2_X1    g04289(.A1(\asqrt[36] ), .A2(new_n4481_), .ZN(new_n4482_));
  XOR2_X1    g04290(.A1(new_n4482_), .A2(new_n4221_), .Z(new_n4483_));
  INV_X1     g04291(.I(new_n4483_), .ZN(new_n4484_));
  AOI21_X1   g04292(.A1(new_n4333_), .A2(new_n4338_), .B(\asqrt[36] ), .ZN(new_n4485_));
  XOR2_X1    g04293(.A1(new_n4485_), .A2(new_n4224_), .Z(new_n4486_));
  AOI21_X1   g04294(.A1(new_n4398_), .A2(new_n4332_), .B(\asqrt[36] ), .ZN(new_n4487_));
  XOR2_X1    g04295(.A1(new_n4487_), .A2(new_n4227_), .Z(new_n4488_));
  XOR2_X1    g04296(.A1(new_n4396_), .A2(\asqrt[51] ), .Z(new_n4489_));
  NOR2_X1    g04297(.A1(\asqrt[36] ), .A2(new_n4489_), .ZN(new_n4490_));
  XOR2_X1    g04298(.A1(new_n4490_), .A2(new_n4229_), .Z(new_n4491_));
  INV_X1     g04299(.I(new_n4491_), .ZN(new_n4492_));
  NOR2_X1    g04300(.A1(new_n4394_), .A2(new_n4327_), .ZN(new_n4493_));
  NOR2_X1    g04301(.A1(\asqrt[36] ), .A2(new_n4493_), .ZN(new_n4494_));
  XOR2_X1    g04302(.A1(new_n4494_), .A2(new_n4233_), .Z(new_n4495_));
  INV_X1     g04303(.I(new_n4495_), .ZN(new_n4496_));
  AOI21_X1   g04304(.A1(new_n4321_), .A2(new_n4326_), .B(\asqrt[36] ), .ZN(new_n4497_));
  XOR2_X1    g04305(.A1(new_n4497_), .A2(new_n4236_), .Z(new_n4498_));
  AOI21_X1   g04306(.A1(new_n4390_), .A2(new_n4320_), .B(\asqrt[36] ), .ZN(new_n4499_));
  XOR2_X1    g04307(.A1(new_n4499_), .A2(new_n4239_), .Z(new_n4500_));
  XOR2_X1    g04308(.A1(new_n4388_), .A2(\asqrt[47] ), .Z(new_n4501_));
  NOR2_X1    g04309(.A1(\asqrt[36] ), .A2(new_n4501_), .ZN(new_n4502_));
  XOR2_X1    g04310(.A1(new_n4502_), .A2(new_n4241_), .Z(new_n4503_));
  INV_X1     g04311(.I(new_n4503_), .ZN(new_n4504_));
  NOR2_X1    g04312(.A1(new_n4386_), .A2(new_n4315_), .ZN(new_n4505_));
  NOR2_X1    g04313(.A1(\asqrt[36] ), .A2(new_n4505_), .ZN(new_n4506_));
  XOR2_X1    g04314(.A1(new_n4506_), .A2(new_n4245_), .Z(new_n4507_));
  INV_X1     g04315(.I(new_n4507_), .ZN(new_n4508_));
  AOI21_X1   g04316(.A1(new_n4309_), .A2(new_n4314_), .B(\asqrt[36] ), .ZN(new_n4509_));
  XOR2_X1    g04317(.A1(new_n4509_), .A2(new_n4248_), .Z(new_n4510_));
  AOI21_X1   g04318(.A1(new_n4382_), .A2(new_n4308_), .B(\asqrt[36] ), .ZN(new_n4511_));
  XOR2_X1    g04319(.A1(new_n4511_), .A2(new_n4251_), .Z(new_n4512_));
  XOR2_X1    g04320(.A1(new_n4380_), .A2(\asqrt[43] ), .Z(new_n4513_));
  NOR2_X1    g04321(.A1(\asqrt[36] ), .A2(new_n4513_), .ZN(new_n4514_));
  XOR2_X1    g04322(.A1(new_n4514_), .A2(new_n4253_), .Z(new_n4515_));
  INV_X1     g04323(.I(new_n4515_), .ZN(new_n4516_));
  NOR2_X1    g04324(.A1(new_n4378_), .A2(new_n4303_), .ZN(new_n4517_));
  NOR2_X1    g04325(.A1(\asqrt[36] ), .A2(new_n4517_), .ZN(new_n4518_));
  XOR2_X1    g04326(.A1(new_n4518_), .A2(new_n4257_), .Z(new_n4519_));
  INV_X1     g04327(.I(new_n4519_), .ZN(new_n4520_));
  AOI21_X1   g04328(.A1(new_n4297_), .A2(new_n4302_), .B(\asqrt[36] ), .ZN(new_n4521_));
  XOR2_X1    g04329(.A1(new_n4521_), .A2(new_n4260_), .Z(new_n4522_));
  AOI21_X1   g04330(.A1(new_n4374_), .A2(new_n4296_), .B(\asqrt[36] ), .ZN(new_n4523_));
  XOR2_X1    g04331(.A1(new_n4523_), .A2(new_n4266_), .Z(new_n4524_));
  AOI21_X1   g04332(.A1(new_n4372_), .A2(new_n4293_), .B(\asqrt[36] ), .ZN(new_n4525_));
  XOR2_X1    g04333(.A1(new_n4525_), .A2(new_n4363_), .Z(new_n4526_));
  INV_X1     g04334(.I(new_n4526_), .ZN(new_n4527_));
  NAND2_X1   g04335(.A1(\asqrt[37] ), .A2(new_n4281_), .ZN(new_n4528_));
  NOR2_X1    g04336(.A1(new_n4288_), .A2(\a[74] ), .ZN(new_n4529_));
  AOI22_X1   g04337(.A1(new_n4528_), .A2(new_n4288_), .B1(\asqrt[37] ), .B2(new_n4529_), .ZN(new_n4530_));
  OAI21_X1   g04338(.A1(new_n4196_), .A2(new_n4281_), .B(new_n4367_), .ZN(new_n4531_));
  AOI21_X1   g04339(.A1(new_n4366_), .A2(new_n4531_), .B(\asqrt[36] ), .ZN(new_n4532_));
  XOR2_X1    g04340(.A1(new_n4532_), .A2(new_n4530_), .Z(new_n4533_));
  INV_X1     g04341(.I(new_n4533_), .ZN(new_n4534_));
  NAND2_X1   g04342(.A1(new_n4438_), .A2(new_n193_), .ZN(new_n4535_));
  NAND3_X1   g04343(.A1(new_n4444_), .A2(\asqrt[37] ), .A3(new_n4446_), .ZN(new_n4536_));
  NOR3_X1    g04344(.A1(new_n4535_), .A2(new_n4460_), .A3(new_n4536_), .ZN(new_n4537_));
  NOR2_X1    g04345(.A1(new_n4461_), .A2(new_n4279_), .ZN(new_n4538_));
  OAI21_X1   g04346(.A1(new_n4538_), .A2(new_n4537_), .B(new_n4281_), .ZN(new_n4539_));
  NOR3_X1    g04347(.A1(new_n4457_), .A2(\asqrt[63] ), .A3(new_n4460_), .ZN(new_n4540_));
  NAND4_X1   g04348(.A1(new_n4540_), .A2(\asqrt[37] ), .A3(new_n4444_), .A4(new_n4446_), .ZN(new_n4541_));
  NAND2_X1   g04349(.A1(\asqrt[36] ), .A2(new_n4278_), .ZN(new_n4542_));
  NAND3_X1   g04350(.A1(new_n4541_), .A2(new_n4542_), .A3(\a[74] ), .ZN(new_n4543_));
  NAND2_X1   g04351(.A1(new_n4543_), .A2(new_n4539_), .ZN(new_n4544_));
  INV_X1     g04352(.I(new_n4544_), .ZN(new_n4545_));
  INV_X1     g04353(.I(\a[72] ), .ZN(new_n4546_));
  NOR2_X1    g04354(.A1(\a[70] ), .A2(\a[71] ), .ZN(new_n4547_));
  NOR3_X1    g04355(.A1(new_n4461_), .A2(new_n4546_), .A3(new_n4547_), .ZN(new_n4548_));
  INV_X1     g04356(.I(new_n4547_), .ZN(new_n4549_));
  AOI21_X1   g04357(.A1(new_n4461_), .A2(\a[72] ), .B(new_n4549_), .ZN(new_n4550_));
  OAI21_X1   g04358(.A1(new_n4548_), .A2(new_n4550_), .B(\asqrt[37] ), .ZN(new_n4551_));
  NAND2_X1   g04359(.A1(new_n4547_), .A2(new_n4546_), .ZN(new_n4552_));
  NAND3_X1   g04360(.A1(new_n4178_), .A2(new_n4180_), .A3(new_n4552_), .ZN(new_n4553_));
  NAND2_X1   g04361(.A1(new_n4267_), .A2(new_n4553_), .ZN(new_n4554_));
  INV_X1     g04362(.I(new_n4554_), .ZN(new_n4555_));
  NOR3_X1    g04363(.A1(new_n4461_), .A2(new_n4546_), .A3(new_n4555_), .ZN(new_n4556_));
  NOR3_X1    g04364(.A1(new_n4461_), .A2(\a[72] ), .A3(\a[73] ), .ZN(new_n4557_));
  INV_X1     g04365(.I(\a[73] ), .ZN(new_n4558_));
  AOI21_X1   g04366(.A1(\asqrt[36] ), .A2(new_n4546_), .B(new_n4558_), .ZN(new_n4559_));
  NOR3_X1    g04367(.A1(new_n4556_), .A2(new_n4557_), .A3(new_n4559_), .ZN(new_n4560_));
  NAND3_X1   g04368(.A1(new_n4551_), .A2(new_n4560_), .A3(new_n3925_), .ZN(new_n4561_));
  AOI21_X1   g04369(.A1(new_n4551_), .A2(new_n4560_), .B(new_n3925_), .ZN(new_n4562_));
  AOI21_X1   g04370(.A1(new_n4545_), .A2(new_n4561_), .B(new_n4562_), .ZN(new_n4563_));
  AOI21_X1   g04371(.A1(new_n4563_), .A2(new_n3681_), .B(new_n4534_), .ZN(new_n4564_));
  NAND2_X1   g04372(.A1(new_n4545_), .A2(new_n4561_), .ZN(new_n4565_));
  NAND3_X1   g04373(.A1(\asqrt[36] ), .A2(\a[72] ), .A3(new_n4549_), .ZN(new_n4566_));
  OAI21_X1   g04374(.A1(\asqrt[36] ), .A2(new_n4546_), .B(new_n4547_), .ZN(new_n4567_));
  AOI21_X1   g04375(.A1(new_n4567_), .A2(new_n4566_), .B(new_n4196_), .ZN(new_n4568_));
  NAND3_X1   g04376(.A1(\asqrt[36] ), .A2(\a[72] ), .A3(new_n4554_), .ZN(new_n4569_));
  NAND3_X1   g04377(.A1(\asqrt[36] ), .A2(new_n4546_), .A3(new_n4558_), .ZN(new_n4570_));
  OAI21_X1   g04378(.A1(new_n4461_), .A2(\a[72] ), .B(\a[73] ), .ZN(new_n4571_));
  NAND3_X1   g04379(.A1(new_n4571_), .A2(new_n4569_), .A3(new_n4570_), .ZN(new_n4572_));
  OAI21_X1   g04380(.A1(new_n4572_), .A2(new_n4568_), .B(\asqrt[38] ), .ZN(new_n4573_));
  AOI21_X1   g04381(.A1(new_n4565_), .A2(new_n4573_), .B(new_n3681_), .ZN(new_n4574_));
  NOR3_X1    g04382(.A1(new_n4564_), .A2(\asqrt[40] ), .A3(new_n4574_), .ZN(new_n4575_));
  OAI21_X1   g04383(.A1(new_n4564_), .A2(new_n4574_), .B(\asqrt[40] ), .ZN(new_n4576_));
  OAI21_X1   g04384(.A1(new_n4527_), .A2(new_n4575_), .B(new_n4576_), .ZN(new_n4577_));
  OAI21_X1   g04385(.A1(new_n4577_), .A2(\asqrt[41] ), .B(new_n4524_), .ZN(new_n4578_));
  NAND2_X1   g04386(.A1(new_n4577_), .A2(\asqrt[41] ), .ZN(new_n4579_));
  NAND3_X1   g04387(.A1(new_n4578_), .A2(new_n4579_), .A3(new_n2960_), .ZN(new_n4580_));
  AOI21_X1   g04388(.A1(new_n4578_), .A2(new_n4579_), .B(new_n2960_), .ZN(new_n4581_));
  AOI21_X1   g04389(.A1(new_n4522_), .A2(new_n4580_), .B(new_n4581_), .ZN(new_n4582_));
  AOI21_X1   g04390(.A1(new_n4582_), .A2(new_n2749_), .B(new_n4520_), .ZN(new_n4583_));
  NAND2_X1   g04391(.A1(new_n4580_), .A2(new_n4522_), .ZN(new_n4584_));
  INV_X1     g04392(.I(new_n4524_), .ZN(new_n4585_));
  NOR3_X1    g04393(.A1(new_n4572_), .A2(new_n4568_), .A3(\asqrt[38] ), .ZN(new_n4586_));
  OAI21_X1   g04394(.A1(new_n4544_), .A2(new_n4586_), .B(new_n4573_), .ZN(new_n4587_));
  OAI21_X1   g04395(.A1(new_n4587_), .A2(\asqrt[39] ), .B(new_n4533_), .ZN(new_n4588_));
  NAND2_X1   g04396(.A1(new_n4587_), .A2(\asqrt[39] ), .ZN(new_n4589_));
  NAND3_X1   g04397(.A1(new_n4588_), .A2(new_n4589_), .A3(new_n3427_), .ZN(new_n4590_));
  AOI21_X1   g04398(.A1(new_n4588_), .A2(new_n4589_), .B(new_n3427_), .ZN(new_n4591_));
  AOI21_X1   g04399(.A1(new_n4526_), .A2(new_n4590_), .B(new_n4591_), .ZN(new_n4592_));
  AOI21_X1   g04400(.A1(new_n4592_), .A2(new_n3195_), .B(new_n4585_), .ZN(new_n4593_));
  NAND2_X1   g04401(.A1(new_n4590_), .A2(new_n4526_), .ZN(new_n4594_));
  AOI21_X1   g04402(.A1(new_n4594_), .A2(new_n4576_), .B(new_n3195_), .ZN(new_n4595_));
  OAI21_X1   g04403(.A1(new_n4593_), .A2(new_n4595_), .B(\asqrt[42] ), .ZN(new_n4596_));
  AOI21_X1   g04404(.A1(new_n4584_), .A2(new_n4596_), .B(new_n2749_), .ZN(new_n4597_));
  NOR3_X1    g04405(.A1(new_n4583_), .A2(\asqrt[44] ), .A3(new_n4597_), .ZN(new_n4598_));
  OAI21_X1   g04406(.A1(new_n4583_), .A2(new_n4597_), .B(\asqrt[44] ), .ZN(new_n4599_));
  OAI21_X1   g04407(.A1(new_n4516_), .A2(new_n4598_), .B(new_n4599_), .ZN(new_n4600_));
  OAI21_X1   g04408(.A1(new_n4600_), .A2(\asqrt[45] ), .B(new_n4512_), .ZN(new_n4601_));
  NAND2_X1   g04409(.A1(new_n4600_), .A2(\asqrt[45] ), .ZN(new_n4602_));
  NAND3_X1   g04410(.A1(new_n4601_), .A2(new_n4602_), .A3(new_n2134_), .ZN(new_n4603_));
  AOI21_X1   g04411(.A1(new_n4601_), .A2(new_n4602_), .B(new_n2134_), .ZN(new_n4604_));
  AOI21_X1   g04412(.A1(new_n4510_), .A2(new_n4603_), .B(new_n4604_), .ZN(new_n4605_));
  AOI21_X1   g04413(.A1(new_n4605_), .A2(new_n1953_), .B(new_n4508_), .ZN(new_n4606_));
  NAND2_X1   g04414(.A1(new_n4603_), .A2(new_n4510_), .ZN(new_n4607_));
  INV_X1     g04415(.I(new_n4512_), .ZN(new_n4608_));
  INV_X1     g04416(.I(new_n4522_), .ZN(new_n4609_));
  NOR3_X1    g04417(.A1(new_n4593_), .A2(\asqrt[42] ), .A3(new_n4595_), .ZN(new_n4610_));
  OAI21_X1   g04418(.A1(new_n4609_), .A2(new_n4610_), .B(new_n4596_), .ZN(new_n4611_));
  OAI21_X1   g04419(.A1(new_n4611_), .A2(\asqrt[43] ), .B(new_n4519_), .ZN(new_n4612_));
  NAND2_X1   g04420(.A1(new_n4611_), .A2(\asqrt[43] ), .ZN(new_n4613_));
  NAND3_X1   g04421(.A1(new_n4612_), .A2(new_n4613_), .A3(new_n2531_), .ZN(new_n4614_));
  AOI21_X1   g04422(.A1(new_n4612_), .A2(new_n4613_), .B(new_n2531_), .ZN(new_n4615_));
  AOI21_X1   g04423(.A1(new_n4515_), .A2(new_n4614_), .B(new_n4615_), .ZN(new_n4616_));
  AOI21_X1   g04424(.A1(new_n4616_), .A2(new_n2332_), .B(new_n4608_), .ZN(new_n4617_));
  NAND2_X1   g04425(.A1(new_n4614_), .A2(new_n4515_), .ZN(new_n4618_));
  AOI21_X1   g04426(.A1(new_n4618_), .A2(new_n4599_), .B(new_n2332_), .ZN(new_n4619_));
  OAI21_X1   g04427(.A1(new_n4617_), .A2(new_n4619_), .B(\asqrt[46] ), .ZN(new_n4620_));
  AOI21_X1   g04428(.A1(new_n4607_), .A2(new_n4620_), .B(new_n1953_), .ZN(new_n4621_));
  NOR3_X1    g04429(.A1(new_n4606_), .A2(\asqrt[48] ), .A3(new_n4621_), .ZN(new_n4622_));
  OAI21_X1   g04430(.A1(new_n4606_), .A2(new_n4621_), .B(\asqrt[48] ), .ZN(new_n4623_));
  OAI21_X1   g04431(.A1(new_n4504_), .A2(new_n4622_), .B(new_n4623_), .ZN(new_n4624_));
  OAI21_X1   g04432(.A1(new_n4624_), .A2(\asqrt[49] ), .B(new_n4500_), .ZN(new_n4625_));
  NAND2_X1   g04433(.A1(new_n4624_), .A2(\asqrt[49] ), .ZN(new_n4626_));
  NAND3_X1   g04434(.A1(new_n4625_), .A2(new_n4626_), .A3(new_n1463_), .ZN(new_n4627_));
  AOI21_X1   g04435(.A1(new_n4625_), .A2(new_n4626_), .B(new_n1463_), .ZN(new_n4628_));
  AOI21_X1   g04436(.A1(new_n4498_), .A2(new_n4627_), .B(new_n4628_), .ZN(new_n4629_));
  AOI21_X1   g04437(.A1(new_n4629_), .A2(new_n1305_), .B(new_n4496_), .ZN(new_n4630_));
  NAND2_X1   g04438(.A1(new_n4627_), .A2(new_n4498_), .ZN(new_n4631_));
  INV_X1     g04439(.I(new_n4500_), .ZN(new_n4632_));
  INV_X1     g04440(.I(new_n4510_), .ZN(new_n4633_));
  NOR3_X1    g04441(.A1(new_n4617_), .A2(\asqrt[46] ), .A3(new_n4619_), .ZN(new_n4634_));
  OAI21_X1   g04442(.A1(new_n4633_), .A2(new_n4634_), .B(new_n4620_), .ZN(new_n4635_));
  OAI21_X1   g04443(.A1(new_n4635_), .A2(\asqrt[47] ), .B(new_n4507_), .ZN(new_n4636_));
  NAND2_X1   g04444(.A1(new_n4635_), .A2(\asqrt[47] ), .ZN(new_n4637_));
  NAND3_X1   g04445(.A1(new_n4636_), .A2(new_n4637_), .A3(new_n1778_), .ZN(new_n4638_));
  AOI21_X1   g04446(.A1(new_n4636_), .A2(new_n4637_), .B(new_n1778_), .ZN(new_n4639_));
  AOI21_X1   g04447(.A1(new_n4503_), .A2(new_n4638_), .B(new_n4639_), .ZN(new_n4640_));
  AOI21_X1   g04448(.A1(new_n4640_), .A2(new_n1632_), .B(new_n4632_), .ZN(new_n4641_));
  NAND2_X1   g04449(.A1(new_n4638_), .A2(new_n4503_), .ZN(new_n4642_));
  AOI21_X1   g04450(.A1(new_n4642_), .A2(new_n4623_), .B(new_n1632_), .ZN(new_n4643_));
  OAI21_X1   g04451(.A1(new_n4641_), .A2(new_n4643_), .B(\asqrt[50] ), .ZN(new_n4644_));
  AOI21_X1   g04452(.A1(new_n4631_), .A2(new_n4644_), .B(new_n1305_), .ZN(new_n4645_));
  NOR3_X1    g04453(.A1(new_n4630_), .A2(\asqrt[52] ), .A3(new_n4645_), .ZN(new_n4646_));
  OAI21_X1   g04454(.A1(new_n4630_), .A2(new_n4645_), .B(\asqrt[52] ), .ZN(new_n4647_));
  OAI21_X1   g04455(.A1(new_n4492_), .A2(new_n4646_), .B(new_n4647_), .ZN(new_n4648_));
  OAI21_X1   g04456(.A1(new_n4648_), .A2(\asqrt[53] ), .B(new_n4488_), .ZN(new_n4649_));
  NAND2_X1   g04457(.A1(new_n4648_), .A2(\asqrt[53] ), .ZN(new_n4650_));
  NAND3_X1   g04458(.A1(new_n4649_), .A2(new_n4650_), .A3(new_n860_), .ZN(new_n4651_));
  AOI21_X1   g04459(.A1(new_n4649_), .A2(new_n4650_), .B(new_n860_), .ZN(new_n4652_));
  AOI21_X1   g04460(.A1(new_n4486_), .A2(new_n4651_), .B(new_n4652_), .ZN(new_n4653_));
  AOI21_X1   g04461(.A1(new_n4653_), .A2(new_n744_), .B(new_n4484_), .ZN(new_n4654_));
  NAND2_X1   g04462(.A1(new_n4651_), .A2(new_n4486_), .ZN(new_n4655_));
  INV_X1     g04463(.I(new_n4488_), .ZN(new_n4656_));
  INV_X1     g04464(.I(new_n4498_), .ZN(new_n4657_));
  NOR3_X1    g04465(.A1(new_n4641_), .A2(\asqrt[50] ), .A3(new_n4643_), .ZN(new_n4658_));
  OAI21_X1   g04466(.A1(new_n4657_), .A2(new_n4658_), .B(new_n4644_), .ZN(new_n4659_));
  OAI21_X1   g04467(.A1(new_n4659_), .A2(\asqrt[51] ), .B(new_n4495_), .ZN(new_n4660_));
  NAND2_X1   g04468(.A1(new_n4659_), .A2(\asqrt[51] ), .ZN(new_n4661_));
  NAND3_X1   g04469(.A1(new_n4660_), .A2(new_n4661_), .A3(new_n1150_), .ZN(new_n4662_));
  AOI21_X1   g04470(.A1(new_n4660_), .A2(new_n4661_), .B(new_n1150_), .ZN(new_n4663_));
  AOI21_X1   g04471(.A1(new_n4491_), .A2(new_n4662_), .B(new_n4663_), .ZN(new_n4664_));
  AOI21_X1   g04472(.A1(new_n4664_), .A2(new_n1006_), .B(new_n4656_), .ZN(new_n4665_));
  NAND2_X1   g04473(.A1(new_n4662_), .A2(new_n4491_), .ZN(new_n4666_));
  AOI21_X1   g04474(.A1(new_n4666_), .A2(new_n4647_), .B(new_n1006_), .ZN(new_n4667_));
  OAI21_X1   g04475(.A1(new_n4665_), .A2(new_n4667_), .B(\asqrt[54] ), .ZN(new_n4668_));
  AOI21_X1   g04476(.A1(new_n4655_), .A2(new_n4668_), .B(new_n744_), .ZN(new_n4669_));
  NOR3_X1    g04477(.A1(new_n4654_), .A2(\asqrt[56] ), .A3(new_n4669_), .ZN(new_n4670_));
  OAI21_X1   g04478(.A1(new_n4654_), .A2(new_n4669_), .B(\asqrt[56] ), .ZN(new_n4671_));
  OAI21_X1   g04479(.A1(new_n4480_), .A2(new_n4670_), .B(new_n4671_), .ZN(new_n4672_));
  OAI21_X1   g04480(.A1(new_n4672_), .A2(\asqrt[57] ), .B(new_n4475_), .ZN(new_n4673_));
  NOR2_X1    g04481(.A1(new_n4670_), .A2(new_n4480_), .ZN(new_n4674_));
  INV_X1     g04482(.I(new_n4486_), .ZN(new_n4675_));
  NOR3_X1    g04483(.A1(new_n4665_), .A2(\asqrt[54] ), .A3(new_n4667_), .ZN(new_n4676_));
  OAI21_X1   g04484(.A1(new_n4675_), .A2(new_n4676_), .B(new_n4668_), .ZN(new_n4677_));
  OAI21_X1   g04485(.A1(new_n4677_), .A2(\asqrt[55] ), .B(new_n4483_), .ZN(new_n4678_));
  NAND2_X1   g04486(.A1(new_n4677_), .A2(\asqrt[55] ), .ZN(new_n4679_));
  AOI21_X1   g04487(.A1(new_n4678_), .A2(new_n4679_), .B(new_n634_), .ZN(new_n4680_));
  OAI21_X1   g04488(.A1(new_n4674_), .A2(new_n4680_), .B(\asqrt[57] ), .ZN(new_n4681_));
  NAND3_X1   g04489(.A1(new_n4673_), .A2(new_n423_), .A3(new_n4681_), .ZN(new_n4682_));
  NAND2_X1   g04490(.A1(new_n4682_), .A2(new_n4473_), .ZN(new_n4683_));
  INV_X1     g04491(.I(new_n4475_), .ZN(new_n4684_));
  NAND3_X1   g04492(.A1(new_n4678_), .A2(new_n4679_), .A3(new_n634_), .ZN(new_n4685_));
  AOI21_X1   g04493(.A1(new_n4479_), .A2(new_n4685_), .B(new_n4680_), .ZN(new_n4686_));
  AOI21_X1   g04494(.A1(new_n4686_), .A2(new_n531_), .B(new_n4684_), .ZN(new_n4687_));
  NAND2_X1   g04495(.A1(new_n4685_), .A2(new_n4479_), .ZN(new_n4688_));
  AOI21_X1   g04496(.A1(new_n4688_), .A2(new_n4671_), .B(new_n531_), .ZN(new_n4689_));
  OAI21_X1   g04497(.A1(new_n4687_), .A2(new_n4689_), .B(\asqrt[58] ), .ZN(new_n4690_));
  NAND3_X1   g04498(.A1(new_n4683_), .A2(new_n337_), .A3(new_n4690_), .ZN(new_n4691_));
  AOI21_X1   g04499(.A1(new_n4683_), .A2(new_n4690_), .B(new_n337_), .ZN(new_n4692_));
  AOI21_X1   g04500(.A1(new_n4471_), .A2(new_n4691_), .B(new_n4692_), .ZN(new_n4693_));
  AOI21_X1   g04501(.A1(new_n4693_), .A2(new_n266_), .B(new_n4468_), .ZN(new_n4694_));
  INV_X1     g04502(.I(new_n4473_), .ZN(new_n4695_));
  NOR3_X1    g04503(.A1(new_n4687_), .A2(\asqrt[58] ), .A3(new_n4689_), .ZN(new_n4696_));
  OAI21_X1   g04504(.A1(new_n4695_), .A2(new_n4696_), .B(new_n4690_), .ZN(new_n4697_));
  OAI21_X1   g04505(.A1(new_n4697_), .A2(\asqrt[59] ), .B(new_n4471_), .ZN(new_n4698_));
  NAND2_X1   g04506(.A1(new_n4697_), .A2(\asqrt[59] ), .ZN(new_n4699_));
  AOI21_X1   g04507(.A1(new_n4698_), .A2(new_n4699_), .B(new_n266_), .ZN(new_n4700_));
  OAI21_X1   g04508(.A1(new_n4694_), .A2(new_n4700_), .B(\asqrt[61] ), .ZN(new_n4701_));
  AOI21_X1   g04509(.A1(new_n4425_), .A2(new_n4420_), .B(\asqrt[36] ), .ZN(new_n4702_));
  XOR2_X1    g04510(.A1(new_n4702_), .A2(new_n4202_), .Z(new_n4703_));
  INV_X1     g04511(.I(new_n4703_), .ZN(new_n4704_));
  NOR3_X1    g04512(.A1(new_n4694_), .A2(\asqrt[61] ), .A3(new_n4700_), .ZN(new_n4705_));
  OAI21_X1   g04513(.A1(new_n4704_), .A2(new_n4705_), .B(new_n4701_), .ZN(new_n4706_));
  NAND3_X1   g04514(.A1(new_n4698_), .A2(new_n4699_), .A3(new_n266_), .ZN(new_n4707_));
  NAND2_X1   g04515(.A1(new_n4707_), .A2(new_n4467_), .ZN(new_n4708_));
  INV_X1     g04516(.I(new_n4471_), .ZN(new_n4709_));
  AOI21_X1   g04517(.A1(new_n4673_), .A2(new_n4681_), .B(new_n423_), .ZN(new_n4710_));
  AOI21_X1   g04518(.A1(new_n4473_), .A2(new_n4682_), .B(new_n4710_), .ZN(new_n4711_));
  AOI21_X1   g04519(.A1(new_n4711_), .A2(new_n337_), .B(new_n4709_), .ZN(new_n4712_));
  OAI21_X1   g04520(.A1(new_n4712_), .A2(new_n4692_), .B(\asqrt[60] ), .ZN(new_n4713_));
  AOI21_X1   g04521(.A1(new_n4708_), .A2(new_n4713_), .B(new_n239_), .ZN(new_n4714_));
  AOI21_X1   g04522(.A1(new_n4467_), .A2(new_n4707_), .B(new_n4700_), .ZN(new_n4715_));
  AOI21_X1   g04523(.A1(new_n4715_), .A2(new_n239_), .B(new_n4704_), .ZN(new_n4716_));
  OAI21_X1   g04524(.A1(new_n4716_), .A2(new_n4714_), .B(new_n201_), .ZN(new_n4717_));
  NOR3_X1    g04525(.A1(new_n4712_), .A2(\asqrt[60] ), .A3(new_n4692_), .ZN(new_n4718_));
  OAI21_X1   g04526(.A1(new_n4468_), .A2(new_n4718_), .B(new_n4713_), .ZN(new_n4719_));
  OAI21_X1   g04527(.A1(new_n4719_), .A2(\asqrt[61] ), .B(new_n4703_), .ZN(new_n4720_));
  NAND3_X1   g04528(.A1(new_n4720_), .A2(\asqrt[62] ), .A3(new_n4701_), .ZN(new_n4721_));
  AOI21_X1   g04529(.A1(new_n4415_), .A2(new_n4421_), .B(\asqrt[36] ), .ZN(new_n4722_));
  XOR2_X1    g04530(.A1(new_n4722_), .A2(new_n4417_), .Z(new_n4723_));
  INV_X1     g04531(.I(new_n4723_), .ZN(new_n4724_));
  AOI22_X1   g04532(.A1(new_n4721_), .A2(new_n4717_), .B1(new_n4706_), .B2(new_n4724_), .ZN(new_n4725_));
  NOR2_X1    g04533(.A1(new_n4434_), .A2(new_n4199_), .ZN(new_n4726_));
  OAI21_X1   g04534(.A1(\asqrt[36] ), .A2(new_n4726_), .B(new_n4441_), .ZN(new_n4727_));
  INV_X1     g04535(.I(new_n4727_), .ZN(new_n4728_));
  OAI21_X1   g04536(.A1(new_n4725_), .A2(new_n4464_), .B(new_n4728_), .ZN(new_n4729_));
  OAI21_X1   g04537(.A1(new_n4706_), .A2(\asqrt[62] ), .B(new_n4723_), .ZN(new_n4730_));
  NAND2_X1   g04538(.A1(new_n4706_), .A2(\asqrt[62] ), .ZN(new_n4731_));
  NAND3_X1   g04539(.A1(new_n4730_), .A2(new_n4731_), .A3(new_n4464_), .ZN(new_n4732_));
  NAND2_X1   g04540(.A1(new_n4461_), .A2(new_n4198_), .ZN(new_n4733_));
  XOR2_X1    g04541(.A1(new_n4434_), .A2(new_n4199_), .Z(new_n4734_));
  NAND3_X1   g04542(.A1(new_n4733_), .A2(\asqrt[63] ), .A3(new_n4734_), .ZN(new_n4735_));
  INV_X1     g04543(.I(new_n4535_), .ZN(new_n4736_));
  NAND4_X1   g04544(.A1(new_n4736_), .A2(new_n4199_), .A3(new_n4441_), .A4(new_n4448_), .ZN(new_n4737_));
  NAND2_X1   g04545(.A1(new_n4735_), .A2(new_n4737_), .ZN(new_n4738_));
  INV_X1     g04546(.I(new_n4738_), .ZN(new_n4739_));
  NAND4_X1   g04547(.A1(new_n4729_), .A2(new_n193_), .A3(new_n4732_), .A4(new_n4739_), .ZN(\asqrt[35] ));
  NOR2_X1    g04548(.A1(new_n4706_), .A2(\asqrt[62] ), .ZN(new_n4741_));
  NOR2_X1    g04549(.A1(new_n4716_), .A2(new_n4714_), .ZN(new_n4742_));
  NOR2_X1    g04550(.A1(new_n4742_), .A2(new_n201_), .ZN(new_n4743_));
  NOR2_X1    g04551(.A1(new_n4741_), .A2(new_n4743_), .ZN(new_n4744_));
  AOI21_X1   g04552(.A1(new_n4720_), .A2(new_n4701_), .B(\asqrt[62] ), .ZN(new_n4745_));
  NOR3_X1    g04553(.A1(new_n4716_), .A2(new_n201_), .A3(new_n4714_), .ZN(new_n4746_));
  OAI22_X1   g04554(.A1(new_n4745_), .A2(new_n4746_), .B1(new_n4742_), .B2(new_n4723_), .ZN(new_n4747_));
  AOI21_X1   g04555(.A1(new_n4747_), .A2(new_n4463_), .B(new_n4727_), .ZN(new_n4748_));
  AOI21_X1   g04556(.A1(new_n4742_), .A2(new_n201_), .B(new_n4724_), .ZN(new_n4749_));
  NOR3_X1    g04557(.A1(new_n4749_), .A2(new_n4743_), .A3(new_n4463_), .ZN(new_n4750_));
  NOR4_X1    g04558(.A1(new_n4748_), .A2(\asqrt[63] ), .A3(new_n4750_), .A4(new_n4738_), .ZN(new_n4751_));
  XOR2_X1    g04559(.A1(new_n4722_), .A2(new_n4417_), .Z(new_n4752_));
  OAI21_X1   g04560(.A1(\asqrt[35] ), .A2(new_n4744_), .B(new_n4752_), .ZN(new_n4753_));
  INV_X1     g04561(.I(new_n4753_), .ZN(new_n4754_));
  AOI21_X1   g04562(.A1(new_n4691_), .A2(new_n4699_), .B(\asqrt[35] ), .ZN(new_n4755_));
  XOR2_X1    g04563(.A1(new_n4755_), .A2(new_n4471_), .Z(new_n4756_));
  INV_X1     g04564(.I(new_n4756_), .ZN(new_n4757_));
  AOI21_X1   g04565(.A1(new_n4682_), .A2(new_n4690_), .B(\asqrt[35] ), .ZN(new_n4758_));
  XOR2_X1    g04566(.A1(new_n4758_), .A2(new_n4473_), .Z(new_n4759_));
  INV_X1     g04567(.I(new_n4759_), .ZN(new_n4760_));
  NAND2_X1   g04568(.A1(new_n4686_), .A2(new_n531_), .ZN(new_n4761_));
  AOI21_X1   g04569(.A1(new_n4761_), .A2(new_n4681_), .B(\asqrt[35] ), .ZN(new_n4762_));
  XOR2_X1    g04570(.A1(new_n4762_), .A2(new_n4475_), .Z(new_n4763_));
  AOI21_X1   g04571(.A1(new_n4685_), .A2(new_n4671_), .B(\asqrt[35] ), .ZN(new_n4764_));
  XOR2_X1    g04572(.A1(new_n4764_), .A2(new_n4479_), .Z(new_n4765_));
  NAND2_X1   g04573(.A1(new_n4653_), .A2(new_n744_), .ZN(new_n4766_));
  AOI21_X1   g04574(.A1(new_n4766_), .A2(new_n4679_), .B(\asqrt[35] ), .ZN(new_n4767_));
  XOR2_X1    g04575(.A1(new_n4767_), .A2(new_n4483_), .Z(new_n4768_));
  INV_X1     g04576(.I(new_n4768_), .ZN(new_n4769_));
  AOI21_X1   g04577(.A1(new_n4651_), .A2(new_n4668_), .B(\asqrt[35] ), .ZN(new_n4770_));
  XOR2_X1    g04578(.A1(new_n4770_), .A2(new_n4486_), .Z(new_n4771_));
  INV_X1     g04579(.I(new_n4771_), .ZN(new_n4772_));
  NAND2_X1   g04580(.A1(new_n4664_), .A2(new_n1006_), .ZN(new_n4773_));
  AOI21_X1   g04581(.A1(new_n4773_), .A2(new_n4650_), .B(\asqrt[35] ), .ZN(new_n4774_));
  XOR2_X1    g04582(.A1(new_n4774_), .A2(new_n4488_), .Z(new_n4775_));
  AOI21_X1   g04583(.A1(new_n4662_), .A2(new_n4647_), .B(\asqrt[35] ), .ZN(new_n4776_));
  XOR2_X1    g04584(.A1(new_n4776_), .A2(new_n4491_), .Z(new_n4777_));
  NAND2_X1   g04585(.A1(new_n4629_), .A2(new_n1305_), .ZN(new_n4778_));
  AOI21_X1   g04586(.A1(new_n4778_), .A2(new_n4661_), .B(\asqrt[35] ), .ZN(new_n4779_));
  XOR2_X1    g04587(.A1(new_n4779_), .A2(new_n4495_), .Z(new_n4780_));
  INV_X1     g04588(.I(new_n4780_), .ZN(new_n4781_));
  AOI21_X1   g04589(.A1(new_n4627_), .A2(new_n4644_), .B(\asqrt[35] ), .ZN(new_n4782_));
  XOR2_X1    g04590(.A1(new_n4782_), .A2(new_n4498_), .Z(new_n4783_));
  INV_X1     g04591(.I(new_n4783_), .ZN(new_n4784_));
  NAND2_X1   g04592(.A1(new_n4640_), .A2(new_n1632_), .ZN(new_n4785_));
  AOI21_X1   g04593(.A1(new_n4785_), .A2(new_n4626_), .B(\asqrt[35] ), .ZN(new_n4786_));
  XOR2_X1    g04594(.A1(new_n4786_), .A2(new_n4500_), .Z(new_n4787_));
  AOI21_X1   g04595(.A1(new_n4638_), .A2(new_n4623_), .B(\asqrt[35] ), .ZN(new_n4788_));
  XOR2_X1    g04596(.A1(new_n4788_), .A2(new_n4503_), .Z(new_n4789_));
  NAND2_X1   g04597(.A1(new_n4605_), .A2(new_n1953_), .ZN(new_n4790_));
  AOI21_X1   g04598(.A1(new_n4790_), .A2(new_n4637_), .B(\asqrt[35] ), .ZN(new_n4791_));
  XOR2_X1    g04599(.A1(new_n4791_), .A2(new_n4507_), .Z(new_n4792_));
  INV_X1     g04600(.I(new_n4792_), .ZN(new_n4793_));
  AOI21_X1   g04601(.A1(new_n4603_), .A2(new_n4620_), .B(\asqrt[35] ), .ZN(new_n4794_));
  XOR2_X1    g04602(.A1(new_n4794_), .A2(new_n4510_), .Z(new_n4795_));
  INV_X1     g04603(.I(new_n4795_), .ZN(new_n4796_));
  NAND2_X1   g04604(.A1(new_n4616_), .A2(new_n2332_), .ZN(new_n4797_));
  AOI21_X1   g04605(.A1(new_n4797_), .A2(new_n4602_), .B(\asqrt[35] ), .ZN(new_n4798_));
  XOR2_X1    g04606(.A1(new_n4798_), .A2(new_n4512_), .Z(new_n4799_));
  AOI21_X1   g04607(.A1(new_n4614_), .A2(new_n4599_), .B(\asqrt[35] ), .ZN(new_n4800_));
  XOR2_X1    g04608(.A1(new_n4800_), .A2(new_n4515_), .Z(new_n4801_));
  NAND2_X1   g04609(.A1(new_n4582_), .A2(new_n2749_), .ZN(new_n4802_));
  AOI21_X1   g04610(.A1(new_n4802_), .A2(new_n4613_), .B(\asqrt[35] ), .ZN(new_n4803_));
  XOR2_X1    g04611(.A1(new_n4803_), .A2(new_n4519_), .Z(new_n4804_));
  INV_X1     g04612(.I(new_n4804_), .ZN(new_n4805_));
  AOI21_X1   g04613(.A1(new_n4580_), .A2(new_n4596_), .B(\asqrt[35] ), .ZN(new_n4806_));
  XOR2_X1    g04614(.A1(new_n4806_), .A2(new_n4522_), .Z(new_n4807_));
  INV_X1     g04615(.I(new_n4807_), .ZN(new_n4808_));
  NAND2_X1   g04616(.A1(new_n4592_), .A2(new_n3195_), .ZN(new_n4809_));
  AOI21_X1   g04617(.A1(new_n4809_), .A2(new_n4579_), .B(\asqrt[35] ), .ZN(new_n4810_));
  XOR2_X1    g04618(.A1(new_n4810_), .A2(new_n4524_), .Z(new_n4811_));
  AOI21_X1   g04619(.A1(new_n4590_), .A2(new_n4576_), .B(\asqrt[35] ), .ZN(new_n4812_));
  XOR2_X1    g04620(.A1(new_n4812_), .A2(new_n4526_), .Z(new_n4813_));
  NAND2_X1   g04621(.A1(new_n4563_), .A2(new_n3681_), .ZN(new_n4814_));
  AOI21_X1   g04622(.A1(new_n4814_), .A2(new_n4589_), .B(\asqrt[35] ), .ZN(new_n4815_));
  XOR2_X1    g04623(.A1(new_n4815_), .A2(new_n4533_), .Z(new_n4816_));
  INV_X1     g04624(.I(new_n4816_), .ZN(new_n4817_));
  AOI21_X1   g04625(.A1(new_n4561_), .A2(new_n4573_), .B(\asqrt[35] ), .ZN(new_n4818_));
  XOR2_X1    g04626(.A1(new_n4818_), .A2(new_n4545_), .Z(new_n4819_));
  INV_X1     g04627(.I(new_n4819_), .ZN(new_n4820_));
  NAND2_X1   g04628(.A1(\asqrt[36] ), .A2(new_n4546_), .ZN(new_n4821_));
  NOR2_X1    g04629(.A1(new_n4558_), .A2(\a[72] ), .ZN(new_n4822_));
  AOI22_X1   g04630(.A1(new_n4821_), .A2(new_n4558_), .B1(\asqrt[36] ), .B2(new_n4822_), .ZN(new_n4823_));
  AOI21_X1   g04631(.A1(\asqrt[36] ), .A2(\a[72] ), .B(new_n4554_), .ZN(new_n4824_));
  OAI21_X1   g04632(.A1(new_n4568_), .A2(new_n4824_), .B(new_n4751_), .ZN(new_n4825_));
  XNOR2_X1   g04633(.A1(new_n4825_), .A2(new_n4823_), .ZN(new_n4826_));
  NAND3_X1   g04634(.A1(new_n4735_), .A2(\asqrt[36] ), .A3(new_n4737_), .ZN(new_n4827_));
  NOR4_X1    g04635(.A1(new_n4748_), .A2(\asqrt[63] ), .A3(new_n4750_), .A4(new_n4827_), .ZN(new_n4828_));
  INV_X1     g04636(.I(new_n4828_), .ZN(new_n4829_));
  NAND2_X1   g04637(.A1(\asqrt[35] ), .A2(new_n4547_), .ZN(new_n4830_));
  AOI21_X1   g04638(.A1(new_n4830_), .A2(new_n4829_), .B(\a[72] ), .ZN(new_n4831_));
  NOR2_X1    g04639(.A1(new_n4751_), .A2(new_n4549_), .ZN(new_n4832_));
  NOR3_X1    g04640(.A1(new_n4832_), .A2(new_n4546_), .A3(new_n4828_), .ZN(new_n4833_));
  NOR2_X1    g04641(.A1(new_n4833_), .A2(new_n4831_), .ZN(new_n4834_));
  INV_X1     g04642(.I(\a[70] ), .ZN(new_n4835_));
  NOR2_X1    g04643(.A1(\a[68] ), .A2(\a[69] ), .ZN(new_n4836_));
  NOR3_X1    g04644(.A1(new_n4751_), .A2(new_n4835_), .A3(new_n4836_), .ZN(new_n4837_));
  INV_X1     g04645(.I(new_n4836_), .ZN(new_n4838_));
  AOI21_X1   g04646(.A1(new_n4751_), .A2(\a[70] ), .B(new_n4838_), .ZN(new_n4839_));
  OAI21_X1   g04647(.A1(new_n4837_), .A2(new_n4839_), .B(\asqrt[36] ), .ZN(new_n4840_));
  NAND2_X1   g04648(.A1(new_n4836_), .A2(new_n4835_), .ZN(new_n4841_));
  NAND3_X1   g04649(.A1(new_n4444_), .A2(new_n4446_), .A3(new_n4841_), .ZN(new_n4842_));
  NAND2_X1   g04650(.A1(new_n4540_), .A2(new_n4842_), .ZN(new_n4843_));
  NAND3_X1   g04651(.A1(\asqrt[35] ), .A2(\a[70] ), .A3(new_n4843_), .ZN(new_n4844_));
  NOR3_X1    g04652(.A1(new_n4751_), .A2(\a[70] ), .A3(\a[71] ), .ZN(new_n4845_));
  INV_X1     g04653(.I(\a[71] ), .ZN(new_n4846_));
  AOI21_X1   g04654(.A1(\asqrt[35] ), .A2(new_n4835_), .B(new_n4846_), .ZN(new_n4847_));
  NOR2_X1    g04655(.A1(new_n4845_), .A2(new_n4847_), .ZN(new_n4848_));
  NAND4_X1   g04656(.A1(new_n4840_), .A2(new_n4848_), .A3(new_n4196_), .A4(new_n4844_), .ZN(new_n4849_));
  NAND2_X1   g04657(.A1(new_n4849_), .A2(new_n4834_), .ZN(new_n4850_));
  NAND3_X1   g04658(.A1(\asqrt[35] ), .A2(\a[70] ), .A3(new_n4838_), .ZN(new_n4851_));
  OAI21_X1   g04659(.A1(\asqrt[35] ), .A2(new_n4835_), .B(new_n4836_), .ZN(new_n4852_));
  AOI21_X1   g04660(.A1(new_n4852_), .A2(new_n4851_), .B(new_n4461_), .ZN(new_n4853_));
  NAND3_X1   g04661(.A1(\asqrt[35] ), .A2(new_n4835_), .A3(new_n4846_), .ZN(new_n4854_));
  OAI21_X1   g04662(.A1(new_n4751_), .A2(\a[70] ), .B(\a[71] ), .ZN(new_n4855_));
  NAND3_X1   g04663(.A1(new_n4844_), .A2(new_n4855_), .A3(new_n4854_), .ZN(new_n4856_));
  OAI21_X1   g04664(.A1(new_n4856_), .A2(new_n4853_), .B(\asqrt[37] ), .ZN(new_n4857_));
  NAND3_X1   g04665(.A1(new_n4850_), .A2(new_n3925_), .A3(new_n4857_), .ZN(new_n4858_));
  AOI21_X1   g04666(.A1(new_n4850_), .A2(new_n4857_), .B(new_n3925_), .ZN(new_n4859_));
  AOI21_X1   g04667(.A1(new_n4826_), .A2(new_n4858_), .B(new_n4859_), .ZN(new_n4860_));
  AOI21_X1   g04668(.A1(new_n4860_), .A2(new_n3681_), .B(new_n4820_), .ZN(new_n4861_));
  OR2_X2     g04669(.A1(new_n4833_), .A2(new_n4831_), .Z(new_n4862_));
  NOR3_X1    g04670(.A1(new_n4856_), .A2(new_n4853_), .A3(\asqrt[37] ), .ZN(new_n4863_));
  OAI21_X1   g04671(.A1(new_n4862_), .A2(new_n4863_), .B(new_n4857_), .ZN(new_n4864_));
  OAI21_X1   g04672(.A1(new_n4864_), .A2(\asqrt[38] ), .B(new_n4826_), .ZN(new_n4865_));
  NAND2_X1   g04673(.A1(new_n4864_), .A2(\asqrt[38] ), .ZN(new_n4866_));
  AOI21_X1   g04674(.A1(new_n4865_), .A2(new_n4866_), .B(new_n3681_), .ZN(new_n4867_));
  NOR3_X1    g04675(.A1(new_n4861_), .A2(\asqrt[40] ), .A3(new_n4867_), .ZN(new_n4868_));
  OAI21_X1   g04676(.A1(new_n4861_), .A2(new_n4867_), .B(\asqrt[40] ), .ZN(new_n4869_));
  OAI21_X1   g04677(.A1(new_n4817_), .A2(new_n4868_), .B(new_n4869_), .ZN(new_n4870_));
  OAI21_X1   g04678(.A1(new_n4870_), .A2(\asqrt[41] ), .B(new_n4813_), .ZN(new_n4871_));
  NAND3_X1   g04679(.A1(new_n4865_), .A2(new_n4866_), .A3(new_n3681_), .ZN(new_n4872_));
  AOI21_X1   g04680(.A1(new_n4819_), .A2(new_n4872_), .B(new_n4867_), .ZN(new_n4873_));
  AOI21_X1   g04681(.A1(new_n4873_), .A2(new_n3427_), .B(new_n4817_), .ZN(new_n4874_));
  NAND2_X1   g04682(.A1(new_n4872_), .A2(new_n4819_), .ZN(new_n4875_));
  INV_X1     g04683(.I(new_n4867_), .ZN(new_n4876_));
  AOI21_X1   g04684(.A1(new_n4875_), .A2(new_n4876_), .B(new_n3427_), .ZN(new_n4877_));
  OAI21_X1   g04685(.A1(new_n4874_), .A2(new_n4877_), .B(\asqrt[41] ), .ZN(new_n4878_));
  NAND3_X1   g04686(.A1(new_n4871_), .A2(new_n2960_), .A3(new_n4878_), .ZN(new_n4879_));
  AOI21_X1   g04687(.A1(new_n4871_), .A2(new_n4878_), .B(new_n2960_), .ZN(new_n4880_));
  AOI21_X1   g04688(.A1(new_n4811_), .A2(new_n4879_), .B(new_n4880_), .ZN(new_n4881_));
  AOI21_X1   g04689(.A1(new_n4881_), .A2(new_n2749_), .B(new_n4808_), .ZN(new_n4882_));
  INV_X1     g04690(.I(new_n4813_), .ZN(new_n4883_));
  NOR3_X1    g04691(.A1(new_n4874_), .A2(\asqrt[41] ), .A3(new_n4877_), .ZN(new_n4884_));
  OAI21_X1   g04692(.A1(new_n4883_), .A2(new_n4884_), .B(new_n4878_), .ZN(new_n4885_));
  OAI21_X1   g04693(.A1(new_n4885_), .A2(\asqrt[42] ), .B(new_n4811_), .ZN(new_n4886_));
  NAND2_X1   g04694(.A1(new_n4885_), .A2(\asqrt[42] ), .ZN(new_n4887_));
  AOI21_X1   g04695(.A1(new_n4886_), .A2(new_n4887_), .B(new_n2749_), .ZN(new_n4888_));
  NOR3_X1    g04696(.A1(new_n4882_), .A2(\asqrt[44] ), .A3(new_n4888_), .ZN(new_n4889_));
  OAI21_X1   g04697(.A1(new_n4882_), .A2(new_n4888_), .B(\asqrt[44] ), .ZN(new_n4890_));
  OAI21_X1   g04698(.A1(new_n4805_), .A2(new_n4889_), .B(new_n4890_), .ZN(new_n4891_));
  OAI21_X1   g04699(.A1(new_n4891_), .A2(\asqrt[45] ), .B(new_n4801_), .ZN(new_n4892_));
  NAND3_X1   g04700(.A1(new_n4886_), .A2(new_n4887_), .A3(new_n2749_), .ZN(new_n4893_));
  AOI21_X1   g04701(.A1(new_n4807_), .A2(new_n4893_), .B(new_n4888_), .ZN(new_n4894_));
  AOI21_X1   g04702(.A1(new_n4894_), .A2(new_n2531_), .B(new_n4805_), .ZN(new_n4895_));
  NAND2_X1   g04703(.A1(new_n4893_), .A2(new_n4807_), .ZN(new_n4896_));
  INV_X1     g04704(.I(new_n4888_), .ZN(new_n4897_));
  AOI21_X1   g04705(.A1(new_n4896_), .A2(new_n4897_), .B(new_n2531_), .ZN(new_n4898_));
  OAI21_X1   g04706(.A1(new_n4895_), .A2(new_n4898_), .B(\asqrt[45] ), .ZN(new_n4899_));
  NAND3_X1   g04707(.A1(new_n4892_), .A2(new_n2134_), .A3(new_n4899_), .ZN(new_n4900_));
  AOI21_X1   g04708(.A1(new_n4892_), .A2(new_n4899_), .B(new_n2134_), .ZN(new_n4901_));
  AOI21_X1   g04709(.A1(new_n4799_), .A2(new_n4900_), .B(new_n4901_), .ZN(new_n4902_));
  AOI21_X1   g04710(.A1(new_n4902_), .A2(new_n1953_), .B(new_n4796_), .ZN(new_n4903_));
  INV_X1     g04711(.I(new_n4801_), .ZN(new_n4904_));
  NOR3_X1    g04712(.A1(new_n4895_), .A2(\asqrt[45] ), .A3(new_n4898_), .ZN(new_n4905_));
  OAI21_X1   g04713(.A1(new_n4904_), .A2(new_n4905_), .B(new_n4899_), .ZN(new_n4906_));
  OAI21_X1   g04714(.A1(new_n4906_), .A2(\asqrt[46] ), .B(new_n4799_), .ZN(new_n4907_));
  NAND2_X1   g04715(.A1(new_n4906_), .A2(\asqrt[46] ), .ZN(new_n4908_));
  AOI21_X1   g04716(.A1(new_n4907_), .A2(new_n4908_), .B(new_n1953_), .ZN(new_n4909_));
  NOR3_X1    g04717(.A1(new_n4903_), .A2(\asqrt[48] ), .A3(new_n4909_), .ZN(new_n4910_));
  OAI21_X1   g04718(.A1(new_n4903_), .A2(new_n4909_), .B(\asqrt[48] ), .ZN(new_n4911_));
  OAI21_X1   g04719(.A1(new_n4793_), .A2(new_n4910_), .B(new_n4911_), .ZN(new_n4912_));
  OAI21_X1   g04720(.A1(new_n4912_), .A2(\asqrt[49] ), .B(new_n4789_), .ZN(new_n4913_));
  NAND3_X1   g04721(.A1(new_n4907_), .A2(new_n4908_), .A3(new_n1953_), .ZN(new_n4914_));
  AOI21_X1   g04722(.A1(new_n4795_), .A2(new_n4914_), .B(new_n4909_), .ZN(new_n4915_));
  AOI21_X1   g04723(.A1(new_n4915_), .A2(new_n1778_), .B(new_n4793_), .ZN(new_n4916_));
  NAND2_X1   g04724(.A1(new_n4914_), .A2(new_n4795_), .ZN(new_n4917_));
  INV_X1     g04725(.I(new_n4909_), .ZN(new_n4918_));
  AOI21_X1   g04726(.A1(new_n4917_), .A2(new_n4918_), .B(new_n1778_), .ZN(new_n4919_));
  OAI21_X1   g04727(.A1(new_n4916_), .A2(new_n4919_), .B(\asqrt[49] ), .ZN(new_n4920_));
  NAND3_X1   g04728(.A1(new_n4913_), .A2(new_n1463_), .A3(new_n4920_), .ZN(new_n4921_));
  AOI21_X1   g04729(.A1(new_n4913_), .A2(new_n4920_), .B(new_n1463_), .ZN(new_n4922_));
  AOI21_X1   g04730(.A1(new_n4787_), .A2(new_n4921_), .B(new_n4922_), .ZN(new_n4923_));
  AOI21_X1   g04731(.A1(new_n4923_), .A2(new_n1305_), .B(new_n4784_), .ZN(new_n4924_));
  INV_X1     g04732(.I(new_n4789_), .ZN(new_n4925_));
  NOR3_X1    g04733(.A1(new_n4916_), .A2(\asqrt[49] ), .A3(new_n4919_), .ZN(new_n4926_));
  OAI21_X1   g04734(.A1(new_n4925_), .A2(new_n4926_), .B(new_n4920_), .ZN(new_n4927_));
  OAI21_X1   g04735(.A1(new_n4927_), .A2(\asqrt[50] ), .B(new_n4787_), .ZN(new_n4928_));
  NAND2_X1   g04736(.A1(new_n4927_), .A2(\asqrt[50] ), .ZN(new_n4929_));
  AOI21_X1   g04737(.A1(new_n4928_), .A2(new_n4929_), .B(new_n1305_), .ZN(new_n4930_));
  NOR3_X1    g04738(.A1(new_n4924_), .A2(\asqrt[52] ), .A3(new_n4930_), .ZN(new_n4931_));
  OAI21_X1   g04739(.A1(new_n4924_), .A2(new_n4930_), .B(\asqrt[52] ), .ZN(new_n4932_));
  OAI21_X1   g04740(.A1(new_n4781_), .A2(new_n4931_), .B(new_n4932_), .ZN(new_n4933_));
  OAI21_X1   g04741(.A1(new_n4933_), .A2(\asqrt[53] ), .B(new_n4777_), .ZN(new_n4934_));
  NAND3_X1   g04742(.A1(new_n4928_), .A2(new_n4929_), .A3(new_n1305_), .ZN(new_n4935_));
  AOI21_X1   g04743(.A1(new_n4783_), .A2(new_n4935_), .B(new_n4930_), .ZN(new_n4936_));
  AOI21_X1   g04744(.A1(new_n4936_), .A2(new_n1150_), .B(new_n4781_), .ZN(new_n4937_));
  NAND2_X1   g04745(.A1(new_n4935_), .A2(new_n4783_), .ZN(new_n4938_));
  INV_X1     g04746(.I(new_n4930_), .ZN(new_n4939_));
  AOI21_X1   g04747(.A1(new_n4938_), .A2(new_n4939_), .B(new_n1150_), .ZN(new_n4940_));
  OAI21_X1   g04748(.A1(new_n4937_), .A2(new_n4940_), .B(\asqrt[53] ), .ZN(new_n4941_));
  NAND3_X1   g04749(.A1(new_n4934_), .A2(new_n860_), .A3(new_n4941_), .ZN(new_n4942_));
  AOI21_X1   g04750(.A1(new_n4934_), .A2(new_n4941_), .B(new_n860_), .ZN(new_n4943_));
  AOI21_X1   g04751(.A1(new_n4775_), .A2(new_n4942_), .B(new_n4943_), .ZN(new_n4944_));
  AOI21_X1   g04752(.A1(new_n4944_), .A2(new_n744_), .B(new_n4772_), .ZN(new_n4945_));
  INV_X1     g04753(.I(new_n4777_), .ZN(new_n4946_));
  NOR3_X1    g04754(.A1(new_n4937_), .A2(\asqrt[53] ), .A3(new_n4940_), .ZN(new_n4947_));
  OAI21_X1   g04755(.A1(new_n4946_), .A2(new_n4947_), .B(new_n4941_), .ZN(new_n4948_));
  OAI21_X1   g04756(.A1(new_n4948_), .A2(\asqrt[54] ), .B(new_n4775_), .ZN(new_n4949_));
  NAND2_X1   g04757(.A1(new_n4948_), .A2(\asqrt[54] ), .ZN(new_n4950_));
  AOI21_X1   g04758(.A1(new_n4949_), .A2(new_n4950_), .B(new_n744_), .ZN(new_n4951_));
  NOR3_X1    g04759(.A1(new_n4945_), .A2(\asqrt[56] ), .A3(new_n4951_), .ZN(new_n4952_));
  OAI21_X1   g04760(.A1(new_n4945_), .A2(new_n4951_), .B(\asqrt[56] ), .ZN(new_n4953_));
  OAI21_X1   g04761(.A1(new_n4769_), .A2(new_n4952_), .B(new_n4953_), .ZN(new_n4954_));
  OAI21_X1   g04762(.A1(new_n4954_), .A2(\asqrt[57] ), .B(new_n4765_), .ZN(new_n4955_));
  NAND3_X1   g04763(.A1(new_n4949_), .A2(new_n4950_), .A3(new_n744_), .ZN(new_n4956_));
  AOI21_X1   g04764(.A1(new_n4771_), .A2(new_n4956_), .B(new_n4951_), .ZN(new_n4957_));
  AOI21_X1   g04765(.A1(new_n4957_), .A2(new_n634_), .B(new_n4769_), .ZN(new_n4958_));
  NAND2_X1   g04766(.A1(new_n4956_), .A2(new_n4771_), .ZN(new_n4959_));
  INV_X1     g04767(.I(new_n4951_), .ZN(new_n4960_));
  AOI21_X1   g04768(.A1(new_n4959_), .A2(new_n4960_), .B(new_n634_), .ZN(new_n4961_));
  OAI21_X1   g04769(.A1(new_n4958_), .A2(new_n4961_), .B(\asqrt[57] ), .ZN(new_n4962_));
  NAND3_X1   g04770(.A1(new_n4955_), .A2(new_n423_), .A3(new_n4962_), .ZN(new_n4963_));
  AOI21_X1   g04771(.A1(new_n4955_), .A2(new_n4962_), .B(new_n423_), .ZN(new_n4964_));
  AOI21_X1   g04772(.A1(new_n4763_), .A2(new_n4963_), .B(new_n4964_), .ZN(new_n4965_));
  AOI21_X1   g04773(.A1(new_n4965_), .A2(new_n337_), .B(new_n4760_), .ZN(new_n4966_));
  NOR2_X1    g04774(.A1(new_n4965_), .A2(new_n337_), .ZN(new_n4967_));
  NOR3_X1    g04775(.A1(new_n4966_), .A2(new_n4967_), .A3(\asqrt[60] ), .ZN(new_n4968_));
  OAI21_X1   g04776(.A1(new_n4966_), .A2(new_n4967_), .B(\asqrt[60] ), .ZN(new_n4969_));
  OAI21_X1   g04777(.A1(new_n4757_), .A2(new_n4968_), .B(new_n4969_), .ZN(new_n4970_));
  NAND2_X1   g04778(.A1(new_n4970_), .A2(\asqrt[61] ), .ZN(new_n4971_));
  AOI21_X1   g04779(.A1(new_n4707_), .A2(new_n4713_), .B(\asqrt[35] ), .ZN(new_n4972_));
  XOR2_X1    g04780(.A1(new_n4972_), .A2(new_n4467_), .Z(new_n4973_));
  OAI21_X1   g04781(.A1(new_n4970_), .A2(\asqrt[61] ), .B(new_n4973_), .ZN(new_n4974_));
  NAND2_X1   g04782(.A1(new_n4974_), .A2(new_n4971_), .ZN(new_n4975_));
  INV_X1     g04783(.I(new_n4765_), .ZN(new_n4976_));
  NOR3_X1    g04784(.A1(new_n4958_), .A2(\asqrt[57] ), .A3(new_n4961_), .ZN(new_n4977_));
  OAI21_X1   g04785(.A1(new_n4976_), .A2(new_n4977_), .B(new_n4962_), .ZN(new_n4978_));
  OAI21_X1   g04786(.A1(new_n4978_), .A2(\asqrt[58] ), .B(new_n4763_), .ZN(new_n4979_));
  NOR2_X1    g04787(.A1(new_n4977_), .A2(new_n4976_), .ZN(new_n4980_));
  INV_X1     g04788(.I(new_n4962_), .ZN(new_n4981_));
  OAI21_X1   g04789(.A1(new_n4980_), .A2(new_n4981_), .B(\asqrt[58] ), .ZN(new_n4982_));
  NAND3_X1   g04790(.A1(new_n4979_), .A2(new_n337_), .A3(new_n4982_), .ZN(new_n4983_));
  NAND2_X1   g04791(.A1(new_n4983_), .A2(new_n4759_), .ZN(new_n4984_));
  INV_X1     g04792(.I(new_n4763_), .ZN(new_n4985_));
  NOR2_X1    g04793(.A1(new_n4980_), .A2(new_n4981_), .ZN(new_n4986_));
  AOI21_X1   g04794(.A1(new_n4986_), .A2(new_n423_), .B(new_n4985_), .ZN(new_n4987_));
  OAI21_X1   g04795(.A1(new_n4987_), .A2(new_n4964_), .B(\asqrt[59] ), .ZN(new_n4988_));
  NAND3_X1   g04796(.A1(new_n4984_), .A2(new_n266_), .A3(new_n4988_), .ZN(new_n4989_));
  NAND2_X1   g04797(.A1(new_n4989_), .A2(new_n4756_), .ZN(new_n4990_));
  AOI21_X1   g04798(.A1(new_n4990_), .A2(new_n4969_), .B(new_n239_), .ZN(new_n4991_));
  AOI21_X1   g04799(.A1(new_n4984_), .A2(new_n4988_), .B(new_n266_), .ZN(new_n4992_));
  AOI21_X1   g04800(.A1(new_n4756_), .A2(new_n4989_), .B(new_n4992_), .ZN(new_n4993_));
  INV_X1     g04801(.I(new_n4973_), .ZN(new_n4994_));
  AOI21_X1   g04802(.A1(new_n4993_), .A2(new_n239_), .B(new_n4994_), .ZN(new_n4995_));
  OAI21_X1   g04803(.A1(new_n4995_), .A2(new_n4991_), .B(new_n201_), .ZN(new_n4996_));
  NAND3_X1   g04804(.A1(new_n4974_), .A2(new_n4971_), .A3(\asqrt[62] ), .ZN(new_n4997_));
  NOR2_X1    g04805(.A1(new_n4705_), .A2(new_n4714_), .ZN(new_n4998_));
  NOR2_X1    g04806(.A1(\asqrt[35] ), .A2(new_n4998_), .ZN(new_n4999_));
  XOR2_X1    g04807(.A1(new_n4999_), .A2(new_n4703_), .Z(new_n5000_));
  INV_X1     g04808(.I(new_n5000_), .ZN(new_n5001_));
  AOI22_X1   g04809(.A1(new_n4997_), .A2(new_n4996_), .B1(new_n4975_), .B2(new_n5001_), .ZN(new_n5002_));
  NOR2_X1    g04810(.A1(new_n4725_), .A2(new_n4464_), .ZN(new_n5003_));
  OAI21_X1   g04811(.A1(\asqrt[35] ), .A2(new_n5003_), .B(new_n4732_), .ZN(new_n5004_));
  INV_X1     g04812(.I(new_n5004_), .ZN(new_n5005_));
  OAI21_X1   g04813(.A1(new_n5002_), .A2(new_n4754_), .B(new_n5005_), .ZN(new_n5006_));
  OAI21_X1   g04814(.A1(new_n4975_), .A2(\asqrt[62] ), .B(new_n5000_), .ZN(new_n5007_));
  NAND2_X1   g04815(.A1(new_n4975_), .A2(\asqrt[62] ), .ZN(new_n5008_));
  NAND3_X1   g04816(.A1(new_n5007_), .A2(new_n5008_), .A3(new_n4754_), .ZN(new_n5009_));
  NAND2_X1   g04817(.A1(new_n4725_), .A2(new_n4463_), .ZN(new_n5010_));
  NAND2_X1   g04818(.A1(new_n4747_), .A2(new_n4464_), .ZN(new_n5011_));
  AOI21_X1   g04819(.A1(new_n5010_), .A2(new_n5011_), .B(new_n193_), .ZN(new_n5012_));
  OAI21_X1   g04820(.A1(\asqrt[35] ), .A2(new_n4464_), .B(new_n5012_), .ZN(new_n5013_));
  NOR2_X1    g04821(.A1(new_n4738_), .A2(new_n4463_), .ZN(new_n5014_));
  NAND4_X1   g04822(.A1(new_n4729_), .A2(new_n193_), .A3(new_n4732_), .A4(new_n5014_), .ZN(new_n5015_));
  NAND2_X1   g04823(.A1(new_n5013_), .A2(new_n5015_), .ZN(new_n5016_));
  INV_X1     g04824(.I(new_n5016_), .ZN(new_n5017_));
  NAND4_X1   g04825(.A1(new_n5006_), .A2(new_n193_), .A3(new_n5009_), .A4(new_n5017_), .ZN(\asqrt[34] ));
  NOR2_X1    g04826(.A1(new_n4975_), .A2(\asqrt[62] ), .ZN(new_n5019_));
  NOR2_X1    g04827(.A1(new_n4995_), .A2(new_n4991_), .ZN(new_n5020_));
  NOR2_X1    g04828(.A1(new_n5020_), .A2(new_n201_), .ZN(new_n5021_));
  NOR2_X1    g04829(.A1(new_n5019_), .A2(new_n5021_), .ZN(new_n5022_));
  AOI21_X1   g04830(.A1(new_n4974_), .A2(new_n4971_), .B(\asqrt[62] ), .ZN(new_n5023_));
  NOR3_X1    g04831(.A1(new_n4995_), .A2(new_n201_), .A3(new_n4991_), .ZN(new_n5024_));
  OAI22_X1   g04832(.A1(new_n5023_), .A2(new_n5024_), .B1(new_n5020_), .B2(new_n5000_), .ZN(new_n5025_));
  AOI21_X1   g04833(.A1(new_n5025_), .A2(new_n4753_), .B(new_n5004_), .ZN(new_n5026_));
  AOI21_X1   g04834(.A1(new_n5020_), .A2(new_n201_), .B(new_n5001_), .ZN(new_n5027_));
  NOR3_X1    g04835(.A1(new_n5027_), .A2(new_n5021_), .A3(new_n4753_), .ZN(new_n5028_));
  NOR4_X1    g04836(.A1(new_n5026_), .A2(\asqrt[63] ), .A3(new_n5028_), .A4(new_n5016_), .ZN(new_n5029_));
  XOR2_X1    g04837(.A1(new_n4999_), .A2(new_n4703_), .Z(new_n5030_));
  OAI21_X1   g04838(.A1(\asqrt[34] ), .A2(new_n5022_), .B(new_n5030_), .ZN(new_n5031_));
  INV_X1     g04839(.I(new_n5031_), .ZN(new_n5032_));
  AOI21_X1   g04840(.A1(new_n4983_), .A2(new_n4988_), .B(\asqrt[34] ), .ZN(new_n5033_));
  XOR2_X1    g04841(.A1(new_n5033_), .A2(new_n4759_), .Z(new_n5034_));
  INV_X1     g04842(.I(new_n5034_), .ZN(new_n5035_));
  AOI21_X1   g04843(.A1(new_n4963_), .A2(new_n4982_), .B(\asqrt[34] ), .ZN(new_n5036_));
  XOR2_X1    g04844(.A1(new_n5036_), .A2(new_n4763_), .Z(new_n5037_));
  INV_X1     g04845(.I(new_n5037_), .ZN(new_n5038_));
  NOR2_X1    g04846(.A1(new_n4981_), .A2(new_n4977_), .ZN(new_n5039_));
  NOR2_X1    g04847(.A1(\asqrt[34] ), .A2(new_n5039_), .ZN(new_n5040_));
  XOR2_X1    g04848(.A1(new_n5040_), .A2(new_n4765_), .Z(new_n5041_));
  NOR2_X1    g04849(.A1(new_n4952_), .A2(new_n4961_), .ZN(new_n5042_));
  NOR2_X1    g04850(.A1(\asqrt[34] ), .A2(new_n5042_), .ZN(new_n5043_));
  XOR2_X1    g04851(.A1(new_n5043_), .A2(new_n4768_), .Z(new_n5044_));
  AOI21_X1   g04852(.A1(new_n4956_), .A2(new_n4960_), .B(\asqrt[34] ), .ZN(new_n5045_));
  XOR2_X1    g04853(.A1(new_n5045_), .A2(new_n4771_), .Z(new_n5046_));
  INV_X1     g04854(.I(new_n5046_), .ZN(new_n5047_));
  AOI21_X1   g04855(.A1(new_n4942_), .A2(new_n4950_), .B(\asqrt[34] ), .ZN(new_n5048_));
  XOR2_X1    g04856(.A1(new_n5048_), .A2(new_n4775_), .Z(new_n5049_));
  INV_X1     g04857(.I(new_n5049_), .ZN(new_n5050_));
  XOR2_X1    g04858(.A1(new_n4933_), .A2(\asqrt[53] ), .Z(new_n5051_));
  NOR2_X1    g04859(.A1(\asqrt[34] ), .A2(new_n5051_), .ZN(new_n5052_));
  XOR2_X1    g04860(.A1(new_n5052_), .A2(new_n4777_), .Z(new_n5053_));
  NOR2_X1    g04861(.A1(new_n4931_), .A2(new_n4940_), .ZN(new_n5054_));
  NOR2_X1    g04862(.A1(\asqrt[34] ), .A2(new_n5054_), .ZN(new_n5055_));
  XOR2_X1    g04863(.A1(new_n5055_), .A2(new_n4780_), .Z(new_n5056_));
  AOI21_X1   g04864(.A1(new_n4935_), .A2(new_n4939_), .B(\asqrt[34] ), .ZN(new_n5057_));
  XOR2_X1    g04865(.A1(new_n5057_), .A2(new_n4783_), .Z(new_n5058_));
  INV_X1     g04866(.I(new_n5058_), .ZN(new_n5059_));
  AOI21_X1   g04867(.A1(new_n4921_), .A2(new_n4929_), .B(\asqrt[34] ), .ZN(new_n5060_));
  XOR2_X1    g04868(.A1(new_n5060_), .A2(new_n4787_), .Z(new_n5061_));
  INV_X1     g04869(.I(new_n5061_), .ZN(new_n5062_));
  XOR2_X1    g04870(.A1(new_n4912_), .A2(\asqrt[49] ), .Z(new_n5063_));
  NOR2_X1    g04871(.A1(\asqrt[34] ), .A2(new_n5063_), .ZN(new_n5064_));
  XOR2_X1    g04872(.A1(new_n5064_), .A2(new_n4789_), .Z(new_n5065_));
  NOR2_X1    g04873(.A1(new_n4910_), .A2(new_n4919_), .ZN(new_n5066_));
  NOR2_X1    g04874(.A1(\asqrt[34] ), .A2(new_n5066_), .ZN(new_n5067_));
  XOR2_X1    g04875(.A1(new_n5067_), .A2(new_n4792_), .Z(new_n5068_));
  AOI21_X1   g04876(.A1(new_n4914_), .A2(new_n4918_), .B(\asqrt[34] ), .ZN(new_n5069_));
  XOR2_X1    g04877(.A1(new_n5069_), .A2(new_n4795_), .Z(new_n5070_));
  INV_X1     g04878(.I(new_n5070_), .ZN(new_n5071_));
  AOI21_X1   g04879(.A1(new_n4900_), .A2(new_n4908_), .B(\asqrt[34] ), .ZN(new_n5072_));
  XOR2_X1    g04880(.A1(new_n5072_), .A2(new_n4799_), .Z(new_n5073_));
  INV_X1     g04881(.I(new_n5073_), .ZN(new_n5074_));
  XOR2_X1    g04882(.A1(new_n4891_), .A2(\asqrt[45] ), .Z(new_n5075_));
  NOR2_X1    g04883(.A1(\asqrt[34] ), .A2(new_n5075_), .ZN(new_n5076_));
  XOR2_X1    g04884(.A1(new_n5076_), .A2(new_n4801_), .Z(new_n5077_));
  NOR2_X1    g04885(.A1(new_n4889_), .A2(new_n4898_), .ZN(new_n5078_));
  NOR2_X1    g04886(.A1(\asqrt[34] ), .A2(new_n5078_), .ZN(new_n5079_));
  XOR2_X1    g04887(.A1(new_n5079_), .A2(new_n4804_), .Z(new_n5080_));
  AOI21_X1   g04888(.A1(new_n4893_), .A2(new_n4897_), .B(\asqrt[34] ), .ZN(new_n5081_));
  XOR2_X1    g04889(.A1(new_n5081_), .A2(new_n4807_), .Z(new_n5082_));
  INV_X1     g04890(.I(new_n5082_), .ZN(new_n5083_));
  AOI21_X1   g04891(.A1(new_n4879_), .A2(new_n4887_), .B(\asqrt[34] ), .ZN(new_n5084_));
  XOR2_X1    g04892(.A1(new_n5084_), .A2(new_n4811_), .Z(new_n5085_));
  INV_X1     g04893(.I(new_n5085_), .ZN(new_n5086_));
  XOR2_X1    g04894(.A1(new_n4870_), .A2(\asqrt[41] ), .Z(new_n5087_));
  NOR2_X1    g04895(.A1(\asqrt[34] ), .A2(new_n5087_), .ZN(new_n5088_));
  XOR2_X1    g04896(.A1(new_n5088_), .A2(new_n4813_), .Z(new_n5089_));
  NOR2_X1    g04897(.A1(new_n4868_), .A2(new_n4877_), .ZN(new_n5090_));
  NOR2_X1    g04898(.A1(\asqrt[34] ), .A2(new_n5090_), .ZN(new_n5091_));
  XOR2_X1    g04899(.A1(new_n5091_), .A2(new_n4816_), .Z(new_n5092_));
  AOI21_X1   g04900(.A1(new_n4872_), .A2(new_n4876_), .B(\asqrt[34] ), .ZN(new_n5093_));
  XOR2_X1    g04901(.A1(new_n5093_), .A2(new_n4819_), .Z(new_n5094_));
  INV_X1     g04902(.I(new_n5094_), .ZN(new_n5095_));
  AOI21_X1   g04903(.A1(new_n4858_), .A2(new_n4866_), .B(\asqrt[34] ), .ZN(new_n5096_));
  XOR2_X1    g04904(.A1(new_n5096_), .A2(new_n4826_), .Z(new_n5097_));
  INV_X1     g04905(.I(new_n5097_), .ZN(new_n5098_));
  AOI21_X1   g04906(.A1(new_n4849_), .A2(new_n4857_), .B(\asqrt[34] ), .ZN(new_n5099_));
  XOR2_X1    g04907(.A1(new_n5099_), .A2(new_n4834_), .Z(new_n5100_));
  NAND2_X1   g04908(.A1(\asqrt[35] ), .A2(new_n4835_), .ZN(new_n5101_));
  NOR2_X1    g04909(.A1(new_n4846_), .A2(\a[70] ), .ZN(new_n5102_));
  AOI22_X1   g04910(.A1(new_n5101_), .A2(new_n4846_), .B1(\asqrt[35] ), .B2(new_n5102_), .ZN(new_n5103_));
  AOI21_X1   g04911(.A1(\asqrt[35] ), .A2(\a[70] ), .B(new_n4843_), .ZN(new_n5104_));
  OAI21_X1   g04912(.A1(new_n4853_), .A2(new_n5104_), .B(new_n5029_), .ZN(new_n5105_));
  XNOR2_X1   g04913(.A1(new_n5105_), .A2(new_n5103_), .ZN(new_n5106_));
  NOR3_X1    g04914(.A1(new_n5026_), .A2(\asqrt[63] ), .A3(new_n5028_), .ZN(new_n5107_));
  NAND4_X1   g04915(.A1(new_n5107_), .A2(\asqrt[35] ), .A3(new_n5013_), .A4(new_n5015_), .ZN(new_n5108_));
  NAND2_X1   g04916(.A1(\asqrt[34] ), .A2(new_n4836_), .ZN(new_n5109_));
  AOI21_X1   g04917(.A1(new_n5108_), .A2(new_n5109_), .B(\a[70] ), .ZN(new_n5110_));
  NAND2_X1   g04918(.A1(new_n5006_), .A2(new_n193_), .ZN(new_n5111_));
  NAND3_X1   g04919(.A1(new_n5013_), .A2(new_n5015_), .A3(\asqrt[35] ), .ZN(new_n5112_));
  NOR3_X1    g04920(.A1(new_n5111_), .A2(new_n5028_), .A3(new_n5112_), .ZN(new_n5113_));
  NOR2_X1    g04921(.A1(new_n5029_), .A2(new_n4838_), .ZN(new_n5114_));
  NOR3_X1    g04922(.A1(new_n5114_), .A2(new_n5113_), .A3(new_n4835_), .ZN(new_n5115_));
  OR2_X2     g04923(.A1(new_n5110_), .A2(new_n5115_), .Z(new_n5116_));
  NOR2_X1    g04924(.A1(\a[66] ), .A2(\a[67] ), .ZN(new_n5117_));
  INV_X1     g04925(.I(new_n5117_), .ZN(new_n5118_));
  NAND3_X1   g04926(.A1(\asqrt[34] ), .A2(\a[68] ), .A3(new_n5118_), .ZN(new_n5119_));
  INV_X1     g04927(.I(\a[68] ), .ZN(new_n5120_));
  OAI21_X1   g04928(.A1(\asqrt[34] ), .A2(new_n5120_), .B(new_n5117_), .ZN(new_n5121_));
  AOI21_X1   g04929(.A1(new_n5121_), .A2(new_n5119_), .B(new_n4751_), .ZN(new_n5122_));
  NOR3_X1    g04930(.A1(new_n4748_), .A2(\asqrt[63] ), .A3(new_n4750_), .ZN(new_n5123_));
  NAND2_X1   g04931(.A1(new_n5117_), .A2(new_n5120_), .ZN(new_n5124_));
  NAND3_X1   g04932(.A1(new_n4735_), .A2(new_n4737_), .A3(new_n5124_), .ZN(new_n5125_));
  NAND2_X1   g04933(.A1(new_n5123_), .A2(new_n5125_), .ZN(new_n5126_));
  NAND3_X1   g04934(.A1(\asqrt[34] ), .A2(\a[68] ), .A3(new_n5126_), .ZN(new_n5127_));
  INV_X1     g04935(.I(\a[69] ), .ZN(new_n5128_));
  NAND3_X1   g04936(.A1(\asqrt[34] ), .A2(new_n5120_), .A3(new_n5128_), .ZN(new_n5129_));
  OAI21_X1   g04937(.A1(new_n5029_), .A2(\a[68] ), .B(\a[69] ), .ZN(new_n5130_));
  NAND3_X1   g04938(.A1(new_n5127_), .A2(new_n5130_), .A3(new_n5129_), .ZN(new_n5131_));
  NOR3_X1    g04939(.A1(new_n5131_), .A2(new_n5122_), .A3(\asqrt[36] ), .ZN(new_n5132_));
  OAI21_X1   g04940(.A1(new_n5131_), .A2(new_n5122_), .B(\asqrt[36] ), .ZN(new_n5133_));
  OAI21_X1   g04941(.A1(new_n5116_), .A2(new_n5132_), .B(new_n5133_), .ZN(new_n5134_));
  OAI21_X1   g04942(.A1(new_n5134_), .A2(\asqrt[37] ), .B(new_n5106_), .ZN(new_n5135_));
  NAND2_X1   g04943(.A1(new_n5134_), .A2(\asqrt[37] ), .ZN(new_n5136_));
  NAND3_X1   g04944(.A1(new_n5135_), .A2(new_n5136_), .A3(new_n3925_), .ZN(new_n5137_));
  AOI21_X1   g04945(.A1(new_n5135_), .A2(new_n5136_), .B(new_n3925_), .ZN(new_n5138_));
  AOI21_X1   g04946(.A1(new_n5100_), .A2(new_n5137_), .B(new_n5138_), .ZN(new_n5139_));
  AOI21_X1   g04947(.A1(new_n5139_), .A2(new_n3681_), .B(new_n5098_), .ZN(new_n5140_));
  NAND2_X1   g04948(.A1(new_n5137_), .A2(new_n5100_), .ZN(new_n5141_));
  INV_X1     g04949(.I(new_n5106_), .ZN(new_n5142_));
  NOR2_X1    g04950(.A1(new_n5110_), .A2(new_n5115_), .ZN(new_n5143_));
  NOR3_X1    g04951(.A1(new_n5029_), .A2(new_n5120_), .A3(new_n5117_), .ZN(new_n5144_));
  AOI21_X1   g04952(.A1(new_n5029_), .A2(\a[68] ), .B(new_n5118_), .ZN(new_n5145_));
  OAI21_X1   g04953(.A1(new_n5144_), .A2(new_n5145_), .B(\asqrt[35] ), .ZN(new_n5146_));
  INV_X1     g04954(.I(new_n5126_), .ZN(new_n5147_));
  NOR3_X1    g04955(.A1(new_n5029_), .A2(new_n5120_), .A3(new_n5147_), .ZN(new_n5148_));
  NOR3_X1    g04956(.A1(new_n5029_), .A2(\a[68] ), .A3(\a[69] ), .ZN(new_n5149_));
  AOI21_X1   g04957(.A1(\asqrt[34] ), .A2(new_n5120_), .B(new_n5128_), .ZN(new_n5150_));
  NOR3_X1    g04958(.A1(new_n5148_), .A2(new_n5149_), .A3(new_n5150_), .ZN(new_n5151_));
  NAND3_X1   g04959(.A1(new_n5151_), .A2(new_n5146_), .A3(new_n4461_), .ZN(new_n5152_));
  AOI21_X1   g04960(.A1(new_n5151_), .A2(new_n5146_), .B(new_n4461_), .ZN(new_n5153_));
  AOI21_X1   g04961(.A1(new_n5143_), .A2(new_n5152_), .B(new_n5153_), .ZN(new_n5154_));
  AOI21_X1   g04962(.A1(new_n5154_), .A2(new_n4196_), .B(new_n5142_), .ZN(new_n5155_));
  NAND2_X1   g04963(.A1(new_n5152_), .A2(new_n5143_), .ZN(new_n5156_));
  AOI21_X1   g04964(.A1(new_n5156_), .A2(new_n5133_), .B(new_n4196_), .ZN(new_n5157_));
  OAI21_X1   g04965(.A1(new_n5155_), .A2(new_n5157_), .B(\asqrt[38] ), .ZN(new_n5158_));
  AOI21_X1   g04966(.A1(new_n5141_), .A2(new_n5158_), .B(new_n3681_), .ZN(new_n5159_));
  NOR3_X1    g04967(.A1(new_n5140_), .A2(\asqrt[40] ), .A3(new_n5159_), .ZN(new_n5160_));
  OAI21_X1   g04968(.A1(new_n5140_), .A2(new_n5159_), .B(\asqrt[40] ), .ZN(new_n5161_));
  OAI21_X1   g04969(.A1(new_n5095_), .A2(new_n5160_), .B(new_n5161_), .ZN(new_n5162_));
  OAI21_X1   g04970(.A1(new_n5162_), .A2(\asqrt[41] ), .B(new_n5092_), .ZN(new_n5163_));
  NAND2_X1   g04971(.A1(new_n5162_), .A2(\asqrt[41] ), .ZN(new_n5164_));
  NAND3_X1   g04972(.A1(new_n5163_), .A2(new_n5164_), .A3(new_n2960_), .ZN(new_n5165_));
  AOI21_X1   g04973(.A1(new_n5163_), .A2(new_n5164_), .B(new_n2960_), .ZN(new_n5166_));
  AOI21_X1   g04974(.A1(new_n5089_), .A2(new_n5165_), .B(new_n5166_), .ZN(new_n5167_));
  AOI21_X1   g04975(.A1(new_n5167_), .A2(new_n2749_), .B(new_n5086_), .ZN(new_n5168_));
  NAND2_X1   g04976(.A1(new_n5165_), .A2(new_n5089_), .ZN(new_n5169_));
  INV_X1     g04977(.I(new_n5092_), .ZN(new_n5170_));
  INV_X1     g04978(.I(new_n5100_), .ZN(new_n5171_));
  NOR3_X1    g04979(.A1(new_n5155_), .A2(\asqrt[38] ), .A3(new_n5157_), .ZN(new_n5172_));
  OAI21_X1   g04980(.A1(new_n5171_), .A2(new_n5172_), .B(new_n5158_), .ZN(new_n5173_));
  OAI21_X1   g04981(.A1(new_n5173_), .A2(\asqrt[39] ), .B(new_n5097_), .ZN(new_n5174_));
  NAND2_X1   g04982(.A1(new_n5173_), .A2(\asqrt[39] ), .ZN(new_n5175_));
  NAND3_X1   g04983(.A1(new_n5174_), .A2(new_n5175_), .A3(new_n3427_), .ZN(new_n5176_));
  AOI21_X1   g04984(.A1(new_n5174_), .A2(new_n5175_), .B(new_n3427_), .ZN(new_n5177_));
  AOI21_X1   g04985(.A1(new_n5094_), .A2(new_n5176_), .B(new_n5177_), .ZN(new_n5178_));
  AOI21_X1   g04986(.A1(new_n5178_), .A2(new_n3195_), .B(new_n5170_), .ZN(new_n5179_));
  NAND2_X1   g04987(.A1(new_n5176_), .A2(new_n5094_), .ZN(new_n5180_));
  AOI21_X1   g04988(.A1(new_n5180_), .A2(new_n5161_), .B(new_n3195_), .ZN(new_n5181_));
  OAI21_X1   g04989(.A1(new_n5179_), .A2(new_n5181_), .B(\asqrt[42] ), .ZN(new_n5182_));
  AOI21_X1   g04990(.A1(new_n5169_), .A2(new_n5182_), .B(new_n2749_), .ZN(new_n5183_));
  NOR3_X1    g04991(.A1(new_n5168_), .A2(\asqrt[44] ), .A3(new_n5183_), .ZN(new_n5184_));
  OAI21_X1   g04992(.A1(new_n5168_), .A2(new_n5183_), .B(\asqrt[44] ), .ZN(new_n5185_));
  OAI21_X1   g04993(.A1(new_n5083_), .A2(new_n5184_), .B(new_n5185_), .ZN(new_n5186_));
  OAI21_X1   g04994(.A1(new_n5186_), .A2(\asqrt[45] ), .B(new_n5080_), .ZN(new_n5187_));
  NAND2_X1   g04995(.A1(new_n5186_), .A2(\asqrt[45] ), .ZN(new_n5188_));
  NAND3_X1   g04996(.A1(new_n5187_), .A2(new_n5188_), .A3(new_n2134_), .ZN(new_n5189_));
  AOI21_X1   g04997(.A1(new_n5187_), .A2(new_n5188_), .B(new_n2134_), .ZN(new_n5190_));
  AOI21_X1   g04998(.A1(new_n5077_), .A2(new_n5189_), .B(new_n5190_), .ZN(new_n5191_));
  AOI21_X1   g04999(.A1(new_n5191_), .A2(new_n1953_), .B(new_n5074_), .ZN(new_n5192_));
  NAND2_X1   g05000(.A1(new_n5189_), .A2(new_n5077_), .ZN(new_n5193_));
  INV_X1     g05001(.I(new_n5080_), .ZN(new_n5194_));
  INV_X1     g05002(.I(new_n5089_), .ZN(new_n5195_));
  NOR3_X1    g05003(.A1(new_n5179_), .A2(\asqrt[42] ), .A3(new_n5181_), .ZN(new_n5196_));
  OAI21_X1   g05004(.A1(new_n5195_), .A2(new_n5196_), .B(new_n5182_), .ZN(new_n5197_));
  OAI21_X1   g05005(.A1(new_n5197_), .A2(\asqrt[43] ), .B(new_n5085_), .ZN(new_n5198_));
  NAND2_X1   g05006(.A1(new_n5197_), .A2(\asqrt[43] ), .ZN(new_n5199_));
  NAND3_X1   g05007(.A1(new_n5198_), .A2(new_n5199_), .A3(new_n2531_), .ZN(new_n5200_));
  AOI21_X1   g05008(.A1(new_n5198_), .A2(new_n5199_), .B(new_n2531_), .ZN(new_n5201_));
  AOI21_X1   g05009(.A1(new_n5082_), .A2(new_n5200_), .B(new_n5201_), .ZN(new_n5202_));
  AOI21_X1   g05010(.A1(new_n5202_), .A2(new_n2332_), .B(new_n5194_), .ZN(new_n5203_));
  NAND2_X1   g05011(.A1(new_n5200_), .A2(new_n5082_), .ZN(new_n5204_));
  AOI21_X1   g05012(.A1(new_n5204_), .A2(new_n5185_), .B(new_n2332_), .ZN(new_n5205_));
  OAI21_X1   g05013(.A1(new_n5203_), .A2(new_n5205_), .B(\asqrt[46] ), .ZN(new_n5206_));
  AOI21_X1   g05014(.A1(new_n5193_), .A2(new_n5206_), .B(new_n1953_), .ZN(new_n5207_));
  NOR3_X1    g05015(.A1(new_n5192_), .A2(\asqrt[48] ), .A3(new_n5207_), .ZN(new_n5208_));
  OAI21_X1   g05016(.A1(new_n5192_), .A2(new_n5207_), .B(\asqrt[48] ), .ZN(new_n5209_));
  OAI21_X1   g05017(.A1(new_n5071_), .A2(new_n5208_), .B(new_n5209_), .ZN(new_n5210_));
  OAI21_X1   g05018(.A1(new_n5210_), .A2(\asqrt[49] ), .B(new_n5068_), .ZN(new_n5211_));
  NAND2_X1   g05019(.A1(new_n5210_), .A2(\asqrt[49] ), .ZN(new_n5212_));
  NAND3_X1   g05020(.A1(new_n5211_), .A2(new_n5212_), .A3(new_n1463_), .ZN(new_n5213_));
  AOI21_X1   g05021(.A1(new_n5211_), .A2(new_n5212_), .B(new_n1463_), .ZN(new_n5214_));
  AOI21_X1   g05022(.A1(new_n5065_), .A2(new_n5213_), .B(new_n5214_), .ZN(new_n5215_));
  AOI21_X1   g05023(.A1(new_n5215_), .A2(new_n1305_), .B(new_n5062_), .ZN(new_n5216_));
  NAND2_X1   g05024(.A1(new_n5213_), .A2(new_n5065_), .ZN(new_n5217_));
  INV_X1     g05025(.I(new_n5068_), .ZN(new_n5218_));
  INV_X1     g05026(.I(new_n5077_), .ZN(new_n5219_));
  NOR3_X1    g05027(.A1(new_n5203_), .A2(\asqrt[46] ), .A3(new_n5205_), .ZN(new_n5220_));
  OAI21_X1   g05028(.A1(new_n5219_), .A2(new_n5220_), .B(new_n5206_), .ZN(new_n5221_));
  OAI21_X1   g05029(.A1(new_n5221_), .A2(\asqrt[47] ), .B(new_n5073_), .ZN(new_n5222_));
  NAND2_X1   g05030(.A1(new_n5221_), .A2(\asqrt[47] ), .ZN(new_n5223_));
  NAND3_X1   g05031(.A1(new_n5222_), .A2(new_n5223_), .A3(new_n1778_), .ZN(new_n5224_));
  AOI21_X1   g05032(.A1(new_n5222_), .A2(new_n5223_), .B(new_n1778_), .ZN(new_n5225_));
  AOI21_X1   g05033(.A1(new_n5070_), .A2(new_n5224_), .B(new_n5225_), .ZN(new_n5226_));
  AOI21_X1   g05034(.A1(new_n5226_), .A2(new_n1632_), .B(new_n5218_), .ZN(new_n5227_));
  NAND2_X1   g05035(.A1(new_n5224_), .A2(new_n5070_), .ZN(new_n5228_));
  AOI21_X1   g05036(.A1(new_n5228_), .A2(new_n5209_), .B(new_n1632_), .ZN(new_n5229_));
  OAI21_X1   g05037(.A1(new_n5227_), .A2(new_n5229_), .B(\asqrt[50] ), .ZN(new_n5230_));
  AOI21_X1   g05038(.A1(new_n5217_), .A2(new_n5230_), .B(new_n1305_), .ZN(new_n5231_));
  NOR3_X1    g05039(.A1(new_n5216_), .A2(\asqrt[52] ), .A3(new_n5231_), .ZN(new_n5232_));
  OAI21_X1   g05040(.A1(new_n5216_), .A2(new_n5231_), .B(\asqrt[52] ), .ZN(new_n5233_));
  OAI21_X1   g05041(.A1(new_n5059_), .A2(new_n5232_), .B(new_n5233_), .ZN(new_n5234_));
  OAI21_X1   g05042(.A1(new_n5234_), .A2(\asqrt[53] ), .B(new_n5056_), .ZN(new_n5235_));
  NAND2_X1   g05043(.A1(new_n5234_), .A2(\asqrt[53] ), .ZN(new_n5236_));
  NAND3_X1   g05044(.A1(new_n5235_), .A2(new_n5236_), .A3(new_n860_), .ZN(new_n5237_));
  AOI21_X1   g05045(.A1(new_n5235_), .A2(new_n5236_), .B(new_n860_), .ZN(new_n5238_));
  AOI21_X1   g05046(.A1(new_n5053_), .A2(new_n5237_), .B(new_n5238_), .ZN(new_n5239_));
  AOI21_X1   g05047(.A1(new_n5239_), .A2(new_n744_), .B(new_n5050_), .ZN(new_n5240_));
  NAND2_X1   g05048(.A1(new_n5237_), .A2(new_n5053_), .ZN(new_n5241_));
  INV_X1     g05049(.I(new_n5056_), .ZN(new_n5242_));
  INV_X1     g05050(.I(new_n5065_), .ZN(new_n5243_));
  NOR3_X1    g05051(.A1(new_n5227_), .A2(\asqrt[50] ), .A3(new_n5229_), .ZN(new_n5244_));
  OAI21_X1   g05052(.A1(new_n5243_), .A2(new_n5244_), .B(new_n5230_), .ZN(new_n5245_));
  OAI21_X1   g05053(.A1(new_n5245_), .A2(\asqrt[51] ), .B(new_n5061_), .ZN(new_n5246_));
  NAND2_X1   g05054(.A1(new_n5245_), .A2(\asqrt[51] ), .ZN(new_n5247_));
  NAND3_X1   g05055(.A1(new_n5246_), .A2(new_n5247_), .A3(new_n1150_), .ZN(new_n5248_));
  AOI21_X1   g05056(.A1(new_n5246_), .A2(new_n5247_), .B(new_n1150_), .ZN(new_n5249_));
  AOI21_X1   g05057(.A1(new_n5058_), .A2(new_n5248_), .B(new_n5249_), .ZN(new_n5250_));
  AOI21_X1   g05058(.A1(new_n5250_), .A2(new_n1006_), .B(new_n5242_), .ZN(new_n5251_));
  NAND2_X1   g05059(.A1(new_n5248_), .A2(new_n5058_), .ZN(new_n5252_));
  AOI21_X1   g05060(.A1(new_n5252_), .A2(new_n5233_), .B(new_n1006_), .ZN(new_n5253_));
  OAI21_X1   g05061(.A1(new_n5251_), .A2(new_n5253_), .B(\asqrt[54] ), .ZN(new_n5254_));
  AOI21_X1   g05062(.A1(new_n5241_), .A2(new_n5254_), .B(new_n744_), .ZN(new_n5255_));
  NOR3_X1    g05063(.A1(new_n5240_), .A2(\asqrt[56] ), .A3(new_n5255_), .ZN(new_n5256_));
  OAI21_X1   g05064(.A1(new_n5240_), .A2(new_n5255_), .B(\asqrt[56] ), .ZN(new_n5257_));
  OAI21_X1   g05065(.A1(new_n5047_), .A2(new_n5256_), .B(new_n5257_), .ZN(new_n5258_));
  OAI21_X1   g05066(.A1(new_n5258_), .A2(\asqrt[57] ), .B(new_n5044_), .ZN(new_n5259_));
  NAND2_X1   g05067(.A1(new_n5258_), .A2(\asqrt[57] ), .ZN(new_n5260_));
  NAND3_X1   g05068(.A1(new_n5259_), .A2(new_n5260_), .A3(new_n423_), .ZN(new_n5261_));
  AOI21_X1   g05069(.A1(new_n5259_), .A2(new_n5260_), .B(new_n423_), .ZN(new_n5262_));
  AOI21_X1   g05070(.A1(new_n5041_), .A2(new_n5261_), .B(new_n5262_), .ZN(new_n5263_));
  AOI21_X1   g05071(.A1(new_n5263_), .A2(new_n337_), .B(new_n5038_), .ZN(new_n5264_));
  NAND2_X1   g05072(.A1(new_n5261_), .A2(new_n5041_), .ZN(new_n5265_));
  INV_X1     g05073(.I(new_n5044_), .ZN(new_n5266_));
  INV_X1     g05074(.I(new_n5053_), .ZN(new_n5267_));
  NOR3_X1    g05075(.A1(new_n5251_), .A2(\asqrt[54] ), .A3(new_n5253_), .ZN(new_n5268_));
  OAI21_X1   g05076(.A1(new_n5267_), .A2(new_n5268_), .B(new_n5254_), .ZN(new_n5269_));
  OAI21_X1   g05077(.A1(new_n5269_), .A2(\asqrt[55] ), .B(new_n5049_), .ZN(new_n5270_));
  NAND2_X1   g05078(.A1(new_n5269_), .A2(\asqrt[55] ), .ZN(new_n5271_));
  NAND3_X1   g05079(.A1(new_n5270_), .A2(new_n5271_), .A3(new_n634_), .ZN(new_n5272_));
  AOI21_X1   g05080(.A1(new_n5270_), .A2(new_n5271_), .B(new_n634_), .ZN(new_n5273_));
  AOI21_X1   g05081(.A1(new_n5046_), .A2(new_n5272_), .B(new_n5273_), .ZN(new_n5274_));
  AOI21_X1   g05082(.A1(new_n5274_), .A2(new_n531_), .B(new_n5266_), .ZN(new_n5275_));
  NAND2_X1   g05083(.A1(new_n5272_), .A2(new_n5046_), .ZN(new_n5276_));
  AOI21_X1   g05084(.A1(new_n5276_), .A2(new_n5257_), .B(new_n531_), .ZN(new_n5277_));
  OAI21_X1   g05085(.A1(new_n5275_), .A2(new_n5277_), .B(\asqrt[58] ), .ZN(new_n5278_));
  AOI21_X1   g05086(.A1(new_n5265_), .A2(new_n5278_), .B(new_n337_), .ZN(new_n5279_));
  NOR3_X1    g05087(.A1(new_n5264_), .A2(\asqrt[60] ), .A3(new_n5279_), .ZN(new_n5280_));
  NOR2_X1    g05088(.A1(new_n5280_), .A2(new_n5035_), .ZN(new_n5281_));
  INV_X1     g05089(.I(new_n5041_), .ZN(new_n5282_));
  NOR3_X1    g05090(.A1(new_n5275_), .A2(\asqrt[58] ), .A3(new_n5277_), .ZN(new_n5283_));
  OAI21_X1   g05091(.A1(new_n5282_), .A2(new_n5283_), .B(new_n5278_), .ZN(new_n5284_));
  OAI21_X1   g05092(.A1(new_n5284_), .A2(\asqrt[59] ), .B(new_n5037_), .ZN(new_n5285_));
  NOR2_X1    g05093(.A1(new_n5283_), .A2(new_n5282_), .ZN(new_n5286_));
  OAI21_X1   g05094(.A1(new_n5286_), .A2(new_n5262_), .B(\asqrt[59] ), .ZN(new_n5287_));
  AOI21_X1   g05095(.A1(new_n5285_), .A2(new_n5287_), .B(new_n266_), .ZN(new_n5288_));
  OAI21_X1   g05096(.A1(new_n5281_), .A2(new_n5288_), .B(\asqrt[61] ), .ZN(new_n5289_));
  OAI21_X1   g05097(.A1(new_n5264_), .A2(new_n5279_), .B(\asqrt[60] ), .ZN(new_n5290_));
  OAI21_X1   g05098(.A1(new_n5035_), .A2(new_n5280_), .B(new_n5290_), .ZN(new_n5291_));
  AOI21_X1   g05099(.A1(new_n4989_), .A2(new_n4969_), .B(\asqrt[34] ), .ZN(new_n5292_));
  XOR2_X1    g05100(.A1(new_n5292_), .A2(new_n4756_), .Z(new_n5293_));
  OAI21_X1   g05101(.A1(new_n5291_), .A2(\asqrt[61] ), .B(new_n5293_), .ZN(new_n5294_));
  NAND2_X1   g05102(.A1(new_n5294_), .A2(new_n5289_), .ZN(new_n5295_));
  NAND3_X1   g05103(.A1(new_n5285_), .A2(new_n266_), .A3(new_n5287_), .ZN(new_n5296_));
  NAND2_X1   g05104(.A1(new_n5296_), .A2(new_n5034_), .ZN(new_n5297_));
  AOI21_X1   g05105(.A1(new_n5297_), .A2(new_n5290_), .B(new_n239_), .ZN(new_n5298_));
  AOI21_X1   g05106(.A1(new_n5034_), .A2(new_n5296_), .B(new_n5288_), .ZN(new_n5299_));
  INV_X1     g05107(.I(new_n5293_), .ZN(new_n5300_));
  AOI21_X1   g05108(.A1(new_n5299_), .A2(new_n239_), .B(new_n5300_), .ZN(new_n5301_));
  OAI21_X1   g05109(.A1(new_n5301_), .A2(new_n5298_), .B(new_n201_), .ZN(new_n5302_));
  NAND3_X1   g05110(.A1(new_n5294_), .A2(\asqrt[62] ), .A3(new_n5289_), .ZN(new_n5303_));
  NAND2_X1   g05111(.A1(new_n4993_), .A2(new_n239_), .ZN(new_n5304_));
  AOI21_X1   g05112(.A1(new_n4971_), .A2(new_n5304_), .B(\asqrt[34] ), .ZN(new_n5305_));
  XOR2_X1    g05113(.A1(new_n5305_), .A2(new_n4973_), .Z(new_n5306_));
  INV_X1     g05114(.I(new_n5306_), .ZN(new_n5307_));
  AOI22_X1   g05115(.A1(new_n5302_), .A2(new_n5303_), .B1(new_n5295_), .B2(new_n5307_), .ZN(new_n5308_));
  NOR2_X1    g05116(.A1(new_n5002_), .A2(new_n4754_), .ZN(new_n5309_));
  OAI21_X1   g05117(.A1(\asqrt[34] ), .A2(new_n5309_), .B(new_n5009_), .ZN(new_n5310_));
  INV_X1     g05118(.I(new_n5310_), .ZN(new_n5311_));
  OAI21_X1   g05119(.A1(new_n5308_), .A2(new_n5032_), .B(new_n5311_), .ZN(new_n5312_));
  OAI21_X1   g05120(.A1(new_n5295_), .A2(\asqrt[62] ), .B(new_n5306_), .ZN(new_n5313_));
  NAND2_X1   g05121(.A1(new_n5295_), .A2(\asqrt[62] ), .ZN(new_n5314_));
  NAND3_X1   g05122(.A1(new_n5313_), .A2(new_n5314_), .A3(new_n5032_), .ZN(new_n5315_));
  NAND2_X1   g05123(.A1(new_n5029_), .A2(new_n4753_), .ZN(new_n5316_));
  XOR2_X1    g05124(.A1(new_n5025_), .A2(new_n4753_), .Z(new_n5317_));
  NAND3_X1   g05125(.A1(new_n5316_), .A2(\asqrt[63] ), .A3(new_n5317_), .ZN(new_n5318_));
  INV_X1     g05126(.I(new_n5111_), .ZN(new_n5319_));
  NAND4_X1   g05127(.A1(new_n5319_), .A2(new_n4754_), .A3(new_n5009_), .A4(new_n5017_), .ZN(new_n5320_));
  NAND2_X1   g05128(.A1(new_n5318_), .A2(new_n5320_), .ZN(new_n5321_));
  INV_X1     g05129(.I(new_n5321_), .ZN(new_n5322_));
  NAND4_X1   g05130(.A1(new_n5312_), .A2(new_n193_), .A3(new_n5315_), .A4(new_n5322_), .ZN(\asqrt[33] ));
  NOR2_X1    g05131(.A1(new_n5295_), .A2(\asqrt[62] ), .ZN(new_n5324_));
  INV_X1     g05132(.I(new_n5314_), .ZN(new_n5325_));
  NOR2_X1    g05133(.A1(new_n5325_), .A2(new_n5324_), .ZN(new_n5326_));
  NAND3_X1   g05134(.A1(new_n5297_), .A2(new_n239_), .A3(new_n5290_), .ZN(new_n5327_));
  AOI21_X1   g05135(.A1(new_n5293_), .A2(new_n5327_), .B(new_n5298_), .ZN(new_n5328_));
  AOI21_X1   g05136(.A1(new_n5294_), .A2(new_n5289_), .B(\asqrt[62] ), .ZN(new_n5329_));
  NOR3_X1    g05137(.A1(new_n5301_), .A2(new_n201_), .A3(new_n5298_), .ZN(new_n5330_));
  OAI22_X1   g05138(.A1(new_n5330_), .A2(new_n5329_), .B1(new_n5328_), .B2(new_n5306_), .ZN(new_n5331_));
  AOI21_X1   g05139(.A1(new_n5331_), .A2(new_n5031_), .B(new_n5310_), .ZN(new_n5332_));
  AOI21_X1   g05140(.A1(new_n5328_), .A2(new_n201_), .B(new_n5307_), .ZN(new_n5333_));
  OAI21_X1   g05141(.A1(new_n5328_), .A2(new_n201_), .B(new_n5032_), .ZN(new_n5334_));
  NOR2_X1    g05142(.A1(new_n5333_), .A2(new_n5334_), .ZN(new_n5335_));
  NOR4_X1    g05143(.A1(new_n5332_), .A2(\asqrt[63] ), .A3(new_n5335_), .A4(new_n5321_), .ZN(new_n5336_));
  XOR2_X1    g05144(.A1(new_n5305_), .A2(new_n4973_), .Z(new_n5337_));
  OAI21_X1   g05145(.A1(\asqrt[33] ), .A2(new_n5326_), .B(new_n5337_), .ZN(new_n5338_));
  INV_X1     g05146(.I(new_n5338_), .ZN(new_n5339_));
  NAND2_X1   g05147(.A1(new_n5263_), .A2(new_n337_), .ZN(new_n5340_));
  AOI21_X1   g05148(.A1(new_n5340_), .A2(new_n5287_), .B(\asqrt[33] ), .ZN(new_n5341_));
  XOR2_X1    g05149(.A1(new_n5341_), .A2(new_n5037_), .Z(new_n5342_));
  INV_X1     g05150(.I(new_n5342_), .ZN(new_n5343_));
  AOI21_X1   g05151(.A1(new_n5261_), .A2(new_n5278_), .B(\asqrt[33] ), .ZN(new_n5344_));
  XOR2_X1    g05152(.A1(new_n5344_), .A2(new_n5041_), .Z(new_n5345_));
  INV_X1     g05153(.I(new_n5345_), .ZN(new_n5346_));
  NAND2_X1   g05154(.A1(new_n5274_), .A2(new_n531_), .ZN(new_n5347_));
  AOI21_X1   g05155(.A1(new_n5347_), .A2(new_n5260_), .B(\asqrt[33] ), .ZN(new_n5348_));
  XOR2_X1    g05156(.A1(new_n5348_), .A2(new_n5044_), .Z(new_n5349_));
  INV_X1     g05157(.I(new_n5349_), .ZN(new_n5350_));
  AOI21_X1   g05158(.A1(new_n5272_), .A2(new_n5257_), .B(\asqrt[33] ), .ZN(new_n5351_));
  XOR2_X1    g05159(.A1(new_n5351_), .A2(new_n5046_), .Z(new_n5352_));
  NAND2_X1   g05160(.A1(new_n5239_), .A2(new_n744_), .ZN(new_n5353_));
  AOI21_X1   g05161(.A1(new_n5353_), .A2(new_n5271_), .B(\asqrt[33] ), .ZN(new_n5354_));
  XOR2_X1    g05162(.A1(new_n5354_), .A2(new_n5049_), .Z(new_n5355_));
  AOI21_X1   g05163(.A1(new_n5237_), .A2(new_n5254_), .B(\asqrt[33] ), .ZN(new_n5356_));
  XOR2_X1    g05164(.A1(new_n5356_), .A2(new_n5053_), .Z(new_n5357_));
  INV_X1     g05165(.I(new_n5357_), .ZN(new_n5358_));
  NAND2_X1   g05166(.A1(new_n5250_), .A2(new_n1006_), .ZN(new_n5359_));
  AOI21_X1   g05167(.A1(new_n5359_), .A2(new_n5236_), .B(\asqrt[33] ), .ZN(new_n5360_));
  XOR2_X1    g05168(.A1(new_n5360_), .A2(new_n5056_), .Z(new_n5361_));
  INV_X1     g05169(.I(new_n5361_), .ZN(new_n5362_));
  AOI21_X1   g05170(.A1(new_n5248_), .A2(new_n5233_), .B(\asqrt[33] ), .ZN(new_n5363_));
  XOR2_X1    g05171(.A1(new_n5363_), .A2(new_n5058_), .Z(new_n5364_));
  NAND2_X1   g05172(.A1(new_n5215_), .A2(new_n1305_), .ZN(new_n5365_));
  AOI21_X1   g05173(.A1(new_n5365_), .A2(new_n5247_), .B(\asqrt[33] ), .ZN(new_n5366_));
  XOR2_X1    g05174(.A1(new_n5366_), .A2(new_n5061_), .Z(new_n5367_));
  AOI21_X1   g05175(.A1(new_n5213_), .A2(new_n5230_), .B(\asqrt[33] ), .ZN(new_n5368_));
  XOR2_X1    g05176(.A1(new_n5368_), .A2(new_n5065_), .Z(new_n5369_));
  INV_X1     g05177(.I(new_n5369_), .ZN(new_n5370_));
  NAND2_X1   g05178(.A1(new_n5226_), .A2(new_n1632_), .ZN(new_n5371_));
  AOI21_X1   g05179(.A1(new_n5371_), .A2(new_n5212_), .B(\asqrt[33] ), .ZN(new_n5372_));
  XOR2_X1    g05180(.A1(new_n5372_), .A2(new_n5068_), .Z(new_n5373_));
  INV_X1     g05181(.I(new_n5373_), .ZN(new_n5374_));
  AOI21_X1   g05182(.A1(new_n5224_), .A2(new_n5209_), .B(\asqrt[33] ), .ZN(new_n5375_));
  XOR2_X1    g05183(.A1(new_n5375_), .A2(new_n5070_), .Z(new_n5376_));
  NAND2_X1   g05184(.A1(new_n5191_), .A2(new_n1953_), .ZN(new_n5377_));
  AOI21_X1   g05185(.A1(new_n5377_), .A2(new_n5223_), .B(\asqrt[33] ), .ZN(new_n5378_));
  XOR2_X1    g05186(.A1(new_n5378_), .A2(new_n5073_), .Z(new_n5379_));
  AOI21_X1   g05187(.A1(new_n5189_), .A2(new_n5206_), .B(\asqrt[33] ), .ZN(new_n5380_));
  XOR2_X1    g05188(.A1(new_n5380_), .A2(new_n5077_), .Z(new_n5381_));
  INV_X1     g05189(.I(new_n5381_), .ZN(new_n5382_));
  NAND2_X1   g05190(.A1(new_n5202_), .A2(new_n2332_), .ZN(new_n5383_));
  AOI21_X1   g05191(.A1(new_n5383_), .A2(new_n5188_), .B(\asqrt[33] ), .ZN(new_n5384_));
  XOR2_X1    g05192(.A1(new_n5384_), .A2(new_n5080_), .Z(new_n5385_));
  INV_X1     g05193(.I(new_n5385_), .ZN(new_n5386_));
  AOI21_X1   g05194(.A1(new_n5200_), .A2(new_n5185_), .B(\asqrt[33] ), .ZN(new_n5387_));
  XOR2_X1    g05195(.A1(new_n5387_), .A2(new_n5082_), .Z(new_n5388_));
  NAND2_X1   g05196(.A1(new_n5167_), .A2(new_n2749_), .ZN(new_n5389_));
  AOI21_X1   g05197(.A1(new_n5389_), .A2(new_n5199_), .B(\asqrt[33] ), .ZN(new_n5390_));
  XOR2_X1    g05198(.A1(new_n5390_), .A2(new_n5085_), .Z(new_n5391_));
  AOI21_X1   g05199(.A1(new_n5165_), .A2(new_n5182_), .B(\asqrt[33] ), .ZN(new_n5392_));
  XOR2_X1    g05200(.A1(new_n5392_), .A2(new_n5089_), .Z(new_n5393_));
  INV_X1     g05201(.I(new_n5393_), .ZN(new_n5394_));
  NAND2_X1   g05202(.A1(new_n5178_), .A2(new_n3195_), .ZN(new_n5395_));
  AOI21_X1   g05203(.A1(new_n5395_), .A2(new_n5164_), .B(\asqrt[33] ), .ZN(new_n5396_));
  XOR2_X1    g05204(.A1(new_n5396_), .A2(new_n5092_), .Z(new_n5397_));
  INV_X1     g05205(.I(new_n5397_), .ZN(new_n5398_));
  AOI21_X1   g05206(.A1(new_n5176_), .A2(new_n5161_), .B(\asqrt[33] ), .ZN(new_n5399_));
  XOR2_X1    g05207(.A1(new_n5399_), .A2(new_n5094_), .Z(new_n5400_));
  NAND2_X1   g05208(.A1(new_n5139_), .A2(new_n3681_), .ZN(new_n5401_));
  AOI21_X1   g05209(.A1(new_n5401_), .A2(new_n5175_), .B(\asqrt[33] ), .ZN(new_n5402_));
  XOR2_X1    g05210(.A1(new_n5402_), .A2(new_n5097_), .Z(new_n5403_));
  AOI21_X1   g05211(.A1(new_n5137_), .A2(new_n5158_), .B(\asqrt[33] ), .ZN(new_n5404_));
  XOR2_X1    g05212(.A1(new_n5404_), .A2(new_n5100_), .Z(new_n5405_));
  INV_X1     g05213(.I(new_n5405_), .ZN(new_n5406_));
  NAND2_X1   g05214(.A1(new_n5154_), .A2(new_n4196_), .ZN(new_n5407_));
  AOI21_X1   g05215(.A1(new_n5407_), .A2(new_n5136_), .B(\asqrt[33] ), .ZN(new_n5408_));
  XOR2_X1    g05216(.A1(new_n5408_), .A2(new_n5106_), .Z(new_n5409_));
  INV_X1     g05217(.I(new_n5409_), .ZN(new_n5410_));
  AOI21_X1   g05218(.A1(new_n5152_), .A2(new_n5133_), .B(\asqrt[33] ), .ZN(new_n5411_));
  XOR2_X1    g05219(.A1(new_n5411_), .A2(new_n5143_), .Z(new_n5412_));
  NAND2_X1   g05220(.A1(\asqrt[34] ), .A2(new_n5120_), .ZN(new_n5413_));
  NOR2_X1    g05221(.A1(new_n5128_), .A2(\a[68] ), .ZN(new_n5414_));
  AOI22_X1   g05222(.A1(new_n5413_), .A2(new_n5128_), .B1(\asqrt[34] ), .B2(new_n5414_), .ZN(new_n5415_));
  OAI21_X1   g05223(.A1(new_n5029_), .A2(new_n5120_), .B(new_n5147_), .ZN(new_n5416_));
  AOI21_X1   g05224(.A1(new_n5146_), .A2(new_n5416_), .B(\asqrt[33] ), .ZN(new_n5417_));
  XOR2_X1    g05225(.A1(new_n5417_), .A2(new_n5415_), .Z(new_n5418_));
  NOR3_X1    g05226(.A1(new_n5332_), .A2(\asqrt[63] ), .A3(new_n5335_), .ZN(new_n5419_));
  NAND3_X1   g05227(.A1(new_n5318_), .A2(\asqrt[34] ), .A3(new_n5320_), .ZN(new_n5420_));
  INV_X1     g05228(.I(new_n5420_), .ZN(new_n5421_));
  NAND2_X1   g05229(.A1(new_n5419_), .A2(new_n5421_), .ZN(new_n5422_));
  NAND2_X1   g05230(.A1(\asqrt[33] ), .A2(new_n5117_), .ZN(new_n5423_));
  AOI21_X1   g05231(.A1(new_n5423_), .A2(new_n5422_), .B(\a[68] ), .ZN(new_n5424_));
  NAND2_X1   g05232(.A1(new_n5312_), .A2(new_n193_), .ZN(new_n5425_));
  NOR3_X1    g05233(.A1(new_n5425_), .A2(new_n5335_), .A3(new_n5420_), .ZN(new_n5426_));
  NOR2_X1    g05234(.A1(new_n5336_), .A2(new_n5118_), .ZN(new_n5427_));
  NOR3_X1    g05235(.A1(new_n5427_), .A2(new_n5426_), .A3(new_n5120_), .ZN(new_n5428_));
  OR2_X2     g05236(.A1(new_n5428_), .A2(new_n5424_), .Z(new_n5429_));
  NOR2_X1    g05237(.A1(\a[64] ), .A2(\a[65] ), .ZN(new_n5430_));
  INV_X1     g05238(.I(new_n5430_), .ZN(new_n5431_));
  NAND3_X1   g05239(.A1(\asqrt[33] ), .A2(\a[66] ), .A3(new_n5431_), .ZN(new_n5432_));
  INV_X1     g05240(.I(\a[66] ), .ZN(new_n5433_));
  OAI21_X1   g05241(.A1(\asqrt[33] ), .A2(new_n5433_), .B(new_n5430_), .ZN(new_n5434_));
  AOI21_X1   g05242(.A1(new_n5434_), .A2(new_n5432_), .B(new_n5029_), .ZN(new_n5435_));
  NAND2_X1   g05243(.A1(new_n5430_), .A2(new_n5433_), .ZN(new_n5436_));
  NAND3_X1   g05244(.A1(new_n5013_), .A2(new_n5015_), .A3(new_n5436_), .ZN(new_n5437_));
  NAND2_X1   g05245(.A1(new_n5107_), .A2(new_n5437_), .ZN(new_n5438_));
  NAND3_X1   g05246(.A1(\asqrt[33] ), .A2(\a[66] ), .A3(new_n5438_), .ZN(new_n5439_));
  INV_X1     g05247(.I(\a[67] ), .ZN(new_n5440_));
  NAND3_X1   g05248(.A1(\asqrt[33] ), .A2(new_n5433_), .A3(new_n5440_), .ZN(new_n5441_));
  OAI21_X1   g05249(.A1(new_n5336_), .A2(\a[66] ), .B(\a[67] ), .ZN(new_n5442_));
  NAND3_X1   g05250(.A1(new_n5439_), .A2(new_n5442_), .A3(new_n5441_), .ZN(new_n5443_));
  NOR3_X1    g05251(.A1(new_n5443_), .A2(new_n5435_), .A3(\asqrt[35] ), .ZN(new_n5444_));
  OAI21_X1   g05252(.A1(new_n5443_), .A2(new_n5435_), .B(\asqrt[35] ), .ZN(new_n5445_));
  OAI21_X1   g05253(.A1(new_n5429_), .A2(new_n5444_), .B(new_n5445_), .ZN(new_n5446_));
  OAI21_X1   g05254(.A1(new_n5446_), .A2(\asqrt[36] ), .B(new_n5418_), .ZN(new_n5447_));
  NAND2_X1   g05255(.A1(new_n5446_), .A2(\asqrt[36] ), .ZN(new_n5448_));
  NAND3_X1   g05256(.A1(new_n5447_), .A2(new_n5448_), .A3(new_n4196_), .ZN(new_n5449_));
  AOI21_X1   g05257(.A1(new_n5447_), .A2(new_n5448_), .B(new_n4196_), .ZN(new_n5450_));
  AOI21_X1   g05258(.A1(new_n5412_), .A2(new_n5449_), .B(new_n5450_), .ZN(new_n5451_));
  AOI21_X1   g05259(.A1(new_n5451_), .A2(new_n3925_), .B(new_n5410_), .ZN(new_n5452_));
  NAND2_X1   g05260(.A1(new_n5449_), .A2(new_n5412_), .ZN(new_n5453_));
  INV_X1     g05261(.I(new_n5450_), .ZN(new_n5454_));
  AOI21_X1   g05262(.A1(new_n5453_), .A2(new_n5454_), .B(new_n3925_), .ZN(new_n5455_));
  NOR3_X1    g05263(.A1(new_n5452_), .A2(\asqrt[39] ), .A3(new_n5455_), .ZN(new_n5456_));
  OAI21_X1   g05264(.A1(new_n5452_), .A2(new_n5455_), .B(\asqrt[39] ), .ZN(new_n5457_));
  OAI21_X1   g05265(.A1(new_n5406_), .A2(new_n5456_), .B(new_n5457_), .ZN(new_n5458_));
  OAI21_X1   g05266(.A1(new_n5458_), .A2(\asqrt[40] ), .B(new_n5403_), .ZN(new_n5459_));
  NAND2_X1   g05267(.A1(new_n5458_), .A2(\asqrt[40] ), .ZN(new_n5460_));
  NAND3_X1   g05268(.A1(new_n5459_), .A2(new_n5460_), .A3(new_n3195_), .ZN(new_n5461_));
  AOI21_X1   g05269(.A1(new_n5459_), .A2(new_n5460_), .B(new_n3195_), .ZN(new_n5462_));
  AOI21_X1   g05270(.A1(new_n5400_), .A2(new_n5461_), .B(new_n5462_), .ZN(new_n5463_));
  AOI21_X1   g05271(.A1(new_n5463_), .A2(new_n2960_), .B(new_n5398_), .ZN(new_n5464_));
  NAND2_X1   g05272(.A1(new_n5461_), .A2(new_n5400_), .ZN(new_n5465_));
  INV_X1     g05273(.I(new_n5462_), .ZN(new_n5466_));
  AOI21_X1   g05274(.A1(new_n5465_), .A2(new_n5466_), .B(new_n2960_), .ZN(new_n5467_));
  NOR3_X1    g05275(.A1(new_n5464_), .A2(\asqrt[43] ), .A3(new_n5467_), .ZN(new_n5468_));
  OAI21_X1   g05276(.A1(new_n5464_), .A2(new_n5467_), .B(\asqrt[43] ), .ZN(new_n5469_));
  OAI21_X1   g05277(.A1(new_n5394_), .A2(new_n5468_), .B(new_n5469_), .ZN(new_n5470_));
  OAI21_X1   g05278(.A1(new_n5470_), .A2(\asqrt[44] ), .B(new_n5391_), .ZN(new_n5471_));
  NAND2_X1   g05279(.A1(new_n5470_), .A2(\asqrt[44] ), .ZN(new_n5472_));
  NAND3_X1   g05280(.A1(new_n5471_), .A2(new_n5472_), .A3(new_n2332_), .ZN(new_n5473_));
  AOI21_X1   g05281(.A1(new_n5471_), .A2(new_n5472_), .B(new_n2332_), .ZN(new_n5474_));
  AOI21_X1   g05282(.A1(new_n5388_), .A2(new_n5473_), .B(new_n5474_), .ZN(new_n5475_));
  AOI21_X1   g05283(.A1(new_n5475_), .A2(new_n2134_), .B(new_n5386_), .ZN(new_n5476_));
  NAND2_X1   g05284(.A1(new_n5473_), .A2(new_n5388_), .ZN(new_n5477_));
  INV_X1     g05285(.I(new_n5474_), .ZN(new_n5478_));
  AOI21_X1   g05286(.A1(new_n5477_), .A2(new_n5478_), .B(new_n2134_), .ZN(new_n5479_));
  NOR3_X1    g05287(.A1(new_n5476_), .A2(\asqrt[47] ), .A3(new_n5479_), .ZN(new_n5480_));
  OAI21_X1   g05288(.A1(new_n5476_), .A2(new_n5479_), .B(\asqrt[47] ), .ZN(new_n5481_));
  OAI21_X1   g05289(.A1(new_n5382_), .A2(new_n5480_), .B(new_n5481_), .ZN(new_n5482_));
  OAI21_X1   g05290(.A1(new_n5482_), .A2(\asqrt[48] ), .B(new_n5379_), .ZN(new_n5483_));
  NAND2_X1   g05291(.A1(new_n5482_), .A2(\asqrt[48] ), .ZN(new_n5484_));
  NAND3_X1   g05292(.A1(new_n5483_), .A2(new_n5484_), .A3(new_n1632_), .ZN(new_n5485_));
  AOI21_X1   g05293(.A1(new_n5483_), .A2(new_n5484_), .B(new_n1632_), .ZN(new_n5486_));
  AOI21_X1   g05294(.A1(new_n5376_), .A2(new_n5485_), .B(new_n5486_), .ZN(new_n5487_));
  AOI21_X1   g05295(.A1(new_n5487_), .A2(new_n1463_), .B(new_n5374_), .ZN(new_n5488_));
  NAND2_X1   g05296(.A1(new_n5485_), .A2(new_n5376_), .ZN(new_n5489_));
  INV_X1     g05297(.I(new_n5486_), .ZN(new_n5490_));
  AOI21_X1   g05298(.A1(new_n5489_), .A2(new_n5490_), .B(new_n1463_), .ZN(new_n5491_));
  NOR3_X1    g05299(.A1(new_n5488_), .A2(\asqrt[51] ), .A3(new_n5491_), .ZN(new_n5492_));
  OAI21_X1   g05300(.A1(new_n5488_), .A2(new_n5491_), .B(\asqrt[51] ), .ZN(new_n5493_));
  OAI21_X1   g05301(.A1(new_n5370_), .A2(new_n5492_), .B(new_n5493_), .ZN(new_n5494_));
  OAI21_X1   g05302(.A1(new_n5494_), .A2(\asqrt[52] ), .B(new_n5367_), .ZN(new_n5495_));
  NAND2_X1   g05303(.A1(new_n5494_), .A2(\asqrt[52] ), .ZN(new_n5496_));
  NAND3_X1   g05304(.A1(new_n5495_), .A2(new_n5496_), .A3(new_n1006_), .ZN(new_n5497_));
  AOI21_X1   g05305(.A1(new_n5495_), .A2(new_n5496_), .B(new_n1006_), .ZN(new_n5498_));
  AOI21_X1   g05306(.A1(new_n5364_), .A2(new_n5497_), .B(new_n5498_), .ZN(new_n5499_));
  AOI21_X1   g05307(.A1(new_n5499_), .A2(new_n860_), .B(new_n5362_), .ZN(new_n5500_));
  NAND2_X1   g05308(.A1(new_n5497_), .A2(new_n5364_), .ZN(new_n5501_));
  INV_X1     g05309(.I(new_n5498_), .ZN(new_n5502_));
  AOI21_X1   g05310(.A1(new_n5501_), .A2(new_n5502_), .B(new_n860_), .ZN(new_n5503_));
  NOR3_X1    g05311(.A1(new_n5500_), .A2(\asqrt[55] ), .A3(new_n5503_), .ZN(new_n5504_));
  OAI21_X1   g05312(.A1(new_n5500_), .A2(new_n5503_), .B(\asqrt[55] ), .ZN(new_n5505_));
  OAI21_X1   g05313(.A1(new_n5358_), .A2(new_n5504_), .B(new_n5505_), .ZN(new_n5506_));
  OAI21_X1   g05314(.A1(new_n5506_), .A2(\asqrt[56] ), .B(new_n5355_), .ZN(new_n5507_));
  NAND2_X1   g05315(.A1(new_n5506_), .A2(\asqrt[56] ), .ZN(new_n5508_));
  NAND3_X1   g05316(.A1(new_n5507_), .A2(new_n5508_), .A3(new_n531_), .ZN(new_n5509_));
  AOI21_X1   g05317(.A1(new_n5507_), .A2(new_n5508_), .B(new_n531_), .ZN(new_n5510_));
  AOI21_X1   g05318(.A1(new_n5352_), .A2(new_n5509_), .B(new_n5510_), .ZN(new_n5511_));
  AOI21_X1   g05319(.A1(new_n5511_), .A2(new_n423_), .B(new_n5350_), .ZN(new_n5512_));
  NAND2_X1   g05320(.A1(new_n5509_), .A2(new_n5352_), .ZN(new_n5513_));
  INV_X1     g05321(.I(new_n5510_), .ZN(new_n5514_));
  AOI21_X1   g05322(.A1(new_n5513_), .A2(new_n5514_), .B(new_n423_), .ZN(new_n5515_));
  NOR3_X1    g05323(.A1(new_n5512_), .A2(\asqrt[59] ), .A3(new_n5515_), .ZN(new_n5516_));
  NOR2_X1    g05324(.A1(new_n5516_), .A2(new_n5346_), .ZN(new_n5517_));
  OAI21_X1   g05325(.A1(new_n5512_), .A2(new_n5515_), .B(\asqrt[59] ), .ZN(new_n5518_));
  INV_X1     g05326(.I(new_n5518_), .ZN(new_n5519_));
  NOR2_X1    g05327(.A1(new_n5517_), .A2(new_n5519_), .ZN(new_n5520_));
  AOI21_X1   g05328(.A1(new_n5520_), .A2(new_n266_), .B(new_n5343_), .ZN(new_n5521_));
  INV_X1     g05329(.I(new_n5352_), .ZN(new_n5522_));
  INV_X1     g05330(.I(new_n5364_), .ZN(new_n5523_));
  INV_X1     g05331(.I(new_n5376_), .ZN(new_n5524_));
  INV_X1     g05332(.I(new_n5388_), .ZN(new_n5525_));
  INV_X1     g05333(.I(new_n5400_), .ZN(new_n5526_));
  INV_X1     g05334(.I(new_n5412_), .ZN(new_n5527_));
  NOR2_X1    g05335(.A1(new_n5428_), .A2(new_n5424_), .ZN(new_n5528_));
  NOR3_X1    g05336(.A1(new_n5336_), .A2(new_n5433_), .A3(new_n5430_), .ZN(new_n5529_));
  AOI21_X1   g05337(.A1(new_n5336_), .A2(\a[66] ), .B(new_n5431_), .ZN(new_n5530_));
  OAI21_X1   g05338(.A1(new_n5529_), .A2(new_n5530_), .B(\asqrt[34] ), .ZN(new_n5531_));
  INV_X1     g05339(.I(new_n5438_), .ZN(new_n5532_));
  NOR3_X1    g05340(.A1(new_n5336_), .A2(new_n5433_), .A3(new_n5532_), .ZN(new_n5533_));
  NOR3_X1    g05341(.A1(new_n5336_), .A2(\a[66] ), .A3(\a[67] ), .ZN(new_n5534_));
  AOI21_X1   g05342(.A1(\asqrt[33] ), .A2(new_n5433_), .B(new_n5440_), .ZN(new_n5535_));
  NOR3_X1    g05343(.A1(new_n5533_), .A2(new_n5534_), .A3(new_n5535_), .ZN(new_n5536_));
  NAND3_X1   g05344(.A1(new_n5536_), .A2(new_n5531_), .A3(new_n4751_), .ZN(new_n5537_));
  NAND2_X1   g05345(.A1(new_n5537_), .A2(new_n5528_), .ZN(new_n5538_));
  NAND3_X1   g05346(.A1(new_n5538_), .A2(new_n4461_), .A3(new_n5445_), .ZN(new_n5539_));
  AOI21_X1   g05347(.A1(new_n5538_), .A2(new_n5445_), .B(new_n4461_), .ZN(new_n5540_));
  AOI21_X1   g05348(.A1(new_n5418_), .A2(new_n5539_), .B(new_n5540_), .ZN(new_n5541_));
  AOI21_X1   g05349(.A1(new_n5541_), .A2(new_n4196_), .B(new_n5527_), .ZN(new_n5542_));
  NOR3_X1    g05350(.A1(new_n5542_), .A2(\asqrt[38] ), .A3(new_n5450_), .ZN(new_n5543_));
  OAI21_X1   g05351(.A1(new_n5542_), .A2(new_n5450_), .B(\asqrt[38] ), .ZN(new_n5544_));
  OAI21_X1   g05352(.A1(new_n5410_), .A2(new_n5543_), .B(new_n5544_), .ZN(new_n5545_));
  OAI21_X1   g05353(.A1(new_n5545_), .A2(\asqrt[39] ), .B(new_n5405_), .ZN(new_n5546_));
  NAND3_X1   g05354(.A1(new_n5546_), .A2(new_n3427_), .A3(new_n5457_), .ZN(new_n5547_));
  AOI21_X1   g05355(.A1(new_n5546_), .A2(new_n5457_), .B(new_n3427_), .ZN(new_n5548_));
  AOI21_X1   g05356(.A1(new_n5403_), .A2(new_n5547_), .B(new_n5548_), .ZN(new_n5549_));
  AOI21_X1   g05357(.A1(new_n5549_), .A2(new_n3195_), .B(new_n5526_), .ZN(new_n5550_));
  NOR3_X1    g05358(.A1(new_n5550_), .A2(\asqrt[42] ), .A3(new_n5462_), .ZN(new_n5551_));
  OAI21_X1   g05359(.A1(new_n5550_), .A2(new_n5462_), .B(\asqrt[42] ), .ZN(new_n5552_));
  OAI21_X1   g05360(.A1(new_n5398_), .A2(new_n5551_), .B(new_n5552_), .ZN(new_n5553_));
  OAI21_X1   g05361(.A1(new_n5553_), .A2(\asqrt[43] ), .B(new_n5393_), .ZN(new_n5554_));
  NAND3_X1   g05362(.A1(new_n5554_), .A2(new_n2531_), .A3(new_n5469_), .ZN(new_n5555_));
  AOI21_X1   g05363(.A1(new_n5554_), .A2(new_n5469_), .B(new_n2531_), .ZN(new_n5556_));
  AOI21_X1   g05364(.A1(new_n5391_), .A2(new_n5555_), .B(new_n5556_), .ZN(new_n5557_));
  AOI21_X1   g05365(.A1(new_n5557_), .A2(new_n2332_), .B(new_n5525_), .ZN(new_n5558_));
  NOR3_X1    g05366(.A1(new_n5558_), .A2(\asqrt[46] ), .A3(new_n5474_), .ZN(new_n5559_));
  OAI21_X1   g05367(.A1(new_n5558_), .A2(new_n5474_), .B(\asqrt[46] ), .ZN(new_n5560_));
  OAI21_X1   g05368(.A1(new_n5386_), .A2(new_n5559_), .B(new_n5560_), .ZN(new_n5561_));
  OAI21_X1   g05369(.A1(new_n5561_), .A2(\asqrt[47] ), .B(new_n5381_), .ZN(new_n5562_));
  NAND3_X1   g05370(.A1(new_n5562_), .A2(new_n1778_), .A3(new_n5481_), .ZN(new_n5563_));
  AOI21_X1   g05371(.A1(new_n5562_), .A2(new_n5481_), .B(new_n1778_), .ZN(new_n5564_));
  AOI21_X1   g05372(.A1(new_n5379_), .A2(new_n5563_), .B(new_n5564_), .ZN(new_n5565_));
  AOI21_X1   g05373(.A1(new_n5565_), .A2(new_n1632_), .B(new_n5524_), .ZN(new_n5566_));
  NOR3_X1    g05374(.A1(new_n5566_), .A2(\asqrt[50] ), .A3(new_n5486_), .ZN(new_n5567_));
  OAI21_X1   g05375(.A1(new_n5566_), .A2(new_n5486_), .B(\asqrt[50] ), .ZN(new_n5568_));
  OAI21_X1   g05376(.A1(new_n5374_), .A2(new_n5567_), .B(new_n5568_), .ZN(new_n5569_));
  OAI21_X1   g05377(.A1(new_n5569_), .A2(\asqrt[51] ), .B(new_n5369_), .ZN(new_n5570_));
  NAND3_X1   g05378(.A1(new_n5570_), .A2(new_n1150_), .A3(new_n5493_), .ZN(new_n5571_));
  AOI21_X1   g05379(.A1(new_n5570_), .A2(new_n5493_), .B(new_n1150_), .ZN(new_n5572_));
  AOI21_X1   g05380(.A1(new_n5367_), .A2(new_n5571_), .B(new_n5572_), .ZN(new_n5573_));
  AOI21_X1   g05381(.A1(new_n5573_), .A2(new_n1006_), .B(new_n5523_), .ZN(new_n5574_));
  NOR3_X1    g05382(.A1(new_n5574_), .A2(\asqrt[54] ), .A3(new_n5498_), .ZN(new_n5575_));
  OAI21_X1   g05383(.A1(new_n5574_), .A2(new_n5498_), .B(\asqrt[54] ), .ZN(new_n5576_));
  OAI21_X1   g05384(.A1(new_n5362_), .A2(new_n5575_), .B(new_n5576_), .ZN(new_n5577_));
  OAI21_X1   g05385(.A1(new_n5577_), .A2(\asqrt[55] ), .B(new_n5357_), .ZN(new_n5578_));
  NAND3_X1   g05386(.A1(new_n5578_), .A2(new_n634_), .A3(new_n5505_), .ZN(new_n5579_));
  AOI21_X1   g05387(.A1(new_n5578_), .A2(new_n5505_), .B(new_n634_), .ZN(new_n5580_));
  AOI21_X1   g05388(.A1(new_n5355_), .A2(new_n5579_), .B(new_n5580_), .ZN(new_n5581_));
  AOI21_X1   g05389(.A1(new_n5581_), .A2(new_n531_), .B(new_n5522_), .ZN(new_n5582_));
  NOR3_X1    g05390(.A1(new_n5582_), .A2(\asqrt[58] ), .A3(new_n5510_), .ZN(new_n5583_));
  OAI21_X1   g05391(.A1(new_n5582_), .A2(new_n5510_), .B(\asqrt[58] ), .ZN(new_n5584_));
  OAI21_X1   g05392(.A1(new_n5350_), .A2(new_n5583_), .B(new_n5584_), .ZN(new_n5585_));
  OAI21_X1   g05393(.A1(new_n5585_), .A2(\asqrt[59] ), .B(new_n5345_), .ZN(new_n5586_));
  AOI21_X1   g05394(.A1(new_n5586_), .A2(new_n5518_), .B(new_n266_), .ZN(new_n5587_));
  OAI21_X1   g05395(.A1(new_n5521_), .A2(new_n5587_), .B(\asqrt[61] ), .ZN(new_n5588_));
  AOI21_X1   g05396(.A1(new_n5296_), .A2(new_n5290_), .B(\asqrt[33] ), .ZN(new_n5589_));
  XOR2_X1    g05397(.A1(new_n5589_), .A2(new_n5034_), .Z(new_n5590_));
  OAI21_X1   g05398(.A1(new_n5346_), .A2(new_n5516_), .B(new_n5518_), .ZN(new_n5591_));
  OAI21_X1   g05399(.A1(new_n5591_), .A2(\asqrt[60] ), .B(new_n5342_), .ZN(new_n5592_));
  OAI21_X1   g05400(.A1(new_n5517_), .A2(new_n5519_), .B(\asqrt[60] ), .ZN(new_n5593_));
  NAND3_X1   g05401(.A1(new_n5592_), .A2(new_n239_), .A3(new_n5593_), .ZN(new_n5594_));
  NAND2_X1   g05402(.A1(new_n5594_), .A2(new_n5590_), .ZN(new_n5595_));
  NAND2_X1   g05403(.A1(new_n5595_), .A2(new_n5588_), .ZN(new_n5596_));
  AOI21_X1   g05404(.A1(new_n5592_), .A2(new_n5593_), .B(new_n239_), .ZN(new_n5597_));
  NAND3_X1   g05405(.A1(new_n5586_), .A2(new_n266_), .A3(new_n5518_), .ZN(new_n5598_));
  AOI21_X1   g05406(.A1(new_n5342_), .A2(new_n5598_), .B(new_n5587_), .ZN(new_n5599_));
  INV_X1     g05407(.I(new_n5590_), .ZN(new_n5600_));
  AOI21_X1   g05408(.A1(new_n5599_), .A2(new_n239_), .B(new_n5600_), .ZN(new_n5601_));
  OAI21_X1   g05409(.A1(new_n5601_), .A2(new_n5597_), .B(new_n201_), .ZN(new_n5602_));
  NAND3_X1   g05410(.A1(new_n5595_), .A2(\asqrt[62] ), .A3(new_n5588_), .ZN(new_n5603_));
  AOI21_X1   g05411(.A1(new_n5289_), .A2(new_n5327_), .B(\asqrt[33] ), .ZN(new_n5604_));
  XOR2_X1    g05412(.A1(new_n5604_), .A2(new_n5293_), .Z(new_n5605_));
  INV_X1     g05413(.I(new_n5605_), .ZN(new_n5606_));
  AOI22_X1   g05414(.A1(new_n5602_), .A2(new_n5603_), .B1(new_n5596_), .B2(new_n5606_), .ZN(new_n5607_));
  NOR2_X1    g05415(.A1(new_n5308_), .A2(new_n5032_), .ZN(new_n5608_));
  OAI21_X1   g05416(.A1(\asqrt[33] ), .A2(new_n5608_), .B(new_n5315_), .ZN(new_n5609_));
  INV_X1     g05417(.I(new_n5609_), .ZN(new_n5610_));
  OAI21_X1   g05418(.A1(new_n5607_), .A2(new_n5339_), .B(new_n5610_), .ZN(new_n5611_));
  OAI21_X1   g05419(.A1(new_n5596_), .A2(\asqrt[62] ), .B(new_n5605_), .ZN(new_n5612_));
  NAND2_X1   g05420(.A1(new_n5596_), .A2(\asqrt[62] ), .ZN(new_n5613_));
  NAND3_X1   g05421(.A1(new_n5612_), .A2(new_n5613_), .A3(new_n5339_), .ZN(new_n5614_));
  NAND2_X1   g05422(.A1(new_n5336_), .A2(new_n5031_), .ZN(new_n5615_));
  XOR2_X1    g05423(.A1(new_n5308_), .A2(new_n5032_), .Z(new_n5616_));
  NAND3_X1   g05424(.A1(new_n5615_), .A2(\asqrt[63] ), .A3(new_n5616_), .ZN(new_n5617_));
  INV_X1     g05425(.I(new_n5425_), .ZN(new_n5618_));
  NAND4_X1   g05426(.A1(new_n5618_), .A2(new_n5032_), .A3(new_n5315_), .A4(new_n5322_), .ZN(new_n5619_));
  NAND2_X1   g05427(.A1(new_n5617_), .A2(new_n5619_), .ZN(new_n5620_));
  INV_X1     g05428(.I(new_n5620_), .ZN(new_n5621_));
  NAND4_X1   g05429(.A1(new_n5611_), .A2(new_n193_), .A3(new_n5614_), .A4(new_n5621_), .ZN(\asqrt[32] ));
  INV_X1     g05430(.I(\a[64] ), .ZN(new_n5623_));
  NAND2_X1   g05431(.A1(\asqrt[32] ), .A2(new_n5623_), .ZN(new_n5624_));
  NOR2_X1    g05432(.A1(new_n194_), .A2(\a[64] ), .ZN(new_n5625_));
  AOI22_X1   g05433(.A1(new_n5624_), .A2(new_n194_), .B1(\asqrt[32] ), .B2(new_n5625_), .ZN(new_n5626_));
  NOR2_X1    g05434(.A1(\a[62] ), .A2(\a[63] ), .ZN(new_n5627_));
  INV_X1     g05435(.I(new_n5627_), .ZN(new_n5628_));
  NAND3_X1   g05436(.A1(\asqrt[32] ), .A2(\a[64] ), .A3(new_n5628_), .ZN(new_n5629_));
  OAI21_X1   g05437(.A1(\asqrt[32] ), .A2(new_n5623_), .B(new_n5627_), .ZN(new_n5630_));
  AOI21_X1   g05438(.A1(new_n5630_), .A2(new_n5629_), .B(new_n5336_), .ZN(new_n5631_));
  NOR2_X1    g05439(.A1(new_n5596_), .A2(\asqrt[62] ), .ZN(new_n5632_));
  INV_X1     g05440(.I(new_n5613_), .ZN(new_n5633_));
  NOR2_X1    g05441(.A1(new_n5633_), .A2(new_n5632_), .ZN(new_n5634_));
  NOR2_X1    g05442(.A1(new_n5601_), .A2(new_n5597_), .ZN(new_n5635_));
  AOI21_X1   g05443(.A1(new_n5595_), .A2(new_n5588_), .B(\asqrt[62] ), .ZN(new_n5636_));
  NOR3_X1    g05444(.A1(new_n5601_), .A2(new_n201_), .A3(new_n5597_), .ZN(new_n5637_));
  OAI22_X1   g05445(.A1(new_n5637_), .A2(new_n5636_), .B1(new_n5635_), .B2(new_n5605_), .ZN(new_n5638_));
  AOI21_X1   g05446(.A1(new_n5638_), .A2(new_n5338_), .B(new_n5609_), .ZN(new_n5639_));
  AOI21_X1   g05447(.A1(new_n5635_), .A2(new_n201_), .B(new_n5606_), .ZN(new_n5640_));
  OAI21_X1   g05448(.A1(new_n5635_), .A2(new_n201_), .B(new_n5339_), .ZN(new_n5641_));
  NOR2_X1    g05449(.A1(new_n5640_), .A2(new_n5641_), .ZN(new_n5642_));
  NOR4_X1    g05450(.A1(new_n5639_), .A2(\asqrt[63] ), .A3(new_n5642_), .A4(new_n5620_), .ZN(new_n5643_));
  XOR2_X1    g05451(.A1(new_n5604_), .A2(new_n5293_), .Z(new_n5644_));
  OAI21_X1   g05452(.A1(\asqrt[32] ), .A2(new_n5634_), .B(new_n5644_), .ZN(new_n5645_));
  NOR2_X1    g05453(.A1(new_n5519_), .A2(new_n5516_), .ZN(new_n5646_));
  NOR2_X1    g05454(.A1(\asqrt[32] ), .A2(new_n5646_), .ZN(new_n5647_));
  XOR2_X1    g05455(.A1(new_n5647_), .A2(new_n5345_), .Z(new_n5648_));
  NOR2_X1    g05456(.A1(new_n5583_), .A2(new_n5515_), .ZN(new_n5649_));
  NOR2_X1    g05457(.A1(\asqrt[32] ), .A2(new_n5649_), .ZN(new_n5650_));
  XOR2_X1    g05458(.A1(new_n5650_), .A2(new_n5349_), .Z(new_n5651_));
  AOI21_X1   g05459(.A1(new_n5509_), .A2(new_n5514_), .B(\asqrt[32] ), .ZN(new_n5652_));
  XOR2_X1    g05460(.A1(new_n5652_), .A2(new_n5352_), .Z(new_n5653_));
  INV_X1     g05461(.I(new_n5653_), .ZN(new_n5654_));
  AOI21_X1   g05462(.A1(new_n5579_), .A2(new_n5508_), .B(\asqrt[32] ), .ZN(new_n5655_));
  XOR2_X1    g05463(.A1(new_n5655_), .A2(new_n5355_), .Z(new_n5656_));
  INV_X1     g05464(.I(new_n5656_), .ZN(new_n5657_));
  INV_X1     g05465(.I(new_n5505_), .ZN(new_n5658_));
  NOR2_X1    g05466(.A1(new_n5658_), .A2(new_n5504_), .ZN(new_n5659_));
  NOR2_X1    g05467(.A1(\asqrt[32] ), .A2(new_n5659_), .ZN(new_n5660_));
  XOR2_X1    g05468(.A1(new_n5660_), .A2(new_n5357_), .Z(new_n5661_));
  NOR2_X1    g05469(.A1(new_n5575_), .A2(new_n5503_), .ZN(new_n5662_));
  NOR2_X1    g05470(.A1(\asqrt[32] ), .A2(new_n5662_), .ZN(new_n5663_));
  XOR2_X1    g05471(.A1(new_n5663_), .A2(new_n5361_), .Z(new_n5664_));
  AOI21_X1   g05472(.A1(new_n5497_), .A2(new_n5502_), .B(\asqrt[32] ), .ZN(new_n5665_));
  XOR2_X1    g05473(.A1(new_n5665_), .A2(new_n5364_), .Z(new_n5666_));
  INV_X1     g05474(.I(new_n5666_), .ZN(new_n5667_));
  AOI21_X1   g05475(.A1(new_n5571_), .A2(new_n5496_), .B(\asqrt[32] ), .ZN(new_n5668_));
  XOR2_X1    g05476(.A1(new_n5668_), .A2(new_n5367_), .Z(new_n5669_));
  INV_X1     g05477(.I(new_n5669_), .ZN(new_n5670_));
  XOR2_X1    g05478(.A1(new_n5569_), .A2(\asqrt[51] ), .Z(new_n5671_));
  NOR2_X1    g05479(.A1(\asqrt[32] ), .A2(new_n5671_), .ZN(new_n5672_));
  XOR2_X1    g05480(.A1(new_n5672_), .A2(new_n5369_), .Z(new_n5673_));
  NOR2_X1    g05481(.A1(new_n5567_), .A2(new_n5491_), .ZN(new_n5674_));
  NOR2_X1    g05482(.A1(\asqrt[32] ), .A2(new_n5674_), .ZN(new_n5675_));
  XOR2_X1    g05483(.A1(new_n5675_), .A2(new_n5373_), .Z(new_n5676_));
  AOI21_X1   g05484(.A1(new_n5485_), .A2(new_n5490_), .B(\asqrt[32] ), .ZN(new_n5677_));
  XOR2_X1    g05485(.A1(new_n5677_), .A2(new_n5376_), .Z(new_n5678_));
  INV_X1     g05486(.I(new_n5678_), .ZN(new_n5679_));
  AOI21_X1   g05487(.A1(new_n5563_), .A2(new_n5484_), .B(\asqrt[32] ), .ZN(new_n5680_));
  XOR2_X1    g05488(.A1(new_n5680_), .A2(new_n5379_), .Z(new_n5681_));
  INV_X1     g05489(.I(new_n5681_), .ZN(new_n5682_));
  XOR2_X1    g05490(.A1(new_n5561_), .A2(\asqrt[47] ), .Z(new_n5683_));
  NOR2_X1    g05491(.A1(\asqrt[32] ), .A2(new_n5683_), .ZN(new_n5684_));
  XOR2_X1    g05492(.A1(new_n5684_), .A2(new_n5381_), .Z(new_n5685_));
  NOR2_X1    g05493(.A1(new_n5559_), .A2(new_n5479_), .ZN(new_n5686_));
  NOR2_X1    g05494(.A1(\asqrt[32] ), .A2(new_n5686_), .ZN(new_n5687_));
  XOR2_X1    g05495(.A1(new_n5687_), .A2(new_n5385_), .Z(new_n5688_));
  AOI21_X1   g05496(.A1(new_n5473_), .A2(new_n5478_), .B(\asqrt[32] ), .ZN(new_n5689_));
  XOR2_X1    g05497(.A1(new_n5689_), .A2(new_n5388_), .Z(new_n5690_));
  INV_X1     g05498(.I(new_n5690_), .ZN(new_n5691_));
  AOI21_X1   g05499(.A1(new_n5555_), .A2(new_n5472_), .B(\asqrt[32] ), .ZN(new_n5692_));
  XOR2_X1    g05500(.A1(new_n5692_), .A2(new_n5391_), .Z(new_n5693_));
  INV_X1     g05501(.I(new_n5693_), .ZN(new_n5694_));
  XOR2_X1    g05502(.A1(new_n5553_), .A2(\asqrt[43] ), .Z(new_n5695_));
  NOR2_X1    g05503(.A1(\asqrt[32] ), .A2(new_n5695_), .ZN(new_n5696_));
  XOR2_X1    g05504(.A1(new_n5696_), .A2(new_n5393_), .Z(new_n5697_));
  NOR2_X1    g05505(.A1(new_n5551_), .A2(new_n5467_), .ZN(new_n5698_));
  NOR2_X1    g05506(.A1(\asqrt[32] ), .A2(new_n5698_), .ZN(new_n5699_));
  XOR2_X1    g05507(.A1(new_n5699_), .A2(new_n5397_), .Z(new_n5700_));
  AOI21_X1   g05508(.A1(new_n5461_), .A2(new_n5466_), .B(\asqrt[32] ), .ZN(new_n5701_));
  XOR2_X1    g05509(.A1(new_n5701_), .A2(new_n5400_), .Z(new_n5702_));
  INV_X1     g05510(.I(new_n5702_), .ZN(new_n5703_));
  AOI21_X1   g05511(.A1(new_n5547_), .A2(new_n5460_), .B(\asqrt[32] ), .ZN(new_n5704_));
  XOR2_X1    g05512(.A1(new_n5704_), .A2(new_n5403_), .Z(new_n5705_));
  INV_X1     g05513(.I(new_n5705_), .ZN(new_n5706_));
  XOR2_X1    g05514(.A1(new_n5545_), .A2(\asqrt[39] ), .Z(new_n5707_));
  NOR2_X1    g05515(.A1(\asqrt[32] ), .A2(new_n5707_), .ZN(new_n5708_));
  XOR2_X1    g05516(.A1(new_n5708_), .A2(new_n5405_), .Z(new_n5709_));
  NOR2_X1    g05517(.A1(new_n5543_), .A2(new_n5455_), .ZN(new_n5710_));
  NOR2_X1    g05518(.A1(\asqrt[32] ), .A2(new_n5710_), .ZN(new_n5711_));
  XOR2_X1    g05519(.A1(new_n5711_), .A2(new_n5409_), .Z(new_n5712_));
  AOI21_X1   g05520(.A1(new_n5449_), .A2(new_n5454_), .B(\asqrt[32] ), .ZN(new_n5713_));
  XOR2_X1    g05521(.A1(new_n5713_), .A2(new_n5412_), .Z(new_n5714_));
  INV_X1     g05522(.I(new_n5714_), .ZN(new_n5715_));
  AOI21_X1   g05523(.A1(new_n5539_), .A2(new_n5448_), .B(\asqrt[32] ), .ZN(new_n5716_));
  XOR2_X1    g05524(.A1(new_n5716_), .A2(new_n5418_), .Z(new_n5717_));
  INV_X1     g05525(.I(new_n5717_), .ZN(new_n5718_));
  AOI21_X1   g05526(.A1(new_n5537_), .A2(new_n5445_), .B(\asqrt[32] ), .ZN(new_n5719_));
  XOR2_X1    g05527(.A1(new_n5719_), .A2(new_n5528_), .Z(new_n5720_));
  NAND2_X1   g05528(.A1(\asqrt[33] ), .A2(new_n5433_), .ZN(new_n5721_));
  NOR2_X1    g05529(.A1(new_n5440_), .A2(\a[66] ), .ZN(new_n5722_));
  AOI22_X1   g05530(.A1(new_n5721_), .A2(new_n5440_), .B1(\asqrt[33] ), .B2(new_n5722_), .ZN(new_n5723_));
  OAI21_X1   g05531(.A1(new_n5336_), .A2(new_n5433_), .B(new_n5532_), .ZN(new_n5724_));
  AOI21_X1   g05532(.A1(new_n5531_), .A2(new_n5724_), .B(\asqrt[32] ), .ZN(new_n5725_));
  XOR2_X1    g05533(.A1(new_n5725_), .A2(new_n5723_), .Z(new_n5726_));
  NAND2_X1   g05534(.A1(new_n5611_), .A2(new_n193_), .ZN(new_n5727_));
  NAND3_X1   g05535(.A1(new_n5617_), .A2(\asqrt[33] ), .A3(new_n5619_), .ZN(new_n5728_));
  NOR3_X1    g05536(.A1(new_n5727_), .A2(new_n5642_), .A3(new_n5728_), .ZN(new_n5729_));
  NOR2_X1    g05537(.A1(new_n5643_), .A2(new_n5431_), .ZN(new_n5730_));
  OAI21_X1   g05538(.A1(new_n5730_), .A2(new_n5729_), .B(new_n5433_), .ZN(new_n5731_));
  NOR3_X1    g05539(.A1(new_n5639_), .A2(\asqrt[63] ), .A3(new_n5642_), .ZN(new_n5732_));
  NAND4_X1   g05540(.A1(new_n5732_), .A2(\asqrt[33] ), .A3(new_n5617_), .A4(new_n5619_), .ZN(new_n5733_));
  NAND2_X1   g05541(.A1(\asqrt[32] ), .A2(new_n5430_), .ZN(new_n5734_));
  NAND3_X1   g05542(.A1(new_n5733_), .A2(new_n5734_), .A3(\a[66] ), .ZN(new_n5735_));
  NAND2_X1   g05543(.A1(new_n5735_), .A2(new_n5731_), .ZN(new_n5736_));
  NAND2_X1   g05544(.A1(new_n5627_), .A2(new_n5623_), .ZN(new_n5737_));
  NAND3_X1   g05545(.A1(new_n5318_), .A2(new_n5320_), .A3(new_n5737_), .ZN(new_n5738_));
  NAND2_X1   g05546(.A1(new_n5419_), .A2(new_n5738_), .ZN(new_n5739_));
  NAND3_X1   g05547(.A1(\asqrt[32] ), .A2(\a[64] ), .A3(new_n5739_), .ZN(new_n5740_));
  NAND3_X1   g05548(.A1(\asqrt[32] ), .A2(new_n5623_), .A3(new_n194_), .ZN(new_n5741_));
  OAI21_X1   g05549(.A1(new_n5643_), .A2(\a[64] ), .B(\a[65] ), .ZN(new_n5742_));
  NAND3_X1   g05550(.A1(new_n5742_), .A2(new_n5740_), .A3(new_n5741_), .ZN(new_n5743_));
  NOR3_X1    g05551(.A1(new_n5743_), .A2(new_n5631_), .A3(\asqrt[34] ), .ZN(new_n5744_));
  OAI21_X1   g05552(.A1(new_n5743_), .A2(new_n5631_), .B(\asqrt[34] ), .ZN(new_n5745_));
  OAI21_X1   g05553(.A1(new_n5736_), .A2(new_n5744_), .B(new_n5745_), .ZN(new_n5746_));
  OAI21_X1   g05554(.A1(new_n5746_), .A2(\asqrt[35] ), .B(new_n5726_), .ZN(new_n5747_));
  NAND2_X1   g05555(.A1(new_n5746_), .A2(\asqrt[35] ), .ZN(new_n5748_));
  NAND3_X1   g05556(.A1(new_n5747_), .A2(new_n5748_), .A3(new_n4461_), .ZN(new_n5749_));
  AOI21_X1   g05557(.A1(new_n5747_), .A2(new_n5748_), .B(new_n4461_), .ZN(new_n5750_));
  AOI21_X1   g05558(.A1(new_n5720_), .A2(new_n5749_), .B(new_n5750_), .ZN(new_n5751_));
  AOI21_X1   g05559(.A1(new_n5751_), .A2(new_n4196_), .B(new_n5718_), .ZN(new_n5752_));
  NAND2_X1   g05560(.A1(new_n5749_), .A2(new_n5720_), .ZN(new_n5753_));
  INV_X1     g05561(.I(new_n5726_), .ZN(new_n5754_));
  INV_X1     g05562(.I(new_n5736_), .ZN(new_n5755_));
  NOR3_X1    g05563(.A1(new_n5643_), .A2(new_n5623_), .A3(new_n5627_), .ZN(new_n5756_));
  AOI21_X1   g05564(.A1(new_n5643_), .A2(\a[64] ), .B(new_n5628_), .ZN(new_n5757_));
  OAI21_X1   g05565(.A1(new_n5756_), .A2(new_n5757_), .B(\asqrt[33] ), .ZN(new_n5758_));
  INV_X1     g05566(.I(new_n5739_), .ZN(new_n5759_));
  NOR3_X1    g05567(.A1(new_n5643_), .A2(new_n5623_), .A3(new_n5759_), .ZN(new_n5760_));
  NOR3_X1    g05568(.A1(new_n5643_), .A2(\a[64] ), .A3(\a[65] ), .ZN(new_n5761_));
  AOI21_X1   g05569(.A1(\asqrt[32] ), .A2(new_n5623_), .B(new_n194_), .ZN(new_n5762_));
  NOR3_X1    g05570(.A1(new_n5760_), .A2(new_n5761_), .A3(new_n5762_), .ZN(new_n5763_));
  NAND3_X1   g05571(.A1(new_n5758_), .A2(new_n5763_), .A3(new_n5029_), .ZN(new_n5764_));
  AOI21_X1   g05572(.A1(new_n5758_), .A2(new_n5763_), .B(new_n5029_), .ZN(new_n5765_));
  AOI21_X1   g05573(.A1(new_n5755_), .A2(new_n5764_), .B(new_n5765_), .ZN(new_n5766_));
  AOI21_X1   g05574(.A1(new_n5766_), .A2(new_n4751_), .B(new_n5754_), .ZN(new_n5767_));
  NAND2_X1   g05575(.A1(new_n5755_), .A2(new_n5764_), .ZN(new_n5768_));
  AOI21_X1   g05576(.A1(new_n5768_), .A2(new_n5745_), .B(new_n4751_), .ZN(new_n5769_));
  OAI21_X1   g05577(.A1(new_n5767_), .A2(new_n5769_), .B(\asqrt[36] ), .ZN(new_n5770_));
  AOI21_X1   g05578(.A1(new_n5753_), .A2(new_n5770_), .B(new_n4196_), .ZN(new_n5771_));
  NOR3_X1    g05579(.A1(new_n5752_), .A2(\asqrt[38] ), .A3(new_n5771_), .ZN(new_n5772_));
  OAI21_X1   g05580(.A1(new_n5752_), .A2(new_n5771_), .B(\asqrt[38] ), .ZN(new_n5773_));
  OAI21_X1   g05581(.A1(new_n5715_), .A2(new_n5772_), .B(new_n5773_), .ZN(new_n5774_));
  OAI21_X1   g05582(.A1(new_n5774_), .A2(\asqrt[39] ), .B(new_n5712_), .ZN(new_n5775_));
  NAND2_X1   g05583(.A1(new_n5774_), .A2(\asqrt[39] ), .ZN(new_n5776_));
  NAND3_X1   g05584(.A1(new_n5775_), .A2(new_n5776_), .A3(new_n3427_), .ZN(new_n5777_));
  AOI21_X1   g05585(.A1(new_n5775_), .A2(new_n5776_), .B(new_n3427_), .ZN(new_n5778_));
  AOI21_X1   g05586(.A1(new_n5709_), .A2(new_n5777_), .B(new_n5778_), .ZN(new_n5779_));
  AOI21_X1   g05587(.A1(new_n5779_), .A2(new_n3195_), .B(new_n5706_), .ZN(new_n5780_));
  NAND2_X1   g05588(.A1(new_n5777_), .A2(new_n5709_), .ZN(new_n5781_));
  INV_X1     g05589(.I(new_n5712_), .ZN(new_n5782_));
  INV_X1     g05590(.I(new_n5720_), .ZN(new_n5783_));
  NOR3_X1    g05591(.A1(new_n5767_), .A2(\asqrt[36] ), .A3(new_n5769_), .ZN(new_n5784_));
  OAI21_X1   g05592(.A1(new_n5783_), .A2(new_n5784_), .B(new_n5770_), .ZN(new_n5785_));
  OAI21_X1   g05593(.A1(new_n5785_), .A2(\asqrt[37] ), .B(new_n5717_), .ZN(new_n5786_));
  NAND2_X1   g05594(.A1(new_n5785_), .A2(\asqrt[37] ), .ZN(new_n5787_));
  NAND3_X1   g05595(.A1(new_n5786_), .A2(new_n5787_), .A3(new_n3925_), .ZN(new_n5788_));
  AOI21_X1   g05596(.A1(new_n5786_), .A2(new_n5787_), .B(new_n3925_), .ZN(new_n5789_));
  AOI21_X1   g05597(.A1(new_n5714_), .A2(new_n5788_), .B(new_n5789_), .ZN(new_n5790_));
  AOI21_X1   g05598(.A1(new_n5790_), .A2(new_n3681_), .B(new_n5782_), .ZN(new_n5791_));
  NAND2_X1   g05599(.A1(new_n5788_), .A2(new_n5714_), .ZN(new_n5792_));
  AOI21_X1   g05600(.A1(new_n5792_), .A2(new_n5773_), .B(new_n3681_), .ZN(new_n5793_));
  OAI21_X1   g05601(.A1(new_n5791_), .A2(new_n5793_), .B(\asqrt[40] ), .ZN(new_n5794_));
  AOI21_X1   g05602(.A1(new_n5781_), .A2(new_n5794_), .B(new_n3195_), .ZN(new_n5795_));
  NOR3_X1    g05603(.A1(new_n5780_), .A2(\asqrt[42] ), .A3(new_n5795_), .ZN(new_n5796_));
  OAI21_X1   g05604(.A1(new_n5780_), .A2(new_n5795_), .B(\asqrt[42] ), .ZN(new_n5797_));
  OAI21_X1   g05605(.A1(new_n5703_), .A2(new_n5796_), .B(new_n5797_), .ZN(new_n5798_));
  OAI21_X1   g05606(.A1(new_n5798_), .A2(\asqrt[43] ), .B(new_n5700_), .ZN(new_n5799_));
  NAND2_X1   g05607(.A1(new_n5798_), .A2(\asqrt[43] ), .ZN(new_n5800_));
  NAND3_X1   g05608(.A1(new_n5799_), .A2(new_n5800_), .A3(new_n2531_), .ZN(new_n5801_));
  AOI21_X1   g05609(.A1(new_n5799_), .A2(new_n5800_), .B(new_n2531_), .ZN(new_n5802_));
  AOI21_X1   g05610(.A1(new_n5697_), .A2(new_n5801_), .B(new_n5802_), .ZN(new_n5803_));
  AOI21_X1   g05611(.A1(new_n5803_), .A2(new_n2332_), .B(new_n5694_), .ZN(new_n5804_));
  NAND2_X1   g05612(.A1(new_n5801_), .A2(new_n5697_), .ZN(new_n5805_));
  INV_X1     g05613(.I(new_n5700_), .ZN(new_n5806_));
  INV_X1     g05614(.I(new_n5709_), .ZN(new_n5807_));
  NOR3_X1    g05615(.A1(new_n5791_), .A2(\asqrt[40] ), .A3(new_n5793_), .ZN(new_n5808_));
  OAI21_X1   g05616(.A1(new_n5807_), .A2(new_n5808_), .B(new_n5794_), .ZN(new_n5809_));
  OAI21_X1   g05617(.A1(new_n5809_), .A2(\asqrt[41] ), .B(new_n5705_), .ZN(new_n5810_));
  NAND2_X1   g05618(.A1(new_n5809_), .A2(\asqrt[41] ), .ZN(new_n5811_));
  NAND3_X1   g05619(.A1(new_n5810_), .A2(new_n5811_), .A3(new_n2960_), .ZN(new_n5812_));
  AOI21_X1   g05620(.A1(new_n5810_), .A2(new_n5811_), .B(new_n2960_), .ZN(new_n5813_));
  AOI21_X1   g05621(.A1(new_n5702_), .A2(new_n5812_), .B(new_n5813_), .ZN(new_n5814_));
  AOI21_X1   g05622(.A1(new_n5814_), .A2(new_n2749_), .B(new_n5806_), .ZN(new_n5815_));
  NAND2_X1   g05623(.A1(new_n5812_), .A2(new_n5702_), .ZN(new_n5816_));
  AOI21_X1   g05624(.A1(new_n5816_), .A2(new_n5797_), .B(new_n2749_), .ZN(new_n5817_));
  OAI21_X1   g05625(.A1(new_n5815_), .A2(new_n5817_), .B(\asqrt[44] ), .ZN(new_n5818_));
  AOI21_X1   g05626(.A1(new_n5805_), .A2(new_n5818_), .B(new_n2332_), .ZN(new_n5819_));
  NOR3_X1    g05627(.A1(new_n5804_), .A2(\asqrt[46] ), .A3(new_n5819_), .ZN(new_n5820_));
  OAI21_X1   g05628(.A1(new_n5804_), .A2(new_n5819_), .B(\asqrt[46] ), .ZN(new_n5821_));
  OAI21_X1   g05629(.A1(new_n5691_), .A2(new_n5820_), .B(new_n5821_), .ZN(new_n5822_));
  OAI21_X1   g05630(.A1(new_n5822_), .A2(\asqrt[47] ), .B(new_n5688_), .ZN(new_n5823_));
  NAND2_X1   g05631(.A1(new_n5822_), .A2(\asqrt[47] ), .ZN(new_n5824_));
  NAND3_X1   g05632(.A1(new_n5823_), .A2(new_n5824_), .A3(new_n1778_), .ZN(new_n5825_));
  AOI21_X1   g05633(.A1(new_n5823_), .A2(new_n5824_), .B(new_n1778_), .ZN(new_n5826_));
  AOI21_X1   g05634(.A1(new_n5685_), .A2(new_n5825_), .B(new_n5826_), .ZN(new_n5827_));
  AOI21_X1   g05635(.A1(new_n5827_), .A2(new_n1632_), .B(new_n5682_), .ZN(new_n5828_));
  NAND2_X1   g05636(.A1(new_n5825_), .A2(new_n5685_), .ZN(new_n5829_));
  INV_X1     g05637(.I(new_n5688_), .ZN(new_n5830_));
  INV_X1     g05638(.I(new_n5697_), .ZN(new_n5831_));
  NOR3_X1    g05639(.A1(new_n5815_), .A2(\asqrt[44] ), .A3(new_n5817_), .ZN(new_n5832_));
  OAI21_X1   g05640(.A1(new_n5831_), .A2(new_n5832_), .B(new_n5818_), .ZN(new_n5833_));
  OAI21_X1   g05641(.A1(new_n5833_), .A2(\asqrt[45] ), .B(new_n5693_), .ZN(new_n5834_));
  NAND2_X1   g05642(.A1(new_n5833_), .A2(\asqrt[45] ), .ZN(new_n5835_));
  NAND3_X1   g05643(.A1(new_n5834_), .A2(new_n5835_), .A3(new_n2134_), .ZN(new_n5836_));
  AOI21_X1   g05644(.A1(new_n5834_), .A2(new_n5835_), .B(new_n2134_), .ZN(new_n5837_));
  AOI21_X1   g05645(.A1(new_n5690_), .A2(new_n5836_), .B(new_n5837_), .ZN(new_n5838_));
  AOI21_X1   g05646(.A1(new_n5838_), .A2(new_n1953_), .B(new_n5830_), .ZN(new_n5839_));
  NAND2_X1   g05647(.A1(new_n5836_), .A2(new_n5690_), .ZN(new_n5840_));
  AOI21_X1   g05648(.A1(new_n5840_), .A2(new_n5821_), .B(new_n1953_), .ZN(new_n5841_));
  OAI21_X1   g05649(.A1(new_n5839_), .A2(new_n5841_), .B(\asqrt[48] ), .ZN(new_n5842_));
  AOI21_X1   g05650(.A1(new_n5829_), .A2(new_n5842_), .B(new_n1632_), .ZN(new_n5843_));
  NOR3_X1    g05651(.A1(new_n5828_), .A2(\asqrt[50] ), .A3(new_n5843_), .ZN(new_n5844_));
  OAI21_X1   g05652(.A1(new_n5828_), .A2(new_n5843_), .B(\asqrt[50] ), .ZN(new_n5845_));
  OAI21_X1   g05653(.A1(new_n5679_), .A2(new_n5844_), .B(new_n5845_), .ZN(new_n5846_));
  OAI21_X1   g05654(.A1(new_n5846_), .A2(\asqrt[51] ), .B(new_n5676_), .ZN(new_n5847_));
  NAND2_X1   g05655(.A1(new_n5846_), .A2(\asqrt[51] ), .ZN(new_n5848_));
  NAND3_X1   g05656(.A1(new_n5847_), .A2(new_n5848_), .A3(new_n1150_), .ZN(new_n5849_));
  AOI21_X1   g05657(.A1(new_n5847_), .A2(new_n5848_), .B(new_n1150_), .ZN(new_n5850_));
  AOI21_X1   g05658(.A1(new_n5673_), .A2(new_n5849_), .B(new_n5850_), .ZN(new_n5851_));
  AOI21_X1   g05659(.A1(new_n5851_), .A2(new_n1006_), .B(new_n5670_), .ZN(new_n5852_));
  NAND2_X1   g05660(.A1(new_n5849_), .A2(new_n5673_), .ZN(new_n5853_));
  INV_X1     g05661(.I(new_n5676_), .ZN(new_n5854_));
  INV_X1     g05662(.I(new_n5685_), .ZN(new_n5855_));
  NOR3_X1    g05663(.A1(new_n5839_), .A2(\asqrt[48] ), .A3(new_n5841_), .ZN(new_n5856_));
  OAI21_X1   g05664(.A1(new_n5855_), .A2(new_n5856_), .B(new_n5842_), .ZN(new_n5857_));
  OAI21_X1   g05665(.A1(new_n5857_), .A2(\asqrt[49] ), .B(new_n5681_), .ZN(new_n5858_));
  NAND2_X1   g05666(.A1(new_n5857_), .A2(\asqrt[49] ), .ZN(new_n5859_));
  NAND3_X1   g05667(.A1(new_n5858_), .A2(new_n5859_), .A3(new_n1463_), .ZN(new_n5860_));
  AOI21_X1   g05668(.A1(new_n5858_), .A2(new_n5859_), .B(new_n1463_), .ZN(new_n5861_));
  AOI21_X1   g05669(.A1(new_n5678_), .A2(new_n5860_), .B(new_n5861_), .ZN(new_n5862_));
  AOI21_X1   g05670(.A1(new_n5862_), .A2(new_n1305_), .B(new_n5854_), .ZN(new_n5863_));
  NAND2_X1   g05671(.A1(new_n5860_), .A2(new_n5678_), .ZN(new_n5864_));
  AOI21_X1   g05672(.A1(new_n5864_), .A2(new_n5845_), .B(new_n1305_), .ZN(new_n5865_));
  OAI21_X1   g05673(.A1(new_n5863_), .A2(new_n5865_), .B(\asqrt[52] ), .ZN(new_n5866_));
  AOI21_X1   g05674(.A1(new_n5853_), .A2(new_n5866_), .B(new_n1006_), .ZN(new_n5867_));
  NOR3_X1    g05675(.A1(new_n5852_), .A2(\asqrt[54] ), .A3(new_n5867_), .ZN(new_n5868_));
  OAI21_X1   g05676(.A1(new_n5852_), .A2(new_n5867_), .B(\asqrt[54] ), .ZN(new_n5869_));
  OAI21_X1   g05677(.A1(new_n5667_), .A2(new_n5868_), .B(new_n5869_), .ZN(new_n5870_));
  OAI21_X1   g05678(.A1(new_n5870_), .A2(\asqrt[55] ), .B(new_n5664_), .ZN(new_n5871_));
  NAND2_X1   g05679(.A1(new_n5870_), .A2(\asqrt[55] ), .ZN(new_n5872_));
  NAND3_X1   g05680(.A1(new_n5871_), .A2(new_n5872_), .A3(new_n634_), .ZN(new_n5873_));
  AOI21_X1   g05681(.A1(new_n5871_), .A2(new_n5872_), .B(new_n634_), .ZN(new_n5874_));
  AOI21_X1   g05682(.A1(new_n5661_), .A2(new_n5873_), .B(new_n5874_), .ZN(new_n5875_));
  AOI21_X1   g05683(.A1(new_n5875_), .A2(new_n531_), .B(new_n5657_), .ZN(new_n5876_));
  NAND2_X1   g05684(.A1(new_n5873_), .A2(new_n5661_), .ZN(new_n5877_));
  INV_X1     g05685(.I(new_n5664_), .ZN(new_n5878_));
  INV_X1     g05686(.I(new_n5673_), .ZN(new_n5879_));
  NOR3_X1    g05687(.A1(new_n5863_), .A2(\asqrt[52] ), .A3(new_n5865_), .ZN(new_n5880_));
  OAI21_X1   g05688(.A1(new_n5879_), .A2(new_n5880_), .B(new_n5866_), .ZN(new_n5881_));
  OAI21_X1   g05689(.A1(new_n5881_), .A2(\asqrt[53] ), .B(new_n5669_), .ZN(new_n5882_));
  NAND2_X1   g05690(.A1(new_n5881_), .A2(\asqrt[53] ), .ZN(new_n5883_));
  NAND3_X1   g05691(.A1(new_n5882_), .A2(new_n5883_), .A3(new_n860_), .ZN(new_n5884_));
  AOI21_X1   g05692(.A1(new_n5882_), .A2(new_n5883_), .B(new_n860_), .ZN(new_n5885_));
  AOI21_X1   g05693(.A1(new_n5666_), .A2(new_n5884_), .B(new_n5885_), .ZN(new_n5886_));
  AOI21_X1   g05694(.A1(new_n5886_), .A2(new_n744_), .B(new_n5878_), .ZN(new_n5887_));
  NAND2_X1   g05695(.A1(new_n5884_), .A2(new_n5666_), .ZN(new_n5888_));
  AOI21_X1   g05696(.A1(new_n5888_), .A2(new_n5869_), .B(new_n744_), .ZN(new_n5889_));
  OAI21_X1   g05697(.A1(new_n5887_), .A2(new_n5889_), .B(\asqrt[56] ), .ZN(new_n5890_));
  AOI21_X1   g05698(.A1(new_n5877_), .A2(new_n5890_), .B(new_n531_), .ZN(new_n5891_));
  NOR3_X1    g05699(.A1(new_n5876_), .A2(\asqrt[58] ), .A3(new_n5891_), .ZN(new_n5892_));
  OAI21_X1   g05700(.A1(new_n5876_), .A2(new_n5891_), .B(\asqrt[58] ), .ZN(new_n5893_));
  OAI21_X1   g05701(.A1(new_n5654_), .A2(new_n5892_), .B(new_n5893_), .ZN(new_n5894_));
  OAI21_X1   g05702(.A1(new_n5894_), .A2(\asqrt[59] ), .B(new_n5651_), .ZN(new_n5895_));
  NAND2_X1   g05703(.A1(new_n5894_), .A2(\asqrt[59] ), .ZN(new_n5896_));
  NAND3_X1   g05704(.A1(new_n5895_), .A2(new_n5896_), .A3(new_n266_), .ZN(new_n5897_));
  NAND2_X1   g05705(.A1(new_n5897_), .A2(new_n5648_), .ZN(new_n5898_));
  INV_X1     g05706(.I(new_n5651_), .ZN(new_n5899_));
  INV_X1     g05707(.I(new_n5661_), .ZN(new_n5900_));
  NOR3_X1    g05708(.A1(new_n5887_), .A2(\asqrt[56] ), .A3(new_n5889_), .ZN(new_n5901_));
  OAI21_X1   g05709(.A1(new_n5900_), .A2(new_n5901_), .B(new_n5890_), .ZN(new_n5902_));
  OAI21_X1   g05710(.A1(new_n5902_), .A2(\asqrt[57] ), .B(new_n5656_), .ZN(new_n5903_));
  NOR2_X1    g05711(.A1(new_n5901_), .A2(new_n5900_), .ZN(new_n5904_));
  OAI21_X1   g05712(.A1(new_n5904_), .A2(new_n5874_), .B(\asqrt[57] ), .ZN(new_n5905_));
  NAND3_X1   g05713(.A1(new_n5903_), .A2(new_n423_), .A3(new_n5905_), .ZN(new_n5906_));
  AOI21_X1   g05714(.A1(new_n5903_), .A2(new_n5905_), .B(new_n423_), .ZN(new_n5907_));
  AOI21_X1   g05715(.A1(new_n5653_), .A2(new_n5906_), .B(new_n5907_), .ZN(new_n5908_));
  AOI21_X1   g05716(.A1(new_n5908_), .A2(new_n337_), .B(new_n5899_), .ZN(new_n5909_));
  NAND2_X1   g05717(.A1(new_n5906_), .A2(new_n5653_), .ZN(new_n5910_));
  AOI21_X1   g05718(.A1(new_n5910_), .A2(new_n5893_), .B(new_n337_), .ZN(new_n5911_));
  OAI21_X1   g05719(.A1(new_n5909_), .A2(new_n5911_), .B(\asqrt[60] ), .ZN(new_n5912_));
  AOI21_X1   g05720(.A1(new_n5898_), .A2(new_n5912_), .B(new_n239_), .ZN(new_n5913_));
  AOI21_X1   g05721(.A1(new_n5895_), .A2(new_n5896_), .B(new_n266_), .ZN(new_n5914_));
  AOI21_X1   g05722(.A1(new_n5648_), .A2(new_n5897_), .B(new_n5914_), .ZN(new_n5915_));
  AOI21_X1   g05723(.A1(new_n5598_), .A2(new_n5593_), .B(\asqrt[32] ), .ZN(new_n5916_));
  XOR2_X1    g05724(.A1(new_n5916_), .A2(new_n5342_), .Z(new_n5917_));
  INV_X1     g05725(.I(new_n5917_), .ZN(new_n5918_));
  AOI21_X1   g05726(.A1(new_n5915_), .A2(new_n239_), .B(new_n5918_), .ZN(new_n5919_));
  NOR2_X1    g05727(.A1(new_n5919_), .A2(new_n5913_), .ZN(new_n5920_));
  INV_X1     g05728(.I(new_n5648_), .ZN(new_n5921_));
  NAND3_X1   g05729(.A1(new_n5910_), .A2(new_n337_), .A3(new_n5893_), .ZN(new_n5922_));
  AOI21_X1   g05730(.A1(new_n5651_), .A2(new_n5922_), .B(new_n5911_), .ZN(new_n5923_));
  AOI21_X1   g05731(.A1(new_n5923_), .A2(new_n266_), .B(new_n5921_), .ZN(new_n5924_));
  OAI21_X1   g05732(.A1(new_n5924_), .A2(new_n5914_), .B(\asqrt[61] ), .ZN(new_n5925_));
  NOR3_X1    g05733(.A1(new_n5909_), .A2(\asqrt[60] ), .A3(new_n5911_), .ZN(new_n5926_));
  OAI21_X1   g05734(.A1(new_n5921_), .A2(new_n5926_), .B(new_n5912_), .ZN(new_n5927_));
  OAI21_X1   g05735(.A1(new_n5927_), .A2(\asqrt[61] ), .B(new_n5917_), .ZN(new_n5928_));
  AOI21_X1   g05736(.A1(new_n5928_), .A2(new_n5925_), .B(\asqrt[62] ), .ZN(new_n5929_));
  NOR3_X1    g05737(.A1(new_n5919_), .A2(new_n201_), .A3(new_n5913_), .ZN(new_n5930_));
  AOI21_X1   g05738(.A1(new_n5588_), .A2(new_n5594_), .B(\asqrt[32] ), .ZN(new_n5931_));
  XOR2_X1    g05739(.A1(new_n5931_), .A2(new_n5590_), .Z(new_n5932_));
  OAI22_X1   g05740(.A1(new_n5929_), .A2(new_n5930_), .B1(new_n5920_), .B2(new_n5932_), .ZN(new_n5933_));
  NOR2_X1    g05741(.A1(new_n5607_), .A2(new_n5339_), .ZN(new_n5934_));
  OAI21_X1   g05742(.A1(\asqrt[32] ), .A2(new_n5934_), .B(new_n5614_), .ZN(new_n5935_));
  AOI21_X1   g05743(.A1(new_n5933_), .A2(new_n5645_), .B(new_n5935_), .ZN(new_n5936_));
  INV_X1     g05744(.I(new_n5932_), .ZN(new_n5937_));
  AOI21_X1   g05745(.A1(new_n5920_), .A2(new_n201_), .B(new_n5937_), .ZN(new_n5938_));
  NOR2_X1    g05746(.A1(new_n5920_), .A2(new_n201_), .ZN(new_n5939_));
  NOR3_X1    g05747(.A1(new_n5938_), .A2(new_n5939_), .A3(new_n5645_), .ZN(new_n5940_));
  NAND2_X1   g05748(.A1(new_n5643_), .A2(new_n5338_), .ZN(new_n5941_));
  XOR2_X1    g05749(.A1(new_n5607_), .A2(new_n5339_), .Z(new_n5942_));
  NAND3_X1   g05750(.A1(new_n5941_), .A2(\asqrt[63] ), .A3(new_n5942_), .ZN(new_n5943_));
  INV_X1     g05751(.I(new_n5727_), .ZN(new_n5944_));
  NAND4_X1   g05752(.A1(new_n5944_), .A2(new_n5339_), .A3(new_n5614_), .A4(new_n5621_), .ZN(new_n5945_));
  NAND2_X1   g05753(.A1(new_n5943_), .A2(new_n5945_), .ZN(new_n5946_));
  NOR4_X1    g05754(.A1(new_n5936_), .A2(\asqrt[63] ), .A3(new_n5940_), .A4(new_n5946_), .ZN(new_n5947_));
  AOI21_X1   g05755(.A1(\asqrt[32] ), .A2(\a[64] ), .B(new_n5739_), .ZN(new_n5948_));
  OAI21_X1   g05756(.A1(new_n5631_), .A2(new_n5948_), .B(new_n5947_), .ZN(new_n5949_));
  XNOR2_X1   g05757(.A1(new_n5949_), .A2(new_n5626_), .ZN(new_n5950_));
  NAND3_X1   g05758(.A1(new_n5943_), .A2(\asqrt[32] ), .A3(new_n5945_), .ZN(new_n5951_));
  NOR4_X1    g05759(.A1(new_n5936_), .A2(\asqrt[63] ), .A3(new_n5940_), .A4(new_n5951_), .ZN(new_n5952_));
  INV_X1     g05760(.I(new_n5952_), .ZN(new_n5953_));
  INV_X1     g05761(.I(new_n5645_), .ZN(new_n5954_));
  NOR3_X1    g05762(.A1(new_n5924_), .A2(\asqrt[61] ), .A3(new_n5914_), .ZN(new_n5955_));
  OAI21_X1   g05763(.A1(new_n5918_), .A2(new_n5955_), .B(new_n5925_), .ZN(new_n5956_));
  OAI21_X1   g05764(.A1(new_n5919_), .A2(new_n5913_), .B(new_n201_), .ZN(new_n5957_));
  NAND3_X1   g05765(.A1(new_n5928_), .A2(\asqrt[62] ), .A3(new_n5925_), .ZN(new_n5958_));
  AOI22_X1   g05766(.A1(new_n5958_), .A2(new_n5957_), .B1(new_n5956_), .B2(new_n5937_), .ZN(new_n5959_));
  INV_X1     g05767(.I(new_n5935_), .ZN(new_n5960_));
  OAI21_X1   g05768(.A1(new_n5959_), .A2(new_n5954_), .B(new_n5960_), .ZN(new_n5961_));
  OAI21_X1   g05769(.A1(new_n5956_), .A2(\asqrt[62] ), .B(new_n5932_), .ZN(new_n5962_));
  NAND2_X1   g05770(.A1(new_n5956_), .A2(\asqrt[62] ), .ZN(new_n5963_));
  NAND3_X1   g05771(.A1(new_n5962_), .A2(new_n5963_), .A3(new_n5954_), .ZN(new_n5964_));
  INV_X1     g05772(.I(new_n5946_), .ZN(new_n5965_));
  NAND4_X1   g05773(.A1(new_n5961_), .A2(new_n193_), .A3(new_n5964_), .A4(new_n5965_), .ZN(\asqrt[31] ));
  NAND2_X1   g05774(.A1(\asqrt[31] ), .A2(new_n5627_), .ZN(new_n5967_));
  AOI21_X1   g05775(.A1(new_n5967_), .A2(new_n5953_), .B(\a[64] ), .ZN(new_n5968_));
  NOR2_X1    g05776(.A1(new_n5947_), .A2(new_n5628_), .ZN(new_n5969_));
  NOR3_X1    g05777(.A1(new_n5969_), .A2(new_n5623_), .A3(new_n5952_), .ZN(new_n5970_));
  NOR2_X1    g05778(.A1(new_n5970_), .A2(new_n5968_), .ZN(new_n5971_));
  INV_X1     g05779(.I(\a[62] ), .ZN(new_n5972_));
  NOR2_X1    g05780(.A1(\a[60] ), .A2(\a[61] ), .ZN(new_n5973_));
  NOR3_X1    g05781(.A1(new_n5947_), .A2(new_n5972_), .A3(new_n5973_), .ZN(new_n5974_));
  INV_X1     g05782(.I(new_n5973_), .ZN(new_n5975_));
  AOI21_X1   g05783(.A1(new_n5947_), .A2(\a[62] ), .B(new_n5975_), .ZN(new_n5976_));
  OAI21_X1   g05784(.A1(new_n5974_), .A2(new_n5976_), .B(\asqrt[32] ), .ZN(new_n5977_));
  NAND2_X1   g05785(.A1(new_n5973_), .A2(new_n5972_), .ZN(new_n5978_));
  NAND3_X1   g05786(.A1(new_n5617_), .A2(new_n5619_), .A3(new_n5978_), .ZN(new_n5979_));
  NAND2_X1   g05787(.A1(new_n5732_), .A2(new_n5979_), .ZN(new_n5980_));
  NAND3_X1   g05788(.A1(\asqrt[31] ), .A2(\a[62] ), .A3(new_n5980_), .ZN(new_n5981_));
  NOR3_X1    g05789(.A1(new_n5947_), .A2(\a[62] ), .A3(\a[63] ), .ZN(new_n5982_));
  INV_X1     g05790(.I(\a[63] ), .ZN(new_n5983_));
  AOI21_X1   g05791(.A1(\asqrt[31] ), .A2(new_n5972_), .B(new_n5983_), .ZN(new_n5984_));
  NOR2_X1    g05792(.A1(new_n5982_), .A2(new_n5984_), .ZN(new_n5985_));
  NAND4_X1   g05793(.A1(new_n5977_), .A2(new_n5985_), .A3(new_n5336_), .A4(new_n5981_), .ZN(new_n5986_));
  NAND2_X1   g05794(.A1(new_n5986_), .A2(new_n5971_), .ZN(new_n5987_));
  NAND3_X1   g05795(.A1(\asqrt[31] ), .A2(\a[62] ), .A3(new_n5975_), .ZN(new_n5988_));
  OAI21_X1   g05796(.A1(\asqrt[31] ), .A2(new_n5972_), .B(new_n5973_), .ZN(new_n5989_));
  AOI21_X1   g05797(.A1(new_n5989_), .A2(new_n5988_), .B(new_n5643_), .ZN(new_n5990_));
  NAND3_X1   g05798(.A1(\asqrt[31] ), .A2(new_n5972_), .A3(new_n5983_), .ZN(new_n5991_));
  OAI21_X1   g05799(.A1(new_n5947_), .A2(\a[62] ), .B(\a[63] ), .ZN(new_n5992_));
  NAND3_X1   g05800(.A1(new_n5981_), .A2(new_n5992_), .A3(new_n5991_), .ZN(new_n5993_));
  OAI21_X1   g05801(.A1(new_n5993_), .A2(new_n5990_), .B(\asqrt[33] ), .ZN(new_n5994_));
  NAND3_X1   g05802(.A1(new_n5987_), .A2(new_n5029_), .A3(new_n5994_), .ZN(new_n5995_));
  OR2_X2     g05803(.A1(new_n5970_), .A2(new_n5968_), .Z(new_n5996_));
  NOR3_X1    g05804(.A1(new_n5993_), .A2(new_n5990_), .A3(\asqrt[33] ), .ZN(new_n5997_));
  OAI21_X1   g05805(.A1(new_n5996_), .A2(new_n5997_), .B(new_n5994_), .ZN(new_n5998_));
  NAND2_X1   g05806(.A1(new_n5998_), .A2(\asqrt[34] ), .ZN(new_n5999_));
  NOR2_X1    g05807(.A1(new_n5956_), .A2(\asqrt[62] ), .ZN(new_n6000_));
  NOR2_X1    g05808(.A1(new_n6000_), .A2(new_n5939_), .ZN(new_n6001_));
  XOR2_X1    g05809(.A1(new_n5931_), .A2(new_n5590_), .Z(new_n6002_));
  OAI21_X1   g05810(.A1(\asqrt[31] ), .A2(new_n6001_), .B(new_n6002_), .ZN(new_n6003_));
  INV_X1     g05811(.I(new_n6003_), .ZN(new_n6004_));
  AOI21_X1   g05812(.A1(new_n5922_), .A2(new_n5896_), .B(\asqrt[31] ), .ZN(new_n6005_));
  XOR2_X1    g05813(.A1(new_n6005_), .A2(new_n5651_), .Z(new_n6006_));
  INV_X1     g05814(.I(new_n6006_), .ZN(new_n6007_));
  AOI21_X1   g05815(.A1(new_n5906_), .A2(new_n5893_), .B(\asqrt[31] ), .ZN(new_n6008_));
  XOR2_X1    g05816(.A1(new_n6008_), .A2(new_n5653_), .Z(new_n6009_));
  INV_X1     g05817(.I(new_n6009_), .ZN(new_n6010_));
  NAND2_X1   g05818(.A1(new_n5875_), .A2(new_n531_), .ZN(new_n6011_));
  AOI21_X1   g05819(.A1(new_n6011_), .A2(new_n5905_), .B(\asqrt[31] ), .ZN(new_n6012_));
  XOR2_X1    g05820(.A1(new_n6012_), .A2(new_n5656_), .Z(new_n6013_));
  AOI21_X1   g05821(.A1(new_n5873_), .A2(new_n5890_), .B(\asqrt[31] ), .ZN(new_n6014_));
  XOR2_X1    g05822(.A1(new_n6014_), .A2(new_n5661_), .Z(new_n6015_));
  NAND2_X1   g05823(.A1(new_n5886_), .A2(new_n744_), .ZN(new_n6016_));
  AOI21_X1   g05824(.A1(new_n6016_), .A2(new_n5872_), .B(\asqrt[31] ), .ZN(new_n6017_));
  XOR2_X1    g05825(.A1(new_n6017_), .A2(new_n5664_), .Z(new_n6018_));
  INV_X1     g05826(.I(new_n6018_), .ZN(new_n6019_));
  AOI21_X1   g05827(.A1(new_n5884_), .A2(new_n5869_), .B(\asqrt[31] ), .ZN(new_n6020_));
  XOR2_X1    g05828(.A1(new_n6020_), .A2(new_n5666_), .Z(new_n6021_));
  INV_X1     g05829(.I(new_n6021_), .ZN(new_n6022_));
  NAND2_X1   g05830(.A1(new_n5851_), .A2(new_n1006_), .ZN(new_n6023_));
  AOI21_X1   g05831(.A1(new_n6023_), .A2(new_n5883_), .B(\asqrt[31] ), .ZN(new_n6024_));
  XOR2_X1    g05832(.A1(new_n6024_), .A2(new_n5669_), .Z(new_n6025_));
  AOI21_X1   g05833(.A1(new_n5849_), .A2(new_n5866_), .B(\asqrt[31] ), .ZN(new_n6026_));
  XOR2_X1    g05834(.A1(new_n6026_), .A2(new_n5673_), .Z(new_n6027_));
  NAND2_X1   g05835(.A1(new_n5862_), .A2(new_n1305_), .ZN(new_n6028_));
  AOI21_X1   g05836(.A1(new_n6028_), .A2(new_n5848_), .B(\asqrt[31] ), .ZN(new_n6029_));
  XOR2_X1    g05837(.A1(new_n6029_), .A2(new_n5676_), .Z(new_n6030_));
  INV_X1     g05838(.I(new_n6030_), .ZN(new_n6031_));
  AOI21_X1   g05839(.A1(new_n5860_), .A2(new_n5845_), .B(\asqrt[31] ), .ZN(new_n6032_));
  XOR2_X1    g05840(.A1(new_n6032_), .A2(new_n5678_), .Z(new_n6033_));
  INV_X1     g05841(.I(new_n6033_), .ZN(new_n6034_));
  NAND2_X1   g05842(.A1(new_n5827_), .A2(new_n1632_), .ZN(new_n6035_));
  AOI21_X1   g05843(.A1(new_n6035_), .A2(new_n5859_), .B(\asqrt[31] ), .ZN(new_n6036_));
  XOR2_X1    g05844(.A1(new_n6036_), .A2(new_n5681_), .Z(new_n6037_));
  AOI21_X1   g05845(.A1(new_n5825_), .A2(new_n5842_), .B(\asqrt[31] ), .ZN(new_n6038_));
  XOR2_X1    g05846(.A1(new_n6038_), .A2(new_n5685_), .Z(new_n6039_));
  NAND2_X1   g05847(.A1(new_n5838_), .A2(new_n1953_), .ZN(new_n6040_));
  AOI21_X1   g05848(.A1(new_n6040_), .A2(new_n5824_), .B(\asqrt[31] ), .ZN(new_n6041_));
  XOR2_X1    g05849(.A1(new_n6041_), .A2(new_n5688_), .Z(new_n6042_));
  INV_X1     g05850(.I(new_n6042_), .ZN(new_n6043_));
  AOI21_X1   g05851(.A1(new_n5836_), .A2(new_n5821_), .B(\asqrt[31] ), .ZN(new_n6044_));
  XOR2_X1    g05852(.A1(new_n6044_), .A2(new_n5690_), .Z(new_n6045_));
  INV_X1     g05853(.I(new_n6045_), .ZN(new_n6046_));
  NAND2_X1   g05854(.A1(new_n5803_), .A2(new_n2332_), .ZN(new_n6047_));
  AOI21_X1   g05855(.A1(new_n6047_), .A2(new_n5835_), .B(\asqrt[31] ), .ZN(new_n6048_));
  XOR2_X1    g05856(.A1(new_n6048_), .A2(new_n5693_), .Z(new_n6049_));
  AOI21_X1   g05857(.A1(new_n5801_), .A2(new_n5818_), .B(\asqrt[31] ), .ZN(new_n6050_));
  XOR2_X1    g05858(.A1(new_n6050_), .A2(new_n5697_), .Z(new_n6051_));
  NAND2_X1   g05859(.A1(new_n5814_), .A2(new_n2749_), .ZN(new_n6052_));
  AOI21_X1   g05860(.A1(new_n6052_), .A2(new_n5800_), .B(\asqrt[31] ), .ZN(new_n6053_));
  XOR2_X1    g05861(.A1(new_n6053_), .A2(new_n5700_), .Z(new_n6054_));
  INV_X1     g05862(.I(new_n6054_), .ZN(new_n6055_));
  AOI21_X1   g05863(.A1(new_n5812_), .A2(new_n5797_), .B(\asqrt[31] ), .ZN(new_n6056_));
  XOR2_X1    g05864(.A1(new_n6056_), .A2(new_n5702_), .Z(new_n6057_));
  INV_X1     g05865(.I(new_n6057_), .ZN(new_n6058_));
  NAND2_X1   g05866(.A1(new_n5779_), .A2(new_n3195_), .ZN(new_n6059_));
  AOI21_X1   g05867(.A1(new_n6059_), .A2(new_n5811_), .B(\asqrt[31] ), .ZN(new_n6060_));
  XOR2_X1    g05868(.A1(new_n6060_), .A2(new_n5705_), .Z(new_n6061_));
  AOI21_X1   g05869(.A1(new_n5777_), .A2(new_n5794_), .B(\asqrt[31] ), .ZN(new_n6062_));
  XOR2_X1    g05870(.A1(new_n6062_), .A2(new_n5709_), .Z(new_n6063_));
  NAND2_X1   g05871(.A1(new_n5790_), .A2(new_n3681_), .ZN(new_n6064_));
  AOI21_X1   g05872(.A1(new_n6064_), .A2(new_n5776_), .B(\asqrt[31] ), .ZN(new_n6065_));
  XOR2_X1    g05873(.A1(new_n6065_), .A2(new_n5712_), .Z(new_n6066_));
  INV_X1     g05874(.I(new_n6066_), .ZN(new_n6067_));
  AOI21_X1   g05875(.A1(new_n5788_), .A2(new_n5773_), .B(\asqrt[31] ), .ZN(new_n6068_));
  XOR2_X1    g05876(.A1(new_n6068_), .A2(new_n5714_), .Z(new_n6069_));
  INV_X1     g05877(.I(new_n6069_), .ZN(new_n6070_));
  NAND2_X1   g05878(.A1(new_n5751_), .A2(new_n4196_), .ZN(new_n6071_));
  AOI21_X1   g05879(.A1(new_n6071_), .A2(new_n5787_), .B(\asqrt[31] ), .ZN(new_n6072_));
  XOR2_X1    g05880(.A1(new_n6072_), .A2(new_n5717_), .Z(new_n6073_));
  AOI21_X1   g05881(.A1(new_n5749_), .A2(new_n5770_), .B(\asqrt[31] ), .ZN(new_n6074_));
  XOR2_X1    g05882(.A1(new_n6074_), .A2(new_n5720_), .Z(new_n6075_));
  NAND2_X1   g05883(.A1(new_n5766_), .A2(new_n4751_), .ZN(new_n6076_));
  AOI21_X1   g05884(.A1(new_n6076_), .A2(new_n5748_), .B(\asqrt[31] ), .ZN(new_n6077_));
  XOR2_X1    g05885(.A1(new_n6077_), .A2(new_n5726_), .Z(new_n6078_));
  INV_X1     g05886(.I(new_n6078_), .ZN(new_n6079_));
  AOI21_X1   g05887(.A1(new_n5764_), .A2(new_n5745_), .B(\asqrt[31] ), .ZN(new_n6080_));
  XOR2_X1    g05888(.A1(new_n6080_), .A2(new_n5755_), .Z(new_n6081_));
  INV_X1     g05889(.I(new_n6081_), .ZN(new_n6082_));
  AOI21_X1   g05890(.A1(new_n5987_), .A2(new_n5994_), .B(new_n5029_), .ZN(new_n6083_));
  AOI21_X1   g05891(.A1(new_n5950_), .A2(new_n5995_), .B(new_n6083_), .ZN(new_n6084_));
  AOI21_X1   g05892(.A1(new_n6084_), .A2(new_n4751_), .B(new_n6082_), .ZN(new_n6085_));
  OAI21_X1   g05893(.A1(new_n5998_), .A2(\asqrt[34] ), .B(new_n5950_), .ZN(new_n6086_));
  AOI21_X1   g05894(.A1(new_n6086_), .A2(new_n5999_), .B(new_n4751_), .ZN(new_n6087_));
  NOR3_X1    g05895(.A1(new_n6085_), .A2(\asqrt[36] ), .A3(new_n6087_), .ZN(new_n6088_));
  OAI21_X1   g05896(.A1(new_n6085_), .A2(new_n6087_), .B(\asqrt[36] ), .ZN(new_n6089_));
  OAI21_X1   g05897(.A1(new_n6079_), .A2(new_n6088_), .B(new_n6089_), .ZN(new_n6090_));
  OAI21_X1   g05898(.A1(new_n6090_), .A2(\asqrt[37] ), .B(new_n6075_), .ZN(new_n6091_));
  NAND3_X1   g05899(.A1(new_n6086_), .A2(new_n5999_), .A3(new_n4751_), .ZN(new_n6092_));
  AOI21_X1   g05900(.A1(new_n6081_), .A2(new_n6092_), .B(new_n6087_), .ZN(new_n6093_));
  AOI21_X1   g05901(.A1(new_n6093_), .A2(new_n4461_), .B(new_n6079_), .ZN(new_n6094_));
  NAND2_X1   g05902(.A1(new_n6092_), .A2(new_n6081_), .ZN(new_n6095_));
  INV_X1     g05903(.I(new_n6087_), .ZN(new_n6096_));
  AOI21_X1   g05904(.A1(new_n6095_), .A2(new_n6096_), .B(new_n4461_), .ZN(new_n6097_));
  OAI21_X1   g05905(.A1(new_n6094_), .A2(new_n6097_), .B(\asqrt[37] ), .ZN(new_n6098_));
  NAND3_X1   g05906(.A1(new_n6091_), .A2(new_n3925_), .A3(new_n6098_), .ZN(new_n6099_));
  AOI21_X1   g05907(.A1(new_n6091_), .A2(new_n6098_), .B(new_n3925_), .ZN(new_n6100_));
  AOI21_X1   g05908(.A1(new_n6073_), .A2(new_n6099_), .B(new_n6100_), .ZN(new_n6101_));
  AOI21_X1   g05909(.A1(new_n6101_), .A2(new_n3681_), .B(new_n6070_), .ZN(new_n6102_));
  INV_X1     g05910(.I(new_n6075_), .ZN(new_n6103_));
  NOR3_X1    g05911(.A1(new_n6094_), .A2(\asqrt[37] ), .A3(new_n6097_), .ZN(new_n6104_));
  OAI21_X1   g05912(.A1(new_n6103_), .A2(new_n6104_), .B(new_n6098_), .ZN(new_n6105_));
  OAI21_X1   g05913(.A1(new_n6105_), .A2(\asqrt[38] ), .B(new_n6073_), .ZN(new_n6106_));
  NAND2_X1   g05914(.A1(new_n6105_), .A2(\asqrt[38] ), .ZN(new_n6107_));
  AOI21_X1   g05915(.A1(new_n6106_), .A2(new_n6107_), .B(new_n3681_), .ZN(new_n6108_));
  NOR3_X1    g05916(.A1(new_n6102_), .A2(\asqrt[40] ), .A3(new_n6108_), .ZN(new_n6109_));
  OAI21_X1   g05917(.A1(new_n6102_), .A2(new_n6108_), .B(\asqrt[40] ), .ZN(new_n6110_));
  OAI21_X1   g05918(.A1(new_n6067_), .A2(new_n6109_), .B(new_n6110_), .ZN(new_n6111_));
  OAI21_X1   g05919(.A1(new_n6111_), .A2(\asqrt[41] ), .B(new_n6063_), .ZN(new_n6112_));
  NAND3_X1   g05920(.A1(new_n6106_), .A2(new_n6107_), .A3(new_n3681_), .ZN(new_n6113_));
  AOI21_X1   g05921(.A1(new_n6069_), .A2(new_n6113_), .B(new_n6108_), .ZN(new_n6114_));
  AOI21_X1   g05922(.A1(new_n6114_), .A2(new_n3427_), .B(new_n6067_), .ZN(new_n6115_));
  NAND2_X1   g05923(.A1(new_n6113_), .A2(new_n6069_), .ZN(new_n6116_));
  INV_X1     g05924(.I(new_n6108_), .ZN(new_n6117_));
  AOI21_X1   g05925(.A1(new_n6116_), .A2(new_n6117_), .B(new_n3427_), .ZN(new_n6118_));
  OAI21_X1   g05926(.A1(new_n6115_), .A2(new_n6118_), .B(\asqrt[41] ), .ZN(new_n6119_));
  NAND3_X1   g05927(.A1(new_n6112_), .A2(new_n2960_), .A3(new_n6119_), .ZN(new_n6120_));
  AOI21_X1   g05928(.A1(new_n6112_), .A2(new_n6119_), .B(new_n2960_), .ZN(new_n6121_));
  AOI21_X1   g05929(.A1(new_n6061_), .A2(new_n6120_), .B(new_n6121_), .ZN(new_n6122_));
  AOI21_X1   g05930(.A1(new_n6122_), .A2(new_n2749_), .B(new_n6058_), .ZN(new_n6123_));
  INV_X1     g05931(.I(new_n6063_), .ZN(new_n6124_));
  NOR3_X1    g05932(.A1(new_n6115_), .A2(\asqrt[41] ), .A3(new_n6118_), .ZN(new_n6125_));
  OAI21_X1   g05933(.A1(new_n6124_), .A2(new_n6125_), .B(new_n6119_), .ZN(new_n6126_));
  OAI21_X1   g05934(.A1(new_n6126_), .A2(\asqrt[42] ), .B(new_n6061_), .ZN(new_n6127_));
  NAND2_X1   g05935(.A1(new_n6126_), .A2(\asqrt[42] ), .ZN(new_n6128_));
  AOI21_X1   g05936(.A1(new_n6127_), .A2(new_n6128_), .B(new_n2749_), .ZN(new_n6129_));
  NOR3_X1    g05937(.A1(new_n6123_), .A2(\asqrt[44] ), .A3(new_n6129_), .ZN(new_n6130_));
  OAI21_X1   g05938(.A1(new_n6123_), .A2(new_n6129_), .B(\asqrt[44] ), .ZN(new_n6131_));
  OAI21_X1   g05939(.A1(new_n6055_), .A2(new_n6130_), .B(new_n6131_), .ZN(new_n6132_));
  OAI21_X1   g05940(.A1(new_n6132_), .A2(\asqrt[45] ), .B(new_n6051_), .ZN(new_n6133_));
  NAND3_X1   g05941(.A1(new_n6127_), .A2(new_n6128_), .A3(new_n2749_), .ZN(new_n6134_));
  AOI21_X1   g05942(.A1(new_n6057_), .A2(new_n6134_), .B(new_n6129_), .ZN(new_n6135_));
  AOI21_X1   g05943(.A1(new_n6135_), .A2(new_n2531_), .B(new_n6055_), .ZN(new_n6136_));
  NAND2_X1   g05944(.A1(new_n6134_), .A2(new_n6057_), .ZN(new_n6137_));
  INV_X1     g05945(.I(new_n6129_), .ZN(new_n6138_));
  AOI21_X1   g05946(.A1(new_n6137_), .A2(new_n6138_), .B(new_n2531_), .ZN(new_n6139_));
  OAI21_X1   g05947(.A1(new_n6136_), .A2(new_n6139_), .B(\asqrt[45] ), .ZN(new_n6140_));
  NAND3_X1   g05948(.A1(new_n6133_), .A2(new_n2134_), .A3(new_n6140_), .ZN(new_n6141_));
  AOI21_X1   g05949(.A1(new_n6133_), .A2(new_n6140_), .B(new_n2134_), .ZN(new_n6142_));
  AOI21_X1   g05950(.A1(new_n6049_), .A2(new_n6141_), .B(new_n6142_), .ZN(new_n6143_));
  AOI21_X1   g05951(.A1(new_n6143_), .A2(new_n1953_), .B(new_n6046_), .ZN(new_n6144_));
  INV_X1     g05952(.I(new_n6051_), .ZN(new_n6145_));
  NOR3_X1    g05953(.A1(new_n6136_), .A2(\asqrt[45] ), .A3(new_n6139_), .ZN(new_n6146_));
  OAI21_X1   g05954(.A1(new_n6145_), .A2(new_n6146_), .B(new_n6140_), .ZN(new_n6147_));
  OAI21_X1   g05955(.A1(new_n6147_), .A2(\asqrt[46] ), .B(new_n6049_), .ZN(new_n6148_));
  NAND2_X1   g05956(.A1(new_n6147_), .A2(\asqrt[46] ), .ZN(new_n6149_));
  AOI21_X1   g05957(.A1(new_n6148_), .A2(new_n6149_), .B(new_n1953_), .ZN(new_n6150_));
  NOR3_X1    g05958(.A1(new_n6144_), .A2(\asqrt[48] ), .A3(new_n6150_), .ZN(new_n6151_));
  OAI21_X1   g05959(.A1(new_n6144_), .A2(new_n6150_), .B(\asqrt[48] ), .ZN(new_n6152_));
  OAI21_X1   g05960(.A1(new_n6043_), .A2(new_n6151_), .B(new_n6152_), .ZN(new_n6153_));
  OAI21_X1   g05961(.A1(new_n6153_), .A2(\asqrt[49] ), .B(new_n6039_), .ZN(new_n6154_));
  NAND3_X1   g05962(.A1(new_n6148_), .A2(new_n6149_), .A3(new_n1953_), .ZN(new_n6155_));
  AOI21_X1   g05963(.A1(new_n6045_), .A2(new_n6155_), .B(new_n6150_), .ZN(new_n6156_));
  AOI21_X1   g05964(.A1(new_n6156_), .A2(new_n1778_), .B(new_n6043_), .ZN(new_n6157_));
  NAND2_X1   g05965(.A1(new_n6155_), .A2(new_n6045_), .ZN(new_n6158_));
  INV_X1     g05966(.I(new_n6150_), .ZN(new_n6159_));
  AOI21_X1   g05967(.A1(new_n6158_), .A2(new_n6159_), .B(new_n1778_), .ZN(new_n6160_));
  OAI21_X1   g05968(.A1(new_n6157_), .A2(new_n6160_), .B(\asqrt[49] ), .ZN(new_n6161_));
  NAND3_X1   g05969(.A1(new_n6154_), .A2(new_n1463_), .A3(new_n6161_), .ZN(new_n6162_));
  AOI21_X1   g05970(.A1(new_n6154_), .A2(new_n6161_), .B(new_n1463_), .ZN(new_n6163_));
  AOI21_X1   g05971(.A1(new_n6037_), .A2(new_n6162_), .B(new_n6163_), .ZN(new_n6164_));
  AOI21_X1   g05972(.A1(new_n6164_), .A2(new_n1305_), .B(new_n6034_), .ZN(new_n6165_));
  INV_X1     g05973(.I(new_n6039_), .ZN(new_n6166_));
  NOR3_X1    g05974(.A1(new_n6157_), .A2(\asqrt[49] ), .A3(new_n6160_), .ZN(new_n6167_));
  OAI21_X1   g05975(.A1(new_n6166_), .A2(new_n6167_), .B(new_n6161_), .ZN(new_n6168_));
  OAI21_X1   g05976(.A1(new_n6168_), .A2(\asqrt[50] ), .B(new_n6037_), .ZN(new_n6169_));
  NAND2_X1   g05977(.A1(new_n6168_), .A2(\asqrt[50] ), .ZN(new_n6170_));
  AOI21_X1   g05978(.A1(new_n6169_), .A2(new_n6170_), .B(new_n1305_), .ZN(new_n6171_));
  NOR3_X1    g05979(.A1(new_n6165_), .A2(\asqrt[52] ), .A3(new_n6171_), .ZN(new_n6172_));
  OAI21_X1   g05980(.A1(new_n6165_), .A2(new_n6171_), .B(\asqrt[52] ), .ZN(new_n6173_));
  OAI21_X1   g05981(.A1(new_n6031_), .A2(new_n6172_), .B(new_n6173_), .ZN(new_n6174_));
  OAI21_X1   g05982(.A1(new_n6174_), .A2(\asqrt[53] ), .B(new_n6027_), .ZN(new_n6175_));
  NAND3_X1   g05983(.A1(new_n6169_), .A2(new_n6170_), .A3(new_n1305_), .ZN(new_n6176_));
  AOI21_X1   g05984(.A1(new_n6033_), .A2(new_n6176_), .B(new_n6171_), .ZN(new_n6177_));
  AOI21_X1   g05985(.A1(new_n6177_), .A2(new_n1150_), .B(new_n6031_), .ZN(new_n6178_));
  NAND2_X1   g05986(.A1(new_n6176_), .A2(new_n6033_), .ZN(new_n6179_));
  INV_X1     g05987(.I(new_n6171_), .ZN(new_n6180_));
  AOI21_X1   g05988(.A1(new_n6179_), .A2(new_n6180_), .B(new_n1150_), .ZN(new_n6181_));
  OAI21_X1   g05989(.A1(new_n6178_), .A2(new_n6181_), .B(\asqrt[53] ), .ZN(new_n6182_));
  NAND3_X1   g05990(.A1(new_n6175_), .A2(new_n860_), .A3(new_n6182_), .ZN(new_n6183_));
  AOI21_X1   g05991(.A1(new_n6175_), .A2(new_n6182_), .B(new_n860_), .ZN(new_n6184_));
  AOI21_X1   g05992(.A1(new_n6025_), .A2(new_n6183_), .B(new_n6184_), .ZN(new_n6185_));
  AOI21_X1   g05993(.A1(new_n6185_), .A2(new_n744_), .B(new_n6022_), .ZN(new_n6186_));
  INV_X1     g05994(.I(new_n6027_), .ZN(new_n6187_));
  NOR3_X1    g05995(.A1(new_n6178_), .A2(\asqrt[53] ), .A3(new_n6181_), .ZN(new_n6188_));
  OAI21_X1   g05996(.A1(new_n6187_), .A2(new_n6188_), .B(new_n6182_), .ZN(new_n6189_));
  OAI21_X1   g05997(.A1(new_n6189_), .A2(\asqrt[54] ), .B(new_n6025_), .ZN(new_n6190_));
  NAND2_X1   g05998(.A1(new_n6189_), .A2(\asqrt[54] ), .ZN(new_n6191_));
  AOI21_X1   g05999(.A1(new_n6190_), .A2(new_n6191_), .B(new_n744_), .ZN(new_n6192_));
  NOR3_X1    g06000(.A1(new_n6186_), .A2(\asqrt[56] ), .A3(new_n6192_), .ZN(new_n6193_));
  OAI21_X1   g06001(.A1(new_n6186_), .A2(new_n6192_), .B(\asqrt[56] ), .ZN(new_n6194_));
  OAI21_X1   g06002(.A1(new_n6019_), .A2(new_n6193_), .B(new_n6194_), .ZN(new_n6195_));
  OAI21_X1   g06003(.A1(new_n6195_), .A2(\asqrt[57] ), .B(new_n6015_), .ZN(new_n6196_));
  NAND3_X1   g06004(.A1(new_n6190_), .A2(new_n6191_), .A3(new_n744_), .ZN(new_n6197_));
  AOI21_X1   g06005(.A1(new_n6021_), .A2(new_n6197_), .B(new_n6192_), .ZN(new_n6198_));
  AOI21_X1   g06006(.A1(new_n6198_), .A2(new_n634_), .B(new_n6019_), .ZN(new_n6199_));
  NAND2_X1   g06007(.A1(new_n6197_), .A2(new_n6021_), .ZN(new_n6200_));
  INV_X1     g06008(.I(new_n6192_), .ZN(new_n6201_));
  AOI21_X1   g06009(.A1(new_n6200_), .A2(new_n6201_), .B(new_n634_), .ZN(new_n6202_));
  OAI21_X1   g06010(.A1(new_n6199_), .A2(new_n6202_), .B(\asqrt[57] ), .ZN(new_n6203_));
  NAND3_X1   g06011(.A1(new_n6196_), .A2(new_n423_), .A3(new_n6203_), .ZN(new_n6204_));
  AOI21_X1   g06012(.A1(new_n6196_), .A2(new_n6203_), .B(new_n423_), .ZN(new_n6205_));
  AOI21_X1   g06013(.A1(new_n6013_), .A2(new_n6204_), .B(new_n6205_), .ZN(new_n6206_));
  AOI21_X1   g06014(.A1(new_n6206_), .A2(new_n337_), .B(new_n6010_), .ZN(new_n6207_));
  NOR2_X1    g06015(.A1(new_n6206_), .A2(new_n337_), .ZN(new_n6208_));
  NOR3_X1    g06016(.A1(new_n6207_), .A2(new_n6208_), .A3(\asqrt[60] ), .ZN(new_n6209_));
  OAI21_X1   g06017(.A1(new_n6207_), .A2(new_n6208_), .B(\asqrt[60] ), .ZN(new_n6210_));
  OAI21_X1   g06018(.A1(new_n6007_), .A2(new_n6209_), .B(new_n6210_), .ZN(new_n6211_));
  NAND2_X1   g06019(.A1(new_n6211_), .A2(\asqrt[61] ), .ZN(new_n6212_));
  AOI21_X1   g06020(.A1(new_n5897_), .A2(new_n5912_), .B(\asqrt[31] ), .ZN(new_n6213_));
  XOR2_X1    g06021(.A1(new_n6213_), .A2(new_n5648_), .Z(new_n6214_));
  OAI21_X1   g06022(.A1(new_n6211_), .A2(\asqrt[61] ), .B(new_n6214_), .ZN(new_n6215_));
  NAND2_X1   g06023(.A1(new_n6215_), .A2(new_n6212_), .ZN(new_n6216_));
  INV_X1     g06024(.I(new_n6015_), .ZN(new_n6217_));
  NOR3_X1    g06025(.A1(new_n6199_), .A2(\asqrt[57] ), .A3(new_n6202_), .ZN(new_n6218_));
  OAI21_X1   g06026(.A1(new_n6217_), .A2(new_n6218_), .B(new_n6203_), .ZN(new_n6219_));
  OAI21_X1   g06027(.A1(new_n6219_), .A2(\asqrt[58] ), .B(new_n6013_), .ZN(new_n6220_));
  NOR2_X1    g06028(.A1(new_n6218_), .A2(new_n6217_), .ZN(new_n6221_));
  INV_X1     g06029(.I(new_n6203_), .ZN(new_n6222_));
  OAI21_X1   g06030(.A1(new_n6221_), .A2(new_n6222_), .B(\asqrt[58] ), .ZN(new_n6223_));
  NAND3_X1   g06031(.A1(new_n6220_), .A2(new_n337_), .A3(new_n6223_), .ZN(new_n6224_));
  NAND2_X1   g06032(.A1(new_n6224_), .A2(new_n6009_), .ZN(new_n6225_));
  INV_X1     g06033(.I(new_n6013_), .ZN(new_n6226_));
  NOR2_X1    g06034(.A1(new_n6221_), .A2(new_n6222_), .ZN(new_n6227_));
  AOI21_X1   g06035(.A1(new_n6227_), .A2(new_n423_), .B(new_n6226_), .ZN(new_n6228_));
  OAI21_X1   g06036(.A1(new_n6228_), .A2(new_n6205_), .B(\asqrt[59] ), .ZN(new_n6229_));
  NAND3_X1   g06037(.A1(new_n6225_), .A2(new_n266_), .A3(new_n6229_), .ZN(new_n6230_));
  NAND2_X1   g06038(.A1(new_n6230_), .A2(new_n6006_), .ZN(new_n6231_));
  AOI21_X1   g06039(.A1(new_n6231_), .A2(new_n6210_), .B(new_n239_), .ZN(new_n6232_));
  AOI21_X1   g06040(.A1(new_n6225_), .A2(new_n6229_), .B(new_n266_), .ZN(new_n6233_));
  AOI21_X1   g06041(.A1(new_n6006_), .A2(new_n6230_), .B(new_n6233_), .ZN(new_n6234_));
  INV_X1     g06042(.I(new_n6214_), .ZN(new_n6235_));
  AOI21_X1   g06043(.A1(new_n6234_), .A2(new_n239_), .B(new_n6235_), .ZN(new_n6236_));
  OAI21_X1   g06044(.A1(new_n6236_), .A2(new_n6232_), .B(new_n201_), .ZN(new_n6237_));
  NAND3_X1   g06045(.A1(new_n6215_), .A2(new_n6212_), .A3(\asqrt[62] ), .ZN(new_n6238_));
  NOR2_X1    g06046(.A1(new_n5955_), .A2(new_n5913_), .ZN(new_n6239_));
  NOR2_X1    g06047(.A1(\asqrt[31] ), .A2(new_n6239_), .ZN(new_n6240_));
  XOR2_X1    g06048(.A1(new_n6240_), .A2(new_n5917_), .Z(new_n6241_));
  INV_X1     g06049(.I(new_n6241_), .ZN(new_n6242_));
  AOI22_X1   g06050(.A1(new_n6238_), .A2(new_n6237_), .B1(new_n6216_), .B2(new_n6242_), .ZN(new_n6243_));
  NOR2_X1    g06051(.A1(new_n5959_), .A2(new_n5954_), .ZN(new_n6244_));
  OAI21_X1   g06052(.A1(\asqrt[31] ), .A2(new_n6244_), .B(new_n5964_), .ZN(new_n6245_));
  INV_X1     g06053(.I(new_n6245_), .ZN(new_n6246_));
  OAI21_X1   g06054(.A1(new_n6243_), .A2(new_n6004_), .B(new_n6246_), .ZN(new_n6247_));
  OAI21_X1   g06055(.A1(new_n6216_), .A2(\asqrt[62] ), .B(new_n6241_), .ZN(new_n6248_));
  NAND2_X1   g06056(.A1(new_n6216_), .A2(\asqrt[62] ), .ZN(new_n6249_));
  NAND3_X1   g06057(.A1(new_n6248_), .A2(new_n6249_), .A3(new_n6004_), .ZN(new_n6250_));
  NAND2_X1   g06058(.A1(new_n5959_), .A2(new_n5645_), .ZN(new_n6251_));
  NAND2_X1   g06059(.A1(new_n5933_), .A2(new_n5954_), .ZN(new_n6252_));
  AOI21_X1   g06060(.A1(new_n6251_), .A2(new_n6252_), .B(new_n193_), .ZN(new_n6253_));
  OAI21_X1   g06061(.A1(\asqrt[31] ), .A2(new_n5954_), .B(new_n6253_), .ZN(new_n6254_));
  NOR2_X1    g06062(.A1(new_n5946_), .A2(new_n5645_), .ZN(new_n6255_));
  NAND4_X1   g06063(.A1(new_n5961_), .A2(new_n193_), .A3(new_n5964_), .A4(new_n6255_), .ZN(new_n6256_));
  NAND2_X1   g06064(.A1(new_n6254_), .A2(new_n6256_), .ZN(new_n6257_));
  INV_X1     g06065(.I(new_n6257_), .ZN(new_n6258_));
  NAND4_X1   g06066(.A1(new_n6247_), .A2(new_n193_), .A3(new_n6250_), .A4(new_n6258_), .ZN(\asqrt[30] ));
  AOI21_X1   g06067(.A1(new_n5995_), .A2(new_n5999_), .B(\asqrt[30] ), .ZN(new_n6260_));
  XOR2_X1    g06068(.A1(new_n6260_), .A2(new_n5950_), .Z(new_n6261_));
  AOI21_X1   g06069(.A1(new_n5986_), .A2(new_n5994_), .B(\asqrt[30] ), .ZN(new_n6262_));
  XOR2_X1    g06070(.A1(new_n6262_), .A2(new_n5971_), .Z(new_n6263_));
  NAND2_X1   g06071(.A1(\asqrt[31] ), .A2(new_n5972_), .ZN(new_n6264_));
  NOR2_X1    g06072(.A1(new_n5983_), .A2(\a[62] ), .ZN(new_n6265_));
  AOI22_X1   g06073(.A1(new_n6264_), .A2(new_n5983_), .B1(\asqrt[31] ), .B2(new_n6265_), .ZN(new_n6266_));
  NOR2_X1    g06074(.A1(new_n6236_), .A2(new_n6232_), .ZN(new_n6267_));
  AOI21_X1   g06075(.A1(new_n6215_), .A2(new_n6212_), .B(\asqrt[62] ), .ZN(new_n6268_));
  NOR3_X1    g06076(.A1(new_n6236_), .A2(new_n201_), .A3(new_n6232_), .ZN(new_n6269_));
  OAI22_X1   g06077(.A1(new_n6268_), .A2(new_n6269_), .B1(new_n6267_), .B2(new_n6241_), .ZN(new_n6270_));
  AOI21_X1   g06078(.A1(new_n6270_), .A2(new_n6003_), .B(new_n6245_), .ZN(new_n6271_));
  AOI21_X1   g06079(.A1(new_n6267_), .A2(new_n201_), .B(new_n6242_), .ZN(new_n6272_));
  NOR2_X1    g06080(.A1(new_n6267_), .A2(new_n201_), .ZN(new_n6273_));
  NOR3_X1    g06081(.A1(new_n6272_), .A2(new_n6273_), .A3(new_n6003_), .ZN(new_n6274_));
  NOR4_X1    g06082(.A1(new_n6271_), .A2(\asqrt[63] ), .A3(new_n6274_), .A4(new_n6257_), .ZN(new_n6275_));
  AOI21_X1   g06083(.A1(\asqrt[31] ), .A2(\a[62] ), .B(new_n5980_), .ZN(new_n6276_));
  OAI21_X1   g06084(.A1(new_n5990_), .A2(new_n6276_), .B(new_n6275_), .ZN(new_n6277_));
  XNOR2_X1   g06085(.A1(new_n6277_), .A2(new_n6266_), .ZN(new_n6278_));
  NOR3_X1    g06086(.A1(new_n6271_), .A2(\asqrt[63] ), .A3(new_n6274_), .ZN(new_n6279_));
  NAND4_X1   g06087(.A1(new_n6279_), .A2(\asqrt[31] ), .A3(new_n6254_), .A4(new_n6256_), .ZN(new_n6280_));
  NAND2_X1   g06088(.A1(\asqrt[30] ), .A2(new_n5973_), .ZN(new_n6281_));
  AOI21_X1   g06089(.A1(new_n6280_), .A2(new_n6281_), .B(\a[62] ), .ZN(new_n6282_));
  NAND2_X1   g06090(.A1(new_n6247_), .A2(new_n193_), .ZN(new_n6283_));
  NAND3_X1   g06091(.A1(new_n6254_), .A2(new_n6256_), .A3(\asqrt[31] ), .ZN(new_n6284_));
  NOR3_X1    g06092(.A1(new_n6283_), .A2(new_n6274_), .A3(new_n6284_), .ZN(new_n6285_));
  NOR2_X1    g06093(.A1(new_n6275_), .A2(new_n5975_), .ZN(new_n6286_));
  NOR3_X1    g06094(.A1(new_n6286_), .A2(new_n6285_), .A3(new_n5972_), .ZN(new_n6287_));
  OR2_X2     g06095(.A1(new_n6282_), .A2(new_n6287_), .Z(new_n6288_));
  NOR2_X1    g06096(.A1(\a[58] ), .A2(\a[59] ), .ZN(new_n6289_));
  INV_X1     g06097(.I(new_n6289_), .ZN(new_n6290_));
  NAND3_X1   g06098(.A1(\asqrt[30] ), .A2(\a[60] ), .A3(new_n6290_), .ZN(new_n6291_));
  INV_X1     g06099(.I(\a[60] ), .ZN(new_n6292_));
  OAI21_X1   g06100(.A1(\asqrt[30] ), .A2(new_n6292_), .B(new_n6289_), .ZN(new_n6293_));
  AOI21_X1   g06101(.A1(new_n6293_), .A2(new_n6291_), .B(new_n5947_), .ZN(new_n6294_));
  NOR3_X1    g06102(.A1(new_n5936_), .A2(\asqrt[63] ), .A3(new_n5940_), .ZN(new_n6295_));
  NAND2_X1   g06103(.A1(new_n6289_), .A2(new_n6292_), .ZN(new_n6296_));
  NAND3_X1   g06104(.A1(new_n5943_), .A2(new_n5945_), .A3(new_n6296_), .ZN(new_n6297_));
  NAND2_X1   g06105(.A1(new_n6295_), .A2(new_n6297_), .ZN(new_n6298_));
  NAND3_X1   g06106(.A1(\asqrt[30] ), .A2(\a[60] ), .A3(new_n6298_), .ZN(new_n6299_));
  INV_X1     g06107(.I(\a[61] ), .ZN(new_n6300_));
  NAND3_X1   g06108(.A1(\asqrt[30] ), .A2(new_n6292_), .A3(new_n6300_), .ZN(new_n6301_));
  OAI21_X1   g06109(.A1(new_n6275_), .A2(\a[60] ), .B(\a[61] ), .ZN(new_n6302_));
  NAND3_X1   g06110(.A1(new_n6299_), .A2(new_n6302_), .A3(new_n6301_), .ZN(new_n6303_));
  NOR3_X1    g06111(.A1(new_n6303_), .A2(new_n6294_), .A3(\asqrt[32] ), .ZN(new_n6304_));
  OAI21_X1   g06112(.A1(new_n6303_), .A2(new_n6294_), .B(\asqrt[32] ), .ZN(new_n6305_));
  OAI21_X1   g06113(.A1(new_n6288_), .A2(new_n6304_), .B(new_n6305_), .ZN(new_n6306_));
  OAI21_X1   g06114(.A1(new_n6306_), .A2(\asqrt[33] ), .B(new_n6278_), .ZN(new_n6307_));
  NAND2_X1   g06115(.A1(new_n6306_), .A2(\asqrt[33] ), .ZN(new_n6308_));
  NAND3_X1   g06116(.A1(new_n6307_), .A2(new_n6308_), .A3(new_n5029_), .ZN(new_n6309_));
  AOI21_X1   g06117(.A1(new_n6307_), .A2(new_n6308_), .B(new_n5029_), .ZN(new_n6310_));
  AOI21_X1   g06118(.A1(new_n6263_), .A2(new_n6309_), .B(new_n6310_), .ZN(new_n6311_));
  NAND2_X1   g06119(.A1(new_n6311_), .A2(new_n4751_), .ZN(new_n6312_));
  INV_X1     g06120(.I(new_n6263_), .ZN(new_n6313_));
  INV_X1     g06121(.I(new_n6278_), .ZN(new_n6314_));
  NOR2_X1    g06122(.A1(new_n6282_), .A2(new_n6287_), .ZN(new_n6315_));
  NOR3_X1    g06123(.A1(new_n6275_), .A2(new_n6292_), .A3(new_n6289_), .ZN(new_n6316_));
  AOI21_X1   g06124(.A1(new_n6275_), .A2(\a[60] ), .B(new_n6290_), .ZN(new_n6317_));
  OAI21_X1   g06125(.A1(new_n6316_), .A2(new_n6317_), .B(\asqrt[31] ), .ZN(new_n6318_));
  INV_X1     g06126(.I(new_n6298_), .ZN(new_n6319_));
  NOR3_X1    g06127(.A1(new_n6275_), .A2(new_n6292_), .A3(new_n6319_), .ZN(new_n6320_));
  NOR3_X1    g06128(.A1(new_n6275_), .A2(\a[60] ), .A3(\a[61] ), .ZN(new_n6321_));
  AOI21_X1   g06129(.A1(\asqrt[30] ), .A2(new_n6292_), .B(new_n6300_), .ZN(new_n6322_));
  NOR3_X1    g06130(.A1(new_n6320_), .A2(new_n6321_), .A3(new_n6322_), .ZN(new_n6323_));
  NAND3_X1   g06131(.A1(new_n6323_), .A2(new_n6318_), .A3(new_n5643_), .ZN(new_n6324_));
  AOI21_X1   g06132(.A1(new_n6323_), .A2(new_n6318_), .B(new_n5643_), .ZN(new_n6325_));
  AOI21_X1   g06133(.A1(new_n6315_), .A2(new_n6324_), .B(new_n6325_), .ZN(new_n6326_));
  AOI21_X1   g06134(.A1(new_n6326_), .A2(new_n5336_), .B(new_n6314_), .ZN(new_n6327_));
  NAND2_X1   g06135(.A1(new_n6324_), .A2(new_n6315_), .ZN(new_n6328_));
  AOI21_X1   g06136(.A1(new_n6328_), .A2(new_n6305_), .B(new_n5336_), .ZN(new_n6329_));
  NOR3_X1    g06137(.A1(new_n6327_), .A2(\asqrt[34] ), .A3(new_n6329_), .ZN(new_n6330_));
  OAI21_X1   g06138(.A1(new_n6327_), .A2(new_n6329_), .B(\asqrt[34] ), .ZN(new_n6331_));
  OAI21_X1   g06139(.A1(new_n6313_), .A2(new_n6330_), .B(new_n6331_), .ZN(new_n6332_));
  NAND2_X1   g06140(.A1(new_n6332_), .A2(\asqrt[35] ), .ZN(new_n6333_));
  NOR2_X1    g06141(.A1(new_n6216_), .A2(\asqrt[62] ), .ZN(new_n6334_));
  NOR2_X1    g06142(.A1(new_n6334_), .A2(new_n6273_), .ZN(new_n6335_));
  XOR2_X1    g06143(.A1(new_n6240_), .A2(new_n5917_), .Z(new_n6336_));
  OAI21_X1   g06144(.A1(\asqrt[30] ), .A2(new_n6335_), .B(new_n6336_), .ZN(new_n6337_));
  INV_X1     g06145(.I(new_n6337_), .ZN(new_n6338_));
  AOI21_X1   g06146(.A1(new_n6224_), .A2(new_n6229_), .B(\asqrt[30] ), .ZN(new_n6339_));
  XOR2_X1    g06147(.A1(new_n6339_), .A2(new_n6009_), .Z(new_n6340_));
  INV_X1     g06148(.I(new_n6340_), .ZN(new_n6341_));
  AOI21_X1   g06149(.A1(new_n6204_), .A2(new_n6223_), .B(\asqrt[30] ), .ZN(new_n6342_));
  XOR2_X1    g06150(.A1(new_n6342_), .A2(new_n6013_), .Z(new_n6343_));
  INV_X1     g06151(.I(new_n6343_), .ZN(new_n6344_));
  NOR2_X1    g06152(.A1(new_n6222_), .A2(new_n6218_), .ZN(new_n6345_));
  NOR2_X1    g06153(.A1(\asqrt[30] ), .A2(new_n6345_), .ZN(new_n6346_));
  XOR2_X1    g06154(.A1(new_n6346_), .A2(new_n6015_), .Z(new_n6347_));
  NOR2_X1    g06155(.A1(new_n6193_), .A2(new_n6202_), .ZN(new_n6348_));
  NOR2_X1    g06156(.A1(\asqrt[30] ), .A2(new_n6348_), .ZN(new_n6349_));
  XOR2_X1    g06157(.A1(new_n6349_), .A2(new_n6018_), .Z(new_n6350_));
  AOI21_X1   g06158(.A1(new_n6197_), .A2(new_n6201_), .B(\asqrt[30] ), .ZN(new_n6351_));
  XOR2_X1    g06159(.A1(new_n6351_), .A2(new_n6021_), .Z(new_n6352_));
  INV_X1     g06160(.I(new_n6352_), .ZN(new_n6353_));
  AOI21_X1   g06161(.A1(new_n6183_), .A2(new_n6191_), .B(\asqrt[30] ), .ZN(new_n6354_));
  XOR2_X1    g06162(.A1(new_n6354_), .A2(new_n6025_), .Z(new_n6355_));
  INV_X1     g06163(.I(new_n6355_), .ZN(new_n6356_));
  XOR2_X1    g06164(.A1(new_n6174_), .A2(\asqrt[53] ), .Z(new_n6357_));
  NOR2_X1    g06165(.A1(\asqrt[30] ), .A2(new_n6357_), .ZN(new_n6358_));
  XOR2_X1    g06166(.A1(new_n6358_), .A2(new_n6027_), .Z(new_n6359_));
  NOR2_X1    g06167(.A1(new_n6172_), .A2(new_n6181_), .ZN(new_n6360_));
  NOR2_X1    g06168(.A1(\asqrt[30] ), .A2(new_n6360_), .ZN(new_n6361_));
  XOR2_X1    g06169(.A1(new_n6361_), .A2(new_n6030_), .Z(new_n6362_));
  AOI21_X1   g06170(.A1(new_n6176_), .A2(new_n6180_), .B(\asqrt[30] ), .ZN(new_n6363_));
  XOR2_X1    g06171(.A1(new_n6363_), .A2(new_n6033_), .Z(new_n6364_));
  INV_X1     g06172(.I(new_n6364_), .ZN(new_n6365_));
  AOI21_X1   g06173(.A1(new_n6162_), .A2(new_n6170_), .B(\asqrt[30] ), .ZN(new_n6366_));
  XOR2_X1    g06174(.A1(new_n6366_), .A2(new_n6037_), .Z(new_n6367_));
  INV_X1     g06175(.I(new_n6367_), .ZN(new_n6368_));
  XOR2_X1    g06176(.A1(new_n6153_), .A2(\asqrt[49] ), .Z(new_n6369_));
  NOR2_X1    g06177(.A1(\asqrt[30] ), .A2(new_n6369_), .ZN(new_n6370_));
  XOR2_X1    g06178(.A1(new_n6370_), .A2(new_n6039_), .Z(new_n6371_));
  NOR2_X1    g06179(.A1(new_n6151_), .A2(new_n6160_), .ZN(new_n6372_));
  NOR2_X1    g06180(.A1(\asqrt[30] ), .A2(new_n6372_), .ZN(new_n6373_));
  XOR2_X1    g06181(.A1(new_n6373_), .A2(new_n6042_), .Z(new_n6374_));
  AOI21_X1   g06182(.A1(new_n6155_), .A2(new_n6159_), .B(\asqrt[30] ), .ZN(new_n6375_));
  XOR2_X1    g06183(.A1(new_n6375_), .A2(new_n6045_), .Z(new_n6376_));
  INV_X1     g06184(.I(new_n6376_), .ZN(new_n6377_));
  AOI21_X1   g06185(.A1(new_n6141_), .A2(new_n6149_), .B(\asqrt[30] ), .ZN(new_n6378_));
  XOR2_X1    g06186(.A1(new_n6378_), .A2(new_n6049_), .Z(new_n6379_));
  INV_X1     g06187(.I(new_n6379_), .ZN(new_n6380_));
  XOR2_X1    g06188(.A1(new_n6132_), .A2(\asqrt[45] ), .Z(new_n6381_));
  NOR2_X1    g06189(.A1(\asqrt[30] ), .A2(new_n6381_), .ZN(new_n6382_));
  XOR2_X1    g06190(.A1(new_n6382_), .A2(new_n6051_), .Z(new_n6383_));
  NOR2_X1    g06191(.A1(new_n6130_), .A2(new_n6139_), .ZN(new_n6384_));
  NOR2_X1    g06192(.A1(\asqrt[30] ), .A2(new_n6384_), .ZN(new_n6385_));
  XOR2_X1    g06193(.A1(new_n6385_), .A2(new_n6054_), .Z(new_n6386_));
  AOI21_X1   g06194(.A1(new_n6134_), .A2(new_n6138_), .B(\asqrt[30] ), .ZN(new_n6387_));
  XOR2_X1    g06195(.A1(new_n6387_), .A2(new_n6057_), .Z(new_n6388_));
  INV_X1     g06196(.I(new_n6388_), .ZN(new_n6389_));
  AOI21_X1   g06197(.A1(new_n6120_), .A2(new_n6128_), .B(\asqrt[30] ), .ZN(new_n6390_));
  XOR2_X1    g06198(.A1(new_n6390_), .A2(new_n6061_), .Z(new_n6391_));
  INV_X1     g06199(.I(new_n6391_), .ZN(new_n6392_));
  XOR2_X1    g06200(.A1(new_n6111_), .A2(\asqrt[41] ), .Z(new_n6393_));
  NOR2_X1    g06201(.A1(\asqrt[30] ), .A2(new_n6393_), .ZN(new_n6394_));
  XOR2_X1    g06202(.A1(new_n6394_), .A2(new_n6063_), .Z(new_n6395_));
  NOR2_X1    g06203(.A1(new_n6109_), .A2(new_n6118_), .ZN(new_n6396_));
  NOR2_X1    g06204(.A1(\asqrt[30] ), .A2(new_n6396_), .ZN(new_n6397_));
  XOR2_X1    g06205(.A1(new_n6397_), .A2(new_n6066_), .Z(new_n6398_));
  AOI21_X1   g06206(.A1(new_n6113_), .A2(new_n6117_), .B(\asqrt[30] ), .ZN(new_n6399_));
  XOR2_X1    g06207(.A1(new_n6399_), .A2(new_n6069_), .Z(new_n6400_));
  INV_X1     g06208(.I(new_n6400_), .ZN(new_n6401_));
  AOI21_X1   g06209(.A1(new_n6099_), .A2(new_n6107_), .B(\asqrt[30] ), .ZN(new_n6402_));
  XOR2_X1    g06210(.A1(new_n6402_), .A2(new_n6073_), .Z(new_n6403_));
  INV_X1     g06211(.I(new_n6403_), .ZN(new_n6404_));
  XOR2_X1    g06212(.A1(new_n6090_), .A2(\asqrt[37] ), .Z(new_n6405_));
  NOR2_X1    g06213(.A1(\asqrt[30] ), .A2(new_n6405_), .ZN(new_n6406_));
  XOR2_X1    g06214(.A1(new_n6406_), .A2(new_n6075_), .Z(new_n6407_));
  NOR2_X1    g06215(.A1(new_n6088_), .A2(new_n6097_), .ZN(new_n6408_));
  NOR2_X1    g06216(.A1(\asqrt[30] ), .A2(new_n6408_), .ZN(new_n6409_));
  XOR2_X1    g06217(.A1(new_n6409_), .A2(new_n6078_), .Z(new_n6410_));
  AOI21_X1   g06218(.A1(new_n6092_), .A2(new_n6096_), .B(\asqrt[30] ), .ZN(new_n6411_));
  XOR2_X1    g06219(.A1(new_n6411_), .A2(new_n6081_), .Z(new_n6412_));
  INV_X1     g06220(.I(new_n6412_), .ZN(new_n6413_));
  INV_X1     g06221(.I(new_n6261_), .ZN(new_n6414_));
  AOI21_X1   g06222(.A1(new_n6311_), .A2(new_n4751_), .B(new_n6414_), .ZN(new_n6415_));
  NAND2_X1   g06223(.A1(new_n6309_), .A2(new_n6263_), .ZN(new_n6416_));
  AOI21_X1   g06224(.A1(new_n6416_), .A2(new_n6331_), .B(new_n4751_), .ZN(new_n6417_));
  NOR3_X1    g06225(.A1(new_n6415_), .A2(\asqrt[36] ), .A3(new_n6417_), .ZN(new_n6418_));
  OAI21_X1   g06226(.A1(new_n6415_), .A2(new_n6417_), .B(\asqrt[36] ), .ZN(new_n6419_));
  OAI21_X1   g06227(.A1(new_n6413_), .A2(new_n6418_), .B(new_n6419_), .ZN(new_n6420_));
  OAI21_X1   g06228(.A1(new_n6420_), .A2(\asqrt[37] ), .B(new_n6410_), .ZN(new_n6421_));
  NAND2_X1   g06229(.A1(new_n6420_), .A2(\asqrt[37] ), .ZN(new_n6422_));
  NAND3_X1   g06230(.A1(new_n6421_), .A2(new_n6422_), .A3(new_n3925_), .ZN(new_n6423_));
  AOI21_X1   g06231(.A1(new_n6421_), .A2(new_n6422_), .B(new_n3925_), .ZN(new_n6424_));
  AOI21_X1   g06232(.A1(new_n6407_), .A2(new_n6423_), .B(new_n6424_), .ZN(new_n6425_));
  AOI21_X1   g06233(.A1(new_n6425_), .A2(new_n3681_), .B(new_n6404_), .ZN(new_n6426_));
  NAND2_X1   g06234(.A1(new_n6423_), .A2(new_n6407_), .ZN(new_n6427_));
  INV_X1     g06235(.I(new_n6410_), .ZN(new_n6428_));
  OAI21_X1   g06236(.A1(new_n6332_), .A2(\asqrt[35] ), .B(new_n6261_), .ZN(new_n6429_));
  NAND3_X1   g06237(.A1(new_n6429_), .A2(new_n6333_), .A3(new_n4461_), .ZN(new_n6430_));
  AOI21_X1   g06238(.A1(new_n6429_), .A2(new_n6333_), .B(new_n4461_), .ZN(new_n6431_));
  AOI21_X1   g06239(.A1(new_n6412_), .A2(new_n6430_), .B(new_n6431_), .ZN(new_n6432_));
  AOI21_X1   g06240(.A1(new_n6432_), .A2(new_n4196_), .B(new_n6428_), .ZN(new_n6433_));
  NAND2_X1   g06241(.A1(new_n6430_), .A2(new_n6412_), .ZN(new_n6434_));
  AOI21_X1   g06242(.A1(new_n6434_), .A2(new_n6419_), .B(new_n4196_), .ZN(new_n6435_));
  OAI21_X1   g06243(.A1(new_n6433_), .A2(new_n6435_), .B(\asqrt[38] ), .ZN(new_n6436_));
  AOI21_X1   g06244(.A1(new_n6427_), .A2(new_n6436_), .B(new_n3681_), .ZN(new_n6437_));
  NOR3_X1    g06245(.A1(new_n6426_), .A2(\asqrt[40] ), .A3(new_n6437_), .ZN(new_n6438_));
  OAI21_X1   g06246(.A1(new_n6426_), .A2(new_n6437_), .B(\asqrt[40] ), .ZN(new_n6439_));
  OAI21_X1   g06247(.A1(new_n6401_), .A2(new_n6438_), .B(new_n6439_), .ZN(new_n6440_));
  OAI21_X1   g06248(.A1(new_n6440_), .A2(\asqrt[41] ), .B(new_n6398_), .ZN(new_n6441_));
  NAND2_X1   g06249(.A1(new_n6440_), .A2(\asqrt[41] ), .ZN(new_n6442_));
  NAND3_X1   g06250(.A1(new_n6441_), .A2(new_n6442_), .A3(new_n2960_), .ZN(new_n6443_));
  AOI21_X1   g06251(.A1(new_n6441_), .A2(new_n6442_), .B(new_n2960_), .ZN(new_n6444_));
  AOI21_X1   g06252(.A1(new_n6395_), .A2(new_n6443_), .B(new_n6444_), .ZN(new_n6445_));
  AOI21_X1   g06253(.A1(new_n6445_), .A2(new_n2749_), .B(new_n6392_), .ZN(new_n6446_));
  NAND2_X1   g06254(.A1(new_n6443_), .A2(new_n6395_), .ZN(new_n6447_));
  INV_X1     g06255(.I(new_n6398_), .ZN(new_n6448_));
  INV_X1     g06256(.I(new_n6407_), .ZN(new_n6449_));
  NOR3_X1    g06257(.A1(new_n6433_), .A2(\asqrt[38] ), .A3(new_n6435_), .ZN(new_n6450_));
  OAI21_X1   g06258(.A1(new_n6449_), .A2(new_n6450_), .B(new_n6436_), .ZN(new_n6451_));
  OAI21_X1   g06259(.A1(new_n6451_), .A2(\asqrt[39] ), .B(new_n6403_), .ZN(new_n6452_));
  NAND2_X1   g06260(.A1(new_n6451_), .A2(\asqrt[39] ), .ZN(new_n6453_));
  NAND3_X1   g06261(.A1(new_n6452_), .A2(new_n6453_), .A3(new_n3427_), .ZN(new_n6454_));
  AOI21_X1   g06262(.A1(new_n6452_), .A2(new_n6453_), .B(new_n3427_), .ZN(new_n6455_));
  AOI21_X1   g06263(.A1(new_n6400_), .A2(new_n6454_), .B(new_n6455_), .ZN(new_n6456_));
  AOI21_X1   g06264(.A1(new_n6456_), .A2(new_n3195_), .B(new_n6448_), .ZN(new_n6457_));
  NAND2_X1   g06265(.A1(new_n6454_), .A2(new_n6400_), .ZN(new_n6458_));
  AOI21_X1   g06266(.A1(new_n6458_), .A2(new_n6439_), .B(new_n3195_), .ZN(new_n6459_));
  OAI21_X1   g06267(.A1(new_n6457_), .A2(new_n6459_), .B(\asqrt[42] ), .ZN(new_n6460_));
  AOI21_X1   g06268(.A1(new_n6447_), .A2(new_n6460_), .B(new_n2749_), .ZN(new_n6461_));
  NOR3_X1    g06269(.A1(new_n6446_), .A2(\asqrt[44] ), .A3(new_n6461_), .ZN(new_n6462_));
  OAI21_X1   g06270(.A1(new_n6446_), .A2(new_n6461_), .B(\asqrt[44] ), .ZN(new_n6463_));
  OAI21_X1   g06271(.A1(new_n6389_), .A2(new_n6462_), .B(new_n6463_), .ZN(new_n6464_));
  OAI21_X1   g06272(.A1(new_n6464_), .A2(\asqrt[45] ), .B(new_n6386_), .ZN(new_n6465_));
  NAND2_X1   g06273(.A1(new_n6464_), .A2(\asqrt[45] ), .ZN(new_n6466_));
  NAND3_X1   g06274(.A1(new_n6465_), .A2(new_n6466_), .A3(new_n2134_), .ZN(new_n6467_));
  AOI21_X1   g06275(.A1(new_n6465_), .A2(new_n6466_), .B(new_n2134_), .ZN(new_n6468_));
  AOI21_X1   g06276(.A1(new_n6383_), .A2(new_n6467_), .B(new_n6468_), .ZN(new_n6469_));
  AOI21_X1   g06277(.A1(new_n6469_), .A2(new_n1953_), .B(new_n6380_), .ZN(new_n6470_));
  NAND2_X1   g06278(.A1(new_n6467_), .A2(new_n6383_), .ZN(new_n6471_));
  INV_X1     g06279(.I(new_n6386_), .ZN(new_n6472_));
  INV_X1     g06280(.I(new_n6395_), .ZN(new_n6473_));
  NOR3_X1    g06281(.A1(new_n6457_), .A2(\asqrt[42] ), .A3(new_n6459_), .ZN(new_n6474_));
  OAI21_X1   g06282(.A1(new_n6473_), .A2(new_n6474_), .B(new_n6460_), .ZN(new_n6475_));
  OAI21_X1   g06283(.A1(new_n6475_), .A2(\asqrt[43] ), .B(new_n6391_), .ZN(new_n6476_));
  NAND2_X1   g06284(.A1(new_n6475_), .A2(\asqrt[43] ), .ZN(new_n6477_));
  NAND3_X1   g06285(.A1(new_n6476_), .A2(new_n6477_), .A3(new_n2531_), .ZN(new_n6478_));
  AOI21_X1   g06286(.A1(new_n6476_), .A2(new_n6477_), .B(new_n2531_), .ZN(new_n6479_));
  AOI21_X1   g06287(.A1(new_n6388_), .A2(new_n6478_), .B(new_n6479_), .ZN(new_n6480_));
  AOI21_X1   g06288(.A1(new_n6480_), .A2(new_n2332_), .B(new_n6472_), .ZN(new_n6481_));
  NAND2_X1   g06289(.A1(new_n6478_), .A2(new_n6388_), .ZN(new_n6482_));
  AOI21_X1   g06290(.A1(new_n6482_), .A2(new_n6463_), .B(new_n2332_), .ZN(new_n6483_));
  OAI21_X1   g06291(.A1(new_n6481_), .A2(new_n6483_), .B(\asqrt[46] ), .ZN(new_n6484_));
  AOI21_X1   g06292(.A1(new_n6471_), .A2(new_n6484_), .B(new_n1953_), .ZN(new_n6485_));
  NOR3_X1    g06293(.A1(new_n6470_), .A2(\asqrt[48] ), .A3(new_n6485_), .ZN(new_n6486_));
  OAI21_X1   g06294(.A1(new_n6470_), .A2(new_n6485_), .B(\asqrt[48] ), .ZN(new_n6487_));
  OAI21_X1   g06295(.A1(new_n6377_), .A2(new_n6486_), .B(new_n6487_), .ZN(new_n6488_));
  OAI21_X1   g06296(.A1(new_n6488_), .A2(\asqrt[49] ), .B(new_n6374_), .ZN(new_n6489_));
  NAND2_X1   g06297(.A1(new_n6488_), .A2(\asqrt[49] ), .ZN(new_n6490_));
  NAND3_X1   g06298(.A1(new_n6489_), .A2(new_n6490_), .A3(new_n1463_), .ZN(new_n6491_));
  AOI21_X1   g06299(.A1(new_n6489_), .A2(new_n6490_), .B(new_n1463_), .ZN(new_n6492_));
  AOI21_X1   g06300(.A1(new_n6371_), .A2(new_n6491_), .B(new_n6492_), .ZN(new_n6493_));
  AOI21_X1   g06301(.A1(new_n6493_), .A2(new_n1305_), .B(new_n6368_), .ZN(new_n6494_));
  NAND2_X1   g06302(.A1(new_n6491_), .A2(new_n6371_), .ZN(new_n6495_));
  INV_X1     g06303(.I(new_n6374_), .ZN(new_n6496_));
  INV_X1     g06304(.I(new_n6383_), .ZN(new_n6497_));
  NOR3_X1    g06305(.A1(new_n6481_), .A2(\asqrt[46] ), .A3(new_n6483_), .ZN(new_n6498_));
  OAI21_X1   g06306(.A1(new_n6497_), .A2(new_n6498_), .B(new_n6484_), .ZN(new_n6499_));
  OAI21_X1   g06307(.A1(new_n6499_), .A2(\asqrt[47] ), .B(new_n6379_), .ZN(new_n6500_));
  NAND2_X1   g06308(.A1(new_n6499_), .A2(\asqrt[47] ), .ZN(new_n6501_));
  NAND3_X1   g06309(.A1(new_n6500_), .A2(new_n6501_), .A3(new_n1778_), .ZN(new_n6502_));
  AOI21_X1   g06310(.A1(new_n6500_), .A2(new_n6501_), .B(new_n1778_), .ZN(new_n6503_));
  AOI21_X1   g06311(.A1(new_n6376_), .A2(new_n6502_), .B(new_n6503_), .ZN(new_n6504_));
  AOI21_X1   g06312(.A1(new_n6504_), .A2(new_n1632_), .B(new_n6496_), .ZN(new_n6505_));
  NAND2_X1   g06313(.A1(new_n6502_), .A2(new_n6376_), .ZN(new_n6506_));
  AOI21_X1   g06314(.A1(new_n6506_), .A2(new_n6487_), .B(new_n1632_), .ZN(new_n6507_));
  OAI21_X1   g06315(.A1(new_n6505_), .A2(new_n6507_), .B(\asqrt[50] ), .ZN(new_n6508_));
  AOI21_X1   g06316(.A1(new_n6495_), .A2(new_n6508_), .B(new_n1305_), .ZN(new_n6509_));
  NOR3_X1    g06317(.A1(new_n6494_), .A2(\asqrt[52] ), .A3(new_n6509_), .ZN(new_n6510_));
  OAI21_X1   g06318(.A1(new_n6494_), .A2(new_n6509_), .B(\asqrt[52] ), .ZN(new_n6511_));
  OAI21_X1   g06319(.A1(new_n6365_), .A2(new_n6510_), .B(new_n6511_), .ZN(new_n6512_));
  OAI21_X1   g06320(.A1(new_n6512_), .A2(\asqrt[53] ), .B(new_n6362_), .ZN(new_n6513_));
  NAND2_X1   g06321(.A1(new_n6512_), .A2(\asqrt[53] ), .ZN(new_n6514_));
  NAND3_X1   g06322(.A1(new_n6513_), .A2(new_n6514_), .A3(new_n860_), .ZN(new_n6515_));
  AOI21_X1   g06323(.A1(new_n6513_), .A2(new_n6514_), .B(new_n860_), .ZN(new_n6516_));
  AOI21_X1   g06324(.A1(new_n6359_), .A2(new_n6515_), .B(new_n6516_), .ZN(new_n6517_));
  AOI21_X1   g06325(.A1(new_n6517_), .A2(new_n744_), .B(new_n6356_), .ZN(new_n6518_));
  NAND2_X1   g06326(.A1(new_n6515_), .A2(new_n6359_), .ZN(new_n6519_));
  INV_X1     g06327(.I(new_n6362_), .ZN(new_n6520_));
  INV_X1     g06328(.I(new_n6371_), .ZN(new_n6521_));
  NOR3_X1    g06329(.A1(new_n6505_), .A2(\asqrt[50] ), .A3(new_n6507_), .ZN(new_n6522_));
  OAI21_X1   g06330(.A1(new_n6521_), .A2(new_n6522_), .B(new_n6508_), .ZN(new_n6523_));
  OAI21_X1   g06331(.A1(new_n6523_), .A2(\asqrt[51] ), .B(new_n6367_), .ZN(new_n6524_));
  NAND2_X1   g06332(.A1(new_n6523_), .A2(\asqrt[51] ), .ZN(new_n6525_));
  NAND3_X1   g06333(.A1(new_n6524_), .A2(new_n6525_), .A3(new_n1150_), .ZN(new_n6526_));
  AOI21_X1   g06334(.A1(new_n6524_), .A2(new_n6525_), .B(new_n1150_), .ZN(new_n6527_));
  AOI21_X1   g06335(.A1(new_n6364_), .A2(new_n6526_), .B(new_n6527_), .ZN(new_n6528_));
  AOI21_X1   g06336(.A1(new_n6528_), .A2(new_n1006_), .B(new_n6520_), .ZN(new_n6529_));
  NAND2_X1   g06337(.A1(new_n6526_), .A2(new_n6364_), .ZN(new_n6530_));
  AOI21_X1   g06338(.A1(new_n6530_), .A2(new_n6511_), .B(new_n1006_), .ZN(new_n6531_));
  OAI21_X1   g06339(.A1(new_n6529_), .A2(new_n6531_), .B(\asqrt[54] ), .ZN(new_n6532_));
  AOI21_X1   g06340(.A1(new_n6519_), .A2(new_n6532_), .B(new_n744_), .ZN(new_n6533_));
  NOR3_X1    g06341(.A1(new_n6518_), .A2(\asqrt[56] ), .A3(new_n6533_), .ZN(new_n6534_));
  OAI21_X1   g06342(.A1(new_n6518_), .A2(new_n6533_), .B(\asqrt[56] ), .ZN(new_n6535_));
  OAI21_X1   g06343(.A1(new_n6353_), .A2(new_n6534_), .B(new_n6535_), .ZN(new_n6536_));
  OAI21_X1   g06344(.A1(new_n6536_), .A2(\asqrt[57] ), .B(new_n6350_), .ZN(new_n6537_));
  NAND2_X1   g06345(.A1(new_n6536_), .A2(\asqrt[57] ), .ZN(new_n6538_));
  NAND3_X1   g06346(.A1(new_n6537_), .A2(new_n6538_), .A3(new_n423_), .ZN(new_n6539_));
  AOI21_X1   g06347(.A1(new_n6537_), .A2(new_n6538_), .B(new_n423_), .ZN(new_n6540_));
  AOI21_X1   g06348(.A1(new_n6347_), .A2(new_n6539_), .B(new_n6540_), .ZN(new_n6541_));
  AOI21_X1   g06349(.A1(new_n6541_), .A2(new_n337_), .B(new_n6344_), .ZN(new_n6542_));
  NAND2_X1   g06350(.A1(new_n6539_), .A2(new_n6347_), .ZN(new_n6543_));
  INV_X1     g06351(.I(new_n6350_), .ZN(new_n6544_));
  INV_X1     g06352(.I(new_n6359_), .ZN(new_n6545_));
  NOR3_X1    g06353(.A1(new_n6529_), .A2(\asqrt[54] ), .A3(new_n6531_), .ZN(new_n6546_));
  OAI21_X1   g06354(.A1(new_n6545_), .A2(new_n6546_), .B(new_n6532_), .ZN(new_n6547_));
  OAI21_X1   g06355(.A1(new_n6547_), .A2(\asqrt[55] ), .B(new_n6355_), .ZN(new_n6548_));
  NAND2_X1   g06356(.A1(new_n6547_), .A2(\asqrt[55] ), .ZN(new_n6549_));
  NAND3_X1   g06357(.A1(new_n6548_), .A2(new_n6549_), .A3(new_n634_), .ZN(new_n6550_));
  AOI21_X1   g06358(.A1(new_n6548_), .A2(new_n6549_), .B(new_n634_), .ZN(new_n6551_));
  AOI21_X1   g06359(.A1(new_n6352_), .A2(new_n6550_), .B(new_n6551_), .ZN(new_n6552_));
  AOI21_X1   g06360(.A1(new_n6552_), .A2(new_n531_), .B(new_n6544_), .ZN(new_n6553_));
  NAND2_X1   g06361(.A1(new_n6550_), .A2(new_n6352_), .ZN(new_n6554_));
  AOI21_X1   g06362(.A1(new_n6554_), .A2(new_n6535_), .B(new_n531_), .ZN(new_n6555_));
  OAI21_X1   g06363(.A1(new_n6553_), .A2(new_n6555_), .B(\asqrt[58] ), .ZN(new_n6556_));
  AOI21_X1   g06364(.A1(new_n6543_), .A2(new_n6556_), .B(new_n337_), .ZN(new_n6557_));
  NOR3_X1    g06365(.A1(new_n6542_), .A2(\asqrt[60] ), .A3(new_n6557_), .ZN(new_n6558_));
  NOR2_X1    g06366(.A1(new_n6558_), .A2(new_n6341_), .ZN(new_n6559_));
  INV_X1     g06367(.I(new_n6347_), .ZN(new_n6560_));
  NOR3_X1    g06368(.A1(new_n6553_), .A2(\asqrt[58] ), .A3(new_n6555_), .ZN(new_n6561_));
  OAI21_X1   g06369(.A1(new_n6560_), .A2(new_n6561_), .B(new_n6556_), .ZN(new_n6562_));
  OAI21_X1   g06370(.A1(new_n6562_), .A2(\asqrt[59] ), .B(new_n6343_), .ZN(new_n6563_));
  NOR2_X1    g06371(.A1(new_n6561_), .A2(new_n6560_), .ZN(new_n6564_));
  OAI21_X1   g06372(.A1(new_n6564_), .A2(new_n6540_), .B(\asqrt[59] ), .ZN(new_n6565_));
  AOI21_X1   g06373(.A1(new_n6563_), .A2(new_n6565_), .B(new_n266_), .ZN(new_n6566_));
  OAI21_X1   g06374(.A1(new_n6559_), .A2(new_n6566_), .B(\asqrt[61] ), .ZN(new_n6567_));
  OAI21_X1   g06375(.A1(new_n6542_), .A2(new_n6557_), .B(\asqrt[60] ), .ZN(new_n6568_));
  OAI21_X1   g06376(.A1(new_n6341_), .A2(new_n6558_), .B(new_n6568_), .ZN(new_n6569_));
  AOI21_X1   g06377(.A1(new_n6230_), .A2(new_n6210_), .B(\asqrt[30] ), .ZN(new_n6570_));
  XOR2_X1    g06378(.A1(new_n6570_), .A2(new_n6006_), .Z(new_n6571_));
  OAI21_X1   g06379(.A1(new_n6569_), .A2(\asqrt[61] ), .B(new_n6571_), .ZN(new_n6572_));
  NAND2_X1   g06380(.A1(new_n6572_), .A2(new_n6567_), .ZN(new_n6573_));
  NAND3_X1   g06381(.A1(new_n6563_), .A2(new_n266_), .A3(new_n6565_), .ZN(new_n6574_));
  NAND2_X1   g06382(.A1(new_n6574_), .A2(new_n6340_), .ZN(new_n6575_));
  AOI21_X1   g06383(.A1(new_n6575_), .A2(new_n6568_), .B(new_n239_), .ZN(new_n6576_));
  AOI21_X1   g06384(.A1(new_n6340_), .A2(new_n6574_), .B(new_n6566_), .ZN(new_n6577_));
  INV_X1     g06385(.I(new_n6571_), .ZN(new_n6578_));
  AOI21_X1   g06386(.A1(new_n6577_), .A2(new_n239_), .B(new_n6578_), .ZN(new_n6579_));
  OAI21_X1   g06387(.A1(new_n6579_), .A2(new_n6576_), .B(new_n201_), .ZN(new_n6580_));
  NAND3_X1   g06388(.A1(new_n6572_), .A2(\asqrt[62] ), .A3(new_n6567_), .ZN(new_n6581_));
  NAND2_X1   g06389(.A1(new_n6234_), .A2(new_n239_), .ZN(new_n6582_));
  AOI21_X1   g06390(.A1(new_n6212_), .A2(new_n6582_), .B(\asqrt[30] ), .ZN(new_n6583_));
  XOR2_X1    g06391(.A1(new_n6583_), .A2(new_n6214_), .Z(new_n6584_));
  INV_X1     g06392(.I(new_n6584_), .ZN(new_n6585_));
  AOI22_X1   g06393(.A1(new_n6580_), .A2(new_n6581_), .B1(new_n6573_), .B2(new_n6585_), .ZN(new_n6586_));
  NOR2_X1    g06394(.A1(new_n6243_), .A2(new_n6004_), .ZN(new_n6587_));
  OAI21_X1   g06395(.A1(\asqrt[30] ), .A2(new_n6587_), .B(new_n6250_), .ZN(new_n6588_));
  INV_X1     g06396(.I(new_n6588_), .ZN(new_n6589_));
  OAI21_X1   g06397(.A1(new_n6586_), .A2(new_n6338_), .B(new_n6589_), .ZN(new_n6590_));
  OAI21_X1   g06398(.A1(new_n6573_), .A2(\asqrt[62] ), .B(new_n6584_), .ZN(new_n6591_));
  NAND2_X1   g06399(.A1(new_n6573_), .A2(\asqrt[62] ), .ZN(new_n6592_));
  NAND3_X1   g06400(.A1(new_n6591_), .A2(new_n6592_), .A3(new_n6338_), .ZN(new_n6593_));
  NAND2_X1   g06401(.A1(new_n6275_), .A2(new_n6003_), .ZN(new_n6594_));
  XOR2_X1    g06402(.A1(new_n6270_), .A2(new_n6003_), .Z(new_n6595_));
  NAND3_X1   g06403(.A1(new_n6594_), .A2(\asqrt[63] ), .A3(new_n6595_), .ZN(new_n6596_));
  INV_X1     g06404(.I(new_n6283_), .ZN(new_n6597_));
  NAND4_X1   g06405(.A1(new_n6597_), .A2(new_n6004_), .A3(new_n6250_), .A4(new_n6258_), .ZN(new_n6598_));
  NAND2_X1   g06406(.A1(new_n6596_), .A2(new_n6598_), .ZN(new_n6599_));
  INV_X1     g06407(.I(new_n6599_), .ZN(new_n6600_));
  NAND4_X1   g06408(.A1(new_n6590_), .A2(new_n193_), .A3(new_n6593_), .A4(new_n6600_), .ZN(\asqrt[29] ));
  AOI21_X1   g06409(.A1(new_n6312_), .A2(new_n6333_), .B(\asqrt[29] ), .ZN(new_n6602_));
  XOR2_X1    g06410(.A1(new_n6602_), .A2(new_n6261_), .Z(new_n6603_));
  AOI21_X1   g06411(.A1(new_n6309_), .A2(new_n6331_), .B(\asqrt[29] ), .ZN(new_n6604_));
  XOR2_X1    g06412(.A1(new_n6604_), .A2(new_n6263_), .Z(new_n6605_));
  NAND2_X1   g06413(.A1(new_n6326_), .A2(new_n5336_), .ZN(new_n6606_));
  AOI21_X1   g06414(.A1(new_n6606_), .A2(new_n6308_), .B(\asqrt[29] ), .ZN(new_n6607_));
  XOR2_X1    g06415(.A1(new_n6607_), .A2(new_n6278_), .Z(new_n6608_));
  INV_X1     g06416(.I(new_n6608_), .ZN(new_n6609_));
  AOI21_X1   g06417(.A1(new_n6324_), .A2(new_n6305_), .B(\asqrt[29] ), .ZN(new_n6610_));
  XOR2_X1    g06418(.A1(new_n6610_), .A2(new_n6315_), .Z(new_n6611_));
  INV_X1     g06419(.I(new_n6611_), .ZN(new_n6612_));
  NAND2_X1   g06420(.A1(\asqrt[30] ), .A2(new_n6292_), .ZN(new_n6613_));
  NOR2_X1    g06421(.A1(new_n6300_), .A2(\a[60] ), .ZN(new_n6614_));
  AOI22_X1   g06422(.A1(new_n6613_), .A2(new_n6300_), .B1(\asqrt[30] ), .B2(new_n6614_), .ZN(new_n6615_));
  OAI21_X1   g06423(.A1(new_n6275_), .A2(new_n6292_), .B(new_n6319_), .ZN(new_n6616_));
  AOI21_X1   g06424(.A1(new_n6318_), .A2(new_n6616_), .B(\asqrt[29] ), .ZN(new_n6617_));
  XOR2_X1    g06425(.A1(new_n6617_), .A2(new_n6615_), .Z(new_n6618_));
  NAND3_X1   g06426(.A1(new_n6575_), .A2(new_n239_), .A3(new_n6568_), .ZN(new_n6619_));
  AOI21_X1   g06427(.A1(new_n6571_), .A2(new_n6619_), .B(new_n6576_), .ZN(new_n6620_));
  AOI21_X1   g06428(.A1(new_n6572_), .A2(new_n6567_), .B(\asqrt[62] ), .ZN(new_n6621_));
  NOR3_X1    g06429(.A1(new_n6579_), .A2(new_n201_), .A3(new_n6576_), .ZN(new_n6622_));
  OAI22_X1   g06430(.A1(new_n6622_), .A2(new_n6621_), .B1(new_n6620_), .B2(new_n6584_), .ZN(new_n6623_));
  AOI21_X1   g06431(.A1(new_n6623_), .A2(new_n6337_), .B(new_n6588_), .ZN(new_n6624_));
  AOI21_X1   g06432(.A1(new_n6620_), .A2(new_n201_), .B(new_n6585_), .ZN(new_n6625_));
  OAI21_X1   g06433(.A1(new_n6620_), .A2(new_n201_), .B(new_n6338_), .ZN(new_n6626_));
  NOR2_X1    g06434(.A1(new_n6625_), .A2(new_n6626_), .ZN(new_n6627_));
  NOR3_X1    g06435(.A1(new_n6624_), .A2(\asqrt[63] ), .A3(new_n6627_), .ZN(new_n6628_));
  NAND3_X1   g06436(.A1(new_n6596_), .A2(\asqrt[30] ), .A3(new_n6598_), .ZN(new_n6629_));
  INV_X1     g06437(.I(new_n6629_), .ZN(new_n6630_));
  NAND2_X1   g06438(.A1(new_n6628_), .A2(new_n6630_), .ZN(new_n6631_));
  NAND2_X1   g06439(.A1(\asqrt[29] ), .A2(new_n6289_), .ZN(new_n6632_));
  AOI21_X1   g06440(.A1(new_n6632_), .A2(new_n6631_), .B(\a[60] ), .ZN(new_n6633_));
  NAND2_X1   g06441(.A1(new_n6590_), .A2(new_n193_), .ZN(new_n6634_));
  NOR3_X1    g06442(.A1(new_n6634_), .A2(new_n6627_), .A3(new_n6629_), .ZN(new_n6635_));
  NOR4_X1    g06443(.A1(new_n6624_), .A2(\asqrt[63] ), .A3(new_n6627_), .A4(new_n6599_), .ZN(new_n6636_));
  NOR2_X1    g06444(.A1(new_n6636_), .A2(new_n6290_), .ZN(new_n6637_));
  NOR3_X1    g06445(.A1(new_n6637_), .A2(new_n6635_), .A3(new_n6292_), .ZN(new_n6638_));
  NOR2_X1    g06446(.A1(new_n6638_), .A2(new_n6633_), .ZN(new_n6639_));
  INV_X1     g06447(.I(\a[58] ), .ZN(new_n6640_));
  NOR2_X1    g06448(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n6641_));
  NOR3_X1    g06449(.A1(new_n6636_), .A2(new_n6640_), .A3(new_n6641_), .ZN(new_n6642_));
  INV_X1     g06450(.I(new_n6641_), .ZN(new_n6643_));
  AOI21_X1   g06451(.A1(new_n6636_), .A2(\a[58] ), .B(new_n6643_), .ZN(new_n6644_));
  OAI21_X1   g06452(.A1(new_n6642_), .A2(new_n6644_), .B(\asqrt[30] ), .ZN(new_n6645_));
  NAND2_X1   g06453(.A1(new_n6641_), .A2(new_n6640_), .ZN(new_n6646_));
  NAND3_X1   g06454(.A1(new_n6254_), .A2(new_n6256_), .A3(new_n6646_), .ZN(new_n6647_));
  NAND2_X1   g06455(.A1(new_n6279_), .A2(new_n6647_), .ZN(new_n6648_));
  INV_X1     g06456(.I(new_n6648_), .ZN(new_n6649_));
  NOR3_X1    g06457(.A1(new_n6636_), .A2(new_n6640_), .A3(new_n6649_), .ZN(new_n6650_));
  NOR3_X1    g06458(.A1(new_n6636_), .A2(\a[58] ), .A3(\a[59] ), .ZN(new_n6651_));
  INV_X1     g06459(.I(\a[59] ), .ZN(new_n6652_));
  AOI21_X1   g06460(.A1(\asqrt[29] ), .A2(new_n6640_), .B(new_n6652_), .ZN(new_n6653_));
  NOR3_X1    g06461(.A1(new_n6650_), .A2(new_n6651_), .A3(new_n6653_), .ZN(new_n6654_));
  NAND3_X1   g06462(.A1(new_n6654_), .A2(new_n6645_), .A3(new_n5947_), .ZN(new_n6655_));
  NAND2_X1   g06463(.A1(new_n6655_), .A2(new_n6639_), .ZN(new_n6656_));
  NAND3_X1   g06464(.A1(\asqrt[29] ), .A2(\a[58] ), .A3(new_n6643_), .ZN(new_n6657_));
  OAI21_X1   g06465(.A1(\asqrt[29] ), .A2(new_n6640_), .B(new_n6641_), .ZN(new_n6658_));
  AOI21_X1   g06466(.A1(new_n6658_), .A2(new_n6657_), .B(new_n6275_), .ZN(new_n6659_));
  NAND3_X1   g06467(.A1(\asqrt[29] ), .A2(\a[58] ), .A3(new_n6648_), .ZN(new_n6660_));
  NAND3_X1   g06468(.A1(\asqrt[29] ), .A2(new_n6640_), .A3(new_n6652_), .ZN(new_n6661_));
  OAI21_X1   g06469(.A1(new_n6636_), .A2(\a[58] ), .B(\a[59] ), .ZN(new_n6662_));
  NAND3_X1   g06470(.A1(new_n6660_), .A2(new_n6662_), .A3(new_n6661_), .ZN(new_n6663_));
  OAI21_X1   g06471(.A1(new_n6663_), .A2(new_n6659_), .B(\asqrt[31] ), .ZN(new_n6664_));
  NAND3_X1   g06472(.A1(new_n6656_), .A2(new_n5643_), .A3(new_n6664_), .ZN(new_n6665_));
  AOI21_X1   g06473(.A1(new_n6656_), .A2(new_n6664_), .B(new_n5643_), .ZN(new_n6666_));
  AOI21_X1   g06474(.A1(new_n6618_), .A2(new_n6665_), .B(new_n6666_), .ZN(new_n6667_));
  AOI21_X1   g06475(.A1(new_n6667_), .A2(new_n5336_), .B(new_n6612_), .ZN(new_n6668_));
  OR2_X2     g06476(.A1(new_n6638_), .A2(new_n6633_), .Z(new_n6669_));
  NOR3_X1    g06477(.A1(new_n6663_), .A2(new_n6659_), .A3(\asqrt[31] ), .ZN(new_n6670_));
  OAI21_X1   g06478(.A1(new_n6669_), .A2(new_n6670_), .B(new_n6664_), .ZN(new_n6671_));
  OAI21_X1   g06479(.A1(new_n6671_), .A2(\asqrt[32] ), .B(new_n6618_), .ZN(new_n6672_));
  NAND2_X1   g06480(.A1(new_n6671_), .A2(\asqrt[32] ), .ZN(new_n6673_));
  AOI21_X1   g06481(.A1(new_n6672_), .A2(new_n6673_), .B(new_n5336_), .ZN(new_n6674_));
  NOR3_X1    g06482(.A1(new_n6668_), .A2(\asqrt[34] ), .A3(new_n6674_), .ZN(new_n6675_));
  OAI21_X1   g06483(.A1(new_n6668_), .A2(new_n6674_), .B(\asqrt[34] ), .ZN(new_n6676_));
  OAI21_X1   g06484(.A1(new_n6609_), .A2(new_n6675_), .B(new_n6676_), .ZN(new_n6677_));
  OAI21_X1   g06485(.A1(new_n6677_), .A2(\asqrt[35] ), .B(new_n6605_), .ZN(new_n6678_));
  NAND3_X1   g06486(.A1(new_n6672_), .A2(new_n6673_), .A3(new_n5336_), .ZN(new_n6679_));
  AOI21_X1   g06487(.A1(new_n6611_), .A2(new_n6679_), .B(new_n6674_), .ZN(new_n6680_));
  AOI21_X1   g06488(.A1(new_n6680_), .A2(new_n5029_), .B(new_n6609_), .ZN(new_n6681_));
  NAND2_X1   g06489(.A1(new_n6679_), .A2(new_n6611_), .ZN(new_n6682_));
  INV_X1     g06490(.I(new_n6674_), .ZN(new_n6683_));
  AOI21_X1   g06491(.A1(new_n6682_), .A2(new_n6683_), .B(new_n5029_), .ZN(new_n6684_));
  OAI21_X1   g06492(.A1(new_n6681_), .A2(new_n6684_), .B(\asqrt[35] ), .ZN(new_n6685_));
  NAND3_X1   g06493(.A1(new_n6678_), .A2(new_n4461_), .A3(new_n6685_), .ZN(new_n6686_));
  INV_X1     g06494(.I(new_n6605_), .ZN(new_n6687_));
  NOR3_X1    g06495(.A1(new_n6681_), .A2(\asqrt[35] ), .A3(new_n6684_), .ZN(new_n6688_));
  OAI21_X1   g06496(.A1(new_n6687_), .A2(new_n6688_), .B(new_n6685_), .ZN(new_n6689_));
  NAND2_X1   g06497(.A1(new_n6689_), .A2(\asqrt[36] ), .ZN(new_n6690_));
  NOR2_X1    g06498(.A1(new_n6573_), .A2(\asqrt[62] ), .ZN(new_n6691_));
  INV_X1     g06499(.I(new_n6592_), .ZN(new_n6692_));
  NOR2_X1    g06500(.A1(new_n6692_), .A2(new_n6691_), .ZN(new_n6693_));
  XOR2_X1    g06501(.A1(new_n6583_), .A2(new_n6214_), .Z(new_n6694_));
  OAI21_X1   g06502(.A1(\asqrt[29] ), .A2(new_n6693_), .B(new_n6694_), .ZN(new_n6695_));
  INV_X1     g06503(.I(new_n6695_), .ZN(new_n6696_));
  NAND2_X1   g06504(.A1(new_n6541_), .A2(new_n337_), .ZN(new_n6697_));
  AOI21_X1   g06505(.A1(new_n6697_), .A2(new_n6565_), .B(\asqrt[29] ), .ZN(new_n6698_));
  XOR2_X1    g06506(.A1(new_n6698_), .A2(new_n6343_), .Z(new_n6699_));
  INV_X1     g06507(.I(new_n6699_), .ZN(new_n6700_));
  AOI21_X1   g06508(.A1(new_n6539_), .A2(new_n6556_), .B(\asqrt[29] ), .ZN(new_n6701_));
  XOR2_X1    g06509(.A1(new_n6701_), .A2(new_n6347_), .Z(new_n6702_));
  INV_X1     g06510(.I(new_n6702_), .ZN(new_n6703_));
  NAND2_X1   g06511(.A1(new_n6552_), .A2(new_n531_), .ZN(new_n6704_));
  AOI21_X1   g06512(.A1(new_n6704_), .A2(new_n6538_), .B(\asqrt[29] ), .ZN(new_n6705_));
  XOR2_X1    g06513(.A1(new_n6705_), .A2(new_n6350_), .Z(new_n6706_));
  INV_X1     g06514(.I(new_n6706_), .ZN(new_n6707_));
  AOI21_X1   g06515(.A1(new_n6550_), .A2(new_n6535_), .B(\asqrt[29] ), .ZN(new_n6708_));
  XOR2_X1    g06516(.A1(new_n6708_), .A2(new_n6352_), .Z(new_n6709_));
  NAND2_X1   g06517(.A1(new_n6517_), .A2(new_n744_), .ZN(new_n6710_));
  AOI21_X1   g06518(.A1(new_n6710_), .A2(new_n6549_), .B(\asqrt[29] ), .ZN(new_n6711_));
  XOR2_X1    g06519(.A1(new_n6711_), .A2(new_n6355_), .Z(new_n6712_));
  AOI21_X1   g06520(.A1(new_n6515_), .A2(new_n6532_), .B(\asqrt[29] ), .ZN(new_n6713_));
  XOR2_X1    g06521(.A1(new_n6713_), .A2(new_n6359_), .Z(new_n6714_));
  INV_X1     g06522(.I(new_n6714_), .ZN(new_n6715_));
  NAND2_X1   g06523(.A1(new_n6528_), .A2(new_n1006_), .ZN(new_n6716_));
  AOI21_X1   g06524(.A1(new_n6716_), .A2(new_n6514_), .B(\asqrt[29] ), .ZN(new_n6717_));
  XOR2_X1    g06525(.A1(new_n6717_), .A2(new_n6362_), .Z(new_n6718_));
  INV_X1     g06526(.I(new_n6718_), .ZN(new_n6719_));
  AOI21_X1   g06527(.A1(new_n6526_), .A2(new_n6511_), .B(\asqrt[29] ), .ZN(new_n6720_));
  XOR2_X1    g06528(.A1(new_n6720_), .A2(new_n6364_), .Z(new_n6721_));
  NAND2_X1   g06529(.A1(new_n6493_), .A2(new_n1305_), .ZN(new_n6722_));
  AOI21_X1   g06530(.A1(new_n6722_), .A2(new_n6525_), .B(\asqrt[29] ), .ZN(new_n6723_));
  XOR2_X1    g06531(.A1(new_n6723_), .A2(new_n6367_), .Z(new_n6724_));
  AOI21_X1   g06532(.A1(new_n6491_), .A2(new_n6508_), .B(\asqrt[29] ), .ZN(new_n6725_));
  XOR2_X1    g06533(.A1(new_n6725_), .A2(new_n6371_), .Z(new_n6726_));
  INV_X1     g06534(.I(new_n6726_), .ZN(new_n6727_));
  NAND2_X1   g06535(.A1(new_n6504_), .A2(new_n1632_), .ZN(new_n6728_));
  AOI21_X1   g06536(.A1(new_n6728_), .A2(new_n6490_), .B(\asqrt[29] ), .ZN(new_n6729_));
  XOR2_X1    g06537(.A1(new_n6729_), .A2(new_n6374_), .Z(new_n6730_));
  INV_X1     g06538(.I(new_n6730_), .ZN(new_n6731_));
  AOI21_X1   g06539(.A1(new_n6502_), .A2(new_n6487_), .B(\asqrt[29] ), .ZN(new_n6732_));
  XOR2_X1    g06540(.A1(new_n6732_), .A2(new_n6376_), .Z(new_n6733_));
  NAND2_X1   g06541(.A1(new_n6469_), .A2(new_n1953_), .ZN(new_n6734_));
  AOI21_X1   g06542(.A1(new_n6734_), .A2(new_n6501_), .B(\asqrt[29] ), .ZN(new_n6735_));
  XOR2_X1    g06543(.A1(new_n6735_), .A2(new_n6379_), .Z(new_n6736_));
  AOI21_X1   g06544(.A1(new_n6467_), .A2(new_n6484_), .B(\asqrt[29] ), .ZN(new_n6737_));
  XOR2_X1    g06545(.A1(new_n6737_), .A2(new_n6383_), .Z(new_n6738_));
  INV_X1     g06546(.I(new_n6738_), .ZN(new_n6739_));
  NAND2_X1   g06547(.A1(new_n6480_), .A2(new_n2332_), .ZN(new_n6740_));
  AOI21_X1   g06548(.A1(new_n6740_), .A2(new_n6466_), .B(\asqrt[29] ), .ZN(new_n6741_));
  XOR2_X1    g06549(.A1(new_n6741_), .A2(new_n6386_), .Z(new_n6742_));
  INV_X1     g06550(.I(new_n6742_), .ZN(new_n6743_));
  AOI21_X1   g06551(.A1(new_n6478_), .A2(new_n6463_), .B(\asqrt[29] ), .ZN(new_n6744_));
  XOR2_X1    g06552(.A1(new_n6744_), .A2(new_n6388_), .Z(new_n6745_));
  NAND2_X1   g06553(.A1(new_n6445_), .A2(new_n2749_), .ZN(new_n6746_));
  AOI21_X1   g06554(.A1(new_n6746_), .A2(new_n6477_), .B(\asqrt[29] ), .ZN(new_n6747_));
  XOR2_X1    g06555(.A1(new_n6747_), .A2(new_n6391_), .Z(new_n6748_));
  AOI21_X1   g06556(.A1(new_n6443_), .A2(new_n6460_), .B(\asqrt[29] ), .ZN(new_n6749_));
  XOR2_X1    g06557(.A1(new_n6749_), .A2(new_n6395_), .Z(new_n6750_));
  INV_X1     g06558(.I(new_n6750_), .ZN(new_n6751_));
  NAND2_X1   g06559(.A1(new_n6456_), .A2(new_n3195_), .ZN(new_n6752_));
  AOI21_X1   g06560(.A1(new_n6752_), .A2(new_n6442_), .B(\asqrt[29] ), .ZN(new_n6753_));
  XOR2_X1    g06561(.A1(new_n6753_), .A2(new_n6398_), .Z(new_n6754_));
  INV_X1     g06562(.I(new_n6754_), .ZN(new_n6755_));
  AOI21_X1   g06563(.A1(new_n6454_), .A2(new_n6439_), .B(\asqrt[29] ), .ZN(new_n6756_));
  XOR2_X1    g06564(.A1(new_n6756_), .A2(new_n6400_), .Z(new_n6757_));
  NAND2_X1   g06565(.A1(new_n6425_), .A2(new_n3681_), .ZN(new_n6758_));
  AOI21_X1   g06566(.A1(new_n6758_), .A2(new_n6453_), .B(\asqrt[29] ), .ZN(new_n6759_));
  XOR2_X1    g06567(.A1(new_n6759_), .A2(new_n6403_), .Z(new_n6760_));
  AOI21_X1   g06568(.A1(new_n6423_), .A2(new_n6436_), .B(\asqrt[29] ), .ZN(new_n6761_));
  XOR2_X1    g06569(.A1(new_n6761_), .A2(new_n6407_), .Z(new_n6762_));
  INV_X1     g06570(.I(new_n6762_), .ZN(new_n6763_));
  NAND2_X1   g06571(.A1(new_n6432_), .A2(new_n4196_), .ZN(new_n6764_));
  AOI21_X1   g06572(.A1(new_n6764_), .A2(new_n6422_), .B(\asqrt[29] ), .ZN(new_n6765_));
  XOR2_X1    g06573(.A1(new_n6765_), .A2(new_n6410_), .Z(new_n6766_));
  INV_X1     g06574(.I(new_n6766_), .ZN(new_n6767_));
  AOI21_X1   g06575(.A1(new_n6430_), .A2(new_n6419_), .B(\asqrt[29] ), .ZN(new_n6768_));
  XOR2_X1    g06576(.A1(new_n6768_), .A2(new_n6412_), .Z(new_n6769_));
  OAI21_X1   g06577(.A1(new_n6689_), .A2(\asqrt[36] ), .B(new_n6603_), .ZN(new_n6770_));
  NAND3_X1   g06578(.A1(new_n6770_), .A2(new_n6690_), .A3(new_n4196_), .ZN(new_n6771_));
  AOI21_X1   g06579(.A1(new_n6770_), .A2(new_n6690_), .B(new_n4196_), .ZN(new_n6772_));
  AOI21_X1   g06580(.A1(new_n6769_), .A2(new_n6771_), .B(new_n6772_), .ZN(new_n6773_));
  AOI21_X1   g06581(.A1(new_n6773_), .A2(new_n3925_), .B(new_n6767_), .ZN(new_n6774_));
  NAND2_X1   g06582(.A1(new_n6771_), .A2(new_n6769_), .ZN(new_n6775_));
  INV_X1     g06583(.I(new_n6772_), .ZN(new_n6776_));
  AOI21_X1   g06584(.A1(new_n6775_), .A2(new_n6776_), .B(new_n3925_), .ZN(new_n6777_));
  NOR3_X1    g06585(.A1(new_n6774_), .A2(\asqrt[39] ), .A3(new_n6777_), .ZN(new_n6778_));
  OAI21_X1   g06586(.A1(new_n6774_), .A2(new_n6777_), .B(\asqrt[39] ), .ZN(new_n6779_));
  OAI21_X1   g06587(.A1(new_n6763_), .A2(new_n6778_), .B(new_n6779_), .ZN(new_n6780_));
  OAI21_X1   g06588(.A1(new_n6780_), .A2(\asqrt[40] ), .B(new_n6760_), .ZN(new_n6781_));
  NAND2_X1   g06589(.A1(new_n6780_), .A2(\asqrt[40] ), .ZN(new_n6782_));
  NAND3_X1   g06590(.A1(new_n6781_), .A2(new_n6782_), .A3(new_n3195_), .ZN(new_n6783_));
  AOI21_X1   g06591(.A1(new_n6781_), .A2(new_n6782_), .B(new_n3195_), .ZN(new_n6784_));
  AOI21_X1   g06592(.A1(new_n6757_), .A2(new_n6783_), .B(new_n6784_), .ZN(new_n6785_));
  AOI21_X1   g06593(.A1(new_n6785_), .A2(new_n2960_), .B(new_n6755_), .ZN(new_n6786_));
  NAND2_X1   g06594(.A1(new_n6783_), .A2(new_n6757_), .ZN(new_n6787_));
  INV_X1     g06595(.I(new_n6784_), .ZN(new_n6788_));
  AOI21_X1   g06596(.A1(new_n6787_), .A2(new_n6788_), .B(new_n2960_), .ZN(new_n6789_));
  NOR3_X1    g06597(.A1(new_n6786_), .A2(\asqrt[43] ), .A3(new_n6789_), .ZN(new_n6790_));
  OAI21_X1   g06598(.A1(new_n6786_), .A2(new_n6789_), .B(\asqrt[43] ), .ZN(new_n6791_));
  OAI21_X1   g06599(.A1(new_n6751_), .A2(new_n6790_), .B(new_n6791_), .ZN(new_n6792_));
  OAI21_X1   g06600(.A1(new_n6792_), .A2(\asqrt[44] ), .B(new_n6748_), .ZN(new_n6793_));
  NAND2_X1   g06601(.A1(new_n6792_), .A2(\asqrt[44] ), .ZN(new_n6794_));
  NAND3_X1   g06602(.A1(new_n6793_), .A2(new_n6794_), .A3(new_n2332_), .ZN(new_n6795_));
  AOI21_X1   g06603(.A1(new_n6793_), .A2(new_n6794_), .B(new_n2332_), .ZN(new_n6796_));
  AOI21_X1   g06604(.A1(new_n6745_), .A2(new_n6795_), .B(new_n6796_), .ZN(new_n6797_));
  AOI21_X1   g06605(.A1(new_n6797_), .A2(new_n2134_), .B(new_n6743_), .ZN(new_n6798_));
  NAND2_X1   g06606(.A1(new_n6795_), .A2(new_n6745_), .ZN(new_n6799_));
  INV_X1     g06607(.I(new_n6796_), .ZN(new_n6800_));
  AOI21_X1   g06608(.A1(new_n6799_), .A2(new_n6800_), .B(new_n2134_), .ZN(new_n6801_));
  NOR3_X1    g06609(.A1(new_n6798_), .A2(\asqrt[47] ), .A3(new_n6801_), .ZN(new_n6802_));
  OAI21_X1   g06610(.A1(new_n6798_), .A2(new_n6801_), .B(\asqrt[47] ), .ZN(new_n6803_));
  OAI21_X1   g06611(.A1(new_n6739_), .A2(new_n6802_), .B(new_n6803_), .ZN(new_n6804_));
  OAI21_X1   g06612(.A1(new_n6804_), .A2(\asqrt[48] ), .B(new_n6736_), .ZN(new_n6805_));
  NAND2_X1   g06613(.A1(new_n6804_), .A2(\asqrt[48] ), .ZN(new_n6806_));
  NAND3_X1   g06614(.A1(new_n6805_), .A2(new_n6806_), .A3(new_n1632_), .ZN(new_n6807_));
  AOI21_X1   g06615(.A1(new_n6805_), .A2(new_n6806_), .B(new_n1632_), .ZN(new_n6808_));
  AOI21_X1   g06616(.A1(new_n6733_), .A2(new_n6807_), .B(new_n6808_), .ZN(new_n6809_));
  AOI21_X1   g06617(.A1(new_n6809_), .A2(new_n1463_), .B(new_n6731_), .ZN(new_n6810_));
  NAND2_X1   g06618(.A1(new_n6807_), .A2(new_n6733_), .ZN(new_n6811_));
  INV_X1     g06619(.I(new_n6808_), .ZN(new_n6812_));
  AOI21_X1   g06620(.A1(new_n6811_), .A2(new_n6812_), .B(new_n1463_), .ZN(new_n6813_));
  NOR3_X1    g06621(.A1(new_n6810_), .A2(\asqrt[51] ), .A3(new_n6813_), .ZN(new_n6814_));
  OAI21_X1   g06622(.A1(new_n6810_), .A2(new_n6813_), .B(\asqrt[51] ), .ZN(new_n6815_));
  OAI21_X1   g06623(.A1(new_n6727_), .A2(new_n6814_), .B(new_n6815_), .ZN(new_n6816_));
  OAI21_X1   g06624(.A1(new_n6816_), .A2(\asqrt[52] ), .B(new_n6724_), .ZN(new_n6817_));
  NAND2_X1   g06625(.A1(new_n6816_), .A2(\asqrt[52] ), .ZN(new_n6818_));
  NAND3_X1   g06626(.A1(new_n6817_), .A2(new_n6818_), .A3(new_n1006_), .ZN(new_n6819_));
  AOI21_X1   g06627(.A1(new_n6817_), .A2(new_n6818_), .B(new_n1006_), .ZN(new_n6820_));
  AOI21_X1   g06628(.A1(new_n6721_), .A2(new_n6819_), .B(new_n6820_), .ZN(new_n6821_));
  AOI21_X1   g06629(.A1(new_n6821_), .A2(new_n860_), .B(new_n6719_), .ZN(new_n6822_));
  NAND2_X1   g06630(.A1(new_n6819_), .A2(new_n6721_), .ZN(new_n6823_));
  INV_X1     g06631(.I(new_n6820_), .ZN(new_n6824_));
  AOI21_X1   g06632(.A1(new_n6823_), .A2(new_n6824_), .B(new_n860_), .ZN(new_n6825_));
  NOR3_X1    g06633(.A1(new_n6822_), .A2(\asqrt[55] ), .A3(new_n6825_), .ZN(new_n6826_));
  OAI21_X1   g06634(.A1(new_n6822_), .A2(new_n6825_), .B(\asqrt[55] ), .ZN(new_n6827_));
  OAI21_X1   g06635(.A1(new_n6715_), .A2(new_n6826_), .B(new_n6827_), .ZN(new_n6828_));
  OAI21_X1   g06636(.A1(new_n6828_), .A2(\asqrt[56] ), .B(new_n6712_), .ZN(new_n6829_));
  NAND2_X1   g06637(.A1(new_n6828_), .A2(\asqrt[56] ), .ZN(new_n6830_));
  NAND3_X1   g06638(.A1(new_n6829_), .A2(new_n6830_), .A3(new_n531_), .ZN(new_n6831_));
  AOI21_X1   g06639(.A1(new_n6829_), .A2(new_n6830_), .B(new_n531_), .ZN(new_n6832_));
  AOI21_X1   g06640(.A1(new_n6709_), .A2(new_n6831_), .B(new_n6832_), .ZN(new_n6833_));
  AOI21_X1   g06641(.A1(new_n6833_), .A2(new_n423_), .B(new_n6707_), .ZN(new_n6834_));
  NAND2_X1   g06642(.A1(new_n6831_), .A2(new_n6709_), .ZN(new_n6835_));
  INV_X1     g06643(.I(new_n6832_), .ZN(new_n6836_));
  AOI21_X1   g06644(.A1(new_n6835_), .A2(new_n6836_), .B(new_n423_), .ZN(new_n6837_));
  NOR3_X1    g06645(.A1(new_n6834_), .A2(\asqrt[59] ), .A3(new_n6837_), .ZN(new_n6838_));
  NOR2_X1    g06646(.A1(new_n6838_), .A2(new_n6703_), .ZN(new_n6839_));
  OAI21_X1   g06647(.A1(new_n6834_), .A2(new_n6837_), .B(\asqrt[59] ), .ZN(new_n6840_));
  INV_X1     g06648(.I(new_n6840_), .ZN(new_n6841_));
  NOR2_X1    g06649(.A1(new_n6839_), .A2(new_n6841_), .ZN(new_n6842_));
  AOI21_X1   g06650(.A1(new_n6842_), .A2(new_n266_), .B(new_n6700_), .ZN(new_n6843_));
  INV_X1     g06651(.I(new_n6709_), .ZN(new_n6844_));
  INV_X1     g06652(.I(new_n6721_), .ZN(new_n6845_));
  INV_X1     g06653(.I(new_n6733_), .ZN(new_n6846_));
  INV_X1     g06654(.I(new_n6745_), .ZN(new_n6847_));
  INV_X1     g06655(.I(new_n6757_), .ZN(new_n6848_));
  INV_X1     g06656(.I(new_n6769_), .ZN(new_n6849_));
  AOI21_X1   g06657(.A1(new_n6678_), .A2(new_n6685_), .B(new_n4461_), .ZN(new_n6850_));
  AOI21_X1   g06658(.A1(new_n6603_), .A2(new_n6686_), .B(new_n6850_), .ZN(new_n6851_));
  AOI21_X1   g06659(.A1(new_n6851_), .A2(new_n4196_), .B(new_n6849_), .ZN(new_n6852_));
  NOR3_X1    g06660(.A1(new_n6852_), .A2(\asqrt[38] ), .A3(new_n6772_), .ZN(new_n6853_));
  OAI21_X1   g06661(.A1(new_n6852_), .A2(new_n6772_), .B(\asqrt[38] ), .ZN(new_n6854_));
  OAI21_X1   g06662(.A1(new_n6767_), .A2(new_n6853_), .B(new_n6854_), .ZN(new_n6855_));
  OAI21_X1   g06663(.A1(new_n6855_), .A2(\asqrt[39] ), .B(new_n6762_), .ZN(new_n6856_));
  NAND3_X1   g06664(.A1(new_n6856_), .A2(new_n3427_), .A3(new_n6779_), .ZN(new_n6857_));
  AOI21_X1   g06665(.A1(new_n6856_), .A2(new_n6779_), .B(new_n3427_), .ZN(new_n6858_));
  AOI21_X1   g06666(.A1(new_n6760_), .A2(new_n6857_), .B(new_n6858_), .ZN(new_n6859_));
  AOI21_X1   g06667(.A1(new_n6859_), .A2(new_n3195_), .B(new_n6848_), .ZN(new_n6860_));
  NOR3_X1    g06668(.A1(new_n6860_), .A2(\asqrt[42] ), .A3(new_n6784_), .ZN(new_n6861_));
  OAI21_X1   g06669(.A1(new_n6860_), .A2(new_n6784_), .B(\asqrt[42] ), .ZN(new_n6862_));
  OAI21_X1   g06670(.A1(new_n6755_), .A2(new_n6861_), .B(new_n6862_), .ZN(new_n6863_));
  OAI21_X1   g06671(.A1(new_n6863_), .A2(\asqrt[43] ), .B(new_n6750_), .ZN(new_n6864_));
  NAND3_X1   g06672(.A1(new_n6864_), .A2(new_n2531_), .A3(new_n6791_), .ZN(new_n6865_));
  AOI21_X1   g06673(.A1(new_n6864_), .A2(new_n6791_), .B(new_n2531_), .ZN(new_n6866_));
  AOI21_X1   g06674(.A1(new_n6748_), .A2(new_n6865_), .B(new_n6866_), .ZN(new_n6867_));
  AOI21_X1   g06675(.A1(new_n6867_), .A2(new_n2332_), .B(new_n6847_), .ZN(new_n6868_));
  NOR3_X1    g06676(.A1(new_n6868_), .A2(\asqrt[46] ), .A3(new_n6796_), .ZN(new_n6869_));
  OAI21_X1   g06677(.A1(new_n6868_), .A2(new_n6796_), .B(\asqrt[46] ), .ZN(new_n6870_));
  OAI21_X1   g06678(.A1(new_n6743_), .A2(new_n6869_), .B(new_n6870_), .ZN(new_n6871_));
  OAI21_X1   g06679(.A1(new_n6871_), .A2(\asqrt[47] ), .B(new_n6738_), .ZN(new_n6872_));
  NAND3_X1   g06680(.A1(new_n6872_), .A2(new_n1778_), .A3(new_n6803_), .ZN(new_n6873_));
  AOI21_X1   g06681(.A1(new_n6872_), .A2(new_n6803_), .B(new_n1778_), .ZN(new_n6874_));
  AOI21_X1   g06682(.A1(new_n6736_), .A2(new_n6873_), .B(new_n6874_), .ZN(new_n6875_));
  AOI21_X1   g06683(.A1(new_n6875_), .A2(new_n1632_), .B(new_n6846_), .ZN(new_n6876_));
  NOR3_X1    g06684(.A1(new_n6876_), .A2(\asqrt[50] ), .A3(new_n6808_), .ZN(new_n6877_));
  OAI21_X1   g06685(.A1(new_n6876_), .A2(new_n6808_), .B(\asqrt[50] ), .ZN(new_n6878_));
  OAI21_X1   g06686(.A1(new_n6731_), .A2(new_n6877_), .B(new_n6878_), .ZN(new_n6879_));
  OAI21_X1   g06687(.A1(new_n6879_), .A2(\asqrt[51] ), .B(new_n6726_), .ZN(new_n6880_));
  NAND3_X1   g06688(.A1(new_n6880_), .A2(new_n1150_), .A3(new_n6815_), .ZN(new_n6881_));
  AOI21_X1   g06689(.A1(new_n6880_), .A2(new_n6815_), .B(new_n1150_), .ZN(new_n6882_));
  AOI21_X1   g06690(.A1(new_n6724_), .A2(new_n6881_), .B(new_n6882_), .ZN(new_n6883_));
  AOI21_X1   g06691(.A1(new_n6883_), .A2(new_n1006_), .B(new_n6845_), .ZN(new_n6884_));
  NOR3_X1    g06692(.A1(new_n6884_), .A2(\asqrt[54] ), .A3(new_n6820_), .ZN(new_n6885_));
  OAI21_X1   g06693(.A1(new_n6884_), .A2(new_n6820_), .B(\asqrt[54] ), .ZN(new_n6886_));
  OAI21_X1   g06694(.A1(new_n6719_), .A2(new_n6885_), .B(new_n6886_), .ZN(new_n6887_));
  OAI21_X1   g06695(.A1(new_n6887_), .A2(\asqrt[55] ), .B(new_n6714_), .ZN(new_n6888_));
  NAND3_X1   g06696(.A1(new_n6888_), .A2(new_n634_), .A3(new_n6827_), .ZN(new_n6889_));
  AOI21_X1   g06697(.A1(new_n6888_), .A2(new_n6827_), .B(new_n634_), .ZN(new_n6890_));
  AOI21_X1   g06698(.A1(new_n6712_), .A2(new_n6889_), .B(new_n6890_), .ZN(new_n6891_));
  AOI21_X1   g06699(.A1(new_n6891_), .A2(new_n531_), .B(new_n6844_), .ZN(new_n6892_));
  NOR3_X1    g06700(.A1(new_n6892_), .A2(\asqrt[58] ), .A3(new_n6832_), .ZN(new_n6893_));
  OAI21_X1   g06701(.A1(new_n6892_), .A2(new_n6832_), .B(\asqrt[58] ), .ZN(new_n6894_));
  OAI21_X1   g06702(.A1(new_n6707_), .A2(new_n6893_), .B(new_n6894_), .ZN(new_n6895_));
  OAI21_X1   g06703(.A1(new_n6895_), .A2(\asqrt[59] ), .B(new_n6702_), .ZN(new_n6896_));
  AOI21_X1   g06704(.A1(new_n6896_), .A2(new_n6840_), .B(new_n266_), .ZN(new_n6897_));
  OAI21_X1   g06705(.A1(new_n6843_), .A2(new_n6897_), .B(\asqrt[61] ), .ZN(new_n6898_));
  AOI21_X1   g06706(.A1(new_n6574_), .A2(new_n6568_), .B(\asqrt[29] ), .ZN(new_n6899_));
  XOR2_X1    g06707(.A1(new_n6899_), .A2(new_n6340_), .Z(new_n6900_));
  OAI21_X1   g06708(.A1(new_n6703_), .A2(new_n6838_), .B(new_n6840_), .ZN(new_n6901_));
  OAI21_X1   g06709(.A1(new_n6901_), .A2(\asqrt[60] ), .B(new_n6699_), .ZN(new_n6902_));
  OAI21_X1   g06710(.A1(new_n6839_), .A2(new_n6841_), .B(\asqrt[60] ), .ZN(new_n6903_));
  NAND3_X1   g06711(.A1(new_n6902_), .A2(new_n239_), .A3(new_n6903_), .ZN(new_n6904_));
  NAND2_X1   g06712(.A1(new_n6904_), .A2(new_n6900_), .ZN(new_n6905_));
  NAND2_X1   g06713(.A1(new_n6905_), .A2(new_n6898_), .ZN(new_n6906_));
  AOI21_X1   g06714(.A1(new_n6902_), .A2(new_n6903_), .B(new_n239_), .ZN(new_n6907_));
  NAND3_X1   g06715(.A1(new_n6896_), .A2(new_n266_), .A3(new_n6840_), .ZN(new_n6908_));
  AOI21_X1   g06716(.A1(new_n6699_), .A2(new_n6908_), .B(new_n6897_), .ZN(new_n6909_));
  INV_X1     g06717(.I(new_n6900_), .ZN(new_n6910_));
  AOI21_X1   g06718(.A1(new_n6909_), .A2(new_n239_), .B(new_n6910_), .ZN(new_n6911_));
  OAI21_X1   g06719(.A1(new_n6911_), .A2(new_n6907_), .B(new_n201_), .ZN(new_n6912_));
  NAND3_X1   g06720(.A1(new_n6905_), .A2(\asqrt[62] ), .A3(new_n6898_), .ZN(new_n6913_));
  AOI21_X1   g06721(.A1(new_n6567_), .A2(new_n6619_), .B(\asqrt[29] ), .ZN(new_n6914_));
  XOR2_X1    g06722(.A1(new_n6914_), .A2(new_n6571_), .Z(new_n6915_));
  INV_X1     g06723(.I(new_n6915_), .ZN(new_n6916_));
  AOI22_X1   g06724(.A1(new_n6912_), .A2(new_n6913_), .B1(new_n6906_), .B2(new_n6916_), .ZN(new_n6917_));
  NOR2_X1    g06725(.A1(new_n6586_), .A2(new_n6338_), .ZN(new_n6918_));
  OAI21_X1   g06726(.A1(\asqrt[29] ), .A2(new_n6918_), .B(new_n6593_), .ZN(new_n6919_));
  INV_X1     g06727(.I(new_n6919_), .ZN(new_n6920_));
  OAI21_X1   g06728(.A1(new_n6917_), .A2(new_n6696_), .B(new_n6920_), .ZN(new_n6921_));
  OAI21_X1   g06729(.A1(new_n6906_), .A2(\asqrt[62] ), .B(new_n6915_), .ZN(new_n6922_));
  NAND2_X1   g06730(.A1(new_n6906_), .A2(\asqrt[62] ), .ZN(new_n6923_));
  NAND3_X1   g06731(.A1(new_n6922_), .A2(new_n6923_), .A3(new_n6696_), .ZN(new_n6924_));
  NAND2_X1   g06732(.A1(new_n6636_), .A2(new_n6337_), .ZN(new_n6925_));
  XOR2_X1    g06733(.A1(new_n6586_), .A2(new_n6338_), .Z(new_n6926_));
  NAND3_X1   g06734(.A1(new_n6925_), .A2(\asqrt[63] ), .A3(new_n6926_), .ZN(new_n6927_));
  INV_X1     g06735(.I(new_n6634_), .ZN(new_n6928_));
  NAND4_X1   g06736(.A1(new_n6928_), .A2(new_n6338_), .A3(new_n6593_), .A4(new_n6600_), .ZN(new_n6929_));
  NAND2_X1   g06737(.A1(new_n6927_), .A2(new_n6929_), .ZN(new_n6930_));
  INV_X1     g06738(.I(new_n6930_), .ZN(new_n6931_));
  NAND4_X1   g06739(.A1(new_n6921_), .A2(new_n193_), .A3(new_n6924_), .A4(new_n6931_), .ZN(\asqrt[28] ));
  AOI21_X1   g06740(.A1(new_n6686_), .A2(new_n6690_), .B(\asqrt[28] ), .ZN(new_n6933_));
  XOR2_X1    g06741(.A1(new_n6933_), .A2(new_n6603_), .Z(new_n6934_));
  XOR2_X1    g06742(.A1(new_n6677_), .A2(\asqrt[35] ), .Z(new_n6935_));
  NOR2_X1    g06743(.A1(\asqrt[28] ), .A2(new_n6935_), .ZN(new_n6936_));
  XOR2_X1    g06744(.A1(new_n6936_), .A2(new_n6605_), .Z(new_n6937_));
  NOR2_X1    g06745(.A1(new_n6675_), .A2(new_n6684_), .ZN(new_n6938_));
  NOR2_X1    g06746(.A1(\asqrt[28] ), .A2(new_n6938_), .ZN(new_n6939_));
  XOR2_X1    g06747(.A1(new_n6939_), .A2(new_n6608_), .Z(new_n6940_));
  AOI21_X1   g06748(.A1(new_n6679_), .A2(new_n6683_), .B(\asqrt[28] ), .ZN(new_n6941_));
  XOR2_X1    g06749(.A1(new_n6941_), .A2(new_n6611_), .Z(new_n6942_));
  INV_X1     g06750(.I(new_n6942_), .ZN(new_n6943_));
  AOI21_X1   g06751(.A1(new_n6665_), .A2(new_n6673_), .B(\asqrt[28] ), .ZN(new_n6944_));
  XOR2_X1    g06752(.A1(new_n6944_), .A2(new_n6618_), .Z(new_n6945_));
  INV_X1     g06753(.I(new_n6945_), .ZN(new_n6946_));
  AOI21_X1   g06754(.A1(new_n6655_), .A2(new_n6664_), .B(\asqrt[28] ), .ZN(new_n6947_));
  XOR2_X1    g06755(.A1(new_n6947_), .A2(new_n6639_), .Z(new_n6948_));
  NAND2_X1   g06756(.A1(\asqrt[29] ), .A2(new_n6640_), .ZN(new_n6949_));
  NOR2_X1    g06757(.A1(new_n6652_), .A2(\a[58] ), .ZN(new_n6950_));
  AOI22_X1   g06758(.A1(new_n6949_), .A2(new_n6652_), .B1(\asqrt[29] ), .B2(new_n6950_), .ZN(new_n6951_));
  OAI21_X1   g06759(.A1(new_n6636_), .A2(new_n6640_), .B(new_n6649_), .ZN(new_n6952_));
  AOI21_X1   g06760(.A1(new_n6645_), .A2(new_n6952_), .B(\asqrt[28] ), .ZN(new_n6953_));
  XOR2_X1    g06761(.A1(new_n6953_), .A2(new_n6951_), .Z(new_n6954_));
  NAND2_X1   g06762(.A1(new_n6921_), .A2(new_n193_), .ZN(new_n6955_));
  NOR2_X1    g06763(.A1(new_n6911_), .A2(new_n6907_), .ZN(new_n6956_));
  AOI21_X1   g06764(.A1(new_n6956_), .A2(new_n201_), .B(new_n6916_), .ZN(new_n6957_));
  OAI21_X1   g06765(.A1(new_n6956_), .A2(new_n201_), .B(new_n6696_), .ZN(new_n6958_));
  NOR2_X1    g06766(.A1(new_n6957_), .A2(new_n6958_), .ZN(new_n6959_));
  NAND3_X1   g06767(.A1(new_n6927_), .A2(\asqrt[29] ), .A3(new_n6929_), .ZN(new_n6960_));
  NOR3_X1    g06768(.A1(new_n6955_), .A2(new_n6959_), .A3(new_n6960_), .ZN(new_n6961_));
  AOI21_X1   g06769(.A1(new_n6905_), .A2(new_n6898_), .B(\asqrt[62] ), .ZN(new_n6962_));
  NOR3_X1    g06770(.A1(new_n6911_), .A2(new_n201_), .A3(new_n6907_), .ZN(new_n6963_));
  OAI22_X1   g06771(.A1(new_n6963_), .A2(new_n6962_), .B1(new_n6956_), .B2(new_n6915_), .ZN(new_n6964_));
  AOI21_X1   g06772(.A1(new_n6964_), .A2(new_n6695_), .B(new_n6919_), .ZN(new_n6965_));
  NOR4_X1    g06773(.A1(new_n6965_), .A2(\asqrt[63] ), .A3(new_n6959_), .A4(new_n6930_), .ZN(new_n6966_));
  NOR2_X1    g06774(.A1(new_n6966_), .A2(new_n6643_), .ZN(new_n6967_));
  OAI21_X1   g06775(.A1(new_n6967_), .A2(new_n6961_), .B(new_n6640_), .ZN(new_n6968_));
  NOR3_X1    g06776(.A1(new_n6965_), .A2(\asqrt[63] ), .A3(new_n6959_), .ZN(new_n6969_));
  NAND4_X1   g06777(.A1(new_n6969_), .A2(\asqrt[29] ), .A3(new_n6927_), .A4(new_n6929_), .ZN(new_n6970_));
  NAND2_X1   g06778(.A1(\asqrt[28] ), .A2(new_n6641_), .ZN(new_n6971_));
  NAND3_X1   g06779(.A1(new_n6970_), .A2(new_n6971_), .A3(\a[58] ), .ZN(new_n6972_));
  NAND2_X1   g06780(.A1(new_n6972_), .A2(new_n6968_), .ZN(new_n6973_));
  NOR2_X1    g06781(.A1(\a[54] ), .A2(\a[55] ), .ZN(new_n6974_));
  INV_X1     g06782(.I(new_n6974_), .ZN(new_n6975_));
  NAND3_X1   g06783(.A1(\asqrt[28] ), .A2(\a[56] ), .A3(new_n6975_), .ZN(new_n6976_));
  INV_X1     g06784(.I(\a[56] ), .ZN(new_n6977_));
  OAI21_X1   g06785(.A1(\asqrt[28] ), .A2(new_n6977_), .B(new_n6974_), .ZN(new_n6978_));
  AOI21_X1   g06786(.A1(new_n6978_), .A2(new_n6976_), .B(new_n6636_), .ZN(new_n6979_));
  NAND2_X1   g06787(.A1(new_n6974_), .A2(new_n6977_), .ZN(new_n6980_));
  NAND3_X1   g06788(.A1(new_n6596_), .A2(new_n6598_), .A3(new_n6980_), .ZN(new_n6981_));
  NAND2_X1   g06789(.A1(new_n6628_), .A2(new_n6981_), .ZN(new_n6982_));
  NAND3_X1   g06790(.A1(\asqrt[28] ), .A2(\a[56] ), .A3(new_n6982_), .ZN(new_n6983_));
  INV_X1     g06791(.I(\a[57] ), .ZN(new_n6984_));
  NAND3_X1   g06792(.A1(\asqrt[28] ), .A2(new_n6977_), .A3(new_n6984_), .ZN(new_n6985_));
  OAI21_X1   g06793(.A1(new_n6966_), .A2(\a[56] ), .B(\a[57] ), .ZN(new_n6986_));
  NAND3_X1   g06794(.A1(new_n6986_), .A2(new_n6983_), .A3(new_n6985_), .ZN(new_n6987_));
  NOR3_X1    g06795(.A1(new_n6987_), .A2(new_n6979_), .A3(\asqrt[30] ), .ZN(new_n6988_));
  OAI21_X1   g06796(.A1(new_n6987_), .A2(new_n6979_), .B(\asqrt[30] ), .ZN(new_n6989_));
  OAI21_X1   g06797(.A1(new_n6973_), .A2(new_n6988_), .B(new_n6989_), .ZN(new_n6990_));
  OAI21_X1   g06798(.A1(new_n6990_), .A2(\asqrt[31] ), .B(new_n6954_), .ZN(new_n6991_));
  NAND2_X1   g06799(.A1(new_n6990_), .A2(\asqrt[31] ), .ZN(new_n6992_));
  NAND3_X1   g06800(.A1(new_n6991_), .A2(new_n6992_), .A3(new_n5643_), .ZN(new_n6993_));
  AOI21_X1   g06801(.A1(new_n6991_), .A2(new_n6992_), .B(new_n5643_), .ZN(new_n6994_));
  AOI21_X1   g06802(.A1(new_n6948_), .A2(new_n6993_), .B(new_n6994_), .ZN(new_n6995_));
  AOI21_X1   g06803(.A1(new_n6995_), .A2(new_n5336_), .B(new_n6946_), .ZN(new_n6996_));
  NAND2_X1   g06804(.A1(new_n6993_), .A2(new_n6948_), .ZN(new_n6997_));
  INV_X1     g06805(.I(new_n6954_), .ZN(new_n6998_));
  INV_X1     g06806(.I(new_n6973_), .ZN(new_n6999_));
  NOR3_X1    g06807(.A1(new_n6966_), .A2(new_n6977_), .A3(new_n6974_), .ZN(new_n7000_));
  AOI21_X1   g06808(.A1(new_n6966_), .A2(\a[56] ), .B(new_n6975_), .ZN(new_n7001_));
  OAI21_X1   g06809(.A1(new_n7000_), .A2(new_n7001_), .B(\asqrt[29] ), .ZN(new_n7002_));
  INV_X1     g06810(.I(new_n6982_), .ZN(new_n7003_));
  NOR3_X1    g06811(.A1(new_n6966_), .A2(new_n6977_), .A3(new_n7003_), .ZN(new_n7004_));
  NOR3_X1    g06812(.A1(new_n6966_), .A2(\a[56] ), .A3(\a[57] ), .ZN(new_n7005_));
  AOI21_X1   g06813(.A1(\asqrt[28] ), .A2(new_n6977_), .B(new_n6984_), .ZN(new_n7006_));
  NOR3_X1    g06814(.A1(new_n7004_), .A2(new_n7005_), .A3(new_n7006_), .ZN(new_n7007_));
  NAND3_X1   g06815(.A1(new_n7002_), .A2(new_n7007_), .A3(new_n6275_), .ZN(new_n7008_));
  AOI21_X1   g06816(.A1(new_n7002_), .A2(new_n7007_), .B(new_n6275_), .ZN(new_n7009_));
  AOI21_X1   g06817(.A1(new_n6999_), .A2(new_n7008_), .B(new_n7009_), .ZN(new_n7010_));
  AOI21_X1   g06818(.A1(new_n7010_), .A2(new_n5947_), .B(new_n6998_), .ZN(new_n7011_));
  NAND2_X1   g06819(.A1(new_n6999_), .A2(new_n7008_), .ZN(new_n7012_));
  AOI21_X1   g06820(.A1(new_n7012_), .A2(new_n6989_), .B(new_n5947_), .ZN(new_n7013_));
  OAI21_X1   g06821(.A1(new_n7011_), .A2(new_n7013_), .B(\asqrt[32] ), .ZN(new_n7014_));
  AOI21_X1   g06822(.A1(new_n6997_), .A2(new_n7014_), .B(new_n5336_), .ZN(new_n7015_));
  NOR3_X1    g06823(.A1(new_n6996_), .A2(\asqrt[34] ), .A3(new_n7015_), .ZN(new_n7016_));
  OAI21_X1   g06824(.A1(new_n6996_), .A2(new_n7015_), .B(\asqrt[34] ), .ZN(new_n7017_));
  OAI21_X1   g06825(.A1(new_n6943_), .A2(new_n7016_), .B(new_n7017_), .ZN(new_n7018_));
  OAI21_X1   g06826(.A1(new_n7018_), .A2(\asqrt[35] ), .B(new_n6940_), .ZN(new_n7019_));
  NAND2_X1   g06827(.A1(new_n7018_), .A2(\asqrt[35] ), .ZN(new_n7020_));
  NAND3_X1   g06828(.A1(new_n7019_), .A2(new_n7020_), .A3(new_n4461_), .ZN(new_n7021_));
  AOI21_X1   g06829(.A1(new_n7019_), .A2(new_n7020_), .B(new_n4461_), .ZN(new_n7022_));
  AOI21_X1   g06830(.A1(new_n6937_), .A2(new_n7021_), .B(new_n7022_), .ZN(new_n7023_));
  NAND2_X1   g06831(.A1(new_n7023_), .A2(new_n4196_), .ZN(new_n7024_));
  INV_X1     g06832(.I(new_n6937_), .ZN(new_n7025_));
  INV_X1     g06833(.I(new_n6940_), .ZN(new_n7026_));
  INV_X1     g06834(.I(new_n6948_), .ZN(new_n7027_));
  NOR3_X1    g06835(.A1(new_n7011_), .A2(\asqrt[32] ), .A3(new_n7013_), .ZN(new_n7028_));
  OAI21_X1   g06836(.A1(new_n7027_), .A2(new_n7028_), .B(new_n7014_), .ZN(new_n7029_));
  OAI21_X1   g06837(.A1(new_n7029_), .A2(\asqrt[33] ), .B(new_n6945_), .ZN(new_n7030_));
  NAND2_X1   g06838(.A1(new_n7029_), .A2(\asqrt[33] ), .ZN(new_n7031_));
  NAND3_X1   g06839(.A1(new_n7030_), .A2(new_n7031_), .A3(new_n5029_), .ZN(new_n7032_));
  AOI21_X1   g06840(.A1(new_n7030_), .A2(new_n7031_), .B(new_n5029_), .ZN(new_n7033_));
  AOI21_X1   g06841(.A1(new_n6942_), .A2(new_n7032_), .B(new_n7033_), .ZN(new_n7034_));
  AOI21_X1   g06842(.A1(new_n7034_), .A2(new_n4751_), .B(new_n7026_), .ZN(new_n7035_));
  NAND2_X1   g06843(.A1(new_n7032_), .A2(new_n6942_), .ZN(new_n7036_));
  AOI21_X1   g06844(.A1(new_n7036_), .A2(new_n7017_), .B(new_n4751_), .ZN(new_n7037_));
  NOR3_X1    g06845(.A1(new_n7035_), .A2(\asqrt[36] ), .A3(new_n7037_), .ZN(new_n7038_));
  OAI21_X1   g06846(.A1(new_n7035_), .A2(new_n7037_), .B(\asqrt[36] ), .ZN(new_n7039_));
  OAI21_X1   g06847(.A1(new_n7025_), .A2(new_n7038_), .B(new_n7039_), .ZN(new_n7040_));
  NAND2_X1   g06848(.A1(new_n7040_), .A2(\asqrt[37] ), .ZN(new_n7041_));
  NOR2_X1    g06849(.A1(new_n6906_), .A2(\asqrt[62] ), .ZN(new_n7042_));
  INV_X1     g06850(.I(new_n6923_), .ZN(new_n7043_));
  NOR2_X1    g06851(.A1(new_n7043_), .A2(new_n7042_), .ZN(new_n7044_));
  XOR2_X1    g06852(.A1(new_n6914_), .A2(new_n6571_), .Z(new_n7045_));
  OAI21_X1   g06853(.A1(\asqrt[28] ), .A2(new_n7044_), .B(new_n7045_), .ZN(new_n7046_));
  INV_X1     g06854(.I(new_n7046_), .ZN(new_n7047_));
  NOR2_X1    g06855(.A1(new_n6841_), .A2(new_n6838_), .ZN(new_n7048_));
  NOR2_X1    g06856(.A1(\asqrt[28] ), .A2(new_n7048_), .ZN(new_n7049_));
  XOR2_X1    g06857(.A1(new_n7049_), .A2(new_n6702_), .Z(new_n7050_));
  INV_X1     g06858(.I(new_n7050_), .ZN(new_n7051_));
  NOR2_X1    g06859(.A1(new_n6893_), .A2(new_n6837_), .ZN(new_n7052_));
  NOR2_X1    g06860(.A1(\asqrt[28] ), .A2(new_n7052_), .ZN(new_n7053_));
  XOR2_X1    g06861(.A1(new_n7053_), .A2(new_n6706_), .Z(new_n7054_));
  AOI21_X1   g06862(.A1(new_n6831_), .A2(new_n6836_), .B(\asqrt[28] ), .ZN(new_n7055_));
  XOR2_X1    g06863(.A1(new_n7055_), .A2(new_n6709_), .Z(new_n7056_));
  AOI21_X1   g06864(.A1(new_n6889_), .A2(new_n6830_), .B(\asqrt[28] ), .ZN(new_n7057_));
  XOR2_X1    g06865(.A1(new_n7057_), .A2(new_n6712_), .Z(new_n7058_));
  INV_X1     g06866(.I(new_n6827_), .ZN(new_n7059_));
  NOR2_X1    g06867(.A1(new_n7059_), .A2(new_n6826_), .ZN(new_n7060_));
  NOR2_X1    g06868(.A1(\asqrt[28] ), .A2(new_n7060_), .ZN(new_n7061_));
  XOR2_X1    g06869(.A1(new_n7061_), .A2(new_n6714_), .Z(new_n7062_));
  INV_X1     g06870(.I(new_n7062_), .ZN(new_n7063_));
  NOR2_X1    g06871(.A1(new_n6885_), .A2(new_n6825_), .ZN(new_n7064_));
  NOR2_X1    g06872(.A1(\asqrt[28] ), .A2(new_n7064_), .ZN(new_n7065_));
  XOR2_X1    g06873(.A1(new_n7065_), .A2(new_n6718_), .Z(new_n7066_));
  INV_X1     g06874(.I(new_n7066_), .ZN(new_n7067_));
  AOI21_X1   g06875(.A1(new_n6819_), .A2(new_n6824_), .B(\asqrt[28] ), .ZN(new_n7068_));
  XOR2_X1    g06876(.A1(new_n7068_), .A2(new_n6721_), .Z(new_n7069_));
  AOI21_X1   g06877(.A1(new_n6881_), .A2(new_n6818_), .B(\asqrt[28] ), .ZN(new_n7070_));
  XOR2_X1    g06878(.A1(new_n7070_), .A2(new_n6724_), .Z(new_n7071_));
  XOR2_X1    g06879(.A1(new_n6879_), .A2(\asqrt[51] ), .Z(new_n7072_));
  NOR2_X1    g06880(.A1(\asqrt[28] ), .A2(new_n7072_), .ZN(new_n7073_));
  XOR2_X1    g06881(.A1(new_n7073_), .A2(new_n6726_), .Z(new_n7074_));
  INV_X1     g06882(.I(new_n7074_), .ZN(new_n7075_));
  NOR2_X1    g06883(.A1(new_n6877_), .A2(new_n6813_), .ZN(new_n7076_));
  NOR2_X1    g06884(.A1(\asqrt[28] ), .A2(new_n7076_), .ZN(new_n7077_));
  XOR2_X1    g06885(.A1(new_n7077_), .A2(new_n6730_), .Z(new_n7078_));
  INV_X1     g06886(.I(new_n7078_), .ZN(new_n7079_));
  AOI21_X1   g06887(.A1(new_n6807_), .A2(new_n6812_), .B(\asqrt[28] ), .ZN(new_n7080_));
  XOR2_X1    g06888(.A1(new_n7080_), .A2(new_n6733_), .Z(new_n7081_));
  AOI21_X1   g06889(.A1(new_n6873_), .A2(new_n6806_), .B(\asqrt[28] ), .ZN(new_n7082_));
  XOR2_X1    g06890(.A1(new_n7082_), .A2(new_n6736_), .Z(new_n7083_));
  XOR2_X1    g06891(.A1(new_n6871_), .A2(\asqrt[47] ), .Z(new_n7084_));
  NOR2_X1    g06892(.A1(\asqrt[28] ), .A2(new_n7084_), .ZN(new_n7085_));
  XOR2_X1    g06893(.A1(new_n7085_), .A2(new_n6738_), .Z(new_n7086_));
  INV_X1     g06894(.I(new_n7086_), .ZN(new_n7087_));
  NOR2_X1    g06895(.A1(new_n6869_), .A2(new_n6801_), .ZN(new_n7088_));
  NOR2_X1    g06896(.A1(\asqrt[28] ), .A2(new_n7088_), .ZN(new_n7089_));
  XOR2_X1    g06897(.A1(new_n7089_), .A2(new_n6742_), .Z(new_n7090_));
  INV_X1     g06898(.I(new_n7090_), .ZN(new_n7091_));
  AOI21_X1   g06899(.A1(new_n6795_), .A2(new_n6800_), .B(\asqrt[28] ), .ZN(new_n7092_));
  XOR2_X1    g06900(.A1(new_n7092_), .A2(new_n6745_), .Z(new_n7093_));
  AOI21_X1   g06901(.A1(new_n6865_), .A2(new_n6794_), .B(\asqrt[28] ), .ZN(new_n7094_));
  XOR2_X1    g06902(.A1(new_n7094_), .A2(new_n6748_), .Z(new_n7095_));
  XOR2_X1    g06903(.A1(new_n6863_), .A2(\asqrt[43] ), .Z(new_n7096_));
  NOR2_X1    g06904(.A1(\asqrt[28] ), .A2(new_n7096_), .ZN(new_n7097_));
  XOR2_X1    g06905(.A1(new_n7097_), .A2(new_n6750_), .Z(new_n7098_));
  INV_X1     g06906(.I(new_n7098_), .ZN(new_n7099_));
  NOR2_X1    g06907(.A1(new_n6861_), .A2(new_n6789_), .ZN(new_n7100_));
  NOR2_X1    g06908(.A1(\asqrt[28] ), .A2(new_n7100_), .ZN(new_n7101_));
  XOR2_X1    g06909(.A1(new_n7101_), .A2(new_n6754_), .Z(new_n7102_));
  INV_X1     g06910(.I(new_n7102_), .ZN(new_n7103_));
  AOI21_X1   g06911(.A1(new_n6783_), .A2(new_n6788_), .B(\asqrt[28] ), .ZN(new_n7104_));
  XOR2_X1    g06912(.A1(new_n7104_), .A2(new_n6757_), .Z(new_n7105_));
  AOI21_X1   g06913(.A1(new_n6857_), .A2(new_n6782_), .B(\asqrt[28] ), .ZN(new_n7106_));
  XOR2_X1    g06914(.A1(new_n7106_), .A2(new_n6760_), .Z(new_n7107_));
  XOR2_X1    g06915(.A1(new_n6855_), .A2(\asqrt[39] ), .Z(new_n7108_));
  NOR2_X1    g06916(.A1(\asqrt[28] ), .A2(new_n7108_), .ZN(new_n7109_));
  XOR2_X1    g06917(.A1(new_n7109_), .A2(new_n6762_), .Z(new_n7110_));
  INV_X1     g06918(.I(new_n7110_), .ZN(new_n7111_));
  NOR2_X1    g06919(.A1(new_n6853_), .A2(new_n6777_), .ZN(new_n7112_));
  NOR2_X1    g06920(.A1(\asqrt[28] ), .A2(new_n7112_), .ZN(new_n7113_));
  XOR2_X1    g06921(.A1(new_n7113_), .A2(new_n6766_), .Z(new_n7114_));
  INV_X1     g06922(.I(new_n7114_), .ZN(new_n7115_));
  AOI21_X1   g06923(.A1(new_n6771_), .A2(new_n6776_), .B(\asqrt[28] ), .ZN(new_n7116_));
  XOR2_X1    g06924(.A1(new_n7116_), .A2(new_n6769_), .Z(new_n7117_));
  OAI21_X1   g06925(.A1(new_n7040_), .A2(\asqrt[37] ), .B(new_n6934_), .ZN(new_n7118_));
  NAND3_X1   g06926(.A1(new_n7118_), .A2(new_n7041_), .A3(new_n3925_), .ZN(new_n7119_));
  AOI21_X1   g06927(.A1(new_n7118_), .A2(new_n7041_), .B(new_n3925_), .ZN(new_n7120_));
  AOI21_X1   g06928(.A1(new_n7117_), .A2(new_n7119_), .B(new_n7120_), .ZN(new_n7121_));
  AOI21_X1   g06929(.A1(new_n7121_), .A2(new_n3681_), .B(new_n7115_), .ZN(new_n7122_));
  NAND2_X1   g06930(.A1(new_n7119_), .A2(new_n7117_), .ZN(new_n7123_));
  INV_X1     g06931(.I(new_n6934_), .ZN(new_n7124_));
  AOI21_X1   g06932(.A1(new_n7023_), .A2(new_n4196_), .B(new_n7124_), .ZN(new_n7125_));
  NAND2_X1   g06933(.A1(new_n7021_), .A2(new_n6937_), .ZN(new_n7126_));
  AOI21_X1   g06934(.A1(new_n7126_), .A2(new_n7039_), .B(new_n4196_), .ZN(new_n7127_));
  OAI21_X1   g06935(.A1(new_n7125_), .A2(new_n7127_), .B(\asqrt[38] ), .ZN(new_n7128_));
  AOI21_X1   g06936(.A1(new_n7123_), .A2(new_n7128_), .B(new_n3681_), .ZN(new_n7129_));
  NOR3_X1    g06937(.A1(new_n7122_), .A2(\asqrt[40] ), .A3(new_n7129_), .ZN(new_n7130_));
  OAI21_X1   g06938(.A1(new_n7122_), .A2(new_n7129_), .B(\asqrt[40] ), .ZN(new_n7131_));
  OAI21_X1   g06939(.A1(new_n7111_), .A2(new_n7130_), .B(new_n7131_), .ZN(new_n7132_));
  OAI21_X1   g06940(.A1(new_n7132_), .A2(\asqrt[41] ), .B(new_n7107_), .ZN(new_n7133_));
  NAND2_X1   g06941(.A1(new_n7132_), .A2(\asqrt[41] ), .ZN(new_n7134_));
  NAND3_X1   g06942(.A1(new_n7133_), .A2(new_n7134_), .A3(new_n2960_), .ZN(new_n7135_));
  AOI21_X1   g06943(.A1(new_n7133_), .A2(new_n7134_), .B(new_n2960_), .ZN(new_n7136_));
  AOI21_X1   g06944(.A1(new_n7105_), .A2(new_n7135_), .B(new_n7136_), .ZN(new_n7137_));
  AOI21_X1   g06945(.A1(new_n7137_), .A2(new_n2749_), .B(new_n7103_), .ZN(new_n7138_));
  NAND2_X1   g06946(.A1(new_n7135_), .A2(new_n7105_), .ZN(new_n7139_));
  INV_X1     g06947(.I(new_n7107_), .ZN(new_n7140_));
  INV_X1     g06948(.I(new_n7117_), .ZN(new_n7141_));
  NOR3_X1    g06949(.A1(new_n7125_), .A2(\asqrt[38] ), .A3(new_n7127_), .ZN(new_n7142_));
  OAI21_X1   g06950(.A1(new_n7141_), .A2(new_n7142_), .B(new_n7128_), .ZN(new_n7143_));
  OAI21_X1   g06951(.A1(new_n7143_), .A2(\asqrt[39] ), .B(new_n7114_), .ZN(new_n7144_));
  NAND2_X1   g06952(.A1(new_n7143_), .A2(\asqrt[39] ), .ZN(new_n7145_));
  NAND3_X1   g06953(.A1(new_n7144_), .A2(new_n7145_), .A3(new_n3427_), .ZN(new_n7146_));
  AOI21_X1   g06954(.A1(new_n7144_), .A2(new_n7145_), .B(new_n3427_), .ZN(new_n7147_));
  AOI21_X1   g06955(.A1(new_n7110_), .A2(new_n7146_), .B(new_n7147_), .ZN(new_n7148_));
  AOI21_X1   g06956(.A1(new_n7148_), .A2(new_n3195_), .B(new_n7140_), .ZN(new_n7149_));
  NAND2_X1   g06957(.A1(new_n7146_), .A2(new_n7110_), .ZN(new_n7150_));
  AOI21_X1   g06958(.A1(new_n7150_), .A2(new_n7131_), .B(new_n3195_), .ZN(new_n7151_));
  OAI21_X1   g06959(.A1(new_n7149_), .A2(new_n7151_), .B(\asqrt[42] ), .ZN(new_n7152_));
  AOI21_X1   g06960(.A1(new_n7139_), .A2(new_n7152_), .B(new_n2749_), .ZN(new_n7153_));
  NOR3_X1    g06961(.A1(new_n7138_), .A2(\asqrt[44] ), .A3(new_n7153_), .ZN(new_n7154_));
  OAI21_X1   g06962(.A1(new_n7138_), .A2(new_n7153_), .B(\asqrt[44] ), .ZN(new_n7155_));
  OAI21_X1   g06963(.A1(new_n7099_), .A2(new_n7154_), .B(new_n7155_), .ZN(new_n7156_));
  OAI21_X1   g06964(.A1(new_n7156_), .A2(\asqrt[45] ), .B(new_n7095_), .ZN(new_n7157_));
  NAND2_X1   g06965(.A1(new_n7156_), .A2(\asqrt[45] ), .ZN(new_n7158_));
  NAND3_X1   g06966(.A1(new_n7157_), .A2(new_n7158_), .A3(new_n2134_), .ZN(new_n7159_));
  AOI21_X1   g06967(.A1(new_n7157_), .A2(new_n7158_), .B(new_n2134_), .ZN(new_n7160_));
  AOI21_X1   g06968(.A1(new_n7093_), .A2(new_n7159_), .B(new_n7160_), .ZN(new_n7161_));
  AOI21_X1   g06969(.A1(new_n7161_), .A2(new_n1953_), .B(new_n7091_), .ZN(new_n7162_));
  NAND2_X1   g06970(.A1(new_n7159_), .A2(new_n7093_), .ZN(new_n7163_));
  INV_X1     g06971(.I(new_n7095_), .ZN(new_n7164_));
  INV_X1     g06972(.I(new_n7105_), .ZN(new_n7165_));
  NOR3_X1    g06973(.A1(new_n7149_), .A2(\asqrt[42] ), .A3(new_n7151_), .ZN(new_n7166_));
  OAI21_X1   g06974(.A1(new_n7165_), .A2(new_n7166_), .B(new_n7152_), .ZN(new_n7167_));
  OAI21_X1   g06975(.A1(new_n7167_), .A2(\asqrt[43] ), .B(new_n7102_), .ZN(new_n7168_));
  NAND2_X1   g06976(.A1(new_n7167_), .A2(\asqrt[43] ), .ZN(new_n7169_));
  NAND3_X1   g06977(.A1(new_n7168_), .A2(new_n7169_), .A3(new_n2531_), .ZN(new_n7170_));
  AOI21_X1   g06978(.A1(new_n7168_), .A2(new_n7169_), .B(new_n2531_), .ZN(new_n7171_));
  AOI21_X1   g06979(.A1(new_n7098_), .A2(new_n7170_), .B(new_n7171_), .ZN(new_n7172_));
  AOI21_X1   g06980(.A1(new_n7172_), .A2(new_n2332_), .B(new_n7164_), .ZN(new_n7173_));
  NAND2_X1   g06981(.A1(new_n7170_), .A2(new_n7098_), .ZN(new_n7174_));
  AOI21_X1   g06982(.A1(new_n7174_), .A2(new_n7155_), .B(new_n2332_), .ZN(new_n7175_));
  OAI21_X1   g06983(.A1(new_n7173_), .A2(new_n7175_), .B(\asqrt[46] ), .ZN(new_n7176_));
  AOI21_X1   g06984(.A1(new_n7163_), .A2(new_n7176_), .B(new_n1953_), .ZN(new_n7177_));
  NOR3_X1    g06985(.A1(new_n7162_), .A2(\asqrt[48] ), .A3(new_n7177_), .ZN(new_n7178_));
  OAI21_X1   g06986(.A1(new_n7162_), .A2(new_n7177_), .B(\asqrt[48] ), .ZN(new_n7179_));
  OAI21_X1   g06987(.A1(new_n7087_), .A2(new_n7178_), .B(new_n7179_), .ZN(new_n7180_));
  OAI21_X1   g06988(.A1(new_n7180_), .A2(\asqrt[49] ), .B(new_n7083_), .ZN(new_n7181_));
  NAND2_X1   g06989(.A1(new_n7180_), .A2(\asqrt[49] ), .ZN(new_n7182_));
  NAND3_X1   g06990(.A1(new_n7181_), .A2(new_n7182_), .A3(new_n1463_), .ZN(new_n7183_));
  AOI21_X1   g06991(.A1(new_n7181_), .A2(new_n7182_), .B(new_n1463_), .ZN(new_n7184_));
  AOI21_X1   g06992(.A1(new_n7081_), .A2(new_n7183_), .B(new_n7184_), .ZN(new_n7185_));
  AOI21_X1   g06993(.A1(new_n7185_), .A2(new_n1305_), .B(new_n7079_), .ZN(new_n7186_));
  NAND2_X1   g06994(.A1(new_n7183_), .A2(new_n7081_), .ZN(new_n7187_));
  INV_X1     g06995(.I(new_n7083_), .ZN(new_n7188_));
  INV_X1     g06996(.I(new_n7093_), .ZN(new_n7189_));
  NOR3_X1    g06997(.A1(new_n7173_), .A2(\asqrt[46] ), .A3(new_n7175_), .ZN(new_n7190_));
  OAI21_X1   g06998(.A1(new_n7189_), .A2(new_n7190_), .B(new_n7176_), .ZN(new_n7191_));
  OAI21_X1   g06999(.A1(new_n7191_), .A2(\asqrt[47] ), .B(new_n7090_), .ZN(new_n7192_));
  NAND2_X1   g07000(.A1(new_n7191_), .A2(\asqrt[47] ), .ZN(new_n7193_));
  NAND3_X1   g07001(.A1(new_n7192_), .A2(new_n7193_), .A3(new_n1778_), .ZN(new_n7194_));
  AOI21_X1   g07002(.A1(new_n7192_), .A2(new_n7193_), .B(new_n1778_), .ZN(new_n7195_));
  AOI21_X1   g07003(.A1(new_n7086_), .A2(new_n7194_), .B(new_n7195_), .ZN(new_n7196_));
  AOI21_X1   g07004(.A1(new_n7196_), .A2(new_n1632_), .B(new_n7188_), .ZN(new_n7197_));
  NAND2_X1   g07005(.A1(new_n7194_), .A2(new_n7086_), .ZN(new_n7198_));
  AOI21_X1   g07006(.A1(new_n7198_), .A2(new_n7179_), .B(new_n1632_), .ZN(new_n7199_));
  OAI21_X1   g07007(.A1(new_n7197_), .A2(new_n7199_), .B(\asqrt[50] ), .ZN(new_n7200_));
  AOI21_X1   g07008(.A1(new_n7187_), .A2(new_n7200_), .B(new_n1305_), .ZN(new_n7201_));
  NOR3_X1    g07009(.A1(new_n7186_), .A2(\asqrt[52] ), .A3(new_n7201_), .ZN(new_n7202_));
  OAI21_X1   g07010(.A1(new_n7186_), .A2(new_n7201_), .B(\asqrt[52] ), .ZN(new_n7203_));
  OAI21_X1   g07011(.A1(new_n7075_), .A2(new_n7202_), .B(new_n7203_), .ZN(new_n7204_));
  OAI21_X1   g07012(.A1(new_n7204_), .A2(\asqrt[53] ), .B(new_n7071_), .ZN(new_n7205_));
  NAND2_X1   g07013(.A1(new_n7204_), .A2(\asqrt[53] ), .ZN(new_n7206_));
  NAND3_X1   g07014(.A1(new_n7205_), .A2(new_n7206_), .A3(new_n860_), .ZN(new_n7207_));
  AOI21_X1   g07015(.A1(new_n7205_), .A2(new_n7206_), .B(new_n860_), .ZN(new_n7208_));
  AOI21_X1   g07016(.A1(new_n7069_), .A2(new_n7207_), .B(new_n7208_), .ZN(new_n7209_));
  AOI21_X1   g07017(.A1(new_n7209_), .A2(new_n744_), .B(new_n7067_), .ZN(new_n7210_));
  NAND2_X1   g07018(.A1(new_n7207_), .A2(new_n7069_), .ZN(new_n7211_));
  INV_X1     g07019(.I(new_n7071_), .ZN(new_n7212_));
  INV_X1     g07020(.I(new_n7081_), .ZN(new_n7213_));
  NOR3_X1    g07021(.A1(new_n7197_), .A2(\asqrt[50] ), .A3(new_n7199_), .ZN(new_n7214_));
  OAI21_X1   g07022(.A1(new_n7213_), .A2(new_n7214_), .B(new_n7200_), .ZN(new_n7215_));
  OAI21_X1   g07023(.A1(new_n7215_), .A2(\asqrt[51] ), .B(new_n7078_), .ZN(new_n7216_));
  NAND2_X1   g07024(.A1(new_n7215_), .A2(\asqrt[51] ), .ZN(new_n7217_));
  NAND3_X1   g07025(.A1(new_n7216_), .A2(new_n7217_), .A3(new_n1150_), .ZN(new_n7218_));
  AOI21_X1   g07026(.A1(new_n7216_), .A2(new_n7217_), .B(new_n1150_), .ZN(new_n7219_));
  AOI21_X1   g07027(.A1(new_n7074_), .A2(new_n7218_), .B(new_n7219_), .ZN(new_n7220_));
  AOI21_X1   g07028(.A1(new_n7220_), .A2(new_n1006_), .B(new_n7212_), .ZN(new_n7221_));
  NAND2_X1   g07029(.A1(new_n7218_), .A2(new_n7074_), .ZN(new_n7222_));
  AOI21_X1   g07030(.A1(new_n7222_), .A2(new_n7203_), .B(new_n1006_), .ZN(new_n7223_));
  OAI21_X1   g07031(.A1(new_n7221_), .A2(new_n7223_), .B(\asqrt[54] ), .ZN(new_n7224_));
  AOI21_X1   g07032(.A1(new_n7211_), .A2(new_n7224_), .B(new_n744_), .ZN(new_n7225_));
  NOR3_X1    g07033(.A1(new_n7210_), .A2(\asqrt[56] ), .A3(new_n7225_), .ZN(new_n7226_));
  OAI21_X1   g07034(.A1(new_n7210_), .A2(new_n7225_), .B(\asqrt[56] ), .ZN(new_n7227_));
  OAI21_X1   g07035(.A1(new_n7063_), .A2(new_n7226_), .B(new_n7227_), .ZN(new_n7228_));
  OAI21_X1   g07036(.A1(new_n7228_), .A2(\asqrt[57] ), .B(new_n7058_), .ZN(new_n7229_));
  NOR2_X1    g07037(.A1(new_n7226_), .A2(new_n7063_), .ZN(new_n7230_));
  INV_X1     g07038(.I(new_n7069_), .ZN(new_n7231_));
  NOR3_X1    g07039(.A1(new_n7221_), .A2(\asqrt[54] ), .A3(new_n7223_), .ZN(new_n7232_));
  OAI21_X1   g07040(.A1(new_n7231_), .A2(new_n7232_), .B(new_n7224_), .ZN(new_n7233_));
  OAI21_X1   g07041(.A1(new_n7233_), .A2(\asqrt[55] ), .B(new_n7066_), .ZN(new_n7234_));
  NAND2_X1   g07042(.A1(new_n7233_), .A2(\asqrt[55] ), .ZN(new_n7235_));
  AOI21_X1   g07043(.A1(new_n7234_), .A2(new_n7235_), .B(new_n634_), .ZN(new_n7236_));
  OAI21_X1   g07044(.A1(new_n7230_), .A2(new_n7236_), .B(\asqrt[57] ), .ZN(new_n7237_));
  NAND3_X1   g07045(.A1(new_n7229_), .A2(new_n423_), .A3(new_n7237_), .ZN(new_n7238_));
  NAND2_X1   g07046(.A1(new_n7238_), .A2(new_n7056_), .ZN(new_n7239_));
  INV_X1     g07047(.I(new_n7058_), .ZN(new_n7240_));
  NAND3_X1   g07048(.A1(new_n7234_), .A2(new_n7235_), .A3(new_n634_), .ZN(new_n7241_));
  AOI21_X1   g07049(.A1(new_n7062_), .A2(new_n7241_), .B(new_n7236_), .ZN(new_n7242_));
  AOI21_X1   g07050(.A1(new_n7242_), .A2(new_n531_), .B(new_n7240_), .ZN(new_n7243_));
  NAND2_X1   g07051(.A1(new_n7241_), .A2(new_n7062_), .ZN(new_n7244_));
  AOI21_X1   g07052(.A1(new_n7244_), .A2(new_n7227_), .B(new_n531_), .ZN(new_n7245_));
  OAI21_X1   g07053(.A1(new_n7243_), .A2(new_n7245_), .B(\asqrt[58] ), .ZN(new_n7246_));
  NAND3_X1   g07054(.A1(new_n7239_), .A2(new_n337_), .A3(new_n7246_), .ZN(new_n7247_));
  AOI21_X1   g07055(.A1(new_n7239_), .A2(new_n7246_), .B(new_n337_), .ZN(new_n7248_));
  AOI21_X1   g07056(.A1(new_n7054_), .A2(new_n7247_), .B(new_n7248_), .ZN(new_n7249_));
  AOI21_X1   g07057(.A1(new_n7249_), .A2(new_n266_), .B(new_n7051_), .ZN(new_n7250_));
  INV_X1     g07058(.I(new_n7056_), .ZN(new_n7251_));
  NOR3_X1    g07059(.A1(new_n7243_), .A2(\asqrt[58] ), .A3(new_n7245_), .ZN(new_n7252_));
  OAI21_X1   g07060(.A1(new_n7251_), .A2(new_n7252_), .B(new_n7246_), .ZN(new_n7253_));
  OAI21_X1   g07061(.A1(new_n7253_), .A2(\asqrt[59] ), .B(new_n7054_), .ZN(new_n7254_));
  NAND2_X1   g07062(.A1(new_n7253_), .A2(\asqrt[59] ), .ZN(new_n7255_));
  AOI21_X1   g07063(.A1(new_n7254_), .A2(new_n7255_), .B(new_n266_), .ZN(new_n7256_));
  OAI21_X1   g07064(.A1(new_n7250_), .A2(new_n7256_), .B(\asqrt[61] ), .ZN(new_n7257_));
  AOI21_X1   g07065(.A1(new_n6908_), .A2(new_n6903_), .B(\asqrt[28] ), .ZN(new_n7258_));
  XOR2_X1    g07066(.A1(new_n7258_), .A2(new_n6699_), .Z(new_n7259_));
  INV_X1     g07067(.I(new_n7259_), .ZN(new_n7260_));
  NOR3_X1    g07068(.A1(new_n7250_), .A2(\asqrt[61] ), .A3(new_n7256_), .ZN(new_n7261_));
  OAI21_X1   g07069(.A1(new_n7260_), .A2(new_n7261_), .B(new_n7257_), .ZN(new_n7262_));
  NAND3_X1   g07070(.A1(new_n7254_), .A2(new_n7255_), .A3(new_n266_), .ZN(new_n7263_));
  NAND2_X1   g07071(.A1(new_n7263_), .A2(new_n7050_), .ZN(new_n7264_));
  INV_X1     g07072(.I(new_n7054_), .ZN(new_n7265_));
  AOI21_X1   g07073(.A1(new_n7229_), .A2(new_n7237_), .B(new_n423_), .ZN(new_n7266_));
  AOI21_X1   g07074(.A1(new_n7056_), .A2(new_n7238_), .B(new_n7266_), .ZN(new_n7267_));
  AOI21_X1   g07075(.A1(new_n7267_), .A2(new_n337_), .B(new_n7265_), .ZN(new_n7268_));
  OAI21_X1   g07076(.A1(new_n7268_), .A2(new_n7248_), .B(\asqrt[60] ), .ZN(new_n7269_));
  AOI21_X1   g07077(.A1(new_n7264_), .A2(new_n7269_), .B(new_n239_), .ZN(new_n7270_));
  AOI21_X1   g07078(.A1(new_n7050_), .A2(new_n7263_), .B(new_n7256_), .ZN(new_n7271_));
  AOI21_X1   g07079(.A1(new_n7271_), .A2(new_n239_), .B(new_n7260_), .ZN(new_n7272_));
  OAI21_X1   g07080(.A1(new_n7272_), .A2(new_n7270_), .B(new_n201_), .ZN(new_n7273_));
  NOR3_X1    g07081(.A1(new_n7268_), .A2(\asqrt[60] ), .A3(new_n7248_), .ZN(new_n7274_));
  OAI21_X1   g07082(.A1(new_n7051_), .A2(new_n7274_), .B(new_n7269_), .ZN(new_n7275_));
  OAI21_X1   g07083(.A1(new_n7275_), .A2(\asqrt[61] ), .B(new_n7259_), .ZN(new_n7276_));
  NAND3_X1   g07084(.A1(new_n7276_), .A2(\asqrt[62] ), .A3(new_n7257_), .ZN(new_n7277_));
  AOI21_X1   g07085(.A1(new_n6898_), .A2(new_n6904_), .B(\asqrt[28] ), .ZN(new_n7278_));
  XOR2_X1    g07086(.A1(new_n7278_), .A2(new_n6900_), .Z(new_n7279_));
  INV_X1     g07087(.I(new_n7279_), .ZN(new_n7280_));
  AOI22_X1   g07088(.A1(new_n7277_), .A2(new_n7273_), .B1(new_n7262_), .B2(new_n7280_), .ZN(new_n7281_));
  NOR2_X1    g07089(.A1(new_n6917_), .A2(new_n6696_), .ZN(new_n7282_));
  OAI21_X1   g07090(.A1(\asqrt[28] ), .A2(new_n7282_), .B(new_n6924_), .ZN(new_n7283_));
  INV_X1     g07091(.I(new_n7283_), .ZN(new_n7284_));
  OAI21_X1   g07092(.A1(new_n7281_), .A2(new_n7047_), .B(new_n7284_), .ZN(new_n7285_));
  OAI21_X1   g07093(.A1(new_n7262_), .A2(\asqrt[62] ), .B(new_n7279_), .ZN(new_n7286_));
  NAND2_X1   g07094(.A1(new_n7262_), .A2(\asqrt[62] ), .ZN(new_n7287_));
  NAND3_X1   g07095(.A1(new_n7286_), .A2(new_n7287_), .A3(new_n7047_), .ZN(new_n7288_));
  NAND2_X1   g07096(.A1(new_n6966_), .A2(new_n6695_), .ZN(new_n7289_));
  XOR2_X1    g07097(.A1(new_n6917_), .A2(new_n6696_), .Z(new_n7290_));
  NAND3_X1   g07098(.A1(new_n7289_), .A2(\asqrt[63] ), .A3(new_n7290_), .ZN(new_n7291_));
  INV_X1     g07099(.I(new_n6955_), .ZN(new_n7292_));
  NAND4_X1   g07100(.A1(new_n7292_), .A2(new_n6696_), .A3(new_n6924_), .A4(new_n6931_), .ZN(new_n7293_));
  NAND2_X1   g07101(.A1(new_n7291_), .A2(new_n7293_), .ZN(new_n7294_));
  INV_X1     g07102(.I(new_n7294_), .ZN(new_n7295_));
  NAND4_X1   g07103(.A1(new_n7285_), .A2(new_n193_), .A3(new_n7288_), .A4(new_n7295_), .ZN(\asqrt[27] ));
  AOI21_X1   g07104(.A1(new_n7024_), .A2(new_n7041_), .B(\asqrt[27] ), .ZN(new_n7297_));
  XOR2_X1    g07105(.A1(new_n7297_), .A2(new_n6934_), .Z(new_n7298_));
  AOI21_X1   g07106(.A1(new_n7021_), .A2(new_n7039_), .B(\asqrt[27] ), .ZN(new_n7299_));
  XOR2_X1    g07107(.A1(new_n7299_), .A2(new_n6937_), .Z(new_n7300_));
  NAND2_X1   g07108(.A1(new_n7034_), .A2(new_n4751_), .ZN(new_n7301_));
  AOI21_X1   g07109(.A1(new_n7301_), .A2(new_n7020_), .B(\asqrt[27] ), .ZN(new_n7302_));
  XOR2_X1    g07110(.A1(new_n7302_), .A2(new_n6940_), .Z(new_n7303_));
  INV_X1     g07111(.I(new_n7303_), .ZN(new_n7304_));
  AOI21_X1   g07112(.A1(new_n7032_), .A2(new_n7017_), .B(\asqrt[27] ), .ZN(new_n7305_));
  XOR2_X1    g07113(.A1(new_n7305_), .A2(new_n6942_), .Z(new_n7306_));
  INV_X1     g07114(.I(new_n7306_), .ZN(new_n7307_));
  NAND2_X1   g07115(.A1(new_n6995_), .A2(new_n5336_), .ZN(new_n7308_));
  AOI21_X1   g07116(.A1(new_n7308_), .A2(new_n7031_), .B(\asqrt[27] ), .ZN(new_n7309_));
  XOR2_X1    g07117(.A1(new_n7309_), .A2(new_n6945_), .Z(new_n7310_));
  AOI21_X1   g07118(.A1(new_n6993_), .A2(new_n7014_), .B(\asqrt[27] ), .ZN(new_n7311_));
  XOR2_X1    g07119(.A1(new_n7311_), .A2(new_n6948_), .Z(new_n7312_));
  NAND2_X1   g07120(.A1(new_n7010_), .A2(new_n5947_), .ZN(new_n7313_));
  AOI21_X1   g07121(.A1(new_n7313_), .A2(new_n6992_), .B(\asqrt[27] ), .ZN(new_n7314_));
  XOR2_X1    g07122(.A1(new_n7314_), .A2(new_n6954_), .Z(new_n7315_));
  INV_X1     g07123(.I(new_n7315_), .ZN(new_n7316_));
  AOI21_X1   g07124(.A1(new_n7008_), .A2(new_n6989_), .B(\asqrt[27] ), .ZN(new_n7317_));
  XOR2_X1    g07125(.A1(new_n7317_), .A2(new_n6999_), .Z(new_n7318_));
  INV_X1     g07126(.I(new_n7318_), .ZN(new_n7319_));
  NAND2_X1   g07127(.A1(\asqrt[28] ), .A2(new_n6977_), .ZN(new_n7320_));
  NOR2_X1    g07128(.A1(new_n6984_), .A2(\a[56] ), .ZN(new_n7321_));
  AOI22_X1   g07129(.A1(new_n7320_), .A2(new_n6984_), .B1(\asqrt[28] ), .B2(new_n7321_), .ZN(new_n7322_));
  NOR2_X1    g07130(.A1(new_n7272_), .A2(new_n7270_), .ZN(new_n7323_));
  AOI21_X1   g07131(.A1(new_n7276_), .A2(new_n7257_), .B(\asqrt[62] ), .ZN(new_n7324_));
  NOR3_X1    g07132(.A1(new_n7272_), .A2(new_n201_), .A3(new_n7270_), .ZN(new_n7325_));
  OAI22_X1   g07133(.A1(new_n7324_), .A2(new_n7325_), .B1(new_n7323_), .B2(new_n7279_), .ZN(new_n7326_));
  AOI21_X1   g07134(.A1(new_n7326_), .A2(new_n7046_), .B(new_n7283_), .ZN(new_n7327_));
  AOI21_X1   g07135(.A1(new_n7323_), .A2(new_n201_), .B(new_n7280_), .ZN(new_n7328_));
  NOR2_X1    g07136(.A1(new_n7323_), .A2(new_n201_), .ZN(new_n7329_));
  NOR3_X1    g07137(.A1(new_n7328_), .A2(new_n7329_), .A3(new_n7046_), .ZN(new_n7330_));
  NOR4_X1    g07138(.A1(new_n7327_), .A2(\asqrt[63] ), .A3(new_n7330_), .A4(new_n7294_), .ZN(new_n7331_));
  AOI21_X1   g07139(.A1(\asqrt[28] ), .A2(\a[56] ), .B(new_n6982_), .ZN(new_n7332_));
  OAI21_X1   g07140(.A1(new_n6979_), .A2(new_n7332_), .B(new_n7331_), .ZN(new_n7333_));
  XNOR2_X1   g07141(.A1(new_n7333_), .A2(new_n7322_), .ZN(new_n7334_));
  NAND3_X1   g07142(.A1(new_n7291_), .A2(\asqrt[28] ), .A3(new_n7293_), .ZN(new_n7335_));
  NOR4_X1    g07143(.A1(new_n7327_), .A2(\asqrt[63] ), .A3(new_n7330_), .A4(new_n7335_), .ZN(new_n7336_));
  INV_X1     g07144(.I(new_n7336_), .ZN(new_n7337_));
  NAND2_X1   g07145(.A1(\asqrt[27] ), .A2(new_n6974_), .ZN(new_n7338_));
  AOI21_X1   g07146(.A1(new_n7338_), .A2(new_n7337_), .B(\a[56] ), .ZN(new_n7339_));
  NOR2_X1    g07147(.A1(new_n7331_), .A2(new_n6975_), .ZN(new_n7340_));
  NOR3_X1    g07148(.A1(new_n7340_), .A2(new_n6977_), .A3(new_n7336_), .ZN(new_n7341_));
  NOR2_X1    g07149(.A1(new_n7341_), .A2(new_n7339_), .ZN(new_n7342_));
  INV_X1     g07150(.I(\a[54] ), .ZN(new_n7343_));
  NOR2_X1    g07151(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n7344_));
  NOR3_X1    g07152(.A1(new_n7331_), .A2(new_n7343_), .A3(new_n7344_), .ZN(new_n7345_));
  INV_X1     g07153(.I(new_n7344_), .ZN(new_n7346_));
  AOI21_X1   g07154(.A1(new_n7331_), .A2(\a[54] ), .B(new_n7346_), .ZN(new_n7347_));
  OAI21_X1   g07155(.A1(new_n7345_), .A2(new_n7347_), .B(\asqrt[28] ), .ZN(new_n7348_));
  NAND2_X1   g07156(.A1(new_n7344_), .A2(new_n7343_), .ZN(new_n7349_));
  NAND3_X1   g07157(.A1(new_n6927_), .A2(new_n6929_), .A3(new_n7349_), .ZN(new_n7350_));
  NAND2_X1   g07158(.A1(new_n6969_), .A2(new_n7350_), .ZN(new_n7351_));
  NAND3_X1   g07159(.A1(\asqrt[27] ), .A2(\a[54] ), .A3(new_n7351_), .ZN(new_n7352_));
  NOR3_X1    g07160(.A1(new_n7331_), .A2(\a[54] ), .A3(\a[55] ), .ZN(new_n7353_));
  INV_X1     g07161(.I(\a[55] ), .ZN(new_n7354_));
  AOI21_X1   g07162(.A1(\asqrt[27] ), .A2(new_n7343_), .B(new_n7354_), .ZN(new_n7355_));
  NOR2_X1    g07163(.A1(new_n7353_), .A2(new_n7355_), .ZN(new_n7356_));
  NAND4_X1   g07164(.A1(new_n7348_), .A2(new_n7356_), .A3(new_n6636_), .A4(new_n7352_), .ZN(new_n7357_));
  NAND2_X1   g07165(.A1(new_n7357_), .A2(new_n7342_), .ZN(new_n7358_));
  NAND3_X1   g07166(.A1(\asqrt[27] ), .A2(\a[54] ), .A3(new_n7346_), .ZN(new_n7359_));
  OAI21_X1   g07167(.A1(\asqrt[27] ), .A2(new_n7343_), .B(new_n7344_), .ZN(new_n7360_));
  AOI21_X1   g07168(.A1(new_n7360_), .A2(new_n7359_), .B(new_n6966_), .ZN(new_n7361_));
  NAND3_X1   g07169(.A1(\asqrt[27] ), .A2(new_n7343_), .A3(new_n7354_), .ZN(new_n7362_));
  OAI21_X1   g07170(.A1(new_n7331_), .A2(\a[54] ), .B(\a[55] ), .ZN(new_n7363_));
  NAND3_X1   g07171(.A1(new_n7352_), .A2(new_n7363_), .A3(new_n7362_), .ZN(new_n7364_));
  OAI21_X1   g07172(.A1(new_n7364_), .A2(new_n7361_), .B(\asqrt[29] ), .ZN(new_n7365_));
  NAND3_X1   g07173(.A1(new_n7358_), .A2(new_n6275_), .A3(new_n7365_), .ZN(new_n7366_));
  AOI21_X1   g07174(.A1(new_n7358_), .A2(new_n7365_), .B(new_n6275_), .ZN(new_n7367_));
  AOI21_X1   g07175(.A1(new_n7334_), .A2(new_n7366_), .B(new_n7367_), .ZN(new_n7368_));
  AOI21_X1   g07176(.A1(new_n7368_), .A2(new_n5947_), .B(new_n7319_), .ZN(new_n7369_));
  OR2_X2     g07177(.A1(new_n7341_), .A2(new_n7339_), .Z(new_n7370_));
  NOR3_X1    g07178(.A1(new_n7364_), .A2(new_n7361_), .A3(\asqrt[29] ), .ZN(new_n7371_));
  OAI21_X1   g07179(.A1(new_n7370_), .A2(new_n7371_), .B(new_n7365_), .ZN(new_n7372_));
  OAI21_X1   g07180(.A1(new_n7372_), .A2(\asqrt[30] ), .B(new_n7334_), .ZN(new_n7373_));
  NAND2_X1   g07181(.A1(new_n7372_), .A2(\asqrt[30] ), .ZN(new_n7374_));
  AOI21_X1   g07182(.A1(new_n7373_), .A2(new_n7374_), .B(new_n5947_), .ZN(new_n7375_));
  NOR3_X1    g07183(.A1(new_n7369_), .A2(\asqrt[32] ), .A3(new_n7375_), .ZN(new_n7376_));
  OAI21_X1   g07184(.A1(new_n7369_), .A2(new_n7375_), .B(\asqrt[32] ), .ZN(new_n7377_));
  OAI21_X1   g07185(.A1(new_n7316_), .A2(new_n7376_), .B(new_n7377_), .ZN(new_n7378_));
  OAI21_X1   g07186(.A1(new_n7378_), .A2(\asqrt[33] ), .B(new_n7312_), .ZN(new_n7379_));
  NAND3_X1   g07187(.A1(new_n7373_), .A2(new_n7374_), .A3(new_n5947_), .ZN(new_n7380_));
  AOI21_X1   g07188(.A1(new_n7318_), .A2(new_n7380_), .B(new_n7375_), .ZN(new_n7381_));
  AOI21_X1   g07189(.A1(new_n7381_), .A2(new_n5643_), .B(new_n7316_), .ZN(new_n7382_));
  NAND2_X1   g07190(.A1(new_n7380_), .A2(new_n7318_), .ZN(new_n7383_));
  INV_X1     g07191(.I(new_n7375_), .ZN(new_n7384_));
  AOI21_X1   g07192(.A1(new_n7383_), .A2(new_n7384_), .B(new_n5643_), .ZN(new_n7385_));
  OAI21_X1   g07193(.A1(new_n7382_), .A2(new_n7385_), .B(\asqrt[33] ), .ZN(new_n7386_));
  NAND3_X1   g07194(.A1(new_n7379_), .A2(new_n5029_), .A3(new_n7386_), .ZN(new_n7387_));
  AOI21_X1   g07195(.A1(new_n7379_), .A2(new_n7386_), .B(new_n5029_), .ZN(new_n7388_));
  AOI21_X1   g07196(.A1(new_n7310_), .A2(new_n7387_), .B(new_n7388_), .ZN(new_n7389_));
  AOI21_X1   g07197(.A1(new_n7389_), .A2(new_n4751_), .B(new_n7307_), .ZN(new_n7390_));
  INV_X1     g07198(.I(new_n7312_), .ZN(new_n7391_));
  NOR3_X1    g07199(.A1(new_n7382_), .A2(\asqrt[33] ), .A3(new_n7385_), .ZN(new_n7392_));
  OAI21_X1   g07200(.A1(new_n7391_), .A2(new_n7392_), .B(new_n7386_), .ZN(new_n7393_));
  OAI21_X1   g07201(.A1(new_n7393_), .A2(\asqrt[34] ), .B(new_n7310_), .ZN(new_n7394_));
  NAND2_X1   g07202(.A1(new_n7393_), .A2(\asqrt[34] ), .ZN(new_n7395_));
  AOI21_X1   g07203(.A1(new_n7394_), .A2(new_n7395_), .B(new_n4751_), .ZN(new_n7396_));
  NOR3_X1    g07204(.A1(new_n7390_), .A2(\asqrt[36] ), .A3(new_n7396_), .ZN(new_n7397_));
  OAI21_X1   g07205(.A1(new_n7390_), .A2(new_n7396_), .B(\asqrt[36] ), .ZN(new_n7398_));
  OAI21_X1   g07206(.A1(new_n7304_), .A2(new_n7397_), .B(new_n7398_), .ZN(new_n7399_));
  OAI21_X1   g07207(.A1(new_n7399_), .A2(\asqrt[37] ), .B(new_n7300_), .ZN(new_n7400_));
  NAND3_X1   g07208(.A1(new_n7394_), .A2(new_n7395_), .A3(new_n4751_), .ZN(new_n7401_));
  AOI21_X1   g07209(.A1(new_n7306_), .A2(new_n7401_), .B(new_n7396_), .ZN(new_n7402_));
  AOI21_X1   g07210(.A1(new_n7402_), .A2(new_n4461_), .B(new_n7304_), .ZN(new_n7403_));
  NAND2_X1   g07211(.A1(new_n7401_), .A2(new_n7306_), .ZN(new_n7404_));
  INV_X1     g07212(.I(new_n7396_), .ZN(new_n7405_));
  AOI21_X1   g07213(.A1(new_n7404_), .A2(new_n7405_), .B(new_n4461_), .ZN(new_n7406_));
  OAI21_X1   g07214(.A1(new_n7403_), .A2(new_n7406_), .B(\asqrt[37] ), .ZN(new_n7407_));
  NAND3_X1   g07215(.A1(new_n7400_), .A2(new_n3925_), .A3(new_n7407_), .ZN(new_n7408_));
  INV_X1     g07216(.I(new_n7300_), .ZN(new_n7409_));
  NOR3_X1    g07217(.A1(new_n7403_), .A2(\asqrt[37] ), .A3(new_n7406_), .ZN(new_n7410_));
  OAI21_X1   g07218(.A1(new_n7409_), .A2(new_n7410_), .B(new_n7407_), .ZN(new_n7411_));
  NAND2_X1   g07219(.A1(new_n7411_), .A2(\asqrt[38] ), .ZN(new_n7412_));
  NOR2_X1    g07220(.A1(new_n7262_), .A2(\asqrt[62] ), .ZN(new_n7413_));
  NOR2_X1    g07221(.A1(new_n7413_), .A2(new_n7329_), .ZN(new_n7414_));
  XOR2_X1    g07222(.A1(new_n7278_), .A2(new_n6900_), .Z(new_n7415_));
  OAI21_X1   g07223(.A1(\asqrt[27] ), .A2(new_n7414_), .B(new_n7415_), .ZN(new_n7416_));
  INV_X1     g07224(.I(new_n7416_), .ZN(new_n7417_));
  AOI21_X1   g07225(.A1(new_n7247_), .A2(new_n7255_), .B(\asqrt[27] ), .ZN(new_n7418_));
  XOR2_X1    g07226(.A1(new_n7418_), .A2(new_n7054_), .Z(new_n7419_));
  INV_X1     g07227(.I(new_n7419_), .ZN(new_n7420_));
  AOI21_X1   g07228(.A1(new_n7238_), .A2(new_n7246_), .B(\asqrt[27] ), .ZN(new_n7421_));
  XOR2_X1    g07229(.A1(new_n7421_), .A2(new_n7056_), .Z(new_n7422_));
  INV_X1     g07230(.I(new_n7422_), .ZN(new_n7423_));
  NAND2_X1   g07231(.A1(new_n7242_), .A2(new_n531_), .ZN(new_n7424_));
  AOI21_X1   g07232(.A1(new_n7424_), .A2(new_n7237_), .B(\asqrt[27] ), .ZN(new_n7425_));
  XOR2_X1    g07233(.A1(new_n7425_), .A2(new_n7058_), .Z(new_n7426_));
  AOI21_X1   g07234(.A1(new_n7241_), .A2(new_n7227_), .B(\asqrt[27] ), .ZN(new_n7427_));
  XOR2_X1    g07235(.A1(new_n7427_), .A2(new_n7062_), .Z(new_n7428_));
  NAND2_X1   g07236(.A1(new_n7209_), .A2(new_n744_), .ZN(new_n7429_));
  AOI21_X1   g07237(.A1(new_n7429_), .A2(new_n7235_), .B(\asqrt[27] ), .ZN(new_n7430_));
  XOR2_X1    g07238(.A1(new_n7430_), .A2(new_n7066_), .Z(new_n7431_));
  INV_X1     g07239(.I(new_n7431_), .ZN(new_n7432_));
  AOI21_X1   g07240(.A1(new_n7207_), .A2(new_n7224_), .B(\asqrt[27] ), .ZN(new_n7433_));
  XOR2_X1    g07241(.A1(new_n7433_), .A2(new_n7069_), .Z(new_n7434_));
  INV_X1     g07242(.I(new_n7434_), .ZN(new_n7435_));
  NAND2_X1   g07243(.A1(new_n7220_), .A2(new_n1006_), .ZN(new_n7436_));
  AOI21_X1   g07244(.A1(new_n7436_), .A2(new_n7206_), .B(\asqrt[27] ), .ZN(new_n7437_));
  XOR2_X1    g07245(.A1(new_n7437_), .A2(new_n7071_), .Z(new_n7438_));
  AOI21_X1   g07246(.A1(new_n7218_), .A2(new_n7203_), .B(\asqrt[27] ), .ZN(new_n7439_));
  XOR2_X1    g07247(.A1(new_n7439_), .A2(new_n7074_), .Z(new_n7440_));
  NAND2_X1   g07248(.A1(new_n7185_), .A2(new_n1305_), .ZN(new_n7441_));
  AOI21_X1   g07249(.A1(new_n7441_), .A2(new_n7217_), .B(\asqrt[27] ), .ZN(new_n7442_));
  XOR2_X1    g07250(.A1(new_n7442_), .A2(new_n7078_), .Z(new_n7443_));
  INV_X1     g07251(.I(new_n7443_), .ZN(new_n7444_));
  AOI21_X1   g07252(.A1(new_n7183_), .A2(new_n7200_), .B(\asqrt[27] ), .ZN(new_n7445_));
  XOR2_X1    g07253(.A1(new_n7445_), .A2(new_n7081_), .Z(new_n7446_));
  INV_X1     g07254(.I(new_n7446_), .ZN(new_n7447_));
  NAND2_X1   g07255(.A1(new_n7196_), .A2(new_n1632_), .ZN(new_n7448_));
  AOI21_X1   g07256(.A1(new_n7448_), .A2(new_n7182_), .B(\asqrt[27] ), .ZN(new_n7449_));
  XOR2_X1    g07257(.A1(new_n7449_), .A2(new_n7083_), .Z(new_n7450_));
  AOI21_X1   g07258(.A1(new_n7194_), .A2(new_n7179_), .B(\asqrt[27] ), .ZN(new_n7451_));
  XOR2_X1    g07259(.A1(new_n7451_), .A2(new_n7086_), .Z(new_n7452_));
  NAND2_X1   g07260(.A1(new_n7161_), .A2(new_n1953_), .ZN(new_n7453_));
  AOI21_X1   g07261(.A1(new_n7453_), .A2(new_n7193_), .B(\asqrt[27] ), .ZN(new_n7454_));
  XOR2_X1    g07262(.A1(new_n7454_), .A2(new_n7090_), .Z(new_n7455_));
  INV_X1     g07263(.I(new_n7455_), .ZN(new_n7456_));
  AOI21_X1   g07264(.A1(new_n7159_), .A2(new_n7176_), .B(\asqrt[27] ), .ZN(new_n7457_));
  XOR2_X1    g07265(.A1(new_n7457_), .A2(new_n7093_), .Z(new_n7458_));
  INV_X1     g07266(.I(new_n7458_), .ZN(new_n7459_));
  NAND2_X1   g07267(.A1(new_n7172_), .A2(new_n2332_), .ZN(new_n7460_));
  AOI21_X1   g07268(.A1(new_n7460_), .A2(new_n7158_), .B(\asqrt[27] ), .ZN(new_n7461_));
  XOR2_X1    g07269(.A1(new_n7461_), .A2(new_n7095_), .Z(new_n7462_));
  AOI21_X1   g07270(.A1(new_n7170_), .A2(new_n7155_), .B(\asqrt[27] ), .ZN(new_n7463_));
  XOR2_X1    g07271(.A1(new_n7463_), .A2(new_n7098_), .Z(new_n7464_));
  NAND2_X1   g07272(.A1(new_n7137_), .A2(new_n2749_), .ZN(new_n7465_));
  AOI21_X1   g07273(.A1(new_n7465_), .A2(new_n7169_), .B(\asqrt[27] ), .ZN(new_n7466_));
  XOR2_X1    g07274(.A1(new_n7466_), .A2(new_n7102_), .Z(new_n7467_));
  INV_X1     g07275(.I(new_n7467_), .ZN(new_n7468_));
  AOI21_X1   g07276(.A1(new_n7135_), .A2(new_n7152_), .B(\asqrt[27] ), .ZN(new_n7469_));
  XOR2_X1    g07277(.A1(new_n7469_), .A2(new_n7105_), .Z(new_n7470_));
  INV_X1     g07278(.I(new_n7470_), .ZN(new_n7471_));
  NAND2_X1   g07279(.A1(new_n7148_), .A2(new_n3195_), .ZN(new_n7472_));
  AOI21_X1   g07280(.A1(new_n7472_), .A2(new_n7134_), .B(\asqrt[27] ), .ZN(new_n7473_));
  XOR2_X1    g07281(.A1(new_n7473_), .A2(new_n7107_), .Z(new_n7474_));
  AOI21_X1   g07282(.A1(new_n7146_), .A2(new_n7131_), .B(\asqrt[27] ), .ZN(new_n7475_));
  XOR2_X1    g07283(.A1(new_n7475_), .A2(new_n7110_), .Z(new_n7476_));
  NAND2_X1   g07284(.A1(new_n7121_), .A2(new_n3681_), .ZN(new_n7477_));
  AOI21_X1   g07285(.A1(new_n7477_), .A2(new_n7145_), .B(\asqrt[27] ), .ZN(new_n7478_));
  XOR2_X1    g07286(.A1(new_n7478_), .A2(new_n7114_), .Z(new_n7479_));
  INV_X1     g07287(.I(new_n7479_), .ZN(new_n7480_));
  AOI21_X1   g07288(.A1(new_n7119_), .A2(new_n7128_), .B(\asqrt[27] ), .ZN(new_n7481_));
  XOR2_X1    g07289(.A1(new_n7481_), .A2(new_n7117_), .Z(new_n7482_));
  INV_X1     g07290(.I(new_n7482_), .ZN(new_n7483_));
  AOI21_X1   g07291(.A1(new_n7400_), .A2(new_n7407_), .B(new_n3925_), .ZN(new_n7484_));
  AOI21_X1   g07292(.A1(new_n7298_), .A2(new_n7408_), .B(new_n7484_), .ZN(new_n7485_));
  AOI21_X1   g07293(.A1(new_n7485_), .A2(new_n3681_), .B(new_n7483_), .ZN(new_n7486_));
  OAI21_X1   g07294(.A1(new_n7411_), .A2(\asqrt[38] ), .B(new_n7298_), .ZN(new_n7487_));
  AOI21_X1   g07295(.A1(new_n7487_), .A2(new_n7412_), .B(new_n3681_), .ZN(new_n7488_));
  NOR3_X1    g07296(.A1(new_n7486_), .A2(\asqrt[40] ), .A3(new_n7488_), .ZN(new_n7489_));
  OAI21_X1   g07297(.A1(new_n7486_), .A2(new_n7488_), .B(\asqrt[40] ), .ZN(new_n7490_));
  OAI21_X1   g07298(.A1(new_n7480_), .A2(new_n7489_), .B(new_n7490_), .ZN(new_n7491_));
  OAI21_X1   g07299(.A1(new_n7491_), .A2(\asqrt[41] ), .B(new_n7476_), .ZN(new_n7492_));
  NAND3_X1   g07300(.A1(new_n7487_), .A2(new_n7412_), .A3(new_n3681_), .ZN(new_n7493_));
  AOI21_X1   g07301(.A1(new_n7482_), .A2(new_n7493_), .B(new_n7488_), .ZN(new_n7494_));
  AOI21_X1   g07302(.A1(new_n7494_), .A2(new_n3427_), .B(new_n7480_), .ZN(new_n7495_));
  NAND2_X1   g07303(.A1(new_n7493_), .A2(new_n7482_), .ZN(new_n7496_));
  INV_X1     g07304(.I(new_n7488_), .ZN(new_n7497_));
  AOI21_X1   g07305(.A1(new_n7496_), .A2(new_n7497_), .B(new_n3427_), .ZN(new_n7498_));
  OAI21_X1   g07306(.A1(new_n7495_), .A2(new_n7498_), .B(\asqrt[41] ), .ZN(new_n7499_));
  NAND3_X1   g07307(.A1(new_n7492_), .A2(new_n2960_), .A3(new_n7499_), .ZN(new_n7500_));
  AOI21_X1   g07308(.A1(new_n7492_), .A2(new_n7499_), .B(new_n2960_), .ZN(new_n7501_));
  AOI21_X1   g07309(.A1(new_n7474_), .A2(new_n7500_), .B(new_n7501_), .ZN(new_n7502_));
  AOI21_X1   g07310(.A1(new_n7502_), .A2(new_n2749_), .B(new_n7471_), .ZN(new_n7503_));
  INV_X1     g07311(.I(new_n7476_), .ZN(new_n7504_));
  NOR3_X1    g07312(.A1(new_n7495_), .A2(\asqrt[41] ), .A3(new_n7498_), .ZN(new_n7505_));
  OAI21_X1   g07313(.A1(new_n7504_), .A2(new_n7505_), .B(new_n7499_), .ZN(new_n7506_));
  OAI21_X1   g07314(.A1(new_n7506_), .A2(\asqrt[42] ), .B(new_n7474_), .ZN(new_n7507_));
  NAND2_X1   g07315(.A1(new_n7506_), .A2(\asqrt[42] ), .ZN(new_n7508_));
  AOI21_X1   g07316(.A1(new_n7507_), .A2(new_n7508_), .B(new_n2749_), .ZN(new_n7509_));
  NOR3_X1    g07317(.A1(new_n7503_), .A2(\asqrt[44] ), .A3(new_n7509_), .ZN(new_n7510_));
  OAI21_X1   g07318(.A1(new_n7503_), .A2(new_n7509_), .B(\asqrt[44] ), .ZN(new_n7511_));
  OAI21_X1   g07319(.A1(new_n7468_), .A2(new_n7510_), .B(new_n7511_), .ZN(new_n7512_));
  OAI21_X1   g07320(.A1(new_n7512_), .A2(\asqrt[45] ), .B(new_n7464_), .ZN(new_n7513_));
  NAND3_X1   g07321(.A1(new_n7507_), .A2(new_n7508_), .A3(new_n2749_), .ZN(new_n7514_));
  AOI21_X1   g07322(.A1(new_n7470_), .A2(new_n7514_), .B(new_n7509_), .ZN(new_n7515_));
  AOI21_X1   g07323(.A1(new_n7515_), .A2(new_n2531_), .B(new_n7468_), .ZN(new_n7516_));
  NAND2_X1   g07324(.A1(new_n7514_), .A2(new_n7470_), .ZN(new_n7517_));
  INV_X1     g07325(.I(new_n7509_), .ZN(new_n7518_));
  AOI21_X1   g07326(.A1(new_n7517_), .A2(new_n7518_), .B(new_n2531_), .ZN(new_n7519_));
  OAI21_X1   g07327(.A1(new_n7516_), .A2(new_n7519_), .B(\asqrt[45] ), .ZN(new_n7520_));
  NAND3_X1   g07328(.A1(new_n7513_), .A2(new_n2134_), .A3(new_n7520_), .ZN(new_n7521_));
  AOI21_X1   g07329(.A1(new_n7513_), .A2(new_n7520_), .B(new_n2134_), .ZN(new_n7522_));
  AOI21_X1   g07330(.A1(new_n7462_), .A2(new_n7521_), .B(new_n7522_), .ZN(new_n7523_));
  AOI21_X1   g07331(.A1(new_n7523_), .A2(new_n1953_), .B(new_n7459_), .ZN(new_n7524_));
  INV_X1     g07332(.I(new_n7464_), .ZN(new_n7525_));
  NOR3_X1    g07333(.A1(new_n7516_), .A2(\asqrt[45] ), .A3(new_n7519_), .ZN(new_n7526_));
  OAI21_X1   g07334(.A1(new_n7525_), .A2(new_n7526_), .B(new_n7520_), .ZN(new_n7527_));
  OAI21_X1   g07335(.A1(new_n7527_), .A2(\asqrt[46] ), .B(new_n7462_), .ZN(new_n7528_));
  NAND2_X1   g07336(.A1(new_n7527_), .A2(\asqrt[46] ), .ZN(new_n7529_));
  AOI21_X1   g07337(.A1(new_n7528_), .A2(new_n7529_), .B(new_n1953_), .ZN(new_n7530_));
  NOR3_X1    g07338(.A1(new_n7524_), .A2(\asqrt[48] ), .A3(new_n7530_), .ZN(new_n7531_));
  OAI21_X1   g07339(.A1(new_n7524_), .A2(new_n7530_), .B(\asqrt[48] ), .ZN(new_n7532_));
  OAI21_X1   g07340(.A1(new_n7456_), .A2(new_n7531_), .B(new_n7532_), .ZN(new_n7533_));
  OAI21_X1   g07341(.A1(new_n7533_), .A2(\asqrt[49] ), .B(new_n7452_), .ZN(new_n7534_));
  NAND3_X1   g07342(.A1(new_n7528_), .A2(new_n7529_), .A3(new_n1953_), .ZN(new_n7535_));
  AOI21_X1   g07343(.A1(new_n7458_), .A2(new_n7535_), .B(new_n7530_), .ZN(new_n7536_));
  AOI21_X1   g07344(.A1(new_n7536_), .A2(new_n1778_), .B(new_n7456_), .ZN(new_n7537_));
  NAND2_X1   g07345(.A1(new_n7535_), .A2(new_n7458_), .ZN(new_n7538_));
  INV_X1     g07346(.I(new_n7530_), .ZN(new_n7539_));
  AOI21_X1   g07347(.A1(new_n7538_), .A2(new_n7539_), .B(new_n1778_), .ZN(new_n7540_));
  OAI21_X1   g07348(.A1(new_n7537_), .A2(new_n7540_), .B(\asqrt[49] ), .ZN(new_n7541_));
  NAND3_X1   g07349(.A1(new_n7534_), .A2(new_n1463_), .A3(new_n7541_), .ZN(new_n7542_));
  AOI21_X1   g07350(.A1(new_n7534_), .A2(new_n7541_), .B(new_n1463_), .ZN(new_n7543_));
  AOI21_X1   g07351(.A1(new_n7450_), .A2(new_n7542_), .B(new_n7543_), .ZN(new_n7544_));
  AOI21_X1   g07352(.A1(new_n7544_), .A2(new_n1305_), .B(new_n7447_), .ZN(new_n7545_));
  INV_X1     g07353(.I(new_n7452_), .ZN(new_n7546_));
  NOR3_X1    g07354(.A1(new_n7537_), .A2(\asqrt[49] ), .A3(new_n7540_), .ZN(new_n7547_));
  OAI21_X1   g07355(.A1(new_n7546_), .A2(new_n7547_), .B(new_n7541_), .ZN(new_n7548_));
  OAI21_X1   g07356(.A1(new_n7548_), .A2(\asqrt[50] ), .B(new_n7450_), .ZN(new_n7549_));
  NAND2_X1   g07357(.A1(new_n7548_), .A2(\asqrt[50] ), .ZN(new_n7550_));
  AOI21_X1   g07358(.A1(new_n7549_), .A2(new_n7550_), .B(new_n1305_), .ZN(new_n7551_));
  NOR3_X1    g07359(.A1(new_n7545_), .A2(\asqrt[52] ), .A3(new_n7551_), .ZN(new_n7552_));
  OAI21_X1   g07360(.A1(new_n7545_), .A2(new_n7551_), .B(\asqrt[52] ), .ZN(new_n7553_));
  OAI21_X1   g07361(.A1(new_n7444_), .A2(new_n7552_), .B(new_n7553_), .ZN(new_n7554_));
  OAI21_X1   g07362(.A1(new_n7554_), .A2(\asqrt[53] ), .B(new_n7440_), .ZN(new_n7555_));
  NAND3_X1   g07363(.A1(new_n7549_), .A2(new_n7550_), .A3(new_n1305_), .ZN(new_n7556_));
  AOI21_X1   g07364(.A1(new_n7446_), .A2(new_n7556_), .B(new_n7551_), .ZN(new_n7557_));
  AOI21_X1   g07365(.A1(new_n7557_), .A2(new_n1150_), .B(new_n7444_), .ZN(new_n7558_));
  NAND2_X1   g07366(.A1(new_n7556_), .A2(new_n7446_), .ZN(new_n7559_));
  INV_X1     g07367(.I(new_n7551_), .ZN(new_n7560_));
  AOI21_X1   g07368(.A1(new_n7559_), .A2(new_n7560_), .B(new_n1150_), .ZN(new_n7561_));
  OAI21_X1   g07369(.A1(new_n7558_), .A2(new_n7561_), .B(\asqrt[53] ), .ZN(new_n7562_));
  NAND3_X1   g07370(.A1(new_n7555_), .A2(new_n860_), .A3(new_n7562_), .ZN(new_n7563_));
  AOI21_X1   g07371(.A1(new_n7555_), .A2(new_n7562_), .B(new_n860_), .ZN(new_n7564_));
  AOI21_X1   g07372(.A1(new_n7438_), .A2(new_n7563_), .B(new_n7564_), .ZN(new_n7565_));
  AOI21_X1   g07373(.A1(new_n7565_), .A2(new_n744_), .B(new_n7435_), .ZN(new_n7566_));
  INV_X1     g07374(.I(new_n7440_), .ZN(new_n7567_));
  NOR3_X1    g07375(.A1(new_n7558_), .A2(\asqrt[53] ), .A3(new_n7561_), .ZN(new_n7568_));
  OAI21_X1   g07376(.A1(new_n7567_), .A2(new_n7568_), .B(new_n7562_), .ZN(new_n7569_));
  OAI21_X1   g07377(.A1(new_n7569_), .A2(\asqrt[54] ), .B(new_n7438_), .ZN(new_n7570_));
  NAND2_X1   g07378(.A1(new_n7569_), .A2(\asqrt[54] ), .ZN(new_n7571_));
  AOI21_X1   g07379(.A1(new_n7570_), .A2(new_n7571_), .B(new_n744_), .ZN(new_n7572_));
  NOR3_X1    g07380(.A1(new_n7566_), .A2(\asqrt[56] ), .A3(new_n7572_), .ZN(new_n7573_));
  OAI21_X1   g07381(.A1(new_n7566_), .A2(new_n7572_), .B(\asqrt[56] ), .ZN(new_n7574_));
  OAI21_X1   g07382(.A1(new_n7432_), .A2(new_n7573_), .B(new_n7574_), .ZN(new_n7575_));
  OAI21_X1   g07383(.A1(new_n7575_), .A2(\asqrt[57] ), .B(new_n7428_), .ZN(new_n7576_));
  NAND3_X1   g07384(.A1(new_n7570_), .A2(new_n7571_), .A3(new_n744_), .ZN(new_n7577_));
  AOI21_X1   g07385(.A1(new_n7434_), .A2(new_n7577_), .B(new_n7572_), .ZN(new_n7578_));
  AOI21_X1   g07386(.A1(new_n7578_), .A2(new_n634_), .B(new_n7432_), .ZN(new_n7579_));
  NAND2_X1   g07387(.A1(new_n7577_), .A2(new_n7434_), .ZN(new_n7580_));
  INV_X1     g07388(.I(new_n7572_), .ZN(new_n7581_));
  AOI21_X1   g07389(.A1(new_n7580_), .A2(new_n7581_), .B(new_n634_), .ZN(new_n7582_));
  OAI21_X1   g07390(.A1(new_n7579_), .A2(new_n7582_), .B(\asqrt[57] ), .ZN(new_n7583_));
  NAND3_X1   g07391(.A1(new_n7576_), .A2(new_n423_), .A3(new_n7583_), .ZN(new_n7584_));
  AOI21_X1   g07392(.A1(new_n7576_), .A2(new_n7583_), .B(new_n423_), .ZN(new_n7585_));
  AOI21_X1   g07393(.A1(new_n7426_), .A2(new_n7584_), .B(new_n7585_), .ZN(new_n7586_));
  AOI21_X1   g07394(.A1(new_n7586_), .A2(new_n337_), .B(new_n7423_), .ZN(new_n7587_));
  NOR2_X1    g07395(.A1(new_n7586_), .A2(new_n337_), .ZN(new_n7588_));
  NOR3_X1    g07396(.A1(new_n7587_), .A2(new_n7588_), .A3(\asqrt[60] ), .ZN(new_n7589_));
  OAI21_X1   g07397(.A1(new_n7587_), .A2(new_n7588_), .B(\asqrt[60] ), .ZN(new_n7590_));
  OAI21_X1   g07398(.A1(new_n7420_), .A2(new_n7589_), .B(new_n7590_), .ZN(new_n7591_));
  NAND2_X1   g07399(.A1(new_n7591_), .A2(\asqrt[61] ), .ZN(new_n7592_));
  AOI21_X1   g07400(.A1(new_n7263_), .A2(new_n7269_), .B(\asqrt[27] ), .ZN(new_n7593_));
  XOR2_X1    g07401(.A1(new_n7593_), .A2(new_n7050_), .Z(new_n7594_));
  OAI21_X1   g07402(.A1(new_n7591_), .A2(\asqrt[61] ), .B(new_n7594_), .ZN(new_n7595_));
  NAND2_X1   g07403(.A1(new_n7595_), .A2(new_n7592_), .ZN(new_n7596_));
  INV_X1     g07404(.I(new_n7428_), .ZN(new_n7597_));
  NOR3_X1    g07405(.A1(new_n7579_), .A2(\asqrt[57] ), .A3(new_n7582_), .ZN(new_n7598_));
  OAI21_X1   g07406(.A1(new_n7597_), .A2(new_n7598_), .B(new_n7583_), .ZN(new_n7599_));
  OAI21_X1   g07407(.A1(new_n7599_), .A2(\asqrt[58] ), .B(new_n7426_), .ZN(new_n7600_));
  NOR2_X1    g07408(.A1(new_n7598_), .A2(new_n7597_), .ZN(new_n7601_));
  INV_X1     g07409(.I(new_n7583_), .ZN(new_n7602_));
  OAI21_X1   g07410(.A1(new_n7601_), .A2(new_n7602_), .B(\asqrt[58] ), .ZN(new_n7603_));
  NAND3_X1   g07411(.A1(new_n7600_), .A2(new_n337_), .A3(new_n7603_), .ZN(new_n7604_));
  NAND2_X1   g07412(.A1(new_n7604_), .A2(new_n7422_), .ZN(new_n7605_));
  INV_X1     g07413(.I(new_n7426_), .ZN(new_n7606_));
  NOR2_X1    g07414(.A1(new_n7601_), .A2(new_n7602_), .ZN(new_n7607_));
  AOI21_X1   g07415(.A1(new_n7607_), .A2(new_n423_), .B(new_n7606_), .ZN(new_n7608_));
  OAI21_X1   g07416(.A1(new_n7608_), .A2(new_n7585_), .B(\asqrt[59] ), .ZN(new_n7609_));
  NAND3_X1   g07417(.A1(new_n7605_), .A2(new_n266_), .A3(new_n7609_), .ZN(new_n7610_));
  NAND2_X1   g07418(.A1(new_n7610_), .A2(new_n7419_), .ZN(new_n7611_));
  AOI21_X1   g07419(.A1(new_n7611_), .A2(new_n7590_), .B(new_n239_), .ZN(new_n7612_));
  AOI21_X1   g07420(.A1(new_n7605_), .A2(new_n7609_), .B(new_n266_), .ZN(new_n7613_));
  AOI21_X1   g07421(.A1(new_n7419_), .A2(new_n7610_), .B(new_n7613_), .ZN(new_n7614_));
  INV_X1     g07422(.I(new_n7594_), .ZN(new_n7615_));
  AOI21_X1   g07423(.A1(new_n7614_), .A2(new_n239_), .B(new_n7615_), .ZN(new_n7616_));
  OAI21_X1   g07424(.A1(new_n7616_), .A2(new_n7612_), .B(new_n201_), .ZN(new_n7617_));
  NAND3_X1   g07425(.A1(new_n7595_), .A2(new_n7592_), .A3(\asqrt[62] ), .ZN(new_n7618_));
  NOR2_X1    g07426(.A1(new_n7261_), .A2(new_n7270_), .ZN(new_n7619_));
  NOR2_X1    g07427(.A1(\asqrt[27] ), .A2(new_n7619_), .ZN(new_n7620_));
  XOR2_X1    g07428(.A1(new_n7620_), .A2(new_n7259_), .Z(new_n7621_));
  INV_X1     g07429(.I(new_n7621_), .ZN(new_n7622_));
  AOI22_X1   g07430(.A1(new_n7618_), .A2(new_n7617_), .B1(new_n7596_), .B2(new_n7622_), .ZN(new_n7623_));
  NOR2_X1    g07431(.A1(new_n7281_), .A2(new_n7047_), .ZN(new_n7624_));
  OAI21_X1   g07432(.A1(\asqrt[27] ), .A2(new_n7624_), .B(new_n7288_), .ZN(new_n7625_));
  INV_X1     g07433(.I(new_n7625_), .ZN(new_n7626_));
  OAI21_X1   g07434(.A1(new_n7623_), .A2(new_n7417_), .B(new_n7626_), .ZN(new_n7627_));
  OAI21_X1   g07435(.A1(new_n7596_), .A2(\asqrt[62] ), .B(new_n7621_), .ZN(new_n7628_));
  NAND2_X1   g07436(.A1(new_n7596_), .A2(\asqrt[62] ), .ZN(new_n7629_));
  NAND3_X1   g07437(.A1(new_n7628_), .A2(new_n7629_), .A3(new_n7417_), .ZN(new_n7630_));
  NAND2_X1   g07438(.A1(new_n7281_), .A2(new_n7046_), .ZN(new_n7631_));
  NAND2_X1   g07439(.A1(new_n7326_), .A2(new_n7047_), .ZN(new_n7632_));
  AOI21_X1   g07440(.A1(new_n7631_), .A2(new_n7632_), .B(new_n193_), .ZN(new_n7633_));
  OAI21_X1   g07441(.A1(\asqrt[27] ), .A2(new_n7047_), .B(new_n7633_), .ZN(new_n7634_));
  NOR2_X1    g07442(.A1(new_n7294_), .A2(new_n7046_), .ZN(new_n7635_));
  NAND4_X1   g07443(.A1(new_n7285_), .A2(new_n193_), .A3(new_n7288_), .A4(new_n7635_), .ZN(new_n7636_));
  NAND2_X1   g07444(.A1(new_n7634_), .A2(new_n7636_), .ZN(new_n7637_));
  INV_X1     g07445(.I(new_n7637_), .ZN(new_n7638_));
  NAND4_X1   g07446(.A1(new_n7627_), .A2(new_n193_), .A3(new_n7630_), .A4(new_n7638_), .ZN(\asqrt[26] ));
  AOI21_X1   g07447(.A1(new_n7408_), .A2(new_n7412_), .B(\asqrt[26] ), .ZN(new_n7640_));
  XOR2_X1    g07448(.A1(new_n7640_), .A2(new_n7298_), .Z(new_n7641_));
  XOR2_X1    g07449(.A1(new_n7399_), .A2(\asqrt[37] ), .Z(new_n7642_));
  NOR2_X1    g07450(.A1(\asqrt[26] ), .A2(new_n7642_), .ZN(new_n7643_));
  XOR2_X1    g07451(.A1(new_n7643_), .A2(new_n7300_), .Z(new_n7644_));
  NOR2_X1    g07452(.A1(new_n7397_), .A2(new_n7406_), .ZN(new_n7645_));
  NOR2_X1    g07453(.A1(\asqrt[26] ), .A2(new_n7645_), .ZN(new_n7646_));
  XOR2_X1    g07454(.A1(new_n7646_), .A2(new_n7303_), .Z(new_n7647_));
  AOI21_X1   g07455(.A1(new_n7401_), .A2(new_n7405_), .B(\asqrt[26] ), .ZN(new_n7648_));
  XOR2_X1    g07456(.A1(new_n7648_), .A2(new_n7306_), .Z(new_n7649_));
  INV_X1     g07457(.I(new_n7649_), .ZN(new_n7650_));
  AOI21_X1   g07458(.A1(new_n7387_), .A2(new_n7395_), .B(\asqrt[26] ), .ZN(new_n7651_));
  XOR2_X1    g07459(.A1(new_n7651_), .A2(new_n7310_), .Z(new_n7652_));
  INV_X1     g07460(.I(new_n7652_), .ZN(new_n7653_));
  XOR2_X1    g07461(.A1(new_n7378_), .A2(\asqrt[33] ), .Z(new_n7654_));
  NOR2_X1    g07462(.A1(\asqrt[26] ), .A2(new_n7654_), .ZN(new_n7655_));
  XOR2_X1    g07463(.A1(new_n7655_), .A2(new_n7312_), .Z(new_n7656_));
  NOR2_X1    g07464(.A1(new_n7376_), .A2(new_n7385_), .ZN(new_n7657_));
  NOR2_X1    g07465(.A1(\asqrt[26] ), .A2(new_n7657_), .ZN(new_n7658_));
  XOR2_X1    g07466(.A1(new_n7658_), .A2(new_n7315_), .Z(new_n7659_));
  AOI21_X1   g07467(.A1(new_n7380_), .A2(new_n7384_), .B(\asqrt[26] ), .ZN(new_n7660_));
  XOR2_X1    g07468(.A1(new_n7660_), .A2(new_n7318_), .Z(new_n7661_));
  INV_X1     g07469(.I(new_n7661_), .ZN(new_n7662_));
  AOI21_X1   g07470(.A1(new_n7366_), .A2(new_n7374_), .B(\asqrt[26] ), .ZN(new_n7663_));
  XOR2_X1    g07471(.A1(new_n7663_), .A2(new_n7334_), .Z(new_n7664_));
  INV_X1     g07472(.I(new_n7664_), .ZN(new_n7665_));
  AOI21_X1   g07473(.A1(new_n7357_), .A2(new_n7365_), .B(\asqrt[26] ), .ZN(new_n7666_));
  XOR2_X1    g07474(.A1(new_n7666_), .A2(new_n7342_), .Z(new_n7667_));
  NAND2_X1   g07475(.A1(\asqrt[27] ), .A2(new_n7343_), .ZN(new_n7668_));
  NOR2_X1    g07476(.A1(new_n7354_), .A2(\a[54] ), .ZN(new_n7669_));
  AOI22_X1   g07477(.A1(new_n7668_), .A2(new_n7354_), .B1(\asqrt[27] ), .B2(new_n7669_), .ZN(new_n7670_));
  AOI21_X1   g07478(.A1(\asqrt[27] ), .A2(\a[54] ), .B(new_n7351_), .ZN(new_n7671_));
  NOR2_X1    g07479(.A1(new_n7361_), .A2(new_n7671_), .ZN(new_n7672_));
  NOR2_X1    g07480(.A1(\asqrt[26] ), .A2(new_n7672_), .ZN(new_n7673_));
  XOR2_X1    g07481(.A1(new_n7673_), .A2(new_n7670_), .Z(new_n7674_));
  NOR2_X1    g07482(.A1(new_n7616_), .A2(new_n7612_), .ZN(new_n7675_));
  AOI21_X1   g07483(.A1(new_n7595_), .A2(new_n7592_), .B(\asqrt[62] ), .ZN(new_n7676_));
  NOR3_X1    g07484(.A1(new_n7616_), .A2(new_n201_), .A3(new_n7612_), .ZN(new_n7677_));
  OAI22_X1   g07485(.A1(new_n7676_), .A2(new_n7677_), .B1(new_n7675_), .B2(new_n7621_), .ZN(new_n7678_));
  AOI21_X1   g07486(.A1(new_n7678_), .A2(new_n7416_), .B(new_n7625_), .ZN(new_n7679_));
  AOI21_X1   g07487(.A1(new_n7675_), .A2(new_n201_), .B(new_n7622_), .ZN(new_n7680_));
  NOR2_X1    g07488(.A1(new_n7675_), .A2(new_n201_), .ZN(new_n7681_));
  NOR3_X1    g07489(.A1(new_n7680_), .A2(new_n7681_), .A3(new_n7416_), .ZN(new_n7682_));
  NOR3_X1    g07490(.A1(new_n7679_), .A2(\asqrt[63] ), .A3(new_n7682_), .ZN(new_n7683_));
  NAND4_X1   g07491(.A1(new_n7683_), .A2(\asqrt[27] ), .A3(new_n7634_), .A4(new_n7636_), .ZN(new_n7684_));
  NAND2_X1   g07492(.A1(\asqrt[26] ), .A2(new_n7344_), .ZN(new_n7685_));
  AOI21_X1   g07493(.A1(new_n7684_), .A2(new_n7685_), .B(\a[54] ), .ZN(new_n7686_));
  NAND2_X1   g07494(.A1(new_n7627_), .A2(new_n193_), .ZN(new_n7687_));
  NAND3_X1   g07495(.A1(new_n7634_), .A2(new_n7636_), .A3(\asqrt[27] ), .ZN(new_n7688_));
  NOR3_X1    g07496(.A1(new_n7687_), .A2(new_n7682_), .A3(new_n7688_), .ZN(new_n7689_));
  NOR4_X1    g07497(.A1(new_n7679_), .A2(\asqrt[63] ), .A3(new_n7682_), .A4(new_n7637_), .ZN(new_n7690_));
  NOR2_X1    g07498(.A1(new_n7690_), .A2(new_n7346_), .ZN(new_n7691_));
  NOR3_X1    g07499(.A1(new_n7691_), .A2(new_n7689_), .A3(new_n7343_), .ZN(new_n7692_));
  OR2_X2     g07500(.A1(new_n7686_), .A2(new_n7692_), .Z(new_n7693_));
  NOR2_X1    g07501(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n7694_));
  INV_X1     g07502(.I(new_n7694_), .ZN(new_n7695_));
  NAND3_X1   g07503(.A1(\asqrt[26] ), .A2(\a[52] ), .A3(new_n7695_), .ZN(new_n7696_));
  INV_X1     g07504(.I(\a[52] ), .ZN(new_n7697_));
  OAI21_X1   g07505(.A1(\asqrt[26] ), .A2(new_n7697_), .B(new_n7694_), .ZN(new_n7698_));
  AOI21_X1   g07506(.A1(new_n7698_), .A2(new_n7696_), .B(new_n7331_), .ZN(new_n7699_));
  NOR3_X1    g07507(.A1(new_n7327_), .A2(\asqrt[63] ), .A3(new_n7330_), .ZN(new_n7700_));
  NAND2_X1   g07508(.A1(new_n7694_), .A2(new_n7697_), .ZN(new_n7701_));
  NAND3_X1   g07509(.A1(new_n7291_), .A2(new_n7293_), .A3(new_n7701_), .ZN(new_n7702_));
  NAND2_X1   g07510(.A1(new_n7700_), .A2(new_n7702_), .ZN(new_n7703_));
  NAND3_X1   g07511(.A1(\asqrt[26] ), .A2(\a[52] ), .A3(new_n7703_), .ZN(new_n7704_));
  INV_X1     g07512(.I(\a[53] ), .ZN(new_n7705_));
  NAND3_X1   g07513(.A1(\asqrt[26] ), .A2(new_n7697_), .A3(new_n7705_), .ZN(new_n7706_));
  OAI21_X1   g07514(.A1(new_n7690_), .A2(\a[52] ), .B(\a[53] ), .ZN(new_n7707_));
  NAND3_X1   g07515(.A1(new_n7704_), .A2(new_n7707_), .A3(new_n7706_), .ZN(new_n7708_));
  NOR3_X1    g07516(.A1(new_n7708_), .A2(new_n7699_), .A3(\asqrt[28] ), .ZN(new_n7709_));
  OAI21_X1   g07517(.A1(new_n7708_), .A2(new_n7699_), .B(\asqrt[28] ), .ZN(new_n7710_));
  OAI21_X1   g07518(.A1(new_n7693_), .A2(new_n7709_), .B(new_n7710_), .ZN(new_n7711_));
  OAI21_X1   g07519(.A1(new_n7711_), .A2(\asqrt[29] ), .B(new_n7674_), .ZN(new_n7712_));
  NAND2_X1   g07520(.A1(new_n7711_), .A2(\asqrt[29] ), .ZN(new_n7713_));
  NAND3_X1   g07521(.A1(new_n7712_), .A2(new_n7713_), .A3(new_n6275_), .ZN(new_n7714_));
  AOI21_X1   g07522(.A1(new_n7712_), .A2(new_n7713_), .B(new_n6275_), .ZN(new_n7715_));
  AOI21_X1   g07523(.A1(new_n7667_), .A2(new_n7714_), .B(new_n7715_), .ZN(new_n7716_));
  AOI21_X1   g07524(.A1(new_n7716_), .A2(new_n5947_), .B(new_n7665_), .ZN(new_n7717_));
  NAND2_X1   g07525(.A1(new_n7714_), .A2(new_n7667_), .ZN(new_n7718_));
  INV_X1     g07526(.I(new_n7674_), .ZN(new_n7719_));
  NOR2_X1    g07527(.A1(new_n7686_), .A2(new_n7692_), .ZN(new_n7720_));
  NOR3_X1    g07528(.A1(new_n7690_), .A2(new_n7697_), .A3(new_n7694_), .ZN(new_n7721_));
  AOI21_X1   g07529(.A1(new_n7690_), .A2(\a[52] ), .B(new_n7695_), .ZN(new_n7722_));
  OAI21_X1   g07530(.A1(new_n7721_), .A2(new_n7722_), .B(\asqrt[27] ), .ZN(new_n7723_));
  INV_X1     g07531(.I(new_n7703_), .ZN(new_n7724_));
  NOR3_X1    g07532(.A1(new_n7690_), .A2(new_n7697_), .A3(new_n7724_), .ZN(new_n7725_));
  NOR3_X1    g07533(.A1(new_n7690_), .A2(\a[52] ), .A3(\a[53] ), .ZN(new_n7726_));
  AOI21_X1   g07534(.A1(\asqrt[26] ), .A2(new_n7697_), .B(new_n7705_), .ZN(new_n7727_));
  NOR3_X1    g07535(.A1(new_n7725_), .A2(new_n7726_), .A3(new_n7727_), .ZN(new_n7728_));
  NAND3_X1   g07536(.A1(new_n7728_), .A2(new_n7723_), .A3(new_n6966_), .ZN(new_n7729_));
  AOI21_X1   g07537(.A1(new_n7728_), .A2(new_n7723_), .B(new_n6966_), .ZN(new_n7730_));
  AOI21_X1   g07538(.A1(new_n7720_), .A2(new_n7729_), .B(new_n7730_), .ZN(new_n7731_));
  AOI21_X1   g07539(.A1(new_n7731_), .A2(new_n6636_), .B(new_n7719_), .ZN(new_n7732_));
  NAND2_X1   g07540(.A1(new_n7729_), .A2(new_n7720_), .ZN(new_n7733_));
  AOI21_X1   g07541(.A1(new_n7733_), .A2(new_n7710_), .B(new_n6636_), .ZN(new_n7734_));
  OAI21_X1   g07542(.A1(new_n7732_), .A2(new_n7734_), .B(\asqrt[30] ), .ZN(new_n7735_));
  AOI21_X1   g07543(.A1(new_n7718_), .A2(new_n7735_), .B(new_n5947_), .ZN(new_n7736_));
  NOR3_X1    g07544(.A1(new_n7717_), .A2(\asqrt[32] ), .A3(new_n7736_), .ZN(new_n7737_));
  OAI21_X1   g07545(.A1(new_n7717_), .A2(new_n7736_), .B(\asqrt[32] ), .ZN(new_n7738_));
  OAI21_X1   g07546(.A1(new_n7662_), .A2(new_n7737_), .B(new_n7738_), .ZN(new_n7739_));
  OAI21_X1   g07547(.A1(new_n7739_), .A2(\asqrt[33] ), .B(new_n7659_), .ZN(new_n7740_));
  NAND2_X1   g07548(.A1(new_n7739_), .A2(\asqrt[33] ), .ZN(new_n7741_));
  NAND3_X1   g07549(.A1(new_n7740_), .A2(new_n7741_), .A3(new_n5029_), .ZN(new_n7742_));
  AOI21_X1   g07550(.A1(new_n7740_), .A2(new_n7741_), .B(new_n5029_), .ZN(new_n7743_));
  AOI21_X1   g07551(.A1(new_n7656_), .A2(new_n7742_), .B(new_n7743_), .ZN(new_n7744_));
  AOI21_X1   g07552(.A1(new_n7744_), .A2(new_n4751_), .B(new_n7653_), .ZN(new_n7745_));
  NAND2_X1   g07553(.A1(new_n7742_), .A2(new_n7656_), .ZN(new_n7746_));
  INV_X1     g07554(.I(new_n7659_), .ZN(new_n7747_));
  INV_X1     g07555(.I(new_n7667_), .ZN(new_n7748_));
  NOR3_X1    g07556(.A1(new_n7732_), .A2(\asqrt[30] ), .A3(new_n7734_), .ZN(new_n7749_));
  OAI21_X1   g07557(.A1(new_n7748_), .A2(new_n7749_), .B(new_n7735_), .ZN(new_n7750_));
  OAI21_X1   g07558(.A1(new_n7750_), .A2(\asqrt[31] ), .B(new_n7664_), .ZN(new_n7751_));
  NAND2_X1   g07559(.A1(new_n7750_), .A2(\asqrt[31] ), .ZN(new_n7752_));
  NAND3_X1   g07560(.A1(new_n7751_), .A2(new_n7752_), .A3(new_n5643_), .ZN(new_n7753_));
  AOI21_X1   g07561(.A1(new_n7751_), .A2(new_n7752_), .B(new_n5643_), .ZN(new_n7754_));
  AOI21_X1   g07562(.A1(new_n7661_), .A2(new_n7753_), .B(new_n7754_), .ZN(new_n7755_));
  AOI21_X1   g07563(.A1(new_n7755_), .A2(new_n5336_), .B(new_n7747_), .ZN(new_n7756_));
  NAND2_X1   g07564(.A1(new_n7753_), .A2(new_n7661_), .ZN(new_n7757_));
  AOI21_X1   g07565(.A1(new_n7757_), .A2(new_n7738_), .B(new_n5336_), .ZN(new_n7758_));
  OAI21_X1   g07566(.A1(new_n7756_), .A2(new_n7758_), .B(\asqrt[34] ), .ZN(new_n7759_));
  AOI21_X1   g07567(.A1(new_n7746_), .A2(new_n7759_), .B(new_n4751_), .ZN(new_n7760_));
  NOR3_X1    g07568(.A1(new_n7745_), .A2(\asqrt[36] ), .A3(new_n7760_), .ZN(new_n7761_));
  OAI21_X1   g07569(.A1(new_n7745_), .A2(new_n7760_), .B(\asqrt[36] ), .ZN(new_n7762_));
  OAI21_X1   g07570(.A1(new_n7650_), .A2(new_n7761_), .B(new_n7762_), .ZN(new_n7763_));
  OAI21_X1   g07571(.A1(new_n7763_), .A2(\asqrt[37] ), .B(new_n7647_), .ZN(new_n7764_));
  NAND2_X1   g07572(.A1(new_n7763_), .A2(\asqrt[37] ), .ZN(new_n7765_));
  NAND3_X1   g07573(.A1(new_n7764_), .A2(new_n7765_), .A3(new_n3925_), .ZN(new_n7766_));
  AOI21_X1   g07574(.A1(new_n7764_), .A2(new_n7765_), .B(new_n3925_), .ZN(new_n7767_));
  AOI21_X1   g07575(.A1(new_n7644_), .A2(new_n7766_), .B(new_n7767_), .ZN(new_n7768_));
  NAND2_X1   g07576(.A1(new_n7768_), .A2(new_n3681_), .ZN(new_n7769_));
  INV_X1     g07577(.I(new_n7644_), .ZN(new_n7770_));
  INV_X1     g07578(.I(new_n7647_), .ZN(new_n7771_));
  INV_X1     g07579(.I(new_n7656_), .ZN(new_n7772_));
  NOR3_X1    g07580(.A1(new_n7756_), .A2(\asqrt[34] ), .A3(new_n7758_), .ZN(new_n7773_));
  OAI21_X1   g07581(.A1(new_n7772_), .A2(new_n7773_), .B(new_n7759_), .ZN(new_n7774_));
  OAI21_X1   g07582(.A1(new_n7774_), .A2(\asqrt[35] ), .B(new_n7652_), .ZN(new_n7775_));
  NAND2_X1   g07583(.A1(new_n7774_), .A2(\asqrt[35] ), .ZN(new_n7776_));
  NAND3_X1   g07584(.A1(new_n7775_), .A2(new_n7776_), .A3(new_n4461_), .ZN(new_n7777_));
  AOI21_X1   g07585(.A1(new_n7775_), .A2(new_n7776_), .B(new_n4461_), .ZN(new_n7778_));
  AOI21_X1   g07586(.A1(new_n7649_), .A2(new_n7777_), .B(new_n7778_), .ZN(new_n7779_));
  AOI21_X1   g07587(.A1(new_n7779_), .A2(new_n4196_), .B(new_n7771_), .ZN(new_n7780_));
  NAND2_X1   g07588(.A1(new_n7777_), .A2(new_n7649_), .ZN(new_n7781_));
  AOI21_X1   g07589(.A1(new_n7781_), .A2(new_n7762_), .B(new_n4196_), .ZN(new_n7782_));
  NOR3_X1    g07590(.A1(new_n7780_), .A2(\asqrt[38] ), .A3(new_n7782_), .ZN(new_n7783_));
  OAI21_X1   g07591(.A1(new_n7780_), .A2(new_n7782_), .B(\asqrt[38] ), .ZN(new_n7784_));
  OAI21_X1   g07592(.A1(new_n7770_), .A2(new_n7783_), .B(new_n7784_), .ZN(new_n7785_));
  NAND2_X1   g07593(.A1(new_n7785_), .A2(\asqrt[39] ), .ZN(new_n7786_));
  NOR2_X1    g07594(.A1(new_n7596_), .A2(\asqrt[62] ), .ZN(new_n7787_));
  NOR2_X1    g07595(.A1(new_n7787_), .A2(new_n7681_), .ZN(new_n7788_));
  XOR2_X1    g07596(.A1(new_n7620_), .A2(new_n7259_), .Z(new_n7789_));
  OAI21_X1   g07597(.A1(\asqrt[26] ), .A2(new_n7788_), .B(new_n7789_), .ZN(new_n7790_));
  INV_X1     g07598(.I(new_n7790_), .ZN(new_n7791_));
  AOI21_X1   g07599(.A1(new_n7604_), .A2(new_n7609_), .B(\asqrt[26] ), .ZN(new_n7792_));
  XOR2_X1    g07600(.A1(new_n7792_), .A2(new_n7422_), .Z(new_n7793_));
  INV_X1     g07601(.I(new_n7793_), .ZN(new_n7794_));
  AOI21_X1   g07602(.A1(new_n7584_), .A2(new_n7603_), .B(\asqrt[26] ), .ZN(new_n7795_));
  XOR2_X1    g07603(.A1(new_n7795_), .A2(new_n7426_), .Z(new_n7796_));
  INV_X1     g07604(.I(new_n7796_), .ZN(new_n7797_));
  NOR2_X1    g07605(.A1(new_n7602_), .A2(new_n7598_), .ZN(new_n7798_));
  NOR2_X1    g07606(.A1(\asqrt[26] ), .A2(new_n7798_), .ZN(new_n7799_));
  XOR2_X1    g07607(.A1(new_n7799_), .A2(new_n7428_), .Z(new_n7800_));
  NOR2_X1    g07608(.A1(new_n7573_), .A2(new_n7582_), .ZN(new_n7801_));
  NOR2_X1    g07609(.A1(\asqrt[26] ), .A2(new_n7801_), .ZN(new_n7802_));
  XOR2_X1    g07610(.A1(new_n7802_), .A2(new_n7431_), .Z(new_n7803_));
  AOI21_X1   g07611(.A1(new_n7577_), .A2(new_n7581_), .B(\asqrt[26] ), .ZN(new_n7804_));
  XOR2_X1    g07612(.A1(new_n7804_), .A2(new_n7434_), .Z(new_n7805_));
  INV_X1     g07613(.I(new_n7805_), .ZN(new_n7806_));
  AOI21_X1   g07614(.A1(new_n7563_), .A2(new_n7571_), .B(\asqrt[26] ), .ZN(new_n7807_));
  XOR2_X1    g07615(.A1(new_n7807_), .A2(new_n7438_), .Z(new_n7808_));
  INV_X1     g07616(.I(new_n7808_), .ZN(new_n7809_));
  XOR2_X1    g07617(.A1(new_n7554_), .A2(\asqrt[53] ), .Z(new_n7810_));
  NOR2_X1    g07618(.A1(\asqrt[26] ), .A2(new_n7810_), .ZN(new_n7811_));
  XOR2_X1    g07619(.A1(new_n7811_), .A2(new_n7440_), .Z(new_n7812_));
  NOR2_X1    g07620(.A1(new_n7552_), .A2(new_n7561_), .ZN(new_n7813_));
  NOR2_X1    g07621(.A1(\asqrt[26] ), .A2(new_n7813_), .ZN(new_n7814_));
  XOR2_X1    g07622(.A1(new_n7814_), .A2(new_n7443_), .Z(new_n7815_));
  AOI21_X1   g07623(.A1(new_n7556_), .A2(new_n7560_), .B(\asqrt[26] ), .ZN(new_n7816_));
  XOR2_X1    g07624(.A1(new_n7816_), .A2(new_n7446_), .Z(new_n7817_));
  INV_X1     g07625(.I(new_n7817_), .ZN(new_n7818_));
  AOI21_X1   g07626(.A1(new_n7542_), .A2(new_n7550_), .B(\asqrt[26] ), .ZN(new_n7819_));
  XOR2_X1    g07627(.A1(new_n7819_), .A2(new_n7450_), .Z(new_n7820_));
  INV_X1     g07628(.I(new_n7820_), .ZN(new_n7821_));
  XOR2_X1    g07629(.A1(new_n7533_), .A2(\asqrt[49] ), .Z(new_n7822_));
  NOR2_X1    g07630(.A1(\asqrt[26] ), .A2(new_n7822_), .ZN(new_n7823_));
  XOR2_X1    g07631(.A1(new_n7823_), .A2(new_n7452_), .Z(new_n7824_));
  NOR2_X1    g07632(.A1(new_n7531_), .A2(new_n7540_), .ZN(new_n7825_));
  NOR2_X1    g07633(.A1(\asqrt[26] ), .A2(new_n7825_), .ZN(new_n7826_));
  XOR2_X1    g07634(.A1(new_n7826_), .A2(new_n7455_), .Z(new_n7827_));
  AOI21_X1   g07635(.A1(new_n7535_), .A2(new_n7539_), .B(\asqrt[26] ), .ZN(new_n7828_));
  XOR2_X1    g07636(.A1(new_n7828_), .A2(new_n7458_), .Z(new_n7829_));
  INV_X1     g07637(.I(new_n7829_), .ZN(new_n7830_));
  AOI21_X1   g07638(.A1(new_n7521_), .A2(new_n7529_), .B(\asqrt[26] ), .ZN(new_n7831_));
  XOR2_X1    g07639(.A1(new_n7831_), .A2(new_n7462_), .Z(new_n7832_));
  INV_X1     g07640(.I(new_n7832_), .ZN(new_n7833_));
  XOR2_X1    g07641(.A1(new_n7512_), .A2(\asqrt[45] ), .Z(new_n7834_));
  NOR2_X1    g07642(.A1(\asqrt[26] ), .A2(new_n7834_), .ZN(new_n7835_));
  XOR2_X1    g07643(.A1(new_n7835_), .A2(new_n7464_), .Z(new_n7836_));
  NOR2_X1    g07644(.A1(new_n7510_), .A2(new_n7519_), .ZN(new_n7837_));
  NOR2_X1    g07645(.A1(\asqrt[26] ), .A2(new_n7837_), .ZN(new_n7838_));
  XOR2_X1    g07646(.A1(new_n7838_), .A2(new_n7467_), .Z(new_n7839_));
  AOI21_X1   g07647(.A1(new_n7514_), .A2(new_n7518_), .B(\asqrt[26] ), .ZN(new_n7840_));
  XOR2_X1    g07648(.A1(new_n7840_), .A2(new_n7470_), .Z(new_n7841_));
  INV_X1     g07649(.I(new_n7841_), .ZN(new_n7842_));
  AOI21_X1   g07650(.A1(new_n7500_), .A2(new_n7508_), .B(\asqrt[26] ), .ZN(new_n7843_));
  XOR2_X1    g07651(.A1(new_n7843_), .A2(new_n7474_), .Z(new_n7844_));
  INV_X1     g07652(.I(new_n7844_), .ZN(new_n7845_));
  XOR2_X1    g07653(.A1(new_n7491_), .A2(\asqrt[41] ), .Z(new_n7846_));
  NOR2_X1    g07654(.A1(\asqrt[26] ), .A2(new_n7846_), .ZN(new_n7847_));
  XOR2_X1    g07655(.A1(new_n7847_), .A2(new_n7476_), .Z(new_n7848_));
  NOR2_X1    g07656(.A1(new_n7489_), .A2(new_n7498_), .ZN(new_n7849_));
  NOR2_X1    g07657(.A1(\asqrt[26] ), .A2(new_n7849_), .ZN(new_n7850_));
  XOR2_X1    g07658(.A1(new_n7850_), .A2(new_n7479_), .Z(new_n7851_));
  AOI21_X1   g07659(.A1(new_n7493_), .A2(new_n7497_), .B(\asqrt[26] ), .ZN(new_n7852_));
  XOR2_X1    g07660(.A1(new_n7852_), .A2(new_n7482_), .Z(new_n7853_));
  INV_X1     g07661(.I(new_n7853_), .ZN(new_n7854_));
  INV_X1     g07662(.I(new_n7641_), .ZN(new_n7855_));
  AOI21_X1   g07663(.A1(new_n7768_), .A2(new_n3681_), .B(new_n7855_), .ZN(new_n7856_));
  NAND2_X1   g07664(.A1(new_n7766_), .A2(new_n7644_), .ZN(new_n7857_));
  AOI21_X1   g07665(.A1(new_n7857_), .A2(new_n7784_), .B(new_n3681_), .ZN(new_n7858_));
  NOR3_X1    g07666(.A1(new_n7856_), .A2(\asqrt[40] ), .A3(new_n7858_), .ZN(new_n7859_));
  OAI21_X1   g07667(.A1(new_n7856_), .A2(new_n7858_), .B(\asqrt[40] ), .ZN(new_n7860_));
  OAI21_X1   g07668(.A1(new_n7854_), .A2(new_n7859_), .B(new_n7860_), .ZN(new_n7861_));
  OAI21_X1   g07669(.A1(new_n7861_), .A2(\asqrt[41] ), .B(new_n7851_), .ZN(new_n7862_));
  NAND2_X1   g07670(.A1(new_n7861_), .A2(\asqrt[41] ), .ZN(new_n7863_));
  NAND3_X1   g07671(.A1(new_n7862_), .A2(new_n7863_), .A3(new_n2960_), .ZN(new_n7864_));
  AOI21_X1   g07672(.A1(new_n7862_), .A2(new_n7863_), .B(new_n2960_), .ZN(new_n7865_));
  AOI21_X1   g07673(.A1(new_n7848_), .A2(new_n7864_), .B(new_n7865_), .ZN(new_n7866_));
  AOI21_X1   g07674(.A1(new_n7866_), .A2(new_n2749_), .B(new_n7845_), .ZN(new_n7867_));
  NAND2_X1   g07675(.A1(new_n7864_), .A2(new_n7848_), .ZN(new_n7868_));
  INV_X1     g07676(.I(new_n7851_), .ZN(new_n7869_));
  OAI21_X1   g07677(.A1(new_n7785_), .A2(\asqrt[39] ), .B(new_n7641_), .ZN(new_n7870_));
  NAND3_X1   g07678(.A1(new_n7870_), .A2(new_n7786_), .A3(new_n3427_), .ZN(new_n7871_));
  AOI21_X1   g07679(.A1(new_n7870_), .A2(new_n7786_), .B(new_n3427_), .ZN(new_n7872_));
  AOI21_X1   g07680(.A1(new_n7853_), .A2(new_n7871_), .B(new_n7872_), .ZN(new_n7873_));
  AOI21_X1   g07681(.A1(new_n7873_), .A2(new_n3195_), .B(new_n7869_), .ZN(new_n7874_));
  NAND2_X1   g07682(.A1(new_n7871_), .A2(new_n7853_), .ZN(new_n7875_));
  AOI21_X1   g07683(.A1(new_n7875_), .A2(new_n7860_), .B(new_n3195_), .ZN(new_n7876_));
  OAI21_X1   g07684(.A1(new_n7874_), .A2(new_n7876_), .B(\asqrt[42] ), .ZN(new_n7877_));
  AOI21_X1   g07685(.A1(new_n7868_), .A2(new_n7877_), .B(new_n2749_), .ZN(new_n7878_));
  NOR3_X1    g07686(.A1(new_n7867_), .A2(\asqrt[44] ), .A3(new_n7878_), .ZN(new_n7879_));
  OAI21_X1   g07687(.A1(new_n7867_), .A2(new_n7878_), .B(\asqrt[44] ), .ZN(new_n7880_));
  OAI21_X1   g07688(.A1(new_n7842_), .A2(new_n7879_), .B(new_n7880_), .ZN(new_n7881_));
  OAI21_X1   g07689(.A1(new_n7881_), .A2(\asqrt[45] ), .B(new_n7839_), .ZN(new_n7882_));
  NAND2_X1   g07690(.A1(new_n7881_), .A2(\asqrt[45] ), .ZN(new_n7883_));
  NAND3_X1   g07691(.A1(new_n7882_), .A2(new_n7883_), .A3(new_n2134_), .ZN(new_n7884_));
  AOI21_X1   g07692(.A1(new_n7882_), .A2(new_n7883_), .B(new_n2134_), .ZN(new_n7885_));
  AOI21_X1   g07693(.A1(new_n7836_), .A2(new_n7884_), .B(new_n7885_), .ZN(new_n7886_));
  AOI21_X1   g07694(.A1(new_n7886_), .A2(new_n1953_), .B(new_n7833_), .ZN(new_n7887_));
  NAND2_X1   g07695(.A1(new_n7884_), .A2(new_n7836_), .ZN(new_n7888_));
  INV_X1     g07696(.I(new_n7839_), .ZN(new_n7889_));
  INV_X1     g07697(.I(new_n7848_), .ZN(new_n7890_));
  NOR3_X1    g07698(.A1(new_n7874_), .A2(\asqrt[42] ), .A3(new_n7876_), .ZN(new_n7891_));
  OAI21_X1   g07699(.A1(new_n7890_), .A2(new_n7891_), .B(new_n7877_), .ZN(new_n7892_));
  OAI21_X1   g07700(.A1(new_n7892_), .A2(\asqrt[43] ), .B(new_n7844_), .ZN(new_n7893_));
  NAND2_X1   g07701(.A1(new_n7892_), .A2(\asqrt[43] ), .ZN(new_n7894_));
  NAND3_X1   g07702(.A1(new_n7893_), .A2(new_n7894_), .A3(new_n2531_), .ZN(new_n7895_));
  AOI21_X1   g07703(.A1(new_n7893_), .A2(new_n7894_), .B(new_n2531_), .ZN(new_n7896_));
  AOI21_X1   g07704(.A1(new_n7841_), .A2(new_n7895_), .B(new_n7896_), .ZN(new_n7897_));
  AOI21_X1   g07705(.A1(new_n7897_), .A2(new_n2332_), .B(new_n7889_), .ZN(new_n7898_));
  NAND2_X1   g07706(.A1(new_n7895_), .A2(new_n7841_), .ZN(new_n7899_));
  AOI21_X1   g07707(.A1(new_n7899_), .A2(new_n7880_), .B(new_n2332_), .ZN(new_n7900_));
  OAI21_X1   g07708(.A1(new_n7898_), .A2(new_n7900_), .B(\asqrt[46] ), .ZN(new_n7901_));
  AOI21_X1   g07709(.A1(new_n7888_), .A2(new_n7901_), .B(new_n1953_), .ZN(new_n7902_));
  NOR3_X1    g07710(.A1(new_n7887_), .A2(\asqrt[48] ), .A3(new_n7902_), .ZN(new_n7903_));
  OAI21_X1   g07711(.A1(new_n7887_), .A2(new_n7902_), .B(\asqrt[48] ), .ZN(new_n7904_));
  OAI21_X1   g07712(.A1(new_n7830_), .A2(new_n7903_), .B(new_n7904_), .ZN(new_n7905_));
  OAI21_X1   g07713(.A1(new_n7905_), .A2(\asqrt[49] ), .B(new_n7827_), .ZN(new_n7906_));
  NAND2_X1   g07714(.A1(new_n7905_), .A2(\asqrt[49] ), .ZN(new_n7907_));
  NAND3_X1   g07715(.A1(new_n7906_), .A2(new_n7907_), .A3(new_n1463_), .ZN(new_n7908_));
  AOI21_X1   g07716(.A1(new_n7906_), .A2(new_n7907_), .B(new_n1463_), .ZN(new_n7909_));
  AOI21_X1   g07717(.A1(new_n7824_), .A2(new_n7908_), .B(new_n7909_), .ZN(new_n7910_));
  AOI21_X1   g07718(.A1(new_n7910_), .A2(new_n1305_), .B(new_n7821_), .ZN(new_n7911_));
  NAND2_X1   g07719(.A1(new_n7908_), .A2(new_n7824_), .ZN(new_n7912_));
  INV_X1     g07720(.I(new_n7827_), .ZN(new_n7913_));
  INV_X1     g07721(.I(new_n7836_), .ZN(new_n7914_));
  NOR3_X1    g07722(.A1(new_n7898_), .A2(\asqrt[46] ), .A3(new_n7900_), .ZN(new_n7915_));
  OAI21_X1   g07723(.A1(new_n7914_), .A2(new_n7915_), .B(new_n7901_), .ZN(new_n7916_));
  OAI21_X1   g07724(.A1(new_n7916_), .A2(\asqrt[47] ), .B(new_n7832_), .ZN(new_n7917_));
  NAND2_X1   g07725(.A1(new_n7916_), .A2(\asqrt[47] ), .ZN(new_n7918_));
  NAND3_X1   g07726(.A1(new_n7917_), .A2(new_n7918_), .A3(new_n1778_), .ZN(new_n7919_));
  AOI21_X1   g07727(.A1(new_n7917_), .A2(new_n7918_), .B(new_n1778_), .ZN(new_n7920_));
  AOI21_X1   g07728(.A1(new_n7829_), .A2(new_n7919_), .B(new_n7920_), .ZN(new_n7921_));
  AOI21_X1   g07729(.A1(new_n7921_), .A2(new_n1632_), .B(new_n7913_), .ZN(new_n7922_));
  NAND2_X1   g07730(.A1(new_n7919_), .A2(new_n7829_), .ZN(new_n7923_));
  AOI21_X1   g07731(.A1(new_n7923_), .A2(new_n7904_), .B(new_n1632_), .ZN(new_n7924_));
  OAI21_X1   g07732(.A1(new_n7922_), .A2(new_n7924_), .B(\asqrt[50] ), .ZN(new_n7925_));
  AOI21_X1   g07733(.A1(new_n7912_), .A2(new_n7925_), .B(new_n1305_), .ZN(new_n7926_));
  NOR3_X1    g07734(.A1(new_n7911_), .A2(\asqrt[52] ), .A3(new_n7926_), .ZN(new_n7927_));
  OAI21_X1   g07735(.A1(new_n7911_), .A2(new_n7926_), .B(\asqrt[52] ), .ZN(new_n7928_));
  OAI21_X1   g07736(.A1(new_n7818_), .A2(new_n7927_), .B(new_n7928_), .ZN(new_n7929_));
  OAI21_X1   g07737(.A1(new_n7929_), .A2(\asqrt[53] ), .B(new_n7815_), .ZN(new_n7930_));
  NAND2_X1   g07738(.A1(new_n7929_), .A2(\asqrt[53] ), .ZN(new_n7931_));
  NAND3_X1   g07739(.A1(new_n7930_), .A2(new_n7931_), .A3(new_n860_), .ZN(new_n7932_));
  AOI21_X1   g07740(.A1(new_n7930_), .A2(new_n7931_), .B(new_n860_), .ZN(new_n7933_));
  AOI21_X1   g07741(.A1(new_n7812_), .A2(new_n7932_), .B(new_n7933_), .ZN(new_n7934_));
  AOI21_X1   g07742(.A1(new_n7934_), .A2(new_n744_), .B(new_n7809_), .ZN(new_n7935_));
  NAND2_X1   g07743(.A1(new_n7932_), .A2(new_n7812_), .ZN(new_n7936_));
  INV_X1     g07744(.I(new_n7815_), .ZN(new_n7937_));
  INV_X1     g07745(.I(new_n7824_), .ZN(new_n7938_));
  NOR3_X1    g07746(.A1(new_n7922_), .A2(\asqrt[50] ), .A3(new_n7924_), .ZN(new_n7939_));
  OAI21_X1   g07747(.A1(new_n7938_), .A2(new_n7939_), .B(new_n7925_), .ZN(new_n7940_));
  OAI21_X1   g07748(.A1(new_n7940_), .A2(\asqrt[51] ), .B(new_n7820_), .ZN(new_n7941_));
  NAND2_X1   g07749(.A1(new_n7940_), .A2(\asqrt[51] ), .ZN(new_n7942_));
  NAND3_X1   g07750(.A1(new_n7941_), .A2(new_n7942_), .A3(new_n1150_), .ZN(new_n7943_));
  AOI21_X1   g07751(.A1(new_n7941_), .A2(new_n7942_), .B(new_n1150_), .ZN(new_n7944_));
  AOI21_X1   g07752(.A1(new_n7817_), .A2(new_n7943_), .B(new_n7944_), .ZN(new_n7945_));
  AOI21_X1   g07753(.A1(new_n7945_), .A2(new_n1006_), .B(new_n7937_), .ZN(new_n7946_));
  NAND2_X1   g07754(.A1(new_n7943_), .A2(new_n7817_), .ZN(new_n7947_));
  AOI21_X1   g07755(.A1(new_n7947_), .A2(new_n7928_), .B(new_n1006_), .ZN(new_n7948_));
  OAI21_X1   g07756(.A1(new_n7946_), .A2(new_n7948_), .B(\asqrt[54] ), .ZN(new_n7949_));
  AOI21_X1   g07757(.A1(new_n7936_), .A2(new_n7949_), .B(new_n744_), .ZN(new_n7950_));
  NOR3_X1    g07758(.A1(new_n7935_), .A2(\asqrt[56] ), .A3(new_n7950_), .ZN(new_n7951_));
  OAI21_X1   g07759(.A1(new_n7935_), .A2(new_n7950_), .B(\asqrt[56] ), .ZN(new_n7952_));
  OAI21_X1   g07760(.A1(new_n7806_), .A2(new_n7951_), .B(new_n7952_), .ZN(new_n7953_));
  OAI21_X1   g07761(.A1(new_n7953_), .A2(\asqrt[57] ), .B(new_n7803_), .ZN(new_n7954_));
  NAND2_X1   g07762(.A1(new_n7953_), .A2(\asqrt[57] ), .ZN(new_n7955_));
  NAND3_X1   g07763(.A1(new_n7954_), .A2(new_n7955_), .A3(new_n423_), .ZN(new_n7956_));
  AOI21_X1   g07764(.A1(new_n7954_), .A2(new_n7955_), .B(new_n423_), .ZN(new_n7957_));
  AOI21_X1   g07765(.A1(new_n7800_), .A2(new_n7956_), .B(new_n7957_), .ZN(new_n7958_));
  AOI21_X1   g07766(.A1(new_n7958_), .A2(new_n337_), .B(new_n7797_), .ZN(new_n7959_));
  NAND2_X1   g07767(.A1(new_n7956_), .A2(new_n7800_), .ZN(new_n7960_));
  INV_X1     g07768(.I(new_n7803_), .ZN(new_n7961_));
  INV_X1     g07769(.I(new_n7812_), .ZN(new_n7962_));
  NOR3_X1    g07770(.A1(new_n7946_), .A2(\asqrt[54] ), .A3(new_n7948_), .ZN(new_n7963_));
  OAI21_X1   g07771(.A1(new_n7962_), .A2(new_n7963_), .B(new_n7949_), .ZN(new_n7964_));
  OAI21_X1   g07772(.A1(new_n7964_), .A2(\asqrt[55] ), .B(new_n7808_), .ZN(new_n7965_));
  NAND2_X1   g07773(.A1(new_n7964_), .A2(\asqrt[55] ), .ZN(new_n7966_));
  NAND3_X1   g07774(.A1(new_n7965_), .A2(new_n7966_), .A3(new_n634_), .ZN(new_n7967_));
  AOI21_X1   g07775(.A1(new_n7965_), .A2(new_n7966_), .B(new_n634_), .ZN(new_n7968_));
  AOI21_X1   g07776(.A1(new_n7805_), .A2(new_n7967_), .B(new_n7968_), .ZN(new_n7969_));
  AOI21_X1   g07777(.A1(new_n7969_), .A2(new_n531_), .B(new_n7961_), .ZN(new_n7970_));
  NAND2_X1   g07778(.A1(new_n7967_), .A2(new_n7805_), .ZN(new_n7971_));
  AOI21_X1   g07779(.A1(new_n7971_), .A2(new_n7952_), .B(new_n531_), .ZN(new_n7972_));
  OAI21_X1   g07780(.A1(new_n7970_), .A2(new_n7972_), .B(\asqrt[58] ), .ZN(new_n7973_));
  AOI21_X1   g07781(.A1(new_n7960_), .A2(new_n7973_), .B(new_n337_), .ZN(new_n7974_));
  NOR3_X1    g07782(.A1(new_n7959_), .A2(\asqrt[60] ), .A3(new_n7974_), .ZN(new_n7975_));
  NOR2_X1    g07783(.A1(new_n7975_), .A2(new_n7794_), .ZN(new_n7976_));
  INV_X1     g07784(.I(new_n7800_), .ZN(new_n7977_));
  NOR3_X1    g07785(.A1(new_n7970_), .A2(\asqrt[58] ), .A3(new_n7972_), .ZN(new_n7978_));
  OAI21_X1   g07786(.A1(new_n7977_), .A2(new_n7978_), .B(new_n7973_), .ZN(new_n7979_));
  OAI21_X1   g07787(.A1(new_n7979_), .A2(\asqrt[59] ), .B(new_n7796_), .ZN(new_n7980_));
  NOR2_X1    g07788(.A1(new_n7978_), .A2(new_n7977_), .ZN(new_n7981_));
  OAI21_X1   g07789(.A1(new_n7981_), .A2(new_n7957_), .B(\asqrt[59] ), .ZN(new_n7982_));
  AOI21_X1   g07790(.A1(new_n7980_), .A2(new_n7982_), .B(new_n266_), .ZN(new_n7983_));
  OAI21_X1   g07791(.A1(new_n7976_), .A2(new_n7983_), .B(\asqrt[61] ), .ZN(new_n7984_));
  OAI21_X1   g07792(.A1(new_n7959_), .A2(new_n7974_), .B(\asqrt[60] ), .ZN(new_n7985_));
  OAI21_X1   g07793(.A1(new_n7794_), .A2(new_n7975_), .B(new_n7985_), .ZN(new_n7986_));
  AOI21_X1   g07794(.A1(new_n7610_), .A2(new_n7590_), .B(\asqrt[26] ), .ZN(new_n7987_));
  XOR2_X1    g07795(.A1(new_n7987_), .A2(new_n7419_), .Z(new_n7988_));
  OAI21_X1   g07796(.A1(new_n7986_), .A2(\asqrt[61] ), .B(new_n7988_), .ZN(new_n7989_));
  NAND2_X1   g07797(.A1(new_n7989_), .A2(new_n7984_), .ZN(new_n7990_));
  NAND3_X1   g07798(.A1(new_n7980_), .A2(new_n266_), .A3(new_n7982_), .ZN(new_n7991_));
  NAND2_X1   g07799(.A1(new_n7991_), .A2(new_n7793_), .ZN(new_n7992_));
  AOI21_X1   g07800(.A1(new_n7992_), .A2(new_n7985_), .B(new_n239_), .ZN(new_n7993_));
  AOI21_X1   g07801(.A1(new_n7793_), .A2(new_n7991_), .B(new_n7983_), .ZN(new_n7994_));
  INV_X1     g07802(.I(new_n7988_), .ZN(new_n7995_));
  AOI21_X1   g07803(.A1(new_n7994_), .A2(new_n239_), .B(new_n7995_), .ZN(new_n7996_));
  OAI21_X1   g07804(.A1(new_n7996_), .A2(new_n7993_), .B(new_n201_), .ZN(new_n7997_));
  NAND3_X1   g07805(.A1(new_n7989_), .A2(\asqrt[62] ), .A3(new_n7984_), .ZN(new_n7998_));
  NAND2_X1   g07806(.A1(new_n7614_), .A2(new_n239_), .ZN(new_n7999_));
  AOI21_X1   g07807(.A1(new_n7592_), .A2(new_n7999_), .B(\asqrt[26] ), .ZN(new_n8000_));
  XOR2_X1    g07808(.A1(new_n8000_), .A2(new_n7594_), .Z(new_n8001_));
  INV_X1     g07809(.I(new_n8001_), .ZN(new_n8002_));
  AOI22_X1   g07810(.A1(new_n7997_), .A2(new_n7998_), .B1(new_n7990_), .B2(new_n8002_), .ZN(new_n8003_));
  NOR2_X1    g07811(.A1(new_n7623_), .A2(new_n7417_), .ZN(new_n8004_));
  OAI21_X1   g07812(.A1(\asqrt[26] ), .A2(new_n8004_), .B(new_n7630_), .ZN(new_n8005_));
  INV_X1     g07813(.I(new_n8005_), .ZN(new_n8006_));
  OAI21_X1   g07814(.A1(new_n8003_), .A2(new_n7791_), .B(new_n8006_), .ZN(new_n8007_));
  OAI21_X1   g07815(.A1(new_n7990_), .A2(\asqrt[62] ), .B(new_n8001_), .ZN(new_n8008_));
  NAND2_X1   g07816(.A1(new_n7990_), .A2(\asqrt[62] ), .ZN(new_n8009_));
  NAND3_X1   g07817(.A1(new_n8008_), .A2(new_n8009_), .A3(new_n7791_), .ZN(new_n8010_));
  NAND2_X1   g07818(.A1(new_n7690_), .A2(new_n7416_), .ZN(new_n8011_));
  XOR2_X1    g07819(.A1(new_n7678_), .A2(new_n7416_), .Z(new_n8012_));
  NAND3_X1   g07820(.A1(new_n8011_), .A2(\asqrt[63] ), .A3(new_n8012_), .ZN(new_n8013_));
  INV_X1     g07821(.I(new_n7687_), .ZN(new_n8014_));
  NAND4_X1   g07822(.A1(new_n8014_), .A2(new_n7417_), .A3(new_n7630_), .A4(new_n7638_), .ZN(new_n8015_));
  NAND2_X1   g07823(.A1(new_n8013_), .A2(new_n8015_), .ZN(new_n8016_));
  INV_X1     g07824(.I(new_n8016_), .ZN(new_n8017_));
  NAND4_X1   g07825(.A1(new_n8007_), .A2(new_n193_), .A3(new_n8010_), .A4(new_n8017_), .ZN(\asqrt[25] ));
  AOI21_X1   g07826(.A1(new_n7769_), .A2(new_n7786_), .B(\asqrt[25] ), .ZN(new_n8019_));
  XOR2_X1    g07827(.A1(new_n8019_), .A2(new_n7641_), .Z(new_n8020_));
  AOI21_X1   g07828(.A1(new_n7766_), .A2(new_n7784_), .B(\asqrt[25] ), .ZN(new_n8021_));
  XOR2_X1    g07829(.A1(new_n8021_), .A2(new_n7644_), .Z(new_n8022_));
  NAND2_X1   g07830(.A1(new_n7779_), .A2(new_n4196_), .ZN(new_n8023_));
  AOI21_X1   g07831(.A1(new_n8023_), .A2(new_n7765_), .B(\asqrt[25] ), .ZN(new_n8024_));
  XOR2_X1    g07832(.A1(new_n8024_), .A2(new_n7647_), .Z(new_n8025_));
  INV_X1     g07833(.I(new_n8025_), .ZN(new_n8026_));
  AOI21_X1   g07834(.A1(new_n7777_), .A2(new_n7762_), .B(\asqrt[25] ), .ZN(new_n8027_));
  XOR2_X1    g07835(.A1(new_n8027_), .A2(new_n7649_), .Z(new_n8028_));
  INV_X1     g07836(.I(new_n8028_), .ZN(new_n8029_));
  NAND2_X1   g07837(.A1(new_n7744_), .A2(new_n4751_), .ZN(new_n8030_));
  AOI21_X1   g07838(.A1(new_n8030_), .A2(new_n7776_), .B(\asqrt[25] ), .ZN(new_n8031_));
  XOR2_X1    g07839(.A1(new_n8031_), .A2(new_n7652_), .Z(new_n8032_));
  AOI21_X1   g07840(.A1(new_n7742_), .A2(new_n7759_), .B(\asqrt[25] ), .ZN(new_n8033_));
  XOR2_X1    g07841(.A1(new_n8033_), .A2(new_n7656_), .Z(new_n8034_));
  NAND2_X1   g07842(.A1(new_n7755_), .A2(new_n5336_), .ZN(new_n8035_));
  AOI21_X1   g07843(.A1(new_n8035_), .A2(new_n7741_), .B(\asqrt[25] ), .ZN(new_n8036_));
  XOR2_X1    g07844(.A1(new_n8036_), .A2(new_n7659_), .Z(new_n8037_));
  INV_X1     g07845(.I(new_n8037_), .ZN(new_n8038_));
  AOI21_X1   g07846(.A1(new_n7753_), .A2(new_n7738_), .B(\asqrt[25] ), .ZN(new_n8039_));
  XOR2_X1    g07847(.A1(new_n8039_), .A2(new_n7661_), .Z(new_n8040_));
  INV_X1     g07848(.I(new_n8040_), .ZN(new_n8041_));
  NAND2_X1   g07849(.A1(new_n7716_), .A2(new_n5947_), .ZN(new_n8042_));
  AOI21_X1   g07850(.A1(new_n8042_), .A2(new_n7752_), .B(\asqrt[25] ), .ZN(new_n8043_));
  XOR2_X1    g07851(.A1(new_n8043_), .A2(new_n7664_), .Z(new_n8044_));
  AOI21_X1   g07852(.A1(new_n7714_), .A2(new_n7735_), .B(\asqrt[25] ), .ZN(new_n8045_));
  XOR2_X1    g07853(.A1(new_n8045_), .A2(new_n7667_), .Z(new_n8046_));
  NAND2_X1   g07854(.A1(new_n7731_), .A2(new_n6636_), .ZN(new_n8047_));
  AOI21_X1   g07855(.A1(new_n8047_), .A2(new_n7713_), .B(\asqrt[25] ), .ZN(new_n8048_));
  XOR2_X1    g07856(.A1(new_n8048_), .A2(new_n7674_), .Z(new_n8049_));
  INV_X1     g07857(.I(new_n8049_), .ZN(new_n8050_));
  AOI21_X1   g07858(.A1(new_n7729_), .A2(new_n7710_), .B(\asqrt[25] ), .ZN(new_n8051_));
  XOR2_X1    g07859(.A1(new_n8051_), .A2(new_n7720_), .Z(new_n8052_));
  INV_X1     g07860(.I(new_n8052_), .ZN(new_n8053_));
  NAND2_X1   g07861(.A1(\asqrt[26] ), .A2(new_n7697_), .ZN(new_n8054_));
  NOR2_X1    g07862(.A1(new_n7705_), .A2(\a[52] ), .ZN(new_n8055_));
  AOI22_X1   g07863(.A1(new_n8054_), .A2(new_n7705_), .B1(\asqrt[26] ), .B2(new_n8055_), .ZN(new_n8056_));
  OAI21_X1   g07864(.A1(new_n7690_), .A2(new_n7697_), .B(new_n7724_), .ZN(new_n8057_));
  AOI21_X1   g07865(.A1(new_n7723_), .A2(new_n8057_), .B(\asqrt[25] ), .ZN(new_n8058_));
  XOR2_X1    g07866(.A1(new_n8058_), .A2(new_n8056_), .Z(new_n8059_));
  NAND3_X1   g07867(.A1(new_n7992_), .A2(new_n239_), .A3(new_n7985_), .ZN(new_n8060_));
  AOI21_X1   g07868(.A1(new_n7988_), .A2(new_n8060_), .B(new_n7993_), .ZN(new_n8061_));
  AOI21_X1   g07869(.A1(new_n7989_), .A2(new_n7984_), .B(\asqrt[62] ), .ZN(new_n8062_));
  NOR3_X1    g07870(.A1(new_n7996_), .A2(new_n201_), .A3(new_n7993_), .ZN(new_n8063_));
  OAI22_X1   g07871(.A1(new_n8063_), .A2(new_n8062_), .B1(new_n8061_), .B2(new_n8001_), .ZN(new_n8064_));
  AOI21_X1   g07872(.A1(new_n8064_), .A2(new_n7790_), .B(new_n8005_), .ZN(new_n8065_));
  AOI21_X1   g07873(.A1(new_n8061_), .A2(new_n201_), .B(new_n8002_), .ZN(new_n8066_));
  OAI21_X1   g07874(.A1(new_n8061_), .A2(new_n201_), .B(new_n7791_), .ZN(new_n8067_));
  NOR2_X1    g07875(.A1(new_n8066_), .A2(new_n8067_), .ZN(new_n8068_));
  NOR3_X1    g07876(.A1(new_n8065_), .A2(\asqrt[63] ), .A3(new_n8068_), .ZN(new_n8069_));
  NAND3_X1   g07877(.A1(new_n8013_), .A2(\asqrt[26] ), .A3(new_n8015_), .ZN(new_n8070_));
  INV_X1     g07878(.I(new_n8070_), .ZN(new_n8071_));
  NAND2_X1   g07879(.A1(new_n8069_), .A2(new_n8071_), .ZN(new_n8072_));
  NAND2_X1   g07880(.A1(\asqrt[25] ), .A2(new_n7694_), .ZN(new_n8073_));
  AOI21_X1   g07881(.A1(new_n8073_), .A2(new_n8072_), .B(\a[52] ), .ZN(new_n8074_));
  NAND2_X1   g07882(.A1(new_n8007_), .A2(new_n193_), .ZN(new_n8075_));
  NOR3_X1    g07883(.A1(new_n8075_), .A2(new_n8068_), .A3(new_n8070_), .ZN(new_n8076_));
  NOR4_X1    g07884(.A1(new_n8065_), .A2(\asqrt[63] ), .A3(new_n8068_), .A4(new_n8016_), .ZN(new_n8077_));
  NOR2_X1    g07885(.A1(new_n8077_), .A2(new_n7695_), .ZN(new_n8078_));
  NOR3_X1    g07886(.A1(new_n8078_), .A2(new_n8076_), .A3(new_n7697_), .ZN(new_n8079_));
  NOR2_X1    g07887(.A1(new_n8079_), .A2(new_n8074_), .ZN(new_n8080_));
  INV_X1     g07888(.I(\a[50] ), .ZN(new_n8081_));
  NOR2_X1    g07889(.A1(\a[48] ), .A2(\a[49] ), .ZN(new_n8082_));
  NOR3_X1    g07890(.A1(new_n8077_), .A2(new_n8081_), .A3(new_n8082_), .ZN(new_n8083_));
  INV_X1     g07891(.I(new_n8082_), .ZN(new_n8084_));
  AOI21_X1   g07892(.A1(new_n8077_), .A2(\a[50] ), .B(new_n8084_), .ZN(new_n8085_));
  OAI21_X1   g07893(.A1(new_n8083_), .A2(new_n8085_), .B(\asqrt[26] ), .ZN(new_n8086_));
  NAND2_X1   g07894(.A1(new_n8082_), .A2(new_n8081_), .ZN(new_n8087_));
  NAND3_X1   g07895(.A1(new_n7634_), .A2(new_n7636_), .A3(new_n8087_), .ZN(new_n8088_));
  NAND2_X1   g07896(.A1(new_n7683_), .A2(new_n8088_), .ZN(new_n8089_));
  INV_X1     g07897(.I(new_n8089_), .ZN(new_n8090_));
  NOR3_X1    g07898(.A1(new_n8077_), .A2(new_n8081_), .A3(new_n8090_), .ZN(new_n8091_));
  NOR3_X1    g07899(.A1(new_n8077_), .A2(\a[50] ), .A3(\a[51] ), .ZN(new_n8092_));
  INV_X1     g07900(.I(\a[51] ), .ZN(new_n8093_));
  AOI21_X1   g07901(.A1(\asqrt[25] ), .A2(new_n8081_), .B(new_n8093_), .ZN(new_n8094_));
  NOR3_X1    g07902(.A1(new_n8091_), .A2(new_n8092_), .A3(new_n8094_), .ZN(new_n8095_));
  NAND3_X1   g07903(.A1(new_n8095_), .A2(new_n8086_), .A3(new_n7331_), .ZN(new_n8096_));
  NAND2_X1   g07904(.A1(new_n8096_), .A2(new_n8080_), .ZN(new_n8097_));
  NAND3_X1   g07905(.A1(\asqrt[25] ), .A2(\a[50] ), .A3(new_n8084_), .ZN(new_n8098_));
  OAI21_X1   g07906(.A1(\asqrt[25] ), .A2(new_n8081_), .B(new_n8082_), .ZN(new_n8099_));
  AOI21_X1   g07907(.A1(new_n8099_), .A2(new_n8098_), .B(new_n7690_), .ZN(new_n8100_));
  NAND3_X1   g07908(.A1(\asqrt[25] ), .A2(\a[50] ), .A3(new_n8089_), .ZN(new_n8101_));
  NAND3_X1   g07909(.A1(\asqrt[25] ), .A2(new_n8081_), .A3(new_n8093_), .ZN(new_n8102_));
  OAI21_X1   g07910(.A1(new_n8077_), .A2(\a[50] ), .B(\a[51] ), .ZN(new_n8103_));
  NAND3_X1   g07911(.A1(new_n8101_), .A2(new_n8103_), .A3(new_n8102_), .ZN(new_n8104_));
  OAI21_X1   g07912(.A1(new_n8104_), .A2(new_n8100_), .B(\asqrt[27] ), .ZN(new_n8105_));
  NAND3_X1   g07913(.A1(new_n8097_), .A2(new_n6966_), .A3(new_n8105_), .ZN(new_n8106_));
  AOI21_X1   g07914(.A1(new_n8097_), .A2(new_n8105_), .B(new_n6966_), .ZN(new_n8107_));
  AOI21_X1   g07915(.A1(new_n8059_), .A2(new_n8106_), .B(new_n8107_), .ZN(new_n8108_));
  AOI21_X1   g07916(.A1(new_n8108_), .A2(new_n6636_), .B(new_n8053_), .ZN(new_n8109_));
  OR2_X2     g07917(.A1(new_n8079_), .A2(new_n8074_), .Z(new_n8110_));
  NOR3_X1    g07918(.A1(new_n8104_), .A2(new_n8100_), .A3(\asqrt[27] ), .ZN(new_n8111_));
  OAI21_X1   g07919(.A1(new_n8110_), .A2(new_n8111_), .B(new_n8105_), .ZN(new_n8112_));
  OAI21_X1   g07920(.A1(new_n8112_), .A2(\asqrt[28] ), .B(new_n8059_), .ZN(new_n8113_));
  NAND2_X1   g07921(.A1(new_n8112_), .A2(\asqrt[28] ), .ZN(new_n8114_));
  AOI21_X1   g07922(.A1(new_n8113_), .A2(new_n8114_), .B(new_n6636_), .ZN(new_n8115_));
  NOR3_X1    g07923(.A1(new_n8109_), .A2(\asqrt[30] ), .A3(new_n8115_), .ZN(new_n8116_));
  OAI21_X1   g07924(.A1(new_n8109_), .A2(new_n8115_), .B(\asqrt[30] ), .ZN(new_n8117_));
  OAI21_X1   g07925(.A1(new_n8050_), .A2(new_n8116_), .B(new_n8117_), .ZN(new_n8118_));
  OAI21_X1   g07926(.A1(new_n8118_), .A2(\asqrt[31] ), .B(new_n8046_), .ZN(new_n8119_));
  NAND3_X1   g07927(.A1(new_n8113_), .A2(new_n8114_), .A3(new_n6636_), .ZN(new_n8120_));
  AOI21_X1   g07928(.A1(new_n8052_), .A2(new_n8120_), .B(new_n8115_), .ZN(new_n8121_));
  AOI21_X1   g07929(.A1(new_n8121_), .A2(new_n6275_), .B(new_n8050_), .ZN(new_n8122_));
  NAND2_X1   g07930(.A1(new_n8120_), .A2(new_n8052_), .ZN(new_n8123_));
  INV_X1     g07931(.I(new_n8115_), .ZN(new_n8124_));
  AOI21_X1   g07932(.A1(new_n8123_), .A2(new_n8124_), .B(new_n6275_), .ZN(new_n8125_));
  OAI21_X1   g07933(.A1(new_n8122_), .A2(new_n8125_), .B(\asqrt[31] ), .ZN(new_n8126_));
  NAND3_X1   g07934(.A1(new_n8119_), .A2(new_n5643_), .A3(new_n8126_), .ZN(new_n8127_));
  AOI21_X1   g07935(.A1(new_n8119_), .A2(new_n8126_), .B(new_n5643_), .ZN(new_n8128_));
  AOI21_X1   g07936(.A1(new_n8044_), .A2(new_n8127_), .B(new_n8128_), .ZN(new_n8129_));
  AOI21_X1   g07937(.A1(new_n8129_), .A2(new_n5336_), .B(new_n8041_), .ZN(new_n8130_));
  INV_X1     g07938(.I(new_n8046_), .ZN(new_n8131_));
  NOR3_X1    g07939(.A1(new_n8122_), .A2(\asqrt[31] ), .A3(new_n8125_), .ZN(new_n8132_));
  OAI21_X1   g07940(.A1(new_n8131_), .A2(new_n8132_), .B(new_n8126_), .ZN(new_n8133_));
  OAI21_X1   g07941(.A1(new_n8133_), .A2(\asqrt[32] ), .B(new_n8044_), .ZN(new_n8134_));
  NAND2_X1   g07942(.A1(new_n8133_), .A2(\asqrt[32] ), .ZN(new_n8135_));
  AOI21_X1   g07943(.A1(new_n8134_), .A2(new_n8135_), .B(new_n5336_), .ZN(new_n8136_));
  NOR3_X1    g07944(.A1(new_n8130_), .A2(\asqrt[34] ), .A3(new_n8136_), .ZN(new_n8137_));
  OAI21_X1   g07945(.A1(new_n8130_), .A2(new_n8136_), .B(\asqrt[34] ), .ZN(new_n8138_));
  OAI21_X1   g07946(.A1(new_n8038_), .A2(new_n8137_), .B(new_n8138_), .ZN(new_n8139_));
  OAI21_X1   g07947(.A1(new_n8139_), .A2(\asqrt[35] ), .B(new_n8034_), .ZN(new_n8140_));
  NAND3_X1   g07948(.A1(new_n8134_), .A2(new_n8135_), .A3(new_n5336_), .ZN(new_n8141_));
  AOI21_X1   g07949(.A1(new_n8040_), .A2(new_n8141_), .B(new_n8136_), .ZN(new_n8142_));
  AOI21_X1   g07950(.A1(new_n8142_), .A2(new_n5029_), .B(new_n8038_), .ZN(new_n8143_));
  NAND2_X1   g07951(.A1(new_n8141_), .A2(new_n8040_), .ZN(new_n8144_));
  INV_X1     g07952(.I(new_n8136_), .ZN(new_n8145_));
  AOI21_X1   g07953(.A1(new_n8144_), .A2(new_n8145_), .B(new_n5029_), .ZN(new_n8146_));
  OAI21_X1   g07954(.A1(new_n8143_), .A2(new_n8146_), .B(\asqrt[35] ), .ZN(new_n8147_));
  NAND3_X1   g07955(.A1(new_n8140_), .A2(new_n4461_), .A3(new_n8147_), .ZN(new_n8148_));
  AOI21_X1   g07956(.A1(new_n8140_), .A2(new_n8147_), .B(new_n4461_), .ZN(new_n8149_));
  AOI21_X1   g07957(.A1(new_n8032_), .A2(new_n8148_), .B(new_n8149_), .ZN(new_n8150_));
  AOI21_X1   g07958(.A1(new_n8150_), .A2(new_n4196_), .B(new_n8029_), .ZN(new_n8151_));
  INV_X1     g07959(.I(new_n8034_), .ZN(new_n8152_));
  NOR3_X1    g07960(.A1(new_n8143_), .A2(\asqrt[35] ), .A3(new_n8146_), .ZN(new_n8153_));
  OAI21_X1   g07961(.A1(new_n8152_), .A2(new_n8153_), .B(new_n8147_), .ZN(new_n8154_));
  OAI21_X1   g07962(.A1(new_n8154_), .A2(\asqrt[36] ), .B(new_n8032_), .ZN(new_n8155_));
  NAND2_X1   g07963(.A1(new_n8154_), .A2(\asqrt[36] ), .ZN(new_n8156_));
  AOI21_X1   g07964(.A1(new_n8155_), .A2(new_n8156_), .B(new_n4196_), .ZN(new_n8157_));
  NOR3_X1    g07965(.A1(new_n8151_), .A2(\asqrt[38] ), .A3(new_n8157_), .ZN(new_n8158_));
  OAI21_X1   g07966(.A1(new_n8151_), .A2(new_n8157_), .B(\asqrt[38] ), .ZN(new_n8159_));
  OAI21_X1   g07967(.A1(new_n8026_), .A2(new_n8158_), .B(new_n8159_), .ZN(new_n8160_));
  OAI21_X1   g07968(.A1(new_n8160_), .A2(\asqrt[39] ), .B(new_n8022_), .ZN(new_n8161_));
  NAND3_X1   g07969(.A1(new_n8155_), .A2(new_n8156_), .A3(new_n4196_), .ZN(new_n8162_));
  AOI21_X1   g07970(.A1(new_n8028_), .A2(new_n8162_), .B(new_n8157_), .ZN(new_n8163_));
  AOI21_X1   g07971(.A1(new_n8163_), .A2(new_n3925_), .B(new_n8026_), .ZN(new_n8164_));
  NAND2_X1   g07972(.A1(new_n8162_), .A2(new_n8028_), .ZN(new_n8165_));
  INV_X1     g07973(.I(new_n8157_), .ZN(new_n8166_));
  AOI21_X1   g07974(.A1(new_n8165_), .A2(new_n8166_), .B(new_n3925_), .ZN(new_n8167_));
  OAI21_X1   g07975(.A1(new_n8164_), .A2(new_n8167_), .B(\asqrt[39] ), .ZN(new_n8168_));
  NAND3_X1   g07976(.A1(new_n8161_), .A2(new_n3427_), .A3(new_n8168_), .ZN(new_n8169_));
  INV_X1     g07977(.I(new_n8022_), .ZN(new_n8170_));
  NOR3_X1    g07978(.A1(new_n8164_), .A2(\asqrt[39] ), .A3(new_n8167_), .ZN(new_n8171_));
  OAI21_X1   g07979(.A1(new_n8170_), .A2(new_n8171_), .B(new_n8168_), .ZN(new_n8172_));
  NAND2_X1   g07980(.A1(new_n8172_), .A2(\asqrt[40] ), .ZN(new_n8173_));
  NOR2_X1    g07981(.A1(new_n7990_), .A2(\asqrt[62] ), .ZN(new_n8174_));
  INV_X1     g07982(.I(new_n8009_), .ZN(new_n8175_));
  NOR2_X1    g07983(.A1(new_n8175_), .A2(new_n8174_), .ZN(new_n8176_));
  XOR2_X1    g07984(.A1(new_n8000_), .A2(new_n7594_), .Z(new_n8177_));
  OAI21_X1   g07985(.A1(\asqrt[25] ), .A2(new_n8176_), .B(new_n8177_), .ZN(new_n8178_));
  INV_X1     g07986(.I(new_n8178_), .ZN(new_n8179_));
  NAND2_X1   g07987(.A1(new_n7958_), .A2(new_n337_), .ZN(new_n8180_));
  AOI21_X1   g07988(.A1(new_n8180_), .A2(new_n7982_), .B(\asqrt[25] ), .ZN(new_n8181_));
  XOR2_X1    g07989(.A1(new_n8181_), .A2(new_n7796_), .Z(new_n8182_));
  INV_X1     g07990(.I(new_n8182_), .ZN(new_n8183_));
  AOI21_X1   g07991(.A1(new_n7956_), .A2(new_n7973_), .B(\asqrt[25] ), .ZN(new_n8184_));
  XOR2_X1    g07992(.A1(new_n8184_), .A2(new_n7800_), .Z(new_n8185_));
  INV_X1     g07993(.I(new_n8185_), .ZN(new_n8186_));
  NAND2_X1   g07994(.A1(new_n7969_), .A2(new_n531_), .ZN(new_n8187_));
  AOI21_X1   g07995(.A1(new_n8187_), .A2(new_n7955_), .B(\asqrt[25] ), .ZN(new_n8188_));
  XOR2_X1    g07996(.A1(new_n8188_), .A2(new_n7803_), .Z(new_n8189_));
  INV_X1     g07997(.I(new_n8189_), .ZN(new_n8190_));
  AOI21_X1   g07998(.A1(new_n7967_), .A2(new_n7952_), .B(\asqrt[25] ), .ZN(new_n8191_));
  XOR2_X1    g07999(.A1(new_n8191_), .A2(new_n7805_), .Z(new_n8192_));
  NAND2_X1   g08000(.A1(new_n7934_), .A2(new_n744_), .ZN(new_n8193_));
  AOI21_X1   g08001(.A1(new_n8193_), .A2(new_n7966_), .B(\asqrt[25] ), .ZN(new_n8194_));
  XOR2_X1    g08002(.A1(new_n8194_), .A2(new_n7808_), .Z(new_n8195_));
  AOI21_X1   g08003(.A1(new_n7932_), .A2(new_n7949_), .B(\asqrt[25] ), .ZN(new_n8196_));
  XOR2_X1    g08004(.A1(new_n8196_), .A2(new_n7812_), .Z(new_n8197_));
  INV_X1     g08005(.I(new_n8197_), .ZN(new_n8198_));
  NAND2_X1   g08006(.A1(new_n7945_), .A2(new_n1006_), .ZN(new_n8199_));
  AOI21_X1   g08007(.A1(new_n8199_), .A2(new_n7931_), .B(\asqrt[25] ), .ZN(new_n8200_));
  XOR2_X1    g08008(.A1(new_n8200_), .A2(new_n7815_), .Z(new_n8201_));
  INV_X1     g08009(.I(new_n8201_), .ZN(new_n8202_));
  AOI21_X1   g08010(.A1(new_n7943_), .A2(new_n7928_), .B(\asqrt[25] ), .ZN(new_n8203_));
  XOR2_X1    g08011(.A1(new_n8203_), .A2(new_n7817_), .Z(new_n8204_));
  NAND2_X1   g08012(.A1(new_n7910_), .A2(new_n1305_), .ZN(new_n8205_));
  AOI21_X1   g08013(.A1(new_n8205_), .A2(new_n7942_), .B(\asqrt[25] ), .ZN(new_n8206_));
  XOR2_X1    g08014(.A1(new_n8206_), .A2(new_n7820_), .Z(new_n8207_));
  AOI21_X1   g08015(.A1(new_n7908_), .A2(new_n7925_), .B(\asqrt[25] ), .ZN(new_n8208_));
  XOR2_X1    g08016(.A1(new_n8208_), .A2(new_n7824_), .Z(new_n8209_));
  INV_X1     g08017(.I(new_n8209_), .ZN(new_n8210_));
  NAND2_X1   g08018(.A1(new_n7921_), .A2(new_n1632_), .ZN(new_n8211_));
  AOI21_X1   g08019(.A1(new_n8211_), .A2(new_n7907_), .B(\asqrt[25] ), .ZN(new_n8212_));
  XOR2_X1    g08020(.A1(new_n8212_), .A2(new_n7827_), .Z(new_n8213_));
  INV_X1     g08021(.I(new_n8213_), .ZN(new_n8214_));
  AOI21_X1   g08022(.A1(new_n7919_), .A2(new_n7904_), .B(\asqrt[25] ), .ZN(new_n8215_));
  XOR2_X1    g08023(.A1(new_n8215_), .A2(new_n7829_), .Z(new_n8216_));
  NAND2_X1   g08024(.A1(new_n7886_), .A2(new_n1953_), .ZN(new_n8217_));
  AOI21_X1   g08025(.A1(new_n8217_), .A2(new_n7918_), .B(\asqrt[25] ), .ZN(new_n8218_));
  XOR2_X1    g08026(.A1(new_n8218_), .A2(new_n7832_), .Z(new_n8219_));
  AOI21_X1   g08027(.A1(new_n7884_), .A2(new_n7901_), .B(\asqrt[25] ), .ZN(new_n8220_));
  XOR2_X1    g08028(.A1(new_n8220_), .A2(new_n7836_), .Z(new_n8221_));
  INV_X1     g08029(.I(new_n8221_), .ZN(new_n8222_));
  NAND2_X1   g08030(.A1(new_n7897_), .A2(new_n2332_), .ZN(new_n8223_));
  AOI21_X1   g08031(.A1(new_n8223_), .A2(new_n7883_), .B(\asqrt[25] ), .ZN(new_n8224_));
  XOR2_X1    g08032(.A1(new_n8224_), .A2(new_n7839_), .Z(new_n8225_));
  INV_X1     g08033(.I(new_n8225_), .ZN(new_n8226_));
  AOI21_X1   g08034(.A1(new_n7895_), .A2(new_n7880_), .B(\asqrt[25] ), .ZN(new_n8227_));
  XOR2_X1    g08035(.A1(new_n8227_), .A2(new_n7841_), .Z(new_n8228_));
  NAND2_X1   g08036(.A1(new_n7866_), .A2(new_n2749_), .ZN(new_n8229_));
  AOI21_X1   g08037(.A1(new_n8229_), .A2(new_n7894_), .B(\asqrt[25] ), .ZN(new_n8230_));
  XOR2_X1    g08038(.A1(new_n8230_), .A2(new_n7844_), .Z(new_n8231_));
  AOI21_X1   g08039(.A1(new_n7864_), .A2(new_n7877_), .B(\asqrt[25] ), .ZN(new_n8232_));
  XOR2_X1    g08040(.A1(new_n8232_), .A2(new_n7848_), .Z(new_n8233_));
  INV_X1     g08041(.I(new_n8233_), .ZN(new_n8234_));
  NAND2_X1   g08042(.A1(new_n7873_), .A2(new_n3195_), .ZN(new_n8235_));
  AOI21_X1   g08043(.A1(new_n8235_), .A2(new_n7863_), .B(\asqrt[25] ), .ZN(new_n8236_));
  XOR2_X1    g08044(.A1(new_n8236_), .A2(new_n7851_), .Z(new_n8237_));
  INV_X1     g08045(.I(new_n8237_), .ZN(new_n8238_));
  AOI21_X1   g08046(.A1(new_n7871_), .A2(new_n7860_), .B(\asqrt[25] ), .ZN(new_n8239_));
  XOR2_X1    g08047(.A1(new_n8239_), .A2(new_n7853_), .Z(new_n8240_));
  OAI21_X1   g08048(.A1(new_n8172_), .A2(\asqrt[40] ), .B(new_n8020_), .ZN(new_n8241_));
  NAND3_X1   g08049(.A1(new_n8241_), .A2(new_n8173_), .A3(new_n3195_), .ZN(new_n8242_));
  AOI21_X1   g08050(.A1(new_n8241_), .A2(new_n8173_), .B(new_n3195_), .ZN(new_n8243_));
  AOI21_X1   g08051(.A1(new_n8240_), .A2(new_n8242_), .B(new_n8243_), .ZN(new_n8244_));
  AOI21_X1   g08052(.A1(new_n8244_), .A2(new_n2960_), .B(new_n8238_), .ZN(new_n8245_));
  NAND2_X1   g08053(.A1(new_n8242_), .A2(new_n8240_), .ZN(new_n8246_));
  INV_X1     g08054(.I(new_n8243_), .ZN(new_n8247_));
  AOI21_X1   g08055(.A1(new_n8246_), .A2(new_n8247_), .B(new_n2960_), .ZN(new_n8248_));
  NOR3_X1    g08056(.A1(new_n8245_), .A2(\asqrt[43] ), .A3(new_n8248_), .ZN(new_n8249_));
  OAI21_X1   g08057(.A1(new_n8245_), .A2(new_n8248_), .B(\asqrt[43] ), .ZN(new_n8250_));
  OAI21_X1   g08058(.A1(new_n8234_), .A2(new_n8249_), .B(new_n8250_), .ZN(new_n8251_));
  OAI21_X1   g08059(.A1(new_n8251_), .A2(\asqrt[44] ), .B(new_n8231_), .ZN(new_n8252_));
  NAND2_X1   g08060(.A1(new_n8251_), .A2(\asqrt[44] ), .ZN(new_n8253_));
  NAND3_X1   g08061(.A1(new_n8252_), .A2(new_n8253_), .A3(new_n2332_), .ZN(new_n8254_));
  AOI21_X1   g08062(.A1(new_n8252_), .A2(new_n8253_), .B(new_n2332_), .ZN(new_n8255_));
  AOI21_X1   g08063(.A1(new_n8228_), .A2(new_n8254_), .B(new_n8255_), .ZN(new_n8256_));
  AOI21_X1   g08064(.A1(new_n8256_), .A2(new_n2134_), .B(new_n8226_), .ZN(new_n8257_));
  NAND2_X1   g08065(.A1(new_n8254_), .A2(new_n8228_), .ZN(new_n8258_));
  INV_X1     g08066(.I(new_n8255_), .ZN(new_n8259_));
  AOI21_X1   g08067(.A1(new_n8258_), .A2(new_n8259_), .B(new_n2134_), .ZN(new_n8260_));
  NOR3_X1    g08068(.A1(new_n8257_), .A2(\asqrt[47] ), .A3(new_n8260_), .ZN(new_n8261_));
  OAI21_X1   g08069(.A1(new_n8257_), .A2(new_n8260_), .B(\asqrt[47] ), .ZN(new_n8262_));
  OAI21_X1   g08070(.A1(new_n8222_), .A2(new_n8261_), .B(new_n8262_), .ZN(new_n8263_));
  OAI21_X1   g08071(.A1(new_n8263_), .A2(\asqrt[48] ), .B(new_n8219_), .ZN(new_n8264_));
  NAND2_X1   g08072(.A1(new_n8263_), .A2(\asqrt[48] ), .ZN(new_n8265_));
  NAND3_X1   g08073(.A1(new_n8264_), .A2(new_n8265_), .A3(new_n1632_), .ZN(new_n8266_));
  AOI21_X1   g08074(.A1(new_n8264_), .A2(new_n8265_), .B(new_n1632_), .ZN(new_n8267_));
  AOI21_X1   g08075(.A1(new_n8216_), .A2(new_n8266_), .B(new_n8267_), .ZN(new_n8268_));
  AOI21_X1   g08076(.A1(new_n8268_), .A2(new_n1463_), .B(new_n8214_), .ZN(new_n8269_));
  NAND2_X1   g08077(.A1(new_n8266_), .A2(new_n8216_), .ZN(new_n8270_));
  INV_X1     g08078(.I(new_n8267_), .ZN(new_n8271_));
  AOI21_X1   g08079(.A1(new_n8270_), .A2(new_n8271_), .B(new_n1463_), .ZN(new_n8272_));
  NOR3_X1    g08080(.A1(new_n8269_), .A2(\asqrt[51] ), .A3(new_n8272_), .ZN(new_n8273_));
  OAI21_X1   g08081(.A1(new_n8269_), .A2(new_n8272_), .B(\asqrt[51] ), .ZN(new_n8274_));
  OAI21_X1   g08082(.A1(new_n8210_), .A2(new_n8273_), .B(new_n8274_), .ZN(new_n8275_));
  OAI21_X1   g08083(.A1(new_n8275_), .A2(\asqrt[52] ), .B(new_n8207_), .ZN(new_n8276_));
  NAND2_X1   g08084(.A1(new_n8275_), .A2(\asqrt[52] ), .ZN(new_n8277_));
  NAND3_X1   g08085(.A1(new_n8276_), .A2(new_n8277_), .A3(new_n1006_), .ZN(new_n8278_));
  AOI21_X1   g08086(.A1(new_n8276_), .A2(new_n8277_), .B(new_n1006_), .ZN(new_n8279_));
  AOI21_X1   g08087(.A1(new_n8204_), .A2(new_n8278_), .B(new_n8279_), .ZN(new_n8280_));
  AOI21_X1   g08088(.A1(new_n8280_), .A2(new_n860_), .B(new_n8202_), .ZN(new_n8281_));
  NAND2_X1   g08089(.A1(new_n8278_), .A2(new_n8204_), .ZN(new_n8282_));
  INV_X1     g08090(.I(new_n8279_), .ZN(new_n8283_));
  AOI21_X1   g08091(.A1(new_n8282_), .A2(new_n8283_), .B(new_n860_), .ZN(new_n8284_));
  NOR3_X1    g08092(.A1(new_n8281_), .A2(\asqrt[55] ), .A3(new_n8284_), .ZN(new_n8285_));
  OAI21_X1   g08093(.A1(new_n8281_), .A2(new_n8284_), .B(\asqrt[55] ), .ZN(new_n8286_));
  OAI21_X1   g08094(.A1(new_n8198_), .A2(new_n8285_), .B(new_n8286_), .ZN(new_n8287_));
  OAI21_X1   g08095(.A1(new_n8287_), .A2(\asqrt[56] ), .B(new_n8195_), .ZN(new_n8288_));
  NAND2_X1   g08096(.A1(new_n8287_), .A2(\asqrt[56] ), .ZN(new_n8289_));
  NAND3_X1   g08097(.A1(new_n8288_), .A2(new_n8289_), .A3(new_n531_), .ZN(new_n8290_));
  AOI21_X1   g08098(.A1(new_n8288_), .A2(new_n8289_), .B(new_n531_), .ZN(new_n8291_));
  AOI21_X1   g08099(.A1(new_n8192_), .A2(new_n8290_), .B(new_n8291_), .ZN(new_n8292_));
  AOI21_X1   g08100(.A1(new_n8292_), .A2(new_n423_), .B(new_n8190_), .ZN(new_n8293_));
  NAND2_X1   g08101(.A1(new_n8290_), .A2(new_n8192_), .ZN(new_n8294_));
  INV_X1     g08102(.I(new_n8291_), .ZN(new_n8295_));
  AOI21_X1   g08103(.A1(new_n8294_), .A2(new_n8295_), .B(new_n423_), .ZN(new_n8296_));
  NOR3_X1    g08104(.A1(new_n8293_), .A2(\asqrt[59] ), .A3(new_n8296_), .ZN(new_n8297_));
  NOR2_X1    g08105(.A1(new_n8297_), .A2(new_n8186_), .ZN(new_n8298_));
  OAI21_X1   g08106(.A1(new_n8293_), .A2(new_n8296_), .B(\asqrt[59] ), .ZN(new_n8299_));
  INV_X1     g08107(.I(new_n8299_), .ZN(new_n8300_));
  NOR2_X1    g08108(.A1(new_n8298_), .A2(new_n8300_), .ZN(new_n8301_));
  AOI21_X1   g08109(.A1(new_n8301_), .A2(new_n266_), .B(new_n8183_), .ZN(new_n8302_));
  INV_X1     g08110(.I(new_n8192_), .ZN(new_n8303_));
  INV_X1     g08111(.I(new_n8204_), .ZN(new_n8304_));
  INV_X1     g08112(.I(new_n8216_), .ZN(new_n8305_));
  INV_X1     g08113(.I(new_n8228_), .ZN(new_n8306_));
  INV_X1     g08114(.I(new_n8240_), .ZN(new_n8307_));
  AOI21_X1   g08115(.A1(new_n8161_), .A2(new_n8168_), .B(new_n3427_), .ZN(new_n8308_));
  AOI21_X1   g08116(.A1(new_n8020_), .A2(new_n8169_), .B(new_n8308_), .ZN(new_n8309_));
  AOI21_X1   g08117(.A1(new_n8309_), .A2(new_n3195_), .B(new_n8307_), .ZN(new_n8310_));
  NOR3_X1    g08118(.A1(new_n8310_), .A2(\asqrt[42] ), .A3(new_n8243_), .ZN(new_n8311_));
  OAI21_X1   g08119(.A1(new_n8310_), .A2(new_n8243_), .B(\asqrt[42] ), .ZN(new_n8312_));
  OAI21_X1   g08120(.A1(new_n8238_), .A2(new_n8311_), .B(new_n8312_), .ZN(new_n8313_));
  OAI21_X1   g08121(.A1(new_n8313_), .A2(\asqrt[43] ), .B(new_n8233_), .ZN(new_n8314_));
  NAND3_X1   g08122(.A1(new_n8314_), .A2(new_n2531_), .A3(new_n8250_), .ZN(new_n8315_));
  AOI21_X1   g08123(.A1(new_n8314_), .A2(new_n8250_), .B(new_n2531_), .ZN(new_n8316_));
  AOI21_X1   g08124(.A1(new_n8231_), .A2(new_n8315_), .B(new_n8316_), .ZN(new_n8317_));
  AOI21_X1   g08125(.A1(new_n8317_), .A2(new_n2332_), .B(new_n8306_), .ZN(new_n8318_));
  NOR3_X1    g08126(.A1(new_n8318_), .A2(\asqrt[46] ), .A3(new_n8255_), .ZN(new_n8319_));
  OAI21_X1   g08127(.A1(new_n8318_), .A2(new_n8255_), .B(\asqrt[46] ), .ZN(new_n8320_));
  OAI21_X1   g08128(.A1(new_n8226_), .A2(new_n8319_), .B(new_n8320_), .ZN(new_n8321_));
  OAI21_X1   g08129(.A1(new_n8321_), .A2(\asqrt[47] ), .B(new_n8221_), .ZN(new_n8322_));
  NAND3_X1   g08130(.A1(new_n8322_), .A2(new_n1778_), .A3(new_n8262_), .ZN(new_n8323_));
  AOI21_X1   g08131(.A1(new_n8322_), .A2(new_n8262_), .B(new_n1778_), .ZN(new_n8324_));
  AOI21_X1   g08132(.A1(new_n8219_), .A2(new_n8323_), .B(new_n8324_), .ZN(new_n8325_));
  AOI21_X1   g08133(.A1(new_n8325_), .A2(new_n1632_), .B(new_n8305_), .ZN(new_n8326_));
  NOR3_X1    g08134(.A1(new_n8326_), .A2(\asqrt[50] ), .A3(new_n8267_), .ZN(new_n8327_));
  OAI21_X1   g08135(.A1(new_n8326_), .A2(new_n8267_), .B(\asqrt[50] ), .ZN(new_n8328_));
  OAI21_X1   g08136(.A1(new_n8214_), .A2(new_n8327_), .B(new_n8328_), .ZN(new_n8329_));
  OAI21_X1   g08137(.A1(new_n8329_), .A2(\asqrt[51] ), .B(new_n8209_), .ZN(new_n8330_));
  NAND3_X1   g08138(.A1(new_n8330_), .A2(new_n1150_), .A3(new_n8274_), .ZN(new_n8331_));
  AOI21_X1   g08139(.A1(new_n8330_), .A2(new_n8274_), .B(new_n1150_), .ZN(new_n8332_));
  AOI21_X1   g08140(.A1(new_n8207_), .A2(new_n8331_), .B(new_n8332_), .ZN(new_n8333_));
  AOI21_X1   g08141(.A1(new_n8333_), .A2(new_n1006_), .B(new_n8304_), .ZN(new_n8334_));
  NOR3_X1    g08142(.A1(new_n8334_), .A2(\asqrt[54] ), .A3(new_n8279_), .ZN(new_n8335_));
  OAI21_X1   g08143(.A1(new_n8334_), .A2(new_n8279_), .B(\asqrt[54] ), .ZN(new_n8336_));
  OAI21_X1   g08144(.A1(new_n8202_), .A2(new_n8335_), .B(new_n8336_), .ZN(new_n8337_));
  OAI21_X1   g08145(.A1(new_n8337_), .A2(\asqrt[55] ), .B(new_n8197_), .ZN(new_n8338_));
  NAND3_X1   g08146(.A1(new_n8338_), .A2(new_n634_), .A3(new_n8286_), .ZN(new_n8339_));
  AOI21_X1   g08147(.A1(new_n8338_), .A2(new_n8286_), .B(new_n634_), .ZN(new_n8340_));
  AOI21_X1   g08148(.A1(new_n8195_), .A2(new_n8339_), .B(new_n8340_), .ZN(new_n8341_));
  AOI21_X1   g08149(.A1(new_n8341_), .A2(new_n531_), .B(new_n8303_), .ZN(new_n8342_));
  NOR3_X1    g08150(.A1(new_n8342_), .A2(\asqrt[58] ), .A3(new_n8291_), .ZN(new_n8343_));
  OAI21_X1   g08151(.A1(new_n8342_), .A2(new_n8291_), .B(\asqrt[58] ), .ZN(new_n8344_));
  OAI21_X1   g08152(.A1(new_n8190_), .A2(new_n8343_), .B(new_n8344_), .ZN(new_n8345_));
  OAI21_X1   g08153(.A1(new_n8345_), .A2(\asqrt[59] ), .B(new_n8185_), .ZN(new_n8346_));
  AOI21_X1   g08154(.A1(new_n8346_), .A2(new_n8299_), .B(new_n266_), .ZN(new_n8347_));
  OAI21_X1   g08155(.A1(new_n8302_), .A2(new_n8347_), .B(\asqrt[61] ), .ZN(new_n8348_));
  AOI21_X1   g08156(.A1(new_n7991_), .A2(new_n7985_), .B(\asqrt[25] ), .ZN(new_n8349_));
  XOR2_X1    g08157(.A1(new_n8349_), .A2(new_n7793_), .Z(new_n8350_));
  OAI21_X1   g08158(.A1(new_n8186_), .A2(new_n8297_), .B(new_n8299_), .ZN(new_n8351_));
  OAI21_X1   g08159(.A1(new_n8351_), .A2(\asqrt[60] ), .B(new_n8182_), .ZN(new_n8352_));
  OAI21_X1   g08160(.A1(new_n8298_), .A2(new_n8300_), .B(\asqrt[60] ), .ZN(new_n8353_));
  NAND3_X1   g08161(.A1(new_n8352_), .A2(new_n239_), .A3(new_n8353_), .ZN(new_n8354_));
  NAND2_X1   g08162(.A1(new_n8354_), .A2(new_n8350_), .ZN(new_n8355_));
  NAND2_X1   g08163(.A1(new_n8355_), .A2(new_n8348_), .ZN(new_n8356_));
  AOI21_X1   g08164(.A1(new_n8352_), .A2(new_n8353_), .B(new_n239_), .ZN(new_n8357_));
  NAND3_X1   g08165(.A1(new_n8346_), .A2(new_n266_), .A3(new_n8299_), .ZN(new_n8358_));
  AOI21_X1   g08166(.A1(new_n8182_), .A2(new_n8358_), .B(new_n8347_), .ZN(new_n8359_));
  INV_X1     g08167(.I(new_n8350_), .ZN(new_n8360_));
  AOI21_X1   g08168(.A1(new_n8359_), .A2(new_n239_), .B(new_n8360_), .ZN(new_n8361_));
  OAI21_X1   g08169(.A1(new_n8361_), .A2(new_n8357_), .B(new_n201_), .ZN(new_n8362_));
  NAND3_X1   g08170(.A1(new_n8355_), .A2(\asqrt[62] ), .A3(new_n8348_), .ZN(new_n8363_));
  AOI21_X1   g08171(.A1(new_n7984_), .A2(new_n8060_), .B(\asqrt[25] ), .ZN(new_n8364_));
  XOR2_X1    g08172(.A1(new_n8364_), .A2(new_n7988_), .Z(new_n8365_));
  INV_X1     g08173(.I(new_n8365_), .ZN(new_n8366_));
  AOI22_X1   g08174(.A1(new_n8362_), .A2(new_n8363_), .B1(new_n8356_), .B2(new_n8366_), .ZN(new_n8367_));
  NOR2_X1    g08175(.A1(new_n8003_), .A2(new_n7791_), .ZN(new_n8368_));
  OAI21_X1   g08176(.A1(\asqrt[25] ), .A2(new_n8368_), .B(new_n8010_), .ZN(new_n8369_));
  INV_X1     g08177(.I(new_n8369_), .ZN(new_n8370_));
  OAI21_X1   g08178(.A1(new_n8367_), .A2(new_n8179_), .B(new_n8370_), .ZN(new_n8371_));
  OAI21_X1   g08179(.A1(new_n8356_), .A2(\asqrt[62] ), .B(new_n8365_), .ZN(new_n8372_));
  NAND2_X1   g08180(.A1(new_n8356_), .A2(\asqrt[62] ), .ZN(new_n8373_));
  NAND3_X1   g08181(.A1(new_n8372_), .A2(new_n8373_), .A3(new_n8179_), .ZN(new_n8374_));
  NAND2_X1   g08182(.A1(new_n8077_), .A2(new_n7790_), .ZN(new_n8375_));
  XOR2_X1    g08183(.A1(new_n8003_), .A2(new_n7791_), .Z(new_n8376_));
  NAND3_X1   g08184(.A1(new_n8375_), .A2(\asqrt[63] ), .A3(new_n8376_), .ZN(new_n8377_));
  INV_X1     g08185(.I(new_n8075_), .ZN(new_n8378_));
  NAND4_X1   g08186(.A1(new_n8378_), .A2(new_n7791_), .A3(new_n8010_), .A4(new_n8017_), .ZN(new_n8379_));
  NAND2_X1   g08187(.A1(new_n8377_), .A2(new_n8379_), .ZN(new_n8380_));
  INV_X1     g08188(.I(new_n8380_), .ZN(new_n8381_));
  NAND4_X1   g08189(.A1(new_n8371_), .A2(new_n193_), .A3(new_n8374_), .A4(new_n8381_), .ZN(\asqrt[24] ));
  AOI21_X1   g08190(.A1(new_n8169_), .A2(new_n8173_), .B(\asqrt[24] ), .ZN(new_n8383_));
  XOR2_X1    g08191(.A1(new_n8383_), .A2(new_n8020_), .Z(new_n8384_));
  XOR2_X1    g08192(.A1(new_n8160_), .A2(\asqrt[39] ), .Z(new_n8385_));
  NOR2_X1    g08193(.A1(\asqrt[24] ), .A2(new_n8385_), .ZN(new_n8386_));
  XOR2_X1    g08194(.A1(new_n8386_), .A2(new_n8022_), .Z(new_n8387_));
  NOR2_X1    g08195(.A1(new_n8158_), .A2(new_n8167_), .ZN(new_n8388_));
  NOR2_X1    g08196(.A1(\asqrt[24] ), .A2(new_n8388_), .ZN(new_n8389_));
  XOR2_X1    g08197(.A1(new_n8389_), .A2(new_n8025_), .Z(new_n8390_));
  AOI21_X1   g08198(.A1(new_n8162_), .A2(new_n8166_), .B(\asqrt[24] ), .ZN(new_n8391_));
  XOR2_X1    g08199(.A1(new_n8391_), .A2(new_n8028_), .Z(new_n8392_));
  INV_X1     g08200(.I(new_n8392_), .ZN(new_n8393_));
  AOI21_X1   g08201(.A1(new_n8148_), .A2(new_n8156_), .B(\asqrt[24] ), .ZN(new_n8394_));
  XOR2_X1    g08202(.A1(new_n8394_), .A2(new_n8032_), .Z(new_n8395_));
  INV_X1     g08203(.I(new_n8395_), .ZN(new_n8396_));
  XOR2_X1    g08204(.A1(new_n8139_), .A2(\asqrt[35] ), .Z(new_n8397_));
  NOR2_X1    g08205(.A1(\asqrt[24] ), .A2(new_n8397_), .ZN(new_n8398_));
  XOR2_X1    g08206(.A1(new_n8398_), .A2(new_n8034_), .Z(new_n8399_));
  NOR2_X1    g08207(.A1(new_n8137_), .A2(new_n8146_), .ZN(new_n8400_));
  NOR2_X1    g08208(.A1(\asqrt[24] ), .A2(new_n8400_), .ZN(new_n8401_));
  XOR2_X1    g08209(.A1(new_n8401_), .A2(new_n8037_), .Z(new_n8402_));
  AOI21_X1   g08210(.A1(new_n8141_), .A2(new_n8145_), .B(\asqrt[24] ), .ZN(new_n8403_));
  XOR2_X1    g08211(.A1(new_n8403_), .A2(new_n8040_), .Z(new_n8404_));
  INV_X1     g08212(.I(new_n8404_), .ZN(new_n8405_));
  AOI21_X1   g08213(.A1(new_n8127_), .A2(new_n8135_), .B(\asqrt[24] ), .ZN(new_n8406_));
  XOR2_X1    g08214(.A1(new_n8406_), .A2(new_n8044_), .Z(new_n8407_));
  INV_X1     g08215(.I(new_n8407_), .ZN(new_n8408_));
  XOR2_X1    g08216(.A1(new_n8118_), .A2(\asqrt[31] ), .Z(new_n8409_));
  NOR2_X1    g08217(.A1(\asqrt[24] ), .A2(new_n8409_), .ZN(new_n8410_));
  XOR2_X1    g08218(.A1(new_n8410_), .A2(new_n8046_), .Z(new_n8411_));
  NOR2_X1    g08219(.A1(new_n8116_), .A2(new_n8125_), .ZN(new_n8412_));
  NOR2_X1    g08220(.A1(\asqrt[24] ), .A2(new_n8412_), .ZN(new_n8413_));
  XOR2_X1    g08221(.A1(new_n8413_), .A2(new_n8049_), .Z(new_n8414_));
  AOI21_X1   g08222(.A1(new_n8120_), .A2(new_n8124_), .B(\asqrt[24] ), .ZN(new_n8415_));
  XOR2_X1    g08223(.A1(new_n8415_), .A2(new_n8052_), .Z(new_n8416_));
  INV_X1     g08224(.I(new_n8416_), .ZN(new_n8417_));
  AOI21_X1   g08225(.A1(new_n8106_), .A2(new_n8114_), .B(\asqrt[24] ), .ZN(new_n8418_));
  XOR2_X1    g08226(.A1(new_n8418_), .A2(new_n8059_), .Z(new_n8419_));
  INV_X1     g08227(.I(new_n8419_), .ZN(new_n8420_));
  AOI21_X1   g08228(.A1(new_n8096_), .A2(new_n8105_), .B(\asqrt[24] ), .ZN(new_n8421_));
  XOR2_X1    g08229(.A1(new_n8421_), .A2(new_n8080_), .Z(new_n8422_));
  NAND2_X1   g08230(.A1(\asqrt[25] ), .A2(new_n8081_), .ZN(new_n8423_));
  NOR2_X1    g08231(.A1(new_n8093_), .A2(\a[50] ), .ZN(new_n8424_));
  AOI22_X1   g08232(.A1(new_n8423_), .A2(new_n8093_), .B1(\asqrt[25] ), .B2(new_n8424_), .ZN(new_n8425_));
  OAI21_X1   g08233(.A1(new_n8077_), .A2(new_n8081_), .B(new_n8090_), .ZN(new_n8426_));
  AOI21_X1   g08234(.A1(new_n8086_), .A2(new_n8426_), .B(\asqrt[24] ), .ZN(new_n8427_));
  XOR2_X1    g08235(.A1(new_n8427_), .A2(new_n8425_), .Z(new_n8428_));
  NAND2_X1   g08236(.A1(new_n8371_), .A2(new_n193_), .ZN(new_n8429_));
  NOR2_X1    g08237(.A1(new_n8361_), .A2(new_n8357_), .ZN(new_n8430_));
  AOI21_X1   g08238(.A1(new_n8430_), .A2(new_n201_), .B(new_n8366_), .ZN(new_n8431_));
  OAI21_X1   g08239(.A1(new_n8430_), .A2(new_n201_), .B(new_n8179_), .ZN(new_n8432_));
  NOR2_X1    g08240(.A1(new_n8431_), .A2(new_n8432_), .ZN(new_n8433_));
  NAND3_X1   g08241(.A1(new_n8377_), .A2(\asqrt[25] ), .A3(new_n8379_), .ZN(new_n8434_));
  NOR3_X1    g08242(.A1(new_n8429_), .A2(new_n8433_), .A3(new_n8434_), .ZN(new_n8435_));
  AOI21_X1   g08243(.A1(new_n8355_), .A2(new_n8348_), .B(\asqrt[62] ), .ZN(new_n8436_));
  NOR3_X1    g08244(.A1(new_n8361_), .A2(new_n201_), .A3(new_n8357_), .ZN(new_n8437_));
  OAI22_X1   g08245(.A1(new_n8437_), .A2(new_n8436_), .B1(new_n8430_), .B2(new_n8365_), .ZN(new_n8438_));
  AOI21_X1   g08246(.A1(new_n8438_), .A2(new_n8178_), .B(new_n8369_), .ZN(new_n8439_));
  NOR4_X1    g08247(.A1(new_n8439_), .A2(\asqrt[63] ), .A3(new_n8433_), .A4(new_n8380_), .ZN(new_n8440_));
  NOR2_X1    g08248(.A1(new_n8440_), .A2(new_n8084_), .ZN(new_n8441_));
  OAI21_X1   g08249(.A1(new_n8441_), .A2(new_n8435_), .B(new_n8081_), .ZN(new_n8442_));
  NOR3_X1    g08250(.A1(new_n8439_), .A2(\asqrt[63] ), .A3(new_n8433_), .ZN(new_n8443_));
  NAND4_X1   g08251(.A1(new_n8443_), .A2(\asqrt[25] ), .A3(new_n8377_), .A4(new_n8379_), .ZN(new_n8444_));
  NAND2_X1   g08252(.A1(\asqrt[24] ), .A2(new_n8082_), .ZN(new_n8445_));
  NAND3_X1   g08253(.A1(new_n8444_), .A2(new_n8445_), .A3(\a[50] ), .ZN(new_n8446_));
  NAND2_X1   g08254(.A1(new_n8446_), .A2(new_n8442_), .ZN(new_n8447_));
  NOR2_X1    g08255(.A1(\a[46] ), .A2(\a[47] ), .ZN(new_n8448_));
  INV_X1     g08256(.I(new_n8448_), .ZN(new_n8449_));
  NAND3_X1   g08257(.A1(\asqrt[24] ), .A2(\a[48] ), .A3(new_n8449_), .ZN(new_n8450_));
  INV_X1     g08258(.I(\a[48] ), .ZN(new_n8451_));
  OAI21_X1   g08259(.A1(\asqrt[24] ), .A2(new_n8451_), .B(new_n8448_), .ZN(new_n8452_));
  AOI21_X1   g08260(.A1(new_n8452_), .A2(new_n8450_), .B(new_n8077_), .ZN(new_n8453_));
  NAND2_X1   g08261(.A1(new_n8448_), .A2(new_n8451_), .ZN(new_n8454_));
  NAND3_X1   g08262(.A1(new_n8013_), .A2(new_n8015_), .A3(new_n8454_), .ZN(new_n8455_));
  NAND2_X1   g08263(.A1(new_n8069_), .A2(new_n8455_), .ZN(new_n8456_));
  NAND3_X1   g08264(.A1(\asqrt[24] ), .A2(\a[48] ), .A3(new_n8456_), .ZN(new_n8457_));
  INV_X1     g08265(.I(\a[49] ), .ZN(new_n8458_));
  NAND3_X1   g08266(.A1(\asqrt[24] ), .A2(new_n8451_), .A3(new_n8458_), .ZN(new_n8459_));
  OAI21_X1   g08267(.A1(new_n8440_), .A2(\a[48] ), .B(\a[49] ), .ZN(new_n8460_));
  NAND3_X1   g08268(.A1(new_n8460_), .A2(new_n8457_), .A3(new_n8459_), .ZN(new_n8461_));
  NOR3_X1    g08269(.A1(new_n8461_), .A2(new_n8453_), .A3(\asqrt[26] ), .ZN(new_n8462_));
  OAI21_X1   g08270(.A1(new_n8461_), .A2(new_n8453_), .B(\asqrt[26] ), .ZN(new_n8463_));
  OAI21_X1   g08271(.A1(new_n8447_), .A2(new_n8462_), .B(new_n8463_), .ZN(new_n8464_));
  OAI21_X1   g08272(.A1(new_n8464_), .A2(\asqrt[27] ), .B(new_n8428_), .ZN(new_n8465_));
  NAND2_X1   g08273(.A1(new_n8464_), .A2(\asqrt[27] ), .ZN(new_n8466_));
  NAND3_X1   g08274(.A1(new_n8465_), .A2(new_n8466_), .A3(new_n6966_), .ZN(new_n8467_));
  AOI21_X1   g08275(.A1(new_n8465_), .A2(new_n8466_), .B(new_n6966_), .ZN(new_n8468_));
  AOI21_X1   g08276(.A1(new_n8422_), .A2(new_n8467_), .B(new_n8468_), .ZN(new_n8469_));
  AOI21_X1   g08277(.A1(new_n8469_), .A2(new_n6636_), .B(new_n8420_), .ZN(new_n8470_));
  NAND2_X1   g08278(.A1(new_n8467_), .A2(new_n8422_), .ZN(new_n8471_));
  INV_X1     g08279(.I(new_n8428_), .ZN(new_n8472_));
  INV_X1     g08280(.I(new_n8447_), .ZN(new_n8473_));
  NOR3_X1    g08281(.A1(new_n8440_), .A2(new_n8451_), .A3(new_n8448_), .ZN(new_n8474_));
  AOI21_X1   g08282(.A1(new_n8440_), .A2(\a[48] ), .B(new_n8449_), .ZN(new_n8475_));
  OAI21_X1   g08283(.A1(new_n8474_), .A2(new_n8475_), .B(\asqrt[25] ), .ZN(new_n8476_));
  INV_X1     g08284(.I(new_n8456_), .ZN(new_n8477_));
  NOR3_X1    g08285(.A1(new_n8440_), .A2(new_n8451_), .A3(new_n8477_), .ZN(new_n8478_));
  NOR3_X1    g08286(.A1(new_n8440_), .A2(\a[48] ), .A3(\a[49] ), .ZN(new_n8479_));
  AOI21_X1   g08287(.A1(\asqrt[24] ), .A2(new_n8451_), .B(new_n8458_), .ZN(new_n8480_));
  NOR3_X1    g08288(.A1(new_n8478_), .A2(new_n8479_), .A3(new_n8480_), .ZN(new_n8481_));
  NAND3_X1   g08289(.A1(new_n8476_), .A2(new_n8481_), .A3(new_n7690_), .ZN(new_n8482_));
  AOI21_X1   g08290(.A1(new_n8476_), .A2(new_n8481_), .B(new_n7690_), .ZN(new_n8483_));
  AOI21_X1   g08291(.A1(new_n8473_), .A2(new_n8482_), .B(new_n8483_), .ZN(new_n8484_));
  AOI21_X1   g08292(.A1(new_n8484_), .A2(new_n7331_), .B(new_n8472_), .ZN(new_n8485_));
  NAND2_X1   g08293(.A1(new_n8473_), .A2(new_n8482_), .ZN(new_n8486_));
  AOI21_X1   g08294(.A1(new_n8486_), .A2(new_n8463_), .B(new_n7331_), .ZN(new_n8487_));
  OAI21_X1   g08295(.A1(new_n8485_), .A2(new_n8487_), .B(\asqrt[28] ), .ZN(new_n8488_));
  AOI21_X1   g08296(.A1(new_n8471_), .A2(new_n8488_), .B(new_n6636_), .ZN(new_n8489_));
  NOR3_X1    g08297(.A1(new_n8470_), .A2(\asqrt[30] ), .A3(new_n8489_), .ZN(new_n8490_));
  OAI21_X1   g08298(.A1(new_n8470_), .A2(new_n8489_), .B(\asqrt[30] ), .ZN(new_n8491_));
  OAI21_X1   g08299(.A1(new_n8417_), .A2(new_n8490_), .B(new_n8491_), .ZN(new_n8492_));
  OAI21_X1   g08300(.A1(new_n8492_), .A2(\asqrt[31] ), .B(new_n8414_), .ZN(new_n8493_));
  NAND2_X1   g08301(.A1(new_n8492_), .A2(\asqrt[31] ), .ZN(new_n8494_));
  NAND3_X1   g08302(.A1(new_n8493_), .A2(new_n8494_), .A3(new_n5643_), .ZN(new_n8495_));
  AOI21_X1   g08303(.A1(new_n8493_), .A2(new_n8494_), .B(new_n5643_), .ZN(new_n8496_));
  AOI21_X1   g08304(.A1(new_n8411_), .A2(new_n8495_), .B(new_n8496_), .ZN(new_n8497_));
  AOI21_X1   g08305(.A1(new_n8497_), .A2(new_n5336_), .B(new_n8408_), .ZN(new_n8498_));
  NAND2_X1   g08306(.A1(new_n8495_), .A2(new_n8411_), .ZN(new_n8499_));
  INV_X1     g08307(.I(new_n8414_), .ZN(new_n8500_));
  INV_X1     g08308(.I(new_n8422_), .ZN(new_n8501_));
  NOR3_X1    g08309(.A1(new_n8485_), .A2(\asqrt[28] ), .A3(new_n8487_), .ZN(new_n8502_));
  OAI21_X1   g08310(.A1(new_n8501_), .A2(new_n8502_), .B(new_n8488_), .ZN(new_n8503_));
  OAI21_X1   g08311(.A1(new_n8503_), .A2(\asqrt[29] ), .B(new_n8419_), .ZN(new_n8504_));
  NAND2_X1   g08312(.A1(new_n8503_), .A2(\asqrt[29] ), .ZN(new_n8505_));
  NAND3_X1   g08313(.A1(new_n8504_), .A2(new_n8505_), .A3(new_n6275_), .ZN(new_n8506_));
  AOI21_X1   g08314(.A1(new_n8504_), .A2(new_n8505_), .B(new_n6275_), .ZN(new_n8507_));
  AOI21_X1   g08315(.A1(new_n8416_), .A2(new_n8506_), .B(new_n8507_), .ZN(new_n8508_));
  AOI21_X1   g08316(.A1(new_n8508_), .A2(new_n5947_), .B(new_n8500_), .ZN(new_n8509_));
  NAND2_X1   g08317(.A1(new_n8506_), .A2(new_n8416_), .ZN(new_n8510_));
  AOI21_X1   g08318(.A1(new_n8510_), .A2(new_n8491_), .B(new_n5947_), .ZN(new_n8511_));
  OAI21_X1   g08319(.A1(new_n8509_), .A2(new_n8511_), .B(\asqrt[32] ), .ZN(new_n8512_));
  AOI21_X1   g08320(.A1(new_n8499_), .A2(new_n8512_), .B(new_n5336_), .ZN(new_n8513_));
  NOR3_X1    g08321(.A1(new_n8498_), .A2(\asqrt[34] ), .A3(new_n8513_), .ZN(new_n8514_));
  OAI21_X1   g08322(.A1(new_n8498_), .A2(new_n8513_), .B(\asqrt[34] ), .ZN(new_n8515_));
  OAI21_X1   g08323(.A1(new_n8405_), .A2(new_n8514_), .B(new_n8515_), .ZN(new_n8516_));
  OAI21_X1   g08324(.A1(new_n8516_), .A2(\asqrt[35] ), .B(new_n8402_), .ZN(new_n8517_));
  NAND2_X1   g08325(.A1(new_n8516_), .A2(\asqrt[35] ), .ZN(new_n8518_));
  NAND3_X1   g08326(.A1(new_n8517_), .A2(new_n8518_), .A3(new_n4461_), .ZN(new_n8519_));
  AOI21_X1   g08327(.A1(new_n8517_), .A2(new_n8518_), .B(new_n4461_), .ZN(new_n8520_));
  AOI21_X1   g08328(.A1(new_n8399_), .A2(new_n8519_), .B(new_n8520_), .ZN(new_n8521_));
  AOI21_X1   g08329(.A1(new_n8521_), .A2(new_n4196_), .B(new_n8396_), .ZN(new_n8522_));
  NAND2_X1   g08330(.A1(new_n8519_), .A2(new_n8399_), .ZN(new_n8523_));
  INV_X1     g08331(.I(new_n8402_), .ZN(new_n8524_));
  INV_X1     g08332(.I(new_n8411_), .ZN(new_n8525_));
  NOR3_X1    g08333(.A1(new_n8509_), .A2(\asqrt[32] ), .A3(new_n8511_), .ZN(new_n8526_));
  OAI21_X1   g08334(.A1(new_n8525_), .A2(new_n8526_), .B(new_n8512_), .ZN(new_n8527_));
  OAI21_X1   g08335(.A1(new_n8527_), .A2(\asqrt[33] ), .B(new_n8407_), .ZN(new_n8528_));
  NAND2_X1   g08336(.A1(new_n8527_), .A2(\asqrt[33] ), .ZN(new_n8529_));
  NAND3_X1   g08337(.A1(new_n8528_), .A2(new_n8529_), .A3(new_n5029_), .ZN(new_n8530_));
  AOI21_X1   g08338(.A1(new_n8528_), .A2(new_n8529_), .B(new_n5029_), .ZN(new_n8531_));
  AOI21_X1   g08339(.A1(new_n8404_), .A2(new_n8530_), .B(new_n8531_), .ZN(new_n8532_));
  AOI21_X1   g08340(.A1(new_n8532_), .A2(new_n4751_), .B(new_n8524_), .ZN(new_n8533_));
  NAND2_X1   g08341(.A1(new_n8530_), .A2(new_n8404_), .ZN(new_n8534_));
  AOI21_X1   g08342(.A1(new_n8534_), .A2(new_n8515_), .B(new_n4751_), .ZN(new_n8535_));
  OAI21_X1   g08343(.A1(new_n8533_), .A2(new_n8535_), .B(\asqrt[36] ), .ZN(new_n8536_));
  AOI21_X1   g08344(.A1(new_n8523_), .A2(new_n8536_), .B(new_n4196_), .ZN(new_n8537_));
  NOR3_X1    g08345(.A1(new_n8522_), .A2(\asqrt[38] ), .A3(new_n8537_), .ZN(new_n8538_));
  OAI21_X1   g08346(.A1(new_n8522_), .A2(new_n8537_), .B(\asqrt[38] ), .ZN(new_n8539_));
  OAI21_X1   g08347(.A1(new_n8393_), .A2(new_n8538_), .B(new_n8539_), .ZN(new_n8540_));
  OAI21_X1   g08348(.A1(new_n8540_), .A2(\asqrt[39] ), .B(new_n8390_), .ZN(new_n8541_));
  NAND2_X1   g08349(.A1(new_n8540_), .A2(\asqrt[39] ), .ZN(new_n8542_));
  NAND3_X1   g08350(.A1(new_n8541_), .A2(new_n8542_), .A3(new_n3427_), .ZN(new_n8543_));
  AOI21_X1   g08351(.A1(new_n8541_), .A2(new_n8542_), .B(new_n3427_), .ZN(new_n8544_));
  AOI21_X1   g08352(.A1(new_n8387_), .A2(new_n8543_), .B(new_n8544_), .ZN(new_n8545_));
  NAND2_X1   g08353(.A1(new_n8545_), .A2(new_n3195_), .ZN(new_n8546_));
  INV_X1     g08354(.I(new_n8387_), .ZN(new_n8547_));
  INV_X1     g08355(.I(new_n8390_), .ZN(new_n8548_));
  INV_X1     g08356(.I(new_n8399_), .ZN(new_n8549_));
  NOR3_X1    g08357(.A1(new_n8533_), .A2(\asqrt[36] ), .A3(new_n8535_), .ZN(new_n8550_));
  OAI21_X1   g08358(.A1(new_n8549_), .A2(new_n8550_), .B(new_n8536_), .ZN(new_n8551_));
  OAI21_X1   g08359(.A1(new_n8551_), .A2(\asqrt[37] ), .B(new_n8395_), .ZN(new_n8552_));
  NAND2_X1   g08360(.A1(new_n8551_), .A2(\asqrt[37] ), .ZN(new_n8553_));
  NAND3_X1   g08361(.A1(new_n8552_), .A2(new_n8553_), .A3(new_n3925_), .ZN(new_n8554_));
  AOI21_X1   g08362(.A1(new_n8552_), .A2(new_n8553_), .B(new_n3925_), .ZN(new_n8555_));
  AOI21_X1   g08363(.A1(new_n8392_), .A2(new_n8554_), .B(new_n8555_), .ZN(new_n8556_));
  AOI21_X1   g08364(.A1(new_n8556_), .A2(new_n3681_), .B(new_n8548_), .ZN(new_n8557_));
  NAND2_X1   g08365(.A1(new_n8554_), .A2(new_n8392_), .ZN(new_n8558_));
  AOI21_X1   g08366(.A1(new_n8558_), .A2(new_n8539_), .B(new_n3681_), .ZN(new_n8559_));
  NOR3_X1    g08367(.A1(new_n8557_), .A2(\asqrt[40] ), .A3(new_n8559_), .ZN(new_n8560_));
  OAI21_X1   g08368(.A1(new_n8557_), .A2(new_n8559_), .B(\asqrt[40] ), .ZN(new_n8561_));
  OAI21_X1   g08369(.A1(new_n8547_), .A2(new_n8560_), .B(new_n8561_), .ZN(new_n8562_));
  NAND2_X1   g08370(.A1(new_n8562_), .A2(\asqrt[41] ), .ZN(new_n8563_));
  NOR2_X1    g08371(.A1(new_n8356_), .A2(\asqrt[62] ), .ZN(new_n8564_));
  INV_X1     g08372(.I(new_n8373_), .ZN(new_n8565_));
  NOR2_X1    g08373(.A1(new_n8565_), .A2(new_n8564_), .ZN(new_n8566_));
  XOR2_X1    g08374(.A1(new_n8364_), .A2(new_n7988_), .Z(new_n8567_));
  OAI21_X1   g08375(.A1(\asqrt[24] ), .A2(new_n8566_), .B(new_n8567_), .ZN(new_n8568_));
  INV_X1     g08376(.I(new_n8568_), .ZN(new_n8569_));
  NOR2_X1    g08377(.A1(new_n8300_), .A2(new_n8297_), .ZN(new_n8570_));
  NOR2_X1    g08378(.A1(\asqrt[24] ), .A2(new_n8570_), .ZN(new_n8571_));
  XOR2_X1    g08379(.A1(new_n8571_), .A2(new_n8185_), .Z(new_n8572_));
  INV_X1     g08380(.I(new_n8572_), .ZN(new_n8573_));
  NOR2_X1    g08381(.A1(new_n8343_), .A2(new_n8296_), .ZN(new_n8574_));
  NOR2_X1    g08382(.A1(\asqrt[24] ), .A2(new_n8574_), .ZN(new_n8575_));
  XOR2_X1    g08383(.A1(new_n8575_), .A2(new_n8189_), .Z(new_n8576_));
  AOI21_X1   g08384(.A1(new_n8290_), .A2(new_n8295_), .B(\asqrt[24] ), .ZN(new_n8577_));
  XOR2_X1    g08385(.A1(new_n8577_), .A2(new_n8192_), .Z(new_n8578_));
  AOI21_X1   g08386(.A1(new_n8339_), .A2(new_n8289_), .B(\asqrt[24] ), .ZN(new_n8579_));
  XOR2_X1    g08387(.A1(new_n8579_), .A2(new_n8195_), .Z(new_n8580_));
  INV_X1     g08388(.I(new_n8286_), .ZN(new_n8581_));
  NOR2_X1    g08389(.A1(new_n8581_), .A2(new_n8285_), .ZN(new_n8582_));
  NOR2_X1    g08390(.A1(\asqrt[24] ), .A2(new_n8582_), .ZN(new_n8583_));
  XOR2_X1    g08391(.A1(new_n8583_), .A2(new_n8197_), .Z(new_n8584_));
  INV_X1     g08392(.I(new_n8584_), .ZN(new_n8585_));
  NOR2_X1    g08393(.A1(new_n8335_), .A2(new_n8284_), .ZN(new_n8586_));
  NOR2_X1    g08394(.A1(\asqrt[24] ), .A2(new_n8586_), .ZN(new_n8587_));
  XOR2_X1    g08395(.A1(new_n8587_), .A2(new_n8201_), .Z(new_n8588_));
  INV_X1     g08396(.I(new_n8588_), .ZN(new_n8589_));
  AOI21_X1   g08397(.A1(new_n8278_), .A2(new_n8283_), .B(\asqrt[24] ), .ZN(new_n8590_));
  XOR2_X1    g08398(.A1(new_n8590_), .A2(new_n8204_), .Z(new_n8591_));
  AOI21_X1   g08399(.A1(new_n8331_), .A2(new_n8277_), .B(\asqrt[24] ), .ZN(new_n8592_));
  XOR2_X1    g08400(.A1(new_n8592_), .A2(new_n8207_), .Z(new_n8593_));
  XOR2_X1    g08401(.A1(new_n8329_), .A2(\asqrt[51] ), .Z(new_n8594_));
  NOR2_X1    g08402(.A1(\asqrt[24] ), .A2(new_n8594_), .ZN(new_n8595_));
  XOR2_X1    g08403(.A1(new_n8595_), .A2(new_n8209_), .Z(new_n8596_));
  INV_X1     g08404(.I(new_n8596_), .ZN(new_n8597_));
  NOR2_X1    g08405(.A1(new_n8327_), .A2(new_n8272_), .ZN(new_n8598_));
  NOR2_X1    g08406(.A1(\asqrt[24] ), .A2(new_n8598_), .ZN(new_n8599_));
  XOR2_X1    g08407(.A1(new_n8599_), .A2(new_n8213_), .Z(new_n8600_));
  INV_X1     g08408(.I(new_n8600_), .ZN(new_n8601_));
  AOI21_X1   g08409(.A1(new_n8266_), .A2(new_n8271_), .B(\asqrt[24] ), .ZN(new_n8602_));
  XOR2_X1    g08410(.A1(new_n8602_), .A2(new_n8216_), .Z(new_n8603_));
  AOI21_X1   g08411(.A1(new_n8323_), .A2(new_n8265_), .B(\asqrt[24] ), .ZN(new_n8604_));
  XOR2_X1    g08412(.A1(new_n8604_), .A2(new_n8219_), .Z(new_n8605_));
  XOR2_X1    g08413(.A1(new_n8321_), .A2(\asqrt[47] ), .Z(new_n8606_));
  NOR2_X1    g08414(.A1(\asqrt[24] ), .A2(new_n8606_), .ZN(new_n8607_));
  XOR2_X1    g08415(.A1(new_n8607_), .A2(new_n8221_), .Z(new_n8608_));
  INV_X1     g08416(.I(new_n8608_), .ZN(new_n8609_));
  NOR2_X1    g08417(.A1(new_n8319_), .A2(new_n8260_), .ZN(new_n8610_));
  NOR2_X1    g08418(.A1(\asqrt[24] ), .A2(new_n8610_), .ZN(new_n8611_));
  XOR2_X1    g08419(.A1(new_n8611_), .A2(new_n8225_), .Z(new_n8612_));
  INV_X1     g08420(.I(new_n8612_), .ZN(new_n8613_));
  AOI21_X1   g08421(.A1(new_n8254_), .A2(new_n8259_), .B(\asqrt[24] ), .ZN(new_n8614_));
  XOR2_X1    g08422(.A1(new_n8614_), .A2(new_n8228_), .Z(new_n8615_));
  AOI21_X1   g08423(.A1(new_n8315_), .A2(new_n8253_), .B(\asqrt[24] ), .ZN(new_n8616_));
  XOR2_X1    g08424(.A1(new_n8616_), .A2(new_n8231_), .Z(new_n8617_));
  XOR2_X1    g08425(.A1(new_n8313_), .A2(\asqrt[43] ), .Z(new_n8618_));
  NOR2_X1    g08426(.A1(\asqrt[24] ), .A2(new_n8618_), .ZN(new_n8619_));
  XOR2_X1    g08427(.A1(new_n8619_), .A2(new_n8233_), .Z(new_n8620_));
  INV_X1     g08428(.I(new_n8620_), .ZN(new_n8621_));
  NOR2_X1    g08429(.A1(new_n8311_), .A2(new_n8248_), .ZN(new_n8622_));
  NOR2_X1    g08430(.A1(\asqrt[24] ), .A2(new_n8622_), .ZN(new_n8623_));
  XOR2_X1    g08431(.A1(new_n8623_), .A2(new_n8237_), .Z(new_n8624_));
  INV_X1     g08432(.I(new_n8624_), .ZN(new_n8625_));
  AOI21_X1   g08433(.A1(new_n8242_), .A2(new_n8247_), .B(\asqrt[24] ), .ZN(new_n8626_));
  XOR2_X1    g08434(.A1(new_n8626_), .A2(new_n8240_), .Z(new_n8627_));
  OAI21_X1   g08435(.A1(new_n8562_), .A2(\asqrt[41] ), .B(new_n8384_), .ZN(new_n8628_));
  NAND3_X1   g08436(.A1(new_n8628_), .A2(new_n8563_), .A3(new_n2960_), .ZN(new_n8629_));
  AOI21_X1   g08437(.A1(new_n8628_), .A2(new_n8563_), .B(new_n2960_), .ZN(new_n8630_));
  AOI21_X1   g08438(.A1(new_n8627_), .A2(new_n8629_), .B(new_n8630_), .ZN(new_n8631_));
  AOI21_X1   g08439(.A1(new_n8631_), .A2(new_n2749_), .B(new_n8625_), .ZN(new_n8632_));
  NAND2_X1   g08440(.A1(new_n8629_), .A2(new_n8627_), .ZN(new_n8633_));
  INV_X1     g08441(.I(new_n8384_), .ZN(new_n8634_));
  AOI21_X1   g08442(.A1(new_n8545_), .A2(new_n3195_), .B(new_n8634_), .ZN(new_n8635_));
  NAND2_X1   g08443(.A1(new_n8543_), .A2(new_n8387_), .ZN(new_n8636_));
  AOI21_X1   g08444(.A1(new_n8636_), .A2(new_n8561_), .B(new_n3195_), .ZN(new_n8637_));
  OAI21_X1   g08445(.A1(new_n8635_), .A2(new_n8637_), .B(\asqrt[42] ), .ZN(new_n8638_));
  AOI21_X1   g08446(.A1(new_n8633_), .A2(new_n8638_), .B(new_n2749_), .ZN(new_n8639_));
  NOR3_X1    g08447(.A1(new_n8632_), .A2(\asqrt[44] ), .A3(new_n8639_), .ZN(new_n8640_));
  OAI21_X1   g08448(.A1(new_n8632_), .A2(new_n8639_), .B(\asqrt[44] ), .ZN(new_n8641_));
  OAI21_X1   g08449(.A1(new_n8621_), .A2(new_n8640_), .B(new_n8641_), .ZN(new_n8642_));
  OAI21_X1   g08450(.A1(new_n8642_), .A2(\asqrt[45] ), .B(new_n8617_), .ZN(new_n8643_));
  NAND2_X1   g08451(.A1(new_n8642_), .A2(\asqrt[45] ), .ZN(new_n8644_));
  NAND3_X1   g08452(.A1(new_n8643_), .A2(new_n8644_), .A3(new_n2134_), .ZN(new_n8645_));
  AOI21_X1   g08453(.A1(new_n8643_), .A2(new_n8644_), .B(new_n2134_), .ZN(new_n8646_));
  AOI21_X1   g08454(.A1(new_n8615_), .A2(new_n8645_), .B(new_n8646_), .ZN(new_n8647_));
  AOI21_X1   g08455(.A1(new_n8647_), .A2(new_n1953_), .B(new_n8613_), .ZN(new_n8648_));
  NAND2_X1   g08456(.A1(new_n8645_), .A2(new_n8615_), .ZN(new_n8649_));
  INV_X1     g08457(.I(new_n8617_), .ZN(new_n8650_));
  INV_X1     g08458(.I(new_n8627_), .ZN(new_n8651_));
  NOR3_X1    g08459(.A1(new_n8635_), .A2(\asqrt[42] ), .A3(new_n8637_), .ZN(new_n8652_));
  OAI21_X1   g08460(.A1(new_n8651_), .A2(new_n8652_), .B(new_n8638_), .ZN(new_n8653_));
  OAI21_X1   g08461(.A1(new_n8653_), .A2(\asqrt[43] ), .B(new_n8624_), .ZN(new_n8654_));
  NAND2_X1   g08462(.A1(new_n8653_), .A2(\asqrt[43] ), .ZN(new_n8655_));
  NAND3_X1   g08463(.A1(new_n8654_), .A2(new_n8655_), .A3(new_n2531_), .ZN(new_n8656_));
  AOI21_X1   g08464(.A1(new_n8654_), .A2(new_n8655_), .B(new_n2531_), .ZN(new_n8657_));
  AOI21_X1   g08465(.A1(new_n8620_), .A2(new_n8656_), .B(new_n8657_), .ZN(new_n8658_));
  AOI21_X1   g08466(.A1(new_n8658_), .A2(new_n2332_), .B(new_n8650_), .ZN(new_n8659_));
  NAND2_X1   g08467(.A1(new_n8656_), .A2(new_n8620_), .ZN(new_n8660_));
  AOI21_X1   g08468(.A1(new_n8660_), .A2(new_n8641_), .B(new_n2332_), .ZN(new_n8661_));
  OAI21_X1   g08469(.A1(new_n8659_), .A2(new_n8661_), .B(\asqrt[46] ), .ZN(new_n8662_));
  AOI21_X1   g08470(.A1(new_n8649_), .A2(new_n8662_), .B(new_n1953_), .ZN(new_n8663_));
  NOR3_X1    g08471(.A1(new_n8648_), .A2(\asqrt[48] ), .A3(new_n8663_), .ZN(new_n8664_));
  OAI21_X1   g08472(.A1(new_n8648_), .A2(new_n8663_), .B(\asqrt[48] ), .ZN(new_n8665_));
  OAI21_X1   g08473(.A1(new_n8609_), .A2(new_n8664_), .B(new_n8665_), .ZN(new_n8666_));
  OAI21_X1   g08474(.A1(new_n8666_), .A2(\asqrt[49] ), .B(new_n8605_), .ZN(new_n8667_));
  NAND2_X1   g08475(.A1(new_n8666_), .A2(\asqrt[49] ), .ZN(new_n8668_));
  NAND3_X1   g08476(.A1(new_n8667_), .A2(new_n8668_), .A3(new_n1463_), .ZN(new_n8669_));
  AOI21_X1   g08477(.A1(new_n8667_), .A2(new_n8668_), .B(new_n1463_), .ZN(new_n8670_));
  AOI21_X1   g08478(.A1(new_n8603_), .A2(new_n8669_), .B(new_n8670_), .ZN(new_n8671_));
  AOI21_X1   g08479(.A1(new_n8671_), .A2(new_n1305_), .B(new_n8601_), .ZN(new_n8672_));
  NAND2_X1   g08480(.A1(new_n8669_), .A2(new_n8603_), .ZN(new_n8673_));
  INV_X1     g08481(.I(new_n8605_), .ZN(new_n8674_));
  INV_X1     g08482(.I(new_n8615_), .ZN(new_n8675_));
  NOR3_X1    g08483(.A1(new_n8659_), .A2(\asqrt[46] ), .A3(new_n8661_), .ZN(new_n8676_));
  OAI21_X1   g08484(.A1(new_n8675_), .A2(new_n8676_), .B(new_n8662_), .ZN(new_n8677_));
  OAI21_X1   g08485(.A1(new_n8677_), .A2(\asqrt[47] ), .B(new_n8612_), .ZN(new_n8678_));
  NAND2_X1   g08486(.A1(new_n8677_), .A2(\asqrt[47] ), .ZN(new_n8679_));
  NAND3_X1   g08487(.A1(new_n8678_), .A2(new_n8679_), .A3(new_n1778_), .ZN(new_n8680_));
  AOI21_X1   g08488(.A1(new_n8678_), .A2(new_n8679_), .B(new_n1778_), .ZN(new_n8681_));
  AOI21_X1   g08489(.A1(new_n8608_), .A2(new_n8680_), .B(new_n8681_), .ZN(new_n8682_));
  AOI21_X1   g08490(.A1(new_n8682_), .A2(new_n1632_), .B(new_n8674_), .ZN(new_n8683_));
  NAND2_X1   g08491(.A1(new_n8680_), .A2(new_n8608_), .ZN(new_n8684_));
  AOI21_X1   g08492(.A1(new_n8684_), .A2(new_n8665_), .B(new_n1632_), .ZN(new_n8685_));
  OAI21_X1   g08493(.A1(new_n8683_), .A2(new_n8685_), .B(\asqrt[50] ), .ZN(new_n8686_));
  AOI21_X1   g08494(.A1(new_n8673_), .A2(new_n8686_), .B(new_n1305_), .ZN(new_n8687_));
  NOR3_X1    g08495(.A1(new_n8672_), .A2(\asqrt[52] ), .A3(new_n8687_), .ZN(new_n8688_));
  OAI21_X1   g08496(.A1(new_n8672_), .A2(new_n8687_), .B(\asqrt[52] ), .ZN(new_n8689_));
  OAI21_X1   g08497(.A1(new_n8597_), .A2(new_n8688_), .B(new_n8689_), .ZN(new_n8690_));
  OAI21_X1   g08498(.A1(new_n8690_), .A2(\asqrt[53] ), .B(new_n8593_), .ZN(new_n8691_));
  NAND2_X1   g08499(.A1(new_n8690_), .A2(\asqrt[53] ), .ZN(new_n8692_));
  NAND3_X1   g08500(.A1(new_n8691_), .A2(new_n8692_), .A3(new_n860_), .ZN(new_n8693_));
  AOI21_X1   g08501(.A1(new_n8691_), .A2(new_n8692_), .B(new_n860_), .ZN(new_n8694_));
  AOI21_X1   g08502(.A1(new_n8591_), .A2(new_n8693_), .B(new_n8694_), .ZN(new_n8695_));
  AOI21_X1   g08503(.A1(new_n8695_), .A2(new_n744_), .B(new_n8589_), .ZN(new_n8696_));
  NAND2_X1   g08504(.A1(new_n8693_), .A2(new_n8591_), .ZN(new_n8697_));
  INV_X1     g08505(.I(new_n8593_), .ZN(new_n8698_));
  INV_X1     g08506(.I(new_n8603_), .ZN(new_n8699_));
  NOR3_X1    g08507(.A1(new_n8683_), .A2(\asqrt[50] ), .A3(new_n8685_), .ZN(new_n8700_));
  OAI21_X1   g08508(.A1(new_n8699_), .A2(new_n8700_), .B(new_n8686_), .ZN(new_n8701_));
  OAI21_X1   g08509(.A1(new_n8701_), .A2(\asqrt[51] ), .B(new_n8600_), .ZN(new_n8702_));
  NAND2_X1   g08510(.A1(new_n8701_), .A2(\asqrt[51] ), .ZN(new_n8703_));
  NAND3_X1   g08511(.A1(new_n8702_), .A2(new_n8703_), .A3(new_n1150_), .ZN(new_n8704_));
  AOI21_X1   g08512(.A1(new_n8702_), .A2(new_n8703_), .B(new_n1150_), .ZN(new_n8705_));
  AOI21_X1   g08513(.A1(new_n8596_), .A2(new_n8704_), .B(new_n8705_), .ZN(new_n8706_));
  AOI21_X1   g08514(.A1(new_n8706_), .A2(new_n1006_), .B(new_n8698_), .ZN(new_n8707_));
  NAND2_X1   g08515(.A1(new_n8704_), .A2(new_n8596_), .ZN(new_n8708_));
  AOI21_X1   g08516(.A1(new_n8708_), .A2(new_n8689_), .B(new_n1006_), .ZN(new_n8709_));
  OAI21_X1   g08517(.A1(new_n8707_), .A2(new_n8709_), .B(\asqrt[54] ), .ZN(new_n8710_));
  AOI21_X1   g08518(.A1(new_n8697_), .A2(new_n8710_), .B(new_n744_), .ZN(new_n8711_));
  NOR3_X1    g08519(.A1(new_n8696_), .A2(\asqrt[56] ), .A3(new_n8711_), .ZN(new_n8712_));
  OAI21_X1   g08520(.A1(new_n8696_), .A2(new_n8711_), .B(\asqrt[56] ), .ZN(new_n8713_));
  OAI21_X1   g08521(.A1(new_n8585_), .A2(new_n8712_), .B(new_n8713_), .ZN(new_n8714_));
  OAI21_X1   g08522(.A1(new_n8714_), .A2(\asqrt[57] ), .B(new_n8580_), .ZN(new_n8715_));
  NOR2_X1    g08523(.A1(new_n8712_), .A2(new_n8585_), .ZN(new_n8716_));
  INV_X1     g08524(.I(new_n8591_), .ZN(new_n8717_));
  NOR3_X1    g08525(.A1(new_n8707_), .A2(\asqrt[54] ), .A3(new_n8709_), .ZN(new_n8718_));
  OAI21_X1   g08526(.A1(new_n8717_), .A2(new_n8718_), .B(new_n8710_), .ZN(new_n8719_));
  OAI21_X1   g08527(.A1(new_n8719_), .A2(\asqrt[55] ), .B(new_n8588_), .ZN(new_n8720_));
  NAND2_X1   g08528(.A1(new_n8719_), .A2(\asqrt[55] ), .ZN(new_n8721_));
  AOI21_X1   g08529(.A1(new_n8720_), .A2(new_n8721_), .B(new_n634_), .ZN(new_n8722_));
  OAI21_X1   g08530(.A1(new_n8716_), .A2(new_n8722_), .B(\asqrt[57] ), .ZN(new_n8723_));
  NAND3_X1   g08531(.A1(new_n8715_), .A2(new_n423_), .A3(new_n8723_), .ZN(new_n8724_));
  NAND2_X1   g08532(.A1(new_n8724_), .A2(new_n8578_), .ZN(new_n8725_));
  INV_X1     g08533(.I(new_n8580_), .ZN(new_n8726_));
  NAND3_X1   g08534(.A1(new_n8720_), .A2(new_n8721_), .A3(new_n634_), .ZN(new_n8727_));
  AOI21_X1   g08535(.A1(new_n8584_), .A2(new_n8727_), .B(new_n8722_), .ZN(new_n8728_));
  AOI21_X1   g08536(.A1(new_n8728_), .A2(new_n531_), .B(new_n8726_), .ZN(new_n8729_));
  NAND2_X1   g08537(.A1(new_n8727_), .A2(new_n8584_), .ZN(new_n8730_));
  AOI21_X1   g08538(.A1(new_n8730_), .A2(new_n8713_), .B(new_n531_), .ZN(new_n8731_));
  OAI21_X1   g08539(.A1(new_n8729_), .A2(new_n8731_), .B(\asqrt[58] ), .ZN(new_n8732_));
  NAND3_X1   g08540(.A1(new_n8725_), .A2(new_n337_), .A3(new_n8732_), .ZN(new_n8733_));
  AOI21_X1   g08541(.A1(new_n8725_), .A2(new_n8732_), .B(new_n337_), .ZN(new_n8734_));
  AOI21_X1   g08542(.A1(new_n8576_), .A2(new_n8733_), .B(new_n8734_), .ZN(new_n8735_));
  AOI21_X1   g08543(.A1(new_n8735_), .A2(new_n266_), .B(new_n8573_), .ZN(new_n8736_));
  INV_X1     g08544(.I(new_n8578_), .ZN(new_n8737_));
  NOR3_X1    g08545(.A1(new_n8729_), .A2(\asqrt[58] ), .A3(new_n8731_), .ZN(new_n8738_));
  OAI21_X1   g08546(.A1(new_n8737_), .A2(new_n8738_), .B(new_n8732_), .ZN(new_n8739_));
  OAI21_X1   g08547(.A1(new_n8739_), .A2(\asqrt[59] ), .B(new_n8576_), .ZN(new_n8740_));
  NAND2_X1   g08548(.A1(new_n8739_), .A2(\asqrt[59] ), .ZN(new_n8741_));
  AOI21_X1   g08549(.A1(new_n8740_), .A2(new_n8741_), .B(new_n266_), .ZN(new_n8742_));
  OAI21_X1   g08550(.A1(new_n8736_), .A2(new_n8742_), .B(\asqrt[61] ), .ZN(new_n8743_));
  AOI21_X1   g08551(.A1(new_n8358_), .A2(new_n8353_), .B(\asqrt[24] ), .ZN(new_n8744_));
  XOR2_X1    g08552(.A1(new_n8744_), .A2(new_n8182_), .Z(new_n8745_));
  INV_X1     g08553(.I(new_n8745_), .ZN(new_n8746_));
  NOR3_X1    g08554(.A1(new_n8736_), .A2(\asqrt[61] ), .A3(new_n8742_), .ZN(new_n8747_));
  OAI21_X1   g08555(.A1(new_n8746_), .A2(new_n8747_), .B(new_n8743_), .ZN(new_n8748_));
  NAND3_X1   g08556(.A1(new_n8740_), .A2(new_n8741_), .A3(new_n266_), .ZN(new_n8749_));
  NAND2_X1   g08557(.A1(new_n8749_), .A2(new_n8572_), .ZN(new_n8750_));
  INV_X1     g08558(.I(new_n8576_), .ZN(new_n8751_));
  AOI21_X1   g08559(.A1(new_n8715_), .A2(new_n8723_), .B(new_n423_), .ZN(new_n8752_));
  AOI21_X1   g08560(.A1(new_n8578_), .A2(new_n8724_), .B(new_n8752_), .ZN(new_n8753_));
  AOI21_X1   g08561(.A1(new_n8753_), .A2(new_n337_), .B(new_n8751_), .ZN(new_n8754_));
  OAI21_X1   g08562(.A1(new_n8754_), .A2(new_n8734_), .B(\asqrt[60] ), .ZN(new_n8755_));
  AOI21_X1   g08563(.A1(new_n8750_), .A2(new_n8755_), .B(new_n239_), .ZN(new_n8756_));
  AOI21_X1   g08564(.A1(new_n8572_), .A2(new_n8749_), .B(new_n8742_), .ZN(new_n8757_));
  AOI21_X1   g08565(.A1(new_n8757_), .A2(new_n239_), .B(new_n8746_), .ZN(new_n8758_));
  OAI21_X1   g08566(.A1(new_n8758_), .A2(new_n8756_), .B(new_n201_), .ZN(new_n8759_));
  NOR3_X1    g08567(.A1(new_n8754_), .A2(\asqrt[60] ), .A3(new_n8734_), .ZN(new_n8760_));
  OAI21_X1   g08568(.A1(new_n8573_), .A2(new_n8760_), .B(new_n8755_), .ZN(new_n8761_));
  OAI21_X1   g08569(.A1(new_n8761_), .A2(\asqrt[61] ), .B(new_n8745_), .ZN(new_n8762_));
  NAND3_X1   g08570(.A1(new_n8762_), .A2(\asqrt[62] ), .A3(new_n8743_), .ZN(new_n8763_));
  AOI21_X1   g08571(.A1(new_n8348_), .A2(new_n8354_), .B(\asqrt[24] ), .ZN(new_n8764_));
  XOR2_X1    g08572(.A1(new_n8764_), .A2(new_n8350_), .Z(new_n8765_));
  INV_X1     g08573(.I(new_n8765_), .ZN(new_n8766_));
  AOI22_X1   g08574(.A1(new_n8763_), .A2(new_n8759_), .B1(new_n8748_), .B2(new_n8766_), .ZN(new_n8767_));
  NOR2_X1    g08575(.A1(new_n8367_), .A2(new_n8179_), .ZN(new_n8768_));
  OAI21_X1   g08576(.A1(\asqrt[24] ), .A2(new_n8768_), .B(new_n8374_), .ZN(new_n8769_));
  INV_X1     g08577(.I(new_n8769_), .ZN(new_n8770_));
  OAI21_X1   g08578(.A1(new_n8767_), .A2(new_n8569_), .B(new_n8770_), .ZN(new_n8771_));
  OAI21_X1   g08579(.A1(new_n8748_), .A2(\asqrt[62] ), .B(new_n8765_), .ZN(new_n8772_));
  NAND2_X1   g08580(.A1(new_n8748_), .A2(\asqrt[62] ), .ZN(new_n8773_));
  NAND3_X1   g08581(.A1(new_n8772_), .A2(new_n8773_), .A3(new_n8569_), .ZN(new_n8774_));
  NAND2_X1   g08582(.A1(new_n8440_), .A2(new_n8178_), .ZN(new_n8775_));
  XOR2_X1    g08583(.A1(new_n8367_), .A2(new_n8179_), .Z(new_n8776_));
  NAND3_X1   g08584(.A1(new_n8775_), .A2(\asqrt[63] ), .A3(new_n8776_), .ZN(new_n8777_));
  INV_X1     g08585(.I(new_n8429_), .ZN(new_n8778_));
  NAND4_X1   g08586(.A1(new_n8778_), .A2(new_n8179_), .A3(new_n8374_), .A4(new_n8381_), .ZN(new_n8779_));
  NAND2_X1   g08587(.A1(new_n8777_), .A2(new_n8779_), .ZN(new_n8780_));
  INV_X1     g08588(.I(new_n8780_), .ZN(new_n8781_));
  NAND4_X1   g08589(.A1(new_n8771_), .A2(new_n193_), .A3(new_n8774_), .A4(new_n8781_), .ZN(\asqrt[23] ));
  AOI21_X1   g08590(.A1(new_n8546_), .A2(new_n8563_), .B(\asqrt[23] ), .ZN(new_n8783_));
  XOR2_X1    g08591(.A1(new_n8783_), .A2(new_n8384_), .Z(new_n8784_));
  AOI21_X1   g08592(.A1(new_n8543_), .A2(new_n8561_), .B(\asqrt[23] ), .ZN(new_n8785_));
  XOR2_X1    g08593(.A1(new_n8785_), .A2(new_n8387_), .Z(new_n8786_));
  NAND2_X1   g08594(.A1(new_n8556_), .A2(new_n3681_), .ZN(new_n8787_));
  AOI21_X1   g08595(.A1(new_n8787_), .A2(new_n8542_), .B(\asqrt[23] ), .ZN(new_n8788_));
  XOR2_X1    g08596(.A1(new_n8788_), .A2(new_n8390_), .Z(new_n8789_));
  INV_X1     g08597(.I(new_n8789_), .ZN(new_n8790_));
  AOI21_X1   g08598(.A1(new_n8554_), .A2(new_n8539_), .B(\asqrt[23] ), .ZN(new_n8791_));
  XOR2_X1    g08599(.A1(new_n8791_), .A2(new_n8392_), .Z(new_n8792_));
  INV_X1     g08600(.I(new_n8792_), .ZN(new_n8793_));
  NAND2_X1   g08601(.A1(new_n8521_), .A2(new_n4196_), .ZN(new_n8794_));
  AOI21_X1   g08602(.A1(new_n8794_), .A2(new_n8553_), .B(\asqrt[23] ), .ZN(new_n8795_));
  XOR2_X1    g08603(.A1(new_n8795_), .A2(new_n8395_), .Z(new_n8796_));
  AOI21_X1   g08604(.A1(new_n8519_), .A2(new_n8536_), .B(\asqrt[23] ), .ZN(new_n8797_));
  XOR2_X1    g08605(.A1(new_n8797_), .A2(new_n8399_), .Z(new_n8798_));
  NAND2_X1   g08606(.A1(new_n8532_), .A2(new_n4751_), .ZN(new_n8799_));
  AOI21_X1   g08607(.A1(new_n8799_), .A2(new_n8518_), .B(\asqrt[23] ), .ZN(new_n8800_));
  XOR2_X1    g08608(.A1(new_n8800_), .A2(new_n8402_), .Z(new_n8801_));
  INV_X1     g08609(.I(new_n8801_), .ZN(new_n8802_));
  AOI21_X1   g08610(.A1(new_n8530_), .A2(new_n8515_), .B(\asqrt[23] ), .ZN(new_n8803_));
  XOR2_X1    g08611(.A1(new_n8803_), .A2(new_n8404_), .Z(new_n8804_));
  INV_X1     g08612(.I(new_n8804_), .ZN(new_n8805_));
  NAND2_X1   g08613(.A1(new_n8497_), .A2(new_n5336_), .ZN(new_n8806_));
  AOI21_X1   g08614(.A1(new_n8806_), .A2(new_n8529_), .B(\asqrt[23] ), .ZN(new_n8807_));
  XOR2_X1    g08615(.A1(new_n8807_), .A2(new_n8407_), .Z(new_n8808_));
  AOI21_X1   g08616(.A1(new_n8495_), .A2(new_n8512_), .B(\asqrt[23] ), .ZN(new_n8809_));
  XOR2_X1    g08617(.A1(new_n8809_), .A2(new_n8411_), .Z(new_n8810_));
  NAND2_X1   g08618(.A1(new_n8508_), .A2(new_n5947_), .ZN(new_n8811_));
  AOI21_X1   g08619(.A1(new_n8811_), .A2(new_n8494_), .B(\asqrt[23] ), .ZN(new_n8812_));
  XOR2_X1    g08620(.A1(new_n8812_), .A2(new_n8414_), .Z(new_n8813_));
  INV_X1     g08621(.I(new_n8813_), .ZN(new_n8814_));
  AOI21_X1   g08622(.A1(new_n8506_), .A2(new_n8491_), .B(\asqrt[23] ), .ZN(new_n8815_));
  XOR2_X1    g08623(.A1(new_n8815_), .A2(new_n8416_), .Z(new_n8816_));
  INV_X1     g08624(.I(new_n8816_), .ZN(new_n8817_));
  NAND2_X1   g08625(.A1(new_n8469_), .A2(new_n6636_), .ZN(new_n8818_));
  AOI21_X1   g08626(.A1(new_n8818_), .A2(new_n8505_), .B(\asqrt[23] ), .ZN(new_n8819_));
  XOR2_X1    g08627(.A1(new_n8819_), .A2(new_n8419_), .Z(new_n8820_));
  AOI21_X1   g08628(.A1(new_n8467_), .A2(new_n8488_), .B(\asqrt[23] ), .ZN(new_n8821_));
  XOR2_X1    g08629(.A1(new_n8821_), .A2(new_n8422_), .Z(new_n8822_));
  NAND2_X1   g08630(.A1(new_n8484_), .A2(new_n7331_), .ZN(new_n8823_));
  AOI21_X1   g08631(.A1(new_n8823_), .A2(new_n8466_), .B(\asqrt[23] ), .ZN(new_n8824_));
  XOR2_X1    g08632(.A1(new_n8824_), .A2(new_n8428_), .Z(new_n8825_));
  INV_X1     g08633(.I(new_n8825_), .ZN(new_n8826_));
  AOI21_X1   g08634(.A1(new_n8482_), .A2(new_n8463_), .B(\asqrt[23] ), .ZN(new_n8827_));
  XOR2_X1    g08635(.A1(new_n8827_), .A2(new_n8473_), .Z(new_n8828_));
  INV_X1     g08636(.I(new_n8828_), .ZN(new_n8829_));
  NAND2_X1   g08637(.A1(\asqrt[24] ), .A2(new_n8451_), .ZN(new_n8830_));
  NOR2_X1    g08638(.A1(new_n8458_), .A2(\a[48] ), .ZN(new_n8831_));
  AOI22_X1   g08639(.A1(new_n8830_), .A2(new_n8458_), .B1(\asqrt[24] ), .B2(new_n8831_), .ZN(new_n8832_));
  OAI21_X1   g08640(.A1(new_n8440_), .A2(new_n8451_), .B(new_n8477_), .ZN(new_n8833_));
  AOI21_X1   g08641(.A1(new_n8476_), .A2(new_n8833_), .B(\asqrt[23] ), .ZN(new_n8834_));
  XOR2_X1    g08642(.A1(new_n8834_), .A2(new_n8832_), .Z(new_n8835_));
  NOR2_X1    g08643(.A1(new_n8758_), .A2(new_n8756_), .ZN(new_n8836_));
  AOI21_X1   g08644(.A1(new_n8762_), .A2(new_n8743_), .B(\asqrt[62] ), .ZN(new_n8837_));
  NOR3_X1    g08645(.A1(new_n8758_), .A2(new_n201_), .A3(new_n8756_), .ZN(new_n8838_));
  OAI22_X1   g08646(.A1(new_n8837_), .A2(new_n8838_), .B1(new_n8836_), .B2(new_n8765_), .ZN(new_n8839_));
  AOI21_X1   g08647(.A1(new_n8839_), .A2(new_n8568_), .B(new_n8769_), .ZN(new_n8840_));
  AOI21_X1   g08648(.A1(new_n8836_), .A2(new_n201_), .B(new_n8766_), .ZN(new_n8841_));
  NOR2_X1    g08649(.A1(new_n8836_), .A2(new_n201_), .ZN(new_n8842_));
  NOR3_X1    g08650(.A1(new_n8841_), .A2(new_n8842_), .A3(new_n8568_), .ZN(new_n8843_));
  NAND3_X1   g08651(.A1(new_n8777_), .A2(\asqrt[24] ), .A3(new_n8779_), .ZN(new_n8844_));
  NOR4_X1    g08652(.A1(new_n8840_), .A2(\asqrt[63] ), .A3(new_n8843_), .A4(new_n8844_), .ZN(new_n8845_));
  INV_X1     g08653(.I(new_n8845_), .ZN(new_n8846_));
  NAND2_X1   g08654(.A1(\asqrt[23] ), .A2(new_n8448_), .ZN(new_n8847_));
  AOI21_X1   g08655(.A1(new_n8847_), .A2(new_n8846_), .B(\a[48] ), .ZN(new_n8848_));
  NOR4_X1    g08656(.A1(new_n8840_), .A2(\asqrt[63] ), .A3(new_n8843_), .A4(new_n8780_), .ZN(new_n8849_));
  NOR2_X1    g08657(.A1(new_n8849_), .A2(new_n8449_), .ZN(new_n8850_));
  NOR3_X1    g08658(.A1(new_n8850_), .A2(new_n8451_), .A3(new_n8845_), .ZN(new_n8851_));
  NOR2_X1    g08659(.A1(new_n8851_), .A2(new_n8848_), .ZN(new_n8852_));
  INV_X1     g08660(.I(\a[46] ), .ZN(new_n8853_));
  NOR2_X1    g08661(.A1(\a[44] ), .A2(\a[45] ), .ZN(new_n8854_));
  NOR3_X1    g08662(.A1(new_n8849_), .A2(new_n8853_), .A3(new_n8854_), .ZN(new_n8855_));
  INV_X1     g08663(.I(new_n8854_), .ZN(new_n8856_));
  AOI21_X1   g08664(.A1(new_n8849_), .A2(\a[46] ), .B(new_n8856_), .ZN(new_n8857_));
  OAI21_X1   g08665(.A1(new_n8855_), .A2(new_n8857_), .B(\asqrt[24] ), .ZN(new_n8858_));
  NAND2_X1   g08666(.A1(new_n8854_), .A2(new_n8853_), .ZN(new_n8859_));
  NAND3_X1   g08667(.A1(new_n8377_), .A2(new_n8379_), .A3(new_n8859_), .ZN(new_n8860_));
  NAND2_X1   g08668(.A1(new_n8443_), .A2(new_n8860_), .ZN(new_n8861_));
  NAND3_X1   g08669(.A1(\asqrt[23] ), .A2(\a[46] ), .A3(new_n8861_), .ZN(new_n8862_));
  NOR3_X1    g08670(.A1(new_n8849_), .A2(\a[46] ), .A3(\a[47] ), .ZN(new_n8863_));
  INV_X1     g08671(.I(\a[47] ), .ZN(new_n8864_));
  AOI21_X1   g08672(.A1(\asqrt[23] ), .A2(new_n8853_), .B(new_n8864_), .ZN(new_n8865_));
  NOR2_X1    g08673(.A1(new_n8863_), .A2(new_n8865_), .ZN(new_n8866_));
  NAND4_X1   g08674(.A1(new_n8858_), .A2(new_n8866_), .A3(new_n8077_), .A4(new_n8862_), .ZN(new_n8867_));
  NAND2_X1   g08675(.A1(new_n8867_), .A2(new_n8852_), .ZN(new_n8868_));
  NAND3_X1   g08676(.A1(\asqrt[23] ), .A2(\a[46] ), .A3(new_n8856_), .ZN(new_n8869_));
  OAI21_X1   g08677(.A1(\asqrt[23] ), .A2(new_n8853_), .B(new_n8854_), .ZN(new_n8870_));
  AOI21_X1   g08678(.A1(new_n8870_), .A2(new_n8869_), .B(new_n8440_), .ZN(new_n8871_));
  NAND3_X1   g08679(.A1(\asqrt[23] ), .A2(new_n8853_), .A3(new_n8864_), .ZN(new_n8872_));
  OAI21_X1   g08680(.A1(new_n8849_), .A2(\a[46] ), .B(\a[47] ), .ZN(new_n8873_));
  NAND3_X1   g08681(.A1(new_n8862_), .A2(new_n8873_), .A3(new_n8872_), .ZN(new_n8874_));
  OAI21_X1   g08682(.A1(new_n8874_), .A2(new_n8871_), .B(\asqrt[25] ), .ZN(new_n8875_));
  NAND3_X1   g08683(.A1(new_n8868_), .A2(new_n7690_), .A3(new_n8875_), .ZN(new_n8876_));
  AOI21_X1   g08684(.A1(new_n8868_), .A2(new_n8875_), .B(new_n7690_), .ZN(new_n8877_));
  AOI21_X1   g08685(.A1(new_n8835_), .A2(new_n8876_), .B(new_n8877_), .ZN(new_n8878_));
  AOI21_X1   g08686(.A1(new_n8878_), .A2(new_n7331_), .B(new_n8829_), .ZN(new_n8879_));
  OR2_X2     g08687(.A1(new_n8851_), .A2(new_n8848_), .Z(new_n8880_));
  NOR3_X1    g08688(.A1(new_n8874_), .A2(new_n8871_), .A3(\asqrt[25] ), .ZN(new_n8881_));
  OAI21_X1   g08689(.A1(new_n8880_), .A2(new_n8881_), .B(new_n8875_), .ZN(new_n8882_));
  OAI21_X1   g08690(.A1(new_n8882_), .A2(\asqrt[26] ), .B(new_n8835_), .ZN(new_n8883_));
  NAND2_X1   g08691(.A1(new_n8882_), .A2(\asqrt[26] ), .ZN(new_n8884_));
  AOI21_X1   g08692(.A1(new_n8883_), .A2(new_n8884_), .B(new_n7331_), .ZN(new_n8885_));
  NOR3_X1    g08693(.A1(new_n8879_), .A2(\asqrt[28] ), .A3(new_n8885_), .ZN(new_n8886_));
  OAI21_X1   g08694(.A1(new_n8879_), .A2(new_n8885_), .B(\asqrt[28] ), .ZN(new_n8887_));
  OAI21_X1   g08695(.A1(new_n8826_), .A2(new_n8886_), .B(new_n8887_), .ZN(new_n8888_));
  OAI21_X1   g08696(.A1(new_n8888_), .A2(\asqrt[29] ), .B(new_n8822_), .ZN(new_n8889_));
  NAND3_X1   g08697(.A1(new_n8883_), .A2(new_n8884_), .A3(new_n7331_), .ZN(new_n8890_));
  AOI21_X1   g08698(.A1(new_n8828_), .A2(new_n8890_), .B(new_n8885_), .ZN(new_n8891_));
  AOI21_X1   g08699(.A1(new_n8891_), .A2(new_n6966_), .B(new_n8826_), .ZN(new_n8892_));
  NAND2_X1   g08700(.A1(new_n8890_), .A2(new_n8828_), .ZN(new_n8893_));
  INV_X1     g08701(.I(new_n8885_), .ZN(new_n8894_));
  AOI21_X1   g08702(.A1(new_n8893_), .A2(new_n8894_), .B(new_n6966_), .ZN(new_n8895_));
  OAI21_X1   g08703(.A1(new_n8892_), .A2(new_n8895_), .B(\asqrt[29] ), .ZN(new_n8896_));
  NAND3_X1   g08704(.A1(new_n8889_), .A2(new_n6275_), .A3(new_n8896_), .ZN(new_n8897_));
  AOI21_X1   g08705(.A1(new_n8889_), .A2(new_n8896_), .B(new_n6275_), .ZN(new_n8898_));
  AOI21_X1   g08706(.A1(new_n8820_), .A2(new_n8897_), .B(new_n8898_), .ZN(new_n8899_));
  AOI21_X1   g08707(.A1(new_n8899_), .A2(new_n5947_), .B(new_n8817_), .ZN(new_n8900_));
  INV_X1     g08708(.I(new_n8822_), .ZN(new_n8901_));
  NOR3_X1    g08709(.A1(new_n8892_), .A2(\asqrt[29] ), .A3(new_n8895_), .ZN(new_n8902_));
  OAI21_X1   g08710(.A1(new_n8901_), .A2(new_n8902_), .B(new_n8896_), .ZN(new_n8903_));
  OAI21_X1   g08711(.A1(new_n8903_), .A2(\asqrt[30] ), .B(new_n8820_), .ZN(new_n8904_));
  NAND2_X1   g08712(.A1(new_n8903_), .A2(\asqrt[30] ), .ZN(new_n8905_));
  AOI21_X1   g08713(.A1(new_n8904_), .A2(new_n8905_), .B(new_n5947_), .ZN(new_n8906_));
  NOR3_X1    g08714(.A1(new_n8900_), .A2(\asqrt[32] ), .A3(new_n8906_), .ZN(new_n8907_));
  OAI21_X1   g08715(.A1(new_n8900_), .A2(new_n8906_), .B(\asqrt[32] ), .ZN(new_n8908_));
  OAI21_X1   g08716(.A1(new_n8814_), .A2(new_n8907_), .B(new_n8908_), .ZN(new_n8909_));
  OAI21_X1   g08717(.A1(new_n8909_), .A2(\asqrt[33] ), .B(new_n8810_), .ZN(new_n8910_));
  NAND3_X1   g08718(.A1(new_n8904_), .A2(new_n8905_), .A3(new_n5947_), .ZN(new_n8911_));
  AOI21_X1   g08719(.A1(new_n8816_), .A2(new_n8911_), .B(new_n8906_), .ZN(new_n8912_));
  AOI21_X1   g08720(.A1(new_n8912_), .A2(new_n5643_), .B(new_n8814_), .ZN(new_n8913_));
  NAND2_X1   g08721(.A1(new_n8911_), .A2(new_n8816_), .ZN(new_n8914_));
  INV_X1     g08722(.I(new_n8906_), .ZN(new_n8915_));
  AOI21_X1   g08723(.A1(new_n8914_), .A2(new_n8915_), .B(new_n5643_), .ZN(new_n8916_));
  OAI21_X1   g08724(.A1(new_n8913_), .A2(new_n8916_), .B(\asqrt[33] ), .ZN(new_n8917_));
  NAND3_X1   g08725(.A1(new_n8910_), .A2(new_n5029_), .A3(new_n8917_), .ZN(new_n8918_));
  AOI21_X1   g08726(.A1(new_n8910_), .A2(new_n8917_), .B(new_n5029_), .ZN(new_n8919_));
  AOI21_X1   g08727(.A1(new_n8808_), .A2(new_n8918_), .B(new_n8919_), .ZN(new_n8920_));
  AOI21_X1   g08728(.A1(new_n8920_), .A2(new_n4751_), .B(new_n8805_), .ZN(new_n8921_));
  INV_X1     g08729(.I(new_n8810_), .ZN(new_n8922_));
  NOR3_X1    g08730(.A1(new_n8913_), .A2(\asqrt[33] ), .A3(new_n8916_), .ZN(new_n8923_));
  OAI21_X1   g08731(.A1(new_n8922_), .A2(new_n8923_), .B(new_n8917_), .ZN(new_n8924_));
  OAI21_X1   g08732(.A1(new_n8924_), .A2(\asqrt[34] ), .B(new_n8808_), .ZN(new_n8925_));
  NAND2_X1   g08733(.A1(new_n8924_), .A2(\asqrt[34] ), .ZN(new_n8926_));
  AOI21_X1   g08734(.A1(new_n8925_), .A2(new_n8926_), .B(new_n4751_), .ZN(new_n8927_));
  NOR3_X1    g08735(.A1(new_n8921_), .A2(\asqrt[36] ), .A3(new_n8927_), .ZN(new_n8928_));
  OAI21_X1   g08736(.A1(new_n8921_), .A2(new_n8927_), .B(\asqrt[36] ), .ZN(new_n8929_));
  OAI21_X1   g08737(.A1(new_n8802_), .A2(new_n8928_), .B(new_n8929_), .ZN(new_n8930_));
  OAI21_X1   g08738(.A1(new_n8930_), .A2(\asqrt[37] ), .B(new_n8798_), .ZN(new_n8931_));
  NAND3_X1   g08739(.A1(new_n8925_), .A2(new_n8926_), .A3(new_n4751_), .ZN(new_n8932_));
  AOI21_X1   g08740(.A1(new_n8804_), .A2(new_n8932_), .B(new_n8927_), .ZN(new_n8933_));
  AOI21_X1   g08741(.A1(new_n8933_), .A2(new_n4461_), .B(new_n8802_), .ZN(new_n8934_));
  NAND2_X1   g08742(.A1(new_n8932_), .A2(new_n8804_), .ZN(new_n8935_));
  INV_X1     g08743(.I(new_n8927_), .ZN(new_n8936_));
  AOI21_X1   g08744(.A1(new_n8935_), .A2(new_n8936_), .B(new_n4461_), .ZN(new_n8937_));
  OAI21_X1   g08745(.A1(new_n8934_), .A2(new_n8937_), .B(\asqrt[37] ), .ZN(new_n8938_));
  NAND3_X1   g08746(.A1(new_n8931_), .A2(new_n3925_), .A3(new_n8938_), .ZN(new_n8939_));
  AOI21_X1   g08747(.A1(new_n8931_), .A2(new_n8938_), .B(new_n3925_), .ZN(new_n8940_));
  AOI21_X1   g08748(.A1(new_n8796_), .A2(new_n8939_), .B(new_n8940_), .ZN(new_n8941_));
  AOI21_X1   g08749(.A1(new_n8941_), .A2(new_n3681_), .B(new_n8793_), .ZN(new_n8942_));
  INV_X1     g08750(.I(new_n8798_), .ZN(new_n8943_));
  NOR3_X1    g08751(.A1(new_n8934_), .A2(\asqrt[37] ), .A3(new_n8937_), .ZN(new_n8944_));
  OAI21_X1   g08752(.A1(new_n8943_), .A2(new_n8944_), .B(new_n8938_), .ZN(new_n8945_));
  OAI21_X1   g08753(.A1(new_n8945_), .A2(\asqrt[38] ), .B(new_n8796_), .ZN(new_n8946_));
  NAND2_X1   g08754(.A1(new_n8945_), .A2(\asqrt[38] ), .ZN(new_n8947_));
  AOI21_X1   g08755(.A1(new_n8946_), .A2(new_n8947_), .B(new_n3681_), .ZN(new_n8948_));
  NOR3_X1    g08756(.A1(new_n8942_), .A2(\asqrt[40] ), .A3(new_n8948_), .ZN(new_n8949_));
  OAI21_X1   g08757(.A1(new_n8942_), .A2(new_n8948_), .B(\asqrt[40] ), .ZN(new_n8950_));
  OAI21_X1   g08758(.A1(new_n8790_), .A2(new_n8949_), .B(new_n8950_), .ZN(new_n8951_));
  OAI21_X1   g08759(.A1(new_n8951_), .A2(\asqrt[41] ), .B(new_n8786_), .ZN(new_n8952_));
  NAND3_X1   g08760(.A1(new_n8946_), .A2(new_n8947_), .A3(new_n3681_), .ZN(new_n8953_));
  AOI21_X1   g08761(.A1(new_n8792_), .A2(new_n8953_), .B(new_n8948_), .ZN(new_n8954_));
  AOI21_X1   g08762(.A1(new_n8954_), .A2(new_n3427_), .B(new_n8790_), .ZN(new_n8955_));
  NAND2_X1   g08763(.A1(new_n8953_), .A2(new_n8792_), .ZN(new_n8956_));
  INV_X1     g08764(.I(new_n8948_), .ZN(new_n8957_));
  AOI21_X1   g08765(.A1(new_n8956_), .A2(new_n8957_), .B(new_n3427_), .ZN(new_n8958_));
  OAI21_X1   g08766(.A1(new_n8955_), .A2(new_n8958_), .B(\asqrt[41] ), .ZN(new_n8959_));
  NAND3_X1   g08767(.A1(new_n8952_), .A2(new_n2960_), .A3(new_n8959_), .ZN(new_n8960_));
  INV_X1     g08768(.I(new_n8786_), .ZN(new_n8961_));
  NOR3_X1    g08769(.A1(new_n8955_), .A2(\asqrt[41] ), .A3(new_n8958_), .ZN(new_n8962_));
  OAI21_X1   g08770(.A1(new_n8961_), .A2(new_n8962_), .B(new_n8959_), .ZN(new_n8963_));
  NAND2_X1   g08771(.A1(new_n8963_), .A2(\asqrt[42] ), .ZN(new_n8964_));
  NOR2_X1    g08772(.A1(new_n8748_), .A2(\asqrt[62] ), .ZN(new_n8965_));
  NOR2_X1    g08773(.A1(new_n8965_), .A2(new_n8842_), .ZN(new_n8966_));
  XOR2_X1    g08774(.A1(new_n8764_), .A2(new_n8350_), .Z(new_n8967_));
  OAI21_X1   g08775(.A1(\asqrt[23] ), .A2(new_n8966_), .B(new_n8967_), .ZN(new_n8968_));
  INV_X1     g08776(.I(new_n8968_), .ZN(new_n8969_));
  AOI21_X1   g08777(.A1(new_n8733_), .A2(new_n8741_), .B(\asqrt[23] ), .ZN(new_n8970_));
  XOR2_X1    g08778(.A1(new_n8970_), .A2(new_n8576_), .Z(new_n8971_));
  INV_X1     g08779(.I(new_n8971_), .ZN(new_n8972_));
  AOI21_X1   g08780(.A1(new_n8724_), .A2(new_n8732_), .B(\asqrt[23] ), .ZN(new_n8973_));
  XOR2_X1    g08781(.A1(new_n8973_), .A2(new_n8578_), .Z(new_n8974_));
  INV_X1     g08782(.I(new_n8974_), .ZN(new_n8975_));
  NAND2_X1   g08783(.A1(new_n8728_), .A2(new_n531_), .ZN(new_n8976_));
  AOI21_X1   g08784(.A1(new_n8976_), .A2(new_n8723_), .B(\asqrt[23] ), .ZN(new_n8977_));
  XOR2_X1    g08785(.A1(new_n8977_), .A2(new_n8580_), .Z(new_n8978_));
  AOI21_X1   g08786(.A1(new_n8727_), .A2(new_n8713_), .B(\asqrt[23] ), .ZN(new_n8979_));
  XOR2_X1    g08787(.A1(new_n8979_), .A2(new_n8584_), .Z(new_n8980_));
  NAND2_X1   g08788(.A1(new_n8695_), .A2(new_n744_), .ZN(new_n8981_));
  AOI21_X1   g08789(.A1(new_n8981_), .A2(new_n8721_), .B(\asqrt[23] ), .ZN(new_n8982_));
  XOR2_X1    g08790(.A1(new_n8982_), .A2(new_n8588_), .Z(new_n8983_));
  INV_X1     g08791(.I(new_n8983_), .ZN(new_n8984_));
  AOI21_X1   g08792(.A1(new_n8693_), .A2(new_n8710_), .B(\asqrt[23] ), .ZN(new_n8985_));
  XOR2_X1    g08793(.A1(new_n8985_), .A2(new_n8591_), .Z(new_n8986_));
  INV_X1     g08794(.I(new_n8986_), .ZN(new_n8987_));
  NAND2_X1   g08795(.A1(new_n8706_), .A2(new_n1006_), .ZN(new_n8988_));
  AOI21_X1   g08796(.A1(new_n8988_), .A2(new_n8692_), .B(\asqrt[23] ), .ZN(new_n8989_));
  XOR2_X1    g08797(.A1(new_n8989_), .A2(new_n8593_), .Z(new_n8990_));
  AOI21_X1   g08798(.A1(new_n8704_), .A2(new_n8689_), .B(\asqrt[23] ), .ZN(new_n8991_));
  XOR2_X1    g08799(.A1(new_n8991_), .A2(new_n8596_), .Z(new_n8992_));
  NAND2_X1   g08800(.A1(new_n8671_), .A2(new_n1305_), .ZN(new_n8993_));
  AOI21_X1   g08801(.A1(new_n8993_), .A2(new_n8703_), .B(\asqrt[23] ), .ZN(new_n8994_));
  XOR2_X1    g08802(.A1(new_n8994_), .A2(new_n8600_), .Z(new_n8995_));
  INV_X1     g08803(.I(new_n8995_), .ZN(new_n8996_));
  AOI21_X1   g08804(.A1(new_n8669_), .A2(new_n8686_), .B(\asqrt[23] ), .ZN(new_n8997_));
  XOR2_X1    g08805(.A1(new_n8997_), .A2(new_n8603_), .Z(new_n8998_));
  INV_X1     g08806(.I(new_n8998_), .ZN(new_n8999_));
  NAND2_X1   g08807(.A1(new_n8682_), .A2(new_n1632_), .ZN(new_n9000_));
  AOI21_X1   g08808(.A1(new_n9000_), .A2(new_n8668_), .B(\asqrt[23] ), .ZN(new_n9001_));
  XOR2_X1    g08809(.A1(new_n9001_), .A2(new_n8605_), .Z(new_n9002_));
  AOI21_X1   g08810(.A1(new_n8680_), .A2(new_n8665_), .B(\asqrt[23] ), .ZN(new_n9003_));
  XOR2_X1    g08811(.A1(new_n9003_), .A2(new_n8608_), .Z(new_n9004_));
  NAND2_X1   g08812(.A1(new_n8647_), .A2(new_n1953_), .ZN(new_n9005_));
  AOI21_X1   g08813(.A1(new_n9005_), .A2(new_n8679_), .B(\asqrt[23] ), .ZN(new_n9006_));
  XOR2_X1    g08814(.A1(new_n9006_), .A2(new_n8612_), .Z(new_n9007_));
  INV_X1     g08815(.I(new_n9007_), .ZN(new_n9008_));
  AOI21_X1   g08816(.A1(new_n8645_), .A2(new_n8662_), .B(\asqrt[23] ), .ZN(new_n9009_));
  XOR2_X1    g08817(.A1(new_n9009_), .A2(new_n8615_), .Z(new_n9010_));
  INV_X1     g08818(.I(new_n9010_), .ZN(new_n9011_));
  NAND2_X1   g08819(.A1(new_n8658_), .A2(new_n2332_), .ZN(new_n9012_));
  AOI21_X1   g08820(.A1(new_n9012_), .A2(new_n8644_), .B(\asqrt[23] ), .ZN(new_n9013_));
  XOR2_X1    g08821(.A1(new_n9013_), .A2(new_n8617_), .Z(new_n9014_));
  AOI21_X1   g08822(.A1(new_n8656_), .A2(new_n8641_), .B(\asqrt[23] ), .ZN(new_n9015_));
  XOR2_X1    g08823(.A1(new_n9015_), .A2(new_n8620_), .Z(new_n9016_));
  NAND2_X1   g08824(.A1(new_n8631_), .A2(new_n2749_), .ZN(new_n9017_));
  AOI21_X1   g08825(.A1(new_n9017_), .A2(new_n8655_), .B(\asqrt[23] ), .ZN(new_n9018_));
  XOR2_X1    g08826(.A1(new_n9018_), .A2(new_n8624_), .Z(new_n9019_));
  INV_X1     g08827(.I(new_n9019_), .ZN(new_n9020_));
  AOI21_X1   g08828(.A1(new_n8629_), .A2(new_n8638_), .B(\asqrt[23] ), .ZN(new_n9021_));
  XOR2_X1    g08829(.A1(new_n9021_), .A2(new_n8627_), .Z(new_n9022_));
  INV_X1     g08830(.I(new_n9022_), .ZN(new_n9023_));
  AOI21_X1   g08831(.A1(new_n8952_), .A2(new_n8959_), .B(new_n2960_), .ZN(new_n9024_));
  AOI21_X1   g08832(.A1(new_n8784_), .A2(new_n8960_), .B(new_n9024_), .ZN(new_n9025_));
  AOI21_X1   g08833(.A1(new_n9025_), .A2(new_n2749_), .B(new_n9023_), .ZN(new_n9026_));
  OAI21_X1   g08834(.A1(new_n8963_), .A2(\asqrt[42] ), .B(new_n8784_), .ZN(new_n9027_));
  AOI21_X1   g08835(.A1(new_n9027_), .A2(new_n8964_), .B(new_n2749_), .ZN(new_n9028_));
  NOR3_X1    g08836(.A1(new_n9026_), .A2(\asqrt[44] ), .A3(new_n9028_), .ZN(new_n9029_));
  OAI21_X1   g08837(.A1(new_n9026_), .A2(new_n9028_), .B(\asqrt[44] ), .ZN(new_n9030_));
  OAI21_X1   g08838(.A1(new_n9020_), .A2(new_n9029_), .B(new_n9030_), .ZN(new_n9031_));
  OAI21_X1   g08839(.A1(new_n9031_), .A2(\asqrt[45] ), .B(new_n9016_), .ZN(new_n9032_));
  NAND3_X1   g08840(.A1(new_n9027_), .A2(new_n8964_), .A3(new_n2749_), .ZN(new_n9033_));
  AOI21_X1   g08841(.A1(new_n9022_), .A2(new_n9033_), .B(new_n9028_), .ZN(new_n9034_));
  AOI21_X1   g08842(.A1(new_n9034_), .A2(new_n2531_), .B(new_n9020_), .ZN(new_n9035_));
  NAND2_X1   g08843(.A1(new_n9033_), .A2(new_n9022_), .ZN(new_n9036_));
  INV_X1     g08844(.I(new_n9028_), .ZN(new_n9037_));
  AOI21_X1   g08845(.A1(new_n9036_), .A2(new_n9037_), .B(new_n2531_), .ZN(new_n9038_));
  OAI21_X1   g08846(.A1(new_n9035_), .A2(new_n9038_), .B(\asqrt[45] ), .ZN(new_n9039_));
  NAND3_X1   g08847(.A1(new_n9032_), .A2(new_n2134_), .A3(new_n9039_), .ZN(new_n9040_));
  AOI21_X1   g08848(.A1(new_n9032_), .A2(new_n9039_), .B(new_n2134_), .ZN(new_n9041_));
  AOI21_X1   g08849(.A1(new_n9014_), .A2(new_n9040_), .B(new_n9041_), .ZN(new_n9042_));
  AOI21_X1   g08850(.A1(new_n9042_), .A2(new_n1953_), .B(new_n9011_), .ZN(new_n9043_));
  INV_X1     g08851(.I(new_n9016_), .ZN(new_n9044_));
  NOR3_X1    g08852(.A1(new_n9035_), .A2(\asqrt[45] ), .A3(new_n9038_), .ZN(new_n9045_));
  OAI21_X1   g08853(.A1(new_n9044_), .A2(new_n9045_), .B(new_n9039_), .ZN(new_n9046_));
  OAI21_X1   g08854(.A1(new_n9046_), .A2(\asqrt[46] ), .B(new_n9014_), .ZN(new_n9047_));
  NAND2_X1   g08855(.A1(new_n9046_), .A2(\asqrt[46] ), .ZN(new_n9048_));
  AOI21_X1   g08856(.A1(new_n9047_), .A2(new_n9048_), .B(new_n1953_), .ZN(new_n9049_));
  NOR3_X1    g08857(.A1(new_n9043_), .A2(\asqrt[48] ), .A3(new_n9049_), .ZN(new_n9050_));
  OAI21_X1   g08858(.A1(new_n9043_), .A2(new_n9049_), .B(\asqrt[48] ), .ZN(new_n9051_));
  OAI21_X1   g08859(.A1(new_n9008_), .A2(new_n9050_), .B(new_n9051_), .ZN(new_n9052_));
  OAI21_X1   g08860(.A1(new_n9052_), .A2(\asqrt[49] ), .B(new_n9004_), .ZN(new_n9053_));
  NAND3_X1   g08861(.A1(new_n9047_), .A2(new_n9048_), .A3(new_n1953_), .ZN(new_n9054_));
  AOI21_X1   g08862(.A1(new_n9010_), .A2(new_n9054_), .B(new_n9049_), .ZN(new_n9055_));
  AOI21_X1   g08863(.A1(new_n9055_), .A2(new_n1778_), .B(new_n9008_), .ZN(new_n9056_));
  NAND2_X1   g08864(.A1(new_n9054_), .A2(new_n9010_), .ZN(new_n9057_));
  INV_X1     g08865(.I(new_n9049_), .ZN(new_n9058_));
  AOI21_X1   g08866(.A1(new_n9057_), .A2(new_n9058_), .B(new_n1778_), .ZN(new_n9059_));
  OAI21_X1   g08867(.A1(new_n9056_), .A2(new_n9059_), .B(\asqrt[49] ), .ZN(new_n9060_));
  NAND3_X1   g08868(.A1(new_n9053_), .A2(new_n1463_), .A3(new_n9060_), .ZN(new_n9061_));
  AOI21_X1   g08869(.A1(new_n9053_), .A2(new_n9060_), .B(new_n1463_), .ZN(new_n9062_));
  AOI21_X1   g08870(.A1(new_n9002_), .A2(new_n9061_), .B(new_n9062_), .ZN(new_n9063_));
  AOI21_X1   g08871(.A1(new_n9063_), .A2(new_n1305_), .B(new_n8999_), .ZN(new_n9064_));
  INV_X1     g08872(.I(new_n9004_), .ZN(new_n9065_));
  NOR3_X1    g08873(.A1(new_n9056_), .A2(\asqrt[49] ), .A3(new_n9059_), .ZN(new_n9066_));
  OAI21_X1   g08874(.A1(new_n9065_), .A2(new_n9066_), .B(new_n9060_), .ZN(new_n9067_));
  OAI21_X1   g08875(.A1(new_n9067_), .A2(\asqrt[50] ), .B(new_n9002_), .ZN(new_n9068_));
  NAND2_X1   g08876(.A1(new_n9067_), .A2(\asqrt[50] ), .ZN(new_n9069_));
  AOI21_X1   g08877(.A1(new_n9068_), .A2(new_n9069_), .B(new_n1305_), .ZN(new_n9070_));
  NOR3_X1    g08878(.A1(new_n9064_), .A2(\asqrt[52] ), .A3(new_n9070_), .ZN(new_n9071_));
  OAI21_X1   g08879(.A1(new_n9064_), .A2(new_n9070_), .B(\asqrt[52] ), .ZN(new_n9072_));
  OAI21_X1   g08880(.A1(new_n8996_), .A2(new_n9071_), .B(new_n9072_), .ZN(new_n9073_));
  OAI21_X1   g08881(.A1(new_n9073_), .A2(\asqrt[53] ), .B(new_n8992_), .ZN(new_n9074_));
  NAND3_X1   g08882(.A1(new_n9068_), .A2(new_n9069_), .A3(new_n1305_), .ZN(new_n9075_));
  AOI21_X1   g08883(.A1(new_n8998_), .A2(new_n9075_), .B(new_n9070_), .ZN(new_n9076_));
  AOI21_X1   g08884(.A1(new_n9076_), .A2(new_n1150_), .B(new_n8996_), .ZN(new_n9077_));
  NAND2_X1   g08885(.A1(new_n9075_), .A2(new_n8998_), .ZN(new_n9078_));
  INV_X1     g08886(.I(new_n9070_), .ZN(new_n9079_));
  AOI21_X1   g08887(.A1(new_n9078_), .A2(new_n9079_), .B(new_n1150_), .ZN(new_n9080_));
  OAI21_X1   g08888(.A1(new_n9077_), .A2(new_n9080_), .B(\asqrt[53] ), .ZN(new_n9081_));
  NAND3_X1   g08889(.A1(new_n9074_), .A2(new_n860_), .A3(new_n9081_), .ZN(new_n9082_));
  AOI21_X1   g08890(.A1(new_n9074_), .A2(new_n9081_), .B(new_n860_), .ZN(new_n9083_));
  AOI21_X1   g08891(.A1(new_n8990_), .A2(new_n9082_), .B(new_n9083_), .ZN(new_n9084_));
  AOI21_X1   g08892(.A1(new_n9084_), .A2(new_n744_), .B(new_n8987_), .ZN(new_n9085_));
  INV_X1     g08893(.I(new_n8992_), .ZN(new_n9086_));
  NOR3_X1    g08894(.A1(new_n9077_), .A2(\asqrt[53] ), .A3(new_n9080_), .ZN(new_n9087_));
  OAI21_X1   g08895(.A1(new_n9086_), .A2(new_n9087_), .B(new_n9081_), .ZN(new_n9088_));
  OAI21_X1   g08896(.A1(new_n9088_), .A2(\asqrt[54] ), .B(new_n8990_), .ZN(new_n9089_));
  NAND2_X1   g08897(.A1(new_n9088_), .A2(\asqrt[54] ), .ZN(new_n9090_));
  AOI21_X1   g08898(.A1(new_n9089_), .A2(new_n9090_), .B(new_n744_), .ZN(new_n9091_));
  NOR3_X1    g08899(.A1(new_n9085_), .A2(\asqrt[56] ), .A3(new_n9091_), .ZN(new_n9092_));
  OAI21_X1   g08900(.A1(new_n9085_), .A2(new_n9091_), .B(\asqrt[56] ), .ZN(new_n9093_));
  OAI21_X1   g08901(.A1(new_n8984_), .A2(new_n9092_), .B(new_n9093_), .ZN(new_n9094_));
  OAI21_X1   g08902(.A1(new_n9094_), .A2(\asqrt[57] ), .B(new_n8980_), .ZN(new_n9095_));
  NAND3_X1   g08903(.A1(new_n9089_), .A2(new_n9090_), .A3(new_n744_), .ZN(new_n9096_));
  AOI21_X1   g08904(.A1(new_n8986_), .A2(new_n9096_), .B(new_n9091_), .ZN(new_n9097_));
  AOI21_X1   g08905(.A1(new_n9097_), .A2(new_n634_), .B(new_n8984_), .ZN(new_n9098_));
  NAND2_X1   g08906(.A1(new_n9096_), .A2(new_n8986_), .ZN(new_n9099_));
  INV_X1     g08907(.I(new_n9091_), .ZN(new_n9100_));
  AOI21_X1   g08908(.A1(new_n9099_), .A2(new_n9100_), .B(new_n634_), .ZN(new_n9101_));
  OAI21_X1   g08909(.A1(new_n9098_), .A2(new_n9101_), .B(\asqrt[57] ), .ZN(new_n9102_));
  NAND3_X1   g08910(.A1(new_n9095_), .A2(new_n423_), .A3(new_n9102_), .ZN(new_n9103_));
  AOI21_X1   g08911(.A1(new_n9095_), .A2(new_n9102_), .B(new_n423_), .ZN(new_n9104_));
  AOI21_X1   g08912(.A1(new_n8978_), .A2(new_n9103_), .B(new_n9104_), .ZN(new_n9105_));
  AOI21_X1   g08913(.A1(new_n9105_), .A2(new_n337_), .B(new_n8975_), .ZN(new_n9106_));
  NOR2_X1    g08914(.A1(new_n9105_), .A2(new_n337_), .ZN(new_n9107_));
  NOR3_X1    g08915(.A1(new_n9106_), .A2(new_n9107_), .A3(\asqrt[60] ), .ZN(new_n9108_));
  OAI21_X1   g08916(.A1(new_n9106_), .A2(new_n9107_), .B(\asqrt[60] ), .ZN(new_n9109_));
  OAI21_X1   g08917(.A1(new_n8972_), .A2(new_n9108_), .B(new_n9109_), .ZN(new_n9110_));
  NAND2_X1   g08918(.A1(new_n9110_), .A2(\asqrt[61] ), .ZN(new_n9111_));
  AOI21_X1   g08919(.A1(new_n8749_), .A2(new_n8755_), .B(\asqrt[23] ), .ZN(new_n9112_));
  XOR2_X1    g08920(.A1(new_n9112_), .A2(new_n8572_), .Z(new_n9113_));
  OAI21_X1   g08921(.A1(new_n9110_), .A2(\asqrt[61] ), .B(new_n9113_), .ZN(new_n9114_));
  NAND2_X1   g08922(.A1(new_n9114_), .A2(new_n9111_), .ZN(new_n9115_));
  INV_X1     g08923(.I(new_n8980_), .ZN(new_n9116_));
  NOR3_X1    g08924(.A1(new_n9098_), .A2(\asqrt[57] ), .A3(new_n9101_), .ZN(new_n9117_));
  OAI21_X1   g08925(.A1(new_n9116_), .A2(new_n9117_), .B(new_n9102_), .ZN(new_n9118_));
  OAI21_X1   g08926(.A1(new_n9118_), .A2(\asqrt[58] ), .B(new_n8978_), .ZN(new_n9119_));
  NOR2_X1    g08927(.A1(new_n9117_), .A2(new_n9116_), .ZN(new_n9120_));
  INV_X1     g08928(.I(new_n9102_), .ZN(new_n9121_));
  OAI21_X1   g08929(.A1(new_n9120_), .A2(new_n9121_), .B(\asqrt[58] ), .ZN(new_n9122_));
  NAND3_X1   g08930(.A1(new_n9119_), .A2(new_n337_), .A3(new_n9122_), .ZN(new_n9123_));
  NAND2_X1   g08931(.A1(new_n9123_), .A2(new_n8974_), .ZN(new_n9124_));
  INV_X1     g08932(.I(new_n8978_), .ZN(new_n9125_));
  NOR2_X1    g08933(.A1(new_n9120_), .A2(new_n9121_), .ZN(new_n9126_));
  AOI21_X1   g08934(.A1(new_n9126_), .A2(new_n423_), .B(new_n9125_), .ZN(new_n9127_));
  OAI21_X1   g08935(.A1(new_n9127_), .A2(new_n9104_), .B(\asqrt[59] ), .ZN(new_n9128_));
  NAND3_X1   g08936(.A1(new_n9124_), .A2(new_n266_), .A3(new_n9128_), .ZN(new_n9129_));
  NAND2_X1   g08937(.A1(new_n9129_), .A2(new_n8971_), .ZN(new_n9130_));
  AOI21_X1   g08938(.A1(new_n9130_), .A2(new_n9109_), .B(new_n239_), .ZN(new_n9131_));
  AOI21_X1   g08939(.A1(new_n9124_), .A2(new_n9128_), .B(new_n266_), .ZN(new_n9132_));
  AOI21_X1   g08940(.A1(new_n8971_), .A2(new_n9129_), .B(new_n9132_), .ZN(new_n9133_));
  INV_X1     g08941(.I(new_n9113_), .ZN(new_n9134_));
  AOI21_X1   g08942(.A1(new_n9133_), .A2(new_n239_), .B(new_n9134_), .ZN(new_n9135_));
  OAI21_X1   g08943(.A1(new_n9135_), .A2(new_n9131_), .B(new_n201_), .ZN(new_n9136_));
  NAND3_X1   g08944(.A1(new_n9114_), .A2(new_n9111_), .A3(\asqrt[62] ), .ZN(new_n9137_));
  NOR2_X1    g08945(.A1(new_n8747_), .A2(new_n8756_), .ZN(new_n9138_));
  NOR2_X1    g08946(.A1(\asqrt[23] ), .A2(new_n9138_), .ZN(new_n9139_));
  XOR2_X1    g08947(.A1(new_n9139_), .A2(new_n8745_), .Z(new_n9140_));
  INV_X1     g08948(.I(new_n9140_), .ZN(new_n9141_));
  AOI22_X1   g08949(.A1(new_n9137_), .A2(new_n9136_), .B1(new_n9115_), .B2(new_n9141_), .ZN(new_n9142_));
  NOR2_X1    g08950(.A1(new_n8767_), .A2(new_n8569_), .ZN(new_n9143_));
  OAI21_X1   g08951(.A1(\asqrt[23] ), .A2(new_n9143_), .B(new_n8774_), .ZN(new_n9144_));
  INV_X1     g08952(.I(new_n9144_), .ZN(new_n9145_));
  OAI21_X1   g08953(.A1(new_n9142_), .A2(new_n8969_), .B(new_n9145_), .ZN(new_n9146_));
  OAI21_X1   g08954(.A1(new_n9115_), .A2(\asqrt[62] ), .B(new_n9140_), .ZN(new_n9147_));
  NAND2_X1   g08955(.A1(new_n9115_), .A2(\asqrt[62] ), .ZN(new_n9148_));
  NAND3_X1   g08956(.A1(new_n9147_), .A2(new_n9148_), .A3(new_n8969_), .ZN(new_n9149_));
  NAND2_X1   g08957(.A1(new_n8767_), .A2(new_n8568_), .ZN(new_n9150_));
  NAND2_X1   g08958(.A1(new_n8839_), .A2(new_n8569_), .ZN(new_n9151_));
  AOI21_X1   g08959(.A1(new_n9150_), .A2(new_n9151_), .B(new_n193_), .ZN(new_n9152_));
  OAI21_X1   g08960(.A1(\asqrt[23] ), .A2(new_n8569_), .B(new_n9152_), .ZN(new_n9153_));
  NOR2_X1    g08961(.A1(new_n8780_), .A2(new_n8568_), .ZN(new_n9154_));
  NAND4_X1   g08962(.A1(new_n8771_), .A2(new_n193_), .A3(new_n8774_), .A4(new_n9154_), .ZN(new_n9155_));
  NAND2_X1   g08963(.A1(new_n9153_), .A2(new_n9155_), .ZN(new_n9156_));
  INV_X1     g08964(.I(new_n9156_), .ZN(new_n9157_));
  NAND4_X1   g08965(.A1(new_n9146_), .A2(new_n193_), .A3(new_n9149_), .A4(new_n9157_), .ZN(\asqrt[22] ));
  AOI21_X1   g08966(.A1(new_n8960_), .A2(new_n8964_), .B(\asqrt[22] ), .ZN(new_n9159_));
  XOR2_X1    g08967(.A1(new_n9159_), .A2(new_n8784_), .Z(new_n9160_));
  XOR2_X1    g08968(.A1(new_n8951_), .A2(\asqrt[41] ), .Z(new_n9161_));
  NOR2_X1    g08969(.A1(\asqrt[22] ), .A2(new_n9161_), .ZN(new_n9162_));
  XOR2_X1    g08970(.A1(new_n9162_), .A2(new_n8786_), .Z(new_n9163_));
  NOR2_X1    g08971(.A1(new_n8949_), .A2(new_n8958_), .ZN(new_n9164_));
  NOR2_X1    g08972(.A1(\asqrt[22] ), .A2(new_n9164_), .ZN(new_n9165_));
  XOR2_X1    g08973(.A1(new_n9165_), .A2(new_n8789_), .Z(new_n9166_));
  AOI21_X1   g08974(.A1(new_n8953_), .A2(new_n8957_), .B(\asqrt[22] ), .ZN(new_n9167_));
  XOR2_X1    g08975(.A1(new_n9167_), .A2(new_n8792_), .Z(new_n9168_));
  INV_X1     g08976(.I(new_n9168_), .ZN(new_n9169_));
  AOI21_X1   g08977(.A1(new_n8939_), .A2(new_n8947_), .B(\asqrt[22] ), .ZN(new_n9170_));
  XOR2_X1    g08978(.A1(new_n9170_), .A2(new_n8796_), .Z(new_n9171_));
  INV_X1     g08979(.I(new_n9171_), .ZN(new_n9172_));
  XOR2_X1    g08980(.A1(new_n8930_), .A2(\asqrt[37] ), .Z(new_n9173_));
  NOR2_X1    g08981(.A1(\asqrt[22] ), .A2(new_n9173_), .ZN(new_n9174_));
  XOR2_X1    g08982(.A1(new_n9174_), .A2(new_n8798_), .Z(new_n9175_));
  NOR2_X1    g08983(.A1(new_n8928_), .A2(new_n8937_), .ZN(new_n9176_));
  NOR2_X1    g08984(.A1(\asqrt[22] ), .A2(new_n9176_), .ZN(new_n9177_));
  XOR2_X1    g08985(.A1(new_n9177_), .A2(new_n8801_), .Z(new_n9178_));
  AOI21_X1   g08986(.A1(new_n8932_), .A2(new_n8936_), .B(\asqrt[22] ), .ZN(new_n9179_));
  XOR2_X1    g08987(.A1(new_n9179_), .A2(new_n8804_), .Z(new_n9180_));
  INV_X1     g08988(.I(new_n9180_), .ZN(new_n9181_));
  AOI21_X1   g08989(.A1(new_n8918_), .A2(new_n8926_), .B(\asqrt[22] ), .ZN(new_n9182_));
  XOR2_X1    g08990(.A1(new_n9182_), .A2(new_n8808_), .Z(new_n9183_));
  INV_X1     g08991(.I(new_n9183_), .ZN(new_n9184_));
  XOR2_X1    g08992(.A1(new_n8909_), .A2(\asqrt[33] ), .Z(new_n9185_));
  NOR2_X1    g08993(.A1(\asqrt[22] ), .A2(new_n9185_), .ZN(new_n9186_));
  XOR2_X1    g08994(.A1(new_n9186_), .A2(new_n8810_), .Z(new_n9187_));
  NOR2_X1    g08995(.A1(new_n8907_), .A2(new_n8916_), .ZN(new_n9188_));
  NOR2_X1    g08996(.A1(\asqrt[22] ), .A2(new_n9188_), .ZN(new_n9189_));
  XOR2_X1    g08997(.A1(new_n9189_), .A2(new_n8813_), .Z(new_n9190_));
  AOI21_X1   g08998(.A1(new_n8911_), .A2(new_n8915_), .B(\asqrt[22] ), .ZN(new_n9191_));
  XOR2_X1    g08999(.A1(new_n9191_), .A2(new_n8816_), .Z(new_n9192_));
  INV_X1     g09000(.I(new_n9192_), .ZN(new_n9193_));
  AOI21_X1   g09001(.A1(new_n8897_), .A2(new_n8905_), .B(\asqrt[22] ), .ZN(new_n9194_));
  XOR2_X1    g09002(.A1(new_n9194_), .A2(new_n8820_), .Z(new_n9195_));
  INV_X1     g09003(.I(new_n9195_), .ZN(new_n9196_));
  XOR2_X1    g09004(.A1(new_n8888_), .A2(\asqrt[29] ), .Z(new_n9197_));
  NOR2_X1    g09005(.A1(\asqrt[22] ), .A2(new_n9197_), .ZN(new_n9198_));
  XOR2_X1    g09006(.A1(new_n9198_), .A2(new_n8822_), .Z(new_n9199_));
  NOR2_X1    g09007(.A1(new_n8886_), .A2(new_n8895_), .ZN(new_n9200_));
  NOR2_X1    g09008(.A1(\asqrt[22] ), .A2(new_n9200_), .ZN(new_n9201_));
  XOR2_X1    g09009(.A1(new_n9201_), .A2(new_n8825_), .Z(new_n9202_));
  AOI21_X1   g09010(.A1(new_n8890_), .A2(new_n8894_), .B(\asqrt[22] ), .ZN(new_n9203_));
  XOR2_X1    g09011(.A1(new_n9203_), .A2(new_n8828_), .Z(new_n9204_));
  INV_X1     g09012(.I(new_n9204_), .ZN(new_n9205_));
  AOI21_X1   g09013(.A1(new_n8876_), .A2(new_n8884_), .B(\asqrt[22] ), .ZN(new_n9206_));
  XOR2_X1    g09014(.A1(new_n9206_), .A2(new_n8835_), .Z(new_n9207_));
  INV_X1     g09015(.I(new_n9207_), .ZN(new_n9208_));
  AOI21_X1   g09016(.A1(new_n8867_), .A2(new_n8875_), .B(\asqrt[22] ), .ZN(new_n9209_));
  XOR2_X1    g09017(.A1(new_n9209_), .A2(new_n8852_), .Z(new_n9210_));
  NAND2_X1   g09018(.A1(\asqrt[23] ), .A2(new_n8853_), .ZN(new_n9211_));
  NOR2_X1    g09019(.A1(new_n8864_), .A2(\a[46] ), .ZN(new_n9212_));
  AOI22_X1   g09020(.A1(new_n9211_), .A2(new_n8864_), .B1(\asqrt[23] ), .B2(new_n9212_), .ZN(new_n9213_));
  AOI21_X1   g09021(.A1(\asqrt[23] ), .A2(\a[46] ), .B(new_n8861_), .ZN(new_n9214_));
  NOR2_X1    g09022(.A1(new_n8871_), .A2(new_n9214_), .ZN(new_n9215_));
  NOR2_X1    g09023(.A1(\asqrt[22] ), .A2(new_n9215_), .ZN(new_n9216_));
  XOR2_X1    g09024(.A1(new_n9216_), .A2(new_n9213_), .Z(new_n9217_));
  NOR2_X1    g09025(.A1(new_n9135_), .A2(new_n9131_), .ZN(new_n9218_));
  AOI21_X1   g09026(.A1(new_n9114_), .A2(new_n9111_), .B(\asqrt[62] ), .ZN(new_n9219_));
  NOR3_X1    g09027(.A1(new_n9135_), .A2(new_n201_), .A3(new_n9131_), .ZN(new_n9220_));
  OAI22_X1   g09028(.A1(new_n9219_), .A2(new_n9220_), .B1(new_n9218_), .B2(new_n9140_), .ZN(new_n9221_));
  AOI21_X1   g09029(.A1(new_n9221_), .A2(new_n8968_), .B(new_n9144_), .ZN(new_n9222_));
  AOI21_X1   g09030(.A1(new_n9218_), .A2(new_n201_), .B(new_n9141_), .ZN(new_n9223_));
  NOR2_X1    g09031(.A1(new_n9218_), .A2(new_n201_), .ZN(new_n9224_));
  NOR3_X1    g09032(.A1(new_n9223_), .A2(new_n9224_), .A3(new_n8968_), .ZN(new_n9225_));
  NOR3_X1    g09033(.A1(new_n9222_), .A2(\asqrt[63] ), .A3(new_n9225_), .ZN(new_n9226_));
  NAND4_X1   g09034(.A1(new_n9226_), .A2(\asqrt[23] ), .A3(new_n9153_), .A4(new_n9155_), .ZN(new_n9227_));
  NAND2_X1   g09035(.A1(\asqrt[22] ), .A2(new_n8854_), .ZN(new_n9228_));
  AOI21_X1   g09036(.A1(new_n9227_), .A2(new_n9228_), .B(\a[46] ), .ZN(new_n9229_));
  NAND2_X1   g09037(.A1(new_n9146_), .A2(new_n193_), .ZN(new_n9230_));
  NAND3_X1   g09038(.A1(new_n9153_), .A2(new_n9155_), .A3(\asqrt[23] ), .ZN(new_n9231_));
  NOR3_X1    g09039(.A1(new_n9230_), .A2(new_n9225_), .A3(new_n9231_), .ZN(new_n9232_));
  NOR4_X1    g09040(.A1(new_n9222_), .A2(\asqrt[63] ), .A3(new_n9225_), .A4(new_n9156_), .ZN(new_n9233_));
  NOR2_X1    g09041(.A1(new_n9233_), .A2(new_n8856_), .ZN(new_n9234_));
  NOR3_X1    g09042(.A1(new_n9234_), .A2(new_n9232_), .A3(new_n8853_), .ZN(new_n9235_));
  OR2_X2     g09043(.A1(new_n9229_), .A2(new_n9235_), .Z(new_n9236_));
  NOR2_X1    g09044(.A1(\a[42] ), .A2(\a[43] ), .ZN(new_n9237_));
  INV_X1     g09045(.I(new_n9237_), .ZN(new_n9238_));
  NAND3_X1   g09046(.A1(\asqrt[22] ), .A2(\a[44] ), .A3(new_n9238_), .ZN(new_n9239_));
  INV_X1     g09047(.I(\a[44] ), .ZN(new_n9240_));
  OAI21_X1   g09048(.A1(\asqrt[22] ), .A2(new_n9240_), .B(new_n9237_), .ZN(new_n9241_));
  AOI21_X1   g09049(.A1(new_n9241_), .A2(new_n9239_), .B(new_n8849_), .ZN(new_n9242_));
  NOR3_X1    g09050(.A1(new_n8840_), .A2(\asqrt[63] ), .A3(new_n8843_), .ZN(new_n9243_));
  NAND2_X1   g09051(.A1(new_n9237_), .A2(new_n9240_), .ZN(new_n9244_));
  NAND3_X1   g09052(.A1(new_n8777_), .A2(new_n8779_), .A3(new_n9244_), .ZN(new_n9245_));
  NAND2_X1   g09053(.A1(new_n9243_), .A2(new_n9245_), .ZN(new_n9246_));
  NAND3_X1   g09054(.A1(\asqrt[22] ), .A2(\a[44] ), .A3(new_n9246_), .ZN(new_n9247_));
  INV_X1     g09055(.I(\a[45] ), .ZN(new_n9248_));
  NAND3_X1   g09056(.A1(\asqrt[22] ), .A2(new_n9240_), .A3(new_n9248_), .ZN(new_n9249_));
  OAI21_X1   g09057(.A1(new_n9233_), .A2(\a[44] ), .B(\a[45] ), .ZN(new_n9250_));
  NAND3_X1   g09058(.A1(new_n9247_), .A2(new_n9250_), .A3(new_n9249_), .ZN(new_n9251_));
  NOR3_X1    g09059(.A1(new_n9251_), .A2(new_n9242_), .A3(\asqrt[24] ), .ZN(new_n9252_));
  OAI21_X1   g09060(.A1(new_n9251_), .A2(new_n9242_), .B(\asqrt[24] ), .ZN(new_n9253_));
  OAI21_X1   g09061(.A1(new_n9236_), .A2(new_n9252_), .B(new_n9253_), .ZN(new_n9254_));
  OAI21_X1   g09062(.A1(new_n9254_), .A2(\asqrt[25] ), .B(new_n9217_), .ZN(new_n9255_));
  NAND2_X1   g09063(.A1(new_n9254_), .A2(\asqrt[25] ), .ZN(new_n9256_));
  NAND3_X1   g09064(.A1(new_n9255_), .A2(new_n9256_), .A3(new_n7690_), .ZN(new_n9257_));
  AOI21_X1   g09065(.A1(new_n9255_), .A2(new_n9256_), .B(new_n7690_), .ZN(new_n9258_));
  AOI21_X1   g09066(.A1(new_n9210_), .A2(new_n9257_), .B(new_n9258_), .ZN(new_n9259_));
  AOI21_X1   g09067(.A1(new_n9259_), .A2(new_n7331_), .B(new_n9208_), .ZN(new_n9260_));
  NAND2_X1   g09068(.A1(new_n9257_), .A2(new_n9210_), .ZN(new_n9261_));
  INV_X1     g09069(.I(new_n9217_), .ZN(new_n9262_));
  NOR2_X1    g09070(.A1(new_n9229_), .A2(new_n9235_), .ZN(new_n9263_));
  NOR3_X1    g09071(.A1(new_n9233_), .A2(new_n9240_), .A3(new_n9237_), .ZN(new_n9264_));
  AOI21_X1   g09072(.A1(new_n9233_), .A2(\a[44] ), .B(new_n9238_), .ZN(new_n9265_));
  OAI21_X1   g09073(.A1(new_n9264_), .A2(new_n9265_), .B(\asqrt[23] ), .ZN(new_n9266_));
  INV_X1     g09074(.I(new_n9246_), .ZN(new_n9267_));
  NOR3_X1    g09075(.A1(new_n9233_), .A2(new_n9240_), .A3(new_n9267_), .ZN(new_n9268_));
  NOR3_X1    g09076(.A1(new_n9233_), .A2(\a[44] ), .A3(\a[45] ), .ZN(new_n9269_));
  AOI21_X1   g09077(.A1(\asqrt[22] ), .A2(new_n9240_), .B(new_n9248_), .ZN(new_n9270_));
  NOR3_X1    g09078(.A1(new_n9268_), .A2(new_n9269_), .A3(new_n9270_), .ZN(new_n9271_));
  NAND3_X1   g09079(.A1(new_n9271_), .A2(new_n9266_), .A3(new_n8440_), .ZN(new_n9272_));
  AOI21_X1   g09080(.A1(new_n9271_), .A2(new_n9266_), .B(new_n8440_), .ZN(new_n9273_));
  AOI21_X1   g09081(.A1(new_n9263_), .A2(new_n9272_), .B(new_n9273_), .ZN(new_n9274_));
  AOI21_X1   g09082(.A1(new_n9274_), .A2(new_n8077_), .B(new_n9262_), .ZN(new_n9275_));
  NAND2_X1   g09083(.A1(new_n9272_), .A2(new_n9263_), .ZN(new_n9276_));
  AOI21_X1   g09084(.A1(new_n9276_), .A2(new_n9253_), .B(new_n8077_), .ZN(new_n9277_));
  OAI21_X1   g09085(.A1(new_n9275_), .A2(new_n9277_), .B(\asqrt[26] ), .ZN(new_n9278_));
  AOI21_X1   g09086(.A1(new_n9261_), .A2(new_n9278_), .B(new_n7331_), .ZN(new_n9279_));
  NOR3_X1    g09087(.A1(new_n9260_), .A2(\asqrt[28] ), .A3(new_n9279_), .ZN(new_n9280_));
  OAI21_X1   g09088(.A1(new_n9260_), .A2(new_n9279_), .B(\asqrt[28] ), .ZN(new_n9281_));
  OAI21_X1   g09089(.A1(new_n9205_), .A2(new_n9280_), .B(new_n9281_), .ZN(new_n9282_));
  OAI21_X1   g09090(.A1(new_n9282_), .A2(\asqrt[29] ), .B(new_n9202_), .ZN(new_n9283_));
  NAND2_X1   g09091(.A1(new_n9282_), .A2(\asqrt[29] ), .ZN(new_n9284_));
  NAND3_X1   g09092(.A1(new_n9283_), .A2(new_n9284_), .A3(new_n6275_), .ZN(new_n9285_));
  AOI21_X1   g09093(.A1(new_n9283_), .A2(new_n9284_), .B(new_n6275_), .ZN(new_n9286_));
  AOI21_X1   g09094(.A1(new_n9199_), .A2(new_n9285_), .B(new_n9286_), .ZN(new_n9287_));
  AOI21_X1   g09095(.A1(new_n9287_), .A2(new_n5947_), .B(new_n9196_), .ZN(new_n9288_));
  NAND2_X1   g09096(.A1(new_n9285_), .A2(new_n9199_), .ZN(new_n9289_));
  INV_X1     g09097(.I(new_n9202_), .ZN(new_n9290_));
  INV_X1     g09098(.I(new_n9210_), .ZN(new_n9291_));
  NOR3_X1    g09099(.A1(new_n9275_), .A2(\asqrt[26] ), .A3(new_n9277_), .ZN(new_n9292_));
  OAI21_X1   g09100(.A1(new_n9291_), .A2(new_n9292_), .B(new_n9278_), .ZN(new_n9293_));
  OAI21_X1   g09101(.A1(new_n9293_), .A2(\asqrt[27] ), .B(new_n9207_), .ZN(new_n9294_));
  NAND2_X1   g09102(.A1(new_n9293_), .A2(\asqrt[27] ), .ZN(new_n9295_));
  NAND3_X1   g09103(.A1(new_n9294_), .A2(new_n9295_), .A3(new_n6966_), .ZN(new_n9296_));
  AOI21_X1   g09104(.A1(new_n9294_), .A2(new_n9295_), .B(new_n6966_), .ZN(new_n9297_));
  AOI21_X1   g09105(.A1(new_n9204_), .A2(new_n9296_), .B(new_n9297_), .ZN(new_n9298_));
  AOI21_X1   g09106(.A1(new_n9298_), .A2(new_n6636_), .B(new_n9290_), .ZN(new_n9299_));
  NAND2_X1   g09107(.A1(new_n9296_), .A2(new_n9204_), .ZN(new_n9300_));
  AOI21_X1   g09108(.A1(new_n9300_), .A2(new_n9281_), .B(new_n6636_), .ZN(new_n9301_));
  OAI21_X1   g09109(.A1(new_n9299_), .A2(new_n9301_), .B(\asqrt[30] ), .ZN(new_n9302_));
  AOI21_X1   g09110(.A1(new_n9289_), .A2(new_n9302_), .B(new_n5947_), .ZN(new_n9303_));
  NOR3_X1    g09111(.A1(new_n9288_), .A2(\asqrt[32] ), .A3(new_n9303_), .ZN(new_n9304_));
  OAI21_X1   g09112(.A1(new_n9288_), .A2(new_n9303_), .B(\asqrt[32] ), .ZN(new_n9305_));
  OAI21_X1   g09113(.A1(new_n9193_), .A2(new_n9304_), .B(new_n9305_), .ZN(new_n9306_));
  OAI21_X1   g09114(.A1(new_n9306_), .A2(\asqrt[33] ), .B(new_n9190_), .ZN(new_n9307_));
  NAND2_X1   g09115(.A1(new_n9306_), .A2(\asqrt[33] ), .ZN(new_n9308_));
  NAND3_X1   g09116(.A1(new_n9307_), .A2(new_n9308_), .A3(new_n5029_), .ZN(new_n9309_));
  AOI21_X1   g09117(.A1(new_n9307_), .A2(new_n9308_), .B(new_n5029_), .ZN(new_n9310_));
  AOI21_X1   g09118(.A1(new_n9187_), .A2(new_n9309_), .B(new_n9310_), .ZN(new_n9311_));
  AOI21_X1   g09119(.A1(new_n9311_), .A2(new_n4751_), .B(new_n9184_), .ZN(new_n9312_));
  NAND2_X1   g09120(.A1(new_n9309_), .A2(new_n9187_), .ZN(new_n9313_));
  INV_X1     g09121(.I(new_n9190_), .ZN(new_n9314_));
  INV_X1     g09122(.I(new_n9199_), .ZN(new_n9315_));
  NOR3_X1    g09123(.A1(new_n9299_), .A2(\asqrt[30] ), .A3(new_n9301_), .ZN(new_n9316_));
  OAI21_X1   g09124(.A1(new_n9315_), .A2(new_n9316_), .B(new_n9302_), .ZN(new_n9317_));
  OAI21_X1   g09125(.A1(new_n9317_), .A2(\asqrt[31] ), .B(new_n9195_), .ZN(new_n9318_));
  NAND2_X1   g09126(.A1(new_n9317_), .A2(\asqrt[31] ), .ZN(new_n9319_));
  NAND3_X1   g09127(.A1(new_n9318_), .A2(new_n9319_), .A3(new_n5643_), .ZN(new_n9320_));
  AOI21_X1   g09128(.A1(new_n9318_), .A2(new_n9319_), .B(new_n5643_), .ZN(new_n9321_));
  AOI21_X1   g09129(.A1(new_n9192_), .A2(new_n9320_), .B(new_n9321_), .ZN(new_n9322_));
  AOI21_X1   g09130(.A1(new_n9322_), .A2(new_n5336_), .B(new_n9314_), .ZN(new_n9323_));
  NAND2_X1   g09131(.A1(new_n9320_), .A2(new_n9192_), .ZN(new_n9324_));
  AOI21_X1   g09132(.A1(new_n9324_), .A2(new_n9305_), .B(new_n5336_), .ZN(new_n9325_));
  OAI21_X1   g09133(.A1(new_n9323_), .A2(new_n9325_), .B(\asqrt[34] ), .ZN(new_n9326_));
  AOI21_X1   g09134(.A1(new_n9313_), .A2(new_n9326_), .B(new_n4751_), .ZN(new_n9327_));
  NOR3_X1    g09135(.A1(new_n9312_), .A2(\asqrt[36] ), .A3(new_n9327_), .ZN(new_n9328_));
  OAI21_X1   g09136(.A1(new_n9312_), .A2(new_n9327_), .B(\asqrt[36] ), .ZN(new_n9329_));
  OAI21_X1   g09137(.A1(new_n9181_), .A2(new_n9328_), .B(new_n9329_), .ZN(new_n9330_));
  OAI21_X1   g09138(.A1(new_n9330_), .A2(\asqrt[37] ), .B(new_n9178_), .ZN(new_n9331_));
  NAND2_X1   g09139(.A1(new_n9330_), .A2(\asqrt[37] ), .ZN(new_n9332_));
  NAND3_X1   g09140(.A1(new_n9331_), .A2(new_n9332_), .A3(new_n3925_), .ZN(new_n9333_));
  AOI21_X1   g09141(.A1(new_n9331_), .A2(new_n9332_), .B(new_n3925_), .ZN(new_n9334_));
  AOI21_X1   g09142(.A1(new_n9175_), .A2(new_n9333_), .B(new_n9334_), .ZN(new_n9335_));
  AOI21_X1   g09143(.A1(new_n9335_), .A2(new_n3681_), .B(new_n9172_), .ZN(new_n9336_));
  NAND2_X1   g09144(.A1(new_n9333_), .A2(new_n9175_), .ZN(new_n9337_));
  INV_X1     g09145(.I(new_n9178_), .ZN(new_n9338_));
  INV_X1     g09146(.I(new_n9187_), .ZN(new_n9339_));
  NOR3_X1    g09147(.A1(new_n9323_), .A2(\asqrt[34] ), .A3(new_n9325_), .ZN(new_n9340_));
  OAI21_X1   g09148(.A1(new_n9339_), .A2(new_n9340_), .B(new_n9326_), .ZN(new_n9341_));
  OAI21_X1   g09149(.A1(new_n9341_), .A2(\asqrt[35] ), .B(new_n9183_), .ZN(new_n9342_));
  NAND2_X1   g09150(.A1(new_n9341_), .A2(\asqrt[35] ), .ZN(new_n9343_));
  NAND3_X1   g09151(.A1(new_n9342_), .A2(new_n9343_), .A3(new_n4461_), .ZN(new_n9344_));
  AOI21_X1   g09152(.A1(new_n9342_), .A2(new_n9343_), .B(new_n4461_), .ZN(new_n9345_));
  AOI21_X1   g09153(.A1(new_n9180_), .A2(new_n9344_), .B(new_n9345_), .ZN(new_n9346_));
  AOI21_X1   g09154(.A1(new_n9346_), .A2(new_n4196_), .B(new_n9338_), .ZN(new_n9347_));
  NAND2_X1   g09155(.A1(new_n9344_), .A2(new_n9180_), .ZN(new_n9348_));
  AOI21_X1   g09156(.A1(new_n9348_), .A2(new_n9329_), .B(new_n4196_), .ZN(new_n9349_));
  OAI21_X1   g09157(.A1(new_n9347_), .A2(new_n9349_), .B(\asqrt[38] ), .ZN(new_n9350_));
  AOI21_X1   g09158(.A1(new_n9337_), .A2(new_n9350_), .B(new_n3681_), .ZN(new_n9351_));
  NOR3_X1    g09159(.A1(new_n9336_), .A2(\asqrt[40] ), .A3(new_n9351_), .ZN(new_n9352_));
  OAI21_X1   g09160(.A1(new_n9336_), .A2(new_n9351_), .B(\asqrt[40] ), .ZN(new_n9353_));
  OAI21_X1   g09161(.A1(new_n9169_), .A2(new_n9352_), .B(new_n9353_), .ZN(new_n9354_));
  OAI21_X1   g09162(.A1(new_n9354_), .A2(\asqrt[41] ), .B(new_n9166_), .ZN(new_n9355_));
  NAND2_X1   g09163(.A1(new_n9354_), .A2(\asqrt[41] ), .ZN(new_n9356_));
  NAND3_X1   g09164(.A1(new_n9355_), .A2(new_n9356_), .A3(new_n2960_), .ZN(new_n9357_));
  AOI21_X1   g09165(.A1(new_n9355_), .A2(new_n9356_), .B(new_n2960_), .ZN(new_n9358_));
  AOI21_X1   g09166(.A1(new_n9163_), .A2(new_n9357_), .B(new_n9358_), .ZN(new_n9359_));
  NAND2_X1   g09167(.A1(new_n9359_), .A2(new_n2749_), .ZN(new_n9360_));
  INV_X1     g09168(.I(new_n9163_), .ZN(new_n9361_));
  INV_X1     g09169(.I(new_n9166_), .ZN(new_n9362_));
  INV_X1     g09170(.I(new_n9175_), .ZN(new_n9363_));
  NOR3_X1    g09171(.A1(new_n9347_), .A2(\asqrt[38] ), .A3(new_n9349_), .ZN(new_n9364_));
  OAI21_X1   g09172(.A1(new_n9363_), .A2(new_n9364_), .B(new_n9350_), .ZN(new_n9365_));
  OAI21_X1   g09173(.A1(new_n9365_), .A2(\asqrt[39] ), .B(new_n9171_), .ZN(new_n9366_));
  NAND2_X1   g09174(.A1(new_n9365_), .A2(\asqrt[39] ), .ZN(new_n9367_));
  NAND3_X1   g09175(.A1(new_n9366_), .A2(new_n9367_), .A3(new_n3427_), .ZN(new_n9368_));
  AOI21_X1   g09176(.A1(new_n9366_), .A2(new_n9367_), .B(new_n3427_), .ZN(new_n9369_));
  AOI21_X1   g09177(.A1(new_n9168_), .A2(new_n9368_), .B(new_n9369_), .ZN(new_n9370_));
  AOI21_X1   g09178(.A1(new_n9370_), .A2(new_n3195_), .B(new_n9362_), .ZN(new_n9371_));
  NAND2_X1   g09179(.A1(new_n9368_), .A2(new_n9168_), .ZN(new_n9372_));
  AOI21_X1   g09180(.A1(new_n9372_), .A2(new_n9353_), .B(new_n3195_), .ZN(new_n9373_));
  NOR3_X1    g09181(.A1(new_n9371_), .A2(\asqrt[42] ), .A3(new_n9373_), .ZN(new_n9374_));
  OAI21_X1   g09182(.A1(new_n9371_), .A2(new_n9373_), .B(\asqrt[42] ), .ZN(new_n9375_));
  OAI21_X1   g09183(.A1(new_n9361_), .A2(new_n9374_), .B(new_n9375_), .ZN(new_n9376_));
  NAND2_X1   g09184(.A1(new_n9376_), .A2(\asqrt[43] ), .ZN(new_n9377_));
  NOR2_X1    g09185(.A1(new_n9115_), .A2(\asqrt[62] ), .ZN(new_n9378_));
  NOR2_X1    g09186(.A1(new_n9378_), .A2(new_n9224_), .ZN(new_n9379_));
  XOR2_X1    g09187(.A1(new_n9139_), .A2(new_n8745_), .Z(new_n9380_));
  OAI21_X1   g09188(.A1(\asqrt[22] ), .A2(new_n9379_), .B(new_n9380_), .ZN(new_n9381_));
  INV_X1     g09189(.I(new_n9381_), .ZN(new_n9382_));
  AOI21_X1   g09190(.A1(new_n9123_), .A2(new_n9128_), .B(\asqrt[22] ), .ZN(new_n9383_));
  XOR2_X1    g09191(.A1(new_n9383_), .A2(new_n8974_), .Z(new_n9384_));
  INV_X1     g09192(.I(new_n9384_), .ZN(new_n9385_));
  AOI21_X1   g09193(.A1(new_n9103_), .A2(new_n9122_), .B(\asqrt[22] ), .ZN(new_n9386_));
  XOR2_X1    g09194(.A1(new_n9386_), .A2(new_n8978_), .Z(new_n9387_));
  INV_X1     g09195(.I(new_n9387_), .ZN(new_n9388_));
  NOR2_X1    g09196(.A1(new_n9121_), .A2(new_n9117_), .ZN(new_n9389_));
  NOR2_X1    g09197(.A1(\asqrt[22] ), .A2(new_n9389_), .ZN(new_n9390_));
  XOR2_X1    g09198(.A1(new_n9390_), .A2(new_n8980_), .Z(new_n9391_));
  NOR2_X1    g09199(.A1(new_n9092_), .A2(new_n9101_), .ZN(new_n9392_));
  NOR2_X1    g09200(.A1(\asqrt[22] ), .A2(new_n9392_), .ZN(new_n9393_));
  XOR2_X1    g09201(.A1(new_n9393_), .A2(new_n8983_), .Z(new_n9394_));
  AOI21_X1   g09202(.A1(new_n9096_), .A2(new_n9100_), .B(\asqrt[22] ), .ZN(new_n9395_));
  XOR2_X1    g09203(.A1(new_n9395_), .A2(new_n8986_), .Z(new_n9396_));
  INV_X1     g09204(.I(new_n9396_), .ZN(new_n9397_));
  AOI21_X1   g09205(.A1(new_n9082_), .A2(new_n9090_), .B(\asqrt[22] ), .ZN(new_n9398_));
  XOR2_X1    g09206(.A1(new_n9398_), .A2(new_n8990_), .Z(new_n9399_));
  INV_X1     g09207(.I(new_n9399_), .ZN(new_n9400_));
  XOR2_X1    g09208(.A1(new_n9073_), .A2(\asqrt[53] ), .Z(new_n9401_));
  NOR2_X1    g09209(.A1(\asqrt[22] ), .A2(new_n9401_), .ZN(new_n9402_));
  XOR2_X1    g09210(.A1(new_n9402_), .A2(new_n8992_), .Z(new_n9403_));
  NOR2_X1    g09211(.A1(new_n9071_), .A2(new_n9080_), .ZN(new_n9404_));
  NOR2_X1    g09212(.A1(\asqrt[22] ), .A2(new_n9404_), .ZN(new_n9405_));
  XOR2_X1    g09213(.A1(new_n9405_), .A2(new_n8995_), .Z(new_n9406_));
  AOI21_X1   g09214(.A1(new_n9075_), .A2(new_n9079_), .B(\asqrt[22] ), .ZN(new_n9407_));
  XOR2_X1    g09215(.A1(new_n9407_), .A2(new_n8998_), .Z(new_n9408_));
  INV_X1     g09216(.I(new_n9408_), .ZN(new_n9409_));
  AOI21_X1   g09217(.A1(new_n9061_), .A2(new_n9069_), .B(\asqrt[22] ), .ZN(new_n9410_));
  XOR2_X1    g09218(.A1(new_n9410_), .A2(new_n9002_), .Z(new_n9411_));
  INV_X1     g09219(.I(new_n9411_), .ZN(new_n9412_));
  XOR2_X1    g09220(.A1(new_n9052_), .A2(\asqrt[49] ), .Z(new_n9413_));
  NOR2_X1    g09221(.A1(\asqrt[22] ), .A2(new_n9413_), .ZN(new_n9414_));
  XOR2_X1    g09222(.A1(new_n9414_), .A2(new_n9004_), .Z(new_n9415_));
  NOR2_X1    g09223(.A1(new_n9050_), .A2(new_n9059_), .ZN(new_n9416_));
  NOR2_X1    g09224(.A1(\asqrt[22] ), .A2(new_n9416_), .ZN(new_n9417_));
  XOR2_X1    g09225(.A1(new_n9417_), .A2(new_n9007_), .Z(new_n9418_));
  AOI21_X1   g09226(.A1(new_n9054_), .A2(new_n9058_), .B(\asqrt[22] ), .ZN(new_n9419_));
  XOR2_X1    g09227(.A1(new_n9419_), .A2(new_n9010_), .Z(new_n9420_));
  INV_X1     g09228(.I(new_n9420_), .ZN(new_n9421_));
  AOI21_X1   g09229(.A1(new_n9040_), .A2(new_n9048_), .B(\asqrt[22] ), .ZN(new_n9422_));
  XOR2_X1    g09230(.A1(new_n9422_), .A2(new_n9014_), .Z(new_n9423_));
  INV_X1     g09231(.I(new_n9423_), .ZN(new_n9424_));
  XOR2_X1    g09232(.A1(new_n9031_), .A2(\asqrt[45] ), .Z(new_n9425_));
  NOR2_X1    g09233(.A1(\asqrt[22] ), .A2(new_n9425_), .ZN(new_n9426_));
  XOR2_X1    g09234(.A1(new_n9426_), .A2(new_n9016_), .Z(new_n9427_));
  NOR2_X1    g09235(.A1(new_n9029_), .A2(new_n9038_), .ZN(new_n9428_));
  NOR2_X1    g09236(.A1(\asqrt[22] ), .A2(new_n9428_), .ZN(new_n9429_));
  XOR2_X1    g09237(.A1(new_n9429_), .A2(new_n9019_), .Z(new_n9430_));
  AOI21_X1   g09238(.A1(new_n9033_), .A2(new_n9037_), .B(\asqrt[22] ), .ZN(new_n9431_));
  XOR2_X1    g09239(.A1(new_n9431_), .A2(new_n9022_), .Z(new_n9432_));
  INV_X1     g09240(.I(new_n9432_), .ZN(new_n9433_));
  INV_X1     g09241(.I(new_n9160_), .ZN(new_n9434_));
  AOI21_X1   g09242(.A1(new_n9359_), .A2(new_n2749_), .B(new_n9434_), .ZN(new_n9435_));
  NAND2_X1   g09243(.A1(new_n9357_), .A2(new_n9163_), .ZN(new_n9436_));
  AOI21_X1   g09244(.A1(new_n9436_), .A2(new_n9375_), .B(new_n2749_), .ZN(new_n9437_));
  NOR3_X1    g09245(.A1(new_n9435_), .A2(\asqrt[44] ), .A3(new_n9437_), .ZN(new_n9438_));
  OAI21_X1   g09246(.A1(new_n9435_), .A2(new_n9437_), .B(\asqrt[44] ), .ZN(new_n9439_));
  OAI21_X1   g09247(.A1(new_n9433_), .A2(new_n9438_), .B(new_n9439_), .ZN(new_n9440_));
  OAI21_X1   g09248(.A1(new_n9440_), .A2(\asqrt[45] ), .B(new_n9430_), .ZN(new_n9441_));
  NAND2_X1   g09249(.A1(new_n9440_), .A2(\asqrt[45] ), .ZN(new_n9442_));
  NAND3_X1   g09250(.A1(new_n9441_), .A2(new_n9442_), .A3(new_n2134_), .ZN(new_n9443_));
  AOI21_X1   g09251(.A1(new_n9441_), .A2(new_n9442_), .B(new_n2134_), .ZN(new_n9444_));
  AOI21_X1   g09252(.A1(new_n9427_), .A2(new_n9443_), .B(new_n9444_), .ZN(new_n9445_));
  AOI21_X1   g09253(.A1(new_n9445_), .A2(new_n1953_), .B(new_n9424_), .ZN(new_n9446_));
  NAND2_X1   g09254(.A1(new_n9443_), .A2(new_n9427_), .ZN(new_n9447_));
  INV_X1     g09255(.I(new_n9430_), .ZN(new_n9448_));
  OAI21_X1   g09256(.A1(new_n9376_), .A2(\asqrt[43] ), .B(new_n9160_), .ZN(new_n9449_));
  NAND3_X1   g09257(.A1(new_n9449_), .A2(new_n9377_), .A3(new_n2531_), .ZN(new_n9450_));
  AOI21_X1   g09258(.A1(new_n9449_), .A2(new_n9377_), .B(new_n2531_), .ZN(new_n9451_));
  AOI21_X1   g09259(.A1(new_n9432_), .A2(new_n9450_), .B(new_n9451_), .ZN(new_n9452_));
  AOI21_X1   g09260(.A1(new_n9452_), .A2(new_n2332_), .B(new_n9448_), .ZN(new_n9453_));
  NAND2_X1   g09261(.A1(new_n9450_), .A2(new_n9432_), .ZN(new_n9454_));
  AOI21_X1   g09262(.A1(new_n9454_), .A2(new_n9439_), .B(new_n2332_), .ZN(new_n9455_));
  OAI21_X1   g09263(.A1(new_n9453_), .A2(new_n9455_), .B(\asqrt[46] ), .ZN(new_n9456_));
  AOI21_X1   g09264(.A1(new_n9447_), .A2(new_n9456_), .B(new_n1953_), .ZN(new_n9457_));
  NOR3_X1    g09265(.A1(new_n9446_), .A2(\asqrt[48] ), .A3(new_n9457_), .ZN(new_n9458_));
  OAI21_X1   g09266(.A1(new_n9446_), .A2(new_n9457_), .B(\asqrt[48] ), .ZN(new_n9459_));
  OAI21_X1   g09267(.A1(new_n9421_), .A2(new_n9458_), .B(new_n9459_), .ZN(new_n9460_));
  OAI21_X1   g09268(.A1(new_n9460_), .A2(\asqrt[49] ), .B(new_n9418_), .ZN(new_n9461_));
  NAND2_X1   g09269(.A1(new_n9460_), .A2(\asqrt[49] ), .ZN(new_n9462_));
  NAND3_X1   g09270(.A1(new_n9461_), .A2(new_n9462_), .A3(new_n1463_), .ZN(new_n9463_));
  AOI21_X1   g09271(.A1(new_n9461_), .A2(new_n9462_), .B(new_n1463_), .ZN(new_n9464_));
  AOI21_X1   g09272(.A1(new_n9415_), .A2(new_n9463_), .B(new_n9464_), .ZN(new_n9465_));
  AOI21_X1   g09273(.A1(new_n9465_), .A2(new_n1305_), .B(new_n9412_), .ZN(new_n9466_));
  NAND2_X1   g09274(.A1(new_n9463_), .A2(new_n9415_), .ZN(new_n9467_));
  INV_X1     g09275(.I(new_n9418_), .ZN(new_n9468_));
  INV_X1     g09276(.I(new_n9427_), .ZN(new_n9469_));
  NOR3_X1    g09277(.A1(new_n9453_), .A2(\asqrt[46] ), .A3(new_n9455_), .ZN(new_n9470_));
  OAI21_X1   g09278(.A1(new_n9469_), .A2(new_n9470_), .B(new_n9456_), .ZN(new_n9471_));
  OAI21_X1   g09279(.A1(new_n9471_), .A2(\asqrt[47] ), .B(new_n9423_), .ZN(new_n9472_));
  NAND2_X1   g09280(.A1(new_n9471_), .A2(\asqrt[47] ), .ZN(new_n9473_));
  NAND3_X1   g09281(.A1(new_n9472_), .A2(new_n9473_), .A3(new_n1778_), .ZN(new_n9474_));
  AOI21_X1   g09282(.A1(new_n9472_), .A2(new_n9473_), .B(new_n1778_), .ZN(new_n9475_));
  AOI21_X1   g09283(.A1(new_n9420_), .A2(new_n9474_), .B(new_n9475_), .ZN(new_n9476_));
  AOI21_X1   g09284(.A1(new_n9476_), .A2(new_n1632_), .B(new_n9468_), .ZN(new_n9477_));
  NAND2_X1   g09285(.A1(new_n9474_), .A2(new_n9420_), .ZN(new_n9478_));
  AOI21_X1   g09286(.A1(new_n9478_), .A2(new_n9459_), .B(new_n1632_), .ZN(new_n9479_));
  OAI21_X1   g09287(.A1(new_n9477_), .A2(new_n9479_), .B(\asqrt[50] ), .ZN(new_n9480_));
  AOI21_X1   g09288(.A1(new_n9467_), .A2(new_n9480_), .B(new_n1305_), .ZN(new_n9481_));
  NOR3_X1    g09289(.A1(new_n9466_), .A2(\asqrt[52] ), .A3(new_n9481_), .ZN(new_n9482_));
  OAI21_X1   g09290(.A1(new_n9466_), .A2(new_n9481_), .B(\asqrt[52] ), .ZN(new_n9483_));
  OAI21_X1   g09291(.A1(new_n9409_), .A2(new_n9482_), .B(new_n9483_), .ZN(new_n9484_));
  OAI21_X1   g09292(.A1(new_n9484_), .A2(\asqrt[53] ), .B(new_n9406_), .ZN(new_n9485_));
  NAND2_X1   g09293(.A1(new_n9484_), .A2(\asqrt[53] ), .ZN(new_n9486_));
  NAND3_X1   g09294(.A1(new_n9485_), .A2(new_n9486_), .A3(new_n860_), .ZN(new_n9487_));
  AOI21_X1   g09295(.A1(new_n9485_), .A2(new_n9486_), .B(new_n860_), .ZN(new_n9488_));
  AOI21_X1   g09296(.A1(new_n9403_), .A2(new_n9487_), .B(new_n9488_), .ZN(new_n9489_));
  AOI21_X1   g09297(.A1(new_n9489_), .A2(new_n744_), .B(new_n9400_), .ZN(new_n9490_));
  NAND2_X1   g09298(.A1(new_n9487_), .A2(new_n9403_), .ZN(new_n9491_));
  INV_X1     g09299(.I(new_n9406_), .ZN(new_n9492_));
  INV_X1     g09300(.I(new_n9415_), .ZN(new_n9493_));
  NOR3_X1    g09301(.A1(new_n9477_), .A2(\asqrt[50] ), .A3(new_n9479_), .ZN(new_n9494_));
  OAI21_X1   g09302(.A1(new_n9493_), .A2(new_n9494_), .B(new_n9480_), .ZN(new_n9495_));
  OAI21_X1   g09303(.A1(new_n9495_), .A2(\asqrt[51] ), .B(new_n9411_), .ZN(new_n9496_));
  NAND2_X1   g09304(.A1(new_n9495_), .A2(\asqrt[51] ), .ZN(new_n9497_));
  NAND3_X1   g09305(.A1(new_n9496_), .A2(new_n9497_), .A3(new_n1150_), .ZN(new_n9498_));
  AOI21_X1   g09306(.A1(new_n9496_), .A2(new_n9497_), .B(new_n1150_), .ZN(new_n9499_));
  AOI21_X1   g09307(.A1(new_n9408_), .A2(new_n9498_), .B(new_n9499_), .ZN(new_n9500_));
  AOI21_X1   g09308(.A1(new_n9500_), .A2(new_n1006_), .B(new_n9492_), .ZN(new_n9501_));
  NAND2_X1   g09309(.A1(new_n9498_), .A2(new_n9408_), .ZN(new_n9502_));
  AOI21_X1   g09310(.A1(new_n9502_), .A2(new_n9483_), .B(new_n1006_), .ZN(new_n9503_));
  OAI21_X1   g09311(.A1(new_n9501_), .A2(new_n9503_), .B(\asqrt[54] ), .ZN(new_n9504_));
  AOI21_X1   g09312(.A1(new_n9491_), .A2(new_n9504_), .B(new_n744_), .ZN(new_n9505_));
  NOR3_X1    g09313(.A1(new_n9490_), .A2(\asqrt[56] ), .A3(new_n9505_), .ZN(new_n9506_));
  OAI21_X1   g09314(.A1(new_n9490_), .A2(new_n9505_), .B(\asqrt[56] ), .ZN(new_n9507_));
  OAI21_X1   g09315(.A1(new_n9397_), .A2(new_n9506_), .B(new_n9507_), .ZN(new_n9508_));
  OAI21_X1   g09316(.A1(new_n9508_), .A2(\asqrt[57] ), .B(new_n9394_), .ZN(new_n9509_));
  NAND2_X1   g09317(.A1(new_n9508_), .A2(\asqrt[57] ), .ZN(new_n9510_));
  NAND3_X1   g09318(.A1(new_n9509_), .A2(new_n9510_), .A3(new_n423_), .ZN(new_n9511_));
  AOI21_X1   g09319(.A1(new_n9509_), .A2(new_n9510_), .B(new_n423_), .ZN(new_n9512_));
  AOI21_X1   g09320(.A1(new_n9391_), .A2(new_n9511_), .B(new_n9512_), .ZN(new_n9513_));
  AOI21_X1   g09321(.A1(new_n9513_), .A2(new_n337_), .B(new_n9388_), .ZN(new_n9514_));
  NAND2_X1   g09322(.A1(new_n9511_), .A2(new_n9391_), .ZN(new_n9515_));
  INV_X1     g09323(.I(new_n9394_), .ZN(new_n9516_));
  INV_X1     g09324(.I(new_n9403_), .ZN(new_n9517_));
  NOR3_X1    g09325(.A1(new_n9501_), .A2(\asqrt[54] ), .A3(new_n9503_), .ZN(new_n9518_));
  OAI21_X1   g09326(.A1(new_n9517_), .A2(new_n9518_), .B(new_n9504_), .ZN(new_n9519_));
  OAI21_X1   g09327(.A1(new_n9519_), .A2(\asqrt[55] ), .B(new_n9399_), .ZN(new_n9520_));
  NAND2_X1   g09328(.A1(new_n9519_), .A2(\asqrt[55] ), .ZN(new_n9521_));
  NAND3_X1   g09329(.A1(new_n9520_), .A2(new_n9521_), .A3(new_n634_), .ZN(new_n9522_));
  AOI21_X1   g09330(.A1(new_n9520_), .A2(new_n9521_), .B(new_n634_), .ZN(new_n9523_));
  AOI21_X1   g09331(.A1(new_n9396_), .A2(new_n9522_), .B(new_n9523_), .ZN(new_n9524_));
  AOI21_X1   g09332(.A1(new_n9524_), .A2(new_n531_), .B(new_n9516_), .ZN(new_n9525_));
  NAND2_X1   g09333(.A1(new_n9522_), .A2(new_n9396_), .ZN(new_n9526_));
  AOI21_X1   g09334(.A1(new_n9526_), .A2(new_n9507_), .B(new_n531_), .ZN(new_n9527_));
  OAI21_X1   g09335(.A1(new_n9525_), .A2(new_n9527_), .B(\asqrt[58] ), .ZN(new_n9528_));
  AOI21_X1   g09336(.A1(new_n9515_), .A2(new_n9528_), .B(new_n337_), .ZN(new_n9529_));
  NOR3_X1    g09337(.A1(new_n9514_), .A2(\asqrt[60] ), .A3(new_n9529_), .ZN(new_n9530_));
  NOR2_X1    g09338(.A1(new_n9530_), .A2(new_n9385_), .ZN(new_n9531_));
  INV_X1     g09339(.I(new_n9391_), .ZN(new_n9532_));
  NOR3_X1    g09340(.A1(new_n9525_), .A2(\asqrt[58] ), .A3(new_n9527_), .ZN(new_n9533_));
  OAI21_X1   g09341(.A1(new_n9532_), .A2(new_n9533_), .B(new_n9528_), .ZN(new_n9534_));
  OAI21_X1   g09342(.A1(new_n9534_), .A2(\asqrt[59] ), .B(new_n9387_), .ZN(new_n9535_));
  NOR2_X1    g09343(.A1(new_n9533_), .A2(new_n9532_), .ZN(new_n9536_));
  OAI21_X1   g09344(.A1(new_n9536_), .A2(new_n9512_), .B(\asqrt[59] ), .ZN(new_n9537_));
  AOI21_X1   g09345(.A1(new_n9535_), .A2(new_n9537_), .B(new_n266_), .ZN(new_n9538_));
  OAI21_X1   g09346(.A1(new_n9531_), .A2(new_n9538_), .B(\asqrt[61] ), .ZN(new_n9539_));
  OAI21_X1   g09347(.A1(new_n9514_), .A2(new_n9529_), .B(\asqrt[60] ), .ZN(new_n9540_));
  OAI21_X1   g09348(.A1(new_n9385_), .A2(new_n9530_), .B(new_n9540_), .ZN(new_n9541_));
  AOI21_X1   g09349(.A1(new_n9129_), .A2(new_n9109_), .B(\asqrt[22] ), .ZN(new_n9542_));
  XOR2_X1    g09350(.A1(new_n9542_), .A2(new_n8971_), .Z(new_n9543_));
  OAI21_X1   g09351(.A1(new_n9541_), .A2(\asqrt[61] ), .B(new_n9543_), .ZN(new_n9544_));
  NAND2_X1   g09352(.A1(new_n9544_), .A2(new_n9539_), .ZN(new_n9545_));
  NAND3_X1   g09353(.A1(new_n9535_), .A2(new_n266_), .A3(new_n9537_), .ZN(new_n9546_));
  NAND2_X1   g09354(.A1(new_n9546_), .A2(new_n9384_), .ZN(new_n9547_));
  AOI21_X1   g09355(.A1(new_n9547_), .A2(new_n9540_), .B(new_n239_), .ZN(new_n9548_));
  AOI21_X1   g09356(.A1(new_n9384_), .A2(new_n9546_), .B(new_n9538_), .ZN(new_n9549_));
  INV_X1     g09357(.I(new_n9543_), .ZN(new_n9550_));
  AOI21_X1   g09358(.A1(new_n9549_), .A2(new_n239_), .B(new_n9550_), .ZN(new_n9551_));
  OAI21_X1   g09359(.A1(new_n9551_), .A2(new_n9548_), .B(new_n201_), .ZN(new_n9552_));
  NAND3_X1   g09360(.A1(new_n9544_), .A2(\asqrt[62] ), .A3(new_n9539_), .ZN(new_n9553_));
  NAND2_X1   g09361(.A1(new_n9133_), .A2(new_n239_), .ZN(new_n9554_));
  AOI21_X1   g09362(.A1(new_n9111_), .A2(new_n9554_), .B(\asqrt[22] ), .ZN(new_n9555_));
  XOR2_X1    g09363(.A1(new_n9555_), .A2(new_n9113_), .Z(new_n9556_));
  INV_X1     g09364(.I(new_n9556_), .ZN(new_n9557_));
  AOI22_X1   g09365(.A1(new_n9552_), .A2(new_n9553_), .B1(new_n9545_), .B2(new_n9557_), .ZN(new_n9558_));
  NOR2_X1    g09366(.A1(new_n9142_), .A2(new_n8969_), .ZN(new_n9559_));
  OAI21_X1   g09367(.A1(\asqrt[22] ), .A2(new_n9559_), .B(new_n9149_), .ZN(new_n9560_));
  INV_X1     g09368(.I(new_n9560_), .ZN(new_n9561_));
  OAI21_X1   g09369(.A1(new_n9558_), .A2(new_n9382_), .B(new_n9561_), .ZN(new_n9562_));
  OAI21_X1   g09370(.A1(new_n9545_), .A2(\asqrt[62] ), .B(new_n9556_), .ZN(new_n9563_));
  NAND2_X1   g09371(.A1(new_n9545_), .A2(\asqrt[62] ), .ZN(new_n9564_));
  NAND3_X1   g09372(.A1(new_n9563_), .A2(new_n9564_), .A3(new_n9382_), .ZN(new_n9565_));
  NAND2_X1   g09373(.A1(new_n9233_), .A2(new_n8968_), .ZN(new_n9566_));
  XOR2_X1    g09374(.A1(new_n9221_), .A2(new_n8968_), .Z(new_n9567_));
  NAND3_X1   g09375(.A1(new_n9566_), .A2(\asqrt[63] ), .A3(new_n9567_), .ZN(new_n9568_));
  INV_X1     g09376(.I(new_n9230_), .ZN(new_n9569_));
  NAND4_X1   g09377(.A1(new_n9569_), .A2(new_n8969_), .A3(new_n9149_), .A4(new_n9157_), .ZN(new_n9570_));
  NAND2_X1   g09378(.A1(new_n9568_), .A2(new_n9570_), .ZN(new_n9571_));
  INV_X1     g09379(.I(new_n9571_), .ZN(new_n9572_));
  NAND4_X1   g09380(.A1(new_n9562_), .A2(new_n193_), .A3(new_n9565_), .A4(new_n9572_), .ZN(\asqrt[21] ));
  AOI21_X1   g09381(.A1(new_n9360_), .A2(new_n9377_), .B(\asqrt[21] ), .ZN(new_n9574_));
  XOR2_X1    g09382(.A1(new_n9574_), .A2(new_n9160_), .Z(new_n9575_));
  AOI21_X1   g09383(.A1(new_n9357_), .A2(new_n9375_), .B(\asqrt[21] ), .ZN(new_n9576_));
  XOR2_X1    g09384(.A1(new_n9576_), .A2(new_n9163_), .Z(new_n9577_));
  NAND2_X1   g09385(.A1(new_n9370_), .A2(new_n3195_), .ZN(new_n9578_));
  AOI21_X1   g09386(.A1(new_n9578_), .A2(new_n9356_), .B(\asqrt[21] ), .ZN(new_n9579_));
  XOR2_X1    g09387(.A1(new_n9579_), .A2(new_n9166_), .Z(new_n9580_));
  INV_X1     g09388(.I(new_n9580_), .ZN(new_n9581_));
  AOI21_X1   g09389(.A1(new_n9368_), .A2(new_n9353_), .B(\asqrt[21] ), .ZN(new_n9582_));
  XOR2_X1    g09390(.A1(new_n9582_), .A2(new_n9168_), .Z(new_n9583_));
  INV_X1     g09391(.I(new_n9583_), .ZN(new_n9584_));
  NAND2_X1   g09392(.A1(new_n9335_), .A2(new_n3681_), .ZN(new_n9585_));
  AOI21_X1   g09393(.A1(new_n9585_), .A2(new_n9367_), .B(\asqrt[21] ), .ZN(new_n9586_));
  XOR2_X1    g09394(.A1(new_n9586_), .A2(new_n9171_), .Z(new_n9587_));
  AOI21_X1   g09395(.A1(new_n9333_), .A2(new_n9350_), .B(\asqrt[21] ), .ZN(new_n9588_));
  XOR2_X1    g09396(.A1(new_n9588_), .A2(new_n9175_), .Z(new_n9589_));
  NAND2_X1   g09397(.A1(new_n9346_), .A2(new_n4196_), .ZN(new_n9590_));
  AOI21_X1   g09398(.A1(new_n9590_), .A2(new_n9332_), .B(\asqrt[21] ), .ZN(new_n9591_));
  XOR2_X1    g09399(.A1(new_n9591_), .A2(new_n9178_), .Z(new_n9592_));
  INV_X1     g09400(.I(new_n9592_), .ZN(new_n9593_));
  AOI21_X1   g09401(.A1(new_n9344_), .A2(new_n9329_), .B(\asqrt[21] ), .ZN(new_n9594_));
  XOR2_X1    g09402(.A1(new_n9594_), .A2(new_n9180_), .Z(new_n9595_));
  INV_X1     g09403(.I(new_n9595_), .ZN(new_n9596_));
  NAND2_X1   g09404(.A1(new_n9311_), .A2(new_n4751_), .ZN(new_n9597_));
  AOI21_X1   g09405(.A1(new_n9597_), .A2(new_n9343_), .B(\asqrt[21] ), .ZN(new_n9598_));
  XOR2_X1    g09406(.A1(new_n9598_), .A2(new_n9183_), .Z(new_n9599_));
  AOI21_X1   g09407(.A1(new_n9309_), .A2(new_n9326_), .B(\asqrt[21] ), .ZN(new_n9600_));
  XOR2_X1    g09408(.A1(new_n9600_), .A2(new_n9187_), .Z(new_n9601_));
  NAND2_X1   g09409(.A1(new_n9322_), .A2(new_n5336_), .ZN(new_n9602_));
  AOI21_X1   g09410(.A1(new_n9602_), .A2(new_n9308_), .B(\asqrt[21] ), .ZN(new_n9603_));
  XOR2_X1    g09411(.A1(new_n9603_), .A2(new_n9190_), .Z(new_n9604_));
  INV_X1     g09412(.I(new_n9604_), .ZN(new_n9605_));
  AOI21_X1   g09413(.A1(new_n9320_), .A2(new_n9305_), .B(\asqrt[21] ), .ZN(new_n9606_));
  XOR2_X1    g09414(.A1(new_n9606_), .A2(new_n9192_), .Z(new_n9607_));
  INV_X1     g09415(.I(new_n9607_), .ZN(new_n9608_));
  NAND2_X1   g09416(.A1(new_n9287_), .A2(new_n5947_), .ZN(new_n9609_));
  AOI21_X1   g09417(.A1(new_n9609_), .A2(new_n9319_), .B(\asqrt[21] ), .ZN(new_n9610_));
  XOR2_X1    g09418(.A1(new_n9610_), .A2(new_n9195_), .Z(new_n9611_));
  AOI21_X1   g09419(.A1(new_n9285_), .A2(new_n9302_), .B(\asqrt[21] ), .ZN(new_n9612_));
  XOR2_X1    g09420(.A1(new_n9612_), .A2(new_n9199_), .Z(new_n9613_));
  NAND2_X1   g09421(.A1(new_n9298_), .A2(new_n6636_), .ZN(new_n9614_));
  AOI21_X1   g09422(.A1(new_n9614_), .A2(new_n9284_), .B(\asqrt[21] ), .ZN(new_n9615_));
  XOR2_X1    g09423(.A1(new_n9615_), .A2(new_n9202_), .Z(new_n9616_));
  INV_X1     g09424(.I(new_n9616_), .ZN(new_n9617_));
  AOI21_X1   g09425(.A1(new_n9296_), .A2(new_n9281_), .B(\asqrt[21] ), .ZN(new_n9618_));
  XOR2_X1    g09426(.A1(new_n9618_), .A2(new_n9204_), .Z(new_n9619_));
  INV_X1     g09427(.I(new_n9619_), .ZN(new_n9620_));
  NAND2_X1   g09428(.A1(new_n9259_), .A2(new_n7331_), .ZN(new_n9621_));
  AOI21_X1   g09429(.A1(new_n9621_), .A2(new_n9295_), .B(\asqrt[21] ), .ZN(new_n9622_));
  XOR2_X1    g09430(.A1(new_n9622_), .A2(new_n9207_), .Z(new_n9623_));
  AOI21_X1   g09431(.A1(new_n9257_), .A2(new_n9278_), .B(\asqrt[21] ), .ZN(new_n9624_));
  XOR2_X1    g09432(.A1(new_n9624_), .A2(new_n9210_), .Z(new_n9625_));
  NAND2_X1   g09433(.A1(new_n9274_), .A2(new_n8077_), .ZN(new_n9626_));
  AOI21_X1   g09434(.A1(new_n9626_), .A2(new_n9256_), .B(\asqrt[21] ), .ZN(new_n9627_));
  XOR2_X1    g09435(.A1(new_n9627_), .A2(new_n9217_), .Z(new_n9628_));
  INV_X1     g09436(.I(new_n9628_), .ZN(new_n9629_));
  AOI21_X1   g09437(.A1(new_n9272_), .A2(new_n9253_), .B(\asqrt[21] ), .ZN(new_n9630_));
  XOR2_X1    g09438(.A1(new_n9630_), .A2(new_n9263_), .Z(new_n9631_));
  INV_X1     g09439(.I(new_n9631_), .ZN(new_n9632_));
  NAND2_X1   g09440(.A1(\asqrt[22] ), .A2(new_n9240_), .ZN(new_n9633_));
  NOR2_X1    g09441(.A1(new_n9248_), .A2(\a[44] ), .ZN(new_n9634_));
  AOI22_X1   g09442(.A1(new_n9633_), .A2(new_n9248_), .B1(\asqrt[22] ), .B2(new_n9634_), .ZN(new_n9635_));
  OAI21_X1   g09443(.A1(new_n9233_), .A2(new_n9240_), .B(new_n9267_), .ZN(new_n9636_));
  AOI21_X1   g09444(.A1(new_n9266_), .A2(new_n9636_), .B(\asqrt[21] ), .ZN(new_n9637_));
  XOR2_X1    g09445(.A1(new_n9637_), .A2(new_n9635_), .Z(new_n9638_));
  NAND3_X1   g09446(.A1(new_n9547_), .A2(new_n239_), .A3(new_n9540_), .ZN(new_n9639_));
  AOI21_X1   g09447(.A1(new_n9543_), .A2(new_n9639_), .B(new_n9548_), .ZN(new_n9640_));
  AOI21_X1   g09448(.A1(new_n9544_), .A2(new_n9539_), .B(\asqrt[62] ), .ZN(new_n9641_));
  NOR3_X1    g09449(.A1(new_n9551_), .A2(new_n201_), .A3(new_n9548_), .ZN(new_n9642_));
  OAI22_X1   g09450(.A1(new_n9642_), .A2(new_n9641_), .B1(new_n9640_), .B2(new_n9556_), .ZN(new_n9643_));
  AOI21_X1   g09451(.A1(new_n9643_), .A2(new_n9381_), .B(new_n9560_), .ZN(new_n9644_));
  AOI21_X1   g09452(.A1(new_n9640_), .A2(new_n201_), .B(new_n9557_), .ZN(new_n9645_));
  OAI21_X1   g09453(.A1(new_n9640_), .A2(new_n201_), .B(new_n9382_), .ZN(new_n9646_));
  NOR2_X1    g09454(.A1(new_n9645_), .A2(new_n9646_), .ZN(new_n9647_));
  NOR3_X1    g09455(.A1(new_n9644_), .A2(\asqrt[63] ), .A3(new_n9647_), .ZN(new_n9648_));
  NAND3_X1   g09456(.A1(new_n9568_), .A2(\asqrt[22] ), .A3(new_n9570_), .ZN(new_n9649_));
  INV_X1     g09457(.I(new_n9649_), .ZN(new_n9650_));
  NAND2_X1   g09458(.A1(new_n9648_), .A2(new_n9650_), .ZN(new_n9651_));
  NAND2_X1   g09459(.A1(\asqrt[21] ), .A2(new_n9237_), .ZN(new_n9652_));
  AOI21_X1   g09460(.A1(new_n9652_), .A2(new_n9651_), .B(\a[44] ), .ZN(new_n9653_));
  NAND2_X1   g09461(.A1(new_n9562_), .A2(new_n193_), .ZN(new_n9654_));
  NOR3_X1    g09462(.A1(new_n9654_), .A2(new_n9647_), .A3(new_n9649_), .ZN(new_n9655_));
  NOR4_X1    g09463(.A1(new_n9644_), .A2(\asqrt[63] ), .A3(new_n9647_), .A4(new_n9571_), .ZN(new_n9656_));
  NOR2_X1    g09464(.A1(new_n9656_), .A2(new_n9238_), .ZN(new_n9657_));
  NOR3_X1    g09465(.A1(new_n9657_), .A2(new_n9655_), .A3(new_n9240_), .ZN(new_n9658_));
  NOR2_X1    g09466(.A1(new_n9658_), .A2(new_n9653_), .ZN(new_n9659_));
  INV_X1     g09467(.I(\a[42] ), .ZN(new_n9660_));
  NOR2_X1    g09468(.A1(\a[40] ), .A2(\a[41] ), .ZN(new_n9661_));
  NOR3_X1    g09469(.A1(new_n9656_), .A2(new_n9660_), .A3(new_n9661_), .ZN(new_n9662_));
  INV_X1     g09470(.I(new_n9661_), .ZN(new_n9663_));
  AOI21_X1   g09471(.A1(new_n9656_), .A2(\a[42] ), .B(new_n9663_), .ZN(new_n9664_));
  OAI21_X1   g09472(.A1(new_n9662_), .A2(new_n9664_), .B(\asqrt[22] ), .ZN(new_n9665_));
  NAND2_X1   g09473(.A1(new_n9661_), .A2(new_n9660_), .ZN(new_n9666_));
  NAND3_X1   g09474(.A1(new_n9153_), .A2(new_n9155_), .A3(new_n9666_), .ZN(new_n9667_));
  NAND2_X1   g09475(.A1(new_n9226_), .A2(new_n9667_), .ZN(new_n9668_));
  INV_X1     g09476(.I(new_n9668_), .ZN(new_n9669_));
  NOR3_X1    g09477(.A1(new_n9656_), .A2(new_n9660_), .A3(new_n9669_), .ZN(new_n9670_));
  NOR3_X1    g09478(.A1(new_n9656_), .A2(\a[42] ), .A3(\a[43] ), .ZN(new_n9671_));
  INV_X1     g09479(.I(\a[43] ), .ZN(new_n9672_));
  AOI21_X1   g09480(.A1(\asqrt[21] ), .A2(new_n9660_), .B(new_n9672_), .ZN(new_n9673_));
  NOR3_X1    g09481(.A1(new_n9670_), .A2(new_n9671_), .A3(new_n9673_), .ZN(new_n9674_));
  NAND3_X1   g09482(.A1(new_n9674_), .A2(new_n9665_), .A3(new_n8849_), .ZN(new_n9675_));
  NAND2_X1   g09483(.A1(new_n9675_), .A2(new_n9659_), .ZN(new_n9676_));
  NAND3_X1   g09484(.A1(\asqrt[21] ), .A2(\a[42] ), .A3(new_n9663_), .ZN(new_n9677_));
  OAI21_X1   g09485(.A1(\asqrt[21] ), .A2(new_n9660_), .B(new_n9661_), .ZN(new_n9678_));
  AOI21_X1   g09486(.A1(new_n9678_), .A2(new_n9677_), .B(new_n9233_), .ZN(new_n9679_));
  NAND3_X1   g09487(.A1(\asqrt[21] ), .A2(\a[42] ), .A3(new_n9668_), .ZN(new_n9680_));
  NAND3_X1   g09488(.A1(\asqrt[21] ), .A2(new_n9660_), .A3(new_n9672_), .ZN(new_n9681_));
  OAI21_X1   g09489(.A1(new_n9656_), .A2(\a[42] ), .B(\a[43] ), .ZN(new_n9682_));
  NAND3_X1   g09490(.A1(new_n9680_), .A2(new_n9682_), .A3(new_n9681_), .ZN(new_n9683_));
  OAI21_X1   g09491(.A1(new_n9683_), .A2(new_n9679_), .B(\asqrt[23] ), .ZN(new_n9684_));
  NAND3_X1   g09492(.A1(new_n9676_), .A2(new_n8440_), .A3(new_n9684_), .ZN(new_n9685_));
  AOI21_X1   g09493(.A1(new_n9676_), .A2(new_n9684_), .B(new_n8440_), .ZN(new_n9686_));
  AOI21_X1   g09494(.A1(new_n9638_), .A2(new_n9685_), .B(new_n9686_), .ZN(new_n9687_));
  AOI21_X1   g09495(.A1(new_n9687_), .A2(new_n8077_), .B(new_n9632_), .ZN(new_n9688_));
  OR2_X2     g09496(.A1(new_n9658_), .A2(new_n9653_), .Z(new_n9689_));
  NOR3_X1    g09497(.A1(new_n9683_), .A2(new_n9679_), .A3(\asqrt[23] ), .ZN(new_n9690_));
  OAI21_X1   g09498(.A1(new_n9689_), .A2(new_n9690_), .B(new_n9684_), .ZN(new_n9691_));
  OAI21_X1   g09499(.A1(new_n9691_), .A2(\asqrt[24] ), .B(new_n9638_), .ZN(new_n9692_));
  NAND2_X1   g09500(.A1(new_n9691_), .A2(\asqrt[24] ), .ZN(new_n9693_));
  AOI21_X1   g09501(.A1(new_n9692_), .A2(new_n9693_), .B(new_n8077_), .ZN(new_n9694_));
  NOR3_X1    g09502(.A1(new_n9688_), .A2(\asqrt[26] ), .A3(new_n9694_), .ZN(new_n9695_));
  OAI21_X1   g09503(.A1(new_n9688_), .A2(new_n9694_), .B(\asqrt[26] ), .ZN(new_n9696_));
  OAI21_X1   g09504(.A1(new_n9629_), .A2(new_n9695_), .B(new_n9696_), .ZN(new_n9697_));
  OAI21_X1   g09505(.A1(new_n9697_), .A2(\asqrt[27] ), .B(new_n9625_), .ZN(new_n9698_));
  NAND3_X1   g09506(.A1(new_n9692_), .A2(new_n9693_), .A3(new_n8077_), .ZN(new_n9699_));
  AOI21_X1   g09507(.A1(new_n9631_), .A2(new_n9699_), .B(new_n9694_), .ZN(new_n9700_));
  AOI21_X1   g09508(.A1(new_n9700_), .A2(new_n7690_), .B(new_n9629_), .ZN(new_n9701_));
  NAND2_X1   g09509(.A1(new_n9699_), .A2(new_n9631_), .ZN(new_n9702_));
  INV_X1     g09510(.I(new_n9694_), .ZN(new_n9703_));
  AOI21_X1   g09511(.A1(new_n9702_), .A2(new_n9703_), .B(new_n7690_), .ZN(new_n9704_));
  OAI21_X1   g09512(.A1(new_n9701_), .A2(new_n9704_), .B(\asqrt[27] ), .ZN(new_n9705_));
  NAND3_X1   g09513(.A1(new_n9698_), .A2(new_n6966_), .A3(new_n9705_), .ZN(new_n9706_));
  AOI21_X1   g09514(.A1(new_n9698_), .A2(new_n9705_), .B(new_n6966_), .ZN(new_n9707_));
  AOI21_X1   g09515(.A1(new_n9623_), .A2(new_n9706_), .B(new_n9707_), .ZN(new_n9708_));
  AOI21_X1   g09516(.A1(new_n9708_), .A2(new_n6636_), .B(new_n9620_), .ZN(new_n9709_));
  INV_X1     g09517(.I(new_n9625_), .ZN(new_n9710_));
  NOR3_X1    g09518(.A1(new_n9701_), .A2(\asqrt[27] ), .A3(new_n9704_), .ZN(new_n9711_));
  OAI21_X1   g09519(.A1(new_n9710_), .A2(new_n9711_), .B(new_n9705_), .ZN(new_n9712_));
  OAI21_X1   g09520(.A1(new_n9712_), .A2(\asqrt[28] ), .B(new_n9623_), .ZN(new_n9713_));
  NAND2_X1   g09521(.A1(new_n9712_), .A2(\asqrt[28] ), .ZN(new_n9714_));
  AOI21_X1   g09522(.A1(new_n9713_), .A2(new_n9714_), .B(new_n6636_), .ZN(new_n9715_));
  NOR3_X1    g09523(.A1(new_n9709_), .A2(\asqrt[30] ), .A3(new_n9715_), .ZN(new_n9716_));
  OAI21_X1   g09524(.A1(new_n9709_), .A2(new_n9715_), .B(\asqrt[30] ), .ZN(new_n9717_));
  OAI21_X1   g09525(.A1(new_n9617_), .A2(new_n9716_), .B(new_n9717_), .ZN(new_n9718_));
  OAI21_X1   g09526(.A1(new_n9718_), .A2(\asqrt[31] ), .B(new_n9613_), .ZN(new_n9719_));
  NAND3_X1   g09527(.A1(new_n9713_), .A2(new_n9714_), .A3(new_n6636_), .ZN(new_n9720_));
  AOI21_X1   g09528(.A1(new_n9619_), .A2(new_n9720_), .B(new_n9715_), .ZN(new_n9721_));
  AOI21_X1   g09529(.A1(new_n9721_), .A2(new_n6275_), .B(new_n9617_), .ZN(new_n9722_));
  NAND2_X1   g09530(.A1(new_n9720_), .A2(new_n9619_), .ZN(new_n9723_));
  INV_X1     g09531(.I(new_n9715_), .ZN(new_n9724_));
  AOI21_X1   g09532(.A1(new_n9723_), .A2(new_n9724_), .B(new_n6275_), .ZN(new_n9725_));
  OAI21_X1   g09533(.A1(new_n9722_), .A2(new_n9725_), .B(\asqrt[31] ), .ZN(new_n9726_));
  NAND3_X1   g09534(.A1(new_n9719_), .A2(new_n5643_), .A3(new_n9726_), .ZN(new_n9727_));
  AOI21_X1   g09535(.A1(new_n9719_), .A2(new_n9726_), .B(new_n5643_), .ZN(new_n9728_));
  AOI21_X1   g09536(.A1(new_n9611_), .A2(new_n9727_), .B(new_n9728_), .ZN(new_n9729_));
  AOI21_X1   g09537(.A1(new_n9729_), .A2(new_n5336_), .B(new_n9608_), .ZN(new_n9730_));
  INV_X1     g09538(.I(new_n9613_), .ZN(new_n9731_));
  NOR3_X1    g09539(.A1(new_n9722_), .A2(\asqrt[31] ), .A3(new_n9725_), .ZN(new_n9732_));
  OAI21_X1   g09540(.A1(new_n9731_), .A2(new_n9732_), .B(new_n9726_), .ZN(new_n9733_));
  OAI21_X1   g09541(.A1(new_n9733_), .A2(\asqrt[32] ), .B(new_n9611_), .ZN(new_n9734_));
  NAND2_X1   g09542(.A1(new_n9733_), .A2(\asqrt[32] ), .ZN(new_n9735_));
  AOI21_X1   g09543(.A1(new_n9734_), .A2(new_n9735_), .B(new_n5336_), .ZN(new_n9736_));
  NOR3_X1    g09544(.A1(new_n9730_), .A2(\asqrt[34] ), .A3(new_n9736_), .ZN(new_n9737_));
  OAI21_X1   g09545(.A1(new_n9730_), .A2(new_n9736_), .B(\asqrt[34] ), .ZN(new_n9738_));
  OAI21_X1   g09546(.A1(new_n9605_), .A2(new_n9737_), .B(new_n9738_), .ZN(new_n9739_));
  OAI21_X1   g09547(.A1(new_n9739_), .A2(\asqrt[35] ), .B(new_n9601_), .ZN(new_n9740_));
  NAND3_X1   g09548(.A1(new_n9734_), .A2(new_n9735_), .A3(new_n5336_), .ZN(new_n9741_));
  AOI21_X1   g09549(.A1(new_n9607_), .A2(new_n9741_), .B(new_n9736_), .ZN(new_n9742_));
  AOI21_X1   g09550(.A1(new_n9742_), .A2(new_n5029_), .B(new_n9605_), .ZN(new_n9743_));
  NAND2_X1   g09551(.A1(new_n9741_), .A2(new_n9607_), .ZN(new_n9744_));
  INV_X1     g09552(.I(new_n9736_), .ZN(new_n9745_));
  AOI21_X1   g09553(.A1(new_n9744_), .A2(new_n9745_), .B(new_n5029_), .ZN(new_n9746_));
  OAI21_X1   g09554(.A1(new_n9743_), .A2(new_n9746_), .B(\asqrt[35] ), .ZN(new_n9747_));
  NAND3_X1   g09555(.A1(new_n9740_), .A2(new_n4461_), .A3(new_n9747_), .ZN(new_n9748_));
  AOI21_X1   g09556(.A1(new_n9740_), .A2(new_n9747_), .B(new_n4461_), .ZN(new_n9749_));
  AOI21_X1   g09557(.A1(new_n9599_), .A2(new_n9748_), .B(new_n9749_), .ZN(new_n9750_));
  AOI21_X1   g09558(.A1(new_n9750_), .A2(new_n4196_), .B(new_n9596_), .ZN(new_n9751_));
  INV_X1     g09559(.I(new_n9601_), .ZN(new_n9752_));
  NOR3_X1    g09560(.A1(new_n9743_), .A2(\asqrt[35] ), .A3(new_n9746_), .ZN(new_n9753_));
  OAI21_X1   g09561(.A1(new_n9752_), .A2(new_n9753_), .B(new_n9747_), .ZN(new_n9754_));
  OAI21_X1   g09562(.A1(new_n9754_), .A2(\asqrt[36] ), .B(new_n9599_), .ZN(new_n9755_));
  NAND2_X1   g09563(.A1(new_n9754_), .A2(\asqrt[36] ), .ZN(new_n9756_));
  AOI21_X1   g09564(.A1(new_n9755_), .A2(new_n9756_), .B(new_n4196_), .ZN(new_n9757_));
  NOR3_X1    g09565(.A1(new_n9751_), .A2(\asqrt[38] ), .A3(new_n9757_), .ZN(new_n9758_));
  OAI21_X1   g09566(.A1(new_n9751_), .A2(new_n9757_), .B(\asqrt[38] ), .ZN(new_n9759_));
  OAI21_X1   g09567(.A1(new_n9593_), .A2(new_n9758_), .B(new_n9759_), .ZN(new_n9760_));
  OAI21_X1   g09568(.A1(new_n9760_), .A2(\asqrt[39] ), .B(new_n9589_), .ZN(new_n9761_));
  NAND3_X1   g09569(.A1(new_n9755_), .A2(new_n9756_), .A3(new_n4196_), .ZN(new_n9762_));
  AOI21_X1   g09570(.A1(new_n9595_), .A2(new_n9762_), .B(new_n9757_), .ZN(new_n9763_));
  AOI21_X1   g09571(.A1(new_n9763_), .A2(new_n3925_), .B(new_n9593_), .ZN(new_n9764_));
  NAND2_X1   g09572(.A1(new_n9762_), .A2(new_n9595_), .ZN(new_n9765_));
  INV_X1     g09573(.I(new_n9757_), .ZN(new_n9766_));
  AOI21_X1   g09574(.A1(new_n9765_), .A2(new_n9766_), .B(new_n3925_), .ZN(new_n9767_));
  OAI21_X1   g09575(.A1(new_n9764_), .A2(new_n9767_), .B(\asqrt[39] ), .ZN(new_n9768_));
  NAND3_X1   g09576(.A1(new_n9761_), .A2(new_n3427_), .A3(new_n9768_), .ZN(new_n9769_));
  AOI21_X1   g09577(.A1(new_n9761_), .A2(new_n9768_), .B(new_n3427_), .ZN(new_n9770_));
  AOI21_X1   g09578(.A1(new_n9587_), .A2(new_n9769_), .B(new_n9770_), .ZN(new_n9771_));
  AOI21_X1   g09579(.A1(new_n9771_), .A2(new_n3195_), .B(new_n9584_), .ZN(new_n9772_));
  INV_X1     g09580(.I(new_n9589_), .ZN(new_n9773_));
  NOR3_X1    g09581(.A1(new_n9764_), .A2(\asqrt[39] ), .A3(new_n9767_), .ZN(new_n9774_));
  OAI21_X1   g09582(.A1(new_n9773_), .A2(new_n9774_), .B(new_n9768_), .ZN(new_n9775_));
  OAI21_X1   g09583(.A1(new_n9775_), .A2(\asqrt[40] ), .B(new_n9587_), .ZN(new_n9776_));
  NAND2_X1   g09584(.A1(new_n9775_), .A2(\asqrt[40] ), .ZN(new_n9777_));
  AOI21_X1   g09585(.A1(new_n9776_), .A2(new_n9777_), .B(new_n3195_), .ZN(new_n9778_));
  NOR3_X1    g09586(.A1(new_n9772_), .A2(\asqrt[42] ), .A3(new_n9778_), .ZN(new_n9779_));
  OAI21_X1   g09587(.A1(new_n9772_), .A2(new_n9778_), .B(\asqrt[42] ), .ZN(new_n9780_));
  OAI21_X1   g09588(.A1(new_n9581_), .A2(new_n9779_), .B(new_n9780_), .ZN(new_n9781_));
  OAI21_X1   g09589(.A1(new_n9781_), .A2(\asqrt[43] ), .B(new_n9577_), .ZN(new_n9782_));
  NAND3_X1   g09590(.A1(new_n9776_), .A2(new_n9777_), .A3(new_n3195_), .ZN(new_n9783_));
  AOI21_X1   g09591(.A1(new_n9583_), .A2(new_n9783_), .B(new_n9778_), .ZN(new_n9784_));
  AOI21_X1   g09592(.A1(new_n9784_), .A2(new_n2960_), .B(new_n9581_), .ZN(new_n9785_));
  NAND2_X1   g09593(.A1(new_n9783_), .A2(new_n9583_), .ZN(new_n9786_));
  INV_X1     g09594(.I(new_n9778_), .ZN(new_n9787_));
  AOI21_X1   g09595(.A1(new_n9786_), .A2(new_n9787_), .B(new_n2960_), .ZN(new_n9788_));
  OAI21_X1   g09596(.A1(new_n9785_), .A2(new_n9788_), .B(\asqrt[43] ), .ZN(new_n9789_));
  NAND3_X1   g09597(.A1(new_n9782_), .A2(new_n2531_), .A3(new_n9789_), .ZN(new_n9790_));
  INV_X1     g09598(.I(new_n9577_), .ZN(new_n9791_));
  NOR3_X1    g09599(.A1(new_n9785_), .A2(\asqrt[43] ), .A3(new_n9788_), .ZN(new_n9792_));
  OAI21_X1   g09600(.A1(new_n9791_), .A2(new_n9792_), .B(new_n9789_), .ZN(new_n9793_));
  NAND2_X1   g09601(.A1(new_n9793_), .A2(\asqrt[44] ), .ZN(new_n9794_));
  NOR2_X1    g09602(.A1(new_n9545_), .A2(\asqrt[62] ), .ZN(new_n9795_));
  INV_X1     g09603(.I(new_n9564_), .ZN(new_n9796_));
  NOR2_X1    g09604(.A1(new_n9796_), .A2(new_n9795_), .ZN(new_n9797_));
  XOR2_X1    g09605(.A1(new_n9555_), .A2(new_n9113_), .Z(new_n9798_));
  OAI21_X1   g09606(.A1(\asqrt[21] ), .A2(new_n9797_), .B(new_n9798_), .ZN(new_n9799_));
  INV_X1     g09607(.I(new_n9799_), .ZN(new_n9800_));
  NAND2_X1   g09608(.A1(new_n9513_), .A2(new_n337_), .ZN(new_n9801_));
  AOI21_X1   g09609(.A1(new_n9801_), .A2(new_n9537_), .B(\asqrt[21] ), .ZN(new_n9802_));
  XOR2_X1    g09610(.A1(new_n9802_), .A2(new_n9387_), .Z(new_n9803_));
  INV_X1     g09611(.I(new_n9803_), .ZN(new_n9804_));
  AOI21_X1   g09612(.A1(new_n9511_), .A2(new_n9528_), .B(\asqrt[21] ), .ZN(new_n9805_));
  XOR2_X1    g09613(.A1(new_n9805_), .A2(new_n9391_), .Z(new_n9806_));
  INV_X1     g09614(.I(new_n9806_), .ZN(new_n9807_));
  NAND2_X1   g09615(.A1(new_n9524_), .A2(new_n531_), .ZN(new_n9808_));
  AOI21_X1   g09616(.A1(new_n9808_), .A2(new_n9510_), .B(\asqrt[21] ), .ZN(new_n9809_));
  XOR2_X1    g09617(.A1(new_n9809_), .A2(new_n9394_), .Z(new_n9810_));
  INV_X1     g09618(.I(new_n9810_), .ZN(new_n9811_));
  AOI21_X1   g09619(.A1(new_n9522_), .A2(new_n9507_), .B(\asqrt[21] ), .ZN(new_n9812_));
  XOR2_X1    g09620(.A1(new_n9812_), .A2(new_n9396_), .Z(new_n9813_));
  NAND2_X1   g09621(.A1(new_n9489_), .A2(new_n744_), .ZN(new_n9814_));
  AOI21_X1   g09622(.A1(new_n9814_), .A2(new_n9521_), .B(\asqrt[21] ), .ZN(new_n9815_));
  XOR2_X1    g09623(.A1(new_n9815_), .A2(new_n9399_), .Z(new_n9816_));
  AOI21_X1   g09624(.A1(new_n9487_), .A2(new_n9504_), .B(\asqrt[21] ), .ZN(new_n9817_));
  XOR2_X1    g09625(.A1(new_n9817_), .A2(new_n9403_), .Z(new_n9818_));
  INV_X1     g09626(.I(new_n9818_), .ZN(new_n9819_));
  NAND2_X1   g09627(.A1(new_n9500_), .A2(new_n1006_), .ZN(new_n9820_));
  AOI21_X1   g09628(.A1(new_n9820_), .A2(new_n9486_), .B(\asqrt[21] ), .ZN(new_n9821_));
  XOR2_X1    g09629(.A1(new_n9821_), .A2(new_n9406_), .Z(new_n9822_));
  INV_X1     g09630(.I(new_n9822_), .ZN(new_n9823_));
  AOI21_X1   g09631(.A1(new_n9498_), .A2(new_n9483_), .B(\asqrt[21] ), .ZN(new_n9824_));
  XOR2_X1    g09632(.A1(new_n9824_), .A2(new_n9408_), .Z(new_n9825_));
  NAND2_X1   g09633(.A1(new_n9465_), .A2(new_n1305_), .ZN(new_n9826_));
  AOI21_X1   g09634(.A1(new_n9826_), .A2(new_n9497_), .B(\asqrt[21] ), .ZN(new_n9827_));
  XOR2_X1    g09635(.A1(new_n9827_), .A2(new_n9411_), .Z(new_n9828_));
  AOI21_X1   g09636(.A1(new_n9463_), .A2(new_n9480_), .B(\asqrt[21] ), .ZN(new_n9829_));
  XOR2_X1    g09637(.A1(new_n9829_), .A2(new_n9415_), .Z(new_n9830_));
  INV_X1     g09638(.I(new_n9830_), .ZN(new_n9831_));
  NAND2_X1   g09639(.A1(new_n9476_), .A2(new_n1632_), .ZN(new_n9832_));
  AOI21_X1   g09640(.A1(new_n9832_), .A2(new_n9462_), .B(\asqrt[21] ), .ZN(new_n9833_));
  XOR2_X1    g09641(.A1(new_n9833_), .A2(new_n9418_), .Z(new_n9834_));
  INV_X1     g09642(.I(new_n9834_), .ZN(new_n9835_));
  AOI21_X1   g09643(.A1(new_n9474_), .A2(new_n9459_), .B(\asqrt[21] ), .ZN(new_n9836_));
  XOR2_X1    g09644(.A1(new_n9836_), .A2(new_n9420_), .Z(new_n9837_));
  NAND2_X1   g09645(.A1(new_n9445_), .A2(new_n1953_), .ZN(new_n9838_));
  AOI21_X1   g09646(.A1(new_n9838_), .A2(new_n9473_), .B(\asqrt[21] ), .ZN(new_n9839_));
  XOR2_X1    g09647(.A1(new_n9839_), .A2(new_n9423_), .Z(new_n9840_));
  AOI21_X1   g09648(.A1(new_n9443_), .A2(new_n9456_), .B(\asqrt[21] ), .ZN(new_n9841_));
  XOR2_X1    g09649(.A1(new_n9841_), .A2(new_n9427_), .Z(new_n9842_));
  INV_X1     g09650(.I(new_n9842_), .ZN(new_n9843_));
  NAND2_X1   g09651(.A1(new_n9452_), .A2(new_n2332_), .ZN(new_n9844_));
  AOI21_X1   g09652(.A1(new_n9844_), .A2(new_n9442_), .B(\asqrt[21] ), .ZN(new_n9845_));
  XOR2_X1    g09653(.A1(new_n9845_), .A2(new_n9430_), .Z(new_n9846_));
  INV_X1     g09654(.I(new_n9846_), .ZN(new_n9847_));
  AOI21_X1   g09655(.A1(new_n9450_), .A2(new_n9439_), .B(\asqrt[21] ), .ZN(new_n9848_));
  XOR2_X1    g09656(.A1(new_n9848_), .A2(new_n9432_), .Z(new_n9849_));
  OAI21_X1   g09657(.A1(new_n9793_), .A2(\asqrt[44] ), .B(new_n9575_), .ZN(new_n9850_));
  NAND3_X1   g09658(.A1(new_n9850_), .A2(new_n9794_), .A3(new_n2332_), .ZN(new_n9851_));
  AOI21_X1   g09659(.A1(new_n9850_), .A2(new_n9794_), .B(new_n2332_), .ZN(new_n9852_));
  AOI21_X1   g09660(.A1(new_n9849_), .A2(new_n9851_), .B(new_n9852_), .ZN(new_n9853_));
  AOI21_X1   g09661(.A1(new_n9853_), .A2(new_n2134_), .B(new_n9847_), .ZN(new_n9854_));
  NAND2_X1   g09662(.A1(new_n9851_), .A2(new_n9849_), .ZN(new_n9855_));
  INV_X1     g09663(.I(new_n9852_), .ZN(new_n9856_));
  AOI21_X1   g09664(.A1(new_n9855_), .A2(new_n9856_), .B(new_n2134_), .ZN(new_n9857_));
  NOR3_X1    g09665(.A1(new_n9854_), .A2(\asqrt[47] ), .A3(new_n9857_), .ZN(new_n9858_));
  OAI21_X1   g09666(.A1(new_n9854_), .A2(new_n9857_), .B(\asqrt[47] ), .ZN(new_n9859_));
  OAI21_X1   g09667(.A1(new_n9843_), .A2(new_n9858_), .B(new_n9859_), .ZN(new_n9860_));
  OAI21_X1   g09668(.A1(new_n9860_), .A2(\asqrt[48] ), .B(new_n9840_), .ZN(new_n9861_));
  NAND2_X1   g09669(.A1(new_n9860_), .A2(\asqrt[48] ), .ZN(new_n9862_));
  NAND3_X1   g09670(.A1(new_n9861_), .A2(new_n9862_), .A3(new_n1632_), .ZN(new_n9863_));
  AOI21_X1   g09671(.A1(new_n9861_), .A2(new_n9862_), .B(new_n1632_), .ZN(new_n9864_));
  AOI21_X1   g09672(.A1(new_n9837_), .A2(new_n9863_), .B(new_n9864_), .ZN(new_n9865_));
  AOI21_X1   g09673(.A1(new_n9865_), .A2(new_n1463_), .B(new_n9835_), .ZN(new_n9866_));
  NAND2_X1   g09674(.A1(new_n9863_), .A2(new_n9837_), .ZN(new_n9867_));
  INV_X1     g09675(.I(new_n9864_), .ZN(new_n9868_));
  AOI21_X1   g09676(.A1(new_n9867_), .A2(new_n9868_), .B(new_n1463_), .ZN(new_n9869_));
  NOR3_X1    g09677(.A1(new_n9866_), .A2(\asqrt[51] ), .A3(new_n9869_), .ZN(new_n9870_));
  OAI21_X1   g09678(.A1(new_n9866_), .A2(new_n9869_), .B(\asqrt[51] ), .ZN(new_n9871_));
  OAI21_X1   g09679(.A1(new_n9831_), .A2(new_n9870_), .B(new_n9871_), .ZN(new_n9872_));
  OAI21_X1   g09680(.A1(new_n9872_), .A2(\asqrt[52] ), .B(new_n9828_), .ZN(new_n9873_));
  NAND2_X1   g09681(.A1(new_n9872_), .A2(\asqrt[52] ), .ZN(new_n9874_));
  NAND3_X1   g09682(.A1(new_n9873_), .A2(new_n9874_), .A3(new_n1006_), .ZN(new_n9875_));
  AOI21_X1   g09683(.A1(new_n9873_), .A2(new_n9874_), .B(new_n1006_), .ZN(new_n9876_));
  AOI21_X1   g09684(.A1(new_n9825_), .A2(new_n9875_), .B(new_n9876_), .ZN(new_n9877_));
  AOI21_X1   g09685(.A1(new_n9877_), .A2(new_n860_), .B(new_n9823_), .ZN(new_n9878_));
  NAND2_X1   g09686(.A1(new_n9875_), .A2(new_n9825_), .ZN(new_n9879_));
  INV_X1     g09687(.I(new_n9876_), .ZN(new_n9880_));
  AOI21_X1   g09688(.A1(new_n9879_), .A2(new_n9880_), .B(new_n860_), .ZN(new_n9881_));
  NOR3_X1    g09689(.A1(new_n9878_), .A2(\asqrt[55] ), .A3(new_n9881_), .ZN(new_n9882_));
  OAI21_X1   g09690(.A1(new_n9878_), .A2(new_n9881_), .B(\asqrt[55] ), .ZN(new_n9883_));
  OAI21_X1   g09691(.A1(new_n9819_), .A2(new_n9882_), .B(new_n9883_), .ZN(new_n9884_));
  OAI21_X1   g09692(.A1(new_n9884_), .A2(\asqrt[56] ), .B(new_n9816_), .ZN(new_n9885_));
  NAND2_X1   g09693(.A1(new_n9884_), .A2(\asqrt[56] ), .ZN(new_n9886_));
  NAND3_X1   g09694(.A1(new_n9885_), .A2(new_n9886_), .A3(new_n531_), .ZN(new_n9887_));
  AOI21_X1   g09695(.A1(new_n9885_), .A2(new_n9886_), .B(new_n531_), .ZN(new_n9888_));
  AOI21_X1   g09696(.A1(new_n9813_), .A2(new_n9887_), .B(new_n9888_), .ZN(new_n9889_));
  AOI21_X1   g09697(.A1(new_n9889_), .A2(new_n423_), .B(new_n9811_), .ZN(new_n9890_));
  NAND2_X1   g09698(.A1(new_n9887_), .A2(new_n9813_), .ZN(new_n9891_));
  INV_X1     g09699(.I(new_n9888_), .ZN(new_n9892_));
  AOI21_X1   g09700(.A1(new_n9891_), .A2(new_n9892_), .B(new_n423_), .ZN(new_n9893_));
  NOR3_X1    g09701(.A1(new_n9890_), .A2(\asqrt[59] ), .A3(new_n9893_), .ZN(new_n9894_));
  NOR2_X1    g09702(.A1(new_n9894_), .A2(new_n9807_), .ZN(new_n9895_));
  OAI21_X1   g09703(.A1(new_n9890_), .A2(new_n9893_), .B(\asqrt[59] ), .ZN(new_n9896_));
  INV_X1     g09704(.I(new_n9896_), .ZN(new_n9897_));
  NOR2_X1    g09705(.A1(new_n9895_), .A2(new_n9897_), .ZN(new_n9898_));
  AOI21_X1   g09706(.A1(new_n9898_), .A2(new_n266_), .B(new_n9804_), .ZN(new_n9899_));
  INV_X1     g09707(.I(new_n9813_), .ZN(new_n9900_));
  INV_X1     g09708(.I(new_n9825_), .ZN(new_n9901_));
  INV_X1     g09709(.I(new_n9837_), .ZN(new_n9902_));
  INV_X1     g09710(.I(new_n9849_), .ZN(new_n9903_));
  AOI21_X1   g09711(.A1(new_n9782_), .A2(new_n9789_), .B(new_n2531_), .ZN(new_n9904_));
  AOI21_X1   g09712(.A1(new_n9575_), .A2(new_n9790_), .B(new_n9904_), .ZN(new_n9905_));
  AOI21_X1   g09713(.A1(new_n9905_), .A2(new_n2332_), .B(new_n9903_), .ZN(new_n9906_));
  NOR3_X1    g09714(.A1(new_n9906_), .A2(\asqrt[46] ), .A3(new_n9852_), .ZN(new_n9907_));
  OAI21_X1   g09715(.A1(new_n9906_), .A2(new_n9852_), .B(\asqrt[46] ), .ZN(new_n9908_));
  OAI21_X1   g09716(.A1(new_n9847_), .A2(new_n9907_), .B(new_n9908_), .ZN(new_n9909_));
  OAI21_X1   g09717(.A1(new_n9909_), .A2(\asqrt[47] ), .B(new_n9842_), .ZN(new_n9910_));
  NAND3_X1   g09718(.A1(new_n9910_), .A2(new_n1778_), .A3(new_n9859_), .ZN(new_n9911_));
  AOI21_X1   g09719(.A1(new_n9910_), .A2(new_n9859_), .B(new_n1778_), .ZN(new_n9912_));
  AOI21_X1   g09720(.A1(new_n9840_), .A2(new_n9911_), .B(new_n9912_), .ZN(new_n9913_));
  AOI21_X1   g09721(.A1(new_n9913_), .A2(new_n1632_), .B(new_n9902_), .ZN(new_n9914_));
  NOR3_X1    g09722(.A1(new_n9914_), .A2(\asqrt[50] ), .A3(new_n9864_), .ZN(new_n9915_));
  OAI21_X1   g09723(.A1(new_n9914_), .A2(new_n9864_), .B(\asqrt[50] ), .ZN(new_n9916_));
  OAI21_X1   g09724(.A1(new_n9835_), .A2(new_n9915_), .B(new_n9916_), .ZN(new_n9917_));
  OAI21_X1   g09725(.A1(new_n9917_), .A2(\asqrt[51] ), .B(new_n9830_), .ZN(new_n9918_));
  NAND3_X1   g09726(.A1(new_n9918_), .A2(new_n1150_), .A3(new_n9871_), .ZN(new_n9919_));
  AOI21_X1   g09727(.A1(new_n9918_), .A2(new_n9871_), .B(new_n1150_), .ZN(new_n9920_));
  AOI21_X1   g09728(.A1(new_n9828_), .A2(new_n9919_), .B(new_n9920_), .ZN(new_n9921_));
  AOI21_X1   g09729(.A1(new_n9921_), .A2(new_n1006_), .B(new_n9901_), .ZN(new_n9922_));
  NOR3_X1    g09730(.A1(new_n9922_), .A2(\asqrt[54] ), .A3(new_n9876_), .ZN(new_n9923_));
  OAI21_X1   g09731(.A1(new_n9922_), .A2(new_n9876_), .B(\asqrt[54] ), .ZN(new_n9924_));
  OAI21_X1   g09732(.A1(new_n9823_), .A2(new_n9923_), .B(new_n9924_), .ZN(new_n9925_));
  OAI21_X1   g09733(.A1(new_n9925_), .A2(\asqrt[55] ), .B(new_n9818_), .ZN(new_n9926_));
  NAND3_X1   g09734(.A1(new_n9926_), .A2(new_n634_), .A3(new_n9883_), .ZN(new_n9927_));
  AOI21_X1   g09735(.A1(new_n9926_), .A2(new_n9883_), .B(new_n634_), .ZN(new_n9928_));
  AOI21_X1   g09736(.A1(new_n9816_), .A2(new_n9927_), .B(new_n9928_), .ZN(new_n9929_));
  AOI21_X1   g09737(.A1(new_n9929_), .A2(new_n531_), .B(new_n9900_), .ZN(new_n9930_));
  NOR3_X1    g09738(.A1(new_n9930_), .A2(\asqrt[58] ), .A3(new_n9888_), .ZN(new_n9931_));
  OAI21_X1   g09739(.A1(new_n9930_), .A2(new_n9888_), .B(\asqrt[58] ), .ZN(new_n9932_));
  OAI21_X1   g09740(.A1(new_n9811_), .A2(new_n9931_), .B(new_n9932_), .ZN(new_n9933_));
  OAI21_X1   g09741(.A1(new_n9933_), .A2(\asqrt[59] ), .B(new_n9806_), .ZN(new_n9934_));
  AOI21_X1   g09742(.A1(new_n9934_), .A2(new_n9896_), .B(new_n266_), .ZN(new_n9935_));
  OAI21_X1   g09743(.A1(new_n9899_), .A2(new_n9935_), .B(\asqrt[61] ), .ZN(new_n9936_));
  AOI21_X1   g09744(.A1(new_n9546_), .A2(new_n9540_), .B(\asqrt[21] ), .ZN(new_n9937_));
  XOR2_X1    g09745(.A1(new_n9937_), .A2(new_n9384_), .Z(new_n9938_));
  OAI21_X1   g09746(.A1(new_n9807_), .A2(new_n9894_), .B(new_n9896_), .ZN(new_n9939_));
  OAI21_X1   g09747(.A1(new_n9939_), .A2(\asqrt[60] ), .B(new_n9803_), .ZN(new_n9940_));
  OAI21_X1   g09748(.A1(new_n9895_), .A2(new_n9897_), .B(\asqrt[60] ), .ZN(new_n9941_));
  NAND3_X1   g09749(.A1(new_n9940_), .A2(new_n239_), .A3(new_n9941_), .ZN(new_n9942_));
  NAND2_X1   g09750(.A1(new_n9942_), .A2(new_n9938_), .ZN(new_n9943_));
  NAND2_X1   g09751(.A1(new_n9943_), .A2(new_n9936_), .ZN(new_n9944_));
  AOI21_X1   g09752(.A1(new_n9940_), .A2(new_n9941_), .B(new_n239_), .ZN(new_n9945_));
  NAND3_X1   g09753(.A1(new_n9934_), .A2(new_n266_), .A3(new_n9896_), .ZN(new_n9946_));
  AOI21_X1   g09754(.A1(new_n9803_), .A2(new_n9946_), .B(new_n9935_), .ZN(new_n9947_));
  INV_X1     g09755(.I(new_n9938_), .ZN(new_n9948_));
  AOI21_X1   g09756(.A1(new_n9947_), .A2(new_n239_), .B(new_n9948_), .ZN(new_n9949_));
  OAI21_X1   g09757(.A1(new_n9949_), .A2(new_n9945_), .B(new_n201_), .ZN(new_n9950_));
  NAND3_X1   g09758(.A1(new_n9943_), .A2(\asqrt[62] ), .A3(new_n9936_), .ZN(new_n9951_));
  AOI21_X1   g09759(.A1(new_n9539_), .A2(new_n9639_), .B(\asqrt[21] ), .ZN(new_n9952_));
  XOR2_X1    g09760(.A1(new_n9952_), .A2(new_n9543_), .Z(new_n9953_));
  INV_X1     g09761(.I(new_n9953_), .ZN(new_n9954_));
  AOI22_X1   g09762(.A1(new_n9950_), .A2(new_n9951_), .B1(new_n9944_), .B2(new_n9954_), .ZN(new_n9955_));
  NOR2_X1    g09763(.A1(new_n9558_), .A2(new_n9382_), .ZN(new_n9956_));
  OAI21_X1   g09764(.A1(\asqrt[21] ), .A2(new_n9956_), .B(new_n9565_), .ZN(new_n9957_));
  INV_X1     g09765(.I(new_n9957_), .ZN(new_n9958_));
  OAI21_X1   g09766(.A1(new_n9955_), .A2(new_n9800_), .B(new_n9958_), .ZN(new_n9959_));
  OAI21_X1   g09767(.A1(new_n9944_), .A2(\asqrt[62] ), .B(new_n9953_), .ZN(new_n9960_));
  NAND2_X1   g09768(.A1(new_n9944_), .A2(\asqrt[62] ), .ZN(new_n9961_));
  NAND3_X1   g09769(.A1(new_n9960_), .A2(new_n9961_), .A3(new_n9800_), .ZN(new_n9962_));
  NAND2_X1   g09770(.A1(new_n9656_), .A2(new_n9381_), .ZN(new_n9963_));
  XOR2_X1    g09771(.A1(new_n9558_), .A2(new_n9382_), .Z(new_n9964_));
  NAND3_X1   g09772(.A1(new_n9963_), .A2(\asqrt[63] ), .A3(new_n9964_), .ZN(new_n9965_));
  INV_X1     g09773(.I(new_n9654_), .ZN(new_n9966_));
  NAND4_X1   g09774(.A1(new_n9966_), .A2(new_n9382_), .A3(new_n9565_), .A4(new_n9572_), .ZN(new_n9967_));
  NAND2_X1   g09775(.A1(new_n9965_), .A2(new_n9967_), .ZN(new_n9968_));
  INV_X1     g09776(.I(new_n9968_), .ZN(new_n9969_));
  NAND4_X1   g09777(.A1(new_n9959_), .A2(new_n193_), .A3(new_n9962_), .A4(new_n9969_), .ZN(\asqrt[20] ));
  AOI21_X1   g09778(.A1(new_n9790_), .A2(new_n9794_), .B(\asqrt[20] ), .ZN(new_n9971_));
  XOR2_X1    g09779(.A1(new_n9971_), .A2(new_n9575_), .Z(new_n9972_));
  XOR2_X1    g09780(.A1(new_n9781_), .A2(\asqrt[43] ), .Z(new_n9973_));
  NOR2_X1    g09781(.A1(\asqrt[20] ), .A2(new_n9973_), .ZN(new_n9974_));
  XOR2_X1    g09782(.A1(new_n9974_), .A2(new_n9577_), .Z(new_n9975_));
  NOR2_X1    g09783(.A1(new_n9779_), .A2(new_n9788_), .ZN(new_n9976_));
  NOR2_X1    g09784(.A1(\asqrt[20] ), .A2(new_n9976_), .ZN(new_n9977_));
  XOR2_X1    g09785(.A1(new_n9977_), .A2(new_n9580_), .Z(new_n9978_));
  AOI21_X1   g09786(.A1(new_n9783_), .A2(new_n9787_), .B(\asqrt[20] ), .ZN(new_n9979_));
  XOR2_X1    g09787(.A1(new_n9979_), .A2(new_n9583_), .Z(new_n9980_));
  INV_X1     g09788(.I(new_n9980_), .ZN(new_n9981_));
  AOI21_X1   g09789(.A1(new_n9769_), .A2(new_n9777_), .B(\asqrt[20] ), .ZN(new_n9982_));
  XOR2_X1    g09790(.A1(new_n9982_), .A2(new_n9587_), .Z(new_n9983_));
  INV_X1     g09791(.I(new_n9983_), .ZN(new_n9984_));
  XOR2_X1    g09792(.A1(new_n9760_), .A2(\asqrt[39] ), .Z(new_n9985_));
  NOR2_X1    g09793(.A1(\asqrt[20] ), .A2(new_n9985_), .ZN(new_n9986_));
  XOR2_X1    g09794(.A1(new_n9986_), .A2(new_n9589_), .Z(new_n9987_));
  NOR2_X1    g09795(.A1(new_n9758_), .A2(new_n9767_), .ZN(new_n9988_));
  NOR2_X1    g09796(.A1(\asqrt[20] ), .A2(new_n9988_), .ZN(new_n9989_));
  XOR2_X1    g09797(.A1(new_n9989_), .A2(new_n9592_), .Z(new_n9990_));
  AOI21_X1   g09798(.A1(new_n9762_), .A2(new_n9766_), .B(\asqrt[20] ), .ZN(new_n9991_));
  XOR2_X1    g09799(.A1(new_n9991_), .A2(new_n9595_), .Z(new_n9992_));
  INV_X1     g09800(.I(new_n9992_), .ZN(new_n9993_));
  AOI21_X1   g09801(.A1(new_n9748_), .A2(new_n9756_), .B(\asqrt[20] ), .ZN(new_n9994_));
  XOR2_X1    g09802(.A1(new_n9994_), .A2(new_n9599_), .Z(new_n9995_));
  INV_X1     g09803(.I(new_n9995_), .ZN(new_n9996_));
  XOR2_X1    g09804(.A1(new_n9739_), .A2(\asqrt[35] ), .Z(new_n9997_));
  NOR2_X1    g09805(.A1(\asqrt[20] ), .A2(new_n9997_), .ZN(new_n9998_));
  XOR2_X1    g09806(.A1(new_n9998_), .A2(new_n9601_), .Z(new_n9999_));
  NOR2_X1    g09807(.A1(new_n9737_), .A2(new_n9746_), .ZN(new_n10000_));
  NOR2_X1    g09808(.A1(\asqrt[20] ), .A2(new_n10000_), .ZN(new_n10001_));
  XOR2_X1    g09809(.A1(new_n10001_), .A2(new_n9604_), .Z(new_n10002_));
  AOI21_X1   g09810(.A1(new_n9741_), .A2(new_n9745_), .B(\asqrt[20] ), .ZN(new_n10003_));
  XOR2_X1    g09811(.A1(new_n10003_), .A2(new_n9607_), .Z(new_n10004_));
  INV_X1     g09812(.I(new_n10004_), .ZN(new_n10005_));
  AOI21_X1   g09813(.A1(new_n9727_), .A2(new_n9735_), .B(\asqrt[20] ), .ZN(new_n10006_));
  XOR2_X1    g09814(.A1(new_n10006_), .A2(new_n9611_), .Z(new_n10007_));
  INV_X1     g09815(.I(new_n10007_), .ZN(new_n10008_));
  XOR2_X1    g09816(.A1(new_n9718_), .A2(\asqrt[31] ), .Z(new_n10009_));
  NOR2_X1    g09817(.A1(\asqrt[20] ), .A2(new_n10009_), .ZN(new_n10010_));
  XOR2_X1    g09818(.A1(new_n10010_), .A2(new_n9613_), .Z(new_n10011_));
  NOR2_X1    g09819(.A1(new_n9716_), .A2(new_n9725_), .ZN(new_n10012_));
  NOR2_X1    g09820(.A1(\asqrt[20] ), .A2(new_n10012_), .ZN(new_n10013_));
  XOR2_X1    g09821(.A1(new_n10013_), .A2(new_n9616_), .Z(new_n10014_));
  AOI21_X1   g09822(.A1(new_n9720_), .A2(new_n9724_), .B(\asqrt[20] ), .ZN(new_n10015_));
  XOR2_X1    g09823(.A1(new_n10015_), .A2(new_n9619_), .Z(new_n10016_));
  INV_X1     g09824(.I(new_n10016_), .ZN(new_n10017_));
  AOI21_X1   g09825(.A1(new_n9706_), .A2(new_n9714_), .B(\asqrt[20] ), .ZN(new_n10018_));
  XOR2_X1    g09826(.A1(new_n10018_), .A2(new_n9623_), .Z(new_n10019_));
  INV_X1     g09827(.I(new_n10019_), .ZN(new_n10020_));
  XOR2_X1    g09828(.A1(new_n9697_), .A2(\asqrt[27] ), .Z(new_n10021_));
  NOR2_X1    g09829(.A1(\asqrt[20] ), .A2(new_n10021_), .ZN(new_n10022_));
  XOR2_X1    g09830(.A1(new_n10022_), .A2(new_n9625_), .Z(new_n10023_));
  NOR2_X1    g09831(.A1(new_n9695_), .A2(new_n9704_), .ZN(new_n10024_));
  NOR2_X1    g09832(.A1(\asqrt[20] ), .A2(new_n10024_), .ZN(new_n10025_));
  XOR2_X1    g09833(.A1(new_n10025_), .A2(new_n9628_), .Z(new_n10026_));
  AOI21_X1   g09834(.A1(new_n9699_), .A2(new_n9703_), .B(\asqrt[20] ), .ZN(new_n10027_));
  XOR2_X1    g09835(.A1(new_n10027_), .A2(new_n9631_), .Z(new_n10028_));
  INV_X1     g09836(.I(new_n10028_), .ZN(new_n10029_));
  AOI21_X1   g09837(.A1(new_n9685_), .A2(new_n9693_), .B(\asqrt[20] ), .ZN(new_n10030_));
  XOR2_X1    g09838(.A1(new_n10030_), .A2(new_n9638_), .Z(new_n10031_));
  INV_X1     g09839(.I(new_n10031_), .ZN(new_n10032_));
  AOI21_X1   g09840(.A1(new_n9675_), .A2(new_n9684_), .B(\asqrt[20] ), .ZN(new_n10033_));
  XOR2_X1    g09841(.A1(new_n10033_), .A2(new_n9659_), .Z(new_n10034_));
  NAND2_X1   g09842(.A1(\asqrt[21] ), .A2(new_n9660_), .ZN(new_n10035_));
  NOR2_X1    g09843(.A1(new_n9672_), .A2(\a[42] ), .ZN(new_n10036_));
  AOI22_X1   g09844(.A1(new_n10035_), .A2(new_n9672_), .B1(\asqrt[21] ), .B2(new_n10036_), .ZN(new_n10037_));
  OAI21_X1   g09845(.A1(new_n9656_), .A2(new_n9660_), .B(new_n9669_), .ZN(new_n10038_));
  AOI21_X1   g09846(.A1(new_n9665_), .A2(new_n10038_), .B(\asqrt[20] ), .ZN(new_n10039_));
  XOR2_X1    g09847(.A1(new_n10039_), .A2(new_n10037_), .Z(new_n10040_));
  NAND2_X1   g09848(.A1(new_n9959_), .A2(new_n193_), .ZN(new_n10041_));
  NOR2_X1    g09849(.A1(new_n9949_), .A2(new_n9945_), .ZN(new_n10042_));
  AOI21_X1   g09850(.A1(new_n10042_), .A2(new_n201_), .B(new_n9954_), .ZN(new_n10043_));
  OAI21_X1   g09851(.A1(new_n10042_), .A2(new_n201_), .B(new_n9800_), .ZN(new_n10044_));
  NOR2_X1    g09852(.A1(new_n10043_), .A2(new_n10044_), .ZN(new_n10045_));
  NAND3_X1   g09853(.A1(new_n9965_), .A2(\asqrt[21] ), .A3(new_n9967_), .ZN(new_n10046_));
  NOR3_X1    g09854(.A1(new_n10041_), .A2(new_n10045_), .A3(new_n10046_), .ZN(new_n10047_));
  AOI21_X1   g09855(.A1(new_n9943_), .A2(new_n9936_), .B(\asqrt[62] ), .ZN(new_n10048_));
  NOR3_X1    g09856(.A1(new_n9949_), .A2(new_n201_), .A3(new_n9945_), .ZN(new_n10049_));
  OAI22_X1   g09857(.A1(new_n10049_), .A2(new_n10048_), .B1(new_n10042_), .B2(new_n9953_), .ZN(new_n10050_));
  AOI21_X1   g09858(.A1(new_n10050_), .A2(new_n9799_), .B(new_n9957_), .ZN(new_n10051_));
  NOR4_X1    g09859(.A1(new_n10051_), .A2(\asqrt[63] ), .A3(new_n10045_), .A4(new_n9968_), .ZN(new_n10052_));
  NOR2_X1    g09860(.A1(new_n10052_), .A2(new_n9663_), .ZN(new_n10053_));
  OAI21_X1   g09861(.A1(new_n10053_), .A2(new_n10047_), .B(new_n9660_), .ZN(new_n10054_));
  NOR3_X1    g09862(.A1(new_n10051_), .A2(\asqrt[63] ), .A3(new_n10045_), .ZN(new_n10055_));
  NAND4_X1   g09863(.A1(new_n10055_), .A2(\asqrt[21] ), .A3(new_n9965_), .A4(new_n9967_), .ZN(new_n10056_));
  NAND2_X1   g09864(.A1(\asqrt[20] ), .A2(new_n9661_), .ZN(new_n10057_));
  NAND3_X1   g09865(.A1(new_n10056_), .A2(new_n10057_), .A3(\a[42] ), .ZN(new_n10058_));
  NAND2_X1   g09866(.A1(new_n10058_), .A2(new_n10054_), .ZN(new_n10059_));
  NOR2_X1    g09867(.A1(\a[38] ), .A2(\a[39] ), .ZN(new_n10060_));
  INV_X1     g09868(.I(new_n10060_), .ZN(new_n10061_));
  NAND3_X1   g09869(.A1(\asqrt[20] ), .A2(\a[40] ), .A3(new_n10061_), .ZN(new_n10062_));
  INV_X1     g09870(.I(\a[40] ), .ZN(new_n10063_));
  OAI21_X1   g09871(.A1(\asqrt[20] ), .A2(new_n10063_), .B(new_n10060_), .ZN(new_n10064_));
  AOI21_X1   g09872(.A1(new_n10064_), .A2(new_n10062_), .B(new_n9656_), .ZN(new_n10065_));
  NAND2_X1   g09873(.A1(new_n10060_), .A2(new_n10063_), .ZN(new_n10066_));
  NAND3_X1   g09874(.A1(new_n9568_), .A2(new_n9570_), .A3(new_n10066_), .ZN(new_n10067_));
  NAND2_X1   g09875(.A1(new_n9648_), .A2(new_n10067_), .ZN(new_n10068_));
  NAND3_X1   g09876(.A1(\asqrt[20] ), .A2(\a[40] ), .A3(new_n10068_), .ZN(new_n10069_));
  INV_X1     g09877(.I(\a[41] ), .ZN(new_n10070_));
  NAND3_X1   g09878(.A1(\asqrt[20] ), .A2(new_n10063_), .A3(new_n10070_), .ZN(new_n10071_));
  OAI21_X1   g09879(.A1(new_n10052_), .A2(\a[40] ), .B(\a[41] ), .ZN(new_n10072_));
  NAND3_X1   g09880(.A1(new_n10072_), .A2(new_n10069_), .A3(new_n10071_), .ZN(new_n10073_));
  NOR3_X1    g09881(.A1(new_n10073_), .A2(new_n10065_), .A3(\asqrt[22] ), .ZN(new_n10074_));
  OAI21_X1   g09882(.A1(new_n10073_), .A2(new_n10065_), .B(\asqrt[22] ), .ZN(new_n10075_));
  OAI21_X1   g09883(.A1(new_n10059_), .A2(new_n10074_), .B(new_n10075_), .ZN(new_n10076_));
  OAI21_X1   g09884(.A1(new_n10076_), .A2(\asqrt[23] ), .B(new_n10040_), .ZN(new_n10077_));
  NAND2_X1   g09885(.A1(new_n10076_), .A2(\asqrt[23] ), .ZN(new_n10078_));
  NAND3_X1   g09886(.A1(new_n10077_), .A2(new_n10078_), .A3(new_n8440_), .ZN(new_n10079_));
  AOI21_X1   g09887(.A1(new_n10077_), .A2(new_n10078_), .B(new_n8440_), .ZN(new_n10080_));
  AOI21_X1   g09888(.A1(new_n10034_), .A2(new_n10079_), .B(new_n10080_), .ZN(new_n10081_));
  AOI21_X1   g09889(.A1(new_n10081_), .A2(new_n8077_), .B(new_n10032_), .ZN(new_n10082_));
  NAND2_X1   g09890(.A1(new_n10079_), .A2(new_n10034_), .ZN(new_n10083_));
  INV_X1     g09891(.I(new_n10040_), .ZN(new_n10084_));
  INV_X1     g09892(.I(new_n10059_), .ZN(new_n10085_));
  NOR3_X1    g09893(.A1(new_n10052_), .A2(new_n10063_), .A3(new_n10060_), .ZN(new_n10086_));
  AOI21_X1   g09894(.A1(new_n10052_), .A2(\a[40] ), .B(new_n10061_), .ZN(new_n10087_));
  OAI21_X1   g09895(.A1(new_n10086_), .A2(new_n10087_), .B(\asqrt[21] ), .ZN(new_n10088_));
  INV_X1     g09896(.I(new_n10068_), .ZN(new_n10089_));
  NOR3_X1    g09897(.A1(new_n10052_), .A2(new_n10063_), .A3(new_n10089_), .ZN(new_n10090_));
  NOR3_X1    g09898(.A1(new_n10052_), .A2(\a[40] ), .A3(\a[41] ), .ZN(new_n10091_));
  AOI21_X1   g09899(.A1(\asqrt[20] ), .A2(new_n10063_), .B(new_n10070_), .ZN(new_n10092_));
  NOR3_X1    g09900(.A1(new_n10090_), .A2(new_n10091_), .A3(new_n10092_), .ZN(new_n10093_));
  NAND3_X1   g09901(.A1(new_n10088_), .A2(new_n10093_), .A3(new_n9233_), .ZN(new_n10094_));
  AOI21_X1   g09902(.A1(new_n10088_), .A2(new_n10093_), .B(new_n9233_), .ZN(new_n10095_));
  AOI21_X1   g09903(.A1(new_n10085_), .A2(new_n10094_), .B(new_n10095_), .ZN(new_n10096_));
  AOI21_X1   g09904(.A1(new_n10096_), .A2(new_n8849_), .B(new_n10084_), .ZN(new_n10097_));
  NAND2_X1   g09905(.A1(new_n10085_), .A2(new_n10094_), .ZN(new_n10098_));
  AOI21_X1   g09906(.A1(new_n10098_), .A2(new_n10075_), .B(new_n8849_), .ZN(new_n10099_));
  OAI21_X1   g09907(.A1(new_n10097_), .A2(new_n10099_), .B(\asqrt[24] ), .ZN(new_n10100_));
  AOI21_X1   g09908(.A1(new_n10083_), .A2(new_n10100_), .B(new_n8077_), .ZN(new_n10101_));
  NOR3_X1    g09909(.A1(new_n10082_), .A2(\asqrt[26] ), .A3(new_n10101_), .ZN(new_n10102_));
  OAI21_X1   g09910(.A1(new_n10082_), .A2(new_n10101_), .B(\asqrt[26] ), .ZN(new_n10103_));
  OAI21_X1   g09911(.A1(new_n10029_), .A2(new_n10102_), .B(new_n10103_), .ZN(new_n10104_));
  OAI21_X1   g09912(.A1(new_n10104_), .A2(\asqrt[27] ), .B(new_n10026_), .ZN(new_n10105_));
  NAND2_X1   g09913(.A1(new_n10104_), .A2(\asqrt[27] ), .ZN(new_n10106_));
  NAND3_X1   g09914(.A1(new_n10105_), .A2(new_n10106_), .A3(new_n6966_), .ZN(new_n10107_));
  AOI21_X1   g09915(.A1(new_n10105_), .A2(new_n10106_), .B(new_n6966_), .ZN(new_n10108_));
  AOI21_X1   g09916(.A1(new_n10023_), .A2(new_n10107_), .B(new_n10108_), .ZN(new_n10109_));
  AOI21_X1   g09917(.A1(new_n10109_), .A2(new_n6636_), .B(new_n10020_), .ZN(new_n10110_));
  NAND2_X1   g09918(.A1(new_n10107_), .A2(new_n10023_), .ZN(new_n10111_));
  INV_X1     g09919(.I(new_n10026_), .ZN(new_n10112_));
  INV_X1     g09920(.I(new_n10034_), .ZN(new_n10113_));
  NOR3_X1    g09921(.A1(new_n10097_), .A2(\asqrt[24] ), .A3(new_n10099_), .ZN(new_n10114_));
  OAI21_X1   g09922(.A1(new_n10113_), .A2(new_n10114_), .B(new_n10100_), .ZN(new_n10115_));
  OAI21_X1   g09923(.A1(new_n10115_), .A2(\asqrt[25] ), .B(new_n10031_), .ZN(new_n10116_));
  NAND2_X1   g09924(.A1(new_n10115_), .A2(\asqrt[25] ), .ZN(new_n10117_));
  NAND3_X1   g09925(.A1(new_n10116_), .A2(new_n10117_), .A3(new_n7690_), .ZN(new_n10118_));
  AOI21_X1   g09926(.A1(new_n10116_), .A2(new_n10117_), .B(new_n7690_), .ZN(new_n10119_));
  AOI21_X1   g09927(.A1(new_n10028_), .A2(new_n10118_), .B(new_n10119_), .ZN(new_n10120_));
  AOI21_X1   g09928(.A1(new_n10120_), .A2(new_n7331_), .B(new_n10112_), .ZN(new_n10121_));
  NAND2_X1   g09929(.A1(new_n10118_), .A2(new_n10028_), .ZN(new_n10122_));
  AOI21_X1   g09930(.A1(new_n10122_), .A2(new_n10103_), .B(new_n7331_), .ZN(new_n10123_));
  OAI21_X1   g09931(.A1(new_n10121_), .A2(new_n10123_), .B(\asqrt[28] ), .ZN(new_n10124_));
  AOI21_X1   g09932(.A1(new_n10111_), .A2(new_n10124_), .B(new_n6636_), .ZN(new_n10125_));
  NOR3_X1    g09933(.A1(new_n10110_), .A2(\asqrt[30] ), .A3(new_n10125_), .ZN(new_n10126_));
  OAI21_X1   g09934(.A1(new_n10110_), .A2(new_n10125_), .B(\asqrt[30] ), .ZN(new_n10127_));
  OAI21_X1   g09935(.A1(new_n10017_), .A2(new_n10126_), .B(new_n10127_), .ZN(new_n10128_));
  OAI21_X1   g09936(.A1(new_n10128_), .A2(\asqrt[31] ), .B(new_n10014_), .ZN(new_n10129_));
  NAND2_X1   g09937(.A1(new_n10128_), .A2(\asqrt[31] ), .ZN(new_n10130_));
  NAND3_X1   g09938(.A1(new_n10129_), .A2(new_n10130_), .A3(new_n5643_), .ZN(new_n10131_));
  AOI21_X1   g09939(.A1(new_n10129_), .A2(new_n10130_), .B(new_n5643_), .ZN(new_n10132_));
  AOI21_X1   g09940(.A1(new_n10011_), .A2(new_n10131_), .B(new_n10132_), .ZN(new_n10133_));
  AOI21_X1   g09941(.A1(new_n10133_), .A2(new_n5336_), .B(new_n10008_), .ZN(new_n10134_));
  NAND2_X1   g09942(.A1(new_n10131_), .A2(new_n10011_), .ZN(new_n10135_));
  INV_X1     g09943(.I(new_n10014_), .ZN(new_n10136_));
  INV_X1     g09944(.I(new_n10023_), .ZN(new_n10137_));
  NOR3_X1    g09945(.A1(new_n10121_), .A2(\asqrt[28] ), .A3(new_n10123_), .ZN(new_n10138_));
  OAI21_X1   g09946(.A1(new_n10137_), .A2(new_n10138_), .B(new_n10124_), .ZN(new_n10139_));
  OAI21_X1   g09947(.A1(new_n10139_), .A2(\asqrt[29] ), .B(new_n10019_), .ZN(new_n10140_));
  NAND2_X1   g09948(.A1(new_n10139_), .A2(\asqrt[29] ), .ZN(new_n10141_));
  NAND3_X1   g09949(.A1(new_n10140_), .A2(new_n10141_), .A3(new_n6275_), .ZN(new_n10142_));
  AOI21_X1   g09950(.A1(new_n10140_), .A2(new_n10141_), .B(new_n6275_), .ZN(new_n10143_));
  AOI21_X1   g09951(.A1(new_n10016_), .A2(new_n10142_), .B(new_n10143_), .ZN(new_n10144_));
  AOI21_X1   g09952(.A1(new_n10144_), .A2(new_n5947_), .B(new_n10136_), .ZN(new_n10145_));
  NAND2_X1   g09953(.A1(new_n10142_), .A2(new_n10016_), .ZN(new_n10146_));
  AOI21_X1   g09954(.A1(new_n10146_), .A2(new_n10127_), .B(new_n5947_), .ZN(new_n10147_));
  OAI21_X1   g09955(.A1(new_n10145_), .A2(new_n10147_), .B(\asqrt[32] ), .ZN(new_n10148_));
  AOI21_X1   g09956(.A1(new_n10135_), .A2(new_n10148_), .B(new_n5336_), .ZN(new_n10149_));
  NOR3_X1    g09957(.A1(new_n10134_), .A2(\asqrt[34] ), .A3(new_n10149_), .ZN(new_n10150_));
  OAI21_X1   g09958(.A1(new_n10134_), .A2(new_n10149_), .B(\asqrt[34] ), .ZN(new_n10151_));
  OAI21_X1   g09959(.A1(new_n10005_), .A2(new_n10150_), .B(new_n10151_), .ZN(new_n10152_));
  OAI21_X1   g09960(.A1(new_n10152_), .A2(\asqrt[35] ), .B(new_n10002_), .ZN(new_n10153_));
  NAND2_X1   g09961(.A1(new_n10152_), .A2(\asqrt[35] ), .ZN(new_n10154_));
  NAND3_X1   g09962(.A1(new_n10153_), .A2(new_n10154_), .A3(new_n4461_), .ZN(new_n10155_));
  AOI21_X1   g09963(.A1(new_n10153_), .A2(new_n10154_), .B(new_n4461_), .ZN(new_n10156_));
  AOI21_X1   g09964(.A1(new_n9999_), .A2(new_n10155_), .B(new_n10156_), .ZN(new_n10157_));
  AOI21_X1   g09965(.A1(new_n10157_), .A2(new_n4196_), .B(new_n9996_), .ZN(new_n10158_));
  NAND2_X1   g09966(.A1(new_n10155_), .A2(new_n9999_), .ZN(new_n10159_));
  INV_X1     g09967(.I(new_n10002_), .ZN(new_n10160_));
  INV_X1     g09968(.I(new_n10011_), .ZN(new_n10161_));
  NOR3_X1    g09969(.A1(new_n10145_), .A2(\asqrt[32] ), .A3(new_n10147_), .ZN(new_n10162_));
  OAI21_X1   g09970(.A1(new_n10161_), .A2(new_n10162_), .B(new_n10148_), .ZN(new_n10163_));
  OAI21_X1   g09971(.A1(new_n10163_), .A2(\asqrt[33] ), .B(new_n10007_), .ZN(new_n10164_));
  NAND2_X1   g09972(.A1(new_n10163_), .A2(\asqrt[33] ), .ZN(new_n10165_));
  NAND3_X1   g09973(.A1(new_n10164_), .A2(new_n10165_), .A3(new_n5029_), .ZN(new_n10166_));
  AOI21_X1   g09974(.A1(new_n10164_), .A2(new_n10165_), .B(new_n5029_), .ZN(new_n10167_));
  AOI21_X1   g09975(.A1(new_n10004_), .A2(new_n10166_), .B(new_n10167_), .ZN(new_n10168_));
  AOI21_X1   g09976(.A1(new_n10168_), .A2(new_n4751_), .B(new_n10160_), .ZN(new_n10169_));
  NAND2_X1   g09977(.A1(new_n10166_), .A2(new_n10004_), .ZN(new_n10170_));
  AOI21_X1   g09978(.A1(new_n10170_), .A2(new_n10151_), .B(new_n4751_), .ZN(new_n10171_));
  OAI21_X1   g09979(.A1(new_n10169_), .A2(new_n10171_), .B(\asqrt[36] ), .ZN(new_n10172_));
  AOI21_X1   g09980(.A1(new_n10159_), .A2(new_n10172_), .B(new_n4196_), .ZN(new_n10173_));
  NOR3_X1    g09981(.A1(new_n10158_), .A2(\asqrt[38] ), .A3(new_n10173_), .ZN(new_n10174_));
  OAI21_X1   g09982(.A1(new_n10158_), .A2(new_n10173_), .B(\asqrt[38] ), .ZN(new_n10175_));
  OAI21_X1   g09983(.A1(new_n9993_), .A2(new_n10174_), .B(new_n10175_), .ZN(new_n10176_));
  OAI21_X1   g09984(.A1(new_n10176_), .A2(\asqrt[39] ), .B(new_n9990_), .ZN(new_n10177_));
  NAND2_X1   g09985(.A1(new_n10176_), .A2(\asqrt[39] ), .ZN(new_n10178_));
  NAND3_X1   g09986(.A1(new_n10177_), .A2(new_n10178_), .A3(new_n3427_), .ZN(new_n10179_));
  AOI21_X1   g09987(.A1(new_n10177_), .A2(new_n10178_), .B(new_n3427_), .ZN(new_n10180_));
  AOI21_X1   g09988(.A1(new_n9987_), .A2(new_n10179_), .B(new_n10180_), .ZN(new_n10181_));
  AOI21_X1   g09989(.A1(new_n10181_), .A2(new_n3195_), .B(new_n9984_), .ZN(new_n10182_));
  NAND2_X1   g09990(.A1(new_n10179_), .A2(new_n9987_), .ZN(new_n10183_));
  INV_X1     g09991(.I(new_n9990_), .ZN(new_n10184_));
  INV_X1     g09992(.I(new_n9999_), .ZN(new_n10185_));
  NOR3_X1    g09993(.A1(new_n10169_), .A2(\asqrt[36] ), .A3(new_n10171_), .ZN(new_n10186_));
  OAI21_X1   g09994(.A1(new_n10185_), .A2(new_n10186_), .B(new_n10172_), .ZN(new_n10187_));
  OAI21_X1   g09995(.A1(new_n10187_), .A2(\asqrt[37] ), .B(new_n9995_), .ZN(new_n10188_));
  NAND2_X1   g09996(.A1(new_n10187_), .A2(\asqrt[37] ), .ZN(new_n10189_));
  NAND3_X1   g09997(.A1(new_n10188_), .A2(new_n10189_), .A3(new_n3925_), .ZN(new_n10190_));
  AOI21_X1   g09998(.A1(new_n10188_), .A2(new_n10189_), .B(new_n3925_), .ZN(new_n10191_));
  AOI21_X1   g09999(.A1(new_n9992_), .A2(new_n10190_), .B(new_n10191_), .ZN(new_n10192_));
  AOI21_X1   g10000(.A1(new_n10192_), .A2(new_n3681_), .B(new_n10184_), .ZN(new_n10193_));
  NAND2_X1   g10001(.A1(new_n10190_), .A2(new_n9992_), .ZN(new_n10194_));
  AOI21_X1   g10002(.A1(new_n10194_), .A2(new_n10175_), .B(new_n3681_), .ZN(new_n10195_));
  OAI21_X1   g10003(.A1(new_n10193_), .A2(new_n10195_), .B(\asqrt[40] ), .ZN(new_n10196_));
  AOI21_X1   g10004(.A1(new_n10183_), .A2(new_n10196_), .B(new_n3195_), .ZN(new_n10197_));
  NOR3_X1    g10005(.A1(new_n10182_), .A2(\asqrt[42] ), .A3(new_n10197_), .ZN(new_n10198_));
  OAI21_X1   g10006(.A1(new_n10182_), .A2(new_n10197_), .B(\asqrt[42] ), .ZN(new_n10199_));
  OAI21_X1   g10007(.A1(new_n9981_), .A2(new_n10198_), .B(new_n10199_), .ZN(new_n10200_));
  OAI21_X1   g10008(.A1(new_n10200_), .A2(\asqrt[43] ), .B(new_n9978_), .ZN(new_n10201_));
  NAND2_X1   g10009(.A1(new_n10200_), .A2(\asqrt[43] ), .ZN(new_n10202_));
  NAND3_X1   g10010(.A1(new_n10201_), .A2(new_n10202_), .A3(new_n2531_), .ZN(new_n10203_));
  AOI21_X1   g10011(.A1(new_n10201_), .A2(new_n10202_), .B(new_n2531_), .ZN(new_n10204_));
  AOI21_X1   g10012(.A1(new_n9975_), .A2(new_n10203_), .B(new_n10204_), .ZN(new_n10205_));
  NAND2_X1   g10013(.A1(new_n10205_), .A2(new_n2332_), .ZN(new_n10206_));
  INV_X1     g10014(.I(new_n9975_), .ZN(new_n10207_));
  INV_X1     g10015(.I(new_n9978_), .ZN(new_n10208_));
  INV_X1     g10016(.I(new_n9987_), .ZN(new_n10209_));
  NOR3_X1    g10017(.A1(new_n10193_), .A2(\asqrt[40] ), .A3(new_n10195_), .ZN(new_n10210_));
  OAI21_X1   g10018(.A1(new_n10209_), .A2(new_n10210_), .B(new_n10196_), .ZN(new_n10211_));
  OAI21_X1   g10019(.A1(new_n10211_), .A2(\asqrt[41] ), .B(new_n9983_), .ZN(new_n10212_));
  NAND2_X1   g10020(.A1(new_n10211_), .A2(\asqrt[41] ), .ZN(new_n10213_));
  NAND3_X1   g10021(.A1(new_n10212_), .A2(new_n10213_), .A3(new_n2960_), .ZN(new_n10214_));
  AOI21_X1   g10022(.A1(new_n10212_), .A2(new_n10213_), .B(new_n2960_), .ZN(new_n10215_));
  AOI21_X1   g10023(.A1(new_n9980_), .A2(new_n10214_), .B(new_n10215_), .ZN(new_n10216_));
  AOI21_X1   g10024(.A1(new_n10216_), .A2(new_n2749_), .B(new_n10208_), .ZN(new_n10217_));
  NAND2_X1   g10025(.A1(new_n10214_), .A2(new_n9980_), .ZN(new_n10218_));
  AOI21_X1   g10026(.A1(new_n10218_), .A2(new_n10199_), .B(new_n2749_), .ZN(new_n10219_));
  NOR3_X1    g10027(.A1(new_n10217_), .A2(\asqrt[44] ), .A3(new_n10219_), .ZN(new_n10220_));
  OAI21_X1   g10028(.A1(new_n10217_), .A2(new_n10219_), .B(\asqrt[44] ), .ZN(new_n10221_));
  OAI21_X1   g10029(.A1(new_n10207_), .A2(new_n10220_), .B(new_n10221_), .ZN(new_n10222_));
  NAND2_X1   g10030(.A1(new_n10222_), .A2(\asqrt[45] ), .ZN(new_n10223_));
  NOR2_X1    g10031(.A1(new_n9944_), .A2(\asqrt[62] ), .ZN(new_n10224_));
  INV_X1     g10032(.I(new_n9961_), .ZN(new_n10225_));
  NOR2_X1    g10033(.A1(new_n10225_), .A2(new_n10224_), .ZN(new_n10226_));
  XOR2_X1    g10034(.A1(new_n9952_), .A2(new_n9543_), .Z(new_n10227_));
  OAI21_X1   g10035(.A1(\asqrt[20] ), .A2(new_n10226_), .B(new_n10227_), .ZN(new_n10228_));
  INV_X1     g10036(.I(new_n10228_), .ZN(new_n10229_));
  NOR2_X1    g10037(.A1(new_n9897_), .A2(new_n9894_), .ZN(new_n10230_));
  NOR2_X1    g10038(.A1(\asqrt[20] ), .A2(new_n10230_), .ZN(new_n10231_));
  XOR2_X1    g10039(.A1(new_n10231_), .A2(new_n9806_), .Z(new_n10232_));
  INV_X1     g10040(.I(new_n10232_), .ZN(new_n10233_));
  NOR2_X1    g10041(.A1(new_n9931_), .A2(new_n9893_), .ZN(new_n10234_));
  NOR2_X1    g10042(.A1(\asqrt[20] ), .A2(new_n10234_), .ZN(new_n10235_));
  XOR2_X1    g10043(.A1(new_n10235_), .A2(new_n9810_), .Z(new_n10236_));
  AOI21_X1   g10044(.A1(new_n9887_), .A2(new_n9892_), .B(\asqrt[20] ), .ZN(new_n10237_));
  XOR2_X1    g10045(.A1(new_n10237_), .A2(new_n9813_), .Z(new_n10238_));
  AOI21_X1   g10046(.A1(new_n9927_), .A2(new_n9886_), .B(\asqrt[20] ), .ZN(new_n10239_));
  XOR2_X1    g10047(.A1(new_n10239_), .A2(new_n9816_), .Z(new_n10240_));
  INV_X1     g10048(.I(new_n9883_), .ZN(new_n10241_));
  NOR2_X1    g10049(.A1(new_n10241_), .A2(new_n9882_), .ZN(new_n10242_));
  NOR2_X1    g10050(.A1(\asqrt[20] ), .A2(new_n10242_), .ZN(new_n10243_));
  XOR2_X1    g10051(.A1(new_n10243_), .A2(new_n9818_), .Z(new_n10244_));
  INV_X1     g10052(.I(new_n10244_), .ZN(new_n10245_));
  NOR2_X1    g10053(.A1(new_n9923_), .A2(new_n9881_), .ZN(new_n10246_));
  NOR2_X1    g10054(.A1(\asqrt[20] ), .A2(new_n10246_), .ZN(new_n10247_));
  XOR2_X1    g10055(.A1(new_n10247_), .A2(new_n9822_), .Z(new_n10248_));
  INV_X1     g10056(.I(new_n10248_), .ZN(new_n10249_));
  AOI21_X1   g10057(.A1(new_n9875_), .A2(new_n9880_), .B(\asqrt[20] ), .ZN(new_n10250_));
  XOR2_X1    g10058(.A1(new_n10250_), .A2(new_n9825_), .Z(new_n10251_));
  AOI21_X1   g10059(.A1(new_n9919_), .A2(new_n9874_), .B(\asqrt[20] ), .ZN(new_n10252_));
  XOR2_X1    g10060(.A1(new_n10252_), .A2(new_n9828_), .Z(new_n10253_));
  XOR2_X1    g10061(.A1(new_n9917_), .A2(\asqrt[51] ), .Z(new_n10254_));
  NOR2_X1    g10062(.A1(\asqrt[20] ), .A2(new_n10254_), .ZN(new_n10255_));
  XOR2_X1    g10063(.A1(new_n10255_), .A2(new_n9830_), .Z(new_n10256_));
  INV_X1     g10064(.I(new_n10256_), .ZN(new_n10257_));
  NOR2_X1    g10065(.A1(new_n9915_), .A2(new_n9869_), .ZN(new_n10258_));
  NOR2_X1    g10066(.A1(\asqrt[20] ), .A2(new_n10258_), .ZN(new_n10259_));
  XOR2_X1    g10067(.A1(new_n10259_), .A2(new_n9834_), .Z(new_n10260_));
  INV_X1     g10068(.I(new_n10260_), .ZN(new_n10261_));
  AOI21_X1   g10069(.A1(new_n9863_), .A2(new_n9868_), .B(\asqrt[20] ), .ZN(new_n10262_));
  XOR2_X1    g10070(.A1(new_n10262_), .A2(new_n9837_), .Z(new_n10263_));
  AOI21_X1   g10071(.A1(new_n9911_), .A2(new_n9862_), .B(\asqrt[20] ), .ZN(new_n10264_));
  XOR2_X1    g10072(.A1(new_n10264_), .A2(new_n9840_), .Z(new_n10265_));
  XOR2_X1    g10073(.A1(new_n9909_), .A2(\asqrt[47] ), .Z(new_n10266_));
  NOR2_X1    g10074(.A1(\asqrt[20] ), .A2(new_n10266_), .ZN(new_n10267_));
  XOR2_X1    g10075(.A1(new_n10267_), .A2(new_n9842_), .Z(new_n10268_));
  INV_X1     g10076(.I(new_n10268_), .ZN(new_n10269_));
  NOR2_X1    g10077(.A1(new_n9907_), .A2(new_n9857_), .ZN(new_n10270_));
  NOR2_X1    g10078(.A1(\asqrt[20] ), .A2(new_n10270_), .ZN(new_n10271_));
  XOR2_X1    g10079(.A1(new_n10271_), .A2(new_n9846_), .Z(new_n10272_));
  INV_X1     g10080(.I(new_n10272_), .ZN(new_n10273_));
  AOI21_X1   g10081(.A1(new_n9851_), .A2(new_n9856_), .B(\asqrt[20] ), .ZN(new_n10274_));
  XOR2_X1    g10082(.A1(new_n10274_), .A2(new_n9849_), .Z(new_n10275_));
  OAI21_X1   g10083(.A1(new_n10222_), .A2(\asqrt[45] ), .B(new_n9972_), .ZN(new_n10276_));
  NAND3_X1   g10084(.A1(new_n10276_), .A2(new_n10223_), .A3(new_n2134_), .ZN(new_n10277_));
  AOI21_X1   g10085(.A1(new_n10276_), .A2(new_n10223_), .B(new_n2134_), .ZN(new_n10278_));
  AOI21_X1   g10086(.A1(new_n10275_), .A2(new_n10277_), .B(new_n10278_), .ZN(new_n10279_));
  AOI21_X1   g10087(.A1(new_n10279_), .A2(new_n1953_), .B(new_n10273_), .ZN(new_n10280_));
  NAND2_X1   g10088(.A1(new_n10277_), .A2(new_n10275_), .ZN(new_n10281_));
  INV_X1     g10089(.I(new_n9972_), .ZN(new_n10282_));
  AOI21_X1   g10090(.A1(new_n10205_), .A2(new_n2332_), .B(new_n10282_), .ZN(new_n10283_));
  NAND2_X1   g10091(.A1(new_n10203_), .A2(new_n9975_), .ZN(new_n10284_));
  AOI21_X1   g10092(.A1(new_n10284_), .A2(new_n10221_), .B(new_n2332_), .ZN(new_n10285_));
  OAI21_X1   g10093(.A1(new_n10283_), .A2(new_n10285_), .B(\asqrt[46] ), .ZN(new_n10286_));
  AOI21_X1   g10094(.A1(new_n10281_), .A2(new_n10286_), .B(new_n1953_), .ZN(new_n10287_));
  NOR3_X1    g10095(.A1(new_n10280_), .A2(\asqrt[48] ), .A3(new_n10287_), .ZN(new_n10288_));
  OAI21_X1   g10096(.A1(new_n10280_), .A2(new_n10287_), .B(\asqrt[48] ), .ZN(new_n10289_));
  OAI21_X1   g10097(.A1(new_n10269_), .A2(new_n10288_), .B(new_n10289_), .ZN(new_n10290_));
  OAI21_X1   g10098(.A1(new_n10290_), .A2(\asqrt[49] ), .B(new_n10265_), .ZN(new_n10291_));
  NAND2_X1   g10099(.A1(new_n10290_), .A2(\asqrt[49] ), .ZN(new_n10292_));
  NAND3_X1   g10100(.A1(new_n10291_), .A2(new_n10292_), .A3(new_n1463_), .ZN(new_n10293_));
  AOI21_X1   g10101(.A1(new_n10291_), .A2(new_n10292_), .B(new_n1463_), .ZN(new_n10294_));
  AOI21_X1   g10102(.A1(new_n10263_), .A2(new_n10293_), .B(new_n10294_), .ZN(new_n10295_));
  AOI21_X1   g10103(.A1(new_n10295_), .A2(new_n1305_), .B(new_n10261_), .ZN(new_n10296_));
  NAND2_X1   g10104(.A1(new_n10293_), .A2(new_n10263_), .ZN(new_n10297_));
  INV_X1     g10105(.I(new_n10265_), .ZN(new_n10298_));
  INV_X1     g10106(.I(new_n10275_), .ZN(new_n10299_));
  NOR3_X1    g10107(.A1(new_n10283_), .A2(\asqrt[46] ), .A3(new_n10285_), .ZN(new_n10300_));
  OAI21_X1   g10108(.A1(new_n10299_), .A2(new_n10300_), .B(new_n10286_), .ZN(new_n10301_));
  OAI21_X1   g10109(.A1(new_n10301_), .A2(\asqrt[47] ), .B(new_n10272_), .ZN(new_n10302_));
  NAND2_X1   g10110(.A1(new_n10301_), .A2(\asqrt[47] ), .ZN(new_n10303_));
  NAND3_X1   g10111(.A1(new_n10302_), .A2(new_n10303_), .A3(new_n1778_), .ZN(new_n10304_));
  AOI21_X1   g10112(.A1(new_n10302_), .A2(new_n10303_), .B(new_n1778_), .ZN(new_n10305_));
  AOI21_X1   g10113(.A1(new_n10268_), .A2(new_n10304_), .B(new_n10305_), .ZN(new_n10306_));
  AOI21_X1   g10114(.A1(new_n10306_), .A2(new_n1632_), .B(new_n10298_), .ZN(new_n10307_));
  NAND2_X1   g10115(.A1(new_n10304_), .A2(new_n10268_), .ZN(new_n10308_));
  AOI21_X1   g10116(.A1(new_n10308_), .A2(new_n10289_), .B(new_n1632_), .ZN(new_n10309_));
  OAI21_X1   g10117(.A1(new_n10307_), .A2(new_n10309_), .B(\asqrt[50] ), .ZN(new_n10310_));
  AOI21_X1   g10118(.A1(new_n10297_), .A2(new_n10310_), .B(new_n1305_), .ZN(new_n10311_));
  NOR3_X1    g10119(.A1(new_n10296_), .A2(\asqrt[52] ), .A3(new_n10311_), .ZN(new_n10312_));
  OAI21_X1   g10120(.A1(new_n10296_), .A2(new_n10311_), .B(\asqrt[52] ), .ZN(new_n10313_));
  OAI21_X1   g10121(.A1(new_n10257_), .A2(new_n10312_), .B(new_n10313_), .ZN(new_n10314_));
  OAI21_X1   g10122(.A1(new_n10314_), .A2(\asqrt[53] ), .B(new_n10253_), .ZN(new_n10315_));
  NAND2_X1   g10123(.A1(new_n10314_), .A2(\asqrt[53] ), .ZN(new_n10316_));
  NAND3_X1   g10124(.A1(new_n10315_), .A2(new_n10316_), .A3(new_n860_), .ZN(new_n10317_));
  AOI21_X1   g10125(.A1(new_n10315_), .A2(new_n10316_), .B(new_n860_), .ZN(new_n10318_));
  AOI21_X1   g10126(.A1(new_n10251_), .A2(new_n10317_), .B(new_n10318_), .ZN(new_n10319_));
  AOI21_X1   g10127(.A1(new_n10319_), .A2(new_n744_), .B(new_n10249_), .ZN(new_n10320_));
  NAND2_X1   g10128(.A1(new_n10317_), .A2(new_n10251_), .ZN(new_n10321_));
  INV_X1     g10129(.I(new_n10253_), .ZN(new_n10322_));
  INV_X1     g10130(.I(new_n10263_), .ZN(new_n10323_));
  NOR3_X1    g10131(.A1(new_n10307_), .A2(\asqrt[50] ), .A3(new_n10309_), .ZN(new_n10324_));
  OAI21_X1   g10132(.A1(new_n10323_), .A2(new_n10324_), .B(new_n10310_), .ZN(new_n10325_));
  OAI21_X1   g10133(.A1(new_n10325_), .A2(\asqrt[51] ), .B(new_n10260_), .ZN(new_n10326_));
  NAND2_X1   g10134(.A1(new_n10325_), .A2(\asqrt[51] ), .ZN(new_n10327_));
  NAND3_X1   g10135(.A1(new_n10326_), .A2(new_n10327_), .A3(new_n1150_), .ZN(new_n10328_));
  AOI21_X1   g10136(.A1(new_n10326_), .A2(new_n10327_), .B(new_n1150_), .ZN(new_n10329_));
  AOI21_X1   g10137(.A1(new_n10256_), .A2(new_n10328_), .B(new_n10329_), .ZN(new_n10330_));
  AOI21_X1   g10138(.A1(new_n10330_), .A2(new_n1006_), .B(new_n10322_), .ZN(new_n10331_));
  NAND2_X1   g10139(.A1(new_n10328_), .A2(new_n10256_), .ZN(new_n10332_));
  AOI21_X1   g10140(.A1(new_n10332_), .A2(new_n10313_), .B(new_n1006_), .ZN(new_n10333_));
  OAI21_X1   g10141(.A1(new_n10331_), .A2(new_n10333_), .B(\asqrt[54] ), .ZN(new_n10334_));
  AOI21_X1   g10142(.A1(new_n10321_), .A2(new_n10334_), .B(new_n744_), .ZN(new_n10335_));
  NOR3_X1    g10143(.A1(new_n10320_), .A2(\asqrt[56] ), .A3(new_n10335_), .ZN(new_n10336_));
  OAI21_X1   g10144(.A1(new_n10320_), .A2(new_n10335_), .B(\asqrt[56] ), .ZN(new_n10337_));
  OAI21_X1   g10145(.A1(new_n10245_), .A2(new_n10336_), .B(new_n10337_), .ZN(new_n10338_));
  OAI21_X1   g10146(.A1(new_n10338_), .A2(\asqrt[57] ), .B(new_n10240_), .ZN(new_n10339_));
  NOR2_X1    g10147(.A1(new_n10336_), .A2(new_n10245_), .ZN(new_n10340_));
  INV_X1     g10148(.I(new_n10251_), .ZN(new_n10341_));
  NOR3_X1    g10149(.A1(new_n10331_), .A2(\asqrt[54] ), .A3(new_n10333_), .ZN(new_n10342_));
  OAI21_X1   g10150(.A1(new_n10341_), .A2(new_n10342_), .B(new_n10334_), .ZN(new_n10343_));
  OAI21_X1   g10151(.A1(new_n10343_), .A2(\asqrt[55] ), .B(new_n10248_), .ZN(new_n10344_));
  NAND2_X1   g10152(.A1(new_n10343_), .A2(\asqrt[55] ), .ZN(new_n10345_));
  AOI21_X1   g10153(.A1(new_n10344_), .A2(new_n10345_), .B(new_n634_), .ZN(new_n10346_));
  OAI21_X1   g10154(.A1(new_n10340_), .A2(new_n10346_), .B(\asqrt[57] ), .ZN(new_n10347_));
  NAND3_X1   g10155(.A1(new_n10339_), .A2(new_n423_), .A3(new_n10347_), .ZN(new_n10348_));
  NAND2_X1   g10156(.A1(new_n10348_), .A2(new_n10238_), .ZN(new_n10349_));
  INV_X1     g10157(.I(new_n10240_), .ZN(new_n10350_));
  NAND3_X1   g10158(.A1(new_n10344_), .A2(new_n10345_), .A3(new_n634_), .ZN(new_n10351_));
  AOI21_X1   g10159(.A1(new_n10244_), .A2(new_n10351_), .B(new_n10346_), .ZN(new_n10352_));
  AOI21_X1   g10160(.A1(new_n10352_), .A2(new_n531_), .B(new_n10350_), .ZN(new_n10353_));
  NAND2_X1   g10161(.A1(new_n10351_), .A2(new_n10244_), .ZN(new_n10354_));
  AOI21_X1   g10162(.A1(new_n10354_), .A2(new_n10337_), .B(new_n531_), .ZN(new_n10355_));
  OAI21_X1   g10163(.A1(new_n10353_), .A2(new_n10355_), .B(\asqrt[58] ), .ZN(new_n10356_));
  NAND3_X1   g10164(.A1(new_n10349_), .A2(new_n337_), .A3(new_n10356_), .ZN(new_n10357_));
  AOI21_X1   g10165(.A1(new_n10349_), .A2(new_n10356_), .B(new_n337_), .ZN(new_n10358_));
  AOI21_X1   g10166(.A1(new_n10236_), .A2(new_n10357_), .B(new_n10358_), .ZN(new_n10359_));
  AOI21_X1   g10167(.A1(new_n10359_), .A2(new_n266_), .B(new_n10233_), .ZN(new_n10360_));
  INV_X1     g10168(.I(new_n10238_), .ZN(new_n10361_));
  NOR3_X1    g10169(.A1(new_n10353_), .A2(\asqrt[58] ), .A3(new_n10355_), .ZN(new_n10362_));
  OAI21_X1   g10170(.A1(new_n10361_), .A2(new_n10362_), .B(new_n10356_), .ZN(new_n10363_));
  OAI21_X1   g10171(.A1(new_n10363_), .A2(\asqrt[59] ), .B(new_n10236_), .ZN(new_n10364_));
  NAND2_X1   g10172(.A1(new_n10363_), .A2(\asqrt[59] ), .ZN(new_n10365_));
  AOI21_X1   g10173(.A1(new_n10364_), .A2(new_n10365_), .B(new_n266_), .ZN(new_n10366_));
  OAI21_X1   g10174(.A1(new_n10360_), .A2(new_n10366_), .B(\asqrt[61] ), .ZN(new_n10367_));
  AOI21_X1   g10175(.A1(new_n9946_), .A2(new_n9941_), .B(\asqrt[20] ), .ZN(new_n10368_));
  XOR2_X1    g10176(.A1(new_n10368_), .A2(new_n9803_), .Z(new_n10369_));
  INV_X1     g10177(.I(new_n10369_), .ZN(new_n10370_));
  NOR3_X1    g10178(.A1(new_n10360_), .A2(\asqrt[61] ), .A3(new_n10366_), .ZN(new_n10371_));
  OAI21_X1   g10179(.A1(new_n10370_), .A2(new_n10371_), .B(new_n10367_), .ZN(new_n10372_));
  NAND3_X1   g10180(.A1(new_n10364_), .A2(new_n10365_), .A3(new_n266_), .ZN(new_n10373_));
  NAND2_X1   g10181(.A1(new_n10373_), .A2(new_n10232_), .ZN(new_n10374_));
  INV_X1     g10182(.I(new_n10236_), .ZN(new_n10375_));
  AOI21_X1   g10183(.A1(new_n10339_), .A2(new_n10347_), .B(new_n423_), .ZN(new_n10376_));
  AOI21_X1   g10184(.A1(new_n10238_), .A2(new_n10348_), .B(new_n10376_), .ZN(new_n10377_));
  AOI21_X1   g10185(.A1(new_n10377_), .A2(new_n337_), .B(new_n10375_), .ZN(new_n10378_));
  OAI21_X1   g10186(.A1(new_n10378_), .A2(new_n10358_), .B(\asqrt[60] ), .ZN(new_n10379_));
  AOI21_X1   g10187(.A1(new_n10374_), .A2(new_n10379_), .B(new_n239_), .ZN(new_n10380_));
  AOI21_X1   g10188(.A1(new_n10232_), .A2(new_n10373_), .B(new_n10366_), .ZN(new_n10381_));
  AOI21_X1   g10189(.A1(new_n10381_), .A2(new_n239_), .B(new_n10370_), .ZN(new_n10382_));
  OAI21_X1   g10190(.A1(new_n10382_), .A2(new_n10380_), .B(new_n201_), .ZN(new_n10383_));
  NOR3_X1    g10191(.A1(new_n10378_), .A2(\asqrt[60] ), .A3(new_n10358_), .ZN(new_n10384_));
  OAI21_X1   g10192(.A1(new_n10233_), .A2(new_n10384_), .B(new_n10379_), .ZN(new_n10385_));
  OAI21_X1   g10193(.A1(new_n10385_), .A2(\asqrt[61] ), .B(new_n10369_), .ZN(new_n10386_));
  NAND3_X1   g10194(.A1(new_n10386_), .A2(\asqrt[62] ), .A3(new_n10367_), .ZN(new_n10387_));
  AOI21_X1   g10195(.A1(new_n9936_), .A2(new_n9942_), .B(\asqrt[20] ), .ZN(new_n10388_));
  XOR2_X1    g10196(.A1(new_n10388_), .A2(new_n9938_), .Z(new_n10389_));
  INV_X1     g10197(.I(new_n10389_), .ZN(new_n10390_));
  AOI22_X1   g10198(.A1(new_n10387_), .A2(new_n10383_), .B1(new_n10372_), .B2(new_n10390_), .ZN(new_n10391_));
  NOR2_X1    g10199(.A1(new_n9955_), .A2(new_n9800_), .ZN(new_n10392_));
  OAI21_X1   g10200(.A1(\asqrt[20] ), .A2(new_n10392_), .B(new_n9962_), .ZN(new_n10393_));
  INV_X1     g10201(.I(new_n10393_), .ZN(new_n10394_));
  OAI21_X1   g10202(.A1(new_n10391_), .A2(new_n10229_), .B(new_n10394_), .ZN(new_n10395_));
  OAI21_X1   g10203(.A1(new_n10372_), .A2(\asqrt[62] ), .B(new_n10389_), .ZN(new_n10396_));
  NAND2_X1   g10204(.A1(new_n10372_), .A2(\asqrt[62] ), .ZN(new_n10397_));
  NAND3_X1   g10205(.A1(new_n10396_), .A2(new_n10397_), .A3(new_n10229_), .ZN(new_n10398_));
  NAND2_X1   g10206(.A1(new_n10052_), .A2(new_n9799_), .ZN(new_n10399_));
  XOR2_X1    g10207(.A1(new_n9955_), .A2(new_n9800_), .Z(new_n10400_));
  NAND3_X1   g10208(.A1(new_n10399_), .A2(\asqrt[63] ), .A3(new_n10400_), .ZN(new_n10401_));
  INV_X1     g10209(.I(new_n10041_), .ZN(new_n10402_));
  NAND4_X1   g10210(.A1(new_n10402_), .A2(new_n9800_), .A3(new_n9962_), .A4(new_n9969_), .ZN(new_n10403_));
  NAND2_X1   g10211(.A1(new_n10401_), .A2(new_n10403_), .ZN(new_n10404_));
  INV_X1     g10212(.I(new_n10404_), .ZN(new_n10405_));
  NAND4_X1   g10213(.A1(new_n10395_), .A2(new_n193_), .A3(new_n10398_), .A4(new_n10405_), .ZN(\asqrt[19] ));
  AOI21_X1   g10214(.A1(new_n10206_), .A2(new_n10223_), .B(\asqrt[19] ), .ZN(new_n10407_));
  XOR2_X1    g10215(.A1(new_n10407_), .A2(new_n9972_), .Z(new_n10408_));
  AOI21_X1   g10216(.A1(new_n10203_), .A2(new_n10221_), .B(\asqrt[19] ), .ZN(new_n10409_));
  XOR2_X1    g10217(.A1(new_n10409_), .A2(new_n9975_), .Z(new_n10410_));
  NAND2_X1   g10218(.A1(new_n10216_), .A2(new_n2749_), .ZN(new_n10411_));
  AOI21_X1   g10219(.A1(new_n10411_), .A2(new_n10202_), .B(\asqrt[19] ), .ZN(new_n10412_));
  XOR2_X1    g10220(.A1(new_n10412_), .A2(new_n9978_), .Z(new_n10413_));
  INV_X1     g10221(.I(new_n10413_), .ZN(new_n10414_));
  AOI21_X1   g10222(.A1(new_n10214_), .A2(new_n10199_), .B(\asqrt[19] ), .ZN(new_n10415_));
  XOR2_X1    g10223(.A1(new_n10415_), .A2(new_n9980_), .Z(new_n10416_));
  INV_X1     g10224(.I(new_n10416_), .ZN(new_n10417_));
  NAND2_X1   g10225(.A1(new_n10181_), .A2(new_n3195_), .ZN(new_n10418_));
  AOI21_X1   g10226(.A1(new_n10418_), .A2(new_n10213_), .B(\asqrt[19] ), .ZN(new_n10419_));
  XOR2_X1    g10227(.A1(new_n10419_), .A2(new_n9983_), .Z(new_n10420_));
  AOI21_X1   g10228(.A1(new_n10179_), .A2(new_n10196_), .B(\asqrt[19] ), .ZN(new_n10421_));
  XOR2_X1    g10229(.A1(new_n10421_), .A2(new_n9987_), .Z(new_n10422_));
  NAND2_X1   g10230(.A1(new_n10192_), .A2(new_n3681_), .ZN(new_n10423_));
  AOI21_X1   g10231(.A1(new_n10423_), .A2(new_n10178_), .B(\asqrt[19] ), .ZN(new_n10424_));
  XOR2_X1    g10232(.A1(new_n10424_), .A2(new_n9990_), .Z(new_n10425_));
  INV_X1     g10233(.I(new_n10425_), .ZN(new_n10426_));
  AOI21_X1   g10234(.A1(new_n10190_), .A2(new_n10175_), .B(\asqrt[19] ), .ZN(new_n10427_));
  XOR2_X1    g10235(.A1(new_n10427_), .A2(new_n9992_), .Z(new_n10428_));
  INV_X1     g10236(.I(new_n10428_), .ZN(new_n10429_));
  NAND2_X1   g10237(.A1(new_n10157_), .A2(new_n4196_), .ZN(new_n10430_));
  AOI21_X1   g10238(.A1(new_n10430_), .A2(new_n10189_), .B(\asqrt[19] ), .ZN(new_n10431_));
  XOR2_X1    g10239(.A1(new_n10431_), .A2(new_n9995_), .Z(new_n10432_));
  AOI21_X1   g10240(.A1(new_n10155_), .A2(new_n10172_), .B(\asqrt[19] ), .ZN(new_n10433_));
  XOR2_X1    g10241(.A1(new_n10433_), .A2(new_n9999_), .Z(new_n10434_));
  NAND2_X1   g10242(.A1(new_n10168_), .A2(new_n4751_), .ZN(new_n10435_));
  AOI21_X1   g10243(.A1(new_n10435_), .A2(new_n10154_), .B(\asqrt[19] ), .ZN(new_n10436_));
  XOR2_X1    g10244(.A1(new_n10436_), .A2(new_n10002_), .Z(new_n10437_));
  INV_X1     g10245(.I(new_n10437_), .ZN(new_n10438_));
  AOI21_X1   g10246(.A1(new_n10166_), .A2(new_n10151_), .B(\asqrt[19] ), .ZN(new_n10439_));
  XOR2_X1    g10247(.A1(new_n10439_), .A2(new_n10004_), .Z(new_n10440_));
  INV_X1     g10248(.I(new_n10440_), .ZN(new_n10441_));
  NAND2_X1   g10249(.A1(new_n10133_), .A2(new_n5336_), .ZN(new_n10442_));
  AOI21_X1   g10250(.A1(new_n10442_), .A2(new_n10165_), .B(\asqrt[19] ), .ZN(new_n10443_));
  XOR2_X1    g10251(.A1(new_n10443_), .A2(new_n10007_), .Z(new_n10444_));
  AOI21_X1   g10252(.A1(new_n10131_), .A2(new_n10148_), .B(\asqrt[19] ), .ZN(new_n10445_));
  XOR2_X1    g10253(.A1(new_n10445_), .A2(new_n10011_), .Z(new_n10446_));
  NAND2_X1   g10254(.A1(new_n10144_), .A2(new_n5947_), .ZN(new_n10447_));
  AOI21_X1   g10255(.A1(new_n10447_), .A2(new_n10130_), .B(\asqrt[19] ), .ZN(new_n10448_));
  XOR2_X1    g10256(.A1(new_n10448_), .A2(new_n10014_), .Z(new_n10449_));
  INV_X1     g10257(.I(new_n10449_), .ZN(new_n10450_));
  AOI21_X1   g10258(.A1(new_n10142_), .A2(new_n10127_), .B(\asqrt[19] ), .ZN(new_n10451_));
  XOR2_X1    g10259(.A1(new_n10451_), .A2(new_n10016_), .Z(new_n10452_));
  INV_X1     g10260(.I(new_n10452_), .ZN(new_n10453_));
  NAND2_X1   g10261(.A1(new_n10109_), .A2(new_n6636_), .ZN(new_n10454_));
  AOI21_X1   g10262(.A1(new_n10454_), .A2(new_n10141_), .B(\asqrt[19] ), .ZN(new_n10455_));
  XOR2_X1    g10263(.A1(new_n10455_), .A2(new_n10019_), .Z(new_n10456_));
  AOI21_X1   g10264(.A1(new_n10107_), .A2(new_n10124_), .B(\asqrt[19] ), .ZN(new_n10457_));
  XOR2_X1    g10265(.A1(new_n10457_), .A2(new_n10023_), .Z(new_n10458_));
  NAND2_X1   g10266(.A1(new_n10120_), .A2(new_n7331_), .ZN(new_n10459_));
  AOI21_X1   g10267(.A1(new_n10459_), .A2(new_n10106_), .B(\asqrt[19] ), .ZN(new_n10460_));
  XOR2_X1    g10268(.A1(new_n10460_), .A2(new_n10026_), .Z(new_n10461_));
  INV_X1     g10269(.I(new_n10461_), .ZN(new_n10462_));
  AOI21_X1   g10270(.A1(new_n10118_), .A2(new_n10103_), .B(\asqrt[19] ), .ZN(new_n10463_));
  XOR2_X1    g10271(.A1(new_n10463_), .A2(new_n10028_), .Z(new_n10464_));
  INV_X1     g10272(.I(new_n10464_), .ZN(new_n10465_));
  NAND2_X1   g10273(.A1(new_n10081_), .A2(new_n8077_), .ZN(new_n10466_));
  AOI21_X1   g10274(.A1(new_n10466_), .A2(new_n10117_), .B(\asqrt[19] ), .ZN(new_n10467_));
  XOR2_X1    g10275(.A1(new_n10467_), .A2(new_n10031_), .Z(new_n10468_));
  AOI21_X1   g10276(.A1(new_n10079_), .A2(new_n10100_), .B(\asqrt[19] ), .ZN(new_n10469_));
  XOR2_X1    g10277(.A1(new_n10469_), .A2(new_n10034_), .Z(new_n10470_));
  NAND2_X1   g10278(.A1(new_n10096_), .A2(new_n8849_), .ZN(new_n10471_));
  AOI21_X1   g10279(.A1(new_n10471_), .A2(new_n10078_), .B(\asqrt[19] ), .ZN(new_n10472_));
  XOR2_X1    g10280(.A1(new_n10472_), .A2(new_n10040_), .Z(new_n10473_));
  INV_X1     g10281(.I(new_n10473_), .ZN(new_n10474_));
  AOI21_X1   g10282(.A1(new_n10094_), .A2(new_n10075_), .B(\asqrt[19] ), .ZN(new_n10475_));
  XOR2_X1    g10283(.A1(new_n10475_), .A2(new_n10085_), .Z(new_n10476_));
  INV_X1     g10284(.I(new_n10476_), .ZN(new_n10477_));
  NAND2_X1   g10285(.A1(\asqrt[20] ), .A2(new_n10063_), .ZN(new_n10478_));
  NOR2_X1    g10286(.A1(new_n10070_), .A2(\a[40] ), .ZN(new_n10479_));
  AOI22_X1   g10287(.A1(new_n10478_), .A2(new_n10070_), .B1(\asqrt[20] ), .B2(new_n10479_), .ZN(new_n10480_));
  OAI21_X1   g10288(.A1(new_n10052_), .A2(new_n10063_), .B(new_n10089_), .ZN(new_n10481_));
  AOI21_X1   g10289(.A1(new_n10088_), .A2(new_n10481_), .B(\asqrt[19] ), .ZN(new_n10482_));
  XOR2_X1    g10290(.A1(new_n10482_), .A2(new_n10480_), .Z(new_n10483_));
  NOR2_X1    g10291(.A1(new_n10382_), .A2(new_n10380_), .ZN(new_n10484_));
  AOI21_X1   g10292(.A1(new_n10386_), .A2(new_n10367_), .B(\asqrt[62] ), .ZN(new_n10485_));
  NOR3_X1    g10293(.A1(new_n10382_), .A2(new_n201_), .A3(new_n10380_), .ZN(new_n10486_));
  OAI22_X1   g10294(.A1(new_n10485_), .A2(new_n10486_), .B1(new_n10484_), .B2(new_n10389_), .ZN(new_n10487_));
  AOI21_X1   g10295(.A1(new_n10487_), .A2(new_n10228_), .B(new_n10393_), .ZN(new_n10488_));
  AOI21_X1   g10296(.A1(new_n10484_), .A2(new_n201_), .B(new_n10390_), .ZN(new_n10489_));
  NOR2_X1    g10297(.A1(new_n10484_), .A2(new_n201_), .ZN(new_n10490_));
  NOR3_X1    g10298(.A1(new_n10489_), .A2(new_n10490_), .A3(new_n10228_), .ZN(new_n10491_));
  NAND3_X1   g10299(.A1(new_n10401_), .A2(\asqrt[20] ), .A3(new_n10403_), .ZN(new_n10492_));
  NOR4_X1    g10300(.A1(new_n10488_), .A2(\asqrt[63] ), .A3(new_n10491_), .A4(new_n10492_), .ZN(new_n10493_));
  INV_X1     g10301(.I(new_n10493_), .ZN(new_n10494_));
  NAND2_X1   g10302(.A1(\asqrt[19] ), .A2(new_n10060_), .ZN(new_n10495_));
  AOI21_X1   g10303(.A1(new_n10495_), .A2(new_n10494_), .B(\a[40] ), .ZN(new_n10496_));
  NOR4_X1    g10304(.A1(new_n10488_), .A2(\asqrt[63] ), .A3(new_n10491_), .A4(new_n10404_), .ZN(new_n10497_));
  NOR2_X1    g10305(.A1(new_n10497_), .A2(new_n10061_), .ZN(new_n10498_));
  NOR3_X1    g10306(.A1(new_n10498_), .A2(new_n10063_), .A3(new_n10493_), .ZN(new_n10499_));
  NOR2_X1    g10307(.A1(new_n10499_), .A2(new_n10496_), .ZN(new_n10500_));
  INV_X1     g10308(.I(\a[38] ), .ZN(new_n10501_));
  NOR2_X1    g10309(.A1(\a[36] ), .A2(\a[37] ), .ZN(new_n10502_));
  NOR3_X1    g10310(.A1(new_n10497_), .A2(new_n10501_), .A3(new_n10502_), .ZN(new_n10503_));
  INV_X1     g10311(.I(new_n10502_), .ZN(new_n10504_));
  AOI21_X1   g10312(.A1(new_n10497_), .A2(\a[38] ), .B(new_n10504_), .ZN(new_n10505_));
  OAI21_X1   g10313(.A1(new_n10503_), .A2(new_n10505_), .B(\asqrt[20] ), .ZN(new_n10506_));
  NAND2_X1   g10314(.A1(new_n10502_), .A2(new_n10501_), .ZN(new_n10507_));
  NAND3_X1   g10315(.A1(new_n9965_), .A2(new_n9967_), .A3(new_n10507_), .ZN(new_n10508_));
  NAND2_X1   g10316(.A1(new_n10055_), .A2(new_n10508_), .ZN(new_n10509_));
  NAND3_X1   g10317(.A1(\asqrt[19] ), .A2(\a[38] ), .A3(new_n10509_), .ZN(new_n10510_));
  NOR3_X1    g10318(.A1(new_n10497_), .A2(\a[38] ), .A3(\a[39] ), .ZN(new_n10511_));
  INV_X1     g10319(.I(\a[39] ), .ZN(new_n10512_));
  AOI21_X1   g10320(.A1(\asqrt[19] ), .A2(new_n10501_), .B(new_n10512_), .ZN(new_n10513_));
  NOR2_X1    g10321(.A1(new_n10511_), .A2(new_n10513_), .ZN(new_n10514_));
  NAND4_X1   g10322(.A1(new_n10506_), .A2(new_n10514_), .A3(new_n9656_), .A4(new_n10510_), .ZN(new_n10515_));
  NAND2_X1   g10323(.A1(new_n10515_), .A2(new_n10500_), .ZN(new_n10516_));
  NAND3_X1   g10324(.A1(\asqrt[19] ), .A2(\a[38] ), .A3(new_n10504_), .ZN(new_n10517_));
  OAI21_X1   g10325(.A1(\asqrt[19] ), .A2(new_n10501_), .B(new_n10502_), .ZN(new_n10518_));
  AOI21_X1   g10326(.A1(new_n10518_), .A2(new_n10517_), .B(new_n10052_), .ZN(new_n10519_));
  NAND3_X1   g10327(.A1(\asqrt[19] ), .A2(new_n10501_), .A3(new_n10512_), .ZN(new_n10520_));
  OAI21_X1   g10328(.A1(new_n10497_), .A2(\a[38] ), .B(\a[39] ), .ZN(new_n10521_));
  NAND3_X1   g10329(.A1(new_n10510_), .A2(new_n10521_), .A3(new_n10520_), .ZN(new_n10522_));
  OAI21_X1   g10330(.A1(new_n10522_), .A2(new_n10519_), .B(\asqrt[21] ), .ZN(new_n10523_));
  NAND3_X1   g10331(.A1(new_n10516_), .A2(new_n9233_), .A3(new_n10523_), .ZN(new_n10524_));
  AOI21_X1   g10332(.A1(new_n10516_), .A2(new_n10523_), .B(new_n9233_), .ZN(new_n10525_));
  AOI21_X1   g10333(.A1(new_n10483_), .A2(new_n10524_), .B(new_n10525_), .ZN(new_n10526_));
  AOI21_X1   g10334(.A1(new_n10526_), .A2(new_n8849_), .B(new_n10477_), .ZN(new_n10527_));
  OR2_X2     g10335(.A1(new_n10499_), .A2(new_n10496_), .Z(new_n10528_));
  NOR3_X1    g10336(.A1(new_n10522_), .A2(new_n10519_), .A3(\asqrt[21] ), .ZN(new_n10529_));
  OAI21_X1   g10337(.A1(new_n10528_), .A2(new_n10529_), .B(new_n10523_), .ZN(new_n10530_));
  OAI21_X1   g10338(.A1(new_n10530_), .A2(\asqrt[22] ), .B(new_n10483_), .ZN(new_n10531_));
  NAND2_X1   g10339(.A1(new_n10530_), .A2(\asqrt[22] ), .ZN(new_n10532_));
  AOI21_X1   g10340(.A1(new_n10531_), .A2(new_n10532_), .B(new_n8849_), .ZN(new_n10533_));
  NOR3_X1    g10341(.A1(new_n10527_), .A2(\asqrt[24] ), .A3(new_n10533_), .ZN(new_n10534_));
  OAI21_X1   g10342(.A1(new_n10527_), .A2(new_n10533_), .B(\asqrt[24] ), .ZN(new_n10535_));
  OAI21_X1   g10343(.A1(new_n10474_), .A2(new_n10534_), .B(new_n10535_), .ZN(new_n10536_));
  OAI21_X1   g10344(.A1(new_n10536_), .A2(\asqrt[25] ), .B(new_n10470_), .ZN(new_n10537_));
  NAND3_X1   g10345(.A1(new_n10531_), .A2(new_n10532_), .A3(new_n8849_), .ZN(new_n10538_));
  AOI21_X1   g10346(.A1(new_n10476_), .A2(new_n10538_), .B(new_n10533_), .ZN(new_n10539_));
  AOI21_X1   g10347(.A1(new_n10539_), .A2(new_n8440_), .B(new_n10474_), .ZN(new_n10540_));
  NAND2_X1   g10348(.A1(new_n10538_), .A2(new_n10476_), .ZN(new_n10541_));
  INV_X1     g10349(.I(new_n10533_), .ZN(new_n10542_));
  AOI21_X1   g10350(.A1(new_n10541_), .A2(new_n10542_), .B(new_n8440_), .ZN(new_n10543_));
  OAI21_X1   g10351(.A1(new_n10540_), .A2(new_n10543_), .B(\asqrt[25] ), .ZN(new_n10544_));
  NAND3_X1   g10352(.A1(new_n10537_), .A2(new_n7690_), .A3(new_n10544_), .ZN(new_n10545_));
  AOI21_X1   g10353(.A1(new_n10537_), .A2(new_n10544_), .B(new_n7690_), .ZN(new_n10546_));
  AOI21_X1   g10354(.A1(new_n10468_), .A2(new_n10545_), .B(new_n10546_), .ZN(new_n10547_));
  AOI21_X1   g10355(.A1(new_n10547_), .A2(new_n7331_), .B(new_n10465_), .ZN(new_n10548_));
  INV_X1     g10356(.I(new_n10470_), .ZN(new_n10549_));
  NOR3_X1    g10357(.A1(new_n10540_), .A2(\asqrt[25] ), .A3(new_n10543_), .ZN(new_n10550_));
  OAI21_X1   g10358(.A1(new_n10549_), .A2(new_n10550_), .B(new_n10544_), .ZN(new_n10551_));
  OAI21_X1   g10359(.A1(new_n10551_), .A2(\asqrt[26] ), .B(new_n10468_), .ZN(new_n10552_));
  NAND2_X1   g10360(.A1(new_n10551_), .A2(\asqrt[26] ), .ZN(new_n10553_));
  AOI21_X1   g10361(.A1(new_n10552_), .A2(new_n10553_), .B(new_n7331_), .ZN(new_n10554_));
  NOR3_X1    g10362(.A1(new_n10548_), .A2(\asqrt[28] ), .A3(new_n10554_), .ZN(new_n10555_));
  OAI21_X1   g10363(.A1(new_n10548_), .A2(new_n10554_), .B(\asqrt[28] ), .ZN(new_n10556_));
  OAI21_X1   g10364(.A1(new_n10462_), .A2(new_n10555_), .B(new_n10556_), .ZN(new_n10557_));
  OAI21_X1   g10365(.A1(new_n10557_), .A2(\asqrt[29] ), .B(new_n10458_), .ZN(new_n10558_));
  NAND3_X1   g10366(.A1(new_n10552_), .A2(new_n10553_), .A3(new_n7331_), .ZN(new_n10559_));
  AOI21_X1   g10367(.A1(new_n10464_), .A2(new_n10559_), .B(new_n10554_), .ZN(new_n10560_));
  AOI21_X1   g10368(.A1(new_n10560_), .A2(new_n6966_), .B(new_n10462_), .ZN(new_n10561_));
  NAND2_X1   g10369(.A1(new_n10559_), .A2(new_n10464_), .ZN(new_n10562_));
  INV_X1     g10370(.I(new_n10554_), .ZN(new_n10563_));
  AOI21_X1   g10371(.A1(new_n10562_), .A2(new_n10563_), .B(new_n6966_), .ZN(new_n10564_));
  OAI21_X1   g10372(.A1(new_n10561_), .A2(new_n10564_), .B(\asqrt[29] ), .ZN(new_n10565_));
  NAND3_X1   g10373(.A1(new_n10558_), .A2(new_n6275_), .A3(new_n10565_), .ZN(new_n10566_));
  AOI21_X1   g10374(.A1(new_n10558_), .A2(new_n10565_), .B(new_n6275_), .ZN(new_n10567_));
  AOI21_X1   g10375(.A1(new_n10456_), .A2(new_n10566_), .B(new_n10567_), .ZN(new_n10568_));
  AOI21_X1   g10376(.A1(new_n10568_), .A2(new_n5947_), .B(new_n10453_), .ZN(new_n10569_));
  INV_X1     g10377(.I(new_n10458_), .ZN(new_n10570_));
  NOR3_X1    g10378(.A1(new_n10561_), .A2(\asqrt[29] ), .A3(new_n10564_), .ZN(new_n10571_));
  OAI21_X1   g10379(.A1(new_n10570_), .A2(new_n10571_), .B(new_n10565_), .ZN(new_n10572_));
  OAI21_X1   g10380(.A1(new_n10572_), .A2(\asqrt[30] ), .B(new_n10456_), .ZN(new_n10573_));
  NAND2_X1   g10381(.A1(new_n10572_), .A2(\asqrt[30] ), .ZN(new_n10574_));
  AOI21_X1   g10382(.A1(new_n10573_), .A2(new_n10574_), .B(new_n5947_), .ZN(new_n10575_));
  NOR3_X1    g10383(.A1(new_n10569_), .A2(\asqrt[32] ), .A3(new_n10575_), .ZN(new_n10576_));
  OAI21_X1   g10384(.A1(new_n10569_), .A2(new_n10575_), .B(\asqrt[32] ), .ZN(new_n10577_));
  OAI21_X1   g10385(.A1(new_n10450_), .A2(new_n10576_), .B(new_n10577_), .ZN(new_n10578_));
  OAI21_X1   g10386(.A1(new_n10578_), .A2(\asqrt[33] ), .B(new_n10446_), .ZN(new_n10579_));
  NAND3_X1   g10387(.A1(new_n10573_), .A2(new_n10574_), .A3(new_n5947_), .ZN(new_n10580_));
  AOI21_X1   g10388(.A1(new_n10452_), .A2(new_n10580_), .B(new_n10575_), .ZN(new_n10581_));
  AOI21_X1   g10389(.A1(new_n10581_), .A2(new_n5643_), .B(new_n10450_), .ZN(new_n10582_));
  NAND2_X1   g10390(.A1(new_n10580_), .A2(new_n10452_), .ZN(new_n10583_));
  INV_X1     g10391(.I(new_n10575_), .ZN(new_n10584_));
  AOI21_X1   g10392(.A1(new_n10583_), .A2(new_n10584_), .B(new_n5643_), .ZN(new_n10585_));
  OAI21_X1   g10393(.A1(new_n10582_), .A2(new_n10585_), .B(\asqrt[33] ), .ZN(new_n10586_));
  NAND3_X1   g10394(.A1(new_n10579_), .A2(new_n5029_), .A3(new_n10586_), .ZN(new_n10587_));
  AOI21_X1   g10395(.A1(new_n10579_), .A2(new_n10586_), .B(new_n5029_), .ZN(new_n10588_));
  AOI21_X1   g10396(.A1(new_n10444_), .A2(new_n10587_), .B(new_n10588_), .ZN(new_n10589_));
  AOI21_X1   g10397(.A1(new_n10589_), .A2(new_n4751_), .B(new_n10441_), .ZN(new_n10590_));
  INV_X1     g10398(.I(new_n10446_), .ZN(new_n10591_));
  NOR3_X1    g10399(.A1(new_n10582_), .A2(\asqrt[33] ), .A3(new_n10585_), .ZN(new_n10592_));
  OAI21_X1   g10400(.A1(new_n10591_), .A2(new_n10592_), .B(new_n10586_), .ZN(new_n10593_));
  OAI21_X1   g10401(.A1(new_n10593_), .A2(\asqrt[34] ), .B(new_n10444_), .ZN(new_n10594_));
  NAND2_X1   g10402(.A1(new_n10593_), .A2(\asqrt[34] ), .ZN(new_n10595_));
  AOI21_X1   g10403(.A1(new_n10594_), .A2(new_n10595_), .B(new_n4751_), .ZN(new_n10596_));
  NOR3_X1    g10404(.A1(new_n10590_), .A2(\asqrt[36] ), .A3(new_n10596_), .ZN(new_n10597_));
  OAI21_X1   g10405(.A1(new_n10590_), .A2(new_n10596_), .B(\asqrt[36] ), .ZN(new_n10598_));
  OAI21_X1   g10406(.A1(new_n10438_), .A2(new_n10597_), .B(new_n10598_), .ZN(new_n10599_));
  OAI21_X1   g10407(.A1(new_n10599_), .A2(\asqrt[37] ), .B(new_n10434_), .ZN(new_n10600_));
  NAND3_X1   g10408(.A1(new_n10594_), .A2(new_n10595_), .A3(new_n4751_), .ZN(new_n10601_));
  AOI21_X1   g10409(.A1(new_n10440_), .A2(new_n10601_), .B(new_n10596_), .ZN(new_n10602_));
  AOI21_X1   g10410(.A1(new_n10602_), .A2(new_n4461_), .B(new_n10438_), .ZN(new_n10603_));
  NAND2_X1   g10411(.A1(new_n10601_), .A2(new_n10440_), .ZN(new_n10604_));
  INV_X1     g10412(.I(new_n10596_), .ZN(new_n10605_));
  AOI21_X1   g10413(.A1(new_n10604_), .A2(new_n10605_), .B(new_n4461_), .ZN(new_n10606_));
  OAI21_X1   g10414(.A1(new_n10603_), .A2(new_n10606_), .B(\asqrt[37] ), .ZN(new_n10607_));
  NAND3_X1   g10415(.A1(new_n10600_), .A2(new_n3925_), .A3(new_n10607_), .ZN(new_n10608_));
  AOI21_X1   g10416(.A1(new_n10600_), .A2(new_n10607_), .B(new_n3925_), .ZN(new_n10609_));
  AOI21_X1   g10417(.A1(new_n10432_), .A2(new_n10608_), .B(new_n10609_), .ZN(new_n10610_));
  AOI21_X1   g10418(.A1(new_n10610_), .A2(new_n3681_), .B(new_n10429_), .ZN(new_n10611_));
  INV_X1     g10419(.I(new_n10434_), .ZN(new_n10612_));
  NOR3_X1    g10420(.A1(new_n10603_), .A2(\asqrt[37] ), .A3(new_n10606_), .ZN(new_n10613_));
  OAI21_X1   g10421(.A1(new_n10612_), .A2(new_n10613_), .B(new_n10607_), .ZN(new_n10614_));
  OAI21_X1   g10422(.A1(new_n10614_), .A2(\asqrt[38] ), .B(new_n10432_), .ZN(new_n10615_));
  NAND2_X1   g10423(.A1(new_n10614_), .A2(\asqrt[38] ), .ZN(new_n10616_));
  AOI21_X1   g10424(.A1(new_n10615_), .A2(new_n10616_), .B(new_n3681_), .ZN(new_n10617_));
  NOR3_X1    g10425(.A1(new_n10611_), .A2(\asqrt[40] ), .A3(new_n10617_), .ZN(new_n10618_));
  OAI21_X1   g10426(.A1(new_n10611_), .A2(new_n10617_), .B(\asqrt[40] ), .ZN(new_n10619_));
  OAI21_X1   g10427(.A1(new_n10426_), .A2(new_n10618_), .B(new_n10619_), .ZN(new_n10620_));
  OAI21_X1   g10428(.A1(new_n10620_), .A2(\asqrt[41] ), .B(new_n10422_), .ZN(new_n10621_));
  NAND3_X1   g10429(.A1(new_n10615_), .A2(new_n10616_), .A3(new_n3681_), .ZN(new_n10622_));
  AOI21_X1   g10430(.A1(new_n10428_), .A2(new_n10622_), .B(new_n10617_), .ZN(new_n10623_));
  AOI21_X1   g10431(.A1(new_n10623_), .A2(new_n3427_), .B(new_n10426_), .ZN(new_n10624_));
  NAND2_X1   g10432(.A1(new_n10622_), .A2(new_n10428_), .ZN(new_n10625_));
  INV_X1     g10433(.I(new_n10617_), .ZN(new_n10626_));
  AOI21_X1   g10434(.A1(new_n10625_), .A2(new_n10626_), .B(new_n3427_), .ZN(new_n10627_));
  OAI21_X1   g10435(.A1(new_n10624_), .A2(new_n10627_), .B(\asqrt[41] ), .ZN(new_n10628_));
  NAND3_X1   g10436(.A1(new_n10621_), .A2(new_n2960_), .A3(new_n10628_), .ZN(new_n10629_));
  AOI21_X1   g10437(.A1(new_n10621_), .A2(new_n10628_), .B(new_n2960_), .ZN(new_n10630_));
  AOI21_X1   g10438(.A1(new_n10420_), .A2(new_n10629_), .B(new_n10630_), .ZN(new_n10631_));
  AOI21_X1   g10439(.A1(new_n10631_), .A2(new_n2749_), .B(new_n10417_), .ZN(new_n10632_));
  INV_X1     g10440(.I(new_n10422_), .ZN(new_n10633_));
  NOR3_X1    g10441(.A1(new_n10624_), .A2(\asqrt[41] ), .A3(new_n10627_), .ZN(new_n10634_));
  OAI21_X1   g10442(.A1(new_n10633_), .A2(new_n10634_), .B(new_n10628_), .ZN(new_n10635_));
  OAI21_X1   g10443(.A1(new_n10635_), .A2(\asqrt[42] ), .B(new_n10420_), .ZN(new_n10636_));
  NAND2_X1   g10444(.A1(new_n10635_), .A2(\asqrt[42] ), .ZN(new_n10637_));
  AOI21_X1   g10445(.A1(new_n10636_), .A2(new_n10637_), .B(new_n2749_), .ZN(new_n10638_));
  NOR3_X1    g10446(.A1(new_n10632_), .A2(\asqrt[44] ), .A3(new_n10638_), .ZN(new_n10639_));
  OAI21_X1   g10447(.A1(new_n10632_), .A2(new_n10638_), .B(\asqrt[44] ), .ZN(new_n10640_));
  OAI21_X1   g10448(.A1(new_n10414_), .A2(new_n10639_), .B(new_n10640_), .ZN(new_n10641_));
  OAI21_X1   g10449(.A1(new_n10641_), .A2(\asqrt[45] ), .B(new_n10410_), .ZN(new_n10642_));
  NAND3_X1   g10450(.A1(new_n10636_), .A2(new_n10637_), .A3(new_n2749_), .ZN(new_n10643_));
  AOI21_X1   g10451(.A1(new_n10416_), .A2(new_n10643_), .B(new_n10638_), .ZN(new_n10644_));
  AOI21_X1   g10452(.A1(new_n10644_), .A2(new_n2531_), .B(new_n10414_), .ZN(new_n10645_));
  NAND2_X1   g10453(.A1(new_n10643_), .A2(new_n10416_), .ZN(new_n10646_));
  INV_X1     g10454(.I(new_n10638_), .ZN(new_n10647_));
  AOI21_X1   g10455(.A1(new_n10646_), .A2(new_n10647_), .B(new_n2531_), .ZN(new_n10648_));
  OAI21_X1   g10456(.A1(new_n10645_), .A2(new_n10648_), .B(\asqrt[45] ), .ZN(new_n10649_));
  NAND3_X1   g10457(.A1(new_n10642_), .A2(new_n2134_), .A3(new_n10649_), .ZN(new_n10650_));
  INV_X1     g10458(.I(new_n10410_), .ZN(new_n10651_));
  NOR3_X1    g10459(.A1(new_n10645_), .A2(\asqrt[45] ), .A3(new_n10648_), .ZN(new_n10652_));
  OAI21_X1   g10460(.A1(new_n10651_), .A2(new_n10652_), .B(new_n10649_), .ZN(new_n10653_));
  NAND2_X1   g10461(.A1(new_n10653_), .A2(\asqrt[46] ), .ZN(new_n10654_));
  NOR2_X1    g10462(.A1(new_n10372_), .A2(\asqrt[62] ), .ZN(new_n10655_));
  NOR2_X1    g10463(.A1(new_n10655_), .A2(new_n10490_), .ZN(new_n10656_));
  XOR2_X1    g10464(.A1(new_n10388_), .A2(new_n9938_), .Z(new_n10657_));
  OAI21_X1   g10465(.A1(\asqrt[19] ), .A2(new_n10656_), .B(new_n10657_), .ZN(new_n10658_));
  INV_X1     g10466(.I(new_n10658_), .ZN(new_n10659_));
  AOI21_X1   g10467(.A1(new_n10357_), .A2(new_n10365_), .B(\asqrt[19] ), .ZN(new_n10660_));
  XOR2_X1    g10468(.A1(new_n10660_), .A2(new_n10236_), .Z(new_n10661_));
  INV_X1     g10469(.I(new_n10661_), .ZN(new_n10662_));
  AOI21_X1   g10470(.A1(new_n10348_), .A2(new_n10356_), .B(\asqrt[19] ), .ZN(new_n10663_));
  XOR2_X1    g10471(.A1(new_n10663_), .A2(new_n10238_), .Z(new_n10664_));
  INV_X1     g10472(.I(new_n10664_), .ZN(new_n10665_));
  NAND2_X1   g10473(.A1(new_n10352_), .A2(new_n531_), .ZN(new_n10666_));
  AOI21_X1   g10474(.A1(new_n10666_), .A2(new_n10347_), .B(\asqrt[19] ), .ZN(new_n10667_));
  XOR2_X1    g10475(.A1(new_n10667_), .A2(new_n10240_), .Z(new_n10668_));
  AOI21_X1   g10476(.A1(new_n10351_), .A2(new_n10337_), .B(\asqrt[19] ), .ZN(new_n10669_));
  XOR2_X1    g10477(.A1(new_n10669_), .A2(new_n10244_), .Z(new_n10670_));
  NAND2_X1   g10478(.A1(new_n10319_), .A2(new_n744_), .ZN(new_n10671_));
  AOI21_X1   g10479(.A1(new_n10671_), .A2(new_n10345_), .B(\asqrt[19] ), .ZN(new_n10672_));
  XOR2_X1    g10480(.A1(new_n10672_), .A2(new_n10248_), .Z(new_n10673_));
  INV_X1     g10481(.I(new_n10673_), .ZN(new_n10674_));
  AOI21_X1   g10482(.A1(new_n10317_), .A2(new_n10334_), .B(\asqrt[19] ), .ZN(new_n10675_));
  XOR2_X1    g10483(.A1(new_n10675_), .A2(new_n10251_), .Z(new_n10676_));
  INV_X1     g10484(.I(new_n10676_), .ZN(new_n10677_));
  NAND2_X1   g10485(.A1(new_n10330_), .A2(new_n1006_), .ZN(new_n10678_));
  AOI21_X1   g10486(.A1(new_n10678_), .A2(new_n10316_), .B(\asqrt[19] ), .ZN(new_n10679_));
  XOR2_X1    g10487(.A1(new_n10679_), .A2(new_n10253_), .Z(new_n10680_));
  AOI21_X1   g10488(.A1(new_n10328_), .A2(new_n10313_), .B(\asqrt[19] ), .ZN(new_n10681_));
  XOR2_X1    g10489(.A1(new_n10681_), .A2(new_n10256_), .Z(new_n10682_));
  NAND2_X1   g10490(.A1(new_n10295_), .A2(new_n1305_), .ZN(new_n10683_));
  AOI21_X1   g10491(.A1(new_n10683_), .A2(new_n10327_), .B(\asqrt[19] ), .ZN(new_n10684_));
  XOR2_X1    g10492(.A1(new_n10684_), .A2(new_n10260_), .Z(new_n10685_));
  INV_X1     g10493(.I(new_n10685_), .ZN(new_n10686_));
  AOI21_X1   g10494(.A1(new_n10293_), .A2(new_n10310_), .B(\asqrt[19] ), .ZN(new_n10687_));
  XOR2_X1    g10495(.A1(new_n10687_), .A2(new_n10263_), .Z(new_n10688_));
  INV_X1     g10496(.I(new_n10688_), .ZN(new_n10689_));
  NAND2_X1   g10497(.A1(new_n10306_), .A2(new_n1632_), .ZN(new_n10690_));
  AOI21_X1   g10498(.A1(new_n10690_), .A2(new_n10292_), .B(\asqrt[19] ), .ZN(new_n10691_));
  XOR2_X1    g10499(.A1(new_n10691_), .A2(new_n10265_), .Z(new_n10692_));
  AOI21_X1   g10500(.A1(new_n10304_), .A2(new_n10289_), .B(\asqrt[19] ), .ZN(new_n10693_));
  XOR2_X1    g10501(.A1(new_n10693_), .A2(new_n10268_), .Z(new_n10694_));
  NAND2_X1   g10502(.A1(new_n10279_), .A2(new_n1953_), .ZN(new_n10695_));
  AOI21_X1   g10503(.A1(new_n10695_), .A2(new_n10303_), .B(\asqrt[19] ), .ZN(new_n10696_));
  XOR2_X1    g10504(.A1(new_n10696_), .A2(new_n10272_), .Z(new_n10697_));
  INV_X1     g10505(.I(new_n10697_), .ZN(new_n10698_));
  AOI21_X1   g10506(.A1(new_n10277_), .A2(new_n10286_), .B(\asqrt[19] ), .ZN(new_n10699_));
  XOR2_X1    g10507(.A1(new_n10699_), .A2(new_n10275_), .Z(new_n10700_));
  INV_X1     g10508(.I(new_n10700_), .ZN(new_n10701_));
  AOI21_X1   g10509(.A1(new_n10642_), .A2(new_n10649_), .B(new_n2134_), .ZN(new_n10702_));
  AOI21_X1   g10510(.A1(new_n10408_), .A2(new_n10650_), .B(new_n10702_), .ZN(new_n10703_));
  AOI21_X1   g10511(.A1(new_n10703_), .A2(new_n1953_), .B(new_n10701_), .ZN(new_n10704_));
  OAI21_X1   g10512(.A1(new_n10653_), .A2(\asqrt[46] ), .B(new_n10408_), .ZN(new_n10705_));
  AOI21_X1   g10513(.A1(new_n10705_), .A2(new_n10654_), .B(new_n1953_), .ZN(new_n10706_));
  NOR3_X1    g10514(.A1(new_n10704_), .A2(\asqrt[48] ), .A3(new_n10706_), .ZN(new_n10707_));
  OAI21_X1   g10515(.A1(new_n10704_), .A2(new_n10706_), .B(\asqrt[48] ), .ZN(new_n10708_));
  OAI21_X1   g10516(.A1(new_n10698_), .A2(new_n10707_), .B(new_n10708_), .ZN(new_n10709_));
  OAI21_X1   g10517(.A1(new_n10709_), .A2(\asqrt[49] ), .B(new_n10694_), .ZN(new_n10710_));
  NAND3_X1   g10518(.A1(new_n10705_), .A2(new_n10654_), .A3(new_n1953_), .ZN(new_n10711_));
  AOI21_X1   g10519(.A1(new_n10700_), .A2(new_n10711_), .B(new_n10706_), .ZN(new_n10712_));
  AOI21_X1   g10520(.A1(new_n10712_), .A2(new_n1778_), .B(new_n10698_), .ZN(new_n10713_));
  NAND2_X1   g10521(.A1(new_n10711_), .A2(new_n10700_), .ZN(new_n10714_));
  INV_X1     g10522(.I(new_n10706_), .ZN(new_n10715_));
  AOI21_X1   g10523(.A1(new_n10714_), .A2(new_n10715_), .B(new_n1778_), .ZN(new_n10716_));
  OAI21_X1   g10524(.A1(new_n10713_), .A2(new_n10716_), .B(\asqrt[49] ), .ZN(new_n10717_));
  NAND3_X1   g10525(.A1(new_n10710_), .A2(new_n1463_), .A3(new_n10717_), .ZN(new_n10718_));
  AOI21_X1   g10526(.A1(new_n10710_), .A2(new_n10717_), .B(new_n1463_), .ZN(new_n10719_));
  AOI21_X1   g10527(.A1(new_n10692_), .A2(new_n10718_), .B(new_n10719_), .ZN(new_n10720_));
  AOI21_X1   g10528(.A1(new_n10720_), .A2(new_n1305_), .B(new_n10689_), .ZN(new_n10721_));
  INV_X1     g10529(.I(new_n10694_), .ZN(new_n10722_));
  NOR3_X1    g10530(.A1(new_n10713_), .A2(\asqrt[49] ), .A3(new_n10716_), .ZN(new_n10723_));
  OAI21_X1   g10531(.A1(new_n10722_), .A2(new_n10723_), .B(new_n10717_), .ZN(new_n10724_));
  OAI21_X1   g10532(.A1(new_n10724_), .A2(\asqrt[50] ), .B(new_n10692_), .ZN(new_n10725_));
  NAND2_X1   g10533(.A1(new_n10724_), .A2(\asqrt[50] ), .ZN(new_n10726_));
  AOI21_X1   g10534(.A1(new_n10725_), .A2(new_n10726_), .B(new_n1305_), .ZN(new_n10727_));
  NOR3_X1    g10535(.A1(new_n10721_), .A2(\asqrt[52] ), .A3(new_n10727_), .ZN(new_n10728_));
  OAI21_X1   g10536(.A1(new_n10721_), .A2(new_n10727_), .B(\asqrt[52] ), .ZN(new_n10729_));
  OAI21_X1   g10537(.A1(new_n10686_), .A2(new_n10728_), .B(new_n10729_), .ZN(new_n10730_));
  OAI21_X1   g10538(.A1(new_n10730_), .A2(\asqrt[53] ), .B(new_n10682_), .ZN(new_n10731_));
  NAND3_X1   g10539(.A1(new_n10725_), .A2(new_n10726_), .A3(new_n1305_), .ZN(new_n10732_));
  AOI21_X1   g10540(.A1(new_n10688_), .A2(new_n10732_), .B(new_n10727_), .ZN(new_n10733_));
  AOI21_X1   g10541(.A1(new_n10733_), .A2(new_n1150_), .B(new_n10686_), .ZN(new_n10734_));
  NAND2_X1   g10542(.A1(new_n10732_), .A2(new_n10688_), .ZN(new_n10735_));
  INV_X1     g10543(.I(new_n10727_), .ZN(new_n10736_));
  AOI21_X1   g10544(.A1(new_n10735_), .A2(new_n10736_), .B(new_n1150_), .ZN(new_n10737_));
  OAI21_X1   g10545(.A1(new_n10734_), .A2(new_n10737_), .B(\asqrt[53] ), .ZN(new_n10738_));
  NAND3_X1   g10546(.A1(new_n10731_), .A2(new_n860_), .A3(new_n10738_), .ZN(new_n10739_));
  AOI21_X1   g10547(.A1(new_n10731_), .A2(new_n10738_), .B(new_n860_), .ZN(new_n10740_));
  AOI21_X1   g10548(.A1(new_n10680_), .A2(new_n10739_), .B(new_n10740_), .ZN(new_n10741_));
  AOI21_X1   g10549(.A1(new_n10741_), .A2(new_n744_), .B(new_n10677_), .ZN(new_n10742_));
  INV_X1     g10550(.I(new_n10682_), .ZN(new_n10743_));
  NOR3_X1    g10551(.A1(new_n10734_), .A2(\asqrt[53] ), .A3(new_n10737_), .ZN(new_n10744_));
  OAI21_X1   g10552(.A1(new_n10743_), .A2(new_n10744_), .B(new_n10738_), .ZN(new_n10745_));
  OAI21_X1   g10553(.A1(new_n10745_), .A2(\asqrt[54] ), .B(new_n10680_), .ZN(new_n10746_));
  NAND2_X1   g10554(.A1(new_n10745_), .A2(\asqrt[54] ), .ZN(new_n10747_));
  AOI21_X1   g10555(.A1(new_n10746_), .A2(new_n10747_), .B(new_n744_), .ZN(new_n10748_));
  NOR3_X1    g10556(.A1(new_n10742_), .A2(\asqrt[56] ), .A3(new_n10748_), .ZN(new_n10749_));
  OAI21_X1   g10557(.A1(new_n10742_), .A2(new_n10748_), .B(\asqrt[56] ), .ZN(new_n10750_));
  OAI21_X1   g10558(.A1(new_n10674_), .A2(new_n10749_), .B(new_n10750_), .ZN(new_n10751_));
  OAI21_X1   g10559(.A1(new_n10751_), .A2(\asqrt[57] ), .B(new_n10670_), .ZN(new_n10752_));
  NAND3_X1   g10560(.A1(new_n10746_), .A2(new_n10747_), .A3(new_n744_), .ZN(new_n10753_));
  AOI21_X1   g10561(.A1(new_n10676_), .A2(new_n10753_), .B(new_n10748_), .ZN(new_n10754_));
  AOI21_X1   g10562(.A1(new_n10754_), .A2(new_n634_), .B(new_n10674_), .ZN(new_n10755_));
  NAND2_X1   g10563(.A1(new_n10753_), .A2(new_n10676_), .ZN(new_n10756_));
  INV_X1     g10564(.I(new_n10748_), .ZN(new_n10757_));
  AOI21_X1   g10565(.A1(new_n10756_), .A2(new_n10757_), .B(new_n634_), .ZN(new_n10758_));
  OAI21_X1   g10566(.A1(new_n10755_), .A2(new_n10758_), .B(\asqrt[57] ), .ZN(new_n10759_));
  NAND3_X1   g10567(.A1(new_n10752_), .A2(new_n423_), .A3(new_n10759_), .ZN(new_n10760_));
  AOI21_X1   g10568(.A1(new_n10752_), .A2(new_n10759_), .B(new_n423_), .ZN(new_n10761_));
  AOI21_X1   g10569(.A1(new_n10668_), .A2(new_n10760_), .B(new_n10761_), .ZN(new_n10762_));
  AOI21_X1   g10570(.A1(new_n10762_), .A2(new_n337_), .B(new_n10665_), .ZN(new_n10763_));
  NOR2_X1    g10571(.A1(new_n10762_), .A2(new_n337_), .ZN(new_n10764_));
  NOR3_X1    g10572(.A1(new_n10763_), .A2(new_n10764_), .A3(\asqrt[60] ), .ZN(new_n10765_));
  OAI21_X1   g10573(.A1(new_n10763_), .A2(new_n10764_), .B(\asqrt[60] ), .ZN(new_n10766_));
  OAI21_X1   g10574(.A1(new_n10662_), .A2(new_n10765_), .B(new_n10766_), .ZN(new_n10767_));
  NAND2_X1   g10575(.A1(new_n10767_), .A2(\asqrt[61] ), .ZN(new_n10768_));
  AOI21_X1   g10576(.A1(new_n10373_), .A2(new_n10379_), .B(\asqrt[19] ), .ZN(new_n10769_));
  XOR2_X1    g10577(.A1(new_n10769_), .A2(new_n10232_), .Z(new_n10770_));
  OAI21_X1   g10578(.A1(new_n10767_), .A2(\asqrt[61] ), .B(new_n10770_), .ZN(new_n10771_));
  NAND2_X1   g10579(.A1(new_n10771_), .A2(new_n10768_), .ZN(new_n10772_));
  INV_X1     g10580(.I(new_n10670_), .ZN(new_n10773_));
  NOR3_X1    g10581(.A1(new_n10755_), .A2(\asqrt[57] ), .A3(new_n10758_), .ZN(new_n10774_));
  OAI21_X1   g10582(.A1(new_n10773_), .A2(new_n10774_), .B(new_n10759_), .ZN(new_n10775_));
  OAI21_X1   g10583(.A1(new_n10775_), .A2(\asqrt[58] ), .B(new_n10668_), .ZN(new_n10776_));
  NOR2_X1    g10584(.A1(new_n10774_), .A2(new_n10773_), .ZN(new_n10777_));
  INV_X1     g10585(.I(new_n10759_), .ZN(new_n10778_));
  OAI21_X1   g10586(.A1(new_n10777_), .A2(new_n10778_), .B(\asqrt[58] ), .ZN(new_n10779_));
  NAND3_X1   g10587(.A1(new_n10776_), .A2(new_n337_), .A3(new_n10779_), .ZN(new_n10780_));
  NAND2_X1   g10588(.A1(new_n10780_), .A2(new_n10664_), .ZN(new_n10781_));
  INV_X1     g10589(.I(new_n10668_), .ZN(new_n10782_));
  NOR2_X1    g10590(.A1(new_n10777_), .A2(new_n10778_), .ZN(new_n10783_));
  AOI21_X1   g10591(.A1(new_n10783_), .A2(new_n423_), .B(new_n10782_), .ZN(new_n10784_));
  OAI21_X1   g10592(.A1(new_n10784_), .A2(new_n10761_), .B(\asqrt[59] ), .ZN(new_n10785_));
  NAND3_X1   g10593(.A1(new_n10781_), .A2(new_n266_), .A3(new_n10785_), .ZN(new_n10786_));
  NAND2_X1   g10594(.A1(new_n10786_), .A2(new_n10661_), .ZN(new_n10787_));
  AOI21_X1   g10595(.A1(new_n10787_), .A2(new_n10766_), .B(new_n239_), .ZN(new_n10788_));
  AOI21_X1   g10596(.A1(new_n10781_), .A2(new_n10785_), .B(new_n266_), .ZN(new_n10789_));
  AOI21_X1   g10597(.A1(new_n10661_), .A2(new_n10786_), .B(new_n10789_), .ZN(new_n10790_));
  INV_X1     g10598(.I(new_n10770_), .ZN(new_n10791_));
  AOI21_X1   g10599(.A1(new_n10790_), .A2(new_n239_), .B(new_n10791_), .ZN(new_n10792_));
  OAI21_X1   g10600(.A1(new_n10792_), .A2(new_n10788_), .B(new_n201_), .ZN(new_n10793_));
  NAND3_X1   g10601(.A1(new_n10771_), .A2(new_n10768_), .A3(\asqrt[62] ), .ZN(new_n10794_));
  NOR2_X1    g10602(.A1(new_n10371_), .A2(new_n10380_), .ZN(new_n10795_));
  NOR2_X1    g10603(.A1(\asqrt[19] ), .A2(new_n10795_), .ZN(new_n10796_));
  XOR2_X1    g10604(.A1(new_n10796_), .A2(new_n10369_), .Z(new_n10797_));
  INV_X1     g10605(.I(new_n10797_), .ZN(new_n10798_));
  AOI22_X1   g10606(.A1(new_n10794_), .A2(new_n10793_), .B1(new_n10772_), .B2(new_n10798_), .ZN(new_n10799_));
  NOR2_X1    g10607(.A1(new_n10391_), .A2(new_n10229_), .ZN(new_n10800_));
  OAI21_X1   g10608(.A1(\asqrt[19] ), .A2(new_n10800_), .B(new_n10398_), .ZN(new_n10801_));
  INV_X1     g10609(.I(new_n10801_), .ZN(new_n10802_));
  OAI21_X1   g10610(.A1(new_n10799_), .A2(new_n10659_), .B(new_n10802_), .ZN(new_n10803_));
  OAI21_X1   g10611(.A1(new_n10772_), .A2(\asqrt[62] ), .B(new_n10797_), .ZN(new_n10804_));
  NAND2_X1   g10612(.A1(new_n10772_), .A2(\asqrt[62] ), .ZN(new_n10805_));
  NAND3_X1   g10613(.A1(new_n10804_), .A2(new_n10805_), .A3(new_n10659_), .ZN(new_n10806_));
  NAND2_X1   g10614(.A1(new_n10391_), .A2(new_n10228_), .ZN(new_n10807_));
  NAND2_X1   g10615(.A1(new_n10487_), .A2(new_n10229_), .ZN(new_n10808_));
  AOI21_X1   g10616(.A1(new_n10807_), .A2(new_n10808_), .B(new_n193_), .ZN(new_n10809_));
  OAI21_X1   g10617(.A1(\asqrt[19] ), .A2(new_n10229_), .B(new_n10809_), .ZN(new_n10810_));
  NOR2_X1    g10618(.A1(new_n10404_), .A2(new_n10228_), .ZN(new_n10811_));
  NAND4_X1   g10619(.A1(new_n10395_), .A2(new_n193_), .A3(new_n10398_), .A4(new_n10811_), .ZN(new_n10812_));
  NAND2_X1   g10620(.A1(new_n10810_), .A2(new_n10812_), .ZN(new_n10813_));
  INV_X1     g10621(.I(new_n10813_), .ZN(new_n10814_));
  NAND4_X1   g10622(.A1(new_n10803_), .A2(new_n193_), .A3(new_n10806_), .A4(new_n10814_), .ZN(\asqrt[18] ));
  AOI21_X1   g10623(.A1(new_n10650_), .A2(new_n10654_), .B(\asqrt[18] ), .ZN(new_n10816_));
  XOR2_X1    g10624(.A1(new_n10816_), .A2(new_n10408_), .Z(new_n10817_));
  XOR2_X1    g10625(.A1(new_n10641_), .A2(\asqrt[45] ), .Z(new_n10818_));
  NOR2_X1    g10626(.A1(\asqrt[18] ), .A2(new_n10818_), .ZN(new_n10819_));
  XOR2_X1    g10627(.A1(new_n10819_), .A2(new_n10410_), .Z(new_n10820_));
  NOR2_X1    g10628(.A1(new_n10639_), .A2(new_n10648_), .ZN(new_n10821_));
  NOR2_X1    g10629(.A1(\asqrt[18] ), .A2(new_n10821_), .ZN(new_n10822_));
  XOR2_X1    g10630(.A1(new_n10822_), .A2(new_n10413_), .Z(new_n10823_));
  AOI21_X1   g10631(.A1(new_n10643_), .A2(new_n10647_), .B(\asqrt[18] ), .ZN(new_n10824_));
  XOR2_X1    g10632(.A1(new_n10824_), .A2(new_n10416_), .Z(new_n10825_));
  INV_X1     g10633(.I(new_n10825_), .ZN(new_n10826_));
  AOI21_X1   g10634(.A1(new_n10629_), .A2(new_n10637_), .B(\asqrt[18] ), .ZN(new_n10827_));
  XOR2_X1    g10635(.A1(new_n10827_), .A2(new_n10420_), .Z(new_n10828_));
  INV_X1     g10636(.I(new_n10828_), .ZN(new_n10829_));
  XOR2_X1    g10637(.A1(new_n10620_), .A2(\asqrt[41] ), .Z(new_n10830_));
  NOR2_X1    g10638(.A1(\asqrt[18] ), .A2(new_n10830_), .ZN(new_n10831_));
  XOR2_X1    g10639(.A1(new_n10831_), .A2(new_n10422_), .Z(new_n10832_));
  NOR2_X1    g10640(.A1(new_n10618_), .A2(new_n10627_), .ZN(new_n10833_));
  NOR2_X1    g10641(.A1(\asqrt[18] ), .A2(new_n10833_), .ZN(new_n10834_));
  XOR2_X1    g10642(.A1(new_n10834_), .A2(new_n10425_), .Z(new_n10835_));
  AOI21_X1   g10643(.A1(new_n10622_), .A2(new_n10626_), .B(\asqrt[18] ), .ZN(new_n10836_));
  XOR2_X1    g10644(.A1(new_n10836_), .A2(new_n10428_), .Z(new_n10837_));
  INV_X1     g10645(.I(new_n10837_), .ZN(new_n10838_));
  AOI21_X1   g10646(.A1(new_n10608_), .A2(new_n10616_), .B(\asqrt[18] ), .ZN(new_n10839_));
  XOR2_X1    g10647(.A1(new_n10839_), .A2(new_n10432_), .Z(new_n10840_));
  INV_X1     g10648(.I(new_n10840_), .ZN(new_n10841_));
  XOR2_X1    g10649(.A1(new_n10599_), .A2(\asqrt[37] ), .Z(new_n10842_));
  NOR2_X1    g10650(.A1(\asqrt[18] ), .A2(new_n10842_), .ZN(new_n10843_));
  XOR2_X1    g10651(.A1(new_n10843_), .A2(new_n10434_), .Z(new_n10844_));
  NOR2_X1    g10652(.A1(new_n10597_), .A2(new_n10606_), .ZN(new_n10845_));
  NOR2_X1    g10653(.A1(\asqrt[18] ), .A2(new_n10845_), .ZN(new_n10846_));
  XOR2_X1    g10654(.A1(new_n10846_), .A2(new_n10437_), .Z(new_n10847_));
  AOI21_X1   g10655(.A1(new_n10601_), .A2(new_n10605_), .B(\asqrt[18] ), .ZN(new_n10848_));
  XOR2_X1    g10656(.A1(new_n10848_), .A2(new_n10440_), .Z(new_n10849_));
  INV_X1     g10657(.I(new_n10849_), .ZN(new_n10850_));
  AOI21_X1   g10658(.A1(new_n10587_), .A2(new_n10595_), .B(\asqrt[18] ), .ZN(new_n10851_));
  XOR2_X1    g10659(.A1(new_n10851_), .A2(new_n10444_), .Z(new_n10852_));
  INV_X1     g10660(.I(new_n10852_), .ZN(new_n10853_));
  XOR2_X1    g10661(.A1(new_n10578_), .A2(\asqrt[33] ), .Z(new_n10854_));
  NOR2_X1    g10662(.A1(\asqrt[18] ), .A2(new_n10854_), .ZN(new_n10855_));
  XOR2_X1    g10663(.A1(new_n10855_), .A2(new_n10446_), .Z(new_n10856_));
  NOR2_X1    g10664(.A1(new_n10576_), .A2(new_n10585_), .ZN(new_n10857_));
  NOR2_X1    g10665(.A1(\asqrt[18] ), .A2(new_n10857_), .ZN(new_n10858_));
  XOR2_X1    g10666(.A1(new_n10858_), .A2(new_n10449_), .Z(new_n10859_));
  AOI21_X1   g10667(.A1(new_n10580_), .A2(new_n10584_), .B(\asqrt[18] ), .ZN(new_n10860_));
  XOR2_X1    g10668(.A1(new_n10860_), .A2(new_n10452_), .Z(new_n10861_));
  INV_X1     g10669(.I(new_n10861_), .ZN(new_n10862_));
  AOI21_X1   g10670(.A1(new_n10566_), .A2(new_n10574_), .B(\asqrt[18] ), .ZN(new_n10863_));
  XOR2_X1    g10671(.A1(new_n10863_), .A2(new_n10456_), .Z(new_n10864_));
  INV_X1     g10672(.I(new_n10864_), .ZN(new_n10865_));
  XOR2_X1    g10673(.A1(new_n10557_), .A2(\asqrt[29] ), .Z(new_n10866_));
  NOR2_X1    g10674(.A1(\asqrt[18] ), .A2(new_n10866_), .ZN(new_n10867_));
  XOR2_X1    g10675(.A1(new_n10867_), .A2(new_n10458_), .Z(new_n10868_));
  NOR2_X1    g10676(.A1(new_n10555_), .A2(new_n10564_), .ZN(new_n10869_));
  NOR2_X1    g10677(.A1(\asqrt[18] ), .A2(new_n10869_), .ZN(new_n10870_));
  XOR2_X1    g10678(.A1(new_n10870_), .A2(new_n10461_), .Z(new_n10871_));
  AOI21_X1   g10679(.A1(new_n10559_), .A2(new_n10563_), .B(\asqrt[18] ), .ZN(new_n10872_));
  XOR2_X1    g10680(.A1(new_n10872_), .A2(new_n10464_), .Z(new_n10873_));
  INV_X1     g10681(.I(new_n10873_), .ZN(new_n10874_));
  AOI21_X1   g10682(.A1(new_n10545_), .A2(new_n10553_), .B(\asqrt[18] ), .ZN(new_n10875_));
  XOR2_X1    g10683(.A1(new_n10875_), .A2(new_n10468_), .Z(new_n10876_));
  INV_X1     g10684(.I(new_n10876_), .ZN(new_n10877_));
  XOR2_X1    g10685(.A1(new_n10536_), .A2(\asqrt[25] ), .Z(new_n10878_));
  NOR2_X1    g10686(.A1(\asqrt[18] ), .A2(new_n10878_), .ZN(new_n10879_));
  XOR2_X1    g10687(.A1(new_n10879_), .A2(new_n10470_), .Z(new_n10880_));
  NOR2_X1    g10688(.A1(new_n10534_), .A2(new_n10543_), .ZN(new_n10881_));
  NOR2_X1    g10689(.A1(\asqrt[18] ), .A2(new_n10881_), .ZN(new_n10882_));
  XOR2_X1    g10690(.A1(new_n10882_), .A2(new_n10473_), .Z(new_n10883_));
  AOI21_X1   g10691(.A1(new_n10538_), .A2(new_n10542_), .B(\asqrt[18] ), .ZN(new_n10884_));
  XOR2_X1    g10692(.A1(new_n10884_), .A2(new_n10476_), .Z(new_n10885_));
  INV_X1     g10693(.I(new_n10885_), .ZN(new_n10886_));
  AOI21_X1   g10694(.A1(new_n10524_), .A2(new_n10532_), .B(\asqrt[18] ), .ZN(new_n10887_));
  XOR2_X1    g10695(.A1(new_n10887_), .A2(new_n10483_), .Z(new_n10888_));
  INV_X1     g10696(.I(new_n10888_), .ZN(new_n10889_));
  AOI21_X1   g10697(.A1(new_n10515_), .A2(new_n10523_), .B(\asqrt[18] ), .ZN(new_n10890_));
  XOR2_X1    g10698(.A1(new_n10890_), .A2(new_n10500_), .Z(new_n10891_));
  NAND2_X1   g10699(.A1(\asqrt[19] ), .A2(new_n10501_), .ZN(new_n10892_));
  NOR2_X1    g10700(.A1(new_n10512_), .A2(\a[38] ), .ZN(new_n10893_));
  AOI22_X1   g10701(.A1(new_n10892_), .A2(new_n10512_), .B1(\asqrt[19] ), .B2(new_n10893_), .ZN(new_n10894_));
  AOI21_X1   g10702(.A1(\asqrt[19] ), .A2(\a[38] ), .B(new_n10509_), .ZN(new_n10895_));
  NOR2_X1    g10703(.A1(new_n10519_), .A2(new_n10895_), .ZN(new_n10896_));
  NOR2_X1    g10704(.A1(\asqrt[18] ), .A2(new_n10896_), .ZN(new_n10897_));
  XOR2_X1    g10705(.A1(new_n10897_), .A2(new_n10894_), .Z(new_n10898_));
  NOR2_X1    g10706(.A1(new_n10792_), .A2(new_n10788_), .ZN(new_n10899_));
  AOI21_X1   g10707(.A1(new_n10771_), .A2(new_n10768_), .B(\asqrt[62] ), .ZN(new_n10900_));
  NOR3_X1    g10708(.A1(new_n10792_), .A2(new_n201_), .A3(new_n10788_), .ZN(new_n10901_));
  OAI22_X1   g10709(.A1(new_n10900_), .A2(new_n10901_), .B1(new_n10899_), .B2(new_n10797_), .ZN(new_n10902_));
  AOI21_X1   g10710(.A1(new_n10902_), .A2(new_n10658_), .B(new_n10801_), .ZN(new_n10903_));
  AOI21_X1   g10711(.A1(new_n10899_), .A2(new_n201_), .B(new_n10798_), .ZN(new_n10904_));
  NOR2_X1    g10712(.A1(new_n10899_), .A2(new_n201_), .ZN(new_n10905_));
  NOR3_X1    g10713(.A1(new_n10904_), .A2(new_n10905_), .A3(new_n10658_), .ZN(new_n10906_));
  NOR3_X1    g10714(.A1(new_n10903_), .A2(\asqrt[63] ), .A3(new_n10906_), .ZN(new_n10907_));
  NAND4_X1   g10715(.A1(new_n10907_), .A2(\asqrt[19] ), .A3(new_n10810_), .A4(new_n10812_), .ZN(new_n10908_));
  NAND2_X1   g10716(.A1(\asqrt[18] ), .A2(new_n10502_), .ZN(new_n10909_));
  AOI21_X1   g10717(.A1(new_n10908_), .A2(new_n10909_), .B(\a[38] ), .ZN(new_n10910_));
  NAND2_X1   g10718(.A1(new_n10803_), .A2(new_n193_), .ZN(new_n10911_));
  NAND3_X1   g10719(.A1(new_n10810_), .A2(new_n10812_), .A3(\asqrt[19] ), .ZN(new_n10912_));
  NOR3_X1    g10720(.A1(new_n10911_), .A2(new_n10906_), .A3(new_n10912_), .ZN(new_n10913_));
  NOR4_X1    g10721(.A1(new_n10903_), .A2(\asqrt[63] ), .A3(new_n10906_), .A4(new_n10813_), .ZN(new_n10914_));
  NOR2_X1    g10722(.A1(new_n10914_), .A2(new_n10504_), .ZN(new_n10915_));
  NOR3_X1    g10723(.A1(new_n10915_), .A2(new_n10913_), .A3(new_n10501_), .ZN(new_n10916_));
  OR2_X2     g10724(.A1(new_n10910_), .A2(new_n10916_), .Z(new_n10917_));
  NOR2_X1    g10725(.A1(\a[34] ), .A2(\a[35] ), .ZN(new_n10918_));
  INV_X1     g10726(.I(new_n10918_), .ZN(new_n10919_));
  NAND3_X1   g10727(.A1(\asqrt[18] ), .A2(\a[36] ), .A3(new_n10919_), .ZN(new_n10920_));
  INV_X1     g10728(.I(\a[36] ), .ZN(new_n10921_));
  OAI21_X1   g10729(.A1(\asqrt[18] ), .A2(new_n10921_), .B(new_n10918_), .ZN(new_n10922_));
  AOI21_X1   g10730(.A1(new_n10922_), .A2(new_n10920_), .B(new_n10497_), .ZN(new_n10923_));
  NOR3_X1    g10731(.A1(new_n10488_), .A2(\asqrt[63] ), .A3(new_n10491_), .ZN(new_n10924_));
  NAND2_X1   g10732(.A1(new_n10918_), .A2(new_n10921_), .ZN(new_n10925_));
  NAND3_X1   g10733(.A1(new_n10401_), .A2(new_n10403_), .A3(new_n10925_), .ZN(new_n10926_));
  NAND2_X1   g10734(.A1(new_n10924_), .A2(new_n10926_), .ZN(new_n10927_));
  NAND3_X1   g10735(.A1(\asqrt[18] ), .A2(\a[36] ), .A3(new_n10927_), .ZN(new_n10928_));
  INV_X1     g10736(.I(\a[37] ), .ZN(new_n10929_));
  NAND3_X1   g10737(.A1(\asqrt[18] ), .A2(new_n10921_), .A3(new_n10929_), .ZN(new_n10930_));
  OAI21_X1   g10738(.A1(new_n10914_), .A2(\a[36] ), .B(\a[37] ), .ZN(new_n10931_));
  NAND3_X1   g10739(.A1(new_n10928_), .A2(new_n10931_), .A3(new_n10930_), .ZN(new_n10932_));
  NOR3_X1    g10740(.A1(new_n10932_), .A2(new_n10923_), .A3(\asqrt[20] ), .ZN(new_n10933_));
  OAI21_X1   g10741(.A1(new_n10932_), .A2(new_n10923_), .B(\asqrt[20] ), .ZN(new_n10934_));
  OAI21_X1   g10742(.A1(new_n10917_), .A2(new_n10933_), .B(new_n10934_), .ZN(new_n10935_));
  OAI21_X1   g10743(.A1(new_n10935_), .A2(\asqrt[21] ), .B(new_n10898_), .ZN(new_n10936_));
  NAND2_X1   g10744(.A1(new_n10935_), .A2(\asqrt[21] ), .ZN(new_n10937_));
  NAND3_X1   g10745(.A1(new_n10936_), .A2(new_n10937_), .A3(new_n9233_), .ZN(new_n10938_));
  AOI21_X1   g10746(.A1(new_n10936_), .A2(new_n10937_), .B(new_n9233_), .ZN(new_n10939_));
  AOI21_X1   g10747(.A1(new_n10891_), .A2(new_n10938_), .B(new_n10939_), .ZN(new_n10940_));
  AOI21_X1   g10748(.A1(new_n10940_), .A2(new_n8849_), .B(new_n10889_), .ZN(new_n10941_));
  NAND2_X1   g10749(.A1(new_n10938_), .A2(new_n10891_), .ZN(new_n10942_));
  INV_X1     g10750(.I(new_n10898_), .ZN(new_n10943_));
  NOR2_X1    g10751(.A1(new_n10910_), .A2(new_n10916_), .ZN(new_n10944_));
  NOR3_X1    g10752(.A1(new_n10914_), .A2(new_n10921_), .A3(new_n10918_), .ZN(new_n10945_));
  AOI21_X1   g10753(.A1(new_n10914_), .A2(\a[36] ), .B(new_n10919_), .ZN(new_n10946_));
  OAI21_X1   g10754(.A1(new_n10945_), .A2(new_n10946_), .B(\asqrt[19] ), .ZN(new_n10947_));
  INV_X1     g10755(.I(new_n10927_), .ZN(new_n10948_));
  NOR3_X1    g10756(.A1(new_n10914_), .A2(new_n10921_), .A3(new_n10948_), .ZN(new_n10949_));
  NOR3_X1    g10757(.A1(new_n10914_), .A2(\a[36] ), .A3(\a[37] ), .ZN(new_n10950_));
  AOI21_X1   g10758(.A1(\asqrt[18] ), .A2(new_n10921_), .B(new_n10929_), .ZN(new_n10951_));
  NOR3_X1    g10759(.A1(new_n10949_), .A2(new_n10950_), .A3(new_n10951_), .ZN(new_n10952_));
  NAND3_X1   g10760(.A1(new_n10952_), .A2(new_n10947_), .A3(new_n10052_), .ZN(new_n10953_));
  AOI21_X1   g10761(.A1(new_n10952_), .A2(new_n10947_), .B(new_n10052_), .ZN(new_n10954_));
  AOI21_X1   g10762(.A1(new_n10944_), .A2(new_n10953_), .B(new_n10954_), .ZN(new_n10955_));
  AOI21_X1   g10763(.A1(new_n10955_), .A2(new_n9656_), .B(new_n10943_), .ZN(new_n10956_));
  NAND2_X1   g10764(.A1(new_n10953_), .A2(new_n10944_), .ZN(new_n10957_));
  AOI21_X1   g10765(.A1(new_n10957_), .A2(new_n10934_), .B(new_n9656_), .ZN(new_n10958_));
  OAI21_X1   g10766(.A1(new_n10956_), .A2(new_n10958_), .B(\asqrt[22] ), .ZN(new_n10959_));
  AOI21_X1   g10767(.A1(new_n10942_), .A2(new_n10959_), .B(new_n8849_), .ZN(new_n10960_));
  NOR3_X1    g10768(.A1(new_n10941_), .A2(\asqrt[24] ), .A3(new_n10960_), .ZN(new_n10961_));
  OAI21_X1   g10769(.A1(new_n10941_), .A2(new_n10960_), .B(\asqrt[24] ), .ZN(new_n10962_));
  OAI21_X1   g10770(.A1(new_n10886_), .A2(new_n10961_), .B(new_n10962_), .ZN(new_n10963_));
  OAI21_X1   g10771(.A1(new_n10963_), .A2(\asqrt[25] ), .B(new_n10883_), .ZN(new_n10964_));
  NAND2_X1   g10772(.A1(new_n10963_), .A2(\asqrt[25] ), .ZN(new_n10965_));
  NAND3_X1   g10773(.A1(new_n10964_), .A2(new_n10965_), .A3(new_n7690_), .ZN(new_n10966_));
  AOI21_X1   g10774(.A1(new_n10964_), .A2(new_n10965_), .B(new_n7690_), .ZN(new_n10967_));
  AOI21_X1   g10775(.A1(new_n10880_), .A2(new_n10966_), .B(new_n10967_), .ZN(new_n10968_));
  AOI21_X1   g10776(.A1(new_n10968_), .A2(new_n7331_), .B(new_n10877_), .ZN(new_n10969_));
  NAND2_X1   g10777(.A1(new_n10966_), .A2(new_n10880_), .ZN(new_n10970_));
  INV_X1     g10778(.I(new_n10883_), .ZN(new_n10971_));
  INV_X1     g10779(.I(new_n10891_), .ZN(new_n10972_));
  NOR3_X1    g10780(.A1(new_n10956_), .A2(\asqrt[22] ), .A3(new_n10958_), .ZN(new_n10973_));
  OAI21_X1   g10781(.A1(new_n10972_), .A2(new_n10973_), .B(new_n10959_), .ZN(new_n10974_));
  OAI21_X1   g10782(.A1(new_n10974_), .A2(\asqrt[23] ), .B(new_n10888_), .ZN(new_n10975_));
  NAND2_X1   g10783(.A1(new_n10974_), .A2(\asqrt[23] ), .ZN(new_n10976_));
  NAND3_X1   g10784(.A1(new_n10975_), .A2(new_n10976_), .A3(new_n8440_), .ZN(new_n10977_));
  AOI21_X1   g10785(.A1(new_n10975_), .A2(new_n10976_), .B(new_n8440_), .ZN(new_n10978_));
  AOI21_X1   g10786(.A1(new_n10885_), .A2(new_n10977_), .B(new_n10978_), .ZN(new_n10979_));
  AOI21_X1   g10787(.A1(new_n10979_), .A2(new_n8077_), .B(new_n10971_), .ZN(new_n10980_));
  NAND2_X1   g10788(.A1(new_n10977_), .A2(new_n10885_), .ZN(new_n10981_));
  AOI21_X1   g10789(.A1(new_n10981_), .A2(new_n10962_), .B(new_n8077_), .ZN(new_n10982_));
  OAI21_X1   g10790(.A1(new_n10980_), .A2(new_n10982_), .B(\asqrt[26] ), .ZN(new_n10983_));
  AOI21_X1   g10791(.A1(new_n10970_), .A2(new_n10983_), .B(new_n7331_), .ZN(new_n10984_));
  NOR3_X1    g10792(.A1(new_n10969_), .A2(\asqrt[28] ), .A3(new_n10984_), .ZN(new_n10985_));
  OAI21_X1   g10793(.A1(new_n10969_), .A2(new_n10984_), .B(\asqrt[28] ), .ZN(new_n10986_));
  OAI21_X1   g10794(.A1(new_n10874_), .A2(new_n10985_), .B(new_n10986_), .ZN(new_n10987_));
  OAI21_X1   g10795(.A1(new_n10987_), .A2(\asqrt[29] ), .B(new_n10871_), .ZN(new_n10988_));
  NAND2_X1   g10796(.A1(new_n10987_), .A2(\asqrt[29] ), .ZN(new_n10989_));
  NAND3_X1   g10797(.A1(new_n10988_), .A2(new_n10989_), .A3(new_n6275_), .ZN(new_n10990_));
  AOI21_X1   g10798(.A1(new_n10988_), .A2(new_n10989_), .B(new_n6275_), .ZN(new_n10991_));
  AOI21_X1   g10799(.A1(new_n10868_), .A2(new_n10990_), .B(new_n10991_), .ZN(new_n10992_));
  AOI21_X1   g10800(.A1(new_n10992_), .A2(new_n5947_), .B(new_n10865_), .ZN(new_n10993_));
  NAND2_X1   g10801(.A1(new_n10990_), .A2(new_n10868_), .ZN(new_n10994_));
  INV_X1     g10802(.I(new_n10871_), .ZN(new_n10995_));
  INV_X1     g10803(.I(new_n10880_), .ZN(new_n10996_));
  NOR3_X1    g10804(.A1(new_n10980_), .A2(\asqrt[26] ), .A3(new_n10982_), .ZN(new_n10997_));
  OAI21_X1   g10805(.A1(new_n10996_), .A2(new_n10997_), .B(new_n10983_), .ZN(new_n10998_));
  OAI21_X1   g10806(.A1(new_n10998_), .A2(\asqrt[27] ), .B(new_n10876_), .ZN(new_n10999_));
  NAND2_X1   g10807(.A1(new_n10998_), .A2(\asqrt[27] ), .ZN(new_n11000_));
  NAND3_X1   g10808(.A1(new_n10999_), .A2(new_n11000_), .A3(new_n6966_), .ZN(new_n11001_));
  AOI21_X1   g10809(.A1(new_n10999_), .A2(new_n11000_), .B(new_n6966_), .ZN(new_n11002_));
  AOI21_X1   g10810(.A1(new_n10873_), .A2(new_n11001_), .B(new_n11002_), .ZN(new_n11003_));
  AOI21_X1   g10811(.A1(new_n11003_), .A2(new_n6636_), .B(new_n10995_), .ZN(new_n11004_));
  NAND2_X1   g10812(.A1(new_n11001_), .A2(new_n10873_), .ZN(new_n11005_));
  AOI21_X1   g10813(.A1(new_n11005_), .A2(new_n10986_), .B(new_n6636_), .ZN(new_n11006_));
  OAI21_X1   g10814(.A1(new_n11004_), .A2(new_n11006_), .B(\asqrt[30] ), .ZN(new_n11007_));
  AOI21_X1   g10815(.A1(new_n10994_), .A2(new_n11007_), .B(new_n5947_), .ZN(new_n11008_));
  NOR3_X1    g10816(.A1(new_n10993_), .A2(\asqrt[32] ), .A3(new_n11008_), .ZN(new_n11009_));
  OAI21_X1   g10817(.A1(new_n10993_), .A2(new_n11008_), .B(\asqrt[32] ), .ZN(new_n11010_));
  OAI21_X1   g10818(.A1(new_n10862_), .A2(new_n11009_), .B(new_n11010_), .ZN(new_n11011_));
  OAI21_X1   g10819(.A1(new_n11011_), .A2(\asqrt[33] ), .B(new_n10859_), .ZN(new_n11012_));
  NAND2_X1   g10820(.A1(new_n11011_), .A2(\asqrt[33] ), .ZN(new_n11013_));
  NAND3_X1   g10821(.A1(new_n11012_), .A2(new_n11013_), .A3(new_n5029_), .ZN(new_n11014_));
  AOI21_X1   g10822(.A1(new_n11012_), .A2(new_n11013_), .B(new_n5029_), .ZN(new_n11015_));
  AOI21_X1   g10823(.A1(new_n10856_), .A2(new_n11014_), .B(new_n11015_), .ZN(new_n11016_));
  AOI21_X1   g10824(.A1(new_n11016_), .A2(new_n4751_), .B(new_n10853_), .ZN(new_n11017_));
  NAND2_X1   g10825(.A1(new_n11014_), .A2(new_n10856_), .ZN(new_n11018_));
  INV_X1     g10826(.I(new_n10859_), .ZN(new_n11019_));
  INV_X1     g10827(.I(new_n10868_), .ZN(new_n11020_));
  NOR3_X1    g10828(.A1(new_n11004_), .A2(\asqrt[30] ), .A3(new_n11006_), .ZN(new_n11021_));
  OAI21_X1   g10829(.A1(new_n11020_), .A2(new_n11021_), .B(new_n11007_), .ZN(new_n11022_));
  OAI21_X1   g10830(.A1(new_n11022_), .A2(\asqrt[31] ), .B(new_n10864_), .ZN(new_n11023_));
  NAND2_X1   g10831(.A1(new_n11022_), .A2(\asqrt[31] ), .ZN(new_n11024_));
  NAND3_X1   g10832(.A1(new_n11023_), .A2(new_n11024_), .A3(new_n5643_), .ZN(new_n11025_));
  AOI21_X1   g10833(.A1(new_n11023_), .A2(new_n11024_), .B(new_n5643_), .ZN(new_n11026_));
  AOI21_X1   g10834(.A1(new_n10861_), .A2(new_n11025_), .B(new_n11026_), .ZN(new_n11027_));
  AOI21_X1   g10835(.A1(new_n11027_), .A2(new_n5336_), .B(new_n11019_), .ZN(new_n11028_));
  NAND2_X1   g10836(.A1(new_n11025_), .A2(new_n10861_), .ZN(new_n11029_));
  AOI21_X1   g10837(.A1(new_n11029_), .A2(new_n11010_), .B(new_n5336_), .ZN(new_n11030_));
  OAI21_X1   g10838(.A1(new_n11028_), .A2(new_n11030_), .B(\asqrt[34] ), .ZN(new_n11031_));
  AOI21_X1   g10839(.A1(new_n11018_), .A2(new_n11031_), .B(new_n4751_), .ZN(new_n11032_));
  NOR3_X1    g10840(.A1(new_n11017_), .A2(\asqrt[36] ), .A3(new_n11032_), .ZN(new_n11033_));
  OAI21_X1   g10841(.A1(new_n11017_), .A2(new_n11032_), .B(\asqrt[36] ), .ZN(new_n11034_));
  OAI21_X1   g10842(.A1(new_n10850_), .A2(new_n11033_), .B(new_n11034_), .ZN(new_n11035_));
  OAI21_X1   g10843(.A1(new_n11035_), .A2(\asqrt[37] ), .B(new_n10847_), .ZN(new_n11036_));
  NAND2_X1   g10844(.A1(new_n11035_), .A2(\asqrt[37] ), .ZN(new_n11037_));
  NAND3_X1   g10845(.A1(new_n11036_), .A2(new_n11037_), .A3(new_n3925_), .ZN(new_n11038_));
  AOI21_X1   g10846(.A1(new_n11036_), .A2(new_n11037_), .B(new_n3925_), .ZN(new_n11039_));
  AOI21_X1   g10847(.A1(new_n10844_), .A2(new_n11038_), .B(new_n11039_), .ZN(new_n11040_));
  AOI21_X1   g10848(.A1(new_n11040_), .A2(new_n3681_), .B(new_n10841_), .ZN(new_n11041_));
  NAND2_X1   g10849(.A1(new_n11038_), .A2(new_n10844_), .ZN(new_n11042_));
  INV_X1     g10850(.I(new_n10847_), .ZN(new_n11043_));
  INV_X1     g10851(.I(new_n10856_), .ZN(new_n11044_));
  NOR3_X1    g10852(.A1(new_n11028_), .A2(\asqrt[34] ), .A3(new_n11030_), .ZN(new_n11045_));
  OAI21_X1   g10853(.A1(new_n11044_), .A2(new_n11045_), .B(new_n11031_), .ZN(new_n11046_));
  OAI21_X1   g10854(.A1(new_n11046_), .A2(\asqrt[35] ), .B(new_n10852_), .ZN(new_n11047_));
  NAND2_X1   g10855(.A1(new_n11046_), .A2(\asqrt[35] ), .ZN(new_n11048_));
  NAND3_X1   g10856(.A1(new_n11047_), .A2(new_n11048_), .A3(new_n4461_), .ZN(new_n11049_));
  AOI21_X1   g10857(.A1(new_n11047_), .A2(new_n11048_), .B(new_n4461_), .ZN(new_n11050_));
  AOI21_X1   g10858(.A1(new_n10849_), .A2(new_n11049_), .B(new_n11050_), .ZN(new_n11051_));
  AOI21_X1   g10859(.A1(new_n11051_), .A2(new_n4196_), .B(new_n11043_), .ZN(new_n11052_));
  NAND2_X1   g10860(.A1(new_n11049_), .A2(new_n10849_), .ZN(new_n11053_));
  AOI21_X1   g10861(.A1(new_n11053_), .A2(new_n11034_), .B(new_n4196_), .ZN(new_n11054_));
  OAI21_X1   g10862(.A1(new_n11052_), .A2(new_n11054_), .B(\asqrt[38] ), .ZN(new_n11055_));
  AOI21_X1   g10863(.A1(new_n11042_), .A2(new_n11055_), .B(new_n3681_), .ZN(new_n11056_));
  NOR3_X1    g10864(.A1(new_n11041_), .A2(\asqrt[40] ), .A3(new_n11056_), .ZN(new_n11057_));
  OAI21_X1   g10865(.A1(new_n11041_), .A2(new_n11056_), .B(\asqrt[40] ), .ZN(new_n11058_));
  OAI21_X1   g10866(.A1(new_n10838_), .A2(new_n11057_), .B(new_n11058_), .ZN(new_n11059_));
  OAI21_X1   g10867(.A1(new_n11059_), .A2(\asqrt[41] ), .B(new_n10835_), .ZN(new_n11060_));
  NAND2_X1   g10868(.A1(new_n11059_), .A2(\asqrt[41] ), .ZN(new_n11061_));
  NAND3_X1   g10869(.A1(new_n11060_), .A2(new_n11061_), .A3(new_n2960_), .ZN(new_n11062_));
  AOI21_X1   g10870(.A1(new_n11060_), .A2(new_n11061_), .B(new_n2960_), .ZN(new_n11063_));
  AOI21_X1   g10871(.A1(new_n10832_), .A2(new_n11062_), .B(new_n11063_), .ZN(new_n11064_));
  AOI21_X1   g10872(.A1(new_n11064_), .A2(new_n2749_), .B(new_n10829_), .ZN(new_n11065_));
  NAND2_X1   g10873(.A1(new_n11062_), .A2(new_n10832_), .ZN(new_n11066_));
  INV_X1     g10874(.I(new_n10835_), .ZN(new_n11067_));
  INV_X1     g10875(.I(new_n10844_), .ZN(new_n11068_));
  NOR3_X1    g10876(.A1(new_n11052_), .A2(\asqrt[38] ), .A3(new_n11054_), .ZN(new_n11069_));
  OAI21_X1   g10877(.A1(new_n11068_), .A2(new_n11069_), .B(new_n11055_), .ZN(new_n11070_));
  OAI21_X1   g10878(.A1(new_n11070_), .A2(\asqrt[39] ), .B(new_n10840_), .ZN(new_n11071_));
  NAND2_X1   g10879(.A1(new_n11070_), .A2(\asqrt[39] ), .ZN(new_n11072_));
  NAND3_X1   g10880(.A1(new_n11071_), .A2(new_n11072_), .A3(new_n3427_), .ZN(new_n11073_));
  AOI21_X1   g10881(.A1(new_n11071_), .A2(new_n11072_), .B(new_n3427_), .ZN(new_n11074_));
  AOI21_X1   g10882(.A1(new_n10837_), .A2(new_n11073_), .B(new_n11074_), .ZN(new_n11075_));
  AOI21_X1   g10883(.A1(new_n11075_), .A2(new_n3195_), .B(new_n11067_), .ZN(new_n11076_));
  NAND2_X1   g10884(.A1(new_n11073_), .A2(new_n10837_), .ZN(new_n11077_));
  AOI21_X1   g10885(.A1(new_n11077_), .A2(new_n11058_), .B(new_n3195_), .ZN(new_n11078_));
  OAI21_X1   g10886(.A1(new_n11076_), .A2(new_n11078_), .B(\asqrt[42] ), .ZN(new_n11079_));
  AOI21_X1   g10887(.A1(new_n11066_), .A2(new_n11079_), .B(new_n2749_), .ZN(new_n11080_));
  NOR3_X1    g10888(.A1(new_n11065_), .A2(\asqrt[44] ), .A3(new_n11080_), .ZN(new_n11081_));
  OAI21_X1   g10889(.A1(new_n11065_), .A2(new_n11080_), .B(\asqrt[44] ), .ZN(new_n11082_));
  OAI21_X1   g10890(.A1(new_n10826_), .A2(new_n11081_), .B(new_n11082_), .ZN(new_n11083_));
  OAI21_X1   g10891(.A1(new_n11083_), .A2(\asqrt[45] ), .B(new_n10823_), .ZN(new_n11084_));
  NAND2_X1   g10892(.A1(new_n11083_), .A2(\asqrt[45] ), .ZN(new_n11085_));
  NAND3_X1   g10893(.A1(new_n11084_), .A2(new_n11085_), .A3(new_n2134_), .ZN(new_n11086_));
  AOI21_X1   g10894(.A1(new_n11084_), .A2(new_n11085_), .B(new_n2134_), .ZN(new_n11087_));
  AOI21_X1   g10895(.A1(new_n10820_), .A2(new_n11086_), .B(new_n11087_), .ZN(new_n11088_));
  NAND2_X1   g10896(.A1(new_n11088_), .A2(new_n1953_), .ZN(new_n11089_));
  INV_X1     g10897(.I(new_n10820_), .ZN(new_n11090_));
  INV_X1     g10898(.I(new_n10823_), .ZN(new_n11091_));
  INV_X1     g10899(.I(new_n10832_), .ZN(new_n11092_));
  NOR3_X1    g10900(.A1(new_n11076_), .A2(\asqrt[42] ), .A3(new_n11078_), .ZN(new_n11093_));
  OAI21_X1   g10901(.A1(new_n11092_), .A2(new_n11093_), .B(new_n11079_), .ZN(new_n11094_));
  OAI21_X1   g10902(.A1(new_n11094_), .A2(\asqrt[43] ), .B(new_n10828_), .ZN(new_n11095_));
  NAND2_X1   g10903(.A1(new_n11094_), .A2(\asqrt[43] ), .ZN(new_n11096_));
  NAND3_X1   g10904(.A1(new_n11095_), .A2(new_n11096_), .A3(new_n2531_), .ZN(new_n11097_));
  AOI21_X1   g10905(.A1(new_n11095_), .A2(new_n11096_), .B(new_n2531_), .ZN(new_n11098_));
  AOI21_X1   g10906(.A1(new_n10825_), .A2(new_n11097_), .B(new_n11098_), .ZN(new_n11099_));
  AOI21_X1   g10907(.A1(new_n11099_), .A2(new_n2332_), .B(new_n11091_), .ZN(new_n11100_));
  NAND2_X1   g10908(.A1(new_n11097_), .A2(new_n10825_), .ZN(new_n11101_));
  AOI21_X1   g10909(.A1(new_n11101_), .A2(new_n11082_), .B(new_n2332_), .ZN(new_n11102_));
  NOR3_X1    g10910(.A1(new_n11100_), .A2(\asqrt[46] ), .A3(new_n11102_), .ZN(new_n11103_));
  OAI21_X1   g10911(.A1(new_n11100_), .A2(new_n11102_), .B(\asqrt[46] ), .ZN(new_n11104_));
  OAI21_X1   g10912(.A1(new_n11090_), .A2(new_n11103_), .B(new_n11104_), .ZN(new_n11105_));
  NAND2_X1   g10913(.A1(new_n11105_), .A2(\asqrt[47] ), .ZN(new_n11106_));
  NOR2_X1    g10914(.A1(new_n10772_), .A2(\asqrt[62] ), .ZN(new_n11107_));
  NOR2_X1    g10915(.A1(new_n11107_), .A2(new_n10905_), .ZN(new_n11108_));
  XOR2_X1    g10916(.A1(new_n10796_), .A2(new_n10369_), .Z(new_n11109_));
  OAI21_X1   g10917(.A1(\asqrt[18] ), .A2(new_n11108_), .B(new_n11109_), .ZN(new_n11110_));
  INV_X1     g10918(.I(new_n11110_), .ZN(new_n11111_));
  AOI21_X1   g10919(.A1(new_n10780_), .A2(new_n10785_), .B(\asqrt[18] ), .ZN(new_n11112_));
  XOR2_X1    g10920(.A1(new_n11112_), .A2(new_n10664_), .Z(new_n11113_));
  INV_X1     g10921(.I(new_n11113_), .ZN(new_n11114_));
  AOI21_X1   g10922(.A1(new_n10760_), .A2(new_n10779_), .B(\asqrt[18] ), .ZN(new_n11115_));
  XOR2_X1    g10923(.A1(new_n11115_), .A2(new_n10668_), .Z(new_n11116_));
  INV_X1     g10924(.I(new_n11116_), .ZN(new_n11117_));
  NOR2_X1    g10925(.A1(new_n10778_), .A2(new_n10774_), .ZN(new_n11118_));
  NOR2_X1    g10926(.A1(\asqrt[18] ), .A2(new_n11118_), .ZN(new_n11119_));
  XOR2_X1    g10927(.A1(new_n11119_), .A2(new_n10670_), .Z(new_n11120_));
  NOR2_X1    g10928(.A1(new_n10749_), .A2(new_n10758_), .ZN(new_n11121_));
  NOR2_X1    g10929(.A1(\asqrt[18] ), .A2(new_n11121_), .ZN(new_n11122_));
  XOR2_X1    g10930(.A1(new_n11122_), .A2(new_n10673_), .Z(new_n11123_));
  AOI21_X1   g10931(.A1(new_n10753_), .A2(new_n10757_), .B(\asqrt[18] ), .ZN(new_n11124_));
  XOR2_X1    g10932(.A1(new_n11124_), .A2(new_n10676_), .Z(new_n11125_));
  INV_X1     g10933(.I(new_n11125_), .ZN(new_n11126_));
  AOI21_X1   g10934(.A1(new_n10739_), .A2(new_n10747_), .B(\asqrt[18] ), .ZN(new_n11127_));
  XOR2_X1    g10935(.A1(new_n11127_), .A2(new_n10680_), .Z(new_n11128_));
  INV_X1     g10936(.I(new_n11128_), .ZN(new_n11129_));
  XOR2_X1    g10937(.A1(new_n10730_), .A2(\asqrt[53] ), .Z(new_n11130_));
  NOR2_X1    g10938(.A1(\asqrt[18] ), .A2(new_n11130_), .ZN(new_n11131_));
  XOR2_X1    g10939(.A1(new_n11131_), .A2(new_n10682_), .Z(new_n11132_));
  NOR2_X1    g10940(.A1(new_n10728_), .A2(new_n10737_), .ZN(new_n11133_));
  NOR2_X1    g10941(.A1(\asqrt[18] ), .A2(new_n11133_), .ZN(new_n11134_));
  XOR2_X1    g10942(.A1(new_n11134_), .A2(new_n10685_), .Z(new_n11135_));
  AOI21_X1   g10943(.A1(new_n10732_), .A2(new_n10736_), .B(\asqrt[18] ), .ZN(new_n11136_));
  XOR2_X1    g10944(.A1(new_n11136_), .A2(new_n10688_), .Z(new_n11137_));
  INV_X1     g10945(.I(new_n11137_), .ZN(new_n11138_));
  AOI21_X1   g10946(.A1(new_n10718_), .A2(new_n10726_), .B(\asqrt[18] ), .ZN(new_n11139_));
  XOR2_X1    g10947(.A1(new_n11139_), .A2(new_n10692_), .Z(new_n11140_));
  INV_X1     g10948(.I(new_n11140_), .ZN(new_n11141_));
  XOR2_X1    g10949(.A1(new_n10709_), .A2(\asqrt[49] ), .Z(new_n11142_));
  NOR2_X1    g10950(.A1(\asqrt[18] ), .A2(new_n11142_), .ZN(new_n11143_));
  XOR2_X1    g10951(.A1(new_n11143_), .A2(new_n10694_), .Z(new_n11144_));
  NOR2_X1    g10952(.A1(new_n10707_), .A2(new_n10716_), .ZN(new_n11145_));
  NOR2_X1    g10953(.A1(\asqrt[18] ), .A2(new_n11145_), .ZN(new_n11146_));
  XOR2_X1    g10954(.A1(new_n11146_), .A2(new_n10697_), .Z(new_n11147_));
  AOI21_X1   g10955(.A1(new_n10711_), .A2(new_n10715_), .B(\asqrt[18] ), .ZN(new_n11148_));
  XOR2_X1    g10956(.A1(new_n11148_), .A2(new_n10700_), .Z(new_n11149_));
  INV_X1     g10957(.I(new_n11149_), .ZN(new_n11150_));
  INV_X1     g10958(.I(new_n10817_), .ZN(new_n11151_));
  AOI21_X1   g10959(.A1(new_n11088_), .A2(new_n1953_), .B(new_n11151_), .ZN(new_n11152_));
  NAND2_X1   g10960(.A1(new_n11086_), .A2(new_n10820_), .ZN(new_n11153_));
  AOI21_X1   g10961(.A1(new_n11153_), .A2(new_n11104_), .B(new_n1953_), .ZN(new_n11154_));
  NOR3_X1    g10962(.A1(new_n11152_), .A2(\asqrt[48] ), .A3(new_n11154_), .ZN(new_n11155_));
  OAI21_X1   g10963(.A1(new_n11152_), .A2(new_n11154_), .B(\asqrt[48] ), .ZN(new_n11156_));
  OAI21_X1   g10964(.A1(new_n11150_), .A2(new_n11155_), .B(new_n11156_), .ZN(new_n11157_));
  OAI21_X1   g10965(.A1(new_n11157_), .A2(\asqrt[49] ), .B(new_n11147_), .ZN(new_n11158_));
  NAND2_X1   g10966(.A1(new_n11157_), .A2(\asqrt[49] ), .ZN(new_n11159_));
  NAND3_X1   g10967(.A1(new_n11158_), .A2(new_n11159_), .A3(new_n1463_), .ZN(new_n11160_));
  AOI21_X1   g10968(.A1(new_n11158_), .A2(new_n11159_), .B(new_n1463_), .ZN(new_n11161_));
  AOI21_X1   g10969(.A1(new_n11144_), .A2(new_n11160_), .B(new_n11161_), .ZN(new_n11162_));
  AOI21_X1   g10970(.A1(new_n11162_), .A2(new_n1305_), .B(new_n11141_), .ZN(new_n11163_));
  NAND2_X1   g10971(.A1(new_n11160_), .A2(new_n11144_), .ZN(new_n11164_));
  INV_X1     g10972(.I(new_n11147_), .ZN(new_n11165_));
  OAI21_X1   g10973(.A1(new_n11105_), .A2(\asqrt[47] ), .B(new_n10817_), .ZN(new_n11166_));
  NAND3_X1   g10974(.A1(new_n11166_), .A2(new_n11106_), .A3(new_n1778_), .ZN(new_n11167_));
  AOI21_X1   g10975(.A1(new_n11166_), .A2(new_n11106_), .B(new_n1778_), .ZN(new_n11168_));
  AOI21_X1   g10976(.A1(new_n11149_), .A2(new_n11167_), .B(new_n11168_), .ZN(new_n11169_));
  AOI21_X1   g10977(.A1(new_n11169_), .A2(new_n1632_), .B(new_n11165_), .ZN(new_n11170_));
  NAND2_X1   g10978(.A1(new_n11167_), .A2(new_n11149_), .ZN(new_n11171_));
  AOI21_X1   g10979(.A1(new_n11171_), .A2(new_n11156_), .B(new_n1632_), .ZN(new_n11172_));
  OAI21_X1   g10980(.A1(new_n11170_), .A2(new_n11172_), .B(\asqrt[50] ), .ZN(new_n11173_));
  AOI21_X1   g10981(.A1(new_n11164_), .A2(new_n11173_), .B(new_n1305_), .ZN(new_n11174_));
  NOR3_X1    g10982(.A1(new_n11163_), .A2(\asqrt[52] ), .A3(new_n11174_), .ZN(new_n11175_));
  OAI21_X1   g10983(.A1(new_n11163_), .A2(new_n11174_), .B(\asqrt[52] ), .ZN(new_n11176_));
  OAI21_X1   g10984(.A1(new_n11138_), .A2(new_n11175_), .B(new_n11176_), .ZN(new_n11177_));
  OAI21_X1   g10985(.A1(new_n11177_), .A2(\asqrt[53] ), .B(new_n11135_), .ZN(new_n11178_));
  NAND2_X1   g10986(.A1(new_n11177_), .A2(\asqrt[53] ), .ZN(new_n11179_));
  NAND3_X1   g10987(.A1(new_n11178_), .A2(new_n11179_), .A3(new_n860_), .ZN(new_n11180_));
  AOI21_X1   g10988(.A1(new_n11178_), .A2(new_n11179_), .B(new_n860_), .ZN(new_n11181_));
  AOI21_X1   g10989(.A1(new_n11132_), .A2(new_n11180_), .B(new_n11181_), .ZN(new_n11182_));
  AOI21_X1   g10990(.A1(new_n11182_), .A2(new_n744_), .B(new_n11129_), .ZN(new_n11183_));
  NAND2_X1   g10991(.A1(new_n11180_), .A2(new_n11132_), .ZN(new_n11184_));
  INV_X1     g10992(.I(new_n11135_), .ZN(new_n11185_));
  INV_X1     g10993(.I(new_n11144_), .ZN(new_n11186_));
  NOR3_X1    g10994(.A1(new_n11170_), .A2(\asqrt[50] ), .A3(new_n11172_), .ZN(new_n11187_));
  OAI21_X1   g10995(.A1(new_n11186_), .A2(new_n11187_), .B(new_n11173_), .ZN(new_n11188_));
  OAI21_X1   g10996(.A1(new_n11188_), .A2(\asqrt[51] ), .B(new_n11140_), .ZN(new_n11189_));
  NAND2_X1   g10997(.A1(new_n11188_), .A2(\asqrt[51] ), .ZN(new_n11190_));
  NAND3_X1   g10998(.A1(new_n11189_), .A2(new_n11190_), .A3(new_n1150_), .ZN(new_n11191_));
  AOI21_X1   g10999(.A1(new_n11189_), .A2(new_n11190_), .B(new_n1150_), .ZN(new_n11192_));
  AOI21_X1   g11000(.A1(new_n11137_), .A2(new_n11191_), .B(new_n11192_), .ZN(new_n11193_));
  AOI21_X1   g11001(.A1(new_n11193_), .A2(new_n1006_), .B(new_n11185_), .ZN(new_n11194_));
  NAND2_X1   g11002(.A1(new_n11191_), .A2(new_n11137_), .ZN(new_n11195_));
  AOI21_X1   g11003(.A1(new_n11195_), .A2(new_n11176_), .B(new_n1006_), .ZN(new_n11196_));
  OAI21_X1   g11004(.A1(new_n11194_), .A2(new_n11196_), .B(\asqrt[54] ), .ZN(new_n11197_));
  AOI21_X1   g11005(.A1(new_n11184_), .A2(new_n11197_), .B(new_n744_), .ZN(new_n11198_));
  NOR3_X1    g11006(.A1(new_n11183_), .A2(\asqrt[56] ), .A3(new_n11198_), .ZN(new_n11199_));
  OAI21_X1   g11007(.A1(new_n11183_), .A2(new_n11198_), .B(\asqrt[56] ), .ZN(new_n11200_));
  OAI21_X1   g11008(.A1(new_n11126_), .A2(new_n11199_), .B(new_n11200_), .ZN(new_n11201_));
  OAI21_X1   g11009(.A1(new_n11201_), .A2(\asqrt[57] ), .B(new_n11123_), .ZN(new_n11202_));
  NAND2_X1   g11010(.A1(new_n11201_), .A2(\asqrt[57] ), .ZN(new_n11203_));
  NAND3_X1   g11011(.A1(new_n11202_), .A2(new_n11203_), .A3(new_n423_), .ZN(new_n11204_));
  AOI21_X1   g11012(.A1(new_n11202_), .A2(new_n11203_), .B(new_n423_), .ZN(new_n11205_));
  AOI21_X1   g11013(.A1(new_n11120_), .A2(new_n11204_), .B(new_n11205_), .ZN(new_n11206_));
  AOI21_X1   g11014(.A1(new_n11206_), .A2(new_n337_), .B(new_n11117_), .ZN(new_n11207_));
  NAND2_X1   g11015(.A1(new_n11204_), .A2(new_n11120_), .ZN(new_n11208_));
  INV_X1     g11016(.I(new_n11123_), .ZN(new_n11209_));
  INV_X1     g11017(.I(new_n11132_), .ZN(new_n11210_));
  NOR3_X1    g11018(.A1(new_n11194_), .A2(\asqrt[54] ), .A3(new_n11196_), .ZN(new_n11211_));
  OAI21_X1   g11019(.A1(new_n11210_), .A2(new_n11211_), .B(new_n11197_), .ZN(new_n11212_));
  OAI21_X1   g11020(.A1(new_n11212_), .A2(\asqrt[55] ), .B(new_n11128_), .ZN(new_n11213_));
  NAND2_X1   g11021(.A1(new_n11212_), .A2(\asqrt[55] ), .ZN(new_n11214_));
  NAND3_X1   g11022(.A1(new_n11213_), .A2(new_n11214_), .A3(new_n634_), .ZN(new_n11215_));
  AOI21_X1   g11023(.A1(new_n11213_), .A2(new_n11214_), .B(new_n634_), .ZN(new_n11216_));
  AOI21_X1   g11024(.A1(new_n11125_), .A2(new_n11215_), .B(new_n11216_), .ZN(new_n11217_));
  AOI21_X1   g11025(.A1(new_n11217_), .A2(new_n531_), .B(new_n11209_), .ZN(new_n11218_));
  NAND2_X1   g11026(.A1(new_n11215_), .A2(new_n11125_), .ZN(new_n11219_));
  AOI21_X1   g11027(.A1(new_n11219_), .A2(new_n11200_), .B(new_n531_), .ZN(new_n11220_));
  OAI21_X1   g11028(.A1(new_n11218_), .A2(new_n11220_), .B(\asqrt[58] ), .ZN(new_n11221_));
  AOI21_X1   g11029(.A1(new_n11208_), .A2(new_n11221_), .B(new_n337_), .ZN(new_n11222_));
  NOR3_X1    g11030(.A1(new_n11207_), .A2(\asqrt[60] ), .A3(new_n11222_), .ZN(new_n11223_));
  NOR2_X1    g11031(.A1(new_n11223_), .A2(new_n11114_), .ZN(new_n11224_));
  INV_X1     g11032(.I(new_n11120_), .ZN(new_n11225_));
  NOR3_X1    g11033(.A1(new_n11218_), .A2(\asqrt[58] ), .A3(new_n11220_), .ZN(new_n11226_));
  OAI21_X1   g11034(.A1(new_n11225_), .A2(new_n11226_), .B(new_n11221_), .ZN(new_n11227_));
  OAI21_X1   g11035(.A1(new_n11227_), .A2(\asqrt[59] ), .B(new_n11116_), .ZN(new_n11228_));
  NOR2_X1    g11036(.A1(new_n11226_), .A2(new_n11225_), .ZN(new_n11229_));
  OAI21_X1   g11037(.A1(new_n11229_), .A2(new_n11205_), .B(\asqrt[59] ), .ZN(new_n11230_));
  AOI21_X1   g11038(.A1(new_n11228_), .A2(new_n11230_), .B(new_n266_), .ZN(new_n11231_));
  OAI21_X1   g11039(.A1(new_n11224_), .A2(new_n11231_), .B(\asqrt[61] ), .ZN(new_n11232_));
  OAI21_X1   g11040(.A1(new_n11207_), .A2(new_n11222_), .B(\asqrt[60] ), .ZN(new_n11233_));
  OAI21_X1   g11041(.A1(new_n11114_), .A2(new_n11223_), .B(new_n11233_), .ZN(new_n11234_));
  AOI21_X1   g11042(.A1(new_n10786_), .A2(new_n10766_), .B(\asqrt[18] ), .ZN(new_n11235_));
  XOR2_X1    g11043(.A1(new_n11235_), .A2(new_n10661_), .Z(new_n11236_));
  OAI21_X1   g11044(.A1(new_n11234_), .A2(\asqrt[61] ), .B(new_n11236_), .ZN(new_n11237_));
  NAND2_X1   g11045(.A1(new_n11237_), .A2(new_n11232_), .ZN(new_n11238_));
  NAND3_X1   g11046(.A1(new_n11228_), .A2(new_n266_), .A3(new_n11230_), .ZN(new_n11239_));
  NAND2_X1   g11047(.A1(new_n11239_), .A2(new_n11113_), .ZN(new_n11240_));
  AOI21_X1   g11048(.A1(new_n11240_), .A2(new_n11233_), .B(new_n239_), .ZN(new_n11241_));
  AOI21_X1   g11049(.A1(new_n11113_), .A2(new_n11239_), .B(new_n11231_), .ZN(new_n11242_));
  INV_X1     g11050(.I(new_n11236_), .ZN(new_n11243_));
  AOI21_X1   g11051(.A1(new_n11242_), .A2(new_n239_), .B(new_n11243_), .ZN(new_n11244_));
  OAI21_X1   g11052(.A1(new_n11244_), .A2(new_n11241_), .B(new_n201_), .ZN(new_n11245_));
  NAND3_X1   g11053(.A1(new_n11237_), .A2(\asqrt[62] ), .A3(new_n11232_), .ZN(new_n11246_));
  NAND2_X1   g11054(.A1(new_n10790_), .A2(new_n239_), .ZN(new_n11247_));
  AOI21_X1   g11055(.A1(new_n10768_), .A2(new_n11247_), .B(\asqrt[18] ), .ZN(new_n11248_));
  XOR2_X1    g11056(.A1(new_n11248_), .A2(new_n10770_), .Z(new_n11249_));
  INV_X1     g11057(.I(new_n11249_), .ZN(new_n11250_));
  AOI22_X1   g11058(.A1(new_n11245_), .A2(new_n11246_), .B1(new_n11238_), .B2(new_n11250_), .ZN(new_n11251_));
  NOR2_X1    g11059(.A1(new_n10799_), .A2(new_n10659_), .ZN(new_n11252_));
  OAI21_X1   g11060(.A1(\asqrt[18] ), .A2(new_n11252_), .B(new_n10806_), .ZN(new_n11253_));
  INV_X1     g11061(.I(new_n11253_), .ZN(new_n11254_));
  OAI21_X1   g11062(.A1(new_n11251_), .A2(new_n11111_), .B(new_n11254_), .ZN(new_n11255_));
  OAI21_X1   g11063(.A1(new_n11238_), .A2(\asqrt[62] ), .B(new_n11249_), .ZN(new_n11256_));
  NAND2_X1   g11064(.A1(new_n11238_), .A2(\asqrt[62] ), .ZN(new_n11257_));
  NAND3_X1   g11065(.A1(new_n11256_), .A2(new_n11257_), .A3(new_n11111_), .ZN(new_n11258_));
  NAND2_X1   g11066(.A1(new_n10914_), .A2(new_n10658_), .ZN(new_n11259_));
  XOR2_X1    g11067(.A1(new_n10902_), .A2(new_n10658_), .Z(new_n11260_));
  NAND3_X1   g11068(.A1(new_n11259_), .A2(\asqrt[63] ), .A3(new_n11260_), .ZN(new_n11261_));
  INV_X1     g11069(.I(new_n10911_), .ZN(new_n11262_));
  NAND4_X1   g11070(.A1(new_n11262_), .A2(new_n10659_), .A3(new_n10806_), .A4(new_n10814_), .ZN(new_n11263_));
  NAND2_X1   g11071(.A1(new_n11261_), .A2(new_n11263_), .ZN(new_n11264_));
  INV_X1     g11072(.I(new_n11264_), .ZN(new_n11265_));
  NAND4_X1   g11073(.A1(new_n11255_), .A2(new_n193_), .A3(new_n11258_), .A4(new_n11265_), .ZN(\asqrt[17] ));
  AOI21_X1   g11074(.A1(new_n11089_), .A2(new_n11106_), .B(\asqrt[17] ), .ZN(new_n11267_));
  XOR2_X1    g11075(.A1(new_n11267_), .A2(new_n10817_), .Z(new_n11268_));
  AOI21_X1   g11076(.A1(new_n11086_), .A2(new_n11104_), .B(\asqrt[17] ), .ZN(new_n11269_));
  XOR2_X1    g11077(.A1(new_n11269_), .A2(new_n10820_), .Z(new_n11270_));
  NAND2_X1   g11078(.A1(new_n11099_), .A2(new_n2332_), .ZN(new_n11271_));
  AOI21_X1   g11079(.A1(new_n11271_), .A2(new_n11085_), .B(\asqrt[17] ), .ZN(new_n11272_));
  XOR2_X1    g11080(.A1(new_n11272_), .A2(new_n10823_), .Z(new_n11273_));
  INV_X1     g11081(.I(new_n11273_), .ZN(new_n11274_));
  AOI21_X1   g11082(.A1(new_n11097_), .A2(new_n11082_), .B(\asqrt[17] ), .ZN(new_n11275_));
  XOR2_X1    g11083(.A1(new_n11275_), .A2(new_n10825_), .Z(new_n11276_));
  INV_X1     g11084(.I(new_n11276_), .ZN(new_n11277_));
  NAND2_X1   g11085(.A1(new_n11064_), .A2(new_n2749_), .ZN(new_n11278_));
  AOI21_X1   g11086(.A1(new_n11278_), .A2(new_n11096_), .B(\asqrt[17] ), .ZN(new_n11279_));
  XOR2_X1    g11087(.A1(new_n11279_), .A2(new_n10828_), .Z(new_n11280_));
  AOI21_X1   g11088(.A1(new_n11062_), .A2(new_n11079_), .B(\asqrt[17] ), .ZN(new_n11281_));
  XOR2_X1    g11089(.A1(new_n11281_), .A2(new_n10832_), .Z(new_n11282_));
  NAND2_X1   g11090(.A1(new_n11075_), .A2(new_n3195_), .ZN(new_n11283_));
  AOI21_X1   g11091(.A1(new_n11283_), .A2(new_n11061_), .B(\asqrt[17] ), .ZN(new_n11284_));
  XOR2_X1    g11092(.A1(new_n11284_), .A2(new_n10835_), .Z(new_n11285_));
  INV_X1     g11093(.I(new_n11285_), .ZN(new_n11286_));
  AOI21_X1   g11094(.A1(new_n11073_), .A2(new_n11058_), .B(\asqrt[17] ), .ZN(new_n11287_));
  XOR2_X1    g11095(.A1(new_n11287_), .A2(new_n10837_), .Z(new_n11288_));
  INV_X1     g11096(.I(new_n11288_), .ZN(new_n11289_));
  NAND2_X1   g11097(.A1(new_n11040_), .A2(new_n3681_), .ZN(new_n11290_));
  AOI21_X1   g11098(.A1(new_n11290_), .A2(new_n11072_), .B(\asqrt[17] ), .ZN(new_n11291_));
  XOR2_X1    g11099(.A1(new_n11291_), .A2(new_n10840_), .Z(new_n11292_));
  AOI21_X1   g11100(.A1(new_n11038_), .A2(new_n11055_), .B(\asqrt[17] ), .ZN(new_n11293_));
  XOR2_X1    g11101(.A1(new_n11293_), .A2(new_n10844_), .Z(new_n11294_));
  NAND2_X1   g11102(.A1(new_n11051_), .A2(new_n4196_), .ZN(new_n11295_));
  AOI21_X1   g11103(.A1(new_n11295_), .A2(new_n11037_), .B(\asqrt[17] ), .ZN(new_n11296_));
  XOR2_X1    g11104(.A1(new_n11296_), .A2(new_n10847_), .Z(new_n11297_));
  INV_X1     g11105(.I(new_n11297_), .ZN(new_n11298_));
  AOI21_X1   g11106(.A1(new_n11049_), .A2(new_n11034_), .B(\asqrt[17] ), .ZN(new_n11299_));
  XOR2_X1    g11107(.A1(new_n11299_), .A2(new_n10849_), .Z(new_n11300_));
  INV_X1     g11108(.I(new_n11300_), .ZN(new_n11301_));
  NAND2_X1   g11109(.A1(new_n11016_), .A2(new_n4751_), .ZN(new_n11302_));
  AOI21_X1   g11110(.A1(new_n11302_), .A2(new_n11048_), .B(\asqrt[17] ), .ZN(new_n11303_));
  XOR2_X1    g11111(.A1(new_n11303_), .A2(new_n10852_), .Z(new_n11304_));
  AOI21_X1   g11112(.A1(new_n11014_), .A2(new_n11031_), .B(\asqrt[17] ), .ZN(new_n11305_));
  XOR2_X1    g11113(.A1(new_n11305_), .A2(new_n10856_), .Z(new_n11306_));
  NAND2_X1   g11114(.A1(new_n11027_), .A2(new_n5336_), .ZN(new_n11307_));
  AOI21_X1   g11115(.A1(new_n11307_), .A2(new_n11013_), .B(\asqrt[17] ), .ZN(new_n11308_));
  XOR2_X1    g11116(.A1(new_n11308_), .A2(new_n10859_), .Z(new_n11309_));
  INV_X1     g11117(.I(new_n11309_), .ZN(new_n11310_));
  AOI21_X1   g11118(.A1(new_n11025_), .A2(new_n11010_), .B(\asqrt[17] ), .ZN(new_n11311_));
  XOR2_X1    g11119(.A1(new_n11311_), .A2(new_n10861_), .Z(new_n11312_));
  INV_X1     g11120(.I(new_n11312_), .ZN(new_n11313_));
  NAND2_X1   g11121(.A1(new_n10992_), .A2(new_n5947_), .ZN(new_n11314_));
  AOI21_X1   g11122(.A1(new_n11314_), .A2(new_n11024_), .B(\asqrt[17] ), .ZN(new_n11315_));
  XOR2_X1    g11123(.A1(new_n11315_), .A2(new_n10864_), .Z(new_n11316_));
  AOI21_X1   g11124(.A1(new_n10990_), .A2(new_n11007_), .B(\asqrt[17] ), .ZN(new_n11317_));
  XOR2_X1    g11125(.A1(new_n11317_), .A2(new_n10868_), .Z(new_n11318_));
  NAND2_X1   g11126(.A1(new_n11003_), .A2(new_n6636_), .ZN(new_n11319_));
  AOI21_X1   g11127(.A1(new_n11319_), .A2(new_n10989_), .B(\asqrt[17] ), .ZN(new_n11320_));
  XOR2_X1    g11128(.A1(new_n11320_), .A2(new_n10871_), .Z(new_n11321_));
  INV_X1     g11129(.I(new_n11321_), .ZN(new_n11322_));
  AOI21_X1   g11130(.A1(new_n11001_), .A2(new_n10986_), .B(\asqrt[17] ), .ZN(new_n11323_));
  XOR2_X1    g11131(.A1(new_n11323_), .A2(new_n10873_), .Z(new_n11324_));
  INV_X1     g11132(.I(new_n11324_), .ZN(new_n11325_));
  NAND2_X1   g11133(.A1(new_n10968_), .A2(new_n7331_), .ZN(new_n11326_));
  AOI21_X1   g11134(.A1(new_n11326_), .A2(new_n11000_), .B(\asqrt[17] ), .ZN(new_n11327_));
  XOR2_X1    g11135(.A1(new_n11327_), .A2(new_n10876_), .Z(new_n11328_));
  AOI21_X1   g11136(.A1(new_n10966_), .A2(new_n10983_), .B(\asqrt[17] ), .ZN(new_n11329_));
  XOR2_X1    g11137(.A1(new_n11329_), .A2(new_n10880_), .Z(new_n11330_));
  NAND2_X1   g11138(.A1(new_n10979_), .A2(new_n8077_), .ZN(new_n11331_));
  AOI21_X1   g11139(.A1(new_n11331_), .A2(new_n10965_), .B(\asqrt[17] ), .ZN(new_n11332_));
  XOR2_X1    g11140(.A1(new_n11332_), .A2(new_n10883_), .Z(new_n11333_));
  INV_X1     g11141(.I(new_n11333_), .ZN(new_n11334_));
  AOI21_X1   g11142(.A1(new_n10977_), .A2(new_n10962_), .B(\asqrt[17] ), .ZN(new_n11335_));
  XOR2_X1    g11143(.A1(new_n11335_), .A2(new_n10885_), .Z(new_n11336_));
  INV_X1     g11144(.I(new_n11336_), .ZN(new_n11337_));
  NAND2_X1   g11145(.A1(new_n10940_), .A2(new_n8849_), .ZN(new_n11338_));
  AOI21_X1   g11146(.A1(new_n11338_), .A2(new_n10976_), .B(\asqrt[17] ), .ZN(new_n11339_));
  XOR2_X1    g11147(.A1(new_n11339_), .A2(new_n10888_), .Z(new_n11340_));
  AOI21_X1   g11148(.A1(new_n10938_), .A2(new_n10959_), .B(\asqrt[17] ), .ZN(new_n11341_));
  XOR2_X1    g11149(.A1(new_n11341_), .A2(new_n10891_), .Z(new_n11342_));
  NAND2_X1   g11150(.A1(new_n10955_), .A2(new_n9656_), .ZN(new_n11343_));
  AOI21_X1   g11151(.A1(new_n11343_), .A2(new_n10937_), .B(\asqrt[17] ), .ZN(new_n11344_));
  XOR2_X1    g11152(.A1(new_n11344_), .A2(new_n10898_), .Z(new_n11345_));
  INV_X1     g11153(.I(new_n11345_), .ZN(new_n11346_));
  AOI21_X1   g11154(.A1(new_n10953_), .A2(new_n10934_), .B(\asqrt[17] ), .ZN(new_n11347_));
  XOR2_X1    g11155(.A1(new_n11347_), .A2(new_n10944_), .Z(new_n11348_));
  INV_X1     g11156(.I(new_n11348_), .ZN(new_n11349_));
  NAND2_X1   g11157(.A1(\asqrt[18] ), .A2(new_n10921_), .ZN(new_n11350_));
  NOR2_X1    g11158(.A1(new_n10929_), .A2(\a[36] ), .ZN(new_n11351_));
  AOI22_X1   g11159(.A1(new_n11350_), .A2(new_n10929_), .B1(\asqrt[18] ), .B2(new_n11351_), .ZN(new_n11352_));
  OAI21_X1   g11160(.A1(new_n10914_), .A2(new_n10921_), .B(new_n10948_), .ZN(new_n11353_));
  AOI21_X1   g11161(.A1(new_n10947_), .A2(new_n11353_), .B(\asqrt[17] ), .ZN(new_n11354_));
  XOR2_X1    g11162(.A1(new_n11354_), .A2(new_n11352_), .Z(new_n11355_));
  NAND3_X1   g11163(.A1(new_n11240_), .A2(new_n239_), .A3(new_n11233_), .ZN(new_n11356_));
  AOI21_X1   g11164(.A1(new_n11236_), .A2(new_n11356_), .B(new_n11241_), .ZN(new_n11357_));
  AOI21_X1   g11165(.A1(new_n11237_), .A2(new_n11232_), .B(\asqrt[62] ), .ZN(new_n11358_));
  NOR3_X1    g11166(.A1(new_n11244_), .A2(new_n201_), .A3(new_n11241_), .ZN(new_n11359_));
  OAI22_X1   g11167(.A1(new_n11359_), .A2(new_n11358_), .B1(new_n11357_), .B2(new_n11249_), .ZN(new_n11360_));
  AOI21_X1   g11168(.A1(new_n11360_), .A2(new_n11110_), .B(new_n11253_), .ZN(new_n11361_));
  AOI21_X1   g11169(.A1(new_n11357_), .A2(new_n201_), .B(new_n11250_), .ZN(new_n11362_));
  OAI21_X1   g11170(.A1(new_n11357_), .A2(new_n201_), .B(new_n11111_), .ZN(new_n11363_));
  NOR2_X1    g11171(.A1(new_n11362_), .A2(new_n11363_), .ZN(new_n11364_));
  NOR3_X1    g11172(.A1(new_n11361_), .A2(\asqrt[63] ), .A3(new_n11364_), .ZN(new_n11365_));
  NAND3_X1   g11173(.A1(new_n11261_), .A2(\asqrt[18] ), .A3(new_n11263_), .ZN(new_n11366_));
  INV_X1     g11174(.I(new_n11366_), .ZN(new_n11367_));
  NAND2_X1   g11175(.A1(new_n11365_), .A2(new_n11367_), .ZN(new_n11368_));
  NAND2_X1   g11176(.A1(\asqrt[17] ), .A2(new_n10918_), .ZN(new_n11369_));
  AOI21_X1   g11177(.A1(new_n11369_), .A2(new_n11368_), .B(\a[36] ), .ZN(new_n11370_));
  NAND2_X1   g11178(.A1(new_n11255_), .A2(new_n193_), .ZN(new_n11371_));
  NOR3_X1    g11179(.A1(new_n11371_), .A2(new_n11364_), .A3(new_n11366_), .ZN(new_n11372_));
  NOR4_X1    g11180(.A1(new_n11361_), .A2(\asqrt[63] ), .A3(new_n11364_), .A4(new_n11264_), .ZN(new_n11373_));
  NOR2_X1    g11181(.A1(new_n11373_), .A2(new_n10919_), .ZN(new_n11374_));
  NOR3_X1    g11182(.A1(new_n11374_), .A2(new_n11372_), .A3(new_n10921_), .ZN(new_n11375_));
  NOR2_X1    g11183(.A1(new_n11375_), .A2(new_n11370_), .ZN(new_n11376_));
  INV_X1     g11184(.I(\a[34] ), .ZN(new_n11377_));
  NOR2_X1    g11185(.A1(\a[32] ), .A2(\a[33] ), .ZN(new_n11378_));
  NOR3_X1    g11186(.A1(new_n11373_), .A2(new_n11377_), .A3(new_n11378_), .ZN(new_n11379_));
  INV_X1     g11187(.I(new_n11378_), .ZN(new_n11380_));
  AOI21_X1   g11188(.A1(new_n11373_), .A2(\a[34] ), .B(new_n11380_), .ZN(new_n11381_));
  OAI21_X1   g11189(.A1(new_n11379_), .A2(new_n11381_), .B(\asqrt[18] ), .ZN(new_n11382_));
  NAND2_X1   g11190(.A1(new_n11378_), .A2(new_n11377_), .ZN(new_n11383_));
  NAND3_X1   g11191(.A1(new_n10810_), .A2(new_n10812_), .A3(new_n11383_), .ZN(new_n11384_));
  NAND2_X1   g11192(.A1(new_n10907_), .A2(new_n11384_), .ZN(new_n11385_));
  INV_X1     g11193(.I(new_n11385_), .ZN(new_n11386_));
  NOR3_X1    g11194(.A1(new_n11373_), .A2(new_n11377_), .A3(new_n11386_), .ZN(new_n11387_));
  NOR3_X1    g11195(.A1(new_n11373_), .A2(\a[34] ), .A3(\a[35] ), .ZN(new_n11388_));
  INV_X1     g11196(.I(\a[35] ), .ZN(new_n11389_));
  AOI21_X1   g11197(.A1(\asqrt[17] ), .A2(new_n11377_), .B(new_n11389_), .ZN(new_n11390_));
  NOR3_X1    g11198(.A1(new_n11387_), .A2(new_n11388_), .A3(new_n11390_), .ZN(new_n11391_));
  NAND3_X1   g11199(.A1(new_n11391_), .A2(new_n11382_), .A3(new_n10497_), .ZN(new_n11392_));
  NAND2_X1   g11200(.A1(new_n11392_), .A2(new_n11376_), .ZN(new_n11393_));
  NAND3_X1   g11201(.A1(\asqrt[17] ), .A2(\a[34] ), .A3(new_n11380_), .ZN(new_n11394_));
  OAI21_X1   g11202(.A1(\asqrt[17] ), .A2(new_n11377_), .B(new_n11378_), .ZN(new_n11395_));
  AOI21_X1   g11203(.A1(new_n11395_), .A2(new_n11394_), .B(new_n10914_), .ZN(new_n11396_));
  NAND3_X1   g11204(.A1(\asqrt[17] ), .A2(\a[34] ), .A3(new_n11385_), .ZN(new_n11397_));
  NAND3_X1   g11205(.A1(\asqrt[17] ), .A2(new_n11377_), .A3(new_n11389_), .ZN(new_n11398_));
  OAI21_X1   g11206(.A1(new_n11373_), .A2(\a[34] ), .B(\a[35] ), .ZN(new_n11399_));
  NAND3_X1   g11207(.A1(new_n11397_), .A2(new_n11399_), .A3(new_n11398_), .ZN(new_n11400_));
  OAI21_X1   g11208(.A1(new_n11400_), .A2(new_n11396_), .B(\asqrt[19] ), .ZN(new_n11401_));
  NAND3_X1   g11209(.A1(new_n11393_), .A2(new_n10052_), .A3(new_n11401_), .ZN(new_n11402_));
  AOI21_X1   g11210(.A1(new_n11393_), .A2(new_n11401_), .B(new_n10052_), .ZN(new_n11403_));
  AOI21_X1   g11211(.A1(new_n11355_), .A2(new_n11402_), .B(new_n11403_), .ZN(new_n11404_));
  AOI21_X1   g11212(.A1(new_n11404_), .A2(new_n9656_), .B(new_n11349_), .ZN(new_n11405_));
  OR2_X2     g11213(.A1(new_n11375_), .A2(new_n11370_), .Z(new_n11406_));
  NOR3_X1    g11214(.A1(new_n11400_), .A2(new_n11396_), .A3(\asqrt[19] ), .ZN(new_n11407_));
  OAI21_X1   g11215(.A1(new_n11406_), .A2(new_n11407_), .B(new_n11401_), .ZN(new_n11408_));
  OAI21_X1   g11216(.A1(new_n11408_), .A2(\asqrt[20] ), .B(new_n11355_), .ZN(new_n11409_));
  NAND2_X1   g11217(.A1(new_n11408_), .A2(\asqrt[20] ), .ZN(new_n11410_));
  AOI21_X1   g11218(.A1(new_n11409_), .A2(new_n11410_), .B(new_n9656_), .ZN(new_n11411_));
  NOR3_X1    g11219(.A1(new_n11405_), .A2(\asqrt[22] ), .A3(new_n11411_), .ZN(new_n11412_));
  OAI21_X1   g11220(.A1(new_n11405_), .A2(new_n11411_), .B(\asqrt[22] ), .ZN(new_n11413_));
  OAI21_X1   g11221(.A1(new_n11346_), .A2(new_n11412_), .B(new_n11413_), .ZN(new_n11414_));
  OAI21_X1   g11222(.A1(new_n11414_), .A2(\asqrt[23] ), .B(new_n11342_), .ZN(new_n11415_));
  NAND3_X1   g11223(.A1(new_n11409_), .A2(new_n11410_), .A3(new_n9656_), .ZN(new_n11416_));
  AOI21_X1   g11224(.A1(new_n11348_), .A2(new_n11416_), .B(new_n11411_), .ZN(new_n11417_));
  AOI21_X1   g11225(.A1(new_n11417_), .A2(new_n9233_), .B(new_n11346_), .ZN(new_n11418_));
  NAND2_X1   g11226(.A1(new_n11416_), .A2(new_n11348_), .ZN(new_n11419_));
  INV_X1     g11227(.I(new_n11411_), .ZN(new_n11420_));
  AOI21_X1   g11228(.A1(new_n11419_), .A2(new_n11420_), .B(new_n9233_), .ZN(new_n11421_));
  OAI21_X1   g11229(.A1(new_n11418_), .A2(new_n11421_), .B(\asqrt[23] ), .ZN(new_n11422_));
  NAND3_X1   g11230(.A1(new_n11415_), .A2(new_n8440_), .A3(new_n11422_), .ZN(new_n11423_));
  AOI21_X1   g11231(.A1(new_n11415_), .A2(new_n11422_), .B(new_n8440_), .ZN(new_n11424_));
  AOI21_X1   g11232(.A1(new_n11340_), .A2(new_n11423_), .B(new_n11424_), .ZN(new_n11425_));
  AOI21_X1   g11233(.A1(new_n11425_), .A2(new_n8077_), .B(new_n11337_), .ZN(new_n11426_));
  INV_X1     g11234(.I(new_n11342_), .ZN(new_n11427_));
  NOR3_X1    g11235(.A1(new_n11418_), .A2(\asqrt[23] ), .A3(new_n11421_), .ZN(new_n11428_));
  OAI21_X1   g11236(.A1(new_n11427_), .A2(new_n11428_), .B(new_n11422_), .ZN(new_n11429_));
  OAI21_X1   g11237(.A1(new_n11429_), .A2(\asqrt[24] ), .B(new_n11340_), .ZN(new_n11430_));
  NAND2_X1   g11238(.A1(new_n11429_), .A2(\asqrt[24] ), .ZN(new_n11431_));
  AOI21_X1   g11239(.A1(new_n11430_), .A2(new_n11431_), .B(new_n8077_), .ZN(new_n11432_));
  NOR3_X1    g11240(.A1(new_n11426_), .A2(\asqrt[26] ), .A3(new_n11432_), .ZN(new_n11433_));
  OAI21_X1   g11241(.A1(new_n11426_), .A2(new_n11432_), .B(\asqrt[26] ), .ZN(new_n11434_));
  OAI21_X1   g11242(.A1(new_n11334_), .A2(new_n11433_), .B(new_n11434_), .ZN(new_n11435_));
  OAI21_X1   g11243(.A1(new_n11435_), .A2(\asqrt[27] ), .B(new_n11330_), .ZN(new_n11436_));
  NAND3_X1   g11244(.A1(new_n11430_), .A2(new_n11431_), .A3(new_n8077_), .ZN(new_n11437_));
  AOI21_X1   g11245(.A1(new_n11336_), .A2(new_n11437_), .B(new_n11432_), .ZN(new_n11438_));
  AOI21_X1   g11246(.A1(new_n11438_), .A2(new_n7690_), .B(new_n11334_), .ZN(new_n11439_));
  NAND2_X1   g11247(.A1(new_n11437_), .A2(new_n11336_), .ZN(new_n11440_));
  INV_X1     g11248(.I(new_n11432_), .ZN(new_n11441_));
  AOI21_X1   g11249(.A1(new_n11440_), .A2(new_n11441_), .B(new_n7690_), .ZN(new_n11442_));
  OAI21_X1   g11250(.A1(new_n11439_), .A2(new_n11442_), .B(\asqrt[27] ), .ZN(new_n11443_));
  NAND3_X1   g11251(.A1(new_n11436_), .A2(new_n6966_), .A3(new_n11443_), .ZN(new_n11444_));
  AOI21_X1   g11252(.A1(new_n11436_), .A2(new_n11443_), .B(new_n6966_), .ZN(new_n11445_));
  AOI21_X1   g11253(.A1(new_n11328_), .A2(new_n11444_), .B(new_n11445_), .ZN(new_n11446_));
  AOI21_X1   g11254(.A1(new_n11446_), .A2(new_n6636_), .B(new_n11325_), .ZN(new_n11447_));
  INV_X1     g11255(.I(new_n11330_), .ZN(new_n11448_));
  NOR3_X1    g11256(.A1(new_n11439_), .A2(\asqrt[27] ), .A3(new_n11442_), .ZN(new_n11449_));
  OAI21_X1   g11257(.A1(new_n11448_), .A2(new_n11449_), .B(new_n11443_), .ZN(new_n11450_));
  OAI21_X1   g11258(.A1(new_n11450_), .A2(\asqrt[28] ), .B(new_n11328_), .ZN(new_n11451_));
  NAND2_X1   g11259(.A1(new_n11450_), .A2(\asqrt[28] ), .ZN(new_n11452_));
  AOI21_X1   g11260(.A1(new_n11451_), .A2(new_n11452_), .B(new_n6636_), .ZN(new_n11453_));
  NOR3_X1    g11261(.A1(new_n11447_), .A2(\asqrt[30] ), .A3(new_n11453_), .ZN(new_n11454_));
  OAI21_X1   g11262(.A1(new_n11447_), .A2(new_n11453_), .B(\asqrt[30] ), .ZN(new_n11455_));
  OAI21_X1   g11263(.A1(new_n11322_), .A2(new_n11454_), .B(new_n11455_), .ZN(new_n11456_));
  OAI21_X1   g11264(.A1(new_n11456_), .A2(\asqrt[31] ), .B(new_n11318_), .ZN(new_n11457_));
  NAND3_X1   g11265(.A1(new_n11451_), .A2(new_n11452_), .A3(new_n6636_), .ZN(new_n11458_));
  AOI21_X1   g11266(.A1(new_n11324_), .A2(new_n11458_), .B(new_n11453_), .ZN(new_n11459_));
  AOI21_X1   g11267(.A1(new_n11459_), .A2(new_n6275_), .B(new_n11322_), .ZN(new_n11460_));
  NAND2_X1   g11268(.A1(new_n11458_), .A2(new_n11324_), .ZN(new_n11461_));
  INV_X1     g11269(.I(new_n11453_), .ZN(new_n11462_));
  AOI21_X1   g11270(.A1(new_n11461_), .A2(new_n11462_), .B(new_n6275_), .ZN(new_n11463_));
  OAI21_X1   g11271(.A1(new_n11460_), .A2(new_n11463_), .B(\asqrt[31] ), .ZN(new_n11464_));
  NAND3_X1   g11272(.A1(new_n11457_), .A2(new_n5643_), .A3(new_n11464_), .ZN(new_n11465_));
  AOI21_X1   g11273(.A1(new_n11457_), .A2(new_n11464_), .B(new_n5643_), .ZN(new_n11466_));
  AOI21_X1   g11274(.A1(new_n11316_), .A2(new_n11465_), .B(new_n11466_), .ZN(new_n11467_));
  AOI21_X1   g11275(.A1(new_n11467_), .A2(new_n5336_), .B(new_n11313_), .ZN(new_n11468_));
  INV_X1     g11276(.I(new_n11318_), .ZN(new_n11469_));
  NOR3_X1    g11277(.A1(new_n11460_), .A2(\asqrt[31] ), .A3(new_n11463_), .ZN(new_n11470_));
  OAI21_X1   g11278(.A1(new_n11469_), .A2(new_n11470_), .B(new_n11464_), .ZN(new_n11471_));
  OAI21_X1   g11279(.A1(new_n11471_), .A2(\asqrt[32] ), .B(new_n11316_), .ZN(new_n11472_));
  NAND2_X1   g11280(.A1(new_n11471_), .A2(\asqrt[32] ), .ZN(new_n11473_));
  AOI21_X1   g11281(.A1(new_n11472_), .A2(new_n11473_), .B(new_n5336_), .ZN(new_n11474_));
  NOR3_X1    g11282(.A1(new_n11468_), .A2(\asqrt[34] ), .A3(new_n11474_), .ZN(new_n11475_));
  OAI21_X1   g11283(.A1(new_n11468_), .A2(new_n11474_), .B(\asqrt[34] ), .ZN(new_n11476_));
  OAI21_X1   g11284(.A1(new_n11310_), .A2(new_n11475_), .B(new_n11476_), .ZN(new_n11477_));
  OAI21_X1   g11285(.A1(new_n11477_), .A2(\asqrt[35] ), .B(new_n11306_), .ZN(new_n11478_));
  NAND3_X1   g11286(.A1(new_n11472_), .A2(new_n11473_), .A3(new_n5336_), .ZN(new_n11479_));
  AOI21_X1   g11287(.A1(new_n11312_), .A2(new_n11479_), .B(new_n11474_), .ZN(new_n11480_));
  AOI21_X1   g11288(.A1(new_n11480_), .A2(new_n5029_), .B(new_n11310_), .ZN(new_n11481_));
  NAND2_X1   g11289(.A1(new_n11479_), .A2(new_n11312_), .ZN(new_n11482_));
  INV_X1     g11290(.I(new_n11474_), .ZN(new_n11483_));
  AOI21_X1   g11291(.A1(new_n11482_), .A2(new_n11483_), .B(new_n5029_), .ZN(new_n11484_));
  OAI21_X1   g11292(.A1(new_n11481_), .A2(new_n11484_), .B(\asqrt[35] ), .ZN(new_n11485_));
  NAND3_X1   g11293(.A1(new_n11478_), .A2(new_n4461_), .A3(new_n11485_), .ZN(new_n11486_));
  AOI21_X1   g11294(.A1(new_n11478_), .A2(new_n11485_), .B(new_n4461_), .ZN(new_n11487_));
  AOI21_X1   g11295(.A1(new_n11304_), .A2(new_n11486_), .B(new_n11487_), .ZN(new_n11488_));
  AOI21_X1   g11296(.A1(new_n11488_), .A2(new_n4196_), .B(new_n11301_), .ZN(new_n11489_));
  INV_X1     g11297(.I(new_n11306_), .ZN(new_n11490_));
  NOR3_X1    g11298(.A1(new_n11481_), .A2(\asqrt[35] ), .A3(new_n11484_), .ZN(new_n11491_));
  OAI21_X1   g11299(.A1(new_n11490_), .A2(new_n11491_), .B(new_n11485_), .ZN(new_n11492_));
  OAI21_X1   g11300(.A1(new_n11492_), .A2(\asqrt[36] ), .B(new_n11304_), .ZN(new_n11493_));
  NAND2_X1   g11301(.A1(new_n11492_), .A2(\asqrt[36] ), .ZN(new_n11494_));
  AOI21_X1   g11302(.A1(new_n11493_), .A2(new_n11494_), .B(new_n4196_), .ZN(new_n11495_));
  NOR3_X1    g11303(.A1(new_n11489_), .A2(\asqrt[38] ), .A3(new_n11495_), .ZN(new_n11496_));
  OAI21_X1   g11304(.A1(new_n11489_), .A2(new_n11495_), .B(\asqrt[38] ), .ZN(new_n11497_));
  OAI21_X1   g11305(.A1(new_n11298_), .A2(new_n11496_), .B(new_n11497_), .ZN(new_n11498_));
  OAI21_X1   g11306(.A1(new_n11498_), .A2(\asqrt[39] ), .B(new_n11294_), .ZN(new_n11499_));
  NAND3_X1   g11307(.A1(new_n11493_), .A2(new_n11494_), .A3(new_n4196_), .ZN(new_n11500_));
  AOI21_X1   g11308(.A1(new_n11300_), .A2(new_n11500_), .B(new_n11495_), .ZN(new_n11501_));
  AOI21_X1   g11309(.A1(new_n11501_), .A2(new_n3925_), .B(new_n11298_), .ZN(new_n11502_));
  NAND2_X1   g11310(.A1(new_n11500_), .A2(new_n11300_), .ZN(new_n11503_));
  INV_X1     g11311(.I(new_n11495_), .ZN(new_n11504_));
  AOI21_X1   g11312(.A1(new_n11503_), .A2(new_n11504_), .B(new_n3925_), .ZN(new_n11505_));
  OAI21_X1   g11313(.A1(new_n11502_), .A2(new_n11505_), .B(\asqrt[39] ), .ZN(new_n11506_));
  NAND3_X1   g11314(.A1(new_n11499_), .A2(new_n3427_), .A3(new_n11506_), .ZN(new_n11507_));
  AOI21_X1   g11315(.A1(new_n11499_), .A2(new_n11506_), .B(new_n3427_), .ZN(new_n11508_));
  AOI21_X1   g11316(.A1(new_n11292_), .A2(new_n11507_), .B(new_n11508_), .ZN(new_n11509_));
  AOI21_X1   g11317(.A1(new_n11509_), .A2(new_n3195_), .B(new_n11289_), .ZN(new_n11510_));
  INV_X1     g11318(.I(new_n11294_), .ZN(new_n11511_));
  NOR3_X1    g11319(.A1(new_n11502_), .A2(\asqrt[39] ), .A3(new_n11505_), .ZN(new_n11512_));
  OAI21_X1   g11320(.A1(new_n11511_), .A2(new_n11512_), .B(new_n11506_), .ZN(new_n11513_));
  OAI21_X1   g11321(.A1(new_n11513_), .A2(\asqrt[40] ), .B(new_n11292_), .ZN(new_n11514_));
  NAND2_X1   g11322(.A1(new_n11513_), .A2(\asqrt[40] ), .ZN(new_n11515_));
  AOI21_X1   g11323(.A1(new_n11514_), .A2(new_n11515_), .B(new_n3195_), .ZN(new_n11516_));
  NOR3_X1    g11324(.A1(new_n11510_), .A2(\asqrt[42] ), .A3(new_n11516_), .ZN(new_n11517_));
  OAI21_X1   g11325(.A1(new_n11510_), .A2(new_n11516_), .B(\asqrt[42] ), .ZN(new_n11518_));
  OAI21_X1   g11326(.A1(new_n11286_), .A2(new_n11517_), .B(new_n11518_), .ZN(new_n11519_));
  OAI21_X1   g11327(.A1(new_n11519_), .A2(\asqrt[43] ), .B(new_n11282_), .ZN(new_n11520_));
  NAND3_X1   g11328(.A1(new_n11514_), .A2(new_n11515_), .A3(new_n3195_), .ZN(new_n11521_));
  AOI21_X1   g11329(.A1(new_n11288_), .A2(new_n11521_), .B(new_n11516_), .ZN(new_n11522_));
  AOI21_X1   g11330(.A1(new_n11522_), .A2(new_n2960_), .B(new_n11286_), .ZN(new_n11523_));
  NAND2_X1   g11331(.A1(new_n11521_), .A2(new_n11288_), .ZN(new_n11524_));
  INV_X1     g11332(.I(new_n11516_), .ZN(new_n11525_));
  AOI21_X1   g11333(.A1(new_n11524_), .A2(new_n11525_), .B(new_n2960_), .ZN(new_n11526_));
  OAI21_X1   g11334(.A1(new_n11523_), .A2(new_n11526_), .B(\asqrt[43] ), .ZN(new_n11527_));
  NAND3_X1   g11335(.A1(new_n11520_), .A2(new_n2531_), .A3(new_n11527_), .ZN(new_n11528_));
  AOI21_X1   g11336(.A1(new_n11520_), .A2(new_n11527_), .B(new_n2531_), .ZN(new_n11529_));
  AOI21_X1   g11337(.A1(new_n11280_), .A2(new_n11528_), .B(new_n11529_), .ZN(new_n11530_));
  AOI21_X1   g11338(.A1(new_n11530_), .A2(new_n2332_), .B(new_n11277_), .ZN(new_n11531_));
  INV_X1     g11339(.I(new_n11282_), .ZN(new_n11532_));
  NOR3_X1    g11340(.A1(new_n11523_), .A2(\asqrt[43] ), .A3(new_n11526_), .ZN(new_n11533_));
  OAI21_X1   g11341(.A1(new_n11532_), .A2(new_n11533_), .B(new_n11527_), .ZN(new_n11534_));
  OAI21_X1   g11342(.A1(new_n11534_), .A2(\asqrt[44] ), .B(new_n11280_), .ZN(new_n11535_));
  NAND2_X1   g11343(.A1(new_n11534_), .A2(\asqrt[44] ), .ZN(new_n11536_));
  AOI21_X1   g11344(.A1(new_n11535_), .A2(new_n11536_), .B(new_n2332_), .ZN(new_n11537_));
  NOR3_X1    g11345(.A1(new_n11531_), .A2(\asqrt[46] ), .A3(new_n11537_), .ZN(new_n11538_));
  OAI21_X1   g11346(.A1(new_n11531_), .A2(new_n11537_), .B(\asqrt[46] ), .ZN(new_n11539_));
  OAI21_X1   g11347(.A1(new_n11274_), .A2(new_n11538_), .B(new_n11539_), .ZN(new_n11540_));
  OAI21_X1   g11348(.A1(new_n11540_), .A2(\asqrt[47] ), .B(new_n11270_), .ZN(new_n11541_));
  NAND3_X1   g11349(.A1(new_n11535_), .A2(new_n11536_), .A3(new_n2332_), .ZN(new_n11542_));
  AOI21_X1   g11350(.A1(new_n11276_), .A2(new_n11542_), .B(new_n11537_), .ZN(new_n11543_));
  AOI21_X1   g11351(.A1(new_n11543_), .A2(new_n2134_), .B(new_n11274_), .ZN(new_n11544_));
  NAND2_X1   g11352(.A1(new_n11542_), .A2(new_n11276_), .ZN(new_n11545_));
  INV_X1     g11353(.I(new_n11537_), .ZN(new_n11546_));
  AOI21_X1   g11354(.A1(new_n11545_), .A2(new_n11546_), .B(new_n2134_), .ZN(new_n11547_));
  OAI21_X1   g11355(.A1(new_n11544_), .A2(new_n11547_), .B(\asqrt[47] ), .ZN(new_n11548_));
  NAND3_X1   g11356(.A1(new_n11541_), .A2(new_n1778_), .A3(new_n11548_), .ZN(new_n11549_));
  INV_X1     g11357(.I(new_n11270_), .ZN(new_n11550_));
  NOR3_X1    g11358(.A1(new_n11544_), .A2(\asqrt[47] ), .A3(new_n11547_), .ZN(new_n11551_));
  OAI21_X1   g11359(.A1(new_n11550_), .A2(new_n11551_), .B(new_n11548_), .ZN(new_n11552_));
  NAND2_X1   g11360(.A1(new_n11552_), .A2(\asqrt[48] ), .ZN(new_n11553_));
  NOR2_X1    g11361(.A1(new_n11238_), .A2(\asqrt[62] ), .ZN(new_n11554_));
  INV_X1     g11362(.I(new_n11257_), .ZN(new_n11555_));
  NOR2_X1    g11363(.A1(new_n11555_), .A2(new_n11554_), .ZN(new_n11556_));
  XOR2_X1    g11364(.A1(new_n11248_), .A2(new_n10770_), .Z(new_n11557_));
  OAI21_X1   g11365(.A1(\asqrt[17] ), .A2(new_n11556_), .B(new_n11557_), .ZN(new_n11558_));
  INV_X1     g11366(.I(new_n11558_), .ZN(new_n11559_));
  NAND2_X1   g11367(.A1(new_n11206_), .A2(new_n337_), .ZN(new_n11560_));
  AOI21_X1   g11368(.A1(new_n11560_), .A2(new_n11230_), .B(\asqrt[17] ), .ZN(new_n11561_));
  XOR2_X1    g11369(.A1(new_n11561_), .A2(new_n11116_), .Z(new_n11562_));
  INV_X1     g11370(.I(new_n11562_), .ZN(new_n11563_));
  AOI21_X1   g11371(.A1(new_n11204_), .A2(new_n11221_), .B(\asqrt[17] ), .ZN(new_n11564_));
  XOR2_X1    g11372(.A1(new_n11564_), .A2(new_n11120_), .Z(new_n11565_));
  INV_X1     g11373(.I(new_n11565_), .ZN(new_n11566_));
  NAND2_X1   g11374(.A1(new_n11217_), .A2(new_n531_), .ZN(new_n11567_));
  AOI21_X1   g11375(.A1(new_n11567_), .A2(new_n11203_), .B(\asqrt[17] ), .ZN(new_n11568_));
  XOR2_X1    g11376(.A1(new_n11568_), .A2(new_n11123_), .Z(new_n11569_));
  INV_X1     g11377(.I(new_n11569_), .ZN(new_n11570_));
  AOI21_X1   g11378(.A1(new_n11215_), .A2(new_n11200_), .B(\asqrt[17] ), .ZN(new_n11571_));
  XOR2_X1    g11379(.A1(new_n11571_), .A2(new_n11125_), .Z(new_n11572_));
  NAND2_X1   g11380(.A1(new_n11182_), .A2(new_n744_), .ZN(new_n11573_));
  AOI21_X1   g11381(.A1(new_n11573_), .A2(new_n11214_), .B(\asqrt[17] ), .ZN(new_n11574_));
  XOR2_X1    g11382(.A1(new_n11574_), .A2(new_n11128_), .Z(new_n11575_));
  AOI21_X1   g11383(.A1(new_n11180_), .A2(new_n11197_), .B(\asqrt[17] ), .ZN(new_n11576_));
  XOR2_X1    g11384(.A1(new_n11576_), .A2(new_n11132_), .Z(new_n11577_));
  INV_X1     g11385(.I(new_n11577_), .ZN(new_n11578_));
  NAND2_X1   g11386(.A1(new_n11193_), .A2(new_n1006_), .ZN(new_n11579_));
  AOI21_X1   g11387(.A1(new_n11579_), .A2(new_n11179_), .B(\asqrt[17] ), .ZN(new_n11580_));
  XOR2_X1    g11388(.A1(new_n11580_), .A2(new_n11135_), .Z(new_n11581_));
  INV_X1     g11389(.I(new_n11581_), .ZN(new_n11582_));
  AOI21_X1   g11390(.A1(new_n11191_), .A2(new_n11176_), .B(\asqrt[17] ), .ZN(new_n11583_));
  XOR2_X1    g11391(.A1(new_n11583_), .A2(new_n11137_), .Z(new_n11584_));
  NAND2_X1   g11392(.A1(new_n11162_), .A2(new_n1305_), .ZN(new_n11585_));
  AOI21_X1   g11393(.A1(new_n11585_), .A2(new_n11190_), .B(\asqrt[17] ), .ZN(new_n11586_));
  XOR2_X1    g11394(.A1(new_n11586_), .A2(new_n11140_), .Z(new_n11587_));
  AOI21_X1   g11395(.A1(new_n11160_), .A2(new_n11173_), .B(\asqrt[17] ), .ZN(new_n11588_));
  XOR2_X1    g11396(.A1(new_n11588_), .A2(new_n11144_), .Z(new_n11589_));
  INV_X1     g11397(.I(new_n11589_), .ZN(new_n11590_));
  NAND2_X1   g11398(.A1(new_n11169_), .A2(new_n1632_), .ZN(new_n11591_));
  AOI21_X1   g11399(.A1(new_n11591_), .A2(new_n11159_), .B(\asqrt[17] ), .ZN(new_n11592_));
  XOR2_X1    g11400(.A1(new_n11592_), .A2(new_n11147_), .Z(new_n11593_));
  INV_X1     g11401(.I(new_n11593_), .ZN(new_n11594_));
  AOI21_X1   g11402(.A1(new_n11167_), .A2(new_n11156_), .B(\asqrt[17] ), .ZN(new_n11595_));
  XOR2_X1    g11403(.A1(new_n11595_), .A2(new_n11149_), .Z(new_n11596_));
  OAI21_X1   g11404(.A1(new_n11552_), .A2(\asqrt[48] ), .B(new_n11268_), .ZN(new_n11597_));
  NAND3_X1   g11405(.A1(new_n11597_), .A2(new_n11553_), .A3(new_n1632_), .ZN(new_n11598_));
  AOI21_X1   g11406(.A1(new_n11597_), .A2(new_n11553_), .B(new_n1632_), .ZN(new_n11599_));
  AOI21_X1   g11407(.A1(new_n11596_), .A2(new_n11598_), .B(new_n11599_), .ZN(new_n11600_));
  AOI21_X1   g11408(.A1(new_n11600_), .A2(new_n1463_), .B(new_n11594_), .ZN(new_n11601_));
  NAND2_X1   g11409(.A1(new_n11598_), .A2(new_n11596_), .ZN(new_n11602_));
  INV_X1     g11410(.I(new_n11599_), .ZN(new_n11603_));
  AOI21_X1   g11411(.A1(new_n11602_), .A2(new_n11603_), .B(new_n1463_), .ZN(new_n11604_));
  NOR3_X1    g11412(.A1(new_n11601_), .A2(\asqrt[51] ), .A3(new_n11604_), .ZN(new_n11605_));
  OAI21_X1   g11413(.A1(new_n11601_), .A2(new_n11604_), .B(\asqrt[51] ), .ZN(new_n11606_));
  OAI21_X1   g11414(.A1(new_n11590_), .A2(new_n11605_), .B(new_n11606_), .ZN(new_n11607_));
  OAI21_X1   g11415(.A1(new_n11607_), .A2(\asqrt[52] ), .B(new_n11587_), .ZN(new_n11608_));
  NAND2_X1   g11416(.A1(new_n11607_), .A2(\asqrt[52] ), .ZN(new_n11609_));
  NAND3_X1   g11417(.A1(new_n11608_), .A2(new_n11609_), .A3(new_n1006_), .ZN(new_n11610_));
  AOI21_X1   g11418(.A1(new_n11608_), .A2(new_n11609_), .B(new_n1006_), .ZN(new_n11611_));
  AOI21_X1   g11419(.A1(new_n11584_), .A2(new_n11610_), .B(new_n11611_), .ZN(new_n11612_));
  AOI21_X1   g11420(.A1(new_n11612_), .A2(new_n860_), .B(new_n11582_), .ZN(new_n11613_));
  NAND2_X1   g11421(.A1(new_n11610_), .A2(new_n11584_), .ZN(new_n11614_));
  INV_X1     g11422(.I(new_n11611_), .ZN(new_n11615_));
  AOI21_X1   g11423(.A1(new_n11614_), .A2(new_n11615_), .B(new_n860_), .ZN(new_n11616_));
  NOR3_X1    g11424(.A1(new_n11613_), .A2(\asqrt[55] ), .A3(new_n11616_), .ZN(new_n11617_));
  OAI21_X1   g11425(.A1(new_n11613_), .A2(new_n11616_), .B(\asqrt[55] ), .ZN(new_n11618_));
  OAI21_X1   g11426(.A1(new_n11578_), .A2(new_n11617_), .B(new_n11618_), .ZN(new_n11619_));
  OAI21_X1   g11427(.A1(new_n11619_), .A2(\asqrt[56] ), .B(new_n11575_), .ZN(new_n11620_));
  NAND2_X1   g11428(.A1(new_n11619_), .A2(\asqrt[56] ), .ZN(new_n11621_));
  NAND3_X1   g11429(.A1(new_n11620_), .A2(new_n11621_), .A3(new_n531_), .ZN(new_n11622_));
  AOI21_X1   g11430(.A1(new_n11620_), .A2(new_n11621_), .B(new_n531_), .ZN(new_n11623_));
  AOI21_X1   g11431(.A1(new_n11572_), .A2(new_n11622_), .B(new_n11623_), .ZN(new_n11624_));
  AOI21_X1   g11432(.A1(new_n11624_), .A2(new_n423_), .B(new_n11570_), .ZN(new_n11625_));
  NAND2_X1   g11433(.A1(new_n11622_), .A2(new_n11572_), .ZN(new_n11626_));
  INV_X1     g11434(.I(new_n11623_), .ZN(new_n11627_));
  AOI21_X1   g11435(.A1(new_n11626_), .A2(new_n11627_), .B(new_n423_), .ZN(new_n11628_));
  NOR3_X1    g11436(.A1(new_n11625_), .A2(\asqrt[59] ), .A3(new_n11628_), .ZN(new_n11629_));
  NOR2_X1    g11437(.A1(new_n11629_), .A2(new_n11566_), .ZN(new_n11630_));
  OAI21_X1   g11438(.A1(new_n11625_), .A2(new_n11628_), .B(\asqrt[59] ), .ZN(new_n11631_));
  INV_X1     g11439(.I(new_n11631_), .ZN(new_n11632_));
  NOR2_X1    g11440(.A1(new_n11630_), .A2(new_n11632_), .ZN(new_n11633_));
  AOI21_X1   g11441(.A1(new_n11633_), .A2(new_n266_), .B(new_n11563_), .ZN(new_n11634_));
  INV_X1     g11442(.I(new_n11572_), .ZN(new_n11635_));
  INV_X1     g11443(.I(new_n11584_), .ZN(new_n11636_));
  INV_X1     g11444(.I(new_n11596_), .ZN(new_n11637_));
  AOI21_X1   g11445(.A1(new_n11541_), .A2(new_n11548_), .B(new_n1778_), .ZN(new_n11638_));
  AOI21_X1   g11446(.A1(new_n11268_), .A2(new_n11549_), .B(new_n11638_), .ZN(new_n11639_));
  AOI21_X1   g11447(.A1(new_n11639_), .A2(new_n1632_), .B(new_n11637_), .ZN(new_n11640_));
  NOR3_X1    g11448(.A1(new_n11640_), .A2(\asqrt[50] ), .A3(new_n11599_), .ZN(new_n11641_));
  OAI21_X1   g11449(.A1(new_n11640_), .A2(new_n11599_), .B(\asqrt[50] ), .ZN(new_n11642_));
  OAI21_X1   g11450(.A1(new_n11594_), .A2(new_n11641_), .B(new_n11642_), .ZN(new_n11643_));
  OAI21_X1   g11451(.A1(new_n11643_), .A2(\asqrt[51] ), .B(new_n11589_), .ZN(new_n11644_));
  NAND3_X1   g11452(.A1(new_n11644_), .A2(new_n1150_), .A3(new_n11606_), .ZN(new_n11645_));
  AOI21_X1   g11453(.A1(new_n11644_), .A2(new_n11606_), .B(new_n1150_), .ZN(new_n11646_));
  AOI21_X1   g11454(.A1(new_n11587_), .A2(new_n11645_), .B(new_n11646_), .ZN(new_n11647_));
  AOI21_X1   g11455(.A1(new_n11647_), .A2(new_n1006_), .B(new_n11636_), .ZN(new_n11648_));
  NOR3_X1    g11456(.A1(new_n11648_), .A2(\asqrt[54] ), .A3(new_n11611_), .ZN(new_n11649_));
  OAI21_X1   g11457(.A1(new_n11648_), .A2(new_n11611_), .B(\asqrt[54] ), .ZN(new_n11650_));
  OAI21_X1   g11458(.A1(new_n11582_), .A2(new_n11649_), .B(new_n11650_), .ZN(new_n11651_));
  OAI21_X1   g11459(.A1(new_n11651_), .A2(\asqrt[55] ), .B(new_n11577_), .ZN(new_n11652_));
  NAND3_X1   g11460(.A1(new_n11652_), .A2(new_n634_), .A3(new_n11618_), .ZN(new_n11653_));
  AOI21_X1   g11461(.A1(new_n11652_), .A2(new_n11618_), .B(new_n634_), .ZN(new_n11654_));
  AOI21_X1   g11462(.A1(new_n11575_), .A2(new_n11653_), .B(new_n11654_), .ZN(new_n11655_));
  AOI21_X1   g11463(.A1(new_n11655_), .A2(new_n531_), .B(new_n11635_), .ZN(new_n11656_));
  NOR3_X1    g11464(.A1(new_n11656_), .A2(\asqrt[58] ), .A3(new_n11623_), .ZN(new_n11657_));
  OAI21_X1   g11465(.A1(new_n11656_), .A2(new_n11623_), .B(\asqrt[58] ), .ZN(new_n11658_));
  OAI21_X1   g11466(.A1(new_n11570_), .A2(new_n11657_), .B(new_n11658_), .ZN(new_n11659_));
  OAI21_X1   g11467(.A1(new_n11659_), .A2(\asqrt[59] ), .B(new_n11565_), .ZN(new_n11660_));
  AOI21_X1   g11468(.A1(new_n11660_), .A2(new_n11631_), .B(new_n266_), .ZN(new_n11661_));
  OAI21_X1   g11469(.A1(new_n11634_), .A2(new_n11661_), .B(\asqrt[61] ), .ZN(new_n11662_));
  AOI21_X1   g11470(.A1(new_n11239_), .A2(new_n11233_), .B(\asqrt[17] ), .ZN(new_n11663_));
  XOR2_X1    g11471(.A1(new_n11663_), .A2(new_n11113_), .Z(new_n11664_));
  OAI21_X1   g11472(.A1(new_n11566_), .A2(new_n11629_), .B(new_n11631_), .ZN(new_n11665_));
  OAI21_X1   g11473(.A1(new_n11665_), .A2(\asqrt[60] ), .B(new_n11562_), .ZN(new_n11666_));
  OAI21_X1   g11474(.A1(new_n11630_), .A2(new_n11632_), .B(\asqrt[60] ), .ZN(new_n11667_));
  NAND3_X1   g11475(.A1(new_n11666_), .A2(new_n239_), .A3(new_n11667_), .ZN(new_n11668_));
  NAND2_X1   g11476(.A1(new_n11668_), .A2(new_n11664_), .ZN(new_n11669_));
  NAND2_X1   g11477(.A1(new_n11669_), .A2(new_n11662_), .ZN(new_n11670_));
  AOI21_X1   g11478(.A1(new_n11666_), .A2(new_n11667_), .B(new_n239_), .ZN(new_n11671_));
  NAND3_X1   g11479(.A1(new_n11660_), .A2(new_n266_), .A3(new_n11631_), .ZN(new_n11672_));
  AOI21_X1   g11480(.A1(new_n11562_), .A2(new_n11672_), .B(new_n11661_), .ZN(new_n11673_));
  INV_X1     g11481(.I(new_n11664_), .ZN(new_n11674_));
  AOI21_X1   g11482(.A1(new_n11673_), .A2(new_n239_), .B(new_n11674_), .ZN(new_n11675_));
  OAI21_X1   g11483(.A1(new_n11675_), .A2(new_n11671_), .B(new_n201_), .ZN(new_n11676_));
  NAND3_X1   g11484(.A1(new_n11669_), .A2(\asqrt[62] ), .A3(new_n11662_), .ZN(new_n11677_));
  AOI21_X1   g11485(.A1(new_n11232_), .A2(new_n11356_), .B(\asqrt[17] ), .ZN(new_n11678_));
  XOR2_X1    g11486(.A1(new_n11678_), .A2(new_n11236_), .Z(new_n11679_));
  INV_X1     g11487(.I(new_n11679_), .ZN(new_n11680_));
  AOI22_X1   g11488(.A1(new_n11676_), .A2(new_n11677_), .B1(new_n11670_), .B2(new_n11680_), .ZN(new_n11681_));
  NOR2_X1    g11489(.A1(new_n11251_), .A2(new_n11111_), .ZN(new_n11682_));
  OAI21_X1   g11490(.A1(\asqrt[17] ), .A2(new_n11682_), .B(new_n11258_), .ZN(new_n11683_));
  INV_X1     g11491(.I(new_n11683_), .ZN(new_n11684_));
  OAI21_X1   g11492(.A1(new_n11681_), .A2(new_n11559_), .B(new_n11684_), .ZN(new_n11685_));
  OAI21_X1   g11493(.A1(new_n11670_), .A2(\asqrt[62] ), .B(new_n11679_), .ZN(new_n11686_));
  NAND2_X1   g11494(.A1(new_n11670_), .A2(\asqrt[62] ), .ZN(new_n11687_));
  NAND3_X1   g11495(.A1(new_n11686_), .A2(new_n11687_), .A3(new_n11559_), .ZN(new_n11688_));
  NAND2_X1   g11496(.A1(new_n11373_), .A2(new_n11110_), .ZN(new_n11689_));
  XOR2_X1    g11497(.A1(new_n11251_), .A2(new_n11111_), .Z(new_n11690_));
  NAND3_X1   g11498(.A1(new_n11689_), .A2(\asqrt[63] ), .A3(new_n11690_), .ZN(new_n11691_));
  INV_X1     g11499(.I(new_n11371_), .ZN(new_n11692_));
  NAND4_X1   g11500(.A1(new_n11692_), .A2(new_n11111_), .A3(new_n11258_), .A4(new_n11265_), .ZN(new_n11693_));
  NAND2_X1   g11501(.A1(new_n11691_), .A2(new_n11693_), .ZN(new_n11694_));
  INV_X1     g11502(.I(new_n11694_), .ZN(new_n11695_));
  NAND4_X1   g11503(.A1(new_n11685_), .A2(new_n193_), .A3(new_n11688_), .A4(new_n11695_), .ZN(\asqrt[16] ));
  AOI21_X1   g11504(.A1(new_n11549_), .A2(new_n11553_), .B(\asqrt[16] ), .ZN(new_n11697_));
  XOR2_X1    g11505(.A1(new_n11697_), .A2(new_n11268_), .Z(new_n11698_));
  XOR2_X1    g11506(.A1(new_n11540_), .A2(\asqrt[47] ), .Z(new_n11699_));
  NOR2_X1    g11507(.A1(\asqrt[16] ), .A2(new_n11699_), .ZN(new_n11700_));
  XOR2_X1    g11508(.A1(new_n11700_), .A2(new_n11270_), .Z(new_n11701_));
  NOR2_X1    g11509(.A1(new_n11538_), .A2(new_n11547_), .ZN(new_n11702_));
  NOR2_X1    g11510(.A1(\asqrt[16] ), .A2(new_n11702_), .ZN(new_n11703_));
  XOR2_X1    g11511(.A1(new_n11703_), .A2(new_n11273_), .Z(new_n11704_));
  AOI21_X1   g11512(.A1(new_n11542_), .A2(new_n11546_), .B(\asqrt[16] ), .ZN(new_n11705_));
  XOR2_X1    g11513(.A1(new_n11705_), .A2(new_n11276_), .Z(new_n11706_));
  INV_X1     g11514(.I(new_n11706_), .ZN(new_n11707_));
  AOI21_X1   g11515(.A1(new_n11528_), .A2(new_n11536_), .B(\asqrt[16] ), .ZN(new_n11708_));
  XOR2_X1    g11516(.A1(new_n11708_), .A2(new_n11280_), .Z(new_n11709_));
  INV_X1     g11517(.I(new_n11709_), .ZN(new_n11710_));
  XOR2_X1    g11518(.A1(new_n11519_), .A2(\asqrt[43] ), .Z(new_n11711_));
  NOR2_X1    g11519(.A1(\asqrt[16] ), .A2(new_n11711_), .ZN(new_n11712_));
  XOR2_X1    g11520(.A1(new_n11712_), .A2(new_n11282_), .Z(new_n11713_));
  NOR2_X1    g11521(.A1(new_n11517_), .A2(new_n11526_), .ZN(new_n11714_));
  NOR2_X1    g11522(.A1(\asqrt[16] ), .A2(new_n11714_), .ZN(new_n11715_));
  XOR2_X1    g11523(.A1(new_n11715_), .A2(new_n11285_), .Z(new_n11716_));
  AOI21_X1   g11524(.A1(new_n11521_), .A2(new_n11525_), .B(\asqrt[16] ), .ZN(new_n11717_));
  XOR2_X1    g11525(.A1(new_n11717_), .A2(new_n11288_), .Z(new_n11718_));
  INV_X1     g11526(.I(new_n11718_), .ZN(new_n11719_));
  AOI21_X1   g11527(.A1(new_n11507_), .A2(new_n11515_), .B(\asqrt[16] ), .ZN(new_n11720_));
  XOR2_X1    g11528(.A1(new_n11720_), .A2(new_n11292_), .Z(new_n11721_));
  INV_X1     g11529(.I(new_n11721_), .ZN(new_n11722_));
  XOR2_X1    g11530(.A1(new_n11498_), .A2(\asqrt[39] ), .Z(new_n11723_));
  NOR2_X1    g11531(.A1(\asqrt[16] ), .A2(new_n11723_), .ZN(new_n11724_));
  XOR2_X1    g11532(.A1(new_n11724_), .A2(new_n11294_), .Z(new_n11725_));
  NOR2_X1    g11533(.A1(new_n11496_), .A2(new_n11505_), .ZN(new_n11726_));
  NOR2_X1    g11534(.A1(\asqrt[16] ), .A2(new_n11726_), .ZN(new_n11727_));
  XOR2_X1    g11535(.A1(new_n11727_), .A2(new_n11297_), .Z(new_n11728_));
  AOI21_X1   g11536(.A1(new_n11500_), .A2(new_n11504_), .B(\asqrt[16] ), .ZN(new_n11729_));
  XOR2_X1    g11537(.A1(new_n11729_), .A2(new_n11300_), .Z(new_n11730_));
  INV_X1     g11538(.I(new_n11730_), .ZN(new_n11731_));
  AOI21_X1   g11539(.A1(new_n11486_), .A2(new_n11494_), .B(\asqrt[16] ), .ZN(new_n11732_));
  XOR2_X1    g11540(.A1(new_n11732_), .A2(new_n11304_), .Z(new_n11733_));
  INV_X1     g11541(.I(new_n11733_), .ZN(new_n11734_));
  XOR2_X1    g11542(.A1(new_n11477_), .A2(\asqrt[35] ), .Z(new_n11735_));
  NOR2_X1    g11543(.A1(\asqrt[16] ), .A2(new_n11735_), .ZN(new_n11736_));
  XOR2_X1    g11544(.A1(new_n11736_), .A2(new_n11306_), .Z(new_n11737_));
  NOR2_X1    g11545(.A1(new_n11475_), .A2(new_n11484_), .ZN(new_n11738_));
  NOR2_X1    g11546(.A1(\asqrt[16] ), .A2(new_n11738_), .ZN(new_n11739_));
  XOR2_X1    g11547(.A1(new_n11739_), .A2(new_n11309_), .Z(new_n11740_));
  AOI21_X1   g11548(.A1(new_n11479_), .A2(new_n11483_), .B(\asqrt[16] ), .ZN(new_n11741_));
  XOR2_X1    g11549(.A1(new_n11741_), .A2(new_n11312_), .Z(new_n11742_));
  INV_X1     g11550(.I(new_n11742_), .ZN(new_n11743_));
  AOI21_X1   g11551(.A1(new_n11465_), .A2(new_n11473_), .B(\asqrt[16] ), .ZN(new_n11744_));
  XOR2_X1    g11552(.A1(new_n11744_), .A2(new_n11316_), .Z(new_n11745_));
  INV_X1     g11553(.I(new_n11745_), .ZN(new_n11746_));
  XOR2_X1    g11554(.A1(new_n11456_), .A2(\asqrt[31] ), .Z(new_n11747_));
  NOR2_X1    g11555(.A1(\asqrt[16] ), .A2(new_n11747_), .ZN(new_n11748_));
  XOR2_X1    g11556(.A1(new_n11748_), .A2(new_n11318_), .Z(new_n11749_));
  NOR2_X1    g11557(.A1(new_n11454_), .A2(new_n11463_), .ZN(new_n11750_));
  NOR2_X1    g11558(.A1(\asqrt[16] ), .A2(new_n11750_), .ZN(new_n11751_));
  XOR2_X1    g11559(.A1(new_n11751_), .A2(new_n11321_), .Z(new_n11752_));
  AOI21_X1   g11560(.A1(new_n11458_), .A2(new_n11462_), .B(\asqrt[16] ), .ZN(new_n11753_));
  XOR2_X1    g11561(.A1(new_n11753_), .A2(new_n11324_), .Z(new_n11754_));
  INV_X1     g11562(.I(new_n11754_), .ZN(new_n11755_));
  AOI21_X1   g11563(.A1(new_n11444_), .A2(new_n11452_), .B(\asqrt[16] ), .ZN(new_n11756_));
  XOR2_X1    g11564(.A1(new_n11756_), .A2(new_n11328_), .Z(new_n11757_));
  INV_X1     g11565(.I(new_n11757_), .ZN(new_n11758_));
  XOR2_X1    g11566(.A1(new_n11435_), .A2(\asqrt[27] ), .Z(new_n11759_));
  NOR2_X1    g11567(.A1(\asqrt[16] ), .A2(new_n11759_), .ZN(new_n11760_));
  XOR2_X1    g11568(.A1(new_n11760_), .A2(new_n11330_), .Z(new_n11761_));
  NOR2_X1    g11569(.A1(new_n11433_), .A2(new_n11442_), .ZN(new_n11762_));
  NOR2_X1    g11570(.A1(\asqrt[16] ), .A2(new_n11762_), .ZN(new_n11763_));
  XOR2_X1    g11571(.A1(new_n11763_), .A2(new_n11333_), .Z(new_n11764_));
  AOI21_X1   g11572(.A1(new_n11437_), .A2(new_n11441_), .B(\asqrt[16] ), .ZN(new_n11765_));
  XOR2_X1    g11573(.A1(new_n11765_), .A2(new_n11336_), .Z(new_n11766_));
  INV_X1     g11574(.I(new_n11766_), .ZN(new_n11767_));
  AOI21_X1   g11575(.A1(new_n11423_), .A2(new_n11431_), .B(\asqrt[16] ), .ZN(new_n11768_));
  XOR2_X1    g11576(.A1(new_n11768_), .A2(new_n11340_), .Z(new_n11769_));
  INV_X1     g11577(.I(new_n11769_), .ZN(new_n11770_));
  XOR2_X1    g11578(.A1(new_n11414_), .A2(\asqrt[23] ), .Z(new_n11771_));
  NOR2_X1    g11579(.A1(\asqrt[16] ), .A2(new_n11771_), .ZN(new_n11772_));
  XOR2_X1    g11580(.A1(new_n11772_), .A2(new_n11342_), .Z(new_n11773_));
  NOR2_X1    g11581(.A1(new_n11412_), .A2(new_n11421_), .ZN(new_n11774_));
  NOR2_X1    g11582(.A1(\asqrt[16] ), .A2(new_n11774_), .ZN(new_n11775_));
  XOR2_X1    g11583(.A1(new_n11775_), .A2(new_n11345_), .Z(new_n11776_));
  AOI21_X1   g11584(.A1(new_n11416_), .A2(new_n11420_), .B(\asqrt[16] ), .ZN(new_n11777_));
  XOR2_X1    g11585(.A1(new_n11777_), .A2(new_n11348_), .Z(new_n11778_));
  INV_X1     g11586(.I(new_n11778_), .ZN(new_n11779_));
  AOI21_X1   g11587(.A1(new_n11402_), .A2(new_n11410_), .B(\asqrt[16] ), .ZN(new_n11780_));
  XOR2_X1    g11588(.A1(new_n11780_), .A2(new_n11355_), .Z(new_n11781_));
  INV_X1     g11589(.I(new_n11781_), .ZN(new_n11782_));
  AOI21_X1   g11590(.A1(new_n11392_), .A2(new_n11401_), .B(\asqrt[16] ), .ZN(new_n11783_));
  XOR2_X1    g11591(.A1(new_n11783_), .A2(new_n11376_), .Z(new_n11784_));
  NAND2_X1   g11592(.A1(\asqrt[17] ), .A2(new_n11377_), .ZN(new_n11785_));
  NOR2_X1    g11593(.A1(new_n11389_), .A2(\a[34] ), .ZN(new_n11786_));
  AOI22_X1   g11594(.A1(new_n11785_), .A2(new_n11389_), .B1(\asqrt[17] ), .B2(new_n11786_), .ZN(new_n11787_));
  OAI21_X1   g11595(.A1(new_n11373_), .A2(new_n11377_), .B(new_n11386_), .ZN(new_n11788_));
  AOI21_X1   g11596(.A1(new_n11382_), .A2(new_n11788_), .B(\asqrt[16] ), .ZN(new_n11789_));
  XOR2_X1    g11597(.A1(new_n11789_), .A2(new_n11787_), .Z(new_n11790_));
  NAND2_X1   g11598(.A1(new_n11685_), .A2(new_n193_), .ZN(new_n11791_));
  NOR2_X1    g11599(.A1(new_n11675_), .A2(new_n11671_), .ZN(new_n11792_));
  AOI21_X1   g11600(.A1(new_n11792_), .A2(new_n201_), .B(new_n11680_), .ZN(new_n11793_));
  OAI21_X1   g11601(.A1(new_n11792_), .A2(new_n201_), .B(new_n11559_), .ZN(new_n11794_));
  NOR2_X1    g11602(.A1(new_n11793_), .A2(new_n11794_), .ZN(new_n11795_));
  NAND3_X1   g11603(.A1(new_n11691_), .A2(\asqrt[17] ), .A3(new_n11693_), .ZN(new_n11796_));
  NOR3_X1    g11604(.A1(new_n11791_), .A2(new_n11795_), .A3(new_n11796_), .ZN(new_n11797_));
  AOI21_X1   g11605(.A1(new_n11669_), .A2(new_n11662_), .B(\asqrt[62] ), .ZN(new_n11798_));
  NOR3_X1    g11606(.A1(new_n11675_), .A2(new_n201_), .A3(new_n11671_), .ZN(new_n11799_));
  OAI22_X1   g11607(.A1(new_n11799_), .A2(new_n11798_), .B1(new_n11792_), .B2(new_n11679_), .ZN(new_n11800_));
  AOI21_X1   g11608(.A1(new_n11800_), .A2(new_n11558_), .B(new_n11683_), .ZN(new_n11801_));
  NOR4_X1    g11609(.A1(new_n11801_), .A2(\asqrt[63] ), .A3(new_n11795_), .A4(new_n11694_), .ZN(new_n11802_));
  NOR2_X1    g11610(.A1(new_n11802_), .A2(new_n11380_), .ZN(new_n11803_));
  OAI21_X1   g11611(.A1(new_n11803_), .A2(new_n11797_), .B(new_n11377_), .ZN(new_n11804_));
  NOR3_X1    g11612(.A1(new_n11801_), .A2(\asqrt[63] ), .A3(new_n11795_), .ZN(new_n11805_));
  NAND4_X1   g11613(.A1(new_n11805_), .A2(\asqrt[17] ), .A3(new_n11691_), .A4(new_n11693_), .ZN(new_n11806_));
  NAND2_X1   g11614(.A1(\asqrt[16] ), .A2(new_n11378_), .ZN(new_n11807_));
  NAND3_X1   g11615(.A1(new_n11806_), .A2(new_n11807_), .A3(\a[34] ), .ZN(new_n11808_));
  NAND2_X1   g11616(.A1(new_n11808_), .A2(new_n11804_), .ZN(new_n11809_));
  NOR2_X1    g11617(.A1(\a[30] ), .A2(\a[31] ), .ZN(new_n11810_));
  INV_X1     g11618(.I(new_n11810_), .ZN(new_n11811_));
  NAND3_X1   g11619(.A1(\asqrt[16] ), .A2(\a[32] ), .A3(new_n11811_), .ZN(new_n11812_));
  INV_X1     g11620(.I(\a[32] ), .ZN(new_n11813_));
  OAI21_X1   g11621(.A1(\asqrt[16] ), .A2(new_n11813_), .B(new_n11810_), .ZN(new_n11814_));
  AOI21_X1   g11622(.A1(new_n11814_), .A2(new_n11812_), .B(new_n11373_), .ZN(new_n11815_));
  NAND2_X1   g11623(.A1(new_n11810_), .A2(new_n11813_), .ZN(new_n11816_));
  NAND3_X1   g11624(.A1(new_n11261_), .A2(new_n11263_), .A3(new_n11816_), .ZN(new_n11817_));
  NAND2_X1   g11625(.A1(new_n11365_), .A2(new_n11817_), .ZN(new_n11818_));
  NAND3_X1   g11626(.A1(\asqrt[16] ), .A2(\a[32] ), .A3(new_n11818_), .ZN(new_n11819_));
  INV_X1     g11627(.I(\a[33] ), .ZN(new_n11820_));
  NAND3_X1   g11628(.A1(\asqrt[16] ), .A2(new_n11813_), .A3(new_n11820_), .ZN(new_n11821_));
  OAI21_X1   g11629(.A1(new_n11802_), .A2(\a[32] ), .B(\a[33] ), .ZN(new_n11822_));
  NAND3_X1   g11630(.A1(new_n11822_), .A2(new_n11819_), .A3(new_n11821_), .ZN(new_n11823_));
  NOR3_X1    g11631(.A1(new_n11823_), .A2(new_n11815_), .A3(\asqrt[18] ), .ZN(new_n11824_));
  OAI21_X1   g11632(.A1(new_n11823_), .A2(new_n11815_), .B(\asqrt[18] ), .ZN(new_n11825_));
  OAI21_X1   g11633(.A1(new_n11809_), .A2(new_n11824_), .B(new_n11825_), .ZN(new_n11826_));
  OAI21_X1   g11634(.A1(new_n11826_), .A2(\asqrt[19] ), .B(new_n11790_), .ZN(new_n11827_));
  NAND2_X1   g11635(.A1(new_n11826_), .A2(\asqrt[19] ), .ZN(new_n11828_));
  NAND3_X1   g11636(.A1(new_n11827_), .A2(new_n11828_), .A3(new_n10052_), .ZN(new_n11829_));
  AOI21_X1   g11637(.A1(new_n11827_), .A2(new_n11828_), .B(new_n10052_), .ZN(new_n11830_));
  AOI21_X1   g11638(.A1(new_n11784_), .A2(new_n11829_), .B(new_n11830_), .ZN(new_n11831_));
  AOI21_X1   g11639(.A1(new_n11831_), .A2(new_n9656_), .B(new_n11782_), .ZN(new_n11832_));
  NAND2_X1   g11640(.A1(new_n11829_), .A2(new_n11784_), .ZN(new_n11833_));
  INV_X1     g11641(.I(new_n11790_), .ZN(new_n11834_));
  INV_X1     g11642(.I(new_n11809_), .ZN(new_n11835_));
  NOR3_X1    g11643(.A1(new_n11802_), .A2(new_n11813_), .A3(new_n11810_), .ZN(new_n11836_));
  AOI21_X1   g11644(.A1(new_n11802_), .A2(\a[32] ), .B(new_n11811_), .ZN(new_n11837_));
  OAI21_X1   g11645(.A1(new_n11836_), .A2(new_n11837_), .B(\asqrt[17] ), .ZN(new_n11838_));
  INV_X1     g11646(.I(new_n11818_), .ZN(new_n11839_));
  NOR3_X1    g11647(.A1(new_n11802_), .A2(new_n11813_), .A3(new_n11839_), .ZN(new_n11840_));
  NOR3_X1    g11648(.A1(new_n11802_), .A2(\a[32] ), .A3(\a[33] ), .ZN(new_n11841_));
  AOI21_X1   g11649(.A1(\asqrt[16] ), .A2(new_n11813_), .B(new_n11820_), .ZN(new_n11842_));
  NOR3_X1    g11650(.A1(new_n11840_), .A2(new_n11841_), .A3(new_n11842_), .ZN(new_n11843_));
  NAND3_X1   g11651(.A1(new_n11838_), .A2(new_n11843_), .A3(new_n10914_), .ZN(new_n11844_));
  AOI21_X1   g11652(.A1(new_n11838_), .A2(new_n11843_), .B(new_n10914_), .ZN(new_n11845_));
  AOI21_X1   g11653(.A1(new_n11835_), .A2(new_n11844_), .B(new_n11845_), .ZN(new_n11846_));
  AOI21_X1   g11654(.A1(new_n11846_), .A2(new_n10497_), .B(new_n11834_), .ZN(new_n11847_));
  NAND2_X1   g11655(.A1(new_n11835_), .A2(new_n11844_), .ZN(new_n11848_));
  AOI21_X1   g11656(.A1(new_n11848_), .A2(new_n11825_), .B(new_n10497_), .ZN(new_n11849_));
  OAI21_X1   g11657(.A1(new_n11847_), .A2(new_n11849_), .B(\asqrt[20] ), .ZN(new_n11850_));
  AOI21_X1   g11658(.A1(new_n11833_), .A2(new_n11850_), .B(new_n9656_), .ZN(new_n11851_));
  NOR3_X1    g11659(.A1(new_n11832_), .A2(\asqrt[22] ), .A3(new_n11851_), .ZN(new_n11852_));
  OAI21_X1   g11660(.A1(new_n11832_), .A2(new_n11851_), .B(\asqrt[22] ), .ZN(new_n11853_));
  OAI21_X1   g11661(.A1(new_n11779_), .A2(new_n11852_), .B(new_n11853_), .ZN(new_n11854_));
  OAI21_X1   g11662(.A1(new_n11854_), .A2(\asqrt[23] ), .B(new_n11776_), .ZN(new_n11855_));
  NAND2_X1   g11663(.A1(new_n11854_), .A2(\asqrt[23] ), .ZN(new_n11856_));
  NAND3_X1   g11664(.A1(new_n11855_), .A2(new_n11856_), .A3(new_n8440_), .ZN(new_n11857_));
  AOI21_X1   g11665(.A1(new_n11855_), .A2(new_n11856_), .B(new_n8440_), .ZN(new_n11858_));
  AOI21_X1   g11666(.A1(new_n11773_), .A2(new_n11857_), .B(new_n11858_), .ZN(new_n11859_));
  AOI21_X1   g11667(.A1(new_n11859_), .A2(new_n8077_), .B(new_n11770_), .ZN(new_n11860_));
  NAND2_X1   g11668(.A1(new_n11857_), .A2(new_n11773_), .ZN(new_n11861_));
  INV_X1     g11669(.I(new_n11776_), .ZN(new_n11862_));
  INV_X1     g11670(.I(new_n11784_), .ZN(new_n11863_));
  NOR3_X1    g11671(.A1(new_n11847_), .A2(\asqrt[20] ), .A3(new_n11849_), .ZN(new_n11864_));
  OAI21_X1   g11672(.A1(new_n11863_), .A2(new_n11864_), .B(new_n11850_), .ZN(new_n11865_));
  OAI21_X1   g11673(.A1(new_n11865_), .A2(\asqrt[21] ), .B(new_n11781_), .ZN(new_n11866_));
  NAND2_X1   g11674(.A1(new_n11865_), .A2(\asqrt[21] ), .ZN(new_n11867_));
  NAND3_X1   g11675(.A1(new_n11866_), .A2(new_n11867_), .A3(new_n9233_), .ZN(new_n11868_));
  AOI21_X1   g11676(.A1(new_n11866_), .A2(new_n11867_), .B(new_n9233_), .ZN(new_n11869_));
  AOI21_X1   g11677(.A1(new_n11778_), .A2(new_n11868_), .B(new_n11869_), .ZN(new_n11870_));
  AOI21_X1   g11678(.A1(new_n11870_), .A2(new_n8849_), .B(new_n11862_), .ZN(new_n11871_));
  NAND2_X1   g11679(.A1(new_n11868_), .A2(new_n11778_), .ZN(new_n11872_));
  AOI21_X1   g11680(.A1(new_n11872_), .A2(new_n11853_), .B(new_n8849_), .ZN(new_n11873_));
  OAI21_X1   g11681(.A1(new_n11871_), .A2(new_n11873_), .B(\asqrt[24] ), .ZN(new_n11874_));
  AOI21_X1   g11682(.A1(new_n11861_), .A2(new_n11874_), .B(new_n8077_), .ZN(new_n11875_));
  NOR3_X1    g11683(.A1(new_n11860_), .A2(\asqrt[26] ), .A3(new_n11875_), .ZN(new_n11876_));
  OAI21_X1   g11684(.A1(new_n11860_), .A2(new_n11875_), .B(\asqrt[26] ), .ZN(new_n11877_));
  OAI21_X1   g11685(.A1(new_n11767_), .A2(new_n11876_), .B(new_n11877_), .ZN(new_n11878_));
  OAI21_X1   g11686(.A1(new_n11878_), .A2(\asqrt[27] ), .B(new_n11764_), .ZN(new_n11879_));
  NAND2_X1   g11687(.A1(new_n11878_), .A2(\asqrt[27] ), .ZN(new_n11880_));
  NAND3_X1   g11688(.A1(new_n11879_), .A2(new_n11880_), .A3(new_n6966_), .ZN(new_n11881_));
  AOI21_X1   g11689(.A1(new_n11879_), .A2(new_n11880_), .B(new_n6966_), .ZN(new_n11882_));
  AOI21_X1   g11690(.A1(new_n11761_), .A2(new_n11881_), .B(new_n11882_), .ZN(new_n11883_));
  AOI21_X1   g11691(.A1(new_n11883_), .A2(new_n6636_), .B(new_n11758_), .ZN(new_n11884_));
  NAND2_X1   g11692(.A1(new_n11881_), .A2(new_n11761_), .ZN(new_n11885_));
  INV_X1     g11693(.I(new_n11764_), .ZN(new_n11886_));
  INV_X1     g11694(.I(new_n11773_), .ZN(new_n11887_));
  NOR3_X1    g11695(.A1(new_n11871_), .A2(\asqrt[24] ), .A3(new_n11873_), .ZN(new_n11888_));
  OAI21_X1   g11696(.A1(new_n11887_), .A2(new_n11888_), .B(new_n11874_), .ZN(new_n11889_));
  OAI21_X1   g11697(.A1(new_n11889_), .A2(\asqrt[25] ), .B(new_n11769_), .ZN(new_n11890_));
  NAND2_X1   g11698(.A1(new_n11889_), .A2(\asqrt[25] ), .ZN(new_n11891_));
  NAND3_X1   g11699(.A1(new_n11890_), .A2(new_n11891_), .A3(new_n7690_), .ZN(new_n11892_));
  AOI21_X1   g11700(.A1(new_n11890_), .A2(new_n11891_), .B(new_n7690_), .ZN(new_n11893_));
  AOI21_X1   g11701(.A1(new_n11766_), .A2(new_n11892_), .B(new_n11893_), .ZN(new_n11894_));
  AOI21_X1   g11702(.A1(new_n11894_), .A2(new_n7331_), .B(new_n11886_), .ZN(new_n11895_));
  NAND2_X1   g11703(.A1(new_n11892_), .A2(new_n11766_), .ZN(new_n11896_));
  AOI21_X1   g11704(.A1(new_n11896_), .A2(new_n11877_), .B(new_n7331_), .ZN(new_n11897_));
  OAI21_X1   g11705(.A1(new_n11895_), .A2(new_n11897_), .B(\asqrt[28] ), .ZN(new_n11898_));
  AOI21_X1   g11706(.A1(new_n11885_), .A2(new_n11898_), .B(new_n6636_), .ZN(new_n11899_));
  NOR3_X1    g11707(.A1(new_n11884_), .A2(\asqrt[30] ), .A3(new_n11899_), .ZN(new_n11900_));
  OAI21_X1   g11708(.A1(new_n11884_), .A2(new_n11899_), .B(\asqrt[30] ), .ZN(new_n11901_));
  OAI21_X1   g11709(.A1(new_n11755_), .A2(new_n11900_), .B(new_n11901_), .ZN(new_n11902_));
  OAI21_X1   g11710(.A1(new_n11902_), .A2(\asqrt[31] ), .B(new_n11752_), .ZN(new_n11903_));
  NAND2_X1   g11711(.A1(new_n11902_), .A2(\asqrt[31] ), .ZN(new_n11904_));
  NAND3_X1   g11712(.A1(new_n11903_), .A2(new_n11904_), .A3(new_n5643_), .ZN(new_n11905_));
  AOI21_X1   g11713(.A1(new_n11903_), .A2(new_n11904_), .B(new_n5643_), .ZN(new_n11906_));
  AOI21_X1   g11714(.A1(new_n11749_), .A2(new_n11905_), .B(new_n11906_), .ZN(new_n11907_));
  AOI21_X1   g11715(.A1(new_n11907_), .A2(new_n5336_), .B(new_n11746_), .ZN(new_n11908_));
  NAND2_X1   g11716(.A1(new_n11905_), .A2(new_n11749_), .ZN(new_n11909_));
  INV_X1     g11717(.I(new_n11752_), .ZN(new_n11910_));
  INV_X1     g11718(.I(new_n11761_), .ZN(new_n11911_));
  NOR3_X1    g11719(.A1(new_n11895_), .A2(\asqrt[28] ), .A3(new_n11897_), .ZN(new_n11912_));
  OAI21_X1   g11720(.A1(new_n11911_), .A2(new_n11912_), .B(new_n11898_), .ZN(new_n11913_));
  OAI21_X1   g11721(.A1(new_n11913_), .A2(\asqrt[29] ), .B(new_n11757_), .ZN(new_n11914_));
  NAND2_X1   g11722(.A1(new_n11913_), .A2(\asqrt[29] ), .ZN(new_n11915_));
  NAND3_X1   g11723(.A1(new_n11914_), .A2(new_n11915_), .A3(new_n6275_), .ZN(new_n11916_));
  AOI21_X1   g11724(.A1(new_n11914_), .A2(new_n11915_), .B(new_n6275_), .ZN(new_n11917_));
  AOI21_X1   g11725(.A1(new_n11754_), .A2(new_n11916_), .B(new_n11917_), .ZN(new_n11918_));
  AOI21_X1   g11726(.A1(new_n11918_), .A2(new_n5947_), .B(new_n11910_), .ZN(new_n11919_));
  NAND2_X1   g11727(.A1(new_n11916_), .A2(new_n11754_), .ZN(new_n11920_));
  AOI21_X1   g11728(.A1(new_n11920_), .A2(new_n11901_), .B(new_n5947_), .ZN(new_n11921_));
  OAI21_X1   g11729(.A1(new_n11919_), .A2(new_n11921_), .B(\asqrt[32] ), .ZN(new_n11922_));
  AOI21_X1   g11730(.A1(new_n11909_), .A2(new_n11922_), .B(new_n5336_), .ZN(new_n11923_));
  NOR3_X1    g11731(.A1(new_n11908_), .A2(\asqrt[34] ), .A3(new_n11923_), .ZN(new_n11924_));
  OAI21_X1   g11732(.A1(new_n11908_), .A2(new_n11923_), .B(\asqrt[34] ), .ZN(new_n11925_));
  OAI21_X1   g11733(.A1(new_n11743_), .A2(new_n11924_), .B(new_n11925_), .ZN(new_n11926_));
  OAI21_X1   g11734(.A1(new_n11926_), .A2(\asqrt[35] ), .B(new_n11740_), .ZN(new_n11927_));
  NAND2_X1   g11735(.A1(new_n11926_), .A2(\asqrt[35] ), .ZN(new_n11928_));
  NAND3_X1   g11736(.A1(new_n11927_), .A2(new_n11928_), .A3(new_n4461_), .ZN(new_n11929_));
  AOI21_X1   g11737(.A1(new_n11927_), .A2(new_n11928_), .B(new_n4461_), .ZN(new_n11930_));
  AOI21_X1   g11738(.A1(new_n11737_), .A2(new_n11929_), .B(new_n11930_), .ZN(new_n11931_));
  AOI21_X1   g11739(.A1(new_n11931_), .A2(new_n4196_), .B(new_n11734_), .ZN(new_n11932_));
  NAND2_X1   g11740(.A1(new_n11929_), .A2(new_n11737_), .ZN(new_n11933_));
  INV_X1     g11741(.I(new_n11740_), .ZN(new_n11934_));
  INV_X1     g11742(.I(new_n11749_), .ZN(new_n11935_));
  NOR3_X1    g11743(.A1(new_n11919_), .A2(\asqrt[32] ), .A3(new_n11921_), .ZN(new_n11936_));
  OAI21_X1   g11744(.A1(new_n11935_), .A2(new_n11936_), .B(new_n11922_), .ZN(new_n11937_));
  OAI21_X1   g11745(.A1(new_n11937_), .A2(\asqrt[33] ), .B(new_n11745_), .ZN(new_n11938_));
  NAND2_X1   g11746(.A1(new_n11937_), .A2(\asqrt[33] ), .ZN(new_n11939_));
  NAND3_X1   g11747(.A1(new_n11938_), .A2(new_n11939_), .A3(new_n5029_), .ZN(new_n11940_));
  AOI21_X1   g11748(.A1(new_n11938_), .A2(new_n11939_), .B(new_n5029_), .ZN(new_n11941_));
  AOI21_X1   g11749(.A1(new_n11742_), .A2(new_n11940_), .B(new_n11941_), .ZN(new_n11942_));
  AOI21_X1   g11750(.A1(new_n11942_), .A2(new_n4751_), .B(new_n11934_), .ZN(new_n11943_));
  NAND2_X1   g11751(.A1(new_n11940_), .A2(new_n11742_), .ZN(new_n11944_));
  AOI21_X1   g11752(.A1(new_n11944_), .A2(new_n11925_), .B(new_n4751_), .ZN(new_n11945_));
  OAI21_X1   g11753(.A1(new_n11943_), .A2(new_n11945_), .B(\asqrt[36] ), .ZN(new_n11946_));
  AOI21_X1   g11754(.A1(new_n11933_), .A2(new_n11946_), .B(new_n4196_), .ZN(new_n11947_));
  NOR3_X1    g11755(.A1(new_n11932_), .A2(\asqrt[38] ), .A3(new_n11947_), .ZN(new_n11948_));
  OAI21_X1   g11756(.A1(new_n11932_), .A2(new_n11947_), .B(\asqrt[38] ), .ZN(new_n11949_));
  OAI21_X1   g11757(.A1(new_n11731_), .A2(new_n11948_), .B(new_n11949_), .ZN(new_n11950_));
  OAI21_X1   g11758(.A1(new_n11950_), .A2(\asqrt[39] ), .B(new_n11728_), .ZN(new_n11951_));
  NAND2_X1   g11759(.A1(new_n11950_), .A2(\asqrt[39] ), .ZN(new_n11952_));
  NAND3_X1   g11760(.A1(new_n11951_), .A2(new_n11952_), .A3(new_n3427_), .ZN(new_n11953_));
  AOI21_X1   g11761(.A1(new_n11951_), .A2(new_n11952_), .B(new_n3427_), .ZN(new_n11954_));
  AOI21_X1   g11762(.A1(new_n11725_), .A2(new_n11953_), .B(new_n11954_), .ZN(new_n11955_));
  AOI21_X1   g11763(.A1(new_n11955_), .A2(new_n3195_), .B(new_n11722_), .ZN(new_n11956_));
  NAND2_X1   g11764(.A1(new_n11953_), .A2(new_n11725_), .ZN(new_n11957_));
  INV_X1     g11765(.I(new_n11728_), .ZN(new_n11958_));
  INV_X1     g11766(.I(new_n11737_), .ZN(new_n11959_));
  NOR3_X1    g11767(.A1(new_n11943_), .A2(\asqrt[36] ), .A3(new_n11945_), .ZN(new_n11960_));
  OAI21_X1   g11768(.A1(new_n11959_), .A2(new_n11960_), .B(new_n11946_), .ZN(new_n11961_));
  OAI21_X1   g11769(.A1(new_n11961_), .A2(\asqrt[37] ), .B(new_n11733_), .ZN(new_n11962_));
  NAND2_X1   g11770(.A1(new_n11961_), .A2(\asqrt[37] ), .ZN(new_n11963_));
  NAND3_X1   g11771(.A1(new_n11962_), .A2(new_n11963_), .A3(new_n3925_), .ZN(new_n11964_));
  AOI21_X1   g11772(.A1(new_n11962_), .A2(new_n11963_), .B(new_n3925_), .ZN(new_n11965_));
  AOI21_X1   g11773(.A1(new_n11730_), .A2(new_n11964_), .B(new_n11965_), .ZN(new_n11966_));
  AOI21_X1   g11774(.A1(new_n11966_), .A2(new_n3681_), .B(new_n11958_), .ZN(new_n11967_));
  NAND2_X1   g11775(.A1(new_n11964_), .A2(new_n11730_), .ZN(new_n11968_));
  AOI21_X1   g11776(.A1(new_n11968_), .A2(new_n11949_), .B(new_n3681_), .ZN(new_n11969_));
  OAI21_X1   g11777(.A1(new_n11967_), .A2(new_n11969_), .B(\asqrt[40] ), .ZN(new_n11970_));
  AOI21_X1   g11778(.A1(new_n11957_), .A2(new_n11970_), .B(new_n3195_), .ZN(new_n11971_));
  NOR3_X1    g11779(.A1(new_n11956_), .A2(\asqrt[42] ), .A3(new_n11971_), .ZN(new_n11972_));
  OAI21_X1   g11780(.A1(new_n11956_), .A2(new_n11971_), .B(\asqrt[42] ), .ZN(new_n11973_));
  OAI21_X1   g11781(.A1(new_n11719_), .A2(new_n11972_), .B(new_n11973_), .ZN(new_n11974_));
  OAI21_X1   g11782(.A1(new_n11974_), .A2(\asqrt[43] ), .B(new_n11716_), .ZN(new_n11975_));
  NAND2_X1   g11783(.A1(new_n11974_), .A2(\asqrt[43] ), .ZN(new_n11976_));
  NAND3_X1   g11784(.A1(new_n11975_), .A2(new_n11976_), .A3(new_n2531_), .ZN(new_n11977_));
  AOI21_X1   g11785(.A1(new_n11975_), .A2(new_n11976_), .B(new_n2531_), .ZN(new_n11978_));
  AOI21_X1   g11786(.A1(new_n11713_), .A2(new_n11977_), .B(new_n11978_), .ZN(new_n11979_));
  AOI21_X1   g11787(.A1(new_n11979_), .A2(new_n2332_), .B(new_n11710_), .ZN(new_n11980_));
  NAND2_X1   g11788(.A1(new_n11977_), .A2(new_n11713_), .ZN(new_n11981_));
  INV_X1     g11789(.I(new_n11716_), .ZN(new_n11982_));
  INV_X1     g11790(.I(new_n11725_), .ZN(new_n11983_));
  NOR3_X1    g11791(.A1(new_n11967_), .A2(\asqrt[40] ), .A3(new_n11969_), .ZN(new_n11984_));
  OAI21_X1   g11792(.A1(new_n11983_), .A2(new_n11984_), .B(new_n11970_), .ZN(new_n11985_));
  OAI21_X1   g11793(.A1(new_n11985_), .A2(\asqrt[41] ), .B(new_n11721_), .ZN(new_n11986_));
  NAND2_X1   g11794(.A1(new_n11985_), .A2(\asqrt[41] ), .ZN(new_n11987_));
  NAND3_X1   g11795(.A1(new_n11986_), .A2(new_n11987_), .A3(new_n2960_), .ZN(new_n11988_));
  AOI21_X1   g11796(.A1(new_n11986_), .A2(new_n11987_), .B(new_n2960_), .ZN(new_n11989_));
  AOI21_X1   g11797(.A1(new_n11718_), .A2(new_n11988_), .B(new_n11989_), .ZN(new_n11990_));
  AOI21_X1   g11798(.A1(new_n11990_), .A2(new_n2749_), .B(new_n11982_), .ZN(new_n11991_));
  NAND2_X1   g11799(.A1(new_n11988_), .A2(new_n11718_), .ZN(new_n11992_));
  AOI21_X1   g11800(.A1(new_n11992_), .A2(new_n11973_), .B(new_n2749_), .ZN(new_n11993_));
  OAI21_X1   g11801(.A1(new_n11991_), .A2(new_n11993_), .B(\asqrt[44] ), .ZN(new_n11994_));
  AOI21_X1   g11802(.A1(new_n11981_), .A2(new_n11994_), .B(new_n2332_), .ZN(new_n11995_));
  NOR3_X1    g11803(.A1(new_n11980_), .A2(\asqrt[46] ), .A3(new_n11995_), .ZN(new_n11996_));
  OAI21_X1   g11804(.A1(new_n11980_), .A2(new_n11995_), .B(\asqrt[46] ), .ZN(new_n11997_));
  OAI21_X1   g11805(.A1(new_n11707_), .A2(new_n11996_), .B(new_n11997_), .ZN(new_n11998_));
  OAI21_X1   g11806(.A1(new_n11998_), .A2(\asqrt[47] ), .B(new_n11704_), .ZN(new_n11999_));
  NAND2_X1   g11807(.A1(new_n11998_), .A2(\asqrt[47] ), .ZN(new_n12000_));
  NAND3_X1   g11808(.A1(new_n11999_), .A2(new_n12000_), .A3(new_n1778_), .ZN(new_n12001_));
  AOI21_X1   g11809(.A1(new_n11999_), .A2(new_n12000_), .B(new_n1778_), .ZN(new_n12002_));
  AOI21_X1   g11810(.A1(new_n11701_), .A2(new_n12001_), .B(new_n12002_), .ZN(new_n12003_));
  NAND2_X1   g11811(.A1(new_n12003_), .A2(new_n1632_), .ZN(new_n12004_));
  INV_X1     g11812(.I(new_n11701_), .ZN(new_n12005_));
  INV_X1     g11813(.I(new_n11704_), .ZN(new_n12006_));
  INV_X1     g11814(.I(new_n11713_), .ZN(new_n12007_));
  NOR3_X1    g11815(.A1(new_n11991_), .A2(\asqrt[44] ), .A3(new_n11993_), .ZN(new_n12008_));
  OAI21_X1   g11816(.A1(new_n12007_), .A2(new_n12008_), .B(new_n11994_), .ZN(new_n12009_));
  OAI21_X1   g11817(.A1(new_n12009_), .A2(\asqrt[45] ), .B(new_n11709_), .ZN(new_n12010_));
  NAND2_X1   g11818(.A1(new_n12009_), .A2(\asqrt[45] ), .ZN(new_n12011_));
  NAND3_X1   g11819(.A1(new_n12010_), .A2(new_n12011_), .A3(new_n2134_), .ZN(new_n12012_));
  AOI21_X1   g11820(.A1(new_n12010_), .A2(new_n12011_), .B(new_n2134_), .ZN(new_n12013_));
  AOI21_X1   g11821(.A1(new_n11706_), .A2(new_n12012_), .B(new_n12013_), .ZN(new_n12014_));
  AOI21_X1   g11822(.A1(new_n12014_), .A2(new_n1953_), .B(new_n12006_), .ZN(new_n12015_));
  NAND2_X1   g11823(.A1(new_n12012_), .A2(new_n11706_), .ZN(new_n12016_));
  AOI21_X1   g11824(.A1(new_n12016_), .A2(new_n11997_), .B(new_n1953_), .ZN(new_n12017_));
  NOR3_X1    g11825(.A1(new_n12015_), .A2(\asqrt[48] ), .A3(new_n12017_), .ZN(new_n12018_));
  OAI21_X1   g11826(.A1(new_n12015_), .A2(new_n12017_), .B(\asqrt[48] ), .ZN(new_n12019_));
  OAI21_X1   g11827(.A1(new_n12005_), .A2(new_n12018_), .B(new_n12019_), .ZN(new_n12020_));
  NAND2_X1   g11828(.A1(new_n12020_), .A2(\asqrt[49] ), .ZN(new_n12021_));
  NOR2_X1    g11829(.A1(new_n11670_), .A2(\asqrt[62] ), .ZN(new_n12022_));
  INV_X1     g11830(.I(new_n11687_), .ZN(new_n12023_));
  NOR2_X1    g11831(.A1(new_n12023_), .A2(new_n12022_), .ZN(new_n12024_));
  XOR2_X1    g11832(.A1(new_n11678_), .A2(new_n11236_), .Z(new_n12025_));
  OAI21_X1   g11833(.A1(\asqrt[16] ), .A2(new_n12024_), .B(new_n12025_), .ZN(new_n12026_));
  INV_X1     g11834(.I(new_n12026_), .ZN(new_n12027_));
  NOR2_X1    g11835(.A1(new_n11632_), .A2(new_n11629_), .ZN(new_n12028_));
  NOR2_X1    g11836(.A1(\asqrt[16] ), .A2(new_n12028_), .ZN(new_n12029_));
  XOR2_X1    g11837(.A1(new_n12029_), .A2(new_n11565_), .Z(new_n12030_));
  INV_X1     g11838(.I(new_n12030_), .ZN(new_n12031_));
  NOR2_X1    g11839(.A1(new_n11657_), .A2(new_n11628_), .ZN(new_n12032_));
  NOR2_X1    g11840(.A1(\asqrt[16] ), .A2(new_n12032_), .ZN(new_n12033_));
  XOR2_X1    g11841(.A1(new_n12033_), .A2(new_n11569_), .Z(new_n12034_));
  AOI21_X1   g11842(.A1(new_n11622_), .A2(new_n11627_), .B(\asqrt[16] ), .ZN(new_n12035_));
  XOR2_X1    g11843(.A1(new_n12035_), .A2(new_n11572_), .Z(new_n12036_));
  AOI21_X1   g11844(.A1(new_n11653_), .A2(new_n11621_), .B(\asqrt[16] ), .ZN(new_n12037_));
  XOR2_X1    g11845(.A1(new_n12037_), .A2(new_n11575_), .Z(new_n12038_));
  INV_X1     g11846(.I(new_n11618_), .ZN(new_n12039_));
  NOR2_X1    g11847(.A1(new_n12039_), .A2(new_n11617_), .ZN(new_n12040_));
  NOR2_X1    g11848(.A1(\asqrt[16] ), .A2(new_n12040_), .ZN(new_n12041_));
  XOR2_X1    g11849(.A1(new_n12041_), .A2(new_n11577_), .Z(new_n12042_));
  INV_X1     g11850(.I(new_n12042_), .ZN(new_n12043_));
  NOR2_X1    g11851(.A1(new_n11649_), .A2(new_n11616_), .ZN(new_n12044_));
  NOR2_X1    g11852(.A1(\asqrt[16] ), .A2(new_n12044_), .ZN(new_n12045_));
  XOR2_X1    g11853(.A1(new_n12045_), .A2(new_n11581_), .Z(new_n12046_));
  INV_X1     g11854(.I(new_n12046_), .ZN(new_n12047_));
  AOI21_X1   g11855(.A1(new_n11610_), .A2(new_n11615_), .B(\asqrt[16] ), .ZN(new_n12048_));
  XOR2_X1    g11856(.A1(new_n12048_), .A2(new_n11584_), .Z(new_n12049_));
  AOI21_X1   g11857(.A1(new_n11645_), .A2(new_n11609_), .B(\asqrt[16] ), .ZN(new_n12050_));
  XOR2_X1    g11858(.A1(new_n12050_), .A2(new_n11587_), .Z(new_n12051_));
  XOR2_X1    g11859(.A1(new_n11643_), .A2(\asqrt[51] ), .Z(new_n12052_));
  NOR2_X1    g11860(.A1(\asqrt[16] ), .A2(new_n12052_), .ZN(new_n12053_));
  XOR2_X1    g11861(.A1(new_n12053_), .A2(new_n11589_), .Z(new_n12054_));
  INV_X1     g11862(.I(new_n12054_), .ZN(new_n12055_));
  NOR2_X1    g11863(.A1(new_n11641_), .A2(new_n11604_), .ZN(new_n12056_));
  NOR2_X1    g11864(.A1(\asqrt[16] ), .A2(new_n12056_), .ZN(new_n12057_));
  XOR2_X1    g11865(.A1(new_n12057_), .A2(new_n11593_), .Z(new_n12058_));
  INV_X1     g11866(.I(new_n12058_), .ZN(new_n12059_));
  AOI21_X1   g11867(.A1(new_n11598_), .A2(new_n11603_), .B(\asqrt[16] ), .ZN(new_n12060_));
  XOR2_X1    g11868(.A1(new_n12060_), .A2(new_n11596_), .Z(new_n12061_));
  OAI21_X1   g11869(.A1(new_n12020_), .A2(\asqrt[49] ), .B(new_n11698_), .ZN(new_n12062_));
  NAND3_X1   g11870(.A1(new_n12062_), .A2(new_n12021_), .A3(new_n1463_), .ZN(new_n12063_));
  AOI21_X1   g11871(.A1(new_n12062_), .A2(new_n12021_), .B(new_n1463_), .ZN(new_n12064_));
  AOI21_X1   g11872(.A1(new_n12061_), .A2(new_n12063_), .B(new_n12064_), .ZN(new_n12065_));
  AOI21_X1   g11873(.A1(new_n12065_), .A2(new_n1305_), .B(new_n12059_), .ZN(new_n12066_));
  NAND2_X1   g11874(.A1(new_n12063_), .A2(new_n12061_), .ZN(new_n12067_));
  INV_X1     g11875(.I(new_n11698_), .ZN(new_n12068_));
  AOI21_X1   g11876(.A1(new_n12003_), .A2(new_n1632_), .B(new_n12068_), .ZN(new_n12069_));
  NAND2_X1   g11877(.A1(new_n12001_), .A2(new_n11701_), .ZN(new_n12070_));
  AOI21_X1   g11878(.A1(new_n12070_), .A2(new_n12019_), .B(new_n1632_), .ZN(new_n12071_));
  OAI21_X1   g11879(.A1(new_n12069_), .A2(new_n12071_), .B(\asqrt[50] ), .ZN(new_n12072_));
  AOI21_X1   g11880(.A1(new_n12067_), .A2(new_n12072_), .B(new_n1305_), .ZN(new_n12073_));
  NOR3_X1    g11881(.A1(new_n12066_), .A2(\asqrt[52] ), .A3(new_n12073_), .ZN(new_n12074_));
  OAI21_X1   g11882(.A1(new_n12066_), .A2(new_n12073_), .B(\asqrt[52] ), .ZN(new_n12075_));
  OAI21_X1   g11883(.A1(new_n12055_), .A2(new_n12074_), .B(new_n12075_), .ZN(new_n12076_));
  OAI21_X1   g11884(.A1(new_n12076_), .A2(\asqrt[53] ), .B(new_n12051_), .ZN(new_n12077_));
  NAND2_X1   g11885(.A1(new_n12076_), .A2(\asqrt[53] ), .ZN(new_n12078_));
  NAND3_X1   g11886(.A1(new_n12077_), .A2(new_n12078_), .A3(new_n860_), .ZN(new_n12079_));
  AOI21_X1   g11887(.A1(new_n12077_), .A2(new_n12078_), .B(new_n860_), .ZN(new_n12080_));
  AOI21_X1   g11888(.A1(new_n12049_), .A2(new_n12079_), .B(new_n12080_), .ZN(new_n12081_));
  AOI21_X1   g11889(.A1(new_n12081_), .A2(new_n744_), .B(new_n12047_), .ZN(new_n12082_));
  NAND2_X1   g11890(.A1(new_n12079_), .A2(new_n12049_), .ZN(new_n12083_));
  INV_X1     g11891(.I(new_n12051_), .ZN(new_n12084_));
  INV_X1     g11892(.I(new_n12061_), .ZN(new_n12085_));
  NOR3_X1    g11893(.A1(new_n12069_), .A2(\asqrt[50] ), .A3(new_n12071_), .ZN(new_n12086_));
  OAI21_X1   g11894(.A1(new_n12085_), .A2(new_n12086_), .B(new_n12072_), .ZN(new_n12087_));
  OAI21_X1   g11895(.A1(new_n12087_), .A2(\asqrt[51] ), .B(new_n12058_), .ZN(new_n12088_));
  NAND2_X1   g11896(.A1(new_n12087_), .A2(\asqrt[51] ), .ZN(new_n12089_));
  NAND3_X1   g11897(.A1(new_n12088_), .A2(new_n12089_), .A3(new_n1150_), .ZN(new_n12090_));
  AOI21_X1   g11898(.A1(new_n12088_), .A2(new_n12089_), .B(new_n1150_), .ZN(new_n12091_));
  AOI21_X1   g11899(.A1(new_n12054_), .A2(new_n12090_), .B(new_n12091_), .ZN(new_n12092_));
  AOI21_X1   g11900(.A1(new_n12092_), .A2(new_n1006_), .B(new_n12084_), .ZN(new_n12093_));
  NAND2_X1   g11901(.A1(new_n12090_), .A2(new_n12054_), .ZN(new_n12094_));
  AOI21_X1   g11902(.A1(new_n12094_), .A2(new_n12075_), .B(new_n1006_), .ZN(new_n12095_));
  OAI21_X1   g11903(.A1(new_n12093_), .A2(new_n12095_), .B(\asqrt[54] ), .ZN(new_n12096_));
  AOI21_X1   g11904(.A1(new_n12083_), .A2(new_n12096_), .B(new_n744_), .ZN(new_n12097_));
  NOR3_X1    g11905(.A1(new_n12082_), .A2(\asqrt[56] ), .A3(new_n12097_), .ZN(new_n12098_));
  OAI21_X1   g11906(.A1(new_n12082_), .A2(new_n12097_), .B(\asqrt[56] ), .ZN(new_n12099_));
  OAI21_X1   g11907(.A1(new_n12043_), .A2(new_n12098_), .B(new_n12099_), .ZN(new_n12100_));
  OAI21_X1   g11908(.A1(new_n12100_), .A2(\asqrt[57] ), .B(new_n12038_), .ZN(new_n12101_));
  NOR2_X1    g11909(.A1(new_n12098_), .A2(new_n12043_), .ZN(new_n12102_));
  INV_X1     g11910(.I(new_n12049_), .ZN(new_n12103_));
  NOR3_X1    g11911(.A1(new_n12093_), .A2(\asqrt[54] ), .A3(new_n12095_), .ZN(new_n12104_));
  OAI21_X1   g11912(.A1(new_n12103_), .A2(new_n12104_), .B(new_n12096_), .ZN(new_n12105_));
  OAI21_X1   g11913(.A1(new_n12105_), .A2(\asqrt[55] ), .B(new_n12046_), .ZN(new_n12106_));
  NAND2_X1   g11914(.A1(new_n12105_), .A2(\asqrt[55] ), .ZN(new_n12107_));
  AOI21_X1   g11915(.A1(new_n12106_), .A2(new_n12107_), .B(new_n634_), .ZN(new_n12108_));
  OAI21_X1   g11916(.A1(new_n12102_), .A2(new_n12108_), .B(\asqrt[57] ), .ZN(new_n12109_));
  NAND3_X1   g11917(.A1(new_n12101_), .A2(new_n423_), .A3(new_n12109_), .ZN(new_n12110_));
  NAND2_X1   g11918(.A1(new_n12110_), .A2(new_n12036_), .ZN(new_n12111_));
  INV_X1     g11919(.I(new_n12038_), .ZN(new_n12112_));
  NAND3_X1   g11920(.A1(new_n12106_), .A2(new_n12107_), .A3(new_n634_), .ZN(new_n12113_));
  AOI21_X1   g11921(.A1(new_n12042_), .A2(new_n12113_), .B(new_n12108_), .ZN(new_n12114_));
  AOI21_X1   g11922(.A1(new_n12114_), .A2(new_n531_), .B(new_n12112_), .ZN(new_n12115_));
  NAND2_X1   g11923(.A1(new_n12113_), .A2(new_n12042_), .ZN(new_n12116_));
  AOI21_X1   g11924(.A1(new_n12116_), .A2(new_n12099_), .B(new_n531_), .ZN(new_n12117_));
  OAI21_X1   g11925(.A1(new_n12115_), .A2(new_n12117_), .B(\asqrt[58] ), .ZN(new_n12118_));
  NAND3_X1   g11926(.A1(new_n12111_), .A2(new_n337_), .A3(new_n12118_), .ZN(new_n12119_));
  AOI21_X1   g11927(.A1(new_n12111_), .A2(new_n12118_), .B(new_n337_), .ZN(new_n12120_));
  AOI21_X1   g11928(.A1(new_n12034_), .A2(new_n12119_), .B(new_n12120_), .ZN(new_n12121_));
  AOI21_X1   g11929(.A1(new_n12121_), .A2(new_n266_), .B(new_n12031_), .ZN(new_n12122_));
  INV_X1     g11930(.I(new_n12036_), .ZN(new_n12123_));
  NOR3_X1    g11931(.A1(new_n12115_), .A2(\asqrt[58] ), .A3(new_n12117_), .ZN(new_n12124_));
  OAI21_X1   g11932(.A1(new_n12123_), .A2(new_n12124_), .B(new_n12118_), .ZN(new_n12125_));
  OAI21_X1   g11933(.A1(new_n12125_), .A2(\asqrt[59] ), .B(new_n12034_), .ZN(new_n12126_));
  NAND2_X1   g11934(.A1(new_n12125_), .A2(\asqrt[59] ), .ZN(new_n12127_));
  AOI21_X1   g11935(.A1(new_n12126_), .A2(new_n12127_), .B(new_n266_), .ZN(new_n12128_));
  OAI21_X1   g11936(.A1(new_n12122_), .A2(new_n12128_), .B(\asqrt[61] ), .ZN(new_n12129_));
  AOI21_X1   g11937(.A1(new_n11672_), .A2(new_n11667_), .B(\asqrt[16] ), .ZN(new_n12130_));
  XOR2_X1    g11938(.A1(new_n12130_), .A2(new_n11562_), .Z(new_n12131_));
  INV_X1     g11939(.I(new_n12131_), .ZN(new_n12132_));
  NOR3_X1    g11940(.A1(new_n12122_), .A2(\asqrt[61] ), .A3(new_n12128_), .ZN(new_n12133_));
  OAI21_X1   g11941(.A1(new_n12132_), .A2(new_n12133_), .B(new_n12129_), .ZN(new_n12134_));
  NAND3_X1   g11942(.A1(new_n12126_), .A2(new_n12127_), .A3(new_n266_), .ZN(new_n12135_));
  NAND2_X1   g11943(.A1(new_n12135_), .A2(new_n12030_), .ZN(new_n12136_));
  INV_X1     g11944(.I(new_n12034_), .ZN(new_n12137_));
  AOI21_X1   g11945(.A1(new_n12101_), .A2(new_n12109_), .B(new_n423_), .ZN(new_n12138_));
  AOI21_X1   g11946(.A1(new_n12036_), .A2(new_n12110_), .B(new_n12138_), .ZN(new_n12139_));
  AOI21_X1   g11947(.A1(new_n12139_), .A2(new_n337_), .B(new_n12137_), .ZN(new_n12140_));
  OAI21_X1   g11948(.A1(new_n12140_), .A2(new_n12120_), .B(\asqrt[60] ), .ZN(new_n12141_));
  AOI21_X1   g11949(.A1(new_n12136_), .A2(new_n12141_), .B(new_n239_), .ZN(new_n12142_));
  AOI21_X1   g11950(.A1(new_n12030_), .A2(new_n12135_), .B(new_n12128_), .ZN(new_n12143_));
  AOI21_X1   g11951(.A1(new_n12143_), .A2(new_n239_), .B(new_n12132_), .ZN(new_n12144_));
  OAI21_X1   g11952(.A1(new_n12144_), .A2(new_n12142_), .B(new_n201_), .ZN(new_n12145_));
  NOR3_X1    g11953(.A1(new_n12140_), .A2(\asqrt[60] ), .A3(new_n12120_), .ZN(new_n12146_));
  OAI21_X1   g11954(.A1(new_n12031_), .A2(new_n12146_), .B(new_n12141_), .ZN(new_n12147_));
  OAI21_X1   g11955(.A1(new_n12147_), .A2(\asqrt[61] ), .B(new_n12131_), .ZN(new_n12148_));
  NAND3_X1   g11956(.A1(new_n12148_), .A2(\asqrt[62] ), .A3(new_n12129_), .ZN(new_n12149_));
  AOI21_X1   g11957(.A1(new_n11662_), .A2(new_n11668_), .B(\asqrt[16] ), .ZN(new_n12150_));
  XOR2_X1    g11958(.A1(new_n12150_), .A2(new_n11664_), .Z(new_n12151_));
  INV_X1     g11959(.I(new_n12151_), .ZN(new_n12152_));
  AOI22_X1   g11960(.A1(new_n12149_), .A2(new_n12145_), .B1(new_n12134_), .B2(new_n12152_), .ZN(new_n12153_));
  NOR2_X1    g11961(.A1(new_n11681_), .A2(new_n11559_), .ZN(new_n12154_));
  OAI21_X1   g11962(.A1(\asqrt[16] ), .A2(new_n12154_), .B(new_n11688_), .ZN(new_n12155_));
  INV_X1     g11963(.I(new_n12155_), .ZN(new_n12156_));
  OAI21_X1   g11964(.A1(new_n12153_), .A2(new_n12027_), .B(new_n12156_), .ZN(new_n12157_));
  OAI21_X1   g11965(.A1(new_n12134_), .A2(\asqrt[62] ), .B(new_n12151_), .ZN(new_n12158_));
  NAND2_X1   g11966(.A1(new_n12134_), .A2(\asqrt[62] ), .ZN(new_n12159_));
  NAND3_X1   g11967(.A1(new_n12158_), .A2(new_n12159_), .A3(new_n12027_), .ZN(new_n12160_));
  NAND2_X1   g11968(.A1(new_n11802_), .A2(new_n11558_), .ZN(new_n12161_));
  XOR2_X1    g11969(.A1(new_n11681_), .A2(new_n11559_), .Z(new_n12162_));
  NAND3_X1   g11970(.A1(new_n12161_), .A2(\asqrt[63] ), .A3(new_n12162_), .ZN(new_n12163_));
  INV_X1     g11971(.I(new_n11791_), .ZN(new_n12164_));
  NAND4_X1   g11972(.A1(new_n12164_), .A2(new_n11559_), .A3(new_n11688_), .A4(new_n11695_), .ZN(new_n12165_));
  NAND2_X1   g11973(.A1(new_n12163_), .A2(new_n12165_), .ZN(new_n12166_));
  INV_X1     g11974(.I(new_n12166_), .ZN(new_n12167_));
  NAND4_X1   g11975(.A1(new_n12157_), .A2(new_n193_), .A3(new_n12160_), .A4(new_n12167_), .ZN(\asqrt[15] ));
  AOI21_X1   g11976(.A1(new_n12004_), .A2(new_n12021_), .B(\asqrt[15] ), .ZN(new_n12169_));
  XOR2_X1    g11977(.A1(new_n12169_), .A2(new_n11698_), .Z(new_n12170_));
  AOI21_X1   g11978(.A1(new_n12001_), .A2(new_n12019_), .B(\asqrt[15] ), .ZN(new_n12171_));
  XOR2_X1    g11979(.A1(new_n12171_), .A2(new_n11701_), .Z(new_n12172_));
  NAND2_X1   g11980(.A1(new_n12014_), .A2(new_n1953_), .ZN(new_n12173_));
  AOI21_X1   g11981(.A1(new_n12173_), .A2(new_n12000_), .B(\asqrt[15] ), .ZN(new_n12174_));
  XOR2_X1    g11982(.A1(new_n12174_), .A2(new_n11704_), .Z(new_n12175_));
  INV_X1     g11983(.I(new_n12175_), .ZN(new_n12176_));
  AOI21_X1   g11984(.A1(new_n12012_), .A2(new_n11997_), .B(\asqrt[15] ), .ZN(new_n12177_));
  XOR2_X1    g11985(.A1(new_n12177_), .A2(new_n11706_), .Z(new_n12178_));
  INV_X1     g11986(.I(new_n12178_), .ZN(new_n12179_));
  NAND2_X1   g11987(.A1(new_n11979_), .A2(new_n2332_), .ZN(new_n12180_));
  AOI21_X1   g11988(.A1(new_n12180_), .A2(new_n12011_), .B(\asqrt[15] ), .ZN(new_n12181_));
  XOR2_X1    g11989(.A1(new_n12181_), .A2(new_n11709_), .Z(new_n12182_));
  AOI21_X1   g11990(.A1(new_n11977_), .A2(new_n11994_), .B(\asqrt[15] ), .ZN(new_n12183_));
  XOR2_X1    g11991(.A1(new_n12183_), .A2(new_n11713_), .Z(new_n12184_));
  NAND2_X1   g11992(.A1(new_n11990_), .A2(new_n2749_), .ZN(new_n12185_));
  AOI21_X1   g11993(.A1(new_n12185_), .A2(new_n11976_), .B(\asqrt[15] ), .ZN(new_n12186_));
  XOR2_X1    g11994(.A1(new_n12186_), .A2(new_n11716_), .Z(new_n12187_));
  INV_X1     g11995(.I(new_n12187_), .ZN(new_n12188_));
  AOI21_X1   g11996(.A1(new_n11988_), .A2(new_n11973_), .B(\asqrt[15] ), .ZN(new_n12189_));
  XOR2_X1    g11997(.A1(new_n12189_), .A2(new_n11718_), .Z(new_n12190_));
  INV_X1     g11998(.I(new_n12190_), .ZN(new_n12191_));
  NAND2_X1   g11999(.A1(new_n11955_), .A2(new_n3195_), .ZN(new_n12192_));
  AOI21_X1   g12000(.A1(new_n12192_), .A2(new_n11987_), .B(\asqrt[15] ), .ZN(new_n12193_));
  XOR2_X1    g12001(.A1(new_n12193_), .A2(new_n11721_), .Z(new_n12194_));
  AOI21_X1   g12002(.A1(new_n11953_), .A2(new_n11970_), .B(\asqrt[15] ), .ZN(new_n12195_));
  XOR2_X1    g12003(.A1(new_n12195_), .A2(new_n11725_), .Z(new_n12196_));
  NAND2_X1   g12004(.A1(new_n11966_), .A2(new_n3681_), .ZN(new_n12197_));
  AOI21_X1   g12005(.A1(new_n12197_), .A2(new_n11952_), .B(\asqrt[15] ), .ZN(new_n12198_));
  XOR2_X1    g12006(.A1(new_n12198_), .A2(new_n11728_), .Z(new_n12199_));
  INV_X1     g12007(.I(new_n12199_), .ZN(new_n12200_));
  AOI21_X1   g12008(.A1(new_n11964_), .A2(new_n11949_), .B(\asqrt[15] ), .ZN(new_n12201_));
  XOR2_X1    g12009(.A1(new_n12201_), .A2(new_n11730_), .Z(new_n12202_));
  INV_X1     g12010(.I(new_n12202_), .ZN(new_n12203_));
  NAND2_X1   g12011(.A1(new_n11931_), .A2(new_n4196_), .ZN(new_n12204_));
  AOI21_X1   g12012(.A1(new_n12204_), .A2(new_n11963_), .B(\asqrt[15] ), .ZN(new_n12205_));
  XOR2_X1    g12013(.A1(new_n12205_), .A2(new_n11733_), .Z(new_n12206_));
  AOI21_X1   g12014(.A1(new_n11929_), .A2(new_n11946_), .B(\asqrt[15] ), .ZN(new_n12207_));
  XOR2_X1    g12015(.A1(new_n12207_), .A2(new_n11737_), .Z(new_n12208_));
  NAND2_X1   g12016(.A1(new_n11942_), .A2(new_n4751_), .ZN(new_n12209_));
  AOI21_X1   g12017(.A1(new_n12209_), .A2(new_n11928_), .B(\asqrt[15] ), .ZN(new_n12210_));
  XOR2_X1    g12018(.A1(new_n12210_), .A2(new_n11740_), .Z(new_n12211_));
  INV_X1     g12019(.I(new_n12211_), .ZN(new_n12212_));
  AOI21_X1   g12020(.A1(new_n11940_), .A2(new_n11925_), .B(\asqrt[15] ), .ZN(new_n12213_));
  XOR2_X1    g12021(.A1(new_n12213_), .A2(new_n11742_), .Z(new_n12214_));
  INV_X1     g12022(.I(new_n12214_), .ZN(new_n12215_));
  NAND2_X1   g12023(.A1(new_n11907_), .A2(new_n5336_), .ZN(new_n12216_));
  AOI21_X1   g12024(.A1(new_n12216_), .A2(new_n11939_), .B(\asqrt[15] ), .ZN(new_n12217_));
  XOR2_X1    g12025(.A1(new_n12217_), .A2(new_n11745_), .Z(new_n12218_));
  AOI21_X1   g12026(.A1(new_n11905_), .A2(new_n11922_), .B(\asqrt[15] ), .ZN(new_n12219_));
  XOR2_X1    g12027(.A1(new_n12219_), .A2(new_n11749_), .Z(new_n12220_));
  NAND2_X1   g12028(.A1(new_n11918_), .A2(new_n5947_), .ZN(new_n12221_));
  AOI21_X1   g12029(.A1(new_n12221_), .A2(new_n11904_), .B(\asqrt[15] ), .ZN(new_n12222_));
  XOR2_X1    g12030(.A1(new_n12222_), .A2(new_n11752_), .Z(new_n12223_));
  INV_X1     g12031(.I(new_n12223_), .ZN(new_n12224_));
  AOI21_X1   g12032(.A1(new_n11916_), .A2(new_n11901_), .B(\asqrt[15] ), .ZN(new_n12225_));
  XOR2_X1    g12033(.A1(new_n12225_), .A2(new_n11754_), .Z(new_n12226_));
  INV_X1     g12034(.I(new_n12226_), .ZN(new_n12227_));
  NAND2_X1   g12035(.A1(new_n11883_), .A2(new_n6636_), .ZN(new_n12228_));
  AOI21_X1   g12036(.A1(new_n12228_), .A2(new_n11915_), .B(\asqrt[15] ), .ZN(new_n12229_));
  XOR2_X1    g12037(.A1(new_n12229_), .A2(new_n11757_), .Z(new_n12230_));
  AOI21_X1   g12038(.A1(new_n11881_), .A2(new_n11898_), .B(\asqrt[15] ), .ZN(new_n12231_));
  XOR2_X1    g12039(.A1(new_n12231_), .A2(new_n11761_), .Z(new_n12232_));
  NAND2_X1   g12040(.A1(new_n11894_), .A2(new_n7331_), .ZN(new_n12233_));
  AOI21_X1   g12041(.A1(new_n12233_), .A2(new_n11880_), .B(\asqrt[15] ), .ZN(new_n12234_));
  XOR2_X1    g12042(.A1(new_n12234_), .A2(new_n11764_), .Z(new_n12235_));
  INV_X1     g12043(.I(new_n12235_), .ZN(new_n12236_));
  AOI21_X1   g12044(.A1(new_n11892_), .A2(new_n11877_), .B(\asqrt[15] ), .ZN(new_n12237_));
  XOR2_X1    g12045(.A1(new_n12237_), .A2(new_n11766_), .Z(new_n12238_));
  INV_X1     g12046(.I(new_n12238_), .ZN(new_n12239_));
  NAND2_X1   g12047(.A1(new_n11859_), .A2(new_n8077_), .ZN(new_n12240_));
  AOI21_X1   g12048(.A1(new_n12240_), .A2(new_n11891_), .B(\asqrt[15] ), .ZN(new_n12241_));
  XOR2_X1    g12049(.A1(new_n12241_), .A2(new_n11769_), .Z(new_n12242_));
  AOI21_X1   g12050(.A1(new_n11857_), .A2(new_n11874_), .B(\asqrt[15] ), .ZN(new_n12243_));
  XOR2_X1    g12051(.A1(new_n12243_), .A2(new_n11773_), .Z(new_n12244_));
  NAND2_X1   g12052(.A1(new_n11870_), .A2(new_n8849_), .ZN(new_n12245_));
  AOI21_X1   g12053(.A1(new_n12245_), .A2(new_n11856_), .B(\asqrt[15] ), .ZN(new_n12246_));
  XOR2_X1    g12054(.A1(new_n12246_), .A2(new_n11776_), .Z(new_n12247_));
  INV_X1     g12055(.I(new_n12247_), .ZN(new_n12248_));
  AOI21_X1   g12056(.A1(new_n11868_), .A2(new_n11853_), .B(\asqrt[15] ), .ZN(new_n12249_));
  XOR2_X1    g12057(.A1(new_n12249_), .A2(new_n11778_), .Z(new_n12250_));
  INV_X1     g12058(.I(new_n12250_), .ZN(new_n12251_));
  NAND2_X1   g12059(.A1(new_n11831_), .A2(new_n9656_), .ZN(new_n12252_));
  AOI21_X1   g12060(.A1(new_n12252_), .A2(new_n11867_), .B(\asqrt[15] ), .ZN(new_n12253_));
  XOR2_X1    g12061(.A1(new_n12253_), .A2(new_n11781_), .Z(new_n12254_));
  AOI21_X1   g12062(.A1(new_n11829_), .A2(new_n11850_), .B(\asqrt[15] ), .ZN(new_n12255_));
  XOR2_X1    g12063(.A1(new_n12255_), .A2(new_n11784_), .Z(new_n12256_));
  NAND2_X1   g12064(.A1(new_n11846_), .A2(new_n10497_), .ZN(new_n12257_));
  AOI21_X1   g12065(.A1(new_n12257_), .A2(new_n11828_), .B(\asqrt[15] ), .ZN(new_n12258_));
  XOR2_X1    g12066(.A1(new_n12258_), .A2(new_n11790_), .Z(new_n12259_));
  INV_X1     g12067(.I(new_n12259_), .ZN(new_n12260_));
  AOI21_X1   g12068(.A1(new_n11844_), .A2(new_n11825_), .B(\asqrt[15] ), .ZN(new_n12261_));
  XOR2_X1    g12069(.A1(new_n12261_), .A2(new_n11835_), .Z(new_n12262_));
  INV_X1     g12070(.I(new_n12262_), .ZN(new_n12263_));
  NAND2_X1   g12071(.A1(\asqrt[16] ), .A2(new_n11813_), .ZN(new_n12264_));
  NOR2_X1    g12072(.A1(new_n11820_), .A2(\a[32] ), .ZN(new_n12265_));
  AOI22_X1   g12073(.A1(new_n12264_), .A2(new_n11820_), .B1(\asqrt[16] ), .B2(new_n12265_), .ZN(new_n12266_));
  OAI21_X1   g12074(.A1(new_n11802_), .A2(new_n11813_), .B(new_n11839_), .ZN(new_n12267_));
  AOI21_X1   g12075(.A1(new_n11838_), .A2(new_n12267_), .B(\asqrt[15] ), .ZN(new_n12268_));
  XOR2_X1    g12076(.A1(new_n12268_), .A2(new_n12266_), .Z(new_n12269_));
  NOR2_X1    g12077(.A1(new_n12144_), .A2(new_n12142_), .ZN(new_n12270_));
  AOI21_X1   g12078(.A1(new_n12148_), .A2(new_n12129_), .B(\asqrt[62] ), .ZN(new_n12271_));
  NOR3_X1    g12079(.A1(new_n12144_), .A2(new_n201_), .A3(new_n12142_), .ZN(new_n12272_));
  OAI22_X1   g12080(.A1(new_n12271_), .A2(new_n12272_), .B1(new_n12270_), .B2(new_n12151_), .ZN(new_n12273_));
  AOI21_X1   g12081(.A1(new_n12273_), .A2(new_n12026_), .B(new_n12155_), .ZN(new_n12274_));
  AOI21_X1   g12082(.A1(new_n12270_), .A2(new_n201_), .B(new_n12152_), .ZN(new_n12275_));
  NOR2_X1    g12083(.A1(new_n12270_), .A2(new_n201_), .ZN(new_n12276_));
  NOR3_X1    g12084(.A1(new_n12275_), .A2(new_n12276_), .A3(new_n12026_), .ZN(new_n12277_));
  NAND3_X1   g12085(.A1(new_n12163_), .A2(\asqrt[16] ), .A3(new_n12165_), .ZN(new_n12278_));
  NOR4_X1    g12086(.A1(new_n12274_), .A2(\asqrt[63] ), .A3(new_n12277_), .A4(new_n12278_), .ZN(new_n12279_));
  INV_X1     g12087(.I(new_n12279_), .ZN(new_n12280_));
  NAND2_X1   g12088(.A1(\asqrt[15] ), .A2(new_n11810_), .ZN(new_n12281_));
  AOI21_X1   g12089(.A1(new_n12281_), .A2(new_n12280_), .B(\a[32] ), .ZN(new_n12282_));
  NOR4_X1    g12090(.A1(new_n12274_), .A2(\asqrt[63] ), .A3(new_n12277_), .A4(new_n12166_), .ZN(new_n12283_));
  NOR2_X1    g12091(.A1(new_n12283_), .A2(new_n11811_), .ZN(new_n12284_));
  NOR3_X1    g12092(.A1(new_n12284_), .A2(new_n11813_), .A3(new_n12279_), .ZN(new_n12285_));
  NOR2_X1    g12093(.A1(new_n12285_), .A2(new_n12282_), .ZN(new_n12286_));
  INV_X1     g12094(.I(\a[30] ), .ZN(new_n12287_));
  NOR2_X1    g12095(.A1(\a[28] ), .A2(\a[29] ), .ZN(new_n12288_));
  NOR3_X1    g12096(.A1(new_n12283_), .A2(new_n12287_), .A3(new_n12288_), .ZN(new_n12289_));
  INV_X1     g12097(.I(new_n12288_), .ZN(new_n12290_));
  AOI21_X1   g12098(.A1(new_n12283_), .A2(\a[30] ), .B(new_n12290_), .ZN(new_n12291_));
  OAI21_X1   g12099(.A1(new_n12289_), .A2(new_n12291_), .B(\asqrt[16] ), .ZN(new_n12292_));
  NAND2_X1   g12100(.A1(new_n12288_), .A2(new_n12287_), .ZN(new_n12293_));
  NAND3_X1   g12101(.A1(new_n11691_), .A2(new_n11693_), .A3(new_n12293_), .ZN(new_n12294_));
  NAND2_X1   g12102(.A1(new_n11805_), .A2(new_n12294_), .ZN(new_n12295_));
  NAND3_X1   g12103(.A1(\asqrt[15] ), .A2(\a[30] ), .A3(new_n12295_), .ZN(new_n12296_));
  NOR3_X1    g12104(.A1(new_n12283_), .A2(\a[30] ), .A3(\a[31] ), .ZN(new_n12297_));
  INV_X1     g12105(.I(\a[31] ), .ZN(new_n12298_));
  AOI21_X1   g12106(.A1(\asqrt[15] ), .A2(new_n12287_), .B(new_n12298_), .ZN(new_n12299_));
  NOR2_X1    g12107(.A1(new_n12297_), .A2(new_n12299_), .ZN(new_n12300_));
  NAND4_X1   g12108(.A1(new_n12292_), .A2(new_n12300_), .A3(new_n11373_), .A4(new_n12296_), .ZN(new_n12301_));
  NAND2_X1   g12109(.A1(new_n12301_), .A2(new_n12286_), .ZN(new_n12302_));
  NAND3_X1   g12110(.A1(\asqrt[15] ), .A2(\a[30] ), .A3(new_n12290_), .ZN(new_n12303_));
  OAI21_X1   g12111(.A1(\asqrt[15] ), .A2(new_n12287_), .B(new_n12288_), .ZN(new_n12304_));
  AOI21_X1   g12112(.A1(new_n12304_), .A2(new_n12303_), .B(new_n11802_), .ZN(new_n12305_));
  NAND3_X1   g12113(.A1(\asqrt[15] ), .A2(new_n12287_), .A3(new_n12298_), .ZN(new_n12306_));
  OAI21_X1   g12114(.A1(new_n12283_), .A2(\a[30] ), .B(\a[31] ), .ZN(new_n12307_));
  NAND3_X1   g12115(.A1(new_n12296_), .A2(new_n12307_), .A3(new_n12306_), .ZN(new_n12308_));
  OAI21_X1   g12116(.A1(new_n12308_), .A2(new_n12305_), .B(\asqrt[17] ), .ZN(new_n12309_));
  NAND3_X1   g12117(.A1(new_n12302_), .A2(new_n10914_), .A3(new_n12309_), .ZN(new_n12310_));
  AOI21_X1   g12118(.A1(new_n12302_), .A2(new_n12309_), .B(new_n10914_), .ZN(new_n12311_));
  AOI21_X1   g12119(.A1(new_n12269_), .A2(new_n12310_), .B(new_n12311_), .ZN(new_n12312_));
  AOI21_X1   g12120(.A1(new_n12312_), .A2(new_n10497_), .B(new_n12263_), .ZN(new_n12313_));
  OR2_X2     g12121(.A1(new_n12285_), .A2(new_n12282_), .Z(new_n12314_));
  NOR3_X1    g12122(.A1(new_n12308_), .A2(new_n12305_), .A3(\asqrt[17] ), .ZN(new_n12315_));
  OAI21_X1   g12123(.A1(new_n12314_), .A2(new_n12315_), .B(new_n12309_), .ZN(new_n12316_));
  OAI21_X1   g12124(.A1(new_n12316_), .A2(\asqrt[18] ), .B(new_n12269_), .ZN(new_n12317_));
  NAND2_X1   g12125(.A1(new_n12316_), .A2(\asqrt[18] ), .ZN(new_n12318_));
  AOI21_X1   g12126(.A1(new_n12317_), .A2(new_n12318_), .B(new_n10497_), .ZN(new_n12319_));
  NOR3_X1    g12127(.A1(new_n12313_), .A2(\asqrt[20] ), .A3(new_n12319_), .ZN(new_n12320_));
  OAI21_X1   g12128(.A1(new_n12313_), .A2(new_n12319_), .B(\asqrt[20] ), .ZN(new_n12321_));
  OAI21_X1   g12129(.A1(new_n12260_), .A2(new_n12320_), .B(new_n12321_), .ZN(new_n12322_));
  OAI21_X1   g12130(.A1(new_n12322_), .A2(\asqrt[21] ), .B(new_n12256_), .ZN(new_n12323_));
  NAND3_X1   g12131(.A1(new_n12317_), .A2(new_n12318_), .A3(new_n10497_), .ZN(new_n12324_));
  AOI21_X1   g12132(.A1(new_n12262_), .A2(new_n12324_), .B(new_n12319_), .ZN(new_n12325_));
  AOI21_X1   g12133(.A1(new_n12325_), .A2(new_n10052_), .B(new_n12260_), .ZN(new_n12326_));
  NAND2_X1   g12134(.A1(new_n12324_), .A2(new_n12262_), .ZN(new_n12327_));
  INV_X1     g12135(.I(new_n12319_), .ZN(new_n12328_));
  AOI21_X1   g12136(.A1(new_n12327_), .A2(new_n12328_), .B(new_n10052_), .ZN(new_n12329_));
  OAI21_X1   g12137(.A1(new_n12326_), .A2(new_n12329_), .B(\asqrt[21] ), .ZN(new_n12330_));
  NAND3_X1   g12138(.A1(new_n12323_), .A2(new_n9233_), .A3(new_n12330_), .ZN(new_n12331_));
  AOI21_X1   g12139(.A1(new_n12323_), .A2(new_n12330_), .B(new_n9233_), .ZN(new_n12332_));
  AOI21_X1   g12140(.A1(new_n12254_), .A2(new_n12331_), .B(new_n12332_), .ZN(new_n12333_));
  AOI21_X1   g12141(.A1(new_n12333_), .A2(new_n8849_), .B(new_n12251_), .ZN(new_n12334_));
  INV_X1     g12142(.I(new_n12256_), .ZN(new_n12335_));
  NOR3_X1    g12143(.A1(new_n12326_), .A2(\asqrt[21] ), .A3(new_n12329_), .ZN(new_n12336_));
  OAI21_X1   g12144(.A1(new_n12335_), .A2(new_n12336_), .B(new_n12330_), .ZN(new_n12337_));
  OAI21_X1   g12145(.A1(new_n12337_), .A2(\asqrt[22] ), .B(new_n12254_), .ZN(new_n12338_));
  NAND2_X1   g12146(.A1(new_n12337_), .A2(\asqrt[22] ), .ZN(new_n12339_));
  AOI21_X1   g12147(.A1(new_n12338_), .A2(new_n12339_), .B(new_n8849_), .ZN(new_n12340_));
  NOR3_X1    g12148(.A1(new_n12334_), .A2(\asqrt[24] ), .A3(new_n12340_), .ZN(new_n12341_));
  OAI21_X1   g12149(.A1(new_n12334_), .A2(new_n12340_), .B(\asqrt[24] ), .ZN(new_n12342_));
  OAI21_X1   g12150(.A1(new_n12248_), .A2(new_n12341_), .B(new_n12342_), .ZN(new_n12343_));
  OAI21_X1   g12151(.A1(new_n12343_), .A2(\asqrt[25] ), .B(new_n12244_), .ZN(new_n12344_));
  NAND3_X1   g12152(.A1(new_n12338_), .A2(new_n12339_), .A3(new_n8849_), .ZN(new_n12345_));
  AOI21_X1   g12153(.A1(new_n12250_), .A2(new_n12345_), .B(new_n12340_), .ZN(new_n12346_));
  AOI21_X1   g12154(.A1(new_n12346_), .A2(new_n8440_), .B(new_n12248_), .ZN(new_n12347_));
  NAND2_X1   g12155(.A1(new_n12345_), .A2(new_n12250_), .ZN(new_n12348_));
  INV_X1     g12156(.I(new_n12340_), .ZN(new_n12349_));
  AOI21_X1   g12157(.A1(new_n12348_), .A2(new_n12349_), .B(new_n8440_), .ZN(new_n12350_));
  OAI21_X1   g12158(.A1(new_n12347_), .A2(new_n12350_), .B(\asqrt[25] ), .ZN(new_n12351_));
  NAND3_X1   g12159(.A1(new_n12344_), .A2(new_n7690_), .A3(new_n12351_), .ZN(new_n12352_));
  AOI21_X1   g12160(.A1(new_n12344_), .A2(new_n12351_), .B(new_n7690_), .ZN(new_n12353_));
  AOI21_X1   g12161(.A1(new_n12242_), .A2(new_n12352_), .B(new_n12353_), .ZN(new_n12354_));
  AOI21_X1   g12162(.A1(new_n12354_), .A2(new_n7331_), .B(new_n12239_), .ZN(new_n12355_));
  INV_X1     g12163(.I(new_n12244_), .ZN(new_n12356_));
  NOR3_X1    g12164(.A1(new_n12347_), .A2(\asqrt[25] ), .A3(new_n12350_), .ZN(new_n12357_));
  OAI21_X1   g12165(.A1(new_n12356_), .A2(new_n12357_), .B(new_n12351_), .ZN(new_n12358_));
  OAI21_X1   g12166(.A1(new_n12358_), .A2(\asqrt[26] ), .B(new_n12242_), .ZN(new_n12359_));
  NAND2_X1   g12167(.A1(new_n12358_), .A2(\asqrt[26] ), .ZN(new_n12360_));
  AOI21_X1   g12168(.A1(new_n12359_), .A2(new_n12360_), .B(new_n7331_), .ZN(new_n12361_));
  NOR3_X1    g12169(.A1(new_n12355_), .A2(\asqrt[28] ), .A3(new_n12361_), .ZN(new_n12362_));
  OAI21_X1   g12170(.A1(new_n12355_), .A2(new_n12361_), .B(\asqrt[28] ), .ZN(new_n12363_));
  OAI21_X1   g12171(.A1(new_n12236_), .A2(new_n12362_), .B(new_n12363_), .ZN(new_n12364_));
  OAI21_X1   g12172(.A1(new_n12364_), .A2(\asqrt[29] ), .B(new_n12232_), .ZN(new_n12365_));
  NAND3_X1   g12173(.A1(new_n12359_), .A2(new_n12360_), .A3(new_n7331_), .ZN(new_n12366_));
  AOI21_X1   g12174(.A1(new_n12238_), .A2(new_n12366_), .B(new_n12361_), .ZN(new_n12367_));
  AOI21_X1   g12175(.A1(new_n12367_), .A2(new_n6966_), .B(new_n12236_), .ZN(new_n12368_));
  NAND2_X1   g12176(.A1(new_n12366_), .A2(new_n12238_), .ZN(new_n12369_));
  INV_X1     g12177(.I(new_n12361_), .ZN(new_n12370_));
  AOI21_X1   g12178(.A1(new_n12369_), .A2(new_n12370_), .B(new_n6966_), .ZN(new_n12371_));
  OAI21_X1   g12179(.A1(new_n12368_), .A2(new_n12371_), .B(\asqrt[29] ), .ZN(new_n12372_));
  NAND3_X1   g12180(.A1(new_n12365_), .A2(new_n6275_), .A3(new_n12372_), .ZN(new_n12373_));
  AOI21_X1   g12181(.A1(new_n12365_), .A2(new_n12372_), .B(new_n6275_), .ZN(new_n12374_));
  AOI21_X1   g12182(.A1(new_n12230_), .A2(new_n12373_), .B(new_n12374_), .ZN(new_n12375_));
  AOI21_X1   g12183(.A1(new_n12375_), .A2(new_n5947_), .B(new_n12227_), .ZN(new_n12376_));
  INV_X1     g12184(.I(new_n12232_), .ZN(new_n12377_));
  NOR3_X1    g12185(.A1(new_n12368_), .A2(\asqrt[29] ), .A3(new_n12371_), .ZN(new_n12378_));
  OAI21_X1   g12186(.A1(new_n12377_), .A2(new_n12378_), .B(new_n12372_), .ZN(new_n12379_));
  OAI21_X1   g12187(.A1(new_n12379_), .A2(\asqrt[30] ), .B(new_n12230_), .ZN(new_n12380_));
  NAND2_X1   g12188(.A1(new_n12379_), .A2(\asqrt[30] ), .ZN(new_n12381_));
  AOI21_X1   g12189(.A1(new_n12380_), .A2(new_n12381_), .B(new_n5947_), .ZN(new_n12382_));
  NOR3_X1    g12190(.A1(new_n12376_), .A2(\asqrt[32] ), .A3(new_n12382_), .ZN(new_n12383_));
  OAI21_X1   g12191(.A1(new_n12376_), .A2(new_n12382_), .B(\asqrt[32] ), .ZN(new_n12384_));
  OAI21_X1   g12192(.A1(new_n12224_), .A2(new_n12383_), .B(new_n12384_), .ZN(new_n12385_));
  OAI21_X1   g12193(.A1(new_n12385_), .A2(\asqrt[33] ), .B(new_n12220_), .ZN(new_n12386_));
  NAND3_X1   g12194(.A1(new_n12380_), .A2(new_n12381_), .A3(new_n5947_), .ZN(new_n12387_));
  AOI21_X1   g12195(.A1(new_n12226_), .A2(new_n12387_), .B(new_n12382_), .ZN(new_n12388_));
  AOI21_X1   g12196(.A1(new_n12388_), .A2(new_n5643_), .B(new_n12224_), .ZN(new_n12389_));
  NAND2_X1   g12197(.A1(new_n12387_), .A2(new_n12226_), .ZN(new_n12390_));
  INV_X1     g12198(.I(new_n12382_), .ZN(new_n12391_));
  AOI21_X1   g12199(.A1(new_n12390_), .A2(new_n12391_), .B(new_n5643_), .ZN(new_n12392_));
  OAI21_X1   g12200(.A1(new_n12389_), .A2(new_n12392_), .B(\asqrt[33] ), .ZN(new_n12393_));
  NAND3_X1   g12201(.A1(new_n12386_), .A2(new_n5029_), .A3(new_n12393_), .ZN(new_n12394_));
  AOI21_X1   g12202(.A1(new_n12386_), .A2(new_n12393_), .B(new_n5029_), .ZN(new_n12395_));
  AOI21_X1   g12203(.A1(new_n12218_), .A2(new_n12394_), .B(new_n12395_), .ZN(new_n12396_));
  AOI21_X1   g12204(.A1(new_n12396_), .A2(new_n4751_), .B(new_n12215_), .ZN(new_n12397_));
  INV_X1     g12205(.I(new_n12220_), .ZN(new_n12398_));
  NOR3_X1    g12206(.A1(new_n12389_), .A2(\asqrt[33] ), .A3(new_n12392_), .ZN(new_n12399_));
  OAI21_X1   g12207(.A1(new_n12398_), .A2(new_n12399_), .B(new_n12393_), .ZN(new_n12400_));
  OAI21_X1   g12208(.A1(new_n12400_), .A2(\asqrt[34] ), .B(new_n12218_), .ZN(new_n12401_));
  NAND2_X1   g12209(.A1(new_n12400_), .A2(\asqrt[34] ), .ZN(new_n12402_));
  AOI21_X1   g12210(.A1(new_n12401_), .A2(new_n12402_), .B(new_n4751_), .ZN(new_n12403_));
  NOR3_X1    g12211(.A1(new_n12397_), .A2(\asqrt[36] ), .A3(new_n12403_), .ZN(new_n12404_));
  OAI21_X1   g12212(.A1(new_n12397_), .A2(new_n12403_), .B(\asqrt[36] ), .ZN(new_n12405_));
  OAI21_X1   g12213(.A1(new_n12212_), .A2(new_n12404_), .B(new_n12405_), .ZN(new_n12406_));
  OAI21_X1   g12214(.A1(new_n12406_), .A2(\asqrt[37] ), .B(new_n12208_), .ZN(new_n12407_));
  NAND3_X1   g12215(.A1(new_n12401_), .A2(new_n12402_), .A3(new_n4751_), .ZN(new_n12408_));
  AOI21_X1   g12216(.A1(new_n12214_), .A2(new_n12408_), .B(new_n12403_), .ZN(new_n12409_));
  AOI21_X1   g12217(.A1(new_n12409_), .A2(new_n4461_), .B(new_n12212_), .ZN(new_n12410_));
  NAND2_X1   g12218(.A1(new_n12408_), .A2(new_n12214_), .ZN(new_n12411_));
  INV_X1     g12219(.I(new_n12403_), .ZN(new_n12412_));
  AOI21_X1   g12220(.A1(new_n12411_), .A2(new_n12412_), .B(new_n4461_), .ZN(new_n12413_));
  OAI21_X1   g12221(.A1(new_n12410_), .A2(new_n12413_), .B(\asqrt[37] ), .ZN(new_n12414_));
  NAND3_X1   g12222(.A1(new_n12407_), .A2(new_n3925_), .A3(new_n12414_), .ZN(new_n12415_));
  AOI21_X1   g12223(.A1(new_n12407_), .A2(new_n12414_), .B(new_n3925_), .ZN(new_n12416_));
  AOI21_X1   g12224(.A1(new_n12206_), .A2(new_n12415_), .B(new_n12416_), .ZN(new_n12417_));
  AOI21_X1   g12225(.A1(new_n12417_), .A2(new_n3681_), .B(new_n12203_), .ZN(new_n12418_));
  INV_X1     g12226(.I(new_n12208_), .ZN(new_n12419_));
  NOR3_X1    g12227(.A1(new_n12410_), .A2(\asqrt[37] ), .A3(new_n12413_), .ZN(new_n12420_));
  OAI21_X1   g12228(.A1(new_n12419_), .A2(new_n12420_), .B(new_n12414_), .ZN(new_n12421_));
  OAI21_X1   g12229(.A1(new_n12421_), .A2(\asqrt[38] ), .B(new_n12206_), .ZN(new_n12422_));
  NAND2_X1   g12230(.A1(new_n12421_), .A2(\asqrt[38] ), .ZN(new_n12423_));
  AOI21_X1   g12231(.A1(new_n12422_), .A2(new_n12423_), .B(new_n3681_), .ZN(new_n12424_));
  NOR3_X1    g12232(.A1(new_n12418_), .A2(\asqrt[40] ), .A3(new_n12424_), .ZN(new_n12425_));
  OAI21_X1   g12233(.A1(new_n12418_), .A2(new_n12424_), .B(\asqrt[40] ), .ZN(new_n12426_));
  OAI21_X1   g12234(.A1(new_n12200_), .A2(new_n12425_), .B(new_n12426_), .ZN(new_n12427_));
  OAI21_X1   g12235(.A1(new_n12427_), .A2(\asqrt[41] ), .B(new_n12196_), .ZN(new_n12428_));
  NAND3_X1   g12236(.A1(new_n12422_), .A2(new_n12423_), .A3(new_n3681_), .ZN(new_n12429_));
  AOI21_X1   g12237(.A1(new_n12202_), .A2(new_n12429_), .B(new_n12424_), .ZN(new_n12430_));
  AOI21_X1   g12238(.A1(new_n12430_), .A2(new_n3427_), .B(new_n12200_), .ZN(new_n12431_));
  NAND2_X1   g12239(.A1(new_n12429_), .A2(new_n12202_), .ZN(new_n12432_));
  INV_X1     g12240(.I(new_n12424_), .ZN(new_n12433_));
  AOI21_X1   g12241(.A1(new_n12432_), .A2(new_n12433_), .B(new_n3427_), .ZN(new_n12434_));
  OAI21_X1   g12242(.A1(new_n12431_), .A2(new_n12434_), .B(\asqrt[41] ), .ZN(new_n12435_));
  NAND3_X1   g12243(.A1(new_n12428_), .A2(new_n2960_), .A3(new_n12435_), .ZN(new_n12436_));
  AOI21_X1   g12244(.A1(new_n12428_), .A2(new_n12435_), .B(new_n2960_), .ZN(new_n12437_));
  AOI21_X1   g12245(.A1(new_n12194_), .A2(new_n12436_), .B(new_n12437_), .ZN(new_n12438_));
  AOI21_X1   g12246(.A1(new_n12438_), .A2(new_n2749_), .B(new_n12191_), .ZN(new_n12439_));
  INV_X1     g12247(.I(new_n12196_), .ZN(new_n12440_));
  NOR3_X1    g12248(.A1(new_n12431_), .A2(\asqrt[41] ), .A3(new_n12434_), .ZN(new_n12441_));
  OAI21_X1   g12249(.A1(new_n12440_), .A2(new_n12441_), .B(new_n12435_), .ZN(new_n12442_));
  OAI21_X1   g12250(.A1(new_n12442_), .A2(\asqrt[42] ), .B(new_n12194_), .ZN(new_n12443_));
  NAND2_X1   g12251(.A1(new_n12442_), .A2(\asqrt[42] ), .ZN(new_n12444_));
  AOI21_X1   g12252(.A1(new_n12443_), .A2(new_n12444_), .B(new_n2749_), .ZN(new_n12445_));
  NOR3_X1    g12253(.A1(new_n12439_), .A2(\asqrt[44] ), .A3(new_n12445_), .ZN(new_n12446_));
  OAI21_X1   g12254(.A1(new_n12439_), .A2(new_n12445_), .B(\asqrt[44] ), .ZN(new_n12447_));
  OAI21_X1   g12255(.A1(new_n12188_), .A2(new_n12446_), .B(new_n12447_), .ZN(new_n12448_));
  OAI21_X1   g12256(.A1(new_n12448_), .A2(\asqrt[45] ), .B(new_n12184_), .ZN(new_n12449_));
  NAND3_X1   g12257(.A1(new_n12443_), .A2(new_n12444_), .A3(new_n2749_), .ZN(new_n12450_));
  AOI21_X1   g12258(.A1(new_n12190_), .A2(new_n12450_), .B(new_n12445_), .ZN(new_n12451_));
  AOI21_X1   g12259(.A1(new_n12451_), .A2(new_n2531_), .B(new_n12188_), .ZN(new_n12452_));
  NAND2_X1   g12260(.A1(new_n12450_), .A2(new_n12190_), .ZN(new_n12453_));
  INV_X1     g12261(.I(new_n12445_), .ZN(new_n12454_));
  AOI21_X1   g12262(.A1(new_n12453_), .A2(new_n12454_), .B(new_n2531_), .ZN(new_n12455_));
  OAI21_X1   g12263(.A1(new_n12452_), .A2(new_n12455_), .B(\asqrt[45] ), .ZN(new_n12456_));
  NAND3_X1   g12264(.A1(new_n12449_), .A2(new_n2134_), .A3(new_n12456_), .ZN(new_n12457_));
  AOI21_X1   g12265(.A1(new_n12449_), .A2(new_n12456_), .B(new_n2134_), .ZN(new_n12458_));
  AOI21_X1   g12266(.A1(new_n12182_), .A2(new_n12457_), .B(new_n12458_), .ZN(new_n12459_));
  AOI21_X1   g12267(.A1(new_n12459_), .A2(new_n1953_), .B(new_n12179_), .ZN(new_n12460_));
  INV_X1     g12268(.I(new_n12184_), .ZN(new_n12461_));
  NOR3_X1    g12269(.A1(new_n12452_), .A2(\asqrt[45] ), .A3(new_n12455_), .ZN(new_n12462_));
  OAI21_X1   g12270(.A1(new_n12461_), .A2(new_n12462_), .B(new_n12456_), .ZN(new_n12463_));
  OAI21_X1   g12271(.A1(new_n12463_), .A2(\asqrt[46] ), .B(new_n12182_), .ZN(new_n12464_));
  NAND2_X1   g12272(.A1(new_n12463_), .A2(\asqrt[46] ), .ZN(new_n12465_));
  AOI21_X1   g12273(.A1(new_n12464_), .A2(new_n12465_), .B(new_n1953_), .ZN(new_n12466_));
  NOR3_X1    g12274(.A1(new_n12460_), .A2(\asqrt[48] ), .A3(new_n12466_), .ZN(new_n12467_));
  OAI21_X1   g12275(.A1(new_n12460_), .A2(new_n12466_), .B(\asqrt[48] ), .ZN(new_n12468_));
  OAI21_X1   g12276(.A1(new_n12176_), .A2(new_n12467_), .B(new_n12468_), .ZN(new_n12469_));
  OAI21_X1   g12277(.A1(new_n12469_), .A2(\asqrt[49] ), .B(new_n12172_), .ZN(new_n12470_));
  NAND3_X1   g12278(.A1(new_n12464_), .A2(new_n12465_), .A3(new_n1953_), .ZN(new_n12471_));
  AOI21_X1   g12279(.A1(new_n12178_), .A2(new_n12471_), .B(new_n12466_), .ZN(new_n12472_));
  AOI21_X1   g12280(.A1(new_n12472_), .A2(new_n1778_), .B(new_n12176_), .ZN(new_n12473_));
  NAND2_X1   g12281(.A1(new_n12471_), .A2(new_n12178_), .ZN(new_n12474_));
  INV_X1     g12282(.I(new_n12466_), .ZN(new_n12475_));
  AOI21_X1   g12283(.A1(new_n12474_), .A2(new_n12475_), .B(new_n1778_), .ZN(new_n12476_));
  OAI21_X1   g12284(.A1(new_n12473_), .A2(new_n12476_), .B(\asqrt[49] ), .ZN(new_n12477_));
  NAND3_X1   g12285(.A1(new_n12470_), .A2(new_n1463_), .A3(new_n12477_), .ZN(new_n12478_));
  INV_X1     g12286(.I(new_n12172_), .ZN(new_n12479_));
  NOR3_X1    g12287(.A1(new_n12473_), .A2(\asqrt[49] ), .A3(new_n12476_), .ZN(new_n12480_));
  OAI21_X1   g12288(.A1(new_n12479_), .A2(new_n12480_), .B(new_n12477_), .ZN(new_n12481_));
  NAND2_X1   g12289(.A1(new_n12481_), .A2(\asqrt[50] ), .ZN(new_n12482_));
  NOR2_X1    g12290(.A1(new_n12134_), .A2(\asqrt[62] ), .ZN(new_n12483_));
  NOR2_X1    g12291(.A1(new_n12483_), .A2(new_n12276_), .ZN(new_n12484_));
  XOR2_X1    g12292(.A1(new_n12150_), .A2(new_n11664_), .Z(new_n12485_));
  OAI21_X1   g12293(.A1(\asqrt[15] ), .A2(new_n12484_), .B(new_n12485_), .ZN(new_n12486_));
  INV_X1     g12294(.I(new_n12486_), .ZN(new_n12487_));
  AOI21_X1   g12295(.A1(new_n12119_), .A2(new_n12127_), .B(\asqrt[15] ), .ZN(new_n12488_));
  XOR2_X1    g12296(.A1(new_n12488_), .A2(new_n12034_), .Z(new_n12489_));
  INV_X1     g12297(.I(new_n12489_), .ZN(new_n12490_));
  AOI21_X1   g12298(.A1(new_n12110_), .A2(new_n12118_), .B(\asqrt[15] ), .ZN(new_n12491_));
  XOR2_X1    g12299(.A1(new_n12491_), .A2(new_n12036_), .Z(new_n12492_));
  INV_X1     g12300(.I(new_n12492_), .ZN(new_n12493_));
  NAND2_X1   g12301(.A1(new_n12114_), .A2(new_n531_), .ZN(new_n12494_));
  AOI21_X1   g12302(.A1(new_n12494_), .A2(new_n12109_), .B(\asqrt[15] ), .ZN(new_n12495_));
  XOR2_X1    g12303(.A1(new_n12495_), .A2(new_n12038_), .Z(new_n12496_));
  AOI21_X1   g12304(.A1(new_n12113_), .A2(new_n12099_), .B(\asqrt[15] ), .ZN(new_n12497_));
  XOR2_X1    g12305(.A1(new_n12497_), .A2(new_n12042_), .Z(new_n12498_));
  NAND2_X1   g12306(.A1(new_n12081_), .A2(new_n744_), .ZN(new_n12499_));
  AOI21_X1   g12307(.A1(new_n12499_), .A2(new_n12107_), .B(\asqrt[15] ), .ZN(new_n12500_));
  XOR2_X1    g12308(.A1(new_n12500_), .A2(new_n12046_), .Z(new_n12501_));
  INV_X1     g12309(.I(new_n12501_), .ZN(new_n12502_));
  AOI21_X1   g12310(.A1(new_n12079_), .A2(new_n12096_), .B(\asqrt[15] ), .ZN(new_n12503_));
  XOR2_X1    g12311(.A1(new_n12503_), .A2(new_n12049_), .Z(new_n12504_));
  INV_X1     g12312(.I(new_n12504_), .ZN(new_n12505_));
  NAND2_X1   g12313(.A1(new_n12092_), .A2(new_n1006_), .ZN(new_n12506_));
  AOI21_X1   g12314(.A1(new_n12506_), .A2(new_n12078_), .B(\asqrt[15] ), .ZN(new_n12507_));
  XOR2_X1    g12315(.A1(new_n12507_), .A2(new_n12051_), .Z(new_n12508_));
  AOI21_X1   g12316(.A1(new_n12090_), .A2(new_n12075_), .B(\asqrt[15] ), .ZN(new_n12509_));
  XOR2_X1    g12317(.A1(new_n12509_), .A2(new_n12054_), .Z(new_n12510_));
  NAND2_X1   g12318(.A1(new_n12065_), .A2(new_n1305_), .ZN(new_n12511_));
  AOI21_X1   g12319(.A1(new_n12511_), .A2(new_n12089_), .B(\asqrt[15] ), .ZN(new_n12512_));
  XOR2_X1    g12320(.A1(new_n12512_), .A2(new_n12058_), .Z(new_n12513_));
  INV_X1     g12321(.I(new_n12513_), .ZN(new_n12514_));
  AOI21_X1   g12322(.A1(new_n12063_), .A2(new_n12072_), .B(\asqrt[15] ), .ZN(new_n12515_));
  XOR2_X1    g12323(.A1(new_n12515_), .A2(new_n12061_), .Z(new_n12516_));
  INV_X1     g12324(.I(new_n12516_), .ZN(new_n12517_));
  AOI21_X1   g12325(.A1(new_n12470_), .A2(new_n12477_), .B(new_n1463_), .ZN(new_n12518_));
  AOI21_X1   g12326(.A1(new_n12170_), .A2(new_n12478_), .B(new_n12518_), .ZN(new_n12519_));
  AOI21_X1   g12327(.A1(new_n12519_), .A2(new_n1305_), .B(new_n12517_), .ZN(new_n12520_));
  OAI21_X1   g12328(.A1(new_n12481_), .A2(\asqrt[50] ), .B(new_n12170_), .ZN(new_n12521_));
  AOI21_X1   g12329(.A1(new_n12521_), .A2(new_n12482_), .B(new_n1305_), .ZN(new_n12522_));
  NOR3_X1    g12330(.A1(new_n12520_), .A2(\asqrt[52] ), .A3(new_n12522_), .ZN(new_n12523_));
  OAI21_X1   g12331(.A1(new_n12520_), .A2(new_n12522_), .B(\asqrt[52] ), .ZN(new_n12524_));
  OAI21_X1   g12332(.A1(new_n12514_), .A2(new_n12523_), .B(new_n12524_), .ZN(new_n12525_));
  OAI21_X1   g12333(.A1(new_n12525_), .A2(\asqrt[53] ), .B(new_n12510_), .ZN(new_n12526_));
  NAND3_X1   g12334(.A1(new_n12521_), .A2(new_n12482_), .A3(new_n1305_), .ZN(new_n12527_));
  AOI21_X1   g12335(.A1(new_n12516_), .A2(new_n12527_), .B(new_n12522_), .ZN(new_n12528_));
  AOI21_X1   g12336(.A1(new_n12528_), .A2(new_n1150_), .B(new_n12514_), .ZN(new_n12529_));
  NAND2_X1   g12337(.A1(new_n12527_), .A2(new_n12516_), .ZN(new_n12530_));
  INV_X1     g12338(.I(new_n12522_), .ZN(new_n12531_));
  AOI21_X1   g12339(.A1(new_n12530_), .A2(new_n12531_), .B(new_n1150_), .ZN(new_n12532_));
  OAI21_X1   g12340(.A1(new_n12529_), .A2(new_n12532_), .B(\asqrt[53] ), .ZN(new_n12533_));
  NAND3_X1   g12341(.A1(new_n12526_), .A2(new_n860_), .A3(new_n12533_), .ZN(new_n12534_));
  AOI21_X1   g12342(.A1(new_n12526_), .A2(new_n12533_), .B(new_n860_), .ZN(new_n12535_));
  AOI21_X1   g12343(.A1(new_n12508_), .A2(new_n12534_), .B(new_n12535_), .ZN(new_n12536_));
  AOI21_X1   g12344(.A1(new_n12536_), .A2(new_n744_), .B(new_n12505_), .ZN(new_n12537_));
  INV_X1     g12345(.I(new_n12510_), .ZN(new_n12538_));
  NOR3_X1    g12346(.A1(new_n12529_), .A2(\asqrt[53] ), .A3(new_n12532_), .ZN(new_n12539_));
  OAI21_X1   g12347(.A1(new_n12538_), .A2(new_n12539_), .B(new_n12533_), .ZN(new_n12540_));
  OAI21_X1   g12348(.A1(new_n12540_), .A2(\asqrt[54] ), .B(new_n12508_), .ZN(new_n12541_));
  NAND2_X1   g12349(.A1(new_n12540_), .A2(\asqrt[54] ), .ZN(new_n12542_));
  AOI21_X1   g12350(.A1(new_n12541_), .A2(new_n12542_), .B(new_n744_), .ZN(new_n12543_));
  NOR3_X1    g12351(.A1(new_n12537_), .A2(\asqrt[56] ), .A3(new_n12543_), .ZN(new_n12544_));
  OAI21_X1   g12352(.A1(new_n12537_), .A2(new_n12543_), .B(\asqrt[56] ), .ZN(new_n12545_));
  OAI21_X1   g12353(.A1(new_n12502_), .A2(new_n12544_), .B(new_n12545_), .ZN(new_n12546_));
  OAI21_X1   g12354(.A1(new_n12546_), .A2(\asqrt[57] ), .B(new_n12498_), .ZN(new_n12547_));
  NAND3_X1   g12355(.A1(new_n12541_), .A2(new_n12542_), .A3(new_n744_), .ZN(new_n12548_));
  AOI21_X1   g12356(.A1(new_n12504_), .A2(new_n12548_), .B(new_n12543_), .ZN(new_n12549_));
  AOI21_X1   g12357(.A1(new_n12549_), .A2(new_n634_), .B(new_n12502_), .ZN(new_n12550_));
  NAND2_X1   g12358(.A1(new_n12548_), .A2(new_n12504_), .ZN(new_n12551_));
  INV_X1     g12359(.I(new_n12543_), .ZN(new_n12552_));
  AOI21_X1   g12360(.A1(new_n12551_), .A2(new_n12552_), .B(new_n634_), .ZN(new_n12553_));
  OAI21_X1   g12361(.A1(new_n12550_), .A2(new_n12553_), .B(\asqrt[57] ), .ZN(new_n12554_));
  NAND3_X1   g12362(.A1(new_n12547_), .A2(new_n423_), .A3(new_n12554_), .ZN(new_n12555_));
  AOI21_X1   g12363(.A1(new_n12547_), .A2(new_n12554_), .B(new_n423_), .ZN(new_n12556_));
  AOI21_X1   g12364(.A1(new_n12496_), .A2(new_n12555_), .B(new_n12556_), .ZN(new_n12557_));
  AOI21_X1   g12365(.A1(new_n12557_), .A2(new_n337_), .B(new_n12493_), .ZN(new_n12558_));
  NOR2_X1    g12366(.A1(new_n12557_), .A2(new_n337_), .ZN(new_n12559_));
  NOR3_X1    g12367(.A1(new_n12558_), .A2(new_n12559_), .A3(\asqrt[60] ), .ZN(new_n12560_));
  OAI21_X1   g12368(.A1(new_n12558_), .A2(new_n12559_), .B(\asqrt[60] ), .ZN(new_n12561_));
  OAI21_X1   g12369(.A1(new_n12490_), .A2(new_n12560_), .B(new_n12561_), .ZN(new_n12562_));
  NAND2_X1   g12370(.A1(new_n12562_), .A2(\asqrt[61] ), .ZN(new_n12563_));
  AOI21_X1   g12371(.A1(new_n12135_), .A2(new_n12141_), .B(\asqrt[15] ), .ZN(new_n12564_));
  XOR2_X1    g12372(.A1(new_n12564_), .A2(new_n12030_), .Z(new_n12565_));
  OAI21_X1   g12373(.A1(new_n12562_), .A2(\asqrt[61] ), .B(new_n12565_), .ZN(new_n12566_));
  NAND2_X1   g12374(.A1(new_n12566_), .A2(new_n12563_), .ZN(new_n12567_));
  INV_X1     g12375(.I(new_n12498_), .ZN(new_n12568_));
  NOR3_X1    g12376(.A1(new_n12550_), .A2(\asqrt[57] ), .A3(new_n12553_), .ZN(new_n12569_));
  OAI21_X1   g12377(.A1(new_n12568_), .A2(new_n12569_), .B(new_n12554_), .ZN(new_n12570_));
  OAI21_X1   g12378(.A1(new_n12570_), .A2(\asqrt[58] ), .B(new_n12496_), .ZN(new_n12571_));
  NOR2_X1    g12379(.A1(new_n12569_), .A2(new_n12568_), .ZN(new_n12572_));
  INV_X1     g12380(.I(new_n12554_), .ZN(new_n12573_));
  OAI21_X1   g12381(.A1(new_n12572_), .A2(new_n12573_), .B(\asqrt[58] ), .ZN(new_n12574_));
  NAND3_X1   g12382(.A1(new_n12571_), .A2(new_n337_), .A3(new_n12574_), .ZN(new_n12575_));
  NAND2_X1   g12383(.A1(new_n12575_), .A2(new_n12492_), .ZN(new_n12576_));
  INV_X1     g12384(.I(new_n12496_), .ZN(new_n12577_));
  NOR2_X1    g12385(.A1(new_n12572_), .A2(new_n12573_), .ZN(new_n12578_));
  AOI21_X1   g12386(.A1(new_n12578_), .A2(new_n423_), .B(new_n12577_), .ZN(new_n12579_));
  OAI21_X1   g12387(.A1(new_n12579_), .A2(new_n12556_), .B(\asqrt[59] ), .ZN(new_n12580_));
  NAND3_X1   g12388(.A1(new_n12576_), .A2(new_n266_), .A3(new_n12580_), .ZN(new_n12581_));
  NAND2_X1   g12389(.A1(new_n12581_), .A2(new_n12489_), .ZN(new_n12582_));
  AOI21_X1   g12390(.A1(new_n12582_), .A2(new_n12561_), .B(new_n239_), .ZN(new_n12583_));
  AOI21_X1   g12391(.A1(new_n12576_), .A2(new_n12580_), .B(new_n266_), .ZN(new_n12584_));
  AOI21_X1   g12392(.A1(new_n12489_), .A2(new_n12581_), .B(new_n12584_), .ZN(new_n12585_));
  INV_X1     g12393(.I(new_n12565_), .ZN(new_n12586_));
  AOI21_X1   g12394(.A1(new_n12585_), .A2(new_n239_), .B(new_n12586_), .ZN(new_n12587_));
  OAI21_X1   g12395(.A1(new_n12587_), .A2(new_n12583_), .B(new_n201_), .ZN(new_n12588_));
  NAND3_X1   g12396(.A1(new_n12566_), .A2(new_n12563_), .A3(\asqrt[62] ), .ZN(new_n12589_));
  NOR2_X1    g12397(.A1(new_n12133_), .A2(new_n12142_), .ZN(new_n12590_));
  NOR2_X1    g12398(.A1(\asqrt[15] ), .A2(new_n12590_), .ZN(new_n12591_));
  XOR2_X1    g12399(.A1(new_n12591_), .A2(new_n12131_), .Z(new_n12592_));
  INV_X1     g12400(.I(new_n12592_), .ZN(new_n12593_));
  AOI22_X1   g12401(.A1(new_n12589_), .A2(new_n12588_), .B1(new_n12567_), .B2(new_n12593_), .ZN(new_n12594_));
  NOR2_X1    g12402(.A1(new_n12153_), .A2(new_n12027_), .ZN(new_n12595_));
  OAI21_X1   g12403(.A1(\asqrt[15] ), .A2(new_n12595_), .B(new_n12160_), .ZN(new_n12596_));
  INV_X1     g12404(.I(new_n12596_), .ZN(new_n12597_));
  OAI21_X1   g12405(.A1(new_n12594_), .A2(new_n12487_), .B(new_n12597_), .ZN(new_n12598_));
  OAI21_X1   g12406(.A1(new_n12567_), .A2(\asqrt[62] ), .B(new_n12592_), .ZN(new_n12599_));
  NAND2_X1   g12407(.A1(new_n12567_), .A2(\asqrt[62] ), .ZN(new_n12600_));
  NAND3_X1   g12408(.A1(new_n12599_), .A2(new_n12600_), .A3(new_n12487_), .ZN(new_n12601_));
  NAND2_X1   g12409(.A1(new_n12153_), .A2(new_n12026_), .ZN(new_n12602_));
  NAND2_X1   g12410(.A1(new_n12273_), .A2(new_n12027_), .ZN(new_n12603_));
  AOI21_X1   g12411(.A1(new_n12602_), .A2(new_n12603_), .B(new_n193_), .ZN(new_n12604_));
  OAI21_X1   g12412(.A1(\asqrt[15] ), .A2(new_n12027_), .B(new_n12604_), .ZN(new_n12605_));
  NOR2_X1    g12413(.A1(new_n12166_), .A2(new_n12026_), .ZN(new_n12606_));
  NAND4_X1   g12414(.A1(new_n12157_), .A2(new_n193_), .A3(new_n12160_), .A4(new_n12606_), .ZN(new_n12607_));
  NAND2_X1   g12415(.A1(new_n12605_), .A2(new_n12607_), .ZN(new_n12608_));
  INV_X1     g12416(.I(new_n12608_), .ZN(new_n12609_));
  NAND4_X1   g12417(.A1(new_n12598_), .A2(new_n193_), .A3(new_n12601_), .A4(new_n12609_), .ZN(\asqrt[14] ));
  AOI21_X1   g12418(.A1(new_n12478_), .A2(new_n12482_), .B(\asqrt[14] ), .ZN(new_n12611_));
  XOR2_X1    g12419(.A1(new_n12611_), .A2(new_n12170_), .Z(new_n12612_));
  XOR2_X1    g12420(.A1(new_n12469_), .A2(\asqrt[49] ), .Z(new_n12613_));
  NOR2_X1    g12421(.A1(\asqrt[14] ), .A2(new_n12613_), .ZN(new_n12614_));
  XOR2_X1    g12422(.A1(new_n12614_), .A2(new_n12172_), .Z(new_n12615_));
  NOR2_X1    g12423(.A1(new_n12467_), .A2(new_n12476_), .ZN(new_n12616_));
  NOR2_X1    g12424(.A1(\asqrt[14] ), .A2(new_n12616_), .ZN(new_n12617_));
  XOR2_X1    g12425(.A1(new_n12617_), .A2(new_n12175_), .Z(new_n12618_));
  AOI21_X1   g12426(.A1(new_n12471_), .A2(new_n12475_), .B(\asqrt[14] ), .ZN(new_n12619_));
  XOR2_X1    g12427(.A1(new_n12619_), .A2(new_n12178_), .Z(new_n12620_));
  INV_X1     g12428(.I(new_n12620_), .ZN(new_n12621_));
  AOI21_X1   g12429(.A1(new_n12457_), .A2(new_n12465_), .B(\asqrt[14] ), .ZN(new_n12622_));
  XOR2_X1    g12430(.A1(new_n12622_), .A2(new_n12182_), .Z(new_n12623_));
  INV_X1     g12431(.I(new_n12623_), .ZN(new_n12624_));
  XOR2_X1    g12432(.A1(new_n12448_), .A2(\asqrt[45] ), .Z(new_n12625_));
  NOR2_X1    g12433(.A1(\asqrt[14] ), .A2(new_n12625_), .ZN(new_n12626_));
  XOR2_X1    g12434(.A1(new_n12626_), .A2(new_n12184_), .Z(new_n12627_));
  NOR2_X1    g12435(.A1(new_n12446_), .A2(new_n12455_), .ZN(new_n12628_));
  NOR2_X1    g12436(.A1(\asqrt[14] ), .A2(new_n12628_), .ZN(new_n12629_));
  XOR2_X1    g12437(.A1(new_n12629_), .A2(new_n12187_), .Z(new_n12630_));
  AOI21_X1   g12438(.A1(new_n12450_), .A2(new_n12454_), .B(\asqrt[14] ), .ZN(new_n12631_));
  XOR2_X1    g12439(.A1(new_n12631_), .A2(new_n12190_), .Z(new_n12632_));
  INV_X1     g12440(.I(new_n12632_), .ZN(new_n12633_));
  AOI21_X1   g12441(.A1(new_n12436_), .A2(new_n12444_), .B(\asqrt[14] ), .ZN(new_n12634_));
  XOR2_X1    g12442(.A1(new_n12634_), .A2(new_n12194_), .Z(new_n12635_));
  INV_X1     g12443(.I(new_n12635_), .ZN(new_n12636_));
  XOR2_X1    g12444(.A1(new_n12427_), .A2(\asqrt[41] ), .Z(new_n12637_));
  NOR2_X1    g12445(.A1(\asqrt[14] ), .A2(new_n12637_), .ZN(new_n12638_));
  XOR2_X1    g12446(.A1(new_n12638_), .A2(new_n12196_), .Z(new_n12639_));
  NOR2_X1    g12447(.A1(new_n12425_), .A2(new_n12434_), .ZN(new_n12640_));
  NOR2_X1    g12448(.A1(\asqrt[14] ), .A2(new_n12640_), .ZN(new_n12641_));
  XOR2_X1    g12449(.A1(new_n12641_), .A2(new_n12199_), .Z(new_n12642_));
  AOI21_X1   g12450(.A1(new_n12429_), .A2(new_n12433_), .B(\asqrt[14] ), .ZN(new_n12643_));
  XOR2_X1    g12451(.A1(new_n12643_), .A2(new_n12202_), .Z(new_n12644_));
  INV_X1     g12452(.I(new_n12644_), .ZN(new_n12645_));
  AOI21_X1   g12453(.A1(new_n12415_), .A2(new_n12423_), .B(\asqrt[14] ), .ZN(new_n12646_));
  XOR2_X1    g12454(.A1(new_n12646_), .A2(new_n12206_), .Z(new_n12647_));
  INV_X1     g12455(.I(new_n12647_), .ZN(new_n12648_));
  XOR2_X1    g12456(.A1(new_n12406_), .A2(\asqrt[37] ), .Z(new_n12649_));
  NOR2_X1    g12457(.A1(\asqrt[14] ), .A2(new_n12649_), .ZN(new_n12650_));
  XOR2_X1    g12458(.A1(new_n12650_), .A2(new_n12208_), .Z(new_n12651_));
  NOR2_X1    g12459(.A1(new_n12404_), .A2(new_n12413_), .ZN(new_n12652_));
  NOR2_X1    g12460(.A1(\asqrt[14] ), .A2(new_n12652_), .ZN(new_n12653_));
  XOR2_X1    g12461(.A1(new_n12653_), .A2(new_n12211_), .Z(new_n12654_));
  AOI21_X1   g12462(.A1(new_n12408_), .A2(new_n12412_), .B(\asqrt[14] ), .ZN(new_n12655_));
  XOR2_X1    g12463(.A1(new_n12655_), .A2(new_n12214_), .Z(new_n12656_));
  INV_X1     g12464(.I(new_n12656_), .ZN(new_n12657_));
  AOI21_X1   g12465(.A1(new_n12394_), .A2(new_n12402_), .B(\asqrt[14] ), .ZN(new_n12658_));
  XOR2_X1    g12466(.A1(new_n12658_), .A2(new_n12218_), .Z(new_n12659_));
  INV_X1     g12467(.I(new_n12659_), .ZN(new_n12660_));
  XOR2_X1    g12468(.A1(new_n12385_), .A2(\asqrt[33] ), .Z(new_n12661_));
  NOR2_X1    g12469(.A1(\asqrt[14] ), .A2(new_n12661_), .ZN(new_n12662_));
  XOR2_X1    g12470(.A1(new_n12662_), .A2(new_n12220_), .Z(new_n12663_));
  NOR2_X1    g12471(.A1(new_n12383_), .A2(new_n12392_), .ZN(new_n12664_));
  NOR2_X1    g12472(.A1(\asqrt[14] ), .A2(new_n12664_), .ZN(new_n12665_));
  XOR2_X1    g12473(.A1(new_n12665_), .A2(new_n12223_), .Z(new_n12666_));
  AOI21_X1   g12474(.A1(new_n12387_), .A2(new_n12391_), .B(\asqrt[14] ), .ZN(new_n12667_));
  XOR2_X1    g12475(.A1(new_n12667_), .A2(new_n12226_), .Z(new_n12668_));
  INV_X1     g12476(.I(new_n12668_), .ZN(new_n12669_));
  AOI21_X1   g12477(.A1(new_n12373_), .A2(new_n12381_), .B(\asqrt[14] ), .ZN(new_n12670_));
  XOR2_X1    g12478(.A1(new_n12670_), .A2(new_n12230_), .Z(new_n12671_));
  INV_X1     g12479(.I(new_n12671_), .ZN(new_n12672_));
  XOR2_X1    g12480(.A1(new_n12364_), .A2(\asqrt[29] ), .Z(new_n12673_));
  NOR2_X1    g12481(.A1(\asqrt[14] ), .A2(new_n12673_), .ZN(new_n12674_));
  XOR2_X1    g12482(.A1(new_n12674_), .A2(new_n12232_), .Z(new_n12675_));
  NOR2_X1    g12483(.A1(new_n12362_), .A2(new_n12371_), .ZN(new_n12676_));
  NOR2_X1    g12484(.A1(\asqrt[14] ), .A2(new_n12676_), .ZN(new_n12677_));
  XOR2_X1    g12485(.A1(new_n12677_), .A2(new_n12235_), .Z(new_n12678_));
  AOI21_X1   g12486(.A1(new_n12366_), .A2(new_n12370_), .B(\asqrt[14] ), .ZN(new_n12679_));
  XOR2_X1    g12487(.A1(new_n12679_), .A2(new_n12238_), .Z(new_n12680_));
  INV_X1     g12488(.I(new_n12680_), .ZN(new_n12681_));
  AOI21_X1   g12489(.A1(new_n12352_), .A2(new_n12360_), .B(\asqrt[14] ), .ZN(new_n12682_));
  XOR2_X1    g12490(.A1(new_n12682_), .A2(new_n12242_), .Z(new_n12683_));
  INV_X1     g12491(.I(new_n12683_), .ZN(new_n12684_));
  XOR2_X1    g12492(.A1(new_n12343_), .A2(\asqrt[25] ), .Z(new_n12685_));
  NOR2_X1    g12493(.A1(\asqrt[14] ), .A2(new_n12685_), .ZN(new_n12686_));
  XOR2_X1    g12494(.A1(new_n12686_), .A2(new_n12244_), .Z(new_n12687_));
  NOR2_X1    g12495(.A1(new_n12341_), .A2(new_n12350_), .ZN(new_n12688_));
  NOR2_X1    g12496(.A1(\asqrt[14] ), .A2(new_n12688_), .ZN(new_n12689_));
  XOR2_X1    g12497(.A1(new_n12689_), .A2(new_n12247_), .Z(new_n12690_));
  AOI21_X1   g12498(.A1(new_n12345_), .A2(new_n12349_), .B(\asqrt[14] ), .ZN(new_n12691_));
  XOR2_X1    g12499(.A1(new_n12691_), .A2(new_n12250_), .Z(new_n12692_));
  INV_X1     g12500(.I(new_n12692_), .ZN(new_n12693_));
  AOI21_X1   g12501(.A1(new_n12331_), .A2(new_n12339_), .B(\asqrt[14] ), .ZN(new_n12694_));
  XOR2_X1    g12502(.A1(new_n12694_), .A2(new_n12254_), .Z(new_n12695_));
  INV_X1     g12503(.I(new_n12695_), .ZN(new_n12696_));
  XOR2_X1    g12504(.A1(new_n12322_), .A2(\asqrt[21] ), .Z(new_n12697_));
  NOR2_X1    g12505(.A1(\asqrt[14] ), .A2(new_n12697_), .ZN(new_n12698_));
  XOR2_X1    g12506(.A1(new_n12698_), .A2(new_n12256_), .Z(new_n12699_));
  NOR2_X1    g12507(.A1(new_n12320_), .A2(new_n12329_), .ZN(new_n12700_));
  NOR2_X1    g12508(.A1(\asqrt[14] ), .A2(new_n12700_), .ZN(new_n12701_));
  XOR2_X1    g12509(.A1(new_n12701_), .A2(new_n12259_), .Z(new_n12702_));
  AOI21_X1   g12510(.A1(new_n12324_), .A2(new_n12328_), .B(\asqrt[14] ), .ZN(new_n12703_));
  XOR2_X1    g12511(.A1(new_n12703_), .A2(new_n12262_), .Z(new_n12704_));
  INV_X1     g12512(.I(new_n12704_), .ZN(new_n12705_));
  AOI21_X1   g12513(.A1(new_n12310_), .A2(new_n12318_), .B(\asqrt[14] ), .ZN(new_n12706_));
  XOR2_X1    g12514(.A1(new_n12706_), .A2(new_n12269_), .Z(new_n12707_));
  INV_X1     g12515(.I(new_n12707_), .ZN(new_n12708_));
  AOI21_X1   g12516(.A1(new_n12301_), .A2(new_n12309_), .B(\asqrt[14] ), .ZN(new_n12709_));
  XOR2_X1    g12517(.A1(new_n12709_), .A2(new_n12286_), .Z(new_n12710_));
  NAND2_X1   g12518(.A1(\asqrt[15] ), .A2(new_n12287_), .ZN(new_n12711_));
  NOR2_X1    g12519(.A1(new_n12298_), .A2(\a[30] ), .ZN(new_n12712_));
  AOI22_X1   g12520(.A1(new_n12711_), .A2(new_n12298_), .B1(\asqrt[15] ), .B2(new_n12712_), .ZN(new_n12713_));
  AOI21_X1   g12521(.A1(\asqrt[15] ), .A2(\a[30] ), .B(new_n12295_), .ZN(new_n12714_));
  NOR2_X1    g12522(.A1(new_n12305_), .A2(new_n12714_), .ZN(new_n12715_));
  NOR2_X1    g12523(.A1(\asqrt[14] ), .A2(new_n12715_), .ZN(new_n12716_));
  XOR2_X1    g12524(.A1(new_n12716_), .A2(new_n12713_), .Z(new_n12717_));
  NOR2_X1    g12525(.A1(new_n12587_), .A2(new_n12583_), .ZN(new_n12718_));
  AOI21_X1   g12526(.A1(new_n12566_), .A2(new_n12563_), .B(\asqrt[62] ), .ZN(new_n12719_));
  NOR3_X1    g12527(.A1(new_n12587_), .A2(new_n201_), .A3(new_n12583_), .ZN(new_n12720_));
  OAI22_X1   g12528(.A1(new_n12719_), .A2(new_n12720_), .B1(new_n12718_), .B2(new_n12592_), .ZN(new_n12721_));
  AOI21_X1   g12529(.A1(new_n12721_), .A2(new_n12486_), .B(new_n12596_), .ZN(new_n12722_));
  AOI21_X1   g12530(.A1(new_n12718_), .A2(new_n201_), .B(new_n12593_), .ZN(new_n12723_));
  NOR2_X1    g12531(.A1(new_n12718_), .A2(new_n201_), .ZN(new_n12724_));
  NOR3_X1    g12532(.A1(new_n12723_), .A2(new_n12724_), .A3(new_n12486_), .ZN(new_n12725_));
  NOR3_X1    g12533(.A1(new_n12722_), .A2(\asqrt[63] ), .A3(new_n12725_), .ZN(new_n12726_));
  NAND4_X1   g12534(.A1(new_n12726_), .A2(\asqrt[15] ), .A3(new_n12605_), .A4(new_n12607_), .ZN(new_n12727_));
  NAND2_X1   g12535(.A1(\asqrt[14] ), .A2(new_n12288_), .ZN(new_n12728_));
  AOI21_X1   g12536(.A1(new_n12727_), .A2(new_n12728_), .B(\a[30] ), .ZN(new_n12729_));
  NAND2_X1   g12537(.A1(new_n12598_), .A2(new_n193_), .ZN(new_n12730_));
  NAND3_X1   g12538(.A1(new_n12605_), .A2(new_n12607_), .A3(\asqrt[15] ), .ZN(new_n12731_));
  NOR3_X1    g12539(.A1(new_n12730_), .A2(new_n12725_), .A3(new_n12731_), .ZN(new_n12732_));
  NOR4_X1    g12540(.A1(new_n12722_), .A2(\asqrt[63] ), .A3(new_n12725_), .A4(new_n12608_), .ZN(new_n12733_));
  NOR2_X1    g12541(.A1(new_n12733_), .A2(new_n12290_), .ZN(new_n12734_));
  NOR3_X1    g12542(.A1(new_n12734_), .A2(new_n12732_), .A3(new_n12287_), .ZN(new_n12735_));
  OR2_X2     g12543(.A1(new_n12729_), .A2(new_n12735_), .Z(new_n12736_));
  NOR2_X1    g12544(.A1(\a[26] ), .A2(\a[27] ), .ZN(new_n12737_));
  INV_X1     g12545(.I(new_n12737_), .ZN(new_n12738_));
  NAND3_X1   g12546(.A1(\asqrt[14] ), .A2(\a[28] ), .A3(new_n12738_), .ZN(new_n12739_));
  INV_X1     g12547(.I(\a[28] ), .ZN(new_n12740_));
  OAI21_X1   g12548(.A1(\asqrt[14] ), .A2(new_n12740_), .B(new_n12737_), .ZN(new_n12741_));
  AOI21_X1   g12549(.A1(new_n12741_), .A2(new_n12739_), .B(new_n12283_), .ZN(new_n12742_));
  NOR3_X1    g12550(.A1(new_n12274_), .A2(\asqrt[63] ), .A3(new_n12277_), .ZN(new_n12743_));
  NAND2_X1   g12551(.A1(new_n12737_), .A2(new_n12740_), .ZN(new_n12744_));
  NAND3_X1   g12552(.A1(new_n12163_), .A2(new_n12165_), .A3(new_n12744_), .ZN(new_n12745_));
  NAND2_X1   g12553(.A1(new_n12743_), .A2(new_n12745_), .ZN(new_n12746_));
  NAND3_X1   g12554(.A1(\asqrt[14] ), .A2(\a[28] ), .A3(new_n12746_), .ZN(new_n12747_));
  INV_X1     g12555(.I(\a[29] ), .ZN(new_n12748_));
  NAND3_X1   g12556(.A1(\asqrt[14] ), .A2(new_n12740_), .A3(new_n12748_), .ZN(new_n12749_));
  OAI21_X1   g12557(.A1(new_n12733_), .A2(\a[28] ), .B(\a[29] ), .ZN(new_n12750_));
  NAND3_X1   g12558(.A1(new_n12747_), .A2(new_n12750_), .A3(new_n12749_), .ZN(new_n12751_));
  NOR3_X1    g12559(.A1(new_n12751_), .A2(new_n12742_), .A3(\asqrt[16] ), .ZN(new_n12752_));
  OAI21_X1   g12560(.A1(new_n12751_), .A2(new_n12742_), .B(\asqrt[16] ), .ZN(new_n12753_));
  OAI21_X1   g12561(.A1(new_n12736_), .A2(new_n12752_), .B(new_n12753_), .ZN(new_n12754_));
  OAI21_X1   g12562(.A1(new_n12754_), .A2(\asqrt[17] ), .B(new_n12717_), .ZN(new_n12755_));
  NAND2_X1   g12563(.A1(new_n12754_), .A2(\asqrt[17] ), .ZN(new_n12756_));
  NAND3_X1   g12564(.A1(new_n12755_), .A2(new_n12756_), .A3(new_n10914_), .ZN(new_n12757_));
  AOI21_X1   g12565(.A1(new_n12755_), .A2(new_n12756_), .B(new_n10914_), .ZN(new_n12758_));
  AOI21_X1   g12566(.A1(new_n12710_), .A2(new_n12757_), .B(new_n12758_), .ZN(new_n12759_));
  AOI21_X1   g12567(.A1(new_n12759_), .A2(new_n10497_), .B(new_n12708_), .ZN(new_n12760_));
  NAND2_X1   g12568(.A1(new_n12757_), .A2(new_n12710_), .ZN(new_n12761_));
  INV_X1     g12569(.I(new_n12717_), .ZN(new_n12762_));
  NOR2_X1    g12570(.A1(new_n12729_), .A2(new_n12735_), .ZN(new_n12763_));
  NOR3_X1    g12571(.A1(new_n12733_), .A2(new_n12740_), .A3(new_n12737_), .ZN(new_n12764_));
  AOI21_X1   g12572(.A1(new_n12733_), .A2(\a[28] ), .B(new_n12738_), .ZN(new_n12765_));
  OAI21_X1   g12573(.A1(new_n12764_), .A2(new_n12765_), .B(\asqrt[15] ), .ZN(new_n12766_));
  INV_X1     g12574(.I(new_n12746_), .ZN(new_n12767_));
  NOR3_X1    g12575(.A1(new_n12733_), .A2(new_n12740_), .A3(new_n12767_), .ZN(new_n12768_));
  NOR3_X1    g12576(.A1(new_n12733_), .A2(\a[28] ), .A3(\a[29] ), .ZN(new_n12769_));
  AOI21_X1   g12577(.A1(\asqrt[14] ), .A2(new_n12740_), .B(new_n12748_), .ZN(new_n12770_));
  NOR3_X1    g12578(.A1(new_n12768_), .A2(new_n12769_), .A3(new_n12770_), .ZN(new_n12771_));
  NAND3_X1   g12579(.A1(new_n12771_), .A2(new_n12766_), .A3(new_n11802_), .ZN(new_n12772_));
  AOI21_X1   g12580(.A1(new_n12771_), .A2(new_n12766_), .B(new_n11802_), .ZN(new_n12773_));
  AOI21_X1   g12581(.A1(new_n12763_), .A2(new_n12772_), .B(new_n12773_), .ZN(new_n12774_));
  AOI21_X1   g12582(.A1(new_n12774_), .A2(new_n11373_), .B(new_n12762_), .ZN(new_n12775_));
  NAND2_X1   g12583(.A1(new_n12772_), .A2(new_n12763_), .ZN(new_n12776_));
  AOI21_X1   g12584(.A1(new_n12776_), .A2(new_n12753_), .B(new_n11373_), .ZN(new_n12777_));
  OAI21_X1   g12585(.A1(new_n12775_), .A2(new_n12777_), .B(\asqrt[18] ), .ZN(new_n12778_));
  AOI21_X1   g12586(.A1(new_n12761_), .A2(new_n12778_), .B(new_n10497_), .ZN(new_n12779_));
  NOR3_X1    g12587(.A1(new_n12760_), .A2(\asqrt[20] ), .A3(new_n12779_), .ZN(new_n12780_));
  OAI21_X1   g12588(.A1(new_n12760_), .A2(new_n12779_), .B(\asqrt[20] ), .ZN(new_n12781_));
  OAI21_X1   g12589(.A1(new_n12705_), .A2(new_n12780_), .B(new_n12781_), .ZN(new_n12782_));
  OAI21_X1   g12590(.A1(new_n12782_), .A2(\asqrt[21] ), .B(new_n12702_), .ZN(new_n12783_));
  NAND2_X1   g12591(.A1(new_n12782_), .A2(\asqrt[21] ), .ZN(new_n12784_));
  NAND3_X1   g12592(.A1(new_n12783_), .A2(new_n12784_), .A3(new_n9233_), .ZN(new_n12785_));
  AOI21_X1   g12593(.A1(new_n12783_), .A2(new_n12784_), .B(new_n9233_), .ZN(new_n12786_));
  AOI21_X1   g12594(.A1(new_n12699_), .A2(new_n12785_), .B(new_n12786_), .ZN(new_n12787_));
  AOI21_X1   g12595(.A1(new_n12787_), .A2(new_n8849_), .B(new_n12696_), .ZN(new_n12788_));
  NAND2_X1   g12596(.A1(new_n12785_), .A2(new_n12699_), .ZN(new_n12789_));
  INV_X1     g12597(.I(new_n12702_), .ZN(new_n12790_));
  INV_X1     g12598(.I(new_n12710_), .ZN(new_n12791_));
  NOR3_X1    g12599(.A1(new_n12775_), .A2(\asqrt[18] ), .A3(new_n12777_), .ZN(new_n12792_));
  OAI21_X1   g12600(.A1(new_n12791_), .A2(new_n12792_), .B(new_n12778_), .ZN(new_n12793_));
  OAI21_X1   g12601(.A1(new_n12793_), .A2(\asqrt[19] ), .B(new_n12707_), .ZN(new_n12794_));
  NAND2_X1   g12602(.A1(new_n12793_), .A2(\asqrt[19] ), .ZN(new_n12795_));
  NAND3_X1   g12603(.A1(new_n12794_), .A2(new_n12795_), .A3(new_n10052_), .ZN(new_n12796_));
  AOI21_X1   g12604(.A1(new_n12794_), .A2(new_n12795_), .B(new_n10052_), .ZN(new_n12797_));
  AOI21_X1   g12605(.A1(new_n12704_), .A2(new_n12796_), .B(new_n12797_), .ZN(new_n12798_));
  AOI21_X1   g12606(.A1(new_n12798_), .A2(new_n9656_), .B(new_n12790_), .ZN(new_n12799_));
  NAND2_X1   g12607(.A1(new_n12796_), .A2(new_n12704_), .ZN(new_n12800_));
  AOI21_X1   g12608(.A1(new_n12800_), .A2(new_n12781_), .B(new_n9656_), .ZN(new_n12801_));
  OAI21_X1   g12609(.A1(new_n12799_), .A2(new_n12801_), .B(\asqrt[22] ), .ZN(new_n12802_));
  AOI21_X1   g12610(.A1(new_n12789_), .A2(new_n12802_), .B(new_n8849_), .ZN(new_n12803_));
  NOR3_X1    g12611(.A1(new_n12788_), .A2(\asqrt[24] ), .A3(new_n12803_), .ZN(new_n12804_));
  OAI21_X1   g12612(.A1(new_n12788_), .A2(new_n12803_), .B(\asqrt[24] ), .ZN(new_n12805_));
  OAI21_X1   g12613(.A1(new_n12693_), .A2(new_n12804_), .B(new_n12805_), .ZN(new_n12806_));
  OAI21_X1   g12614(.A1(new_n12806_), .A2(\asqrt[25] ), .B(new_n12690_), .ZN(new_n12807_));
  NAND2_X1   g12615(.A1(new_n12806_), .A2(\asqrt[25] ), .ZN(new_n12808_));
  NAND3_X1   g12616(.A1(new_n12807_), .A2(new_n12808_), .A3(new_n7690_), .ZN(new_n12809_));
  AOI21_X1   g12617(.A1(new_n12807_), .A2(new_n12808_), .B(new_n7690_), .ZN(new_n12810_));
  AOI21_X1   g12618(.A1(new_n12687_), .A2(new_n12809_), .B(new_n12810_), .ZN(new_n12811_));
  AOI21_X1   g12619(.A1(new_n12811_), .A2(new_n7331_), .B(new_n12684_), .ZN(new_n12812_));
  NAND2_X1   g12620(.A1(new_n12809_), .A2(new_n12687_), .ZN(new_n12813_));
  INV_X1     g12621(.I(new_n12690_), .ZN(new_n12814_));
  INV_X1     g12622(.I(new_n12699_), .ZN(new_n12815_));
  NOR3_X1    g12623(.A1(new_n12799_), .A2(\asqrt[22] ), .A3(new_n12801_), .ZN(new_n12816_));
  OAI21_X1   g12624(.A1(new_n12815_), .A2(new_n12816_), .B(new_n12802_), .ZN(new_n12817_));
  OAI21_X1   g12625(.A1(new_n12817_), .A2(\asqrt[23] ), .B(new_n12695_), .ZN(new_n12818_));
  NAND2_X1   g12626(.A1(new_n12817_), .A2(\asqrt[23] ), .ZN(new_n12819_));
  NAND3_X1   g12627(.A1(new_n12818_), .A2(new_n12819_), .A3(new_n8440_), .ZN(new_n12820_));
  AOI21_X1   g12628(.A1(new_n12818_), .A2(new_n12819_), .B(new_n8440_), .ZN(new_n12821_));
  AOI21_X1   g12629(.A1(new_n12692_), .A2(new_n12820_), .B(new_n12821_), .ZN(new_n12822_));
  AOI21_X1   g12630(.A1(new_n12822_), .A2(new_n8077_), .B(new_n12814_), .ZN(new_n12823_));
  NAND2_X1   g12631(.A1(new_n12820_), .A2(new_n12692_), .ZN(new_n12824_));
  AOI21_X1   g12632(.A1(new_n12824_), .A2(new_n12805_), .B(new_n8077_), .ZN(new_n12825_));
  OAI21_X1   g12633(.A1(new_n12823_), .A2(new_n12825_), .B(\asqrt[26] ), .ZN(new_n12826_));
  AOI21_X1   g12634(.A1(new_n12813_), .A2(new_n12826_), .B(new_n7331_), .ZN(new_n12827_));
  NOR3_X1    g12635(.A1(new_n12812_), .A2(\asqrt[28] ), .A3(new_n12827_), .ZN(new_n12828_));
  OAI21_X1   g12636(.A1(new_n12812_), .A2(new_n12827_), .B(\asqrt[28] ), .ZN(new_n12829_));
  OAI21_X1   g12637(.A1(new_n12681_), .A2(new_n12828_), .B(new_n12829_), .ZN(new_n12830_));
  OAI21_X1   g12638(.A1(new_n12830_), .A2(\asqrt[29] ), .B(new_n12678_), .ZN(new_n12831_));
  NAND2_X1   g12639(.A1(new_n12830_), .A2(\asqrt[29] ), .ZN(new_n12832_));
  NAND3_X1   g12640(.A1(new_n12831_), .A2(new_n12832_), .A3(new_n6275_), .ZN(new_n12833_));
  AOI21_X1   g12641(.A1(new_n12831_), .A2(new_n12832_), .B(new_n6275_), .ZN(new_n12834_));
  AOI21_X1   g12642(.A1(new_n12675_), .A2(new_n12833_), .B(new_n12834_), .ZN(new_n12835_));
  AOI21_X1   g12643(.A1(new_n12835_), .A2(new_n5947_), .B(new_n12672_), .ZN(new_n12836_));
  NAND2_X1   g12644(.A1(new_n12833_), .A2(new_n12675_), .ZN(new_n12837_));
  INV_X1     g12645(.I(new_n12678_), .ZN(new_n12838_));
  INV_X1     g12646(.I(new_n12687_), .ZN(new_n12839_));
  NOR3_X1    g12647(.A1(new_n12823_), .A2(\asqrt[26] ), .A3(new_n12825_), .ZN(new_n12840_));
  OAI21_X1   g12648(.A1(new_n12839_), .A2(new_n12840_), .B(new_n12826_), .ZN(new_n12841_));
  OAI21_X1   g12649(.A1(new_n12841_), .A2(\asqrt[27] ), .B(new_n12683_), .ZN(new_n12842_));
  NAND2_X1   g12650(.A1(new_n12841_), .A2(\asqrt[27] ), .ZN(new_n12843_));
  NAND3_X1   g12651(.A1(new_n12842_), .A2(new_n12843_), .A3(new_n6966_), .ZN(new_n12844_));
  AOI21_X1   g12652(.A1(new_n12842_), .A2(new_n12843_), .B(new_n6966_), .ZN(new_n12845_));
  AOI21_X1   g12653(.A1(new_n12680_), .A2(new_n12844_), .B(new_n12845_), .ZN(new_n12846_));
  AOI21_X1   g12654(.A1(new_n12846_), .A2(new_n6636_), .B(new_n12838_), .ZN(new_n12847_));
  NAND2_X1   g12655(.A1(new_n12844_), .A2(new_n12680_), .ZN(new_n12848_));
  AOI21_X1   g12656(.A1(new_n12848_), .A2(new_n12829_), .B(new_n6636_), .ZN(new_n12849_));
  OAI21_X1   g12657(.A1(new_n12847_), .A2(new_n12849_), .B(\asqrt[30] ), .ZN(new_n12850_));
  AOI21_X1   g12658(.A1(new_n12837_), .A2(new_n12850_), .B(new_n5947_), .ZN(new_n12851_));
  NOR3_X1    g12659(.A1(new_n12836_), .A2(\asqrt[32] ), .A3(new_n12851_), .ZN(new_n12852_));
  OAI21_X1   g12660(.A1(new_n12836_), .A2(new_n12851_), .B(\asqrt[32] ), .ZN(new_n12853_));
  OAI21_X1   g12661(.A1(new_n12669_), .A2(new_n12852_), .B(new_n12853_), .ZN(new_n12854_));
  OAI21_X1   g12662(.A1(new_n12854_), .A2(\asqrt[33] ), .B(new_n12666_), .ZN(new_n12855_));
  NAND2_X1   g12663(.A1(new_n12854_), .A2(\asqrt[33] ), .ZN(new_n12856_));
  NAND3_X1   g12664(.A1(new_n12855_), .A2(new_n12856_), .A3(new_n5029_), .ZN(new_n12857_));
  AOI21_X1   g12665(.A1(new_n12855_), .A2(new_n12856_), .B(new_n5029_), .ZN(new_n12858_));
  AOI21_X1   g12666(.A1(new_n12663_), .A2(new_n12857_), .B(new_n12858_), .ZN(new_n12859_));
  AOI21_X1   g12667(.A1(new_n12859_), .A2(new_n4751_), .B(new_n12660_), .ZN(new_n12860_));
  NAND2_X1   g12668(.A1(new_n12857_), .A2(new_n12663_), .ZN(new_n12861_));
  INV_X1     g12669(.I(new_n12666_), .ZN(new_n12862_));
  INV_X1     g12670(.I(new_n12675_), .ZN(new_n12863_));
  NOR3_X1    g12671(.A1(new_n12847_), .A2(\asqrt[30] ), .A3(new_n12849_), .ZN(new_n12864_));
  OAI21_X1   g12672(.A1(new_n12863_), .A2(new_n12864_), .B(new_n12850_), .ZN(new_n12865_));
  OAI21_X1   g12673(.A1(new_n12865_), .A2(\asqrt[31] ), .B(new_n12671_), .ZN(new_n12866_));
  NAND2_X1   g12674(.A1(new_n12865_), .A2(\asqrt[31] ), .ZN(new_n12867_));
  NAND3_X1   g12675(.A1(new_n12866_), .A2(new_n12867_), .A3(new_n5643_), .ZN(new_n12868_));
  AOI21_X1   g12676(.A1(new_n12866_), .A2(new_n12867_), .B(new_n5643_), .ZN(new_n12869_));
  AOI21_X1   g12677(.A1(new_n12668_), .A2(new_n12868_), .B(new_n12869_), .ZN(new_n12870_));
  AOI21_X1   g12678(.A1(new_n12870_), .A2(new_n5336_), .B(new_n12862_), .ZN(new_n12871_));
  NAND2_X1   g12679(.A1(new_n12868_), .A2(new_n12668_), .ZN(new_n12872_));
  AOI21_X1   g12680(.A1(new_n12872_), .A2(new_n12853_), .B(new_n5336_), .ZN(new_n12873_));
  OAI21_X1   g12681(.A1(new_n12871_), .A2(new_n12873_), .B(\asqrt[34] ), .ZN(new_n12874_));
  AOI21_X1   g12682(.A1(new_n12861_), .A2(new_n12874_), .B(new_n4751_), .ZN(new_n12875_));
  NOR3_X1    g12683(.A1(new_n12860_), .A2(\asqrt[36] ), .A3(new_n12875_), .ZN(new_n12876_));
  OAI21_X1   g12684(.A1(new_n12860_), .A2(new_n12875_), .B(\asqrt[36] ), .ZN(new_n12877_));
  OAI21_X1   g12685(.A1(new_n12657_), .A2(new_n12876_), .B(new_n12877_), .ZN(new_n12878_));
  OAI21_X1   g12686(.A1(new_n12878_), .A2(\asqrt[37] ), .B(new_n12654_), .ZN(new_n12879_));
  NAND2_X1   g12687(.A1(new_n12878_), .A2(\asqrt[37] ), .ZN(new_n12880_));
  NAND3_X1   g12688(.A1(new_n12879_), .A2(new_n12880_), .A3(new_n3925_), .ZN(new_n12881_));
  AOI21_X1   g12689(.A1(new_n12879_), .A2(new_n12880_), .B(new_n3925_), .ZN(new_n12882_));
  AOI21_X1   g12690(.A1(new_n12651_), .A2(new_n12881_), .B(new_n12882_), .ZN(new_n12883_));
  AOI21_X1   g12691(.A1(new_n12883_), .A2(new_n3681_), .B(new_n12648_), .ZN(new_n12884_));
  NAND2_X1   g12692(.A1(new_n12881_), .A2(new_n12651_), .ZN(new_n12885_));
  INV_X1     g12693(.I(new_n12654_), .ZN(new_n12886_));
  INV_X1     g12694(.I(new_n12663_), .ZN(new_n12887_));
  NOR3_X1    g12695(.A1(new_n12871_), .A2(\asqrt[34] ), .A3(new_n12873_), .ZN(new_n12888_));
  OAI21_X1   g12696(.A1(new_n12887_), .A2(new_n12888_), .B(new_n12874_), .ZN(new_n12889_));
  OAI21_X1   g12697(.A1(new_n12889_), .A2(\asqrt[35] ), .B(new_n12659_), .ZN(new_n12890_));
  NAND2_X1   g12698(.A1(new_n12889_), .A2(\asqrt[35] ), .ZN(new_n12891_));
  NAND3_X1   g12699(.A1(new_n12890_), .A2(new_n12891_), .A3(new_n4461_), .ZN(new_n12892_));
  AOI21_X1   g12700(.A1(new_n12890_), .A2(new_n12891_), .B(new_n4461_), .ZN(new_n12893_));
  AOI21_X1   g12701(.A1(new_n12656_), .A2(new_n12892_), .B(new_n12893_), .ZN(new_n12894_));
  AOI21_X1   g12702(.A1(new_n12894_), .A2(new_n4196_), .B(new_n12886_), .ZN(new_n12895_));
  NAND2_X1   g12703(.A1(new_n12892_), .A2(new_n12656_), .ZN(new_n12896_));
  AOI21_X1   g12704(.A1(new_n12896_), .A2(new_n12877_), .B(new_n4196_), .ZN(new_n12897_));
  OAI21_X1   g12705(.A1(new_n12895_), .A2(new_n12897_), .B(\asqrt[38] ), .ZN(new_n12898_));
  AOI21_X1   g12706(.A1(new_n12885_), .A2(new_n12898_), .B(new_n3681_), .ZN(new_n12899_));
  NOR3_X1    g12707(.A1(new_n12884_), .A2(\asqrt[40] ), .A3(new_n12899_), .ZN(new_n12900_));
  OAI21_X1   g12708(.A1(new_n12884_), .A2(new_n12899_), .B(\asqrt[40] ), .ZN(new_n12901_));
  OAI21_X1   g12709(.A1(new_n12645_), .A2(new_n12900_), .B(new_n12901_), .ZN(new_n12902_));
  OAI21_X1   g12710(.A1(new_n12902_), .A2(\asqrt[41] ), .B(new_n12642_), .ZN(new_n12903_));
  NAND2_X1   g12711(.A1(new_n12902_), .A2(\asqrt[41] ), .ZN(new_n12904_));
  NAND3_X1   g12712(.A1(new_n12903_), .A2(new_n12904_), .A3(new_n2960_), .ZN(new_n12905_));
  AOI21_X1   g12713(.A1(new_n12903_), .A2(new_n12904_), .B(new_n2960_), .ZN(new_n12906_));
  AOI21_X1   g12714(.A1(new_n12639_), .A2(new_n12905_), .B(new_n12906_), .ZN(new_n12907_));
  AOI21_X1   g12715(.A1(new_n12907_), .A2(new_n2749_), .B(new_n12636_), .ZN(new_n12908_));
  NAND2_X1   g12716(.A1(new_n12905_), .A2(new_n12639_), .ZN(new_n12909_));
  INV_X1     g12717(.I(new_n12642_), .ZN(new_n12910_));
  INV_X1     g12718(.I(new_n12651_), .ZN(new_n12911_));
  NOR3_X1    g12719(.A1(new_n12895_), .A2(\asqrt[38] ), .A3(new_n12897_), .ZN(new_n12912_));
  OAI21_X1   g12720(.A1(new_n12911_), .A2(new_n12912_), .B(new_n12898_), .ZN(new_n12913_));
  OAI21_X1   g12721(.A1(new_n12913_), .A2(\asqrt[39] ), .B(new_n12647_), .ZN(new_n12914_));
  NAND2_X1   g12722(.A1(new_n12913_), .A2(\asqrt[39] ), .ZN(new_n12915_));
  NAND3_X1   g12723(.A1(new_n12914_), .A2(new_n12915_), .A3(new_n3427_), .ZN(new_n12916_));
  AOI21_X1   g12724(.A1(new_n12914_), .A2(new_n12915_), .B(new_n3427_), .ZN(new_n12917_));
  AOI21_X1   g12725(.A1(new_n12644_), .A2(new_n12916_), .B(new_n12917_), .ZN(new_n12918_));
  AOI21_X1   g12726(.A1(new_n12918_), .A2(new_n3195_), .B(new_n12910_), .ZN(new_n12919_));
  NAND2_X1   g12727(.A1(new_n12916_), .A2(new_n12644_), .ZN(new_n12920_));
  AOI21_X1   g12728(.A1(new_n12920_), .A2(new_n12901_), .B(new_n3195_), .ZN(new_n12921_));
  OAI21_X1   g12729(.A1(new_n12919_), .A2(new_n12921_), .B(\asqrt[42] ), .ZN(new_n12922_));
  AOI21_X1   g12730(.A1(new_n12909_), .A2(new_n12922_), .B(new_n2749_), .ZN(new_n12923_));
  NOR3_X1    g12731(.A1(new_n12908_), .A2(\asqrt[44] ), .A3(new_n12923_), .ZN(new_n12924_));
  OAI21_X1   g12732(.A1(new_n12908_), .A2(new_n12923_), .B(\asqrt[44] ), .ZN(new_n12925_));
  OAI21_X1   g12733(.A1(new_n12633_), .A2(new_n12924_), .B(new_n12925_), .ZN(new_n12926_));
  OAI21_X1   g12734(.A1(new_n12926_), .A2(\asqrt[45] ), .B(new_n12630_), .ZN(new_n12927_));
  NAND2_X1   g12735(.A1(new_n12926_), .A2(\asqrt[45] ), .ZN(new_n12928_));
  NAND3_X1   g12736(.A1(new_n12927_), .A2(new_n12928_), .A3(new_n2134_), .ZN(new_n12929_));
  AOI21_X1   g12737(.A1(new_n12927_), .A2(new_n12928_), .B(new_n2134_), .ZN(new_n12930_));
  AOI21_X1   g12738(.A1(new_n12627_), .A2(new_n12929_), .B(new_n12930_), .ZN(new_n12931_));
  AOI21_X1   g12739(.A1(new_n12931_), .A2(new_n1953_), .B(new_n12624_), .ZN(new_n12932_));
  NAND2_X1   g12740(.A1(new_n12929_), .A2(new_n12627_), .ZN(new_n12933_));
  INV_X1     g12741(.I(new_n12630_), .ZN(new_n12934_));
  INV_X1     g12742(.I(new_n12639_), .ZN(new_n12935_));
  NOR3_X1    g12743(.A1(new_n12919_), .A2(\asqrt[42] ), .A3(new_n12921_), .ZN(new_n12936_));
  OAI21_X1   g12744(.A1(new_n12935_), .A2(new_n12936_), .B(new_n12922_), .ZN(new_n12937_));
  OAI21_X1   g12745(.A1(new_n12937_), .A2(\asqrt[43] ), .B(new_n12635_), .ZN(new_n12938_));
  NAND2_X1   g12746(.A1(new_n12937_), .A2(\asqrt[43] ), .ZN(new_n12939_));
  NAND3_X1   g12747(.A1(new_n12938_), .A2(new_n12939_), .A3(new_n2531_), .ZN(new_n12940_));
  AOI21_X1   g12748(.A1(new_n12938_), .A2(new_n12939_), .B(new_n2531_), .ZN(new_n12941_));
  AOI21_X1   g12749(.A1(new_n12632_), .A2(new_n12940_), .B(new_n12941_), .ZN(new_n12942_));
  AOI21_X1   g12750(.A1(new_n12942_), .A2(new_n2332_), .B(new_n12934_), .ZN(new_n12943_));
  NAND2_X1   g12751(.A1(new_n12940_), .A2(new_n12632_), .ZN(new_n12944_));
  AOI21_X1   g12752(.A1(new_n12944_), .A2(new_n12925_), .B(new_n2332_), .ZN(new_n12945_));
  OAI21_X1   g12753(.A1(new_n12943_), .A2(new_n12945_), .B(\asqrt[46] ), .ZN(new_n12946_));
  AOI21_X1   g12754(.A1(new_n12933_), .A2(new_n12946_), .B(new_n1953_), .ZN(new_n12947_));
  NOR3_X1    g12755(.A1(new_n12932_), .A2(\asqrt[48] ), .A3(new_n12947_), .ZN(new_n12948_));
  OAI21_X1   g12756(.A1(new_n12932_), .A2(new_n12947_), .B(\asqrt[48] ), .ZN(new_n12949_));
  OAI21_X1   g12757(.A1(new_n12621_), .A2(new_n12948_), .B(new_n12949_), .ZN(new_n12950_));
  OAI21_X1   g12758(.A1(new_n12950_), .A2(\asqrt[49] ), .B(new_n12618_), .ZN(new_n12951_));
  NAND2_X1   g12759(.A1(new_n12950_), .A2(\asqrt[49] ), .ZN(new_n12952_));
  NAND3_X1   g12760(.A1(new_n12951_), .A2(new_n12952_), .A3(new_n1463_), .ZN(new_n12953_));
  AOI21_X1   g12761(.A1(new_n12951_), .A2(new_n12952_), .B(new_n1463_), .ZN(new_n12954_));
  AOI21_X1   g12762(.A1(new_n12615_), .A2(new_n12953_), .B(new_n12954_), .ZN(new_n12955_));
  NAND2_X1   g12763(.A1(new_n12955_), .A2(new_n1305_), .ZN(new_n12956_));
  INV_X1     g12764(.I(new_n12615_), .ZN(new_n12957_));
  INV_X1     g12765(.I(new_n12618_), .ZN(new_n12958_));
  INV_X1     g12766(.I(new_n12627_), .ZN(new_n12959_));
  NOR3_X1    g12767(.A1(new_n12943_), .A2(\asqrt[46] ), .A3(new_n12945_), .ZN(new_n12960_));
  OAI21_X1   g12768(.A1(new_n12959_), .A2(new_n12960_), .B(new_n12946_), .ZN(new_n12961_));
  OAI21_X1   g12769(.A1(new_n12961_), .A2(\asqrt[47] ), .B(new_n12623_), .ZN(new_n12962_));
  NAND2_X1   g12770(.A1(new_n12961_), .A2(\asqrt[47] ), .ZN(new_n12963_));
  NAND3_X1   g12771(.A1(new_n12962_), .A2(new_n12963_), .A3(new_n1778_), .ZN(new_n12964_));
  AOI21_X1   g12772(.A1(new_n12962_), .A2(new_n12963_), .B(new_n1778_), .ZN(new_n12965_));
  AOI21_X1   g12773(.A1(new_n12620_), .A2(new_n12964_), .B(new_n12965_), .ZN(new_n12966_));
  AOI21_X1   g12774(.A1(new_n12966_), .A2(new_n1632_), .B(new_n12958_), .ZN(new_n12967_));
  NAND2_X1   g12775(.A1(new_n12964_), .A2(new_n12620_), .ZN(new_n12968_));
  AOI21_X1   g12776(.A1(new_n12968_), .A2(new_n12949_), .B(new_n1632_), .ZN(new_n12969_));
  NOR3_X1    g12777(.A1(new_n12967_), .A2(\asqrt[50] ), .A3(new_n12969_), .ZN(new_n12970_));
  OAI21_X1   g12778(.A1(new_n12967_), .A2(new_n12969_), .B(\asqrt[50] ), .ZN(new_n12971_));
  OAI21_X1   g12779(.A1(new_n12957_), .A2(new_n12970_), .B(new_n12971_), .ZN(new_n12972_));
  NAND2_X1   g12780(.A1(new_n12972_), .A2(\asqrt[51] ), .ZN(new_n12973_));
  NOR2_X1    g12781(.A1(new_n12567_), .A2(\asqrt[62] ), .ZN(new_n12974_));
  NOR2_X1    g12782(.A1(new_n12974_), .A2(new_n12724_), .ZN(new_n12975_));
  XOR2_X1    g12783(.A1(new_n12591_), .A2(new_n12131_), .Z(new_n12976_));
  OAI21_X1   g12784(.A1(\asqrt[14] ), .A2(new_n12975_), .B(new_n12976_), .ZN(new_n12977_));
  INV_X1     g12785(.I(new_n12977_), .ZN(new_n12978_));
  AOI21_X1   g12786(.A1(new_n12575_), .A2(new_n12580_), .B(\asqrt[14] ), .ZN(new_n12979_));
  XOR2_X1    g12787(.A1(new_n12979_), .A2(new_n12492_), .Z(new_n12980_));
  INV_X1     g12788(.I(new_n12980_), .ZN(new_n12981_));
  AOI21_X1   g12789(.A1(new_n12555_), .A2(new_n12574_), .B(\asqrt[14] ), .ZN(new_n12982_));
  XOR2_X1    g12790(.A1(new_n12982_), .A2(new_n12496_), .Z(new_n12983_));
  INV_X1     g12791(.I(new_n12983_), .ZN(new_n12984_));
  NOR2_X1    g12792(.A1(new_n12573_), .A2(new_n12569_), .ZN(new_n12985_));
  NOR2_X1    g12793(.A1(\asqrt[14] ), .A2(new_n12985_), .ZN(new_n12986_));
  XOR2_X1    g12794(.A1(new_n12986_), .A2(new_n12498_), .Z(new_n12987_));
  NOR2_X1    g12795(.A1(new_n12544_), .A2(new_n12553_), .ZN(new_n12988_));
  NOR2_X1    g12796(.A1(\asqrt[14] ), .A2(new_n12988_), .ZN(new_n12989_));
  XOR2_X1    g12797(.A1(new_n12989_), .A2(new_n12501_), .Z(new_n12990_));
  AOI21_X1   g12798(.A1(new_n12548_), .A2(new_n12552_), .B(\asqrt[14] ), .ZN(new_n12991_));
  XOR2_X1    g12799(.A1(new_n12991_), .A2(new_n12504_), .Z(new_n12992_));
  INV_X1     g12800(.I(new_n12992_), .ZN(new_n12993_));
  AOI21_X1   g12801(.A1(new_n12534_), .A2(new_n12542_), .B(\asqrt[14] ), .ZN(new_n12994_));
  XOR2_X1    g12802(.A1(new_n12994_), .A2(new_n12508_), .Z(new_n12995_));
  INV_X1     g12803(.I(new_n12995_), .ZN(new_n12996_));
  XOR2_X1    g12804(.A1(new_n12525_), .A2(\asqrt[53] ), .Z(new_n12997_));
  NOR2_X1    g12805(.A1(\asqrt[14] ), .A2(new_n12997_), .ZN(new_n12998_));
  XOR2_X1    g12806(.A1(new_n12998_), .A2(new_n12510_), .Z(new_n12999_));
  NOR2_X1    g12807(.A1(new_n12523_), .A2(new_n12532_), .ZN(new_n13000_));
  NOR2_X1    g12808(.A1(\asqrt[14] ), .A2(new_n13000_), .ZN(new_n13001_));
  XOR2_X1    g12809(.A1(new_n13001_), .A2(new_n12513_), .Z(new_n13002_));
  AOI21_X1   g12810(.A1(new_n12527_), .A2(new_n12531_), .B(\asqrt[14] ), .ZN(new_n13003_));
  XOR2_X1    g12811(.A1(new_n13003_), .A2(new_n12516_), .Z(new_n13004_));
  INV_X1     g12812(.I(new_n13004_), .ZN(new_n13005_));
  INV_X1     g12813(.I(new_n12612_), .ZN(new_n13006_));
  AOI21_X1   g12814(.A1(new_n12955_), .A2(new_n1305_), .B(new_n13006_), .ZN(new_n13007_));
  NAND2_X1   g12815(.A1(new_n12953_), .A2(new_n12615_), .ZN(new_n13008_));
  AOI21_X1   g12816(.A1(new_n13008_), .A2(new_n12971_), .B(new_n1305_), .ZN(new_n13009_));
  NOR3_X1    g12817(.A1(new_n13007_), .A2(\asqrt[52] ), .A3(new_n13009_), .ZN(new_n13010_));
  OAI21_X1   g12818(.A1(new_n13007_), .A2(new_n13009_), .B(\asqrt[52] ), .ZN(new_n13011_));
  OAI21_X1   g12819(.A1(new_n13005_), .A2(new_n13010_), .B(new_n13011_), .ZN(new_n13012_));
  OAI21_X1   g12820(.A1(new_n13012_), .A2(\asqrt[53] ), .B(new_n13002_), .ZN(new_n13013_));
  NAND2_X1   g12821(.A1(new_n13012_), .A2(\asqrt[53] ), .ZN(new_n13014_));
  NAND3_X1   g12822(.A1(new_n13013_), .A2(new_n13014_), .A3(new_n860_), .ZN(new_n13015_));
  AOI21_X1   g12823(.A1(new_n13013_), .A2(new_n13014_), .B(new_n860_), .ZN(new_n13016_));
  AOI21_X1   g12824(.A1(new_n12999_), .A2(new_n13015_), .B(new_n13016_), .ZN(new_n13017_));
  AOI21_X1   g12825(.A1(new_n13017_), .A2(new_n744_), .B(new_n12996_), .ZN(new_n13018_));
  NAND2_X1   g12826(.A1(new_n13015_), .A2(new_n12999_), .ZN(new_n13019_));
  INV_X1     g12827(.I(new_n13002_), .ZN(new_n13020_));
  OAI21_X1   g12828(.A1(new_n12972_), .A2(\asqrt[51] ), .B(new_n12612_), .ZN(new_n13021_));
  NAND3_X1   g12829(.A1(new_n13021_), .A2(new_n12973_), .A3(new_n1150_), .ZN(new_n13022_));
  AOI21_X1   g12830(.A1(new_n13021_), .A2(new_n12973_), .B(new_n1150_), .ZN(new_n13023_));
  AOI21_X1   g12831(.A1(new_n13004_), .A2(new_n13022_), .B(new_n13023_), .ZN(new_n13024_));
  AOI21_X1   g12832(.A1(new_n13024_), .A2(new_n1006_), .B(new_n13020_), .ZN(new_n13025_));
  NAND2_X1   g12833(.A1(new_n13022_), .A2(new_n13004_), .ZN(new_n13026_));
  AOI21_X1   g12834(.A1(new_n13026_), .A2(new_n13011_), .B(new_n1006_), .ZN(new_n13027_));
  OAI21_X1   g12835(.A1(new_n13025_), .A2(new_n13027_), .B(\asqrt[54] ), .ZN(new_n13028_));
  AOI21_X1   g12836(.A1(new_n13019_), .A2(new_n13028_), .B(new_n744_), .ZN(new_n13029_));
  NOR3_X1    g12837(.A1(new_n13018_), .A2(\asqrt[56] ), .A3(new_n13029_), .ZN(new_n13030_));
  OAI21_X1   g12838(.A1(new_n13018_), .A2(new_n13029_), .B(\asqrt[56] ), .ZN(new_n13031_));
  OAI21_X1   g12839(.A1(new_n12993_), .A2(new_n13030_), .B(new_n13031_), .ZN(new_n13032_));
  OAI21_X1   g12840(.A1(new_n13032_), .A2(\asqrt[57] ), .B(new_n12990_), .ZN(new_n13033_));
  NAND2_X1   g12841(.A1(new_n13032_), .A2(\asqrt[57] ), .ZN(new_n13034_));
  NAND3_X1   g12842(.A1(new_n13033_), .A2(new_n13034_), .A3(new_n423_), .ZN(new_n13035_));
  AOI21_X1   g12843(.A1(new_n13033_), .A2(new_n13034_), .B(new_n423_), .ZN(new_n13036_));
  AOI21_X1   g12844(.A1(new_n12987_), .A2(new_n13035_), .B(new_n13036_), .ZN(new_n13037_));
  AOI21_X1   g12845(.A1(new_n13037_), .A2(new_n337_), .B(new_n12984_), .ZN(new_n13038_));
  NAND2_X1   g12846(.A1(new_n13035_), .A2(new_n12987_), .ZN(new_n13039_));
  INV_X1     g12847(.I(new_n12990_), .ZN(new_n13040_));
  INV_X1     g12848(.I(new_n12999_), .ZN(new_n13041_));
  NOR3_X1    g12849(.A1(new_n13025_), .A2(\asqrt[54] ), .A3(new_n13027_), .ZN(new_n13042_));
  OAI21_X1   g12850(.A1(new_n13041_), .A2(new_n13042_), .B(new_n13028_), .ZN(new_n13043_));
  OAI21_X1   g12851(.A1(new_n13043_), .A2(\asqrt[55] ), .B(new_n12995_), .ZN(new_n13044_));
  NAND2_X1   g12852(.A1(new_n13043_), .A2(\asqrt[55] ), .ZN(new_n13045_));
  NAND3_X1   g12853(.A1(new_n13044_), .A2(new_n13045_), .A3(new_n634_), .ZN(new_n13046_));
  AOI21_X1   g12854(.A1(new_n13044_), .A2(new_n13045_), .B(new_n634_), .ZN(new_n13047_));
  AOI21_X1   g12855(.A1(new_n12992_), .A2(new_n13046_), .B(new_n13047_), .ZN(new_n13048_));
  AOI21_X1   g12856(.A1(new_n13048_), .A2(new_n531_), .B(new_n13040_), .ZN(new_n13049_));
  NAND2_X1   g12857(.A1(new_n13046_), .A2(new_n12992_), .ZN(new_n13050_));
  AOI21_X1   g12858(.A1(new_n13050_), .A2(new_n13031_), .B(new_n531_), .ZN(new_n13051_));
  OAI21_X1   g12859(.A1(new_n13049_), .A2(new_n13051_), .B(\asqrt[58] ), .ZN(new_n13052_));
  AOI21_X1   g12860(.A1(new_n13039_), .A2(new_n13052_), .B(new_n337_), .ZN(new_n13053_));
  NOR3_X1    g12861(.A1(new_n13038_), .A2(\asqrt[60] ), .A3(new_n13053_), .ZN(new_n13054_));
  NOR2_X1    g12862(.A1(new_n13054_), .A2(new_n12981_), .ZN(new_n13055_));
  INV_X1     g12863(.I(new_n12987_), .ZN(new_n13056_));
  NOR3_X1    g12864(.A1(new_n13049_), .A2(\asqrt[58] ), .A3(new_n13051_), .ZN(new_n13057_));
  OAI21_X1   g12865(.A1(new_n13056_), .A2(new_n13057_), .B(new_n13052_), .ZN(new_n13058_));
  OAI21_X1   g12866(.A1(new_n13058_), .A2(\asqrt[59] ), .B(new_n12983_), .ZN(new_n13059_));
  NOR2_X1    g12867(.A1(new_n13057_), .A2(new_n13056_), .ZN(new_n13060_));
  OAI21_X1   g12868(.A1(new_n13060_), .A2(new_n13036_), .B(\asqrt[59] ), .ZN(new_n13061_));
  AOI21_X1   g12869(.A1(new_n13059_), .A2(new_n13061_), .B(new_n266_), .ZN(new_n13062_));
  OAI21_X1   g12870(.A1(new_n13055_), .A2(new_n13062_), .B(\asqrt[61] ), .ZN(new_n13063_));
  OAI21_X1   g12871(.A1(new_n13038_), .A2(new_n13053_), .B(\asqrt[60] ), .ZN(new_n13064_));
  OAI21_X1   g12872(.A1(new_n12981_), .A2(new_n13054_), .B(new_n13064_), .ZN(new_n13065_));
  AOI21_X1   g12873(.A1(new_n12581_), .A2(new_n12561_), .B(\asqrt[14] ), .ZN(new_n13066_));
  XOR2_X1    g12874(.A1(new_n13066_), .A2(new_n12489_), .Z(new_n13067_));
  OAI21_X1   g12875(.A1(new_n13065_), .A2(\asqrt[61] ), .B(new_n13067_), .ZN(new_n13068_));
  NAND2_X1   g12876(.A1(new_n13068_), .A2(new_n13063_), .ZN(new_n13069_));
  NAND3_X1   g12877(.A1(new_n13059_), .A2(new_n266_), .A3(new_n13061_), .ZN(new_n13070_));
  NAND2_X1   g12878(.A1(new_n13070_), .A2(new_n12980_), .ZN(new_n13071_));
  AOI21_X1   g12879(.A1(new_n13071_), .A2(new_n13064_), .B(new_n239_), .ZN(new_n13072_));
  AOI21_X1   g12880(.A1(new_n12980_), .A2(new_n13070_), .B(new_n13062_), .ZN(new_n13073_));
  INV_X1     g12881(.I(new_n13067_), .ZN(new_n13074_));
  AOI21_X1   g12882(.A1(new_n13073_), .A2(new_n239_), .B(new_n13074_), .ZN(new_n13075_));
  OAI21_X1   g12883(.A1(new_n13075_), .A2(new_n13072_), .B(new_n201_), .ZN(new_n13076_));
  NAND3_X1   g12884(.A1(new_n13068_), .A2(\asqrt[62] ), .A3(new_n13063_), .ZN(new_n13077_));
  NAND2_X1   g12885(.A1(new_n12585_), .A2(new_n239_), .ZN(new_n13078_));
  AOI21_X1   g12886(.A1(new_n12563_), .A2(new_n13078_), .B(\asqrt[14] ), .ZN(new_n13079_));
  XOR2_X1    g12887(.A1(new_n13079_), .A2(new_n12565_), .Z(new_n13080_));
  INV_X1     g12888(.I(new_n13080_), .ZN(new_n13081_));
  AOI22_X1   g12889(.A1(new_n13076_), .A2(new_n13077_), .B1(new_n13069_), .B2(new_n13081_), .ZN(new_n13082_));
  NOR2_X1    g12890(.A1(new_n12594_), .A2(new_n12487_), .ZN(new_n13083_));
  OAI21_X1   g12891(.A1(\asqrt[14] ), .A2(new_n13083_), .B(new_n12601_), .ZN(new_n13084_));
  INV_X1     g12892(.I(new_n13084_), .ZN(new_n13085_));
  OAI21_X1   g12893(.A1(new_n13082_), .A2(new_n12978_), .B(new_n13085_), .ZN(new_n13086_));
  OAI21_X1   g12894(.A1(new_n13069_), .A2(\asqrt[62] ), .B(new_n13080_), .ZN(new_n13087_));
  NAND2_X1   g12895(.A1(new_n13069_), .A2(\asqrt[62] ), .ZN(new_n13088_));
  NAND3_X1   g12896(.A1(new_n13087_), .A2(new_n13088_), .A3(new_n12978_), .ZN(new_n13089_));
  NAND2_X1   g12897(.A1(new_n12733_), .A2(new_n12486_), .ZN(new_n13090_));
  XOR2_X1    g12898(.A1(new_n12721_), .A2(new_n12486_), .Z(new_n13091_));
  NAND3_X1   g12899(.A1(new_n13090_), .A2(\asqrt[63] ), .A3(new_n13091_), .ZN(new_n13092_));
  INV_X1     g12900(.I(new_n12730_), .ZN(new_n13093_));
  NAND4_X1   g12901(.A1(new_n13093_), .A2(new_n12487_), .A3(new_n12601_), .A4(new_n12609_), .ZN(new_n13094_));
  NAND2_X1   g12902(.A1(new_n13092_), .A2(new_n13094_), .ZN(new_n13095_));
  INV_X1     g12903(.I(new_n13095_), .ZN(new_n13096_));
  NAND4_X1   g12904(.A1(new_n13086_), .A2(new_n193_), .A3(new_n13089_), .A4(new_n13096_), .ZN(\asqrt[13] ));
  AOI21_X1   g12905(.A1(new_n12956_), .A2(new_n12973_), .B(\asqrt[13] ), .ZN(new_n13098_));
  XOR2_X1    g12906(.A1(new_n13098_), .A2(new_n12612_), .Z(new_n13099_));
  AOI21_X1   g12907(.A1(new_n12953_), .A2(new_n12971_), .B(\asqrt[13] ), .ZN(new_n13100_));
  XOR2_X1    g12908(.A1(new_n13100_), .A2(new_n12615_), .Z(new_n13101_));
  NAND2_X1   g12909(.A1(new_n12966_), .A2(new_n1632_), .ZN(new_n13102_));
  AOI21_X1   g12910(.A1(new_n13102_), .A2(new_n12952_), .B(\asqrt[13] ), .ZN(new_n13103_));
  XOR2_X1    g12911(.A1(new_n13103_), .A2(new_n12618_), .Z(new_n13104_));
  INV_X1     g12912(.I(new_n13104_), .ZN(new_n13105_));
  AOI21_X1   g12913(.A1(new_n12964_), .A2(new_n12949_), .B(\asqrt[13] ), .ZN(new_n13106_));
  XOR2_X1    g12914(.A1(new_n13106_), .A2(new_n12620_), .Z(new_n13107_));
  INV_X1     g12915(.I(new_n13107_), .ZN(new_n13108_));
  NAND2_X1   g12916(.A1(new_n12931_), .A2(new_n1953_), .ZN(new_n13109_));
  AOI21_X1   g12917(.A1(new_n13109_), .A2(new_n12963_), .B(\asqrt[13] ), .ZN(new_n13110_));
  XOR2_X1    g12918(.A1(new_n13110_), .A2(new_n12623_), .Z(new_n13111_));
  AOI21_X1   g12919(.A1(new_n12929_), .A2(new_n12946_), .B(\asqrt[13] ), .ZN(new_n13112_));
  XOR2_X1    g12920(.A1(new_n13112_), .A2(new_n12627_), .Z(new_n13113_));
  NAND2_X1   g12921(.A1(new_n12942_), .A2(new_n2332_), .ZN(new_n13114_));
  AOI21_X1   g12922(.A1(new_n13114_), .A2(new_n12928_), .B(\asqrt[13] ), .ZN(new_n13115_));
  XOR2_X1    g12923(.A1(new_n13115_), .A2(new_n12630_), .Z(new_n13116_));
  INV_X1     g12924(.I(new_n13116_), .ZN(new_n13117_));
  AOI21_X1   g12925(.A1(new_n12940_), .A2(new_n12925_), .B(\asqrt[13] ), .ZN(new_n13118_));
  XOR2_X1    g12926(.A1(new_n13118_), .A2(new_n12632_), .Z(new_n13119_));
  INV_X1     g12927(.I(new_n13119_), .ZN(new_n13120_));
  NAND2_X1   g12928(.A1(new_n12907_), .A2(new_n2749_), .ZN(new_n13121_));
  AOI21_X1   g12929(.A1(new_n13121_), .A2(new_n12939_), .B(\asqrt[13] ), .ZN(new_n13122_));
  XOR2_X1    g12930(.A1(new_n13122_), .A2(new_n12635_), .Z(new_n13123_));
  AOI21_X1   g12931(.A1(new_n12905_), .A2(new_n12922_), .B(\asqrt[13] ), .ZN(new_n13124_));
  XOR2_X1    g12932(.A1(new_n13124_), .A2(new_n12639_), .Z(new_n13125_));
  NAND2_X1   g12933(.A1(new_n12918_), .A2(new_n3195_), .ZN(new_n13126_));
  AOI21_X1   g12934(.A1(new_n13126_), .A2(new_n12904_), .B(\asqrt[13] ), .ZN(new_n13127_));
  XOR2_X1    g12935(.A1(new_n13127_), .A2(new_n12642_), .Z(new_n13128_));
  INV_X1     g12936(.I(new_n13128_), .ZN(new_n13129_));
  AOI21_X1   g12937(.A1(new_n12916_), .A2(new_n12901_), .B(\asqrt[13] ), .ZN(new_n13130_));
  XOR2_X1    g12938(.A1(new_n13130_), .A2(new_n12644_), .Z(new_n13131_));
  INV_X1     g12939(.I(new_n13131_), .ZN(new_n13132_));
  NAND2_X1   g12940(.A1(new_n12883_), .A2(new_n3681_), .ZN(new_n13133_));
  AOI21_X1   g12941(.A1(new_n13133_), .A2(new_n12915_), .B(\asqrt[13] ), .ZN(new_n13134_));
  XOR2_X1    g12942(.A1(new_n13134_), .A2(new_n12647_), .Z(new_n13135_));
  AOI21_X1   g12943(.A1(new_n12881_), .A2(new_n12898_), .B(\asqrt[13] ), .ZN(new_n13136_));
  XOR2_X1    g12944(.A1(new_n13136_), .A2(new_n12651_), .Z(new_n13137_));
  NAND2_X1   g12945(.A1(new_n12894_), .A2(new_n4196_), .ZN(new_n13138_));
  AOI21_X1   g12946(.A1(new_n13138_), .A2(new_n12880_), .B(\asqrt[13] ), .ZN(new_n13139_));
  XOR2_X1    g12947(.A1(new_n13139_), .A2(new_n12654_), .Z(new_n13140_));
  INV_X1     g12948(.I(new_n13140_), .ZN(new_n13141_));
  AOI21_X1   g12949(.A1(new_n12892_), .A2(new_n12877_), .B(\asqrt[13] ), .ZN(new_n13142_));
  XOR2_X1    g12950(.A1(new_n13142_), .A2(new_n12656_), .Z(new_n13143_));
  INV_X1     g12951(.I(new_n13143_), .ZN(new_n13144_));
  NAND2_X1   g12952(.A1(new_n12859_), .A2(new_n4751_), .ZN(new_n13145_));
  AOI21_X1   g12953(.A1(new_n13145_), .A2(new_n12891_), .B(\asqrt[13] ), .ZN(new_n13146_));
  XOR2_X1    g12954(.A1(new_n13146_), .A2(new_n12659_), .Z(new_n13147_));
  AOI21_X1   g12955(.A1(new_n12857_), .A2(new_n12874_), .B(\asqrt[13] ), .ZN(new_n13148_));
  XOR2_X1    g12956(.A1(new_n13148_), .A2(new_n12663_), .Z(new_n13149_));
  NAND2_X1   g12957(.A1(new_n12870_), .A2(new_n5336_), .ZN(new_n13150_));
  AOI21_X1   g12958(.A1(new_n13150_), .A2(new_n12856_), .B(\asqrt[13] ), .ZN(new_n13151_));
  XOR2_X1    g12959(.A1(new_n13151_), .A2(new_n12666_), .Z(new_n13152_));
  INV_X1     g12960(.I(new_n13152_), .ZN(new_n13153_));
  AOI21_X1   g12961(.A1(new_n12868_), .A2(new_n12853_), .B(\asqrt[13] ), .ZN(new_n13154_));
  XOR2_X1    g12962(.A1(new_n13154_), .A2(new_n12668_), .Z(new_n13155_));
  INV_X1     g12963(.I(new_n13155_), .ZN(new_n13156_));
  NAND2_X1   g12964(.A1(new_n12835_), .A2(new_n5947_), .ZN(new_n13157_));
  AOI21_X1   g12965(.A1(new_n13157_), .A2(new_n12867_), .B(\asqrt[13] ), .ZN(new_n13158_));
  XOR2_X1    g12966(.A1(new_n13158_), .A2(new_n12671_), .Z(new_n13159_));
  AOI21_X1   g12967(.A1(new_n12833_), .A2(new_n12850_), .B(\asqrt[13] ), .ZN(new_n13160_));
  XOR2_X1    g12968(.A1(new_n13160_), .A2(new_n12675_), .Z(new_n13161_));
  NAND2_X1   g12969(.A1(new_n12846_), .A2(new_n6636_), .ZN(new_n13162_));
  AOI21_X1   g12970(.A1(new_n13162_), .A2(new_n12832_), .B(\asqrt[13] ), .ZN(new_n13163_));
  XOR2_X1    g12971(.A1(new_n13163_), .A2(new_n12678_), .Z(new_n13164_));
  INV_X1     g12972(.I(new_n13164_), .ZN(new_n13165_));
  AOI21_X1   g12973(.A1(new_n12844_), .A2(new_n12829_), .B(\asqrt[13] ), .ZN(new_n13166_));
  XOR2_X1    g12974(.A1(new_n13166_), .A2(new_n12680_), .Z(new_n13167_));
  INV_X1     g12975(.I(new_n13167_), .ZN(new_n13168_));
  NAND2_X1   g12976(.A1(new_n12811_), .A2(new_n7331_), .ZN(new_n13169_));
  AOI21_X1   g12977(.A1(new_n13169_), .A2(new_n12843_), .B(\asqrt[13] ), .ZN(new_n13170_));
  XOR2_X1    g12978(.A1(new_n13170_), .A2(new_n12683_), .Z(new_n13171_));
  AOI21_X1   g12979(.A1(new_n12809_), .A2(new_n12826_), .B(\asqrt[13] ), .ZN(new_n13172_));
  XOR2_X1    g12980(.A1(new_n13172_), .A2(new_n12687_), .Z(new_n13173_));
  NAND2_X1   g12981(.A1(new_n12822_), .A2(new_n8077_), .ZN(new_n13174_));
  AOI21_X1   g12982(.A1(new_n13174_), .A2(new_n12808_), .B(\asqrt[13] ), .ZN(new_n13175_));
  XOR2_X1    g12983(.A1(new_n13175_), .A2(new_n12690_), .Z(new_n13176_));
  INV_X1     g12984(.I(new_n13176_), .ZN(new_n13177_));
  AOI21_X1   g12985(.A1(new_n12820_), .A2(new_n12805_), .B(\asqrt[13] ), .ZN(new_n13178_));
  XOR2_X1    g12986(.A1(new_n13178_), .A2(new_n12692_), .Z(new_n13179_));
  INV_X1     g12987(.I(new_n13179_), .ZN(new_n13180_));
  NAND2_X1   g12988(.A1(new_n12787_), .A2(new_n8849_), .ZN(new_n13181_));
  AOI21_X1   g12989(.A1(new_n13181_), .A2(new_n12819_), .B(\asqrt[13] ), .ZN(new_n13182_));
  XOR2_X1    g12990(.A1(new_n13182_), .A2(new_n12695_), .Z(new_n13183_));
  AOI21_X1   g12991(.A1(new_n12785_), .A2(new_n12802_), .B(\asqrt[13] ), .ZN(new_n13184_));
  XOR2_X1    g12992(.A1(new_n13184_), .A2(new_n12699_), .Z(new_n13185_));
  NAND2_X1   g12993(.A1(new_n12798_), .A2(new_n9656_), .ZN(new_n13186_));
  AOI21_X1   g12994(.A1(new_n13186_), .A2(new_n12784_), .B(\asqrt[13] ), .ZN(new_n13187_));
  XOR2_X1    g12995(.A1(new_n13187_), .A2(new_n12702_), .Z(new_n13188_));
  INV_X1     g12996(.I(new_n13188_), .ZN(new_n13189_));
  AOI21_X1   g12997(.A1(new_n12796_), .A2(new_n12781_), .B(\asqrt[13] ), .ZN(new_n13190_));
  XOR2_X1    g12998(.A1(new_n13190_), .A2(new_n12704_), .Z(new_n13191_));
  INV_X1     g12999(.I(new_n13191_), .ZN(new_n13192_));
  NAND2_X1   g13000(.A1(new_n12759_), .A2(new_n10497_), .ZN(new_n13193_));
  AOI21_X1   g13001(.A1(new_n13193_), .A2(new_n12795_), .B(\asqrt[13] ), .ZN(new_n13194_));
  XOR2_X1    g13002(.A1(new_n13194_), .A2(new_n12707_), .Z(new_n13195_));
  AOI21_X1   g13003(.A1(new_n12757_), .A2(new_n12778_), .B(\asqrt[13] ), .ZN(new_n13196_));
  XOR2_X1    g13004(.A1(new_n13196_), .A2(new_n12710_), .Z(new_n13197_));
  NAND2_X1   g13005(.A1(new_n12774_), .A2(new_n11373_), .ZN(new_n13198_));
  AOI21_X1   g13006(.A1(new_n13198_), .A2(new_n12756_), .B(\asqrt[13] ), .ZN(new_n13199_));
  XOR2_X1    g13007(.A1(new_n13199_), .A2(new_n12717_), .Z(new_n13200_));
  INV_X1     g13008(.I(new_n13200_), .ZN(new_n13201_));
  AOI21_X1   g13009(.A1(new_n12772_), .A2(new_n12753_), .B(\asqrt[13] ), .ZN(new_n13202_));
  XOR2_X1    g13010(.A1(new_n13202_), .A2(new_n12763_), .Z(new_n13203_));
  INV_X1     g13011(.I(new_n13203_), .ZN(new_n13204_));
  NAND2_X1   g13012(.A1(\asqrt[14] ), .A2(new_n12740_), .ZN(new_n13205_));
  NOR2_X1    g13013(.A1(new_n12748_), .A2(\a[28] ), .ZN(new_n13206_));
  AOI22_X1   g13014(.A1(new_n13205_), .A2(new_n12748_), .B1(\asqrt[14] ), .B2(new_n13206_), .ZN(new_n13207_));
  OAI21_X1   g13015(.A1(new_n12733_), .A2(new_n12740_), .B(new_n12767_), .ZN(new_n13208_));
  AOI21_X1   g13016(.A1(new_n12766_), .A2(new_n13208_), .B(\asqrt[13] ), .ZN(new_n13209_));
  XOR2_X1    g13017(.A1(new_n13209_), .A2(new_n13207_), .Z(new_n13210_));
  NAND3_X1   g13018(.A1(new_n13071_), .A2(new_n239_), .A3(new_n13064_), .ZN(new_n13211_));
  AOI21_X1   g13019(.A1(new_n13067_), .A2(new_n13211_), .B(new_n13072_), .ZN(new_n13212_));
  AOI21_X1   g13020(.A1(new_n13068_), .A2(new_n13063_), .B(\asqrt[62] ), .ZN(new_n13213_));
  NOR3_X1    g13021(.A1(new_n13075_), .A2(new_n201_), .A3(new_n13072_), .ZN(new_n13214_));
  OAI22_X1   g13022(.A1(new_n13214_), .A2(new_n13213_), .B1(new_n13212_), .B2(new_n13080_), .ZN(new_n13215_));
  AOI21_X1   g13023(.A1(new_n13215_), .A2(new_n12977_), .B(new_n13084_), .ZN(new_n13216_));
  AOI21_X1   g13024(.A1(new_n13212_), .A2(new_n201_), .B(new_n13081_), .ZN(new_n13217_));
  OAI21_X1   g13025(.A1(new_n13212_), .A2(new_n201_), .B(new_n12978_), .ZN(new_n13218_));
  NOR2_X1    g13026(.A1(new_n13217_), .A2(new_n13218_), .ZN(new_n13219_));
  NOR3_X1    g13027(.A1(new_n13216_), .A2(\asqrt[63] ), .A3(new_n13219_), .ZN(new_n13220_));
  NAND3_X1   g13028(.A1(new_n13092_), .A2(\asqrt[14] ), .A3(new_n13094_), .ZN(new_n13221_));
  INV_X1     g13029(.I(new_n13221_), .ZN(new_n13222_));
  NAND2_X1   g13030(.A1(new_n13220_), .A2(new_n13222_), .ZN(new_n13223_));
  NAND2_X1   g13031(.A1(\asqrt[13] ), .A2(new_n12737_), .ZN(new_n13224_));
  AOI21_X1   g13032(.A1(new_n13224_), .A2(new_n13223_), .B(\a[28] ), .ZN(new_n13225_));
  NAND2_X1   g13033(.A1(new_n13086_), .A2(new_n193_), .ZN(new_n13226_));
  NOR3_X1    g13034(.A1(new_n13226_), .A2(new_n13219_), .A3(new_n13221_), .ZN(new_n13227_));
  NOR4_X1    g13035(.A1(new_n13216_), .A2(\asqrt[63] ), .A3(new_n13219_), .A4(new_n13095_), .ZN(new_n13228_));
  NOR2_X1    g13036(.A1(new_n13228_), .A2(new_n12738_), .ZN(new_n13229_));
  NOR3_X1    g13037(.A1(new_n13229_), .A2(new_n13227_), .A3(new_n12740_), .ZN(new_n13230_));
  NOR2_X1    g13038(.A1(new_n13230_), .A2(new_n13225_), .ZN(new_n13231_));
  INV_X1     g13039(.I(\a[26] ), .ZN(new_n13232_));
  NOR2_X1    g13040(.A1(\a[24] ), .A2(\a[25] ), .ZN(new_n13233_));
  NOR3_X1    g13041(.A1(new_n13228_), .A2(new_n13232_), .A3(new_n13233_), .ZN(new_n13234_));
  INV_X1     g13042(.I(new_n13233_), .ZN(new_n13235_));
  AOI21_X1   g13043(.A1(new_n13228_), .A2(\a[26] ), .B(new_n13235_), .ZN(new_n13236_));
  OAI21_X1   g13044(.A1(new_n13234_), .A2(new_n13236_), .B(\asqrt[14] ), .ZN(new_n13237_));
  NAND2_X1   g13045(.A1(new_n13233_), .A2(new_n13232_), .ZN(new_n13238_));
  NAND3_X1   g13046(.A1(new_n12605_), .A2(new_n12607_), .A3(new_n13238_), .ZN(new_n13239_));
  NAND2_X1   g13047(.A1(new_n12726_), .A2(new_n13239_), .ZN(new_n13240_));
  INV_X1     g13048(.I(new_n13240_), .ZN(new_n13241_));
  NOR3_X1    g13049(.A1(new_n13228_), .A2(new_n13232_), .A3(new_n13241_), .ZN(new_n13242_));
  NOR3_X1    g13050(.A1(new_n13228_), .A2(\a[26] ), .A3(\a[27] ), .ZN(new_n13243_));
  INV_X1     g13051(.I(\a[27] ), .ZN(new_n13244_));
  AOI21_X1   g13052(.A1(\asqrt[13] ), .A2(new_n13232_), .B(new_n13244_), .ZN(new_n13245_));
  NOR3_X1    g13053(.A1(new_n13242_), .A2(new_n13243_), .A3(new_n13245_), .ZN(new_n13246_));
  NAND3_X1   g13054(.A1(new_n13246_), .A2(new_n13237_), .A3(new_n12283_), .ZN(new_n13247_));
  NAND2_X1   g13055(.A1(new_n13247_), .A2(new_n13231_), .ZN(new_n13248_));
  NAND3_X1   g13056(.A1(\asqrt[13] ), .A2(\a[26] ), .A3(new_n13235_), .ZN(new_n13249_));
  OAI21_X1   g13057(.A1(\asqrt[13] ), .A2(new_n13232_), .B(new_n13233_), .ZN(new_n13250_));
  AOI21_X1   g13058(.A1(new_n13250_), .A2(new_n13249_), .B(new_n12733_), .ZN(new_n13251_));
  NAND3_X1   g13059(.A1(\asqrt[13] ), .A2(\a[26] ), .A3(new_n13240_), .ZN(new_n13252_));
  NAND3_X1   g13060(.A1(\asqrt[13] ), .A2(new_n13232_), .A3(new_n13244_), .ZN(new_n13253_));
  OAI21_X1   g13061(.A1(new_n13228_), .A2(\a[26] ), .B(\a[27] ), .ZN(new_n13254_));
  NAND3_X1   g13062(.A1(new_n13252_), .A2(new_n13254_), .A3(new_n13253_), .ZN(new_n13255_));
  OAI21_X1   g13063(.A1(new_n13255_), .A2(new_n13251_), .B(\asqrt[15] ), .ZN(new_n13256_));
  NAND3_X1   g13064(.A1(new_n13248_), .A2(new_n11802_), .A3(new_n13256_), .ZN(new_n13257_));
  AOI21_X1   g13065(.A1(new_n13248_), .A2(new_n13256_), .B(new_n11802_), .ZN(new_n13258_));
  AOI21_X1   g13066(.A1(new_n13210_), .A2(new_n13257_), .B(new_n13258_), .ZN(new_n13259_));
  AOI21_X1   g13067(.A1(new_n13259_), .A2(new_n11373_), .B(new_n13204_), .ZN(new_n13260_));
  OR2_X2     g13068(.A1(new_n13230_), .A2(new_n13225_), .Z(new_n13261_));
  NOR3_X1    g13069(.A1(new_n13255_), .A2(new_n13251_), .A3(\asqrt[15] ), .ZN(new_n13262_));
  OAI21_X1   g13070(.A1(new_n13261_), .A2(new_n13262_), .B(new_n13256_), .ZN(new_n13263_));
  OAI21_X1   g13071(.A1(new_n13263_), .A2(\asqrt[16] ), .B(new_n13210_), .ZN(new_n13264_));
  NAND2_X1   g13072(.A1(new_n13263_), .A2(\asqrt[16] ), .ZN(new_n13265_));
  AOI21_X1   g13073(.A1(new_n13264_), .A2(new_n13265_), .B(new_n11373_), .ZN(new_n13266_));
  NOR3_X1    g13074(.A1(new_n13260_), .A2(\asqrt[18] ), .A3(new_n13266_), .ZN(new_n13267_));
  OAI21_X1   g13075(.A1(new_n13260_), .A2(new_n13266_), .B(\asqrt[18] ), .ZN(new_n13268_));
  OAI21_X1   g13076(.A1(new_n13201_), .A2(new_n13267_), .B(new_n13268_), .ZN(new_n13269_));
  OAI21_X1   g13077(.A1(new_n13269_), .A2(\asqrt[19] ), .B(new_n13197_), .ZN(new_n13270_));
  NAND3_X1   g13078(.A1(new_n13264_), .A2(new_n13265_), .A3(new_n11373_), .ZN(new_n13271_));
  AOI21_X1   g13079(.A1(new_n13203_), .A2(new_n13271_), .B(new_n13266_), .ZN(new_n13272_));
  AOI21_X1   g13080(.A1(new_n13272_), .A2(new_n10914_), .B(new_n13201_), .ZN(new_n13273_));
  NAND2_X1   g13081(.A1(new_n13271_), .A2(new_n13203_), .ZN(new_n13274_));
  INV_X1     g13082(.I(new_n13266_), .ZN(new_n13275_));
  AOI21_X1   g13083(.A1(new_n13274_), .A2(new_n13275_), .B(new_n10914_), .ZN(new_n13276_));
  OAI21_X1   g13084(.A1(new_n13273_), .A2(new_n13276_), .B(\asqrt[19] ), .ZN(new_n13277_));
  NAND3_X1   g13085(.A1(new_n13270_), .A2(new_n10052_), .A3(new_n13277_), .ZN(new_n13278_));
  AOI21_X1   g13086(.A1(new_n13270_), .A2(new_n13277_), .B(new_n10052_), .ZN(new_n13279_));
  AOI21_X1   g13087(.A1(new_n13195_), .A2(new_n13278_), .B(new_n13279_), .ZN(new_n13280_));
  AOI21_X1   g13088(.A1(new_n13280_), .A2(new_n9656_), .B(new_n13192_), .ZN(new_n13281_));
  INV_X1     g13089(.I(new_n13197_), .ZN(new_n13282_));
  NOR3_X1    g13090(.A1(new_n13273_), .A2(\asqrt[19] ), .A3(new_n13276_), .ZN(new_n13283_));
  OAI21_X1   g13091(.A1(new_n13282_), .A2(new_n13283_), .B(new_n13277_), .ZN(new_n13284_));
  OAI21_X1   g13092(.A1(new_n13284_), .A2(\asqrt[20] ), .B(new_n13195_), .ZN(new_n13285_));
  NAND2_X1   g13093(.A1(new_n13284_), .A2(\asqrt[20] ), .ZN(new_n13286_));
  AOI21_X1   g13094(.A1(new_n13285_), .A2(new_n13286_), .B(new_n9656_), .ZN(new_n13287_));
  NOR3_X1    g13095(.A1(new_n13281_), .A2(\asqrt[22] ), .A3(new_n13287_), .ZN(new_n13288_));
  OAI21_X1   g13096(.A1(new_n13281_), .A2(new_n13287_), .B(\asqrt[22] ), .ZN(new_n13289_));
  OAI21_X1   g13097(.A1(new_n13189_), .A2(new_n13288_), .B(new_n13289_), .ZN(new_n13290_));
  OAI21_X1   g13098(.A1(new_n13290_), .A2(\asqrt[23] ), .B(new_n13185_), .ZN(new_n13291_));
  NAND3_X1   g13099(.A1(new_n13285_), .A2(new_n13286_), .A3(new_n9656_), .ZN(new_n13292_));
  AOI21_X1   g13100(.A1(new_n13191_), .A2(new_n13292_), .B(new_n13287_), .ZN(new_n13293_));
  AOI21_X1   g13101(.A1(new_n13293_), .A2(new_n9233_), .B(new_n13189_), .ZN(new_n13294_));
  NAND2_X1   g13102(.A1(new_n13292_), .A2(new_n13191_), .ZN(new_n13295_));
  INV_X1     g13103(.I(new_n13287_), .ZN(new_n13296_));
  AOI21_X1   g13104(.A1(new_n13295_), .A2(new_n13296_), .B(new_n9233_), .ZN(new_n13297_));
  OAI21_X1   g13105(.A1(new_n13294_), .A2(new_n13297_), .B(\asqrt[23] ), .ZN(new_n13298_));
  NAND3_X1   g13106(.A1(new_n13291_), .A2(new_n8440_), .A3(new_n13298_), .ZN(new_n13299_));
  AOI21_X1   g13107(.A1(new_n13291_), .A2(new_n13298_), .B(new_n8440_), .ZN(new_n13300_));
  AOI21_X1   g13108(.A1(new_n13183_), .A2(new_n13299_), .B(new_n13300_), .ZN(new_n13301_));
  AOI21_X1   g13109(.A1(new_n13301_), .A2(new_n8077_), .B(new_n13180_), .ZN(new_n13302_));
  INV_X1     g13110(.I(new_n13185_), .ZN(new_n13303_));
  NOR3_X1    g13111(.A1(new_n13294_), .A2(\asqrt[23] ), .A3(new_n13297_), .ZN(new_n13304_));
  OAI21_X1   g13112(.A1(new_n13303_), .A2(new_n13304_), .B(new_n13298_), .ZN(new_n13305_));
  OAI21_X1   g13113(.A1(new_n13305_), .A2(\asqrt[24] ), .B(new_n13183_), .ZN(new_n13306_));
  NAND2_X1   g13114(.A1(new_n13305_), .A2(\asqrt[24] ), .ZN(new_n13307_));
  AOI21_X1   g13115(.A1(new_n13306_), .A2(new_n13307_), .B(new_n8077_), .ZN(new_n13308_));
  NOR3_X1    g13116(.A1(new_n13302_), .A2(\asqrt[26] ), .A3(new_n13308_), .ZN(new_n13309_));
  OAI21_X1   g13117(.A1(new_n13302_), .A2(new_n13308_), .B(\asqrt[26] ), .ZN(new_n13310_));
  OAI21_X1   g13118(.A1(new_n13177_), .A2(new_n13309_), .B(new_n13310_), .ZN(new_n13311_));
  OAI21_X1   g13119(.A1(new_n13311_), .A2(\asqrt[27] ), .B(new_n13173_), .ZN(new_n13312_));
  NAND3_X1   g13120(.A1(new_n13306_), .A2(new_n13307_), .A3(new_n8077_), .ZN(new_n13313_));
  AOI21_X1   g13121(.A1(new_n13179_), .A2(new_n13313_), .B(new_n13308_), .ZN(new_n13314_));
  AOI21_X1   g13122(.A1(new_n13314_), .A2(new_n7690_), .B(new_n13177_), .ZN(new_n13315_));
  NAND2_X1   g13123(.A1(new_n13313_), .A2(new_n13179_), .ZN(new_n13316_));
  INV_X1     g13124(.I(new_n13308_), .ZN(new_n13317_));
  AOI21_X1   g13125(.A1(new_n13316_), .A2(new_n13317_), .B(new_n7690_), .ZN(new_n13318_));
  OAI21_X1   g13126(.A1(new_n13315_), .A2(new_n13318_), .B(\asqrt[27] ), .ZN(new_n13319_));
  NAND3_X1   g13127(.A1(new_n13312_), .A2(new_n6966_), .A3(new_n13319_), .ZN(new_n13320_));
  AOI21_X1   g13128(.A1(new_n13312_), .A2(new_n13319_), .B(new_n6966_), .ZN(new_n13321_));
  AOI21_X1   g13129(.A1(new_n13171_), .A2(new_n13320_), .B(new_n13321_), .ZN(new_n13322_));
  AOI21_X1   g13130(.A1(new_n13322_), .A2(new_n6636_), .B(new_n13168_), .ZN(new_n13323_));
  INV_X1     g13131(.I(new_n13173_), .ZN(new_n13324_));
  NOR3_X1    g13132(.A1(new_n13315_), .A2(\asqrt[27] ), .A3(new_n13318_), .ZN(new_n13325_));
  OAI21_X1   g13133(.A1(new_n13324_), .A2(new_n13325_), .B(new_n13319_), .ZN(new_n13326_));
  OAI21_X1   g13134(.A1(new_n13326_), .A2(\asqrt[28] ), .B(new_n13171_), .ZN(new_n13327_));
  NAND2_X1   g13135(.A1(new_n13326_), .A2(\asqrt[28] ), .ZN(new_n13328_));
  AOI21_X1   g13136(.A1(new_n13327_), .A2(new_n13328_), .B(new_n6636_), .ZN(new_n13329_));
  NOR3_X1    g13137(.A1(new_n13323_), .A2(\asqrt[30] ), .A3(new_n13329_), .ZN(new_n13330_));
  OAI21_X1   g13138(.A1(new_n13323_), .A2(new_n13329_), .B(\asqrt[30] ), .ZN(new_n13331_));
  OAI21_X1   g13139(.A1(new_n13165_), .A2(new_n13330_), .B(new_n13331_), .ZN(new_n13332_));
  OAI21_X1   g13140(.A1(new_n13332_), .A2(\asqrt[31] ), .B(new_n13161_), .ZN(new_n13333_));
  NAND3_X1   g13141(.A1(new_n13327_), .A2(new_n13328_), .A3(new_n6636_), .ZN(new_n13334_));
  AOI21_X1   g13142(.A1(new_n13167_), .A2(new_n13334_), .B(new_n13329_), .ZN(new_n13335_));
  AOI21_X1   g13143(.A1(new_n13335_), .A2(new_n6275_), .B(new_n13165_), .ZN(new_n13336_));
  NAND2_X1   g13144(.A1(new_n13334_), .A2(new_n13167_), .ZN(new_n13337_));
  INV_X1     g13145(.I(new_n13329_), .ZN(new_n13338_));
  AOI21_X1   g13146(.A1(new_n13337_), .A2(new_n13338_), .B(new_n6275_), .ZN(new_n13339_));
  OAI21_X1   g13147(.A1(new_n13336_), .A2(new_n13339_), .B(\asqrt[31] ), .ZN(new_n13340_));
  NAND3_X1   g13148(.A1(new_n13333_), .A2(new_n5643_), .A3(new_n13340_), .ZN(new_n13341_));
  AOI21_X1   g13149(.A1(new_n13333_), .A2(new_n13340_), .B(new_n5643_), .ZN(new_n13342_));
  AOI21_X1   g13150(.A1(new_n13159_), .A2(new_n13341_), .B(new_n13342_), .ZN(new_n13343_));
  AOI21_X1   g13151(.A1(new_n13343_), .A2(new_n5336_), .B(new_n13156_), .ZN(new_n13344_));
  INV_X1     g13152(.I(new_n13161_), .ZN(new_n13345_));
  NOR3_X1    g13153(.A1(new_n13336_), .A2(\asqrt[31] ), .A3(new_n13339_), .ZN(new_n13346_));
  OAI21_X1   g13154(.A1(new_n13345_), .A2(new_n13346_), .B(new_n13340_), .ZN(new_n13347_));
  OAI21_X1   g13155(.A1(new_n13347_), .A2(\asqrt[32] ), .B(new_n13159_), .ZN(new_n13348_));
  NAND2_X1   g13156(.A1(new_n13347_), .A2(\asqrt[32] ), .ZN(new_n13349_));
  AOI21_X1   g13157(.A1(new_n13348_), .A2(new_n13349_), .B(new_n5336_), .ZN(new_n13350_));
  NOR3_X1    g13158(.A1(new_n13344_), .A2(\asqrt[34] ), .A3(new_n13350_), .ZN(new_n13351_));
  OAI21_X1   g13159(.A1(new_n13344_), .A2(new_n13350_), .B(\asqrt[34] ), .ZN(new_n13352_));
  OAI21_X1   g13160(.A1(new_n13153_), .A2(new_n13351_), .B(new_n13352_), .ZN(new_n13353_));
  OAI21_X1   g13161(.A1(new_n13353_), .A2(\asqrt[35] ), .B(new_n13149_), .ZN(new_n13354_));
  NAND3_X1   g13162(.A1(new_n13348_), .A2(new_n13349_), .A3(new_n5336_), .ZN(new_n13355_));
  AOI21_X1   g13163(.A1(new_n13155_), .A2(new_n13355_), .B(new_n13350_), .ZN(new_n13356_));
  AOI21_X1   g13164(.A1(new_n13356_), .A2(new_n5029_), .B(new_n13153_), .ZN(new_n13357_));
  NAND2_X1   g13165(.A1(new_n13355_), .A2(new_n13155_), .ZN(new_n13358_));
  INV_X1     g13166(.I(new_n13350_), .ZN(new_n13359_));
  AOI21_X1   g13167(.A1(new_n13358_), .A2(new_n13359_), .B(new_n5029_), .ZN(new_n13360_));
  OAI21_X1   g13168(.A1(new_n13357_), .A2(new_n13360_), .B(\asqrt[35] ), .ZN(new_n13361_));
  NAND3_X1   g13169(.A1(new_n13354_), .A2(new_n4461_), .A3(new_n13361_), .ZN(new_n13362_));
  AOI21_X1   g13170(.A1(new_n13354_), .A2(new_n13361_), .B(new_n4461_), .ZN(new_n13363_));
  AOI21_X1   g13171(.A1(new_n13147_), .A2(new_n13362_), .B(new_n13363_), .ZN(new_n13364_));
  AOI21_X1   g13172(.A1(new_n13364_), .A2(new_n4196_), .B(new_n13144_), .ZN(new_n13365_));
  INV_X1     g13173(.I(new_n13149_), .ZN(new_n13366_));
  NOR3_X1    g13174(.A1(new_n13357_), .A2(\asqrt[35] ), .A3(new_n13360_), .ZN(new_n13367_));
  OAI21_X1   g13175(.A1(new_n13366_), .A2(new_n13367_), .B(new_n13361_), .ZN(new_n13368_));
  OAI21_X1   g13176(.A1(new_n13368_), .A2(\asqrt[36] ), .B(new_n13147_), .ZN(new_n13369_));
  NAND2_X1   g13177(.A1(new_n13368_), .A2(\asqrt[36] ), .ZN(new_n13370_));
  AOI21_X1   g13178(.A1(new_n13369_), .A2(new_n13370_), .B(new_n4196_), .ZN(new_n13371_));
  NOR3_X1    g13179(.A1(new_n13365_), .A2(\asqrt[38] ), .A3(new_n13371_), .ZN(new_n13372_));
  OAI21_X1   g13180(.A1(new_n13365_), .A2(new_n13371_), .B(\asqrt[38] ), .ZN(new_n13373_));
  OAI21_X1   g13181(.A1(new_n13141_), .A2(new_n13372_), .B(new_n13373_), .ZN(new_n13374_));
  OAI21_X1   g13182(.A1(new_n13374_), .A2(\asqrt[39] ), .B(new_n13137_), .ZN(new_n13375_));
  NAND3_X1   g13183(.A1(new_n13369_), .A2(new_n13370_), .A3(new_n4196_), .ZN(new_n13376_));
  AOI21_X1   g13184(.A1(new_n13143_), .A2(new_n13376_), .B(new_n13371_), .ZN(new_n13377_));
  AOI21_X1   g13185(.A1(new_n13377_), .A2(new_n3925_), .B(new_n13141_), .ZN(new_n13378_));
  NAND2_X1   g13186(.A1(new_n13376_), .A2(new_n13143_), .ZN(new_n13379_));
  INV_X1     g13187(.I(new_n13371_), .ZN(new_n13380_));
  AOI21_X1   g13188(.A1(new_n13379_), .A2(new_n13380_), .B(new_n3925_), .ZN(new_n13381_));
  OAI21_X1   g13189(.A1(new_n13378_), .A2(new_n13381_), .B(\asqrt[39] ), .ZN(new_n13382_));
  NAND3_X1   g13190(.A1(new_n13375_), .A2(new_n3427_), .A3(new_n13382_), .ZN(new_n13383_));
  AOI21_X1   g13191(.A1(new_n13375_), .A2(new_n13382_), .B(new_n3427_), .ZN(new_n13384_));
  AOI21_X1   g13192(.A1(new_n13135_), .A2(new_n13383_), .B(new_n13384_), .ZN(new_n13385_));
  AOI21_X1   g13193(.A1(new_n13385_), .A2(new_n3195_), .B(new_n13132_), .ZN(new_n13386_));
  INV_X1     g13194(.I(new_n13137_), .ZN(new_n13387_));
  NOR3_X1    g13195(.A1(new_n13378_), .A2(\asqrt[39] ), .A3(new_n13381_), .ZN(new_n13388_));
  OAI21_X1   g13196(.A1(new_n13387_), .A2(new_n13388_), .B(new_n13382_), .ZN(new_n13389_));
  OAI21_X1   g13197(.A1(new_n13389_), .A2(\asqrt[40] ), .B(new_n13135_), .ZN(new_n13390_));
  NAND2_X1   g13198(.A1(new_n13389_), .A2(\asqrt[40] ), .ZN(new_n13391_));
  AOI21_X1   g13199(.A1(new_n13390_), .A2(new_n13391_), .B(new_n3195_), .ZN(new_n13392_));
  NOR3_X1    g13200(.A1(new_n13386_), .A2(\asqrt[42] ), .A3(new_n13392_), .ZN(new_n13393_));
  OAI21_X1   g13201(.A1(new_n13386_), .A2(new_n13392_), .B(\asqrt[42] ), .ZN(new_n13394_));
  OAI21_X1   g13202(.A1(new_n13129_), .A2(new_n13393_), .B(new_n13394_), .ZN(new_n13395_));
  OAI21_X1   g13203(.A1(new_n13395_), .A2(\asqrt[43] ), .B(new_n13125_), .ZN(new_n13396_));
  NAND3_X1   g13204(.A1(new_n13390_), .A2(new_n13391_), .A3(new_n3195_), .ZN(new_n13397_));
  AOI21_X1   g13205(.A1(new_n13131_), .A2(new_n13397_), .B(new_n13392_), .ZN(new_n13398_));
  AOI21_X1   g13206(.A1(new_n13398_), .A2(new_n2960_), .B(new_n13129_), .ZN(new_n13399_));
  NAND2_X1   g13207(.A1(new_n13397_), .A2(new_n13131_), .ZN(new_n13400_));
  INV_X1     g13208(.I(new_n13392_), .ZN(new_n13401_));
  AOI21_X1   g13209(.A1(new_n13400_), .A2(new_n13401_), .B(new_n2960_), .ZN(new_n13402_));
  OAI21_X1   g13210(.A1(new_n13399_), .A2(new_n13402_), .B(\asqrt[43] ), .ZN(new_n13403_));
  NAND3_X1   g13211(.A1(new_n13396_), .A2(new_n2531_), .A3(new_n13403_), .ZN(new_n13404_));
  AOI21_X1   g13212(.A1(new_n13396_), .A2(new_n13403_), .B(new_n2531_), .ZN(new_n13405_));
  AOI21_X1   g13213(.A1(new_n13123_), .A2(new_n13404_), .B(new_n13405_), .ZN(new_n13406_));
  AOI21_X1   g13214(.A1(new_n13406_), .A2(new_n2332_), .B(new_n13120_), .ZN(new_n13407_));
  INV_X1     g13215(.I(new_n13125_), .ZN(new_n13408_));
  NOR3_X1    g13216(.A1(new_n13399_), .A2(\asqrt[43] ), .A3(new_n13402_), .ZN(new_n13409_));
  OAI21_X1   g13217(.A1(new_n13408_), .A2(new_n13409_), .B(new_n13403_), .ZN(new_n13410_));
  OAI21_X1   g13218(.A1(new_n13410_), .A2(\asqrt[44] ), .B(new_n13123_), .ZN(new_n13411_));
  NAND2_X1   g13219(.A1(new_n13410_), .A2(\asqrt[44] ), .ZN(new_n13412_));
  AOI21_X1   g13220(.A1(new_n13411_), .A2(new_n13412_), .B(new_n2332_), .ZN(new_n13413_));
  NOR3_X1    g13221(.A1(new_n13407_), .A2(\asqrt[46] ), .A3(new_n13413_), .ZN(new_n13414_));
  OAI21_X1   g13222(.A1(new_n13407_), .A2(new_n13413_), .B(\asqrt[46] ), .ZN(new_n13415_));
  OAI21_X1   g13223(.A1(new_n13117_), .A2(new_n13414_), .B(new_n13415_), .ZN(new_n13416_));
  OAI21_X1   g13224(.A1(new_n13416_), .A2(\asqrt[47] ), .B(new_n13113_), .ZN(new_n13417_));
  NAND3_X1   g13225(.A1(new_n13411_), .A2(new_n13412_), .A3(new_n2332_), .ZN(new_n13418_));
  AOI21_X1   g13226(.A1(new_n13119_), .A2(new_n13418_), .B(new_n13413_), .ZN(new_n13419_));
  AOI21_X1   g13227(.A1(new_n13419_), .A2(new_n2134_), .B(new_n13117_), .ZN(new_n13420_));
  NAND2_X1   g13228(.A1(new_n13418_), .A2(new_n13119_), .ZN(new_n13421_));
  INV_X1     g13229(.I(new_n13413_), .ZN(new_n13422_));
  AOI21_X1   g13230(.A1(new_n13421_), .A2(new_n13422_), .B(new_n2134_), .ZN(new_n13423_));
  OAI21_X1   g13231(.A1(new_n13420_), .A2(new_n13423_), .B(\asqrt[47] ), .ZN(new_n13424_));
  NAND3_X1   g13232(.A1(new_n13417_), .A2(new_n1778_), .A3(new_n13424_), .ZN(new_n13425_));
  AOI21_X1   g13233(.A1(new_n13417_), .A2(new_n13424_), .B(new_n1778_), .ZN(new_n13426_));
  AOI21_X1   g13234(.A1(new_n13111_), .A2(new_n13425_), .B(new_n13426_), .ZN(new_n13427_));
  AOI21_X1   g13235(.A1(new_n13427_), .A2(new_n1632_), .B(new_n13108_), .ZN(new_n13428_));
  INV_X1     g13236(.I(new_n13113_), .ZN(new_n13429_));
  NOR3_X1    g13237(.A1(new_n13420_), .A2(\asqrt[47] ), .A3(new_n13423_), .ZN(new_n13430_));
  OAI21_X1   g13238(.A1(new_n13429_), .A2(new_n13430_), .B(new_n13424_), .ZN(new_n13431_));
  OAI21_X1   g13239(.A1(new_n13431_), .A2(\asqrt[48] ), .B(new_n13111_), .ZN(new_n13432_));
  NAND2_X1   g13240(.A1(new_n13431_), .A2(\asqrt[48] ), .ZN(new_n13433_));
  AOI21_X1   g13241(.A1(new_n13432_), .A2(new_n13433_), .B(new_n1632_), .ZN(new_n13434_));
  NOR3_X1    g13242(.A1(new_n13428_), .A2(\asqrt[50] ), .A3(new_n13434_), .ZN(new_n13435_));
  OAI21_X1   g13243(.A1(new_n13428_), .A2(new_n13434_), .B(\asqrt[50] ), .ZN(new_n13436_));
  OAI21_X1   g13244(.A1(new_n13105_), .A2(new_n13435_), .B(new_n13436_), .ZN(new_n13437_));
  OAI21_X1   g13245(.A1(new_n13437_), .A2(\asqrt[51] ), .B(new_n13101_), .ZN(new_n13438_));
  NAND3_X1   g13246(.A1(new_n13432_), .A2(new_n13433_), .A3(new_n1632_), .ZN(new_n13439_));
  AOI21_X1   g13247(.A1(new_n13107_), .A2(new_n13439_), .B(new_n13434_), .ZN(new_n13440_));
  AOI21_X1   g13248(.A1(new_n13440_), .A2(new_n1463_), .B(new_n13105_), .ZN(new_n13441_));
  NAND2_X1   g13249(.A1(new_n13439_), .A2(new_n13107_), .ZN(new_n13442_));
  INV_X1     g13250(.I(new_n13434_), .ZN(new_n13443_));
  AOI21_X1   g13251(.A1(new_n13442_), .A2(new_n13443_), .B(new_n1463_), .ZN(new_n13444_));
  OAI21_X1   g13252(.A1(new_n13441_), .A2(new_n13444_), .B(\asqrt[51] ), .ZN(new_n13445_));
  NAND3_X1   g13253(.A1(new_n13438_), .A2(new_n1150_), .A3(new_n13445_), .ZN(new_n13446_));
  INV_X1     g13254(.I(new_n13101_), .ZN(new_n13447_));
  NOR3_X1    g13255(.A1(new_n13441_), .A2(\asqrt[51] ), .A3(new_n13444_), .ZN(new_n13448_));
  OAI21_X1   g13256(.A1(new_n13447_), .A2(new_n13448_), .B(new_n13445_), .ZN(new_n13449_));
  NAND2_X1   g13257(.A1(new_n13449_), .A2(\asqrt[52] ), .ZN(new_n13450_));
  NOR2_X1    g13258(.A1(new_n13069_), .A2(\asqrt[62] ), .ZN(new_n13451_));
  INV_X1     g13259(.I(new_n13088_), .ZN(new_n13452_));
  NOR2_X1    g13260(.A1(new_n13452_), .A2(new_n13451_), .ZN(new_n13453_));
  XOR2_X1    g13261(.A1(new_n13079_), .A2(new_n12565_), .Z(new_n13454_));
  OAI21_X1   g13262(.A1(\asqrt[13] ), .A2(new_n13453_), .B(new_n13454_), .ZN(new_n13455_));
  INV_X1     g13263(.I(new_n13455_), .ZN(new_n13456_));
  NAND2_X1   g13264(.A1(new_n13037_), .A2(new_n337_), .ZN(new_n13457_));
  AOI21_X1   g13265(.A1(new_n13457_), .A2(new_n13061_), .B(\asqrt[13] ), .ZN(new_n13458_));
  XOR2_X1    g13266(.A1(new_n13458_), .A2(new_n12983_), .Z(new_n13459_));
  INV_X1     g13267(.I(new_n13459_), .ZN(new_n13460_));
  AOI21_X1   g13268(.A1(new_n13035_), .A2(new_n13052_), .B(\asqrt[13] ), .ZN(new_n13461_));
  XOR2_X1    g13269(.A1(new_n13461_), .A2(new_n12987_), .Z(new_n13462_));
  INV_X1     g13270(.I(new_n13462_), .ZN(new_n13463_));
  NAND2_X1   g13271(.A1(new_n13048_), .A2(new_n531_), .ZN(new_n13464_));
  AOI21_X1   g13272(.A1(new_n13464_), .A2(new_n13034_), .B(\asqrt[13] ), .ZN(new_n13465_));
  XOR2_X1    g13273(.A1(new_n13465_), .A2(new_n12990_), .Z(new_n13466_));
  INV_X1     g13274(.I(new_n13466_), .ZN(new_n13467_));
  AOI21_X1   g13275(.A1(new_n13046_), .A2(new_n13031_), .B(\asqrt[13] ), .ZN(new_n13468_));
  XOR2_X1    g13276(.A1(new_n13468_), .A2(new_n12992_), .Z(new_n13469_));
  NAND2_X1   g13277(.A1(new_n13017_), .A2(new_n744_), .ZN(new_n13470_));
  AOI21_X1   g13278(.A1(new_n13470_), .A2(new_n13045_), .B(\asqrt[13] ), .ZN(new_n13471_));
  XOR2_X1    g13279(.A1(new_n13471_), .A2(new_n12995_), .Z(new_n13472_));
  AOI21_X1   g13280(.A1(new_n13015_), .A2(new_n13028_), .B(\asqrt[13] ), .ZN(new_n13473_));
  XOR2_X1    g13281(.A1(new_n13473_), .A2(new_n12999_), .Z(new_n13474_));
  INV_X1     g13282(.I(new_n13474_), .ZN(new_n13475_));
  NAND2_X1   g13283(.A1(new_n13024_), .A2(new_n1006_), .ZN(new_n13476_));
  AOI21_X1   g13284(.A1(new_n13476_), .A2(new_n13014_), .B(\asqrt[13] ), .ZN(new_n13477_));
  XOR2_X1    g13285(.A1(new_n13477_), .A2(new_n13002_), .Z(new_n13478_));
  INV_X1     g13286(.I(new_n13478_), .ZN(new_n13479_));
  AOI21_X1   g13287(.A1(new_n13022_), .A2(new_n13011_), .B(\asqrt[13] ), .ZN(new_n13480_));
  XOR2_X1    g13288(.A1(new_n13480_), .A2(new_n13004_), .Z(new_n13481_));
  OAI21_X1   g13289(.A1(new_n13449_), .A2(\asqrt[52] ), .B(new_n13099_), .ZN(new_n13482_));
  NAND3_X1   g13290(.A1(new_n13482_), .A2(new_n13450_), .A3(new_n1006_), .ZN(new_n13483_));
  AOI21_X1   g13291(.A1(new_n13482_), .A2(new_n13450_), .B(new_n1006_), .ZN(new_n13484_));
  AOI21_X1   g13292(.A1(new_n13481_), .A2(new_n13483_), .B(new_n13484_), .ZN(new_n13485_));
  AOI21_X1   g13293(.A1(new_n13485_), .A2(new_n860_), .B(new_n13479_), .ZN(new_n13486_));
  NAND2_X1   g13294(.A1(new_n13483_), .A2(new_n13481_), .ZN(new_n13487_));
  INV_X1     g13295(.I(new_n13484_), .ZN(new_n13488_));
  AOI21_X1   g13296(.A1(new_n13487_), .A2(new_n13488_), .B(new_n860_), .ZN(new_n13489_));
  NOR3_X1    g13297(.A1(new_n13486_), .A2(\asqrt[55] ), .A3(new_n13489_), .ZN(new_n13490_));
  OAI21_X1   g13298(.A1(new_n13486_), .A2(new_n13489_), .B(\asqrt[55] ), .ZN(new_n13491_));
  OAI21_X1   g13299(.A1(new_n13475_), .A2(new_n13490_), .B(new_n13491_), .ZN(new_n13492_));
  OAI21_X1   g13300(.A1(new_n13492_), .A2(\asqrt[56] ), .B(new_n13472_), .ZN(new_n13493_));
  NAND2_X1   g13301(.A1(new_n13492_), .A2(\asqrt[56] ), .ZN(new_n13494_));
  NAND3_X1   g13302(.A1(new_n13493_), .A2(new_n13494_), .A3(new_n531_), .ZN(new_n13495_));
  AOI21_X1   g13303(.A1(new_n13493_), .A2(new_n13494_), .B(new_n531_), .ZN(new_n13496_));
  AOI21_X1   g13304(.A1(new_n13469_), .A2(new_n13495_), .B(new_n13496_), .ZN(new_n13497_));
  AOI21_X1   g13305(.A1(new_n13497_), .A2(new_n423_), .B(new_n13467_), .ZN(new_n13498_));
  NAND2_X1   g13306(.A1(new_n13495_), .A2(new_n13469_), .ZN(new_n13499_));
  INV_X1     g13307(.I(new_n13496_), .ZN(new_n13500_));
  AOI21_X1   g13308(.A1(new_n13499_), .A2(new_n13500_), .B(new_n423_), .ZN(new_n13501_));
  NOR3_X1    g13309(.A1(new_n13498_), .A2(\asqrt[59] ), .A3(new_n13501_), .ZN(new_n13502_));
  NOR2_X1    g13310(.A1(new_n13502_), .A2(new_n13463_), .ZN(new_n13503_));
  OAI21_X1   g13311(.A1(new_n13498_), .A2(new_n13501_), .B(\asqrt[59] ), .ZN(new_n13504_));
  INV_X1     g13312(.I(new_n13504_), .ZN(new_n13505_));
  NOR2_X1    g13313(.A1(new_n13503_), .A2(new_n13505_), .ZN(new_n13506_));
  AOI21_X1   g13314(.A1(new_n13506_), .A2(new_n266_), .B(new_n13460_), .ZN(new_n13507_));
  INV_X1     g13315(.I(new_n13469_), .ZN(new_n13508_));
  INV_X1     g13316(.I(new_n13481_), .ZN(new_n13509_));
  AOI21_X1   g13317(.A1(new_n13438_), .A2(new_n13445_), .B(new_n1150_), .ZN(new_n13510_));
  AOI21_X1   g13318(.A1(new_n13099_), .A2(new_n13446_), .B(new_n13510_), .ZN(new_n13511_));
  AOI21_X1   g13319(.A1(new_n13511_), .A2(new_n1006_), .B(new_n13509_), .ZN(new_n13512_));
  NOR3_X1    g13320(.A1(new_n13512_), .A2(\asqrt[54] ), .A3(new_n13484_), .ZN(new_n13513_));
  OAI21_X1   g13321(.A1(new_n13512_), .A2(new_n13484_), .B(\asqrt[54] ), .ZN(new_n13514_));
  OAI21_X1   g13322(.A1(new_n13479_), .A2(new_n13513_), .B(new_n13514_), .ZN(new_n13515_));
  OAI21_X1   g13323(.A1(new_n13515_), .A2(\asqrt[55] ), .B(new_n13474_), .ZN(new_n13516_));
  NAND3_X1   g13324(.A1(new_n13516_), .A2(new_n634_), .A3(new_n13491_), .ZN(new_n13517_));
  AOI21_X1   g13325(.A1(new_n13516_), .A2(new_n13491_), .B(new_n634_), .ZN(new_n13518_));
  AOI21_X1   g13326(.A1(new_n13472_), .A2(new_n13517_), .B(new_n13518_), .ZN(new_n13519_));
  AOI21_X1   g13327(.A1(new_n13519_), .A2(new_n531_), .B(new_n13508_), .ZN(new_n13520_));
  NOR3_X1    g13328(.A1(new_n13520_), .A2(\asqrt[58] ), .A3(new_n13496_), .ZN(new_n13521_));
  OAI21_X1   g13329(.A1(new_n13520_), .A2(new_n13496_), .B(\asqrt[58] ), .ZN(new_n13522_));
  OAI21_X1   g13330(.A1(new_n13467_), .A2(new_n13521_), .B(new_n13522_), .ZN(new_n13523_));
  OAI21_X1   g13331(.A1(new_n13523_), .A2(\asqrt[59] ), .B(new_n13462_), .ZN(new_n13524_));
  AOI21_X1   g13332(.A1(new_n13524_), .A2(new_n13504_), .B(new_n266_), .ZN(new_n13525_));
  OAI21_X1   g13333(.A1(new_n13507_), .A2(new_n13525_), .B(\asqrt[61] ), .ZN(new_n13526_));
  AOI21_X1   g13334(.A1(new_n13070_), .A2(new_n13064_), .B(\asqrt[13] ), .ZN(new_n13527_));
  XOR2_X1    g13335(.A1(new_n13527_), .A2(new_n12980_), .Z(new_n13528_));
  OAI21_X1   g13336(.A1(new_n13463_), .A2(new_n13502_), .B(new_n13504_), .ZN(new_n13529_));
  OAI21_X1   g13337(.A1(new_n13529_), .A2(\asqrt[60] ), .B(new_n13459_), .ZN(new_n13530_));
  OAI21_X1   g13338(.A1(new_n13503_), .A2(new_n13505_), .B(\asqrt[60] ), .ZN(new_n13531_));
  NAND3_X1   g13339(.A1(new_n13530_), .A2(new_n239_), .A3(new_n13531_), .ZN(new_n13532_));
  NAND2_X1   g13340(.A1(new_n13532_), .A2(new_n13528_), .ZN(new_n13533_));
  NAND2_X1   g13341(.A1(new_n13533_), .A2(new_n13526_), .ZN(new_n13534_));
  AOI21_X1   g13342(.A1(new_n13530_), .A2(new_n13531_), .B(new_n239_), .ZN(new_n13535_));
  NAND3_X1   g13343(.A1(new_n13524_), .A2(new_n266_), .A3(new_n13504_), .ZN(new_n13536_));
  AOI21_X1   g13344(.A1(new_n13459_), .A2(new_n13536_), .B(new_n13525_), .ZN(new_n13537_));
  INV_X1     g13345(.I(new_n13528_), .ZN(new_n13538_));
  AOI21_X1   g13346(.A1(new_n13537_), .A2(new_n239_), .B(new_n13538_), .ZN(new_n13539_));
  OAI21_X1   g13347(.A1(new_n13539_), .A2(new_n13535_), .B(new_n201_), .ZN(new_n13540_));
  NAND3_X1   g13348(.A1(new_n13533_), .A2(\asqrt[62] ), .A3(new_n13526_), .ZN(new_n13541_));
  AOI21_X1   g13349(.A1(new_n13063_), .A2(new_n13211_), .B(\asqrt[13] ), .ZN(new_n13542_));
  XOR2_X1    g13350(.A1(new_n13542_), .A2(new_n13067_), .Z(new_n13543_));
  INV_X1     g13351(.I(new_n13543_), .ZN(new_n13544_));
  AOI22_X1   g13352(.A1(new_n13540_), .A2(new_n13541_), .B1(new_n13534_), .B2(new_n13544_), .ZN(new_n13545_));
  NOR2_X1    g13353(.A1(new_n13082_), .A2(new_n12978_), .ZN(new_n13546_));
  OAI21_X1   g13354(.A1(\asqrt[13] ), .A2(new_n13546_), .B(new_n13089_), .ZN(new_n13547_));
  INV_X1     g13355(.I(new_n13547_), .ZN(new_n13548_));
  OAI21_X1   g13356(.A1(new_n13545_), .A2(new_n13456_), .B(new_n13548_), .ZN(new_n13549_));
  OAI21_X1   g13357(.A1(new_n13534_), .A2(\asqrt[62] ), .B(new_n13543_), .ZN(new_n13550_));
  NAND2_X1   g13358(.A1(new_n13534_), .A2(\asqrt[62] ), .ZN(new_n13551_));
  NAND3_X1   g13359(.A1(new_n13550_), .A2(new_n13551_), .A3(new_n13456_), .ZN(new_n13552_));
  NAND2_X1   g13360(.A1(new_n13228_), .A2(new_n12977_), .ZN(new_n13553_));
  XOR2_X1    g13361(.A1(new_n13082_), .A2(new_n12978_), .Z(new_n13554_));
  NAND3_X1   g13362(.A1(new_n13553_), .A2(\asqrt[63] ), .A3(new_n13554_), .ZN(new_n13555_));
  INV_X1     g13363(.I(new_n13226_), .ZN(new_n13556_));
  NAND4_X1   g13364(.A1(new_n13556_), .A2(new_n12978_), .A3(new_n13089_), .A4(new_n13096_), .ZN(new_n13557_));
  NAND2_X1   g13365(.A1(new_n13555_), .A2(new_n13557_), .ZN(new_n13558_));
  INV_X1     g13366(.I(new_n13558_), .ZN(new_n13559_));
  NAND4_X1   g13367(.A1(new_n13549_), .A2(new_n193_), .A3(new_n13552_), .A4(new_n13559_), .ZN(\asqrt[12] ));
  AOI21_X1   g13368(.A1(new_n13446_), .A2(new_n13450_), .B(\asqrt[12] ), .ZN(new_n13561_));
  XOR2_X1    g13369(.A1(new_n13561_), .A2(new_n13099_), .Z(new_n13562_));
  XOR2_X1    g13370(.A1(new_n13437_), .A2(\asqrt[51] ), .Z(new_n13563_));
  NOR2_X1    g13371(.A1(\asqrt[12] ), .A2(new_n13563_), .ZN(new_n13564_));
  XOR2_X1    g13372(.A1(new_n13564_), .A2(new_n13101_), .Z(new_n13565_));
  NOR2_X1    g13373(.A1(new_n13435_), .A2(new_n13444_), .ZN(new_n13566_));
  NOR2_X1    g13374(.A1(\asqrt[12] ), .A2(new_n13566_), .ZN(new_n13567_));
  XOR2_X1    g13375(.A1(new_n13567_), .A2(new_n13104_), .Z(new_n13568_));
  AOI21_X1   g13376(.A1(new_n13439_), .A2(new_n13443_), .B(\asqrt[12] ), .ZN(new_n13569_));
  XOR2_X1    g13377(.A1(new_n13569_), .A2(new_n13107_), .Z(new_n13570_));
  INV_X1     g13378(.I(new_n13570_), .ZN(new_n13571_));
  AOI21_X1   g13379(.A1(new_n13425_), .A2(new_n13433_), .B(\asqrt[12] ), .ZN(new_n13572_));
  XOR2_X1    g13380(.A1(new_n13572_), .A2(new_n13111_), .Z(new_n13573_));
  INV_X1     g13381(.I(new_n13573_), .ZN(new_n13574_));
  XOR2_X1    g13382(.A1(new_n13416_), .A2(\asqrt[47] ), .Z(new_n13575_));
  NOR2_X1    g13383(.A1(\asqrt[12] ), .A2(new_n13575_), .ZN(new_n13576_));
  XOR2_X1    g13384(.A1(new_n13576_), .A2(new_n13113_), .Z(new_n13577_));
  NOR2_X1    g13385(.A1(new_n13414_), .A2(new_n13423_), .ZN(new_n13578_));
  NOR2_X1    g13386(.A1(\asqrt[12] ), .A2(new_n13578_), .ZN(new_n13579_));
  XOR2_X1    g13387(.A1(new_n13579_), .A2(new_n13116_), .Z(new_n13580_));
  AOI21_X1   g13388(.A1(new_n13418_), .A2(new_n13422_), .B(\asqrt[12] ), .ZN(new_n13581_));
  XOR2_X1    g13389(.A1(new_n13581_), .A2(new_n13119_), .Z(new_n13582_));
  INV_X1     g13390(.I(new_n13582_), .ZN(new_n13583_));
  AOI21_X1   g13391(.A1(new_n13404_), .A2(new_n13412_), .B(\asqrt[12] ), .ZN(new_n13584_));
  XOR2_X1    g13392(.A1(new_n13584_), .A2(new_n13123_), .Z(new_n13585_));
  INV_X1     g13393(.I(new_n13585_), .ZN(new_n13586_));
  XOR2_X1    g13394(.A1(new_n13395_), .A2(\asqrt[43] ), .Z(new_n13587_));
  NOR2_X1    g13395(.A1(\asqrt[12] ), .A2(new_n13587_), .ZN(new_n13588_));
  XOR2_X1    g13396(.A1(new_n13588_), .A2(new_n13125_), .Z(new_n13589_));
  NOR2_X1    g13397(.A1(new_n13393_), .A2(new_n13402_), .ZN(new_n13590_));
  NOR2_X1    g13398(.A1(\asqrt[12] ), .A2(new_n13590_), .ZN(new_n13591_));
  XOR2_X1    g13399(.A1(new_n13591_), .A2(new_n13128_), .Z(new_n13592_));
  AOI21_X1   g13400(.A1(new_n13397_), .A2(new_n13401_), .B(\asqrt[12] ), .ZN(new_n13593_));
  XOR2_X1    g13401(.A1(new_n13593_), .A2(new_n13131_), .Z(new_n13594_));
  INV_X1     g13402(.I(new_n13594_), .ZN(new_n13595_));
  AOI21_X1   g13403(.A1(new_n13383_), .A2(new_n13391_), .B(\asqrt[12] ), .ZN(new_n13596_));
  XOR2_X1    g13404(.A1(new_n13596_), .A2(new_n13135_), .Z(new_n13597_));
  INV_X1     g13405(.I(new_n13597_), .ZN(new_n13598_));
  XOR2_X1    g13406(.A1(new_n13374_), .A2(\asqrt[39] ), .Z(new_n13599_));
  NOR2_X1    g13407(.A1(\asqrt[12] ), .A2(new_n13599_), .ZN(new_n13600_));
  XOR2_X1    g13408(.A1(new_n13600_), .A2(new_n13137_), .Z(new_n13601_));
  NOR2_X1    g13409(.A1(new_n13372_), .A2(new_n13381_), .ZN(new_n13602_));
  NOR2_X1    g13410(.A1(\asqrt[12] ), .A2(new_n13602_), .ZN(new_n13603_));
  XOR2_X1    g13411(.A1(new_n13603_), .A2(new_n13140_), .Z(new_n13604_));
  AOI21_X1   g13412(.A1(new_n13376_), .A2(new_n13380_), .B(\asqrt[12] ), .ZN(new_n13605_));
  XOR2_X1    g13413(.A1(new_n13605_), .A2(new_n13143_), .Z(new_n13606_));
  INV_X1     g13414(.I(new_n13606_), .ZN(new_n13607_));
  AOI21_X1   g13415(.A1(new_n13362_), .A2(new_n13370_), .B(\asqrt[12] ), .ZN(new_n13608_));
  XOR2_X1    g13416(.A1(new_n13608_), .A2(new_n13147_), .Z(new_n13609_));
  INV_X1     g13417(.I(new_n13609_), .ZN(new_n13610_));
  XOR2_X1    g13418(.A1(new_n13353_), .A2(\asqrt[35] ), .Z(new_n13611_));
  NOR2_X1    g13419(.A1(\asqrt[12] ), .A2(new_n13611_), .ZN(new_n13612_));
  XOR2_X1    g13420(.A1(new_n13612_), .A2(new_n13149_), .Z(new_n13613_));
  NOR2_X1    g13421(.A1(new_n13351_), .A2(new_n13360_), .ZN(new_n13614_));
  NOR2_X1    g13422(.A1(\asqrt[12] ), .A2(new_n13614_), .ZN(new_n13615_));
  XOR2_X1    g13423(.A1(new_n13615_), .A2(new_n13152_), .Z(new_n13616_));
  AOI21_X1   g13424(.A1(new_n13355_), .A2(new_n13359_), .B(\asqrt[12] ), .ZN(new_n13617_));
  XOR2_X1    g13425(.A1(new_n13617_), .A2(new_n13155_), .Z(new_n13618_));
  INV_X1     g13426(.I(new_n13618_), .ZN(new_n13619_));
  AOI21_X1   g13427(.A1(new_n13341_), .A2(new_n13349_), .B(\asqrt[12] ), .ZN(new_n13620_));
  XOR2_X1    g13428(.A1(new_n13620_), .A2(new_n13159_), .Z(new_n13621_));
  INV_X1     g13429(.I(new_n13621_), .ZN(new_n13622_));
  XOR2_X1    g13430(.A1(new_n13332_), .A2(\asqrt[31] ), .Z(new_n13623_));
  NOR2_X1    g13431(.A1(\asqrt[12] ), .A2(new_n13623_), .ZN(new_n13624_));
  XOR2_X1    g13432(.A1(new_n13624_), .A2(new_n13161_), .Z(new_n13625_));
  NOR2_X1    g13433(.A1(new_n13330_), .A2(new_n13339_), .ZN(new_n13626_));
  NOR2_X1    g13434(.A1(\asqrt[12] ), .A2(new_n13626_), .ZN(new_n13627_));
  XOR2_X1    g13435(.A1(new_n13627_), .A2(new_n13164_), .Z(new_n13628_));
  AOI21_X1   g13436(.A1(new_n13334_), .A2(new_n13338_), .B(\asqrt[12] ), .ZN(new_n13629_));
  XOR2_X1    g13437(.A1(new_n13629_), .A2(new_n13167_), .Z(new_n13630_));
  INV_X1     g13438(.I(new_n13630_), .ZN(new_n13631_));
  AOI21_X1   g13439(.A1(new_n13320_), .A2(new_n13328_), .B(\asqrt[12] ), .ZN(new_n13632_));
  XOR2_X1    g13440(.A1(new_n13632_), .A2(new_n13171_), .Z(new_n13633_));
  INV_X1     g13441(.I(new_n13633_), .ZN(new_n13634_));
  XOR2_X1    g13442(.A1(new_n13311_), .A2(\asqrt[27] ), .Z(new_n13635_));
  NOR2_X1    g13443(.A1(\asqrt[12] ), .A2(new_n13635_), .ZN(new_n13636_));
  XOR2_X1    g13444(.A1(new_n13636_), .A2(new_n13173_), .Z(new_n13637_));
  NOR2_X1    g13445(.A1(new_n13309_), .A2(new_n13318_), .ZN(new_n13638_));
  NOR2_X1    g13446(.A1(\asqrt[12] ), .A2(new_n13638_), .ZN(new_n13639_));
  XOR2_X1    g13447(.A1(new_n13639_), .A2(new_n13176_), .Z(new_n13640_));
  AOI21_X1   g13448(.A1(new_n13313_), .A2(new_n13317_), .B(\asqrt[12] ), .ZN(new_n13641_));
  XOR2_X1    g13449(.A1(new_n13641_), .A2(new_n13179_), .Z(new_n13642_));
  INV_X1     g13450(.I(new_n13642_), .ZN(new_n13643_));
  AOI21_X1   g13451(.A1(new_n13299_), .A2(new_n13307_), .B(\asqrt[12] ), .ZN(new_n13644_));
  XOR2_X1    g13452(.A1(new_n13644_), .A2(new_n13183_), .Z(new_n13645_));
  INV_X1     g13453(.I(new_n13645_), .ZN(new_n13646_));
  XOR2_X1    g13454(.A1(new_n13290_), .A2(\asqrt[23] ), .Z(new_n13647_));
  NOR2_X1    g13455(.A1(\asqrt[12] ), .A2(new_n13647_), .ZN(new_n13648_));
  XOR2_X1    g13456(.A1(new_n13648_), .A2(new_n13185_), .Z(new_n13649_));
  NOR2_X1    g13457(.A1(new_n13288_), .A2(new_n13297_), .ZN(new_n13650_));
  NOR2_X1    g13458(.A1(\asqrt[12] ), .A2(new_n13650_), .ZN(new_n13651_));
  XOR2_X1    g13459(.A1(new_n13651_), .A2(new_n13188_), .Z(new_n13652_));
  AOI21_X1   g13460(.A1(new_n13292_), .A2(new_n13296_), .B(\asqrt[12] ), .ZN(new_n13653_));
  XOR2_X1    g13461(.A1(new_n13653_), .A2(new_n13191_), .Z(new_n13654_));
  INV_X1     g13462(.I(new_n13654_), .ZN(new_n13655_));
  AOI21_X1   g13463(.A1(new_n13278_), .A2(new_n13286_), .B(\asqrt[12] ), .ZN(new_n13656_));
  XOR2_X1    g13464(.A1(new_n13656_), .A2(new_n13195_), .Z(new_n13657_));
  INV_X1     g13465(.I(new_n13657_), .ZN(new_n13658_));
  XOR2_X1    g13466(.A1(new_n13269_), .A2(\asqrt[19] ), .Z(new_n13659_));
  NOR2_X1    g13467(.A1(\asqrt[12] ), .A2(new_n13659_), .ZN(new_n13660_));
  XOR2_X1    g13468(.A1(new_n13660_), .A2(new_n13197_), .Z(new_n13661_));
  NOR2_X1    g13469(.A1(new_n13267_), .A2(new_n13276_), .ZN(new_n13662_));
  NOR2_X1    g13470(.A1(\asqrt[12] ), .A2(new_n13662_), .ZN(new_n13663_));
  XOR2_X1    g13471(.A1(new_n13663_), .A2(new_n13200_), .Z(new_n13664_));
  AOI21_X1   g13472(.A1(new_n13271_), .A2(new_n13275_), .B(\asqrt[12] ), .ZN(new_n13665_));
  XOR2_X1    g13473(.A1(new_n13665_), .A2(new_n13203_), .Z(new_n13666_));
  INV_X1     g13474(.I(new_n13666_), .ZN(new_n13667_));
  AOI21_X1   g13475(.A1(new_n13257_), .A2(new_n13265_), .B(\asqrt[12] ), .ZN(new_n13668_));
  XOR2_X1    g13476(.A1(new_n13668_), .A2(new_n13210_), .Z(new_n13669_));
  INV_X1     g13477(.I(new_n13669_), .ZN(new_n13670_));
  AOI21_X1   g13478(.A1(new_n13247_), .A2(new_n13256_), .B(\asqrt[12] ), .ZN(new_n13671_));
  XOR2_X1    g13479(.A1(new_n13671_), .A2(new_n13231_), .Z(new_n13672_));
  NAND2_X1   g13480(.A1(\asqrt[13] ), .A2(new_n13232_), .ZN(new_n13673_));
  NOR2_X1    g13481(.A1(new_n13244_), .A2(\a[26] ), .ZN(new_n13674_));
  AOI22_X1   g13482(.A1(new_n13673_), .A2(new_n13244_), .B1(\asqrt[13] ), .B2(new_n13674_), .ZN(new_n13675_));
  OAI21_X1   g13483(.A1(new_n13228_), .A2(new_n13232_), .B(new_n13241_), .ZN(new_n13676_));
  AOI21_X1   g13484(.A1(new_n13237_), .A2(new_n13676_), .B(\asqrt[12] ), .ZN(new_n13677_));
  XOR2_X1    g13485(.A1(new_n13677_), .A2(new_n13675_), .Z(new_n13678_));
  NAND2_X1   g13486(.A1(new_n13549_), .A2(new_n193_), .ZN(new_n13679_));
  NOR2_X1    g13487(.A1(new_n13539_), .A2(new_n13535_), .ZN(new_n13680_));
  AOI21_X1   g13488(.A1(new_n13680_), .A2(new_n201_), .B(new_n13544_), .ZN(new_n13681_));
  OAI21_X1   g13489(.A1(new_n13680_), .A2(new_n201_), .B(new_n13456_), .ZN(new_n13682_));
  NOR2_X1    g13490(.A1(new_n13681_), .A2(new_n13682_), .ZN(new_n13683_));
  NAND3_X1   g13491(.A1(new_n13555_), .A2(\asqrt[13] ), .A3(new_n13557_), .ZN(new_n13684_));
  NOR3_X1    g13492(.A1(new_n13679_), .A2(new_n13683_), .A3(new_n13684_), .ZN(new_n13685_));
  AOI21_X1   g13493(.A1(new_n13533_), .A2(new_n13526_), .B(\asqrt[62] ), .ZN(new_n13686_));
  NOR3_X1    g13494(.A1(new_n13539_), .A2(new_n201_), .A3(new_n13535_), .ZN(new_n13687_));
  OAI22_X1   g13495(.A1(new_n13687_), .A2(new_n13686_), .B1(new_n13680_), .B2(new_n13543_), .ZN(new_n13688_));
  AOI21_X1   g13496(.A1(new_n13688_), .A2(new_n13455_), .B(new_n13547_), .ZN(new_n13689_));
  NOR4_X1    g13497(.A1(new_n13689_), .A2(\asqrt[63] ), .A3(new_n13683_), .A4(new_n13558_), .ZN(new_n13690_));
  NOR2_X1    g13498(.A1(new_n13690_), .A2(new_n13235_), .ZN(new_n13691_));
  OAI21_X1   g13499(.A1(new_n13691_), .A2(new_n13685_), .B(new_n13232_), .ZN(new_n13692_));
  NOR3_X1    g13500(.A1(new_n13689_), .A2(\asqrt[63] ), .A3(new_n13683_), .ZN(new_n13693_));
  NAND4_X1   g13501(.A1(new_n13693_), .A2(\asqrt[13] ), .A3(new_n13555_), .A4(new_n13557_), .ZN(new_n13694_));
  NAND2_X1   g13502(.A1(\asqrt[12] ), .A2(new_n13233_), .ZN(new_n13695_));
  NAND3_X1   g13503(.A1(new_n13694_), .A2(new_n13695_), .A3(\a[26] ), .ZN(new_n13696_));
  NAND2_X1   g13504(.A1(new_n13696_), .A2(new_n13692_), .ZN(new_n13697_));
  NOR2_X1    g13505(.A1(\a[22] ), .A2(\a[23] ), .ZN(new_n13698_));
  INV_X1     g13506(.I(new_n13698_), .ZN(new_n13699_));
  NAND3_X1   g13507(.A1(\asqrt[12] ), .A2(\a[24] ), .A3(new_n13699_), .ZN(new_n13700_));
  INV_X1     g13508(.I(\a[24] ), .ZN(new_n13701_));
  OAI21_X1   g13509(.A1(\asqrt[12] ), .A2(new_n13701_), .B(new_n13698_), .ZN(new_n13702_));
  AOI21_X1   g13510(.A1(new_n13702_), .A2(new_n13700_), .B(new_n13228_), .ZN(new_n13703_));
  NAND2_X1   g13511(.A1(new_n13698_), .A2(new_n13701_), .ZN(new_n13704_));
  NAND3_X1   g13512(.A1(new_n13092_), .A2(new_n13094_), .A3(new_n13704_), .ZN(new_n13705_));
  NAND2_X1   g13513(.A1(new_n13220_), .A2(new_n13705_), .ZN(new_n13706_));
  NAND3_X1   g13514(.A1(\asqrt[12] ), .A2(\a[24] ), .A3(new_n13706_), .ZN(new_n13707_));
  INV_X1     g13515(.I(\a[25] ), .ZN(new_n13708_));
  NAND3_X1   g13516(.A1(\asqrt[12] ), .A2(new_n13701_), .A3(new_n13708_), .ZN(new_n13709_));
  OAI21_X1   g13517(.A1(new_n13690_), .A2(\a[24] ), .B(\a[25] ), .ZN(new_n13710_));
  NAND3_X1   g13518(.A1(new_n13710_), .A2(new_n13707_), .A3(new_n13709_), .ZN(new_n13711_));
  NOR3_X1    g13519(.A1(new_n13711_), .A2(new_n13703_), .A3(\asqrt[14] ), .ZN(new_n13712_));
  OAI21_X1   g13520(.A1(new_n13711_), .A2(new_n13703_), .B(\asqrt[14] ), .ZN(new_n13713_));
  OAI21_X1   g13521(.A1(new_n13697_), .A2(new_n13712_), .B(new_n13713_), .ZN(new_n13714_));
  OAI21_X1   g13522(.A1(new_n13714_), .A2(\asqrt[15] ), .B(new_n13678_), .ZN(new_n13715_));
  NAND2_X1   g13523(.A1(new_n13714_), .A2(\asqrt[15] ), .ZN(new_n13716_));
  NAND3_X1   g13524(.A1(new_n13715_), .A2(new_n13716_), .A3(new_n11802_), .ZN(new_n13717_));
  AOI21_X1   g13525(.A1(new_n13715_), .A2(new_n13716_), .B(new_n11802_), .ZN(new_n13718_));
  AOI21_X1   g13526(.A1(new_n13672_), .A2(new_n13717_), .B(new_n13718_), .ZN(new_n13719_));
  AOI21_X1   g13527(.A1(new_n13719_), .A2(new_n11373_), .B(new_n13670_), .ZN(new_n13720_));
  NAND2_X1   g13528(.A1(new_n13717_), .A2(new_n13672_), .ZN(new_n13721_));
  INV_X1     g13529(.I(new_n13678_), .ZN(new_n13722_));
  INV_X1     g13530(.I(new_n13697_), .ZN(new_n13723_));
  NOR3_X1    g13531(.A1(new_n13690_), .A2(new_n13701_), .A3(new_n13698_), .ZN(new_n13724_));
  AOI21_X1   g13532(.A1(new_n13690_), .A2(\a[24] ), .B(new_n13699_), .ZN(new_n13725_));
  OAI21_X1   g13533(.A1(new_n13724_), .A2(new_n13725_), .B(\asqrt[13] ), .ZN(new_n13726_));
  INV_X1     g13534(.I(new_n13706_), .ZN(new_n13727_));
  NOR3_X1    g13535(.A1(new_n13690_), .A2(new_n13701_), .A3(new_n13727_), .ZN(new_n13728_));
  NOR3_X1    g13536(.A1(new_n13690_), .A2(\a[24] ), .A3(\a[25] ), .ZN(new_n13729_));
  AOI21_X1   g13537(.A1(\asqrt[12] ), .A2(new_n13701_), .B(new_n13708_), .ZN(new_n13730_));
  NOR3_X1    g13538(.A1(new_n13728_), .A2(new_n13729_), .A3(new_n13730_), .ZN(new_n13731_));
  NAND3_X1   g13539(.A1(new_n13726_), .A2(new_n13731_), .A3(new_n12733_), .ZN(new_n13732_));
  AOI21_X1   g13540(.A1(new_n13726_), .A2(new_n13731_), .B(new_n12733_), .ZN(new_n13733_));
  AOI21_X1   g13541(.A1(new_n13723_), .A2(new_n13732_), .B(new_n13733_), .ZN(new_n13734_));
  AOI21_X1   g13542(.A1(new_n13734_), .A2(new_n12283_), .B(new_n13722_), .ZN(new_n13735_));
  NAND2_X1   g13543(.A1(new_n13723_), .A2(new_n13732_), .ZN(new_n13736_));
  AOI21_X1   g13544(.A1(new_n13736_), .A2(new_n13713_), .B(new_n12283_), .ZN(new_n13737_));
  OAI21_X1   g13545(.A1(new_n13735_), .A2(new_n13737_), .B(\asqrt[16] ), .ZN(new_n13738_));
  AOI21_X1   g13546(.A1(new_n13721_), .A2(new_n13738_), .B(new_n11373_), .ZN(new_n13739_));
  NOR3_X1    g13547(.A1(new_n13720_), .A2(\asqrt[18] ), .A3(new_n13739_), .ZN(new_n13740_));
  OAI21_X1   g13548(.A1(new_n13720_), .A2(new_n13739_), .B(\asqrt[18] ), .ZN(new_n13741_));
  OAI21_X1   g13549(.A1(new_n13667_), .A2(new_n13740_), .B(new_n13741_), .ZN(new_n13742_));
  OAI21_X1   g13550(.A1(new_n13742_), .A2(\asqrt[19] ), .B(new_n13664_), .ZN(new_n13743_));
  NAND2_X1   g13551(.A1(new_n13742_), .A2(\asqrt[19] ), .ZN(new_n13744_));
  NAND3_X1   g13552(.A1(new_n13743_), .A2(new_n13744_), .A3(new_n10052_), .ZN(new_n13745_));
  AOI21_X1   g13553(.A1(new_n13743_), .A2(new_n13744_), .B(new_n10052_), .ZN(new_n13746_));
  AOI21_X1   g13554(.A1(new_n13661_), .A2(new_n13745_), .B(new_n13746_), .ZN(new_n13747_));
  AOI21_X1   g13555(.A1(new_n13747_), .A2(new_n9656_), .B(new_n13658_), .ZN(new_n13748_));
  NAND2_X1   g13556(.A1(new_n13745_), .A2(new_n13661_), .ZN(new_n13749_));
  INV_X1     g13557(.I(new_n13664_), .ZN(new_n13750_));
  INV_X1     g13558(.I(new_n13672_), .ZN(new_n13751_));
  NOR3_X1    g13559(.A1(new_n13735_), .A2(\asqrt[16] ), .A3(new_n13737_), .ZN(new_n13752_));
  OAI21_X1   g13560(.A1(new_n13751_), .A2(new_n13752_), .B(new_n13738_), .ZN(new_n13753_));
  OAI21_X1   g13561(.A1(new_n13753_), .A2(\asqrt[17] ), .B(new_n13669_), .ZN(new_n13754_));
  NAND2_X1   g13562(.A1(new_n13753_), .A2(\asqrt[17] ), .ZN(new_n13755_));
  NAND3_X1   g13563(.A1(new_n13754_), .A2(new_n13755_), .A3(new_n10914_), .ZN(new_n13756_));
  AOI21_X1   g13564(.A1(new_n13754_), .A2(new_n13755_), .B(new_n10914_), .ZN(new_n13757_));
  AOI21_X1   g13565(.A1(new_n13666_), .A2(new_n13756_), .B(new_n13757_), .ZN(new_n13758_));
  AOI21_X1   g13566(.A1(new_n13758_), .A2(new_n10497_), .B(new_n13750_), .ZN(new_n13759_));
  NAND2_X1   g13567(.A1(new_n13756_), .A2(new_n13666_), .ZN(new_n13760_));
  AOI21_X1   g13568(.A1(new_n13760_), .A2(new_n13741_), .B(new_n10497_), .ZN(new_n13761_));
  OAI21_X1   g13569(.A1(new_n13759_), .A2(new_n13761_), .B(\asqrt[20] ), .ZN(new_n13762_));
  AOI21_X1   g13570(.A1(new_n13749_), .A2(new_n13762_), .B(new_n9656_), .ZN(new_n13763_));
  NOR3_X1    g13571(.A1(new_n13748_), .A2(\asqrt[22] ), .A3(new_n13763_), .ZN(new_n13764_));
  OAI21_X1   g13572(.A1(new_n13748_), .A2(new_n13763_), .B(\asqrt[22] ), .ZN(new_n13765_));
  OAI21_X1   g13573(.A1(new_n13655_), .A2(new_n13764_), .B(new_n13765_), .ZN(new_n13766_));
  OAI21_X1   g13574(.A1(new_n13766_), .A2(\asqrt[23] ), .B(new_n13652_), .ZN(new_n13767_));
  NAND2_X1   g13575(.A1(new_n13766_), .A2(\asqrt[23] ), .ZN(new_n13768_));
  NAND3_X1   g13576(.A1(new_n13767_), .A2(new_n13768_), .A3(new_n8440_), .ZN(new_n13769_));
  AOI21_X1   g13577(.A1(new_n13767_), .A2(new_n13768_), .B(new_n8440_), .ZN(new_n13770_));
  AOI21_X1   g13578(.A1(new_n13649_), .A2(new_n13769_), .B(new_n13770_), .ZN(new_n13771_));
  AOI21_X1   g13579(.A1(new_n13771_), .A2(new_n8077_), .B(new_n13646_), .ZN(new_n13772_));
  NAND2_X1   g13580(.A1(new_n13769_), .A2(new_n13649_), .ZN(new_n13773_));
  INV_X1     g13581(.I(new_n13652_), .ZN(new_n13774_));
  INV_X1     g13582(.I(new_n13661_), .ZN(new_n13775_));
  NOR3_X1    g13583(.A1(new_n13759_), .A2(\asqrt[20] ), .A3(new_n13761_), .ZN(new_n13776_));
  OAI21_X1   g13584(.A1(new_n13775_), .A2(new_n13776_), .B(new_n13762_), .ZN(new_n13777_));
  OAI21_X1   g13585(.A1(new_n13777_), .A2(\asqrt[21] ), .B(new_n13657_), .ZN(new_n13778_));
  NAND2_X1   g13586(.A1(new_n13777_), .A2(\asqrt[21] ), .ZN(new_n13779_));
  NAND3_X1   g13587(.A1(new_n13778_), .A2(new_n13779_), .A3(new_n9233_), .ZN(new_n13780_));
  AOI21_X1   g13588(.A1(new_n13778_), .A2(new_n13779_), .B(new_n9233_), .ZN(new_n13781_));
  AOI21_X1   g13589(.A1(new_n13654_), .A2(new_n13780_), .B(new_n13781_), .ZN(new_n13782_));
  AOI21_X1   g13590(.A1(new_n13782_), .A2(new_n8849_), .B(new_n13774_), .ZN(new_n13783_));
  NAND2_X1   g13591(.A1(new_n13780_), .A2(new_n13654_), .ZN(new_n13784_));
  AOI21_X1   g13592(.A1(new_n13784_), .A2(new_n13765_), .B(new_n8849_), .ZN(new_n13785_));
  OAI21_X1   g13593(.A1(new_n13783_), .A2(new_n13785_), .B(\asqrt[24] ), .ZN(new_n13786_));
  AOI21_X1   g13594(.A1(new_n13773_), .A2(new_n13786_), .B(new_n8077_), .ZN(new_n13787_));
  NOR3_X1    g13595(.A1(new_n13772_), .A2(\asqrt[26] ), .A3(new_n13787_), .ZN(new_n13788_));
  OAI21_X1   g13596(.A1(new_n13772_), .A2(new_n13787_), .B(\asqrt[26] ), .ZN(new_n13789_));
  OAI21_X1   g13597(.A1(new_n13643_), .A2(new_n13788_), .B(new_n13789_), .ZN(new_n13790_));
  OAI21_X1   g13598(.A1(new_n13790_), .A2(\asqrt[27] ), .B(new_n13640_), .ZN(new_n13791_));
  NAND2_X1   g13599(.A1(new_n13790_), .A2(\asqrt[27] ), .ZN(new_n13792_));
  NAND3_X1   g13600(.A1(new_n13791_), .A2(new_n13792_), .A3(new_n6966_), .ZN(new_n13793_));
  AOI21_X1   g13601(.A1(new_n13791_), .A2(new_n13792_), .B(new_n6966_), .ZN(new_n13794_));
  AOI21_X1   g13602(.A1(new_n13637_), .A2(new_n13793_), .B(new_n13794_), .ZN(new_n13795_));
  AOI21_X1   g13603(.A1(new_n13795_), .A2(new_n6636_), .B(new_n13634_), .ZN(new_n13796_));
  NAND2_X1   g13604(.A1(new_n13793_), .A2(new_n13637_), .ZN(new_n13797_));
  INV_X1     g13605(.I(new_n13640_), .ZN(new_n13798_));
  INV_X1     g13606(.I(new_n13649_), .ZN(new_n13799_));
  NOR3_X1    g13607(.A1(new_n13783_), .A2(\asqrt[24] ), .A3(new_n13785_), .ZN(new_n13800_));
  OAI21_X1   g13608(.A1(new_n13799_), .A2(new_n13800_), .B(new_n13786_), .ZN(new_n13801_));
  OAI21_X1   g13609(.A1(new_n13801_), .A2(\asqrt[25] ), .B(new_n13645_), .ZN(new_n13802_));
  NAND2_X1   g13610(.A1(new_n13801_), .A2(\asqrt[25] ), .ZN(new_n13803_));
  NAND3_X1   g13611(.A1(new_n13802_), .A2(new_n13803_), .A3(new_n7690_), .ZN(new_n13804_));
  AOI21_X1   g13612(.A1(new_n13802_), .A2(new_n13803_), .B(new_n7690_), .ZN(new_n13805_));
  AOI21_X1   g13613(.A1(new_n13642_), .A2(new_n13804_), .B(new_n13805_), .ZN(new_n13806_));
  AOI21_X1   g13614(.A1(new_n13806_), .A2(new_n7331_), .B(new_n13798_), .ZN(new_n13807_));
  NAND2_X1   g13615(.A1(new_n13804_), .A2(new_n13642_), .ZN(new_n13808_));
  AOI21_X1   g13616(.A1(new_n13808_), .A2(new_n13789_), .B(new_n7331_), .ZN(new_n13809_));
  OAI21_X1   g13617(.A1(new_n13807_), .A2(new_n13809_), .B(\asqrt[28] ), .ZN(new_n13810_));
  AOI21_X1   g13618(.A1(new_n13797_), .A2(new_n13810_), .B(new_n6636_), .ZN(new_n13811_));
  NOR3_X1    g13619(.A1(new_n13796_), .A2(\asqrt[30] ), .A3(new_n13811_), .ZN(new_n13812_));
  OAI21_X1   g13620(.A1(new_n13796_), .A2(new_n13811_), .B(\asqrt[30] ), .ZN(new_n13813_));
  OAI21_X1   g13621(.A1(new_n13631_), .A2(new_n13812_), .B(new_n13813_), .ZN(new_n13814_));
  OAI21_X1   g13622(.A1(new_n13814_), .A2(\asqrt[31] ), .B(new_n13628_), .ZN(new_n13815_));
  NAND2_X1   g13623(.A1(new_n13814_), .A2(\asqrt[31] ), .ZN(new_n13816_));
  NAND3_X1   g13624(.A1(new_n13815_), .A2(new_n13816_), .A3(new_n5643_), .ZN(new_n13817_));
  AOI21_X1   g13625(.A1(new_n13815_), .A2(new_n13816_), .B(new_n5643_), .ZN(new_n13818_));
  AOI21_X1   g13626(.A1(new_n13625_), .A2(new_n13817_), .B(new_n13818_), .ZN(new_n13819_));
  AOI21_X1   g13627(.A1(new_n13819_), .A2(new_n5336_), .B(new_n13622_), .ZN(new_n13820_));
  NAND2_X1   g13628(.A1(new_n13817_), .A2(new_n13625_), .ZN(new_n13821_));
  INV_X1     g13629(.I(new_n13628_), .ZN(new_n13822_));
  INV_X1     g13630(.I(new_n13637_), .ZN(new_n13823_));
  NOR3_X1    g13631(.A1(new_n13807_), .A2(\asqrt[28] ), .A3(new_n13809_), .ZN(new_n13824_));
  OAI21_X1   g13632(.A1(new_n13823_), .A2(new_n13824_), .B(new_n13810_), .ZN(new_n13825_));
  OAI21_X1   g13633(.A1(new_n13825_), .A2(\asqrt[29] ), .B(new_n13633_), .ZN(new_n13826_));
  NAND2_X1   g13634(.A1(new_n13825_), .A2(\asqrt[29] ), .ZN(new_n13827_));
  NAND3_X1   g13635(.A1(new_n13826_), .A2(new_n13827_), .A3(new_n6275_), .ZN(new_n13828_));
  AOI21_X1   g13636(.A1(new_n13826_), .A2(new_n13827_), .B(new_n6275_), .ZN(new_n13829_));
  AOI21_X1   g13637(.A1(new_n13630_), .A2(new_n13828_), .B(new_n13829_), .ZN(new_n13830_));
  AOI21_X1   g13638(.A1(new_n13830_), .A2(new_n5947_), .B(new_n13822_), .ZN(new_n13831_));
  NAND2_X1   g13639(.A1(new_n13828_), .A2(new_n13630_), .ZN(new_n13832_));
  AOI21_X1   g13640(.A1(new_n13832_), .A2(new_n13813_), .B(new_n5947_), .ZN(new_n13833_));
  OAI21_X1   g13641(.A1(new_n13831_), .A2(new_n13833_), .B(\asqrt[32] ), .ZN(new_n13834_));
  AOI21_X1   g13642(.A1(new_n13821_), .A2(new_n13834_), .B(new_n5336_), .ZN(new_n13835_));
  NOR3_X1    g13643(.A1(new_n13820_), .A2(\asqrt[34] ), .A3(new_n13835_), .ZN(new_n13836_));
  OAI21_X1   g13644(.A1(new_n13820_), .A2(new_n13835_), .B(\asqrt[34] ), .ZN(new_n13837_));
  OAI21_X1   g13645(.A1(new_n13619_), .A2(new_n13836_), .B(new_n13837_), .ZN(new_n13838_));
  OAI21_X1   g13646(.A1(new_n13838_), .A2(\asqrt[35] ), .B(new_n13616_), .ZN(new_n13839_));
  NAND2_X1   g13647(.A1(new_n13838_), .A2(\asqrt[35] ), .ZN(new_n13840_));
  NAND3_X1   g13648(.A1(new_n13839_), .A2(new_n13840_), .A3(new_n4461_), .ZN(new_n13841_));
  AOI21_X1   g13649(.A1(new_n13839_), .A2(new_n13840_), .B(new_n4461_), .ZN(new_n13842_));
  AOI21_X1   g13650(.A1(new_n13613_), .A2(new_n13841_), .B(new_n13842_), .ZN(new_n13843_));
  AOI21_X1   g13651(.A1(new_n13843_), .A2(new_n4196_), .B(new_n13610_), .ZN(new_n13844_));
  NAND2_X1   g13652(.A1(new_n13841_), .A2(new_n13613_), .ZN(new_n13845_));
  INV_X1     g13653(.I(new_n13616_), .ZN(new_n13846_));
  INV_X1     g13654(.I(new_n13625_), .ZN(new_n13847_));
  NOR3_X1    g13655(.A1(new_n13831_), .A2(\asqrt[32] ), .A3(new_n13833_), .ZN(new_n13848_));
  OAI21_X1   g13656(.A1(new_n13847_), .A2(new_n13848_), .B(new_n13834_), .ZN(new_n13849_));
  OAI21_X1   g13657(.A1(new_n13849_), .A2(\asqrt[33] ), .B(new_n13621_), .ZN(new_n13850_));
  NAND2_X1   g13658(.A1(new_n13849_), .A2(\asqrt[33] ), .ZN(new_n13851_));
  NAND3_X1   g13659(.A1(new_n13850_), .A2(new_n13851_), .A3(new_n5029_), .ZN(new_n13852_));
  AOI21_X1   g13660(.A1(new_n13850_), .A2(new_n13851_), .B(new_n5029_), .ZN(new_n13853_));
  AOI21_X1   g13661(.A1(new_n13618_), .A2(new_n13852_), .B(new_n13853_), .ZN(new_n13854_));
  AOI21_X1   g13662(.A1(new_n13854_), .A2(new_n4751_), .B(new_n13846_), .ZN(new_n13855_));
  NAND2_X1   g13663(.A1(new_n13852_), .A2(new_n13618_), .ZN(new_n13856_));
  AOI21_X1   g13664(.A1(new_n13856_), .A2(new_n13837_), .B(new_n4751_), .ZN(new_n13857_));
  OAI21_X1   g13665(.A1(new_n13855_), .A2(new_n13857_), .B(\asqrt[36] ), .ZN(new_n13858_));
  AOI21_X1   g13666(.A1(new_n13845_), .A2(new_n13858_), .B(new_n4196_), .ZN(new_n13859_));
  NOR3_X1    g13667(.A1(new_n13844_), .A2(\asqrt[38] ), .A3(new_n13859_), .ZN(new_n13860_));
  OAI21_X1   g13668(.A1(new_n13844_), .A2(new_n13859_), .B(\asqrt[38] ), .ZN(new_n13861_));
  OAI21_X1   g13669(.A1(new_n13607_), .A2(new_n13860_), .B(new_n13861_), .ZN(new_n13862_));
  OAI21_X1   g13670(.A1(new_n13862_), .A2(\asqrt[39] ), .B(new_n13604_), .ZN(new_n13863_));
  NAND2_X1   g13671(.A1(new_n13862_), .A2(\asqrt[39] ), .ZN(new_n13864_));
  NAND3_X1   g13672(.A1(new_n13863_), .A2(new_n13864_), .A3(new_n3427_), .ZN(new_n13865_));
  AOI21_X1   g13673(.A1(new_n13863_), .A2(new_n13864_), .B(new_n3427_), .ZN(new_n13866_));
  AOI21_X1   g13674(.A1(new_n13601_), .A2(new_n13865_), .B(new_n13866_), .ZN(new_n13867_));
  AOI21_X1   g13675(.A1(new_n13867_), .A2(new_n3195_), .B(new_n13598_), .ZN(new_n13868_));
  NAND2_X1   g13676(.A1(new_n13865_), .A2(new_n13601_), .ZN(new_n13869_));
  INV_X1     g13677(.I(new_n13604_), .ZN(new_n13870_));
  INV_X1     g13678(.I(new_n13613_), .ZN(new_n13871_));
  NOR3_X1    g13679(.A1(new_n13855_), .A2(\asqrt[36] ), .A3(new_n13857_), .ZN(new_n13872_));
  OAI21_X1   g13680(.A1(new_n13871_), .A2(new_n13872_), .B(new_n13858_), .ZN(new_n13873_));
  OAI21_X1   g13681(.A1(new_n13873_), .A2(\asqrt[37] ), .B(new_n13609_), .ZN(new_n13874_));
  NAND2_X1   g13682(.A1(new_n13873_), .A2(\asqrt[37] ), .ZN(new_n13875_));
  NAND3_X1   g13683(.A1(new_n13874_), .A2(new_n13875_), .A3(new_n3925_), .ZN(new_n13876_));
  AOI21_X1   g13684(.A1(new_n13874_), .A2(new_n13875_), .B(new_n3925_), .ZN(new_n13877_));
  AOI21_X1   g13685(.A1(new_n13606_), .A2(new_n13876_), .B(new_n13877_), .ZN(new_n13878_));
  AOI21_X1   g13686(.A1(new_n13878_), .A2(new_n3681_), .B(new_n13870_), .ZN(new_n13879_));
  NAND2_X1   g13687(.A1(new_n13876_), .A2(new_n13606_), .ZN(new_n13880_));
  AOI21_X1   g13688(.A1(new_n13880_), .A2(new_n13861_), .B(new_n3681_), .ZN(new_n13881_));
  OAI21_X1   g13689(.A1(new_n13879_), .A2(new_n13881_), .B(\asqrt[40] ), .ZN(new_n13882_));
  AOI21_X1   g13690(.A1(new_n13869_), .A2(new_n13882_), .B(new_n3195_), .ZN(new_n13883_));
  NOR3_X1    g13691(.A1(new_n13868_), .A2(\asqrt[42] ), .A3(new_n13883_), .ZN(new_n13884_));
  OAI21_X1   g13692(.A1(new_n13868_), .A2(new_n13883_), .B(\asqrt[42] ), .ZN(new_n13885_));
  OAI21_X1   g13693(.A1(new_n13595_), .A2(new_n13884_), .B(new_n13885_), .ZN(new_n13886_));
  OAI21_X1   g13694(.A1(new_n13886_), .A2(\asqrt[43] ), .B(new_n13592_), .ZN(new_n13887_));
  NAND2_X1   g13695(.A1(new_n13886_), .A2(\asqrt[43] ), .ZN(new_n13888_));
  NAND3_X1   g13696(.A1(new_n13887_), .A2(new_n13888_), .A3(new_n2531_), .ZN(new_n13889_));
  AOI21_X1   g13697(.A1(new_n13887_), .A2(new_n13888_), .B(new_n2531_), .ZN(new_n13890_));
  AOI21_X1   g13698(.A1(new_n13589_), .A2(new_n13889_), .B(new_n13890_), .ZN(new_n13891_));
  AOI21_X1   g13699(.A1(new_n13891_), .A2(new_n2332_), .B(new_n13586_), .ZN(new_n13892_));
  NAND2_X1   g13700(.A1(new_n13889_), .A2(new_n13589_), .ZN(new_n13893_));
  INV_X1     g13701(.I(new_n13592_), .ZN(new_n13894_));
  INV_X1     g13702(.I(new_n13601_), .ZN(new_n13895_));
  NOR3_X1    g13703(.A1(new_n13879_), .A2(\asqrt[40] ), .A3(new_n13881_), .ZN(new_n13896_));
  OAI21_X1   g13704(.A1(new_n13895_), .A2(new_n13896_), .B(new_n13882_), .ZN(new_n13897_));
  OAI21_X1   g13705(.A1(new_n13897_), .A2(\asqrt[41] ), .B(new_n13597_), .ZN(new_n13898_));
  NAND2_X1   g13706(.A1(new_n13897_), .A2(\asqrt[41] ), .ZN(new_n13899_));
  NAND3_X1   g13707(.A1(new_n13898_), .A2(new_n13899_), .A3(new_n2960_), .ZN(new_n13900_));
  AOI21_X1   g13708(.A1(new_n13898_), .A2(new_n13899_), .B(new_n2960_), .ZN(new_n13901_));
  AOI21_X1   g13709(.A1(new_n13594_), .A2(new_n13900_), .B(new_n13901_), .ZN(new_n13902_));
  AOI21_X1   g13710(.A1(new_n13902_), .A2(new_n2749_), .B(new_n13894_), .ZN(new_n13903_));
  NAND2_X1   g13711(.A1(new_n13900_), .A2(new_n13594_), .ZN(new_n13904_));
  AOI21_X1   g13712(.A1(new_n13904_), .A2(new_n13885_), .B(new_n2749_), .ZN(new_n13905_));
  OAI21_X1   g13713(.A1(new_n13903_), .A2(new_n13905_), .B(\asqrt[44] ), .ZN(new_n13906_));
  AOI21_X1   g13714(.A1(new_n13893_), .A2(new_n13906_), .B(new_n2332_), .ZN(new_n13907_));
  NOR3_X1    g13715(.A1(new_n13892_), .A2(\asqrt[46] ), .A3(new_n13907_), .ZN(new_n13908_));
  OAI21_X1   g13716(.A1(new_n13892_), .A2(new_n13907_), .B(\asqrt[46] ), .ZN(new_n13909_));
  OAI21_X1   g13717(.A1(new_n13583_), .A2(new_n13908_), .B(new_n13909_), .ZN(new_n13910_));
  OAI21_X1   g13718(.A1(new_n13910_), .A2(\asqrt[47] ), .B(new_n13580_), .ZN(new_n13911_));
  NAND2_X1   g13719(.A1(new_n13910_), .A2(\asqrt[47] ), .ZN(new_n13912_));
  NAND3_X1   g13720(.A1(new_n13911_), .A2(new_n13912_), .A3(new_n1778_), .ZN(new_n13913_));
  AOI21_X1   g13721(.A1(new_n13911_), .A2(new_n13912_), .B(new_n1778_), .ZN(new_n13914_));
  AOI21_X1   g13722(.A1(new_n13577_), .A2(new_n13913_), .B(new_n13914_), .ZN(new_n13915_));
  AOI21_X1   g13723(.A1(new_n13915_), .A2(new_n1632_), .B(new_n13574_), .ZN(new_n13916_));
  NAND2_X1   g13724(.A1(new_n13913_), .A2(new_n13577_), .ZN(new_n13917_));
  INV_X1     g13725(.I(new_n13580_), .ZN(new_n13918_));
  INV_X1     g13726(.I(new_n13589_), .ZN(new_n13919_));
  NOR3_X1    g13727(.A1(new_n13903_), .A2(\asqrt[44] ), .A3(new_n13905_), .ZN(new_n13920_));
  OAI21_X1   g13728(.A1(new_n13919_), .A2(new_n13920_), .B(new_n13906_), .ZN(new_n13921_));
  OAI21_X1   g13729(.A1(new_n13921_), .A2(\asqrt[45] ), .B(new_n13585_), .ZN(new_n13922_));
  NAND2_X1   g13730(.A1(new_n13921_), .A2(\asqrt[45] ), .ZN(new_n13923_));
  NAND3_X1   g13731(.A1(new_n13922_), .A2(new_n13923_), .A3(new_n2134_), .ZN(new_n13924_));
  AOI21_X1   g13732(.A1(new_n13922_), .A2(new_n13923_), .B(new_n2134_), .ZN(new_n13925_));
  AOI21_X1   g13733(.A1(new_n13582_), .A2(new_n13924_), .B(new_n13925_), .ZN(new_n13926_));
  AOI21_X1   g13734(.A1(new_n13926_), .A2(new_n1953_), .B(new_n13918_), .ZN(new_n13927_));
  NAND2_X1   g13735(.A1(new_n13924_), .A2(new_n13582_), .ZN(new_n13928_));
  AOI21_X1   g13736(.A1(new_n13928_), .A2(new_n13909_), .B(new_n1953_), .ZN(new_n13929_));
  OAI21_X1   g13737(.A1(new_n13927_), .A2(new_n13929_), .B(\asqrt[48] ), .ZN(new_n13930_));
  AOI21_X1   g13738(.A1(new_n13917_), .A2(new_n13930_), .B(new_n1632_), .ZN(new_n13931_));
  NOR3_X1    g13739(.A1(new_n13916_), .A2(\asqrt[50] ), .A3(new_n13931_), .ZN(new_n13932_));
  OAI21_X1   g13740(.A1(new_n13916_), .A2(new_n13931_), .B(\asqrt[50] ), .ZN(new_n13933_));
  OAI21_X1   g13741(.A1(new_n13571_), .A2(new_n13932_), .B(new_n13933_), .ZN(new_n13934_));
  OAI21_X1   g13742(.A1(new_n13934_), .A2(\asqrt[51] ), .B(new_n13568_), .ZN(new_n13935_));
  NAND2_X1   g13743(.A1(new_n13934_), .A2(\asqrt[51] ), .ZN(new_n13936_));
  NAND3_X1   g13744(.A1(new_n13935_), .A2(new_n13936_), .A3(new_n1150_), .ZN(new_n13937_));
  AOI21_X1   g13745(.A1(new_n13935_), .A2(new_n13936_), .B(new_n1150_), .ZN(new_n13938_));
  AOI21_X1   g13746(.A1(new_n13565_), .A2(new_n13937_), .B(new_n13938_), .ZN(new_n13939_));
  NAND2_X1   g13747(.A1(new_n13939_), .A2(new_n1006_), .ZN(new_n13940_));
  INV_X1     g13748(.I(new_n13565_), .ZN(new_n13941_));
  INV_X1     g13749(.I(new_n13568_), .ZN(new_n13942_));
  INV_X1     g13750(.I(new_n13577_), .ZN(new_n13943_));
  NOR3_X1    g13751(.A1(new_n13927_), .A2(\asqrt[48] ), .A3(new_n13929_), .ZN(new_n13944_));
  OAI21_X1   g13752(.A1(new_n13943_), .A2(new_n13944_), .B(new_n13930_), .ZN(new_n13945_));
  OAI21_X1   g13753(.A1(new_n13945_), .A2(\asqrt[49] ), .B(new_n13573_), .ZN(new_n13946_));
  NAND2_X1   g13754(.A1(new_n13945_), .A2(\asqrt[49] ), .ZN(new_n13947_));
  NAND3_X1   g13755(.A1(new_n13946_), .A2(new_n13947_), .A3(new_n1463_), .ZN(new_n13948_));
  AOI21_X1   g13756(.A1(new_n13946_), .A2(new_n13947_), .B(new_n1463_), .ZN(new_n13949_));
  AOI21_X1   g13757(.A1(new_n13570_), .A2(new_n13948_), .B(new_n13949_), .ZN(new_n13950_));
  AOI21_X1   g13758(.A1(new_n13950_), .A2(new_n1305_), .B(new_n13942_), .ZN(new_n13951_));
  NAND2_X1   g13759(.A1(new_n13948_), .A2(new_n13570_), .ZN(new_n13952_));
  AOI21_X1   g13760(.A1(new_n13952_), .A2(new_n13933_), .B(new_n1305_), .ZN(new_n13953_));
  NOR3_X1    g13761(.A1(new_n13951_), .A2(\asqrt[52] ), .A3(new_n13953_), .ZN(new_n13954_));
  OAI21_X1   g13762(.A1(new_n13951_), .A2(new_n13953_), .B(\asqrt[52] ), .ZN(new_n13955_));
  OAI21_X1   g13763(.A1(new_n13941_), .A2(new_n13954_), .B(new_n13955_), .ZN(new_n13956_));
  NAND2_X1   g13764(.A1(new_n13956_), .A2(\asqrt[53] ), .ZN(new_n13957_));
  NOR2_X1    g13765(.A1(new_n13534_), .A2(\asqrt[62] ), .ZN(new_n13958_));
  INV_X1     g13766(.I(new_n13551_), .ZN(new_n13959_));
  NOR2_X1    g13767(.A1(new_n13959_), .A2(new_n13958_), .ZN(new_n13960_));
  XOR2_X1    g13768(.A1(new_n13542_), .A2(new_n13067_), .Z(new_n13961_));
  OAI21_X1   g13769(.A1(\asqrt[12] ), .A2(new_n13960_), .B(new_n13961_), .ZN(new_n13962_));
  INV_X1     g13770(.I(new_n13962_), .ZN(new_n13963_));
  NOR2_X1    g13771(.A1(new_n13505_), .A2(new_n13502_), .ZN(new_n13964_));
  NOR2_X1    g13772(.A1(\asqrt[12] ), .A2(new_n13964_), .ZN(new_n13965_));
  XOR2_X1    g13773(.A1(new_n13965_), .A2(new_n13462_), .Z(new_n13966_));
  INV_X1     g13774(.I(new_n13966_), .ZN(new_n13967_));
  NOR2_X1    g13775(.A1(new_n13521_), .A2(new_n13501_), .ZN(new_n13968_));
  NOR2_X1    g13776(.A1(\asqrt[12] ), .A2(new_n13968_), .ZN(new_n13969_));
  XOR2_X1    g13777(.A1(new_n13969_), .A2(new_n13466_), .Z(new_n13970_));
  AOI21_X1   g13778(.A1(new_n13495_), .A2(new_n13500_), .B(\asqrt[12] ), .ZN(new_n13971_));
  XOR2_X1    g13779(.A1(new_n13971_), .A2(new_n13469_), .Z(new_n13972_));
  AOI21_X1   g13780(.A1(new_n13517_), .A2(new_n13494_), .B(\asqrt[12] ), .ZN(new_n13973_));
  XOR2_X1    g13781(.A1(new_n13973_), .A2(new_n13472_), .Z(new_n13974_));
  INV_X1     g13782(.I(new_n13491_), .ZN(new_n13975_));
  NOR2_X1    g13783(.A1(new_n13975_), .A2(new_n13490_), .ZN(new_n13976_));
  NOR2_X1    g13784(.A1(\asqrt[12] ), .A2(new_n13976_), .ZN(new_n13977_));
  XOR2_X1    g13785(.A1(new_n13977_), .A2(new_n13474_), .Z(new_n13978_));
  INV_X1     g13786(.I(new_n13978_), .ZN(new_n13979_));
  NOR2_X1    g13787(.A1(new_n13513_), .A2(new_n13489_), .ZN(new_n13980_));
  NOR2_X1    g13788(.A1(\asqrt[12] ), .A2(new_n13980_), .ZN(new_n13981_));
  XOR2_X1    g13789(.A1(new_n13981_), .A2(new_n13478_), .Z(new_n13982_));
  INV_X1     g13790(.I(new_n13982_), .ZN(new_n13983_));
  AOI21_X1   g13791(.A1(new_n13483_), .A2(new_n13488_), .B(\asqrt[12] ), .ZN(new_n13984_));
  XOR2_X1    g13792(.A1(new_n13984_), .A2(new_n13481_), .Z(new_n13985_));
  OAI21_X1   g13793(.A1(new_n13956_), .A2(\asqrt[53] ), .B(new_n13562_), .ZN(new_n13986_));
  NAND3_X1   g13794(.A1(new_n13986_), .A2(new_n13957_), .A3(new_n860_), .ZN(new_n13987_));
  AOI21_X1   g13795(.A1(new_n13986_), .A2(new_n13957_), .B(new_n860_), .ZN(new_n13988_));
  AOI21_X1   g13796(.A1(new_n13985_), .A2(new_n13987_), .B(new_n13988_), .ZN(new_n13989_));
  AOI21_X1   g13797(.A1(new_n13989_), .A2(new_n744_), .B(new_n13983_), .ZN(new_n13990_));
  NAND2_X1   g13798(.A1(new_n13987_), .A2(new_n13985_), .ZN(new_n13991_));
  INV_X1     g13799(.I(new_n13562_), .ZN(new_n13992_));
  AOI21_X1   g13800(.A1(new_n13939_), .A2(new_n1006_), .B(new_n13992_), .ZN(new_n13993_));
  NAND2_X1   g13801(.A1(new_n13937_), .A2(new_n13565_), .ZN(new_n13994_));
  AOI21_X1   g13802(.A1(new_n13994_), .A2(new_n13955_), .B(new_n1006_), .ZN(new_n13995_));
  OAI21_X1   g13803(.A1(new_n13993_), .A2(new_n13995_), .B(\asqrt[54] ), .ZN(new_n13996_));
  AOI21_X1   g13804(.A1(new_n13991_), .A2(new_n13996_), .B(new_n744_), .ZN(new_n13997_));
  NOR3_X1    g13805(.A1(new_n13990_), .A2(\asqrt[56] ), .A3(new_n13997_), .ZN(new_n13998_));
  OAI21_X1   g13806(.A1(new_n13990_), .A2(new_n13997_), .B(\asqrt[56] ), .ZN(new_n13999_));
  OAI21_X1   g13807(.A1(new_n13979_), .A2(new_n13998_), .B(new_n13999_), .ZN(new_n14000_));
  OAI21_X1   g13808(.A1(new_n14000_), .A2(\asqrt[57] ), .B(new_n13974_), .ZN(new_n14001_));
  NOR2_X1    g13809(.A1(new_n13998_), .A2(new_n13979_), .ZN(new_n14002_));
  INV_X1     g13810(.I(new_n13985_), .ZN(new_n14003_));
  NOR3_X1    g13811(.A1(new_n13993_), .A2(\asqrt[54] ), .A3(new_n13995_), .ZN(new_n14004_));
  OAI21_X1   g13812(.A1(new_n14003_), .A2(new_n14004_), .B(new_n13996_), .ZN(new_n14005_));
  OAI21_X1   g13813(.A1(new_n14005_), .A2(\asqrt[55] ), .B(new_n13982_), .ZN(new_n14006_));
  NAND2_X1   g13814(.A1(new_n14005_), .A2(\asqrt[55] ), .ZN(new_n14007_));
  AOI21_X1   g13815(.A1(new_n14006_), .A2(new_n14007_), .B(new_n634_), .ZN(new_n14008_));
  OAI21_X1   g13816(.A1(new_n14002_), .A2(new_n14008_), .B(\asqrt[57] ), .ZN(new_n14009_));
  NAND3_X1   g13817(.A1(new_n14001_), .A2(new_n423_), .A3(new_n14009_), .ZN(new_n14010_));
  NAND2_X1   g13818(.A1(new_n14010_), .A2(new_n13972_), .ZN(new_n14011_));
  INV_X1     g13819(.I(new_n13974_), .ZN(new_n14012_));
  NAND3_X1   g13820(.A1(new_n14006_), .A2(new_n14007_), .A3(new_n634_), .ZN(new_n14013_));
  AOI21_X1   g13821(.A1(new_n13978_), .A2(new_n14013_), .B(new_n14008_), .ZN(new_n14014_));
  AOI21_X1   g13822(.A1(new_n14014_), .A2(new_n531_), .B(new_n14012_), .ZN(new_n14015_));
  NAND2_X1   g13823(.A1(new_n14013_), .A2(new_n13978_), .ZN(new_n14016_));
  AOI21_X1   g13824(.A1(new_n14016_), .A2(new_n13999_), .B(new_n531_), .ZN(new_n14017_));
  OAI21_X1   g13825(.A1(new_n14015_), .A2(new_n14017_), .B(\asqrt[58] ), .ZN(new_n14018_));
  NAND3_X1   g13826(.A1(new_n14011_), .A2(new_n337_), .A3(new_n14018_), .ZN(new_n14019_));
  AOI21_X1   g13827(.A1(new_n14011_), .A2(new_n14018_), .B(new_n337_), .ZN(new_n14020_));
  AOI21_X1   g13828(.A1(new_n13970_), .A2(new_n14019_), .B(new_n14020_), .ZN(new_n14021_));
  AOI21_X1   g13829(.A1(new_n14021_), .A2(new_n266_), .B(new_n13967_), .ZN(new_n14022_));
  INV_X1     g13830(.I(new_n13972_), .ZN(new_n14023_));
  NOR3_X1    g13831(.A1(new_n14015_), .A2(\asqrt[58] ), .A3(new_n14017_), .ZN(new_n14024_));
  OAI21_X1   g13832(.A1(new_n14023_), .A2(new_n14024_), .B(new_n14018_), .ZN(new_n14025_));
  OAI21_X1   g13833(.A1(new_n14025_), .A2(\asqrt[59] ), .B(new_n13970_), .ZN(new_n14026_));
  NAND2_X1   g13834(.A1(new_n14025_), .A2(\asqrt[59] ), .ZN(new_n14027_));
  AOI21_X1   g13835(.A1(new_n14026_), .A2(new_n14027_), .B(new_n266_), .ZN(new_n14028_));
  OAI21_X1   g13836(.A1(new_n14022_), .A2(new_n14028_), .B(\asqrt[61] ), .ZN(new_n14029_));
  AOI21_X1   g13837(.A1(new_n13536_), .A2(new_n13531_), .B(\asqrt[12] ), .ZN(new_n14030_));
  XOR2_X1    g13838(.A1(new_n14030_), .A2(new_n13459_), .Z(new_n14031_));
  INV_X1     g13839(.I(new_n14031_), .ZN(new_n14032_));
  NOR3_X1    g13840(.A1(new_n14022_), .A2(\asqrt[61] ), .A3(new_n14028_), .ZN(new_n14033_));
  OAI21_X1   g13841(.A1(new_n14032_), .A2(new_n14033_), .B(new_n14029_), .ZN(new_n14034_));
  NAND3_X1   g13842(.A1(new_n14026_), .A2(new_n14027_), .A3(new_n266_), .ZN(new_n14035_));
  NAND2_X1   g13843(.A1(new_n14035_), .A2(new_n13966_), .ZN(new_n14036_));
  INV_X1     g13844(.I(new_n13970_), .ZN(new_n14037_));
  AOI21_X1   g13845(.A1(new_n14001_), .A2(new_n14009_), .B(new_n423_), .ZN(new_n14038_));
  AOI21_X1   g13846(.A1(new_n13972_), .A2(new_n14010_), .B(new_n14038_), .ZN(new_n14039_));
  AOI21_X1   g13847(.A1(new_n14039_), .A2(new_n337_), .B(new_n14037_), .ZN(new_n14040_));
  OAI21_X1   g13848(.A1(new_n14040_), .A2(new_n14020_), .B(\asqrt[60] ), .ZN(new_n14041_));
  AOI21_X1   g13849(.A1(new_n14036_), .A2(new_n14041_), .B(new_n239_), .ZN(new_n14042_));
  AOI21_X1   g13850(.A1(new_n13966_), .A2(new_n14035_), .B(new_n14028_), .ZN(new_n14043_));
  AOI21_X1   g13851(.A1(new_n14043_), .A2(new_n239_), .B(new_n14032_), .ZN(new_n14044_));
  OAI21_X1   g13852(.A1(new_n14044_), .A2(new_n14042_), .B(new_n201_), .ZN(new_n14045_));
  NOR3_X1    g13853(.A1(new_n14040_), .A2(\asqrt[60] ), .A3(new_n14020_), .ZN(new_n14046_));
  OAI21_X1   g13854(.A1(new_n13967_), .A2(new_n14046_), .B(new_n14041_), .ZN(new_n14047_));
  OAI21_X1   g13855(.A1(new_n14047_), .A2(\asqrt[61] ), .B(new_n14031_), .ZN(new_n14048_));
  NAND3_X1   g13856(.A1(new_n14048_), .A2(\asqrt[62] ), .A3(new_n14029_), .ZN(new_n14049_));
  AOI21_X1   g13857(.A1(new_n13526_), .A2(new_n13532_), .B(\asqrt[12] ), .ZN(new_n14050_));
  XOR2_X1    g13858(.A1(new_n14050_), .A2(new_n13528_), .Z(new_n14051_));
  INV_X1     g13859(.I(new_n14051_), .ZN(new_n14052_));
  AOI22_X1   g13860(.A1(new_n14049_), .A2(new_n14045_), .B1(new_n14034_), .B2(new_n14052_), .ZN(new_n14053_));
  NOR2_X1    g13861(.A1(new_n13545_), .A2(new_n13456_), .ZN(new_n14054_));
  OAI21_X1   g13862(.A1(\asqrt[12] ), .A2(new_n14054_), .B(new_n13552_), .ZN(new_n14055_));
  INV_X1     g13863(.I(new_n14055_), .ZN(new_n14056_));
  OAI21_X1   g13864(.A1(new_n14053_), .A2(new_n13963_), .B(new_n14056_), .ZN(new_n14057_));
  OAI21_X1   g13865(.A1(new_n14034_), .A2(\asqrt[62] ), .B(new_n14051_), .ZN(new_n14058_));
  NAND2_X1   g13866(.A1(new_n14034_), .A2(\asqrt[62] ), .ZN(new_n14059_));
  NAND3_X1   g13867(.A1(new_n14058_), .A2(new_n14059_), .A3(new_n13963_), .ZN(new_n14060_));
  NAND2_X1   g13868(.A1(new_n13690_), .A2(new_n13455_), .ZN(new_n14061_));
  XOR2_X1    g13869(.A1(new_n13545_), .A2(new_n13456_), .Z(new_n14062_));
  NAND3_X1   g13870(.A1(new_n14061_), .A2(\asqrt[63] ), .A3(new_n14062_), .ZN(new_n14063_));
  INV_X1     g13871(.I(new_n13679_), .ZN(new_n14064_));
  NAND4_X1   g13872(.A1(new_n14064_), .A2(new_n13456_), .A3(new_n13552_), .A4(new_n13559_), .ZN(new_n14065_));
  NAND2_X1   g13873(.A1(new_n14063_), .A2(new_n14065_), .ZN(new_n14066_));
  INV_X1     g13874(.I(new_n14066_), .ZN(new_n14067_));
  NAND4_X1   g13875(.A1(new_n14057_), .A2(new_n193_), .A3(new_n14060_), .A4(new_n14067_), .ZN(\asqrt[11] ));
  AOI21_X1   g13876(.A1(new_n13940_), .A2(new_n13957_), .B(\asqrt[11] ), .ZN(new_n14069_));
  XOR2_X1    g13877(.A1(new_n14069_), .A2(new_n13562_), .Z(new_n14070_));
  AOI21_X1   g13878(.A1(new_n13937_), .A2(new_n13955_), .B(\asqrt[11] ), .ZN(new_n14071_));
  XOR2_X1    g13879(.A1(new_n14071_), .A2(new_n13565_), .Z(new_n14072_));
  NAND2_X1   g13880(.A1(new_n13950_), .A2(new_n1305_), .ZN(new_n14073_));
  AOI21_X1   g13881(.A1(new_n14073_), .A2(new_n13936_), .B(\asqrt[11] ), .ZN(new_n14074_));
  XOR2_X1    g13882(.A1(new_n14074_), .A2(new_n13568_), .Z(new_n14075_));
  INV_X1     g13883(.I(new_n14075_), .ZN(new_n14076_));
  AOI21_X1   g13884(.A1(new_n13948_), .A2(new_n13933_), .B(\asqrt[11] ), .ZN(new_n14077_));
  XOR2_X1    g13885(.A1(new_n14077_), .A2(new_n13570_), .Z(new_n14078_));
  INV_X1     g13886(.I(new_n14078_), .ZN(new_n14079_));
  NAND2_X1   g13887(.A1(new_n13915_), .A2(new_n1632_), .ZN(new_n14080_));
  AOI21_X1   g13888(.A1(new_n14080_), .A2(new_n13947_), .B(\asqrt[11] ), .ZN(new_n14081_));
  XOR2_X1    g13889(.A1(new_n14081_), .A2(new_n13573_), .Z(new_n14082_));
  AOI21_X1   g13890(.A1(new_n13913_), .A2(new_n13930_), .B(\asqrt[11] ), .ZN(new_n14083_));
  XOR2_X1    g13891(.A1(new_n14083_), .A2(new_n13577_), .Z(new_n14084_));
  NAND2_X1   g13892(.A1(new_n13926_), .A2(new_n1953_), .ZN(new_n14085_));
  AOI21_X1   g13893(.A1(new_n14085_), .A2(new_n13912_), .B(\asqrt[11] ), .ZN(new_n14086_));
  XOR2_X1    g13894(.A1(new_n14086_), .A2(new_n13580_), .Z(new_n14087_));
  INV_X1     g13895(.I(new_n14087_), .ZN(new_n14088_));
  AOI21_X1   g13896(.A1(new_n13924_), .A2(new_n13909_), .B(\asqrt[11] ), .ZN(new_n14089_));
  XOR2_X1    g13897(.A1(new_n14089_), .A2(new_n13582_), .Z(new_n14090_));
  INV_X1     g13898(.I(new_n14090_), .ZN(new_n14091_));
  NAND2_X1   g13899(.A1(new_n13891_), .A2(new_n2332_), .ZN(new_n14092_));
  AOI21_X1   g13900(.A1(new_n14092_), .A2(new_n13923_), .B(\asqrt[11] ), .ZN(new_n14093_));
  XOR2_X1    g13901(.A1(new_n14093_), .A2(new_n13585_), .Z(new_n14094_));
  AOI21_X1   g13902(.A1(new_n13889_), .A2(new_n13906_), .B(\asqrt[11] ), .ZN(new_n14095_));
  XOR2_X1    g13903(.A1(new_n14095_), .A2(new_n13589_), .Z(new_n14096_));
  NAND2_X1   g13904(.A1(new_n13902_), .A2(new_n2749_), .ZN(new_n14097_));
  AOI21_X1   g13905(.A1(new_n14097_), .A2(new_n13888_), .B(\asqrt[11] ), .ZN(new_n14098_));
  XOR2_X1    g13906(.A1(new_n14098_), .A2(new_n13592_), .Z(new_n14099_));
  INV_X1     g13907(.I(new_n14099_), .ZN(new_n14100_));
  AOI21_X1   g13908(.A1(new_n13900_), .A2(new_n13885_), .B(\asqrt[11] ), .ZN(new_n14101_));
  XOR2_X1    g13909(.A1(new_n14101_), .A2(new_n13594_), .Z(new_n14102_));
  INV_X1     g13910(.I(new_n14102_), .ZN(new_n14103_));
  NAND2_X1   g13911(.A1(new_n13867_), .A2(new_n3195_), .ZN(new_n14104_));
  AOI21_X1   g13912(.A1(new_n14104_), .A2(new_n13899_), .B(\asqrt[11] ), .ZN(new_n14105_));
  XOR2_X1    g13913(.A1(new_n14105_), .A2(new_n13597_), .Z(new_n14106_));
  AOI21_X1   g13914(.A1(new_n13865_), .A2(new_n13882_), .B(\asqrt[11] ), .ZN(new_n14107_));
  XOR2_X1    g13915(.A1(new_n14107_), .A2(new_n13601_), .Z(new_n14108_));
  NAND2_X1   g13916(.A1(new_n13878_), .A2(new_n3681_), .ZN(new_n14109_));
  AOI21_X1   g13917(.A1(new_n14109_), .A2(new_n13864_), .B(\asqrt[11] ), .ZN(new_n14110_));
  XOR2_X1    g13918(.A1(new_n14110_), .A2(new_n13604_), .Z(new_n14111_));
  INV_X1     g13919(.I(new_n14111_), .ZN(new_n14112_));
  AOI21_X1   g13920(.A1(new_n13876_), .A2(new_n13861_), .B(\asqrt[11] ), .ZN(new_n14113_));
  XOR2_X1    g13921(.A1(new_n14113_), .A2(new_n13606_), .Z(new_n14114_));
  INV_X1     g13922(.I(new_n14114_), .ZN(new_n14115_));
  NAND2_X1   g13923(.A1(new_n13843_), .A2(new_n4196_), .ZN(new_n14116_));
  AOI21_X1   g13924(.A1(new_n14116_), .A2(new_n13875_), .B(\asqrt[11] ), .ZN(new_n14117_));
  XOR2_X1    g13925(.A1(new_n14117_), .A2(new_n13609_), .Z(new_n14118_));
  AOI21_X1   g13926(.A1(new_n13841_), .A2(new_n13858_), .B(\asqrt[11] ), .ZN(new_n14119_));
  XOR2_X1    g13927(.A1(new_n14119_), .A2(new_n13613_), .Z(new_n14120_));
  NAND2_X1   g13928(.A1(new_n13854_), .A2(new_n4751_), .ZN(new_n14121_));
  AOI21_X1   g13929(.A1(new_n14121_), .A2(new_n13840_), .B(\asqrt[11] ), .ZN(new_n14122_));
  XOR2_X1    g13930(.A1(new_n14122_), .A2(new_n13616_), .Z(new_n14123_));
  INV_X1     g13931(.I(new_n14123_), .ZN(new_n14124_));
  AOI21_X1   g13932(.A1(new_n13852_), .A2(new_n13837_), .B(\asqrt[11] ), .ZN(new_n14125_));
  XOR2_X1    g13933(.A1(new_n14125_), .A2(new_n13618_), .Z(new_n14126_));
  INV_X1     g13934(.I(new_n14126_), .ZN(new_n14127_));
  NAND2_X1   g13935(.A1(new_n13819_), .A2(new_n5336_), .ZN(new_n14128_));
  AOI21_X1   g13936(.A1(new_n14128_), .A2(new_n13851_), .B(\asqrt[11] ), .ZN(new_n14129_));
  XOR2_X1    g13937(.A1(new_n14129_), .A2(new_n13621_), .Z(new_n14130_));
  AOI21_X1   g13938(.A1(new_n13817_), .A2(new_n13834_), .B(\asqrt[11] ), .ZN(new_n14131_));
  XOR2_X1    g13939(.A1(new_n14131_), .A2(new_n13625_), .Z(new_n14132_));
  NAND2_X1   g13940(.A1(new_n13830_), .A2(new_n5947_), .ZN(new_n14133_));
  AOI21_X1   g13941(.A1(new_n14133_), .A2(new_n13816_), .B(\asqrt[11] ), .ZN(new_n14134_));
  XOR2_X1    g13942(.A1(new_n14134_), .A2(new_n13628_), .Z(new_n14135_));
  INV_X1     g13943(.I(new_n14135_), .ZN(new_n14136_));
  AOI21_X1   g13944(.A1(new_n13828_), .A2(new_n13813_), .B(\asqrt[11] ), .ZN(new_n14137_));
  XOR2_X1    g13945(.A1(new_n14137_), .A2(new_n13630_), .Z(new_n14138_));
  INV_X1     g13946(.I(new_n14138_), .ZN(new_n14139_));
  NAND2_X1   g13947(.A1(new_n13795_), .A2(new_n6636_), .ZN(new_n14140_));
  AOI21_X1   g13948(.A1(new_n14140_), .A2(new_n13827_), .B(\asqrt[11] ), .ZN(new_n14141_));
  XOR2_X1    g13949(.A1(new_n14141_), .A2(new_n13633_), .Z(new_n14142_));
  AOI21_X1   g13950(.A1(new_n13793_), .A2(new_n13810_), .B(\asqrt[11] ), .ZN(new_n14143_));
  XOR2_X1    g13951(.A1(new_n14143_), .A2(new_n13637_), .Z(new_n14144_));
  NAND2_X1   g13952(.A1(new_n13806_), .A2(new_n7331_), .ZN(new_n14145_));
  AOI21_X1   g13953(.A1(new_n14145_), .A2(new_n13792_), .B(\asqrt[11] ), .ZN(new_n14146_));
  XOR2_X1    g13954(.A1(new_n14146_), .A2(new_n13640_), .Z(new_n14147_));
  INV_X1     g13955(.I(new_n14147_), .ZN(new_n14148_));
  AOI21_X1   g13956(.A1(new_n13804_), .A2(new_n13789_), .B(\asqrt[11] ), .ZN(new_n14149_));
  XOR2_X1    g13957(.A1(new_n14149_), .A2(new_n13642_), .Z(new_n14150_));
  INV_X1     g13958(.I(new_n14150_), .ZN(new_n14151_));
  NAND2_X1   g13959(.A1(new_n13771_), .A2(new_n8077_), .ZN(new_n14152_));
  AOI21_X1   g13960(.A1(new_n14152_), .A2(new_n13803_), .B(\asqrt[11] ), .ZN(new_n14153_));
  XOR2_X1    g13961(.A1(new_n14153_), .A2(new_n13645_), .Z(new_n14154_));
  AOI21_X1   g13962(.A1(new_n13769_), .A2(new_n13786_), .B(\asqrt[11] ), .ZN(new_n14155_));
  XOR2_X1    g13963(.A1(new_n14155_), .A2(new_n13649_), .Z(new_n14156_));
  NAND2_X1   g13964(.A1(new_n13782_), .A2(new_n8849_), .ZN(new_n14157_));
  AOI21_X1   g13965(.A1(new_n14157_), .A2(new_n13768_), .B(\asqrt[11] ), .ZN(new_n14158_));
  XOR2_X1    g13966(.A1(new_n14158_), .A2(new_n13652_), .Z(new_n14159_));
  INV_X1     g13967(.I(new_n14159_), .ZN(new_n14160_));
  AOI21_X1   g13968(.A1(new_n13780_), .A2(new_n13765_), .B(\asqrt[11] ), .ZN(new_n14161_));
  XOR2_X1    g13969(.A1(new_n14161_), .A2(new_n13654_), .Z(new_n14162_));
  INV_X1     g13970(.I(new_n14162_), .ZN(new_n14163_));
  NAND2_X1   g13971(.A1(new_n13747_), .A2(new_n9656_), .ZN(new_n14164_));
  AOI21_X1   g13972(.A1(new_n14164_), .A2(new_n13779_), .B(\asqrt[11] ), .ZN(new_n14165_));
  XOR2_X1    g13973(.A1(new_n14165_), .A2(new_n13657_), .Z(new_n14166_));
  AOI21_X1   g13974(.A1(new_n13745_), .A2(new_n13762_), .B(\asqrt[11] ), .ZN(new_n14167_));
  XOR2_X1    g13975(.A1(new_n14167_), .A2(new_n13661_), .Z(new_n14168_));
  NAND2_X1   g13976(.A1(new_n13758_), .A2(new_n10497_), .ZN(new_n14169_));
  AOI21_X1   g13977(.A1(new_n14169_), .A2(new_n13744_), .B(\asqrt[11] ), .ZN(new_n14170_));
  XOR2_X1    g13978(.A1(new_n14170_), .A2(new_n13664_), .Z(new_n14171_));
  INV_X1     g13979(.I(new_n14171_), .ZN(new_n14172_));
  AOI21_X1   g13980(.A1(new_n13756_), .A2(new_n13741_), .B(\asqrt[11] ), .ZN(new_n14173_));
  XOR2_X1    g13981(.A1(new_n14173_), .A2(new_n13666_), .Z(new_n14174_));
  INV_X1     g13982(.I(new_n14174_), .ZN(new_n14175_));
  NAND2_X1   g13983(.A1(new_n13719_), .A2(new_n11373_), .ZN(new_n14176_));
  AOI21_X1   g13984(.A1(new_n14176_), .A2(new_n13755_), .B(\asqrt[11] ), .ZN(new_n14177_));
  XOR2_X1    g13985(.A1(new_n14177_), .A2(new_n13669_), .Z(new_n14178_));
  AOI21_X1   g13986(.A1(new_n13717_), .A2(new_n13738_), .B(\asqrt[11] ), .ZN(new_n14179_));
  XOR2_X1    g13987(.A1(new_n14179_), .A2(new_n13672_), .Z(new_n14180_));
  NAND2_X1   g13988(.A1(new_n13734_), .A2(new_n12283_), .ZN(new_n14181_));
  AOI21_X1   g13989(.A1(new_n14181_), .A2(new_n13716_), .B(\asqrt[11] ), .ZN(new_n14182_));
  XOR2_X1    g13990(.A1(new_n14182_), .A2(new_n13678_), .Z(new_n14183_));
  INV_X1     g13991(.I(new_n14183_), .ZN(new_n14184_));
  AOI21_X1   g13992(.A1(new_n13732_), .A2(new_n13713_), .B(\asqrt[11] ), .ZN(new_n14185_));
  XOR2_X1    g13993(.A1(new_n14185_), .A2(new_n13723_), .Z(new_n14186_));
  INV_X1     g13994(.I(new_n14186_), .ZN(new_n14187_));
  NAND2_X1   g13995(.A1(\asqrt[12] ), .A2(new_n13701_), .ZN(new_n14188_));
  NOR2_X1    g13996(.A1(new_n13708_), .A2(\a[24] ), .ZN(new_n14189_));
  AOI22_X1   g13997(.A1(new_n14188_), .A2(new_n13708_), .B1(\asqrt[12] ), .B2(new_n14189_), .ZN(new_n14190_));
  OAI21_X1   g13998(.A1(new_n13690_), .A2(new_n13701_), .B(new_n13727_), .ZN(new_n14191_));
  AOI21_X1   g13999(.A1(new_n13726_), .A2(new_n14191_), .B(\asqrt[11] ), .ZN(new_n14192_));
  XOR2_X1    g14000(.A1(new_n14192_), .A2(new_n14190_), .Z(new_n14193_));
  NOR2_X1    g14001(.A1(new_n14044_), .A2(new_n14042_), .ZN(new_n14194_));
  AOI21_X1   g14002(.A1(new_n14048_), .A2(new_n14029_), .B(\asqrt[62] ), .ZN(new_n14195_));
  NOR3_X1    g14003(.A1(new_n14044_), .A2(new_n201_), .A3(new_n14042_), .ZN(new_n14196_));
  OAI22_X1   g14004(.A1(new_n14195_), .A2(new_n14196_), .B1(new_n14194_), .B2(new_n14051_), .ZN(new_n14197_));
  AOI21_X1   g14005(.A1(new_n14197_), .A2(new_n13962_), .B(new_n14055_), .ZN(new_n14198_));
  AOI21_X1   g14006(.A1(new_n14194_), .A2(new_n201_), .B(new_n14052_), .ZN(new_n14199_));
  NOR2_X1    g14007(.A1(new_n14194_), .A2(new_n201_), .ZN(new_n14200_));
  NOR3_X1    g14008(.A1(new_n14199_), .A2(new_n14200_), .A3(new_n13962_), .ZN(new_n14201_));
  NAND3_X1   g14009(.A1(new_n14063_), .A2(\asqrt[12] ), .A3(new_n14065_), .ZN(new_n14202_));
  NOR4_X1    g14010(.A1(new_n14198_), .A2(\asqrt[63] ), .A3(new_n14201_), .A4(new_n14202_), .ZN(new_n14203_));
  INV_X1     g14011(.I(new_n14203_), .ZN(new_n14204_));
  NAND2_X1   g14012(.A1(\asqrt[11] ), .A2(new_n13698_), .ZN(new_n14205_));
  AOI21_X1   g14013(.A1(new_n14205_), .A2(new_n14204_), .B(\a[24] ), .ZN(new_n14206_));
  NOR4_X1    g14014(.A1(new_n14198_), .A2(\asqrt[63] ), .A3(new_n14201_), .A4(new_n14066_), .ZN(new_n14207_));
  NOR2_X1    g14015(.A1(new_n14207_), .A2(new_n13699_), .ZN(new_n14208_));
  NOR3_X1    g14016(.A1(new_n14208_), .A2(new_n13701_), .A3(new_n14203_), .ZN(new_n14209_));
  NOR2_X1    g14017(.A1(new_n14209_), .A2(new_n14206_), .ZN(new_n14210_));
  INV_X1     g14018(.I(\a[22] ), .ZN(new_n14211_));
  NOR2_X1    g14019(.A1(\a[20] ), .A2(\a[21] ), .ZN(new_n14212_));
  NOR3_X1    g14020(.A1(new_n14207_), .A2(new_n14211_), .A3(new_n14212_), .ZN(new_n14213_));
  INV_X1     g14021(.I(new_n14212_), .ZN(new_n14214_));
  AOI21_X1   g14022(.A1(new_n14207_), .A2(\a[22] ), .B(new_n14214_), .ZN(new_n14215_));
  OAI21_X1   g14023(.A1(new_n14213_), .A2(new_n14215_), .B(\asqrt[12] ), .ZN(new_n14216_));
  NAND2_X1   g14024(.A1(new_n14212_), .A2(new_n14211_), .ZN(new_n14217_));
  NAND3_X1   g14025(.A1(new_n13555_), .A2(new_n13557_), .A3(new_n14217_), .ZN(new_n14218_));
  NAND2_X1   g14026(.A1(new_n13693_), .A2(new_n14218_), .ZN(new_n14219_));
  NAND3_X1   g14027(.A1(\asqrt[11] ), .A2(\a[22] ), .A3(new_n14219_), .ZN(new_n14220_));
  NOR3_X1    g14028(.A1(new_n14207_), .A2(\a[22] ), .A3(\a[23] ), .ZN(new_n14221_));
  INV_X1     g14029(.I(\a[23] ), .ZN(new_n14222_));
  AOI21_X1   g14030(.A1(\asqrt[11] ), .A2(new_n14211_), .B(new_n14222_), .ZN(new_n14223_));
  NOR2_X1    g14031(.A1(new_n14221_), .A2(new_n14223_), .ZN(new_n14224_));
  NAND4_X1   g14032(.A1(new_n14216_), .A2(new_n14224_), .A3(new_n13228_), .A4(new_n14220_), .ZN(new_n14225_));
  NAND2_X1   g14033(.A1(new_n14225_), .A2(new_n14210_), .ZN(new_n14226_));
  NAND3_X1   g14034(.A1(\asqrt[11] ), .A2(\a[22] ), .A3(new_n14214_), .ZN(new_n14227_));
  OAI21_X1   g14035(.A1(\asqrt[11] ), .A2(new_n14211_), .B(new_n14212_), .ZN(new_n14228_));
  AOI21_X1   g14036(.A1(new_n14228_), .A2(new_n14227_), .B(new_n13690_), .ZN(new_n14229_));
  NAND3_X1   g14037(.A1(\asqrt[11] ), .A2(new_n14211_), .A3(new_n14222_), .ZN(new_n14230_));
  OAI21_X1   g14038(.A1(new_n14207_), .A2(\a[22] ), .B(\a[23] ), .ZN(new_n14231_));
  NAND3_X1   g14039(.A1(new_n14220_), .A2(new_n14231_), .A3(new_n14230_), .ZN(new_n14232_));
  OAI21_X1   g14040(.A1(new_n14232_), .A2(new_n14229_), .B(\asqrt[13] ), .ZN(new_n14233_));
  NAND3_X1   g14041(.A1(new_n14226_), .A2(new_n12733_), .A3(new_n14233_), .ZN(new_n14234_));
  AOI21_X1   g14042(.A1(new_n14226_), .A2(new_n14233_), .B(new_n12733_), .ZN(new_n14235_));
  AOI21_X1   g14043(.A1(new_n14193_), .A2(new_n14234_), .B(new_n14235_), .ZN(new_n14236_));
  AOI21_X1   g14044(.A1(new_n14236_), .A2(new_n12283_), .B(new_n14187_), .ZN(new_n14237_));
  OR2_X2     g14045(.A1(new_n14209_), .A2(new_n14206_), .Z(new_n14238_));
  NOR3_X1    g14046(.A1(new_n14232_), .A2(new_n14229_), .A3(\asqrt[13] ), .ZN(new_n14239_));
  OAI21_X1   g14047(.A1(new_n14238_), .A2(new_n14239_), .B(new_n14233_), .ZN(new_n14240_));
  OAI21_X1   g14048(.A1(new_n14240_), .A2(\asqrt[14] ), .B(new_n14193_), .ZN(new_n14241_));
  NAND2_X1   g14049(.A1(new_n14240_), .A2(\asqrt[14] ), .ZN(new_n14242_));
  AOI21_X1   g14050(.A1(new_n14241_), .A2(new_n14242_), .B(new_n12283_), .ZN(new_n14243_));
  NOR3_X1    g14051(.A1(new_n14237_), .A2(\asqrt[16] ), .A3(new_n14243_), .ZN(new_n14244_));
  OAI21_X1   g14052(.A1(new_n14237_), .A2(new_n14243_), .B(\asqrt[16] ), .ZN(new_n14245_));
  OAI21_X1   g14053(.A1(new_n14184_), .A2(new_n14244_), .B(new_n14245_), .ZN(new_n14246_));
  OAI21_X1   g14054(.A1(new_n14246_), .A2(\asqrt[17] ), .B(new_n14180_), .ZN(new_n14247_));
  NAND3_X1   g14055(.A1(new_n14241_), .A2(new_n14242_), .A3(new_n12283_), .ZN(new_n14248_));
  AOI21_X1   g14056(.A1(new_n14186_), .A2(new_n14248_), .B(new_n14243_), .ZN(new_n14249_));
  AOI21_X1   g14057(.A1(new_n14249_), .A2(new_n11802_), .B(new_n14184_), .ZN(new_n14250_));
  NAND2_X1   g14058(.A1(new_n14248_), .A2(new_n14186_), .ZN(new_n14251_));
  INV_X1     g14059(.I(new_n14243_), .ZN(new_n14252_));
  AOI21_X1   g14060(.A1(new_n14251_), .A2(new_n14252_), .B(new_n11802_), .ZN(new_n14253_));
  OAI21_X1   g14061(.A1(new_n14250_), .A2(new_n14253_), .B(\asqrt[17] ), .ZN(new_n14254_));
  NAND3_X1   g14062(.A1(new_n14247_), .A2(new_n10914_), .A3(new_n14254_), .ZN(new_n14255_));
  AOI21_X1   g14063(.A1(new_n14247_), .A2(new_n14254_), .B(new_n10914_), .ZN(new_n14256_));
  AOI21_X1   g14064(.A1(new_n14178_), .A2(new_n14255_), .B(new_n14256_), .ZN(new_n14257_));
  AOI21_X1   g14065(.A1(new_n14257_), .A2(new_n10497_), .B(new_n14175_), .ZN(new_n14258_));
  INV_X1     g14066(.I(new_n14180_), .ZN(new_n14259_));
  NOR3_X1    g14067(.A1(new_n14250_), .A2(\asqrt[17] ), .A3(new_n14253_), .ZN(new_n14260_));
  OAI21_X1   g14068(.A1(new_n14259_), .A2(new_n14260_), .B(new_n14254_), .ZN(new_n14261_));
  OAI21_X1   g14069(.A1(new_n14261_), .A2(\asqrt[18] ), .B(new_n14178_), .ZN(new_n14262_));
  NAND2_X1   g14070(.A1(new_n14261_), .A2(\asqrt[18] ), .ZN(new_n14263_));
  AOI21_X1   g14071(.A1(new_n14262_), .A2(new_n14263_), .B(new_n10497_), .ZN(new_n14264_));
  NOR3_X1    g14072(.A1(new_n14258_), .A2(\asqrt[20] ), .A3(new_n14264_), .ZN(new_n14265_));
  OAI21_X1   g14073(.A1(new_n14258_), .A2(new_n14264_), .B(\asqrt[20] ), .ZN(new_n14266_));
  OAI21_X1   g14074(.A1(new_n14172_), .A2(new_n14265_), .B(new_n14266_), .ZN(new_n14267_));
  OAI21_X1   g14075(.A1(new_n14267_), .A2(\asqrt[21] ), .B(new_n14168_), .ZN(new_n14268_));
  NAND3_X1   g14076(.A1(new_n14262_), .A2(new_n14263_), .A3(new_n10497_), .ZN(new_n14269_));
  AOI21_X1   g14077(.A1(new_n14174_), .A2(new_n14269_), .B(new_n14264_), .ZN(new_n14270_));
  AOI21_X1   g14078(.A1(new_n14270_), .A2(new_n10052_), .B(new_n14172_), .ZN(new_n14271_));
  NAND2_X1   g14079(.A1(new_n14269_), .A2(new_n14174_), .ZN(new_n14272_));
  INV_X1     g14080(.I(new_n14264_), .ZN(new_n14273_));
  AOI21_X1   g14081(.A1(new_n14272_), .A2(new_n14273_), .B(new_n10052_), .ZN(new_n14274_));
  OAI21_X1   g14082(.A1(new_n14271_), .A2(new_n14274_), .B(\asqrt[21] ), .ZN(new_n14275_));
  NAND3_X1   g14083(.A1(new_n14268_), .A2(new_n9233_), .A3(new_n14275_), .ZN(new_n14276_));
  AOI21_X1   g14084(.A1(new_n14268_), .A2(new_n14275_), .B(new_n9233_), .ZN(new_n14277_));
  AOI21_X1   g14085(.A1(new_n14166_), .A2(new_n14276_), .B(new_n14277_), .ZN(new_n14278_));
  AOI21_X1   g14086(.A1(new_n14278_), .A2(new_n8849_), .B(new_n14163_), .ZN(new_n14279_));
  INV_X1     g14087(.I(new_n14168_), .ZN(new_n14280_));
  NOR3_X1    g14088(.A1(new_n14271_), .A2(\asqrt[21] ), .A3(new_n14274_), .ZN(new_n14281_));
  OAI21_X1   g14089(.A1(new_n14280_), .A2(new_n14281_), .B(new_n14275_), .ZN(new_n14282_));
  OAI21_X1   g14090(.A1(new_n14282_), .A2(\asqrt[22] ), .B(new_n14166_), .ZN(new_n14283_));
  NAND2_X1   g14091(.A1(new_n14282_), .A2(\asqrt[22] ), .ZN(new_n14284_));
  AOI21_X1   g14092(.A1(new_n14283_), .A2(new_n14284_), .B(new_n8849_), .ZN(new_n14285_));
  NOR3_X1    g14093(.A1(new_n14279_), .A2(\asqrt[24] ), .A3(new_n14285_), .ZN(new_n14286_));
  OAI21_X1   g14094(.A1(new_n14279_), .A2(new_n14285_), .B(\asqrt[24] ), .ZN(new_n14287_));
  OAI21_X1   g14095(.A1(new_n14160_), .A2(new_n14286_), .B(new_n14287_), .ZN(new_n14288_));
  OAI21_X1   g14096(.A1(new_n14288_), .A2(\asqrt[25] ), .B(new_n14156_), .ZN(new_n14289_));
  NAND3_X1   g14097(.A1(new_n14283_), .A2(new_n14284_), .A3(new_n8849_), .ZN(new_n14290_));
  AOI21_X1   g14098(.A1(new_n14162_), .A2(new_n14290_), .B(new_n14285_), .ZN(new_n14291_));
  AOI21_X1   g14099(.A1(new_n14291_), .A2(new_n8440_), .B(new_n14160_), .ZN(new_n14292_));
  NAND2_X1   g14100(.A1(new_n14290_), .A2(new_n14162_), .ZN(new_n14293_));
  INV_X1     g14101(.I(new_n14285_), .ZN(new_n14294_));
  AOI21_X1   g14102(.A1(new_n14293_), .A2(new_n14294_), .B(new_n8440_), .ZN(new_n14295_));
  OAI21_X1   g14103(.A1(new_n14292_), .A2(new_n14295_), .B(\asqrt[25] ), .ZN(new_n14296_));
  NAND3_X1   g14104(.A1(new_n14289_), .A2(new_n7690_), .A3(new_n14296_), .ZN(new_n14297_));
  AOI21_X1   g14105(.A1(new_n14289_), .A2(new_n14296_), .B(new_n7690_), .ZN(new_n14298_));
  AOI21_X1   g14106(.A1(new_n14154_), .A2(new_n14297_), .B(new_n14298_), .ZN(new_n14299_));
  AOI21_X1   g14107(.A1(new_n14299_), .A2(new_n7331_), .B(new_n14151_), .ZN(new_n14300_));
  INV_X1     g14108(.I(new_n14156_), .ZN(new_n14301_));
  NOR3_X1    g14109(.A1(new_n14292_), .A2(\asqrt[25] ), .A3(new_n14295_), .ZN(new_n14302_));
  OAI21_X1   g14110(.A1(new_n14301_), .A2(new_n14302_), .B(new_n14296_), .ZN(new_n14303_));
  OAI21_X1   g14111(.A1(new_n14303_), .A2(\asqrt[26] ), .B(new_n14154_), .ZN(new_n14304_));
  NAND2_X1   g14112(.A1(new_n14303_), .A2(\asqrt[26] ), .ZN(new_n14305_));
  AOI21_X1   g14113(.A1(new_n14304_), .A2(new_n14305_), .B(new_n7331_), .ZN(new_n14306_));
  NOR3_X1    g14114(.A1(new_n14300_), .A2(\asqrt[28] ), .A3(new_n14306_), .ZN(new_n14307_));
  OAI21_X1   g14115(.A1(new_n14300_), .A2(new_n14306_), .B(\asqrt[28] ), .ZN(new_n14308_));
  OAI21_X1   g14116(.A1(new_n14148_), .A2(new_n14307_), .B(new_n14308_), .ZN(new_n14309_));
  OAI21_X1   g14117(.A1(new_n14309_), .A2(\asqrt[29] ), .B(new_n14144_), .ZN(new_n14310_));
  NAND3_X1   g14118(.A1(new_n14304_), .A2(new_n14305_), .A3(new_n7331_), .ZN(new_n14311_));
  AOI21_X1   g14119(.A1(new_n14150_), .A2(new_n14311_), .B(new_n14306_), .ZN(new_n14312_));
  AOI21_X1   g14120(.A1(new_n14312_), .A2(new_n6966_), .B(new_n14148_), .ZN(new_n14313_));
  NAND2_X1   g14121(.A1(new_n14311_), .A2(new_n14150_), .ZN(new_n14314_));
  INV_X1     g14122(.I(new_n14306_), .ZN(new_n14315_));
  AOI21_X1   g14123(.A1(new_n14314_), .A2(new_n14315_), .B(new_n6966_), .ZN(new_n14316_));
  OAI21_X1   g14124(.A1(new_n14313_), .A2(new_n14316_), .B(\asqrt[29] ), .ZN(new_n14317_));
  NAND3_X1   g14125(.A1(new_n14310_), .A2(new_n6275_), .A3(new_n14317_), .ZN(new_n14318_));
  AOI21_X1   g14126(.A1(new_n14310_), .A2(new_n14317_), .B(new_n6275_), .ZN(new_n14319_));
  AOI21_X1   g14127(.A1(new_n14142_), .A2(new_n14318_), .B(new_n14319_), .ZN(new_n14320_));
  AOI21_X1   g14128(.A1(new_n14320_), .A2(new_n5947_), .B(new_n14139_), .ZN(new_n14321_));
  INV_X1     g14129(.I(new_n14144_), .ZN(new_n14322_));
  NOR3_X1    g14130(.A1(new_n14313_), .A2(\asqrt[29] ), .A3(new_n14316_), .ZN(new_n14323_));
  OAI21_X1   g14131(.A1(new_n14322_), .A2(new_n14323_), .B(new_n14317_), .ZN(new_n14324_));
  OAI21_X1   g14132(.A1(new_n14324_), .A2(\asqrt[30] ), .B(new_n14142_), .ZN(new_n14325_));
  NAND2_X1   g14133(.A1(new_n14324_), .A2(\asqrt[30] ), .ZN(new_n14326_));
  AOI21_X1   g14134(.A1(new_n14325_), .A2(new_n14326_), .B(new_n5947_), .ZN(new_n14327_));
  NOR3_X1    g14135(.A1(new_n14321_), .A2(\asqrt[32] ), .A3(new_n14327_), .ZN(new_n14328_));
  OAI21_X1   g14136(.A1(new_n14321_), .A2(new_n14327_), .B(\asqrt[32] ), .ZN(new_n14329_));
  OAI21_X1   g14137(.A1(new_n14136_), .A2(new_n14328_), .B(new_n14329_), .ZN(new_n14330_));
  OAI21_X1   g14138(.A1(new_n14330_), .A2(\asqrt[33] ), .B(new_n14132_), .ZN(new_n14331_));
  NAND3_X1   g14139(.A1(new_n14325_), .A2(new_n14326_), .A3(new_n5947_), .ZN(new_n14332_));
  AOI21_X1   g14140(.A1(new_n14138_), .A2(new_n14332_), .B(new_n14327_), .ZN(new_n14333_));
  AOI21_X1   g14141(.A1(new_n14333_), .A2(new_n5643_), .B(new_n14136_), .ZN(new_n14334_));
  NAND2_X1   g14142(.A1(new_n14332_), .A2(new_n14138_), .ZN(new_n14335_));
  INV_X1     g14143(.I(new_n14327_), .ZN(new_n14336_));
  AOI21_X1   g14144(.A1(new_n14335_), .A2(new_n14336_), .B(new_n5643_), .ZN(new_n14337_));
  OAI21_X1   g14145(.A1(new_n14334_), .A2(new_n14337_), .B(\asqrt[33] ), .ZN(new_n14338_));
  NAND3_X1   g14146(.A1(new_n14331_), .A2(new_n5029_), .A3(new_n14338_), .ZN(new_n14339_));
  AOI21_X1   g14147(.A1(new_n14331_), .A2(new_n14338_), .B(new_n5029_), .ZN(new_n14340_));
  AOI21_X1   g14148(.A1(new_n14130_), .A2(new_n14339_), .B(new_n14340_), .ZN(new_n14341_));
  AOI21_X1   g14149(.A1(new_n14341_), .A2(new_n4751_), .B(new_n14127_), .ZN(new_n14342_));
  INV_X1     g14150(.I(new_n14132_), .ZN(new_n14343_));
  NOR3_X1    g14151(.A1(new_n14334_), .A2(\asqrt[33] ), .A3(new_n14337_), .ZN(new_n14344_));
  OAI21_X1   g14152(.A1(new_n14343_), .A2(new_n14344_), .B(new_n14338_), .ZN(new_n14345_));
  OAI21_X1   g14153(.A1(new_n14345_), .A2(\asqrt[34] ), .B(new_n14130_), .ZN(new_n14346_));
  NAND2_X1   g14154(.A1(new_n14345_), .A2(\asqrt[34] ), .ZN(new_n14347_));
  AOI21_X1   g14155(.A1(new_n14346_), .A2(new_n14347_), .B(new_n4751_), .ZN(new_n14348_));
  NOR3_X1    g14156(.A1(new_n14342_), .A2(\asqrt[36] ), .A3(new_n14348_), .ZN(new_n14349_));
  OAI21_X1   g14157(.A1(new_n14342_), .A2(new_n14348_), .B(\asqrt[36] ), .ZN(new_n14350_));
  OAI21_X1   g14158(.A1(new_n14124_), .A2(new_n14349_), .B(new_n14350_), .ZN(new_n14351_));
  OAI21_X1   g14159(.A1(new_n14351_), .A2(\asqrt[37] ), .B(new_n14120_), .ZN(new_n14352_));
  NAND3_X1   g14160(.A1(new_n14346_), .A2(new_n14347_), .A3(new_n4751_), .ZN(new_n14353_));
  AOI21_X1   g14161(.A1(new_n14126_), .A2(new_n14353_), .B(new_n14348_), .ZN(new_n14354_));
  AOI21_X1   g14162(.A1(new_n14354_), .A2(new_n4461_), .B(new_n14124_), .ZN(new_n14355_));
  NAND2_X1   g14163(.A1(new_n14353_), .A2(new_n14126_), .ZN(new_n14356_));
  INV_X1     g14164(.I(new_n14348_), .ZN(new_n14357_));
  AOI21_X1   g14165(.A1(new_n14356_), .A2(new_n14357_), .B(new_n4461_), .ZN(new_n14358_));
  OAI21_X1   g14166(.A1(new_n14355_), .A2(new_n14358_), .B(\asqrt[37] ), .ZN(new_n14359_));
  NAND3_X1   g14167(.A1(new_n14352_), .A2(new_n3925_), .A3(new_n14359_), .ZN(new_n14360_));
  AOI21_X1   g14168(.A1(new_n14352_), .A2(new_n14359_), .B(new_n3925_), .ZN(new_n14361_));
  AOI21_X1   g14169(.A1(new_n14118_), .A2(new_n14360_), .B(new_n14361_), .ZN(new_n14362_));
  AOI21_X1   g14170(.A1(new_n14362_), .A2(new_n3681_), .B(new_n14115_), .ZN(new_n14363_));
  INV_X1     g14171(.I(new_n14120_), .ZN(new_n14364_));
  NOR3_X1    g14172(.A1(new_n14355_), .A2(\asqrt[37] ), .A3(new_n14358_), .ZN(new_n14365_));
  OAI21_X1   g14173(.A1(new_n14364_), .A2(new_n14365_), .B(new_n14359_), .ZN(new_n14366_));
  OAI21_X1   g14174(.A1(new_n14366_), .A2(\asqrt[38] ), .B(new_n14118_), .ZN(new_n14367_));
  NAND2_X1   g14175(.A1(new_n14366_), .A2(\asqrt[38] ), .ZN(new_n14368_));
  AOI21_X1   g14176(.A1(new_n14367_), .A2(new_n14368_), .B(new_n3681_), .ZN(new_n14369_));
  NOR3_X1    g14177(.A1(new_n14363_), .A2(\asqrt[40] ), .A3(new_n14369_), .ZN(new_n14370_));
  OAI21_X1   g14178(.A1(new_n14363_), .A2(new_n14369_), .B(\asqrt[40] ), .ZN(new_n14371_));
  OAI21_X1   g14179(.A1(new_n14112_), .A2(new_n14370_), .B(new_n14371_), .ZN(new_n14372_));
  OAI21_X1   g14180(.A1(new_n14372_), .A2(\asqrt[41] ), .B(new_n14108_), .ZN(new_n14373_));
  NAND3_X1   g14181(.A1(new_n14367_), .A2(new_n14368_), .A3(new_n3681_), .ZN(new_n14374_));
  AOI21_X1   g14182(.A1(new_n14114_), .A2(new_n14374_), .B(new_n14369_), .ZN(new_n14375_));
  AOI21_X1   g14183(.A1(new_n14375_), .A2(new_n3427_), .B(new_n14112_), .ZN(new_n14376_));
  NAND2_X1   g14184(.A1(new_n14374_), .A2(new_n14114_), .ZN(new_n14377_));
  INV_X1     g14185(.I(new_n14369_), .ZN(new_n14378_));
  AOI21_X1   g14186(.A1(new_n14377_), .A2(new_n14378_), .B(new_n3427_), .ZN(new_n14379_));
  OAI21_X1   g14187(.A1(new_n14376_), .A2(new_n14379_), .B(\asqrt[41] ), .ZN(new_n14380_));
  NAND3_X1   g14188(.A1(new_n14373_), .A2(new_n2960_), .A3(new_n14380_), .ZN(new_n14381_));
  AOI21_X1   g14189(.A1(new_n14373_), .A2(new_n14380_), .B(new_n2960_), .ZN(new_n14382_));
  AOI21_X1   g14190(.A1(new_n14106_), .A2(new_n14381_), .B(new_n14382_), .ZN(new_n14383_));
  AOI21_X1   g14191(.A1(new_n14383_), .A2(new_n2749_), .B(new_n14103_), .ZN(new_n14384_));
  INV_X1     g14192(.I(new_n14108_), .ZN(new_n14385_));
  NOR3_X1    g14193(.A1(new_n14376_), .A2(\asqrt[41] ), .A3(new_n14379_), .ZN(new_n14386_));
  OAI21_X1   g14194(.A1(new_n14385_), .A2(new_n14386_), .B(new_n14380_), .ZN(new_n14387_));
  OAI21_X1   g14195(.A1(new_n14387_), .A2(\asqrt[42] ), .B(new_n14106_), .ZN(new_n14388_));
  NAND2_X1   g14196(.A1(new_n14387_), .A2(\asqrt[42] ), .ZN(new_n14389_));
  AOI21_X1   g14197(.A1(new_n14388_), .A2(new_n14389_), .B(new_n2749_), .ZN(new_n14390_));
  NOR3_X1    g14198(.A1(new_n14384_), .A2(\asqrt[44] ), .A3(new_n14390_), .ZN(new_n14391_));
  OAI21_X1   g14199(.A1(new_n14384_), .A2(new_n14390_), .B(\asqrt[44] ), .ZN(new_n14392_));
  OAI21_X1   g14200(.A1(new_n14100_), .A2(new_n14391_), .B(new_n14392_), .ZN(new_n14393_));
  OAI21_X1   g14201(.A1(new_n14393_), .A2(\asqrt[45] ), .B(new_n14096_), .ZN(new_n14394_));
  NAND3_X1   g14202(.A1(new_n14388_), .A2(new_n14389_), .A3(new_n2749_), .ZN(new_n14395_));
  AOI21_X1   g14203(.A1(new_n14102_), .A2(new_n14395_), .B(new_n14390_), .ZN(new_n14396_));
  AOI21_X1   g14204(.A1(new_n14396_), .A2(new_n2531_), .B(new_n14100_), .ZN(new_n14397_));
  NAND2_X1   g14205(.A1(new_n14395_), .A2(new_n14102_), .ZN(new_n14398_));
  INV_X1     g14206(.I(new_n14390_), .ZN(new_n14399_));
  AOI21_X1   g14207(.A1(new_n14398_), .A2(new_n14399_), .B(new_n2531_), .ZN(new_n14400_));
  OAI21_X1   g14208(.A1(new_n14397_), .A2(new_n14400_), .B(\asqrt[45] ), .ZN(new_n14401_));
  NAND3_X1   g14209(.A1(new_n14394_), .A2(new_n2134_), .A3(new_n14401_), .ZN(new_n14402_));
  AOI21_X1   g14210(.A1(new_n14394_), .A2(new_n14401_), .B(new_n2134_), .ZN(new_n14403_));
  AOI21_X1   g14211(.A1(new_n14094_), .A2(new_n14402_), .B(new_n14403_), .ZN(new_n14404_));
  AOI21_X1   g14212(.A1(new_n14404_), .A2(new_n1953_), .B(new_n14091_), .ZN(new_n14405_));
  INV_X1     g14213(.I(new_n14096_), .ZN(new_n14406_));
  NOR3_X1    g14214(.A1(new_n14397_), .A2(\asqrt[45] ), .A3(new_n14400_), .ZN(new_n14407_));
  OAI21_X1   g14215(.A1(new_n14406_), .A2(new_n14407_), .B(new_n14401_), .ZN(new_n14408_));
  OAI21_X1   g14216(.A1(new_n14408_), .A2(\asqrt[46] ), .B(new_n14094_), .ZN(new_n14409_));
  NAND2_X1   g14217(.A1(new_n14408_), .A2(\asqrt[46] ), .ZN(new_n14410_));
  AOI21_X1   g14218(.A1(new_n14409_), .A2(new_n14410_), .B(new_n1953_), .ZN(new_n14411_));
  NOR3_X1    g14219(.A1(new_n14405_), .A2(\asqrt[48] ), .A3(new_n14411_), .ZN(new_n14412_));
  OAI21_X1   g14220(.A1(new_n14405_), .A2(new_n14411_), .B(\asqrt[48] ), .ZN(new_n14413_));
  OAI21_X1   g14221(.A1(new_n14088_), .A2(new_n14412_), .B(new_n14413_), .ZN(new_n14414_));
  OAI21_X1   g14222(.A1(new_n14414_), .A2(\asqrt[49] ), .B(new_n14084_), .ZN(new_n14415_));
  NAND3_X1   g14223(.A1(new_n14409_), .A2(new_n14410_), .A3(new_n1953_), .ZN(new_n14416_));
  AOI21_X1   g14224(.A1(new_n14090_), .A2(new_n14416_), .B(new_n14411_), .ZN(new_n14417_));
  AOI21_X1   g14225(.A1(new_n14417_), .A2(new_n1778_), .B(new_n14088_), .ZN(new_n14418_));
  NAND2_X1   g14226(.A1(new_n14416_), .A2(new_n14090_), .ZN(new_n14419_));
  INV_X1     g14227(.I(new_n14411_), .ZN(new_n14420_));
  AOI21_X1   g14228(.A1(new_n14419_), .A2(new_n14420_), .B(new_n1778_), .ZN(new_n14421_));
  OAI21_X1   g14229(.A1(new_n14418_), .A2(new_n14421_), .B(\asqrt[49] ), .ZN(new_n14422_));
  NAND3_X1   g14230(.A1(new_n14415_), .A2(new_n1463_), .A3(new_n14422_), .ZN(new_n14423_));
  AOI21_X1   g14231(.A1(new_n14415_), .A2(new_n14422_), .B(new_n1463_), .ZN(new_n14424_));
  AOI21_X1   g14232(.A1(new_n14082_), .A2(new_n14423_), .B(new_n14424_), .ZN(new_n14425_));
  AOI21_X1   g14233(.A1(new_n14425_), .A2(new_n1305_), .B(new_n14079_), .ZN(new_n14426_));
  INV_X1     g14234(.I(new_n14084_), .ZN(new_n14427_));
  NOR3_X1    g14235(.A1(new_n14418_), .A2(\asqrt[49] ), .A3(new_n14421_), .ZN(new_n14428_));
  OAI21_X1   g14236(.A1(new_n14427_), .A2(new_n14428_), .B(new_n14422_), .ZN(new_n14429_));
  OAI21_X1   g14237(.A1(new_n14429_), .A2(\asqrt[50] ), .B(new_n14082_), .ZN(new_n14430_));
  NAND2_X1   g14238(.A1(new_n14429_), .A2(\asqrt[50] ), .ZN(new_n14431_));
  AOI21_X1   g14239(.A1(new_n14430_), .A2(new_n14431_), .B(new_n1305_), .ZN(new_n14432_));
  NOR3_X1    g14240(.A1(new_n14426_), .A2(\asqrt[52] ), .A3(new_n14432_), .ZN(new_n14433_));
  OAI21_X1   g14241(.A1(new_n14426_), .A2(new_n14432_), .B(\asqrt[52] ), .ZN(new_n14434_));
  OAI21_X1   g14242(.A1(new_n14076_), .A2(new_n14433_), .B(new_n14434_), .ZN(new_n14435_));
  OAI21_X1   g14243(.A1(new_n14435_), .A2(\asqrt[53] ), .B(new_n14072_), .ZN(new_n14436_));
  NAND3_X1   g14244(.A1(new_n14430_), .A2(new_n14431_), .A3(new_n1305_), .ZN(new_n14437_));
  AOI21_X1   g14245(.A1(new_n14078_), .A2(new_n14437_), .B(new_n14432_), .ZN(new_n14438_));
  AOI21_X1   g14246(.A1(new_n14438_), .A2(new_n1150_), .B(new_n14076_), .ZN(new_n14439_));
  NAND2_X1   g14247(.A1(new_n14437_), .A2(new_n14078_), .ZN(new_n14440_));
  INV_X1     g14248(.I(new_n14432_), .ZN(new_n14441_));
  AOI21_X1   g14249(.A1(new_n14440_), .A2(new_n14441_), .B(new_n1150_), .ZN(new_n14442_));
  OAI21_X1   g14250(.A1(new_n14439_), .A2(new_n14442_), .B(\asqrt[53] ), .ZN(new_n14443_));
  NAND3_X1   g14251(.A1(new_n14436_), .A2(new_n860_), .A3(new_n14443_), .ZN(new_n14444_));
  INV_X1     g14252(.I(new_n14072_), .ZN(new_n14445_));
  NOR3_X1    g14253(.A1(new_n14439_), .A2(\asqrt[53] ), .A3(new_n14442_), .ZN(new_n14446_));
  OAI21_X1   g14254(.A1(new_n14445_), .A2(new_n14446_), .B(new_n14443_), .ZN(new_n14447_));
  NAND2_X1   g14255(.A1(new_n14447_), .A2(\asqrt[54] ), .ZN(new_n14448_));
  NOR2_X1    g14256(.A1(new_n14034_), .A2(\asqrt[62] ), .ZN(new_n14449_));
  NOR2_X1    g14257(.A1(new_n14449_), .A2(new_n14200_), .ZN(new_n14450_));
  XOR2_X1    g14258(.A1(new_n14050_), .A2(new_n13528_), .Z(new_n14451_));
  OAI21_X1   g14259(.A1(\asqrt[11] ), .A2(new_n14450_), .B(new_n14451_), .ZN(new_n14452_));
  INV_X1     g14260(.I(new_n14452_), .ZN(new_n14453_));
  AOI21_X1   g14261(.A1(new_n14019_), .A2(new_n14027_), .B(\asqrt[11] ), .ZN(new_n14454_));
  XOR2_X1    g14262(.A1(new_n14454_), .A2(new_n13970_), .Z(new_n14455_));
  INV_X1     g14263(.I(new_n14455_), .ZN(new_n14456_));
  AOI21_X1   g14264(.A1(new_n14010_), .A2(new_n14018_), .B(\asqrt[11] ), .ZN(new_n14457_));
  XOR2_X1    g14265(.A1(new_n14457_), .A2(new_n13972_), .Z(new_n14458_));
  INV_X1     g14266(.I(new_n14458_), .ZN(new_n14459_));
  NAND2_X1   g14267(.A1(new_n14014_), .A2(new_n531_), .ZN(new_n14460_));
  AOI21_X1   g14268(.A1(new_n14460_), .A2(new_n14009_), .B(\asqrt[11] ), .ZN(new_n14461_));
  XOR2_X1    g14269(.A1(new_n14461_), .A2(new_n13974_), .Z(new_n14462_));
  AOI21_X1   g14270(.A1(new_n14013_), .A2(new_n13999_), .B(\asqrt[11] ), .ZN(new_n14463_));
  XOR2_X1    g14271(.A1(new_n14463_), .A2(new_n13978_), .Z(new_n14464_));
  NAND2_X1   g14272(.A1(new_n13989_), .A2(new_n744_), .ZN(new_n14465_));
  AOI21_X1   g14273(.A1(new_n14465_), .A2(new_n14007_), .B(\asqrt[11] ), .ZN(new_n14466_));
  XOR2_X1    g14274(.A1(new_n14466_), .A2(new_n13982_), .Z(new_n14467_));
  INV_X1     g14275(.I(new_n14467_), .ZN(new_n14468_));
  AOI21_X1   g14276(.A1(new_n13987_), .A2(new_n13996_), .B(\asqrt[11] ), .ZN(new_n14469_));
  XOR2_X1    g14277(.A1(new_n14469_), .A2(new_n13985_), .Z(new_n14470_));
  INV_X1     g14278(.I(new_n14470_), .ZN(new_n14471_));
  AOI21_X1   g14279(.A1(new_n14436_), .A2(new_n14443_), .B(new_n860_), .ZN(new_n14472_));
  AOI21_X1   g14280(.A1(new_n14070_), .A2(new_n14444_), .B(new_n14472_), .ZN(new_n14473_));
  AOI21_X1   g14281(.A1(new_n14473_), .A2(new_n744_), .B(new_n14471_), .ZN(new_n14474_));
  OAI21_X1   g14282(.A1(new_n14447_), .A2(\asqrt[54] ), .B(new_n14070_), .ZN(new_n14475_));
  AOI21_X1   g14283(.A1(new_n14475_), .A2(new_n14448_), .B(new_n744_), .ZN(new_n14476_));
  NOR3_X1    g14284(.A1(new_n14474_), .A2(\asqrt[56] ), .A3(new_n14476_), .ZN(new_n14477_));
  OAI21_X1   g14285(.A1(new_n14474_), .A2(new_n14476_), .B(\asqrt[56] ), .ZN(new_n14478_));
  OAI21_X1   g14286(.A1(new_n14468_), .A2(new_n14477_), .B(new_n14478_), .ZN(new_n14479_));
  OAI21_X1   g14287(.A1(new_n14479_), .A2(\asqrt[57] ), .B(new_n14464_), .ZN(new_n14480_));
  NAND3_X1   g14288(.A1(new_n14475_), .A2(new_n14448_), .A3(new_n744_), .ZN(new_n14481_));
  AOI21_X1   g14289(.A1(new_n14470_), .A2(new_n14481_), .B(new_n14476_), .ZN(new_n14482_));
  AOI21_X1   g14290(.A1(new_n14482_), .A2(new_n634_), .B(new_n14468_), .ZN(new_n14483_));
  NAND2_X1   g14291(.A1(new_n14481_), .A2(new_n14470_), .ZN(new_n14484_));
  INV_X1     g14292(.I(new_n14476_), .ZN(new_n14485_));
  AOI21_X1   g14293(.A1(new_n14484_), .A2(new_n14485_), .B(new_n634_), .ZN(new_n14486_));
  OAI21_X1   g14294(.A1(new_n14483_), .A2(new_n14486_), .B(\asqrt[57] ), .ZN(new_n14487_));
  NAND3_X1   g14295(.A1(new_n14480_), .A2(new_n423_), .A3(new_n14487_), .ZN(new_n14488_));
  AOI21_X1   g14296(.A1(new_n14480_), .A2(new_n14487_), .B(new_n423_), .ZN(new_n14489_));
  AOI21_X1   g14297(.A1(new_n14462_), .A2(new_n14488_), .B(new_n14489_), .ZN(new_n14490_));
  AOI21_X1   g14298(.A1(new_n14490_), .A2(new_n337_), .B(new_n14459_), .ZN(new_n14491_));
  NOR2_X1    g14299(.A1(new_n14490_), .A2(new_n337_), .ZN(new_n14492_));
  NOR3_X1    g14300(.A1(new_n14491_), .A2(new_n14492_), .A3(\asqrt[60] ), .ZN(new_n14493_));
  OAI21_X1   g14301(.A1(new_n14491_), .A2(new_n14492_), .B(\asqrt[60] ), .ZN(new_n14494_));
  OAI21_X1   g14302(.A1(new_n14456_), .A2(new_n14493_), .B(new_n14494_), .ZN(new_n14495_));
  NAND2_X1   g14303(.A1(new_n14495_), .A2(\asqrt[61] ), .ZN(new_n14496_));
  AOI21_X1   g14304(.A1(new_n14035_), .A2(new_n14041_), .B(\asqrt[11] ), .ZN(new_n14497_));
  XOR2_X1    g14305(.A1(new_n14497_), .A2(new_n13966_), .Z(new_n14498_));
  OAI21_X1   g14306(.A1(new_n14495_), .A2(\asqrt[61] ), .B(new_n14498_), .ZN(new_n14499_));
  NAND2_X1   g14307(.A1(new_n14499_), .A2(new_n14496_), .ZN(new_n14500_));
  INV_X1     g14308(.I(new_n14464_), .ZN(new_n14501_));
  NOR3_X1    g14309(.A1(new_n14483_), .A2(\asqrt[57] ), .A3(new_n14486_), .ZN(new_n14502_));
  OAI21_X1   g14310(.A1(new_n14501_), .A2(new_n14502_), .B(new_n14487_), .ZN(new_n14503_));
  OAI21_X1   g14311(.A1(new_n14503_), .A2(\asqrt[58] ), .B(new_n14462_), .ZN(new_n14504_));
  NOR2_X1    g14312(.A1(new_n14502_), .A2(new_n14501_), .ZN(new_n14505_));
  INV_X1     g14313(.I(new_n14487_), .ZN(new_n14506_));
  OAI21_X1   g14314(.A1(new_n14505_), .A2(new_n14506_), .B(\asqrt[58] ), .ZN(new_n14507_));
  NAND3_X1   g14315(.A1(new_n14504_), .A2(new_n337_), .A3(new_n14507_), .ZN(new_n14508_));
  NAND2_X1   g14316(.A1(new_n14508_), .A2(new_n14458_), .ZN(new_n14509_));
  INV_X1     g14317(.I(new_n14462_), .ZN(new_n14510_));
  NOR2_X1    g14318(.A1(new_n14505_), .A2(new_n14506_), .ZN(new_n14511_));
  AOI21_X1   g14319(.A1(new_n14511_), .A2(new_n423_), .B(new_n14510_), .ZN(new_n14512_));
  OAI21_X1   g14320(.A1(new_n14512_), .A2(new_n14489_), .B(\asqrt[59] ), .ZN(new_n14513_));
  NAND3_X1   g14321(.A1(new_n14509_), .A2(new_n266_), .A3(new_n14513_), .ZN(new_n14514_));
  NAND2_X1   g14322(.A1(new_n14514_), .A2(new_n14455_), .ZN(new_n14515_));
  AOI21_X1   g14323(.A1(new_n14515_), .A2(new_n14494_), .B(new_n239_), .ZN(new_n14516_));
  AOI21_X1   g14324(.A1(new_n14509_), .A2(new_n14513_), .B(new_n266_), .ZN(new_n14517_));
  AOI21_X1   g14325(.A1(new_n14455_), .A2(new_n14514_), .B(new_n14517_), .ZN(new_n14518_));
  INV_X1     g14326(.I(new_n14498_), .ZN(new_n14519_));
  AOI21_X1   g14327(.A1(new_n14518_), .A2(new_n239_), .B(new_n14519_), .ZN(new_n14520_));
  OAI21_X1   g14328(.A1(new_n14520_), .A2(new_n14516_), .B(new_n201_), .ZN(new_n14521_));
  NAND3_X1   g14329(.A1(new_n14499_), .A2(new_n14496_), .A3(\asqrt[62] ), .ZN(new_n14522_));
  NOR2_X1    g14330(.A1(new_n14033_), .A2(new_n14042_), .ZN(new_n14523_));
  NOR2_X1    g14331(.A1(\asqrt[11] ), .A2(new_n14523_), .ZN(new_n14524_));
  XOR2_X1    g14332(.A1(new_n14524_), .A2(new_n14031_), .Z(new_n14525_));
  INV_X1     g14333(.I(new_n14525_), .ZN(new_n14526_));
  AOI22_X1   g14334(.A1(new_n14522_), .A2(new_n14521_), .B1(new_n14500_), .B2(new_n14526_), .ZN(new_n14527_));
  NOR2_X1    g14335(.A1(new_n14053_), .A2(new_n13963_), .ZN(new_n14528_));
  OAI21_X1   g14336(.A1(\asqrt[11] ), .A2(new_n14528_), .B(new_n14060_), .ZN(new_n14529_));
  INV_X1     g14337(.I(new_n14529_), .ZN(new_n14530_));
  OAI21_X1   g14338(.A1(new_n14527_), .A2(new_n14453_), .B(new_n14530_), .ZN(new_n14531_));
  OAI21_X1   g14339(.A1(new_n14500_), .A2(\asqrt[62] ), .B(new_n14525_), .ZN(new_n14532_));
  NAND2_X1   g14340(.A1(new_n14500_), .A2(\asqrt[62] ), .ZN(new_n14533_));
  NAND3_X1   g14341(.A1(new_n14532_), .A2(new_n14533_), .A3(new_n14453_), .ZN(new_n14534_));
  NAND2_X1   g14342(.A1(new_n14053_), .A2(new_n13962_), .ZN(new_n14535_));
  NAND2_X1   g14343(.A1(new_n14197_), .A2(new_n13963_), .ZN(new_n14536_));
  AOI21_X1   g14344(.A1(new_n14535_), .A2(new_n14536_), .B(new_n193_), .ZN(new_n14537_));
  OAI21_X1   g14345(.A1(\asqrt[11] ), .A2(new_n13963_), .B(new_n14537_), .ZN(new_n14538_));
  NOR2_X1    g14346(.A1(new_n14066_), .A2(new_n13962_), .ZN(new_n14539_));
  NAND4_X1   g14347(.A1(new_n14057_), .A2(new_n193_), .A3(new_n14060_), .A4(new_n14539_), .ZN(new_n14540_));
  NAND2_X1   g14348(.A1(new_n14538_), .A2(new_n14540_), .ZN(new_n14541_));
  INV_X1     g14349(.I(new_n14541_), .ZN(new_n14542_));
  NAND4_X1   g14350(.A1(new_n14531_), .A2(new_n193_), .A3(new_n14534_), .A4(new_n14542_), .ZN(\asqrt[10] ));
  AOI21_X1   g14351(.A1(new_n14444_), .A2(new_n14448_), .B(\asqrt[10] ), .ZN(new_n14544_));
  XOR2_X1    g14352(.A1(new_n14544_), .A2(new_n14070_), .Z(new_n14545_));
  XOR2_X1    g14353(.A1(new_n14435_), .A2(\asqrt[53] ), .Z(new_n14546_));
  NOR2_X1    g14354(.A1(\asqrt[10] ), .A2(new_n14546_), .ZN(new_n14547_));
  XOR2_X1    g14355(.A1(new_n14547_), .A2(new_n14072_), .Z(new_n14548_));
  NOR2_X1    g14356(.A1(new_n14433_), .A2(new_n14442_), .ZN(new_n14549_));
  NOR2_X1    g14357(.A1(\asqrt[10] ), .A2(new_n14549_), .ZN(new_n14550_));
  XOR2_X1    g14358(.A1(new_n14550_), .A2(new_n14075_), .Z(new_n14551_));
  AOI21_X1   g14359(.A1(new_n14437_), .A2(new_n14441_), .B(\asqrt[10] ), .ZN(new_n14552_));
  XOR2_X1    g14360(.A1(new_n14552_), .A2(new_n14078_), .Z(new_n14553_));
  INV_X1     g14361(.I(new_n14553_), .ZN(new_n14554_));
  AOI21_X1   g14362(.A1(new_n14423_), .A2(new_n14431_), .B(\asqrt[10] ), .ZN(new_n14555_));
  XOR2_X1    g14363(.A1(new_n14555_), .A2(new_n14082_), .Z(new_n14556_));
  INV_X1     g14364(.I(new_n14556_), .ZN(new_n14557_));
  XOR2_X1    g14365(.A1(new_n14414_), .A2(\asqrt[49] ), .Z(new_n14558_));
  NOR2_X1    g14366(.A1(\asqrt[10] ), .A2(new_n14558_), .ZN(new_n14559_));
  XOR2_X1    g14367(.A1(new_n14559_), .A2(new_n14084_), .Z(new_n14560_));
  NOR2_X1    g14368(.A1(new_n14412_), .A2(new_n14421_), .ZN(new_n14561_));
  NOR2_X1    g14369(.A1(\asqrt[10] ), .A2(new_n14561_), .ZN(new_n14562_));
  XOR2_X1    g14370(.A1(new_n14562_), .A2(new_n14087_), .Z(new_n14563_));
  AOI21_X1   g14371(.A1(new_n14416_), .A2(new_n14420_), .B(\asqrt[10] ), .ZN(new_n14564_));
  XOR2_X1    g14372(.A1(new_n14564_), .A2(new_n14090_), .Z(new_n14565_));
  INV_X1     g14373(.I(new_n14565_), .ZN(new_n14566_));
  AOI21_X1   g14374(.A1(new_n14402_), .A2(new_n14410_), .B(\asqrt[10] ), .ZN(new_n14567_));
  XOR2_X1    g14375(.A1(new_n14567_), .A2(new_n14094_), .Z(new_n14568_));
  INV_X1     g14376(.I(new_n14568_), .ZN(new_n14569_));
  XOR2_X1    g14377(.A1(new_n14393_), .A2(\asqrt[45] ), .Z(new_n14570_));
  NOR2_X1    g14378(.A1(\asqrt[10] ), .A2(new_n14570_), .ZN(new_n14571_));
  XOR2_X1    g14379(.A1(new_n14571_), .A2(new_n14096_), .Z(new_n14572_));
  NOR2_X1    g14380(.A1(new_n14391_), .A2(new_n14400_), .ZN(new_n14573_));
  NOR2_X1    g14381(.A1(\asqrt[10] ), .A2(new_n14573_), .ZN(new_n14574_));
  XOR2_X1    g14382(.A1(new_n14574_), .A2(new_n14099_), .Z(new_n14575_));
  AOI21_X1   g14383(.A1(new_n14395_), .A2(new_n14399_), .B(\asqrt[10] ), .ZN(new_n14576_));
  XOR2_X1    g14384(.A1(new_n14576_), .A2(new_n14102_), .Z(new_n14577_));
  INV_X1     g14385(.I(new_n14577_), .ZN(new_n14578_));
  AOI21_X1   g14386(.A1(new_n14381_), .A2(new_n14389_), .B(\asqrt[10] ), .ZN(new_n14579_));
  XOR2_X1    g14387(.A1(new_n14579_), .A2(new_n14106_), .Z(new_n14580_));
  INV_X1     g14388(.I(new_n14580_), .ZN(new_n14581_));
  XOR2_X1    g14389(.A1(new_n14372_), .A2(\asqrt[41] ), .Z(new_n14582_));
  NOR2_X1    g14390(.A1(\asqrt[10] ), .A2(new_n14582_), .ZN(new_n14583_));
  XOR2_X1    g14391(.A1(new_n14583_), .A2(new_n14108_), .Z(new_n14584_));
  NOR2_X1    g14392(.A1(new_n14370_), .A2(new_n14379_), .ZN(new_n14585_));
  NOR2_X1    g14393(.A1(\asqrt[10] ), .A2(new_n14585_), .ZN(new_n14586_));
  XOR2_X1    g14394(.A1(new_n14586_), .A2(new_n14111_), .Z(new_n14587_));
  AOI21_X1   g14395(.A1(new_n14374_), .A2(new_n14378_), .B(\asqrt[10] ), .ZN(new_n14588_));
  XOR2_X1    g14396(.A1(new_n14588_), .A2(new_n14114_), .Z(new_n14589_));
  INV_X1     g14397(.I(new_n14589_), .ZN(new_n14590_));
  AOI21_X1   g14398(.A1(new_n14360_), .A2(new_n14368_), .B(\asqrt[10] ), .ZN(new_n14591_));
  XOR2_X1    g14399(.A1(new_n14591_), .A2(new_n14118_), .Z(new_n14592_));
  INV_X1     g14400(.I(new_n14592_), .ZN(new_n14593_));
  XOR2_X1    g14401(.A1(new_n14351_), .A2(\asqrt[37] ), .Z(new_n14594_));
  NOR2_X1    g14402(.A1(\asqrt[10] ), .A2(new_n14594_), .ZN(new_n14595_));
  XOR2_X1    g14403(.A1(new_n14595_), .A2(new_n14120_), .Z(new_n14596_));
  NOR2_X1    g14404(.A1(new_n14349_), .A2(new_n14358_), .ZN(new_n14597_));
  NOR2_X1    g14405(.A1(\asqrt[10] ), .A2(new_n14597_), .ZN(new_n14598_));
  XOR2_X1    g14406(.A1(new_n14598_), .A2(new_n14123_), .Z(new_n14599_));
  AOI21_X1   g14407(.A1(new_n14353_), .A2(new_n14357_), .B(\asqrt[10] ), .ZN(new_n14600_));
  XOR2_X1    g14408(.A1(new_n14600_), .A2(new_n14126_), .Z(new_n14601_));
  INV_X1     g14409(.I(new_n14601_), .ZN(new_n14602_));
  AOI21_X1   g14410(.A1(new_n14339_), .A2(new_n14347_), .B(\asqrt[10] ), .ZN(new_n14603_));
  XOR2_X1    g14411(.A1(new_n14603_), .A2(new_n14130_), .Z(new_n14604_));
  INV_X1     g14412(.I(new_n14604_), .ZN(new_n14605_));
  XOR2_X1    g14413(.A1(new_n14330_), .A2(\asqrt[33] ), .Z(new_n14606_));
  NOR2_X1    g14414(.A1(\asqrt[10] ), .A2(new_n14606_), .ZN(new_n14607_));
  XOR2_X1    g14415(.A1(new_n14607_), .A2(new_n14132_), .Z(new_n14608_));
  NOR2_X1    g14416(.A1(new_n14328_), .A2(new_n14337_), .ZN(new_n14609_));
  NOR2_X1    g14417(.A1(\asqrt[10] ), .A2(new_n14609_), .ZN(new_n14610_));
  XOR2_X1    g14418(.A1(new_n14610_), .A2(new_n14135_), .Z(new_n14611_));
  AOI21_X1   g14419(.A1(new_n14332_), .A2(new_n14336_), .B(\asqrt[10] ), .ZN(new_n14612_));
  XOR2_X1    g14420(.A1(new_n14612_), .A2(new_n14138_), .Z(new_n14613_));
  INV_X1     g14421(.I(new_n14613_), .ZN(new_n14614_));
  AOI21_X1   g14422(.A1(new_n14318_), .A2(new_n14326_), .B(\asqrt[10] ), .ZN(new_n14615_));
  XOR2_X1    g14423(.A1(new_n14615_), .A2(new_n14142_), .Z(new_n14616_));
  INV_X1     g14424(.I(new_n14616_), .ZN(new_n14617_));
  XOR2_X1    g14425(.A1(new_n14309_), .A2(\asqrt[29] ), .Z(new_n14618_));
  NOR2_X1    g14426(.A1(\asqrt[10] ), .A2(new_n14618_), .ZN(new_n14619_));
  XOR2_X1    g14427(.A1(new_n14619_), .A2(new_n14144_), .Z(new_n14620_));
  NOR2_X1    g14428(.A1(new_n14307_), .A2(new_n14316_), .ZN(new_n14621_));
  NOR2_X1    g14429(.A1(\asqrt[10] ), .A2(new_n14621_), .ZN(new_n14622_));
  XOR2_X1    g14430(.A1(new_n14622_), .A2(new_n14147_), .Z(new_n14623_));
  AOI21_X1   g14431(.A1(new_n14311_), .A2(new_n14315_), .B(\asqrt[10] ), .ZN(new_n14624_));
  XOR2_X1    g14432(.A1(new_n14624_), .A2(new_n14150_), .Z(new_n14625_));
  INV_X1     g14433(.I(new_n14625_), .ZN(new_n14626_));
  AOI21_X1   g14434(.A1(new_n14297_), .A2(new_n14305_), .B(\asqrt[10] ), .ZN(new_n14627_));
  XOR2_X1    g14435(.A1(new_n14627_), .A2(new_n14154_), .Z(new_n14628_));
  INV_X1     g14436(.I(new_n14628_), .ZN(new_n14629_));
  XOR2_X1    g14437(.A1(new_n14288_), .A2(\asqrt[25] ), .Z(new_n14630_));
  NOR2_X1    g14438(.A1(\asqrt[10] ), .A2(new_n14630_), .ZN(new_n14631_));
  XOR2_X1    g14439(.A1(new_n14631_), .A2(new_n14156_), .Z(new_n14632_));
  NOR2_X1    g14440(.A1(new_n14286_), .A2(new_n14295_), .ZN(new_n14633_));
  NOR2_X1    g14441(.A1(\asqrt[10] ), .A2(new_n14633_), .ZN(new_n14634_));
  XOR2_X1    g14442(.A1(new_n14634_), .A2(new_n14159_), .Z(new_n14635_));
  AOI21_X1   g14443(.A1(new_n14290_), .A2(new_n14294_), .B(\asqrt[10] ), .ZN(new_n14636_));
  XOR2_X1    g14444(.A1(new_n14636_), .A2(new_n14162_), .Z(new_n14637_));
  INV_X1     g14445(.I(new_n14637_), .ZN(new_n14638_));
  AOI21_X1   g14446(.A1(new_n14276_), .A2(new_n14284_), .B(\asqrt[10] ), .ZN(new_n14639_));
  XOR2_X1    g14447(.A1(new_n14639_), .A2(new_n14166_), .Z(new_n14640_));
  INV_X1     g14448(.I(new_n14640_), .ZN(new_n14641_));
  XOR2_X1    g14449(.A1(new_n14267_), .A2(\asqrt[21] ), .Z(new_n14642_));
  NOR2_X1    g14450(.A1(\asqrt[10] ), .A2(new_n14642_), .ZN(new_n14643_));
  XOR2_X1    g14451(.A1(new_n14643_), .A2(new_n14168_), .Z(new_n14644_));
  NOR2_X1    g14452(.A1(new_n14265_), .A2(new_n14274_), .ZN(new_n14645_));
  NOR2_X1    g14453(.A1(\asqrt[10] ), .A2(new_n14645_), .ZN(new_n14646_));
  XOR2_X1    g14454(.A1(new_n14646_), .A2(new_n14171_), .Z(new_n14647_));
  AOI21_X1   g14455(.A1(new_n14269_), .A2(new_n14273_), .B(\asqrt[10] ), .ZN(new_n14648_));
  XOR2_X1    g14456(.A1(new_n14648_), .A2(new_n14174_), .Z(new_n14649_));
  INV_X1     g14457(.I(new_n14649_), .ZN(new_n14650_));
  AOI21_X1   g14458(.A1(new_n14255_), .A2(new_n14263_), .B(\asqrt[10] ), .ZN(new_n14651_));
  XOR2_X1    g14459(.A1(new_n14651_), .A2(new_n14178_), .Z(new_n14652_));
  INV_X1     g14460(.I(new_n14652_), .ZN(new_n14653_));
  XOR2_X1    g14461(.A1(new_n14246_), .A2(\asqrt[17] ), .Z(new_n14654_));
  NOR2_X1    g14462(.A1(\asqrt[10] ), .A2(new_n14654_), .ZN(new_n14655_));
  XOR2_X1    g14463(.A1(new_n14655_), .A2(new_n14180_), .Z(new_n14656_));
  NOR2_X1    g14464(.A1(new_n14244_), .A2(new_n14253_), .ZN(new_n14657_));
  NOR2_X1    g14465(.A1(\asqrt[10] ), .A2(new_n14657_), .ZN(new_n14658_));
  XOR2_X1    g14466(.A1(new_n14658_), .A2(new_n14183_), .Z(new_n14659_));
  AOI21_X1   g14467(.A1(new_n14248_), .A2(new_n14252_), .B(\asqrt[10] ), .ZN(new_n14660_));
  XOR2_X1    g14468(.A1(new_n14660_), .A2(new_n14186_), .Z(new_n14661_));
  INV_X1     g14469(.I(new_n14661_), .ZN(new_n14662_));
  AOI21_X1   g14470(.A1(new_n14234_), .A2(new_n14242_), .B(\asqrt[10] ), .ZN(new_n14663_));
  XOR2_X1    g14471(.A1(new_n14663_), .A2(new_n14193_), .Z(new_n14664_));
  INV_X1     g14472(.I(new_n14664_), .ZN(new_n14665_));
  AOI21_X1   g14473(.A1(new_n14225_), .A2(new_n14233_), .B(\asqrt[10] ), .ZN(new_n14666_));
  XOR2_X1    g14474(.A1(new_n14666_), .A2(new_n14210_), .Z(new_n14667_));
  NAND2_X1   g14475(.A1(\asqrt[11] ), .A2(new_n14211_), .ZN(new_n14668_));
  NOR2_X1    g14476(.A1(new_n14222_), .A2(\a[22] ), .ZN(new_n14669_));
  AOI22_X1   g14477(.A1(new_n14668_), .A2(new_n14222_), .B1(\asqrt[11] ), .B2(new_n14669_), .ZN(new_n14670_));
  AOI21_X1   g14478(.A1(\asqrt[11] ), .A2(\a[22] ), .B(new_n14219_), .ZN(new_n14671_));
  NOR2_X1    g14479(.A1(new_n14229_), .A2(new_n14671_), .ZN(new_n14672_));
  NOR2_X1    g14480(.A1(\asqrt[10] ), .A2(new_n14672_), .ZN(new_n14673_));
  XOR2_X1    g14481(.A1(new_n14673_), .A2(new_n14670_), .Z(new_n14674_));
  NOR2_X1    g14482(.A1(new_n14520_), .A2(new_n14516_), .ZN(new_n14675_));
  AOI21_X1   g14483(.A1(new_n14499_), .A2(new_n14496_), .B(\asqrt[62] ), .ZN(new_n14676_));
  NOR3_X1    g14484(.A1(new_n14520_), .A2(new_n201_), .A3(new_n14516_), .ZN(new_n14677_));
  OAI22_X1   g14485(.A1(new_n14676_), .A2(new_n14677_), .B1(new_n14675_), .B2(new_n14525_), .ZN(new_n14678_));
  AOI21_X1   g14486(.A1(new_n14678_), .A2(new_n14452_), .B(new_n14529_), .ZN(new_n14679_));
  AOI21_X1   g14487(.A1(new_n14675_), .A2(new_n201_), .B(new_n14526_), .ZN(new_n14680_));
  NOR2_X1    g14488(.A1(new_n14675_), .A2(new_n201_), .ZN(new_n14681_));
  NOR3_X1    g14489(.A1(new_n14680_), .A2(new_n14681_), .A3(new_n14452_), .ZN(new_n14682_));
  NOR3_X1    g14490(.A1(new_n14679_), .A2(\asqrt[63] ), .A3(new_n14682_), .ZN(new_n14683_));
  NAND4_X1   g14491(.A1(new_n14683_), .A2(\asqrt[11] ), .A3(new_n14538_), .A4(new_n14540_), .ZN(new_n14684_));
  NAND2_X1   g14492(.A1(\asqrt[10] ), .A2(new_n14212_), .ZN(new_n14685_));
  AOI21_X1   g14493(.A1(new_n14684_), .A2(new_n14685_), .B(\a[22] ), .ZN(new_n14686_));
  NAND2_X1   g14494(.A1(new_n14531_), .A2(new_n193_), .ZN(new_n14687_));
  NAND3_X1   g14495(.A1(new_n14538_), .A2(new_n14540_), .A3(\asqrt[11] ), .ZN(new_n14688_));
  NOR3_X1    g14496(.A1(new_n14687_), .A2(new_n14682_), .A3(new_n14688_), .ZN(new_n14689_));
  NOR4_X1    g14497(.A1(new_n14679_), .A2(\asqrt[63] ), .A3(new_n14682_), .A4(new_n14541_), .ZN(new_n14690_));
  NOR2_X1    g14498(.A1(new_n14690_), .A2(new_n14214_), .ZN(new_n14691_));
  NOR3_X1    g14499(.A1(new_n14691_), .A2(new_n14689_), .A3(new_n14211_), .ZN(new_n14692_));
  OR2_X2     g14500(.A1(new_n14686_), .A2(new_n14692_), .Z(new_n14693_));
  NOR2_X1    g14501(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n14694_));
  INV_X1     g14502(.I(new_n14694_), .ZN(new_n14695_));
  NAND3_X1   g14503(.A1(\asqrt[10] ), .A2(\a[20] ), .A3(new_n14695_), .ZN(new_n14696_));
  INV_X1     g14504(.I(\a[20] ), .ZN(new_n14697_));
  OAI21_X1   g14505(.A1(\asqrt[10] ), .A2(new_n14697_), .B(new_n14694_), .ZN(new_n14698_));
  AOI21_X1   g14506(.A1(new_n14698_), .A2(new_n14696_), .B(new_n14207_), .ZN(new_n14699_));
  NOR3_X1    g14507(.A1(new_n14198_), .A2(\asqrt[63] ), .A3(new_n14201_), .ZN(new_n14700_));
  NAND2_X1   g14508(.A1(new_n14694_), .A2(new_n14697_), .ZN(new_n14701_));
  NAND3_X1   g14509(.A1(new_n14063_), .A2(new_n14065_), .A3(new_n14701_), .ZN(new_n14702_));
  NAND2_X1   g14510(.A1(new_n14700_), .A2(new_n14702_), .ZN(new_n14703_));
  NAND3_X1   g14511(.A1(\asqrt[10] ), .A2(\a[20] ), .A3(new_n14703_), .ZN(new_n14704_));
  INV_X1     g14512(.I(\a[21] ), .ZN(new_n14705_));
  NAND3_X1   g14513(.A1(\asqrt[10] ), .A2(new_n14697_), .A3(new_n14705_), .ZN(new_n14706_));
  OAI21_X1   g14514(.A1(new_n14690_), .A2(\a[20] ), .B(\a[21] ), .ZN(new_n14707_));
  NAND3_X1   g14515(.A1(new_n14704_), .A2(new_n14707_), .A3(new_n14706_), .ZN(new_n14708_));
  NOR3_X1    g14516(.A1(new_n14708_), .A2(new_n14699_), .A3(\asqrt[12] ), .ZN(new_n14709_));
  OAI21_X1   g14517(.A1(new_n14708_), .A2(new_n14699_), .B(\asqrt[12] ), .ZN(new_n14710_));
  OAI21_X1   g14518(.A1(new_n14693_), .A2(new_n14709_), .B(new_n14710_), .ZN(new_n14711_));
  OAI21_X1   g14519(.A1(new_n14711_), .A2(\asqrt[13] ), .B(new_n14674_), .ZN(new_n14712_));
  NAND2_X1   g14520(.A1(new_n14711_), .A2(\asqrt[13] ), .ZN(new_n14713_));
  NAND3_X1   g14521(.A1(new_n14712_), .A2(new_n14713_), .A3(new_n12733_), .ZN(new_n14714_));
  AOI21_X1   g14522(.A1(new_n14712_), .A2(new_n14713_), .B(new_n12733_), .ZN(new_n14715_));
  AOI21_X1   g14523(.A1(new_n14667_), .A2(new_n14714_), .B(new_n14715_), .ZN(new_n14716_));
  AOI21_X1   g14524(.A1(new_n14716_), .A2(new_n12283_), .B(new_n14665_), .ZN(new_n14717_));
  NAND2_X1   g14525(.A1(new_n14714_), .A2(new_n14667_), .ZN(new_n14718_));
  INV_X1     g14526(.I(new_n14674_), .ZN(new_n14719_));
  NOR2_X1    g14527(.A1(new_n14686_), .A2(new_n14692_), .ZN(new_n14720_));
  NOR3_X1    g14528(.A1(new_n14690_), .A2(new_n14697_), .A3(new_n14694_), .ZN(new_n14721_));
  AOI21_X1   g14529(.A1(new_n14690_), .A2(\a[20] ), .B(new_n14695_), .ZN(new_n14722_));
  OAI21_X1   g14530(.A1(new_n14721_), .A2(new_n14722_), .B(\asqrt[11] ), .ZN(new_n14723_));
  INV_X1     g14531(.I(new_n14703_), .ZN(new_n14724_));
  NOR3_X1    g14532(.A1(new_n14690_), .A2(new_n14697_), .A3(new_n14724_), .ZN(new_n14725_));
  NOR3_X1    g14533(.A1(new_n14690_), .A2(\a[20] ), .A3(\a[21] ), .ZN(new_n14726_));
  AOI21_X1   g14534(.A1(\asqrt[10] ), .A2(new_n14697_), .B(new_n14705_), .ZN(new_n14727_));
  NOR3_X1    g14535(.A1(new_n14725_), .A2(new_n14726_), .A3(new_n14727_), .ZN(new_n14728_));
  NAND3_X1   g14536(.A1(new_n14728_), .A2(new_n14723_), .A3(new_n13690_), .ZN(new_n14729_));
  AOI21_X1   g14537(.A1(new_n14728_), .A2(new_n14723_), .B(new_n13690_), .ZN(new_n14730_));
  AOI21_X1   g14538(.A1(new_n14720_), .A2(new_n14729_), .B(new_n14730_), .ZN(new_n14731_));
  AOI21_X1   g14539(.A1(new_n14731_), .A2(new_n13228_), .B(new_n14719_), .ZN(new_n14732_));
  NAND2_X1   g14540(.A1(new_n14729_), .A2(new_n14720_), .ZN(new_n14733_));
  AOI21_X1   g14541(.A1(new_n14733_), .A2(new_n14710_), .B(new_n13228_), .ZN(new_n14734_));
  OAI21_X1   g14542(.A1(new_n14732_), .A2(new_n14734_), .B(\asqrt[14] ), .ZN(new_n14735_));
  AOI21_X1   g14543(.A1(new_n14718_), .A2(new_n14735_), .B(new_n12283_), .ZN(new_n14736_));
  NOR3_X1    g14544(.A1(new_n14717_), .A2(\asqrt[16] ), .A3(new_n14736_), .ZN(new_n14737_));
  OAI21_X1   g14545(.A1(new_n14717_), .A2(new_n14736_), .B(\asqrt[16] ), .ZN(new_n14738_));
  OAI21_X1   g14546(.A1(new_n14662_), .A2(new_n14737_), .B(new_n14738_), .ZN(new_n14739_));
  OAI21_X1   g14547(.A1(new_n14739_), .A2(\asqrt[17] ), .B(new_n14659_), .ZN(new_n14740_));
  NAND2_X1   g14548(.A1(new_n14739_), .A2(\asqrt[17] ), .ZN(new_n14741_));
  NAND3_X1   g14549(.A1(new_n14740_), .A2(new_n14741_), .A3(new_n10914_), .ZN(new_n14742_));
  AOI21_X1   g14550(.A1(new_n14740_), .A2(new_n14741_), .B(new_n10914_), .ZN(new_n14743_));
  AOI21_X1   g14551(.A1(new_n14656_), .A2(new_n14742_), .B(new_n14743_), .ZN(new_n14744_));
  AOI21_X1   g14552(.A1(new_n14744_), .A2(new_n10497_), .B(new_n14653_), .ZN(new_n14745_));
  NAND2_X1   g14553(.A1(new_n14742_), .A2(new_n14656_), .ZN(new_n14746_));
  INV_X1     g14554(.I(new_n14659_), .ZN(new_n14747_));
  INV_X1     g14555(.I(new_n14667_), .ZN(new_n14748_));
  NOR3_X1    g14556(.A1(new_n14732_), .A2(\asqrt[14] ), .A3(new_n14734_), .ZN(new_n14749_));
  OAI21_X1   g14557(.A1(new_n14748_), .A2(new_n14749_), .B(new_n14735_), .ZN(new_n14750_));
  OAI21_X1   g14558(.A1(new_n14750_), .A2(\asqrt[15] ), .B(new_n14664_), .ZN(new_n14751_));
  NAND2_X1   g14559(.A1(new_n14750_), .A2(\asqrt[15] ), .ZN(new_n14752_));
  NAND3_X1   g14560(.A1(new_n14751_), .A2(new_n14752_), .A3(new_n11802_), .ZN(new_n14753_));
  AOI21_X1   g14561(.A1(new_n14751_), .A2(new_n14752_), .B(new_n11802_), .ZN(new_n14754_));
  AOI21_X1   g14562(.A1(new_n14661_), .A2(new_n14753_), .B(new_n14754_), .ZN(new_n14755_));
  AOI21_X1   g14563(.A1(new_n14755_), .A2(new_n11373_), .B(new_n14747_), .ZN(new_n14756_));
  NAND2_X1   g14564(.A1(new_n14753_), .A2(new_n14661_), .ZN(new_n14757_));
  AOI21_X1   g14565(.A1(new_n14757_), .A2(new_n14738_), .B(new_n11373_), .ZN(new_n14758_));
  OAI21_X1   g14566(.A1(new_n14756_), .A2(new_n14758_), .B(\asqrt[18] ), .ZN(new_n14759_));
  AOI21_X1   g14567(.A1(new_n14746_), .A2(new_n14759_), .B(new_n10497_), .ZN(new_n14760_));
  NOR3_X1    g14568(.A1(new_n14745_), .A2(\asqrt[20] ), .A3(new_n14760_), .ZN(new_n14761_));
  OAI21_X1   g14569(.A1(new_n14745_), .A2(new_n14760_), .B(\asqrt[20] ), .ZN(new_n14762_));
  OAI21_X1   g14570(.A1(new_n14650_), .A2(new_n14761_), .B(new_n14762_), .ZN(new_n14763_));
  OAI21_X1   g14571(.A1(new_n14763_), .A2(\asqrt[21] ), .B(new_n14647_), .ZN(new_n14764_));
  NAND2_X1   g14572(.A1(new_n14763_), .A2(\asqrt[21] ), .ZN(new_n14765_));
  NAND3_X1   g14573(.A1(new_n14764_), .A2(new_n14765_), .A3(new_n9233_), .ZN(new_n14766_));
  AOI21_X1   g14574(.A1(new_n14764_), .A2(new_n14765_), .B(new_n9233_), .ZN(new_n14767_));
  AOI21_X1   g14575(.A1(new_n14644_), .A2(new_n14766_), .B(new_n14767_), .ZN(new_n14768_));
  AOI21_X1   g14576(.A1(new_n14768_), .A2(new_n8849_), .B(new_n14641_), .ZN(new_n14769_));
  NAND2_X1   g14577(.A1(new_n14766_), .A2(new_n14644_), .ZN(new_n14770_));
  INV_X1     g14578(.I(new_n14647_), .ZN(new_n14771_));
  INV_X1     g14579(.I(new_n14656_), .ZN(new_n14772_));
  NOR3_X1    g14580(.A1(new_n14756_), .A2(\asqrt[18] ), .A3(new_n14758_), .ZN(new_n14773_));
  OAI21_X1   g14581(.A1(new_n14772_), .A2(new_n14773_), .B(new_n14759_), .ZN(new_n14774_));
  OAI21_X1   g14582(.A1(new_n14774_), .A2(\asqrt[19] ), .B(new_n14652_), .ZN(new_n14775_));
  NAND2_X1   g14583(.A1(new_n14774_), .A2(\asqrt[19] ), .ZN(new_n14776_));
  NAND3_X1   g14584(.A1(new_n14775_), .A2(new_n14776_), .A3(new_n10052_), .ZN(new_n14777_));
  AOI21_X1   g14585(.A1(new_n14775_), .A2(new_n14776_), .B(new_n10052_), .ZN(new_n14778_));
  AOI21_X1   g14586(.A1(new_n14649_), .A2(new_n14777_), .B(new_n14778_), .ZN(new_n14779_));
  AOI21_X1   g14587(.A1(new_n14779_), .A2(new_n9656_), .B(new_n14771_), .ZN(new_n14780_));
  NAND2_X1   g14588(.A1(new_n14777_), .A2(new_n14649_), .ZN(new_n14781_));
  AOI21_X1   g14589(.A1(new_n14781_), .A2(new_n14762_), .B(new_n9656_), .ZN(new_n14782_));
  OAI21_X1   g14590(.A1(new_n14780_), .A2(new_n14782_), .B(\asqrt[22] ), .ZN(new_n14783_));
  AOI21_X1   g14591(.A1(new_n14770_), .A2(new_n14783_), .B(new_n8849_), .ZN(new_n14784_));
  NOR3_X1    g14592(.A1(new_n14769_), .A2(\asqrt[24] ), .A3(new_n14784_), .ZN(new_n14785_));
  OAI21_X1   g14593(.A1(new_n14769_), .A2(new_n14784_), .B(\asqrt[24] ), .ZN(new_n14786_));
  OAI21_X1   g14594(.A1(new_n14638_), .A2(new_n14785_), .B(new_n14786_), .ZN(new_n14787_));
  OAI21_X1   g14595(.A1(new_n14787_), .A2(\asqrt[25] ), .B(new_n14635_), .ZN(new_n14788_));
  NAND2_X1   g14596(.A1(new_n14787_), .A2(\asqrt[25] ), .ZN(new_n14789_));
  NAND3_X1   g14597(.A1(new_n14788_), .A2(new_n14789_), .A3(new_n7690_), .ZN(new_n14790_));
  AOI21_X1   g14598(.A1(new_n14788_), .A2(new_n14789_), .B(new_n7690_), .ZN(new_n14791_));
  AOI21_X1   g14599(.A1(new_n14632_), .A2(new_n14790_), .B(new_n14791_), .ZN(new_n14792_));
  AOI21_X1   g14600(.A1(new_n14792_), .A2(new_n7331_), .B(new_n14629_), .ZN(new_n14793_));
  NAND2_X1   g14601(.A1(new_n14790_), .A2(new_n14632_), .ZN(new_n14794_));
  INV_X1     g14602(.I(new_n14635_), .ZN(new_n14795_));
  INV_X1     g14603(.I(new_n14644_), .ZN(new_n14796_));
  NOR3_X1    g14604(.A1(new_n14780_), .A2(\asqrt[22] ), .A3(new_n14782_), .ZN(new_n14797_));
  OAI21_X1   g14605(.A1(new_n14796_), .A2(new_n14797_), .B(new_n14783_), .ZN(new_n14798_));
  OAI21_X1   g14606(.A1(new_n14798_), .A2(\asqrt[23] ), .B(new_n14640_), .ZN(new_n14799_));
  NAND2_X1   g14607(.A1(new_n14798_), .A2(\asqrt[23] ), .ZN(new_n14800_));
  NAND3_X1   g14608(.A1(new_n14799_), .A2(new_n14800_), .A3(new_n8440_), .ZN(new_n14801_));
  AOI21_X1   g14609(.A1(new_n14799_), .A2(new_n14800_), .B(new_n8440_), .ZN(new_n14802_));
  AOI21_X1   g14610(.A1(new_n14637_), .A2(new_n14801_), .B(new_n14802_), .ZN(new_n14803_));
  AOI21_X1   g14611(.A1(new_n14803_), .A2(new_n8077_), .B(new_n14795_), .ZN(new_n14804_));
  NAND2_X1   g14612(.A1(new_n14801_), .A2(new_n14637_), .ZN(new_n14805_));
  AOI21_X1   g14613(.A1(new_n14805_), .A2(new_n14786_), .B(new_n8077_), .ZN(new_n14806_));
  OAI21_X1   g14614(.A1(new_n14804_), .A2(new_n14806_), .B(\asqrt[26] ), .ZN(new_n14807_));
  AOI21_X1   g14615(.A1(new_n14794_), .A2(new_n14807_), .B(new_n7331_), .ZN(new_n14808_));
  NOR3_X1    g14616(.A1(new_n14793_), .A2(\asqrt[28] ), .A3(new_n14808_), .ZN(new_n14809_));
  OAI21_X1   g14617(.A1(new_n14793_), .A2(new_n14808_), .B(\asqrt[28] ), .ZN(new_n14810_));
  OAI21_X1   g14618(.A1(new_n14626_), .A2(new_n14809_), .B(new_n14810_), .ZN(new_n14811_));
  OAI21_X1   g14619(.A1(new_n14811_), .A2(\asqrt[29] ), .B(new_n14623_), .ZN(new_n14812_));
  NAND2_X1   g14620(.A1(new_n14811_), .A2(\asqrt[29] ), .ZN(new_n14813_));
  NAND3_X1   g14621(.A1(new_n14812_), .A2(new_n14813_), .A3(new_n6275_), .ZN(new_n14814_));
  AOI21_X1   g14622(.A1(new_n14812_), .A2(new_n14813_), .B(new_n6275_), .ZN(new_n14815_));
  AOI21_X1   g14623(.A1(new_n14620_), .A2(new_n14814_), .B(new_n14815_), .ZN(new_n14816_));
  AOI21_X1   g14624(.A1(new_n14816_), .A2(new_n5947_), .B(new_n14617_), .ZN(new_n14817_));
  NAND2_X1   g14625(.A1(new_n14814_), .A2(new_n14620_), .ZN(new_n14818_));
  INV_X1     g14626(.I(new_n14623_), .ZN(new_n14819_));
  INV_X1     g14627(.I(new_n14632_), .ZN(new_n14820_));
  NOR3_X1    g14628(.A1(new_n14804_), .A2(\asqrt[26] ), .A3(new_n14806_), .ZN(new_n14821_));
  OAI21_X1   g14629(.A1(new_n14820_), .A2(new_n14821_), .B(new_n14807_), .ZN(new_n14822_));
  OAI21_X1   g14630(.A1(new_n14822_), .A2(\asqrt[27] ), .B(new_n14628_), .ZN(new_n14823_));
  NAND2_X1   g14631(.A1(new_n14822_), .A2(\asqrt[27] ), .ZN(new_n14824_));
  NAND3_X1   g14632(.A1(new_n14823_), .A2(new_n14824_), .A3(new_n6966_), .ZN(new_n14825_));
  AOI21_X1   g14633(.A1(new_n14823_), .A2(new_n14824_), .B(new_n6966_), .ZN(new_n14826_));
  AOI21_X1   g14634(.A1(new_n14625_), .A2(new_n14825_), .B(new_n14826_), .ZN(new_n14827_));
  AOI21_X1   g14635(.A1(new_n14827_), .A2(new_n6636_), .B(new_n14819_), .ZN(new_n14828_));
  NAND2_X1   g14636(.A1(new_n14825_), .A2(new_n14625_), .ZN(new_n14829_));
  AOI21_X1   g14637(.A1(new_n14829_), .A2(new_n14810_), .B(new_n6636_), .ZN(new_n14830_));
  OAI21_X1   g14638(.A1(new_n14828_), .A2(new_n14830_), .B(\asqrt[30] ), .ZN(new_n14831_));
  AOI21_X1   g14639(.A1(new_n14818_), .A2(new_n14831_), .B(new_n5947_), .ZN(new_n14832_));
  NOR3_X1    g14640(.A1(new_n14817_), .A2(\asqrt[32] ), .A3(new_n14832_), .ZN(new_n14833_));
  OAI21_X1   g14641(.A1(new_n14817_), .A2(new_n14832_), .B(\asqrt[32] ), .ZN(new_n14834_));
  OAI21_X1   g14642(.A1(new_n14614_), .A2(new_n14833_), .B(new_n14834_), .ZN(new_n14835_));
  OAI21_X1   g14643(.A1(new_n14835_), .A2(\asqrt[33] ), .B(new_n14611_), .ZN(new_n14836_));
  NAND2_X1   g14644(.A1(new_n14835_), .A2(\asqrt[33] ), .ZN(new_n14837_));
  NAND3_X1   g14645(.A1(new_n14836_), .A2(new_n14837_), .A3(new_n5029_), .ZN(new_n14838_));
  AOI21_X1   g14646(.A1(new_n14836_), .A2(new_n14837_), .B(new_n5029_), .ZN(new_n14839_));
  AOI21_X1   g14647(.A1(new_n14608_), .A2(new_n14838_), .B(new_n14839_), .ZN(new_n14840_));
  AOI21_X1   g14648(.A1(new_n14840_), .A2(new_n4751_), .B(new_n14605_), .ZN(new_n14841_));
  NAND2_X1   g14649(.A1(new_n14838_), .A2(new_n14608_), .ZN(new_n14842_));
  INV_X1     g14650(.I(new_n14611_), .ZN(new_n14843_));
  INV_X1     g14651(.I(new_n14620_), .ZN(new_n14844_));
  NOR3_X1    g14652(.A1(new_n14828_), .A2(\asqrt[30] ), .A3(new_n14830_), .ZN(new_n14845_));
  OAI21_X1   g14653(.A1(new_n14844_), .A2(new_n14845_), .B(new_n14831_), .ZN(new_n14846_));
  OAI21_X1   g14654(.A1(new_n14846_), .A2(\asqrt[31] ), .B(new_n14616_), .ZN(new_n14847_));
  NAND2_X1   g14655(.A1(new_n14846_), .A2(\asqrt[31] ), .ZN(new_n14848_));
  NAND3_X1   g14656(.A1(new_n14847_), .A2(new_n14848_), .A3(new_n5643_), .ZN(new_n14849_));
  AOI21_X1   g14657(.A1(new_n14847_), .A2(new_n14848_), .B(new_n5643_), .ZN(new_n14850_));
  AOI21_X1   g14658(.A1(new_n14613_), .A2(new_n14849_), .B(new_n14850_), .ZN(new_n14851_));
  AOI21_X1   g14659(.A1(new_n14851_), .A2(new_n5336_), .B(new_n14843_), .ZN(new_n14852_));
  NAND2_X1   g14660(.A1(new_n14849_), .A2(new_n14613_), .ZN(new_n14853_));
  AOI21_X1   g14661(.A1(new_n14853_), .A2(new_n14834_), .B(new_n5336_), .ZN(new_n14854_));
  OAI21_X1   g14662(.A1(new_n14852_), .A2(new_n14854_), .B(\asqrt[34] ), .ZN(new_n14855_));
  AOI21_X1   g14663(.A1(new_n14842_), .A2(new_n14855_), .B(new_n4751_), .ZN(new_n14856_));
  NOR3_X1    g14664(.A1(new_n14841_), .A2(\asqrt[36] ), .A3(new_n14856_), .ZN(new_n14857_));
  OAI21_X1   g14665(.A1(new_n14841_), .A2(new_n14856_), .B(\asqrt[36] ), .ZN(new_n14858_));
  OAI21_X1   g14666(.A1(new_n14602_), .A2(new_n14857_), .B(new_n14858_), .ZN(new_n14859_));
  OAI21_X1   g14667(.A1(new_n14859_), .A2(\asqrt[37] ), .B(new_n14599_), .ZN(new_n14860_));
  NAND2_X1   g14668(.A1(new_n14859_), .A2(\asqrt[37] ), .ZN(new_n14861_));
  NAND3_X1   g14669(.A1(new_n14860_), .A2(new_n14861_), .A3(new_n3925_), .ZN(new_n14862_));
  AOI21_X1   g14670(.A1(new_n14860_), .A2(new_n14861_), .B(new_n3925_), .ZN(new_n14863_));
  AOI21_X1   g14671(.A1(new_n14596_), .A2(new_n14862_), .B(new_n14863_), .ZN(new_n14864_));
  AOI21_X1   g14672(.A1(new_n14864_), .A2(new_n3681_), .B(new_n14593_), .ZN(new_n14865_));
  NAND2_X1   g14673(.A1(new_n14862_), .A2(new_n14596_), .ZN(new_n14866_));
  INV_X1     g14674(.I(new_n14599_), .ZN(new_n14867_));
  INV_X1     g14675(.I(new_n14608_), .ZN(new_n14868_));
  NOR3_X1    g14676(.A1(new_n14852_), .A2(\asqrt[34] ), .A3(new_n14854_), .ZN(new_n14869_));
  OAI21_X1   g14677(.A1(new_n14868_), .A2(new_n14869_), .B(new_n14855_), .ZN(new_n14870_));
  OAI21_X1   g14678(.A1(new_n14870_), .A2(\asqrt[35] ), .B(new_n14604_), .ZN(new_n14871_));
  NAND2_X1   g14679(.A1(new_n14870_), .A2(\asqrt[35] ), .ZN(new_n14872_));
  NAND3_X1   g14680(.A1(new_n14871_), .A2(new_n14872_), .A3(new_n4461_), .ZN(new_n14873_));
  AOI21_X1   g14681(.A1(new_n14871_), .A2(new_n14872_), .B(new_n4461_), .ZN(new_n14874_));
  AOI21_X1   g14682(.A1(new_n14601_), .A2(new_n14873_), .B(new_n14874_), .ZN(new_n14875_));
  AOI21_X1   g14683(.A1(new_n14875_), .A2(new_n4196_), .B(new_n14867_), .ZN(new_n14876_));
  NAND2_X1   g14684(.A1(new_n14873_), .A2(new_n14601_), .ZN(new_n14877_));
  AOI21_X1   g14685(.A1(new_n14877_), .A2(new_n14858_), .B(new_n4196_), .ZN(new_n14878_));
  OAI21_X1   g14686(.A1(new_n14876_), .A2(new_n14878_), .B(\asqrt[38] ), .ZN(new_n14879_));
  AOI21_X1   g14687(.A1(new_n14866_), .A2(new_n14879_), .B(new_n3681_), .ZN(new_n14880_));
  NOR3_X1    g14688(.A1(new_n14865_), .A2(\asqrt[40] ), .A3(new_n14880_), .ZN(new_n14881_));
  OAI21_X1   g14689(.A1(new_n14865_), .A2(new_n14880_), .B(\asqrt[40] ), .ZN(new_n14882_));
  OAI21_X1   g14690(.A1(new_n14590_), .A2(new_n14881_), .B(new_n14882_), .ZN(new_n14883_));
  OAI21_X1   g14691(.A1(new_n14883_), .A2(\asqrt[41] ), .B(new_n14587_), .ZN(new_n14884_));
  NAND2_X1   g14692(.A1(new_n14883_), .A2(\asqrt[41] ), .ZN(new_n14885_));
  NAND3_X1   g14693(.A1(new_n14884_), .A2(new_n14885_), .A3(new_n2960_), .ZN(new_n14886_));
  AOI21_X1   g14694(.A1(new_n14884_), .A2(new_n14885_), .B(new_n2960_), .ZN(new_n14887_));
  AOI21_X1   g14695(.A1(new_n14584_), .A2(new_n14886_), .B(new_n14887_), .ZN(new_n14888_));
  AOI21_X1   g14696(.A1(new_n14888_), .A2(new_n2749_), .B(new_n14581_), .ZN(new_n14889_));
  NAND2_X1   g14697(.A1(new_n14886_), .A2(new_n14584_), .ZN(new_n14890_));
  INV_X1     g14698(.I(new_n14587_), .ZN(new_n14891_));
  INV_X1     g14699(.I(new_n14596_), .ZN(new_n14892_));
  NOR3_X1    g14700(.A1(new_n14876_), .A2(\asqrt[38] ), .A3(new_n14878_), .ZN(new_n14893_));
  OAI21_X1   g14701(.A1(new_n14892_), .A2(new_n14893_), .B(new_n14879_), .ZN(new_n14894_));
  OAI21_X1   g14702(.A1(new_n14894_), .A2(\asqrt[39] ), .B(new_n14592_), .ZN(new_n14895_));
  NAND2_X1   g14703(.A1(new_n14894_), .A2(\asqrt[39] ), .ZN(new_n14896_));
  NAND3_X1   g14704(.A1(new_n14895_), .A2(new_n14896_), .A3(new_n3427_), .ZN(new_n14897_));
  AOI21_X1   g14705(.A1(new_n14895_), .A2(new_n14896_), .B(new_n3427_), .ZN(new_n14898_));
  AOI21_X1   g14706(.A1(new_n14589_), .A2(new_n14897_), .B(new_n14898_), .ZN(new_n14899_));
  AOI21_X1   g14707(.A1(new_n14899_), .A2(new_n3195_), .B(new_n14891_), .ZN(new_n14900_));
  NAND2_X1   g14708(.A1(new_n14897_), .A2(new_n14589_), .ZN(new_n14901_));
  AOI21_X1   g14709(.A1(new_n14901_), .A2(new_n14882_), .B(new_n3195_), .ZN(new_n14902_));
  OAI21_X1   g14710(.A1(new_n14900_), .A2(new_n14902_), .B(\asqrt[42] ), .ZN(new_n14903_));
  AOI21_X1   g14711(.A1(new_n14890_), .A2(new_n14903_), .B(new_n2749_), .ZN(new_n14904_));
  NOR3_X1    g14712(.A1(new_n14889_), .A2(\asqrt[44] ), .A3(new_n14904_), .ZN(new_n14905_));
  OAI21_X1   g14713(.A1(new_n14889_), .A2(new_n14904_), .B(\asqrt[44] ), .ZN(new_n14906_));
  OAI21_X1   g14714(.A1(new_n14578_), .A2(new_n14905_), .B(new_n14906_), .ZN(new_n14907_));
  OAI21_X1   g14715(.A1(new_n14907_), .A2(\asqrt[45] ), .B(new_n14575_), .ZN(new_n14908_));
  NAND2_X1   g14716(.A1(new_n14907_), .A2(\asqrt[45] ), .ZN(new_n14909_));
  NAND3_X1   g14717(.A1(new_n14908_), .A2(new_n14909_), .A3(new_n2134_), .ZN(new_n14910_));
  AOI21_X1   g14718(.A1(new_n14908_), .A2(new_n14909_), .B(new_n2134_), .ZN(new_n14911_));
  AOI21_X1   g14719(.A1(new_n14572_), .A2(new_n14910_), .B(new_n14911_), .ZN(new_n14912_));
  AOI21_X1   g14720(.A1(new_n14912_), .A2(new_n1953_), .B(new_n14569_), .ZN(new_n14913_));
  NAND2_X1   g14721(.A1(new_n14910_), .A2(new_n14572_), .ZN(new_n14914_));
  INV_X1     g14722(.I(new_n14575_), .ZN(new_n14915_));
  INV_X1     g14723(.I(new_n14584_), .ZN(new_n14916_));
  NOR3_X1    g14724(.A1(new_n14900_), .A2(\asqrt[42] ), .A3(new_n14902_), .ZN(new_n14917_));
  OAI21_X1   g14725(.A1(new_n14916_), .A2(new_n14917_), .B(new_n14903_), .ZN(new_n14918_));
  OAI21_X1   g14726(.A1(new_n14918_), .A2(\asqrt[43] ), .B(new_n14580_), .ZN(new_n14919_));
  NAND2_X1   g14727(.A1(new_n14918_), .A2(\asqrt[43] ), .ZN(new_n14920_));
  NAND3_X1   g14728(.A1(new_n14919_), .A2(new_n14920_), .A3(new_n2531_), .ZN(new_n14921_));
  AOI21_X1   g14729(.A1(new_n14919_), .A2(new_n14920_), .B(new_n2531_), .ZN(new_n14922_));
  AOI21_X1   g14730(.A1(new_n14577_), .A2(new_n14921_), .B(new_n14922_), .ZN(new_n14923_));
  AOI21_X1   g14731(.A1(new_n14923_), .A2(new_n2332_), .B(new_n14915_), .ZN(new_n14924_));
  NAND2_X1   g14732(.A1(new_n14921_), .A2(new_n14577_), .ZN(new_n14925_));
  AOI21_X1   g14733(.A1(new_n14925_), .A2(new_n14906_), .B(new_n2332_), .ZN(new_n14926_));
  OAI21_X1   g14734(.A1(new_n14924_), .A2(new_n14926_), .B(\asqrt[46] ), .ZN(new_n14927_));
  AOI21_X1   g14735(.A1(new_n14914_), .A2(new_n14927_), .B(new_n1953_), .ZN(new_n14928_));
  NOR3_X1    g14736(.A1(new_n14913_), .A2(\asqrt[48] ), .A3(new_n14928_), .ZN(new_n14929_));
  OAI21_X1   g14737(.A1(new_n14913_), .A2(new_n14928_), .B(\asqrt[48] ), .ZN(new_n14930_));
  OAI21_X1   g14738(.A1(new_n14566_), .A2(new_n14929_), .B(new_n14930_), .ZN(new_n14931_));
  OAI21_X1   g14739(.A1(new_n14931_), .A2(\asqrt[49] ), .B(new_n14563_), .ZN(new_n14932_));
  NAND2_X1   g14740(.A1(new_n14931_), .A2(\asqrt[49] ), .ZN(new_n14933_));
  NAND3_X1   g14741(.A1(new_n14932_), .A2(new_n14933_), .A3(new_n1463_), .ZN(new_n14934_));
  AOI21_X1   g14742(.A1(new_n14932_), .A2(new_n14933_), .B(new_n1463_), .ZN(new_n14935_));
  AOI21_X1   g14743(.A1(new_n14560_), .A2(new_n14934_), .B(new_n14935_), .ZN(new_n14936_));
  AOI21_X1   g14744(.A1(new_n14936_), .A2(new_n1305_), .B(new_n14557_), .ZN(new_n14937_));
  NAND2_X1   g14745(.A1(new_n14934_), .A2(new_n14560_), .ZN(new_n14938_));
  INV_X1     g14746(.I(new_n14563_), .ZN(new_n14939_));
  INV_X1     g14747(.I(new_n14572_), .ZN(new_n14940_));
  NOR3_X1    g14748(.A1(new_n14924_), .A2(\asqrt[46] ), .A3(new_n14926_), .ZN(new_n14941_));
  OAI21_X1   g14749(.A1(new_n14940_), .A2(new_n14941_), .B(new_n14927_), .ZN(new_n14942_));
  OAI21_X1   g14750(.A1(new_n14942_), .A2(\asqrt[47] ), .B(new_n14568_), .ZN(new_n14943_));
  NAND2_X1   g14751(.A1(new_n14942_), .A2(\asqrt[47] ), .ZN(new_n14944_));
  NAND3_X1   g14752(.A1(new_n14943_), .A2(new_n14944_), .A3(new_n1778_), .ZN(new_n14945_));
  AOI21_X1   g14753(.A1(new_n14943_), .A2(new_n14944_), .B(new_n1778_), .ZN(new_n14946_));
  AOI21_X1   g14754(.A1(new_n14565_), .A2(new_n14945_), .B(new_n14946_), .ZN(new_n14947_));
  AOI21_X1   g14755(.A1(new_n14947_), .A2(new_n1632_), .B(new_n14939_), .ZN(new_n14948_));
  NAND2_X1   g14756(.A1(new_n14945_), .A2(new_n14565_), .ZN(new_n14949_));
  AOI21_X1   g14757(.A1(new_n14949_), .A2(new_n14930_), .B(new_n1632_), .ZN(new_n14950_));
  OAI21_X1   g14758(.A1(new_n14948_), .A2(new_n14950_), .B(\asqrt[50] ), .ZN(new_n14951_));
  AOI21_X1   g14759(.A1(new_n14938_), .A2(new_n14951_), .B(new_n1305_), .ZN(new_n14952_));
  NOR3_X1    g14760(.A1(new_n14937_), .A2(\asqrt[52] ), .A3(new_n14952_), .ZN(new_n14953_));
  OAI21_X1   g14761(.A1(new_n14937_), .A2(new_n14952_), .B(\asqrt[52] ), .ZN(new_n14954_));
  OAI21_X1   g14762(.A1(new_n14554_), .A2(new_n14953_), .B(new_n14954_), .ZN(new_n14955_));
  OAI21_X1   g14763(.A1(new_n14955_), .A2(\asqrt[53] ), .B(new_n14551_), .ZN(new_n14956_));
  NAND2_X1   g14764(.A1(new_n14955_), .A2(\asqrt[53] ), .ZN(new_n14957_));
  NAND3_X1   g14765(.A1(new_n14956_), .A2(new_n14957_), .A3(new_n860_), .ZN(new_n14958_));
  AOI21_X1   g14766(.A1(new_n14956_), .A2(new_n14957_), .B(new_n860_), .ZN(new_n14959_));
  AOI21_X1   g14767(.A1(new_n14548_), .A2(new_n14958_), .B(new_n14959_), .ZN(new_n14960_));
  NAND2_X1   g14768(.A1(new_n14960_), .A2(new_n744_), .ZN(new_n14961_));
  INV_X1     g14769(.I(new_n14548_), .ZN(new_n14962_));
  INV_X1     g14770(.I(new_n14551_), .ZN(new_n14963_));
  INV_X1     g14771(.I(new_n14560_), .ZN(new_n14964_));
  NOR3_X1    g14772(.A1(new_n14948_), .A2(\asqrt[50] ), .A3(new_n14950_), .ZN(new_n14965_));
  OAI21_X1   g14773(.A1(new_n14964_), .A2(new_n14965_), .B(new_n14951_), .ZN(new_n14966_));
  OAI21_X1   g14774(.A1(new_n14966_), .A2(\asqrt[51] ), .B(new_n14556_), .ZN(new_n14967_));
  NAND2_X1   g14775(.A1(new_n14966_), .A2(\asqrt[51] ), .ZN(new_n14968_));
  NAND3_X1   g14776(.A1(new_n14967_), .A2(new_n14968_), .A3(new_n1150_), .ZN(new_n14969_));
  AOI21_X1   g14777(.A1(new_n14967_), .A2(new_n14968_), .B(new_n1150_), .ZN(new_n14970_));
  AOI21_X1   g14778(.A1(new_n14553_), .A2(new_n14969_), .B(new_n14970_), .ZN(new_n14971_));
  AOI21_X1   g14779(.A1(new_n14971_), .A2(new_n1006_), .B(new_n14963_), .ZN(new_n14972_));
  NAND2_X1   g14780(.A1(new_n14969_), .A2(new_n14553_), .ZN(new_n14973_));
  AOI21_X1   g14781(.A1(new_n14973_), .A2(new_n14954_), .B(new_n1006_), .ZN(new_n14974_));
  NOR3_X1    g14782(.A1(new_n14972_), .A2(\asqrt[54] ), .A3(new_n14974_), .ZN(new_n14975_));
  OAI21_X1   g14783(.A1(new_n14972_), .A2(new_n14974_), .B(\asqrt[54] ), .ZN(new_n14976_));
  OAI21_X1   g14784(.A1(new_n14962_), .A2(new_n14975_), .B(new_n14976_), .ZN(new_n14977_));
  NAND2_X1   g14785(.A1(new_n14977_), .A2(\asqrt[55] ), .ZN(new_n14978_));
  NOR2_X1    g14786(.A1(new_n14500_), .A2(\asqrt[62] ), .ZN(new_n14979_));
  NOR2_X1    g14787(.A1(new_n14979_), .A2(new_n14681_), .ZN(new_n14980_));
  XOR2_X1    g14788(.A1(new_n14524_), .A2(new_n14031_), .Z(new_n14981_));
  OAI21_X1   g14789(.A1(\asqrt[10] ), .A2(new_n14980_), .B(new_n14981_), .ZN(new_n14982_));
  INV_X1     g14790(.I(new_n14982_), .ZN(new_n14983_));
  AOI21_X1   g14791(.A1(new_n14508_), .A2(new_n14513_), .B(\asqrt[10] ), .ZN(new_n14984_));
  XOR2_X1    g14792(.A1(new_n14984_), .A2(new_n14458_), .Z(new_n14985_));
  INV_X1     g14793(.I(new_n14985_), .ZN(new_n14986_));
  AOI21_X1   g14794(.A1(new_n14488_), .A2(new_n14507_), .B(\asqrt[10] ), .ZN(new_n14987_));
  XOR2_X1    g14795(.A1(new_n14987_), .A2(new_n14462_), .Z(new_n14988_));
  INV_X1     g14796(.I(new_n14988_), .ZN(new_n14989_));
  NOR2_X1    g14797(.A1(new_n14506_), .A2(new_n14502_), .ZN(new_n14990_));
  NOR2_X1    g14798(.A1(\asqrt[10] ), .A2(new_n14990_), .ZN(new_n14991_));
  XOR2_X1    g14799(.A1(new_n14991_), .A2(new_n14464_), .Z(new_n14992_));
  NOR2_X1    g14800(.A1(new_n14477_), .A2(new_n14486_), .ZN(new_n14993_));
  NOR2_X1    g14801(.A1(\asqrt[10] ), .A2(new_n14993_), .ZN(new_n14994_));
  XOR2_X1    g14802(.A1(new_n14994_), .A2(new_n14467_), .Z(new_n14995_));
  AOI21_X1   g14803(.A1(new_n14481_), .A2(new_n14485_), .B(\asqrt[10] ), .ZN(new_n14996_));
  XOR2_X1    g14804(.A1(new_n14996_), .A2(new_n14470_), .Z(new_n14997_));
  INV_X1     g14805(.I(new_n14997_), .ZN(new_n14998_));
  INV_X1     g14806(.I(new_n14545_), .ZN(new_n14999_));
  AOI21_X1   g14807(.A1(new_n14960_), .A2(new_n744_), .B(new_n14999_), .ZN(new_n15000_));
  NAND2_X1   g14808(.A1(new_n14958_), .A2(new_n14548_), .ZN(new_n15001_));
  AOI21_X1   g14809(.A1(new_n15001_), .A2(new_n14976_), .B(new_n744_), .ZN(new_n15002_));
  NOR3_X1    g14810(.A1(new_n15000_), .A2(\asqrt[56] ), .A3(new_n15002_), .ZN(new_n15003_));
  OAI21_X1   g14811(.A1(new_n15000_), .A2(new_n15002_), .B(\asqrt[56] ), .ZN(new_n15004_));
  OAI21_X1   g14812(.A1(new_n14998_), .A2(new_n15003_), .B(new_n15004_), .ZN(new_n15005_));
  OAI21_X1   g14813(.A1(new_n15005_), .A2(\asqrt[57] ), .B(new_n14995_), .ZN(new_n15006_));
  NAND2_X1   g14814(.A1(new_n15005_), .A2(\asqrt[57] ), .ZN(new_n15007_));
  NAND3_X1   g14815(.A1(new_n15006_), .A2(new_n15007_), .A3(new_n423_), .ZN(new_n15008_));
  AOI21_X1   g14816(.A1(new_n15006_), .A2(new_n15007_), .B(new_n423_), .ZN(new_n15009_));
  AOI21_X1   g14817(.A1(new_n14992_), .A2(new_n15008_), .B(new_n15009_), .ZN(new_n15010_));
  AOI21_X1   g14818(.A1(new_n15010_), .A2(new_n337_), .B(new_n14989_), .ZN(new_n15011_));
  NAND2_X1   g14819(.A1(new_n15008_), .A2(new_n14992_), .ZN(new_n15012_));
  INV_X1     g14820(.I(new_n14995_), .ZN(new_n15013_));
  OAI21_X1   g14821(.A1(new_n14977_), .A2(\asqrt[55] ), .B(new_n14545_), .ZN(new_n15014_));
  NAND3_X1   g14822(.A1(new_n15014_), .A2(new_n14978_), .A3(new_n634_), .ZN(new_n15015_));
  AOI21_X1   g14823(.A1(new_n15014_), .A2(new_n14978_), .B(new_n634_), .ZN(new_n15016_));
  AOI21_X1   g14824(.A1(new_n14997_), .A2(new_n15015_), .B(new_n15016_), .ZN(new_n15017_));
  AOI21_X1   g14825(.A1(new_n15017_), .A2(new_n531_), .B(new_n15013_), .ZN(new_n15018_));
  NAND2_X1   g14826(.A1(new_n15015_), .A2(new_n14997_), .ZN(new_n15019_));
  AOI21_X1   g14827(.A1(new_n15019_), .A2(new_n15004_), .B(new_n531_), .ZN(new_n15020_));
  OAI21_X1   g14828(.A1(new_n15018_), .A2(new_n15020_), .B(\asqrt[58] ), .ZN(new_n15021_));
  AOI21_X1   g14829(.A1(new_n15012_), .A2(new_n15021_), .B(new_n337_), .ZN(new_n15022_));
  NOR3_X1    g14830(.A1(new_n15011_), .A2(\asqrt[60] ), .A3(new_n15022_), .ZN(new_n15023_));
  NOR2_X1    g14831(.A1(new_n15023_), .A2(new_n14986_), .ZN(new_n15024_));
  INV_X1     g14832(.I(new_n14992_), .ZN(new_n15025_));
  NOR3_X1    g14833(.A1(new_n15018_), .A2(\asqrt[58] ), .A3(new_n15020_), .ZN(new_n15026_));
  OAI21_X1   g14834(.A1(new_n15025_), .A2(new_n15026_), .B(new_n15021_), .ZN(new_n15027_));
  OAI21_X1   g14835(.A1(new_n15027_), .A2(\asqrt[59] ), .B(new_n14988_), .ZN(new_n15028_));
  NOR2_X1    g14836(.A1(new_n15026_), .A2(new_n15025_), .ZN(new_n15029_));
  OAI21_X1   g14837(.A1(new_n15029_), .A2(new_n15009_), .B(\asqrt[59] ), .ZN(new_n15030_));
  AOI21_X1   g14838(.A1(new_n15028_), .A2(new_n15030_), .B(new_n266_), .ZN(new_n15031_));
  OAI21_X1   g14839(.A1(new_n15024_), .A2(new_n15031_), .B(\asqrt[61] ), .ZN(new_n15032_));
  OAI21_X1   g14840(.A1(new_n15011_), .A2(new_n15022_), .B(\asqrt[60] ), .ZN(new_n15033_));
  OAI21_X1   g14841(.A1(new_n14986_), .A2(new_n15023_), .B(new_n15033_), .ZN(new_n15034_));
  AOI21_X1   g14842(.A1(new_n14514_), .A2(new_n14494_), .B(\asqrt[10] ), .ZN(new_n15035_));
  XOR2_X1    g14843(.A1(new_n15035_), .A2(new_n14455_), .Z(new_n15036_));
  OAI21_X1   g14844(.A1(new_n15034_), .A2(\asqrt[61] ), .B(new_n15036_), .ZN(new_n15037_));
  NAND2_X1   g14845(.A1(new_n15037_), .A2(new_n15032_), .ZN(new_n15038_));
  NAND3_X1   g14846(.A1(new_n15028_), .A2(new_n266_), .A3(new_n15030_), .ZN(new_n15039_));
  NAND2_X1   g14847(.A1(new_n15039_), .A2(new_n14985_), .ZN(new_n15040_));
  AOI21_X1   g14848(.A1(new_n15040_), .A2(new_n15033_), .B(new_n239_), .ZN(new_n15041_));
  AOI21_X1   g14849(.A1(new_n14985_), .A2(new_n15039_), .B(new_n15031_), .ZN(new_n15042_));
  INV_X1     g14850(.I(new_n15036_), .ZN(new_n15043_));
  AOI21_X1   g14851(.A1(new_n15042_), .A2(new_n239_), .B(new_n15043_), .ZN(new_n15044_));
  OAI21_X1   g14852(.A1(new_n15044_), .A2(new_n15041_), .B(new_n201_), .ZN(new_n15045_));
  NAND3_X1   g14853(.A1(new_n15037_), .A2(\asqrt[62] ), .A3(new_n15032_), .ZN(new_n15046_));
  NAND2_X1   g14854(.A1(new_n14518_), .A2(new_n239_), .ZN(new_n15047_));
  AOI21_X1   g14855(.A1(new_n14496_), .A2(new_n15047_), .B(\asqrt[10] ), .ZN(new_n15048_));
  XOR2_X1    g14856(.A1(new_n15048_), .A2(new_n14498_), .Z(new_n15049_));
  INV_X1     g14857(.I(new_n15049_), .ZN(new_n15050_));
  AOI22_X1   g14858(.A1(new_n15045_), .A2(new_n15046_), .B1(new_n15038_), .B2(new_n15050_), .ZN(new_n15051_));
  NOR2_X1    g14859(.A1(new_n14527_), .A2(new_n14453_), .ZN(new_n15052_));
  OAI21_X1   g14860(.A1(\asqrt[10] ), .A2(new_n15052_), .B(new_n14534_), .ZN(new_n15053_));
  INV_X1     g14861(.I(new_n15053_), .ZN(new_n15054_));
  OAI21_X1   g14862(.A1(new_n15051_), .A2(new_n14983_), .B(new_n15054_), .ZN(new_n15055_));
  OAI21_X1   g14863(.A1(new_n15038_), .A2(\asqrt[62] ), .B(new_n15049_), .ZN(new_n15056_));
  NAND2_X1   g14864(.A1(new_n15038_), .A2(\asqrt[62] ), .ZN(new_n15057_));
  NAND3_X1   g14865(.A1(new_n15056_), .A2(new_n15057_), .A3(new_n14983_), .ZN(new_n15058_));
  NAND2_X1   g14866(.A1(new_n14690_), .A2(new_n14452_), .ZN(new_n15059_));
  XOR2_X1    g14867(.A1(new_n14678_), .A2(new_n14452_), .Z(new_n15060_));
  NAND3_X1   g14868(.A1(new_n15059_), .A2(\asqrt[63] ), .A3(new_n15060_), .ZN(new_n15061_));
  INV_X1     g14869(.I(new_n14687_), .ZN(new_n15062_));
  NAND4_X1   g14870(.A1(new_n15062_), .A2(new_n14453_), .A3(new_n14534_), .A4(new_n14542_), .ZN(new_n15063_));
  NAND2_X1   g14871(.A1(new_n15061_), .A2(new_n15063_), .ZN(new_n15064_));
  INV_X1     g14872(.I(new_n15064_), .ZN(new_n15065_));
  NAND4_X1   g14873(.A1(new_n15055_), .A2(new_n193_), .A3(new_n15058_), .A4(new_n15065_), .ZN(\asqrt[9] ));
  AOI21_X1   g14874(.A1(new_n14961_), .A2(new_n14978_), .B(\asqrt[9] ), .ZN(new_n15067_));
  XOR2_X1    g14875(.A1(new_n15067_), .A2(new_n14545_), .Z(new_n15068_));
  AOI21_X1   g14876(.A1(new_n14958_), .A2(new_n14976_), .B(\asqrt[9] ), .ZN(new_n15069_));
  XOR2_X1    g14877(.A1(new_n15069_), .A2(new_n14548_), .Z(new_n15070_));
  NAND2_X1   g14878(.A1(new_n14971_), .A2(new_n1006_), .ZN(new_n15071_));
  AOI21_X1   g14879(.A1(new_n15071_), .A2(new_n14957_), .B(\asqrt[9] ), .ZN(new_n15072_));
  XOR2_X1    g14880(.A1(new_n15072_), .A2(new_n14551_), .Z(new_n15073_));
  INV_X1     g14881(.I(new_n15073_), .ZN(new_n15074_));
  AOI21_X1   g14882(.A1(new_n14969_), .A2(new_n14954_), .B(\asqrt[9] ), .ZN(new_n15075_));
  XOR2_X1    g14883(.A1(new_n15075_), .A2(new_n14553_), .Z(new_n15076_));
  INV_X1     g14884(.I(new_n15076_), .ZN(new_n15077_));
  NAND2_X1   g14885(.A1(new_n14936_), .A2(new_n1305_), .ZN(new_n15078_));
  AOI21_X1   g14886(.A1(new_n15078_), .A2(new_n14968_), .B(\asqrt[9] ), .ZN(new_n15079_));
  XOR2_X1    g14887(.A1(new_n15079_), .A2(new_n14556_), .Z(new_n15080_));
  AOI21_X1   g14888(.A1(new_n14934_), .A2(new_n14951_), .B(\asqrt[9] ), .ZN(new_n15081_));
  XOR2_X1    g14889(.A1(new_n15081_), .A2(new_n14560_), .Z(new_n15082_));
  NAND2_X1   g14890(.A1(new_n14947_), .A2(new_n1632_), .ZN(new_n15083_));
  AOI21_X1   g14891(.A1(new_n15083_), .A2(new_n14933_), .B(\asqrt[9] ), .ZN(new_n15084_));
  XOR2_X1    g14892(.A1(new_n15084_), .A2(new_n14563_), .Z(new_n15085_));
  INV_X1     g14893(.I(new_n15085_), .ZN(new_n15086_));
  AOI21_X1   g14894(.A1(new_n14945_), .A2(new_n14930_), .B(\asqrt[9] ), .ZN(new_n15087_));
  XOR2_X1    g14895(.A1(new_n15087_), .A2(new_n14565_), .Z(new_n15088_));
  INV_X1     g14896(.I(new_n15088_), .ZN(new_n15089_));
  NAND2_X1   g14897(.A1(new_n14912_), .A2(new_n1953_), .ZN(new_n15090_));
  AOI21_X1   g14898(.A1(new_n15090_), .A2(new_n14944_), .B(\asqrt[9] ), .ZN(new_n15091_));
  XOR2_X1    g14899(.A1(new_n15091_), .A2(new_n14568_), .Z(new_n15092_));
  AOI21_X1   g14900(.A1(new_n14910_), .A2(new_n14927_), .B(\asqrt[9] ), .ZN(new_n15093_));
  XOR2_X1    g14901(.A1(new_n15093_), .A2(new_n14572_), .Z(new_n15094_));
  NAND2_X1   g14902(.A1(new_n14923_), .A2(new_n2332_), .ZN(new_n15095_));
  AOI21_X1   g14903(.A1(new_n15095_), .A2(new_n14909_), .B(\asqrt[9] ), .ZN(new_n15096_));
  XOR2_X1    g14904(.A1(new_n15096_), .A2(new_n14575_), .Z(new_n15097_));
  INV_X1     g14905(.I(new_n15097_), .ZN(new_n15098_));
  AOI21_X1   g14906(.A1(new_n14921_), .A2(new_n14906_), .B(\asqrt[9] ), .ZN(new_n15099_));
  XOR2_X1    g14907(.A1(new_n15099_), .A2(new_n14577_), .Z(new_n15100_));
  INV_X1     g14908(.I(new_n15100_), .ZN(new_n15101_));
  NAND2_X1   g14909(.A1(new_n14888_), .A2(new_n2749_), .ZN(new_n15102_));
  AOI21_X1   g14910(.A1(new_n15102_), .A2(new_n14920_), .B(\asqrt[9] ), .ZN(new_n15103_));
  XOR2_X1    g14911(.A1(new_n15103_), .A2(new_n14580_), .Z(new_n15104_));
  AOI21_X1   g14912(.A1(new_n14886_), .A2(new_n14903_), .B(\asqrt[9] ), .ZN(new_n15105_));
  XOR2_X1    g14913(.A1(new_n15105_), .A2(new_n14584_), .Z(new_n15106_));
  NAND2_X1   g14914(.A1(new_n14899_), .A2(new_n3195_), .ZN(new_n15107_));
  AOI21_X1   g14915(.A1(new_n15107_), .A2(new_n14885_), .B(\asqrt[9] ), .ZN(new_n15108_));
  XOR2_X1    g14916(.A1(new_n15108_), .A2(new_n14587_), .Z(new_n15109_));
  INV_X1     g14917(.I(new_n15109_), .ZN(new_n15110_));
  AOI21_X1   g14918(.A1(new_n14897_), .A2(new_n14882_), .B(\asqrt[9] ), .ZN(new_n15111_));
  XOR2_X1    g14919(.A1(new_n15111_), .A2(new_n14589_), .Z(new_n15112_));
  INV_X1     g14920(.I(new_n15112_), .ZN(new_n15113_));
  NAND2_X1   g14921(.A1(new_n14864_), .A2(new_n3681_), .ZN(new_n15114_));
  AOI21_X1   g14922(.A1(new_n15114_), .A2(new_n14896_), .B(\asqrt[9] ), .ZN(new_n15115_));
  XOR2_X1    g14923(.A1(new_n15115_), .A2(new_n14592_), .Z(new_n15116_));
  AOI21_X1   g14924(.A1(new_n14862_), .A2(new_n14879_), .B(\asqrt[9] ), .ZN(new_n15117_));
  XOR2_X1    g14925(.A1(new_n15117_), .A2(new_n14596_), .Z(new_n15118_));
  NAND2_X1   g14926(.A1(new_n14875_), .A2(new_n4196_), .ZN(new_n15119_));
  AOI21_X1   g14927(.A1(new_n15119_), .A2(new_n14861_), .B(\asqrt[9] ), .ZN(new_n15120_));
  XOR2_X1    g14928(.A1(new_n15120_), .A2(new_n14599_), .Z(new_n15121_));
  INV_X1     g14929(.I(new_n15121_), .ZN(new_n15122_));
  AOI21_X1   g14930(.A1(new_n14873_), .A2(new_n14858_), .B(\asqrt[9] ), .ZN(new_n15123_));
  XOR2_X1    g14931(.A1(new_n15123_), .A2(new_n14601_), .Z(new_n15124_));
  INV_X1     g14932(.I(new_n15124_), .ZN(new_n15125_));
  NAND2_X1   g14933(.A1(new_n14840_), .A2(new_n4751_), .ZN(new_n15126_));
  AOI21_X1   g14934(.A1(new_n15126_), .A2(new_n14872_), .B(\asqrt[9] ), .ZN(new_n15127_));
  XOR2_X1    g14935(.A1(new_n15127_), .A2(new_n14604_), .Z(new_n15128_));
  AOI21_X1   g14936(.A1(new_n14838_), .A2(new_n14855_), .B(\asqrt[9] ), .ZN(new_n15129_));
  XOR2_X1    g14937(.A1(new_n15129_), .A2(new_n14608_), .Z(new_n15130_));
  NAND2_X1   g14938(.A1(new_n14851_), .A2(new_n5336_), .ZN(new_n15131_));
  AOI21_X1   g14939(.A1(new_n15131_), .A2(new_n14837_), .B(\asqrt[9] ), .ZN(new_n15132_));
  XOR2_X1    g14940(.A1(new_n15132_), .A2(new_n14611_), .Z(new_n15133_));
  INV_X1     g14941(.I(new_n15133_), .ZN(new_n15134_));
  AOI21_X1   g14942(.A1(new_n14849_), .A2(new_n14834_), .B(\asqrt[9] ), .ZN(new_n15135_));
  XOR2_X1    g14943(.A1(new_n15135_), .A2(new_n14613_), .Z(new_n15136_));
  INV_X1     g14944(.I(new_n15136_), .ZN(new_n15137_));
  NAND2_X1   g14945(.A1(new_n14816_), .A2(new_n5947_), .ZN(new_n15138_));
  AOI21_X1   g14946(.A1(new_n15138_), .A2(new_n14848_), .B(\asqrt[9] ), .ZN(new_n15139_));
  XOR2_X1    g14947(.A1(new_n15139_), .A2(new_n14616_), .Z(new_n15140_));
  AOI21_X1   g14948(.A1(new_n14814_), .A2(new_n14831_), .B(\asqrt[9] ), .ZN(new_n15141_));
  XOR2_X1    g14949(.A1(new_n15141_), .A2(new_n14620_), .Z(new_n15142_));
  NAND2_X1   g14950(.A1(new_n14827_), .A2(new_n6636_), .ZN(new_n15143_));
  AOI21_X1   g14951(.A1(new_n15143_), .A2(new_n14813_), .B(\asqrt[9] ), .ZN(new_n15144_));
  XOR2_X1    g14952(.A1(new_n15144_), .A2(new_n14623_), .Z(new_n15145_));
  INV_X1     g14953(.I(new_n15145_), .ZN(new_n15146_));
  AOI21_X1   g14954(.A1(new_n14825_), .A2(new_n14810_), .B(\asqrt[9] ), .ZN(new_n15147_));
  XOR2_X1    g14955(.A1(new_n15147_), .A2(new_n14625_), .Z(new_n15148_));
  INV_X1     g14956(.I(new_n15148_), .ZN(new_n15149_));
  NAND2_X1   g14957(.A1(new_n14792_), .A2(new_n7331_), .ZN(new_n15150_));
  AOI21_X1   g14958(.A1(new_n15150_), .A2(new_n14824_), .B(\asqrt[9] ), .ZN(new_n15151_));
  XOR2_X1    g14959(.A1(new_n15151_), .A2(new_n14628_), .Z(new_n15152_));
  AOI21_X1   g14960(.A1(new_n14790_), .A2(new_n14807_), .B(\asqrt[9] ), .ZN(new_n15153_));
  XOR2_X1    g14961(.A1(new_n15153_), .A2(new_n14632_), .Z(new_n15154_));
  NAND2_X1   g14962(.A1(new_n14803_), .A2(new_n8077_), .ZN(new_n15155_));
  AOI21_X1   g14963(.A1(new_n15155_), .A2(new_n14789_), .B(\asqrt[9] ), .ZN(new_n15156_));
  XOR2_X1    g14964(.A1(new_n15156_), .A2(new_n14635_), .Z(new_n15157_));
  INV_X1     g14965(.I(new_n15157_), .ZN(new_n15158_));
  AOI21_X1   g14966(.A1(new_n14801_), .A2(new_n14786_), .B(\asqrt[9] ), .ZN(new_n15159_));
  XOR2_X1    g14967(.A1(new_n15159_), .A2(new_n14637_), .Z(new_n15160_));
  INV_X1     g14968(.I(new_n15160_), .ZN(new_n15161_));
  NAND2_X1   g14969(.A1(new_n14768_), .A2(new_n8849_), .ZN(new_n15162_));
  AOI21_X1   g14970(.A1(new_n15162_), .A2(new_n14800_), .B(\asqrt[9] ), .ZN(new_n15163_));
  XOR2_X1    g14971(.A1(new_n15163_), .A2(new_n14640_), .Z(new_n15164_));
  AOI21_X1   g14972(.A1(new_n14766_), .A2(new_n14783_), .B(\asqrt[9] ), .ZN(new_n15165_));
  XOR2_X1    g14973(.A1(new_n15165_), .A2(new_n14644_), .Z(new_n15166_));
  NAND2_X1   g14974(.A1(new_n14779_), .A2(new_n9656_), .ZN(new_n15167_));
  AOI21_X1   g14975(.A1(new_n15167_), .A2(new_n14765_), .B(\asqrt[9] ), .ZN(new_n15168_));
  XOR2_X1    g14976(.A1(new_n15168_), .A2(new_n14647_), .Z(new_n15169_));
  INV_X1     g14977(.I(new_n15169_), .ZN(new_n15170_));
  AOI21_X1   g14978(.A1(new_n14777_), .A2(new_n14762_), .B(\asqrt[9] ), .ZN(new_n15171_));
  XOR2_X1    g14979(.A1(new_n15171_), .A2(new_n14649_), .Z(new_n15172_));
  INV_X1     g14980(.I(new_n15172_), .ZN(new_n15173_));
  NAND2_X1   g14981(.A1(new_n14744_), .A2(new_n10497_), .ZN(new_n15174_));
  AOI21_X1   g14982(.A1(new_n15174_), .A2(new_n14776_), .B(\asqrt[9] ), .ZN(new_n15175_));
  XOR2_X1    g14983(.A1(new_n15175_), .A2(new_n14652_), .Z(new_n15176_));
  AOI21_X1   g14984(.A1(new_n14742_), .A2(new_n14759_), .B(\asqrt[9] ), .ZN(new_n15177_));
  XOR2_X1    g14985(.A1(new_n15177_), .A2(new_n14656_), .Z(new_n15178_));
  NAND2_X1   g14986(.A1(new_n14755_), .A2(new_n11373_), .ZN(new_n15179_));
  AOI21_X1   g14987(.A1(new_n15179_), .A2(new_n14741_), .B(\asqrt[9] ), .ZN(new_n15180_));
  XOR2_X1    g14988(.A1(new_n15180_), .A2(new_n14659_), .Z(new_n15181_));
  INV_X1     g14989(.I(new_n15181_), .ZN(new_n15182_));
  AOI21_X1   g14990(.A1(new_n14753_), .A2(new_n14738_), .B(\asqrt[9] ), .ZN(new_n15183_));
  XOR2_X1    g14991(.A1(new_n15183_), .A2(new_n14661_), .Z(new_n15184_));
  INV_X1     g14992(.I(new_n15184_), .ZN(new_n15185_));
  NAND2_X1   g14993(.A1(new_n14716_), .A2(new_n12283_), .ZN(new_n15186_));
  AOI21_X1   g14994(.A1(new_n15186_), .A2(new_n14752_), .B(\asqrt[9] ), .ZN(new_n15187_));
  XOR2_X1    g14995(.A1(new_n15187_), .A2(new_n14664_), .Z(new_n15188_));
  AOI21_X1   g14996(.A1(new_n14714_), .A2(new_n14735_), .B(\asqrt[9] ), .ZN(new_n15189_));
  XOR2_X1    g14997(.A1(new_n15189_), .A2(new_n14667_), .Z(new_n15190_));
  NAND2_X1   g14998(.A1(new_n14731_), .A2(new_n13228_), .ZN(new_n15191_));
  AOI21_X1   g14999(.A1(new_n15191_), .A2(new_n14713_), .B(\asqrt[9] ), .ZN(new_n15192_));
  XOR2_X1    g15000(.A1(new_n15192_), .A2(new_n14674_), .Z(new_n15193_));
  INV_X1     g15001(.I(new_n15193_), .ZN(new_n15194_));
  AOI21_X1   g15002(.A1(new_n14729_), .A2(new_n14710_), .B(\asqrt[9] ), .ZN(new_n15195_));
  XOR2_X1    g15003(.A1(new_n15195_), .A2(new_n14720_), .Z(new_n15196_));
  INV_X1     g15004(.I(new_n15196_), .ZN(new_n15197_));
  NAND2_X1   g15005(.A1(\asqrt[10] ), .A2(new_n14697_), .ZN(new_n15198_));
  NOR2_X1    g15006(.A1(new_n14705_), .A2(\a[20] ), .ZN(new_n15199_));
  AOI22_X1   g15007(.A1(new_n15198_), .A2(new_n14705_), .B1(\asqrt[10] ), .B2(new_n15199_), .ZN(new_n15200_));
  OAI21_X1   g15008(.A1(new_n14690_), .A2(new_n14697_), .B(new_n14724_), .ZN(new_n15201_));
  AOI21_X1   g15009(.A1(new_n14723_), .A2(new_n15201_), .B(\asqrt[9] ), .ZN(new_n15202_));
  XOR2_X1    g15010(.A1(new_n15202_), .A2(new_n15200_), .Z(new_n15203_));
  NAND3_X1   g15011(.A1(new_n15040_), .A2(new_n239_), .A3(new_n15033_), .ZN(new_n15204_));
  AOI21_X1   g15012(.A1(new_n15036_), .A2(new_n15204_), .B(new_n15041_), .ZN(new_n15205_));
  AOI21_X1   g15013(.A1(new_n15037_), .A2(new_n15032_), .B(\asqrt[62] ), .ZN(new_n15206_));
  NOR3_X1    g15014(.A1(new_n15044_), .A2(new_n201_), .A3(new_n15041_), .ZN(new_n15207_));
  OAI22_X1   g15015(.A1(new_n15207_), .A2(new_n15206_), .B1(new_n15205_), .B2(new_n15049_), .ZN(new_n15208_));
  AOI21_X1   g15016(.A1(new_n15208_), .A2(new_n14982_), .B(new_n15053_), .ZN(new_n15209_));
  AOI21_X1   g15017(.A1(new_n15205_), .A2(new_n201_), .B(new_n15050_), .ZN(new_n15210_));
  OAI21_X1   g15018(.A1(new_n15205_), .A2(new_n201_), .B(new_n14983_), .ZN(new_n15211_));
  NOR2_X1    g15019(.A1(new_n15210_), .A2(new_n15211_), .ZN(new_n15212_));
  NOR3_X1    g15020(.A1(new_n15209_), .A2(\asqrt[63] ), .A3(new_n15212_), .ZN(new_n15213_));
  NAND3_X1   g15021(.A1(new_n15061_), .A2(\asqrt[10] ), .A3(new_n15063_), .ZN(new_n15214_));
  INV_X1     g15022(.I(new_n15214_), .ZN(new_n15215_));
  NAND2_X1   g15023(.A1(new_n15213_), .A2(new_n15215_), .ZN(new_n15216_));
  NAND2_X1   g15024(.A1(\asqrt[9] ), .A2(new_n14694_), .ZN(new_n15217_));
  AOI21_X1   g15025(.A1(new_n15217_), .A2(new_n15216_), .B(\a[20] ), .ZN(new_n15218_));
  NAND2_X1   g15026(.A1(new_n15055_), .A2(new_n193_), .ZN(new_n15219_));
  NOR3_X1    g15027(.A1(new_n15219_), .A2(new_n15212_), .A3(new_n15214_), .ZN(new_n15220_));
  NOR4_X1    g15028(.A1(new_n15209_), .A2(\asqrt[63] ), .A3(new_n15212_), .A4(new_n15064_), .ZN(new_n15221_));
  NOR2_X1    g15029(.A1(new_n15221_), .A2(new_n14695_), .ZN(new_n15222_));
  NOR3_X1    g15030(.A1(new_n15222_), .A2(new_n15220_), .A3(new_n14697_), .ZN(new_n15223_));
  NOR2_X1    g15031(.A1(new_n15223_), .A2(new_n15218_), .ZN(new_n15224_));
  INV_X1     g15032(.I(\a[18] ), .ZN(new_n15225_));
  NOR2_X1    g15033(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n15226_));
  NOR3_X1    g15034(.A1(new_n15221_), .A2(new_n15225_), .A3(new_n15226_), .ZN(new_n15227_));
  INV_X1     g15035(.I(new_n15226_), .ZN(new_n15228_));
  AOI21_X1   g15036(.A1(new_n15221_), .A2(\a[18] ), .B(new_n15228_), .ZN(new_n15229_));
  OAI21_X1   g15037(.A1(new_n15227_), .A2(new_n15229_), .B(\asqrt[10] ), .ZN(new_n15230_));
  NAND2_X1   g15038(.A1(new_n15226_), .A2(new_n15225_), .ZN(new_n15231_));
  NAND3_X1   g15039(.A1(new_n14538_), .A2(new_n14540_), .A3(new_n15231_), .ZN(new_n15232_));
  NAND2_X1   g15040(.A1(new_n14683_), .A2(new_n15232_), .ZN(new_n15233_));
  INV_X1     g15041(.I(new_n15233_), .ZN(new_n15234_));
  NOR3_X1    g15042(.A1(new_n15221_), .A2(new_n15225_), .A3(new_n15234_), .ZN(new_n15235_));
  NOR3_X1    g15043(.A1(new_n15221_), .A2(\a[18] ), .A3(\a[19] ), .ZN(new_n15236_));
  INV_X1     g15044(.I(\a[19] ), .ZN(new_n15237_));
  AOI21_X1   g15045(.A1(\asqrt[9] ), .A2(new_n15225_), .B(new_n15237_), .ZN(new_n15238_));
  NOR3_X1    g15046(.A1(new_n15235_), .A2(new_n15236_), .A3(new_n15238_), .ZN(new_n15239_));
  NAND3_X1   g15047(.A1(new_n15239_), .A2(new_n15230_), .A3(new_n14207_), .ZN(new_n15240_));
  NAND2_X1   g15048(.A1(new_n15240_), .A2(new_n15224_), .ZN(new_n15241_));
  NAND3_X1   g15049(.A1(\asqrt[9] ), .A2(\a[18] ), .A3(new_n15228_), .ZN(new_n15242_));
  OAI21_X1   g15050(.A1(\asqrt[9] ), .A2(new_n15225_), .B(new_n15226_), .ZN(new_n15243_));
  AOI21_X1   g15051(.A1(new_n15243_), .A2(new_n15242_), .B(new_n14690_), .ZN(new_n15244_));
  NAND3_X1   g15052(.A1(\asqrt[9] ), .A2(\a[18] ), .A3(new_n15233_), .ZN(new_n15245_));
  NAND3_X1   g15053(.A1(\asqrt[9] ), .A2(new_n15225_), .A3(new_n15237_), .ZN(new_n15246_));
  OAI21_X1   g15054(.A1(new_n15221_), .A2(\a[18] ), .B(\a[19] ), .ZN(new_n15247_));
  NAND3_X1   g15055(.A1(new_n15245_), .A2(new_n15247_), .A3(new_n15246_), .ZN(new_n15248_));
  OAI21_X1   g15056(.A1(new_n15248_), .A2(new_n15244_), .B(\asqrt[11] ), .ZN(new_n15249_));
  NAND3_X1   g15057(.A1(new_n15241_), .A2(new_n13690_), .A3(new_n15249_), .ZN(new_n15250_));
  AOI21_X1   g15058(.A1(new_n15241_), .A2(new_n15249_), .B(new_n13690_), .ZN(new_n15251_));
  AOI21_X1   g15059(.A1(new_n15203_), .A2(new_n15250_), .B(new_n15251_), .ZN(new_n15252_));
  AOI21_X1   g15060(.A1(new_n15252_), .A2(new_n13228_), .B(new_n15197_), .ZN(new_n15253_));
  OR2_X2     g15061(.A1(new_n15223_), .A2(new_n15218_), .Z(new_n15254_));
  NOR3_X1    g15062(.A1(new_n15248_), .A2(new_n15244_), .A3(\asqrt[11] ), .ZN(new_n15255_));
  OAI21_X1   g15063(.A1(new_n15254_), .A2(new_n15255_), .B(new_n15249_), .ZN(new_n15256_));
  OAI21_X1   g15064(.A1(new_n15256_), .A2(\asqrt[12] ), .B(new_n15203_), .ZN(new_n15257_));
  NAND2_X1   g15065(.A1(new_n15256_), .A2(\asqrt[12] ), .ZN(new_n15258_));
  AOI21_X1   g15066(.A1(new_n15257_), .A2(new_n15258_), .B(new_n13228_), .ZN(new_n15259_));
  NOR3_X1    g15067(.A1(new_n15253_), .A2(\asqrt[14] ), .A3(new_n15259_), .ZN(new_n15260_));
  OAI21_X1   g15068(.A1(new_n15253_), .A2(new_n15259_), .B(\asqrt[14] ), .ZN(new_n15261_));
  OAI21_X1   g15069(.A1(new_n15194_), .A2(new_n15260_), .B(new_n15261_), .ZN(new_n15262_));
  OAI21_X1   g15070(.A1(new_n15262_), .A2(\asqrt[15] ), .B(new_n15190_), .ZN(new_n15263_));
  NAND3_X1   g15071(.A1(new_n15257_), .A2(new_n15258_), .A3(new_n13228_), .ZN(new_n15264_));
  AOI21_X1   g15072(.A1(new_n15196_), .A2(new_n15264_), .B(new_n15259_), .ZN(new_n15265_));
  AOI21_X1   g15073(.A1(new_n15265_), .A2(new_n12733_), .B(new_n15194_), .ZN(new_n15266_));
  NAND2_X1   g15074(.A1(new_n15264_), .A2(new_n15196_), .ZN(new_n15267_));
  INV_X1     g15075(.I(new_n15259_), .ZN(new_n15268_));
  AOI21_X1   g15076(.A1(new_n15267_), .A2(new_n15268_), .B(new_n12733_), .ZN(new_n15269_));
  OAI21_X1   g15077(.A1(new_n15266_), .A2(new_n15269_), .B(\asqrt[15] ), .ZN(new_n15270_));
  NAND3_X1   g15078(.A1(new_n15263_), .A2(new_n11802_), .A3(new_n15270_), .ZN(new_n15271_));
  AOI21_X1   g15079(.A1(new_n15263_), .A2(new_n15270_), .B(new_n11802_), .ZN(new_n15272_));
  AOI21_X1   g15080(.A1(new_n15188_), .A2(new_n15271_), .B(new_n15272_), .ZN(new_n15273_));
  AOI21_X1   g15081(.A1(new_n15273_), .A2(new_n11373_), .B(new_n15185_), .ZN(new_n15274_));
  INV_X1     g15082(.I(new_n15190_), .ZN(new_n15275_));
  NOR3_X1    g15083(.A1(new_n15266_), .A2(\asqrt[15] ), .A3(new_n15269_), .ZN(new_n15276_));
  OAI21_X1   g15084(.A1(new_n15275_), .A2(new_n15276_), .B(new_n15270_), .ZN(new_n15277_));
  OAI21_X1   g15085(.A1(new_n15277_), .A2(\asqrt[16] ), .B(new_n15188_), .ZN(new_n15278_));
  NAND2_X1   g15086(.A1(new_n15277_), .A2(\asqrt[16] ), .ZN(new_n15279_));
  AOI21_X1   g15087(.A1(new_n15278_), .A2(new_n15279_), .B(new_n11373_), .ZN(new_n15280_));
  NOR3_X1    g15088(.A1(new_n15274_), .A2(\asqrt[18] ), .A3(new_n15280_), .ZN(new_n15281_));
  OAI21_X1   g15089(.A1(new_n15274_), .A2(new_n15280_), .B(\asqrt[18] ), .ZN(new_n15282_));
  OAI21_X1   g15090(.A1(new_n15182_), .A2(new_n15281_), .B(new_n15282_), .ZN(new_n15283_));
  OAI21_X1   g15091(.A1(new_n15283_), .A2(\asqrt[19] ), .B(new_n15178_), .ZN(new_n15284_));
  NAND3_X1   g15092(.A1(new_n15278_), .A2(new_n15279_), .A3(new_n11373_), .ZN(new_n15285_));
  AOI21_X1   g15093(.A1(new_n15184_), .A2(new_n15285_), .B(new_n15280_), .ZN(new_n15286_));
  AOI21_X1   g15094(.A1(new_n15286_), .A2(new_n10914_), .B(new_n15182_), .ZN(new_n15287_));
  NAND2_X1   g15095(.A1(new_n15285_), .A2(new_n15184_), .ZN(new_n15288_));
  INV_X1     g15096(.I(new_n15280_), .ZN(new_n15289_));
  AOI21_X1   g15097(.A1(new_n15288_), .A2(new_n15289_), .B(new_n10914_), .ZN(new_n15290_));
  OAI21_X1   g15098(.A1(new_n15287_), .A2(new_n15290_), .B(\asqrt[19] ), .ZN(new_n15291_));
  NAND3_X1   g15099(.A1(new_n15284_), .A2(new_n10052_), .A3(new_n15291_), .ZN(new_n15292_));
  AOI21_X1   g15100(.A1(new_n15284_), .A2(new_n15291_), .B(new_n10052_), .ZN(new_n15293_));
  AOI21_X1   g15101(.A1(new_n15176_), .A2(new_n15292_), .B(new_n15293_), .ZN(new_n15294_));
  AOI21_X1   g15102(.A1(new_n15294_), .A2(new_n9656_), .B(new_n15173_), .ZN(new_n15295_));
  INV_X1     g15103(.I(new_n15178_), .ZN(new_n15296_));
  NOR3_X1    g15104(.A1(new_n15287_), .A2(\asqrt[19] ), .A3(new_n15290_), .ZN(new_n15297_));
  OAI21_X1   g15105(.A1(new_n15296_), .A2(new_n15297_), .B(new_n15291_), .ZN(new_n15298_));
  OAI21_X1   g15106(.A1(new_n15298_), .A2(\asqrt[20] ), .B(new_n15176_), .ZN(new_n15299_));
  NAND2_X1   g15107(.A1(new_n15298_), .A2(\asqrt[20] ), .ZN(new_n15300_));
  AOI21_X1   g15108(.A1(new_n15299_), .A2(new_n15300_), .B(new_n9656_), .ZN(new_n15301_));
  NOR3_X1    g15109(.A1(new_n15295_), .A2(\asqrt[22] ), .A3(new_n15301_), .ZN(new_n15302_));
  OAI21_X1   g15110(.A1(new_n15295_), .A2(new_n15301_), .B(\asqrt[22] ), .ZN(new_n15303_));
  OAI21_X1   g15111(.A1(new_n15170_), .A2(new_n15302_), .B(new_n15303_), .ZN(new_n15304_));
  OAI21_X1   g15112(.A1(new_n15304_), .A2(\asqrt[23] ), .B(new_n15166_), .ZN(new_n15305_));
  NAND3_X1   g15113(.A1(new_n15299_), .A2(new_n15300_), .A3(new_n9656_), .ZN(new_n15306_));
  AOI21_X1   g15114(.A1(new_n15172_), .A2(new_n15306_), .B(new_n15301_), .ZN(new_n15307_));
  AOI21_X1   g15115(.A1(new_n15307_), .A2(new_n9233_), .B(new_n15170_), .ZN(new_n15308_));
  NAND2_X1   g15116(.A1(new_n15306_), .A2(new_n15172_), .ZN(new_n15309_));
  INV_X1     g15117(.I(new_n15301_), .ZN(new_n15310_));
  AOI21_X1   g15118(.A1(new_n15309_), .A2(new_n15310_), .B(new_n9233_), .ZN(new_n15311_));
  OAI21_X1   g15119(.A1(new_n15308_), .A2(new_n15311_), .B(\asqrt[23] ), .ZN(new_n15312_));
  NAND3_X1   g15120(.A1(new_n15305_), .A2(new_n8440_), .A3(new_n15312_), .ZN(new_n15313_));
  AOI21_X1   g15121(.A1(new_n15305_), .A2(new_n15312_), .B(new_n8440_), .ZN(new_n15314_));
  AOI21_X1   g15122(.A1(new_n15164_), .A2(new_n15313_), .B(new_n15314_), .ZN(new_n15315_));
  AOI21_X1   g15123(.A1(new_n15315_), .A2(new_n8077_), .B(new_n15161_), .ZN(new_n15316_));
  INV_X1     g15124(.I(new_n15166_), .ZN(new_n15317_));
  NOR3_X1    g15125(.A1(new_n15308_), .A2(\asqrt[23] ), .A3(new_n15311_), .ZN(new_n15318_));
  OAI21_X1   g15126(.A1(new_n15317_), .A2(new_n15318_), .B(new_n15312_), .ZN(new_n15319_));
  OAI21_X1   g15127(.A1(new_n15319_), .A2(\asqrt[24] ), .B(new_n15164_), .ZN(new_n15320_));
  NAND2_X1   g15128(.A1(new_n15319_), .A2(\asqrt[24] ), .ZN(new_n15321_));
  AOI21_X1   g15129(.A1(new_n15320_), .A2(new_n15321_), .B(new_n8077_), .ZN(new_n15322_));
  NOR3_X1    g15130(.A1(new_n15316_), .A2(\asqrt[26] ), .A3(new_n15322_), .ZN(new_n15323_));
  OAI21_X1   g15131(.A1(new_n15316_), .A2(new_n15322_), .B(\asqrt[26] ), .ZN(new_n15324_));
  OAI21_X1   g15132(.A1(new_n15158_), .A2(new_n15323_), .B(new_n15324_), .ZN(new_n15325_));
  OAI21_X1   g15133(.A1(new_n15325_), .A2(\asqrt[27] ), .B(new_n15154_), .ZN(new_n15326_));
  NAND3_X1   g15134(.A1(new_n15320_), .A2(new_n15321_), .A3(new_n8077_), .ZN(new_n15327_));
  AOI21_X1   g15135(.A1(new_n15160_), .A2(new_n15327_), .B(new_n15322_), .ZN(new_n15328_));
  AOI21_X1   g15136(.A1(new_n15328_), .A2(new_n7690_), .B(new_n15158_), .ZN(new_n15329_));
  NAND2_X1   g15137(.A1(new_n15327_), .A2(new_n15160_), .ZN(new_n15330_));
  INV_X1     g15138(.I(new_n15322_), .ZN(new_n15331_));
  AOI21_X1   g15139(.A1(new_n15330_), .A2(new_n15331_), .B(new_n7690_), .ZN(new_n15332_));
  OAI21_X1   g15140(.A1(new_n15329_), .A2(new_n15332_), .B(\asqrt[27] ), .ZN(new_n15333_));
  NAND3_X1   g15141(.A1(new_n15326_), .A2(new_n6966_), .A3(new_n15333_), .ZN(new_n15334_));
  AOI21_X1   g15142(.A1(new_n15326_), .A2(new_n15333_), .B(new_n6966_), .ZN(new_n15335_));
  AOI21_X1   g15143(.A1(new_n15152_), .A2(new_n15334_), .B(new_n15335_), .ZN(new_n15336_));
  AOI21_X1   g15144(.A1(new_n15336_), .A2(new_n6636_), .B(new_n15149_), .ZN(new_n15337_));
  INV_X1     g15145(.I(new_n15154_), .ZN(new_n15338_));
  NOR3_X1    g15146(.A1(new_n15329_), .A2(\asqrt[27] ), .A3(new_n15332_), .ZN(new_n15339_));
  OAI21_X1   g15147(.A1(new_n15338_), .A2(new_n15339_), .B(new_n15333_), .ZN(new_n15340_));
  OAI21_X1   g15148(.A1(new_n15340_), .A2(\asqrt[28] ), .B(new_n15152_), .ZN(new_n15341_));
  NAND2_X1   g15149(.A1(new_n15340_), .A2(\asqrt[28] ), .ZN(new_n15342_));
  AOI21_X1   g15150(.A1(new_n15341_), .A2(new_n15342_), .B(new_n6636_), .ZN(new_n15343_));
  NOR3_X1    g15151(.A1(new_n15337_), .A2(\asqrt[30] ), .A3(new_n15343_), .ZN(new_n15344_));
  OAI21_X1   g15152(.A1(new_n15337_), .A2(new_n15343_), .B(\asqrt[30] ), .ZN(new_n15345_));
  OAI21_X1   g15153(.A1(new_n15146_), .A2(new_n15344_), .B(new_n15345_), .ZN(new_n15346_));
  OAI21_X1   g15154(.A1(new_n15346_), .A2(\asqrt[31] ), .B(new_n15142_), .ZN(new_n15347_));
  NAND3_X1   g15155(.A1(new_n15341_), .A2(new_n15342_), .A3(new_n6636_), .ZN(new_n15348_));
  AOI21_X1   g15156(.A1(new_n15148_), .A2(new_n15348_), .B(new_n15343_), .ZN(new_n15349_));
  AOI21_X1   g15157(.A1(new_n15349_), .A2(new_n6275_), .B(new_n15146_), .ZN(new_n15350_));
  NAND2_X1   g15158(.A1(new_n15348_), .A2(new_n15148_), .ZN(new_n15351_));
  INV_X1     g15159(.I(new_n15343_), .ZN(new_n15352_));
  AOI21_X1   g15160(.A1(new_n15351_), .A2(new_n15352_), .B(new_n6275_), .ZN(new_n15353_));
  OAI21_X1   g15161(.A1(new_n15350_), .A2(new_n15353_), .B(\asqrt[31] ), .ZN(new_n15354_));
  NAND3_X1   g15162(.A1(new_n15347_), .A2(new_n5643_), .A3(new_n15354_), .ZN(new_n15355_));
  AOI21_X1   g15163(.A1(new_n15347_), .A2(new_n15354_), .B(new_n5643_), .ZN(new_n15356_));
  AOI21_X1   g15164(.A1(new_n15140_), .A2(new_n15355_), .B(new_n15356_), .ZN(new_n15357_));
  AOI21_X1   g15165(.A1(new_n15357_), .A2(new_n5336_), .B(new_n15137_), .ZN(new_n15358_));
  INV_X1     g15166(.I(new_n15142_), .ZN(new_n15359_));
  NOR3_X1    g15167(.A1(new_n15350_), .A2(\asqrt[31] ), .A3(new_n15353_), .ZN(new_n15360_));
  OAI21_X1   g15168(.A1(new_n15359_), .A2(new_n15360_), .B(new_n15354_), .ZN(new_n15361_));
  OAI21_X1   g15169(.A1(new_n15361_), .A2(\asqrt[32] ), .B(new_n15140_), .ZN(new_n15362_));
  NAND2_X1   g15170(.A1(new_n15361_), .A2(\asqrt[32] ), .ZN(new_n15363_));
  AOI21_X1   g15171(.A1(new_n15362_), .A2(new_n15363_), .B(new_n5336_), .ZN(new_n15364_));
  NOR3_X1    g15172(.A1(new_n15358_), .A2(\asqrt[34] ), .A3(new_n15364_), .ZN(new_n15365_));
  OAI21_X1   g15173(.A1(new_n15358_), .A2(new_n15364_), .B(\asqrt[34] ), .ZN(new_n15366_));
  OAI21_X1   g15174(.A1(new_n15134_), .A2(new_n15365_), .B(new_n15366_), .ZN(new_n15367_));
  OAI21_X1   g15175(.A1(new_n15367_), .A2(\asqrt[35] ), .B(new_n15130_), .ZN(new_n15368_));
  NAND3_X1   g15176(.A1(new_n15362_), .A2(new_n15363_), .A3(new_n5336_), .ZN(new_n15369_));
  AOI21_X1   g15177(.A1(new_n15136_), .A2(new_n15369_), .B(new_n15364_), .ZN(new_n15370_));
  AOI21_X1   g15178(.A1(new_n15370_), .A2(new_n5029_), .B(new_n15134_), .ZN(new_n15371_));
  NAND2_X1   g15179(.A1(new_n15369_), .A2(new_n15136_), .ZN(new_n15372_));
  INV_X1     g15180(.I(new_n15364_), .ZN(new_n15373_));
  AOI21_X1   g15181(.A1(new_n15372_), .A2(new_n15373_), .B(new_n5029_), .ZN(new_n15374_));
  OAI21_X1   g15182(.A1(new_n15371_), .A2(new_n15374_), .B(\asqrt[35] ), .ZN(new_n15375_));
  NAND3_X1   g15183(.A1(new_n15368_), .A2(new_n4461_), .A3(new_n15375_), .ZN(new_n15376_));
  AOI21_X1   g15184(.A1(new_n15368_), .A2(new_n15375_), .B(new_n4461_), .ZN(new_n15377_));
  AOI21_X1   g15185(.A1(new_n15128_), .A2(new_n15376_), .B(new_n15377_), .ZN(new_n15378_));
  AOI21_X1   g15186(.A1(new_n15378_), .A2(new_n4196_), .B(new_n15125_), .ZN(new_n15379_));
  INV_X1     g15187(.I(new_n15130_), .ZN(new_n15380_));
  NOR3_X1    g15188(.A1(new_n15371_), .A2(\asqrt[35] ), .A3(new_n15374_), .ZN(new_n15381_));
  OAI21_X1   g15189(.A1(new_n15380_), .A2(new_n15381_), .B(new_n15375_), .ZN(new_n15382_));
  OAI21_X1   g15190(.A1(new_n15382_), .A2(\asqrt[36] ), .B(new_n15128_), .ZN(new_n15383_));
  NAND2_X1   g15191(.A1(new_n15382_), .A2(\asqrt[36] ), .ZN(new_n15384_));
  AOI21_X1   g15192(.A1(new_n15383_), .A2(new_n15384_), .B(new_n4196_), .ZN(new_n15385_));
  NOR3_X1    g15193(.A1(new_n15379_), .A2(\asqrt[38] ), .A3(new_n15385_), .ZN(new_n15386_));
  OAI21_X1   g15194(.A1(new_n15379_), .A2(new_n15385_), .B(\asqrt[38] ), .ZN(new_n15387_));
  OAI21_X1   g15195(.A1(new_n15122_), .A2(new_n15386_), .B(new_n15387_), .ZN(new_n15388_));
  OAI21_X1   g15196(.A1(new_n15388_), .A2(\asqrt[39] ), .B(new_n15118_), .ZN(new_n15389_));
  NAND3_X1   g15197(.A1(new_n15383_), .A2(new_n15384_), .A3(new_n4196_), .ZN(new_n15390_));
  AOI21_X1   g15198(.A1(new_n15124_), .A2(new_n15390_), .B(new_n15385_), .ZN(new_n15391_));
  AOI21_X1   g15199(.A1(new_n15391_), .A2(new_n3925_), .B(new_n15122_), .ZN(new_n15392_));
  NAND2_X1   g15200(.A1(new_n15390_), .A2(new_n15124_), .ZN(new_n15393_));
  INV_X1     g15201(.I(new_n15385_), .ZN(new_n15394_));
  AOI21_X1   g15202(.A1(new_n15393_), .A2(new_n15394_), .B(new_n3925_), .ZN(new_n15395_));
  OAI21_X1   g15203(.A1(new_n15392_), .A2(new_n15395_), .B(\asqrt[39] ), .ZN(new_n15396_));
  NAND3_X1   g15204(.A1(new_n15389_), .A2(new_n3427_), .A3(new_n15396_), .ZN(new_n15397_));
  AOI21_X1   g15205(.A1(new_n15389_), .A2(new_n15396_), .B(new_n3427_), .ZN(new_n15398_));
  AOI21_X1   g15206(.A1(new_n15116_), .A2(new_n15397_), .B(new_n15398_), .ZN(new_n15399_));
  AOI21_X1   g15207(.A1(new_n15399_), .A2(new_n3195_), .B(new_n15113_), .ZN(new_n15400_));
  INV_X1     g15208(.I(new_n15118_), .ZN(new_n15401_));
  NOR3_X1    g15209(.A1(new_n15392_), .A2(\asqrt[39] ), .A3(new_n15395_), .ZN(new_n15402_));
  OAI21_X1   g15210(.A1(new_n15401_), .A2(new_n15402_), .B(new_n15396_), .ZN(new_n15403_));
  OAI21_X1   g15211(.A1(new_n15403_), .A2(\asqrt[40] ), .B(new_n15116_), .ZN(new_n15404_));
  NAND2_X1   g15212(.A1(new_n15403_), .A2(\asqrt[40] ), .ZN(new_n15405_));
  AOI21_X1   g15213(.A1(new_n15404_), .A2(new_n15405_), .B(new_n3195_), .ZN(new_n15406_));
  NOR3_X1    g15214(.A1(new_n15400_), .A2(\asqrt[42] ), .A3(new_n15406_), .ZN(new_n15407_));
  OAI21_X1   g15215(.A1(new_n15400_), .A2(new_n15406_), .B(\asqrt[42] ), .ZN(new_n15408_));
  OAI21_X1   g15216(.A1(new_n15110_), .A2(new_n15407_), .B(new_n15408_), .ZN(new_n15409_));
  OAI21_X1   g15217(.A1(new_n15409_), .A2(\asqrt[43] ), .B(new_n15106_), .ZN(new_n15410_));
  NAND3_X1   g15218(.A1(new_n15404_), .A2(new_n15405_), .A3(new_n3195_), .ZN(new_n15411_));
  AOI21_X1   g15219(.A1(new_n15112_), .A2(new_n15411_), .B(new_n15406_), .ZN(new_n15412_));
  AOI21_X1   g15220(.A1(new_n15412_), .A2(new_n2960_), .B(new_n15110_), .ZN(new_n15413_));
  NAND2_X1   g15221(.A1(new_n15411_), .A2(new_n15112_), .ZN(new_n15414_));
  INV_X1     g15222(.I(new_n15406_), .ZN(new_n15415_));
  AOI21_X1   g15223(.A1(new_n15414_), .A2(new_n15415_), .B(new_n2960_), .ZN(new_n15416_));
  OAI21_X1   g15224(.A1(new_n15413_), .A2(new_n15416_), .B(\asqrt[43] ), .ZN(new_n15417_));
  NAND3_X1   g15225(.A1(new_n15410_), .A2(new_n2531_), .A3(new_n15417_), .ZN(new_n15418_));
  AOI21_X1   g15226(.A1(new_n15410_), .A2(new_n15417_), .B(new_n2531_), .ZN(new_n15419_));
  AOI21_X1   g15227(.A1(new_n15104_), .A2(new_n15418_), .B(new_n15419_), .ZN(new_n15420_));
  AOI21_X1   g15228(.A1(new_n15420_), .A2(new_n2332_), .B(new_n15101_), .ZN(new_n15421_));
  INV_X1     g15229(.I(new_n15106_), .ZN(new_n15422_));
  NOR3_X1    g15230(.A1(new_n15413_), .A2(\asqrt[43] ), .A3(new_n15416_), .ZN(new_n15423_));
  OAI21_X1   g15231(.A1(new_n15422_), .A2(new_n15423_), .B(new_n15417_), .ZN(new_n15424_));
  OAI21_X1   g15232(.A1(new_n15424_), .A2(\asqrt[44] ), .B(new_n15104_), .ZN(new_n15425_));
  NAND2_X1   g15233(.A1(new_n15424_), .A2(\asqrt[44] ), .ZN(new_n15426_));
  AOI21_X1   g15234(.A1(new_n15425_), .A2(new_n15426_), .B(new_n2332_), .ZN(new_n15427_));
  NOR3_X1    g15235(.A1(new_n15421_), .A2(\asqrt[46] ), .A3(new_n15427_), .ZN(new_n15428_));
  OAI21_X1   g15236(.A1(new_n15421_), .A2(new_n15427_), .B(\asqrt[46] ), .ZN(new_n15429_));
  OAI21_X1   g15237(.A1(new_n15098_), .A2(new_n15428_), .B(new_n15429_), .ZN(new_n15430_));
  OAI21_X1   g15238(.A1(new_n15430_), .A2(\asqrt[47] ), .B(new_n15094_), .ZN(new_n15431_));
  NAND3_X1   g15239(.A1(new_n15425_), .A2(new_n15426_), .A3(new_n2332_), .ZN(new_n15432_));
  AOI21_X1   g15240(.A1(new_n15100_), .A2(new_n15432_), .B(new_n15427_), .ZN(new_n15433_));
  AOI21_X1   g15241(.A1(new_n15433_), .A2(new_n2134_), .B(new_n15098_), .ZN(new_n15434_));
  NAND2_X1   g15242(.A1(new_n15432_), .A2(new_n15100_), .ZN(new_n15435_));
  INV_X1     g15243(.I(new_n15427_), .ZN(new_n15436_));
  AOI21_X1   g15244(.A1(new_n15435_), .A2(new_n15436_), .B(new_n2134_), .ZN(new_n15437_));
  OAI21_X1   g15245(.A1(new_n15434_), .A2(new_n15437_), .B(\asqrt[47] ), .ZN(new_n15438_));
  NAND3_X1   g15246(.A1(new_n15431_), .A2(new_n1778_), .A3(new_n15438_), .ZN(new_n15439_));
  AOI21_X1   g15247(.A1(new_n15431_), .A2(new_n15438_), .B(new_n1778_), .ZN(new_n15440_));
  AOI21_X1   g15248(.A1(new_n15092_), .A2(new_n15439_), .B(new_n15440_), .ZN(new_n15441_));
  AOI21_X1   g15249(.A1(new_n15441_), .A2(new_n1632_), .B(new_n15089_), .ZN(new_n15442_));
  INV_X1     g15250(.I(new_n15094_), .ZN(new_n15443_));
  NOR3_X1    g15251(.A1(new_n15434_), .A2(\asqrt[47] ), .A3(new_n15437_), .ZN(new_n15444_));
  OAI21_X1   g15252(.A1(new_n15443_), .A2(new_n15444_), .B(new_n15438_), .ZN(new_n15445_));
  OAI21_X1   g15253(.A1(new_n15445_), .A2(\asqrt[48] ), .B(new_n15092_), .ZN(new_n15446_));
  NAND2_X1   g15254(.A1(new_n15445_), .A2(\asqrt[48] ), .ZN(new_n15447_));
  AOI21_X1   g15255(.A1(new_n15446_), .A2(new_n15447_), .B(new_n1632_), .ZN(new_n15448_));
  NOR3_X1    g15256(.A1(new_n15442_), .A2(\asqrt[50] ), .A3(new_n15448_), .ZN(new_n15449_));
  OAI21_X1   g15257(.A1(new_n15442_), .A2(new_n15448_), .B(\asqrt[50] ), .ZN(new_n15450_));
  OAI21_X1   g15258(.A1(new_n15086_), .A2(new_n15449_), .B(new_n15450_), .ZN(new_n15451_));
  OAI21_X1   g15259(.A1(new_n15451_), .A2(\asqrt[51] ), .B(new_n15082_), .ZN(new_n15452_));
  NAND3_X1   g15260(.A1(new_n15446_), .A2(new_n15447_), .A3(new_n1632_), .ZN(new_n15453_));
  AOI21_X1   g15261(.A1(new_n15088_), .A2(new_n15453_), .B(new_n15448_), .ZN(new_n15454_));
  AOI21_X1   g15262(.A1(new_n15454_), .A2(new_n1463_), .B(new_n15086_), .ZN(new_n15455_));
  NAND2_X1   g15263(.A1(new_n15453_), .A2(new_n15088_), .ZN(new_n15456_));
  INV_X1     g15264(.I(new_n15448_), .ZN(new_n15457_));
  AOI21_X1   g15265(.A1(new_n15456_), .A2(new_n15457_), .B(new_n1463_), .ZN(new_n15458_));
  OAI21_X1   g15266(.A1(new_n15455_), .A2(new_n15458_), .B(\asqrt[51] ), .ZN(new_n15459_));
  NAND3_X1   g15267(.A1(new_n15452_), .A2(new_n1150_), .A3(new_n15459_), .ZN(new_n15460_));
  AOI21_X1   g15268(.A1(new_n15452_), .A2(new_n15459_), .B(new_n1150_), .ZN(new_n15461_));
  AOI21_X1   g15269(.A1(new_n15080_), .A2(new_n15460_), .B(new_n15461_), .ZN(new_n15462_));
  AOI21_X1   g15270(.A1(new_n15462_), .A2(new_n1006_), .B(new_n15077_), .ZN(new_n15463_));
  INV_X1     g15271(.I(new_n15082_), .ZN(new_n15464_));
  NOR3_X1    g15272(.A1(new_n15455_), .A2(\asqrt[51] ), .A3(new_n15458_), .ZN(new_n15465_));
  OAI21_X1   g15273(.A1(new_n15464_), .A2(new_n15465_), .B(new_n15459_), .ZN(new_n15466_));
  OAI21_X1   g15274(.A1(new_n15466_), .A2(\asqrt[52] ), .B(new_n15080_), .ZN(new_n15467_));
  NAND2_X1   g15275(.A1(new_n15466_), .A2(\asqrt[52] ), .ZN(new_n15468_));
  AOI21_X1   g15276(.A1(new_n15467_), .A2(new_n15468_), .B(new_n1006_), .ZN(new_n15469_));
  NOR3_X1    g15277(.A1(new_n15463_), .A2(\asqrt[54] ), .A3(new_n15469_), .ZN(new_n15470_));
  OAI21_X1   g15278(.A1(new_n15463_), .A2(new_n15469_), .B(\asqrt[54] ), .ZN(new_n15471_));
  OAI21_X1   g15279(.A1(new_n15074_), .A2(new_n15470_), .B(new_n15471_), .ZN(new_n15472_));
  OAI21_X1   g15280(.A1(new_n15472_), .A2(\asqrt[55] ), .B(new_n15070_), .ZN(new_n15473_));
  NAND3_X1   g15281(.A1(new_n15467_), .A2(new_n15468_), .A3(new_n1006_), .ZN(new_n15474_));
  AOI21_X1   g15282(.A1(new_n15076_), .A2(new_n15474_), .B(new_n15469_), .ZN(new_n15475_));
  AOI21_X1   g15283(.A1(new_n15475_), .A2(new_n860_), .B(new_n15074_), .ZN(new_n15476_));
  NAND2_X1   g15284(.A1(new_n15474_), .A2(new_n15076_), .ZN(new_n15477_));
  INV_X1     g15285(.I(new_n15469_), .ZN(new_n15478_));
  AOI21_X1   g15286(.A1(new_n15477_), .A2(new_n15478_), .B(new_n860_), .ZN(new_n15479_));
  OAI21_X1   g15287(.A1(new_n15476_), .A2(new_n15479_), .B(\asqrt[55] ), .ZN(new_n15480_));
  NAND3_X1   g15288(.A1(new_n15473_), .A2(new_n634_), .A3(new_n15480_), .ZN(new_n15481_));
  INV_X1     g15289(.I(new_n15070_), .ZN(new_n15482_));
  NOR3_X1    g15290(.A1(new_n15476_), .A2(\asqrt[55] ), .A3(new_n15479_), .ZN(new_n15483_));
  OAI21_X1   g15291(.A1(new_n15482_), .A2(new_n15483_), .B(new_n15480_), .ZN(new_n15484_));
  NAND2_X1   g15292(.A1(new_n15484_), .A2(\asqrt[56] ), .ZN(new_n15485_));
  NOR2_X1    g15293(.A1(new_n15038_), .A2(\asqrt[62] ), .ZN(new_n15486_));
  INV_X1     g15294(.I(new_n15057_), .ZN(new_n15487_));
  NOR2_X1    g15295(.A1(new_n15487_), .A2(new_n15486_), .ZN(new_n15488_));
  XOR2_X1    g15296(.A1(new_n15048_), .A2(new_n14498_), .Z(new_n15489_));
  OAI21_X1   g15297(.A1(\asqrt[9] ), .A2(new_n15488_), .B(new_n15489_), .ZN(new_n15490_));
  INV_X1     g15298(.I(new_n15490_), .ZN(new_n15491_));
  NAND2_X1   g15299(.A1(new_n15010_), .A2(new_n337_), .ZN(new_n15492_));
  AOI21_X1   g15300(.A1(new_n15492_), .A2(new_n15030_), .B(\asqrt[9] ), .ZN(new_n15493_));
  XOR2_X1    g15301(.A1(new_n15493_), .A2(new_n14988_), .Z(new_n15494_));
  INV_X1     g15302(.I(new_n15494_), .ZN(new_n15495_));
  AOI21_X1   g15303(.A1(new_n15008_), .A2(new_n15021_), .B(\asqrt[9] ), .ZN(new_n15496_));
  XOR2_X1    g15304(.A1(new_n15496_), .A2(new_n14992_), .Z(new_n15497_));
  INV_X1     g15305(.I(new_n15497_), .ZN(new_n15498_));
  NAND2_X1   g15306(.A1(new_n15017_), .A2(new_n531_), .ZN(new_n15499_));
  AOI21_X1   g15307(.A1(new_n15499_), .A2(new_n15007_), .B(\asqrt[9] ), .ZN(new_n15500_));
  XOR2_X1    g15308(.A1(new_n15500_), .A2(new_n14995_), .Z(new_n15501_));
  INV_X1     g15309(.I(new_n15501_), .ZN(new_n15502_));
  AOI21_X1   g15310(.A1(new_n15015_), .A2(new_n15004_), .B(\asqrt[9] ), .ZN(new_n15503_));
  XOR2_X1    g15311(.A1(new_n15503_), .A2(new_n14997_), .Z(new_n15504_));
  OAI21_X1   g15312(.A1(new_n15484_), .A2(\asqrt[56] ), .B(new_n15068_), .ZN(new_n15505_));
  NAND3_X1   g15313(.A1(new_n15505_), .A2(new_n15485_), .A3(new_n531_), .ZN(new_n15506_));
  AOI21_X1   g15314(.A1(new_n15505_), .A2(new_n15485_), .B(new_n531_), .ZN(new_n15507_));
  AOI21_X1   g15315(.A1(new_n15504_), .A2(new_n15506_), .B(new_n15507_), .ZN(new_n15508_));
  AOI21_X1   g15316(.A1(new_n15508_), .A2(new_n423_), .B(new_n15502_), .ZN(new_n15509_));
  NAND2_X1   g15317(.A1(new_n15506_), .A2(new_n15504_), .ZN(new_n15510_));
  INV_X1     g15318(.I(new_n15507_), .ZN(new_n15511_));
  AOI21_X1   g15319(.A1(new_n15510_), .A2(new_n15511_), .B(new_n423_), .ZN(new_n15512_));
  NOR3_X1    g15320(.A1(new_n15509_), .A2(\asqrt[59] ), .A3(new_n15512_), .ZN(new_n15513_));
  NOR2_X1    g15321(.A1(new_n15513_), .A2(new_n15498_), .ZN(new_n15514_));
  OAI21_X1   g15322(.A1(new_n15509_), .A2(new_n15512_), .B(\asqrt[59] ), .ZN(new_n15515_));
  INV_X1     g15323(.I(new_n15515_), .ZN(new_n15516_));
  NOR2_X1    g15324(.A1(new_n15514_), .A2(new_n15516_), .ZN(new_n15517_));
  AOI21_X1   g15325(.A1(new_n15517_), .A2(new_n266_), .B(new_n15495_), .ZN(new_n15518_));
  INV_X1     g15326(.I(new_n15504_), .ZN(new_n15519_));
  AOI21_X1   g15327(.A1(new_n15473_), .A2(new_n15480_), .B(new_n634_), .ZN(new_n15520_));
  AOI21_X1   g15328(.A1(new_n15068_), .A2(new_n15481_), .B(new_n15520_), .ZN(new_n15521_));
  AOI21_X1   g15329(.A1(new_n15521_), .A2(new_n531_), .B(new_n15519_), .ZN(new_n15522_));
  NOR3_X1    g15330(.A1(new_n15522_), .A2(\asqrt[58] ), .A3(new_n15507_), .ZN(new_n15523_));
  OAI21_X1   g15331(.A1(new_n15522_), .A2(new_n15507_), .B(\asqrt[58] ), .ZN(new_n15524_));
  OAI21_X1   g15332(.A1(new_n15502_), .A2(new_n15523_), .B(new_n15524_), .ZN(new_n15525_));
  OAI21_X1   g15333(.A1(new_n15525_), .A2(\asqrt[59] ), .B(new_n15497_), .ZN(new_n15526_));
  AOI21_X1   g15334(.A1(new_n15526_), .A2(new_n15515_), .B(new_n266_), .ZN(new_n15527_));
  OAI21_X1   g15335(.A1(new_n15518_), .A2(new_n15527_), .B(\asqrt[61] ), .ZN(new_n15528_));
  AOI21_X1   g15336(.A1(new_n15039_), .A2(new_n15033_), .B(\asqrt[9] ), .ZN(new_n15529_));
  XOR2_X1    g15337(.A1(new_n15529_), .A2(new_n14985_), .Z(new_n15530_));
  OAI21_X1   g15338(.A1(new_n15498_), .A2(new_n15513_), .B(new_n15515_), .ZN(new_n15531_));
  OAI21_X1   g15339(.A1(new_n15531_), .A2(\asqrt[60] ), .B(new_n15494_), .ZN(new_n15532_));
  OAI21_X1   g15340(.A1(new_n15514_), .A2(new_n15516_), .B(\asqrt[60] ), .ZN(new_n15533_));
  NAND3_X1   g15341(.A1(new_n15532_), .A2(new_n239_), .A3(new_n15533_), .ZN(new_n15534_));
  NAND2_X1   g15342(.A1(new_n15534_), .A2(new_n15530_), .ZN(new_n15535_));
  NAND2_X1   g15343(.A1(new_n15535_), .A2(new_n15528_), .ZN(new_n15536_));
  AOI21_X1   g15344(.A1(new_n15532_), .A2(new_n15533_), .B(new_n239_), .ZN(new_n15537_));
  NAND3_X1   g15345(.A1(new_n15526_), .A2(new_n266_), .A3(new_n15515_), .ZN(new_n15538_));
  AOI21_X1   g15346(.A1(new_n15494_), .A2(new_n15538_), .B(new_n15527_), .ZN(new_n15539_));
  INV_X1     g15347(.I(new_n15530_), .ZN(new_n15540_));
  AOI21_X1   g15348(.A1(new_n15539_), .A2(new_n239_), .B(new_n15540_), .ZN(new_n15541_));
  OAI21_X1   g15349(.A1(new_n15541_), .A2(new_n15537_), .B(new_n201_), .ZN(new_n15542_));
  NAND3_X1   g15350(.A1(new_n15535_), .A2(\asqrt[62] ), .A3(new_n15528_), .ZN(new_n15543_));
  AOI21_X1   g15351(.A1(new_n15032_), .A2(new_n15204_), .B(\asqrt[9] ), .ZN(new_n15544_));
  XOR2_X1    g15352(.A1(new_n15544_), .A2(new_n15036_), .Z(new_n15545_));
  INV_X1     g15353(.I(new_n15545_), .ZN(new_n15546_));
  AOI22_X1   g15354(.A1(new_n15542_), .A2(new_n15543_), .B1(new_n15536_), .B2(new_n15546_), .ZN(new_n15547_));
  NOR2_X1    g15355(.A1(new_n15051_), .A2(new_n14983_), .ZN(new_n15548_));
  OAI21_X1   g15356(.A1(\asqrt[9] ), .A2(new_n15548_), .B(new_n15058_), .ZN(new_n15549_));
  INV_X1     g15357(.I(new_n15549_), .ZN(new_n15550_));
  OAI21_X1   g15358(.A1(new_n15547_), .A2(new_n15491_), .B(new_n15550_), .ZN(new_n15551_));
  OAI21_X1   g15359(.A1(new_n15536_), .A2(\asqrt[62] ), .B(new_n15545_), .ZN(new_n15552_));
  NAND2_X1   g15360(.A1(new_n15536_), .A2(\asqrt[62] ), .ZN(new_n15553_));
  NAND3_X1   g15361(.A1(new_n15552_), .A2(new_n15553_), .A3(new_n15491_), .ZN(new_n15554_));
  NAND2_X1   g15362(.A1(new_n15221_), .A2(new_n14982_), .ZN(new_n15555_));
  XOR2_X1    g15363(.A1(new_n15051_), .A2(new_n14983_), .Z(new_n15556_));
  NAND3_X1   g15364(.A1(new_n15555_), .A2(\asqrt[63] ), .A3(new_n15556_), .ZN(new_n15557_));
  INV_X1     g15365(.I(new_n15219_), .ZN(new_n15558_));
  NAND4_X1   g15366(.A1(new_n15558_), .A2(new_n14983_), .A3(new_n15058_), .A4(new_n15065_), .ZN(new_n15559_));
  NAND2_X1   g15367(.A1(new_n15557_), .A2(new_n15559_), .ZN(new_n15560_));
  INV_X1     g15368(.I(new_n15560_), .ZN(new_n15561_));
  NAND4_X1   g15369(.A1(new_n15551_), .A2(new_n193_), .A3(new_n15554_), .A4(new_n15561_), .ZN(\asqrt[8] ));
  AOI21_X1   g15370(.A1(new_n15481_), .A2(new_n15485_), .B(\asqrt[8] ), .ZN(new_n15563_));
  XOR2_X1    g15371(.A1(new_n15563_), .A2(new_n15068_), .Z(new_n15564_));
  INV_X1     g15372(.I(new_n15480_), .ZN(new_n15565_));
  NOR2_X1    g15373(.A1(new_n15565_), .A2(new_n15483_), .ZN(new_n15566_));
  NOR2_X1    g15374(.A1(\asqrt[8] ), .A2(new_n15566_), .ZN(new_n15567_));
  XOR2_X1    g15375(.A1(new_n15567_), .A2(new_n15070_), .Z(new_n15568_));
  NOR2_X1    g15376(.A1(new_n15470_), .A2(new_n15479_), .ZN(new_n15569_));
  NOR2_X1    g15377(.A1(\asqrt[8] ), .A2(new_n15569_), .ZN(new_n15570_));
  XOR2_X1    g15378(.A1(new_n15570_), .A2(new_n15073_), .Z(new_n15571_));
  AOI21_X1   g15379(.A1(new_n15474_), .A2(new_n15478_), .B(\asqrt[8] ), .ZN(new_n15572_));
  XOR2_X1    g15380(.A1(new_n15572_), .A2(new_n15076_), .Z(new_n15573_));
  INV_X1     g15381(.I(new_n15573_), .ZN(new_n15574_));
  AOI21_X1   g15382(.A1(new_n15460_), .A2(new_n15468_), .B(\asqrt[8] ), .ZN(new_n15575_));
  XOR2_X1    g15383(.A1(new_n15575_), .A2(new_n15080_), .Z(new_n15576_));
  INV_X1     g15384(.I(new_n15576_), .ZN(new_n15577_));
  XOR2_X1    g15385(.A1(new_n15451_), .A2(\asqrt[51] ), .Z(new_n15578_));
  NOR2_X1    g15386(.A1(\asqrt[8] ), .A2(new_n15578_), .ZN(new_n15579_));
  XOR2_X1    g15387(.A1(new_n15579_), .A2(new_n15082_), .Z(new_n15580_));
  NOR2_X1    g15388(.A1(new_n15449_), .A2(new_n15458_), .ZN(new_n15581_));
  NOR2_X1    g15389(.A1(\asqrt[8] ), .A2(new_n15581_), .ZN(new_n15582_));
  XOR2_X1    g15390(.A1(new_n15582_), .A2(new_n15085_), .Z(new_n15583_));
  AOI21_X1   g15391(.A1(new_n15453_), .A2(new_n15457_), .B(\asqrt[8] ), .ZN(new_n15584_));
  XOR2_X1    g15392(.A1(new_n15584_), .A2(new_n15088_), .Z(new_n15585_));
  INV_X1     g15393(.I(new_n15585_), .ZN(new_n15586_));
  AOI21_X1   g15394(.A1(new_n15439_), .A2(new_n15447_), .B(\asqrt[8] ), .ZN(new_n15587_));
  XOR2_X1    g15395(.A1(new_n15587_), .A2(new_n15092_), .Z(new_n15588_));
  INV_X1     g15396(.I(new_n15588_), .ZN(new_n15589_));
  XOR2_X1    g15397(.A1(new_n15430_), .A2(\asqrt[47] ), .Z(new_n15590_));
  NOR2_X1    g15398(.A1(\asqrt[8] ), .A2(new_n15590_), .ZN(new_n15591_));
  XOR2_X1    g15399(.A1(new_n15591_), .A2(new_n15094_), .Z(new_n15592_));
  NOR2_X1    g15400(.A1(new_n15428_), .A2(new_n15437_), .ZN(new_n15593_));
  NOR2_X1    g15401(.A1(\asqrt[8] ), .A2(new_n15593_), .ZN(new_n15594_));
  XOR2_X1    g15402(.A1(new_n15594_), .A2(new_n15097_), .Z(new_n15595_));
  AOI21_X1   g15403(.A1(new_n15432_), .A2(new_n15436_), .B(\asqrt[8] ), .ZN(new_n15596_));
  XOR2_X1    g15404(.A1(new_n15596_), .A2(new_n15100_), .Z(new_n15597_));
  INV_X1     g15405(.I(new_n15597_), .ZN(new_n15598_));
  AOI21_X1   g15406(.A1(new_n15418_), .A2(new_n15426_), .B(\asqrt[8] ), .ZN(new_n15599_));
  XOR2_X1    g15407(.A1(new_n15599_), .A2(new_n15104_), .Z(new_n15600_));
  INV_X1     g15408(.I(new_n15600_), .ZN(new_n15601_));
  XOR2_X1    g15409(.A1(new_n15409_), .A2(\asqrt[43] ), .Z(new_n15602_));
  NOR2_X1    g15410(.A1(\asqrt[8] ), .A2(new_n15602_), .ZN(new_n15603_));
  XOR2_X1    g15411(.A1(new_n15603_), .A2(new_n15106_), .Z(new_n15604_));
  NOR2_X1    g15412(.A1(new_n15407_), .A2(new_n15416_), .ZN(new_n15605_));
  NOR2_X1    g15413(.A1(\asqrt[8] ), .A2(new_n15605_), .ZN(new_n15606_));
  XOR2_X1    g15414(.A1(new_n15606_), .A2(new_n15109_), .Z(new_n15607_));
  AOI21_X1   g15415(.A1(new_n15411_), .A2(new_n15415_), .B(\asqrt[8] ), .ZN(new_n15608_));
  XOR2_X1    g15416(.A1(new_n15608_), .A2(new_n15112_), .Z(new_n15609_));
  INV_X1     g15417(.I(new_n15609_), .ZN(new_n15610_));
  AOI21_X1   g15418(.A1(new_n15397_), .A2(new_n15405_), .B(\asqrt[8] ), .ZN(new_n15611_));
  XOR2_X1    g15419(.A1(new_n15611_), .A2(new_n15116_), .Z(new_n15612_));
  INV_X1     g15420(.I(new_n15612_), .ZN(new_n15613_));
  XOR2_X1    g15421(.A1(new_n15388_), .A2(\asqrt[39] ), .Z(new_n15614_));
  NOR2_X1    g15422(.A1(\asqrt[8] ), .A2(new_n15614_), .ZN(new_n15615_));
  XOR2_X1    g15423(.A1(new_n15615_), .A2(new_n15118_), .Z(new_n15616_));
  NOR2_X1    g15424(.A1(new_n15386_), .A2(new_n15395_), .ZN(new_n15617_));
  NOR2_X1    g15425(.A1(\asqrt[8] ), .A2(new_n15617_), .ZN(new_n15618_));
  XOR2_X1    g15426(.A1(new_n15618_), .A2(new_n15121_), .Z(new_n15619_));
  AOI21_X1   g15427(.A1(new_n15390_), .A2(new_n15394_), .B(\asqrt[8] ), .ZN(new_n15620_));
  XOR2_X1    g15428(.A1(new_n15620_), .A2(new_n15124_), .Z(new_n15621_));
  INV_X1     g15429(.I(new_n15621_), .ZN(new_n15622_));
  AOI21_X1   g15430(.A1(new_n15376_), .A2(new_n15384_), .B(\asqrt[8] ), .ZN(new_n15623_));
  XOR2_X1    g15431(.A1(new_n15623_), .A2(new_n15128_), .Z(new_n15624_));
  INV_X1     g15432(.I(new_n15624_), .ZN(new_n15625_));
  XOR2_X1    g15433(.A1(new_n15367_), .A2(\asqrt[35] ), .Z(new_n15626_));
  NOR2_X1    g15434(.A1(\asqrt[8] ), .A2(new_n15626_), .ZN(new_n15627_));
  XOR2_X1    g15435(.A1(new_n15627_), .A2(new_n15130_), .Z(new_n15628_));
  NOR2_X1    g15436(.A1(new_n15365_), .A2(new_n15374_), .ZN(new_n15629_));
  NOR2_X1    g15437(.A1(\asqrt[8] ), .A2(new_n15629_), .ZN(new_n15630_));
  XOR2_X1    g15438(.A1(new_n15630_), .A2(new_n15133_), .Z(new_n15631_));
  AOI21_X1   g15439(.A1(new_n15369_), .A2(new_n15373_), .B(\asqrt[8] ), .ZN(new_n15632_));
  XOR2_X1    g15440(.A1(new_n15632_), .A2(new_n15136_), .Z(new_n15633_));
  INV_X1     g15441(.I(new_n15633_), .ZN(new_n15634_));
  AOI21_X1   g15442(.A1(new_n15355_), .A2(new_n15363_), .B(\asqrt[8] ), .ZN(new_n15635_));
  XOR2_X1    g15443(.A1(new_n15635_), .A2(new_n15140_), .Z(new_n15636_));
  INV_X1     g15444(.I(new_n15636_), .ZN(new_n15637_));
  XOR2_X1    g15445(.A1(new_n15346_), .A2(\asqrt[31] ), .Z(new_n15638_));
  NOR2_X1    g15446(.A1(\asqrt[8] ), .A2(new_n15638_), .ZN(new_n15639_));
  XOR2_X1    g15447(.A1(new_n15639_), .A2(new_n15142_), .Z(new_n15640_));
  NOR2_X1    g15448(.A1(new_n15344_), .A2(new_n15353_), .ZN(new_n15641_));
  NOR2_X1    g15449(.A1(\asqrt[8] ), .A2(new_n15641_), .ZN(new_n15642_));
  XOR2_X1    g15450(.A1(new_n15642_), .A2(new_n15145_), .Z(new_n15643_));
  AOI21_X1   g15451(.A1(new_n15348_), .A2(new_n15352_), .B(\asqrt[8] ), .ZN(new_n15644_));
  XOR2_X1    g15452(.A1(new_n15644_), .A2(new_n15148_), .Z(new_n15645_));
  INV_X1     g15453(.I(new_n15645_), .ZN(new_n15646_));
  AOI21_X1   g15454(.A1(new_n15334_), .A2(new_n15342_), .B(\asqrt[8] ), .ZN(new_n15647_));
  XOR2_X1    g15455(.A1(new_n15647_), .A2(new_n15152_), .Z(new_n15648_));
  INV_X1     g15456(.I(new_n15648_), .ZN(new_n15649_));
  XOR2_X1    g15457(.A1(new_n15325_), .A2(\asqrt[27] ), .Z(new_n15650_));
  NOR2_X1    g15458(.A1(\asqrt[8] ), .A2(new_n15650_), .ZN(new_n15651_));
  XOR2_X1    g15459(.A1(new_n15651_), .A2(new_n15154_), .Z(new_n15652_));
  NOR2_X1    g15460(.A1(new_n15323_), .A2(new_n15332_), .ZN(new_n15653_));
  NOR2_X1    g15461(.A1(\asqrt[8] ), .A2(new_n15653_), .ZN(new_n15654_));
  XOR2_X1    g15462(.A1(new_n15654_), .A2(new_n15157_), .Z(new_n15655_));
  AOI21_X1   g15463(.A1(new_n15327_), .A2(new_n15331_), .B(\asqrt[8] ), .ZN(new_n15656_));
  XOR2_X1    g15464(.A1(new_n15656_), .A2(new_n15160_), .Z(new_n15657_));
  INV_X1     g15465(.I(new_n15657_), .ZN(new_n15658_));
  AOI21_X1   g15466(.A1(new_n15313_), .A2(new_n15321_), .B(\asqrt[8] ), .ZN(new_n15659_));
  XOR2_X1    g15467(.A1(new_n15659_), .A2(new_n15164_), .Z(new_n15660_));
  INV_X1     g15468(.I(new_n15660_), .ZN(new_n15661_));
  XOR2_X1    g15469(.A1(new_n15304_), .A2(\asqrt[23] ), .Z(new_n15662_));
  NOR2_X1    g15470(.A1(\asqrt[8] ), .A2(new_n15662_), .ZN(new_n15663_));
  XOR2_X1    g15471(.A1(new_n15663_), .A2(new_n15166_), .Z(new_n15664_));
  NOR2_X1    g15472(.A1(new_n15302_), .A2(new_n15311_), .ZN(new_n15665_));
  NOR2_X1    g15473(.A1(\asqrt[8] ), .A2(new_n15665_), .ZN(new_n15666_));
  XOR2_X1    g15474(.A1(new_n15666_), .A2(new_n15169_), .Z(new_n15667_));
  AOI21_X1   g15475(.A1(new_n15306_), .A2(new_n15310_), .B(\asqrt[8] ), .ZN(new_n15668_));
  XOR2_X1    g15476(.A1(new_n15668_), .A2(new_n15172_), .Z(new_n15669_));
  INV_X1     g15477(.I(new_n15669_), .ZN(new_n15670_));
  AOI21_X1   g15478(.A1(new_n15292_), .A2(new_n15300_), .B(\asqrt[8] ), .ZN(new_n15671_));
  XOR2_X1    g15479(.A1(new_n15671_), .A2(new_n15176_), .Z(new_n15672_));
  INV_X1     g15480(.I(new_n15672_), .ZN(new_n15673_));
  XOR2_X1    g15481(.A1(new_n15283_), .A2(\asqrt[19] ), .Z(new_n15674_));
  NOR2_X1    g15482(.A1(\asqrt[8] ), .A2(new_n15674_), .ZN(new_n15675_));
  XOR2_X1    g15483(.A1(new_n15675_), .A2(new_n15178_), .Z(new_n15676_));
  NOR2_X1    g15484(.A1(new_n15281_), .A2(new_n15290_), .ZN(new_n15677_));
  NOR2_X1    g15485(.A1(\asqrt[8] ), .A2(new_n15677_), .ZN(new_n15678_));
  XOR2_X1    g15486(.A1(new_n15678_), .A2(new_n15181_), .Z(new_n15679_));
  AOI21_X1   g15487(.A1(new_n15285_), .A2(new_n15289_), .B(\asqrt[8] ), .ZN(new_n15680_));
  XOR2_X1    g15488(.A1(new_n15680_), .A2(new_n15184_), .Z(new_n15681_));
  INV_X1     g15489(.I(new_n15681_), .ZN(new_n15682_));
  AOI21_X1   g15490(.A1(new_n15271_), .A2(new_n15279_), .B(\asqrt[8] ), .ZN(new_n15683_));
  XOR2_X1    g15491(.A1(new_n15683_), .A2(new_n15188_), .Z(new_n15684_));
  INV_X1     g15492(.I(new_n15684_), .ZN(new_n15685_));
  XOR2_X1    g15493(.A1(new_n15262_), .A2(\asqrt[15] ), .Z(new_n15686_));
  NOR2_X1    g15494(.A1(\asqrt[8] ), .A2(new_n15686_), .ZN(new_n15687_));
  XOR2_X1    g15495(.A1(new_n15687_), .A2(new_n15190_), .Z(new_n15688_));
  NOR2_X1    g15496(.A1(new_n15260_), .A2(new_n15269_), .ZN(new_n15689_));
  NOR2_X1    g15497(.A1(\asqrt[8] ), .A2(new_n15689_), .ZN(new_n15690_));
  XOR2_X1    g15498(.A1(new_n15690_), .A2(new_n15193_), .Z(new_n15691_));
  AOI21_X1   g15499(.A1(new_n15264_), .A2(new_n15268_), .B(\asqrt[8] ), .ZN(new_n15692_));
  XOR2_X1    g15500(.A1(new_n15692_), .A2(new_n15196_), .Z(new_n15693_));
  INV_X1     g15501(.I(new_n15693_), .ZN(new_n15694_));
  AOI21_X1   g15502(.A1(new_n15250_), .A2(new_n15258_), .B(\asqrt[8] ), .ZN(new_n15695_));
  XOR2_X1    g15503(.A1(new_n15695_), .A2(new_n15203_), .Z(new_n15696_));
  INV_X1     g15504(.I(new_n15696_), .ZN(new_n15697_));
  AOI21_X1   g15505(.A1(new_n15240_), .A2(new_n15249_), .B(\asqrt[8] ), .ZN(new_n15698_));
  XOR2_X1    g15506(.A1(new_n15698_), .A2(new_n15224_), .Z(new_n15699_));
  NAND2_X1   g15507(.A1(\asqrt[9] ), .A2(new_n15225_), .ZN(new_n15700_));
  NOR2_X1    g15508(.A1(new_n15237_), .A2(\a[18] ), .ZN(new_n15701_));
  AOI22_X1   g15509(.A1(new_n15700_), .A2(new_n15237_), .B1(\asqrt[9] ), .B2(new_n15701_), .ZN(new_n15702_));
  OAI21_X1   g15510(.A1(new_n15221_), .A2(new_n15225_), .B(new_n15234_), .ZN(new_n15703_));
  AOI21_X1   g15511(.A1(new_n15230_), .A2(new_n15703_), .B(\asqrt[8] ), .ZN(new_n15704_));
  XOR2_X1    g15512(.A1(new_n15704_), .A2(new_n15702_), .Z(new_n15705_));
  NAND2_X1   g15513(.A1(new_n15551_), .A2(new_n193_), .ZN(new_n15706_));
  NOR2_X1    g15514(.A1(new_n15541_), .A2(new_n15537_), .ZN(new_n15707_));
  AOI21_X1   g15515(.A1(new_n15707_), .A2(new_n201_), .B(new_n15546_), .ZN(new_n15708_));
  OAI21_X1   g15516(.A1(new_n15707_), .A2(new_n201_), .B(new_n15491_), .ZN(new_n15709_));
  NOR2_X1    g15517(.A1(new_n15708_), .A2(new_n15709_), .ZN(new_n15710_));
  NAND3_X1   g15518(.A1(new_n15557_), .A2(\asqrt[9] ), .A3(new_n15559_), .ZN(new_n15711_));
  NOR3_X1    g15519(.A1(new_n15706_), .A2(new_n15710_), .A3(new_n15711_), .ZN(new_n15712_));
  AOI21_X1   g15520(.A1(new_n15535_), .A2(new_n15528_), .B(\asqrt[62] ), .ZN(new_n15713_));
  NOR3_X1    g15521(.A1(new_n15541_), .A2(new_n201_), .A3(new_n15537_), .ZN(new_n15714_));
  OAI22_X1   g15522(.A1(new_n15714_), .A2(new_n15713_), .B1(new_n15707_), .B2(new_n15545_), .ZN(new_n15715_));
  AOI21_X1   g15523(.A1(new_n15715_), .A2(new_n15490_), .B(new_n15549_), .ZN(new_n15716_));
  NOR4_X1    g15524(.A1(new_n15716_), .A2(\asqrt[63] ), .A3(new_n15710_), .A4(new_n15560_), .ZN(new_n15717_));
  NOR2_X1    g15525(.A1(new_n15717_), .A2(new_n15228_), .ZN(new_n15718_));
  OAI21_X1   g15526(.A1(new_n15718_), .A2(new_n15712_), .B(new_n15225_), .ZN(new_n15719_));
  NOR3_X1    g15527(.A1(new_n15716_), .A2(\asqrt[63] ), .A3(new_n15710_), .ZN(new_n15720_));
  NAND4_X1   g15528(.A1(new_n15720_), .A2(\asqrt[9] ), .A3(new_n15557_), .A4(new_n15559_), .ZN(new_n15721_));
  NAND2_X1   g15529(.A1(\asqrt[8] ), .A2(new_n15226_), .ZN(new_n15722_));
  NAND3_X1   g15530(.A1(new_n15721_), .A2(new_n15722_), .A3(\a[18] ), .ZN(new_n15723_));
  NAND2_X1   g15531(.A1(new_n15723_), .A2(new_n15719_), .ZN(new_n15724_));
  NOR2_X1    g15532(.A1(\a[14] ), .A2(\a[15] ), .ZN(new_n15725_));
  INV_X1     g15533(.I(new_n15725_), .ZN(new_n15726_));
  NAND3_X1   g15534(.A1(\asqrt[8] ), .A2(\a[16] ), .A3(new_n15726_), .ZN(new_n15727_));
  INV_X1     g15535(.I(\a[16] ), .ZN(new_n15728_));
  OAI21_X1   g15536(.A1(\asqrt[8] ), .A2(new_n15728_), .B(new_n15725_), .ZN(new_n15729_));
  AOI21_X1   g15537(.A1(new_n15729_), .A2(new_n15727_), .B(new_n15221_), .ZN(new_n15730_));
  NAND2_X1   g15538(.A1(new_n15725_), .A2(new_n15728_), .ZN(new_n15731_));
  NAND3_X1   g15539(.A1(new_n15061_), .A2(new_n15063_), .A3(new_n15731_), .ZN(new_n15732_));
  NAND2_X1   g15540(.A1(new_n15213_), .A2(new_n15732_), .ZN(new_n15733_));
  NAND3_X1   g15541(.A1(\asqrt[8] ), .A2(\a[16] ), .A3(new_n15733_), .ZN(new_n15734_));
  INV_X1     g15542(.I(\a[17] ), .ZN(new_n15735_));
  NAND3_X1   g15543(.A1(\asqrt[8] ), .A2(new_n15728_), .A3(new_n15735_), .ZN(new_n15736_));
  OAI21_X1   g15544(.A1(new_n15717_), .A2(\a[16] ), .B(\a[17] ), .ZN(new_n15737_));
  NAND3_X1   g15545(.A1(new_n15737_), .A2(new_n15734_), .A3(new_n15736_), .ZN(new_n15738_));
  NOR3_X1    g15546(.A1(new_n15738_), .A2(new_n15730_), .A3(\asqrt[10] ), .ZN(new_n15739_));
  OAI21_X1   g15547(.A1(new_n15738_), .A2(new_n15730_), .B(\asqrt[10] ), .ZN(new_n15740_));
  OAI21_X1   g15548(.A1(new_n15724_), .A2(new_n15739_), .B(new_n15740_), .ZN(new_n15741_));
  OAI21_X1   g15549(.A1(new_n15741_), .A2(\asqrt[11] ), .B(new_n15705_), .ZN(new_n15742_));
  NAND2_X1   g15550(.A1(new_n15741_), .A2(\asqrt[11] ), .ZN(new_n15743_));
  NAND3_X1   g15551(.A1(new_n15742_), .A2(new_n15743_), .A3(new_n13690_), .ZN(new_n15744_));
  AOI21_X1   g15552(.A1(new_n15742_), .A2(new_n15743_), .B(new_n13690_), .ZN(new_n15745_));
  AOI21_X1   g15553(.A1(new_n15699_), .A2(new_n15744_), .B(new_n15745_), .ZN(new_n15746_));
  AOI21_X1   g15554(.A1(new_n15746_), .A2(new_n13228_), .B(new_n15697_), .ZN(new_n15747_));
  NAND2_X1   g15555(.A1(new_n15744_), .A2(new_n15699_), .ZN(new_n15748_));
  INV_X1     g15556(.I(new_n15705_), .ZN(new_n15749_));
  INV_X1     g15557(.I(new_n15724_), .ZN(new_n15750_));
  NOR3_X1    g15558(.A1(new_n15717_), .A2(new_n15728_), .A3(new_n15725_), .ZN(new_n15751_));
  AOI21_X1   g15559(.A1(new_n15717_), .A2(\a[16] ), .B(new_n15726_), .ZN(new_n15752_));
  OAI21_X1   g15560(.A1(new_n15751_), .A2(new_n15752_), .B(\asqrt[9] ), .ZN(new_n15753_));
  INV_X1     g15561(.I(new_n15733_), .ZN(new_n15754_));
  NOR3_X1    g15562(.A1(new_n15717_), .A2(new_n15728_), .A3(new_n15754_), .ZN(new_n15755_));
  NOR3_X1    g15563(.A1(new_n15717_), .A2(\a[16] ), .A3(\a[17] ), .ZN(new_n15756_));
  AOI21_X1   g15564(.A1(\asqrt[8] ), .A2(new_n15728_), .B(new_n15735_), .ZN(new_n15757_));
  NOR3_X1    g15565(.A1(new_n15755_), .A2(new_n15756_), .A3(new_n15757_), .ZN(new_n15758_));
  NAND3_X1   g15566(.A1(new_n15753_), .A2(new_n15758_), .A3(new_n14690_), .ZN(new_n15759_));
  AOI21_X1   g15567(.A1(new_n15753_), .A2(new_n15758_), .B(new_n14690_), .ZN(new_n15760_));
  AOI21_X1   g15568(.A1(new_n15750_), .A2(new_n15759_), .B(new_n15760_), .ZN(new_n15761_));
  AOI21_X1   g15569(.A1(new_n15761_), .A2(new_n14207_), .B(new_n15749_), .ZN(new_n15762_));
  NAND2_X1   g15570(.A1(new_n15750_), .A2(new_n15759_), .ZN(new_n15763_));
  AOI21_X1   g15571(.A1(new_n15763_), .A2(new_n15740_), .B(new_n14207_), .ZN(new_n15764_));
  OAI21_X1   g15572(.A1(new_n15762_), .A2(new_n15764_), .B(\asqrt[12] ), .ZN(new_n15765_));
  AOI21_X1   g15573(.A1(new_n15748_), .A2(new_n15765_), .B(new_n13228_), .ZN(new_n15766_));
  NOR3_X1    g15574(.A1(new_n15747_), .A2(\asqrt[14] ), .A3(new_n15766_), .ZN(new_n15767_));
  OAI21_X1   g15575(.A1(new_n15747_), .A2(new_n15766_), .B(\asqrt[14] ), .ZN(new_n15768_));
  OAI21_X1   g15576(.A1(new_n15694_), .A2(new_n15767_), .B(new_n15768_), .ZN(new_n15769_));
  OAI21_X1   g15577(.A1(new_n15769_), .A2(\asqrt[15] ), .B(new_n15691_), .ZN(new_n15770_));
  NAND2_X1   g15578(.A1(new_n15769_), .A2(\asqrt[15] ), .ZN(new_n15771_));
  NAND3_X1   g15579(.A1(new_n15770_), .A2(new_n15771_), .A3(new_n11802_), .ZN(new_n15772_));
  AOI21_X1   g15580(.A1(new_n15770_), .A2(new_n15771_), .B(new_n11802_), .ZN(new_n15773_));
  AOI21_X1   g15581(.A1(new_n15688_), .A2(new_n15772_), .B(new_n15773_), .ZN(new_n15774_));
  AOI21_X1   g15582(.A1(new_n15774_), .A2(new_n11373_), .B(new_n15685_), .ZN(new_n15775_));
  NAND2_X1   g15583(.A1(new_n15772_), .A2(new_n15688_), .ZN(new_n15776_));
  INV_X1     g15584(.I(new_n15691_), .ZN(new_n15777_));
  INV_X1     g15585(.I(new_n15699_), .ZN(new_n15778_));
  NOR3_X1    g15586(.A1(new_n15762_), .A2(\asqrt[12] ), .A3(new_n15764_), .ZN(new_n15779_));
  OAI21_X1   g15587(.A1(new_n15778_), .A2(new_n15779_), .B(new_n15765_), .ZN(new_n15780_));
  OAI21_X1   g15588(.A1(new_n15780_), .A2(\asqrt[13] ), .B(new_n15696_), .ZN(new_n15781_));
  NAND2_X1   g15589(.A1(new_n15780_), .A2(\asqrt[13] ), .ZN(new_n15782_));
  NAND3_X1   g15590(.A1(new_n15781_), .A2(new_n15782_), .A3(new_n12733_), .ZN(new_n15783_));
  AOI21_X1   g15591(.A1(new_n15781_), .A2(new_n15782_), .B(new_n12733_), .ZN(new_n15784_));
  AOI21_X1   g15592(.A1(new_n15693_), .A2(new_n15783_), .B(new_n15784_), .ZN(new_n15785_));
  AOI21_X1   g15593(.A1(new_n15785_), .A2(new_n12283_), .B(new_n15777_), .ZN(new_n15786_));
  NAND2_X1   g15594(.A1(new_n15783_), .A2(new_n15693_), .ZN(new_n15787_));
  AOI21_X1   g15595(.A1(new_n15787_), .A2(new_n15768_), .B(new_n12283_), .ZN(new_n15788_));
  OAI21_X1   g15596(.A1(new_n15786_), .A2(new_n15788_), .B(\asqrt[16] ), .ZN(new_n15789_));
  AOI21_X1   g15597(.A1(new_n15776_), .A2(new_n15789_), .B(new_n11373_), .ZN(new_n15790_));
  NOR3_X1    g15598(.A1(new_n15775_), .A2(\asqrt[18] ), .A3(new_n15790_), .ZN(new_n15791_));
  OAI21_X1   g15599(.A1(new_n15775_), .A2(new_n15790_), .B(\asqrt[18] ), .ZN(new_n15792_));
  OAI21_X1   g15600(.A1(new_n15682_), .A2(new_n15791_), .B(new_n15792_), .ZN(new_n15793_));
  OAI21_X1   g15601(.A1(new_n15793_), .A2(\asqrt[19] ), .B(new_n15679_), .ZN(new_n15794_));
  NAND2_X1   g15602(.A1(new_n15793_), .A2(\asqrt[19] ), .ZN(new_n15795_));
  NAND3_X1   g15603(.A1(new_n15794_), .A2(new_n15795_), .A3(new_n10052_), .ZN(new_n15796_));
  AOI21_X1   g15604(.A1(new_n15794_), .A2(new_n15795_), .B(new_n10052_), .ZN(new_n15797_));
  AOI21_X1   g15605(.A1(new_n15676_), .A2(new_n15796_), .B(new_n15797_), .ZN(new_n15798_));
  AOI21_X1   g15606(.A1(new_n15798_), .A2(new_n9656_), .B(new_n15673_), .ZN(new_n15799_));
  NAND2_X1   g15607(.A1(new_n15796_), .A2(new_n15676_), .ZN(new_n15800_));
  INV_X1     g15608(.I(new_n15679_), .ZN(new_n15801_));
  INV_X1     g15609(.I(new_n15688_), .ZN(new_n15802_));
  NOR3_X1    g15610(.A1(new_n15786_), .A2(\asqrt[16] ), .A3(new_n15788_), .ZN(new_n15803_));
  OAI21_X1   g15611(.A1(new_n15802_), .A2(new_n15803_), .B(new_n15789_), .ZN(new_n15804_));
  OAI21_X1   g15612(.A1(new_n15804_), .A2(\asqrt[17] ), .B(new_n15684_), .ZN(new_n15805_));
  NAND2_X1   g15613(.A1(new_n15804_), .A2(\asqrt[17] ), .ZN(new_n15806_));
  NAND3_X1   g15614(.A1(new_n15805_), .A2(new_n15806_), .A3(new_n10914_), .ZN(new_n15807_));
  AOI21_X1   g15615(.A1(new_n15805_), .A2(new_n15806_), .B(new_n10914_), .ZN(new_n15808_));
  AOI21_X1   g15616(.A1(new_n15681_), .A2(new_n15807_), .B(new_n15808_), .ZN(new_n15809_));
  AOI21_X1   g15617(.A1(new_n15809_), .A2(new_n10497_), .B(new_n15801_), .ZN(new_n15810_));
  NAND2_X1   g15618(.A1(new_n15807_), .A2(new_n15681_), .ZN(new_n15811_));
  AOI21_X1   g15619(.A1(new_n15811_), .A2(new_n15792_), .B(new_n10497_), .ZN(new_n15812_));
  OAI21_X1   g15620(.A1(new_n15810_), .A2(new_n15812_), .B(\asqrt[20] ), .ZN(new_n15813_));
  AOI21_X1   g15621(.A1(new_n15800_), .A2(new_n15813_), .B(new_n9656_), .ZN(new_n15814_));
  NOR3_X1    g15622(.A1(new_n15799_), .A2(\asqrt[22] ), .A3(new_n15814_), .ZN(new_n15815_));
  OAI21_X1   g15623(.A1(new_n15799_), .A2(new_n15814_), .B(\asqrt[22] ), .ZN(new_n15816_));
  OAI21_X1   g15624(.A1(new_n15670_), .A2(new_n15815_), .B(new_n15816_), .ZN(new_n15817_));
  OAI21_X1   g15625(.A1(new_n15817_), .A2(\asqrt[23] ), .B(new_n15667_), .ZN(new_n15818_));
  NAND2_X1   g15626(.A1(new_n15817_), .A2(\asqrt[23] ), .ZN(new_n15819_));
  NAND3_X1   g15627(.A1(new_n15818_), .A2(new_n15819_), .A3(new_n8440_), .ZN(new_n15820_));
  AOI21_X1   g15628(.A1(new_n15818_), .A2(new_n15819_), .B(new_n8440_), .ZN(new_n15821_));
  AOI21_X1   g15629(.A1(new_n15664_), .A2(new_n15820_), .B(new_n15821_), .ZN(new_n15822_));
  AOI21_X1   g15630(.A1(new_n15822_), .A2(new_n8077_), .B(new_n15661_), .ZN(new_n15823_));
  NAND2_X1   g15631(.A1(new_n15820_), .A2(new_n15664_), .ZN(new_n15824_));
  INV_X1     g15632(.I(new_n15667_), .ZN(new_n15825_));
  INV_X1     g15633(.I(new_n15676_), .ZN(new_n15826_));
  NOR3_X1    g15634(.A1(new_n15810_), .A2(\asqrt[20] ), .A3(new_n15812_), .ZN(new_n15827_));
  OAI21_X1   g15635(.A1(new_n15826_), .A2(new_n15827_), .B(new_n15813_), .ZN(new_n15828_));
  OAI21_X1   g15636(.A1(new_n15828_), .A2(\asqrt[21] ), .B(new_n15672_), .ZN(new_n15829_));
  NAND2_X1   g15637(.A1(new_n15828_), .A2(\asqrt[21] ), .ZN(new_n15830_));
  NAND3_X1   g15638(.A1(new_n15829_), .A2(new_n15830_), .A3(new_n9233_), .ZN(new_n15831_));
  AOI21_X1   g15639(.A1(new_n15829_), .A2(new_n15830_), .B(new_n9233_), .ZN(new_n15832_));
  AOI21_X1   g15640(.A1(new_n15669_), .A2(new_n15831_), .B(new_n15832_), .ZN(new_n15833_));
  AOI21_X1   g15641(.A1(new_n15833_), .A2(new_n8849_), .B(new_n15825_), .ZN(new_n15834_));
  NAND2_X1   g15642(.A1(new_n15831_), .A2(new_n15669_), .ZN(new_n15835_));
  AOI21_X1   g15643(.A1(new_n15835_), .A2(new_n15816_), .B(new_n8849_), .ZN(new_n15836_));
  OAI21_X1   g15644(.A1(new_n15834_), .A2(new_n15836_), .B(\asqrt[24] ), .ZN(new_n15837_));
  AOI21_X1   g15645(.A1(new_n15824_), .A2(new_n15837_), .B(new_n8077_), .ZN(new_n15838_));
  NOR3_X1    g15646(.A1(new_n15823_), .A2(\asqrt[26] ), .A3(new_n15838_), .ZN(new_n15839_));
  OAI21_X1   g15647(.A1(new_n15823_), .A2(new_n15838_), .B(\asqrt[26] ), .ZN(new_n15840_));
  OAI21_X1   g15648(.A1(new_n15658_), .A2(new_n15839_), .B(new_n15840_), .ZN(new_n15841_));
  OAI21_X1   g15649(.A1(new_n15841_), .A2(\asqrt[27] ), .B(new_n15655_), .ZN(new_n15842_));
  NAND2_X1   g15650(.A1(new_n15841_), .A2(\asqrt[27] ), .ZN(new_n15843_));
  NAND3_X1   g15651(.A1(new_n15842_), .A2(new_n15843_), .A3(new_n6966_), .ZN(new_n15844_));
  AOI21_X1   g15652(.A1(new_n15842_), .A2(new_n15843_), .B(new_n6966_), .ZN(new_n15845_));
  AOI21_X1   g15653(.A1(new_n15652_), .A2(new_n15844_), .B(new_n15845_), .ZN(new_n15846_));
  AOI21_X1   g15654(.A1(new_n15846_), .A2(new_n6636_), .B(new_n15649_), .ZN(new_n15847_));
  NAND2_X1   g15655(.A1(new_n15844_), .A2(new_n15652_), .ZN(new_n15848_));
  INV_X1     g15656(.I(new_n15655_), .ZN(new_n15849_));
  INV_X1     g15657(.I(new_n15664_), .ZN(new_n15850_));
  NOR3_X1    g15658(.A1(new_n15834_), .A2(\asqrt[24] ), .A3(new_n15836_), .ZN(new_n15851_));
  OAI21_X1   g15659(.A1(new_n15850_), .A2(new_n15851_), .B(new_n15837_), .ZN(new_n15852_));
  OAI21_X1   g15660(.A1(new_n15852_), .A2(\asqrt[25] ), .B(new_n15660_), .ZN(new_n15853_));
  NAND2_X1   g15661(.A1(new_n15852_), .A2(\asqrt[25] ), .ZN(new_n15854_));
  NAND3_X1   g15662(.A1(new_n15853_), .A2(new_n15854_), .A3(new_n7690_), .ZN(new_n15855_));
  AOI21_X1   g15663(.A1(new_n15853_), .A2(new_n15854_), .B(new_n7690_), .ZN(new_n15856_));
  AOI21_X1   g15664(.A1(new_n15657_), .A2(new_n15855_), .B(new_n15856_), .ZN(new_n15857_));
  AOI21_X1   g15665(.A1(new_n15857_), .A2(new_n7331_), .B(new_n15849_), .ZN(new_n15858_));
  NAND2_X1   g15666(.A1(new_n15855_), .A2(new_n15657_), .ZN(new_n15859_));
  AOI21_X1   g15667(.A1(new_n15859_), .A2(new_n15840_), .B(new_n7331_), .ZN(new_n15860_));
  OAI21_X1   g15668(.A1(new_n15858_), .A2(new_n15860_), .B(\asqrt[28] ), .ZN(new_n15861_));
  AOI21_X1   g15669(.A1(new_n15848_), .A2(new_n15861_), .B(new_n6636_), .ZN(new_n15862_));
  NOR3_X1    g15670(.A1(new_n15847_), .A2(\asqrt[30] ), .A3(new_n15862_), .ZN(new_n15863_));
  OAI21_X1   g15671(.A1(new_n15847_), .A2(new_n15862_), .B(\asqrt[30] ), .ZN(new_n15864_));
  OAI21_X1   g15672(.A1(new_n15646_), .A2(new_n15863_), .B(new_n15864_), .ZN(new_n15865_));
  OAI21_X1   g15673(.A1(new_n15865_), .A2(\asqrt[31] ), .B(new_n15643_), .ZN(new_n15866_));
  NAND2_X1   g15674(.A1(new_n15865_), .A2(\asqrt[31] ), .ZN(new_n15867_));
  NAND3_X1   g15675(.A1(new_n15866_), .A2(new_n15867_), .A3(new_n5643_), .ZN(new_n15868_));
  AOI21_X1   g15676(.A1(new_n15866_), .A2(new_n15867_), .B(new_n5643_), .ZN(new_n15869_));
  AOI21_X1   g15677(.A1(new_n15640_), .A2(new_n15868_), .B(new_n15869_), .ZN(new_n15870_));
  AOI21_X1   g15678(.A1(new_n15870_), .A2(new_n5336_), .B(new_n15637_), .ZN(new_n15871_));
  NAND2_X1   g15679(.A1(new_n15868_), .A2(new_n15640_), .ZN(new_n15872_));
  INV_X1     g15680(.I(new_n15643_), .ZN(new_n15873_));
  INV_X1     g15681(.I(new_n15652_), .ZN(new_n15874_));
  NOR3_X1    g15682(.A1(new_n15858_), .A2(\asqrt[28] ), .A3(new_n15860_), .ZN(new_n15875_));
  OAI21_X1   g15683(.A1(new_n15874_), .A2(new_n15875_), .B(new_n15861_), .ZN(new_n15876_));
  OAI21_X1   g15684(.A1(new_n15876_), .A2(\asqrt[29] ), .B(new_n15648_), .ZN(new_n15877_));
  NAND2_X1   g15685(.A1(new_n15876_), .A2(\asqrt[29] ), .ZN(new_n15878_));
  NAND3_X1   g15686(.A1(new_n15877_), .A2(new_n15878_), .A3(new_n6275_), .ZN(new_n15879_));
  AOI21_X1   g15687(.A1(new_n15877_), .A2(new_n15878_), .B(new_n6275_), .ZN(new_n15880_));
  AOI21_X1   g15688(.A1(new_n15645_), .A2(new_n15879_), .B(new_n15880_), .ZN(new_n15881_));
  AOI21_X1   g15689(.A1(new_n15881_), .A2(new_n5947_), .B(new_n15873_), .ZN(new_n15882_));
  NAND2_X1   g15690(.A1(new_n15879_), .A2(new_n15645_), .ZN(new_n15883_));
  AOI21_X1   g15691(.A1(new_n15883_), .A2(new_n15864_), .B(new_n5947_), .ZN(new_n15884_));
  OAI21_X1   g15692(.A1(new_n15882_), .A2(new_n15884_), .B(\asqrt[32] ), .ZN(new_n15885_));
  AOI21_X1   g15693(.A1(new_n15872_), .A2(new_n15885_), .B(new_n5336_), .ZN(new_n15886_));
  NOR3_X1    g15694(.A1(new_n15871_), .A2(\asqrt[34] ), .A3(new_n15886_), .ZN(new_n15887_));
  OAI21_X1   g15695(.A1(new_n15871_), .A2(new_n15886_), .B(\asqrt[34] ), .ZN(new_n15888_));
  OAI21_X1   g15696(.A1(new_n15634_), .A2(new_n15887_), .B(new_n15888_), .ZN(new_n15889_));
  OAI21_X1   g15697(.A1(new_n15889_), .A2(\asqrt[35] ), .B(new_n15631_), .ZN(new_n15890_));
  NAND2_X1   g15698(.A1(new_n15889_), .A2(\asqrt[35] ), .ZN(new_n15891_));
  NAND3_X1   g15699(.A1(new_n15890_), .A2(new_n15891_), .A3(new_n4461_), .ZN(new_n15892_));
  AOI21_X1   g15700(.A1(new_n15890_), .A2(new_n15891_), .B(new_n4461_), .ZN(new_n15893_));
  AOI21_X1   g15701(.A1(new_n15628_), .A2(new_n15892_), .B(new_n15893_), .ZN(new_n15894_));
  AOI21_X1   g15702(.A1(new_n15894_), .A2(new_n4196_), .B(new_n15625_), .ZN(new_n15895_));
  NAND2_X1   g15703(.A1(new_n15892_), .A2(new_n15628_), .ZN(new_n15896_));
  INV_X1     g15704(.I(new_n15631_), .ZN(new_n15897_));
  INV_X1     g15705(.I(new_n15640_), .ZN(new_n15898_));
  NOR3_X1    g15706(.A1(new_n15882_), .A2(\asqrt[32] ), .A3(new_n15884_), .ZN(new_n15899_));
  OAI21_X1   g15707(.A1(new_n15898_), .A2(new_n15899_), .B(new_n15885_), .ZN(new_n15900_));
  OAI21_X1   g15708(.A1(new_n15900_), .A2(\asqrt[33] ), .B(new_n15636_), .ZN(new_n15901_));
  NAND2_X1   g15709(.A1(new_n15900_), .A2(\asqrt[33] ), .ZN(new_n15902_));
  NAND3_X1   g15710(.A1(new_n15901_), .A2(new_n15902_), .A3(new_n5029_), .ZN(new_n15903_));
  AOI21_X1   g15711(.A1(new_n15901_), .A2(new_n15902_), .B(new_n5029_), .ZN(new_n15904_));
  AOI21_X1   g15712(.A1(new_n15633_), .A2(new_n15903_), .B(new_n15904_), .ZN(new_n15905_));
  AOI21_X1   g15713(.A1(new_n15905_), .A2(new_n4751_), .B(new_n15897_), .ZN(new_n15906_));
  NAND2_X1   g15714(.A1(new_n15903_), .A2(new_n15633_), .ZN(new_n15907_));
  AOI21_X1   g15715(.A1(new_n15907_), .A2(new_n15888_), .B(new_n4751_), .ZN(new_n15908_));
  OAI21_X1   g15716(.A1(new_n15906_), .A2(new_n15908_), .B(\asqrt[36] ), .ZN(new_n15909_));
  AOI21_X1   g15717(.A1(new_n15896_), .A2(new_n15909_), .B(new_n4196_), .ZN(new_n15910_));
  NOR3_X1    g15718(.A1(new_n15895_), .A2(\asqrt[38] ), .A3(new_n15910_), .ZN(new_n15911_));
  OAI21_X1   g15719(.A1(new_n15895_), .A2(new_n15910_), .B(\asqrt[38] ), .ZN(new_n15912_));
  OAI21_X1   g15720(.A1(new_n15622_), .A2(new_n15911_), .B(new_n15912_), .ZN(new_n15913_));
  OAI21_X1   g15721(.A1(new_n15913_), .A2(\asqrt[39] ), .B(new_n15619_), .ZN(new_n15914_));
  NAND2_X1   g15722(.A1(new_n15913_), .A2(\asqrt[39] ), .ZN(new_n15915_));
  NAND3_X1   g15723(.A1(new_n15914_), .A2(new_n15915_), .A3(new_n3427_), .ZN(new_n15916_));
  AOI21_X1   g15724(.A1(new_n15914_), .A2(new_n15915_), .B(new_n3427_), .ZN(new_n15917_));
  AOI21_X1   g15725(.A1(new_n15616_), .A2(new_n15916_), .B(new_n15917_), .ZN(new_n15918_));
  AOI21_X1   g15726(.A1(new_n15918_), .A2(new_n3195_), .B(new_n15613_), .ZN(new_n15919_));
  NAND2_X1   g15727(.A1(new_n15916_), .A2(new_n15616_), .ZN(new_n15920_));
  INV_X1     g15728(.I(new_n15619_), .ZN(new_n15921_));
  INV_X1     g15729(.I(new_n15628_), .ZN(new_n15922_));
  NOR3_X1    g15730(.A1(new_n15906_), .A2(\asqrt[36] ), .A3(new_n15908_), .ZN(new_n15923_));
  OAI21_X1   g15731(.A1(new_n15922_), .A2(new_n15923_), .B(new_n15909_), .ZN(new_n15924_));
  OAI21_X1   g15732(.A1(new_n15924_), .A2(\asqrt[37] ), .B(new_n15624_), .ZN(new_n15925_));
  NAND2_X1   g15733(.A1(new_n15924_), .A2(\asqrt[37] ), .ZN(new_n15926_));
  NAND3_X1   g15734(.A1(new_n15925_), .A2(new_n15926_), .A3(new_n3925_), .ZN(new_n15927_));
  AOI21_X1   g15735(.A1(new_n15925_), .A2(new_n15926_), .B(new_n3925_), .ZN(new_n15928_));
  AOI21_X1   g15736(.A1(new_n15621_), .A2(new_n15927_), .B(new_n15928_), .ZN(new_n15929_));
  AOI21_X1   g15737(.A1(new_n15929_), .A2(new_n3681_), .B(new_n15921_), .ZN(new_n15930_));
  NAND2_X1   g15738(.A1(new_n15927_), .A2(new_n15621_), .ZN(new_n15931_));
  AOI21_X1   g15739(.A1(new_n15931_), .A2(new_n15912_), .B(new_n3681_), .ZN(new_n15932_));
  OAI21_X1   g15740(.A1(new_n15930_), .A2(new_n15932_), .B(\asqrt[40] ), .ZN(new_n15933_));
  AOI21_X1   g15741(.A1(new_n15920_), .A2(new_n15933_), .B(new_n3195_), .ZN(new_n15934_));
  NOR3_X1    g15742(.A1(new_n15919_), .A2(\asqrt[42] ), .A3(new_n15934_), .ZN(new_n15935_));
  OAI21_X1   g15743(.A1(new_n15919_), .A2(new_n15934_), .B(\asqrt[42] ), .ZN(new_n15936_));
  OAI21_X1   g15744(.A1(new_n15610_), .A2(new_n15935_), .B(new_n15936_), .ZN(new_n15937_));
  OAI21_X1   g15745(.A1(new_n15937_), .A2(\asqrt[43] ), .B(new_n15607_), .ZN(new_n15938_));
  NAND2_X1   g15746(.A1(new_n15937_), .A2(\asqrt[43] ), .ZN(new_n15939_));
  NAND3_X1   g15747(.A1(new_n15938_), .A2(new_n15939_), .A3(new_n2531_), .ZN(new_n15940_));
  AOI21_X1   g15748(.A1(new_n15938_), .A2(new_n15939_), .B(new_n2531_), .ZN(new_n15941_));
  AOI21_X1   g15749(.A1(new_n15604_), .A2(new_n15940_), .B(new_n15941_), .ZN(new_n15942_));
  AOI21_X1   g15750(.A1(new_n15942_), .A2(new_n2332_), .B(new_n15601_), .ZN(new_n15943_));
  NAND2_X1   g15751(.A1(new_n15940_), .A2(new_n15604_), .ZN(new_n15944_));
  INV_X1     g15752(.I(new_n15607_), .ZN(new_n15945_));
  INV_X1     g15753(.I(new_n15616_), .ZN(new_n15946_));
  NOR3_X1    g15754(.A1(new_n15930_), .A2(\asqrt[40] ), .A3(new_n15932_), .ZN(new_n15947_));
  OAI21_X1   g15755(.A1(new_n15946_), .A2(new_n15947_), .B(new_n15933_), .ZN(new_n15948_));
  OAI21_X1   g15756(.A1(new_n15948_), .A2(\asqrt[41] ), .B(new_n15612_), .ZN(new_n15949_));
  NAND2_X1   g15757(.A1(new_n15948_), .A2(\asqrt[41] ), .ZN(new_n15950_));
  NAND3_X1   g15758(.A1(new_n15949_), .A2(new_n15950_), .A3(new_n2960_), .ZN(new_n15951_));
  AOI21_X1   g15759(.A1(new_n15949_), .A2(new_n15950_), .B(new_n2960_), .ZN(new_n15952_));
  AOI21_X1   g15760(.A1(new_n15609_), .A2(new_n15951_), .B(new_n15952_), .ZN(new_n15953_));
  AOI21_X1   g15761(.A1(new_n15953_), .A2(new_n2749_), .B(new_n15945_), .ZN(new_n15954_));
  NAND2_X1   g15762(.A1(new_n15951_), .A2(new_n15609_), .ZN(new_n15955_));
  AOI21_X1   g15763(.A1(new_n15955_), .A2(new_n15936_), .B(new_n2749_), .ZN(new_n15956_));
  OAI21_X1   g15764(.A1(new_n15954_), .A2(new_n15956_), .B(\asqrt[44] ), .ZN(new_n15957_));
  AOI21_X1   g15765(.A1(new_n15944_), .A2(new_n15957_), .B(new_n2332_), .ZN(new_n15958_));
  NOR3_X1    g15766(.A1(new_n15943_), .A2(\asqrt[46] ), .A3(new_n15958_), .ZN(new_n15959_));
  OAI21_X1   g15767(.A1(new_n15943_), .A2(new_n15958_), .B(\asqrt[46] ), .ZN(new_n15960_));
  OAI21_X1   g15768(.A1(new_n15598_), .A2(new_n15959_), .B(new_n15960_), .ZN(new_n15961_));
  OAI21_X1   g15769(.A1(new_n15961_), .A2(\asqrt[47] ), .B(new_n15595_), .ZN(new_n15962_));
  NAND2_X1   g15770(.A1(new_n15961_), .A2(\asqrt[47] ), .ZN(new_n15963_));
  NAND3_X1   g15771(.A1(new_n15962_), .A2(new_n15963_), .A3(new_n1778_), .ZN(new_n15964_));
  AOI21_X1   g15772(.A1(new_n15962_), .A2(new_n15963_), .B(new_n1778_), .ZN(new_n15965_));
  AOI21_X1   g15773(.A1(new_n15592_), .A2(new_n15964_), .B(new_n15965_), .ZN(new_n15966_));
  AOI21_X1   g15774(.A1(new_n15966_), .A2(new_n1632_), .B(new_n15589_), .ZN(new_n15967_));
  NAND2_X1   g15775(.A1(new_n15964_), .A2(new_n15592_), .ZN(new_n15968_));
  INV_X1     g15776(.I(new_n15595_), .ZN(new_n15969_));
  INV_X1     g15777(.I(new_n15604_), .ZN(new_n15970_));
  NOR3_X1    g15778(.A1(new_n15954_), .A2(\asqrt[44] ), .A3(new_n15956_), .ZN(new_n15971_));
  OAI21_X1   g15779(.A1(new_n15970_), .A2(new_n15971_), .B(new_n15957_), .ZN(new_n15972_));
  OAI21_X1   g15780(.A1(new_n15972_), .A2(\asqrt[45] ), .B(new_n15600_), .ZN(new_n15973_));
  NAND2_X1   g15781(.A1(new_n15972_), .A2(\asqrt[45] ), .ZN(new_n15974_));
  NAND3_X1   g15782(.A1(new_n15973_), .A2(new_n15974_), .A3(new_n2134_), .ZN(new_n15975_));
  AOI21_X1   g15783(.A1(new_n15973_), .A2(new_n15974_), .B(new_n2134_), .ZN(new_n15976_));
  AOI21_X1   g15784(.A1(new_n15597_), .A2(new_n15975_), .B(new_n15976_), .ZN(new_n15977_));
  AOI21_X1   g15785(.A1(new_n15977_), .A2(new_n1953_), .B(new_n15969_), .ZN(new_n15978_));
  NAND2_X1   g15786(.A1(new_n15975_), .A2(new_n15597_), .ZN(new_n15979_));
  AOI21_X1   g15787(.A1(new_n15979_), .A2(new_n15960_), .B(new_n1953_), .ZN(new_n15980_));
  OAI21_X1   g15788(.A1(new_n15978_), .A2(new_n15980_), .B(\asqrt[48] ), .ZN(new_n15981_));
  AOI21_X1   g15789(.A1(new_n15968_), .A2(new_n15981_), .B(new_n1632_), .ZN(new_n15982_));
  NOR3_X1    g15790(.A1(new_n15967_), .A2(\asqrt[50] ), .A3(new_n15982_), .ZN(new_n15983_));
  OAI21_X1   g15791(.A1(new_n15967_), .A2(new_n15982_), .B(\asqrt[50] ), .ZN(new_n15984_));
  OAI21_X1   g15792(.A1(new_n15586_), .A2(new_n15983_), .B(new_n15984_), .ZN(new_n15985_));
  OAI21_X1   g15793(.A1(new_n15985_), .A2(\asqrt[51] ), .B(new_n15583_), .ZN(new_n15986_));
  NAND2_X1   g15794(.A1(new_n15985_), .A2(\asqrt[51] ), .ZN(new_n15987_));
  NAND3_X1   g15795(.A1(new_n15986_), .A2(new_n15987_), .A3(new_n1150_), .ZN(new_n15988_));
  AOI21_X1   g15796(.A1(new_n15986_), .A2(new_n15987_), .B(new_n1150_), .ZN(new_n15989_));
  AOI21_X1   g15797(.A1(new_n15580_), .A2(new_n15988_), .B(new_n15989_), .ZN(new_n15990_));
  AOI21_X1   g15798(.A1(new_n15990_), .A2(new_n1006_), .B(new_n15577_), .ZN(new_n15991_));
  NAND2_X1   g15799(.A1(new_n15988_), .A2(new_n15580_), .ZN(new_n15992_));
  INV_X1     g15800(.I(new_n15583_), .ZN(new_n15993_));
  INV_X1     g15801(.I(new_n15592_), .ZN(new_n15994_));
  NOR3_X1    g15802(.A1(new_n15978_), .A2(\asqrt[48] ), .A3(new_n15980_), .ZN(new_n15995_));
  OAI21_X1   g15803(.A1(new_n15994_), .A2(new_n15995_), .B(new_n15981_), .ZN(new_n15996_));
  OAI21_X1   g15804(.A1(new_n15996_), .A2(\asqrt[49] ), .B(new_n15588_), .ZN(new_n15997_));
  NAND2_X1   g15805(.A1(new_n15996_), .A2(\asqrt[49] ), .ZN(new_n15998_));
  NAND3_X1   g15806(.A1(new_n15997_), .A2(new_n15998_), .A3(new_n1463_), .ZN(new_n15999_));
  AOI21_X1   g15807(.A1(new_n15997_), .A2(new_n15998_), .B(new_n1463_), .ZN(new_n16000_));
  AOI21_X1   g15808(.A1(new_n15585_), .A2(new_n15999_), .B(new_n16000_), .ZN(new_n16001_));
  AOI21_X1   g15809(.A1(new_n16001_), .A2(new_n1305_), .B(new_n15993_), .ZN(new_n16002_));
  NAND2_X1   g15810(.A1(new_n15999_), .A2(new_n15585_), .ZN(new_n16003_));
  AOI21_X1   g15811(.A1(new_n16003_), .A2(new_n15984_), .B(new_n1305_), .ZN(new_n16004_));
  OAI21_X1   g15812(.A1(new_n16002_), .A2(new_n16004_), .B(\asqrt[52] ), .ZN(new_n16005_));
  AOI21_X1   g15813(.A1(new_n15992_), .A2(new_n16005_), .B(new_n1006_), .ZN(new_n16006_));
  NOR3_X1    g15814(.A1(new_n15991_), .A2(\asqrt[54] ), .A3(new_n16006_), .ZN(new_n16007_));
  OAI21_X1   g15815(.A1(new_n15991_), .A2(new_n16006_), .B(\asqrt[54] ), .ZN(new_n16008_));
  OAI21_X1   g15816(.A1(new_n15574_), .A2(new_n16007_), .B(new_n16008_), .ZN(new_n16009_));
  OAI21_X1   g15817(.A1(new_n16009_), .A2(\asqrt[55] ), .B(new_n15571_), .ZN(new_n16010_));
  NAND2_X1   g15818(.A1(new_n16009_), .A2(\asqrt[55] ), .ZN(new_n16011_));
  NAND3_X1   g15819(.A1(new_n16010_), .A2(new_n16011_), .A3(new_n634_), .ZN(new_n16012_));
  AOI21_X1   g15820(.A1(new_n16010_), .A2(new_n16011_), .B(new_n634_), .ZN(new_n16013_));
  AOI21_X1   g15821(.A1(new_n15568_), .A2(new_n16012_), .B(new_n16013_), .ZN(new_n16014_));
  NAND2_X1   g15822(.A1(new_n16014_), .A2(new_n531_), .ZN(new_n16015_));
  INV_X1     g15823(.I(new_n15568_), .ZN(new_n16016_));
  INV_X1     g15824(.I(new_n15571_), .ZN(new_n16017_));
  INV_X1     g15825(.I(new_n15580_), .ZN(new_n16018_));
  NOR3_X1    g15826(.A1(new_n16002_), .A2(\asqrt[52] ), .A3(new_n16004_), .ZN(new_n16019_));
  OAI21_X1   g15827(.A1(new_n16018_), .A2(new_n16019_), .B(new_n16005_), .ZN(new_n16020_));
  OAI21_X1   g15828(.A1(new_n16020_), .A2(\asqrt[53] ), .B(new_n15576_), .ZN(new_n16021_));
  NAND2_X1   g15829(.A1(new_n16020_), .A2(\asqrt[53] ), .ZN(new_n16022_));
  NAND3_X1   g15830(.A1(new_n16021_), .A2(new_n16022_), .A3(new_n860_), .ZN(new_n16023_));
  AOI21_X1   g15831(.A1(new_n16021_), .A2(new_n16022_), .B(new_n860_), .ZN(new_n16024_));
  AOI21_X1   g15832(.A1(new_n15573_), .A2(new_n16023_), .B(new_n16024_), .ZN(new_n16025_));
  AOI21_X1   g15833(.A1(new_n16025_), .A2(new_n744_), .B(new_n16017_), .ZN(new_n16026_));
  NAND2_X1   g15834(.A1(new_n16023_), .A2(new_n15573_), .ZN(new_n16027_));
  AOI21_X1   g15835(.A1(new_n16027_), .A2(new_n16008_), .B(new_n744_), .ZN(new_n16028_));
  NOR3_X1    g15836(.A1(new_n16026_), .A2(\asqrt[56] ), .A3(new_n16028_), .ZN(new_n16029_));
  NOR2_X1    g15837(.A1(new_n16029_), .A2(new_n16016_), .ZN(new_n16030_));
  OAI21_X1   g15838(.A1(new_n16030_), .A2(new_n16013_), .B(\asqrt[57] ), .ZN(new_n16031_));
  NOR2_X1    g15839(.A1(new_n15536_), .A2(\asqrt[62] ), .ZN(new_n16032_));
  INV_X1     g15840(.I(new_n15553_), .ZN(new_n16033_));
  NOR2_X1    g15841(.A1(new_n16033_), .A2(new_n16032_), .ZN(new_n16034_));
  XOR2_X1    g15842(.A1(new_n15544_), .A2(new_n15036_), .Z(new_n16035_));
  OAI21_X1   g15843(.A1(\asqrt[8] ), .A2(new_n16034_), .B(new_n16035_), .ZN(new_n16036_));
  INV_X1     g15844(.I(new_n16036_), .ZN(new_n16037_));
  NOR2_X1    g15845(.A1(new_n15516_), .A2(new_n15513_), .ZN(new_n16038_));
  NOR2_X1    g15846(.A1(\asqrt[8] ), .A2(new_n16038_), .ZN(new_n16039_));
  XOR2_X1    g15847(.A1(new_n16039_), .A2(new_n15497_), .Z(new_n16040_));
  INV_X1     g15848(.I(new_n16040_), .ZN(new_n16041_));
  NOR2_X1    g15849(.A1(new_n15523_), .A2(new_n15512_), .ZN(new_n16042_));
  NOR2_X1    g15850(.A1(\asqrt[8] ), .A2(new_n16042_), .ZN(new_n16043_));
  XOR2_X1    g15851(.A1(new_n16043_), .A2(new_n15501_), .Z(new_n16044_));
  AOI21_X1   g15852(.A1(new_n15506_), .A2(new_n15511_), .B(\asqrt[8] ), .ZN(new_n16045_));
  XOR2_X1    g15853(.A1(new_n16045_), .A2(new_n15504_), .Z(new_n16046_));
  OAI21_X1   g15854(.A1(new_n16026_), .A2(new_n16028_), .B(\asqrt[56] ), .ZN(new_n16047_));
  OAI21_X1   g15855(.A1(new_n16016_), .A2(new_n16029_), .B(new_n16047_), .ZN(new_n16048_));
  OAI21_X1   g15856(.A1(new_n16048_), .A2(\asqrt[57] ), .B(new_n15564_), .ZN(new_n16049_));
  NAND3_X1   g15857(.A1(new_n16049_), .A2(new_n423_), .A3(new_n16031_), .ZN(new_n16050_));
  NAND2_X1   g15858(.A1(new_n16050_), .A2(new_n16046_), .ZN(new_n16051_));
  INV_X1     g15859(.I(new_n15564_), .ZN(new_n16052_));
  AOI21_X1   g15860(.A1(new_n16014_), .A2(new_n531_), .B(new_n16052_), .ZN(new_n16053_));
  NAND2_X1   g15861(.A1(new_n16012_), .A2(new_n15568_), .ZN(new_n16054_));
  AOI21_X1   g15862(.A1(new_n16054_), .A2(new_n16047_), .B(new_n531_), .ZN(new_n16055_));
  OAI21_X1   g15863(.A1(new_n16053_), .A2(new_n16055_), .B(\asqrt[58] ), .ZN(new_n16056_));
  NAND3_X1   g15864(.A1(new_n16051_), .A2(new_n337_), .A3(new_n16056_), .ZN(new_n16057_));
  AOI21_X1   g15865(.A1(new_n16051_), .A2(new_n16056_), .B(new_n337_), .ZN(new_n16058_));
  AOI21_X1   g15866(.A1(new_n16044_), .A2(new_n16057_), .B(new_n16058_), .ZN(new_n16059_));
  AOI21_X1   g15867(.A1(new_n16059_), .A2(new_n266_), .B(new_n16041_), .ZN(new_n16060_));
  INV_X1     g15868(.I(new_n16046_), .ZN(new_n16061_));
  NOR3_X1    g15869(.A1(new_n16053_), .A2(\asqrt[58] ), .A3(new_n16055_), .ZN(new_n16062_));
  OAI21_X1   g15870(.A1(new_n16061_), .A2(new_n16062_), .B(new_n16056_), .ZN(new_n16063_));
  OAI21_X1   g15871(.A1(new_n16063_), .A2(\asqrt[59] ), .B(new_n16044_), .ZN(new_n16064_));
  NAND2_X1   g15872(.A1(new_n16063_), .A2(\asqrt[59] ), .ZN(new_n16065_));
  AOI21_X1   g15873(.A1(new_n16064_), .A2(new_n16065_), .B(new_n266_), .ZN(new_n16066_));
  OAI21_X1   g15874(.A1(new_n16060_), .A2(new_n16066_), .B(\asqrt[61] ), .ZN(new_n16067_));
  AOI21_X1   g15875(.A1(new_n15538_), .A2(new_n15533_), .B(\asqrt[8] ), .ZN(new_n16068_));
  XOR2_X1    g15876(.A1(new_n16068_), .A2(new_n15494_), .Z(new_n16069_));
  INV_X1     g15877(.I(new_n16069_), .ZN(new_n16070_));
  NOR3_X1    g15878(.A1(new_n16060_), .A2(\asqrt[61] ), .A3(new_n16066_), .ZN(new_n16071_));
  OAI21_X1   g15879(.A1(new_n16070_), .A2(new_n16071_), .B(new_n16067_), .ZN(new_n16072_));
  NAND3_X1   g15880(.A1(new_n16064_), .A2(new_n16065_), .A3(new_n266_), .ZN(new_n16073_));
  NAND2_X1   g15881(.A1(new_n16073_), .A2(new_n16040_), .ZN(new_n16074_));
  INV_X1     g15882(.I(new_n16044_), .ZN(new_n16075_));
  AOI21_X1   g15883(.A1(new_n16049_), .A2(new_n16031_), .B(new_n423_), .ZN(new_n16076_));
  AOI21_X1   g15884(.A1(new_n16046_), .A2(new_n16050_), .B(new_n16076_), .ZN(new_n16077_));
  AOI21_X1   g15885(.A1(new_n16077_), .A2(new_n337_), .B(new_n16075_), .ZN(new_n16078_));
  OAI21_X1   g15886(.A1(new_n16078_), .A2(new_n16058_), .B(\asqrt[60] ), .ZN(new_n16079_));
  AOI21_X1   g15887(.A1(new_n16074_), .A2(new_n16079_), .B(new_n239_), .ZN(new_n16080_));
  AOI21_X1   g15888(.A1(new_n16040_), .A2(new_n16073_), .B(new_n16066_), .ZN(new_n16081_));
  AOI21_X1   g15889(.A1(new_n16081_), .A2(new_n239_), .B(new_n16070_), .ZN(new_n16082_));
  OAI21_X1   g15890(.A1(new_n16082_), .A2(new_n16080_), .B(new_n201_), .ZN(new_n16083_));
  NOR3_X1    g15891(.A1(new_n16078_), .A2(\asqrt[60] ), .A3(new_n16058_), .ZN(new_n16084_));
  OAI21_X1   g15892(.A1(new_n16041_), .A2(new_n16084_), .B(new_n16079_), .ZN(new_n16085_));
  OAI21_X1   g15893(.A1(new_n16085_), .A2(\asqrt[61] ), .B(new_n16069_), .ZN(new_n16086_));
  NAND3_X1   g15894(.A1(new_n16086_), .A2(\asqrt[62] ), .A3(new_n16067_), .ZN(new_n16087_));
  AOI21_X1   g15895(.A1(new_n15528_), .A2(new_n15534_), .B(\asqrt[8] ), .ZN(new_n16088_));
  XOR2_X1    g15896(.A1(new_n16088_), .A2(new_n15530_), .Z(new_n16089_));
  INV_X1     g15897(.I(new_n16089_), .ZN(new_n16090_));
  AOI22_X1   g15898(.A1(new_n16087_), .A2(new_n16083_), .B1(new_n16072_), .B2(new_n16090_), .ZN(new_n16091_));
  NOR2_X1    g15899(.A1(new_n15547_), .A2(new_n15491_), .ZN(new_n16092_));
  OAI21_X1   g15900(.A1(\asqrt[8] ), .A2(new_n16092_), .B(new_n15554_), .ZN(new_n16093_));
  INV_X1     g15901(.I(new_n16093_), .ZN(new_n16094_));
  OAI21_X1   g15902(.A1(new_n16091_), .A2(new_n16037_), .B(new_n16094_), .ZN(new_n16095_));
  OAI21_X1   g15903(.A1(new_n16072_), .A2(\asqrt[62] ), .B(new_n16089_), .ZN(new_n16096_));
  NAND2_X1   g15904(.A1(new_n16072_), .A2(\asqrt[62] ), .ZN(new_n16097_));
  NAND3_X1   g15905(.A1(new_n16096_), .A2(new_n16097_), .A3(new_n16037_), .ZN(new_n16098_));
  NAND2_X1   g15906(.A1(new_n15717_), .A2(new_n15490_), .ZN(new_n16099_));
  XOR2_X1    g15907(.A1(new_n15547_), .A2(new_n15491_), .Z(new_n16100_));
  NAND3_X1   g15908(.A1(new_n16099_), .A2(\asqrt[63] ), .A3(new_n16100_), .ZN(new_n16101_));
  INV_X1     g15909(.I(new_n15706_), .ZN(new_n16102_));
  NAND4_X1   g15910(.A1(new_n16102_), .A2(new_n15491_), .A3(new_n15554_), .A4(new_n15561_), .ZN(new_n16103_));
  NAND2_X1   g15911(.A1(new_n16101_), .A2(new_n16103_), .ZN(new_n16104_));
  INV_X1     g15912(.I(new_n16104_), .ZN(new_n16105_));
  NAND4_X1   g15913(.A1(new_n16095_), .A2(new_n193_), .A3(new_n16098_), .A4(new_n16105_), .ZN(\asqrt[7] ));
  AOI21_X1   g15914(.A1(new_n16015_), .A2(new_n16031_), .B(\asqrt[7] ), .ZN(new_n16107_));
  XOR2_X1    g15915(.A1(new_n16107_), .A2(new_n15564_), .Z(new_n16108_));
  AOI21_X1   g15916(.A1(new_n16012_), .A2(new_n16047_), .B(\asqrt[7] ), .ZN(new_n16109_));
  XOR2_X1    g15917(.A1(new_n16109_), .A2(new_n15568_), .Z(new_n16110_));
  NAND2_X1   g15918(.A1(new_n16025_), .A2(new_n744_), .ZN(new_n16111_));
  AOI21_X1   g15919(.A1(new_n16111_), .A2(new_n16011_), .B(\asqrt[7] ), .ZN(new_n16112_));
  XOR2_X1    g15920(.A1(new_n16112_), .A2(new_n15571_), .Z(new_n16113_));
  INV_X1     g15921(.I(new_n16113_), .ZN(new_n16114_));
  AOI21_X1   g15922(.A1(new_n16023_), .A2(new_n16008_), .B(\asqrt[7] ), .ZN(new_n16115_));
  XOR2_X1    g15923(.A1(new_n16115_), .A2(new_n15573_), .Z(new_n16116_));
  INV_X1     g15924(.I(new_n16116_), .ZN(new_n16117_));
  NAND2_X1   g15925(.A1(new_n15990_), .A2(new_n1006_), .ZN(new_n16118_));
  AOI21_X1   g15926(.A1(new_n16118_), .A2(new_n16022_), .B(\asqrt[7] ), .ZN(new_n16119_));
  XOR2_X1    g15927(.A1(new_n16119_), .A2(new_n15576_), .Z(new_n16120_));
  AOI21_X1   g15928(.A1(new_n15988_), .A2(new_n16005_), .B(\asqrt[7] ), .ZN(new_n16121_));
  XOR2_X1    g15929(.A1(new_n16121_), .A2(new_n15580_), .Z(new_n16122_));
  NAND2_X1   g15930(.A1(new_n16001_), .A2(new_n1305_), .ZN(new_n16123_));
  AOI21_X1   g15931(.A1(new_n16123_), .A2(new_n15987_), .B(\asqrt[7] ), .ZN(new_n16124_));
  XOR2_X1    g15932(.A1(new_n16124_), .A2(new_n15583_), .Z(new_n16125_));
  INV_X1     g15933(.I(new_n16125_), .ZN(new_n16126_));
  AOI21_X1   g15934(.A1(new_n15999_), .A2(new_n15984_), .B(\asqrt[7] ), .ZN(new_n16127_));
  XOR2_X1    g15935(.A1(new_n16127_), .A2(new_n15585_), .Z(new_n16128_));
  INV_X1     g15936(.I(new_n16128_), .ZN(new_n16129_));
  NAND2_X1   g15937(.A1(new_n15966_), .A2(new_n1632_), .ZN(new_n16130_));
  AOI21_X1   g15938(.A1(new_n16130_), .A2(new_n15998_), .B(\asqrt[7] ), .ZN(new_n16131_));
  XOR2_X1    g15939(.A1(new_n16131_), .A2(new_n15588_), .Z(new_n16132_));
  AOI21_X1   g15940(.A1(new_n15964_), .A2(new_n15981_), .B(\asqrt[7] ), .ZN(new_n16133_));
  XOR2_X1    g15941(.A1(new_n16133_), .A2(new_n15592_), .Z(new_n16134_));
  NAND2_X1   g15942(.A1(new_n15977_), .A2(new_n1953_), .ZN(new_n16135_));
  AOI21_X1   g15943(.A1(new_n16135_), .A2(new_n15963_), .B(\asqrt[7] ), .ZN(new_n16136_));
  XOR2_X1    g15944(.A1(new_n16136_), .A2(new_n15595_), .Z(new_n16137_));
  INV_X1     g15945(.I(new_n16137_), .ZN(new_n16138_));
  AOI21_X1   g15946(.A1(new_n15975_), .A2(new_n15960_), .B(\asqrt[7] ), .ZN(new_n16139_));
  XOR2_X1    g15947(.A1(new_n16139_), .A2(new_n15597_), .Z(new_n16140_));
  INV_X1     g15948(.I(new_n16140_), .ZN(new_n16141_));
  NAND2_X1   g15949(.A1(new_n15942_), .A2(new_n2332_), .ZN(new_n16142_));
  AOI21_X1   g15950(.A1(new_n16142_), .A2(new_n15974_), .B(\asqrt[7] ), .ZN(new_n16143_));
  XOR2_X1    g15951(.A1(new_n16143_), .A2(new_n15600_), .Z(new_n16144_));
  AOI21_X1   g15952(.A1(new_n15940_), .A2(new_n15957_), .B(\asqrt[7] ), .ZN(new_n16145_));
  XOR2_X1    g15953(.A1(new_n16145_), .A2(new_n15604_), .Z(new_n16146_));
  NAND2_X1   g15954(.A1(new_n15953_), .A2(new_n2749_), .ZN(new_n16147_));
  AOI21_X1   g15955(.A1(new_n16147_), .A2(new_n15939_), .B(\asqrt[7] ), .ZN(new_n16148_));
  XOR2_X1    g15956(.A1(new_n16148_), .A2(new_n15607_), .Z(new_n16149_));
  INV_X1     g15957(.I(new_n16149_), .ZN(new_n16150_));
  AOI21_X1   g15958(.A1(new_n15951_), .A2(new_n15936_), .B(\asqrt[7] ), .ZN(new_n16151_));
  XOR2_X1    g15959(.A1(new_n16151_), .A2(new_n15609_), .Z(new_n16152_));
  INV_X1     g15960(.I(new_n16152_), .ZN(new_n16153_));
  NAND2_X1   g15961(.A1(new_n15918_), .A2(new_n3195_), .ZN(new_n16154_));
  AOI21_X1   g15962(.A1(new_n16154_), .A2(new_n15950_), .B(\asqrt[7] ), .ZN(new_n16155_));
  XOR2_X1    g15963(.A1(new_n16155_), .A2(new_n15612_), .Z(new_n16156_));
  AOI21_X1   g15964(.A1(new_n15916_), .A2(new_n15933_), .B(\asqrt[7] ), .ZN(new_n16157_));
  XOR2_X1    g15965(.A1(new_n16157_), .A2(new_n15616_), .Z(new_n16158_));
  NAND2_X1   g15966(.A1(new_n15929_), .A2(new_n3681_), .ZN(new_n16159_));
  AOI21_X1   g15967(.A1(new_n16159_), .A2(new_n15915_), .B(\asqrt[7] ), .ZN(new_n16160_));
  XOR2_X1    g15968(.A1(new_n16160_), .A2(new_n15619_), .Z(new_n16161_));
  INV_X1     g15969(.I(new_n16161_), .ZN(new_n16162_));
  AOI21_X1   g15970(.A1(new_n15927_), .A2(new_n15912_), .B(\asqrt[7] ), .ZN(new_n16163_));
  XOR2_X1    g15971(.A1(new_n16163_), .A2(new_n15621_), .Z(new_n16164_));
  INV_X1     g15972(.I(new_n16164_), .ZN(new_n16165_));
  NAND2_X1   g15973(.A1(new_n15894_), .A2(new_n4196_), .ZN(new_n16166_));
  AOI21_X1   g15974(.A1(new_n16166_), .A2(new_n15926_), .B(\asqrt[7] ), .ZN(new_n16167_));
  XOR2_X1    g15975(.A1(new_n16167_), .A2(new_n15624_), .Z(new_n16168_));
  AOI21_X1   g15976(.A1(new_n15892_), .A2(new_n15909_), .B(\asqrt[7] ), .ZN(new_n16169_));
  XOR2_X1    g15977(.A1(new_n16169_), .A2(new_n15628_), .Z(new_n16170_));
  NAND2_X1   g15978(.A1(new_n15905_), .A2(new_n4751_), .ZN(new_n16171_));
  AOI21_X1   g15979(.A1(new_n16171_), .A2(new_n15891_), .B(\asqrt[7] ), .ZN(new_n16172_));
  XOR2_X1    g15980(.A1(new_n16172_), .A2(new_n15631_), .Z(new_n16173_));
  INV_X1     g15981(.I(new_n16173_), .ZN(new_n16174_));
  AOI21_X1   g15982(.A1(new_n15903_), .A2(new_n15888_), .B(\asqrt[7] ), .ZN(new_n16175_));
  XOR2_X1    g15983(.A1(new_n16175_), .A2(new_n15633_), .Z(new_n16176_));
  INV_X1     g15984(.I(new_n16176_), .ZN(new_n16177_));
  NAND2_X1   g15985(.A1(new_n15870_), .A2(new_n5336_), .ZN(new_n16178_));
  AOI21_X1   g15986(.A1(new_n16178_), .A2(new_n15902_), .B(\asqrt[7] ), .ZN(new_n16179_));
  XOR2_X1    g15987(.A1(new_n16179_), .A2(new_n15636_), .Z(new_n16180_));
  AOI21_X1   g15988(.A1(new_n15868_), .A2(new_n15885_), .B(\asqrt[7] ), .ZN(new_n16181_));
  XOR2_X1    g15989(.A1(new_n16181_), .A2(new_n15640_), .Z(new_n16182_));
  NAND2_X1   g15990(.A1(new_n15881_), .A2(new_n5947_), .ZN(new_n16183_));
  AOI21_X1   g15991(.A1(new_n16183_), .A2(new_n15867_), .B(\asqrt[7] ), .ZN(new_n16184_));
  XOR2_X1    g15992(.A1(new_n16184_), .A2(new_n15643_), .Z(new_n16185_));
  INV_X1     g15993(.I(new_n16185_), .ZN(new_n16186_));
  AOI21_X1   g15994(.A1(new_n15879_), .A2(new_n15864_), .B(\asqrt[7] ), .ZN(new_n16187_));
  XOR2_X1    g15995(.A1(new_n16187_), .A2(new_n15645_), .Z(new_n16188_));
  INV_X1     g15996(.I(new_n16188_), .ZN(new_n16189_));
  NAND2_X1   g15997(.A1(new_n15846_), .A2(new_n6636_), .ZN(new_n16190_));
  AOI21_X1   g15998(.A1(new_n16190_), .A2(new_n15878_), .B(\asqrt[7] ), .ZN(new_n16191_));
  XOR2_X1    g15999(.A1(new_n16191_), .A2(new_n15648_), .Z(new_n16192_));
  AOI21_X1   g16000(.A1(new_n15844_), .A2(new_n15861_), .B(\asqrt[7] ), .ZN(new_n16193_));
  XOR2_X1    g16001(.A1(new_n16193_), .A2(new_n15652_), .Z(new_n16194_));
  NAND2_X1   g16002(.A1(new_n15857_), .A2(new_n7331_), .ZN(new_n16195_));
  AOI21_X1   g16003(.A1(new_n16195_), .A2(new_n15843_), .B(\asqrt[7] ), .ZN(new_n16196_));
  XOR2_X1    g16004(.A1(new_n16196_), .A2(new_n15655_), .Z(new_n16197_));
  INV_X1     g16005(.I(new_n16197_), .ZN(new_n16198_));
  AOI21_X1   g16006(.A1(new_n15855_), .A2(new_n15840_), .B(\asqrt[7] ), .ZN(new_n16199_));
  XOR2_X1    g16007(.A1(new_n16199_), .A2(new_n15657_), .Z(new_n16200_));
  INV_X1     g16008(.I(new_n16200_), .ZN(new_n16201_));
  NAND2_X1   g16009(.A1(new_n15822_), .A2(new_n8077_), .ZN(new_n16202_));
  AOI21_X1   g16010(.A1(new_n16202_), .A2(new_n15854_), .B(\asqrt[7] ), .ZN(new_n16203_));
  XOR2_X1    g16011(.A1(new_n16203_), .A2(new_n15660_), .Z(new_n16204_));
  AOI21_X1   g16012(.A1(new_n15820_), .A2(new_n15837_), .B(\asqrt[7] ), .ZN(new_n16205_));
  XOR2_X1    g16013(.A1(new_n16205_), .A2(new_n15664_), .Z(new_n16206_));
  NAND2_X1   g16014(.A1(new_n15833_), .A2(new_n8849_), .ZN(new_n16207_));
  AOI21_X1   g16015(.A1(new_n16207_), .A2(new_n15819_), .B(\asqrt[7] ), .ZN(new_n16208_));
  XOR2_X1    g16016(.A1(new_n16208_), .A2(new_n15667_), .Z(new_n16209_));
  INV_X1     g16017(.I(new_n16209_), .ZN(new_n16210_));
  AOI21_X1   g16018(.A1(new_n15831_), .A2(new_n15816_), .B(\asqrt[7] ), .ZN(new_n16211_));
  XOR2_X1    g16019(.A1(new_n16211_), .A2(new_n15669_), .Z(new_n16212_));
  INV_X1     g16020(.I(new_n16212_), .ZN(new_n16213_));
  NAND2_X1   g16021(.A1(new_n15798_), .A2(new_n9656_), .ZN(new_n16214_));
  AOI21_X1   g16022(.A1(new_n16214_), .A2(new_n15830_), .B(\asqrt[7] ), .ZN(new_n16215_));
  XOR2_X1    g16023(.A1(new_n16215_), .A2(new_n15672_), .Z(new_n16216_));
  AOI21_X1   g16024(.A1(new_n15796_), .A2(new_n15813_), .B(\asqrt[7] ), .ZN(new_n16217_));
  XOR2_X1    g16025(.A1(new_n16217_), .A2(new_n15676_), .Z(new_n16218_));
  NAND2_X1   g16026(.A1(new_n15809_), .A2(new_n10497_), .ZN(new_n16219_));
  AOI21_X1   g16027(.A1(new_n16219_), .A2(new_n15795_), .B(\asqrt[7] ), .ZN(new_n16220_));
  XOR2_X1    g16028(.A1(new_n16220_), .A2(new_n15679_), .Z(new_n16221_));
  INV_X1     g16029(.I(new_n16221_), .ZN(new_n16222_));
  AOI21_X1   g16030(.A1(new_n15807_), .A2(new_n15792_), .B(\asqrt[7] ), .ZN(new_n16223_));
  XOR2_X1    g16031(.A1(new_n16223_), .A2(new_n15681_), .Z(new_n16224_));
  INV_X1     g16032(.I(new_n16224_), .ZN(new_n16225_));
  NAND2_X1   g16033(.A1(new_n15774_), .A2(new_n11373_), .ZN(new_n16226_));
  AOI21_X1   g16034(.A1(new_n16226_), .A2(new_n15806_), .B(\asqrt[7] ), .ZN(new_n16227_));
  XOR2_X1    g16035(.A1(new_n16227_), .A2(new_n15684_), .Z(new_n16228_));
  AOI21_X1   g16036(.A1(new_n15772_), .A2(new_n15789_), .B(\asqrt[7] ), .ZN(new_n16229_));
  XOR2_X1    g16037(.A1(new_n16229_), .A2(new_n15688_), .Z(new_n16230_));
  NAND2_X1   g16038(.A1(new_n15785_), .A2(new_n12283_), .ZN(new_n16231_));
  AOI21_X1   g16039(.A1(new_n16231_), .A2(new_n15771_), .B(\asqrt[7] ), .ZN(new_n16232_));
  XOR2_X1    g16040(.A1(new_n16232_), .A2(new_n15691_), .Z(new_n16233_));
  INV_X1     g16041(.I(new_n16233_), .ZN(new_n16234_));
  AOI21_X1   g16042(.A1(new_n15783_), .A2(new_n15768_), .B(\asqrt[7] ), .ZN(new_n16235_));
  XOR2_X1    g16043(.A1(new_n16235_), .A2(new_n15693_), .Z(new_n16236_));
  INV_X1     g16044(.I(new_n16236_), .ZN(new_n16237_));
  NAND2_X1   g16045(.A1(new_n15746_), .A2(new_n13228_), .ZN(new_n16238_));
  AOI21_X1   g16046(.A1(new_n16238_), .A2(new_n15782_), .B(\asqrt[7] ), .ZN(new_n16239_));
  XOR2_X1    g16047(.A1(new_n16239_), .A2(new_n15696_), .Z(new_n16240_));
  AOI21_X1   g16048(.A1(new_n15744_), .A2(new_n15765_), .B(\asqrt[7] ), .ZN(new_n16241_));
  XOR2_X1    g16049(.A1(new_n16241_), .A2(new_n15699_), .Z(new_n16242_));
  NAND2_X1   g16050(.A1(new_n15761_), .A2(new_n14207_), .ZN(new_n16243_));
  AOI21_X1   g16051(.A1(new_n16243_), .A2(new_n15743_), .B(\asqrt[7] ), .ZN(new_n16244_));
  XOR2_X1    g16052(.A1(new_n16244_), .A2(new_n15705_), .Z(new_n16245_));
  INV_X1     g16053(.I(new_n16245_), .ZN(new_n16246_));
  AOI21_X1   g16054(.A1(new_n15759_), .A2(new_n15740_), .B(\asqrt[7] ), .ZN(new_n16247_));
  XOR2_X1    g16055(.A1(new_n16247_), .A2(new_n15750_), .Z(new_n16248_));
  INV_X1     g16056(.I(new_n16248_), .ZN(new_n16249_));
  NAND2_X1   g16057(.A1(\asqrt[8] ), .A2(new_n15728_), .ZN(new_n16250_));
  NOR2_X1    g16058(.A1(new_n15735_), .A2(\a[16] ), .ZN(new_n16251_));
  AOI22_X1   g16059(.A1(new_n16250_), .A2(new_n15735_), .B1(\asqrt[8] ), .B2(new_n16251_), .ZN(new_n16252_));
  OAI21_X1   g16060(.A1(new_n15717_), .A2(new_n15728_), .B(new_n15754_), .ZN(new_n16253_));
  AOI21_X1   g16061(.A1(new_n15753_), .A2(new_n16253_), .B(\asqrt[7] ), .ZN(new_n16254_));
  XOR2_X1    g16062(.A1(new_n16254_), .A2(new_n16252_), .Z(new_n16255_));
  NOR2_X1    g16063(.A1(new_n16082_), .A2(new_n16080_), .ZN(new_n16256_));
  AOI21_X1   g16064(.A1(new_n16086_), .A2(new_n16067_), .B(\asqrt[62] ), .ZN(new_n16257_));
  NOR3_X1    g16065(.A1(new_n16082_), .A2(new_n201_), .A3(new_n16080_), .ZN(new_n16258_));
  OAI22_X1   g16066(.A1(new_n16257_), .A2(new_n16258_), .B1(new_n16256_), .B2(new_n16089_), .ZN(new_n16259_));
  AOI21_X1   g16067(.A1(new_n16259_), .A2(new_n16036_), .B(new_n16093_), .ZN(new_n16260_));
  AOI21_X1   g16068(.A1(new_n16256_), .A2(new_n201_), .B(new_n16090_), .ZN(new_n16261_));
  NOR2_X1    g16069(.A1(new_n16256_), .A2(new_n201_), .ZN(new_n16262_));
  NOR3_X1    g16070(.A1(new_n16261_), .A2(new_n16262_), .A3(new_n16036_), .ZN(new_n16263_));
  NAND3_X1   g16071(.A1(new_n16101_), .A2(\asqrt[8] ), .A3(new_n16103_), .ZN(new_n16264_));
  NOR4_X1    g16072(.A1(new_n16260_), .A2(\asqrt[63] ), .A3(new_n16263_), .A4(new_n16264_), .ZN(new_n16265_));
  INV_X1     g16073(.I(new_n16265_), .ZN(new_n16266_));
  NAND2_X1   g16074(.A1(\asqrt[7] ), .A2(new_n15725_), .ZN(new_n16267_));
  AOI21_X1   g16075(.A1(new_n16267_), .A2(new_n16266_), .B(\a[16] ), .ZN(new_n16268_));
  NOR4_X1    g16076(.A1(new_n16260_), .A2(\asqrt[63] ), .A3(new_n16263_), .A4(new_n16104_), .ZN(new_n16269_));
  NOR2_X1    g16077(.A1(new_n16269_), .A2(new_n15726_), .ZN(new_n16270_));
  NOR3_X1    g16078(.A1(new_n16270_), .A2(new_n15728_), .A3(new_n16265_), .ZN(new_n16271_));
  NOR2_X1    g16079(.A1(new_n16271_), .A2(new_n16268_), .ZN(new_n16272_));
  INV_X1     g16080(.I(\a[14] ), .ZN(new_n16273_));
  NOR2_X1    g16081(.A1(\a[12] ), .A2(\a[13] ), .ZN(new_n16274_));
  NOR3_X1    g16082(.A1(new_n16269_), .A2(new_n16273_), .A3(new_n16274_), .ZN(new_n16275_));
  INV_X1     g16083(.I(new_n16274_), .ZN(new_n16276_));
  AOI21_X1   g16084(.A1(new_n16269_), .A2(\a[14] ), .B(new_n16276_), .ZN(new_n16277_));
  OAI21_X1   g16085(.A1(new_n16275_), .A2(new_n16277_), .B(\asqrt[8] ), .ZN(new_n16278_));
  NAND2_X1   g16086(.A1(new_n16274_), .A2(new_n16273_), .ZN(new_n16279_));
  NAND3_X1   g16087(.A1(new_n15557_), .A2(new_n15559_), .A3(new_n16279_), .ZN(new_n16280_));
  NAND2_X1   g16088(.A1(new_n15720_), .A2(new_n16280_), .ZN(new_n16281_));
  NAND3_X1   g16089(.A1(\asqrt[7] ), .A2(\a[14] ), .A3(new_n16281_), .ZN(new_n16282_));
  NOR3_X1    g16090(.A1(new_n16269_), .A2(\a[14] ), .A3(\a[15] ), .ZN(new_n16283_));
  INV_X1     g16091(.I(\a[15] ), .ZN(new_n16284_));
  AOI21_X1   g16092(.A1(\asqrt[7] ), .A2(new_n16273_), .B(new_n16284_), .ZN(new_n16285_));
  NOR2_X1    g16093(.A1(new_n16283_), .A2(new_n16285_), .ZN(new_n16286_));
  NAND4_X1   g16094(.A1(new_n16278_), .A2(new_n16286_), .A3(new_n15221_), .A4(new_n16282_), .ZN(new_n16287_));
  NAND2_X1   g16095(.A1(new_n16287_), .A2(new_n16272_), .ZN(new_n16288_));
  NAND3_X1   g16096(.A1(\asqrt[7] ), .A2(\a[14] ), .A3(new_n16276_), .ZN(new_n16289_));
  OAI21_X1   g16097(.A1(\asqrt[7] ), .A2(new_n16273_), .B(new_n16274_), .ZN(new_n16290_));
  AOI21_X1   g16098(.A1(new_n16290_), .A2(new_n16289_), .B(new_n15717_), .ZN(new_n16291_));
  NAND3_X1   g16099(.A1(\asqrt[7] ), .A2(new_n16273_), .A3(new_n16284_), .ZN(new_n16292_));
  OAI21_X1   g16100(.A1(new_n16269_), .A2(\a[14] ), .B(\a[15] ), .ZN(new_n16293_));
  NAND3_X1   g16101(.A1(new_n16282_), .A2(new_n16293_), .A3(new_n16292_), .ZN(new_n16294_));
  OAI21_X1   g16102(.A1(new_n16294_), .A2(new_n16291_), .B(\asqrt[9] ), .ZN(new_n16295_));
  NAND3_X1   g16103(.A1(new_n16288_), .A2(new_n14690_), .A3(new_n16295_), .ZN(new_n16296_));
  AOI21_X1   g16104(.A1(new_n16288_), .A2(new_n16295_), .B(new_n14690_), .ZN(new_n16297_));
  AOI21_X1   g16105(.A1(new_n16255_), .A2(new_n16296_), .B(new_n16297_), .ZN(new_n16298_));
  AOI21_X1   g16106(.A1(new_n16298_), .A2(new_n14207_), .B(new_n16249_), .ZN(new_n16299_));
  OR2_X2     g16107(.A1(new_n16271_), .A2(new_n16268_), .Z(new_n16300_));
  NOR3_X1    g16108(.A1(new_n16294_), .A2(new_n16291_), .A3(\asqrt[9] ), .ZN(new_n16301_));
  OAI21_X1   g16109(.A1(new_n16300_), .A2(new_n16301_), .B(new_n16295_), .ZN(new_n16302_));
  OAI21_X1   g16110(.A1(new_n16302_), .A2(\asqrt[10] ), .B(new_n16255_), .ZN(new_n16303_));
  NAND2_X1   g16111(.A1(new_n16302_), .A2(\asqrt[10] ), .ZN(new_n16304_));
  AOI21_X1   g16112(.A1(new_n16303_), .A2(new_n16304_), .B(new_n14207_), .ZN(new_n16305_));
  NOR3_X1    g16113(.A1(new_n16299_), .A2(\asqrt[12] ), .A3(new_n16305_), .ZN(new_n16306_));
  OAI21_X1   g16114(.A1(new_n16299_), .A2(new_n16305_), .B(\asqrt[12] ), .ZN(new_n16307_));
  OAI21_X1   g16115(.A1(new_n16246_), .A2(new_n16306_), .B(new_n16307_), .ZN(new_n16308_));
  OAI21_X1   g16116(.A1(new_n16308_), .A2(\asqrt[13] ), .B(new_n16242_), .ZN(new_n16309_));
  NAND3_X1   g16117(.A1(new_n16303_), .A2(new_n16304_), .A3(new_n14207_), .ZN(new_n16310_));
  AOI21_X1   g16118(.A1(new_n16248_), .A2(new_n16310_), .B(new_n16305_), .ZN(new_n16311_));
  AOI21_X1   g16119(.A1(new_n16311_), .A2(new_n13690_), .B(new_n16246_), .ZN(new_n16312_));
  NAND2_X1   g16120(.A1(new_n16310_), .A2(new_n16248_), .ZN(new_n16313_));
  INV_X1     g16121(.I(new_n16305_), .ZN(new_n16314_));
  AOI21_X1   g16122(.A1(new_n16313_), .A2(new_n16314_), .B(new_n13690_), .ZN(new_n16315_));
  OAI21_X1   g16123(.A1(new_n16312_), .A2(new_n16315_), .B(\asqrt[13] ), .ZN(new_n16316_));
  NAND3_X1   g16124(.A1(new_n16309_), .A2(new_n12733_), .A3(new_n16316_), .ZN(new_n16317_));
  AOI21_X1   g16125(.A1(new_n16309_), .A2(new_n16316_), .B(new_n12733_), .ZN(new_n16318_));
  AOI21_X1   g16126(.A1(new_n16240_), .A2(new_n16317_), .B(new_n16318_), .ZN(new_n16319_));
  AOI21_X1   g16127(.A1(new_n16319_), .A2(new_n12283_), .B(new_n16237_), .ZN(new_n16320_));
  INV_X1     g16128(.I(new_n16242_), .ZN(new_n16321_));
  NOR3_X1    g16129(.A1(new_n16312_), .A2(\asqrt[13] ), .A3(new_n16315_), .ZN(new_n16322_));
  OAI21_X1   g16130(.A1(new_n16321_), .A2(new_n16322_), .B(new_n16316_), .ZN(new_n16323_));
  OAI21_X1   g16131(.A1(new_n16323_), .A2(\asqrt[14] ), .B(new_n16240_), .ZN(new_n16324_));
  NAND2_X1   g16132(.A1(new_n16323_), .A2(\asqrt[14] ), .ZN(new_n16325_));
  AOI21_X1   g16133(.A1(new_n16324_), .A2(new_n16325_), .B(new_n12283_), .ZN(new_n16326_));
  NOR3_X1    g16134(.A1(new_n16320_), .A2(\asqrt[16] ), .A3(new_n16326_), .ZN(new_n16327_));
  OAI21_X1   g16135(.A1(new_n16320_), .A2(new_n16326_), .B(\asqrt[16] ), .ZN(new_n16328_));
  OAI21_X1   g16136(.A1(new_n16234_), .A2(new_n16327_), .B(new_n16328_), .ZN(new_n16329_));
  OAI21_X1   g16137(.A1(new_n16329_), .A2(\asqrt[17] ), .B(new_n16230_), .ZN(new_n16330_));
  NAND3_X1   g16138(.A1(new_n16324_), .A2(new_n16325_), .A3(new_n12283_), .ZN(new_n16331_));
  AOI21_X1   g16139(.A1(new_n16236_), .A2(new_n16331_), .B(new_n16326_), .ZN(new_n16332_));
  AOI21_X1   g16140(.A1(new_n16332_), .A2(new_n11802_), .B(new_n16234_), .ZN(new_n16333_));
  NAND2_X1   g16141(.A1(new_n16331_), .A2(new_n16236_), .ZN(new_n16334_));
  INV_X1     g16142(.I(new_n16326_), .ZN(new_n16335_));
  AOI21_X1   g16143(.A1(new_n16334_), .A2(new_n16335_), .B(new_n11802_), .ZN(new_n16336_));
  OAI21_X1   g16144(.A1(new_n16333_), .A2(new_n16336_), .B(\asqrt[17] ), .ZN(new_n16337_));
  NAND3_X1   g16145(.A1(new_n16330_), .A2(new_n10914_), .A3(new_n16337_), .ZN(new_n16338_));
  AOI21_X1   g16146(.A1(new_n16330_), .A2(new_n16337_), .B(new_n10914_), .ZN(new_n16339_));
  AOI21_X1   g16147(.A1(new_n16228_), .A2(new_n16338_), .B(new_n16339_), .ZN(new_n16340_));
  AOI21_X1   g16148(.A1(new_n16340_), .A2(new_n10497_), .B(new_n16225_), .ZN(new_n16341_));
  INV_X1     g16149(.I(new_n16230_), .ZN(new_n16342_));
  NOR3_X1    g16150(.A1(new_n16333_), .A2(\asqrt[17] ), .A3(new_n16336_), .ZN(new_n16343_));
  OAI21_X1   g16151(.A1(new_n16342_), .A2(new_n16343_), .B(new_n16337_), .ZN(new_n16344_));
  OAI21_X1   g16152(.A1(new_n16344_), .A2(\asqrt[18] ), .B(new_n16228_), .ZN(new_n16345_));
  NAND2_X1   g16153(.A1(new_n16344_), .A2(\asqrt[18] ), .ZN(new_n16346_));
  AOI21_X1   g16154(.A1(new_n16345_), .A2(new_n16346_), .B(new_n10497_), .ZN(new_n16347_));
  NOR3_X1    g16155(.A1(new_n16341_), .A2(\asqrt[20] ), .A3(new_n16347_), .ZN(new_n16348_));
  OAI21_X1   g16156(.A1(new_n16341_), .A2(new_n16347_), .B(\asqrt[20] ), .ZN(new_n16349_));
  OAI21_X1   g16157(.A1(new_n16222_), .A2(new_n16348_), .B(new_n16349_), .ZN(new_n16350_));
  OAI21_X1   g16158(.A1(new_n16350_), .A2(\asqrt[21] ), .B(new_n16218_), .ZN(new_n16351_));
  NAND3_X1   g16159(.A1(new_n16345_), .A2(new_n16346_), .A3(new_n10497_), .ZN(new_n16352_));
  AOI21_X1   g16160(.A1(new_n16224_), .A2(new_n16352_), .B(new_n16347_), .ZN(new_n16353_));
  AOI21_X1   g16161(.A1(new_n16353_), .A2(new_n10052_), .B(new_n16222_), .ZN(new_n16354_));
  NAND2_X1   g16162(.A1(new_n16352_), .A2(new_n16224_), .ZN(new_n16355_));
  INV_X1     g16163(.I(new_n16347_), .ZN(new_n16356_));
  AOI21_X1   g16164(.A1(new_n16355_), .A2(new_n16356_), .B(new_n10052_), .ZN(new_n16357_));
  OAI21_X1   g16165(.A1(new_n16354_), .A2(new_n16357_), .B(\asqrt[21] ), .ZN(new_n16358_));
  NAND3_X1   g16166(.A1(new_n16351_), .A2(new_n9233_), .A3(new_n16358_), .ZN(new_n16359_));
  AOI21_X1   g16167(.A1(new_n16351_), .A2(new_n16358_), .B(new_n9233_), .ZN(new_n16360_));
  AOI21_X1   g16168(.A1(new_n16216_), .A2(new_n16359_), .B(new_n16360_), .ZN(new_n16361_));
  AOI21_X1   g16169(.A1(new_n16361_), .A2(new_n8849_), .B(new_n16213_), .ZN(new_n16362_));
  INV_X1     g16170(.I(new_n16218_), .ZN(new_n16363_));
  NOR3_X1    g16171(.A1(new_n16354_), .A2(\asqrt[21] ), .A3(new_n16357_), .ZN(new_n16364_));
  OAI21_X1   g16172(.A1(new_n16363_), .A2(new_n16364_), .B(new_n16358_), .ZN(new_n16365_));
  OAI21_X1   g16173(.A1(new_n16365_), .A2(\asqrt[22] ), .B(new_n16216_), .ZN(new_n16366_));
  NAND2_X1   g16174(.A1(new_n16365_), .A2(\asqrt[22] ), .ZN(new_n16367_));
  AOI21_X1   g16175(.A1(new_n16366_), .A2(new_n16367_), .B(new_n8849_), .ZN(new_n16368_));
  NOR3_X1    g16176(.A1(new_n16362_), .A2(\asqrt[24] ), .A3(new_n16368_), .ZN(new_n16369_));
  OAI21_X1   g16177(.A1(new_n16362_), .A2(new_n16368_), .B(\asqrt[24] ), .ZN(new_n16370_));
  OAI21_X1   g16178(.A1(new_n16210_), .A2(new_n16369_), .B(new_n16370_), .ZN(new_n16371_));
  OAI21_X1   g16179(.A1(new_n16371_), .A2(\asqrt[25] ), .B(new_n16206_), .ZN(new_n16372_));
  NAND3_X1   g16180(.A1(new_n16366_), .A2(new_n16367_), .A3(new_n8849_), .ZN(new_n16373_));
  AOI21_X1   g16181(.A1(new_n16212_), .A2(new_n16373_), .B(new_n16368_), .ZN(new_n16374_));
  AOI21_X1   g16182(.A1(new_n16374_), .A2(new_n8440_), .B(new_n16210_), .ZN(new_n16375_));
  NAND2_X1   g16183(.A1(new_n16373_), .A2(new_n16212_), .ZN(new_n16376_));
  INV_X1     g16184(.I(new_n16368_), .ZN(new_n16377_));
  AOI21_X1   g16185(.A1(new_n16376_), .A2(new_n16377_), .B(new_n8440_), .ZN(new_n16378_));
  OAI21_X1   g16186(.A1(new_n16375_), .A2(new_n16378_), .B(\asqrt[25] ), .ZN(new_n16379_));
  NAND3_X1   g16187(.A1(new_n16372_), .A2(new_n7690_), .A3(new_n16379_), .ZN(new_n16380_));
  AOI21_X1   g16188(.A1(new_n16372_), .A2(new_n16379_), .B(new_n7690_), .ZN(new_n16381_));
  AOI21_X1   g16189(.A1(new_n16204_), .A2(new_n16380_), .B(new_n16381_), .ZN(new_n16382_));
  AOI21_X1   g16190(.A1(new_n16382_), .A2(new_n7331_), .B(new_n16201_), .ZN(new_n16383_));
  INV_X1     g16191(.I(new_n16206_), .ZN(new_n16384_));
  NOR3_X1    g16192(.A1(new_n16375_), .A2(\asqrt[25] ), .A3(new_n16378_), .ZN(new_n16385_));
  OAI21_X1   g16193(.A1(new_n16384_), .A2(new_n16385_), .B(new_n16379_), .ZN(new_n16386_));
  OAI21_X1   g16194(.A1(new_n16386_), .A2(\asqrt[26] ), .B(new_n16204_), .ZN(new_n16387_));
  NAND2_X1   g16195(.A1(new_n16386_), .A2(\asqrt[26] ), .ZN(new_n16388_));
  AOI21_X1   g16196(.A1(new_n16387_), .A2(new_n16388_), .B(new_n7331_), .ZN(new_n16389_));
  NOR3_X1    g16197(.A1(new_n16383_), .A2(\asqrt[28] ), .A3(new_n16389_), .ZN(new_n16390_));
  OAI21_X1   g16198(.A1(new_n16383_), .A2(new_n16389_), .B(\asqrt[28] ), .ZN(new_n16391_));
  OAI21_X1   g16199(.A1(new_n16198_), .A2(new_n16390_), .B(new_n16391_), .ZN(new_n16392_));
  OAI21_X1   g16200(.A1(new_n16392_), .A2(\asqrt[29] ), .B(new_n16194_), .ZN(new_n16393_));
  NAND3_X1   g16201(.A1(new_n16387_), .A2(new_n16388_), .A3(new_n7331_), .ZN(new_n16394_));
  AOI21_X1   g16202(.A1(new_n16200_), .A2(new_n16394_), .B(new_n16389_), .ZN(new_n16395_));
  AOI21_X1   g16203(.A1(new_n16395_), .A2(new_n6966_), .B(new_n16198_), .ZN(new_n16396_));
  NAND2_X1   g16204(.A1(new_n16394_), .A2(new_n16200_), .ZN(new_n16397_));
  INV_X1     g16205(.I(new_n16389_), .ZN(new_n16398_));
  AOI21_X1   g16206(.A1(new_n16397_), .A2(new_n16398_), .B(new_n6966_), .ZN(new_n16399_));
  OAI21_X1   g16207(.A1(new_n16396_), .A2(new_n16399_), .B(\asqrt[29] ), .ZN(new_n16400_));
  NAND3_X1   g16208(.A1(new_n16393_), .A2(new_n6275_), .A3(new_n16400_), .ZN(new_n16401_));
  AOI21_X1   g16209(.A1(new_n16393_), .A2(new_n16400_), .B(new_n6275_), .ZN(new_n16402_));
  AOI21_X1   g16210(.A1(new_n16192_), .A2(new_n16401_), .B(new_n16402_), .ZN(new_n16403_));
  AOI21_X1   g16211(.A1(new_n16403_), .A2(new_n5947_), .B(new_n16189_), .ZN(new_n16404_));
  INV_X1     g16212(.I(new_n16194_), .ZN(new_n16405_));
  NOR3_X1    g16213(.A1(new_n16396_), .A2(\asqrt[29] ), .A3(new_n16399_), .ZN(new_n16406_));
  OAI21_X1   g16214(.A1(new_n16405_), .A2(new_n16406_), .B(new_n16400_), .ZN(new_n16407_));
  OAI21_X1   g16215(.A1(new_n16407_), .A2(\asqrt[30] ), .B(new_n16192_), .ZN(new_n16408_));
  NAND2_X1   g16216(.A1(new_n16407_), .A2(\asqrt[30] ), .ZN(new_n16409_));
  AOI21_X1   g16217(.A1(new_n16408_), .A2(new_n16409_), .B(new_n5947_), .ZN(new_n16410_));
  NOR3_X1    g16218(.A1(new_n16404_), .A2(\asqrt[32] ), .A3(new_n16410_), .ZN(new_n16411_));
  OAI21_X1   g16219(.A1(new_n16404_), .A2(new_n16410_), .B(\asqrt[32] ), .ZN(new_n16412_));
  OAI21_X1   g16220(.A1(new_n16186_), .A2(new_n16411_), .B(new_n16412_), .ZN(new_n16413_));
  OAI21_X1   g16221(.A1(new_n16413_), .A2(\asqrt[33] ), .B(new_n16182_), .ZN(new_n16414_));
  NAND3_X1   g16222(.A1(new_n16408_), .A2(new_n16409_), .A3(new_n5947_), .ZN(new_n16415_));
  AOI21_X1   g16223(.A1(new_n16188_), .A2(new_n16415_), .B(new_n16410_), .ZN(new_n16416_));
  AOI21_X1   g16224(.A1(new_n16416_), .A2(new_n5643_), .B(new_n16186_), .ZN(new_n16417_));
  NAND2_X1   g16225(.A1(new_n16415_), .A2(new_n16188_), .ZN(new_n16418_));
  INV_X1     g16226(.I(new_n16410_), .ZN(new_n16419_));
  AOI21_X1   g16227(.A1(new_n16418_), .A2(new_n16419_), .B(new_n5643_), .ZN(new_n16420_));
  OAI21_X1   g16228(.A1(new_n16417_), .A2(new_n16420_), .B(\asqrt[33] ), .ZN(new_n16421_));
  NAND3_X1   g16229(.A1(new_n16414_), .A2(new_n5029_), .A3(new_n16421_), .ZN(new_n16422_));
  AOI21_X1   g16230(.A1(new_n16414_), .A2(new_n16421_), .B(new_n5029_), .ZN(new_n16423_));
  AOI21_X1   g16231(.A1(new_n16180_), .A2(new_n16422_), .B(new_n16423_), .ZN(new_n16424_));
  AOI21_X1   g16232(.A1(new_n16424_), .A2(new_n4751_), .B(new_n16177_), .ZN(new_n16425_));
  INV_X1     g16233(.I(new_n16182_), .ZN(new_n16426_));
  NOR3_X1    g16234(.A1(new_n16417_), .A2(\asqrt[33] ), .A3(new_n16420_), .ZN(new_n16427_));
  OAI21_X1   g16235(.A1(new_n16426_), .A2(new_n16427_), .B(new_n16421_), .ZN(new_n16428_));
  OAI21_X1   g16236(.A1(new_n16428_), .A2(\asqrt[34] ), .B(new_n16180_), .ZN(new_n16429_));
  NAND2_X1   g16237(.A1(new_n16428_), .A2(\asqrt[34] ), .ZN(new_n16430_));
  AOI21_X1   g16238(.A1(new_n16429_), .A2(new_n16430_), .B(new_n4751_), .ZN(new_n16431_));
  NOR3_X1    g16239(.A1(new_n16425_), .A2(\asqrt[36] ), .A3(new_n16431_), .ZN(new_n16432_));
  OAI21_X1   g16240(.A1(new_n16425_), .A2(new_n16431_), .B(\asqrt[36] ), .ZN(new_n16433_));
  OAI21_X1   g16241(.A1(new_n16174_), .A2(new_n16432_), .B(new_n16433_), .ZN(new_n16434_));
  OAI21_X1   g16242(.A1(new_n16434_), .A2(\asqrt[37] ), .B(new_n16170_), .ZN(new_n16435_));
  NAND3_X1   g16243(.A1(new_n16429_), .A2(new_n16430_), .A3(new_n4751_), .ZN(new_n16436_));
  AOI21_X1   g16244(.A1(new_n16176_), .A2(new_n16436_), .B(new_n16431_), .ZN(new_n16437_));
  AOI21_X1   g16245(.A1(new_n16437_), .A2(new_n4461_), .B(new_n16174_), .ZN(new_n16438_));
  NAND2_X1   g16246(.A1(new_n16436_), .A2(new_n16176_), .ZN(new_n16439_));
  INV_X1     g16247(.I(new_n16431_), .ZN(new_n16440_));
  AOI21_X1   g16248(.A1(new_n16439_), .A2(new_n16440_), .B(new_n4461_), .ZN(new_n16441_));
  OAI21_X1   g16249(.A1(new_n16438_), .A2(new_n16441_), .B(\asqrt[37] ), .ZN(new_n16442_));
  NAND3_X1   g16250(.A1(new_n16435_), .A2(new_n3925_), .A3(new_n16442_), .ZN(new_n16443_));
  AOI21_X1   g16251(.A1(new_n16435_), .A2(new_n16442_), .B(new_n3925_), .ZN(new_n16444_));
  AOI21_X1   g16252(.A1(new_n16168_), .A2(new_n16443_), .B(new_n16444_), .ZN(new_n16445_));
  AOI21_X1   g16253(.A1(new_n16445_), .A2(new_n3681_), .B(new_n16165_), .ZN(new_n16446_));
  INV_X1     g16254(.I(new_n16170_), .ZN(new_n16447_));
  NOR3_X1    g16255(.A1(new_n16438_), .A2(\asqrt[37] ), .A3(new_n16441_), .ZN(new_n16448_));
  OAI21_X1   g16256(.A1(new_n16447_), .A2(new_n16448_), .B(new_n16442_), .ZN(new_n16449_));
  OAI21_X1   g16257(.A1(new_n16449_), .A2(\asqrt[38] ), .B(new_n16168_), .ZN(new_n16450_));
  NAND2_X1   g16258(.A1(new_n16449_), .A2(\asqrt[38] ), .ZN(new_n16451_));
  AOI21_X1   g16259(.A1(new_n16450_), .A2(new_n16451_), .B(new_n3681_), .ZN(new_n16452_));
  NOR3_X1    g16260(.A1(new_n16446_), .A2(\asqrt[40] ), .A3(new_n16452_), .ZN(new_n16453_));
  OAI21_X1   g16261(.A1(new_n16446_), .A2(new_n16452_), .B(\asqrt[40] ), .ZN(new_n16454_));
  OAI21_X1   g16262(.A1(new_n16162_), .A2(new_n16453_), .B(new_n16454_), .ZN(new_n16455_));
  OAI21_X1   g16263(.A1(new_n16455_), .A2(\asqrt[41] ), .B(new_n16158_), .ZN(new_n16456_));
  NAND3_X1   g16264(.A1(new_n16450_), .A2(new_n16451_), .A3(new_n3681_), .ZN(new_n16457_));
  AOI21_X1   g16265(.A1(new_n16164_), .A2(new_n16457_), .B(new_n16452_), .ZN(new_n16458_));
  AOI21_X1   g16266(.A1(new_n16458_), .A2(new_n3427_), .B(new_n16162_), .ZN(new_n16459_));
  NAND2_X1   g16267(.A1(new_n16457_), .A2(new_n16164_), .ZN(new_n16460_));
  INV_X1     g16268(.I(new_n16452_), .ZN(new_n16461_));
  AOI21_X1   g16269(.A1(new_n16460_), .A2(new_n16461_), .B(new_n3427_), .ZN(new_n16462_));
  OAI21_X1   g16270(.A1(new_n16459_), .A2(new_n16462_), .B(\asqrt[41] ), .ZN(new_n16463_));
  NAND3_X1   g16271(.A1(new_n16456_), .A2(new_n2960_), .A3(new_n16463_), .ZN(new_n16464_));
  AOI21_X1   g16272(.A1(new_n16456_), .A2(new_n16463_), .B(new_n2960_), .ZN(new_n16465_));
  AOI21_X1   g16273(.A1(new_n16156_), .A2(new_n16464_), .B(new_n16465_), .ZN(new_n16466_));
  AOI21_X1   g16274(.A1(new_n16466_), .A2(new_n2749_), .B(new_n16153_), .ZN(new_n16467_));
  INV_X1     g16275(.I(new_n16158_), .ZN(new_n16468_));
  NOR3_X1    g16276(.A1(new_n16459_), .A2(\asqrt[41] ), .A3(new_n16462_), .ZN(new_n16469_));
  OAI21_X1   g16277(.A1(new_n16468_), .A2(new_n16469_), .B(new_n16463_), .ZN(new_n16470_));
  OAI21_X1   g16278(.A1(new_n16470_), .A2(\asqrt[42] ), .B(new_n16156_), .ZN(new_n16471_));
  NAND2_X1   g16279(.A1(new_n16470_), .A2(\asqrt[42] ), .ZN(new_n16472_));
  AOI21_X1   g16280(.A1(new_n16471_), .A2(new_n16472_), .B(new_n2749_), .ZN(new_n16473_));
  NOR3_X1    g16281(.A1(new_n16467_), .A2(\asqrt[44] ), .A3(new_n16473_), .ZN(new_n16474_));
  OAI21_X1   g16282(.A1(new_n16467_), .A2(new_n16473_), .B(\asqrt[44] ), .ZN(new_n16475_));
  OAI21_X1   g16283(.A1(new_n16150_), .A2(new_n16474_), .B(new_n16475_), .ZN(new_n16476_));
  OAI21_X1   g16284(.A1(new_n16476_), .A2(\asqrt[45] ), .B(new_n16146_), .ZN(new_n16477_));
  NAND3_X1   g16285(.A1(new_n16471_), .A2(new_n16472_), .A3(new_n2749_), .ZN(new_n16478_));
  AOI21_X1   g16286(.A1(new_n16152_), .A2(new_n16478_), .B(new_n16473_), .ZN(new_n16479_));
  AOI21_X1   g16287(.A1(new_n16479_), .A2(new_n2531_), .B(new_n16150_), .ZN(new_n16480_));
  NAND2_X1   g16288(.A1(new_n16478_), .A2(new_n16152_), .ZN(new_n16481_));
  INV_X1     g16289(.I(new_n16473_), .ZN(new_n16482_));
  AOI21_X1   g16290(.A1(new_n16481_), .A2(new_n16482_), .B(new_n2531_), .ZN(new_n16483_));
  OAI21_X1   g16291(.A1(new_n16480_), .A2(new_n16483_), .B(\asqrt[45] ), .ZN(new_n16484_));
  NAND3_X1   g16292(.A1(new_n16477_), .A2(new_n2134_), .A3(new_n16484_), .ZN(new_n16485_));
  AOI21_X1   g16293(.A1(new_n16477_), .A2(new_n16484_), .B(new_n2134_), .ZN(new_n16486_));
  AOI21_X1   g16294(.A1(new_n16144_), .A2(new_n16485_), .B(new_n16486_), .ZN(new_n16487_));
  AOI21_X1   g16295(.A1(new_n16487_), .A2(new_n1953_), .B(new_n16141_), .ZN(new_n16488_));
  INV_X1     g16296(.I(new_n16146_), .ZN(new_n16489_));
  NOR3_X1    g16297(.A1(new_n16480_), .A2(\asqrt[45] ), .A3(new_n16483_), .ZN(new_n16490_));
  OAI21_X1   g16298(.A1(new_n16489_), .A2(new_n16490_), .B(new_n16484_), .ZN(new_n16491_));
  OAI21_X1   g16299(.A1(new_n16491_), .A2(\asqrt[46] ), .B(new_n16144_), .ZN(new_n16492_));
  NAND2_X1   g16300(.A1(new_n16491_), .A2(\asqrt[46] ), .ZN(new_n16493_));
  AOI21_X1   g16301(.A1(new_n16492_), .A2(new_n16493_), .B(new_n1953_), .ZN(new_n16494_));
  NOR3_X1    g16302(.A1(new_n16488_), .A2(\asqrt[48] ), .A3(new_n16494_), .ZN(new_n16495_));
  OAI21_X1   g16303(.A1(new_n16488_), .A2(new_n16494_), .B(\asqrt[48] ), .ZN(new_n16496_));
  OAI21_X1   g16304(.A1(new_n16138_), .A2(new_n16495_), .B(new_n16496_), .ZN(new_n16497_));
  OAI21_X1   g16305(.A1(new_n16497_), .A2(\asqrt[49] ), .B(new_n16134_), .ZN(new_n16498_));
  NAND3_X1   g16306(.A1(new_n16492_), .A2(new_n16493_), .A3(new_n1953_), .ZN(new_n16499_));
  AOI21_X1   g16307(.A1(new_n16140_), .A2(new_n16499_), .B(new_n16494_), .ZN(new_n16500_));
  AOI21_X1   g16308(.A1(new_n16500_), .A2(new_n1778_), .B(new_n16138_), .ZN(new_n16501_));
  NAND2_X1   g16309(.A1(new_n16499_), .A2(new_n16140_), .ZN(new_n16502_));
  INV_X1     g16310(.I(new_n16494_), .ZN(new_n16503_));
  AOI21_X1   g16311(.A1(new_n16502_), .A2(new_n16503_), .B(new_n1778_), .ZN(new_n16504_));
  OAI21_X1   g16312(.A1(new_n16501_), .A2(new_n16504_), .B(\asqrt[49] ), .ZN(new_n16505_));
  NAND3_X1   g16313(.A1(new_n16498_), .A2(new_n1463_), .A3(new_n16505_), .ZN(new_n16506_));
  AOI21_X1   g16314(.A1(new_n16498_), .A2(new_n16505_), .B(new_n1463_), .ZN(new_n16507_));
  AOI21_X1   g16315(.A1(new_n16132_), .A2(new_n16506_), .B(new_n16507_), .ZN(new_n16508_));
  AOI21_X1   g16316(.A1(new_n16508_), .A2(new_n1305_), .B(new_n16129_), .ZN(new_n16509_));
  INV_X1     g16317(.I(new_n16134_), .ZN(new_n16510_));
  NOR3_X1    g16318(.A1(new_n16501_), .A2(\asqrt[49] ), .A3(new_n16504_), .ZN(new_n16511_));
  OAI21_X1   g16319(.A1(new_n16510_), .A2(new_n16511_), .B(new_n16505_), .ZN(new_n16512_));
  OAI21_X1   g16320(.A1(new_n16512_), .A2(\asqrt[50] ), .B(new_n16132_), .ZN(new_n16513_));
  NAND2_X1   g16321(.A1(new_n16512_), .A2(\asqrt[50] ), .ZN(new_n16514_));
  AOI21_X1   g16322(.A1(new_n16513_), .A2(new_n16514_), .B(new_n1305_), .ZN(new_n16515_));
  NOR3_X1    g16323(.A1(new_n16509_), .A2(\asqrt[52] ), .A3(new_n16515_), .ZN(new_n16516_));
  OAI21_X1   g16324(.A1(new_n16509_), .A2(new_n16515_), .B(\asqrt[52] ), .ZN(new_n16517_));
  OAI21_X1   g16325(.A1(new_n16126_), .A2(new_n16516_), .B(new_n16517_), .ZN(new_n16518_));
  OAI21_X1   g16326(.A1(new_n16518_), .A2(\asqrt[53] ), .B(new_n16122_), .ZN(new_n16519_));
  NAND3_X1   g16327(.A1(new_n16513_), .A2(new_n16514_), .A3(new_n1305_), .ZN(new_n16520_));
  AOI21_X1   g16328(.A1(new_n16128_), .A2(new_n16520_), .B(new_n16515_), .ZN(new_n16521_));
  AOI21_X1   g16329(.A1(new_n16521_), .A2(new_n1150_), .B(new_n16126_), .ZN(new_n16522_));
  NAND2_X1   g16330(.A1(new_n16520_), .A2(new_n16128_), .ZN(new_n16523_));
  INV_X1     g16331(.I(new_n16515_), .ZN(new_n16524_));
  AOI21_X1   g16332(.A1(new_n16523_), .A2(new_n16524_), .B(new_n1150_), .ZN(new_n16525_));
  OAI21_X1   g16333(.A1(new_n16522_), .A2(new_n16525_), .B(\asqrt[53] ), .ZN(new_n16526_));
  NAND3_X1   g16334(.A1(new_n16519_), .A2(new_n860_), .A3(new_n16526_), .ZN(new_n16527_));
  AOI21_X1   g16335(.A1(new_n16519_), .A2(new_n16526_), .B(new_n860_), .ZN(new_n16528_));
  AOI21_X1   g16336(.A1(new_n16120_), .A2(new_n16527_), .B(new_n16528_), .ZN(new_n16529_));
  AOI21_X1   g16337(.A1(new_n16529_), .A2(new_n744_), .B(new_n16117_), .ZN(new_n16530_));
  INV_X1     g16338(.I(new_n16122_), .ZN(new_n16531_));
  NOR3_X1    g16339(.A1(new_n16522_), .A2(\asqrt[53] ), .A3(new_n16525_), .ZN(new_n16532_));
  OAI21_X1   g16340(.A1(new_n16531_), .A2(new_n16532_), .B(new_n16526_), .ZN(new_n16533_));
  OAI21_X1   g16341(.A1(new_n16533_), .A2(\asqrt[54] ), .B(new_n16120_), .ZN(new_n16534_));
  NAND2_X1   g16342(.A1(new_n16533_), .A2(\asqrt[54] ), .ZN(new_n16535_));
  AOI21_X1   g16343(.A1(new_n16534_), .A2(new_n16535_), .B(new_n744_), .ZN(new_n16536_));
  NOR3_X1    g16344(.A1(new_n16530_), .A2(\asqrt[56] ), .A3(new_n16536_), .ZN(new_n16537_));
  OAI21_X1   g16345(.A1(new_n16530_), .A2(new_n16536_), .B(\asqrt[56] ), .ZN(new_n16538_));
  OAI21_X1   g16346(.A1(new_n16114_), .A2(new_n16537_), .B(new_n16538_), .ZN(new_n16539_));
  OAI21_X1   g16347(.A1(new_n16539_), .A2(\asqrt[57] ), .B(new_n16110_), .ZN(new_n16540_));
  NAND3_X1   g16348(.A1(new_n16534_), .A2(new_n16535_), .A3(new_n744_), .ZN(new_n16541_));
  AOI21_X1   g16349(.A1(new_n16116_), .A2(new_n16541_), .B(new_n16536_), .ZN(new_n16542_));
  AOI21_X1   g16350(.A1(new_n16542_), .A2(new_n634_), .B(new_n16114_), .ZN(new_n16543_));
  NAND2_X1   g16351(.A1(new_n16541_), .A2(new_n16116_), .ZN(new_n16544_));
  INV_X1     g16352(.I(new_n16536_), .ZN(new_n16545_));
  AOI21_X1   g16353(.A1(new_n16544_), .A2(new_n16545_), .B(new_n634_), .ZN(new_n16546_));
  OAI21_X1   g16354(.A1(new_n16543_), .A2(new_n16546_), .B(\asqrt[57] ), .ZN(new_n16547_));
  NAND3_X1   g16355(.A1(new_n16540_), .A2(new_n423_), .A3(new_n16547_), .ZN(new_n16548_));
  INV_X1     g16356(.I(new_n16110_), .ZN(new_n16549_));
  NOR3_X1    g16357(.A1(new_n16543_), .A2(\asqrt[57] ), .A3(new_n16546_), .ZN(new_n16550_));
  NOR2_X1    g16358(.A1(new_n16550_), .A2(new_n16549_), .ZN(new_n16551_));
  INV_X1     g16359(.I(new_n16547_), .ZN(new_n16552_));
  OAI21_X1   g16360(.A1(new_n16551_), .A2(new_n16552_), .B(\asqrt[58] ), .ZN(new_n16553_));
  NAND2_X1   g16361(.A1(new_n16256_), .A2(new_n201_), .ZN(new_n16554_));
  AOI21_X1   g16362(.A1(new_n16554_), .A2(new_n16097_), .B(\asqrt[7] ), .ZN(new_n16555_));
  XOR2_X1    g16363(.A1(new_n16555_), .A2(new_n16089_), .Z(new_n16556_));
  INV_X1     g16364(.I(new_n16556_), .ZN(new_n16557_));
  AOI21_X1   g16365(.A1(new_n16057_), .A2(new_n16065_), .B(\asqrt[7] ), .ZN(new_n16558_));
  XOR2_X1    g16366(.A1(new_n16558_), .A2(new_n16044_), .Z(new_n16559_));
  INV_X1     g16367(.I(new_n16559_), .ZN(new_n16560_));
  AOI21_X1   g16368(.A1(new_n16050_), .A2(new_n16056_), .B(\asqrt[7] ), .ZN(new_n16561_));
  XOR2_X1    g16369(.A1(new_n16561_), .A2(new_n16046_), .Z(new_n16562_));
  INV_X1     g16370(.I(new_n16562_), .ZN(new_n16563_));
  AOI21_X1   g16371(.A1(new_n16540_), .A2(new_n16547_), .B(new_n423_), .ZN(new_n16564_));
  AOI21_X1   g16372(.A1(new_n16108_), .A2(new_n16548_), .B(new_n16564_), .ZN(new_n16565_));
  AOI21_X1   g16373(.A1(new_n16565_), .A2(new_n337_), .B(new_n16563_), .ZN(new_n16566_));
  NOR2_X1    g16374(.A1(new_n16565_), .A2(new_n337_), .ZN(new_n16567_));
  NOR3_X1    g16375(.A1(new_n16566_), .A2(new_n16567_), .A3(\asqrt[60] ), .ZN(new_n16568_));
  OAI21_X1   g16376(.A1(new_n16566_), .A2(new_n16567_), .B(\asqrt[60] ), .ZN(new_n16569_));
  OAI21_X1   g16377(.A1(new_n16560_), .A2(new_n16568_), .B(new_n16569_), .ZN(new_n16570_));
  NAND2_X1   g16378(.A1(new_n16570_), .A2(\asqrt[61] ), .ZN(new_n16571_));
  AOI21_X1   g16379(.A1(new_n16073_), .A2(new_n16079_), .B(\asqrt[7] ), .ZN(new_n16572_));
  XOR2_X1    g16380(.A1(new_n16572_), .A2(new_n16040_), .Z(new_n16573_));
  OAI21_X1   g16381(.A1(new_n16570_), .A2(\asqrt[61] ), .B(new_n16573_), .ZN(new_n16574_));
  NAND2_X1   g16382(.A1(new_n16574_), .A2(new_n16571_), .ZN(new_n16575_));
  OAI21_X1   g16383(.A1(new_n16549_), .A2(new_n16550_), .B(new_n16547_), .ZN(new_n16576_));
  OAI21_X1   g16384(.A1(new_n16576_), .A2(\asqrt[58] ), .B(new_n16108_), .ZN(new_n16577_));
  NAND3_X1   g16385(.A1(new_n16577_), .A2(new_n337_), .A3(new_n16553_), .ZN(new_n16578_));
  NAND2_X1   g16386(.A1(new_n16578_), .A2(new_n16562_), .ZN(new_n16579_));
  INV_X1     g16387(.I(new_n16108_), .ZN(new_n16580_));
  NOR2_X1    g16388(.A1(new_n16551_), .A2(new_n16552_), .ZN(new_n16581_));
  AOI21_X1   g16389(.A1(new_n16581_), .A2(new_n423_), .B(new_n16580_), .ZN(new_n16582_));
  OAI21_X1   g16390(.A1(new_n16582_), .A2(new_n16564_), .B(\asqrt[59] ), .ZN(new_n16583_));
  NAND3_X1   g16391(.A1(new_n16579_), .A2(new_n266_), .A3(new_n16583_), .ZN(new_n16584_));
  NAND2_X1   g16392(.A1(new_n16584_), .A2(new_n16559_), .ZN(new_n16585_));
  AOI21_X1   g16393(.A1(new_n16585_), .A2(new_n16569_), .B(new_n239_), .ZN(new_n16586_));
  AOI21_X1   g16394(.A1(new_n16579_), .A2(new_n16583_), .B(new_n266_), .ZN(new_n16587_));
  AOI21_X1   g16395(.A1(new_n16559_), .A2(new_n16584_), .B(new_n16587_), .ZN(new_n16588_));
  INV_X1     g16396(.I(new_n16573_), .ZN(new_n16589_));
  AOI21_X1   g16397(.A1(new_n16588_), .A2(new_n239_), .B(new_n16589_), .ZN(new_n16590_));
  OAI21_X1   g16398(.A1(new_n16590_), .A2(new_n16586_), .B(new_n201_), .ZN(new_n16591_));
  NAND3_X1   g16399(.A1(new_n16574_), .A2(new_n16571_), .A3(\asqrt[62] ), .ZN(new_n16592_));
  NOR2_X1    g16400(.A1(new_n16071_), .A2(new_n16080_), .ZN(new_n16593_));
  NOR2_X1    g16401(.A1(\asqrt[7] ), .A2(new_n16593_), .ZN(new_n16594_));
  XOR2_X1    g16402(.A1(new_n16594_), .A2(new_n16069_), .Z(new_n16595_));
  INV_X1     g16403(.I(new_n16595_), .ZN(new_n16596_));
  AOI22_X1   g16404(.A1(new_n16592_), .A2(new_n16591_), .B1(new_n16575_), .B2(new_n16596_), .ZN(new_n16597_));
  NOR2_X1    g16405(.A1(new_n16091_), .A2(new_n16037_), .ZN(new_n16598_));
  OAI21_X1   g16406(.A1(\asqrt[7] ), .A2(new_n16598_), .B(new_n16098_), .ZN(new_n16599_));
  INV_X1     g16407(.I(new_n16599_), .ZN(new_n16600_));
  OAI21_X1   g16408(.A1(new_n16597_), .A2(new_n16557_), .B(new_n16600_), .ZN(new_n16601_));
  OAI21_X1   g16409(.A1(new_n16575_), .A2(\asqrt[62] ), .B(new_n16595_), .ZN(new_n16602_));
  NAND2_X1   g16410(.A1(new_n16575_), .A2(\asqrt[62] ), .ZN(new_n16603_));
  NAND3_X1   g16411(.A1(new_n16602_), .A2(new_n16603_), .A3(new_n16557_), .ZN(new_n16604_));
  XOR2_X1    g16412(.A1(new_n16259_), .A2(new_n16037_), .Z(new_n16605_));
  NOR2_X1    g16413(.A1(new_n16605_), .A2(new_n193_), .ZN(new_n16606_));
  OAI21_X1   g16414(.A1(new_n16037_), .A2(\asqrt[7] ), .B(new_n16606_), .ZN(new_n16607_));
  NOR2_X1    g16415(.A1(new_n16104_), .A2(new_n16036_), .ZN(new_n16608_));
  NAND4_X1   g16416(.A1(new_n16095_), .A2(new_n193_), .A3(new_n16098_), .A4(new_n16608_), .ZN(new_n16609_));
  NAND2_X1   g16417(.A1(new_n16607_), .A2(new_n16609_), .ZN(new_n16610_));
  INV_X1     g16418(.I(new_n16610_), .ZN(new_n16611_));
  NAND4_X1   g16419(.A1(new_n16601_), .A2(new_n193_), .A3(new_n16604_), .A4(new_n16611_), .ZN(\asqrt[6] ));
  AOI21_X1   g16420(.A1(new_n16548_), .A2(new_n16553_), .B(\asqrt[6] ), .ZN(new_n16613_));
  XOR2_X1    g16421(.A1(new_n16613_), .A2(new_n16108_), .Z(new_n16614_));
  NOR2_X1    g16422(.A1(new_n16552_), .A2(new_n16550_), .ZN(new_n16615_));
  NOR2_X1    g16423(.A1(\asqrt[6] ), .A2(new_n16615_), .ZN(new_n16616_));
  XOR2_X1    g16424(.A1(new_n16616_), .A2(new_n16110_), .Z(new_n16617_));
  NOR2_X1    g16425(.A1(new_n16537_), .A2(new_n16546_), .ZN(new_n16618_));
  NOR2_X1    g16426(.A1(\asqrt[6] ), .A2(new_n16618_), .ZN(new_n16619_));
  XOR2_X1    g16427(.A1(new_n16619_), .A2(new_n16113_), .Z(new_n16620_));
  AOI21_X1   g16428(.A1(new_n16541_), .A2(new_n16545_), .B(\asqrt[6] ), .ZN(new_n16621_));
  XOR2_X1    g16429(.A1(new_n16621_), .A2(new_n16116_), .Z(new_n16622_));
  INV_X1     g16430(.I(new_n16622_), .ZN(new_n16623_));
  AOI21_X1   g16431(.A1(new_n16527_), .A2(new_n16535_), .B(\asqrt[6] ), .ZN(new_n16624_));
  XOR2_X1    g16432(.A1(new_n16624_), .A2(new_n16120_), .Z(new_n16625_));
  INV_X1     g16433(.I(new_n16625_), .ZN(new_n16626_));
  XOR2_X1    g16434(.A1(new_n16518_), .A2(\asqrt[53] ), .Z(new_n16627_));
  NOR2_X1    g16435(.A1(\asqrt[6] ), .A2(new_n16627_), .ZN(new_n16628_));
  XOR2_X1    g16436(.A1(new_n16628_), .A2(new_n16122_), .Z(new_n16629_));
  NOR2_X1    g16437(.A1(new_n16516_), .A2(new_n16525_), .ZN(new_n16630_));
  NOR2_X1    g16438(.A1(\asqrt[6] ), .A2(new_n16630_), .ZN(new_n16631_));
  XOR2_X1    g16439(.A1(new_n16631_), .A2(new_n16125_), .Z(new_n16632_));
  AOI21_X1   g16440(.A1(new_n16520_), .A2(new_n16524_), .B(\asqrt[6] ), .ZN(new_n16633_));
  XOR2_X1    g16441(.A1(new_n16633_), .A2(new_n16128_), .Z(new_n16634_));
  INV_X1     g16442(.I(new_n16634_), .ZN(new_n16635_));
  AOI21_X1   g16443(.A1(new_n16506_), .A2(new_n16514_), .B(\asqrt[6] ), .ZN(new_n16636_));
  XOR2_X1    g16444(.A1(new_n16636_), .A2(new_n16132_), .Z(new_n16637_));
  INV_X1     g16445(.I(new_n16637_), .ZN(new_n16638_));
  XOR2_X1    g16446(.A1(new_n16497_), .A2(\asqrt[49] ), .Z(new_n16639_));
  NOR2_X1    g16447(.A1(\asqrt[6] ), .A2(new_n16639_), .ZN(new_n16640_));
  XOR2_X1    g16448(.A1(new_n16640_), .A2(new_n16134_), .Z(new_n16641_));
  NOR2_X1    g16449(.A1(new_n16495_), .A2(new_n16504_), .ZN(new_n16642_));
  NOR2_X1    g16450(.A1(\asqrt[6] ), .A2(new_n16642_), .ZN(new_n16643_));
  XOR2_X1    g16451(.A1(new_n16643_), .A2(new_n16137_), .Z(new_n16644_));
  AOI21_X1   g16452(.A1(new_n16499_), .A2(new_n16503_), .B(\asqrt[6] ), .ZN(new_n16645_));
  XOR2_X1    g16453(.A1(new_n16645_), .A2(new_n16140_), .Z(new_n16646_));
  INV_X1     g16454(.I(new_n16646_), .ZN(new_n16647_));
  AOI21_X1   g16455(.A1(new_n16485_), .A2(new_n16493_), .B(\asqrt[6] ), .ZN(new_n16648_));
  XOR2_X1    g16456(.A1(new_n16648_), .A2(new_n16144_), .Z(new_n16649_));
  INV_X1     g16457(.I(new_n16649_), .ZN(new_n16650_));
  XOR2_X1    g16458(.A1(new_n16476_), .A2(\asqrt[45] ), .Z(new_n16651_));
  NOR2_X1    g16459(.A1(\asqrt[6] ), .A2(new_n16651_), .ZN(new_n16652_));
  XOR2_X1    g16460(.A1(new_n16652_), .A2(new_n16146_), .Z(new_n16653_));
  NOR2_X1    g16461(.A1(new_n16474_), .A2(new_n16483_), .ZN(new_n16654_));
  NOR2_X1    g16462(.A1(\asqrt[6] ), .A2(new_n16654_), .ZN(new_n16655_));
  XOR2_X1    g16463(.A1(new_n16655_), .A2(new_n16149_), .Z(new_n16656_));
  AOI21_X1   g16464(.A1(new_n16478_), .A2(new_n16482_), .B(\asqrt[6] ), .ZN(new_n16657_));
  XOR2_X1    g16465(.A1(new_n16657_), .A2(new_n16152_), .Z(new_n16658_));
  INV_X1     g16466(.I(new_n16658_), .ZN(new_n16659_));
  AOI21_X1   g16467(.A1(new_n16464_), .A2(new_n16472_), .B(\asqrt[6] ), .ZN(new_n16660_));
  XOR2_X1    g16468(.A1(new_n16660_), .A2(new_n16156_), .Z(new_n16661_));
  INV_X1     g16469(.I(new_n16661_), .ZN(new_n16662_));
  XOR2_X1    g16470(.A1(new_n16455_), .A2(\asqrt[41] ), .Z(new_n16663_));
  NOR2_X1    g16471(.A1(\asqrt[6] ), .A2(new_n16663_), .ZN(new_n16664_));
  XOR2_X1    g16472(.A1(new_n16664_), .A2(new_n16158_), .Z(new_n16665_));
  NOR2_X1    g16473(.A1(new_n16453_), .A2(new_n16462_), .ZN(new_n16666_));
  NOR2_X1    g16474(.A1(\asqrt[6] ), .A2(new_n16666_), .ZN(new_n16667_));
  XOR2_X1    g16475(.A1(new_n16667_), .A2(new_n16161_), .Z(new_n16668_));
  AOI21_X1   g16476(.A1(new_n16457_), .A2(new_n16461_), .B(\asqrt[6] ), .ZN(new_n16669_));
  XOR2_X1    g16477(.A1(new_n16669_), .A2(new_n16164_), .Z(new_n16670_));
  INV_X1     g16478(.I(new_n16670_), .ZN(new_n16671_));
  AOI21_X1   g16479(.A1(new_n16443_), .A2(new_n16451_), .B(\asqrt[6] ), .ZN(new_n16672_));
  XOR2_X1    g16480(.A1(new_n16672_), .A2(new_n16168_), .Z(new_n16673_));
  INV_X1     g16481(.I(new_n16673_), .ZN(new_n16674_));
  XOR2_X1    g16482(.A1(new_n16434_), .A2(\asqrt[37] ), .Z(new_n16675_));
  NOR2_X1    g16483(.A1(\asqrt[6] ), .A2(new_n16675_), .ZN(new_n16676_));
  XOR2_X1    g16484(.A1(new_n16676_), .A2(new_n16170_), .Z(new_n16677_));
  NOR2_X1    g16485(.A1(new_n16432_), .A2(new_n16441_), .ZN(new_n16678_));
  NOR2_X1    g16486(.A1(\asqrt[6] ), .A2(new_n16678_), .ZN(new_n16679_));
  XOR2_X1    g16487(.A1(new_n16679_), .A2(new_n16173_), .Z(new_n16680_));
  AOI21_X1   g16488(.A1(new_n16436_), .A2(new_n16440_), .B(\asqrt[6] ), .ZN(new_n16681_));
  XOR2_X1    g16489(.A1(new_n16681_), .A2(new_n16176_), .Z(new_n16682_));
  INV_X1     g16490(.I(new_n16682_), .ZN(new_n16683_));
  AOI21_X1   g16491(.A1(new_n16422_), .A2(new_n16430_), .B(\asqrt[6] ), .ZN(new_n16684_));
  XOR2_X1    g16492(.A1(new_n16684_), .A2(new_n16180_), .Z(new_n16685_));
  INV_X1     g16493(.I(new_n16685_), .ZN(new_n16686_));
  XOR2_X1    g16494(.A1(new_n16413_), .A2(\asqrt[33] ), .Z(new_n16687_));
  NOR2_X1    g16495(.A1(\asqrt[6] ), .A2(new_n16687_), .ZN(new_n16688_));
  XOR2_X1    g16496(.A1(new_n16688_), .A2(new_n16182_), .Z(new_n16689_));
  NOR2_X1    g16497(.A1(new_n16411_), .A2(new_n16420_), .ZN(new_n16690_));
  NOR2_X1    g16498(.A1(\asqrt[6] ), .A2(new_n16690_), .ZN(new_n16691_));
  XOR2_X1    g16499(.A1(new_n16691_), .A2(new_n16185_), .Z(new_n16692_));
  AOI21_X1   g16500(.A1(new_n16415_), .A2(new_n16419_), .B(\asqrt[6] ), .ZN(new_n16693_));
  XOR2_X1    g16501(.A1(new_n16693_), .A2(new_n16188_), .Z(new_n16694_));
  INV_X1     g16502(.I(new_n16694_), .ZN(new_n16695_));
  AOI21_X1   g16503(.A1(new_n16401_), .A2(new_n16409_), .B(\asqrt[6] ), .ZN(new_n16696_));
  XOR2_X1    g16504(.A1(new_n16696_), .A2(new_n16192_), .Z(new_n16697_));
  INV_X1     g16505(.I(new_n16697_), .ZN(new_n16698_));
  XOR2_X1    g16506(.A1(new_n16392_), .A2(\asqrt[29] ), .Z(new_n16699_));
  NOR2_X1    g16507(.A1(\asqrt[6] ), .A2(new_n16699_), .ZN(new_n16700_));
  XOR2_X1    g16508(.A1(new_n16700_), .A2(new_n16194_), .Z(new_n16701_));
  NOR2_X1    g16509(.A1(new_n16390_), .A2(new_n16399_), .ZN(new_n16702_));
  NOR2_X1    g16510(.A1(\asqrt[6] ), .A2(new_n16702_), .ZN(new_n16703_));
  XOR2_X1    g16511(.A1(new_n16703_), .A2(new_n16197_), .Z(new_n16704_));
  AOI21_X1   g16512(.A1(new_n16394_), .A2(new_n16398_), .B(\asqrt[6] ), .ZN(new_n16705_));
  XOR2_X1    g16513(.A1(new_n16705_), .A2(new_n16200_), .Z(new_n16706_));
  INV_X1     g16514(.I(new_n16706_), .ZN(new_n16707_));
  AOI21_X1   g16515(.A1(new_n16380_), .A2(new_n16388_), .B(\asqrt[6] ), .ZN(new_n16708_));
  XOR2_X1    g16516(.A1(new_n16708_), .A2(new_n16204_), .Z(new_n16709_));
  INV_X1     g16517(.I(new_n16709_), .ZN(new_n16710_));
  XOR2_X1    g16518(.A1(new_n16371_), .A2(\asqrt[25] ), .Z(new_n16711_));
  NOR2_X1    g16519(.A1(\asqrt[6] ), .A2(new_n16711_), .ZN(new_n16712_));
  XOR2_X1    g16520(.A1(new_n16712_), .A2(new_n16206_), .Z(new_n16713_));
  NOR2_X1    g16521(.A1(new_n16369_), .A2(new_n16378_), .ZN(new_n16714_));
  NOR2_X1    g16522(.A1(\asqrt[6] ), .A2(new_n16714_), .ZN(new_n16715_));
  XOR2_X1    g16523(.A1(new_n16715_), .A2(new_n16209_), .Z(new_n16716_));
  AOI21_X1   g16524(.A1(new_n16373_), .A2(new_n16377_), .B(\asqrt[6] ), .ZN(new_n16717_));
  XOR2_X1    g16525(.A1(new_n16717_), .A2(new_n16212_), .Z(new_n16718_));
  INV_X1     g16526(.I(new_n16718_), .ZN(new_n16719_));
  AOI21_X1   g16527(.A1(new_n16359_), .A2(new_n16367_), .B(\asqrt[6] ), .ZN(new_n16720_));
  XOR2_X1    g16528(.A1(new_n16720_), .A2(new_n16216_), .Z(new_n16721_));
  INV_X1     g16529(.I(new_n16721_), .ZN(new_n16722_));
  XOR2_X1    g16530(.A1(new_n16350_), .A2(\asqrt[21] ), .Z(new_n16723_));
  NOR2_X1    g16531(.A1(\asqrt[6] ), .A2(new_n16723_), .ZN(new_n16724_));
  XOR2_X1    g16532(.A1(new_n16724_), .A2(new_n16218_), .Z(new_n16725_));
  NOR2_X1    g16533(.A1(new_n16348_), .A2(new_n16357_), .ZN(new_n16726_));
  NOR2_X1    g16534(.A1(\asqrt[6] ), .A2(new_n16726_), .ZN(new_n16727_));
  XOR2_X1    g16535(.A1(new_n16727_), .A2(new_n16221_), .Z(new_n16728_));
  AOI21_X1   g16536(.A1(new_n16352_), .A2(new_n16356_), .B(\asqrt[6] ), .ZN(new_n16729_));
  XOR2_X1    g16537(.A1(new_n16729_), .A2(new_n16224_), .Z(new_n16730_));
  INV_X1     g16538(.I(new_n16730_), .ZN(new_n16731_));
  AOI21_X1   g16539(.A1(new_n16338_), .A2(new_n16346_), .B(\asqrt[6] ), .ZN(new_n16732_));
  XOR2_X1    g16540(.A1(new_n16732_), .A2(new_n16228_), .Z(new_n16733_));
  INV_X1     g16541(.I(new_n16733_), .ZN(new_n16734_));
  XOR2_X1    g16542(.A1(new_n16329_), .A2(\asqrt[17] ), .Z(new_n16735_));
  NOR2_X1    g16543(.A1(\asqrt[6] ), .A2(new_n16735_), .ZN(new_n16736_));
  XOR2_X1    g16544(.A1(new_n16736_), .A2(new_n16230_), .Z(new_n16737_));
  NOR2_X1    g16545(.A1(new_n16327_), .A2(new_n16336_), .ZN(new_n16738_));
  NOR2_X1    g16546(.A1(\asqrt[6] ), .A2(new_n16738_), .ZN(new_n16739_));
  XOR2_X1    g16547(.A1(new_n16739_), .A2(new_n16233_), .Z(new_n16740_));
  AOI21_X1   g16548(.A1(new_n16331_), .A2(new_n16335_), .B(\asqrt[6] ), .ZN(new_n16741_));
  XOR2_X1    g16549(.A1(new_n16741_), .A2(new_n16236_), .Z(new_n16742_));
  INV_X1     g16550(.I(new_n16742_), .ZN(new_n16743_));
  AOI21_X1   g16551(.A1(new_n16317_), .A2(new_n16325_), .B(\asqrt[6] ), .ZN(new_n16744_));
  XOR2_X1    g16552(.A1(new_n16744_), .A2(new_n16240_), .Z(new_n16745_));
  INV_X1     g16553(.I(new_n16745_), .ZN(new_n16746_));
  XOR2_X1    g16554(.A1(new_n16308_), .A2(\asqrt[13] ), .Z(new_n16747_));
  NOR2_X1    g16555(.A1(\asqrt[6] ), .A2(new_n16747_), .ZN(new_n16748_));
  XOR2_X1    g16556(.A1(new_n16748_), .A2(new_n16242_), .Z(new_n16749_));
  NOR2_X1    g16557(.A1(new_n16306_), .A2(new_n16315_), .ZN(new_n16750_));
  NOR2_X1    g16558(.A1(\asqrt[6] ), .A2(new_n16750_), .ZN(new_n16751_));
  XOR2_X1    g16559(.A1(new_n16751_), .A2(new_n16245_), .Z(new_n16752_));
  AOI21_X1   g16560(.A1(new_n16310_), .A2(new_n16314_), .B(\asqrt[6] ), .ZN(new_n16753_));
  XOR2_X1    g16561(.A1(new_n16753_), .A2(new_n16248_), .Z(new_n16754_));
  INV_X1     g16562(.I(new_n16754_), .ZN(new_n16755_));
  AOI21_X1   g16563(.A1(new_n16296_), .A2(new_n16304_), .B(\asqrt[6] ), .ZN(new_n16756_));
  XOR2_X1    g16564(.A1(new_n16756_), .A2(new_n16255_), .Z(new_n16757_));
  INV_X1     g16565(.I(new_n16757_), .ZN(new_n16758_));
  AOI21_X1   g16566(.A1(new_n16287_), .A2(new_n16295_), .B(\asqrt[6] ), .ZN(new_n16759_));
  XOR2_X1    g16567(.A1(new_n16759_), .A2(new_n16272_), .Z(new_n16760_));
  NAND2_X1   g16568(.A1(\asqrt[7] ), .A2(new_n16273_), .ZN(new_n16761_));
  NOR2_X1    g16569(.A1(new_n16284_), .A2(\a[14] ), .ZN(new_n16762_));
  AOI22_X1   g16570(.A1(new_n16761_), .A2(new_n16284_), .B1(\asqrt[7] ), .B2(new_n16762_), .ZN(new_n16763_));
  AOI21_X1   g16571(.A1(\asqrt[7] ), .A2(\a[14] ), .B(new_n16281_), .ZN(new_n16764_));
  NOR2_X1    g16572(.A1(new_n16291_), .A2(new_n16764_), .ZN(new_n16765_));
  NOR2_X1    g16573(.A1(\asqrt[6] ), .A2(new_n16765_), .ZN(new_n16766_));
  XOR2_X1    g16574(.A1(new_n16766_), .A2(new_n16763_), .Z(new_n16767_));
  NAND2_X1   g16575(.A1(new_n16601_), .A2(new_n193_), .ZN(new_n16768_));
  NOR2_X1    g16576(.A1(new_n16590_), .A2(new_n16586_), .ZN(new_n16769_));
  NAND2_X1   g16577(.A1(new_n16769_), .A2(new_n201_), .ZN(new_n16770_));
  OAI21_X1   g16578(.A1(new_n16769_), .A2(new_n201_), .B(new_n16557_), .ZN(new_n16771_));
  AOI21_X1   g16579(.A1(new_n16595_), .A2(new_n16770_), .B(new_n16771_), .ZN(new_n16772_));
  NAND3_X1   g16580(.A1(new_n16607_), .A2(\asqrt[7] ), .A3(new_n16609_), .ZN(new_n16773_));
  NOR3_X1    g16581(.A1(new_n16768_), .A2(new_n16772_), .A3(new_n16773_), .ZN(new_n16774_));
  AOI21_X1   g16582(.A1(new_n16574_), .A2(new_n16571_), .B(\asqrt[62] ), .ZN(new_n16775_));
  NOR3_X1    g16583(.A1(new_n16590_), .A2(new_n201_), .A3(new_n16586_), .ZN(new_n16776_));
  OAI22_X1   g16584(.A1(new_n16775_), .A2(new_n16776_), .B1(new_n16769_), .B2(new_n16595_), .ZN(new_n16777_));
  AOI21_X1   g16585(.A1(new_n16777_), .A2(new_n16556_), .B(new_n16599_), .ZN(new_n16778_));
  NOR4_X1    g16586(.A1(new_n16778_), .A2(\asqrt[63] ), .A3(new_n16772_), .A4(new_n16610_), .ZN(new_n16779_));
  NOR2_X1    g16587(.A1(new_n16779_), .A2(new_n16276_), .ZN(new_n16780_));
  OAI21_X1   g16588(.A1(new_n16780_), .A2(new_n16774_), .B(new_n16273_), .ZN(new_n16781_));
  NOR3_X1    g16589(.A1(new_n16780_), .A2(new_n16774_), .A3(new_n16273_), .ZN(new_n16782_));
  INV_X1     g16590(.I(new_n16782_), .ZN(new_n16783_));
  NAND2_X1   g16591(.A1(new_n16783_), .A2(new_n16781_), .ZN(new_n16784_));
  NOR2_X1    g16592(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n16785_));
  INV_X1     g16593(.I(new_n16785_), .ZN(new_n16786_));
  NAND3_X1   g16594(.A1(\asqrt[6] ), .A2(\a[12] ), .A3(new_n16786_), .ZN(new_n16787_));
  INV_X1     g16595(.I(\a[12] ), .ZN(new_n16788_));
  OAI21_X1   g16596(.A1(\asqrt[6] ), .A2(new_n16788_), .B(new_n16785_), .ZN(new_n16789_));
  AOI21_X1   g16597(.A1(new_n16789_), .A2(new_n16787_), .B(new_n16269_), .ZN(new_n16790_));
  NOR3_X1    g16598(.A1(new_n16260_), .A2(\asqrt[63] ), .A3(new_n16263_), .ZN(new_n16791_));
  NAND2_X1   g16599(.A1(new_n16785_), .A2(new_n16788_), .ZN(new_n16792_));
  NAND3_X1   g16600(.A1(new_n16101_), .A2(new_n16103_), .A3(new_n16792_), .ZN(new_n16793_));
  NAND2_X1   g16601(.A1(new_n16791_), .A2(new_n16793_), .ZN(new_n16794_));
  NAND3_X1   g16602(.A1(\asqrt[6] ), .A2(\a[12] ), .A3(new_n16794_), .ZN(new_n16795_));
  INV_X1     g16603(.I(\a[13] ), .ZN(new_n16796_));
  NAND3_X1   g16604(.A1(\asqrt[6] ), .A2(new_n16788_), .A3(new_n16796_), .ZN(new_n16797_));
  OAI21_X1   g16605(.A1(new_n16779_), .A2(\a[12] ), .B(\a[13] ), .ZN(new_n16798_));
  NAND3_X1   g16606(.A1(new_n16795_), .A2(new_n16798_), .A3(new_n16797_), .ZN(new_n16799_));
  NOR3_X1    g16607(.A1(new_n16799_), .A2(new_n16790_), .A3(\asqrt[8] ), .ZN(new_n16800_));
  OAI21_X1   g16608(.A1(new_n16799_), .A2(new_n16790_), .B(\asqrt[8] ), .ZN(new_n16801_));
  OAI21_X1   g16609(.A1(new_n16784_), .A2(new_n16800_), .B(new_n16801_), .ZN(new_n16802_));
  OAI21_X1   g16610(.A1(new_n16802_), .A2(\asqrt[9] ), .B(new_n16767_), .ZN(new_n16803_));
  NAND2_X1   g16611(.A1(new_n16802_), .A2(\asqrt[9] ), .ZN(new_n16804_));
  NAND3_X1   g16612(.A1(new_n16803_), .A2(new_n16804_), .A3(new_n14690_), .ZN(new_n16805_));
  AOI21_X1   g16613(.A1(new_n16803_), .A2(new_n16804_), .B(new_n14690_), .ZN(new_n16806_));
  AOI21_X1   g16614(.A1(new_n16760_), .A2(new_n16805_), .B(new_n16806_), .ZN(new_n16807_));
  AOI21_X1   g16615(.A1(new_n16807_), .A2(new_n14207_), .B(new_n16758_), .ZN(new_n16808_));
  NAND2_X1   g16616(.A1(new_n16805_), .A2(new_n16760_), .ZN(new_n16809_));
  INV_X1     g16617(.I(new_n16767_), .ZN(new_n16810_));
  INV_X1     g16618(.I(new_n16781_), .ZN(new_n16811_));
  NOR2_X1    g16619(.A1(new_n16811_), .A2(new_n16782_), .ZN(new_n16812_));
  NOR3_X1    g16620(.A1(new_n16779_), .A2(new_n16788_), .A3(new_n16785_), .ZN(new_n16813_));
  AOI21_X1   g16621(.A1(new_n16779_), .A2(\a[12] ), .B(new_n16786_), .ZN(new_n16814_));
  OAI21_X1   g16622(.A1(new_n16813_), .A2(new_n16814_), .B(\asqrt[7] ), .ZN(new_n16815_));
  INV_X1     g16623(.I(new_n16794_), .ZN(new_n16816_));
  NOR3_X1    g16624(.A1(new_n16779_), .A2(new_n16788_), .A3(new_n16816_), .ZN(new_n16817_));
  NOR3_X1    g16625(.A1(new_n16779_), .A2(\a[12] ), .A3(\a[13] ), .ZN(new_n16818_));
  AOI21_X1   g16626(.A1(\asqrt[6] ), .A2(new_n16788_), .B(new_n16796_), .ZN(new_n16819_));
  NOR3_X1    g16627(.A1(new_n16817_), .A2(new_n16818_), .A3(new_n16819_), .ZN(new_n16820_));
  NAND3_X1   g16628(.A1(new_n16820_), .A2(new_n16815_), .A3(new_n15717_), .ZN(new_n16821_));
  AOI21_X1   g16629(.A1(new_n16820_), .A2(new_n16815_), .B(new_n15717_), .ZN(new_n16822_));
  AOI21_X1   g16630(.A1(new_n16812_), .A2(new_n16821_), .B(new_n16822_), .ZN(new_n16823_));
  AOI21_X1   g16631(.A1(new_n16823_), .A2(new_n15221_), .B(new_n16810_), .ZN(new_n16824_));
  NAND2_X1   g16632(.A1(new_n16812_), .A2(new_n16821_), .ZN(new_n16825_));
  AOI21_X1   g16633(.A1(new_n16825_), .A2(new_n16801_), .B(new_n15221_), .ZN(new_n16826_));
  OAI21_X1   g16634(.A1(new_n16824_), .A2(new_n16826_), .B(\asqrt[10] ), .ZN(new_n16827_));
  AOI21_X1   g16635(.A1(new_n16809_), .A2(new_n16827_), .B(new_n14207_), .ZN(new_n16828_));
  NOR3_X1    g16636(.A1(new_n16808_), .A2(\asqrt[12] ), .A3(new_n16828_), .ZN(new_n16829_));
  OAI21_X1   g16637(.A1(new_n16808_), .A2(new_n16828_), .B(\asqrt[12] ), .ZN(new_n16830_));
  OAI21_X1   g16638(.A1(new_n16755_), .A2(new_n16829_), .B(new_n16830_), .ZN(new_n16831_));
  OAI21_X1   g16639(.A1(new_n16831_), .A2(\asqrt[13] ), .B(new_n16752_), .ZN(new_n16832_));
  NAND2_X1   g16640(.A1(new_n16831_), .A2(\asqrt[13] ), .ZN(new_n16833_));
  NAND3_X1   g16641(.A1(new_n16832_), .A2(new_n16833_), .A3(new_n12733_), .ZN(new_n16834_));
  AOI21_X1   g16642(.A1(new_n16832_), .A2(new_n16833_), .B(new_n12733_), .ZN(new_n16835_));
  AOI21_X1   g16643(.A1(new_n16749_), .A2(new_n16834_), .B(new_n16835_), .ZN(new_n16836_));
  AOI21_X1   g16644(.A1(new_n16836_), .A2(new_n12283_), .B(new_n16746_), .ZN(new_n16837_));
  NAND2_X1   g16645(.A1(new_n16834_), .A2(new_n16749_), .ZN(new_n16838_));
  INV_X1     g16646(.I(new_n16752_), .ZN(new_n16839_));
  INV_X1     g16647(.I(new_n16760_), .ZN(new_n16840_));
  NOR3_X1    g16648(.A1(new_n16824_), .A2(\asqrt[10] ), .A3(new_n16826_), .ZN(new_n16841_));
  OAI21_X1   g16649(.A1(new_n16840_), .A2(new_n16841_), .B(new_n16827_), .ZN(new_n16842_));
  OAI21_X1   g16650(.A1(new_n16842_), .A2(\asqrt[11] ), .B(new_n16757_), .ZN(new_n16843_));
  NAND2_X1   g16651(.A1(new_n16842_), .A2(\asqrt[11] ), .ZN(new_n16844_));
  NAND3_X1   g16652(.A1(new_n16843_), .A2(new_n16844_), .A3(new_n13690_), .ZN(new_n16845_));
  AOI21_X1   g16653(.A1(new_n16843_), .A2(new_n16844_), .B(new_n13690_), .ZN(new_n16846_));
  AOI21_X1   g16654(.A1(new_n16754_), .A2(new_n16845_), .B(new_n16846_), .ZN(new_n16847_));
  AOI21_X1   g16655(.A1(new_n16847_), .A2(new_n13228_), .B(new_n16839_), .ZN(new_n16848_));
  NAND2_X1   g16656(.A1(new_n16845_), .A2(new_n16754_), .ZN(new_n16849_));
  AOI21_X1   g16657(.A1(new_n16849_), .A2(new_n16830_), .B(new_n13228_), .ZN(new_n16850_));
  OAI21_X1   g16658(.A1(new_n16848_), .A2(new_n16850_), .B(\asqrt[14] ), .ZN(new_n16851_));
  AOI21_X1   g16659(.A1(new_n16838_), .A2(new_n16851_), .B(new_n12283_), .ZN(new_n16852_));
  NOR3_X1    g16660(.A1(new_n16837_), .A2(\asqrt[16] ), .A3(new_n16852_), .ZN(new_n16853_));
  OAI21_X1   g16661(.A1(new_n16837_), .A2(new_n16852_), .B(\asqrt[16] ), .ZN(new_n16854_));
  OAI21_X1   g16662(.A1(new_n16743_), .A2(new_n16853_), .B(new_n16854_), .ZN(new_n16855_));
  OAI21_X1   g16663(.A1(new_n16855_), .A2(\asqrt[17] ), .B(new_n16740_), .ZN(new_n16856_));
  NAND2_X1   g16664(.A1(new_n16855_), .A2(\asqrt[17] ), .ZN(new_n16857_));
  NAND3_X1   g16665(.A1(new_n16856_), .A2(new_n16857_), .A3(new_n10914_), .ZN(new_n16858_));
  AOI21_X1   g16666(.A1(new_n16856_), .A2(new_n16857_), .B(new_n10914_), .ZN(new_n16859_));
  AOI21_X1   g16667(.A1(new_n16737_), .A2(new_n16858_), .B(new_n16859_), .ZN(new_n16860_));
  AOI21_X1   g16668(.A1(new_n16860_), .A2(new_n10497_), .B(new_n16734_), .ZN(new_n16861_));
  NAND2_X1   g16669(.A1(new_n16858_), .A2(new_n16737_), .ZN(new_n16862_));
  INV_X1     g16670(.I(new_n16740_), .ZN(new_n16863_));
  INV_X1     g16671(.I(new_n16749_), .ZN(new_n16864_));
  NOR3_X1    g16672(.A1(new_n16848_), .A2(\asqrt[14] ), .A3(new_n16850_), .ZN(new_n16865_));
  OAI21_X1   g16673(.A1(new_n16864_), .A2(new_n16865_), .B(new_n16851_), .ZN(new_n16866_));
  OAI21_X1   g16674(.A1(new_n16866_), .A2(\asqrt[15] ), .B(new_n16745_), .ZN(new_n16867_));
  NAND2_X1   g16675(.A1(new_n16866_), .A2(\asqrt[15] ), .ZN(new_n16868_));
  NAND3_X1   g16676(.A1(new_n16867_), .A2(new_n16868_), .A3(new_n11802_), .ZN(new_n16869_));
  AOI21_X1   g16677(.A1(new_n16867_), .A2(new_n16868_), .B(new_n11802_), .ZN(new_n16870_));
  AOI21_X1   g16678(.A1(new_n16742_), .A2(new_n16869_), .B(new_n16870_), .ZN(new_n16871_));
  AOI21_X1   g16679(.A1(new_n16871_), .A2(new_n11373_), .B(new_n16863_), .ZN(new_n16872_));
  NAND2_X1   g16680(.A1(new_n16869_), .A2(new_n16742_), .ZN(new_n16873_));
  AOI21_X1   g16681(.A1(new_n16873_), .A2(new_n16854_), .B(new_n11373_), .ZN(new_n16874_));
  OAI21_X1   g16682(.A1(new_n16872_), .A2(new_n16874_), .B(\asqrt[18] ), .ZN(new_n16875_));
  AOI21_X1   g16683(.A1(new_n16862_), .A2(new_n16875_), .B(new_n10497_), .ZN(new_n16876_));
  NOR3_X1    g16684(.A1(new_n16861_), .A2(\asqrt[20] ), .A3(new_n16876_), .ZN(new_n16877_));
  OAI21_X1   g16685(.A1(new_n16861_), .A2(new_n16876_), .B(\asqrt[20] ), .ZN(new_n16878_));
  OAI21_X1   g16686(.A1(new_n16731_), .A2(new_n16877_), .B(new_n16878_), .ZN(new_n16879_));
  OAI21_X1   g16687(.A1(new_n16879_), .A2(\asqrt[21] ), .B(new_n16728_), .ZN(new_n16880_));
  NAND2_X1   g16688(.A1(new_n16879_), .A2(\asqrt[21] ), .ZN(new_n16881_));
  NAND3_X1   g16689(.A1(new_n16880_), .A2(new_n16881_), .A3(new_n9233_), .ZN(new_n16882_));
  AOI21_X1   g16690(.A1(new_n16880_), .A2(new_n16881_), .B(new_n9233_), .ZN(new_n16883_));
  AOI21_X1   g16691(.A1(new_n16725_), .A2(new_n16882_), .B(new_n16883_), .ZN(new_n16884_));
  AOI21_X1   g16692(.A1(new_n16884_), .A2(new_n8849_), .B(new_n16722_), .ZN(new_n16885_));
  NAND2_X1   g16693(.A1(new_n16882_), .A2(new_n16725_), .ZN(new_n16886_));
  INV_X1     g16694(.I(new_n16728_), .ZN(new_n16887_));
  INV_X1     g16695(.I(new_n16737_), .ZN(new_n16888_));
  NOR3_X1    g16696(.A1(new_n16872_), .A2(\asqrt[18] ), .A3(new_n16874_), .ZN(new_n16889_));
  OAI21_X1   g16697(.A1(new_n16888_), .A2(new_n16889_), .B(new_n16875_), .ZN(new_n16890_));
  OAI21_X1   g16698(.A1(new_n16890_), .A2(\asqrt[19] ), .B(new_n16733_), .ZN(new_n16891_));
  NAND2_X1   g16699(.A1(new_n16890_), .A2(\asqrt[19] ), .ZN(new_n16892_));
  NAND3_X1   g16700(.A1(new_n16891_), .A2(new_n16892_), .A3(new_n10052_), .ZN(new_n16893_));
  AOI21_X1   g16701(.A1(new_n16891_), .A2(new_n16892_), .B(new_n10052_), .ZN(new_n16894_));
  AOI21_X1   g16702(.A1(new_n16730_), .A2(new_n16893_), .B(new_n16894_), .ZN(new_n16895_));
  AOI21_X1   g16703(.A1(new_n16895_), .A2(new_n9656_), .B(new_n16887_), .ZN(new_n16896_));
  NAND2_X1   g16704(.A1(new_n16893_), .A2(new_n16730_), .ZN(new_n16897_));
  AOI21_X1   g16705(.A1(new_n16897_), .A2(new_n16878_), .B(new_n9656_), .ZN(new_n16898_));
  OAI21_X1   g16706(.A1(new_n16896_), .A2(new_n16898_), .B(\asqrt[22] ), .ZN(new_n16899_));
  AOI21_X1   g16707(.A1(new_n16886_), .A2(new_n16899_), .B(new_n8849_), .ZN(new_n16900_));
  NOR3_X1    g16708(.A1(new_n16885_), .A2(\asqrt[24] ), .A3(new_n16900_), .ZN(new_n16901_));
  OAI21_X1   g16709(.A1(new_n16885_), .A2(new_n16900_), .B(\asqrt[24] ), .ZN(new_n16902_));
  OAI21_X1   g16710(.A1(new_n16719_), .A2(new_n16901_), .B(new_n16902_), .ZN(new_n16903_));
  OAI21_X1   g16711(.A1(new_n16903_), .A2(\asqrt[25] ), .B(new_n16716_), .ZN(new_n16904_));
  NAND2_X1   g16712(.A1(new_n16903_), .A2(\asqrt[25] ), .ZN(new_n16905_));
  NAND3_X1   g16713(.A1(new_n16904_), .A2(new_n16905_), .A3(new_n7690_), .ZN(new_n16906_));
  AOI21_X1   g16714(.A1(new_n16904_), .A2(new_n16905_), .B(new_n7690_), .ZN(new_n16907_));
  AOI21_X1   g16715(.A1(new_n16713_), .A2(new_n16906_), .B(new_n16907_), .ZN(new_n16908_));
  AOI21_X1   g16716(.A1(new_n16908_), .A2(new_n7331_), .B(new_n16710_), .ZN(new_n16909_));
  NAND2_X1   g16717(.A1(new_n16906_), .A2(new_n16713_), .ZN(new_n16910_));
  INV_X1     g16718(.I(new_n16716_), .ZN(new_n16911_));
  INV_X1     g16719(.I(new_n16725_), .ZN(new_n16912_));
  NOR3_X1    g16720(.A1(new_n16896_), .A2(\asqrt[22] ), .A3(new_n16898_), .ZN(new_n16913_));
  OAI21_X1   g16721(.A1(new_n16912_), .A2(new_n16913_), .B(new_n16899_), .ZN(new_n16914_));
  OAI21_X1   g16722(.A1(new_n16914_), .A2(\asqrt[23] ), .B(new_n16721_), .ZN(new_n16915_));
  NAND2_X1   g16723(.A1(new_n16914_), .A2(\asqrt[23] ), .ZN(new_n16916_));
  NAND3_X1   g16724(.A1(new_n16915_), .A2(new_n16916_), .A3(new_n8440_), .ZN(new_n16917_));
  AOI21_X1   g16725(.A1(new_n16915_), .A2(new_n16916_), .B(new_n8440_), .ZN(new_n16918_));
  AOI21_X1   g16726(.A1(new_n16718_), .A2(new_n16917_), .B(new_n16918_), .ZN(new_n16919_));
  AOI21_X1   g16727(.A1(new_n16919_), .A2(new_n8077_), .B(new_n16911_), .ZN(new_n16920_));
  NAND2_X1   g16728(.A1(new_n16917_), .A2(new_n16718_), .ZN(new_n16921_));
  AOI21_X1   g16729(.A1(new_n16921_), .A2(new_n16902_), .B(new_n8077_), .ZN(new_n16922_));
  OAI21_X1   g16730(.A1(new_n16920_), .A2(new_n16922_), .B(\asqrt[26] ), .ZN(new_n16923_));
  AOI21_X1   g16731(.A1(new_n16910_), .A2(new_n16923_), .B(new_n7331_), .ZN(new_n16924_));
  NOR3_X1    g16732(.A1(new_n16909_), .A2(\asqrt[28] ), .A3(new_n16924_), .ZN(new_n16925_));
  OAI21_X1   g16733(.A1(new_n16909_), .A2(new_n16924_), .B(\asqrt[28] ), .ZN(new_n16926_));
  OAI21_X1   g16734(.A1(new_n16707_), .A2(new_n16925_), .B(new_n16926_), .ZN(new_n16927_));
  OAI21_X1   g16735(.A1(new_n16927_), .A2(\asqrt[29] ), .B(new_n16704_), .ZN(new_n16928_));
  NAND2_X1   g16736(.A1(new_n16927_), .A2(\asqrt[29] ), .ZN(new_n16929_));
  NAND3_X1   g16737(.A1(new_n16928_), .A2(new_n16929_), .A3(new_n6275_), .ZN(new_n16930_));
  AOI21_X1   g16738(.A1(new_n16928_), .A2(new_n16929_), .B(new_n6275_), .ZN(new_n16931_));
  AOI21_X1   g16739(.A1(new_n16701_), .A2(new_n16930_), .B(new_n16931_), .ZN(new_n16932_));
  AOI21_X1   g16740(.A1(new_n16932_), .A2(new_n5947_), .B(new_n16698_), .ZN(new_n16933_));
  NAND2_X1   g16741(.A1(new_n16930_), .A2(new_n16701_), .ZN(new_n16934_));
  INV_X1     g16742(.I(new_n16704_), .ZN(new_n16935_));
  INV_X1     g16743(.I(new_n16713_), .ZN(new_n16936_));
  NOR3_X1    g16744(.A1(new_n16920_), .A2(\asqrt[26] ), .A3(new_n16922_), .ZN(new_n16937_));
  OAI21_X1   g16745(.A1(new_n16936_), .A2(new_n16937_), .B(new_n16923_), .ZN(new_n16938_));
  OAI21_X1   g16746(.A1(new_n16938_), .A2(\asqrt[27] ), .B(new_n16709_), .ZN(new_n16939_));
  NAND2_X1   g16747(.A1(new_n16938_), .A2(\asqrt[27] ), .ZN(new_n16940_));
  NAND3_X1   g16748(.A1(new_n16939_), .A2(new_n16940_), .A3(new_n6966_), .ZN(new_n16941_));
  AOI21_X1   g16749(.A1(new_n16939_), .A2(new_n16940_), .B(new_n6966_), .ZN(new_n16942_));
  AOI21_X1   g16750(.A1(new_n16706_), .A2(new_n16941_), .B(new_n16942_), .ZN(new_n16943_));
  AOI21_X1   g16751(.A1(new_n16943_), .A2(new_n6636_), .B(new_n16935_), .ZN(new_n16944_));
  NAND2_X1   g16752(.A1(new_n16941_), .A2(new_n16706_), .ZN(new_n16945_));
  AOI21_X1   g16753(.A1(new_n16945_), .A2(new_n16926_), .B(new_n6636_), .ZN(new_n16946_));
  OAI21_X1   g16754(.A1(new_n16944_), .A2(new_n16946_), .B(\asqrt[30] ), .ZN(new_n16947_));
  AOI21_X1   g16755(.A1(new_n16934_), .A2(new_n16947_), .B(new_n5947_), .ZN(new_n16948_));
  NOR3_X1    g16756(.A1(new_n16933_), .A2(\asqrt[32] ), .A3(new_n16948_), .ZN(new_n16949_));
  OAI21_X1   g16757(.A1(new_n16933_), .A2(new_n16948_), .B(\asqrt[32] ), .ZN(new_n16950_));
  OAI21_X1   g16758(.A1(new_n16695_), .A2(new_n16949_), .B(new_n16950_), .ZN(new_n16951_));
  OAI21_X1   g16759(.A1(new_n16951_), .A2(\asqrt[33] ), .B(new_n16692_), .ZN(new_n16952_));
  NAND2_X1   g16760(.A1(new_n16951_), .A2(\asqrt[33] ), .ZN(new_n16953_));
  NAND3_X1   g16761(.A1(new_n16952_), .A2(new_n16953_), .A3(new_n5029_), .ZN(new_n16954_));
  AOI21_X1   g16762(.A1(new_n16952_), .A2(new_n16953_), .B(new_n5029_), .ZN(new_n16955_));
  AOI21_X1   g16763(.A1(new_n16689_), .A2(new_n16954_), .B(new_n16955_), .ZN(new_n16956_));
  AOI21_X1   g16764(.A1(new_n16956_), .A2(new_n4751_), .B(new_n16686_), .ZN(new_n16957_));
  NAND2_X1   g16765(.A1(new_n16954_), .A2(new_n16689_), .ZN(new_n16958_));
  INV_X1     g16766(.I(new_n16692_), .ZN(new_n16959_));
  INV_X1     g16767(.I(new_n16701_), .ZN(new_n16960_));
  NOR3_X1    g16768(.A1(new_n16944_), .A2(\asqrt[30] ), .A3(new_n16946_), .ZN(new_n16961_));
  OAI21_X1   g16769(.A1(new_n16960_), .A2(new_n16961_), .B(new_n16947_), .ZN(new_n16962_));
  OAI21_X1   g16770(.A1(new_n16962_), .A2(\asqrt[31] ), .B(new_n16697_), .ZN(new_n16963_));
  NAND2_X1   g16771(.A1(new_n16962_), .A2(\asqrt[31] ), .ZN(new_n16964_));
  NAND3_X1   g16772(.A1(new_n16963_), .A2(new_n16964_), .A3(new_n5643_), .ZN(new_n16965_));
  AOI21_X1   g16773(.A1(new_n16963_), .A2(new_n16964_), .B(new_n5643_), .ZN(new_n16966_));
  AOI21_X1   g16774(.A1(new_n16694_), .A2(new_n16965_), .B(new_n16966_), .ZN(new_n16967_));
  AOI21_X1   g16775(.A1(new_n16967_), .A2(new_n5336_), .B(new_n16959_), .ZN(new_n16968_));
  NAND2_X1   g16776(.A1(new_n16965_), .A2(new_n16694_), .ZN(new_n16969_));
  AOI21_X1   g16777(.A1(new_n16969_), .A2(new_n16950_), .B(new_n5336_), .ZN(new_n16970_));
  OAI21_X1   g16778(.A1(new_n16968_), .A2(new_n16970_), .B(\asqrt[34] ), .ZN(new_n16971_));
  AOI21_X1   g16779(.A1(new_n16958_), .A2(new_n16971_), .B(new_n4751_), .ZN(new_n16972_));
  NOR3_X1    g16780(.A1(new_n16957_), .A2(\asqrt[36] ), .A3(new_n16972_), .ZN(new_n16973_));
  OAI21_X1   g16781(.A1(new_n16957_), .A2(new_n16972_), .B(\asqrt[36] ), .ZN(new_n16974_));
  OAI21_X1   g16782(.A1(new_n16683_), .A2(new_n16973_), .B(new_n16974_), .ZN(new_n16975_));
  OAI21_X1   g16783(.A1(new_n16975_), .A2(\asqrt[37] ), .B(new_n16680_), .ZN(new_n16976_));
  NAND2_X1   g16784(.A1(new_n16975_), .A2(\asqrt[37] ), .ZN(new_n16977_));
  NAND3_X1   g16785(.A1(new_n16976_), .A2(new_n16977_), .A3(new_n3925_), .ZN(new_n16978_));
  AOI21_X1   g16786(.A1(new_n16976_), .A2(new_n16977_), .B(new_n3925_), .ZN(new_n16979_));
  AOI21_X1   g16787(.A1(new_n16677_), .A2(new_n16978_), .B(new_n16979_), .ZN(new_n16980_));
  AOI21_X1   g16788(.A1(new_n16980_), .A2(new_n3681_), .B(new_n16674_), .ZN(new_n16981_));
  NAND2_X1   g16789(.A1(new_n16978_), .A2(new_n16677_), .ZN(new_n16982_));
  INV_X1     g16790(.I(new_n16680_), .ZN(new_n16983_));
  INV_X1     g16791(.I(new_n16689_), .ZN(new_n16984_));
  NOR3_X1    g16792(.A1(new_n16968_), .A2(\asqrt[34] ), .A3(new_n16970_), .ZN(new_n16985_));
  OAI21_X1   g16793(.A1(new_n16984_), .A2(new_n16985_), .B(new_n16971_), .ZN(new_n16986_));
  OAI21_X1   g16794(.A1(new_n16986_), .A2(\asqrt[35] ), .B(new_n16685_), .ZN(new_n16987_));
  NAND2_X1   g16795(.A1(new_n16986_), .A2(\asqrt[35] ), .ZN(new_n16988_));
  NAND3_X1   g16796(.A1(new_n16987_), .A2(new_n16988_), .A3(new_n4461_), .ZN(new_n16989_));
  AOI21_X1   g16797(.A1(new_n16987_), .A2(new_n16988_), .B(new_n4461_), .ZN(new_n16990_));
  AOI21_X1   g16798(.A1(new_n16682_), .A2(new_n16989_), .B(new_n16990_), .ZN(new_n16991_));
  AOI21_X1   g16799(.A1(new_n16991_), .A2(new_n4196_), .B(new_n16983_), .ZN(new_n16992_));
  NAND2_X1   g16800(.A1(new_n16989_), .A2(new_n16682_), .ZN(new_n16993_));
  AOI21_X1   g16801(.A1(new_n16993_), .A2(new_n16974_), .B(new_n4196_), .ZN(new_n16994_));
  OAI21_X1   g16802(.A1(new_n16992_), .A2(new_n16994_), .B(\asqrt[38] ), .ZN(new_n16995_));
  AOI21_X1   g16803(.A1(new_n16982_), .A2(new_n16995_), .B(new_n3681_), .ZN(new_n16996_));
  NOR3_X1    g16804(.A1(new_n16981_), .A2(\asqrt[40] ), .A3(new_n16996_), .ZN(new_n16997_));
  OAI21_X1   g16805(.A1(new_n16981_), .A2(new_n16996_), .B(\asqrt[40] ), .ZN(new_n16998_));
  OAI21_X1   g16806(.A1(new_n16671_), .A2(new_n16997_), .B(new_n16998_), .ZN(new_n16999_));
  OAI21_X1   g16807(.A1(new_n16999_), .A2(\asqrt[41] ), .B(new_n16668_), .ZN(new_n17000_));
  NAND2_X1   g16808(.A1(new_n16999_), .A2(\asqrt[41] ), .ZN(new_n17001_));
  NAND3_X1   g16809(.A1(new_n17000_), .A2(new_n17001_), .A3(new_n2960_), .ZN(new_n17002_));
  AOI21_X1   g16810(.A1(new_n17000_), .A2(new_n17001_), .B(new_n2960_), .ZN(new_n17003_));
  AOI21_X1   g16811(.A1(new_n16665_), .A2(new_n17002_), .B(new_n17003_), .ZN(new_n17004_));
  AOI21_X1   g16812(.A1(new_n17004_), .A2(new_n2749_), .B(new_n16662_), .ZN(new_n17005_));
  NAND2_X1   g16813(.A1(new_n17002_), .A2(new_n16665_), .ZN(new_n17006_));
  INV_X1     g16814(.I(new_n16668_), .ZN(new_n17007_));
  INV_X1     g16815(.I(new_n16677_), .ZN(new_n17008_));
  NOR3_X1    g16816(.A1(new_n16992_), .A2(\asqrt[38] ), .A3(new_n16994_), .ZN(new_n17009_));
  OAI21_X1   g16817(.A1(new_n17008_), .A2(new_n17009_), .B(new_n16995_), .ZN(new_n17010_));
  OAI21_X1   g16818(.A1(new_n17010_), .A2(\asqrt[39] ), .B(new_n16673_), .ZN(new_n17011_));
  NAND2_X1   g16819(.A1(new_n17010_), .A2(\asqrt[39] ), .ZN(new_n17012_));
  NAND3_X1   g16820(.A1(new_n17011_), .A2(new_n17012_), .A3(new_n3427_), .ZN(new_n17013_));
  AOI21_X1   g16821(.A1(new_n17011_), .A2(new_n17012_), .B(new_n3427_), .ZN(new_n17014_));
  AOI21_X1   g16822(.A1(new_n16670_), .A2(new_n17013_), .B(new_n17014_), .ZN(new_n17015_));
  AOI21_X1   g16823(.A1(new_n17015_), .A2(new_n3195_), .B(new_n17007_), .ZN(new_n17016_));
  NAND2_X1   g16824(.A1(new_n17013_), .A2(new_n16670_), .ZN(new_n17017_));
  AOI21_X1   g16825(.A1(new_n17017_), .A2(new_n16998_), .B(new_n3195_), .ZN(new_n17018_));
  OAI21_X1   g16826(.A1(new_n17016_), .A2(new_n17018_), .B(\asqrt[42] ), .ZN(new_n17019_));
  AOI21_X1   g16827(.A1(new_n17006_), .A2(new_n17019_), .B(new_n2749_), .ZN(new_n17020_));
  NOR3_X1    g16828(.A1(new_n17005_), .A2(\asqrt[44] ), .A3(new_n17020_), .ZN(new_n17021_));
  OAI21_X1   g16829(.A1(new_n17005_), .A2(new_n17020_), .B(\asqrt[44] ), .ZN(new_n17022_));
  OAI21_X1   g16830(.A1(new_n16659_), .A2(new_n17021_), .B(new_n17022_), .ZN(new_n17023_));
  OAI21_X1   g16831(.A1(new_n17023_), .A2(\asqrt[45] ), .B(new_n16656_), .ZN(new_n17024_));
  NAND2_X1   g16832(.A1(new_n17023_), .A2(\asqrt[45] ), .ZN(new_n17025_));
  NAND3_X1   g16833(.A1(new_n17024_), .A2(new_n17025_), .A3(new_n2134_), .ZN(new_n17026_));
  AOI21_X1   g16834(.A1(new_n17024_), .A2(new_n17025_), .B(new_n2134_), .ZN(new_n17027_));
  AOI21_X1   g16835(.A1(new_n16653_), .A2(new_n17026_), .B(new_n17027_), .ZN(new_n17028_));
  AOI21_X1   g16836(.A1(new_n17028_), .A2(new_n1953_), .B(new_n16650_), .ZN(new_n17029_));
  NAND2_X1   g16837(.A1(new_n17026_), .A2(new_n16653_), .ZN(new_n17030_));
  INV_X1     g16838(.I(new_n16656_), .ZN(new_n17031_));
  INV_X1     g16839(.I(new_n16665_), .ZN(new_n17032_));
  NOR3_X1    g16840(.A1(new_n17016_), .A2(\asqrt[42] ), .A3(new_n17018_), .ZN(new_n17033_));
  OAI21_X1   g16841(.A1(new_n17032_), .A2(new_n17033_), .B(new_n17019_), .ZN(new_n17034_));
  OAI21_X1   g16842(.A1(new_n17034_), .A2(\asqrt[43] ), .B(new_n16661_), .ZN(new_n17035_));
  NAND2_X1   g16843(.A1(new_n17034_), .A2(\asqrt[43] ), .ZN(new_n17036_));
  NAND3_X1   g16844(.A1(new_n17035_), .A2(new_n17036_), .A3(new_n2531_), .ZN(new_n17037_));
  AOI21_X1   g16845(.A1(new_n17035_), .A2(new_n17036_), .B(new_n2531_), .ZN(new_n17038_));
  AOI21_X1   g16846(.A1(new_n16658_), .A2(new_n17037_), .B(new_n17038_), .ZN(new_n17039_));
  AOI21_X1   g16847(.A1(new_n17039_), .A2(new_n2332_), .B(new_n17031_), .ZN(new_n17040_));
  NAND2_X1   g16848(.A1(new_n17037_), .A2(new_n16658_), .ZN(new_n17041_));
  AOI21_X1   g16849(.A1(new_n17041_), .A2(new_n17022_), .B(new_n2332_), .ZN(new_n17042_));
  OAI21_X1   g16850(.A1(new_n17040_), .A2(new_n17042_), .B(\asqrt[46] ), .ZN(new_n17043_));
  AOI21_X1   g16851(.A1(new_n17030_), .A2(new_n17043_), .B(new_n1953_), .ZN(new_n17044_));
  NOR3_X1    g16852(.A1(new_n17029_), .A2(\asqrt[48] ), .A3(new_n17044_), .ZN(new_n17045_));
  OAI21_X1   g16853(.A1(new_n17029_), .A2(new_n17044_), .B(\asqrt[48] ), .ZN(new_n17046_));
  OAI21_X1   g16854(.A1(new_n16647_), .A2(new_n17045_), .B(new_n17046_), .ZN(new_n17047_));
  OAI21_X1   g16855(.A1(new_n17047_), .A2(\asqrt[49] ), .B(new_n16644_), .ZN(new_n17048_));
  NAND2_X1   g16856(.A1(new_n17047_), .A2(\asqrt[49] ), .ZN(new_n17049_));
  NAND3_X1   g16857(.A1(new_n17048_), .A2(new_n17049_), .A3(new_n1463_), .ZN(new_n17050_));
  AOI21_X1   g16858(.A1(new_n17048_), .A2(new_n17049_), .B(new_n1463_), .ZN(new_n17051_));
  AOI21_X1   g16859(.A1(new_n16641_), .A2(new_n17050_), .B(new_n17051_), .ZN(new_n17052_));
  AOI21_X1   g16860(.A1(new_n17052_), .A2(new_n1305_), .B(new_n16638_), .ZN(new_n17053_));
  NAND2_X1   g16861(.A1(new_n17050_), .A2(new_n16641_), .ZN(new_n17054_));
  INV_X1     g16862(.I(new_n16644_), .ZN(new_n17055_));
  INV_X1     g16863(.I(new_n16653_), .ZN(new_n17056_));
  NOR3_X1    g16864(.A1(new_n17040_), .A2(\asqrt[46] ), .A3(new_n17042_), .ZN(new_n17057_));
  OAI21_X1   g16865(.A1(new_n17056_), .A2(new_n17057_), .B(new_n17043_), .ZN(new_n17058_));
  OAI21_X1   g16866(.A1(new_n17058_), .A2(\asqrt[47] ), .B(new_n16649_), .ZN(new_n17059_));
  NAND2_X1   g16867(.A1(new_n17058_), .A2(\asqrt[47] ), .ZN(new_n17060_));
  NAND3_X1   g16868(.A1(new_n17059_), .A2(new_n17060_), .A3(new_n1778_), .ZN(new_n17061_));
  AOI21_X1   g16869(.A1(new_n17059_), .A2(new_n17060_), .B(new_n1778_), .ZN(new_n17062_));
  AOI21_X1   g16870(.A1(new_n16646_), .A2(new_n17061_), .B(new_n17062_), .ZN(new_n17063_));
  AOI21_X1   g16871(.A1(new_n17063_), .A2(new_n1632_), .B(new_n17055_), .ZN(new_n17064_));
  NAND2_X1   g16872(.A1(new_n17061_), .A2(new_n16646_), .ZN(new_n17065_));
  AOI21_X1   g16873(.A1(new_n17065_), .A2(new_n17046_), .B(new_n1632_), .ZN(new_n17066_));
  OAI21_X1   g16874(.A1(new_n17064_), .A2(new_n17066_), .B(\asqrt[50] ), .ZN(new_n17067_));
  AOI21_X1   g16875(.A1(new_n17054_), .A2(new_n17067_), .B(new_n1305_), .ZN(new_n17068_));
  NOR3_X1    g16876(.A1(new_n17053_), .A2(\asqrt[52] ), .A3(new_n17068_), .ZN(new_n17069_));
  OAI21_X1   g16877(.A1(new_n17053_), .A2(new_n17068_), .B(\asqrt[52] ), .ZN(new_n17070_));
  OAI21_X1   g16878(.A1(new_n16635_), .A2(new_n17069_), .B(new_n17070_), .ZN(new_n17071_));
  OAI21_X1   g16879(.A1(new_n17071_), .A2(\asqrt[53] ), .B(new_n16632_), .ZN(new_n17072_));
  NAND2_X1   g16880(.A1(new_n17071_), .A2(\asqrt[53] ), .ZN(new_n17073_));
  NAND3_X1   g16881(.A1(new_n17072_), .A2(new_n17073_), .A3(new_n860_), .ZN(new_n17074_));
  AOI21_X1   g16882(.A1(new_n17072_), .A2(new_n17073_), .B(new_n860_), .ZN(new_n17075_));
  AOI21_X1   g16883(.A1(new_n16629_), .A2(new_n17074_), .B(new_n17075_), .ZN(new_n17076_));
  AOI21_X1   g16884(.A1(new_n17076_), .A2(new_n744_), .B(new_n16626_), .ZN(new_n17077_));
  NAND2_X1   g16885(.A1(new_n17074_), .A2(new_n16629_), .ZN(new_n17078_));
  INV_X1     g16886(.I(new_n16632_), .ZN(new_n17079_));
  INV_X1     g16887(.I(new_n16641_), .ZN(new_n17080_));
  NOR3_X1    g16888(.A1(new_n17064_), .A2(\asqrt[50] ), .A3(new_n17066_), .ZN(new_n17081_));
  OAI21_X1   g16889(.A1(new_n17080_), .A2(new_n17081_), .B(new_n17067_), .ZN(new_n17082_));
  OAI21_X1   g16890(.A1(new_n17082_), .A2(\asqrt[51] ), .B(new_n16637_), .ZN(new_n17083_));
  NAND2_X1   g16891(.A1(new_n17082_), .A2(\asqrt[51] ), .ZN(new_n17084_));
  NAND3_X1   g16892(.A1(new_n17083_), .A2(new_n17084_), .A3(new_n1150_), .ZN(new_n17085_));
  AOI21_X1   g16893(.A1(new_n17083_), .A2(new_n17084_), .B(new_n1150_), .ZN(new_n17086_));
  AOI21_X1   g16894(.A1(new_n16634_), .A2(new_n17085_), .B(new_n17086_), .ZN(new_n17087_));
  AOI21_X1   g16895(.A1(new_n17087_), .A2(new_n1006_), .B(new_n17079_), .ZN(new_n17088_));
  NAND2_X1   g16896(.A1(new_n17085_), .A2(new_n16634_), .ZN(new_n17089_));
  AOI21_X1   g16897(.A1(new_n17089_), .A2(new_n17070_), .B(new_n1006_), .ZN(new_n17090_));
  OAI21_X1   g16898(.A1(new_n17088_), .A2(new_n17090_), .B(\asqrt[54] ), .ZN(new_n17091_));
  AOI21_X1   g16899(.A1(new_n17078_), .A2(new_n17091_), .B(new_n744_), .ZN(new_n17092_));
  NOR3_X1    g16900(.A1(new_n17077_), .A2(\asqrt[56] ), .A3(new_n17092_), .ZN(new_n17093_));
  OAI21_X1   g16901(.A1(new_n17077_), .A2(new_n17092_), .B(\asqrt[56] ), .ZN(new_n17094_));
  OAI21_X1   g16902(.A1(new_n16623_), .A2(new_n17093_), .B(new_n17094_), .ZN(new_n17095_));
  OAI21_X1   g16903(.A1(new_n17095_), .A2(\asqrt[57] ), .B(new_n16620_), .ZN(new_n17096_));
  NAND2_X1   g16904(.A1(new_n17095_), .A2(\asqrt[57] ), .ZN(new_n17097_));
  NAND3_X1   g16905(.A1(new_n17096_), .A2(new_n17097_), .A3(new_n423_), .ZN(new_n17098_));
  AOI21_X1   g16906(.A1(new_n17096_), .A2(new_n17097_), .B(new_n423_), .ZN(new_n17099_));
  AOI21_X1   g16907(.A1(new_n16617_), .A2(new_n17098_), .B(new_n17099_), .ZN(new_n17100_));
  NAND2_X1   g16908(.A1(new_n17100_), .A2(new_n337_), .ZN(new_n17101_));
  INV_X1     g16909(.I(new_n16617_), .ZN(new_n17102_));
  INV_X1     g16910(.I(new_n16620_), .ZN(new_n17103_));
  INV_X1     g16911(.I(new_n16629_), .ZN(new_n17104_));
  NOR3_X1    g16912(.A1(new_n17088_), .A2(\asqrt[54] ), .A3(new_n17090_), .ZN(new_n17105_));
  OAI21_X1   g16913(.A1(new_n17104_), .A2(new_n17105_), .B(new_n17091_), .ZN(new_n17106_));
  OAI21_X1   g16914(.A1(new_n17106_), .A2(\asqrt[55] ), .B(new_n16625_), .ZN(new_n17107_));
  NAND2_X1   g16915(.A1(new_n17106_), .A2(\asqrt[55] ), .ZN(new_n17108_));
  NAND3_X1   g16916(.A1(new_n17107_), .A2(new_n17108_), .A3(new_n634_), .ZN(new_n17109_));
  AOI21_X1   g16917(.A1(new_n17107_), .A2(new_n17108_), .B(new_n634_), .ZN(new_n17110_));
  AOI21_X1   g16918(.A1(new_n16622_), .A2(new_n17109_), .B(new_n17110_), .ZN(new_n17111_));
  AOI21_X1   g16919(.A1(new_n17111_), .A2(new_n531_), .B(new_n17103_), .ZN(new_n17112_));
  NAND2_X1   g16920(.A1(new_n17109_), .A2(new_n16622_), .ZN(new_n17113_));
  AOI21_X1   g16921(.A1(new_n17113_), .A2(new_n17094_), .B(new_n531_), .ZN(new_n17114_));
  NOR3_X1    g16922(.A1(new_n17112_), .A2(\asqrt[58] ), .A3(new_n17114_), .ZN(new_n17115_));
  NOR2_X1    g16923(.A1(new_n17115_), .A2(new_n17102_), .ZN(new_n17116_));
  OAI21_X1   g16924(.A1(new_n17116_), .A2(new_n17099_), .B(\asqrt[59] ), .ZN(new_n17117_));
  NOR2_X1    g16925(.A1(\asqrt[6] ), .A2(new_n16557_), .ZN(new_n17118_));
  NOR2_X1    g16926(.A1(new_n16777_), .A2(new_n16557_), .ZN(new_n17119_));
  NOR2_X1    g16927(.A1(new_n16597_), .A2(new_n16556_), .ZN(new_n17120_));
  OAI21_X1   g16928(.A1(new_n17120_), .A2(new_n17119_), .B(\asqrt[63] ), .ZN(new_n17121_));
  NOR2_X1    g16929(.A1(new_n17118_), .A2(new_n17121_), .ZN(new_n17122_));
  INV_X1     g16930(.I(new_n17122_), .ZN(new_n17123_));
  AOI21_X1   g16931(.A1(new_n16770_), .A2(new_n16603_), .B(\asqrt[6] ), .ZN(new_n17124_));
  XOR2_X1    g16932(.A1(new_n17124_), .A2(new_n16595_), .Z(new_n17125_));
  INV_X1     g16933(.I(new_n17125_), .ZN(new_n17126_));
  AOI21_X1   g16934(.A1(new_n16578_), .A2(new_n16583_), .B(\asqrt[6] ), .ZN(new_n17127_));
  XOR2_X1    g16935(.A1(new_n17127_), .A2(new_n16562_), .Z(new_n17128_));
  INV_X1     g16936(.I(new_n17128_), .ZN(new_n17129_));
  INV_X1     g16937(.I(new_n16614_), .ZN(new_n17130_));
  AOI21_X1   g16938(.A1(new_n17100_), .A2(new_n337_), .B(new_n17130_), .ZN(new_n17131_));
  NAND2_X1   g16939(.A1(new_n17098_), .A2(new_n16617_), .ZN(new_n17132_));
  OAI21_X1   g16940(.A1(new_n17112_), .A2(new_n17114_), .B(\asqrt[58] ), .ZN(new_n17133_));
  AOI21_X1   g16941(.A1(new_n17132_), .A2(new_n17133_), .B(new_n337_), .ZN(new_n17134_));
  NOR3_X1    g16942(.A1(new_n17131_), .A2(\asqrt[60] ), .A3(new_n17134_), .ZN(new_n17135_));
  NOR2_X1    g16943(.A1(new_n17135_), .A2(new_n17129_), .ZN(new_n17136_));
  OAI21_X1   g16944(.A1(new_n17102_), .A2(new_n17115_), .B(new_n17133_), .ZN(new_n17137_));
  OAI21_X1   g16945(.A1(new_n17137_), .A2(\asqrt[59] ), .B(new_n16614_), .ZN(new_n17138_));
  AOI21_X1   g16946(.A1(new_n17138_), .A2(new_n17117_), .B(new_n266_), .ZN(new_n17139_));
  OAI21_X1   g16947(.A1(new_n17136_), .A2(new_n17139_), .B(\asqrt[61] ), .ZN(new_n17140_));
  OAI21_X1   g16948(.A1(new_n17131_), .A2(new_n17134_), .B(\asqrt[60] ), .ZN(new_n17141_));
  OAI21_X1   g16949(.A1(new_n17129_), .A2(new_n17135_), .B(new_n17141_), .ZN(new_n17142_));
  AOI21_X1   g16950(.A1(new_n16584_), .A2(new_n16569_), .B(\asqrt[6] ), .ZN(new_n17143_));
  XOR2_X1    g16951(.A1(new_n17143_), .A2(new_n16559_), .Z(new_n17144_));
  OAI21_X1   g16952(.A1(new_n17142_), .A2(\asqrt[61] ), .B(new_n17144_), .ZN(new_n17145_));
  NAND2_X1   g16953(.A1(new_n17145_), .A2(new_n17140_), .ZN(new_n17146_));
  NAND3_X1   g16954(.A1(new_n17138_), .A2(new_n266_), .A3(new_n17117_), .ZN(new_n17147_));
  NAND2_X1   g16955(.A1(new_n17147_), .A2(new_n17128_), .ZN(new_n17148_));
  AOI21_X1   g16956(.A1(new_n17148_), .A2(new_n17141_), .B(new_n239_), .ZN(new_n17149_));
  AOI21_X1   g16957(.A1(new_n17128_), .A2(new_n17147_), .B(new_n17139_), .ZN(new_n17150_));
  INV_X1     g16958(.I(new_n17144_), .ZN(new_n17151_));
  AOI21_X1   g16959(.A1(new_n17150_), .A2(new_n239_), .B(new_n17151_), .ZN(new_n17152_));
  OAI21_X1   g16960(.A1(new_n17152_), .A2(new_n17149_), .B(new_n201_), .ZN(new_n17153_));
  NAND3_X1   g16961(.A1(new_n17145_), .A2(\asqrt[62] ), .A3(new_n17140_), .ZN(new_n17154_));
  NAND2_X1   g16962(.A1(new_n16588_), .A2(new_n239_), .ZN(new_n17155_));
  AOI21_X1   g16963(.A1(new_n16571_), .A2(new_n17155_), .B(\asqrt[6] ), .ZN(new_n17156_));
  XOR2_X1    g16964(.A1(new_n17156_), .A2(new_n16573_), .Z(new_n17157_));
  INV_X1     g16965(.I(new_n17157_), .ZN(new_n17158_));
  AOI22_X1   g16966(.A1(new_n17153_), .A2(new_n17154_), .B1(new_n17146_), .B2(new_n17158_), .ZN(new_n17159_));
  NOR2_X1    g16967(.A1(new_n16597_), .A2(new_n16557_), .ZN(new_n17160_));
  OAI21_X1   g16968(.A1(\asqrt[6] ), .A2(new_n17160_), .B(new_n16604_), .ZN(new_n17161_));
  INV_X1     g16969(.I(new_n17161_), .ZN(new_n17162_));
  OAI21_X1   g16970(.A1(new_n17159_), .A2(new_n17126_), .B(new_n17162_), .ZN(new_n17163_));
  OAI21_X1   g16971(.A1(new_n17146_), .A2(\asqrt[62] ), .B(new_n17157_), .ZN(new_n17164_));
  NAND2_X1   g16972(.A1(new_n17146_), .A2(\asqrt[62] ), .ZN(new_n17165_));
  NAND3_X1   g16973(.A1(new_n17164_), .A2(new_n17165_), .A3(new_n17126_), .ZN(new_n17166_));
  NAND4_X1   g16974(.A1(new_n17163_), .A2(new_n193_), .A3(new_n17123_), .A4(new_n17166_), .ZN(\asqrt[5] ));
  AOI21_X1   g16975(.A1(new_n17101_), .A2(new_n17117_), .B(\asqrt[5] ), .ZN(new_n17168_));
  XOR2_X1    g16976(.A1(new_n17168_), .A2(new_n16614_), .Z(new_n17169_));
  AOI21_X1   g16977(.A1(new_n17098_), .A2(new_n17133_), .B(\asqrt[5] ), .ZN(new_n17170_));
  XOR2_X1    g16978(.A1(new_n17170_), .A2(new_n16617_), .Z(new_n17171_));
  NAND2_X1   g16979(.A1(new_n17111_), .A2(new_n531_), .ZN(new_n17172_));
  AOI21_X1   g16980(.A1(new_n17172_), .A2(new_n17097_), .B(\asqrt[5] ), .ZN(new_n17173_));
  XOR2_X1    g16981(.A1(new_n17173_), .A2(new_n16620_), .Z(new_n17174_));
  INV_X1     g16982(.I(new_n17174_), .ZN(new_n17175_));
  AOI21_X1   g16983(.A1(new_n17109_), .A2(new_n17094_), .B(\asqrt[5] ), .ZN(new_n17176_));
  XOR2_X1    g16984(.A1(new_n17176_), .A2(new_n16622_), .Z(new_n17177_));
  INV_X1     g16985(.I(new_n17177_), .ZN(new_n17178_));
  NAND2_X1   g16986(.A1(new_n17076_), .A2(new_n744_), .ZN(new_n17179_));
  AOI21_X1   g16987(.A1(new_n17179_), .A2(new_n17108_), .B(\asqrt[5] ), .ZN(new_n17180_));
  XOR2_X1    g16988(.A1(new_n17180_), .A2(new_n16625_), .Z(new_n17181_));
  AOI21_X1   g16989(.A1(new_n17074_), .A2(new_n17091_), .B(\asqrt[5] ), .ZN(new_n17182_));
  XOR2_X1    g16990(.A1(new_n17182_), .A2(new_n16629_), .Z(new_n17183_));
  NAND2_X1   g16991(.A1(new_n17087_), .A2(new_n1006_), .ZN(new_n17184_));
  AOI21_X1   g16992(.A1(new_n17184_), .A2(new_n17073_), .B(\asqrt[5] ), .ZN(new_n17185_));
  XOR2_X1    g16993(.A1(new_n17185_), .A2(new_n16632_), .Z(new_n17186_));
  INV_X1     g16994(.I(new_n17186_), .ZN(new_n17187_));
  AOI21_X1   g16995(.A1(new_n17085_), .A2(new_n17070_), .B(\asqrt[5] ), .ZN(new_n17188_));
  XOR2_X1    g16996(.A1(new_n17188_), .A2(new_n16634_), .Z(new_n17189_));
  INV_X1     g16997(.I(new_n17189_), .ZN(new_n17190_));
  NAND2_X1   g16998(.A1(new_n17052_), .A2(new_n1305_), .ZN(new_n17191_));
  AOI21_X1   g16999(.A1(new_n17191_), .A2(new_n17084_), .B(\asqrt[5] ), .ZN(new_n17192_));
  XOR2_X1    g17000(.A1(new_n17192_), .A2(new_n16637_), .Z(new_n17193_));
  AOI21_X1   g17001(.A1(new_n17050_), .A2(new_n17067_), .B(\asqrt[5] ), .ZN(new_n17194_));
  XOR2_X1    g17002(.A1(new_n17194_), .A2(new_n16641_), .Z(new_n17195_));
  NAND2_X1   g17003(.A1(new_n17063_), .A2(new_n1632_), .ZN(new_n17196_));
  AOI21_X1   g17004(.A1(new_n17196_), .A2(new_n17049_), .B(\asqrt[5] ), .ZN(new_n17197_));
  XOR2_X1    g17005(.A1(new_n17197_), .A2(new_n16644_), .Z(new_n17198_));
  INV_X1     g17006(.I(new_n17198_), .ZN(new_n17199_));
  AOI21_X1   g17007(.A1(new_n17061_), .A2(new_n17046_), .B(\asqrt[5] ), .ZN(new_n17200_));
  XOR2_X1    g17008(.A1(new_n17200_), .A2(new_n16646_), .Z(new_n17201_));
  INV_X1     g17009(.I(new_n17201_), .ZN(new_n17202_));
  NAND2_X1   g17010(.A1(new_n17028_), .A2(new_n1953_), .ZN(new_n17203_));
  AOI21_X1   g17011(.A1(new_n17203_), .A2(new_n17060_), .B(\asqrt[5] ), .ZN(new_n17204_));
  XOR2_X1    g17012(.A1(new_n17204_), .A2(new_n16649_), .Z(new_n17205_));
  AOI21_X1   g17013(.A1(new_n17026_), .A2(new_n17043_), .B(\asqrt[5] ), .ZN(new_n17206_));
  XOR2_X1    g17014(.A1(new_n17206_), .A2(new_n16653_), .Z(new_n17207_));
  NAND2_X1   g17015(.A1(new_n17039_), .A2(new_n2332_), .ZN(new_n17208_));
  AOI21_X1   g17016(.A1(new_n17208_), .A2(new_n17025_), .B(\asqrt[5] ), .ZN(new_n17209_));
  XOR2_X1    g17017(.A1(new_n17209_), .A2(new_n16656_), .Z(new_n17210_));
  INV_X1     g17018(.I(new_n17210_), .ZN(new_n17211_));
  AOI21_X1   g17019(.A1(new_n17037_), .A2(new_n17022_), .B(\asqrt[5] ), .ZN(new_n17212_));
  XOR2_X1    g17020(.A1(new_n17212_), .A2(new_n16658_), .Z(new_n17213_));
  INV_X1     g17021(.I(new_n17213_), .ZN(new_n17214_));
  NAND2_X1   g17022(.A1(new_n17004_), .A2(new_n2749_), .ZN(new_n17215_));
  AOI21_X1   g17023(.A1(new_n17215_), .A2(new_n17036_), .B(\asqrt[5] ), .ZN(new_n17216_));
  XOR2_X1    g17024(.A1(new_n17216_), .A2(new_n16661_), .Z(new_n17217_));
  AOI21_X1   g17025(.A1(new_n17002_), .A2(new_n17019_), .B(\asqrt[5] ), .ZN(new_n17218_));
  XOR2_X1    g17026(.A1(new_n17218_), .A2(new_n16665_), .Z(new_n17219_));
  NAND2_X1   g17027(.A1(new_n17015_), .A2(new_n3195_), .ZN(new_n17220_));
  AOI21_X1   g17028(.A1(new_n17220_), .A2(new_n17001_), .B(\asqrt[5] ), .ZN(new_n17221_));
  XOR2_X1    g17029(.A1(new_n17221_), .A2(new_n16668_), .Z(new_n17222_));
  INV_X1     g17030(.I(new_n17222_), .ZN(new_n17223_));
  AOI21_X1   g17031(.A1(new_n17013_), .A2(new_n16998_), .B(\asqrt[5] ), .ZN(new_n17224_));
  XOR2_X1    g17032(.A1(new_n17224_), .A2(new_n16670_), .Z(new_n17225_));
  INV_X1     g17033(.I(new_n17225_), .ZN(new_n17226_));
  NAND2_X1   g17034(.A1(new_n16980_), .A2(new_n3681_), .ZN(new_n17227_));
  AOI21_X1   g17035(.A1(new_n17227_), .A2(new_n17012_), .B(\asqrt[5] ), .ZN(new_n17228_));
  XOR2_X1    g17036(.A1(new_n17228_), .A2(new_n16673_), .Z(new_n17229_));
  AOI21_X1   g17037(.A1(new_n16978_), .A2(new_n16995_), .B(\asqrt[5] ), .ZN(new_n17230_));
  XOR2_X1    g17038(.A1(new_n17230_), .A2(new_n16677_), .Z(new_n17231_));
  NAND2_X1   g17039(.A1(new_n16991_), .A2(new_n4196_), .ZN(new_n17232_));
  AOI21_X1   g17040(.A1(new_n17232_), .A2(new_n16977_), .B(\asqrt[5] ), .ZN(new_n17233_));
  XOR2_X1    g17041(.A1(new_n17233_), .A2(new_n16680_), .Z(new_n17234_));
  INV_X1     g17042(.I(new_n17234_), .ZN(new_n17235_));
  AOI21_X1   g17043(.A1(new_n16989_), .A2(new_n16974_), .B(\asqrt[5] ), .ZN(new_n17236_));
  XOR2_X1    g17044(.A1(new_n17236_), .A2(new_n16682_), .Z(new_n17237_));
  INV_X1     g17045(.I(new_n17237_), .ZN(new_n17238_));
  NAND2_X1   g17046(.A1(new_n16956_), .A2(new_n4751_), .ZN(new_n17239_));
  AOI21_X1   g17047(.A1(new_n17239_), .A2(new_n16988_), .B(\asqrt[5] ), .ZN(new_n17240_));
  XOR2_X1    g17048(.A1(new_n17240_), .A2(new_n16685_), .Z(new_n17241_));
  AOI21_X1   g17049(.A1(new_n16954_), .A2(new_n16971_), .B(\asqrt[5] ), .ZN(new_n17242_));
  XOR2_X1    g17050(.A1(new_n17242_), .A2(new_n16689_), .Z(new_n17243_));
  NAND2_X1   g17051(.A1(new_n16967_), .A2(new_n5336_), .ZN(new_n17244_));
  AOI21_X1   g17052(.A1(new_n17244_), .A2(new_n16953_), .B(\asqrt[5] ), .ZN(new_n17245_));
  XOR2_X1    g17053(.A1(new_n17245_), .A2(new_n16692_), .Z(new_n17246_));
  INV_X1     g17054(.I(new_n17246_), .ZN(new_n17247_));
  AOI21_X1   g17055(.A1(new_n16965_), .A2(new_n16950_), .B(\asqrt[5] ), .ZN(new_n17248_));
  XOR2_X1    g17056(.A1(new_n17248_), .A2(new_n16694_), .Z(new_n17249_));
  INV_X1     g17057(.I(new_n17249_), .ZN(new_n17250_));
  NAND2_X1   g17058(.A1(new_n16932_), .A2(new_n5947_), .ZN(new_n17251_));
  AOI21_X1   g17059(.A1(new_n17251_), .A2(new_n16964_), .B(\asqrt[5] ), .ZN(new_n17252_));
  XOR2_X1    g17060(.A1(new_n17252_), .A2(new_n16697_), .Z(new_n17253_));
  AOI21_X1   g17061(.A1(new_n16930_), .A2(new_n16947_), .B(\asqrt[5] ), .ZN(new_n17254_));
  XOR2_X1    g17062(.A1(new_n17254_), .A2(new_n16701_), .Z(new_n17255_));
  NAND2_X1   g17063(.A1(new_n16943_), .A2(new_n6636_), .ZN(new_n17256_));
  AOI21_X1   g17064(.A1(new_n17256_), .A2(new_n16929_), .B(\asqrt[5] ), .ZN(new_n17257_));
  XOR2_X1    g17065(.A1(new_n17257_), .A2(new_n16704_), .Z(new_n17258_));
  INV_X1     g17066(.I(new_n17258_), .ZN(new_n17259_));
  AOI21_X1   g17067(.A1(new_n16941_), .A2(new_n16926_), .B(\asqrt[5] ), .ZN(new_n17260_));
  XOR2_X1    g17068(.A1(new_n17260_), .A2(new_n16706_), .Z(new_n17261_));
  INV_X1     g17069(.I(new_n17261_), .ZN(new_n17262_));
  NAND2_X1   g17070(.A1(new_n16908_), .A2(new_n7331_), .ZN(new_n17263_));
  AOI21_X1   g17071(.A1(new_n17263_), .A2(new_n16940_), .B(\asqrt[5] ), .ZN(new_n17264_));
  XOR2_X1    g17072(.A1(new_n17264_), .A2(new_n16709_), .Z(new_n17265_));
  AOI21_X1   g17073(.A1(new_n16906_), .A2(new_n16923_), .B(\asqrt[5] ), .ZN(new_n17266_));
  XOR2_X1    g17074(.A1(new_n17266_), .A2(new_n16713_), .Z(new_n17267_));
  NAND2_X1   g17075(.A1(new_n16919_), .A2(new_n8077_), .ZN(new_n17268_));
  AOI21_X1   g17076(.A1(new_n17268_), .A2(new_n16905_), .B(\asqrt[5] ), .ZN(new_n17269_));
  XOR2_X1    g17077(.A1(new_n17269_), .A2(new_n16716_), .Z(new_n17270_));
  INV_X1     g17078(.I(new_n17270_), .ZN(new_n17271_));
  AOI21_X1   g17079(.A1(new_n16917_), .A2(new_n16902_), .B(\asqrt[5] ), .ZN(new_n17272_));
  XOR2_X1    g17080(.A1(new_n17272_), .A2(new_n16718_), .Z(new_n17273_));
  INV_X1     g17081(.I(new_n17273_), .ZN(new_n17274_));
  NAND2_X1   g17082(.A1(new_n16884_), .A2(new_n8849_), .ZN(new_n17275_));
  AOI21_X1   g17083(.A1(new_n17275_), .A2(new_n16916_), .B(\asqrt[5] ), .ZN(new_n17276_));
  XOR2_X1    g17084(.A1(new_n17276_), .A2(new_n16721_), .Z(new_n17277_));
  AOI21_X1   g17085(.A1(new_n16882_), .A2(new_n16899_), .B(\asqrt[5] ), .ZN(new_n17278_));
  XOR2_X1    g17086(.A1(new_n17278_), .A2(new_n16725_), .Z(new_n17279_));
  NAND2_X1   g17087(.A1(new_n16895_), .A2(new_n9656_), .ZN(new_n17280_));
  AOI21_X1   g17088(.A1(new_n17280_), .A2(new_n16881_), .B(\asqrt[5] ), .ZN(new_n17281_));
  XOR2_X1    g17089(.A1(new_n17281_), .A2(new_n16728_), .Z(new_n17282_));
  INV_X1     g17090(.I(new_n17282_), .ZN(new_n17283_));
  AOI21_X1   g17091(.A1(new_n16893_), .A2(new_n16878_), .B(\asqrt[5] ), .ZN(new_n17284_));
  XOR2_X1    g17092(.A1(new_n17284_), .A2(new_n16730_), .Z(new_n17285_));
  INV_X1     g17093(.I(new_n17285_), .ZN(new_n17286_));
  NAND2_X1   g17094(.A1(new_n16860_), .A2(new_n10497_), .ZN(new_n17287_));
  AOI21_X1   g17095(.A1(new_n17287_), .A2(new_n16892_), .B(\asqrt[5] ), .ZN(new_n17288_));
  XOR2_X1    g17096(.A1(new_n17288_), .A2(new_n16733_), .Z(new_n17289_));
  AOI21_X1   g17097(.A1(new_n16858_), .A2(new_n16875_), .B(\asqrt[5] ), .ZN(new_n17290_));
  XOR2_X1    g17098(.A1(new_n17290_), .A2(new_n16737_), .Z(new_n17291_));
  NAND2_X1   g17099(.A1(new_n16871_), .A2(new_n11373_), .ZN(new_n17292_));
  AOI21_X1   g17100(.A1(new_n17292_), .A2(new_n16857_), .B(\asqrt[5] ), .ZN(new_n17293_));
  XOR2_X1    g17101(.A1(new_n17293_), .A2(new_n16740_), .Z(new_n17294_));
  INV_X1     g17102(.I(new_n17294_), .ZN(new_n17295_));
  AOI21_X1   g17103(.A1(new_n16869_), .A2(new_n16854_), .B(\asqrt[5] ), .ZN(new_n17296_));
  XOR2_X1    g17104(.A1(new_n17296_), .A2(new_n16742_), .Z(new_n17297_));
  INV_X1     g17105(.I(new_n17297_), .ZN(new_n17298_));
  NAND2_X1   g17106(.A1(new_n16836_), .A2(new_n12283_), .ZN(new_n17299_));
  AOI21_X1   g17107(.A1(new_n17299_), .A2(new_n16868_), .B(\asqrt[5] ), .ZN(new_n17300_));
  XOR2_X1    g17108(.A1(new_n17300_), .A2(new_n16745_), .Z(new_n17301_));
  AOI21_X1   g17109(.A1(new_n16834_), .A2(new_n16851_), .B(\asqrt[5] ), .ZN(new_n17302_));
  XOR2_X1    g17110(.A1(new_n17302_), .A2(new_n16749_), .Z(new_n17303_));
  NAND2_X1   g17111(.A1(new_n16847_), .A2(new_n13228_), .ZN(new_n17304_));
  AOI21_X1   g17112(.A1(new_n17304_), .A2(new_n16833_), .B(\asqrt[5] ), .ZN(new_n17305_));
  XOR2_X1    g17113(.A1(new_n17305_), .A2(new_n16752_), .Z(new_n17306_));
  INV_X1     g17114(.I(new_n17306_), .ZN(new_n17307_));
  AOI21_X1   g17115(.A1(new_n16845_), .A2(new_n16830_), .B(\asqrt[5] ), .ZN(new_n17308_));
  XOR2_X1    g17116(.A1(new_n17308_), .A2(new_n16754_), .Z(new_n17309_));
  INV_X1     g17117(.I(new_n17309_), .ZN(new_n17310_));
  NAND2_X1   g17118(.A1(new_n16807_), .A2(new_n14207_), .ZN(new_n17311_));
  AOI21_X1   g17119(.A1(new_n17311_), .A2(new_n16844_), .B(\asqrt[5] ), .ZN(new_n17312_));
  XOR2_X1    g17120(.A1(new_n17312_), .A2(new_n16757_), .Z(new_n17313_));
  AOI21_X1   g17121(.A1(new_n16805_), .A2(new_n16827_), .B(\asqrt[5] ), .ZN(new_n17314_));
  XOR2_X1    g17122(.A1(new_n17314_), .A2(new_n16760_), .Z(new_n17315_));
  NAND2_X1   g17123(.A1(new_n16823_), .A2(new_n15221_), .ZN(new_n17316_));
  AOI21_X1   g17124(.A1(new_n17316_), .A2(new_n16804_), .B(\asqrt[5] ), .ZN(new_n17317_));
  XOR2_X1    g17125(.A1(new_n17317_), .A2(new_n16767_), .Z(new_n17318_));
  INV_X1     g17126(.I(new_n17318_), .ZN(new_n17319_));
  AOI21_X1   g17127(.A1(new_n16821_), .A2(new_n16801_), .B(\asqrt[5] ), .ZN(new_n17320_));
  XOR2_X1    g17128(.A1(new_n17320_), .A2(new_n16812_), .Z(new_n17321_));
  INV_X1     g17129(.I(new_n17321_), .ZN(new_n17322_));
  NAND2_X1   g17130(.A1(\asqrt[6] ), .A2(new_n16788_), .ZN(new_n17323_));
  NOR2_X1    g17131(.A1(new_n16796_), .A2(\a[12] ), .ZN(new_n17324_));
  AOI22_X1   g17132(.A1(new_n17323_), .A2(new_n16796_), .B1(\asqrt[6] ), .B2(new_n17324_), .ZN(new_n17325_));
  OAI21_X1   g17133(.A1(new_n16779_), .A2(new_n16788_), .B(new_n16816_), .ZN(new_n17326_));
  AOI21_X1   g17134(.A1(new_n16815_), .A2(new_n17326_), .B(\asqrt[5] ), .ZN(new_n17327_));
  XOR2_X1    g17135(.A1(new_n17327_), .A2(new_n17325_), .Z(new_n17328_));
  NOR2_X1    g17136(.A1(new_n17122_), .A2(new_n16779_), .ZN(new_n17329_));
  NAND4_X1   g17137(.A1(new_n17163_), .A2(new_n193_), .A3(new_n17166_), .A4(new_n17329_), .ZN(new_n17330_));
  NAND2_X1   g17138(.A1(\asqrt[5] ), .A2(new_n16785_), .ZN(new_n17331_));
  AOI21_X1   g17139(.A1(new_n17331_), .A2(new_n17330_), .B(\a[12] ), .ZN(new_n17332_));
  NAND3_X1   g17140(.A1(new_n17148_), .A2(new_n239_), .A3(new_n17141_), .ZN(new_n17333_));
  AOI21_X1   g17141(.A1(new_n17144_), .A2(new_n17333_), .B(new_n17149_), .ZN(new_n17334_));
  AOI21_X1   g17142(.A1(new_n17145_), .A2(new_n17140_), .B(\asqrt[62] ), .ZN(new_n17335_));
  NOR3_X1    g17143(.A1(new_n17152_), .A2(new_n201_), .A3(new_n17149_), .ZN(new_n17336_));
  OAI22_X1   g17144(.A1(new_n17336_), .A2(new_n17335_), .B1(new_n17334_), .B2(new_n17157_), .ZN(new_n17337_));
  AOI21_X1   g17145(.A1(new_n17337_), .A2(new_n17125_), .B(new_n17161_), .ZN(new_n17338_));
  AOI21_X1   g17146(.A1(new_n17334_), .A2(new_n201_), .B(new_n17158_), .ZN(new_n17339_));
  OAI21_X1   g17147(.A1(new_n17334_), .A2(new_n201_), .B(new_n17126_), .ZN(new_n17340_));
  NOR2_X1    g17148(.A1(new_n17339_), .A2(new_n17340_), .ZN(new_n17341_));
  NOR4_X1    g17149(.A1(new_n17338_), .A2(\asqrt[63] ), .A3(new_n17122_), .A4(new_n17341_), .ZN(new_n17342_));
  OAI21_X1   g17150(.A1(new_n16786_), .A2(new_n17342_), .B(new_n17330_), .ZN(new_n17343_));
  NOR2_X1    g17151(.A1(new_n17343_), .A2(new_n16788_), .ZN(new_n17344_));
  NOR2_X1    g17152(.A1(new_n17344_), .A2(new_n17332_), .ZN(new_n17345_));
  INV_X1     g17153(.I(\a[10] ), .ZN(new_n17346_));
  NOR2_X1    g17154(.A1(\a[8] ), .A2(\a[9] ), .ZN(new_n17347_));
  NOR3_X1    g17155(.A1(new_n17342_), .A2(new_n17346_), .A3(new_n17347_), .ZN(new_n17348_));
  INV_X1     g17156(.I(new_n17347_), .ZN(new_n17349_));
  AOI21_X1   g17157(.A1(new_n17342_), .A2(\a[10] ), .B(new_n17349_), .ZN(new_n17350_));
  OAI21_X1   g17158(.A1(new_n17348_), .A2(new_n17350_), .B(\asqrt[6] ), .ZN(new_n17351_));
  INV_X1     g17159(.I(\a[11] ), .ZN(new_n17352_));
  AOI21_X1   g17160(.A1(\asqrt[5] ), .A2(new_n17346_), .B(new_n17352_), .ZN(new_n17353_));
  NOR3_X1    g17161(.A1(new_n17342_), .A2(\a[10] ), .A3(\a[11] ), .ZN(new_n17354_));
  INV_X1     g17162(.I(new_n16768_), .ZN(new_n17355_));
  NAND2_X1   g17163(.A1(new_n17347_), .A2(new_n17346_), .ZN(new_n17356_));
  NAND3_X1   g17164(.A1(new_n16607_), .A2(new_n16609_), .A3(new_n17356_), .ZN(new_n17357_));
  NOR2_X1    g17165(.A1(new_n16772_), .A2(new_n17357_), .ZN(new_n17358_));
  AOI21_X1   g17166(.A1(new_n17355_), .A2(new_n17358_), .B(new_n17346_), .ZN(new_n17359_));
  INV_X1     g17167(.I(new_n17359_), .ZN(new_n17360_));
  NOR2_X1    g17168(.A1(new_n17342_), .A2(new_n17360_), .ZN(new_n17361_));
  NOR3_X1    g17169(.A1(new_n17354_), .A2(new_n17353_), .A3(new_n17361_), .ZN(new_n17362_));
  NAND3_X1   g17170(.A1(new_n17351_), .A2(new_n17362_), .A3(new_n16269_), .ZN(new_n17363_));
  NAND2_X1   g17171(.A1(new_n17363_), .A2(new_n17345_), .ZN(new_n17364_));
  NAND3_X1   g17172(.A1(\asqrt[5] ), .A2(\a[10] ), .A3(new_n17349_), .ZN(new_n17365_));
  OAI21_X1   g17173(.A1(\asqrt[5] ), .A2(new_n17346_), .B(new_n17347_), .ZN(new_n17366_));
  AOI21_X1   g17174(.A1(new_n17366_), .A2(new_n17365_), .B(new_n16779_), .ZN(new_n17367_));
  OAI21_X1   g17175(.A1(new_n17342_), .A2(\a[10] ), .B(\a[11] ), .ZN(new_n17368_));
  NAND3_X1   g17176(.A1(\asqrt[5] ), .A2(new_n17346_), .A3(new_n17352_), .ZN(new_n17369_));
  NAND2_X1   g17177(.A1(\asqrt[5] ), .A2(new_n17359_), .ZN(new_n17370_));
  NAND3_X1   g17178(.A1(new_n17368_), .A2(new_n17369_), .A3(new_n17370_), .ZN(new_n17371_));
  OAI21_X1   g17179(.A1(new_n17367_), .A2(new_n17371_), .B(\asqrt[7] ), .ZN(new_n17372_));
  NAND3_X1   g17180(.A1(new_n17364_), .A2(new_n15717_), .A3(new_n17372_), .ZN(new_n17373_));
  AOI21_X1   g17181(.A1(new_n17364_), .A2(new_n17372_), .B(new_n15717_), .ZN(new_n17374_));
  AOI21_X1   g17182(.A1(new_n17328_), .A2(new_n17373_), .B(new_n17374_), .ZN(new_n17375_));
  AOI21_X1   g17183(.A1(new_n17375_), .A2(new_n15221_), .B(new_n17322_), .ZN(new_n17376_));
  XOR2_X1    g17184(.A1(new_n17343_), .A2(\a[12] ), .Z(new_n17377_));
  NOR3_X1    g17185(.A1(new_n17367_), .A2(new_n17371_), .A3(\asqrt[7] ), .ZN(new_n17378_));
  OAI21_X1   g17186(.A1(new_n17377_), .A2(new_n17378_), .B(new_n17372_), .ZN(new_n17379_));
  OAI21_X1   g17187(.A1(new_n17379_), .A2(\asqrt[8] ), .B(new_n17328_), .ZN(new_n17380_));
  NAND2_X1   g17188(.A1(new_n17379_), .A2(\asqrt[8] ), .ZN(new_n17381_));
  AOI21_X1   g17189(.A1(new_n17380_), .A2(new_n17381_), .B(new_n15221_), .ZN(new_n17382_));
  NOR3_X1    g17190(.A1(new_n17376_), .A2(\asqrt[10] ), .A3(new_n17382_), .ZN(new_n17383_));
  OAI21_X1   g17191(.A1(new_n17376_), .A2(new_n17382_), .B(\asqrt[10] ), .ZN(new_n17384_));
  OAI21_X1   g17192(.A1(new_n17319_), .A2(new_n17383_), .B(new_n17384_), .ZN(new_n17385_));
  OAI21_X1   g17193(.A1(new_n17385_), .A2(\asqrt[11] ), .B(new_n17315_), .ZN(new_n17386_));
  NAND3_X1   g17194(.A1(new_n17380_), .A2(new_n17381_), .A3(new_n15221_), .ZN(new_n17387_));
  AOI21_X1   g17195(.A1(new_n17321_), .A2(new_n17387_), .B(new_n17382_), .ZN(new_n17388_));
  AOI21_X1   g17196(.A1(new_n17388_), .A2(new_n14690_), .B(new_n17319_), .ZN(new_n17389_));
  NAND2_X1   g17197(.A1(new_n17387_), .A2(new_n17321_), .ZN(new_n17390_));
  INV_X1     g17198(.I(new_n17382_), .ZN(new_n17391_));
  AOI21_X1   g17199(.A1(new_n17390_), .A2(new_n17391_), .B(new_n14690_), .ZN(new_n17392_));
  OAI21_X1   g17200(.A1(new_n17389_), .A2(new_n17392_), .B(\asqrt[11] ), .ZN(new_n17393_));
  NAND3_X1   g17201(.A1(new_n17386_), .A2(new_n13690_), .A3(new_n17393_), .ZN(new_n17394_));
  AOI21_X1   g17202(.A1(new_n17386_), .A2(new_n17393_), .B(new_n13690_), .ZN(new_n17395_));
  AOI21_X1   g17203(.A1(new_n17313_), .A2(new_n17394_), .B(new_n17395_), .ZN(new_n17396_));
  AOI21_X1   g17204(.A1(new_n17396_), .A2(new_n13228_), .B(new_n17310_), .ZN(new_n17397_));
  INV_X1     g17205(.I(new_n17315_), .ZN(new_n17398_));
  NOR3_X1    g17206(.A1(new_n17389_), .A2(\asqrt[11] ), .A3(new_n17392_), .ZN(new_n17399_));
  OAI21_X1   g17207(.A1(new_n17398_), .A2(new_n17399_), .B(new_n17393_), .ZN(new_n17400_));
  OAI21_X1   g17208(.A1(new_n17400_), .A2(\asqrt[12] ), .B(new_n17313_), .ZN(new_n17401_));
  NAND2_X1   g17209(.A1(new_n17400_), .A2(\asqrt[12] ), .ZN(new_n17402_));
  AOI21_X1   g17210(.A1(new_n17401_), .A2(new_n17402_), .B(new_n13228_), .ZN(new_n17403_));
  NOR3_X1    g17211(.A1(new_n17397_), .A2(\asqrt[14] ), .A3(new_n17403_), .ZN(new_n17404_));
  OAI21_X1   g17212(.A1(new_n17397_), .A2(new_n17403_), .B(\asqrt[14] ), .ZN(new_n17405_));
  OAI21_X1   g17213(.A1(new_n17307_), .A2(new_n17404_), .B(new_n17405_), .ZN(new_n17406_));
  OAI21_X1   g17214(.A1(new_n17406_), .A2(\asqrt[15] ), .B(new_n17303_), .ZN(new_n17407_));
  NAND3_X1   g17215(.A1(new_n17401_), .A2(new_n17402_), .A3(new_n13228_), .ZN(new_n17408_));
  AOI21_X1   g17216(.A1(new_n17309_), .A2(new_n17408_), .B(new_n17403_), .ZN(new_n17409_));
  AOI21_X1   g17217(.A1(new_n17409_), .A2(new_n12733_), .B(new_n17307_), .ZN(new_n17410_));
  NAND2_X1   g17218(.A1(new_n17408_), .A2(new_n17309_), .ZN(new_n17411_));
  INV_X1     g17219(.I(new_n17403_), .ZN(new_n17412_));
  AOI21_X1   g17220(.A1(new_n17411_), .A2(new_n17412_), .B(new_n12733_), .ZN(new_n17413_));
  OAI21_X1   g17221(.A1(new_n17410_), .A2(new_n17413_), .B(\asqrt[15] ), .ZN(new_n17414_));
  NAND3_X1   g17222(.A1(new_n17407_), .A2(new_n11802_), .A3(new_n17414_), .ZN(new_n17415_));
  AOI21_X1   g17223(.A1(new_n17407_), .A2(new_n17414_), .B(new_n11802_), .ZN(new_n17416_));
  AOI21_X1   g17224(.A1(new_n17301_), .A2(new_n17415_), .B(new_n17416_), .ZN(new_n17417_));
  AOI21_X1   g17225(.A1(new_n17417_), .A2(new_n11373_), .B(new_n17298_), .ZN(new_n17418_));
  INV_X1     g17226(.I(new_n17303_), .ZN(new_n17419_));
  NOR3_X1    g17227(.A1(new_n17410_), .A2(\asqrt[15] ), .A3(new_n17413_), .ZN(new_n17420_));
  OAI21_X1   g17228(.A1(new_n17419_), .A2(new_n17420_), .B(new_n17414_), .ZN(new_n17421_));
  OAI21_X1   g17229(.A1(new_n17421_), .A2(\asqrt[16] ), .B(new_n17301_), .ZN(new_n17422_));
  NAND2_X1   g17230(.A1(new_n17421_), .A2(\asqrt[16] ), .ZN(new_n17423_));
  AOI21_X1   g17231(.A1(new_n17422_), .A2(new_n17423_), .B(new_n11373_), .ZN(new_n17424_));
  NOR3_X1    g17232(.A1(new_n17418_), .A2(\asqrt[18] ), .A3(new_n17424_), .ZN(new_n17425_));
  OAI21_X1   g17233(.A1(new_n17418_), .A2(new_n17424_), .B(\asqrt[18] ), .ZN(new_n17426_));
  OAI21_X1   g17234(.A1(new_n17295_), .A2(new_n17425_), .B(new_n17426_), .ZN(new_n17427_));
  OAI21_X1   g17235(.A1(new_n17427_), .A2(\asqrt[19] ), .B(new_n17291_), .ZN(new_n17428_));
  NAND3_X1   g17236(.A1(new_n17422_), .A2(new_n17423_), .A3(new_n11373_), .ZN(new_n17429_));
  AOI21_X1   g17237(.A1(new_n17297_), .A2(new_n17429_), .B(new_n17424_), .ZN(new_n17430_));
  AOI21_X1   g17238(.A1(new_n17430_), .A2(new_n10914_), .B(new_n17295_), .ZN(new_n17431_));
  NAND2_X1   g17239(.A1(new_n17429_), .A2(new_n17297_), .ZN(new_n17432_));
  INV_X1     g17240(.I(new_n17424_), .ZN(new_n17433_));
  AOI21_X1   g17241(.A1(new_n17432_), .A2(new_n17433_), .B(new_n10914_), .ZN(new_n17434_));
  OAI21_X1   g17242(.A1(new_n17431_), .A2(new_n17434_), .B(\asqrt[19] ), .ZN(new_n17435_));
  NAND3_X1   g17243(.A1(new_n17428_), .A2(new_n10052_), .A3(new_n17435_), .ZN(new_n17436_));
  AOI21_X1   g17244(.A1(new_n17428_), .A2(new_n17435_), .B(new_n10052_), .ZN(new_n17437_));
  AOI21_X1   g17245(.A1(new_n17289_), .A2(new_n17436_), .B(new_n17437_), .ZN(new_n17438_));
  AOI21_X1   g17246(.A1(new_n17438_), .A2(new_n9656_), .B(new_n17286_), .ZN(new_n17439_));
  INV_X1     g17247(.I(new_n17291_), .ZN(new_n17440_));
  NOR3_X1    g17248(.A1(new_n17431_), .A2(\asqrt[19] ), .A3(new_n17434_), .ZN(new_n17441_));
  OAI21_X1   g17249(.A1(new_n17440_), .A2(new_n17441_), .B(new_n17435_), .ZN(new_n17442_));
  OAI21_X1   g17250(.A1(new_n17442_), .A2(\asqrt[20] ), .B(new_n17289_), .ZN(new_n17443_));
  NAND2_X1   g17251(.A1(new_n17442_), .A2(\asqrt[20] ), .ZN(new_n17444_));
  AOI21_X1   g17252(.A1(new_n17443_), .A2(new_n17444_), .B(new_n9656_), .ZN(new_n17445_));
  NOR3_X1    g17253(.A1(new_n17439_), .A2(\asqrt[22] ), .A3(new_n17445_), .ZN(new_n17446_));
  OAI21_X1   g17254(.A1(new_n17439_), .A2(new_n17445_), .B(\asqrt[22] ), .ZN(new_n17447_));
  OAI21_X1   g17255(.A1(new_n17283_), .A2(new_n17446_), .B(new_n17447_), .ZN(new_n17448_));
  OAI21_X1   g17256(.A1(new_n17448_), .A2(\asqrt[23] ), .B(new_n17279_), .ZN(new_n17449_));
  NAND3_X1   g17257(.A1(new_n17443_), .A2(new_n17444_), .A3(new_n9656_), .ZN(new_n17450_));
  AOI21_X1   g17258(.A1(new_n17285_), .A2(new_n17450_), .B(new_n17445_), .ZN(new_n17451_));
  AOI21_X1   g17259(.A1(new_n17451_), .A2(new_n9233_), .B(new_n17283_), .ZN(new_n17452_));
  NAND2_X1   g17260(.A1(new_n17450_), .A2(new_n17285_), .ZN(new_n17453_));
  INV_X1     g17261(.I(new_n17445_), .ZN(new_n17454_));
  AOI21_X1   g17262(.A1(new_n17453_), .A2(new_n17454_), .B(new_n9233_), .ZN(new_n17455_));
  OAI21_X1   g17263(.A1(new_n17452_), .A2(new_n17455_), .B(\asqrt[23] ), .ZN(new_n17456_));
  NAND3_X1   g17264(.A1(new_n17449_), .A2(new_n8440_), .A3(new_n17456_), .ZN(new_n17457_));
  AOI21_X1   g17265(.A1(new_n17449_), .A2(new_n17456_), .B(new_n8440_), .ZN(new_n17458_));
  AOI21_X1   g17266(.A1(new_n17277_), .A2(new_n17457_), .B(new_n17458_), .ZN(new_n17459_));
  AOI21_X1   g17267(.A1(new_n17459_), .A2(new_n8077_), .B(new_n17274_), .ZN(new_n17460_));
  INV_X1     g17268(.I(new_n17279_), .ZN(new_n17461_));
  NOR3_X1    g17269(.A1(new_n17452_), .A2(\asqrt[23] ), .A3(new_n17455_), .ZN(new_n17462_));
  OAI21_X1   g17270(.A1(new_n17461_), .A2(new_n17462_), .B(new_n17456_), .ZN(new_n17463_));
  OAI21_X1   g17271(.A1(new_n17463_), .A2(\asqrt[24] ), .B(new_n17277_), .ZN(new_n17464_));
  NAND2_X1   g17272(.A1(new_n17463_), .A2(\asqrt[24] ), .ZN(new_n17465_));
  AOI21_X1   g17273(.A1(new_n17464_), .A2(new_n17465_), .B(new_n8077_), .ZN(new_n17466_));
  NOR3_X1    g17274(.A1(new_n17460_), .A2(\asqrt[26] ), .A3(new_n17466_), .ZN(new_n17467_));
  OAI21_X1   g17275(.A1(new_n17460_), .A2(new_n17466_), .B(\asqrt[26] ), .ZN(new_n17468_));
  OAI21_X1   g17276(.A1(new_n17271_), .A2(new_n17467_), .B(new_n17468_), .ZN(new_n17469_));
  OAI21_X1   g17277(.A1(new_n17469_), .A2(\asqrt[27] ), .B(new_n17267_), .ZN(new_n17470_));
  NAND3_X1   g17278(.A1(new_n17464_), .A2(new_n17465_), .A3(new_n8077_), .ZN(new_n17471_));
  AOI21_X1   g17279(.A1(new_n17273_), .A2(new_n17471_), .B(new_n17466_), .ZN(new_n17472_));
  AOI21_X1   g17280(.A1(new_n17472_), .A2(new_n7690_), .B(new_n17271_), .ZN(new_n17473_));
  NAND2_X1   g17281(.A1(new_n17471_), .A2(new_n17273_), .ZN(new_n17474_));
  INV_X1     g17282(.I(new_n17466_), .ZN(new_n17475_));
  AOI21_X1   g17283(.A1(new_n17474_), .A2(new_n17475_), .B(new_n7690_), .ZN(new_n17476_));
  OAI21_X1   g17284(.A1(new_n17473_), .A2(new_n17476_), .B(\asqrt[27] ), .ZN(new_n17477_));
  NAND3_X1   g17285(.A1(new_n17470_), .A2(new_n6966_), .A3(new_n17477_), .ZN(new_n17478_));
  AOI21_X1   g17286(.A1(new_n17470_), .A2(new_n17477_), .B(new_n6966_), .ZN(new_n17479_));
  AOI21_X1   g17287(.A1(new_n17265_), .A2(new_n17478_), .B(new_n17479_), .ZN(new_n17480_));
  AOI21_X1   g17288(.A1(new_n17480_), .A2(new_n6636_), .B(new_n17262_), .ZN(new_n17481_));
  INV_X1     g17289(.I(new_n17267_), .ZN(new_n17482_));
  NOR3_X1    g17290(.A1(new_n17473_), .A2(\asqrt[27] ), .A3(new_n17476_), .ZN(new_n17483_));
  OAI21_X1   g17291(.A1(new_n17482_), .A2(new_n17483_), .B(new_n17477_), .ZN(new_n17484_));
  OAI21_X1   g17292(.A1(new_n17484_), .A2(\asqrt[28] ), .B(new_n17265_), .ZN(new_n17485_));
  NAND2_X1   g17293(.A1(new_n17484_), .A2(\asqrt[28] ), .ZN(new_n17486_));
  AOI21_X1   g17294(.A1(new_n17485_), .A2(new_n17486_), .B(new_n6636_), .ZN(new_n17487_));
  NOR3_X1    g17295(.A1(new_n17481_), .A2(\asqrt[30] ), .A3(new_n17487_), .ZN(new_n17488_));
  OAI21_X1   g17296(.A1(new_n17481_), .A2(new_n17487_), .B(\asqrt[30] ), .ZN(new_n17489_));
  OAI21_X1   g17297(.A1(new_n17259_), .A2(new_n17488_), .B(new_n17489_), .ZN(new_n17490_));
  OAI21_X1   g17298(.A1(new_n17490_), .A2(\asqrt[31] ), .B(new_n17255_), .ZN(new_n17491_));
  NAND3_X1   g17299(.A1(new_n17485_), .A2(new_n17486_), .A3(new_n6636_), .ZN(new_n17492_));
  AOI21_X1   g17300(.A1(new_n17261_), .A2(new_n17492_), .B(new_n17487_), .ZN(new_n17493_));
  AOI21_X1   g17301(.A1(new_n17493_), .A2(new_n6275_), .B(new_n17259_), .ZN(new_n17494_));
  NAND2_X1   g17302(.A1(new_n17492_), .A2(new_n17261_), .ZN(new_n17495_));
  INV_X1     g17303(.I(new_n17487_), .ZN(new_n17496_));
  AOI21_X1   g17304(.A1(new_n17495_), .A2(new_n17496_), .B(new_n6275_), .ZN(new_n17497_));
  OAI21_X1   g17305(.A1(new_n17494_), .A2(new_n17497_), .B(\asqrt[31] ), .ZN(new_n17498_));
  NAND3_X1   g17306(.A1(new_n17491_), .A2(new_n5643_), .A3(new_n17498_), .ZN(new_n17499_));
  AOI21_X1   g17307(.A1(new_n17491_), .A2(new_n17498_), .B(new_n5643_), .ZN(new_n17500_));
  AOI21_X1   g17308(.A1(new_n17253_), .A2(new_n17499_), .B(new_n17500_), .ZN(new_n17501_));
  AOI21_X1   g17309(.A1(new_n17501_), .A2(new_n5336_), .B(new_n17250_), .ZN(new_n17502_));
  INV_X1     g17310(.I(new_n17255_), .ZN(new_n17503_));
  NOR3_X1    g17311(.A1(new_n17494_), .A2(\asqrt[31] ), .A3(new_n17497_), .ZN(new_n17504_));
  OAI21_X1   g17312(.A1(new_n17503_), .A2(new_n17504_), .B(new_n17498_), .ZN(new_n17505_));
  OAI21_X1   g17313(.A1(new_n17505_), .A2(\asqrt[32] ), .B(new_n17253_), .ZN(new_n17506_));
  NAND2_X1   g17314(.A1(new_n17505_), .A2(\asqrt[32] ), .ZN(new_n17507_));
  AOI21_X1   g17315(.A1(new_n17506_), .A2(new_n17507_), .B(new_n5336_), .ZN(new_n17508_));
  NOR3_X1    g17316(.A1(new_n17502_), .A2(\asqrt[34] ), .A3(new_n17508_), .ZN(new_n17509_));
  OAI21_X1   g17317(.A1(new_n17502_), .A2(new_n17508_), .B(\asqrt[34] ), .ZN(new_n17510_));
  OAI21_X1   g17318(.A1(new_n17247_), .A2(new_n17509_), .B(new_n17510_), .ZN(new_n17511_));
  OAI21_X1   g17319(.A1(new_n17511_), .A2(\asqrt[35] ), .B(new_n17243_), .ZN(new_n17512_));
  NAND3_X1   g17320(.A1(new_n17506_), .A2(new_n17507_), .A3(new_n5336_), .ZN(new_n17513_));
  AOI21_X1   g17321(.A1(new_n17249_), .A2(new_n17513_), .B(new_n17508_), .ZN(new_n17514_));
  AOI21_X1   g17322(.A1(new_n17514_), .A2(new_n5029_), .B(new_n17247_), .ZN(new_n17515_));
  NAND2_X1   g17323(.A1(new_n17513_), .A2(new_n17249_), .ZN(new_n17516_));
  INV_X1     g17324(.I(new_n17508_), .ZN(new_n17517_));
  AOI21_X1   g17325(.A1(new_n17516_), .A2(new_n17517_), .B(new_n5029_), .ZN(new_n17518_));
  OAI21_X1   g17326(.A1(new_n17515_), .A2(new_n17518_), .B(\asqrt[35] ), .ZN(new_n17519_));
  NAND3_X1   g17327(.A1(new_n17512_), .A2(new_n4461_), .A3(new_n17519_), .ZN(new_n17520_));
  AOI21_X1   g17328(.A1(new_n17512_), .A2(new_n17519_), .B(new_n4461_), .ZN(new_n17521_));
  AOI21_X1   g17329(.A1(new_n17241_), .A2(new_n17520_), .B(new_n17521_), .ZN(new_n17522_));
  AOI21_X1   g17330(.A1(new_n17522_), .A2(new_n4196_), .B(new_n17238_), .ZN(new_n17523_));
  INV_X1     g17331(.I(new_n17243_), .ZN(new_n17524_));
  NOR3_X1    g17332(.A1(new_n17515_), .A2(\asqrt[35] ), .A3(new_n17518_), .ZN(new_n17525_));
  OAI21_X1   g17333(.A1(new_n17524_), .A2(new_n17525_), .B(new_n17519_), .ZN(new_n17526_));
  OAI21_X1   g17334(.A1(new_n17526_), .A2(\asqrt[36] ), .B(new_n17241_), .ZN(new_n17527_));
  NAND2_X1   g17335(.A1(new_n17526_), .A2(\asqrt[36] ), .ZN(new_n17528_));
  AOI21_X1   g17336(.A1(new_n17527_), .A2(new_n17528_), .B(new_n4196_), .ZN(new_n17529_));
  NOR3_X1    g17337(.A1(new_n17523_), .A2(\asqrt[38] ), .A3(new_n17529_), .ZN(new_n17530_));
  OAI21_X1   g17338(.A1(new_n17523_), .A2(new_n17529_), .B(\asqrt[38] ), .ZN(new_n17531_));
  OAI21_X1   g17339(.A1(new_n17235_), .A2(new_n17530_), .B(new_n17531_), .ZN(new_n17532_));
  OAI21_X1   g17340(.A1(new_n17532_), .A2(\asqrt[39] ), .B(new_n17231_), .ZN(new_n17533_));
  NAND3_X1   g17341(.A1(new_n17527_), .A2(new_n17528_), .A3(new_n4196_), .ZN(new_n17534_));
  AOI21_X1   g17342(.A1(new_n17237_), .A2(new_n17534_), .B(new_n17529_), .ZN(new_n17535_));
  AOI21_X1   g17343(.A1(new_n17535_), .A2(new_n3925_), .B(new_n17235_), .ZN(new_n17536_));
  NAND2_X1   g17344(.A1(new_n17534_), .A2(new_n17237_), .ZN(new_n17537_));
  INV_X1     g17345(.I(new_n17529_), .ZN(new_n17538_));
  AOI21_X1   g17346(.A1(new_n17537_), .A2(new_n17538_), .B(new_n3925_), .ZN(new_n17539_));
  OAI21_X1   g17347(.A1(new_n17536_), .A2(new_n17539_), .B(\asqrt[39] ), .ZN(new_n17540_));
  NAND3_X1   g17348(.A1(new_n17533_), .A2(new_n3427_), .A3(new_n17540_), .ZN(new_n17541_));
  AOI21_X1   g17349(.A1(new_n17533_), .A2(new_n17540_), .B(new_n3427_), .ZN(new_n17542_));
  AOI21_X1   g17350(.A1(new_n17229_), .A2(new_n17541_), .B(new_n17542_), .ZN(new_n17543_));
  AOI21_X1   g17351(.A1(new_n17543_), .A2(new_n3195_), .B(new_n17226_), .ZN(new_n17544_));
  INV_X1     g17352(.I(new_n17231_), .ZN(new_n17545_));
  NOR3_X1    g17353(.A1(new_n17536_), .A2(\asqrt[39] ), .A3(new_n17539_), .ZN(new_n17546_));
  OAI21_X1   g17354(.A1(new_n17545_), .A2(new_n17546_), .B(new_n17540_), .ZN(new_n17547_));
  OAI21_X1   g17355(.A1(new_n17547_), .A2(\asqrt[40] ), .B(new_n17229_), .ZN(new_n17548_));
  NAND2_X1   g17356(.A1(new_n17547_), .A2(\asqrt[40] ), .ZN(new_n17549_));
  AOI21_X1   g17357(.A1(new_n17548_), .A2(new_n17549_), .B(new_n3195_), .ZN(new_n17550_));
  NOR3_X1    g17358(.A1(new_n17544_), .A2(\asqrt[42] ), .A3(new_n17550_), .ZN(new_n17551_));
  OAI21_X1   g17359(.A1(new_n17544_), .A2(new_n17550_), .B(\asqrt[42] ), .ZN(new_n17552_));
  OAI21_X1   g17360(.A1(new_n17223_), .A2(new_n17551_), .B(new_n17552_), .ZN(new_n17553_));
  OAI21_X1   g17361(.A1(new_n17553_), .A2(\asqrt[43] ), .B(new_n17219_), .ZN(new_n17554_));
  NAND3_X1   g17362(.A1(new_n17548_), .A2(new_n17549_), .A3(new_n3195_), .ZN(new_n17555_));
  AOI21_X1   g17363(.A1(new_n17225_), .A2(new_n17555_), .B(new_n17550_), .ZN(new_n17556_));
  AOI21_X1   g17364(.A1(new_n17556_), .A2(new_n2960_), .B(new_n17223_), .ZN(new_n17557_));
  NAND2_X1   g17365(.A1(new_n17555_), .A2(new_n17225_), .ZN(new_n17558_));
  INV_X1     g17366(.I(new_n17550_), .ZN(new_n17559_));
  AOI21_X1   g17367(.A1(new_n17558_), .A2(new_n17559_), .B(new_n2960_), .ZN(new_n17560_));
  OAI21_X1   g17368(.A1(new_n17557_), .A2(new_n17560_), .B(\asqrt[43] ), .ZN(new_n17561_));
  NAND3_X1   g17369(.A1(new_n17554_), .A2(new_n2531_), .A3(new_n17561_), .ZN(new_n17562_));
  AOI21_X1   g17370(.A1(new_n17554_), .A2(new_n17561_), .B(new_n2531_), .ZN(new_n17563_));
  AOI21_X1   g17371(.A1(new_n17217_), .A2(new_n17562_), .B(new_n17563_), .ZN(new_n17564_));
  AOI21_X1   g17372(.A1(new_n17564_), .A2(new_n2332_), .B(new_n17214_), .ZN(new_n17565_));
  INV_X1     g17373(.I(new_n17219_), .ZN(new_n17566_));
  NOR3_X1    g17374(.A1(new_n17557_), .A2(\asqrt[43] ), .A3(new_n17560_), .ZN(new_n17567_));
  OAI21_X1   g17375(.A1(new_n17566_), .A2(new_n17567_), .B(new_n17561_), .ZN(new_n17568_));
  OAI21_X1   g17376(.A1(new_n17568_), .A2(\asqrt[44] ), .B(new_n17217_), .ZN(new_n17569_));
  NAND2_X1   g17377(.A1(new_n17568_), .A2(\asqrt[44] ), .ZN(new_n17570_));
  AOI21_X1   g17378(.A1(new_n17569_), .A2(new_n17570_), .B(new_n2332_), .ZN(new_n17571_));
  NOR3_X1    g17379(.A1(new_n17565_), .A2(\asqrt[46] ), .A3(new_n17571_), .ZN(new_n17572_));
  OAI21_X1   g17380(.A1(new_n17565_), .A2(new_n17571_), .B(\asqrt[46] ), .ZN(new_n17573_));
  OAI21_X1   g17381(.A1(new_n17211_), .A2(new_n17572_), .B(new_n17573_), .ZN(new_n17574_));
  OAI21_X1   g17382(.A1(new_n17574_), .A2(\asqrt[47] ), .B(new_n17207_), .ZN(new_n17575_));
  NAND3_X1   g17383(.A1(new_n17569_), .A2(new_n17570_), .A3(new_n2332_), .ZN(new_n17576_));
  AOI21_X1   g17384(.A1(new_n17213_), .A2(new_n17576_), .B(new_n17571_), .ZN(new_n17577_));
  AOI21_X1   g17385(.A1(new_n17577_), .A2(new_n2134_), .B(new_n17211_), .ZN(new_n17578_));
  NAND2_X1   g17386(.A1(new_n17576_), .A2(new_n17213_), .ZN(new_n17579_));
  INV_X1     g17387(.I(new_n17571_), .ZN(new_n17580_));
  AOI21_X1   g17388(.A1(new_n17579_), .A2(new_n17580_), .B(new_n2134_), .ZN(new_n17581_));
  OAI21_X1   g17389(.A1(new_n17578_), .A2(new_n17581_), .B(\asqrt[47] ), .ZN(new_n17582_));
  NAND3_X1   g17390(.A1(new_n17575_), .A2(new_n1778_), .A3(new_n17582_), .ZN(new_n17583_));
  AOI21_X1   g17391(.A1(new_n17575_), .A2(new_n17582_), .B(new_n1778_), .ZN(new_n17584_));
  AOI21_X1   g17392(.A1(new_n17205_), .A2(new_n17583_), .B(new_n17584_), .ZN(new_n17585_));
  AOI21_X1   g17393(.A1(new_n17585_), .A2(new_n1632_), .B(new_n17202_), .ZN(new_n17586_));
  INV_X1     g17394(.I(new_n17207_), .ZN(new_n17587_));
  NOR3_X1    g17395(.A1(new_n17578_), .A2(\asqrt[47] ), .A3(new_n17581_), .ZN(new_n17588_));
  OAI21_X1   g17396(.A1(new_n17587_), .A2(new_n17588_), .B(new_n17582_), .ZN(new_n17589_));
  OAI21_X1   g17397(.A1(new_n17589_), .A2(\asqrt[48] ), .B(new_n17205_), .ZN(new_n17590_));
  NAND2_X1   g17398(.A1(new_n17589_), .A2(\asqrt[48] ), .ZN(new_n17591_));
  AOI21_X1   g17399(.A1(new_n17590_), .A2(new_n17591_), .B(new_n1632_), .ZN(new_n17592_));
  NOR3_X1    g17400(.A1(new_n17586_), .A2(\asqrt[50] ), .A3(new_n17592_), .ZN(new_n17593_));
  OAI21_X1   g17401(.A1(new_n17586_), .A2(new_n17592_), .B(\asqrt[50] ), .ZN(new_n17594_));
  OAI21_X1   g17402(.A1(new_n17199_), .A2(new_n17593_), .B(new_n17594_), .ZN(new_n17595_));
  OAI21_X1   g17403(.A1(new_n17595_), .A2(\asqrt[51] ), .B(new_n17195_), .ZN(new_n17596_));
  NAND3_X1   g17404(.A1(new_n17590_), .A2(new_n17591_), .A3(new_n1632_), .ZN(new_n17597_));
  AOI21_X1   g17405(.A1(new_n17201_), .A2(new_n17597_), .B(new_n17592_), .ZN(new_n17598_));
  AOI21_X1   g17406(.A1(new_n17598_), .A2(new_n1463_), .B(new_n17199_), .ZN(new_n17599_));
  NAND2_X1   g17407(.A1(new_n17597_), .A2(new_n17201_), .ZN(new_n17600_));
  INV_X1     g17408(.I(new_n17592_), .ZN(new_n17601_));
  AOI21_X1   g17409(.A1(new_n17600_), .A2(new_n17601_), .B(new_n1463_), .ZN(new_n17602_));
  OAI21_X1   g17410(.A1(new_n17599_), .A2(new_n17602_), .B(\asqrt[51] ), .ZN(new_n17603_));
  NAND3_X1   g17411(.A1(new_n17596_), .A2(new_n1150_), .A3(new_n17603_), .ZN(new_n17604_));
  AOI21_X1   g17412(.A1(new_n17596_), .A2(new_n17603_), .B(new_n1150_), .ZN(new_n17605_));
  AOI21_X1   g17413(.A1(new_n17193_), .A2(new_n17604_), .B(new_n17605_), .ZN(new_n17606_));
  AOI21_X1   g17414(.A1(new_n17606_), .A2(new_n1006_), .B(new_n17190_), .ZN(new_n17607_));
  INV_X1     g17415(.I(new_n17195_), .ZN(new_n17608_));
  NOR3_X1    g17416(.A1(new_n17599_), .A2(\asqrt[51] ), .A3(new_n17602_), .ZN(new_n17609_));
  OAI21_X1   g17417(.A1(new_n17608_), .A2(new_n17609_), .B(new_n17603_), .ZN(new_n17610_));
  OAI21_X1   g17418(.A1(new_n17610_), .A2(\asqrt[52] ), .B(new_n17193_), .ZN(new_n17611_));
  NAND2_X1   g17419(.A1(new_n17610_), .A2(\asqrt[52] ), .ZN(new_n17612_));
  AOI21_X1   g17420(.A1(new_n17611_), .A2(new_n17612_), .B(new_n1006_), .ZN(new_n17613_));
  NOR3_X1    g17421(.A1(new_n17607_), .A2(\asqrt[54] ), .A3(new_n17613_), .ZN(new_n17614_));
  OAI21_X1   g17422(.A1(new_n17607_), .A2(new_n17613_), .B(\asqrt[54] ), .ZN(new_n17615_));
  OAI21_X1   g17423(.A1(new_n17187_), .A2(new_n17614_), .B(new_n17615_), .ZN(new_n17616_));
  OAI21_X1   g17424(.A1(new_n17616_), .A2(\asqrt[55] ), .B(new_n17183_), .ZN(new_n17617_));
  NAND3_X1   g17425(.A1(new_n17611_), .A2(new_n17612_), .A3(new_n1006_), .ZN(new_n17618_));
  AOI21_X1   g17426(.A1(new_n17189_), .A2(new_n17618_), .B(new_n17613_), .ZN(new_n17619_));
  AOI21_X1   g17427(.A1(new_n17619_), .A2(new_n860_), .B(new_n17187_), .ZN(new_n17620_));
  NAND2_X1   g17428(.A1(new_n17618_), .A2(new_n17189_), .ZN(new_n17621_));
  INV_X1     g17429(.I(new_n17613_), .ZN(new_n17622_));
  AOI21_X1   g17430(.A1(new_n17621_), .A2(new_n17622_), .B(new_n860_), .ZN(new_n17623_));
  OAI21_X1   g17431(.A1(new_n17620_), .A2(new_n17623_), .B(\asqrt[55] ), .ZN(new_n17624_));
  NAND3_X1   g17432(.A1(new_n17617_), .A2(new_n634_), .A3(new_n17624_), .ZN(new_n17625_));
  AOI21_X1   g17433(.A1(new_n17617_), .A2(new_n17624_), .B(new_n634_), .ZN(new_n17626_));
  AOI21_X1   g17434(.A1(new_n17181_), .A2(new_n17625_), .B(new_n17626_), .ZN(new_n17627_));
  AOI21_X1   g17435(.A1(new_n17627_), .A2(new_n531_), .B(new_n17178_), .ZN(new_n17628_));
  INV_X1     g17436(.I(new_n17183_), .ZN(new_n17629_));
  NOR3_X1    g17437(.A1(new_n17620_), .A2(\asqrt[55] ), .A3(new_n17623_), .ZN(new_n17630_));
  OAI21_X1   g17438(.A1(new_n17629_), .A2(new_n17630_), .B(new_n17624_), .ZN(new_n17631_));
  OAI21_X1   g17439(.A1(new_n17631_), .A2(\asqrt[56] ), .B(new_n17181_), .ZN(new_n17632_));
  NAND2_X1   g17440(.A1(new_n17631_), .A2(\asqrt[56] ), .ZN(new_n17633_));
  AOI21_X1   g17441(.A1(new_n17632_), .A2(new_n17633_), .B(new_n531_), .ZN(new_n17634_));
  NOR3_X1    g17442(.A1(new_n17628_), .A2(\asqrt[58] ), .A3(new_n17634_), .ZN(new_n17635_));
  OAI21_X1   g17443(.A1(new_n17628_), .A2(new_n17634_), .B(\asqrt[58] ), .ZN(new_n17636_));
  OAI21_X1   g17444(.A1(new_n17175_), .A2(new_n17635_), .B(new_n17636_), .ZN(new_n17637_));
  OAI21_X1   g17445(.A1(new_n17637_), .A2(\asqrt[59] ), .B(new_n17171_), .ZN(new_n17638_));
  NAND3_X1   g17446(.A1(new_n17632_), .A2(new_n17633_), .A3(new_n531_), .ZN(new_n17639_));
  AOI21_X1   g17447(.A1(new_n17177_), .A2(new_n17639_), .B(new_n17634_), .ZN(new_n17640_));
  AOI21_X1   g17448(.A1(new_n17640_), .A2(new_n423_), .B(new_n17175_), .ZN(new_n17641_));
  NAND2_X1   g17449(.A1(new_n17639_), .A2(new_n17177_), .ZN(new_n17642_));
  INV_X1     g17450(.I(new_n17634_), .ZN(new_n17643_));
  AOI21_X1   g17451(.A1(new_n17642_), .A2(new_n17643_), .B(new_n423_), .ZN(new_n17644_));
  OAI21_X1   g17452(.A1(new_n17641_), .A2(new_n17644_), .B(\asqrt[59] ), .ZN(new_n17645_));
  NAND3_X1   g17453(.A1(new_n17638_), .A2(new_n266_), .A3(new_n17645_), .ZN(new_n17646_));
  INV_X1     g17454(.I(new_n17171_), .ZN(new_n17647_));
  NOR3_X1    g17455(.A1(new_n17641_), .A2(\asqrt[59] ), .A3(new_n17644_), .ZN(new_n17648_));
  NOR2_X1    g17456(.A1(new_n17648_), .A2(new_n17647_), .ZN(new_n17649_));
  INV_X1     g17457(.I(new_n17645_), .ZN(new_n17650_));
  OAI21_X1   g17458(.A1(new_n17649_), .A2(new_n17650_), .B(\asqrt[60] ), .ZN(new_n17651_));
  NOR2_X1    g17459(.A1(\asqrt[5] ), .A2(new_n17126_), .ZN(new_n17652_));
  NOR2_X1    g17460(.A1(new_n17337_), .A2(new_n17126_), .ZN(new_n17653_));
  NOR2_X1    g17461(.A1(new_n17159_), .A2(new_n17125_), .ZN(new_n17654_));
  OAI21_X1   g17462(.A1(new_n17653_), .A2(new_n17654_), .B(\asqrt[63] ), .ZN(new_n17655_));
  NOR2_X1    g17463(.A1(new_n17652_), .A2(new_n17655_), .ZN(new_n17656_));
  INV_X1     g17464(.I(new_n17656_), .ZN(new_n17657_));
  NAND2_X1   g17465(.A1(new_n17334_), .A2(new_n201_), .ZN(new_n17658_));
  AOI21_X1   g17466(.A1(new_n17658_), .A2(new_n17165_), .B(\asqrt[5] ), .ZN(new_n17659_));
  XOR2_X1    g17467(.A1(new_n17659_), .A2(new_n17157_), .Z(new_n17660_));
  INV_X1     g17468(.I(new_n17660_), .ZN(new_n17661_));
  INV_X1     g17469(.I(new_n17169_), .ZN(new_n17662_));
  NOR2_X1    g17470(.A1(new_n17649_), .A2(new_n17650_), .ZN(new_n17663_));
  AOI21_X1   g17471(.A1(new_n17663_), .A2(new_n266_), .B(new_n17662_), .ZN(new_n17664_));
  AOI21_X1   g17472(.A1(new_n17638_), .A2(new_n17645_), .B(new_n266_), .ZN(new_n17665_));
  OAI21_X1   g17473(.A1(new_n17664_), .A2(new_n17665_), .B(\asqrt[61] ), .ZN(new_n17666_));
  AOI21_X1   g17474(.A1(new_n17147_), .A2(new_n17141_), .B(\asqrt[5] ), .ZN(new_n17667_));
  XOR2_X1    g17475(.A1(new_n17667_), .A2(new_n17128_), .Z(new_n17668_));
  OAI21_X1   g17476(.A1(new_n17647_), .A2(new_n17648_), .B(new_n17645_), .ZN(new_n17669_));
  OAI21_X1   g17477(.A1(new_n17669_), .A2(\asqrt[60] ), .B(new_n17169_), .ZN(new_n17670_));
  NAND3_X1   g17478(.A1(new_n17670_), .A2(new_n239_), .A3(new_n17651_), .ZN(new_n17671_));
  NAND2_X1   g17479(.A1(new_n17671_), .A2(new_n17668_), .ZN(new_n17672_));
  NAND2_X1   g17480(.A1(new_n17672_), .A2(new_n17666_), .ZN(new_n17673_));
  AOI21_X1   g17481(.A1(new_n17670_), .A2(new_n17651_), .B(new_n239_), .ZN(new_n17674_));
  AOI21_X1   g17482(.A1(new_n17169_), .A2(new_n17646_), .B(new_n17665_), .ZN(new_n17675_));
  INV_X1     g17483(.I(new_n17668_), .ZN(new_n17676_));
  AOI21_X1   g17484(.A1(new_n17675_), .A2(new_n239_), .B(new_n17676_), .ZN(new_n17677_));
  OAI21_X1   g17485(.A1(new_n17677_), .A2(new_n17674_), .B(new_n201_), .ZN(new_n17678_));
  NAND3_X1   g17486(.A1(new_n17672_), .A2(\asqrt[62] ), .A3(new_n17666_), .ZN(new_n17679_));
  AOI21_X1   g17487(.A1(new_n17140_), .A2(new_n17333_), .B(\asqrt[5] ), .ZN(new_n17680_));
  XOR2_X1    g17488(.A1(new_n17680_), .A2(new_n17144_), .Z(new_n17681_));
  INV_X1     g17489(.I(new_n17681_), .ZN(new_n17682_));
  AOI22_X1   g17490(.A1(new_n17678_), .A2(new_n17679_), .B1(new_n17673_), .B2(new_n17682_), .ZN(new_n17683_));
  NOR2_X1    g17491(.A1(new_n17159_), .A2(new_n17126_), .ZN(new_n17684_));
  OAI21_X1   g17492(.A1(\asqrt[5] ), .A2(new_n17684_), .B(new_n17166_), .ZN(new_n17685_));
  INV_X1     g17493(.I(new_n17685_), .ZN(new_n17686_));
  OAI21_X1   g17494(.A1(new_n17683_), .A2(new_n17661_), .B(new_n17686_), .ZN(new_n17687_));
  OAI21_X1   g17495(.A1(new_n17673_), .A2(\asqrt[62] ), .B(new_n17681_), .ZN(new_n17688_));
  NAND2_X1   g17496(.A1(new_n17673_), .A2(\asqrt[62] ), .ZN(new_n17689_));
  NAND3_X1   g17497(.A1(new_n17688_), .A2(new_n17689_), .A3(new_n17661_), .ZN(new_n17690_));
  NAND4_X1   g17498(.A1(new_n17687_), .A2(new_n193_), .A3(new_n17657_), .A4(new_n17690_), .ZN(\asqrt[4] ));
  AOI21_X1   g17499(.A1(new_n17646_), .A2(new_n17651_), .B(\asqrt[4] ), .ZN(new_n17692_));
  XOR2_X1    g17500(.A1(new_n17692_), .A2(new_n17169_), .Z(new_n17693_));
  INV_X1     g17501(.I(new_n17693_), .ZN(new_n17694_));
  NOR2_X1    g17502(.A1(new_n17650_), .A2(new_n17648_), .ZN(new_n17695_));
  NOR2_X1    g17503(.A1(\asqrt[4] ), .A2(new_n17695_), .ZN(new_n17696_));
  XOR2_X1    g17504(.A1(new_n17696_), .A2(new_n17171_), .Z(new_n17697_));
  NOR2_X1    g17505(.A1(new_n17635_), .A2(new_n17644_), .ZN(new_n17698_));
  NOR2_X1    g17506(.A1(\asqrt[4] ), .A2(new_n17698_), .ZN(new_n17699_));
  XOR2_X1    g17507(.A1(new_n17699_), .A2(new_n17174_), .Z(new_n17700_));
  AOI21_X1   g17508(.A1(new_n17639_), .A2(new_n17643_), .B(\asqrt[4] ), .ZN(new_n17701_));
  XOR2_X1    g17509(.A1(new_n17701_), .A2(new_n17177_), .Z(new_n17702_));
  INV_X1     g17510(.I(new_n17702_), .ZN(new_n17703_));
  AOI21_X1   g17511(.A1(new_n17625_), .A2(new_n17633_), .B(\asqrt[4] ), .ZN(new_n17704_));
  XOR2_X1    g17512(.A1(new_n17704_), .A2(new_n17181_), .Z(new_n17705_));
  INV_X1     g17513(.I(new_n17705_), .ZN(new_n17706_));
  INV_X1     g17514(.I(new_n17624_), .ZN(new_n17707_));
  NOR2_X1    g17515(.A1(new_n17707_), .A2(new_n17630_), .ZN(new_n17708_));
  NOR2_X1    g17516(.A1(\asqrt[4] ), .A2(new_n17708_), .ZN(new_n17709_));
  XOR2_X1    g17517(.A1(new_n17709_), .A2(new_n17183_), .Z(new_n17710_));
  NOR2_X1    g17518(.A1(new_n17614_), .A2(new_n17623_), .ZN(new_n17711_));
  NOR2_X1    g17519(.A1(\asqrt[4] ), .A2(new_n17711_), .ZN(new_n17712_));
  XOR2_X1    g17520(.A1(new_n17712_), .A2(new_n17186_), .Z(new_n17713_));
  AOI21_X1   g17521(.A1(new_n17618_), .A2(new_n17622_), .B(\asqrt[4] ), .ZN(new_n17714_));
  XOR2_X1    g17522(.A1(new_n17714_), .A2(new_n17189_), .Z(new_n17715_));
  INV_X1     g17523(.I(new_n17715_), .ZN(new_n17716_));
  AOI21_X1   g17524(.A1(new_n17604_), .A2(new_n17612_), .B(\asqrt[4] ), .ZN(new_n17717_));
  XOR2_X1    g17525(.A1(new_n17717_), .A2(new_n17193_), .Z(new_n17718_));
  INV_X1     g17526(.I(new_n17718_), .ZN(new_n17719_));
  XOR2_X1    g17527(.A1(new_n17595_), .A2(\asqrt[51] ), .Z(new_n17720_));
  NOR2_X1    g17528(.A1(\asqrt[4] ), .A2(new_n17720_), .ZN(new_n17721_));
  XOR2_X1    g17529(.A1(new_n17721_), .A2(new_n17195_), .Z(new_n17722_));
  NOR2_X1    g17530(.A1(new_n17593_), .A2(new_n17602_), .ZN(new_n17723_));
  NOR2_X1    g17531(.A1(\asqrt[4] ), .A2(new_n17723_), .ZN(new_n17724_));
  XOR2_X1    g17532(.A1(new_n17724_), .A2(new_n17198_), .Z(new_n17725_));
  AOI21_X1   g17533(.A1(new_n17597_), .A2(new_n17601_), .B(\asqrt[4] ), .ZN(new_n17726_));
  XOR2_X1    g17534(.A1(new_n17726_), .A2(new_n17201_), .Z(new_n17727_));
  INV_X1     g17535(.I(new_n17727_), .ZN(new_n17728_));
  AOI21_X1   g17536(.A1(new_n17583_), .A2(new_n17591_), .B(\asqrt[4] ), .ZN(new_n17729_));
  XOR2_X1    g17537(.A1(new_n17729_), .A2(new_n17205_), .Z(new_n17730_));
  INV_X1     g17538(.I(new_n17730_), .ZN(new_n17731_));
  XOR2_X1    g17539(.A1(new_n17574_), .A2(\asqrt[47] ), .Z(new_n17732_));
  NOR2_X1    g17540(.A1(\asqrt[4] ), .A2(new_n17732_), .ZN(new_n17733_));
  XOR2_X1    g17541(.A1(new_n17733_), .A2(new_n17207_), .Z(new_n17734_));
  NOR2_X1    g17542(.A1(new_n17572_), .A2(new_n17581_), .ZN(new_n17735_));
  NOR2_X1    g17543(.A1(\asqrt[4] ), .A2(new_n17735_), .ZN(new_n17736_));
  XOR2_X1    g17544(.A1(new_n17736_), .A2(new_n17210_), .Z(new_n17737_));
  AOI21_X1   g17545(.A1(new_n17576_), .A2(new_n17580_), .B(\asqrt[4] ), .ZN(new_n17738_));
  XOR2_X1    g17546(.A1(new_n17738_), .A2(new_n17213_), .Z(new_n17739_));
  INV_X1     g17547(.I(new_n17739_), .ZN(new_n17740_));
  AOI21_X1   g17548(.A1(new_n17562_), .A2(new_n17570_), .B(\asqrt[4] ), .ZN(new_n17741_));
  XOR2_X1    g17549(.A1(new_n17741_), .A2(new_n17217_), .Z(new_n17742_));
  INV_X1     g17550(.I(new_n17742_), .ZN(new_n17743_));
  XOR2_X1    g17551(.A1(new_n17553_), .A2(\asqrt[43] ), .Z(new_n17744_));
  NOR2_X1    g17552(.A1(\asqrt[4] ), .A2(new_n17744_), .ZN(new_n17745_));
  XOR2_X1    g17553(.A1(new_n17745_), .A2(new_n17219_), .Z(new_n17746_));
  NOR2_X1    g17554(.A1(new_n17551_), .A2(new_n17560_), .ZN(new_n17747_));
  NOR2_X1    g17555(.A1(\asqrt[4] ), .A2(new_n17747_), .ZN(new_n17748_));
  XOR2_X1    g17556(.A1(new_n17748_), .A2(new_n17222_), .Z(new_n17749_));
  AOI21_X1   g17557(.A1(new_n17555_), .A2(new_n17559_), .B(\asqrt[4] ), .ZN(new_n17750_));
  XOR2_X1    g17558(.A1(new_n17750_), .A2(new_n17225_), .Z(new_n17751_));
  INV_X1     g17559(.I(new_n17751_), .ZN(new_n17752_));
  AOI21_X1   g17560(.A1(new_n17541_), .A2(new_n17549_), .B(\asqrt[4] ), .ZN(new_n17753_));
  XOR2_X1    g17561(.A1(new_n17753_), .A2(new_n17229_), .Z(new_n17754_));
  INV_X1     g17562(.I(new_n17754_), .ZN(new_n17755_));
  XOR2_X1    g17563(.A1(new_n17532_), .A2(\asqrt[39] ), .Z(new_n17756_));
  NOR2_X1    g17564(.A1(\asqrt[4] ), .A2(new_n17756_), .ZN(new_n17757_));
  XOR2_X1    g17565(.A1(new_n17757_), .A2(new_n17231_), .Z(new_n17758_));
  NOR2_X1    g17566(.A1(new_n17530_), .A2(new_n17539_), .ZN(new_n17759_));
  NOR2_X1    g17567(.A1(\asqrt[4] ), .A2(new_n17759_), .ZN(new_n17760_));
  XOR2_X1    g17568(.A1(new_n17760_), .A2(new_n17234_), .Z(new_n17761_));
  AOI21_X1   g17569(.A1(new_n17534_), .A2(new_n17538_), .B(\asqrt[4] ), .ZN(new_n17762_));
  XOR2_X1    g17570(.A1(new_n17762_), .A2(new_n17237_), .Z(new_n17763_));
  INV_X1     g17571(.I(new_n17763_), .ZN(new_n17764_));
  AOI21_X1   g17572(.A1(new_n17520_), .A2(new_n17528_), .B(\asqrt[4] ), .ZN(new_n17765_));
  XOR2_X1    g17573(.A1(new_n17765_), .A2(new_n17241_), .Z(new_n17766_));
  INV_X1     g17574(.I(new_n17766_), .ZN(new_n17767_));
  XOR2_X1    g17575(.A1(new_n17511_), .A2(\asqrt[35] ), .Z(new_n17768_));
  NOR2_X1    g17576(.A1(\asqrt[4] ), .A2(new_n17768_), .ZN(new_n17769_));
  XOR2_X1    g17577(.A1(new_n17769_), .A2(new_n17243_), .Z(new_n17770_));
  NOR2_X1    g17578(.A1(new_n17509_), .A2(new_n17518_), .ZN(new_n17771_));
  NOR2_X1    g17579(.A1(\asqrt[4] ), .A2(new_n17771_), .ZN(new_n17772_));
  XOR2_X1    g17580(.A1(new_n17772_), .A2(new_n17246_), .Z(new_n17773_));
  AOI21_X1   g17581(.A1(new_n17513_), .A2(new_n17517_), .B(\asqrt[4] ), .ZN(new_n17774_));
  XOR2_X1    g17582(.A1(new_n17774_), .A2(new_n17249_), .Z(new_n17775_));
  INV_X1     g17583(.I(new_n17775_), .ZN(new_n17776_));
  AOI21_X1   g17584(.A1(new_n17499_), .A2(new_n17507_), .B(\asqrt[4] ), .ZN(new_n17777_));
  XOR2_X1    g17585(.A1(new_n17777_), .A2(new_n17253_), .Z(new_n17778_));
  INV_X1     g17586(.I(new_n17778_), .ZN(new_n17779_));
  XOR2_X1    g17587(.A1(new_n17490_), .A2(\asqrt[31] ), .Z(new_n17780_));
  NOR2_X1    g17588(.A1(\asqrt[4] ), .A2(new_n17780_), .ZN(new_n17781_));
  XOR2_X1    g17589(.A1(new_n17781_), .A2(new_n17255_), .Z(new_n17782_));
  NOR2_X1    g17590(.A1(new_n17488_), .A2(new_n17497_), .ZN(new_n17783_));
  NOR2_X1    g17591(.A1(\asqrt[4] ), .A2(new_n17783_), .ZN(new_n17784_));
  XOR2_X1    g17592(.A1(new_n17784_), .A2(new_n17258_), .Z(new_n17785_));
  AOI21_X1   g17593(.A1(new_n17492_), .A2(new_n17496_), .B(\asqrt[4] ), .ZN(new_n17786_));
  XOR2_X1    g17594(.A1(new_n17786_), .A2(new_n17261_), .Z(new_n17787_));
  INV_X1     g17595(.I(new_n17787_), .ZN(new_n17788_));
  AOI21_X1   g17596(.A1(new_n17478_), .A2(new_n17486_), .B(\asqrt[4] ), .ZN(new_n17789_));
  XOR2_X1    g17597(.A1(new_n17789_), .A2(new_n17265_), .Z(new_n17790_));
  INV_X1     g17598(.I(new_n17790_), .ZN(new_n17791_));
  XOR2_X1    g17599(.A1(new_n17469_), .A2(\asqrt[27] ), .Z(new_n17792_));
  NOR2_X1    g17600(.A1(\asqrt[4] ), .A2(new_n17792_), .ZN(new_n17793_));
  XOR2_X1    g17601(.A1(new_n17793_), .A2(new_n17267_), .Z(new_n17794_));
  NOR2_X1    g17602(.A1(new_n17467_), .A2(new_n17476_), .ZN(new_n17795_));
  NOR2_X1    g17603(.A1(\asqrt[4] ), .A2(new_n17795_), .ZN(new_n17796_));
  XOR2_X1    g17604(.A1(new_n17796_), .A2(new_n17270_), .Z(new_n17797_));
  AOI21_X1   g17605(.A1(new_n17471_), .A2(new_n17475_), .B(\asqrt[4] ), .ZN(new_n17798_));
  XOR2_X1    g17606(.A1(new_n17798_), .A2(new_n17273_), .Z(new_n17799_));
  INV_X1     g17607(.I(new_n17799_), .ZN(new_n17800_));
  AOI21_X1   g17608(.A1(new_n17457_), .A2(new_n17465_), .B(\asqrt[4] ), .ZN(new_n17801_));
  XOR2_X1    g17609(.A1(new_n17801_), .A2(new_n17277_), .Z(new_n17802_));
  INV_X1     g17610(.I(new_n17802_), .ZN(new_n17803_));
  XOR2_X1    g17611(.A1(new_n17448_), .A2(\asqrt[23] ), .Z(new_n17804_));
  NOR2_X1    g17612(.A1(\asqrt[4] ), .A2(new_n17804_), .ZN(new_n17805_));
  XOR2_X1    g17613(.A1(new_n17805_), .A2(new_n17279_), .Z(new_n17806_));
  NOR2_X1    g17614(.A1(new_n17446_), .A2(new_n17455_), .ZN(new_n17807_));
  NOR2_X1    g17615(.A1(\asqrt[4] ), .A2(new_n17807_), .ZN(new_n17808_));
  XOR2_X1    g17616(.A1(new_n17808_), .A2(new_n17282_), .Z(new_n17809_));
  AOI21_X1   g17617(.A1(new_n17450_), .A2(new_n17454_), .B(\asqrt[4] ), .ZN(new_n17810_));
  XOR2_X1    g17618(.A1(new_n17810_), .A2(new_n17285_), .Z(new_n17811_));
  INV_X1     g17619(.I(new_n17811_), .ZN(new_n17812_));
  AOI21_X1   g17620(.A1(new_n17436_), .A2(new_n17444_), .B(\asqrt[4] ), .ZN(new_n17813_));
  XOR2_X1    g17621(.A1(new_n17813_), .A2(new_n17289_), .Z(new_n17814_));
  INV_X1     g17622(.I(new_n17814_), .ZN(new_n17815_));
  XOR2_X1    g17623(.A1(new_n17427_), .A2(\asqrt[19] ), .Z(new_n17816_));
  NOR2_X1    g17624(.A1(\asqrt[4] ), .A2(new_n17816_), .ZN(new_n17817_));
  XOR2_X1    g17625(.A1(new_n17817_), .A2(new_n17291_), .Z(new_n17818_));
  NOR2_X1    g17626(.A1(new_n17425_), .A2(new_n17434_), .ZN(new_n17819_));
  NOR2_X1    g17627(.A1(\asqrt[4] ), .A2(new_n17819_), .ZN(new_n17820_));
  XOR2_X1    g17628(.A1(new_n17820_), .A2(new_n17294_), .Z(new_n17821_));
  AOI21_X1   g17629(.A1(new_n17429_), .A2(new_n17433_), .B(\asqrt[4] ), .ZN(new_n17822_));
  XOR2_X1    g17630(.A1(new_n17822_), .A2(new_n17297_), .Z(new_n17823_));
  INV_X1     g17631(.I(new_n17823_), .ZN(new_n17824_));
  AOI21_X1   g17632(.A1(new_n17415_), .A2(new_n17423_), .B(\asqrt[4] ), .ZN(new_n17825_));
  XOR2_X1    g17633(.A1(new_n17825_), .A2(new_n17301_), .Z(new_n17826_));
  INV_X1     g17634(.I(new_n17826_), .ZN(new_n17827_));
  XOR2_X1    g17635(.A1(new_n17406_), .A2(\asqrt[15] ), .Z(new_n17828_));
  NOR2_X1    g17636(.A1(\asqrt[4] ), .A2(new_n17828_), .ZN(new_n17829_));
  XOR2_X1    g17637(.A1(new_n17829_), .A2(new_n17303_), .Z(new_n17830_));
  NOR2_X1    g17638(.A1(new_n17404_), .A2(new_n17413_), .ZN(new_n17831_));
  NOR2_X1    g17639(.A1(\asqrt[4] ), .A2(new_n17831_), .ZN(new_n17832_));
  XOR2_X1    g17640(.A1(new_n17832_), .A2(new_n17306_), .Z(new_n17833_));
  AOI21_X1   g17641(.A1(new_n17408_), .A2(new_n17412_), .B(\asqrt[4] ), .ZN(new_n17834_));
  XOR2_X1    g17642(.A1(new_n17834_), .A2(new_n17309_), .Z(new_n17835_));
  INV_X1     g17643(.I(new_n17835_), .ZN(new_n17836_));
  AOI21_X1   g17644(.A1(new_n17394_), .A2(new_n17402_), .B(\asqrt[4] ), .ZN(new_n17837_));
  XOR2_X1    g17645(.A1(new_n17837_), .A2(new_n17313_), .Z(new_n17838_));
  INV_X1     g17646(.I(new_n17838_), .ZN(new_n17839_));
  XOR2_X1    g17647(.A1(new_n17385_), .A2(\asqrt[11] ), .Z(new_n17840_));
  NOR2_X1    g17648(.A1(\asqrt[4] ), .A2(new_n17840_), .ZN(new_n17841_));
  XOR2_X1    g17649(.A1(new_n17841_), .A2(new_n17315_), .Z(new_n17842_));
  NOR2_X1    g17650(.A1(new_n17383_), .A2(new_n17392_), .ZN(new_n17843_));
  NOR2_X1    g17651(.A1(\asqrt[4] ), .A2(new_n17843_), .ZN(new_n17844_));
  XOR2_X1    g17652(.A1(new_n17844_), .A2(new_n17318_), .Z(new_n17845_));
  AOI21_X1   g17653(.A1(new_n17387_), .A2(new_n17391_), .B(\asqrt[4] ), .ZN(new_n17846_));
  XOR2_X1    g17654(.A1(new_n17846_), .A2(new_n17321_), .Z(new_n17847_));
  INV_X1     g17655(.I(new_n17847_), .ZN(new_n17848_));
  AOI21_X1   g17656(.A1(new_n17373_), .A2(new_n17381_), .B(\asqrt[4] ), .ZN(new_n17849_));
  XOR2_X1    g17657(.A1(new_n17849_), .A2(new_n17328_), .Z(new_n17850_));
  INV_X1     g17658(.I(new_n17850_), .ZN(new_n17851_));
  AOI21_X1   g17659(.A1(new_n17363_), .A2(new_n17372_), .B(\asqrt[4] ), .ZN(new_n17852_));
  XOR2_X1    g17660(.A1(new_n17852_), .A2(new_n17345_), .Z(new_n17853_));
  NOR2_X1    g17661(.A1(new_n17342_), .A2(\a[10] ), .ZN(new_n17854_));
  INV_X1     g17662(.I(new_n17854_), .ZN(new_n17855_));
  NOR2_X1    g17663(.A1(new_n17352_), .A2(\a[10] ), .ZN(new_n17856_));
  AOI22_X1   g17664(.A1(new_n17855_), .A2(new_n17352_), .B1(\asqrt[5] ), .B2(new_n17856_), .ZN(new_n17857_));
  INV_X1     g17665(.I(new_n17857_), .ZN(new_n17858_));
  AOI21_X1   g17666(.A1(new_n17668_), .A2(new_n17671_), .B(new_n17674_), .ZN(new_n17859_));
  AOI21_X1   g17667(.A1(new_n17672_), .A2(new_n17666_), .B(\asqrt[62] ), .ZN(new_n17860_));
  NOR3_X1    g17668(.A1(new_n17677_), .A2(new_n201_), .A3(new_n17674_), .ZN(new_n17861_));
  OAI22_X1   g17669(.A1(new_n17861_), .A2(new_n17860_), .B1(new_n17859_), .B2(new_n17681_), .ZN(new_n17862_));
  AOI21_X1   g17670(.A1(new_n17862_), .A2(new_n17660_), .B(new_n17685_), .ZN(new_n17863_));
  NAND2_X1   g17671(.A1(new_n17859_), .A2(new_n201_), .ZN(new_n17864_));
  OAI21_X1   g17672(.A1(new_n17859_), .A2(new_n201_), .B(new_n17661_), .ZN(new_n17865_));
  AOI21_X1   g17673(.A1(new_n17681_), .A2(new_n17864_), .B(new_n17865_), .ZN(new_n17866_));
  NOR4_X1    g17674(.A1(new_n17863_), .A2(\asqrt[63] ), .A3(new_n17656_), .A4(new_n17866_), .ZN(new_n17867_));
  NOR2_X1    g17675(.A1(new_n17367_), .A2(new_n17361_), .ZN(new_n17868_));
  NOR2_X1    g17676(.A1(new_n17867_), .A2(new_n17868_), .ZN(new_n17869_));
  NOR2_X1    g17677(.A1(new_n17869_), .A2(new_n17858_), .ZN(new_n17870_));
  NOR3_X1    g17678(.A1(new_n17867_), .A2(new_n17857_), .A3(new_n17868_), .ZN(new_n17871_));
  NOR2_X1    g17679(.A1(new_n17870_), .A2(new_n17871_), .ZN(new_n17872_));
  NOR2_X1    g17680(.A1(new_n17656_), .A2(new_n17342_), .ZN(new_n17873_));
  NAND4_X1   g17681(.A1(new_n17687_), .A2(new_n193_), .A3(new_n17690_), .A4(new_n17873_), .ZN(new_n17874_));
  NAND2_X1   g17682(.A1(\asqrt[4] ), .A2(new_n17347_), .ZN(new_n17875_));
  AOI21_X1   g17683(.A1(new_n17875_), .A2(new_n17874_), .B(\a[10] ), .ZN(new_n17876_));
  INV_X1     g17684(.I(new_n17876_), .ZN(new_n17877_));
  NAND3_X1   g17685(.A1(new_n17875_), .A2(\a[10] ), .A3(new_n17874_), .ZN(new_n17878_));
  NAND2_X1   g17686(.A1(new_n17877_), .A2(new_n17878_), .ZN(new_n17879_));
  NOR2_X1    g17687(.A1(\a[6] ), .A2(\a[7] ), .ZN(new_n17880_));
  INV_X1     g17688(.I(new_n17880_), .ZN(new_n17881_));
  NAND3_X1   g17689(.A1(\asqrt[4] ), .A2(\a[8] ), .A3(new_n17881_), .ZN(new_n17882_));
  INV_X1     g17690(.I(\a[8] ), .ZN(new_n17883_));
  OAI21_X1   g17691(.A1(\asqrt[4] ), .A2(new_n17883_), .B(new_n17880_), .ZN(new_n17884_));
  AOI21_X1   g17692(.A1(new_n17884_), .A2(new_n17882_), .B(new_n17342_), .ZN(new_n17885_));
  OAI21_X1   g17693(.A1(new_n17867_), .A2(\a[8] ), .B(\a[9] ), .ZN(new_n17886_));
  INV_X1     g17694(.I(\a[9] ), .ZN(new_n17887_));
  NAND3_X1   g17695(.A1(\asqrt[4] ), .A2(new_n17883_), .A3(new_n17887_), .ZN(new_n17888_));
  NOR3_X1    g17696(.A1(new_n17338_), .A2(\asqrt[63] ), .A3(new_n17341_), .ZN(new_n17889_));
  AOI21_X1   g17697(.A1(new_n17889_), .A2(new_n17123_), .B(new_n17883_), .ZN(new_n17890_));
  NAND2_X1   g17698(.A1(\asqrt[4] ), .A2(new_n17890_), .ZN(new_n17891_));
  NAND3_X1   g17699(.A1(new_n17886_), .A2(new_n17888_), .A3(new_n17891_), .ZN(new_n17892_));
  NOR3_X1    g17700(.A1(new_n17885_), .A2(new_n17892_), .A3(\asqrt[6] ), .ZN(new_n17893_));
  OAI21_X1   g17701(.A1(new_n17885_), .A2(new_n17892_), .B(\asqrt[6] ), .ZN(new_n17894_));
  OAI21_X1   g17702(.A1(new_n17879_), .A2(new_n17893_), .B(new_n17894_), .ZN(new_n17895_));
  OAI21_X1   g17703(.A1(new_n17895_), .A2(\asqrt[7] ), .B(new_n17872_), .ZN(new_n17896_));
  NAND2_X1   g17704(.A1(new_n17895_), .A2(\asqrt[7] ), .ZN(new_n17897_));
  NAND3_X1   g17705(.A1(new_n17896_), .A2(new_n17897_), .A3(new_n15717_), .ZN(new_n17898_));
  AOI21_X1   g17706(.A1(new_n17896_), .A2(new_n17897_), .B(new_n15717_), .ZN(new_n17899_));
  AOI21_X1   g17707(.A1(new_n17853_), .A2(new_n17898_), .B(new_n17899_), .ZN(new_n17900_));
  AOI21_X1   g17708(.A1(new_n17900_), .A2(new_n15221_), .B(new_n17851_), .ZN(new_n17901_));
  NAND2_X1   g17709(.A1(new_n17898_), .A2(new_n17853_), .ZN(new_n17902_));
  INV_X1     g17710(.I(new_n17872_), .ZN(new_n17903_));
  INV_X1     g17711(.I(new_n17878_), .ZN(new_n17904_));
  NOR2_X1    g17712(.A1(new_n17904_), .A2(new_n17876_), .ZN(new_n17905_));
  NOR3_X1    g17713(.A1(new_n17867_), .A2(new_n17883_), .A3(new_n17880_), .ZN(new_n17906_));
  AOI21_X1   g17714(.A1(new_n17867_), .A2(\a[8] ), .B(new_n17881_), .ZN(new_n17907_));
  OAI21_X1   g17715(.A1(new_n17906_), .A2(new_n17907_), .B(\asqrt[5] ), .ZN(new_n17908_));
  AOI21_X1   g17716(.A1(\asqrt[4] ), .A2(new_n17883_), .B(new_n17887_), .ZN(new_n17909_));
  NOR3_X1    g17717(.A1(new_n17867_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n17910_));
  INV_X1     g17718(.I(new_n17890_), .ZN(new_n17911_));
  NOR2_X1    g17719(.A1(new_n17867_), .A2(new_n17911_), .ZN(new_n17912_));
  NOR3_X1    g17720(.A1(new_n17910_), .A2(new_n17909_), .A3(new_n17912_), .ZN(new_n17913_));
  NAND3_X1   g17721(.A1(new_n17908_), .A2(new_n17913_), .A3(new_n16779_), .ZN(new_n17914_));
  AOI21_X1   g17722(.A1(new_n17908_), .A2(new_n17913_), .B(new_n16779_), .ZN(new_n17915_));
  AOI21_X1   g17723(.A1(new_n17905_), .A2(new_n17914_), .B(new_n17915_), .ZN(new_n17916_));
  AOI21_X1   g17724(.A1(new_n17916_), .A2(new_n16269_), .B(new_n17903_), .ZN(new_n17917_));
  NOR2_X1    g17725(.A1(new_n17916_), .A2(new_n16269_), .ZN(new_n17918_));
  OAI21_X1   g17726(.A1(new_n17917_), .A2(new_n17918_), .B(\asqrt[8] ), .ZN(new_n17919_));
  AOI21_X1   g17727(.A1(new_n17902_), .A2(new_n17919_), .B(new_n15221_), .ZN(new_n17920_));
  NOR3_X1    g17728(.A1(new_n17901_), .A2(\asqrt[10] ), .A3(new_n17920_), .ZN(new_n17921_));
  OAI21_X1   g17729(.A1(new_n17901_), .A2(new_n17920_), .B(\asqrt[10] ), .ZN(new_n17922_));
  OAI21_X1   g17730(.A1(new_n17848_), .A2(new_n17921_), .B(new_n17922_), .ZN(new_n17923_));
  OAI21_X1   g17731(.A1(new_n17923_), .A2(\asqrt[11] ), .B(new_n17845_), .ZN(new_n17924_));
  NAND2_X1   g17732(.A1(new_n17923_), .A2(\asqrt[11] ), .ZN(new_n17925_));
  NAND3_X1   g17733(.A1(new_n17924_), .A2(new_n17925_), .A3(new_n13690_), .ZN(new_n17926_));
  AOI21_X1   g17734(.A1(new_n17924_), .A2(new_n17925_), .B(new_n13690_), .ZN(new_n17927_));
  AOI21_X1   g17735(.A1(new_n17842_), .A2(new_n17926_), .B(new_n17927_), .ZN(new_n17928_));
  AOI21_X1   g17736(.A1(new_n17928_), .A2(new_n13228_), .B(new_n17839_), .ZN(new_n17929_));
  NAND2_X1   g17737(.A1(new_n17926_), .A2(new_n17842_), .ZN(new_n17930_));
  INV_X1     g17738(.I(new_n17845_), .ZN(new_n17931_));
  INV_X1     g17739(.I(new_n17853_), .ZN(new_n17932_));
  NOR3_X1    g17740(.A1(new_n17917_), .A2(new_n17918_), .A3(\asqrt[8] ), .ZN(new_n17933_));
  OAI21_X1   g17741(.A1(new_n17932_), .A2(new_n17933_), .B(new_n17919_), .ZN(new_n17934_));
  OAI21_X1   g17742(.A1(new_n17934_), .A2(\asqrt[9] ), .B(new_n17850_), .ZN(new_n17935_));
  NAND2_X1   g17743(.A1(new_n17934_), .A2(\asqrt[9] ), .ZN(new_n17936_));
  NAND3_X1   g17744(.A1(new_n17935_), .A2(new_n17936_), .A3(new_n14690_), .ZN(new_n17937_));
  AOI21_X1   g17745(.A1(new_n17935_), .A2(new_n17936_), .B(new_n14690_), .ZN(new_n17938_));
  AOI21_X1   g17746(.A1(new_n17847_), .A2(new_n17937_), .B(new_n17938_), .ZN(new_n17939_));
  AOI21_X1   g17747(.A1(new_n17939_), .A2(new_n14207_), .B(new_n17931_), .ZN(new_n17940_));
  NOR2_X1    g17748(.A1(new_n17939_), .A2(new_n14207_), .ZN(new_n17941_));
  OAI21_X1   g17749(.A1(new_n17940_), .A2(new_n17941_), .B(\asqrt[12] ), .ZN(new_n17942_));
  AOI21_X1   g17750(.A1(new_n17930_), .A2(new_n17942_), .B(new_n13228_), .ZN(new_n17943_));
  NOR3_X1    g17751(.A1(new_n17929_), .A2(\asqrt[14] ), .A3(new_n17943_), .ZN(new_n17944_));
  OAI21_X1   g17752(.A1(new_n17929_), .A2(new_n17943_), .B(\asqrt[14] ), .ZN(new_n17945_));
  OAI21_X1   g17753(.A1(new_n17836_), .A2(new_n17944_), .B(new_n17945_), .ZN(new_n17946_));
  OAI21_X1   g17754(.A1(new_n17946_), .A2(\asqrt[15] ), .B(new_n17833_), .ZN(new_n17947_));
  NAND2_X1   g17755(.A1(new_n17946_), .A2(\asqrt[15] ), .ZN(new_n17948_));
  NAND3_X1   g17756(.A1(new_n17947_), .A2(new_n17948_), .A3(new_n11802_), .ZN(new_n17949_));
  AOI21_X1   g17757(.A1(new_n17947_), .A2(new_n17948_), .B(new_n11802_), .ZN(new_n17950_));
  AOI21_X1   g17758(.A1(new_n17830_), .A2(new_n17949_), .B(new_n17950_), .ZN(new_n17951_));
  AOI21_X1   g17759(.A1(new_n17951_), .A2(new_n11373_), .B(new_n17827_), .ZN(new_n17952_));
  NAND2_X1   g17760(.A1(new_n17949_), .A2(new_n17830_), .ZN(new_n17953_));
  INV_X1     g17761(.I(new_n17833_), .ZN(new_n17954_));
  INV_X1     g17762(.I(new_n17842_), .ZN(new_n17955_));
  NOR3_X1    g17763(.A1(new_n17940_), .A2(new_n17941_), .A3(\asqrt[12] ), .ZN(new_n17956_));
  OAI21_X1   g17764(.A1(new_n17955_), .A2(new_n17956_), .B(new_n17942_), .ZN(new_n17957_));
  OAI21_X1   g17765(.A1(new_n17957_), .A2(\asqrt[13] ), .B(new_n17838_), .ZN(new_n17958_));
  NAND2_X1   g17766(.A1(new_n17957_), .A2(\asqrt[13] ), .ZN(new_n17959_));
  NAND3_X1   g17767(.A1(new_n17958_), .A2(new_n17959_), .A3(new_n12733_), .ZN(new_n17960_));
  AOI21_X1   g17768(.A1(new_n17958_), .A2(new_n17959_), .B(new_n12733_), .ZN(new_n17961_));
  AOI21_X1   g17769(.A1(new_n17835_), .A2(new_n17960_), .B(new_n17961_), .ZN(new_n17962_));
  AOI21_X1   g17770(.A1(new_n17962_), .A2(new_n12283_), .B(new_n17954_), .ZN(new_n17963_));
  NOR2_X1    g17771(.A1(new_n17962_), .A2(new_n12283_), .ZN(new_n17964_));
  OAI21_X1   g17772(.A1(new_n17963_), .A2(new_n17964_), .B(\asqrt[16] ), .ZN(new_n17965_));
  AOI21_X1   g17773(.A1(new_n17953_), .A2(new_n17965_), .B(new_n11373_), .ZN(new_n17966_));
  NOR3_X1    g17774(.A1(new_n17952_), .A2(\asqrt[18] ), .A3(new_n17966_), .ZN(new_n17967_));
  OAI21_X1   g17775(.A1(new_n17952_), .A2(new_n17966_), .B(\asqrt[18] ), .ZN(new_n17968_));
  OAI21_X1   g17776(.A1(new_n17824_), .A2(new_n17967_), .B(new_n17968_), .ZN(new_n17969_));
  OAI21_X1   g17777(.A1(new_n17969_), .A2(\asqrt[19] ), .B(new_n17821_), .ZN(new_n17970_));
  NAND2_X1   g17778(.A1(new_n17969_), .A2(\asqrt[19] ), .ZN(new_n17971_));
  NAND3_X1   g17779(.A1(new_n17970_), .A2(new_n17971_), .A3(new_n10052_), .ZN(new_n17972_));
  AOI21_X1   g17780(.A1(new_n17970_), .A2(new_n17971_), .B(new_n10052_), .ZN(new_n17973_));
  AOI21_X1   g17781(.A1(new_n17818_), .A2(new_n17972_), .B(new_n17973_), .ZN(new_n17974_));
  AOI21_X1   g17782(.A1(new_n17974_), .A2(new_n9656_), .B(new_n17815_), .ZN(new_n17975_));
  NAND2_X1   g17783(.A1(new_n17972_), .A2(new_n17818_), .ZN(new_n17976_));
  INV_X1     g17784(.I(new_n17821_), .ZN(new_n17977_));
  INV_X1     g17785(.I(new_n17830_), .ZN(new_n17978_));
  NOR3_X1    g17786(.A1(new_n17963_), .A2(new_n17964_), .A3(\asqrt[16] ), .ZN(new_n17979_));
  OAI21_X1   g17787(.A1(new_n17978_), .A2(new_n17979_), .B(new_n17965_), .ZN(new_n17980_));
  OAI21_X1   g17788(.A1(new_n17980_), .A2(\asqrt[17] ), .B(new_n17826_), .ZN(new_n17981_));
  NAND2_X1   g17789(.A1(new_n17980_), .A2(\asqrt[17] ), .ZN(new_n17982_));
  NAND3_X1   g17790(.A1(new_n17981_), .A2(new_n17982_), .A3(new_n10914_), .ZN(new_n17983_));
  AOI21_X1   g17791(.A1(new_n17981_), .A2(new_n17982_), .B(new_n10914_), .ZN(new_n17984_));
  AOI21_X1   g17792(.A1(new_n17823_), .A2(new_n17983_), .B(new_n17984_), .ZN(new_n17985_));
  AOI21_X1   g17793(.A1(new_n17985_), .A2(new_n10497_), .B(new_n17977_), .ZN(new_n17986_));
  NOR2_X1    g17794(.A1(new_n17985_), .A2(new_n10497_), .ZN(new_n17987_));
  OAI21_X1   g17795(.A1(new_n17986_), .A2(new_n17987_), .B(\asqrt[20] ), .ZN(new_n17988_));
  AOI21_X1   g17796(.A1(new_n17976_), .A2(new_n17988_), .B(new_n9656_), .ZN(new_n17989_));
  NOR3_X1    g17797(.A1(new_n17975_), .A2(\asqrt[22] ), .A3(new_n17989_), .ZN(new_n17990_));
  OAI21_X1   g17798(.A1(new_n17975_), .A2(new_n17989_), .B(\asqrt[22] ), .ZN(new_n17991_));
  OAI21_X1   g17799(.A1(new_n17812_), .A2(new_n17990_), .B(new_n17991_), .ZN(new_n17992_));
  OAI21_X1   g17800(.A1(new_n17992_), .A2(\asqrt[23] ), .B(new_n17809_), .ZN(new_n17993_));
  NAND2_X1   g17801(.A1(new_n17992_), .A2(\asqrt[23] ), .ZN(new_n17994_));
  NAND3_X1   g17802(.A1(new_n17993_), .A2(new_n17994_), .A3(new_n8440_), .ZN(new_n17995_));
  AOI21_X1   g17803(.A1(new_n17993_), .A2(new_n17994_), .B(new_n8440_), .ZN(new_n17996_));
  AOI21_X1   g17804(.A1(new_n17806_), .A2(new_n17995_), .B(new_n17996_), .ZN(new_n17997_));
  AOI21_X1   g17805(.A1(new_n17997_), .A2(new_n8077_), .B(new_n17803_), .ZN(new_n17998_));
  NAND2_X1   g17806(.A1(new_n17995_), .A2(new_n17806_), .ZN(new_n17999_));
  INV_X1     g17807(.I(new_n17809_), .ZN(new_n18000_));
  INV_X1     g17808(.I(new_n17818_), .ZN(new_n18001_));
  NOR3_X1    g17809(.A1(new_n17986_), .A2(new_n17987_), .A3(\asqrt[20] ), .ZN(new_n18002_));
  OAI21_X1   g17810(.A1(new_n18001_), .A2(new_n18002_), .B(new_n17988_), .ZN(new_n18003_));
  OAI21_X1   g17811(.A1(new_n18003_), .A2(\asqrt[21] ), .B(new_n17814_), .ZN(new_n18004_));
  NAND2_X1   g17812(.A1(new_n18003_), .A2(\asqrt[21] ), .ZN(new_n18005_));
  NAND3_X1   g17813(.A1(new_n18004_), .A2(new_n18005_), .A3(new_n9233_), .ZN(new_n18006_));
  AOI21_X1   g17814(.A1(new_n18004_), .A2(new_n18005_), .B(new_n9233_), .ZN(new_n18007_));
  AOI21_X1   g17815(.A1(new_n17811_), .A2(new_n18006_), .B(new_n18007_), .ZN(new_n18008_));
  AOI21_X1   g17816(.A1(new_n18008_), .A2(new_n8849_), .B(new_n18000_), .ZN(new_n18009_));
  NOR2_X1    g17817(.A1(new_n18008_), .A2(new_n8849_), .ZN(new_n18010_));
  OAI21_X1   g17818(.A1(new_n18009_), .A2(new_n18010_), .B(\asqrt[24] ), .ZN(new_n18011_));
  AOI21_X1   g17819(.A1(new_n17999_), .A2(new_n18011_), .B(new_n8077_), .ZN(new_n18012_));
  NOR3_X1    g17820(.A1(new_n17998_), .A2(\asqrt[26] ), .A3(new_n18012_), .ZN(new_n18013_));
  OAI21_X1   g17821(.A1(new_n17998_), .A2(new_n18012_), .B(\asqrt[26] ), .ZN(new_n18014_));
  OAI21_X1   g17822(.A1(new_n17800_), .A2(new_n18013_), .B(new_n18014_), .ZN(new_n18015_));
  OAI21_X1   g17823(.A1(new_n18015_), .A2(\asqrt[27] ), .B(new_n17797_), .ZN(new_n18016_));
  NAND2_X1   g17824(.A1(new_n18015_), .A2(\asqrt[27] ), .ZN(new_n18017_));
  NAND3_X1   g17825(.A1(new_n18016_), .A2(new_n18017_), .A3(new_n6966_), .ZN(new_n18018_));
  AOI21_X1   g17826(.A1(new_n18016_), .A2(new_n18017_), .B(new_n6966_), .ZN(new_n18019_));
  AOI21_X1   g17827(.A1(new_n17794_), .A2(new_n18018_), .B(new_n18019_), .ZN(new_n18020_));
  AOI21_X1   g17828(.A1(new_n18020_), .A2(new_n6636_), .B(new_n17791_), .ZN(new_n18021_));
  NAND2_X1   g17829(.A1(new_n18018_), .A2(new_n17794_), .ZN(new_n18022_));
  INV_X1     g17830(.I(new_n17797_), .ZN(new_n18023_));
  INV_X1     g17831(.I(new_n17806_), .ZN(new_n18024_));
  NOR3_X1    g17832(.A1(new_n18009_), .A2(new_n18010_), .A3(\asqrt[24] ), .ZN(new_n18025_));
  OAI21_X1   g17833(.A1(new_n18024_), .A2(new_n18025_), .B(new_n18011_), .ZN(new_n18026_));
  OAI21_X1   g17834(.A1(new_n18026_), .A2(\asqrt[25] ), .B(new_n17802_), .ZN(new_n18027_));
  NAND2_X1   g17835(.A1(new_n18026_), .A2(\asqrt[25] ), .ZN(new_n18028_));
  NAND3_X1   g17836(.A1(new_n18027_), .A2(new_n18028_), .A3(new_n7690_), .ZN(new_n18029_));
  AOI21_X1   g17837(.A1(new_n18027_), .A2(new_n18028_), .B(new_n7690_), .ZN(new_n18030_));
  AOI21_X1   g17838(.A1(new_n17799_), .A2(new_n18029_), .B(new_n18030_), .ZN(new_n18031_));
  AOI21_X1   g17839(.A1(new_n18031_), .A2(new_n7331_), .B(new_n18023_), .ZN(new_n18032_));
  NOR2_X1    g17840(.A1(new_n18031_), .A2(new_n7331_), .ZN(new_n18033_));
  OAI21_X1   g17841(.A1(new_n18032_), .A2(new_n18033_), .B(\asqrt[28] ), .ZN(new_n18034_));
  AOI21_X1   g17842(.A1(new_n18022_), .A2(new_n18034_), .B(new_n6636_), .ZN(new_n18035_));
  NOR3_X1    g17843(.A1(new_n18021_), .A2(\asqrt[30] ), .A3(new_n18035_), .ZN(new_n18036_));
  OAI21_X1   g17844(.A1(new_n18021_), .A2(new_n18035_), .B(\asqrt[30] ), .ZN(new_n18037_));
  OAI21_X1   g17845(.A1(new_n17788_), .A2(new_n18036_), .B(new_n18037_), .ZN(new_n18038_));
  OAI21_X1   g17846(.A1(new_n18038_), .A2(\asqrt[31] ), .B(new_n17785_), .ZN(new_n18039_));
  NAND2_X1   g17847(.A1(new_n18038_), .A2(\asqrt[31] ), .ZN(new_n18040_));
  NAND3_X1   g17848(.A1(new_n18039_), .A2(new_n18040_), .A3(new_n5643_), .ZN(new_n18041_));
  AOI21_X1   g17849(.A1(new_n18039_), .A2(new_n18040_), .B(new_n5643_), .ZN(new_n18042_));
  AOI21_X1   g17850(.A1(new_n17782_), .A2(new_n18041_), .B(new_n18042_), .ZN(new_n18043_));
  AOI21_X1   g17851(.A1(new_n18043_), .A2(new_n5336_), .B(new_n17779_), .ZN(new_n18044_));
  NAND2_X1   g17852(.A1(new_n18041_), .A2(new_n17782_), .ZN(new_n18045_));
  INV_X1     g17853(.I(new_n17785_), .ZN(new_n18046_));
  INV_X1     g17854(.I(new_n17794_), .ZN(new_n18047_));
  NOR3_X1    g17855(.A1(new_n18032_), .A2(new_n18033_), .A3(\asqrt[28] ), .ZN(new_n18048_));
  OAI21_X1   g17856(.A1(new_n18047_), .A2(new_n18048_), .B(new_n18034_), .ZN(new_n18049_));
  OAI21_X1   g17857(.A1(new_n18049_), .A2(\asqrt[29] ), .B(new_n17790_), .ZN(new_n18050_));
  NAND2_X1   g17858(.A1(new_n18049_), .A2(\asqrt[29] ), .ZN(new_n18051_));
  NAND3_X1   g17859(.A1(new_n18050_), .A2(new_n18051_), .A3(new_n6275_), .ZN(new_n18052_));
  AOI21_X1   g17860(.A1(new_n18050_), .A2(new_n18051_), .B(new_n6275_), .ZN(new_n18053_));
  AOI21_X1   g17861(.A1(new_n17787_), .A2(new_n18052_), .B(new_n18053_), .ZN(new_n18054_));
  AOI21_X1   g17862(.A1(new_n18054_), .A2(new_n5947_), .B(new_n18046_), .ZN(new_n18055_));
  NOR2_X1    g17863(.A1(new_n18054_), .A2(new_n5947_), .ZN(new_n18056_));
  OAI21_X1   g17864(.A1(new_n18055_), .A2(new_n18056_), .B(\asqrt[32] ), .ZN(new_n18057_));
  AOI21_X1   g17865(.A1(new_n18045_), .A2(new_n18057_), .B(new_n5336_), .ZN(new_n18058_));
  NOR3_X1    g17866(.A1(new_n18044_), .A2(\asqrt[34] ), .A3(new_n18058_), .ZN(new_n18059_));
  OAI21_X1   g17867(.A1(new_n18044_), .A2(new_n18058_), .B(\asqrt[34] ), .ZN(new_n18060_));
  OAI21_X1   g17868(.A1(new_n17776_), .A2(new_n18059_), .B(new_n18060_), .ZN(new_n18061_));
  OAI21_X1   g17869(.A1(new_n18061_), .A2(\asqrt[35] ), .B(new_n17773_), .ZN(new_n18062_));
  NAND2_X1   g17870(.A1(new_n18061_), .A2(\asqrt[35] ), .ZN(new_n18063_));
  NAND3_X1   g17871(.A1(new_n18062_), .A2(new_n18063_), .A3(new_n4461_), .ZN(new_n18064_));
  AOI21_X1   g17872(.A1(new_n18062_), .A2(new_n18063_), .B(new_n4461_), .ZN(new_n18065_));
  AOI21_X1   g17873(.A1(new_n17770_), .A2(new_n18064_), .B(new_n18065_), .ZN(new_n18066_));
  AOI21_X1   g17874(.A1(new_n18066_), .A2(new_n4196_), .B(new_n17767_), .ZN(new_n18067_));
  NAND2_X1   g17875(.A1(new_n18064_), .A2(new_n17770_), .ZN(new_n18068_));
  INV_X1     g17876(.I(new_n17773_), .ZN(new_n18069_));
  INV_X1     g17877(.I(new_n17782_), .ZN(new_n18070_));
  NOR3_X1    g17878(.A1(new_n18055_), .A2(new_n18056_), .A3(\asqrt[32] ), .ZN(new_n18071_));
  OAI21_X1   g17879(.A1(new_n18070_), .A2(new_n18071_), .B(new_n18057_), .ZN(new_n18072_));
  OAI21_X1   g17880(.A1(new_n18072_), .A2(\asqrt[33] ), .B(new_n17778_), .ZN(new_n18073_));
  NAND2_X1   g17881(.A1(new_n18072_), .A2(\asqrt[33] ), .ZN(new_n18074_));
  NAND3_X1   g17882(.A1(new_n18073_), .A2(new_n18074_), .A3(new_n5029_), .ZN(new_n18075_));
  AOI21_X1   g17883(.A1(new_n18073_), .A2(new_n18074_), .B(new_n5029_), .ZN(new_n18076_));
  AOI21_X1   g17884(.A1(new_n17775_), .A2(new_n18075_), .B(new_n18076_), .ZN(new_n18077_));
  AOI21_X1   g17885(.A1(new_n18077_), .A2(new_n4751_), .B(new_n18069_), .ZN(new_n18078_));
  NOR2_X1    g17886(.A1(new_n18077_), .A2(new_n4751_), .ZN(new_n18079_));
  OAI21_X1   g17887(.A1(new_n18078_), .A2(new_n18079_), .B(\asqrt[36] ), .ZN(new_n18080_));
  AOI21_X1   g17888(.A1(new_n18068_), .A2(new_n18080_), .B(new_n4196_), .ZN(new_n18081_));
  NOR3_X1    g17889(.A1(new_n18067_), .A2(\asqrt[38] ), .A3(new_n18081_), .ZN(new_n18082_));
  OAI21_X1   g17890(.A1(new_n18067_), .A2(new_n18081_), .B(\asqrt[38] ), .ZN(new_n18083_));
  OAI21_X1   g17891(.A1(new_n17764_), .A2(new_n18082_), .B(new_n18083_), .ZN(new_n18084_));
  OAI21_X1   g17892(.A1(new_n18084_), .A2(\asqrt[39] ), .B(new_n17761_), .ZN(new_n18085_));
  NAND2_X1   g17893(.A1(new_n18084_), .A2(\asqrt[39] ), .ZN(new_n18086_));
  NAND3_X1   g17894(.A1(new_n18085_), .A2(new_n18086_), .A3(new_n3427_), .ZN(new_n18087_));
  AOI21_X1   g17895(.A1(new_n18085_), .A2(new_n18086_), .B(new_n3427_), .ZN(new_n18088_));
  AOI21_X1   g17896(.A1(new_n17758_), .A2(new_n18087_), .B(new_n18088_), .ZN(new_n18089_));
  AOI21_X1   g17897(.A1(new_n18089_), .A2(new_n3195_), .B(new_n17755_), .ZN(new_n18090_));
  NAND2_X1   g17898(.A1(new_n18087_), .A2(new_n17758_), .ZN(new_n18091_));
  INV_X1     g17899(.I(new_n17761_), .ZN(new_n18092_));
  INV_X1     g17900(.I(new_n17770_), .ZN(new_n18093_));
  NOR3_X1    g17901(.A1(new_n18078_), .A2(new_n18079_), .A3(\asqrt[36] ), .ZN(new_n18094_));
  OAI21_X1   g17902(.A1(new_n18093_), .A2(new_n18094_), .B(new_n18080_), .ZN(new_n18095_));
  OAI21_X1   g17903(.A1(new_n18095_), .A2(\asqrt[37] ), .B(new_n17766_), .ZN(new_n18096_));
  NAND2_X1   g17904(.A1(new_n18095_), .A2(\asqrt[37] ), .ZN(new_n18097_));
  NAND3_X1   g17905(.A1(new_n18096_), .A2(new_n18097_), .A3(new_n3925_), .ZN(new_n18098_));
  AOI21_X1   g17906(.A1(new_n18096_), .A2(new_n18097_), .B(new_n3925_), .ZN(new_n18099_));
  AOI21_X1   g17907(.A1(new_n17763_), .A2(new_n18098_), .B(new_n18099_), .ZN(new_n18100_));
  AOI21_X1   g17908(.A1(new_n18100_), .A2(new_n3681_), .B(new_n18092_), .ZN(new_n18101_));
  NOR2_X1    g17909(.A1(new_n18100_), .A2(new_n3681_), .ZN(new_n18102_));
  OAI21_X1   g17910(.A1(new_n18101_), .A2(new_n18102_), .B(\asqrt[40] ), .ZN(new_n18103_));
  AOI21_X1   g17911(.A1(new_n18091_), .A2(new_n18103_), .B(new_n3195_), .ZN(new_n18104_));
  NOR3_X1    g17912(.A1(new_n18090_), .A2(\asqrt[42] ), .A3(new_n18104_), .ZN(new_n18105_));
  OAI21_X1   g17913(.A1(new_n18090_), .A2(new_n18104_), .B(\asqrt[42] ), .ZN(new_n18106_));
  OAI21_X1   g17914(.A1(new_n17752_), .A2(new_n18105_), .B(new_n18106_), .ZN(new_n18107_));
  OAI21_X1   g17915(.A1(new_n18107_), .A2(\asqrt[43] ), .B(new_n17749_), .ZN(new_n18108_));
  NAND2_X1   g17916(.A1(new_n18107_), .A2(\asqrt[43] ), .ZN(new_n18109_));
  NAND3_X1   g17917(.A1(new_n18108_), .A2(new_n18109_), .A3(new_n2531_), .ZN(new_n18110_));
  AOI21_X1   g17918(.A1(new_n18108_), .A2(new_n18109_), .B(new_n2531_), .ZN(new_n18111_));
  AOI21_X1   g17919(.A1(new_n17746_), .A2(new_n18110_), .B(new_n18111_), .ZN(new_n18112_));
  AOI21_X1   g17920(.A1(new_n18112_), .A2(new_n2332_), .B(new_n17743_), .ZN(new_n18113_));
  NAND2_X1   g17921(.A1(new_n18110_), .A2(new_n17746_), .ZN(new_n18114_));
  INV_X1     g17922(.I(new_n17749_), .ZN(new_n18115_));
  INV_X1     g17923(.I(new_n17758_), .ZN(new_n18116_));
  NOR3_X1    g17924(.A1(new_n18101_), .A2(new_n18102_), .A3(\asqrt[40] ), .ZN(new_n18117_));
  OAI21_X1   g17925(.A1(new_n18116_), .A2(new_n18117_), .B(new_n18103_), .ZN(new_n18118_));
  OAI21_X1   g17926(.A1(new_n18118_), .A2(\asqrt[41] ), .B(new_n17754_), .ZN(new_n18119_));
  NAND2_X1   g17927(.A1(new_n18118_), .A2(\asqrt[41] ), .ZN(new_n18120_));
  NAND3_X1   g17928(.A1(new_n18119_), .A2(new_n18120_), .A3(new_n2960_), .ZN(new_n18121_));
  AOI21_X1   g17929(.A1(new_n18119_), .A2(new_n18120_), .B(new_n2960_), .ZN(new_n18122_));
  AOI21_X1   g17930(.A1(new_n17751_), .A2(new_n18121_), .B(new_n18122_), .ZN(new_n18123_));
  AOI21_X1   g17931(.A1(new_n18123_), .A2(new_n2749_), .B(new_n18115_), .ZN(new_n18124_));
  NOR2_X1    g17932(.A1(new_n18123_), .A2(new_n2749_), .ZN(new_n18125_));
  OAI21_X1   g17933(.A1(new_n18124_), .A2(new_n18125_), .B(\asqrt[44] ), .ZN(new_n18126_));
  AOI21_X1   g17934(.A1(new_n18114_), .A2(new_n18126_), .B(new_n2332_), .ZN(new_n18127_));
  NOR3_X1    g17935(.A1(new_n18113_), .A2(\asqrt[46] ), .A3(new_n18127_), .ZN(new_n18128_));
  OAI21_X1   g17936(.A1(new_n18113_), .A2(new_n18127_), .B(\asqrt[46] ), .ZN(new_n18129_));
  OAI21_X1   g17937(.A1(new_n17740_), .A2(new_n18128_), .B(new_n18129_), .ZN(new_n18130_));
  OAI21_X1   g17938(.A1(new_n18130_), .A2(\asqrt[47] ), .B(new_n17737_), .ZN(new_n18131_));
  NAND2_X1   g17939(.A1(new_n18130_), .A2(\asqrt[47] ), .ZN(new_n18132_));
  NAND3_X1   g17940(.A1(new_n18131_), .A2(new_n18132_), .A3(new_n1778_), .ZN(new_n18133_));
  AOI21_X1   g17941(.A1(new_n18131_), .A2(new_n18132_), .B(new_n1778_), .ZN(new_n18134_));
  AOI21_X1   g17942(.A1(new_n17734_), .A2(new_n18133_), .B(new_n18134_), .ZN(new_n18135_));
  AOI21_X1   g17943(.A1(new_n18135_), .A2(new_n1632_), .B(new_n17731_), .ZN(new_n18136_));
  NAND2_X1   g17944(.A1(new_n18133_), .A2(new_n17734_), .ZN(new_n18137_));
  INV_X1     g17945(.I(new_n17737_), .ZN(new_n18138_));
  INV_X1     g17946(.I(new_n17746_), .ZN(new_n18139_));
  NOR3_X1    g17947(.A1(new_n18124_), .A2(new_n18125_), .A3(\asqrt[44] ), .ZN(new_n18140_));
  OAI21_X1   g17948(.A1(new_n18139_), .A2(new_n18140_), .B(new_n18126_), .ZN(new_n18141_));
  OAI21_X1   g17949(.A1(new_n18141_), .A2(\asqrt[45] ), .B(new_n17742_), .ZN(new_n18142_));
  NAND2_X1   g17950(.A1(new_n18141_), .A2(\asqrt[45] ), .ZN(new_n18143_));
  NAND3_X1   g17951(.A1(new_n18142_), .A2(new_n18143_), .A3(new_n2134_), .ZN(new_n18144_));
  AOI21_X1   g17952(.A1(new_n18142_), .A2(new_n18143_), .B(new_n2134_), .ZN(new_n18145_));
  AOI21_X1   g17953(.A1(new_n17739_), .A2(new_n18144_), .B(new_n18145_), .ZN(new_n18146_));
  AOI21_X1   g17954(.A1(new_n18146_), .A2(new_n1953_), .B(new_n18138_), .ZN(new_n18147_));
  NOR2_X1    g17955(.A1(new_n18146_), .A2(new_n1953_), .ZN(new_n18148_));
  OAI21_X1   g17956(.A1(new_n18147_), .A2(new_n18148_), .B(\asqrt[48] ), .ZN(new_n18149_));
  AOI21_X1   g17957(.A1(new_n18137_), .A2(new_n18149_), .B(new_n1632_), .ZN(new_n18150_));
  NOR3_X1    g17958(.A1(new_n18136_), .A2(\asqrt[50] ), .A3(new_n18150_), .ZN(new_n18151_));
  OAI21_X1   g17959(.A1(new_n18136_), .A2(new_n18150_), .B(\asqrt[50] ), .ZN(new_n18152_));
  OAI21_X1   g17960(.A1(new_n17728_), .A2(new_n18151_), .B(new_n18152_), .ZN(new_n18153_));
  OAI21_X1   g17961(.A1(new_n18153_), .A2(\asqrt[51] ), .B(new_n17725_), .ZN(new_n18154_));
  NAND2_X1   g17962(.A1(new_n18153_), .A2(\asqrt[51] ), .ZN(new_n18155_));
  NAND3_X1   g17963(.A1(new_n18154_), .A2(new_n18155_), .A3(new_n1150_), .ZN(new_n18156_));
  AOI21_X1   g17964(.A1(new_n18154_), .A2(new_n18155_), .B(new_n1150_), .ZN(new_n18157_));
  AOI21_X1   g17965(.A1(new_n17722_), .A2(new_n18156_), .B(new_n18157_), .ZN(new_n18158_));
  AOI21_X1   g17966(.A1(new_n18158_), .A2(new_n1006_), .B(new_n17719_), .ZN(new_n18159_));
  NAND2_X1   g17967(.A1(new_n18156_), .A2(new_n17722_), .ZN(new_n18160_));
  INV_X1     g17968(.I(new_n17725_), .ZN(new_n18161_));
  INV_X1     g17969(.I(new_n17734_), .ZN(new_n18162_));
  NOR3_X1    g17970(.A1(new_n18147_), .A2(new_n18148_), .A3(\asqrt[48] ), .ZN(new_n18163_));
  OAI21_X1   g17971(.A1(new_n18162_), .A2(new_n18163_), .B(new_n18149_), .ZN(new_n18164_));
  OAI21_X1   g17972(.A1(new_n18164_), .A2(\asqrt[49] ), .B(new_n17730_), .ZN(new_n18165_));
  NAND2_X1   g17973(.A1(new_n18164_), .A2(\asqrt[49] ), .ZN(new_n18166_));
  NAND3_X1   g17974(.A1(new_n18165_), .A2(new_n18166_), .A3(new_n1463_), .ZN(new_n18167_));
  AOI21_X1   g17975(.A1(new_n18165_), .A2(new_n18166_), .B(new_n1463_), .ZN(new_n18168_));
  AOI21_X1   g17976(.A1(new_n17727_), .A2(new_n18167_), .B(new_n18168_), .ZN(new_n18169_));
  AOI21_X1   g17977(.A1(new_n18169_), .A2(new_n1305_), .B(new_n18161_), .ZN(new_n18170_));
  NOR2_X1    g17978(.A1(new_n18169_), .A2(new_n1305_), .ZN(new_n18171_));
  OAI21_X1   g17979(.A1(new_n18170_), .A2(new_n18171_), .B(\asqrt[52] ), .ZN(new_n18172_));
  AOI21_X1   g17980(.A1(new_n18160_), .A2(new_n18172_), .B(new_n1006_), .ZN(new_n18173_));
  NOR3_X1    g17981(.A1(new_n18159_), .A2(\asqrt[54] ), .A3(new_n18173_), .ZN(new_n18174_));
  OAI21_X1   g17982(.A1(new_n18159_), .A2(new_n18173_), .B(\asqrt[54] ), .ZN(new_n18175_));
  OAI21_X1   g17983(.A1(new_n17716_), .A2(new_n18174_), .B(new_n18175_), .ZN(new_n18176_));
  OAI21_X1   g17984(.A1(new_n18176_), .A2(\asqrt[55] ), .B(new_n17713_), .ZN(new_n18177_));
  NAND2_X1   g17985(.A1(new_n18176_), .A2(\asqrt[55] ), .ZN(new_n18178_));
  NAND3_X1   g17986(.A1(new_n18177_), .A2(new_n18178_), .A3(new_n634_), .ZN(new_n18179_));
  AOI21_X1   g17987(.A1(new_n18177_), .A2(new_n18178_), .B(new_n634_), .ZN(new_n18180_));
  AOI21_X1   g17988(.A1(new_n17710_), .A2(new_n18179_), .B(new_n18180_), .ZN(new_n18181_));
  AOI21_X1   g17989(.A1(new_n18181_), .A2(new_n531_), .B(new_n17706_), .ZN(new_n18182_));
  NAND2_X1   g17990(.A1(new_n18179_), .A2(new_n17710_), .ZN(new_n18183_));
  INV_X1     g17991(.I(new_n17713_), .ZN(new_n18184_));
  INV_X1     g17992(.I(new_n17722_), .ZN(new_n18185_));
  NOR3_X1    g17993(.A1(new_n18170_), .A2(new_n18171_), .A3(\asqrt[52] ), .ZN(new_n18186_));
  OAI21_X1   g17994(.A1(new_n18185_), .A2(new_n18186_), .B(new_n18172_), .ZN(new_n18187_));
  OAI21_X1   g17995(.A1(new_n18187_), .A2(\asqrt[53] ), .B(new_n17718_), .ZN(new_n18188_));
  NAND2_X1   g17996(.A1(new_n18187_), .A2(\asqrt[53] ), .ZN(new_n18189_));
  NAND3_X1   g17997(.A1(new_n18188_), .A2(new_n18189_), .A3(new_n860_), .ZN(new_n18190_));
  AOI21_X1   g17998(.A1(new_n18188_), .A2(new_n18189_), .B(new_n860_), .ZN(new_n18191_));
  AOI21_X1   g17999(.A1(new_n17715_), .A2(new_n18190_), .B(new_n18191_), .ZN(new_n18192_));
  AOI21_X1   g18000(.A1(new_n18192_), .A2(new_n744_), .B(new_n18184_), .ZN(new_n18193_));
  NOR2_X1    g18001(.A1(new_n18192_), .A2(new_n744_), .ZN(new_n18194_));
  OAI21_X1   g18002(.A1(new_n18193_), .A2(new_n18194_), .B(\asqrt[56] ), .ZN(new_n18195_));
  AOI21_X1   g18003(.A1(new_n18183_), .A2(new_n18195_), .B(new_n531_), .ZN(new_n18196_));
  NOR3_X1    g18004(.A1(new_n18182_), .A2(\asqrt[58] ), .A3(new_n18196_), .ZN(new_n18197_));
  OAI21_X1   g18005(.A1(new_n18182_), .A2(new_n18196_), .B(\asqrt[58] ), .ZN(new_n18198_));
  OAI21_X1   g18006(.A1(new_n17703_), .A2(new_n18197_), .B(new_n18198_), .ZN(new_n18199_));
  OAI21_X1   g18007(.A1(new_n18199_), .A2(\asqrt[59] ), .B(new_n17700_), .ZN(new_n18200_));
  NAND2_X1   g18008(.A1(new_n18199_), .A2(\asqrt[59] ), .ZN(new_n18201_));
  NAND3_X1   g18009(.A1(new_n18200_), .A2(new_n18201_), .A3(new_n266_), .ZN(new_n18202_));
  NAND2_X1   g18010(.A1(new_n18202_), .A2(new_n17697_), .ZN(new_n18203_));
  INV_X1     g18011(.I(new_n17700_), .ZN(new_n18204_));
  INV_X1     g18012(.I(new_n17710_), .ZN(new_n18205_));
  NOR3_X1    g18013(.A1(new_n18193_), .A2(new_n18194_), .A3(\asqrt[56] ), .ZN(new_n18206_));
  OAI21_X1   g18014(.A1(new_n18205_), .A2(new_n18206_), .B(new_n18195_), .ZN(new_n18207_));
  OAI21_X1   g18015(.A1(new_n18207_), .A2(\asqrt[57] ), .B(new_n17705_), .ZN(new_n18208_));
  NOR2_X1    g18016(.A1(new_n18206_), .A2(new_n18205_), .ZN(new_n18209_));
  OAI21_X1   g18017(.A1(new_n18209_), .A2(new_n18180_), .B(\asqrt[57] ), .ZN(new_n18210_));
  NAND3_X1   g18018(.A1(new_n18208_), .A2(new_n423_), .A3(new_n18210_), .ZN(new_n18211_));
  AOI21_X1   g18019(.A1(new_n18208_), .A2(new_n18210_), .B(new_n423_), .ZN(new_n18212_));
  AOI21_X1   g18020(.A1(new_n17702_), .A2(new_n18211_), .B(new_n18212_), .ZN(new_n18213_));
  AOI21_X1   g18021(.A1(new_n18213_), .A2(new_n337_), .B(new_n18204_), .ZN(new_n18214_));
  NAND2_X1   g18022(.A1(new_n18211_), .A2(new_n17702_), .ZN(new_n18215_));
  AOI21_X1   g18023(.A1(new_n18215_), .A2(new_n18198_), .B(new_n337_), .ZN(new_n18216_));
  OAI21_X1   g18024(.A1(new_n18214_), .A2(new_n18216_), .B(\asqrt[60] ), .ZN(new_n18217_));
  AOI21_X1   g18025(.A1(new_n18203_), .A2(new_n18217_), .B(new_n239_), .ZN(new_n18218_));
  INV_X1     g18026(.I(new_n17697_), .ZN(new_n18219_));
  NAND3_X1   g18027(.A1(new_n18215_), .A2(new_n337_), .A3(new_n18198_), .ZN(new_n18220_));
  AOI21_X1   g18028(.A1(new_n17700_), .A2(new_n18220_), .B(new_n18216_), .ZN(new_n18221_));
  AOI21_X1   g18029(.A1(new_n18221_), .A2(new_n266_), .B(new_n18219_), .ZN(new_n18222_));
  AOI21_X1   g18030(.A1(new_n18200_), .A2(new_n18201_), .B(new_n266_), .ZN(new_n18223_));
  NOR3_X1    g18031(.A1(new_n18222_), .A2(\asqrt[61] ), .A3(new_n18223_), .ZN(new_n18224_));
  AOI21_X1   g18032(.A1(new_n17864_), .A2(new_n17689_), .B(\asqrt[4] ), .ZN(new_n18225_));
  XOR2_X1    g18033(.A1(new_n18225_), .A2(new_n17681_), .Z(new_n18226_));
  AOI21_X1   g18034(.A1(new_n17697_), .A2(new_n18202_), .B(new_n18223_), .ZN(new_n18227_));
  AOI21_X1   g18035(.A1(new_n18227_), .A2(new_n239_), .B(new_n17694_), .ZN(new_n18228_));
  NOR2_X1    g18036(.A1(new_n18228_), .A2(new_n18218_), .ZN(new_n18229_));
  OAI21_X1   g18037(.A1(new_n18222_), .A2(new_n18223_), .B(\asqrt[61] ), .ZN(new_n18230_));
  NOR3_X1    g18038(.A1(new_n18214_), .A2(\asqrt[60] ), .A3(new_n18216_), .ZN(new_n18231_));
  OAI21_X1   g18039(.A1(new_n18219_), .A2(new_n18231_), .B(new_n18217_), .ZN(new_n18232_));
  OAI21_X1   g18040(.A1(new_n18232_), .A2(\asqrt[61] ), .B(new_n17693_), .ZN(new_n18233_));
  AOI21_X1   g18041(.A1(new_n18233_), .A2(new_n18230_), .B(\asqrt[62] ), .ZN(new_n18234_));
  NOR3_X1    g18042(.A1(new_n18228_), .A2(new_n201_), .A3(new_n18218_), .ZN(new_n18235_));
  AOI21_X1   g18043(.A1(new_n17666_), .A2(new_n17671_), .B(\asqrt[4] ), .ZN(new_n18236_));
  XOR2_X1    g18044(.A1(new_n18236_), .A2(new_n17668_), .Z(new_n18237_));
  OAI22_X1   g18045(.A1(new_n18234_), .A2(new_n18235_), .B1(new_n18229_), .B2(new_n18237_), .ZN(new_n18238_));
  NOR2_X1    g18046(.A1(new_n17683_), .A2(new_n17661_), .ZN(new_n18239_));
  OAI21_X1   g18047(.A1(\asqrt[4] ), .A2(new_n18239_), .B(new_n17690_), .ZN(new_n18240_));
  AOI21_X1   g18048(.A1(new_n18238_), .A2(new_n18226_), .B(new_n18240_), .ZN(new_n18241_));
  NOR2_X1    g18049(.A1(\asqrt[4] ), .A2(new_n17661_), .ZN(new_n18242_));
  NOR2_X1    g18050(.A1(new_n17862_), .A2(new_n17661_), .ZN(new_n18243_));
  NOR2_X1    g18051(.A1(new_n17683_), .A2(new_n17660_), .ZN(new_n18244_));
  OAI21_X1   g18052(.A1(new_n18243_), .A2(new_n18244_), .B(\asqrt[63] ), .ZN(new_n18245_));
  NOR2_X1    g18053(.A1(new_n18242_), .A2(new_n18245_), .ZN(new_n18246_));
  INV_X1     g18054(.I(new_n18246_), .ZN(new_n18247_));
  INV_X1     g18055(.I(new_n18237_), .ZN(new_n18248_));
  AOI21_X1   g18056(.A1(new_n18229_), .A2(new_n201_), .B(new_n18248_), .ZN(new_n18249_));
  INV_X1     g18057(.I(new_n18226_), .ZN(new_n18250_));
  OAI21_X1   g18058(.A1(new_n18229_), .A2(new_n201_), .B(new_n18250_), .ZN(new_n18251_));
  OAI21_X1   g18059(.A1(new_n18249_), .A2(new_n18251_), .B(new_n18247_), .ZN(new_n18252_));
  NOR3_X1    g18060(.A1(new_n18241_), .A2(\asqrt[63] ), .A3(new_n18252_), .ZN(new_n18253_));
  OAI21_X1   g18061(.A1(new_n18218_), .A2(new_n18224_), .B(new_n18253_), .ZN(new_n18254_));
  XOR2_X1    g18062(.A1(new_n18254_), .A2(new_n17694_), .Z(new_n18255_));
  INV_X1     g18063(.I(new_n18255_), .ZN(new_n18256_));
  XOR2_X1    g18064(.A1(new_n18229_), .A2(\asqrt[62] ), .Z(new_n18257_));
  NAND2_X1   g18065(.A1(new_n18253_), .A2(new_n18257_), .ZN(new_n18258_));
  XOR2_X1    g18066(.A1(new_n18258_), .A2(new_n18248_), .Z(new_n18259_));
  NAND2_X1   g18067(.A1(new_n18201_), .A2(new_n18220_), .ZN(new_n18260_));
  NAND2_X1   g18068(.A1(new_n18253_), .A2(new_n18260_), .ZN(new_n18261_));
  XOR2_X1    g18069(.A1(new_n18261_), .A2(new_n18204_), .Z(new_n18262_));
  OAI21_X1   g18070(.A1(new_n18197_), .A2(new_n18212_), .B(new_n18253_), .ZN(new_n18263_));
  XOR2_X1    g18071(.A1(new_n18263_), .A2(new_n17703_), .Z(new_n18264_));
  NOR2_X1    g18072(.A1(new_n18207_), .A2(\asqrt[57] ), .ZN(new_n18265_));
  OAI21_X1   g18073(.A1(new_n18265_), .A2(new_n18196_), .B(new_n18253_), .ZN(new_n18266_));
  XOR2_X1    g18074(.A1(new_n18266_), .A2(new_n17706_), .Z(new_n18267_));
  OAI21_X1   g18075(.A1(new_n18206_), .A2(new_n18180_), .B(new_n18253_), .ZN(new_n18268_));
  XOR2_X1    g18076(.A1(new_n18268_), .A2(new_n18205_), .Z(new_n18269_));
  INV_X1     g18077(.I(new_n18269_), .ZN(new_n18270_));
  NAND2_X1   g18078(.A1(new_n18192_), .A2(new_n744_), .ZN(new_n18271_));
  NAND2_X1   g18079(.A1(new_n18271_), .A2(new_n18178_), .ZN(new_n18272_));
  NAND2_X1   g18080(.A1(new_n18253_), .A2(new_n18272_), .ZN(new_n18273_));
  XOR2_X1    g18081(.A1(new_n18273_), .A2(new_n18184_), .Z(new_n18274_));
  INV_X1     g18082(.I(new_n18274_), .ZN(new_n18275_));
  OAI21_X1   g18083(.A1(new_n18174_), .A2(new_n18191_), .B(new_n18253_), .ZN(new_n18276_));
  XOR2_X1    g18084(.A1(new_n18276_), .A2(new_n17716_), .Z(new_n18277_));
  NOR2_X1    g18085(.A1(new_n18187_), .A2(\asqrt[53] ), .ZN(new_n18278_));
  OAI21_X1   g18086(.A1(new_n18278_), .A2(new_n18173_), .B(new_n18253_), .ZN(new_n18279_));
  XOR2_X1    g18087(.A1(new_n18279_), .A2(new_n17719_), .Z(new_n18280_));
  OAI21_X1   g18088(.A1(new_n18186_), .A2(new_n18157_), .B(new_n18253_), .ZN(new_n18281_));
  XOR2_X1    g18089(.A1(new_n18281_), .A2(new_n18185_), .Z(new_n18282_));
  INV_X1     g18090(.I(new_n18282_), .ZN(new_n18283_));
  NAND2_X1   g18091(.A1(new_n18169_), .A2(new_n1305_), .ZN(new_n18284_));
  NAND2_X1   g18092(.A1(new_n18284_), .A2(new_n18155_), .ZN(new_n18285_));
  NAND2_X1   g18093(.A1(new_n18253_), .A2(new_n18285_), .ZN(new_n18286_));
  XOR2_X1    g18094(.A1(new_n18286_), .A2(new_n18161_), .Z(new_n18287_));
  INV_X1     g18095(.I(new_n18287_), .ZN(new_n18288_));
  OAI21_X1   g18096(.A1(new_n18151_), .A2(new_n18168_), .B(new_n18253_), .ZN(new_n18289_));
  XOR2_X1    g18097(.A1(new_n18289_), .A2(new_n17728_), .Z(new_n18290_));
  NOR2_X1    g18098(.A1(new_n18164_), .A2(\asqrt[49] ), .ZN(new_n18291_));
  OAI21_X1   g18099(.A1(new_n18291_), .A2(new_n18150_), .B(new_n18253_), .ZN(new_n18292_));
  XOR2_X1    g18100(.A1(new_n18292_), .A2(new_n17731_), .Z(new_n18293_));
  OAI21_X1   g18101(.A1(new_n18163_), .A2(new_n18134_), .B(new_n18253_), .ZN(new_n18294_));
  XOR2_X1    g18102(.A1(new_n18294_), .A2(new_n18162_), .Z(new_n18295_));
  INV_X1     g18103(.I(new_n18295_), .ZN(new_n18296_));
  NAND2_X1   g18104(.A1(new_n18146_), .A2(new_n1953_), .ZN(new_n18297_));
  OAI21_X1   g18105(.A1(new_n17694_), .A2(new_n18224_), .B(new_n18230_), .ZN(new_n18298_));
  OAI21_X1   g18106(.A1(new_n18228_), .A2(new_n18218_), .B(new_n201_), .ZN(new_n18299_));
  NAND3_X1   g18107(.A1(new_n18233_), .A2(\asqrt[62] ), .A3(new_n18230_), .ZN(new_n18300_));
  AOI22_X1   g18108(.A1(new_n18300_), .A2(new_n18299_), .B1(new_n18298_), .B2(new_n18248_), .ZN(new_n18301_));
  INV_X1     g18109(.I(new_n18240_), .ZN(new_n18302_));
  OAI21_X1   g18110(.A1(new_n18301_), .A2(new_n18250_), .B(new_n18302_), .ZN(new_n18303_));
  OAI21_X1   g18111(.A1(new_n18298_), .A2(\asqrt[62] ), .B(new_n18237_), .ZN(new_n18304_));
  AOI21_X1   g18112(.A1(new_n18298_), .A2(\asqrt[62] ), .B(new_n18226_), .ZN(new_n18305_));
  AOI21_X1   g18113(.A1(new_n18305_), .A2(new_n18304_), .B(new_n18246_), .ZN(new_n18306_));
  NAND3_X1   g18114(.A1(new_n18303_), .A2(new_n193_), .A3(new_n18306_), .ZN(\asqrt[3] ));
  AOI21_X1   g18115(.A1(new_n18297_), .A2(new_n18132_), .B(\asqrt[3] ), .ZN(new_n18308_));
  XOR2_X1    g18116(.A1(new_n18308_), .A2(new_n17737_), .Z(new_n18309_));
  INV_X1     g18117(.I(new_n18309_), .ZN(new_n18310_));
  OAI21_X1   g18118(.A1(new_n18128_), .A2(new_n18145_), .B(new_n18253_), .ZN(new_n18311_));
  XOR2_X1    g18119(.A1(new_n18311_), .A2(new_n17740_), .Z(new_n18312_));
  NOR2_X1    g18120(.A1(new_n18141_), .A2(\asqrt[45] ), .ZN(new_n18313_));
  OAI21_X1   g18121(.A1(new_n18313_), .A2(new_n18127_), .B(new_n18253_), .ZN(new_n18314_));
  XOR2_X1    g18122(.A1(new_n18314_), .A2(new_n17743_), .Z(new_n18315_));
  OAI21_X1   g18123(.A1(new_n18140_), .A2(new_n18111_), .B(new_n18253_), .ZN(new_n18316_));
  XOR2_X1    g18124(.A1(new_n18316_), .A2(new_n18139_), .Z(new_n18317_));
  INV_X1     g18125(.I(new_n18317_), .ZN(new_n18318_));
  NAND2_X1   g18126(.A1(new_n18123_), .A2(new_n2749_), .ZN(new_n18319_));
  AOI21_X1   g18127(.A1(new_n18319_), .A2(new_n18109_), .B(\asqrt[3] ), .ZN(new_n18320_));
  XOR2_X1    g18128(.A1(new_n18320_), .A2(new_n17749_), .Z(new_n18321_));
  INV_X1     g18129(.I(new_n18321_), .ZN(new_n18322_));
  OAI21_X1   g18130(.A1(new_n18105_), .A2(new_n18122_), .B(new_n18253_), .ZN(new_n18323_));
  XOR2_X1    g18131(.A1(new_n18323_), .A2(new_n17752_), .Z(new_n18324_));
  NOR2_X1    g18132(.A1(new_n18118_), .A2(\asqrt[41] ), .ZN(new_n18325_));
  OAI21_X1   g18133(.A1(new_n18325_), .A2(new_n18104_), .B(new_n18253_), .ZN(new_n18326_));
  XOR2_X1    g18134(.A1(new_n18326_), .A2(new_n17755_), .Z(new_n18327_));
  OAI21_X1   g18135(.A1(new_n18117_), .A2(new_n18088_), .B(new_n18253_), .ZN(new_n18328_));
  XOR2_X1    g18136(.A1(new_n18328_), .A2(new_n18116_), .Z(new_n18329_));
  INV_X1     g18137(.I(new_n18329_), .ZN(new_n18330_));
  NAND2_X1   g18138(.A1(new_n18100_), .A2(new_n3681_), .ZN(new_n18331_));
  AOI21_X1   g18139(.A1(new_n18331_), .A2(new_n18086_), .B(\asqrt[3] ), .ZN(new_n18332_));
  XOR2_X1    g18140(.A1(new_n18332_), .A2(new_n17761_), .Z(new_n18333_));
  INV_X1     g18141(.I(new_n18333_), .ZN(new_n18334_));
  OAI21_X1   g18142(.A1(new_n18082_), .A2(new_n18099_), .B(new_n18253_), .ZN(new_n18335_));
  XOR2_X1    g18143(.A1(new_n18335_), .A2(new_n17764_), .Z(new_n18336_));
  NOR2_X1    g18144(.A1(new_n18095_), .A2(\asqrt[37] ), .ZN(new_n18337_));
  OAI21_X1   g18145(.A1(new_n18337_), .A2(new_n18081_), .B(new_n18253_), .ZN(new_n18338_));
  XOR2_X1    g18146(.A1(new_n18338_), .A2(new_n17767_), .Z(new_n18339_));
  OAI21_X1   g18147(.A1(new_n18094_), .A2(new_n18065_), .B(new_n18253_), .ZN(new_n18340_));
  XOR2_X1    g18148(.A1(new_n18340_), .A2(new_n18093_), .Z(new_n18341_));
  INV_X1     g18149(.I(new_n18341_), .ZN(new_n18342_));
  NAND2_X1   g18150(.A1(new_n18077_), .A2(new_n4751_), .ZN(new_n18343_));
  AOI21_X1   g18151(.A1(new_n18343_), .A2(new_n18063_), .B(\asqrt[3] ), .ZN(new_n18344_));
  XOR2_X1    g18152(.A1(new_n18344_), .A2(new_n17773_), .Z(new_n18345_));
  INV_X1     g18153(.I(new_n18345_), .ZN(new_n18346_));
  OAI21_X1   g18154(.A1(new_n18059_), .A2(new_n18076_), .B(new_n18253_), .ZN(new_n18347_));
  XOR2_X1    g18155(.A1(new_n18347_), .A2(new_n17776_), .Z(new_n18348_));
  NOR2_X1    g18156(.A1(new_n18072_), .A2(\asqrt[33] ), .ZN(new_n18349_));
  OAI21_X1   g18157(.A1(new_n18349_), .A2(new_n18058_), .B(new_n18253_), .ZN(new_n18350_));
  XOR2_X1    g18158(.A1(new_n18350_), .A2(new_n17779_), .Z(new_n18351_));
  OAI21_X1   g18159(.A1(new_n18071_), .A2(new_n18042_), .B(new_n18253_), .ZN(new_n18352_));
  XOR2_X1    g18160(.A1(new_n18352_), .A2(new_n18070_), .Z(new_n18353_));
  INV_X1     g18161(.I(new_n18353_), .ZN(new_n18354_));
  NAND2_X1   g18162(.A1(new_n18054_), .A2(new_n5947_), .ZN(new_n18355_));
  AOI21_X1   g18163(.A1(new_n18355_), .A2(new_n18040_), .B(\asqrt[3] ), .ZN(new_n18356_));
  XOR2_X1    g18164(.A1(new_n18356_), .A2(new_n17785_), .Z(new_n18357_));
  INV_X1     g18165(.I(new_n18357_), .ZN(new_n18358_));
  OAI21_X1   g18166(.A1(new_n18036_), .A2(new_n18053_), .B(new_n18253_), .ZN(new_n18359_));
  XOR2_X1    g18167(.A1(new_n18359_), .A2(new_n17788_), .Z(new_n18360_));
  NOR2_X1    g18168(.A1(new_n18049_), .A2(\asqrt[29] ), .ZN(new_n18361_));
  OAI21_X1   g18169(.A1(new_n18361_), .A2(new_n18035_), .B(new_n18253_), .ZN(new_n18362_));
  XOR2_X1    g18170(.A1(new_n18362_), .A2(new_n17791_), .Z(new_n18363_));
  OAI21_X1   g18171(.A1(new_n18048_), .A2(new_n18019_), .B(new_n18253_), .ZN(new_n18364_));
  XOR2_X1    g18172(.A1(new_n18364_), .A2(new_n18047_), .Z(new_n18365_));
  INV_X1     g18173(.I(new_n18365_), .ZN(new_n18366_));
  NAND2_X1   g18174(.A1(new_n18031_), .A2(new_n7331_), .ZN(new_n18367_));
  AOI21_X1   g18175(.A1(new_n18367_), .A2(new_n18017_), .B(\asqrt[3] ), .ZN(new_n18368_));
  XOR2_X1    g18176(.A1(new_n18368_), .A2(new_n17797_), .Z(new_n18369_));
  INV_X1     g18177(.I(new_n18369_), .ZN(new_n18370_));
  OAI21_X1   g18178(.A1(new_n18013_), .A2(new_n18030_), .B(new_n18253_), .ZN(new_n18371_));
  XOR2_X1    g18179(.A1(new_n18371_), .A2(new_n17800_), .Z(new_n18372_));
  NOR2_X1    g18180(.A1(new_n18026_), .A2(\asqrt[25] ), .ZN(new_n18373_));
  OAI21_X1   g18181(.A1(new_n18373_), .A2(new_n18012_), .B(new_n18253_), .ZN(new_n18374_));
  XOR2_X1    g18182(.A1(new_n18374_), .A2(new_n17803_), .Z(new_n18375_));
  OAI21_X1   g18183(.A1(new_n18025_), .A2(new_n17996_), .B(new_n18253_), .ZN(new_n18376_));
  XOR2_X1    g18184(.A1(new_n18376_), .A2(new_n18024_), .Z(new_n18377_));
  INV_X1     g18185(.I(new_n18377_), .ZN(new_n18378_));
  NAND2_X1   g18186(.A1(new_n18008_), .A2(new_n8849_), .ZN(new_n18379_));
  AOI21_X1   g18187(.A1(new_n18379_), .A2(new_n17994_), .B(\asqrt[3] ), .ZN(new_n18380_));
  XOR2_X1    g18188(.A1(new_n18380_), .A2(new_n17809_), .Z(new_n18381_));
  INV_X1     g18189(.I(new_n18381_), .ZN(new_n18382_));
  OAI21_X1   g18190(.A1(new_n17990_), .A2(new_n18007_), .B(new_n18253_), .ZN(new_n18383_));
  XOR2_X1    g18191(.A1(new_n18383_), .A2(new_n17812_), .Z(new_n18384_));
  NOR2_X1    g18192(.A1(new_n18003_), .A2(\asqrt[21] ), .ZN(new_n18385_));
  OAI21_X1   g18193(.A1(new_n18385_), .A2(new_n17989_), .B(new_n18253_), .ZN(new_n18386_));
  XOR2_X1    g18194(.A1(new_n18386_), .A2(new_n17815_), .Z(new_n18387_));
  OAI21_X1   g18195(.A1(new_n18002_), .A2(new_n17973_), .B(new_n18253_), .ZN(new_n18388_));
  XOR2_X1    g18196(.A1(new_n18388_), .A2(new_n18001_), .Z(new_n18389_));
  INV_X1     g18197(.I(new_n18389_), .ZN(new_n18390_));
  NAND2_X1   g18198(.A1(new_n17985_), .A2(new_n10497_), .ZN(new_n18391_));
  AOI21_X1   g18199(.A1(new_n18391_), .A2(new_n17971_), .B(\asqrt[3] ), .ZN(new_n18392_));
  XOR2_X1    g18200(.A1(new_n18392_), .A2(new_n17821_), .Z(new_n18393_));
  INV_X1     g18201(.I(new_n18393_), .ZN(new_n18394_));
  OAI21_X1   g18202(.A1(new_n17967_), .A2(new_n17984_), .B(new_n18253_), .ZN(new_n18395_));
  XOR2_X1    g18203(.A1(new_n18395_), .A2(new_n17824_), .Z(new_n18396_));
  NOR2_X1    g18204(.A1(new_n17980_), .A2(\asqrt[17] ), .ZN(new_n18397_));
  OAI21_X1   g18205(.A1(new_n18397_), .A2(new_n17966_), .B(new_n18253_), .ZN(new_n18398_));
  XOR2_X1    g18206(.A1(new_n18398_), .A2(new_n17827_), .Z(new_n18399_));
  OAI21_X1   g18207(.A1(new_n17979_), .A2(new_n17950_), .B(new_n18253_), .ZN(new_n18400_));
  XOR2_X1    g18208(.A1(new_n18400_), .A2(new_n17978_), .Z(new_n18401_));
  INV_X1     g18209(.I(new_n18401_), .ZN(new_n18402_));
  NAND2_X1   g18210(.A1(new_n17962_), .A2(new_n12283_), .ZN(new_n18403_));
  AOI21_X1   g18211(.A1(new_n18403_), .A2(new_n17948_), .B(\asqrt[3] ), .ZN(new_n18404_));
  XOR2_X1    g18212(.A1(new_n18404_), .A2(new_n17833_), .Z(new_n18405_));
  INV_X1     g18213(.I(new_n18405_), .ZN(new_n18406_));
  OAI21_X1   g18214(.A1(new_n17944_), .A2(new_n17961_), .B(new_n18253_), .ZN(new_n18407_));
  XOR2_X1    g18215(.A1(new_n18407_), .A2(new_n17836_), .Z(new_n18408_));
  NOR2_X1    g18216(.A1(new_n17957_), .A2(\asqrt[13] ), .ZN(new_n18409_));
  OAI21_X1   g18217(.A1(new_n18409_), .A2(new_n17943_), .B(new_n18253_), .ZN(new_n18410_));
  XOR2_X1    g18218(.A1(new_n18410_), .A2(new_n17839_), .Z(new_n18411_));
  OAI21_X1   g18219(.A1(new_n17956_), .A2(new_n17927_), .B(new_n18253_), .ZN(new_n18412_));
  XOR2_X1    g18220(.A1(new_n18412_), .A2(new_n17955_), .Z(new_n18413_));
  INV_X1     g18221(.I(new_n18413_), .ZN(new_n18414_));
  NAND2_X1   g18222(.A1(new_n17939_), .A2(new_n14207_), .ZN(new_n18415_));
  AOI21_X1   g18223(.A1(new_n18415_), .A2(new_n17925_), .B(\asqrt[3] ), .ZN(new_n18416_));
  XOR2_X1    g18224(.A1(new_n18416_), .A2(new_n17845_), .Z(new_n18417_));
  INV_X1     g18225(.I(new_n18417_), .ZN(new_n18418_));
  OAI21_X1   g18226(.A1(new_n17921_), .A2(new_n17938_), .B(new_n18253_), .ZN(new_n18419_));
  XOR2_X1    g18227(.A1(new_n18419_), .A2(new_n17848_), .Z(new_n18420_));
  NOR2_X1    g18228(.A1(new_n17934_), .A2(\asqrt[9] ), .ZN(new_n18421_));
  OAI21_X1   g18229(.A1(new_n18421_), .A2(new_n17920_), .B(new_n18253_), .ZN(new_n18422_));
  XOR2_X1    g18230(.A1(new_n18422_), .A2(new_n17851_), .Z(new_n18423_));
  OAI21_X1   g18231(.A1(new_n17933_), .A2(new_n17899_), .B(new_n18253_), .ZN(new_n18424_));
  XOR2_X1    g18232(.A1(new_n18424_), .A2(new_n17932_), .Z(new_n18425_));
  INV_X1     g18233(.I(new_n18425_), .ZN(new_n18426_));
  NOR2_X1    g18234(.A1(new_n17895_), .A2(\asqrt[7] ), .ZN(new_n18427_));
  OAI21_X1   g18235(.A1(new_n18427_), .A2(new_n17918_), .B(new_n18253_), .ZN(new_n18428_));
  XOR2_X1    g18236(.A1(new_n18428_), .A2(new_n17903_), .Z(new_n18429_));
  INV_X1     g18237(.I(new_n18429_), .ZN(new_n18430_));
  OAI21_X1   g18238(.A1(new_n17893_), .A2(new_n17915_), .B(new_n18253_), .ZN(new_n18431_));
  XOR2_X1    g18239(.A1(new_n18431_), .A2(new_n17879_), .Z(new_n18432_));
  NOR2_X1    g18240(.A1(new_n17867_), .A2(\a[8] ), .ZN(new_n18433_));
  INV_X1     g18241(.I(new_n18433_), .ZN(new_n18434_));
  NOR2_X1    g18242(.A1(new_n17887_), .A2(\a[8] ), .ZN(new_n18435_));
  AOI22_X1   g18243(.A1(new_n18434_), .A2(new_n17887_), .B1(\asqrt[4] ), .B2(new_n18435_), .ZN(new_n18436_));
  NOR2_X1    g18244(.A1(new_n17885_), .A2(new_n17912_), .ZN(new_n18437_));
  INV_X1     g18245(.I(new_n18437_), .ZN(new_n18438_));
  NAND2_X1   g18246(.A1(\asqrt[3] ), .A2(new_n18438_), .ZN(new_n18439_));
  NOR2_X1    g18247(.A1(new_n18437_), .A2(new_n18436_), .ZN(new_n18440_));
  AOI22_X1   g18248(.A1(new_n18439_), .A2(new_n18436_), .B1(\asqrt[3] ), .B2(new_n18440_), .ZN(new_n18441_));
  NOR2_X1    g18249(.A1(new_n18249_), .A2(new_n18251_), .ZN(new_n18442_));
  INV_X1     g18250(.I(new_n18442_), .ZN(new_n18443_));
  NOR2_X1    g18251(.A1(new_n18246_), .A2(new_n17867_), .ZN(new_n18444_));
  NAND4_X1   g18252(.A1(new_n18303_), .A2(new_n193_), .A3(new_n18443_), .A4(new_n18444_), .ZN(new_n18445_));
  NAND2_X1   g18253(.A1(\asqrt[3] ), .A2(new_n17880_), .ZN(new_n18446_));
  AOI21_X1   g18254(.A1(new_n18446_), .A2(new_n18445_), .B(\a[8] ), .ZN(new_n18447_));
  INV_X1     g18255(.I(new_n18447_), .ZN(new_n18448_));
  NAND3_X1   g18256(.A1(new_n18446_), .A2(\a[8] ), .A3(new_n18445_), .ZN(new_n18449_));
  NAND2_X1   g18257(.A1(new_n18448_), .A2(new_n18449_), .ZN(new_n18450_));
  NOR2_X1    g18258(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n18451_));
  INV_X1     g18259(.I(new_n18451_), .ZN(new_n18452_));
  NAND3_X1   g18260(.A1(\asqrt[3] ), .A2(\a[6] ), .A3(new_n18452_), .ZN(new_n18453_));
  INV_X1     g18261(.I(\a[6] ), .ZN(new_n18454_));
  OAI21_X1   g18262(.A1(\asqrt[3] ), .A2(new_n18454_), .B(new_n18451_), .ZN(new_n18455_));
  AOI21_X1   g18263(.A1(new_n18455_), .A2(new_n18453_), .B(new_n17867_), .ZN(new_n18456_));
  OAI21_X1   g18264(.A1(new_n18253_), .A2(\a[6] ), .B(\a[7] ), .ZN(new_n18457_));
  INV_X1     g18265(.I(\a[7] ), .ZN(new_n18458_));
  NAND3_X1   g18266(.A1(\asqrt[3] ), .A2(new_n18454_), .A3(new_n18458_), .ZN(new_n18459_));
  NOR3_X1    g18267(.A1(new_n17863_), .A2(\asqrt[63] ), .A3(new_n17866_), .ZN(new_n18460_));
  AOI21_X1   g18268(.A1(new_n18460_), .A2(new_n17657_), .B(new_n18454_), .ZN(new_n18461_));
  NAND2_X1   g18269(.A1(\asqrt[3] ), .A2(new_n18461_), .ZN(new_n18462_));
  NAND3_X1   g18270(.A1(new_n18457_), .A2(new_n18459_), .A3(new_n18462_), .ZN(new_n18463_));
  NOR3_X1    g18271(.A1(new_n18456_), .A2(new_n18463_), .A3(\asqrt[5] ), .ZN(new_n18464_));
  OAI21_X1   g18272(.A1(new_n18456_), .A2(new_n18463_), .B(\asqrt[5] ), .ZN(new_n18465_));
  OAI21_X1   g18273(.A1(new_n18450_), .A2(new_n18464_), .B(new_n18465_), .ZN(new_n18466_));
  OAI21_X1   g18274(.A1(new_n18466_), .A2(\asqrt[6] ), .B(new_n18441_), .ZN(new_n18467_));
  NAND2_X1   g18275(.A1(new_n18466_), .A2(\asqrt[6] ), .ZN(new_n18468_));
  NAND3_X1   g18276(.A1(new_n18467_), .A2(new_n18468_), .A3(new_n16269_), .ZN(new_n18469_));
  AOI21_X1   g18277(.A1(new_n18467_), .A2(new_n18468_), .B(new_n16269_), .ZN(new_n18470_));
  AOI21_X1   g18278(.A1(new_n18432_), .A2(new_n18469_), .B(new_n18470_), .ZN(new_n18471_));
  AOI21_X1   g18279(.A1(new_n18471_), .A2(new_n15717_), .B(new_n18430_), .ZN(new_n18472_));
  NAND2_X1   g18280(.A1(new_n18469_), .A2(new_n18432_), .ZN(new_n18473_));
  INV_X1     g18281(.I(new_n18470_), .ZN(new_n18474_));
  AOI21_X1   g18282(.A1(new_n18473_), .A2(new_n18474_), .B(new_n15717_), .ZN(new_n18475_));
  NOR3_X1    g18283(.A1(new_n18472_), .A2(\asqrt[9] ), .A3(new_n18475_), .ZN(new_n18476_));
  OAI21_X1   g18284(.A1(new_n18472_), .A2(new_n18475_), .B(\asqrt[9] ), .ZN(new_n18477_));
  OAI21_X1   g18285(.A1(new_n18426_), .A2(new_n18476_), .B(new_n18477_), .ZN(new_n18478_));
  OAI21_X1   g18286(.A1(new_n18478_), .A2(\asqrt[10] ), .B(new_n18423_), .ZN(new_n18479_));
  NAND2_X1   g18287(.A1(new_n18478_), .A2(\asqrt[10] ), .ZN(new_n18480_));
  NAND3_X1   g18288(.A1(new_n18479_), .A2(new_n18480_), .A3(new_n14207_), .ZN(new_n18481_));
  AOI21_X1   g18289(.A1(new_n18479_), .A2(new_n18480_), .B(new_n14207_), .ZN(new_n18482_));
  AOI21_X1   g18290(.A1(new_n18420_), .A2(new_n18481_), .B(new_n18482_), .ZN(new_n18483_));
  AOI21_X1   g18291(.A1(new_n18483_), .A2(new_n13690_), .B(new_n18418_), .ZN(new_n18484_));
  NAND2_X1   g18292(.A1(new_n18481_), .A2(new_n18420_), .ZN(new_n18485_));
  INV_X1     g18293(.I(new_n18482_), .ZN(new_n18486_));
  AOI21_X1   g18294(.A1(new_n18485_), .A2(new_n18486_), .B(new_n13690_), .ZN(new_n18487_));
  NOR3_X1    g18295(.A1(new_n18484_), .A2(\asqrt[13] ), .A3(new_n18487_), .ZN(new_n18488_));
  OAI21_X1   g18296(.A1(new_n18484_), .A2(new_n18487_), .B(\asqrt[13] ), .ZN(new_n18489_));
  OAI21_X1   g18297(.A1(new_n18414_), .A2(new_n18488_), .B(new_n18489_), .ZN(new_n18490_));
  OAI21_X1   g18298(.A1(new_n18490_), .A2(\asqrt[14] ), .B(new_n18411_), .ZN(new_n18491_));
  NAND2_X1   g18299(.A1(new_n18490_), .A2(\asqrt[14] ), .ZN(new_n18492_));
  NAND3_X1   g18300(.A1(new_n18491_), .A2(new_n18492_), .A3(new_n12283_), .ZN(new_n18493_));
  AOI21_X1   g18301(.A1(new_n18491_), .A2(new_n18492_), .B(new_n12283_), .ZN(new_n18494_));
  AOI21_X1   g18302(.A1(new_n18408_), .A2(new_n18493_), .B(new_n18494_), .ZN(new_n18495_));
  AOI21_X1   g18303(.A1(new_n18495_), .A2(new_n11802_), .B(new_n18406_), .ZN(new_n18496_));
  NAND2_X1   g18304(.A1(new_n18493_), .A2(new_n18408_), .ZN(new_n18497_));
  INV_X1     g18305(.I(new_n18494_), .ZN(new_n18498_));
  AOI21_X1   g18306(.A1(new_n18497_), .A2(new_n18498_), .B(new_n11802_), .ZN(new_n18499_));
  NOR3_X1    g18307(.A1(new_n18496_), .A2(\asqrt[17] ), .A3(new_n18499_), .ZN(new_n18500_));
  OAI21_X1   g18308(.A1(new_n18496_), .A2(new_n18499_), .B(\asqrt[17] ), .ZN(new_n18501_));
  OAI21_X1   g18309(.A1(new_n18402_), .A2(new_n18500_), .B(new_n18501_), .ZN(new_n18502_));
  OAI21_X1   g18310(.A1(new_n18502_), .A2(\asqrt[18] ), .B(new_n18399_), .ZN(new_n18503_));
  NAND2_X1   g18311(.A1(new_n18502_), .A2(\asqrt[18] ), .ZN(new_n18504_));
  NAND3_X1   g18312(.A1(new_n18503_), .A2(new_n18504_), .A3(new_n10497_), .ZN(new_n18505_));
  AOI21_X1   g18313(.A1(new_n18503_), .A2(new_n18504_), .B(new_n10497_), .ZN(new_n18506_));
  AOI21_X1   g18314(.A1(new_n18396_), .A2(new_n18505_), .B(new_n18506_), .ZN(new_n18507_));
  AOI21_X1   g18315(.A1(new_n18507_), .A2(new_n10052_), .B(new_n18394_), .ZN(new_n18508_));
  NAND2_X1   g18316(.A1(new_n18505_), .A2(new_n18396_), .ZN(new_n18509_));
  INV_X1     g18317(.I(new_n18506_), .ZN(new_n18510_));
  AOI21_X1   g18318(.A1(new_n18509_), .A2(new_n18510_), .B(new_n10052_), .ZN(new_n18511_));
  NOR3_X1    g18319(.A1(new_n18508_), .A2(\asqrt[21] ), .A3(new_n18511_), .ZN(new_n18512_));
  OAI21_X1   g18320(.A1(new_n18508_), .A2(new_n18511_), .B(\asqrt[21] ), .ZN(new_n18513_));
  OAI21_X1   g18321(.A1(new_n18390_), .A2(new_n18512_), .B(new_n18513_), .ZN(new_n18514_));
  OAI21_X1   g18322(.A1(new_n18514_), .A2(\asqrt[22] ), .B(new_n18387_), .ZN(new_n18515_));
  NAND2_X1   g18323(.A1(new_n18514_), .A2(\asqrt[22] ), .ZN(new_n18516_));
  NAND3_X1   g18324(.A1(new_n18515_), .A2(new_n18516_), .A3(new_n8849_), .ZN(new_n18517_));
  AOI21_X1   g18325(.A1(new_n18515_), .A2(new_n18516_), .B(new_n8849_), .ZN(new_n18518_));
  AOI21_X1   g18326(.A1(new_n18384_), .A2(new_n18517_), .B(new_n18518_), .ZN(new_n18519_));
  AOI21_X1   g18327(.A1(new_n18519_), .A2(new_n8440_), .B(new_n18382_), .ZN(new_n18520_));
  NAND2_X1   g18328(.A1(new_n18517_), .A2(new_n18384_), .ZN(new_n18521_));
  INV_X1     g18329(.I(new_n18518_), .ZN(new_n18522_));
  AOI21_X1   g18330(.A1(new_n18521_), .A2(new_n18522_), .B(new_n8440_), .ZN(new_n18523_));
  NOR3_X1    g18331(.A1(new_n18520_), .A2(\asqrt[25] ), .A3(new_n18523_), .ZN(new_n18524_));
  OAI21_X1   g18332(.A1(new_n18520_), .A2(new_n18523_), .B(\asqrt[25] ), .ZN(new_n18525_));
  OAI21_X1   g18333(.A1(new_n18378_), .A2(new_n18524_), .B(new_n18525_), .ZN(new_n18526_));
  OAI21_X1   g18334(.A1(new_n18526_), .A2(\asqrt[26] ), .B(new_n18375_), .ZN(new_n18527_));
  NAND2_X1   g18335(.A1(new_n18526_), .A2(\asqrt[26] ), .ZN(new_n18528_));
  NAND3_X1   g18336(.A1(new_n18527_), .A2(new_n18528_), .A3(new_n7331_), .ZN(new_n18529_));
  AOI21_X1   g18337(.A1(new_n18527_), .A2(new_n18528_), .B(new_n7331_), .ZN(new_n18530_));
  AOI21_X1   g18338(.A1(new_n18372_), .A2(new_n18529_), .B(new_n18530_), .ZN(new_n18531_));
  AOI21_X1   g18339(.A1(new_n18531_), .A2(new_n6966_), .B(new_n18370_), .ZN(new_n18532_));
  NAND2_X1   g18340(.A1(new_n18529_), .A2(new_n18372_), .ZN(new_n18533_));
  INV_X1     g18341(.I(new_n18530_), .ZN(new_n18534_));
  AOI21_X1   g18342(.A1(new_n18533_), .A2(new_n18534_), .B(new_n6966_), .ZN(new_n18535_));
  NOR3_X1    g18343(.A1(new_n18532_), .A2(\asqrt[29] ), .A3(new_n18535_), .ZN(new_n18536_));
  OAI21_X1   g18344(.A1(new_n18532_), .A2(new_n18535_), .B(\asqrt[29] ), .ZN(new_n18537_));
  OAI21_X1   g18345(.A1(new_n18366_), .A2(new_n18536_), .B(new_n18537_), .ZN(new_n18538_));
  OAI21_X1   g18346(.A1(new_n18538_), .A2(\asqrt[30] ), .B(new_n18363_), .ZN(new_n18539_));
  NAND2_X1   g18347(.A1(new_n18538_), .A2(\asqrt[30] ), .ZN(new_n18540_));
  NAND3_X1   g18348(.A1(new_n18539_), .A2(new_n18540_), .A3(new_n5947_), .ZN(new_n18541_));
  AOI21_X1   g18349(.A1(new_n18539_), .A2(new_n18540_), .B(new_n5947_), .ZN(new_n18542_));
  AOI21_X1   g18350(.A1(new_n18360_), .A2(new_n18541_), .B(new_n18542_), .ZN(new_n18543_));
  AOI21_X1   g18351(.A1(new_n18543_), .A2(new_n5643_), .B(new_n18358_), .ZN(new_n18544_));
  NAND2_X1   g18352(.A1(new_n18541_), .A2(new_n18360_), .ZN(new_n18545_));
  INV_X1     g18353(.I(new_n18542_), .ZN(new_n18546_));
  AOI21_X1   g18354(.A1(new_n18545_), .A2(new_n18546_), .B(new_n5643_), .ZN(new_n18547_));
  NOR3_X1    g18355(.A1(new_n18544_), .A2(\asqrt[33] ), .A3(new_n18547_), .ZN(new_n18548_));
  OAI21_X1   g18356(.A1(new_n18544_), .A2(new_n18547_), .B(\asqrt[33] ), .ZN(new_n18549_));
  OAI21_X1   g18357(.A1(new_n18354_), .A2(new_n18548_), .B(new_n18549_), .ZN(new_n18550_));
  OAI21_X1   g18358(.A1(new_n18550_), .A2(\asqrt[34] ), .B(new_n18351_), .ZN(new_n18551_));
  NAND2_X1   g18359(.A1(new_n18550_), .A2(\asqrt[34] ), .ZN(new_n18552_));
  NAND3_X1   g18360(.A1(new_n18551_), .A2(new_n18552_), .A3(new_n4751_), .ZN(new_n18553_));
  AOI21_X1   g18361(.A1(new_n18551_), .A2(new_n18552_), .B(new_n4751_), .ZN(new_n18554_));
  AOI21_X1   g18362(.A1(new_n18348_), .A2(new_n18553_), .B(new_n18554_), .ZN(new_n18555_));
  AOI21_X1   g18363(.A1(new_n18555_), .A2(new_n4461_), .B(new_n18346_), .ZN(new_n18556_));
  NAND2_X1   g18364(.A1(new_n18553_), .A2(new_n18348_), .ZN(new_n18557_));
  INV_X1     g18365(.I(new_n18554_), .ZN(new_n18558_));
  AOI21_X1   g18366(.A1(new_n18557_), .A2(new_n18558_), .B(new_n4461_), .ZN(new_n18559_));
  NOR3_X1    g18367(.A1(new_n18556_), .A2(\asqrt[37] ), .A3(new_n18559_), .ZN(new_n18560_));
  OAI21_X1   g18368(.A1(new_n18556_), .A2(new_n18559_), .B(\asqrt[37] ), .ZN(new_n18561_));
  OAI21_X1   g18369(.A1(new_n18342_), .A2(new_n18560_), .B(new_n18561_), .ZN(new_n18562_));
  OAI21_X1   g18370(.A1(new_n18562_), .A2(\asqrt[38] ), .B(new_n18339_), .ZN(new_n18563_));
  NAND2_X1   g18371(.A1(new_n18562_), .A2(\asqrt[38] ), .ZN(new_n18564_));
  NAND3_X1   g18372(.A1(new_n18563_), .A2(new_n18564_), .A3(new_n3681_), .ZN(new_n18565_));
  AOI21_X1   g18373(.A1(new_n18563_), .A2(new_n18564_), .B(new_n3681_), .ZN(new_n18566_));
  AOI21_X1   g18374(.A1(new_n18336_), .A2(new_n18565_), .B(new_n18566_), .ZN(new_n18567_));
  AOI21_X1   g18375(.A1(new_n18567_), .A2(new_n3427_), .B(new_n18334_), .ZN(new_n18568_));
  NAND2_X1   g18376(.A1(new_n18565_), .A2(new_n18336_), .ZN(new_n18569_));
  INV_X1     g18377(.I(new_n18566_), .ZN(new_n18570_));
  AOI21_X1   g18378(.A1(new_n18569_), .A2(new_n18570_), .B(new_n3427_), .ZN(new_n18571_));
  NOR3_X1    g18379(.A1(new_n18568_), .A2(\asqrt[41] ), .A3(new_n18571_), .ZN(new_n18572_));
  OAI21_X1   g18380(.A1(new_n18568_), .A2(new_n18571_), .B(\asqrt[41] ), .ZN(new_n18573_));
  OAI21_X1   g18381(.A1(new_n18330_), .A2(new_n18572_), .B(new_n18573_), .ZN(new_n18574_));
  OAI21_X1   g18382(.A1(new_n18574_), .A2(\asqrt[42] ), .B(new_n18327_), .ZN(new_n18575_));
  NAND2_X1   g18383(.A1(new_n18574_), .A2(\asqrt[42] ), .ZN(new_n18576_));
  NAND3_X1   g18384(.A1(new_n18575_), .A2(new_n18576_), .A3(new_n2749_), .ZN(new_n18577_));
  AOI21_X1   g18385(.A1(new_n18575_), .A2(new_n18576_), .B(new_n2749_), .ZN(new_n18578_));
  AOI21_X1   g18386(.A1(new_n18324_), .A2(new_n18577_), .B(new_n18578_), .ZN(new_n18579_));
  AOI21_X1   g18387(.A1(new_n18579_), .A2(new_n2531_), .B(new_n18322_), .ZN(new_n18580_));
  NAND2_X1   g18388(.A1(new_n18577_), .A2(new_n18324_), .ZN(new_n18581_));
  INV_X1     g18389(.I(new_n18578_), .ZN(new_n18582_));
  AOI21_X1   g18390(.A1(new_n18581_), .A2(new_n18582_), .B(new_n2531_), .ZN(new_n18583_));
  NOR3_X1    g18391(.A1(new_n18580_), .A2(\asqrt[45] ), .A3(new_n18583_), .ZN(new_n18584_));
  OAI21_X1   g18392(.A1(new_n18580_), .A2(new_n18583_), .B(\asqrt[45] ), .ZN(new_n18585_));
  OAI21_X1   g18393(.A1(new_n18318_), .A2(new_n18584_), .B(new_n18585_), .ZN(new_n18586_));
  OAI21_X1   g18394(.A1(new_n18586_), .A2(\asqrt[46] ), .B(new_n18315_), .ZN(new_n18587_));
  NAND2_X1   g18395(.A1(new_n18586_), .A2(\asqrt[46] ), .ZN(new_n18588_));
  NAND3_X1   g18396(.A1(new_n18587_), .A2(new_n18588_), .A3(new_n1953_), .ZN(new_n18589_));
  AOI21_X1   g18397(.A1(new_n18587_), .A2(new_n18588_), .B(new_n1953_), .ZN(new_n18590_));
  AOI21_X1   g18398(.A1(new_n18312_), .A2(new_n18589_), .B(new_n18590_), .ZN(new_n18591_));
  AOI21_X1   g18399(.A1(new_n18591_), .A2(new_n1778_), .B(new_n18310_), .ZN(new_n18592_));
  NAND2_X1   g18400(.A1(new_n18589_), .A2(new_n18312_), .ZN(new_n18593_));
  INV_X1     g18401(.I(new_n18590_), .ZN(new_n18594_));
  AOI21_X1   g18402(.A1(new_n18593_), .A2(new_n18594_), .B(new_n1778_), .ZN(new_n18595_));
  NOR3_X1    g18403(.A1(new_n18592_), .A2(\asqrt[49] ), .A3(new_n18595_), .ZN(new_n18596_));
  OAI21_X1   g18404(.A1(new_n18592_), .A2(new_n18595_), .B(\asqrt[49] ), .ZN(new_n18597_));
  OAI21_X1   g18405(.A1(new_n18296_), .A2(new_n18596_), .B(new_n18597_), .ZN(new_n18598_));
  OAI21_X1   g18406(.A1(new_n18598_), .A2(\asqrt[50] ), .B(new_n18293_), .ZN(new_n18599_));
  NAND2_X1   g18407(.A1(new_n18598_), .A2(\asqrt[50] ), .ZN(new_n18600_));
  NAND3_X1   g18408(.A1(new_n18599_), .A2(new_n18600_), .A3(new_n1305_), .ZN(new_n18601_));
  AOI21_X1   g18409(.A1(new_n18599_), .A2(new_n18600_), .B(new_n1305_), .ZN(new_n18602_));
  AOI21_X1   g18410(.A1(new_n18290_), .A2(new_n18601_), .B(new_n18602_), .ZN(new_n18603_));
  AOI21_X1   g18411(.A1(new_n18603_), .A2(new_n1150_), .B(new_n18288_), .ZN(new_n18604_));
  NAND2_X1   g18412(.A1(new_n18601_), .A2(new_n18290_), .ZN(new_n18605_));
  INV_X1     g18413(.I(new_n18602_), .ZN(new_n18606_));
  AOI21_X1   g18414(.A1(new_n18605_), .A2(new_n18606_), .B(new_n1150_), .ZN(new_n18607_));
  NOR3_X1    g18415(.A1(new_n18604_), .A2(\asqrt[53] ), .A3(new_n18607_), .ZN(new_n18608_));
  OAI21_X1   g18416(.A1(new_n18604_), .A2(new_n18607_), .B(\asqrt[53] ), .ZN(new_n18609_));
  OAI21_X1   g18417(.A1(new_n18283_), .A2(new_n18608_), .B(new_n18609_), .ZN(new_n18610_));
  OAI21_X1   g18418(.A1(new_n18610_), .A2(\asqrt[54] ), .B(new_n18280_), .ZN(new_n18611_));
  NAND2_X1   g18419(.A1(new_n18610_), .A2(\asqrt[54] ), .ZN(new_n18612_));
  NAND3_X1   g18420(.A1(new_n18611_), .A2(new_n18612_), .A3(new_n744_), .ZN(new_n18613_));
  AOI21_X1   g18421(.A1(new_n18611_), .A2(new_n18612_), .B(new_n744_), .ZN(new_n18614_));
  AOI21_X1   g18422(.A1(new_n18277_), .A2(new_n18613_), .B(new_n18614_), .ZN(new_n18615_));
  AOI21_X1   g18423(.A1(new_n18615_), .A2(new_n634_), .B(new_n18275_), .ZN(new_n18616_));
  NAND2_X1   g18424(.A1(new_n18613_), .A2(new_n18277_), .ZN(new_n18617_));
  INV_X1     g18425(.I(new_n18614_), .ZN(new_n18618_));
  AOI21_X1   g18426(.A1(new_n18617_), .A2(new_n18618_), .B(new_n634_), .ZN(new_n18619_));
  NOR3_X1    g18427(.A1(new_n18616_), .A2(\asqrt[57] ), .A3(new_n18619_), .ZN(new_n18620_));
  OAI21_X1   g18428(.A1(new_n18616_), .A2(new_n18619_), .B(\asqrt[57] ), .ZN(new_n18621_));
  OAI21_X1   g18429(.A1(new_n18270_), .A2(new_n18620_), .B(new_n18621_), .ZN(new_n18622_));
  OAI21_X1   g18430(.A1(new_n18622_), .A2(\asqrt[58] ), .B(new_n18267_), .ZN(new_n18623_));
  NOR2_X1    g18431(.A1(new_n18620_), .A2(new_n18270_), .ZN(new_n18624_));
  INV_X1     g18432(.I(new_n18621_), .ZN(new_n18625_));
  OAI21_X1   g18433(.A1(new_n18624_), .A2(new_n18625_), .B(\asqrt[58] ), .ZN(new_n18626_));
  NAND3_X1   g18434(.A1(new_n18623_), .A2(new_n337_), .A3(new_n18626_), .ZN(new_n18627_));
  NAND2_X1   g18435(.A1(new_n18627_), .A2(new_n18264_), .ZN(new_n18628_));
  INV_X1     g18436(.I(new_n18267_), .ZN(new_n18629_));
  NOR2_X1    g18437(.A1(new_n18624_), .A2(new_n18625_), .ZN(new_n18630_));
  AOI21_X1   g18438(.A1(new_n18630_), .A2(new_n423_), .B(new_n18629_), .ZN(new_n18631_));
  INV_X1     g18439(.I(new_n18277_), .ZN(new_n18632_));
  INV_X1     g18440(.I(new_n18290_), .ZN(new_n18633_));
  INV_X1     g18441(.I(new_n18312_), .ZN(new_n18634_));
  INV_X1     g18442(.I(new_n18324_), .ZN(new_n18635_));
  INV_X1     g18443(.I(new_n18336_), .ZN(new_n18636_));
  INV_X1     g18444(.I(new_n18348_), .ZN(new_n18637_));
  INV_X1     g18445(.I(new_n18360_), .ZN(new_n18638_));
  INV_X1     g18446(.I(new_n18372_), .ZN(new_n18639_));
  INV_X1     g18447(.I(new_n18384_), .ZN(new_n18640_));
  INV_X1     g18448(.I(new_n18396_), .ZN(new_n18641_));
  INV_X1     g18449(.I(new_n18408_), .ZN(new_n18642_));
  INV_X1     g18450(.I(new_n18420_), .ZN(new_n18643_));
  INV_X1     g18451(.I(new_n18432_), .ZN(new_n18644_));
  INV_X1     g18452(.I(new_n18445_), .ZN(new_n18645_));
  NOR2_X1    g18453(.A1(new_n18253_), .A2(new_n17881_), .ZN(new_n18646_));
  NOR3_X1    g18454(.A1(new_n18645_), .A2(new_n18646_), .A3(new_n17883_), .ZN(new_n18647_));
  NOR2_X1    g18455(.A1(new_n18647_), .A2(new_n18447_), .ZN(new_n18648_));
  NOR3_X1    g18456(.A1(new_n18253_), .A2(new_n18454_), .A3(new_n18451_), .ZN(new_n18649_));
  AOI21_X1   g18457(.A1(new_n18253_), .A2(\a[6] ), .B(new_n18452_), .ZN(new_n18650_));
  OAI21_X1   g18458(.A1(new_n18649_), .A2(new_n18650_), .B(\asqrt[4] ), .ZN(new_n18651_));
  NOR3_X1    g18459(.A1(new_n18253_), .A2(\a[6] ), .A3(\a[7] ), .ZN(new_n18652_));
  INV_X1     g18460(.I(new_n18461_), .ZN(new_n18653_));
  NOR2_X1    g18461(.A1(new_n18253_), .A2(new_n18653_), .ZN(new_n18654_));
  NOR2_X1    g18462(.A1(new_n18652_), .A2(new_n18654_), .ZN(new_n18655_));
  NAND4_X1   g18463(.A1(new_n18651_), .A2(new_n17342_), .A3(new_n18655_), .A4(new_n18457_), .ZN(new_n18656_));
  NAND2_X1   g18464(.A1(new_n18656_), .A2(new_n18648_), .ZN(new_n18657_));
  NAND3_X1   g18465(.A1(new_n18657_), .A2(new_n16779_), .A3(new_n18465_), .ZN(new_n18658_));
  AOI21_X1   g18466(.A1(new_n18657_), .A2(new_n18465_), .B(new_n16779_), .ZN(new_n18659_));
  AOI21_X1   g18467(.A1(new_n18441_), .A2(new_n18658_), .B(new_n18659_), .ZN(new_n18660_));
  AOI21_X1   g18468(.A1(new_n18660_), .A2(new_n16269_), .B(new_n18644_), .ZN(new_n18661_));
  NOR3_X1    g18469(.A1(new_n18661_), .A2(\asqrt[8] ), .A3(new_n18470_), .ZN(new_n18662_));
  OAI21_X1   g18470(.A1(new_n18661_), .A2(new_n18470_), .B(\asqrt[8] ), .ZN(new_n18663_));
  OAI21_X1   g18471(.A1(new_n18430_), .A2(new_n18662_), .B(new_n18663_), .ZN(new_n18664_));
  OAI21_X1   g18472(.A1(new_n18664_), .A2(\asqrt[9] ), .B(new_n18425_), .ZN(new_n18665_));
  NAND3_X1   g18473(.A1(new_n18665_), .A2(new_n14690_), .A3(new_n18477_), .ZN(new_n18666_));
  AOI21_X1   g18474(.A1(new_n18665_), .A2(new_n18477_), .B(new_n14690_), .ZN(new_n18667_));
  AOI21_X1   g18475(.A1(new_n18423_), .A2(new_n18666_), .B(new_n18667_), .ZN(new_n18668_));
  AOI21_X1   g18476(.A1(new_n18668_), .A2(new_n14207_), .B(new_n18643_), .ZN(new_n18669_));
  NOR3_X1    g18477(.A1(new_n18669_), .A2(\asqrt[12] ), .A3(new_n18482_), .ZN(new_n18670_));
  OAI21_X1   g18478(.A1(new_n18669_), .A2(new_n18482_), .B(\asqrt[12] ), .ZN(new_n18671_));
  OAI21_X1   g18479(.A1(new_n18418_), .A2(new_n18670_), .B(new_n18671_), .ZN(new_n18672_));
  OAI21_X1   g18480(.A1(new_n18672_), .A2(\asqrt[13] ), .B(new_n18413_), .ZN(new_n18673_));
  NAND3_X1   g18481(.A1(new_n18673_), .A2(new_n12733_), .A3(new_n18489_), .ZN(new_n18674_));
  AOI21_X1   g18482(.A1(new_n18673_), .A2(new_n18489_), .B(new_n12733_), .ZN(new_n18675_));
  AOI21_X1   g18483(.A1(new_n18411_), .A2(new_n18674_), .B(new_n18675_), .ZN(new_n18676_));
  AOI21_X1   g18484(.A1(new_n18676_), .A2(new_n12283_), .B(new_n18642_), .ZN(new_n18677_));
  NOR3_X1    g18485(.A1(new_n18677_), .A2(\asqrt[16] ), .A3(new_n18494_), .ZN(new_n18678_));
  OAI21_X1   g18486(.A1(new_n18677_), .A2(new_n18494_), .B(\asqrt[16] ), .ZN(new_n18679_));
  OAI21_X1   g18487(.A1(new_n18406_), .A2(new_n18678_), .B(new_n18679_), .ZN(new_n18680_));
  OAI21_X1   g18488(.A1(new_n18680_), .A2(\asqrt[17] ), .B(new_n18401_), .ZN(new_n18681_));
  NAND3_X1   g18489(.A1(new_n18681_), .A2(new_n10914_), .A3(new_n18501_), .ZN(new_n18682_));
  AOI21_X1   g18490(.A1(new_n18681_), .A2(new_n18501_), .B(new_n10914_), .ZN(new_n18683_));
  AOI21_X1   g18491(.A1(new_n18399_), .A2(new_n18682_), .B(new_n18683_), .ZN(new_n18684_));
  AOI21_X1   g18492(.A1(new_n18684_), .A2(new_n10497_), .B(new_n18641_), .ZN(new_n18685_));
  NOR3_X1    g18493(.A1(new_n18685_), .A2(\asqrt[20] ), .A3(new_n18506_), .ZN(new_n18686_));
  OAI21_X1   g18494(.A1(new_n18685_), .A2(new_n18506_), .B(\asqrt[20] ), .ZN(new_n18687_));
  OAI21_X1   g18495(.A1(new_n18394_), .A2(new_n18686_), .B(new_n18687_), .ZN(new_n18688_));
  OAI21_X1   g18496(.A1(new_n18688_), .A2(\asqrt[21] ), .B(new_n18389_), .ZN(new_n18689_));
  NAND3_X1   g18497(.A1(new_n18689_), .A2(new_n9233_), .A3(new_n18513_), .ZN(new_n18690_));
  AOI21_X1   g18498(.A1(new_n18689_), .A2(new_n18513_), .B(new_n9233_), .ZN(new_n18691_));
  AOI21_X1   g18499(.A1(new_n18387_), .A2(new_n18690_), .B(new_n18691_), .ZN(new_n18692_));
  AOI21_X1   g18500(.A1(new_n18692_), .A2(new_n8849_), .B(new_n18640_), .ZN(new_n18693_));
  NOR3_X1    g18501(.A1(new_n18693_), .A2(\asqrt[24] ), .A3(new_n18518_), .ZN(new_n18694_));
  OAI21_X1   g18502(.A1(new_n18693_), .A2(new_n18518_), .B(\asqrt[24] ), .ZN(new_n18695_));
  OAI21_X1   g18503(.A1(new_n18382_), .A2(new_n18694_), .B(new_n18695_), .ZN(new_n18696_));
  OAI21_X1   g18504(.A1(new_n18696_), .A2(\asqrt[25] ), .B(new_n18377_), .ZN(new_n18697_));
  NAND3_X1   g18505(.A1(new_n18697_), .A2(new_n7690_), .A3(new_n18525_), .ZN(new_n18698_));
  AOI21_X1   g18506(.A1(new_n18697_), .A2(new_n18525_), .B(new_n7690_), .ZN(new_n18699_));
  AOI21_X1   g18507(.A1(new_n18375_), .A2(new_n18698_), .B(new_n18699_), .ZN(new_n18700_));
  AOI21_X1   g18508(.A1(new_n18700_), .A2(new_n7331_), .B(new_n18639_), .ZN(new_n18701_));
  NOR3_X1    g18509(.A1(new_n18701_), .A2(\asqrt[28] ), .A3(new_n18530_), .ZN(new_n18702_));
  OAI21_X1   g18510(.A1(new_n18701_), .A2(new_n18530_), .B(\asqrt[28] ), .ZN(new_n18703_));
  OAI21_X1   g18511(.A1(new_n18370_), .A2(new_n18702_), .B(new_n18703_), .ZN(new_n18704_));
  OAI21_X1   g18512(.A1(new_n18704_), .A2(\asqrt[29] ), .B(new_n18365_), .ZN(new_n18705_));
  NAND3_X1   g18513(.A1(new_n18705_), .A2(new_n6275_), .A3(new_n18537_), .ZN(new_n18706_));
  AOI21_X1   g18514(.A1(new_n18705_), .A2(new_n18537_), .B(new_n6275_), .ZN(new_n18707_));
  AOI21_X1   g18515(.A1(new_n18363_), .A2(new_n18706_), .B(new_n18707_), .ZN(new_n18708_));
  AOI21_X1   g18516(.A1(new_n18708_), .A2(new_n5947_), .B(new_n18638_), .ZN(new_n18709_));
  NOR3_X1    g18517(.A1(new_n18709_), .A2(\asqrt[32] ), .A3(new_n18542_), .ZN(new_n18710_));
  OAI21_X1   g18518(.A1(new_n18709_), .A2(new_n18542_), .B(\asqrt[32] ), .ZN(new_n18711_));
  OAI21_X1   g18519(.A1(new_n18358_), .A2(new_n18710_), .B(new_n18711_), .ZN(new_n18712_));
  OAI21_X1   g18520(.A1(new_n18712_), .A2(\asqrt[33] ), .B(new_n18353_), .ZN(new_n18713_));
  NAND3_X1   g18521(.A1(new_n18713_), .A2(new_n5029_), .A3(new_n18549_), .ZN(new_n18714_));
  AOI21_X1   g18522(.A1(new_n18713_), .A2(new_n18549_), .B(new_n5029_), .ZN(new_n18715_));
  AOI21_X1   g18523(.A1(new_n18351_), .A2(new_n18714_), .B(new_n18715_), .ZN(new_n18716_));
  AOI21_X1   g18524(.A1(new_n18716_), .A2(new_n4751_), .B(new_n18637_), .ZN(new_n18717_));
  NOR3_X1    g18525(.A1(new_n18717_), .A2(\asqrt[36] ), .A3(new_n18554_), .ZN(new_n18718_));
  OAI21_X1   g18526(.A1(new_n18717_), .A2(new_n18554_), .B(\asqrt[36] ), .ZN(new_n18719_));
  OAI21_X1   g18527(.A1(new_n18346_), .A2(new_n18718_), .B(new_n18719_), .ZN(new_n18720_));
  OAI21_X1   g18528(.A1(new_n18720_), .A2(\asqrt[37] ), .B(new_n18341_), .ZN(new_n18721_));
  NAND3_X1   g18529(.A1(new_n18721_), .A2(new_n3925_), .A3(new_n18561_), .ZN(new_n18722_));
  AOI21_X1   g18530(.A1(new_n18721_), .A2(new_n18561_), .B(new_n3925_), .ZN(new_n18723_));
  AOI21_X1   g18531(.A1(new_n18339_), .A2(new_n18722_), .B(new_n18723_), .ZN(new_n18724_));
  AOI21_X1   g18532(.A1(new_n18724_), .A2(new_n3681_), .B(new_n18636_), .ZN(new_n18725_));
  NOR3_X1    g18533(.A1(new_n18725_), .A2(\asqrt[40] ), .A3(new_n18566_), .ZN(new_n18726_));
  OAI21_X1   g18534(.A1(new_n18725_), .A2(new_n18566_), .B(\asqrt[40] ), .ZN(new_n18727_));
  OAI21_X1   g18535(.A1(new_n18334_), .A2(new_n18726_), .B(new_n18727_), .ZN(new_n18728_));
  OAI21_X1   g18536(.A1(new_n18728_), .A2(\asqrt[41] ), .B(new_n18329_), .ZN(new_n18729_));
  NAND3_X1   g18537(.A1(new_n18729_), .A2(new_n2960_), .A3(new_n18573_), .ZN(new_n18730_));
  AOI21_X1   g18538(.A1(new_n18729_), .A2(new_n18573_), .B(new_n2960_), .ZN(new_n18731_));
  AOI21_X1   g18539(.A1(new_n18327_), .A2(new_n18730_), .B(new_n18731_), .ZN(new_n18732_));
  AOI21_X1   g18540(.A1(new_n18732_), .A2(new_n2749_), .B(new_n18635_), .ZN(new_n18733_));
  NOR3_X1    g18541(.A1(new_n18733_), .A2(\asqrt[44] ), .A3(new_n18578_), .ZN(new_n18734_));
  OAI21_X1   g18542(.A1(new_n18733_), .A2(new_n18578_), .B(\asqrt[44] ), .ZN(new_n18735_));
  OAI21_X1   g18543(.A1(new_n18322_), .A2(new_n18734_), .B(new_n18735_), .ZN(new_n18736_));
  OAI21_X1   g18544(.A1(new_n18736_), .A2(\asqrt[45] ), .B(new_n18317_), .ZN(new_n18737_));
  NAND3_X1   g18545(.A1(new_n18737_), .A2(new_n2134_), .A3(new_n18585_), .ZN(new_n18738_));
  AOI21_X1   g18546(.A1(new_n18737_), .A2(new_n18585_), .B(new_n2134_), .ZN(new_n18739_));
  AOI21_X1   g18547(.A1(new_n18315_), .A2(new_n18738_), .B(new_n18739_), .ZN(new_n18740_));
  AOI21_X1   g18548(.A1(new_n18740_), .A2(new_n1953_), .B(new_n18634_), .ZN(new_n18741_));
  NOR3_X1    g18549(.A1(new_n18741_), .A2(\asqrt[48] ), .A3(new_n18590_), .ZN(new_n18742_));
  OAI21_X1   g18550(.A1(new_n18741_), .A2(new_n18590_), .B(\asqrt[48] ), .ZN(new_n18743_));
  OAI21_X1   g18551(.A1(new_n18310_), .A2(new_n18742_), .B(new_n18743_), .ZN(new_n18744_));
  OAI21_X1   g18552(.A1(new_n18744_), .A2(\asqrt[49] ), .B(new_n18295_), .ZN(new_n18745_));
  NAND3_X1   g18553(.A1(new_n18745_), .A2(new_n1463_), .A3(new_n18597_), .ZN(new_n18746_));
  AOI21_X1   g18554(.A1(new_n18745_), .A2(new_n18597_), .B(new_n1463_), .ZN(new_n18747_));
  AOI21_X1   g18555(.A1(new_n18293_), .A2(new_n18746_), .B(new_n18747_), .ZN(new_n18748_));
  AOI21_X1   g18556(.A1(new_n18748_), .A2(new_n1305_), .B(new_n18633_), .ZN(new_n18749_));
  NOR3_X1    g18557(.A1(new_n18749_), .A2(\asqrt[52] ), .A3(new_n18602_), .ZN(new_n18750_));
  OAI21_X1   g18558(.A1(new_n18749_), .A2(new_n18602_), .B(\asqrt[52] ), .ZN(new_n18751_));
  OAI21_X1   g18559(.A1(new_n18288_), .A2(new_n18750_), .B(new_n18751_), .ZN(new_n18752_));
  OAI21_X1   g18560(.A1(new_n18752_), .A2(\asqrt[53] ), .B(new_n18282_), .ZN(new_n18753_));
  NAND3_X1   g18561(.A1(new_n18753_), .A2(new_n860_), .A3(new_n18609_), .ZN(new_n18754_));
  AOI21_X1   g18562(.A1(new_n18753_), .A2(new_n18609_), .B(new_n860_), .ZN(new_n18755_));
  AOI21_X1   g18563(.A1(new_n18280_), .A2(new_n18754_), .B(new_n18755_), .ZN(new_n18756_));
  AOI21_X1   g18564(.A1(new_n18756_), .A2(new_n744_), .B(new_n18632_), .ZN(new_n18757_));
  NOR3_X1    g18565(.A1(new_n18757_), .A2(\asqrt[56] ), .A3(new_n18614_), .ZN(new_n18758_));
  OAI21_X1   g18566(.A1(new_n18757_), .A2(new_n18614_), .B(\asqrt[56] ), .ZN(new_n18759_));
  OAI21_X1   g18567(.A1(new_n18275_), .A2(new_n18758_), .B(new_n18759_), .ZN(new_n18760_));
  OAI21_X1   g18568(.A1(new_n18760_), .A2(\asqrt[57] ), .B(new_n18269_), .ZN(new_n18761_));
  AOI21_X1   g18569(.A1(new_n18761_), .A2(new_n18621_), .B(new_n423_), .ZN(new_n18762_));
  OAI21_X1   g18570(.A1(new_n18631_), .A2(new_n18762_), .B(\asqrt[59] ), .ZN(new_n18763_));
  NAND3_X1   g18571(.A1(new_n18628_), .A2(new_n266_), .A3(new_n18763_), .ZN(new_n18764_));
  NAND2_X1   g18572(.A1(new_n18764_), .A2(new_n18262_), .ZN(new_n18765_));
  INV_X1     g18573(.I(new_n18264_), .ZN(new_n18766_));
  NAND3_X1   g18574(.A1(new_n18761_), .A2(new_n423_), .A3(new_n18621_), .ZN(new_n18767_));
  AOI21_X1   g18575(.A1(new_n18267_), .A2(new_n18767_), .B(new_n18762_), .ZN(new_n18768_));
  AOI21_X1   g18576(.A1(new_n18768_), .A2(new_n337_), .B(new_n18766_), .ZN(new_n18769_));
  AOI21_X1   g18577(.A1(new_n18623_), .A2(new_n18626_), .B(new_n337_), .ZN(new_n18770_));
  OAI21_X1   g18578(.A1(new_n18769_), .A2(new_n18770_), .B(\asqrt[60] ), .ZN(new_n18771_));
  AOI21_X1   g18579(.A1(new_n18765_), .A2(new_n18771_), .B(new_n239_), .ZN(new_n18772_));
  AOI21_X1   g18580(.A1(new_n18628_), .A2(new_n18763_), .B(new_n266_), .ZN(new_n18773_));
  AOI21_X1   g18581(.A1(new_n18262_), .A2(new_n18764_), .B(new_n18773_), .ZN(new_n18774_));
  OAI21_X1   g18582(.A1(new_n18231_), .A2(new_n18223_), .B(new_n18253_), .ZN(new_n18775_));
  XOR2_X1    g18583(.A1(new_n18775_), .A2(new_n18219_), .Z(new_n18776_));
  INV_X1     g18584(.I(new_n18776_), .ZN(new_n18777_));
  AOI21_X1   g18585(.A1(new_n18774_), .A2(new_n239_), .B(new_n18777_), .ZN(new_n18778_));
  NOR2_X1    g18586(.A1(new_n18778_), .A2(new_n18772_), .ZN(new_n18779_));
  INV_X1     g18587(.I(new_n18262_), .ZN(new_n18780_));
  AOI21_X1   g18588(.A1(new_n18264_), .A2(new_n18627_), .B(new_n18770_), .ZN(new_n18781_));
  AOI21_X1   g18589(.A1(new_n18781_), .A2(new_n266_), .B(new_n18780_), .ZN(new_n18782_));
  OAI21_X1   g18590(.A1(new_n18782_), .A2(new_n18773_), .B(\asqrt[61] ), .ZN(new_n18783_));
  NOR3_X1    g18591(.A1(new_n18769_), .A2(\asqrt[60] ), .A3(new_n18770_), .ZN(new_n18784_));
  OAI21_X1   g18592(.A1(new_n18780_), .A2(new_n18784_), .B(new_n18771_), .ZN(new_n18785_));
  OAI21_X1   g18593(.A1(new_n18785_), .A2(\asqrt[61] ), .B(new_n18776_), .ZN(new_n18786_));
  AOI21_X1   g18594(.A1(new_n18786_), .A2(new_n18783_), .B(\asqrt[62] ), .ZN(new_n18787_));
  NOR3_X1    g18595(.A1(new_n18778_), .A2(new_n201_), .A3(new_n18772_), .ZN(new_n18788_));
  OAI22_X1   g18596(.A1(new_n18787_), .A2(new_n18788_), .B1(new_n18779_), .B2(new_n18255_), .ZN(new_n18789_));
  NOR2_X1    g18597(.A1(new_n18301_), .A2(new_n18250_), .ZN(new_n18790_));
  OAI21_X1   g18598(.A1(\asqrt[3] ), .A2(new_n18790_), .B(new_n18443_), .ZN(new_n18791_));
  AOI21_X1   g18599(.A1(new_n18789_), .A2(new_n18259_), .B(new_n18791_), .ZN(new_n18792_));
  NAND2_X1   g18600(.A1(new_n18253_), .A2(new_n18226_), .ZN(new_n18793_));
  NAND2_X1   g18601(.A1(new_n18301_), .A2(new_n18226_), .ZN(new_n18794_));
  NAND2_X1   g18602(.A1(new_n18238_), .A2(new_n18250_), .ZN(new_n18795_));
  AOI21_X1   g18603(.A1(new_n18794_), .A2(new_n18795_), .B(new_n193_), .ZN(new_n18796_));
  NAND2_X1   g18604(.A1(new_n18793_), .A2(new_n18796_), .ZN(new_n18797_));
  AOI21_X1   g18605(.A1(new_n18779_), .A2(new_n201_), .B(new_n18256_), .ZN(new_n18798_));
  INV_X1     g18606(.I(new_n18259_), .ZN(new_n18799_));
  OAI21_X1   g18607(.A1(new_n18779_), .A2(new_n201_), .B(new_n18799_), .ZN(new_n18800_));
  OAI21_X1   g18608(.A1(new_n18798_), .A2(new_n18800_), .B(new_n18797_), .ZN(new_n18801_));
  NOR3_X1    g18609(.A1(new_n18792_), .A2(\asqrt[63] ), .A3(new_n18801_), .ZN(new_n18802_));
  NOR3_X1    g18610(.A1(new_n18782_), .A2(\asqrt[61] ), .A3(new_n18773_), .ZN(new_n18803_));
  OAI21_X1   g18611(.A1(new_n18777_), .A2(new_n18803_), .B(new_n18783_), .ZN(new_n18804_));
  XOR2_X1    g18612(.A1(new_n18804_), .A2(new_n201_), .Z(new_n18805_));
  NAND2_X1   g18613(.A1(new_n18802_), .A2(new_n18805_), .ZN(new_n18806_));
  XOR2_X1    g18614(.A1(new_n18806_), .A2(new_n18256_), .Z(new_n18807_));
  INV_X1     g18615(.I(new_n18807_), .ZN(new_n18808_));
  NAND2_X1   g18616(.A1(new_n18763_), .A2(new_n18627_), .ZN(new_n18809_));
  NAND2_X1   g18617(.A1(new_n18802_), .A2(new_n18809_), .ZN(new_n18810_));
  XOR2_X1    g18618(.A1(new_n18810_), .A2(new_n18766_), .Z(new_n18811_));
  INV_X1     g18619(.I(new_n18811_), .ZN(new_n18812_));
  NAND2_X1   g18620(.A1(new_n18767_), .A2(new_n18626_), .ZN(new_n18813_));
  NAND2_X1   g18621(.A1(new_n18802_), .A2(new_n18813_), .ZN(new_n18814_));
  XOR2_X1    g18622(.A1(new_n18814_), .A2(new_n18629_), .Z(new_n18815_));
  INV_X1     g18623(.I(new_n18815_), .ZN(new_n18816_));
  OAI21_X1   g18624(.A1(new_n18620_), .A2(new_n18625_), .B(new_n18802_), .ZN(new_n18817_));
  XOR2_X1    g18625(.A1(new_n18817_), .A2(new_n18270_), .Z(new_n18818_));
  OAI21_X1   g18626(.A1(new_n18758_), .A2(new_n18619_), .B(new_n18802_), .ZN(new_n18819_));
  XOR2_X1    g18627(.A1(new_n18819_), .A2(new_n18275_), .Z(new_n18820_));
  NAND2_X1   g18628(.A1(new_n18618_), .A2(new_n18613_), .ZN(new_n18821_));
  NAND2_X1   g18629(.A1(new_n18802_), .A2(new_n18821_), .ZN(new_n18822_));
  XOR2_X1    g18630(.A1(new_n18822_), .A2(new_n18632_), .Z(new_n18823_));
  INV_X1     g18631(.I(new_n18823_), .ZN(new_n18824_));
  INV_X1     g18632(.I(new_n18280_), .ZN(new_n18825_));
  NAND2_X1   g18633(.A1(new_n18612_), .A2(new_n18754_), .ZN(new_n18826_));
  NAND2_X1   g18634(.A1(new_n18802_), .A2(new_n18826_), .ZN(new_n18827_));
  XOR2_X1    g18635(.A1(new_n18827_), .A2(new_n18825_), .Z(new_n18828_));
  INV_X1     g18636(.I(new_n18828_), .ZN(new_n18829_));
  INV_X1     g18637(.I(new_n18609_), .ZN(new_n18830_));
  OAI21_X1   g18638(.A1(new_n18608_), .A2(new_n18830_), .B(new_n18802_), .ZN(new_n18831_));
  XOR2_X1    g18639(.A1(new_n18831_), .A2(new_n18283_), .Z(new_n18832_));
  OAI21_X1   g18640(.A1(new_n18750_), .A2(new_n18607_), .B(new_n18802_), .ZN(new_n18833_));
  XOR2_X1    g18641(.A1(new_n18833_), .A2(new_n18288_), .Z(new_n18834_));
  NAND2_X1   g18642(.A1(new_n18606_), .A2(new_n18601_), .ZN(new_n18835_));
  NAND2_X1   g18643(.A1(new_n18802_), .A2(new_n18835_), .ZN(new_n18836_));
  XOR2_X1    g18644(.A1(new_n18836_), .A2(new_n18633_), .Z(new_n18837_));
  INV_X1     g18645(.I(new_n18837_), .ZN(new_n18838_));
  INV_X1     g18646(.I(new_n18293_), .ZN(new_n18839_));
  NAND2_X1   g18647(.A1(new_n18600_), .A2(new_n18746_), .ZN(new_n18840_));
  NAND2_X1   g18648(.A1(new_n18802_), .A2(new_n18840_), .ZN(new_n18841_));
  XOR2_X1    g18649(.A1(new_n18841_), .A2(new_n18839_), .Z(new_n18842_));
  INV_X1     g18650(.I(new_n18842_), .ZN(new_n18843_));
  XOR2_X1    g18651(.A1(new_n18744_), .A2(new_n1632_), .Z(new_n18844_));
  NAND2_X1   g18652(.A1(new_n18802_), .A2(new_n18844_), .ZN(new_n18845_));
  XOR2_X1    g18653(.A1(new_n18845_), .A2(new_n18296_), .Z(new_n18846_));
  OAI21_X1   g18654(.A1(new_n18742_), .A2(new_n18595_), .B(new_n18802_), .ZN(new_n18847_));
  XOR2_X1    g18655(.A1(new_n18847_), .A2(new_n18310_), .Z(new_n18848_));
  NAND2_X1   g18656(.A1(new_n18594_), .A2(new_n18589_), .ZN(new_n18849_));
  NAND2_X1   g18657(.A1(new_n18802_), .A2(new_n18849_), .ZN(new_n18850_));
  XOR2_X1    g18658(.A1(new_n18850_), .A2(new_n18634_), .Z(new_n18851_));
  INV_X1     g18659(.I(new_n18851_), .ZN(new_n18852_));
  INV_X1     g18660(.I(new_n18315_), .ZN(new_n18853_));
  NAND2_X1   g18661(.A1(new_n18588_), .A2(new_n18738_), .ZN(new_n18854_));
  NAND2_X1   g18662(.A1(new_n18802_), .A2(new_n18854_), .ZN(new_n18855_));
  XOR2_X1    g18663(.A1(new_n18855_), .A2(new_n18853_), .Z(new_n18856_));
  INV_X1     g18664(.I(new_n18856_), .ZN(new_n18857_));
  XOR2_X1    g18665(.A1(new_n18736_), .A2(new_n2332_), .Z(new_n18858_));
  NAND2_X1   g18666(.A1(new_n18802_), .A2(new_n18858_), .ZN(new_n18859_));
  XOR2_X1    g18667(.A1(new_n18859_), .A2(new_n18318_), .Z(new_n18860_));
  OAI21_X1   g18668(.A1(new_n18734_), .A2(new_n18583_), .B(new_n18802_), .ZN(new_n18861_));
  XOR2_X1    g18669(.A1(new_n18861_), .A2(new_n18322_), .Z(new_n18862_));
  NAND2_X1   g18670(.A1(new_n18582_), .A2(new_n18577_), .ZN(new_n18863_));
  NAND2_X1   g18671(.A1(new_n18802_), .A2(new_n18863_), .ZN(new_n18864_));
  XOR2_X1    g18672(.A1(new_n18864_), .A2(new_n18635_), .Z(new_n18865_));
  INV_X1     g18673(.I(new_n18865_), .ZN(new_n18866_));
  INV_X1     g18674(.I(new_n18327_), .ZN(new_n18867_));
  NAND2_X1   g18675(.A1(new_n18576_), .A2(new_n18730_), .ZN(new_n18868_));
  NAND2_X1   g18676(.A1(new_n18802_), .A2(new_n18868_), .ZN(new_n18869_));
  XOR2_X1    g18677(.A1(new_n18869_), .A2(new_n18867_), .Z(new_n18870_));
  INV_X1     g18678(.I(new_n18870_), .ZN(new_n18871_));
  XOR2_X1    g18679(.A1(new_n18728_), .A2(new_n3195_), .Z(new_n18872_));
  NAND2_X1   g18680(.A1(new_n18802_), .A2(new_n18872_), .ZN(new_n18873_));
  XOR2_X1    g18681(.A1(new_n18873_), .A2(new_n18330_), .Z(new_n18874_));
  OAI21_X1   g18682(.A1(new_n18726_), .A2(new_n18571_), .B(new_n18802_), .ZN(new_n18875_));
  XOR2_X1    g18683(.A1(new_n18875_), .A2(new_n18334_), .Z(new_n18876_));
  NAND2_X1   g18684(.A1(new_n18570_), .A2(new_n18565_), .ZN(new_n18877_));
  NAND2_X1   g18685(.A1(new_n18802_), .A2(new_n18877_), .ZN(new_n18878_));
  XOR2_X1    g18686(.A1(new_n18878_), .A2(new_n18636_), .Z(new_n18879_));
  INV_X1     g18687(.I(new_n18879_), .ZN(new_n18880_));
  INV_X1     g18688(.I(new_n18339_), .ZN(new_n18881_));
  NAND2_X1   g18689(.A1(new_n18564_), .A2(new_n18722_), .ZN(new_n18882_));
  NAND2_X1   g18690(.A1(new_n18802_), .A2(new_n18882_), .ZN(new_n18883_));
  XOR2_X1    g18691(.A1(new_n18883_), .A2(new_n18881_), .Z(new_n18884_));
  INV_X1     g18692(.I(new_n18884_), .ZN(new_n18885_));
  XOR2_X1    g18693(.A1(new_n18720_), .A2(new_n4196_), .Z(new_n18886_));
  NAND2_X1   g18694(.A1(new_n18802_), .A2(new_n18886_), .ZN(new_n18887_));
  XOR2_X1    g18695(.A1(new_n18887_), .A2(new_n18342_), .Z(new_n18888_));
  OAI21_X1   g18696(.A1(new_n18718_), .A2(new_n18559_), .B(new_n18802_), .ZN(new_n18889_));
  XOR2_X1    g18697(.A1(new_n18889_), .A2(new_n18346_), .Z(new_n18890_));
  NAND2_X1   g18698(.A1(new_n18558_), .A2(new_n18553_), .ZN(new_n18891_));
  NAND2_X1   g18699(.A1(new_n18802_), .A2(new_n18891_), .ZN(new_n18892_));
  XOR2_X1    g18700(.A1(new_n18892_), .A2(new_n18637_), .Z(new_n18893_));
  INV_X1     g18701(.I(new_n18893_), .ZN(new_n18894_));
  INV_X1     g18702(.I(new_n18351_), .ZN(new_n18895_));
  NAND2_X1   g18703(.A1(new_n18552_), .A2(new_n18714_), .ZN(new_n18896_));
  NAND2_X1   g18704(.A1(new_n18802_), .A2(new_n18896_), .ZN(new_n18897_));
  XOR2_X1    g18705(.A1(new_n18897_), .A2(new_n18895_), .Z(new_n18898_));
  INV_X1     g18706(.I(new_n18898_), .ZN(new_n18899_));
  XOR2_X1    g18707(.A1(new_n18712_), .A2(new_n5336_), .Z(new_n18900_));
  NAND2_X1   g18708(.A1(new_n18802_), .A2(new_n18900_), .ZN(new_n18901_));
  XOR2_X1    g18709(.A1(new_n18901_), .A2(new_n18354_), .Z(new_n18902_));
  OAI21_X1   g18710(.A1(new_n18710_), .A2(new_n18547_), .B(new_n18802_), .ZN(new_n18903_));
  XOR2_X1    g18711(.A1(new_n18903_), .A2(new_n18358_), .Z(new_n18904_));
  NAND2_X1   g18712(.A1(new_n18546_), .A2(new_n18541_), .ZN(new_n18905_));
  NAND2_X1   g18713(.A1(new_n18802_), .A2(new_n18905_), .ZN(new_n18906_));
  XOR2_X1    g18714(.A1(new_n18906_), .A2(new_n18638_), .Z(new_n18907_));
  INV_X1     g18715(.I(new_n18907_), .ZN(new_n18908_));
  INV_X1     g18716(.I(new_n18363_), .ZN(new_n18909_));
  NAND2_X1   g18717(.A1(new_n18540_), .A2(new_n18706_), .ZN(new_n18910_));
  NAND2_X1   g18718(.A1(new_n18802_), .A2(new_n18910_), .ZN(new_n18911_));
  XOR2_X1    g18719(.A1(new_n18911_), .A2(new_n18909_), .Z(new_n18912_));
  INV_X1     g18720(.I(new_n18912_), .ZN(new_n18913_));
  XOR2_X1    g18721(.A1(new_n18704_), .A2(new_n6636_), .Z(new_n18914_));
  NAND2_X1   g18722(.A1(new_n18802_), .A2(new_n18914_), .ZN(new_n18915_));
  XOR2_X1    g18723(.A1(new_n18915_), .A2(new_n18366_), .Z(new_n18916_));
  OAI21_X1   g18724(.A1(new_n18702_), .A2(new_n18535_), .B(new_n18802_), .ZN(new_n18917_));
  XOR2_X1    g18725(.A1(new_n18917_), .A2(new_n18370_), .Z(new_n18918_));
  NAND2_X1   g18726(.A1(new_n18534_), .A2(new_n18529_), .ZN(new_n18919_));
  NAND2_X1   g18727(.A1(new_n18802_), .A2(new_n18919_), .ZN(new_n18920_));
  XOR2_X1    g18728(.A1(new_n18920_), .A2(new_n18639_), .Z(new_n18921_));
  INV_X1     g18729(.I(new_n18921_), .ZN(new_n18922_));
  INV_X1     g18730(.I(new_n18375_), .ZN(new_n18923_));
  NAND2_X1   g18731(.A1(new_n18528_), .A2(new_n18698_), .ZN(new_n18924_));
  NAND2_X1   g18732(.A1(new_n18802_), .A2(new_n18924_), .ZN(new_n18925_));
  XOR2_X1    g18733(.A1(new_n18925_), .A2(new_n18923_), .Z(new_n18926_));
  INV_X1     g18734(.I(new_n18926_), .ZN(new_n18927_));
  XOR2_X1    g18735(.A1(new_n18696_), .A2(new_n8077_), .Z(new_n18928_));
  NAND2_X1   g18736(.A1(new_n18802_), .A2(new_n18928_), .ZN(new_n18929_));
  XOR2_X1    g18737(.A1(new_n18929_), .A2(new_n18378_), .Z(new_n18930_));
  OAI21_X1   g18738(.A1(new_n18694_), .A2(new_n18523_), .B(new_n18802_), .ZN(new_n18931_));
  XOR2_X1    g18739(.A1(new_n18931_), .A2(new_n18382_), .Z(new_n18932_));
  NAND2_X1   g18740(.A1(new_n18522_), .A2(new_n18517_), .ZN(new_n18933_));
  NAND2_X1   g18741(.A1(new_n18802_), .A2(new_n18933_), .ZN(new_n18934_));
  XOR2_X1    g18742(.A1(new_n18934_), .A2(new_n18640_), .Z(new_n18935_));
  INV_X1     g18743(.I(new_n18935_), .ZN(new_n18936_));
  INV_X1     g18744(.I(new_n18387_), .ZN(new_n18937_));
  NAND2_X1   g18745(.A1(new_n18516_), .A2(new_n18690_), .ZN(new_n18938_));
  NAND2_X1   g18746(.A1(new_n18802_), .A2(new_n18938_), .ZN(new_n18939_));
  XOR2_X1    g18747(.A1(new_n18939_), .A2(new_n18937_), .Z(new_n18940_));
  INV_X1     g18748(.I(new_n18940_), .ZN(new_n18941_));
  XOR2_X1    g18749(.A1(new_n18688_), .A2(new_n9656_), .Z(new_n18942_));
  NAND2_X1   g18750(.A1(new_n18802_), .A2(new_n18942_), .ZN(new_n18943_));
  XOR2_X1    g18751(.A1(new_n18943_), .A2(new_n18390_), .Z(new_n18944_));
  OAI21_X1   g18752(.A1(new_n18686_), .A2(new_n18511_), .B(new_n18802_), .ZN(new_n18945_));
  XOR2_X1    g18753(.A1(new_n18945_), .A2(new_n18394_), .Z(new_n18946_));
  NAND2_X1   g18754(.A1(new_n18510_), .A2(new_n18505_), .ZN(new_n18947_));
  NAND2_X1   g18755(.A1(new_n18802_), .A2(new_n18947_), .ZN(new_n18948_));
  XOR2_X1    g18756(.A1(new_n18948_), .A2(new_n18641_), .Z(new_n18949_));
  INV_X1     g18757(.I(new_n18949_), .ZN(new_n18950_));
  INV_X1     g18758(.I(new_n18399_), .ZN(new_n18951_));
  NAND2_X1   g18759(.A1(new_n18504_), .A2(new_n18682_), .ZN(new_n18952_));
  NAND2_X1   g18760(.A1(new_n18802_), .A2(new_n18952_), .ZN(new_n18953_));
  XOR2_X1    g18761(.A1(new_n18953_), .A2(new_n18951_), .Z(new_n18954_));
  INV_X1     g18762(.I(new_n18954_), .ZN(new_n18955_));
  XOR2_X1    g18763(.A1(new_n18680_), .A2(new_n11373_), .Z(new_n18956_));
  NAND2_X1   g18764(.A1(new_n18802_), .A2(new_n18956_), .ZN(new_n18957_));
  XOR2_X1    g18765(.A1(new_n18957_), .A2(new_n18402_), .Z(new_n18958_));
  OAI21_X1   g18766(.A1(new_n18678_), .A2(new_n18499_), .B(new_n18802_), .ZN(new_n18959_));
  XOR2_X1    g18767(.A1(new_n18959_), .A2(new_n18406_), .Z(new_n18960_));
  NAND2_X1   g18768(.A1(new_n18498_), .A2(new_n18493_), .ZN(new_n18961_));
  NAND2_X1   g18769(.A1(new_n18802_), .A2(new_n18961_), .ZN(new_n18962_));
  XOR2_X1    g18770(.A1(new_n18962_), .A2(new_n18642_), .Z(new_n18963_));
  INV_X1     g18771(.I(new_n18963_), .ZN(new_n18964_));
  INV_X1     g18772(.I(new_n18411_), .ZN(new_n18965_));
  NAND2_X1   g18773(.A1(new_n18492_), .A2(new_n18674_), .ZN(new_n18966_));
  NAND2_X1   g18774(.A1(new_n18802_), .A2(new_n18966_), .ZN(new_n18967_));
  XOR2_X1    g18775(.A1(new_n18967_), .A2(new_n18965_), .Z(new_n18968_));
  INV_X1     g18776(.I(new_n18968_), .ZN(new_n18969_));
  XOR2_X1    g18777(.A1(new_n18672_), .A2(new_n13228_), .Z(new_n18970_));
  NAND2_X1   g18778(.A1(new_n18802_), .A2(new_n18970_), .ZN(new_n18971_));
  XOR2_X1    g18779(.A1(new_n18971_), .A2(new_n18414_), .Z(new_n18972_));
  OAI21_X1   g18780(.A1(new_n18670_), .A2(new_n18487_), .B(new_n18802_), .ZN(new_n18973_));
  XOR2_X1    g18781(.A1(new_n18973_), .A2(new_n18418_), .Z(new_n18974_));
  NAND2_X1   g18782(.A1(new_n18486_), .A2(new_n18481_), .ZN(new_n18975_));
  NAND2_X1   g18783(.A1(new_n18802_), .A2(new_n18975_), .ZN(new_n18976_));
  XOR2_X1    g18784(.A1(new_n18976_), .A2(new_n18643_), .Z(new_n18977_));
  INV_X1     g18785(.I(new_n18977_), .ZN(new_n18978_));
  INV_X1     g18786(.I(new_n18423_), .ZN(new_n18979_));
  NAND2_X1   g18787(.A1(new_n18480_), .A2(new_n18666_), .ZN(new_n18980_));
  NAND2_X1   g18788(.A1(new_n18802_), .A2(new_n18980_), .ZN(new_n18981_));
  XOR2_X1    g18789(.A1(new_n18981_), .A2(new_n18979_), .Z(new_n18982_));
  INV_X1     g18790(.I(new_n18982_), .ZN(new_n18983_));
  XOR2_X1    g18791(.A1(new_n18664_), .A2(new_n15221_), .Z(new_n18984_));
  NAND2_X1   g18792(.A1(new_n18802_), .A2(new_n18984_), .ZN(new_n18985_));
  XOR2_X1    g18793(.A1(new_n18985_), .A2(new_n18426_), .Z(new_n18986_));
  OAI21_X1   g18794(.A1(new_n18662_), .A2(new_n18475_), .B(new_n18802_), .ZN(new_n18987_));
  XOR2_X1    g18795(.A1(new_n18987_), .A2(new_n18430_), .Z(new_n18988_));
  NAND2_X1   g18796(.A1(new_n18474_), .A2(new_n18469_), .ZN(new_n18989_));
  NAND2_X1   g18797(.A1(new_n18802_), .A2(new_n18989_), .ZN(new_n18990_));
  XOR2_X1    g18798(.A1(new_n18990_), .A2(new_n18644_), .Z(new_n18991_));
  INV_X1     g18799(.I(new_n18991_), .ZN(new_n18992_));
  NAND2_X1   g18800(.A1(new_n18468_), .A2(new_n18658_), .ZN(new_n18993_));
  NAND2_X1   g18801(.A1(new_n18802_), .A2(new_n18993_), .ZN(new_n18994_));
  XNOR2_X1   g18802(.A1(new_n18994_), .A2(new_n18441_), .ZN(new_n18995_));
  INV_X1     g18803(.I(new_n18995_), .ZN(new_n18996_));
  NAND2_X1   g18804(.A1(new_n18656_), .A2(new_n18465_), .ZN(new_n18997_));
  NAND2_X1   g18805(.A1(new_n18802_), .A2(new_n18997_), .ZN(new_n18998_));
  XOR2_X1    g18806(.A1(new_n18998_), .A2(new_n18450_), .Z(new_n18999_));
  NOR2_X1    g18807(.A1(new_n18253_), .A2(\a[6] ), .ZN(new_n19000_));
  INV_X1     g18808(.I(new_n19000_), .ZN(new_n19001_));
  NOR2_X1    g18809(.A1(new_n18458_), .A2(\a[6] ), .ZN(new_n19002_));
  AOI22_X1   g18810(.A1(new_n19001_), .A2(new_n18458_), .B1(\asqrt[3] ), .B2(new_n19002_), .ZN(new_n19003_));
  INV_X1     g18811(.I(new_n19003_), .ZN(new_n19004_));
  NOR2_X1    g18812(.A1(new_n18456_), .A2(new_n18654_), .ZN(new_n19005_));
  NOR2_X1    g18813(.A1(new_n18802_), .A2(new_n19005_), .ZN(new_n19006_));
  NOR2_X1    g18814(.A1(new_n19006_), .A2(new_n19004_), .ZN(new_n19007_));
  NOR3_X1    g18815(.A1(new_n18802_), .A2(new_n19003_), .A3(new_n19005_), .ZN(new_n19008_));
  NOR2_X1    g18816(.A1(new_n19007_), .A2(new_n19008_), .ZN(new_n19009_));
  OAI21_X1   g18817(.A1(new_n18778_), .A2(new_n18772_), .B(new_n201_), .ZN(new_n19010_));
  NAND3_X1   g18818(.A1(new_n18786_), .A2(\asqrt[62] ), .A3(new_n18783_), .ZN(new_n19011_));
  AOI22_X1   g18819(.A1(new_n19011_), .A2(new_n19010_), .B1(new_n18256_), .B2(new_n18804_), .ZN(new_n19012_));
  INV_X1     g18820(.I(new_n18791_), .ZN(new_n19013_));
  OAI21_X1   g18821(.A1(new_n19012_), .A2(new_n18799_), .B(new_n19013_), .ZN(new_n19014_));
  NAND2_X1   g18822(.A1(new_n19014_), .A2(new_n193_), .ZN(new_n19015_));
  NOR2_X1    g18823(.A1(new_n18798_), .A2(new_n18800_), .ZN(new_n19016_));
  NAND2_X1   g18824(.A1(new_n18797_), .A2(\asqrt[3] ), .ZN(new_n19017_));
  NOR3_X1    g18825(.A1(new_n19015_), .A2(new_n19016_), .A3(new_n19017_), .ZN(new_n19018_));
  NOR2_X1    g18826(.A1(new_n18802_), .A2(new_n18452_), .ZN(new_n19019_));
  OAI21_X1   g18827(.A1(new_n19019_), .A2(new_n19018_), .B(new_n18454_), .ZN(new_n19020_));
  NOR3_X1    g18828(.A1(new_n19019_), .A2(new_n19018_), .A3(new_n18454_), .ZN(new_n19021_));
  INV_X1     g18829(.I(new_n19021_), .ZN(new_n19022_));
  NAND2_X1   g18830(.A1(new_n19022_), .A2(new_n19020_), .ZN(new_n19023_));
  OAI21_X1   g18831(.A1(new_n18804_), .A2(\asqrt[62] ), .B(new_n18255_), .ZN(new_n19024_));
  AOI21_X1   g18832(.A1(new_n18804_), .A2(\asqrt[62] ), .B(new_n18259_), .ZN(new_n19025_));
  AOI22_X1   g18833(.A1(new_n19025_), .A2(new_n19024_), .B1(new_n18793_), .B2(new_n18796_), .ZN(new_n19026_));
  NAND3_X1   g18834(.A1(new_n19014_), .A2(new_n193_), .A3(new_n19026_), .ZN(\asqrt[2] ));
  NOR2_X1    g18835(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n19028_));
  INV_X1     g18836(.I(new_n19028_), .ZN(new_n19029_));
  NAND3_X1   g18837(.A1(\asqrt[2] ), .A2(\a[4] ), .A3(new_n19029_), .ZN(new_n19030_));
  INV_X1     g18838(.I(\a[4] ), .ZN(new_n19031_));
  OAI21_X1   g18839(.A1(\asqrt[2] ), .A2(new_n19031_), .B(new_n19028_), .ZN(new_n19032_));
  AOI21_X1   g18840(.A1(new_n19032_), .A2(new_n19030_), .B(new_n18253_), .ZN(new_n19033_));
  NAND2_X1   g18841(.A1(new_n18303_), .A2(new_n193_), .ZN(new_n19034_));
  AOI21_X1   g18842(.A1(new_n19031_), .A2(new_n19028_), .B(new_n18246_), .ZN(new_n19035_));
  AOI21_X1   g18843(.A1(new_n18443_), .A2(new_n19035_), .B(new_n19034_), .ZN(new_n19036_));
  INV_X1     g18844(.I(new_n19036_), .ZN(new_n19037_));
  NAND3_X1   g18845(.A1(\asqrt[2] ), .A2(\a[4] ), .A3(new_n19037_), .ZN(new_n19038_));
  INV_X1     g18846(.I(\a[5] ), .ZN(new_n19039_));
  NAND3_X1   g18847(.A1(\asqrt[2] ), .A2(new_n19031_), .A3(new_n19039_), .ZN(new_n19040_));
  OAI21_X1   g18848(.A1(new_n18802_), .A2(\a[4] ), .B(\a[5] ), .ZN(new_n19041_));
  NAND3_X1   g18849(.A1(new_n19038_), .A2(new_n19041_), .A3(new_n19040_), .ZN(new_n19042_));
  NOR3_X1    g18850(.A1(new_n19042_), .A2(new_n19033_), .A3(\asqrt[4] ), .ZN(new_n19043_));
  OAI21_X1   g18851(.A1(new_n19042_), .A2(new_n19033_), .B(\asqrt[4] ), .ZN(new_n19044_));
  OAI21_X1   g18852(.A1(new_n19023_), .A2(new_n19043_), .B(new_n19044_), .ZN(new_n19045_));
  OAI21_X1   g18853(.A1(new_n19045_), .A2(\asqrt[5] ), .B(new_n19009_), .ZN(new_n19046_));
  NAND2_X1   g18854(.A1(new_n19045_), .A2(\asqrt[5] ), .ZN(new_n19047_));
  NAND3_X1   g18855(.A1(new_n19046_), .A2(new_n19047_), .A3(new_n16779_), .ZN(new_n19048_));
  AOI21_X1   g18856(.A1(new_n19046_), .A2(new_n19047_), .B(new_n16779_), .ZN(new_n19049_));
  AOI21_X1   g18857(.A1(new_n18999_), .A2(new_n19048_), .B(new_n19049_), .ZN(new_n19050_));
  AOI21_X1   g18858(.A1(new_n19050_), .A2(new_n16269_), .B(new_n18996_), .ZN(new_n19051_));
  NAND2_X1   g18859(.A1(new_n19048_), .A2(new_n18999_), .ZN(new_n19052_));
  INV_X1     g18860(.I(new_n19009_), .ZN(new_n19053_));
  INV_X1     g18861(.I(new_n19020_), .ZN(new_n19054_));
  NOR2_X1    g18862(.A1(new_n19054_), .A2(new_n19021_), .ZN(new_n19055_));
  NOR3_X1    g18863(.A1(new_n18802_), .A2(new_n19031_), .A3(new_n19028_), .ZN(new_n19056_));
  AOI21_X1   g18864(.A1(new_n18802_), .A2(\a[4] ), .B(new_n19029_), .ZN(new_n19057_));
  OAI21_X1   g18865(.A1(new_n19056_), .A2(new_n19057_), .B(\asqrt[3] ), .ZN(new_n19058_));
  NOR3_X1    g18866(.A1(new_n18802_), .A2(new_n19031_), .A3(new_n19036_), .ZN(new_n19059_));
  NOR3_X1    g18867(.A1(new_n18802_), .A2(\a[4] ), .A3(\a[5] ), .ZN(new_n19060_));
  AOI21_X1   g18868(.A1(\asqrt[2] ), .A2(new_n19031_), .B(new_n19039_), .ZN(new_n19061_));
  NOR3_X1    g18869(.A1(new_n19059_), .A2(new_n19060_), .A3(new_n19061_), .ZN(new_n19062_));
  NAND3_X1   g18870(.A1(new_n19062_), .A2(new_n19058_), .A3(new_n17867_), .ZN(new_n19063_));
  AOI21_X1   g18871(.A1(new_n19062_), .A2(new_n19058_), .B(new_n17867_), .ZN(new_n19064_));
  AOI21_X1   g18872(.A1(new_n19055_), .A2(new_n19063_), .B(new_n19064_), .ZN(new_n19065_));
  AOI21_X1   g18873(.A1(new_n19065_), .A2(new_n17342_), .B(new_n19053_), .ZN(new_n19066_));
  NAND2_X1   g18874(.A1(new_n19055_), .A2(new_n19063_), .ZN(new_n19067_));
  AOI21_X1   g18875(.A1(new_n19067_), .A2(new_n19044_), .B(new_n17342_), .ZN(new_n19068_));
  OAI21_X1   g18876(.A1(new_n19066_), .A2(new_n19068_), .B(\asqrt[6] ), .ZN(new_n19069_));
  AOI21_X1   g18877(.A1(new_n19052_), .A2(new_n19069_), .B(new_n16269_), .ZN(new_n19070_));
  NOR3_X1    g18878(.A1(new_n19051_), .A2(\asqrt[8] ), .A3(new_n19070_), .ZN(new_n19071_));
  OAI21_X1   g18879(.A1(new_n19051_), .A2(new_n19070_), .B(\asqrt[8] ), .ZN(new_n19072_));
  OAI21_X1   g18880(.A1(new_n18992_), .A2(new_n19071_), .B(new_n19072_), .ZN(new_n19073_));
  OAI21_X1   g18881(.A1(new_n19073_), .A2(\asqrt[9] ), .B(new_n18988_), .ZN(new_n19074_));
  NAND2_X1   g18882(.A1(new_n19073_), .A2(\asqrt[9] ), .ZN(new_n19075_));
  NAND3_X1   g18883(.A1(new_n19074_), .A2(new_n19075_), .A3(new_n14690_), .ZN(new_n19076_));
  AOI21_X1   g18884(.A1(new_n19074_), .A2(new_n19075_), .B(new_n14690_), .ZN(new_n19077_));
  AOI21_X1   g18885(.A1(new_n18986_), .A2(new_n19076_), .B(new_n19077_), .ZN(new_n19078_));
  AOI21_X1   g18886(.A1(new_n19078_), .A2(new_n14207_), .B(new_n18983_), .ZN(new_n19079_));
  NAND2_X1   g18887(.A1(new_n19076_), .A2(new_n18986_), .ZN(new_n19080_));
  INV_X1     g18888(.I(new_n18988_), .ZN(new_n19081_));
  INV_X1     g18889(.I(new_n18999_), .ZN(new_n19082_));
  NOR3_X1    g18890(.A1(new_n19066_), .A2(\asqrt[6] ), .A3(new_n19068_), .ZN(new_n19083_));
  OAI21_X1   g18891(.A1(new_n19082_), .A2(new_n19083_), .B(new_n19069_), .ZN(new_n19084_));
  OAI21_X1   g18892(.A1(new_n19084_), .A2(\asqrt[7] ), .B(new_n18995_), .ZN(new_n19085_));
  NAND2_X1   g18893(.A1(new_n19084_), .A2(\asqrt[7] ), .ZN(new_n19086_));
  NAND3_X1   g18894(.A1(new_n19085_), .A2(new_n19086_), .A3(new_n15717_), .ZN(new_n19087_));
  AOI21_X1   g18895(.A1(new_n19085_), .A2(new_n19086_), .B(new_n15717_), .ZN(new_n19088_));
  AOI21_X1   g18896(.A1(new_n18991_), .A2(new_n19087_), .B(new_n19088_), .ZN(new_n19089_));
  AOI21_X1   g18897(.A1(new_n19089_), .A2(new_n15221_), .B(new_n19081_), .ZN(new_n19090_));
  NAND2_X1   g18898(.A1(new_n19087_), .A2(new_n18991_), .ZN(new_n19091_));
  AOI21_X1   g18899(.A1(new_n19091_), .A2(new_n19072_), .B(new_n15221_), .ZN(new_n19092_));
  OAI21_X1   g18900(.A1(new_n19090_), .A2(new_n19092_), .B(\asqrt[10] ), .ZN(new_n19093_));
  AOI21_X1   g18901(.A1(new_n19080_), .A2(new_n19093_), .B(new_n14207_), .ZN(new_n19094_));
  NOR3_X1    g18902(.A1(new_n19079_), .A2(\asqrt[12] ), .A3(new_n19094_), .ZN(new_n19095_));
  OAI21_X1   g18903(.A1(new_n19079_), .A2(new_n19094_), .B(\asqrt[12] ), .ZN(new_n19096_));
  OAI21_X1   g18904(.A1(new_n18978_), .A2(new_n19095_), .B(new_n19096_), .ZN(new_n19097_));
  OAI21_X1   g18905(.A1(new_n19097_), .A2(\asqrt[13] ), .B(new_n18974_), .ZN(new_n19098_));
  NAND2_X1   g18906(.A1(new_n19097_), .A2(\asqrt[13] ), .ZN(new_n19099_));
  NAND3_X1   g18907(.A1(new_n19098_), .A2(new_n19099_), .A3(new_n12733_), .ZN(new_n19100_));
  AOI21_X1   g18908(.A1(new_n19098_), .A2(new_n19099_), .B(new_n12733_), .ZN(new_n19101_));
  AOI21_X1   g18909(.A1(new_n18972_), .A2(new_n19100_), .B(new_n19101_), .ZN(new_n19102_));
  AOI21_X1   g18910(.A1(new_n19102_), .A2(new_n12283_), .B(new_n18969_), .ZN(new_n19103_));
  NAND2_X1   g18911(.A1(new_n19100_), .A2(new_n18972_), .ZN(new_n19104_));
  INV_X1     g18912(.I(new_n18974_), .ZN(new_n19105_));
  INV_X1     g18913(.I(new_n18986_), .ZN(new_n19106_));
  NOR3_X1    g18914(.A1(new_n19090_), .A2(\asqrt[10] ), .A3(new_n19092_), .ZN(new_n19107_));
  OAI21_X1   g18915(.A1(new_n19106_), .A2(new_n19107_), .B(new_n19093_), .ZN(new_n19108_));
  OAI21_X1   g18916(.A1(new_n19108_), .A2(\asqrt[11] ), .B(new_n18982_), .ZN(new_n19109_));
  NAND2_X1   g18917(.A1(new_n19108_), .A2(\asqrt[11] ), .ZN(new_n19110_));
  NAND3_X1   g18918(.A1(new_n19109_), .A2(new_n19110_), .A3(new_n13690_), .ZN(new_n19111_));
  AOI21_X1   g18919(.A1(new_n19109_), .A2(new_n19110_), .B(new_n13690_), .ZN(new_n19112_));
  AOI21_X1   g18920(.A1(new_n18977_), .A2(new_n19111_), .B(new_n19112_), .ZN(new_n19113_));
  AOI21_X1   g18921(.A1(new_n19113_), .A2(new_n13228_), .B(new_n19105_), .ZN(new_n19114_));
  NAND2_X1   g18922(.A1(new_n19111_), .A2(new_n18977_), .ZN(new_n19115_));
  AOI21_X1   g18923(.A1(new_n19115_), .A2(new_n19096_), .B(new_n13228_), .ZN(new_n19116_));
  OAI21_X1   g18924(.A1(new_n19114_), .A2(new_n19116_), .B(\asqrt[14] ), .ZN(new_n19117_));
  AOI21_X1   g18925(.A1(new_n19104_), .A2(new_n19117_), .B(new_n12283_), .ZN(new_n19118_));
  NOR3_X1    g18926(.A1(new_n19103_), .A2(\asqrt[16] ), .A3(new_n19118_), .ZN(new_n19119_));
  OAI21_X1   g18927(.A1(new_n19103_), .A2(new_n19118_), .B(\asqrt[16] ), .ZN(new_n19120_));
  OAI21_X1   g18928(.A1(new_n18964_), .A2(new_n19119_), .B(new_n19120_), .ZN(new_n19121_));
  OAI21_X1   g18929(.A1(new_n19121_), .A2(\asqrt[17] ), .B(new_n18960_), .ZN(new_n19122_));
  NAND2_X1   g18930(.A1(new_n19121_), .A2(\asqrt[17] ), .ZN(new_n19123_));
  NAND3_X1   g18931(.A1(new_n19122_), .A2(new_n19123_), .A3(new_n10914_), .ZN(new_n19124_));
  AOI21_X1   g18932(.A1(new_n19122_), .A2(new_n19123_), .B(new_n10914_), .ZN(new_n19125_));
  AOI21_X1   g18933(.A1(new_n18958_), .A2(new_n19124_), .B(new_n19125_), .ZN(new_n19126_));
  AOI21_X1   g18934(.A1(new_n19126_), .A2(new_n10497_), .B(new_n18955_), .ZN(new_n19127_));
  NAND2_X1   g18935(.A1(new_n19124_), .A2(new_n18958_), .ZN(new_n19128_));
  INV_X1     g18936(.I(new_n18960_), .ZN(new_n19129_));
  INV_X1     g18937(.I(new_n18972_), .ZN(new_n19130_));
  NOR3_X1    g18938(.A1(new_n19114_), .A2(\asqrt[14] ), .A3(new_n19116_), .ZN(new_n19131_));
  OAI21_X1   g18939(.A1(new_n19130_), .A2(new_n19131_), .B(new_n19117_), .ZN(new_n19132_));
  OAI21_X1   g18940(.A1(new_n19132_), .A2(\asqrt[15] ), .B(new_n18968_), .ZN(new_n19133_));
  NAND2_X1   g18941(.A1(new_n19132_), .A2(\asqrt[15] ), .ZN(new_n19134_));
  NAND3_X1   g18942(.A1(new_n19133_), .A2(new_n19134_), .A3(new_n11802_), .ZN(new_n19135_));
  AOI21_X1   g18943(.A1(new_n19133_), .A2(new_n19134_), .B(new_n11802_), .ZN(new_n19136_));
  AOI21_X1   g18944(.A1(new_n18963_), .A2(new_n19135_), .B(new_n19136_), .ZN(new_n19137_));
  AOI21_X1   g18945(.A1(new_n19137_), .A2(new_n11373_), .B(new_n19129_), .ZN(new_n19138_));
  NAND2_X1   g18946(.A1(new_n19135_), .A2(new_n18963_), .ZN(new_n19139_));
  AOI21_X1   g18947(.A1(new_n19139_), .A2(new_n19120_), .B(new_n11373_), .ZN(new_n19140_));
  OAI21_X1   g18948(.A1(new_n19138_), .A2(new_n19140_), .B(\asqrt[18] ), .ZN(new_n19141_));
  AOI21_X1   g18949(.A1(new_n19128_), .A2(new_n19141_), .B(new_n10497_), .ZN(new_n19142_));
  NOR3_X1    g18950(.A1(new_n19127_), .A2(\asqrt[20] ), .A3(new_n19142_), .ZN(new_n19143_));
  OAI21_X1   g18951(.A1(new_n19127_), .A2(new_n19142_), .B(\asqrt[20] ), .ZN(new_n19144_));
  OAI21_X1   g18952(.A1(new_n18950_), .A2(new_n19143_), .B(new_n19144_), .ZN(new_n19145_));
  OAI21_X1   g18953(.A1(new_n19145_), .A2(\asqrt[21] ), .B(new_n18946_), .ZN(new_n19146_));
  NAND2_X1   g18954(.A1(new_n19145_), .A2(\asqrt[21] ), .ZN(new_n19147_));
  NAND3_X1   g18955(.A1(new_n19146_), .A2(new_n19147_), .A3(new_n9233_), .ZN(new_n19148_));
  AOI21_X1   g18956(.A1(new_n19146_), .A2(new_n19147_), .B(new_n9233_), .ZN(new_n19149_));
  AOI21_X1   g18957(.A1(new_n18944_), .A2(new_n19148_), .B(new_n19149_), .ZN(new_n19150_));
  AOI21_X1   g18958(.A1(new_n19150_), .A2(new_n8849_), .B(new_n18941_), .ZN(new_n19151_));
  NAND2_X1   g18959(.A1(new_n19148_), .A2(new_n18944_), .ZN(new_n19152_));
  INV_X1     g18960(.I(new_n18946_), .ZN(new_n19153_));
  INV_X1     g18961(.I(new_n18958_), .ZN(new_n19154_));
  NOR3_X1    g18962(.A1(new_n19138_), .A2(\asqrt[18] ), .A3(new_n19140_), .ZN(new_n19155_));
  OAI21_X1   g18963(.A1(new_n19154_), .A2(new_n19155_), .B(new_n19141_), .ZN(new_n19156_));
  OAI21_X1   g18964(.A1(new_n19156_), .A2(\asqrt[19] ), .B(new_n18954_), .ZN(new_n19157_));
  NAND2_X1   g18965(.A1(new_n19156_), .A2(\asqrt[19] ), .ZN(new_n19158_));
  NAND3_X1   g18966(.A1(new_n19157_), .A2(new_n19158_), .A3(new_n10052_), .ZN(new_n19159_));
  AOI21_X1   g18967(.A1(new_n19157_), .A2(new_n19158_), .B(new_n10052_), .ZN(new_n19160_));
  AOI21_X1   g18968(.A1(new_n18949_), .A2(new_n19159_), .B(new_n19160_), .ZN(new_n19161_));
  AOI21_X1   g18969(.A1(new_n19161_), .A2(new_n9656_), .B(new_n19153_), .ZN(new_n19162_));
  NAND2_X1   g18970(.A1(new_n19159_), .A2(new_n18949_), .ZN(new_n19163_));
  AOI21_X1   g18971(.A1(new_n19163_), .A2(new_n19144_), .B(new_n9656_), .ZN(new_n19164_));
  OAI21_X1   g18972(.A1(new_n19162_), .A2(new_n19164_), .B(\asqrt[22] ), .ZN(new_n19165_));
  AOI21_X1   g18973(.A1(new_n19152_), .A2(new_n19165_), .B(new_n8849_), .ZN(new_n19166_));
  NOR3_X1    g18974(.A1(new_n19151_), .A2(\asqrt[24] ), .A3(new_n19166_), .ZN(new_n19167_));
  OAI21_X1   g18975(.A1(new_n19151_), .A2(new_n19166_), .B(\asqrt[24] ), .ZN(new_n19168_));
  OAI21_X1   g18976(.A1(new_n18936_), .A2(new_n19167_), .B(new_n19168_), .ZN(new_n19169_));
  OAI21_X1   g18977(.A1(new_n19169_), .A2(\asqrt[25] ), .B(new_n18932_), .ZN(new_n19170_));
  NAND2_X1   g18978(.A1(new_n19169_), .A2(\asqrt[25] ), .ZN(new_n19171_));
  NAND3_X1   g18979(.A1(new_n19170_), .A2(new_n19171_), .A3(new_n7690_), .ZN(new_n19172_));
  AOI21_X1   g18980(.A1(new_n19170_), .A2(new_n19171_), .B(new_n7690_), .ZN(new_n19173_));
  AOI21_X1   g18981(.A1(new_n18930_), .A2(new_n19172_), .B(new_n19173_), .ZN(new_n19174_));
  AOI21_X1   g18982(.A1(new_n19174_), .A2(new_n7331_), .B(new_n18927_), .ZN(new_n19175_));
  NAND2_X1   g18983(.A1(new_n19172_), .A2(new_n18930_), .ZN(new_n19176_));
  INV_X1     g18984(.I(new_n18932_), .ZN(new_n19177_));
  INV_X1     g18985(.I(new_n18944_), .ZN(new_n19178_));
  NOR3_X1    g18986(.A1(new_n19162_), .A2(\asqrt[22] ), .A3(new_n19164_), .ZN(new_n19179_));
  OAI21_X1   g18987(.A1(new_n19178_), .A2(new_n19179_), .B(new_n19165_), .ZN(new_n19180_));
  OAI21_X1   g18988(.A1(new_n19180_), .A2(\asqrt[23] ), .B(new_n18940_), .ZN(new_n19181_));
  NAND2_X1   g18989(.A1(new_n19180_), .A2(\asqrt[23] ), .ZN(new_n19182_));
  NAND3_X1   g18990(.A1(new_n19181_), .A2(new_n19182_), .A3(new_n8440_), .ZN(new_n19183_));
  AOI21_X1   g18991(.A1(new_n19181_), .A2(new_n19182_), .B(new_n8440_), .ZN(new_n19184_));
  AOI21_X1   g18992(.A1(new_n18935_), .A2(new_n19183_), .B(new_n19184_), .ZN(new_n19185_));
  AOI21_X1   g18993(.A1(new_n19185_), .A2(new_n8077_), .B(new_n19177_), .ZN(new_n19186_));
  NAND2_X1   g18994(.A1(new_n19183_), .A2(new_n18935_), .ZN(new_n19187_));
  AOI21_X1   g18995(.A1(new_n19187_), .A2(new_n19168_), .B(new_n8077_), .ZN(new_n19188_));
  OAI21_X1   g18996(.A1(new_n19186_), .A2(new_n19188_), .B(\asqrt[26] ), .ZN(new_n19189_));
  AOI21_X1   g18997(.A1(new_n19176_), .A2(new_n19189_), .B(new_n7331_), .ZN(new_n19190_));
  NOR3_X1    g18998(.A1(new_n19175_), .A2(\asqrt[28] ), .A3(new_n19190_), .ZN(new_n19191_));
  OAI21_X1   g18999(.A1(new_n19175_), .A2(new_n19190_), .B(\asqrt[28] ), .ZN(new_n19192_));
  OAI21_X1   g19000(.A1(new_n18922_), .A2(new_n19191_), .B(new_n19192_), .ZN(new_n19193_));
  OAI21_X1   g19001(.A1(new_n19193_), .A2(\asqrt[29] ), .B(new_n18918_), .ZN(new_n19194_));
  NAND2_X1   g19002(.A1(new_n19193_), .A2(\asqrt[29] ), .ZN(new_n19195_));
  NAND3_X1   g19003(.A1(new_n19194_), .A2(new_n19195_), .A3(new_n6275_), .ZN(new_n19196_));
  AOI21_X1   g19004(.A1(new_n19194_), .A2(new_n19195_), .B(new_n6275_), .ZN(new_n19197_));
  AOI21_X1   g19005(.A1(new_n18916_), .A2(new_n19196_), .B(new_n19197_), .ZN(new_n19198_));
  AOI21_X1   g19006(.A1(new_n19198_), .A2(new_n5947_), .B(new_n18913_), .ZN(new_n19199_));
  NAND2_X1   g19007(.A1(new_n19196_), .A2(new_n18916_), .ZN(new_n19200_));
  INV_X1     g19008(.I(new_n18918_), .ZN(new_n19201_));
  INV_X1     g19009(.I(new_n18930_), .ZN(new_n19202_));
  NOR3_X1    g19010(.A1(new_n19186_), .A2(\asqrt[26] ), .A3(new_n19188_), .ZN(new_n19203_));
  OAI21_X1   g19011(.A1(new_n19202_), .A2(new_n19203_), .B(new_n19189_), .ZN(new_n19204_));
  OAI21_X1   g19012(.A1(new_n19204_), .A2(\asqrt[27] ), .B(new_n18926_), .ZN(new_n19205_));
  NAND2_X1   g19013(.A1(new_n19204_), .A2(\asqrt[27] ), .ZN(new_n19206_));
  NAND3_X1   g19014(.A1(new_n19205_), .A2(new_n19206_), .A3(new_n6966_), .ZN(new_n19207_));
  AOI21_X1   g19015(.A1(new_n19205_), .A2(new_n19206_), .B(new_n6966_), .ZN(new_n19208_));
  AOI21_X1   g19016(.A1(new_n18921_), .A2(new_n19207_), .B(new_n19208_), .ZN(new_n19209_));
  AOI21_X1   g19017(.A1(new_n19209_), .A2(new_n6636_), .B(new_n19201_), .ZN(new_n19210_));
  NAND2_X1   g19018(.A1(new_n19207_), .A2(new_n18921_), .ZN(new_n19211_));
  AOI21_X1   g19019(.A1(new_n19211_), .A2(new_n19192_), .B(new_n6636_), .ZN(new_n19212_));
  OAI21_X1   g19020(.A1(new_n19210_), .A2(new_n19212_), .B(\asqrt[30] ), .ZN(new_n19213_));
  AOI21_X1   g19021(.A1(new_n19200_), .A2(new_n19213_), .B(new_n5947_), .ZN(new_n19214_));
  NOR3_X1    g19022(.A1(new_n19199_), .A2(\asqrt[32] ), .A3(new_n19214_), .ZN(new_n19215_));
  OAI21_X1   g19023(.A1(new_n19199_), .A2(new_n19214_), .B(\asqrt[32] ), .ZN(new_n19216_));
  OAI21_X1   g19024(.A1(new_n18908_), .A2(new_n19215_), .B(new_n19216_), .ZN(new_n19217_));
  OAI21_X1   g19025(.A1(new_n19217_), .A2(\asqrt[33] ), .B(new_n18904_), .ZN(new_n19218_));
  NAND2_X1   g19026(.A1(new_n19217_), .A2(\asqrt[33] ), .ZN(new_n19219_));
  NAND3_X1   g19027(.A1(new_n19218_), .A2(new_n19219_), .A3(new_n5029_), .ZN(new_n19220_));
  AOI21_X1   g19028(.A1(new_n19218_), .A2(new_n19219_), .B(new_n5029_), .ZN(new_n19221_));
  AOI21_X1   g19029(.A1(new_n18902_), .A2(new_n19220_), .B(new_n19221_), .ZN(new_n19222_));
  AOI21_X1   g19030(.A1(new_n19222_), .A2(new_n4751_), .B(new_n18899_), .ZN(new_n19223_));
  NAND2_X1   g19031(.A1(new_n19220_), .A2(new_n18902_), .ZN(new_n19224_));
  INV_X1     g19032(.I(new_n18904_), .ZN(new_n19225_));
  INV_X1     g19033(.I(new_n18916_), .ZN(new_n19226_));
  NOR3_X1    g19034(.A1(new_n19210_), .A2(\asqrt[30] ), .A3(new_n19212_), .ZN(new_n19227_));
  OAI21_X1   g19035(.A1(new_n19226_), .A2(new_n19227_), .B(new_n19213_), .ZN(new_n19228_));
  OAI21_X1   g19036(.A1(new_n19228_), .A2(\asqrt[31] ), .B(new_n18912_), .ZN(new_n19229_));
  NAND2_X1   g19037(.A1(new_n19228_), .A2(\asqrt[31] ), .ZN(new_n19230_));
  NAND3_X1   g19038(.A1(new_n19229_), .A2(new_n19230_), .A3(new_n5643_), .ZN(new_n19231_));
  AOI21_X1   g19039(.A1(new_n19229_), .A2(new_n19230_), .B(new_n5643_), .ZN(new_n19232_));
  AOI21_X1   g19040(.A1(new_n18907_), .A2(new_n19231_), .B(new_n19232_), .ZN(new_n19233_));
  AOI21_X1   g19041(.A1(new_n19233_), .A2(new_n5336_), .B(new_n19225_), .ZN(new_n19234_));
  NAND2_X1   g19042(.A1(new_n19231_), .A2(new_n18907_), .ZN(new_n19235_));
  AOI21_X1   g19043(.A1(new_n19235_), .A2(new_n19216_), .B(new_n5336_), .ZN(new_n19236_));
  OAI21_X1   g19044(.A1(new_n19234_), .A2(new_n19236_), .B(\asqrt[34] ), .ZN(new_n19237_));
  AOI21_X1   g19045(.A1(new_n19224_), .A2(new_n19237_), .B(new_n4751_), .ZN(new_n19238_));
  NOR3_X1    g19046(.A1(new_n19223_), .A2(\asqrt[36] ), .A3(new_n19238_), .ZN(new_n19239_));
  OAI21_X1   g19047(.A1(new_n19223_), .A2(new_n19238_), .B(\asqrt[36] ), .ZN(new_n19240_));
  OAI21_X1   g19048(.A1(new_n18894_), .A2(new_n19239_), .B(new_n19240_), .ZN(new_n19241_));
  OAI21_X1   g19049(.A1(new_n19241_), .A2(\asqrt[37] ), .B(new_n18890_), .ZN(new_n19242_));
  NAND2_X1   g19050(.A1(new_n19241_), .A2(\asqrt[37] ), .ZN(new_n19243_));
  NAND3_X1   g19051(.A1(new_n19242_), .A2(new_n19243_), .A3(new_n3925_), .ZN(new_n19244_));
  AOI21_X1   g19052(.A1(new_n19242_), .A2(new_n19243_), .B(new_n3925_), .ZN(new_n19245_));
  AOI21_X1   g19053(.A1(new_n18888_), .A2(new_n19244_), .B(new_n19245_), .ZN(new_n19246_));
  AOI21_X1   g19054(.A1(new_n19246_), .A2(new_n3681_), .B(new_n18885_), .ZN(new_n19247_));
  NAND2_X1   g19055(.A1(new_n19244_), .A2(new_n18888_), .ZN(new_n19248_));
  INV_X1     g19056(.I(new_n18890_), .ZN(new_n19249_));
  INV_X1     g19057(.I(new_n18902_), .ZN(new_n19250_));
  NOR3_X1    g19058(.A1(new_n19234_), .A2(\asqrt[34] ), .A3(new_n19236_), .ZN(new_n19251_));
  OAI21_X1   g19059(.A1(new_n19250_), .A2(new_n19251_), .B(new_n19237_), .ZN(new_n19252_));
  OAI21_X1   g19060(.A1(new_n19252_), .A2(\asqrt[35] ), .B(new_n18898_), .ZN(new_n19253_));
  NAND2_X1   g19061(.A1(new_n19252_), .A2(\asqrt[35] ), .ZN(new_n19254_));
  NAND3_X1   g19062(.A1(new_n19253_), .A2(new_n19254_), .A3(new_n4461_), .ZN(new_n19255_));
  AOI21_X1   g19063(.A1(new_n19253_), .A2(new_n19254_), .B(new_n4461_), .ZN(new_n19256_));
  AOI21_X1   g19064(.A1(new_n18893_), .A2(new_n19255_), .B(new_n19256_), .ZN(new_n19257_));
  AOI21_X1   g19065(.A1(new_n19257_), .A2(new_n4196_), .B(new_n19249_), .ZN(new_n19258_));
  NAND2_X1   g19066(.A1(new_n19255_), .A2(new_n18893_), .ZN(new_n19259_));
  AOI21_X1   g19067(.A1(new_n19259_), .A2(new_n19240_), .B(new_n4196_), .ZN(new_n19260_));
  OAI21_X1   g19068(.A1(new_n19258_), .A2(new_n19260_), .B(\asqrt[38] ), .ZN(new_n19261_));
  AOI21_X1   g19069(.A1(new_n19248_), .A2(new_n19261_), .B(new_n3681_), .ZN(new_n19262_));
  NOR3_X1    g19070(.A1(new_n19247_), .A2(\asqrt[40] ), .A3(new_n19262_), .ZN(new_n19263_));
  OAI21_X1   g19071(.A1(new_n19247_), .A2(new_n19262_), .B(\asqrt[40] ), .ZN(new_n19264_));
  OAI21_X1   g19072(.A1(new_n18880_), .A2(new_n19263_), .B(new_n19264_), .ZN(new_n19265_));
  OAI21_X1   g19073(.A1(new_n19265_), .A2(\asqrt[41] ), .B(new_n18876_), .ZN(new_n19266_));
  NAND2_X1   g19074(.A1(new_n19265_), .A2(\asqrt[41] ), .ZN(new_n19267_));
  NAND3_X1   g19075(.A1(new_n19266_), .A2(new_n19267_), .A3(new_n2960_), .ZN(new_n19268_));
  AOI21_X1   g19076(.A1(new_n19266_), .A2(new_n19267_), .B(new_n2960_), .ZN(new_n19269_));
  AOI21_X1   g19077(.A1(new_n18874_), .A2(new_n19268_), .B(new_n19269_), .ZN(new_n19270_));
  AOI21_X1   g19078(.A1(new_n19270_), .A2(new_n2749_), .B(new_n18871_), .ZN(new_n19271_));
  NAND2_X1   g19079(.A1(new_n19268_), .A2(new_n18874_), .ZN(new_n19272_));
  INV_X1     g19080(.I(new_n18876_), .ZN(new_n19273_));
  INV_X1     g19081(.I(new_n18888_), .ZN(new_n19274_));
  NOR3_X1    g19082(.A1(new_n19258_), .A2(\asqrt[38] ), .A3(new_n19260_), .ZN(new_n19275_));
  OAI21_X1   g19083(.A1(new_n19274_), .A2(new_n19275_), .B(new_n19261_), .ZN(new_n19276_));
  OAI21_X1   g19084(.A1(new_n19276_), .A2(\asqrt[39] ), .B(new_n18884_), .ZN(new_n19277_));
  NAND2_X1   g19085(.A1(new_n19276_), .A2(\asqrt[39] ), .ZN(new_n19278_));
  NAND3_X1   g19086(.A1(new_n19277_), .A2(new_n19278_), .A3(new_n3427_), .ZN(new_n19279_));
  AOI21_X1   g19087(.A1(new_n19277_), .A2(new_n19278_), .B(new_n3427_), .ZN(new_n19280_));
  AOI21_X1   g19088(.A1(new_n18879_), .A2(new_n19279_), .B(new_n19280_), .ZN(new_n19281_));
  AOI21_X1   g19089(.A1(new_n19281_), .A2(new_n3195_), .B(new_n19273_), .ZN(new_n19282_));
  NAND2_X1   g19090(.A1(new_n19279_), .A2(new_n18879_), .ZN(new_n19283_));
  AOI21_X1   g19091(.A1(new_n19283_), .A2(new_n19264_), .B(new_n3195_), .ZN(new_n19284_));
  OAI21_X1   g19092(.A1(new_n19282_), .A2(new_n19284_), .B(\asqrt[42] ), .ZN(new_n19285_));
  AOI21_X1   g19093(.A1(new_n19272_), .A2(new_n19285_), .B(new_n2749_), .ZN(new_n19286_));
  NOR3_X1    g19094(.A1(new_n19271_), .A2(\asqrt[44] ), .A3(new_n19286_), .ZN(new_n19287_));
  OAI21_X1   g19095(.A1(new_n19271_), .A2(new_n19286_), .B(\asqrt[44] ), .ZN(new_n19288_));
  OAI21_X1   g19096(.A1(new_n18866_), .A2(new_n19287_), .B(new_n19288_), .ZN(new_n19289_));
  OAI21_X1   g19097(.A1(new_n19289_), .A2(\asqrt[45] ), .B(new_n18862_), .ZN(new_n19290_));
  NAND2_X1   g19098(.A1(new_n19289_), .A2(\asqrt[45] ), .ZN(new_n19291_));
  NAND3_X1   g19099(.A1(new_n19290_), .A2(new_n19291_), .A3(new_n2134_), .ZN(new_n19292_));
  AOI21_X1   g19100(.A1(new_n19290_), .A2(new_n19291_), .B(new_n2134_), .ZN(new_n19293_));
  AOI21_X1   g19101(.A1(new_n18860_), .A2(new_n19292_), .B(new_n19293_), .ZN(new_n19294_));
  AOI21_X1   g19102(.A1(new_n19294_), .A2(new_n1953_), .B(new_n18857_), .ZN(new_n19295_));
  NAND2_X1   g19103(.A1(new_n19292_), .A2(new_n18860_), .ZN(new_n19296_));
  INV_X1     g19104(.I(new_n18862_), .ZN(new_n19297_));
  INV_X1     g19105(.I(new_n18874_), .ZN(new_n19298_));
  NOR3_X1    g19106(.A1(new_n19282_), .A2(\asqrt[42] ), .A3(new_n19284_), .ZN(new_n19299_));
  OAI21_X1   g19107(.A1(new_n19298_), .A2(new_n19299_), .B(new_n19285_), .ZN(new_n19300_));
  OAI21_X1   g19108(.A1(new_n19300_), .A2(\asqrt[43] ), .B(new_n18870_), .ZN(new_n19301_));
  NAND2_X1   g19109(.A1(new_n19300_), .A2(\asqrt[43] ), .ZN(new_n19302_));
  NAND3_X1   g19110(.A1(new_n19301_), .A2(new_n19302_), .A3(new_n2531_), .ZN(new_n19303_));
  AOI21_X1   g19111(.A1(new_n19301_), .A2(new_n19302_), .B(new_n2531_), .ZN(new_n19304_));
  AOI21_X1   g19112(.A1(new_n18865_), .A2(new_n19303_), .B(new_n19304_), .ZN(new_n19305_));
  AOI21_X1   g19113(.A1(new_n19305_), .A2(new_n2332_), .B(new_n19297_), .ZN(new_n19306_));
  NAND2_X1   g19114(.A1(new_n19303_), .A2(new_n18865_), .ZN(new_n19307_));
  AOI21_X1   g19115(.A1(new_n19307_), .A2(new_n19288_), .B(new_n2332_), .ZN(new_n19308_));
  OAI21_X1   g19116(.A1(new_n19306_), .A2(new_n19308_), .B(\asqrt[46] ), .ZN(new_n19309_));
  AOI21_X1   g19117(.A1(new_n19296_), .A2(new_n19309_), .B(new_n1953_), .ZN(new_n19310_));
  NOR3_X1    g19118(.A1(new_n19295_), .A2(\asqrt[48] ), .A3(new_n19310_), .ZN(new_n19311_));
  OAI21_X1   g19119(.A1(new_n19295_), .A2(new_n19310_), .B(\asqrt[48] ), .ZN(new_n19312_));
  OAI21_X1   g19120(.A1(new_n18852_), .A2(new_n19311_), .B(new_n19312_), .ZN(new_n19313_));
  OAI21_X1   g19121(.A1(new_n19313_), .A2(\asqrt[49] ), .B(new_n18848_), .ZN(new_n19314_));
  NAND2_X1   g19122(.A1(new_n19313_), .A2(\asqrt[49] ), .ZN(new_n19315_));
  NAND3_X1   g19123(.A1(new_n19314_), .A2(new_n19315_), .A3(new_n1463_), .ZN(new_n19316_));
  AOI21_X1   g19124(.A1(new_n19314_), .A2(new_n19315_), .B(new_n1463_), .ZN(new_n19317_));
  AOI21_X1   g19125(.A1(new_n18846_), .A2(new_n19316_), .B(new_n19317_), .ZN(new_n19318_));
  AOI21_X1   g19126(.A1(new_n19318_), .A2(new_n1305_), .B(new_n18843_), .ZN(new_n19319_));
  NAND2_X1   g19127(.A1(new_n19316_), .A2(new_n18846_), .ZN(new_n19320_));
  INV_X1     g19128(.I(new_n18848_), .ZN(new_n19321_));
  INV_X1     g19129(.I(new_n18860_), .ZN(new_n19322_));
  NOR3_X1    g19130(.A1(new_n19306_), .A2(\asqrt[46] ), .A3(new_n19308_), .ZN(new_n19323_));
  OAI21_X1   g19131(.A1(new_n19322_), .A2(new_n19323_), .B(new_n19309_), .ZN(new_n19324_));
  OAI21_X1   g19132(.A1(new_n19324_), .A2(\asqrt[47] ), .B(new_n18856_), .ZN(new_n19325_));
  NAND2_X1   g19133(.A1(new_n19324_), .A2(\asqrt[47] ), .ZN(new_n19326_));
  NAND3_X1   g19134(.A1(new_n19325_), .A2(new_n19326_), .A3(new_n1778_), .ZN(new_n19327_));
  AOI21_X1   g19135(.A1(new_n19325_), .A2(new_n19326_), .B(new_n1778_), .ZN(new_n19328_));
  AOI21_X1   g19136(.A1(new_n18851_), .A2(new_n19327_), .B(new_n19328_), .ZN(new_n19329_));
  AOI21_X1   g19137(.A1(new_n19329_), .A2(new_n1632_), .B(new_n19321_), .ZN(new_n19330_));
  NAND2_X1   g19138(.A1(new_n19327_), .A2(new_n18851_), .ZN(new_n19331_));
  AOI21_X1   g19139(.A1(new_n19331_), .A2(new_n19312_), .B(new_n1632_), .ZN(new_n19332_));
  OAI21_X1   g19140(.A1(new_n19330_), .A2(new_n19332_), .B(\asqrt[50] ), .ZN(new_n19333_));
  AOI21_X1   g19141(.A1(new_n19320_), .A2(new_n19333_), .B(new_n1305_), .ZN(new_n19334_));
  NOR3_X1    g19142(.A1(new_n19319_), .A2(\asqrt[52] ), .A3(new_n19334_), .ZN(new_n19335_));
  OAI21_X1   g19143(.A1(new_n19319_), .A2(new_n19334_), .B(\asqrt[52] ), .ZN(new_n19336_));
  OAI21_X1   g19144(.A1(new_n18838_), .A2(new_n19335_), .B(new_n19336_), .ZN(new_n19337_));
  OAI21_X1   g19145(.A1(new_n19337_), .A2(\asqrt[53] ), .B(new_n18834_), .ZN(new_n19338_));
  NAND2_X1   g19146(.A1(new_n19337_), .A2(\asqrt[53] ), .ZN(new_n19339_));
  NAND3_X1   g19147(.A1(new_n19338_), .A2(new_n19339_), .A3(new_n860_), .ZN(new_n19340_));
  AOI21_X1   g19148(.A1(new_n19338_), .A2(new_n19339_), .B(new_n860_), .ZN(new_n19341_));
  AOI21_X1   g19149(.A1(new_n18832_), .A2(new_n19340_), .B(new_n19341_), .ZN(new_n19342_));
  AOI21_X1   g19150(.A1(new_n19342_), .A2(new_n744_), .B(new_n18829_), .ZN(new_n19343_));
  NAND2_X1   g19151(.A1(new_n19340_), .A2(new_n18832_), .ZN(new_n19344_));
  INV_X1     g19152(.I(new_n18834_), .ZN(new_n19345_));
  INV_X1     g19153(.I(new_n18846_), .ZN(new_n19346_));
  NOR3_X1    g19154(.A1(new_n19330_), .A2(\asqrt[50] ), .A3(new_n19332_), .ZN(new_n19347_));
  OAI21_X1   g19155(.A1(new_n19346_), .A2(new_n19347_), .B(new_n19333_), .ZN(new_n19348_));
  OAI21_X1   g19156(.A1(new_n19348_), .A2(\asqrt[51] ), .B(new_n18842_), .ZN(new_n19349_));
  NAND2_X1   g19157(.A1(new_n19348_), .A2(\asqrt[51] ), .ZN(new_n19350_));
  NAND3_X1   g19158(.A1(new_n19349_), .A2(new_n19350_), .A3(new_n1150_), .ZN(new_n19351_));
  AOI21_X1   g19159(.A1(new_n19349_), .A2(new_n19350_), .B(new_n1150_), .ZN(new_n19352_));
  AOI21_X1   g19160(.A1(new_n18837_), .A2(new_n19351_), .B(new_n19352_), .ZN(new_n19353_));
  AOI21_X1   g19161(.A1(new_n19353_), .A2(new_n1006_), .B(new_n19345_), .ZN(new_n19354_));
  NAND2_X1   g19162(.A1(new_n19351_), .A2(new_n18837_), .ZN(new_n19355_));
  AOI21_X1   g19163(.A1(new_n19355_), .A2(new_n19336_), .B(new_n1006_), .ZN(new_n19356_));
  OAI21_X1   g19164(.A1(new_n19354_), .A2(new_n19356_), .B(\asqrt[54] ), .ZN(new_n19357_));
  AOI21_X1   g19165(.A1(new_n19344_), .A2(new_n19357_), .B(new_n744_), .ZN(new_n19358_));
  NOR3_X1    g19166(.A1(new_n19343_), .A2(\asqrt[56] ), .A3(new_n19358_), .ZN(new_n19359_));
  OAI21_X1   g19167(.A1(new_n19343_), .A2(new_n19358_), .B(\asqrt[56] ), .ZN(new_n19360_));
  OAI21_X1   g19168(.A1(new_n18824_), .A2(new_n19359_), .B(new_n19360_), .ZN(new_n19361_));
  OAI21_X1   g19169(.A1(new_n19361_), .A2(\asqrt[57] ), .B(new_n18820_), .ZN(new_n19362_));
  NAND2_X1   g19170(.A1(new_n19361_), .A2(\asqrt[57] ), .ZN(new_n19363_));
  NAND3_X1   g19171(.A1(new_n19362_), .A2(new_n19363_), .A3(new_n423_), .ZN(new_n19364_));
  AOI21_X1   g19172(.A1(new_n19362_), .A2(new_n19363_), .B(new_n423_), .ZN(new_n19365_));
  AOI21_X1   g19173(.A1(new_n18818_), .A2(new_n19364_), .B(new_n19365_), .ZN(new_n19366_));
  AOI21_X1   g19174(.A1(new_n19366_), .A2(new_n337_), .B(new_n18816_), .ZN(new_n19367_));
  NAND2_X1   g19175(.A1(new_n19364_), .A2(new_n18818_), .ZN(new_n19368_));
  INV_X1     g19176(.I(new_n18820_), .ZN(new_n19369_));
  INV_X1     g19177(.I(new_n18832_), .ZN(new_n19370_));
  NOR3_X1    g19178(.A1(new_n19354_), .A2(\asqrt[54] ), .A3(new_n19356_), .ZN(new_n19371_));
  OAI21_X1   g19179(.A1(new_n19370_), .A2(new_n19371_), .B(new_n19357_), .ZN(new_n19372_));
  OAI21_X1   g19180(.A1(new_n19372_), .A2(\asqrt[55] ), .B(new_n18828_), .ZN(new_n19373_));
  NAND2_X1   g19181(.A1(new_n19372_), .A2(\asqrt[55] ), .ZN(new_n19374_));
  NAND3_X1   g19182(.A1(new_n19373_), .A2(new_n19374_), .A3(new_n634_), .ZN(new_n19375_));
  AOI21_X1   g19183(.A1(new_n19373_), .A2(new_n19374_), .B(new_n634_), .ZN(new_n19376_));
  AOI21_X1   g19184(.A1(new_n18823_), .A2(new_n19375_), .B(new_n19376_), .ZN(new_n19377_));
  AOI21_X1   g19185(.A1(new_n19377_), .A2(new_n531_), .B(new_n19369_), .ZN(new_n19378_));
  NAND2_X1   g19186(.A1(new_n19375_), .A2(new_n18823_), .ZN(new_n19379_));
  AOI21_X1   g19187(.A1(new_n19379_), .A2(new_n19360_), .B(new_n531_), .ZN(new_n19380_));
  OAI21_X1   g19188(.A1(new_n19378_), .A2(new_n19380_), .B(\asqrt[58] ), .ZN(new_n19381_));
  AOI21_X1   g19189(.A1(new_n19368_), .A2(new_n19381_), .B(new_n337_), .ZN(new_n19382_));
  NOR3_X1    g19190(.A1(new_n19367_), .A2(\asqrt[60] ), .A3(new_n19382_), .ZN(new_n19383_));
  NOR2_X1    g19191(.A1(new_n19383_), .A2(new_n18812_), .ZN(new_n19384_));
  INV_X1     g19192(.I(new_n18818_), .ZN(new_n19385_));
  NOR3_X1    g19193(.A1(new_n19378_), .A2(\asqrt[58] ), .A3(new_n19380_), .ZN(new_n19386_));
  OAI21_X1   g19194(.A1(new_n19385_), .A2(new_n19386_), .B(new_n19381_), .ZN(new_n19387_));
  OAI21_X1   g19195(.A1(new_n19387_), .A2(\asqrt[59] ), .B(new_n18815_), .ZN(new_n19388_));
  NAND2_X1   g19196(.A1(new_n19387_), .A2(\asqrt[59] ), .ZN(new_n19389_));
  AOI21_X1   g19197(.A1(new_n19388_), .A2(new_n19389_), .B(new_n266_), .ZN(new_n19390_));
  OAI21_X1   g19198(.A1(new_n19384_), .A2(new_n19390_), .B(\asqrt[61] ), .ZN(new_n19391_));
  OAI21_X1   g19199(.A1(new_n19367_), .A2(new_n19382_), .B(\asqrt[60] ), .ZN(new_n19392_));
  OAI21_X1   g19200(.A1(new_n18812_), .A2(new_n19383_), .B(new_n19392_), .ZN(new_n19393_));
  OAI21_X1   g19201(.A1(new_n18784_), .A2(new_n18773_), .B(new_n18802_), .ZN(new_n19394_));
  XOR2_X1    g19202(.A1(new_n19394_), .A2(new_n18780_), .Z(new_n19395_));
  OAI21_X1   g19203(.A1(new_n19393_), .A2(\asqrt[61] ), .B(new_n19395_), .ZN(new_n19396_));
  NAND2_X1   g19204(.A1(new_n19396_), .A2(new_n19391_), .ZN(new_n19397_));
  NAND3_X1   g19205(.A1(new_n19388_), .A2(new_n19389_), .A3(new_n266_), .ZN(new_n19398_));
  NAND2_X1   g19206(.A1(new_n19398_), .A2(new_n18811_), .ZN(new_n19399_));
  AOI21_X1   g19207(.A1(new_n19399_), .A2(new_n19392_), .B(new_n239_), .ZN(new_n19400_));
  AOI21_X1   g19208(.A1(new_n18811_), .A2(new_n19398_), .B(new_n19390_), .ZN(new_n19401_));
  INV_X1     g19209(.I(new_n19395_), .ZN(new_n19402_));
  AOI21_X1   g19210(.A1(new_n19401_), .A2(new_n239_), .B(new_n19402_), .ZN(new_n19403_));
  OAI21_X1   g19211(.A1(new_n19403_), .A2(new_n19400_), .B(new_n201_), .ZN(new_n19404_));
  NAND3_X1   g19212(.A1(new_n19396_), .A2(\asqrt[62] ), .A3(new_n19391_), .ZN(new_n19405_));
  OAI21_X1   g19213(.A1(new_n18772_), .A2(new_n18803_), .B(new_n18802_), .ZN(new_n19406_));
  XOR2_X1    g19214(.A1(new_n19406_), .A2(new_n18777_), .Z(new_n19407_));
  INV_X1     g19215(.I(new_n19407_), .ZN(new_n19408_));
  AOI22_X1   g19216(.A1(new_n19404_), .A2(new_n19405_), .B1(new_n19397_), .B2(new_n19408_), .ZN(new_n19409_));
  NAND2_X1   g19217(.A1(new_n18789_), .A2(new_n18259_), .ZN(new_n19410_));
  AOI21_X1   g19218(.A1(new_n18802_), .A2(new_n19410_), .B(new_n19016_), .ZN(new_n19411_));
  OAI21_X1   g19219(.A1(new_n19409_), .A2(new_n18808_), .B(new_n19411_), .ZN(new_n19412_));
  NAND2_X1   g19220(.A1(new_n18802_), .A2(new_n18259_), .ZN(new_n19413_));
  NAND2_X1   g19221(.A1(new_n19012_), .A2(new_n18259_), .ZN(new_n19414_));
  NAND2_X1   g19222(.A1(new_n18789_), .A2(new_n18799_), .ZN(new_n19415_));
  AOI21_X1   g19223(.A1(new_n19414_), .A2(new_n19415_), .B(new_n193_), .ZN(new_n19416_));
  NAND2_X1   g19224(.A1(new_n19413_), .A2(new_n19416_), .ZN(new_n19417_));
  NAND3_X1   g19225(.A1(new_n19396_), .A2(new_n201_), .A3(new_n19391_), .ZN(new_n19418_));
  AOI21_X1   g19226(.A1(new_n19396_), .A2(new_n19391_), .B(new_n201_), .ZN(new_n19419_));
  AOI21_X1   g19227(.A1(new_n19407_), .A2(new_n19418_), .B(new_n19419_), .ZN(new_n19420_));
  OAI21_X1   g19228(.A1(new_n19420_), .A2(new_n18808_), .B(new_n19417_), .ZN(new_n19421_));
  NAND3_X1   g19229(.A1(new_n19412_), .A2(new_n19421_), .A3(new_n193_), .ZN(\asqrt[1] ));
  NOR2_X1    g19230(.A1(\asqrt[1] ), .A2(new_n18808_), .ZN(new_n19423_));
  XOR2_X1    g19231(.A1(new_n19409_), .A2(new_n18807_), .Z(new_n19424_));
  NOR3_X1    g19232(.A1(new_n19423_), .A2(new_n193_), .A3(new_n19424_), .ZN(new_n19425_));
  NOR2_X1    g19233(.A1(new_n18802_), .A2(\a[4] ), .ZN(new_n19426_));
  INV_X1     g19234(.I(new_n19426_), .ZN(new_n19427_));
  NOR2_X1    g19235(.A1(new_n19039_), .A2(\a[4] ), .ZN(new_n19428_));
  AOI22_X1   g19236(.A1(new_n19427_), .A2(new_n19039_), .B1(\asqrt[2] ), .B2(new_n19428_), .ZN(new_n19429_));
  INV_X1     g19237(.I(new_n19429_), .ZN(new_n19430_));
  NAND2_X1   g19238(.A1(\asqrt[2] ), .A2(\a[4] ), .ZN(new_n19431_));
  AOI21_X1   g19239(.A1(new_n19036_), .A2(new_n19431_), .B(new_n19033_), .ZN(new_n19432_));
  NOR3_X1    g19240(.A1(\asqrt[1] ), .A2(new_n19430_), .A3(new_n19432_), .ZN(new_n19433_));
  NOR2_X1    g19241(.A1(new_n19403_), .A2(new_n19400_), .ZN(new_n19434_));
  AOI21_X1   g19242(.A1(new_n19396_), .A2(new_n19391_), .B(\asqrt[62] ), .ZN(new_n19435_));
  NOR3_X1    g19243(.A1(new_n19403_), .A2(new_n201_), .A3(new_n19400_), .ZN(new_n19436_));
  OAI22_X1   g19244(.A1(new_n19436_), .A2(new_n19435_), .B1(new_n19434_), .B2(new_n19407_), .ZN(new_n19437_));
  INV_X1     g19245(.I(new_n19411_), .ZN(new_n19438_));
  AOI21_X1   g19246(.A1(new_n19437_), .A2(new_n18807_), .B(new_n19438_), .ZN(new_n19439_));
  INV_X1     g19247(.I(new_n19417_), .ZN(new_n19440_));
  NOR3_X1    g19248(.A1(new_n19403_), .A2(\asqrt[62] ), .A3(new_n19400_), .ZN(new_n19441_));
  OAI21_X1   g19249(.A1(new_n19403_), .A2(new_n19400_), .B(\asqrt[62] ), .ZN(new_n19442_));
  OAI21_X1   g19250(.A1(new_n19408_), .A2(new_n19441_), .B(new_n19442_), .ZN(new_n19443_));
  AOI21_X1   g19251(.A1(new_n19443_), .A2(new_n18807_), .B(new_n19440_), .ZN(new_n19444_));
  NOR3_X1    g19252(.A1(new_n19439_), .A2(new_n19444_), .A3(\asqrt[63] ), .ZN(new_n19445_));
  INV_X1     g19253(.I(new_n19432_), .ZN(new_n19446_));
  AOI21_X1   g19254(.A1(new_n19445_), .A2(new_n19446_), .B(new_n19429_), .ZN(new_n19447_));
  NOR2_X1    g19255(.A1(new_n19447_), .A2(new_n19433_), .ZN(new_n19448_));
  INV_X1     g19256(.I(\a[2] ), .ZN(new_n19449_));
  OAI21_X1   g19257(.A1(\a[0] ), .A2(\a[1] ), .B(new_n19449_), .ZN(new_n19450_));
  INV_X1     g19258(.I(new_n19450_), .ZN(new_n19451_));
  NOR2_X1    g19259(.A1(new_n19440_), .A2(new_n19449_), .ZN(new_n19452_));
  INV_X1     g19260(.I(new_n19452_), .ZN(new_n19453_));
  NAND3_X1   g19261(.A1(new_n19443_), .A2(new_n18807_), .A3(new_n19453_), .ZN(new_n19454_));
  NOR3_X1    g19262(.A1(new_n19439_), .A2(new_n19454_), .A3(\asqrt[63] ), .ZN(new_n19455_));
  OAI21_X1   g19263(.A1(new_n19455_), .A2(new_n19451_), .B(\asqrt[2] ), .ZN(new_n19456_));
  NOR3_X1    g19264(.A1(new_n19420_), .A2(new_n18808_), .A3(new_n19452_), .ZN(new_n19457_));
  NAND3_X1   g19265(.A1(new_n19412_), .A2(new_n19457_), .A3(new_n193_), .ZN(new_n19458_));
  NAND3_X1   g19266(.A1(new_n19458_), .A2(new_n18802_), .A3(new_n19450_), .ZN(new_n19459_));
  NAND2_X1   g19267(.A1(\asqrt[1] ), .A2(new_n19028_), .ZN(new_n19460_));
  OAI21_X1   g19268(.A1(new_n19445_), .A2(\a[2] ), .B(\a[3] ), .ZN(new_n19461_));
  NAND2_X1   g19269(.A1(new_n19461_), .A2(new_n19460_), .ZN(new_n19462_));
  AOI22_X1   g19270(.A1(new_n19462_), .A2(\asqrt[2] ), .B1(new_n19456_), .B2(new_n19459_), .ZN(new_n19463_));
  NAND2_X1   g19271(.A1(new_n19437_), .A2(new_n18807_), .ZN(new_n19464_));
  AOI21_X1   g19272(.A1(new_n19464_), .A2(new_n19411_), .B(\asqrt[63] ), .ZN(new_n19465_));
  AOI21_X1   g19273(.A1(new_n19465_), .A2(new_n19421_), .B(new_n19029_), .ZN(new_n19466_));
  NAND2_X1   g19274(.A1(new_n19420_), .A2(new_n18808_), .ZN(new_n19467_));
  INV_X1     g19275(.I(new_n19467_), .ZN(new_n19468_));
  NAND2_X1   g19276(.A1(new_n19417_), .A2(\asqrt[2] ), .ZN(new_n19469_));
  NOR4_X1    g19277(.A1(new_n19468_), .A2(\asqrt[63] ), .A3(new_n19439_), .A4(new_n19469_), .ZN(new_n19470_));
  OAI21_X1   g19278(.A1(new_n19466_), .A2(new_n19470_), .B(new_n19031_), .ZN(new_n19471_));
  INV_X1     g19279(.I(new_n19471_), .ZN(new_n19472_));
  NOR3_X1    g19280(.A1(new_n19466_), .A2(new_n19470_), .A3(new_n19031_), .ZN(new_n19473_));
  NOR3_X1    g19281(.A1(new_n19463_), .A2(\asqrt[3] ), .A3(new_n19448_), .ZN(new_n19474_));
  OR2_X2     g19282(.A1(new_n19474_), .A2(\asqrt[4] ), .Z(new_n19475_));
  OAI21_X1   g19283(.A1(new_n19043_), .A2(new_n19064_), .B(new_n19445_), .ZN(new_n19476_));
  XOR2_X1    g19284(.A1(new_n19476_), .A2(new_n19023_), .Z(new_n19477_));
  INV_X1     g19285(.I(new_n19477_), .ZN(new_n19478_));
  NAND3_X1   g19286(.A1(new_n19458_), .A2(new_n18802_), .A3(new_n19450_), .ZN(new_n19479_));
  NAND2_X1   g19287(.A1(new_n19456_), .A2(new_n19459_), .ZN(new_n19480_));
  INV_X1     g19288(.I(\a[3] ), .ZN(new_n19481_));
  AOI21_X1   g19289(.A1(\asqrt[1] ), .A2(new_n19449_), .B(new_n19481_), .ZN(new_n19482_));
  NOR2_X1    g19290(.A1(new_n19482_), .A2(new_n19466_), .ZN(new_n19483_));
  NAND2_X1   g19291(.A1(new_n19480_), .A2(new_n19483_), .ZN(new_n19484_));
  NAND3_X1   g19292(.A1(new_n19484_), .A2(\asqrt[3] ), .A3(new_n19479_), .ZN(new_n19485_));
  NAND2_X1   g19293(.A1(new_n19463_), .A2(new_n18253_), .ZN(new_n19486_));
  NAND2_X1   g19294(.A1(new_n19486_), .A2(new_n19485_), .ZN(new_n19487_));
  NOR2_X1    g19295(.A1(new_n19470_), .A2(new_n19031_), .ZN(new_n19488_));
  NAND2_X1   g19296(.A1(new_n19488_), .A2(new_n19460_), .ZN(new_n19489_));
  NAND3_X1   g19297(.A1(new_n19489_), .A2(new_n19448_), .A3(new_n19471_), .ZN(new_n19490_));
  AOI21_X1   g19298(.A1(\asqrt[3] ), .A2(new_n19463_), .B(new_n19490_), .ZN(new_n19491_));
  AOI21_X1   g19299(.A1(new_n19487_), .A2(new_n19491_), .B(new_n19478_), .ZN(new_n19492_));
  OAI21_X1   g19300(.A1(new_n19492_), .A2(new_n19475_), .B(new_n17342_), .ZN(new_n19493_));
  NOR2_X1    g19301(.A1(new_n19045_), .A2(\asqrt[5] ), .ZN(new_n19494_));
  OAI21_X1   g19302(.A1(new_n19494_), .A2(new_n19068_), .B(new_n19445_), .ZN(new_n19495_));
  XOR2_X1    g19303(.A1(new_n19495_), .A2(new_n19053_), .Z(new_n19496_));
  INV_X1     g19304(.I(new_n19496_), .ZN(new_n19497_));
  AOI21_X1   g19305(.A1(new_n19492_), .A2(new_n19475_), .B(new_n19497_), .ZN(new_n19498_));
  OAI21_X1   g19306(.A1(new_n19498_), .A2(new_n19493_), .B(new_n16779_), .ZN(new_n19499_));
  OAI21_X1   g19307(.A1(new_n19083_), .A2(new_n19049_), .B(new_n19445_), .ZN(new_n19500_));
  XOR2_X1    g19308(.A1(new_n19500_), .A2(new_n19082_), .Z(new_n19501_));
  INV_X1     g19309(.I(new_n19501_), .ZN(new_n19502_));
  AOI21_X1   g19310(.A1(new_n19498_), .A2(new_n19493_), .B(new_n19502_), .ZN(new_n19503_));
  OAI21_X1   g19311(.A1(new_n19503_), .A2(new_n19499_), .B(new_n16269_), .ZN(new_n19504_));
  NOR2_X1    g19312(.A1(new_n19084_), .A2(\asqrt[7] ), .ZN(new_n19505_));
  OAI21_X1   g19313(.A1(new_n19505_), .A2(new_n19070_), .B(new_n19445_), .ZN(new_n19506_));
  XOR2_X1    g19314(.A1(new_n19506_), .A2(new_n18996_), .Z(new_n19507_));
  INV_X1     g19315(.I(new_n19507_), .ZN(new_n19508_));
  AOI21_X1   g19316(.A1(new_n19503_), .A2(new_n19499_), .B(new_n19508_), .ZN(new_n19509_));
  OAI21_X1   g19317(.A1(new_n19509_), .A2(new_n19504_), .B(new_n15717_), .ZN(new_n19510_));
  OAI21_X1   g19318(.A1(new_n19071_), .A2(new_n19088_), .B(new_n19445_), .ZN(new_n19511_));
  XOR2_X1    g19319(.A1(new_n19511_), .A2(new_n18992_), .Z(new_n19512_));
  INV_X1     g19320(.I(new_n19512_), .ZN(new_n19513_));
  AOI21_X1   g19321(.A1(new_n19509_), .A2(new_n19504_), .B(new_n19513_), .ZN(new_n19514_));
  OAI21_X1   g19322(.A1(new_n19514_), .A2(new_n19510_), .B(new_n15221_), .ZN(new_n19515_));
  NOR2_X1    g19323(.A1(new_n19073_), .A2(\asqrt[9] ), .ZN(new_n19516_));
  OAI21_X1   g19324(.A1(new_n19516_), .A2(new_n19092_), .B(new_n19445_), .ZN(new_n19517_));
  XOR2_X1    g19325(.A1(new_n19517_), .A2(new_n19081_), .Z(new_n19518_));
  INV_X1     g19326(.I(new_n19518_), .ZN(new_n19519_));
  AOI21_X1   g19327(.A1(new_n19514_), .A2(new_n19510_), .B(new_n19519_), .ZN(new_n19520_));
  OAI21_X1   g19328(.A1(new_n19520_), .A2(new_n19515_), .B(new_n14690_), .ZN(new_n19521_));
  OAI21_X1   g19329(.A1(new_n19107_), .A2(new_n19077_), .B(new_n19445_), .ZN(new_n19522_));
  XOR2_X1    g19330(.A1(new_n19522_), .A2(new_n19106_), .Z(new_n19523_));
  INV_X1     g19331(.I(new_n19523_), .ZN(new_n19524_));
  AOI21_X1   g19332(.A1(new_n19520_), .A2(new_n19515_), .B(new_n19524_), .ZN(new_n19525_));
  OAI21_X1   g19333(.A1(new_n19525_), .A2(new_n19521_), .B(new_n14207_), .ZN(new_n19526_));
  NOR2_X1    g19334(.A1(new_n19108_), .A2(\asqrt[11] ), .ZN(new_n19527_));
  OAI21_X1   g19335(.A1(new_n19527_), .A2(new_n19094_), .B(new_n19445_), .ZN(new_n19528_));
  XOR2_X1    g19336(.A1(new_n19528_), .A2(new_n18983_), .Z(new_n19529_));
  INV_X1     g19337(.I(new_n19529_), .ZN(new_n19530_));
  AOI21_X1   g19338(.A1(new_n19525_), .A2(new_n19521_), .B(new_n19530_), .ZN(new_n19531_));
  OAI21_X1   g19339(.A1(new_n19531_), .A2(new_n19526_), .B(new_n13690_), .ZN(new_n19532_));
  OAI21_X1   g19340(.A1(new_n19095_), .A2(new_n19112_), .B(new_n19445_), .ZN(new_n19533_));
  XOR2_X1    g19341(.A1(new_n19533_), .A2(new_n18978_), .Z(new_n19534_));
  INV_X1     g19342(.I(new_n19534_), .ZN(new_n19535_));
  AOI21_X1   g19343(.A1(new_n19531_), .A2(new_n19526_), .B(new_n19535_), .ZN(new_n19536_));
  OAI21_X1   g19344(.A1(new_n19536_), .A2(new_n19532_), .B(new_n13228_), .ZN(new_n19537_));
  NOR2_X1    g19345(.A1(new_n19097_), .A2(\asqrt[13] ), .ZN(new_n19538_));
  OAI21_X1   g19346(.A1(new_n19538_), .A2(new_n19116_), .B(new_n19445_), .ZN(new_n19539_));
  XOR2_X1    g19347(.A1(new_n19539_), .A2(new_n19105_), .Z(new_n19540_));
  INV_X1     g19348(.I(new_n19540_), .ZN(new_n19541_));
  AOI21_X1   g19349(.A1(new_n19536_), .A2(new_n19532_), .B(new_n19541_), .ZN(new_n19542_));
  OAI21_X1   g19350(.A1(new_n19542_), .A2(new_n19537_), .B(new_n12733_), .ZN(new_n19543_));
  OAI21_X1   g19351(.A1(new_n19131_), .A2(new_n19101_), .B(new_n19445_), .ZN(new_n19544_));
  XOR2_X1    g19352(.A1(new_n19544_), .A2(new_n19130_), .Z(new_n19545_));
  INV_X1     g19353(.I(new_n19545_), .ZN(new_n19546_));
  AOI21_X1   g19354(.A1(new_n19542_), .A2(new_n19537_), .B(new_n19546_), .ZN(new_n19547_));
  OAI21_X1   g19355(.A1(new_n19547_), .A2(new_n19543_), .B(new_n12283_), .ZN(new_n19548_));
  NOR2_X1    g19356(.A1(new_n19132_), .A2(\asqrt[15] ), .ZN(new_n19549_));
  OAI21_X1   g19357(.A1(new_n19549_), .A2(new_n19118_), .B(new_n19445_), .ZN(new_n19550_));
  XOR2_X1    g19358(.A1(new_n19550_), .A2(new_n18969_), .Z(new_n19551_));
  INV_X1     g19359(.I(new_n19551_), .ZN(new_n19552_));
  AOI21_X1   g19360(.A1(new_n19547_), .A2(new_n19543_), .B(new_n19552_), .ZN(new_n19553_));
  OAI21_X1   g19361(.A1(new_n19553_), .A2(new_n19548_), .B(new_n11802_), .ZN(new_n19554_));
  OAI21_X1   g19362(.A1(new_n19119_), .A2(new_n19136_), .B(new_n19445_), .ZN(new_n19555_));
  XOR2_X1    g19363(.A1(new_n19555_), .A2(new_n18964_), .Z(new_n19556_));
  INV_X1     g19364(.I(new_n19556_), .ZN(new_n19557_));
  AOI21_X1   g19365(.A1(new_n19553_), .A2(new_n19548_), .B(new_n19557_), .ZN(new_n19558_));
  OAI21_X1   g19366(.A1(new_n19558_), .A2(new_n19554_), .B(new_n11373_), .ZN(new_n19559_));
  NOR2_X1    g19367(.A1(new_n19121_), .A2(\asqrt[17] ), .ZN(new_n19560_));
  OAI21_X1   g19368(.A1(new_n19560_), .A2(new_n19140_), .B(new_n19445_), .ZN(new_n19561_));
  XOR2_X1    g19369(.A1(new_n19561_), .A2(new_n19129_), .Z(new_n19562_));
  INV_X1     g19370(.I(new_n19562_), .ZN(new_n19563_));
  AOI21_X1   g19371(.A1(new_n19558_), .A2(new_n19554_), .B(new_n19563_), .ZN(new_n19564_));
  OAI21_X1   g19372(.A1(new_n19564_), .A2(new_n19559_), .B(new_n10914_), .ZN(new_n19565_));
  OAI21_X1   g19373(.A1(new_n19155_), .A2(new_n19125_), .B(new_n19445_), .ZN(new_n19566_));
  XOR2_X1    g19374(.A1(new_n19566_), .A2(new_n19154_), .Z(new_n19567_));
  INV_X1     g19375(.I(new_n19567_), .ZN(new_n19568_));
  AOI21_X1   g19376(.A1(new_n19564_), .A2(new_n19559_), .B(new_n19568_), .ZN(new_n19569_));
  OAI21_X1   g19377(.A1(new_n19569_), .A2(new_n19565_), .B(new_n10497_), .ZN(new_n19570_));
  NOR2_X1    g19378(.A1(new_n19156_), .A2(\asqrt[19] ), .ZN(new_n19571_));
  OAI21_X1   g19379(.A1(new_n19571_), .A2(new_n19142_), .B(new_n19445_), .ZN(new_n19572_));
  XOR2_X1    g19380(.A1(new_n19572_), .A2(new_n18955_), .Z(new_n19573_));
  INV_X1     g19381(.I(new_n19573_), .ZN(new_n19574_));
  AOI21_X1   g19382(.A1(new_n19569_), .A2(new_n19565_), .B(new_n19574_), .ZN(new_n19575_));
  OAI21_X1   g19383(.A1(new_n19575_), .A2(new_n19570_), .B(new_n10052_), .ZN(new_n19576_));
  OAI21_X1   g19384(.A1(new_n19143_), .A2(new_n19160_), .B(new_n19445_), .ZN(new_n19577_));
  XOR2_X1    g19385(.A1(new_n19577_), .A2(new_n18950_), .Z(new_n19578_));
  INV_X1     g19386(.I(new_n19578_), .ZN(new_n19579_));
  AOI21_X1   g19387(.A1(new_n19575_), .A2(new_n19570_), .B(new_n19579_), .ZN(new_n19580_));
  OAI21_X1   g19388(.A1(new_n19580_), .A2(new_n19576_), .B(new_n9656_), .ZN(new_n19581_));
  NOR2_X1    g19389(.A1(new_n19145_), .A2(\asqrt[21] ), .ZN(new_n19582_));
  OAI21_X1   g19390(.A1(new_n19582_), .A2(new_n19164_), .B(new_n19445_), .ZN(new_n19583_));
  XOR2_X1    g19391(.A1(new_n19583_), .A2(new_n19153_), .Z(new_n19584_));
  INV_X1     g19392(.I(new_n19584_), .ZN(new_n19585_));
  AOI21_X1   g19393(.A1(new_n19580_), .A2(new_n19576_), .B(new_n19585_), .ZN(new_n19586_));
  OAI21_X1   g19394(.A1(new_n19586_), .A2(new_n19581_), .B(new_n9233_), .ZN(new_n19587_));
  OAI21_X1   g19395(.A1(new_n19179_), .A2(new_n19149_), .B(new_n19445_), .ZN(new_n19588_));
  XOR2_X1    g19396(.A1(new_n19588_), .A2(new_n19178_), .Z(new_n19589_));
  INV_X1     g19397(.I(new_n19589_), .ZN(new_n19590_));
  AOI21_X1   g19398(.A1(new_n19586_), .A2(new_n19581_), .B(new_n19590_), .ZN(new_n19591_));
  OAI21_X1   g19399(.A1(new_n19591_), .A2(new_n19587_), .B(new_n8849_), .ZN(new_n19592_));
  NOR2_X1    g19400(.A1(new_n19180_), .A2(\asqrt[23] ), .ZN(new_n19593_));
  OAI21_X1   g19401(.A1(new_n19593_), .A2(new_n19166_), .B(new_n19445_), .ZN(new_n19594_));
  XOR2_X1    g19402(.A1(new_n19594_), .A2(new_n18941_), .Z(new_n19595_));
  INV_X1     g19403(.I(new_n19595_), .ZN(new_n19596_));
  AOI21_X1   g19404(.A1(new_n19591_), .A2(new_n19587_), .B(new_n19596_), .ZN(new_n19597_));
  OAI21_X1   g19405(.A1(new_n19597_), .A2(new_n19592_), .B(new_n8440_), .ZN(new_n19598_));
  OAI21_X1   g19406(.A1(new_n19167_), .A2(new_n19184_), .B(new_n19445_), .ZN(new_n19599_));
  XOR2_X1    g19407(.A1(new_n19599_), .A2(new_n18936_), .Z(new_n19600_));
  INV_X1     g19408(.I(new_n19600_), .ZN(new_n19601_));
  AOI21_X1   g19409(.A1(new_n19597_), .A2(new_n19592_), .B(new_n19601_), .ZN(new_n19602_));
  OAI21_X1   g19410(.A1(new_n19602_), .A2(new_n19598_), .B(new_n8077_), .ZN(new_n19603_));
  NOR2_X1    g19411(.A1(new_n19169_), .A2(\asqrt[25] ), .ZN(new_n19604_));
  OAI21_X1   g19412(.A1(new_n19604_), .A2(new_n19188_), .B(new_n19445_), .ZN(new_n19605_));
  XOR2_X1    g19413(.A1(new_n19605_), .A2(new_n19177_), .Z(new_n19606_));
  INV_X1     g19414(.I(new_n19606_), .ZN(new_n19607_));
  AOI21_X1   g19415(.A1(new_n19602_), .A2(new_n19598_), .B(new_n19607_), .ZN(new_n19608_));
  OAI21_X1   g19416(.A1(new_n19608_), .A2(new_n19603_), .B(new_n7690_), .ZN(new_n19609_));
  OAI21_X1   g19417(.A1(new_n19203_), .A2(new_n19173_), .B(new_n19445_), .ZN(new_n19610_));
  XOR2_X1    g19418(.A1(new_n19610_), .A2(new_n19202_), .Z(new_n19611_));
  INV_X1     g19419(.I(new_n19611_), .ZN(new_n19612_));
  AOI21_X1   g19420(.A1(new_n19608_), .A2(new_n19603_), .B(new_n19612_), .ZN(new_n19613_));
  OAI21_X1   g19421(.A1(new_n19613_), .A2(new_n19609_), .B(new_n7331_), .ZN(new_n19614_));
  NOR2_X1    g19422(.A1(new_n19204_), .A2(\asqrt[27] ), .ZN(new_n19615_));
  OAI21_X1   g19423(.A1(new_n19615_), .A2(new_n19190_), .B(new_n19445_), .ZN(new_n19616_));
  XOR2_X1    g19424(.A1(new_n19616_), .A2(new_n18927_), .Z(new_n19617_));
  INV_X1     g19425(.I(new_n19617_), .ZN(new_n19618_));
  AOI21_X1   g19426(.A1(new_n19613_), .A2(new_n19609_), .B(new_n19618_), .ZN(new_n19619_));
  OAI21_X1   g19427(.A1(new_n19619_), .A2(new_n19614_), .B(new_n6966_), .ZN(new_n19620_));
  OAI21_X1   g19428(.A1(new_n19191_), .A2(new_n19208_), .B(new_n19445_), .ZN(new_n19621_));
  XOR2_X1    g19429(.A1(new_n19621_), .A2(new_n18922_), .Z(new_n19622_));
  INV_X1     g19430(.I(new_n19622_), .ZN(new_n19623_));
  AOI21_X1   g19431(.A1(new_n19619_), .A2(new_n19614_), .B(new_n19623_), .ZN(new_n19624_));
  OAI21_X1   g19432(.A1(new_n19624_), .A2(new_n19620_), .B(new_n6636_), .ZN(new_n19625_));
  NOR2_X1    g19433(.A1(new_n19193_), .A2(\asqrt[29] ), .ZN(new_n19626_));
  OAI21_X1   g19434(.A1(new_n19626_), .A2(new_n19212_), .B(new_n19445_), .ZN(new_n19627_));
  XOR2_X1    g19435(.A1(new_n19627_), .A2(new_n19201_), .Z(new_n19628_));
  INV_X1     g19436(.I(new_n19628_), .ZN(new_n19629_));
  AOI21_X1   g19437(.A1(new_n19624_), .A2(new_n19620_), .B(new_n19629_), .ZN(new_n19630_));
  OAI21_X1   g19438(.A1(new_n19630_), .A2(new_n19625_), .B(new_n6275_), .ZN(new_n19631_));
  OAI21_X1   g19439(.A1(new_n19227_), .A2(new_n19197_), .B(new_n19445_), .ZN(new_n19632_));
  XOR2_X1    g19440(.A1(new_n19632_), .A2(new_n19226_), .Z(new_n19633_));
  INV_X1     g19441(.I(new_n19633_), .ZN(new_n19634_));
  AOI21_X1   g19442(.A1(new_n19630_), .A2(new_n19625_), .B(new_n19634_), .ZN(new_n19635_));
  OAI21_X1   g19443(.A1(new_n19635_), .A2(new_n19631_), .B(new_n5947_), .ZN(new_n19636_));
  NOR2_X1    g19444(.A1(new_n19228_), .A2(\asqrt[31] ), .ZN(new_n19637_));
  OAI21_X1   g19445(.A1(new_n19637_), .A2(new_n19214_), .B(new_n19445_), .ZN(new_n19638_));
  XOR2_X1    g19446(.A1(new_n19638_), .A2(new_n18913_), .Z(new_n19639_));
  INV_X1     g19447(.I(new_n19639_), .ZN(new_n19640_));
  AOI21_X1   g19448(.A1(new_n19635_), .A2(new_n19631_), .B(new_n19640_), .ZN(new_n19641_));
  OAI21_X1   g19449(.A1(new_n19641_), .A2(new_n19636_), .B(new_n5643_), .ZN(new_n19642_));
  OAI21_X1   g19450(.A1(new_n19215_), .A2(new_n19232_), .B(new_n19445_), .ZN(new_n19643_));
  XOR2_X1    g19451(.A1(new_n19643_), .A2(new_n18908_), .Z(new_n19644_));
  INV_X1     g19452(.I(new_n19644_), .ZN(new_n19645_));
  AOI21_X1   g19453(.A1(new_n19641_), .A2(new_n19636_), .B(new_n19645_), .ZN(new_n19646_));
  OAI21_X1   g19454(.A1(new_n19646_), .A2(new_n19642_), .B(new_n5336_), .ZN(new_n19647_));
  NOR2_X1    g19455(.A1(new_n19217_), .A2(\asqrt[33] ), .ZN(new_n19648_));
  OAI21_X1   g19456(.A1(new_n19648_), .A2(new_n19236_), .B(new_n19445_), .ZN(new_n19649_));
  XOR2_X1    g19457(.A1(new_n19649_), .A2(new_n19225_), .Z(new_n19650_));
  INV_X1     g19458(.I(new_n19650_), .ZN(new_n19651_));
  AOI21_X1   g19459(.A1(new_n19646_), .A2(new_n19642_), .B(new_n19651_), .ZN(new_n19652_));
  OAI21_X1   g19460(.A1(new_n19652_), .A2(new_n19647_), .B(new_n5029_), .ZN(new_n19653_));
  OAI21_X1   g19461(.A1(new_n19251_), .A2(new_n19221_), .B(new_n19445_), .ZN(new_n19654_));
  XOR2_X1    g19462(.A1(new_n19654_), .A2(new_n19250_), .Z(new_n19655_));
  INV_X1     g19463(.I(new_n19655_), .ZN(new_n19656_));
  AOI21_X1   g19464(.A1(new_n19652_), .A2(new_n19647_), .B(new_n19656_), .ZN(new_n19657_));
  OAI21_X1   g19465(.A1(new_n19657_), .A2(new_n19653_), .B(new_n4751_), .ZN(new_n19658_));
  NOR2_X1    g19466(.A1(new_n19252_), .A2(\asqrt[35] ), .ZN(new_n19659_));
  OAI21_X1   g19467(.A1(new_n19659_), .A2(new_n19238_), .B(new_n19445_), .ZN(new_n19660_));
  XOR2_X1    g19468(.A1(new_n19660_), .A2(new_n18899_), .Z(new_n19661_));
  INV_X1     g19469(.I(new_n19661_), .ZN(new_n19662_));
  AOI21_X1   g19470(.A1(new_n19657_), .A2(new_n19653_), .B(new_n19662_), .ZN(new_n19663_));
  OAI21_X1   g19471(.A1(new_n19663_), .A2(new_n19658_), .B(new_n4461_), .ZN(new_n19664_));
  OAI21_X1   g19472(.A1(new_n19239_), .A2(new_n19256_), .B(new_n19445_), .ZN(new_n19665_));
  XOR2_X1    g19473(.A1(new_n19665_), .A2(new_n18894_), .Z(new_n19666_));
  INV_X1     g19474(.I(new_n19666_), .ZN(new_n19667_));
  AOI21_X1   g19475(.A1(new_n19663_), .A2(new_n19658_), .B(new_n19667_), .ZN(new_n19668_));
  OAI21_X1   g19476(.A1(new_n19668_), .A2(new_n19664_), .B(new_n4196_), .ZN(new_n19669_));
  NOR2_X1    g19477(.A1(new_n19241_), .A2(\asqrt[37] ), .ZN(new_n19670_));
  OAI21_X1   g19478(.A1(new_n19670_), .A2(new_n19260_), .B(new_n19445_), .ZN(new_n19671_));
  XOR2_X1    g19479(.A1(new_n19671_), .A2(new_n19249_), .Z(new_n19672_));
  INV_X1     g19480(.I(new_n19672_), .ZN(new_n19673_));
  AOI21_X1   g19481(.A1(new_n19668_), .A2(new_n19664_), .B(new_n19673_), .ZN(new_n19674_));
  OAI21_X1   g19482(.A1(new_n19674_), .A2(new_n19669_), .B(new_n3925_), .ZN(new_n19675_));
  OAI21_X1   g19483(.A1(new_n19275_), .A2(new_n19245_), .B(new_n19445_), .ZN(new_n19676_));
  XOR2_X1    g19484(.A1(new_n19676_), .A2(new_n19274_), .Z(new_n19677_));
  INV_X1     g19485(.I(new_n19677_), .ZN(new_n19678_));
  AOI21_X1   g19486(.A1(new_n19674_), .A2(new_n19669_), .B(new_n19678_), .ZN(new_n19679_));
  OAI21_X1   g19487(.A1(new_n19679_), .A2(new_n19675_), .B(new_n3681_), .ZN(new_n19680_));
  NOR2_X1    g19488(.A1(new_n19276_), .A2(\asqrt[39] ), .ZN(new_n19681_));
  OAI21_X1   g19489(.A1(new_n19681_), .A2(new_n19262_), .B(new_n19445_), .ZN(new_n19682_));
  XOR2_X1    g19490(.A1(new_n19682_), .A2(new_n18885_), .Z(new_n19683_));
  INV_X1     g19491(.I(new_n19683_), .ZN(new_n19684_));
  AOI21_X1   g19492(.A1(new_n19679_), .A2(new_n19675_), .B(new_n19684_), .ZN(new_n19685_));
  OAI21_X1   g19493(.A1(new_n19685_), .A2(new_n19680_), .B(new_n3427_), .ZN(new_n19686_));
  OAI21_X1   g19494(.A1(new_n19263_), .A2(new_n19280_), .B(new_n19445_), .ZN(new_n19687_));
  XOR2_X1    g19495(.A1(new_n19687_), .A2(new_n18880_), .Z(new_n19688_));
  INV_X1     g19496(.I(new_n19688_), .ZN(new_n19689_));
  AOI21_X1   g19497(.A1(new_n19685_), .A2(new_n19680_), .B(new_n19689_), .ZN(new_n19690_));
  OAI21_X1   g19498(.A1(new_n19690_), .A2(new_n19686_), .B(new_n3195_), .ZN(new_n19691_));
  NOR2_X1    g19499(.A1(new_n19265_), .A2(\asqrt[41] ), .ZN(new_n19692_));
  OAI21_X1   g19500(.A1(new_n19692_), .A2(new_n19284_), .B(new_n19445_), .ZN(new_n19693_));
  XOR2_X1    g19501(.A1(new_n19693_), .A2(new_n19273_), .Z(new_n19694_));
  INV_X1     g19502(.I(new_n19694_), .ZN(new_n19695_));
  AOI21_X1   g19503(.A1(new_n19690_), .A2(new_n19686_), .B(new_n19695_), .ZN(new_n19696_));
  OAI21_X1   g19504(.A1(new_n19696_), .A2(new_n19691_), .B(new_n2960_), .ZN(new_n19697_));
  OAI21_X1   g19505(.A1(new_n19299_), .A2(new_n19269_), .B(new_n19445_), .ZN(new_n19698_));
  XOR2_X1    g19506(.A1(new_n19698_), .A2(new_n19298_), .Z(new_n19699_));
  INV_X1     g19507(.I(new_n19699_), .ZN(new_n19700_));
  AOI21_X1   g19508(.A1(new_n19696_), .A2(new_n19691_), .B(new_n19700_), .ZN(new_n19701_));
  OAI21_X1   g19509(.A1(new_n19701_), .A2(new_n19697_), .B(new_n2749_), .ZN(new_n19702_));
  NOR2_X1    g19510(.A1(new_n19300_), .A2(\asqrt[43] ), .ZN(new_n19703_));
  OAI21_X1   g19511(.A1(new_n19703_), .A2(new_n19286_), .B(new_n19445_), .ZN(new_n19704_));
  XOR2_X1    g19512(.A1(new_n19704_), .A2(new_n18871_), .Z(new_n19705_));
  INV_X1     g19513(.I(new_n19705_), .ZN(new_n19706_));
  AOI21_X1   g19514(.A1(new_n19701_), .A2(new_n19697_), .B(new_n19706_), .ZN(new_n19707_));
  OAI21_X1   g19515(.A1(new_n19707_), .A2(new_n19702_), .B(new_n2531_), .ZN(new_n19708_));
  OAI21_X1   g19516(.A1(new_n19287_), .A2(new_n19304_), .B(new_n19445_), .ZN(new_n19709_));
  XOR2_X1    g19517(.A1(new_n19709_), .A2(new_n18866_), .Z(new_n19710_));
  INV_X1     g19518(.I(new_n19710_), .ZN(new_n19711_));
  AOI21_X1   g19519(.A1(new_n19707_), .A2(new_n19702_), .B(new_n19711_), .ZN(new_n19712_));
  OAI21_X1   g19520(.A1(new_n19712_), .A2(new_n19708_), .B(new_n2332_), .ZN(new_n19713_));
  NOR2_X1    g19521(.A1(new_n19289_), .A2(\asqrt[45] ), .ZN(new_n19714_));
  OAI21_X1   g19522(.A1(new_n19714_), .A2(new_n19308_), .B(new_n19445_), .ZN(new_n19715_));
  XOR2_X1    g19523(.A1(new_n19715_), .A2(new_n19297_), .Z(new_n19716_));
  INV_X1     g19524(.I(new_n19716_), .ZN(new_n19717_));
  AOI21_X1   g19525(.A1(new_n19712_), .A2(new_n19708_), .B(new_n19717_), .ZN(new_n19718_));
  OAI21_X1   g19526(.A1(new_n19718_), .A2(new_n19713_), .B(new_n2134_), .ZN(new_n19719_));
  OAI21_X1   g19527(.A1(new_n19323_), .A2(new_n19293_), .B(new_n19445_), .ZN(new_n19720_));
  XOR2_X1    g19528(.A1(new_n19720_), .A2(new_n19322_), .Z(new_n19721_));
  INV_X1     g19529(.I(new_n19721_), .ZN(new_n19722_));
  AOI21_X1   g19530(.A1(new_n19718_), .A2(new_n19713_), .B(new_n19722_), .ZN(new_n19723_));
  OAI21_X1   g19531(.A1(new_n19723_), .A2(new_n19719_), .B(new_n1953_), .ZN(new_n19724_));
  NOR2_X1    g19532(.A1(new_n19324_), .A2(\asqrt[47] ), .ZN(new_n19725_));
  OAI21_X1   g19533(.A1(new_n19725_), .A2(new_n19310_), .B(new_n19445_), .ZN(new_n19726_));
  XOR2_X1    g19534(.A1(new_n19726_), .A2(new_n18857_), .Z(new_n19727_));
  INV_X1     g19535(.I(new_n19727_), .ZN(new_n19728_));
  AOI21_X1   g19536(.A1(new_n19723_), .A2(new_n19719_), .B(new_n19728_), .ZN(new_n19729_));
  OAI21_X1   g19537(.A1(new_n19729_), .A2(new_n19724_), .B(new_n1778_), .ZN(new_n19730_));
  OAI21_X1   g19538(.A1(new_n19311_), .A2(new_n19328_), .B(new_n19445_), .ZN(new_n19731_));
  XOR2_X1    g19539(.A1(new_n19731_), .A2(new_n18852_), .Z(new_n19732_));
  INV_X1     g19540(.I(new_n19732_), .ZN(new_n19733_));
  AOI21_X1   g19541(.A1(new_n19729_), .A2(new_n19724_), .B(new_n19733_), .ZN(new_n19734_));
  OAI21_X1   g19542(.A1(new_n19734_), .A2(new_n19730_), .B(new_n1632_), .ZN(new_n19735_));
  NOR2_X1    g19543(.A1(new_n19313_), .A2(\asqrt[49] ), .ZN(new_n19736_));
  OAI21_X1   g19544(.A1(new_n19736_), .A2(new_n19332_), .B(new_n19445_), .ZN(new_n19737_));
  XOR2_X1    g19545(.A1(new_n19737_), .A2(new_n19321_), .Z(new_n19738_));
  INV_X1     g19546(.I(new_n19738_), .ZN(new_n19739_));
  AOI21_X1   g19547(.A1(new_n19734_), .A2(new_n19730_), .B(new_n19739_), .ZN(new_n19740_));
  OAI21_X1   g19548(.A1(new_n19740_), .A2(new_n19735_), .B(new_n1463_), .ZN(new_n19741_));
  OAI21_X1   g19549(.A1(new_n19347_), .A2(new_n19317_), .B(new_n19445_), .ZN(new_n19742_));
  XOR2_X1    g19550(.A1(new_n19742_), .A2(new_n19346_), .Z(new_n19743_));
  INV_X1     g19551(.I(new_n19743_), .ZN(new_n19744_));
  AOI21_X1   g19552(.A1(new_n19740_), .A2(new_n19735_), .B(new_n19744_), .ZN(new_n19745_));
  OAI21_X1   g19553(.A1(new_n19745_), .A2(new_n19741_), .B(new_n1305_), .ZN(new_n19746_));
  NOR2_X1    g19554(.A1(new_n19348_), .A2(\asqrt[51] ), .ZN(new_n19747_));
  OAI21_X1   g19555(.A1(new_n19747_), .A2(new_n19334_), .B(new_n19445_), .ZN(new_n19748_));
  XOR2_X1    g19556(.A1(new_n19748_), .A2(new_n18843_), .Z(new_n19749_));
  INV_X1     g19557(.I(new_n19749_), .ZN(new_n19750_));
  AOI21_X1   g19558(.A1(new_n19745_), .A2(new_n19741_), .B(new_n19750_), .ZN(new_n19751_));
  OAI21_X1   g19559(.A1(new_n19751_), .A2(new_n19746_), .B(new_n1150_), .ZN(new_n19752_));
  OAI21_X1   g19560(.A1(new_n19335_), .A2(new_n19352_), .B(new_n19445_), .ZN(new_n19753_));
  XOR2_X1    g19561(.A1(new_n19753_), .A2(new_n18838_), .Z(new_n19754_));
  INV_X1     g19562(.I(new_n19754_), .ZN(new_n19755_));
  AOI21_X1   g19563(.A1(new_n19751_), .A2(new_n19746_), .B(new_n19755_), .ZN(new_n19756_));
  OAI21_X1   g19564(.A1(new_n19756_), .A2(new_n19752_), .B(new_n1006_), .ZN(new_n19757_));
  NOR2_X1    g19565(.A1(new_n19337_), .A2(\asqrt[53] ), .ZN(new_n19758_));
  OAI21_X1   g19566(.A1(new_n19758_), .A2(new_n19356_), .B(new_n19445_), .ZN(new_n19759_));
  XOR2_X1    g19567(.A1(new_n19759_), .A2(new_n19345_), .Z(new_n19760_));
  INV_X1     g19568(.I(new_n19760_), .ZN(new_n19761_));
  AOI21_X1   g19569(.A1(new_n19756_), .A2(new_n19752_), .B(new_n19761_), .ZN(new_n19762_));
  OAI21_X1   g19570(.A1(new_n19762_), .A2(new_n19757_), .B(new_n860_), .ZN(new_n19763_));
  OAI21_X1   g19571(.A1(new_n19371_), .A2(new_n19341_), .B(new_n19445_), .ZN(new_n19764_));
  XOR2_X1    g19572(.A1(new_n19764_), .A2(new_n19370_), .Z(new_n19765_));
  INV_X1     g19573(.I(new_n19765_), .ZN(new_n19766_));
  AOI21_X1   g19574(.A1(new_n19762_), .A2(new_n19757_), .B(new_n19766_), .ZN(new_n19767_));
  OAI21_X1   g19575(.A1(new_n19767_), .A2(new_n19763_), .B(new_n744_), .ZN(new_n19768_));
  NOR2_X1    g19576(.A1(new_n19372_), .A2(\asqrt[55] ), .ZN(new_n19769_));
  OAI21_X1   g19577(.A1(new_n19769_), .A2(new_n19358_), .B(new_n19445_), .ZN(new_n19770_));
  XOR2_X1    g19578(.A1(new_n19770_), .A2(new_n18829_), .Z(new_n19771_));
  INV_X1     g19579(.I(new_n19771_), .ZN(new_n19772_));
  AOI21_X1   g19580(.A1(new_n19767_), .A2(new_n19763_), .B(new_n19772_), .ZN(new_n19773_));
  OAI21_X1   g19581(.A1(new_n19773_), .A2(new_n19768_), .B(new_n634_), .ZN(new_n19774_));
  OAI21_X1   g19582(.A1(new_n19359_), .A2(new_n19376_), .B(new_n19445_), .ZN(new_n19775_));
  XOR2_X1    g19583(.A1(new_n19775_), .A2(new_n18824_), .Z(new_n19776_));
  INV_X1     g19584(.I(new_n19776_), .ZN(new_n19777_));
  AOI21_X1   g19585(.A1(new_n19773_), .A2(new_n19768_), .B(new_n19777_), .ZN(new_n19778_));
  OAI21_X1   g19586(.A1(new_n19778_), .A2(new_n19774_), .B(new_n531_), .ZN(new_n19779_));
  NOR2_X1    g19587(.A1(new_n19361_), .A2(\asqrt[57] ), .ZN(new_n19780_));
  OAI21_X1   g19588(.A1(new_n19780_), .A2(new_n19380_), .B(new_n19445_), .ZN(new_n19781_));
  XOR2_X1    g19589(.A1(new_n19781_), .A2(new_n19369_), .Z(new_n19782_));
  INV_X1     g19590(.I(new_n19782_), .ZN(new_n19783_));
  AOI21_X1   g19591(.A1(new_n19778_), .A2(new_n19774_), .B(new_n19783_), .ZN(new_n19784_));
  OAI21_X1   g19592(.A1(new_n19784_), .A2(new_n19779_), .B(new_n423_), .ZN(new_n19785_));
  OAI21_X1   g19593(.A1(new_n19386_), .A2(new_n19365_), .B(new_n19445_), .ZN(new_n19786_));
  XOR2_X1    g19594(.A1(new_n19786_), .A2(new_n19385_), .Z(new_n19787_));
  INV_X1     g19595(.I(new_n19787_), .ZN(new_n19788_));
  AOI21_X1   g19596(.A1(new_n19784_), .A2(new_n19779_), .B(new_n19788_), .ZN(new_n19789_));
  OAI21_X1   g19597(.A1(new_n19789_), .A2(new_n19785_), .B(new_n337_), .ZN(new_n19790_));
  NOR2_X1    g19598(.A1(new_n19387_), .A2(\asqrt[59] ), .ZN(new_n19791_));
  OAI21_X1   g19599(.A1(new_n19791_), .A2(new_n19382_), .B(new_n19445_), .ZN(new_n19792_));
  XOR2_X1    g19600(.A1(new_n19792_), .A2(new_n18816_), .Z(new_n19793_));
  INV_X1     g19601(.I(new_n19793_), .ZN(new_n19794_));
  AOI21_X1   g19602(.A1(new_n19789_), .A2(new_n19785_), .B(new_n19794_), .ZN(new_n19795_));
  OAI21_X1   g19603(.A1(new_n19795_), .A2(new_n19790_), .B(new_n266_), .ZN(new_n19796_));
  OAI21_X1   g19604(.A1(new_n19383_), .A2(new_n19390_), .B(new_n19445_), .ZN(new_n19797_));
  XOR2_X1    g19605(.A1(new_n19797_), .A2(new_n18812_), .Z(new_n19798_));
  INV_X1     g19606(.I(new_n19798_), .ZN(new_n19799_));
  AOI21_X1   g19607(.A1(new_n19795_), .A2(new_n19790_), .B(new_n19799_), .ZN(new_n19800_));
  OAI21_X1   g19608(.A1(new_n19800_), .A2(new_n19796_), .B(new_n239_), .ZN(new_n19801_));
  NOR2_X1    g19609(.A1(new_n19393_), .A2(\asqrt[61] ), .ZN(new_n19802_));
  OAI21_X1   g19610(.A1(new_n19400_), .A2(new_n19802_), .B(new_n19445_), .ZN(new_n19803_));
  XOR2_X1    g19611(.A1(new_n19803_), .A2(new_n19402_), .Z(new_n19804_));
  INV_X1     g19612(.I(new_n19804_), .ZN(new_n19805_));
  AOI21_X1   g19613(.A1(new_n19800_), .A2(new_n19796_), .B(new_n19805_), .ZN(new_n19806_));
  OAI21_X1   g19614(.A1(new_n19806_), .A2(new_n19801_), .B(new_n201_), .ZN(new_n19807_));
  AOI21_X1   g19615(.A1(new_n19418_), .A2(new_n19442_), .B(\asqrt[1] ), .ZN(new_n19808_));
  XOR2_X1    g19616(.A1(new_n19808_), .A2(new_n19408_), .Z(new_n19809_));
  AOI21_X1   g19617(.A1(new_n19806_), .A2(new_n19801_), .B(new_n19809_), .ZN(new_n19810_));
  AOI21_X1   g19618(.A1(new_n19810_), .A2(new_n19807_), .B(new_n19425_), .ZN(new_n19811_));
  NOR2_X1    g19619(.A1(new_n19474_), .A2(\asqrt[4] ), .ZN(new_n19812_));
  NOR2_X1    g19620(.A1(new_n19463_), .A2(new_n18253_), .ZN(new_n19813_));
  AOI21_X1   g19621(.A1(new_n19484_), .A2(new_n19479_), .B(\asqrt[3] ), .ZN(new_n19814_));
  NOR2_X1    g19622(.A1(new_n19813_), .A2(new_n19814_), .ZN(new_n19815_));
  NAND2_X1   g19623(.A1(new_n19463_), .A2(\asqrt[3] ), .ZN(new_n19816_));
  NOR4_X1    g19624(.A1(new_n19472_), .A2(new_n19473_), .A3(new_n19433_), .A4(new_n19447_), .ZN(new_n19817_));
  NAND2_X1   g19625(.A1(new_n19816_), .A2(new_n19817_), .ZN(new_n19818_));
  OAI21_X1   g19626(.A1(new_n19815_), .A2(new_n19818_), .B(new_n19477_), .ZN(new_n19819_));
  AOI21_X1   g19627(.A1(new_n19819_), .A2(new_n19812_), .B(\asqrt[5] ), .ZN(new_n19820_));
  OAI21_X1   g19628(.A1(new_n19819_), .A2(new_n19812_), .B(new_n19496_), .ZN(new_n19821_));
  AOI21_X1   g19629(.A1(new_n19820_), .A2(new_n19821_), .B(\asqrt[6] ), .ZN(new_n19822_));
  OAI21_X1   g19630(.A1(new_n19820_), .A2(new_n19821_), .B(new_n19501_), .ZN(new_n19823_));
  AOI21_X1   g19631(.A1(new_n19822_), .A2(new_n19823_), .B(\asqrt[7] ), .ZN(new_n19824_));
  OAI21_X1   g19632(.A1(new_n19822_), .A2(new_n19823_), .B(new_n19507_), .ZN(new_n19825_));
  AOI21_X1   g19633(.A1(new_n19824_), .A2(new_n19825_), .B(\asqrt[8] ), .ZN(new_n19826_));
  OAI21_X1   g19634(.A1(new_n19824_), .A2(new_n19825_), .B(new_n19512_), .ZN(new_n19827_));
  AOI21_X1   g19635(.A1(new_n19826_), .A2(new_n19827_), .B(\asqrt[9] ), .ZN(new_n19828_));
  OAI21_X1   g19636(.A1(new_n19826_), .A2(new_n19827_), .B(new_n19518_), .ZN(new_n19829_));
  AOI21_X1   g19637(.A1(new_n19828_), .A2(new_n19829_), .B(\asqrt[10] ), .ZN(new_n19830_));
  OAI21_X1   g19638(.A1(new_n19828_), .A2(new_n19829_), .B(new_n19523_), .ZN(new_n19831_));
  AOI21_X1   g19639(.A1(new_n19830_), .A2(new_n19831_), .B(\asqrt[11] ), .ZN(new_n19832_));
  OAI21_X1   g19640(.A1(new_n19830_), .A2(new_n19831_), .B(new_n19529_), .ZN(new_n19833_));
  AOI21_X1   g19641(.A1(new_n19832_), .A2(new_n19833_), .B(\asqrt[12] ), .ZN(new_n19834_));
  OAI21_X1   g19642(.A1(new_n19832_), .A2(new_n19833_), .B(new_n19534_), .ZN(new_n19835_));
  AOI21_X1   g19643(.A1(new_n19834_), .A2(new_n19835_), .B(\asqrt[13] ), .ZN(new_n19836_));
  OAI21_X1   g19644(.A1(new_n19834_), .A2(new_n19835_), .B(new_n19540_), .ZN(new_n19837_));
  AOI21_X1   g19645(.A1(new_n19836_), .A2(new_n19837_), .B(\asqrt[14] ), .ZN(new_n19838_));
  OAI21_X1   g19646(.A1(new_n19836_), .A2(new_n19837_), .B(new_n19545_), .ZN(new_n19839_));
  AOI21_X1   g19647(.A1(new_n19838_), .A2(new_n19839_), .B(\asqrt[15] ), .ZN(new_n19840_));
  OAI21_X1   g19648(.A1(new_n19838_), .A2(new_n19839_), .B(new_n19551_), .ZN(new_n19841_));
  AOI21_X1   g19649(.A1(new_n19840_), .A2(new_n19841_), .B(\asqrt[16] ), .ZN(new_n19842_));
  OAI21_X1   g19650(.A1(new_n19840_), .A2(new_n19841_), .B(new_n19556_), .ZN(new_n19843_));
  AOI21_X1   g19651(.A1(new_n19842_), .A2(new_n19843_), .B(\asqrt[17] ), .ZN(new_n19844_));
  OAI21_X1   g19652(.A1(new_n19842_), .A2(new_n19843_), .B(new_n19562_), .ZN(new_n19845_));
  AOI21_X1   g19653(.A1(new_n19844_), .A2(new_n19845_), .B(\asqrt[18] ), .ZN(new_n19846_));
  OAI21_X1   g19654(.A1(new_n19844_), .A2(new_n19845_), .B(new_n19567_), .ZN(new_n19847_));
  AOI21_X1   g19655(.A1(new_n19846_), .A2(new_n19847_), .B(\asqrt[19] ), .ZN(new_n19848_));
  OAI21_X1   g19656(.A1(new_n19846_), .A2(new_n19847_), .B(new_n19573_), .ZN(new_n19849_));
  AOI21_X1   g19657(.A1(new_n19848_), .A2(new_n19849_), .B(\asqrt[20] ), .ZN(new_n19850_));
  OAI21_X1   g19658(.A1(new_n19848_), .A2(new_n19849_), .B(new_n19578_), .ZN(new_n19851_));
  AOI21_X1   g19659(.A1(new_n19850_), .A2(new_n19851_), .B(\asqrt[21] ), .ZN(new_n19852_));
  OAI21_X1   g19660(.A1(new_n19850_), .A2(new_n19851_), .B(new_n19584_), .ZN(new_n19853_));
  AOI21_X1   g19661(.A1(new_n19852_), .A2(new_n19853_), .B(\asqrt[22] ), .ZN(new_n19854_));
  OAI21_X1   g19662(.A1(new_n19852_), .A2(new_n19853_), .B(new_n19589_), .ZN(new_n19855_));
  AOI21_X1   g19663(.A1(new_n19854_), .A2(new_n19855_), .B(\asqrt[23] ), .ZN(new_n19856_));
  OAI21_X1   g19664(.A1(new_n19854_), .A2(new_n19855_), .B(new_n19595_), .ZN(new_n19857_));
  AOI21_X1   g19665(.A1(new_n19856_), .A2(new_n19857_), .B(\asqrt[24] ), .ZN(new_n19858_));
  OAI21_X1   g19666(.A1(new_n19856_), .A2(new_n19857_), .B(new_n19600_), .ZN(new_n19859_));
  AOI21_X1   g19667(.A1(new_n19858_), .A2(new_n19859_), .B(\asqrt[25] ), .ZN(new_n19860_));
  OAI21_X1   g19668(.A1(new_n19858_), .A2(new_n19859_), .B(new_n19606_), .ZN(new_n19861_));
  AOI21_X1   g19669(.A1(new_n19860_), .A2(new_n19861_), .B(\asqrt[26] ), .ZN(new_n19862_));
  OAI21_X1   g19670(.A1(new_n19860_), .A2(new_n19861_), .B(new_n19611_), .ZN(new_n19863_));
  AOI21_X1   g19671(.A1(new_n19862_), .A2(new_n19863_), .B(\asqrt[27] ), .ZN(new_n19864_));
  OAI21_X1   g19672(.A1(new_n19862_), .A2(new_n19863_), .B(new_n19617_), .ZN(new_n19865_));
  AOI21_X1   g19673(.A1(new_n19864_), .A2(new_n19865_), .B(\asqrt[28] ), .ZN(new_n19866_));
  OAI21_X1   g19674(.A1(new_n19864_), .A2(new_n19865_), .B(new_n19622_), .ZN(new_n19867_));
  AOI21_X1   g19675(.A1(new_n19866_), .A2(new_n19867_), .B(\asqrt[29] ), .ZN(new_n19868_));
  OAI21_X1   g19676(.A1(new_n19866_), .A2(new_n19867_), .B(new_n19628_), .ZN(new_n19869_));
  AOI21_X1   g19677(.A1(new_n19868_), .A2(new_n19869_), .B(\asqrt[30] ), .ZN(new_n19870_));
  OAI21_X1   g19678(.A1(new_n19868_), .A2(new_n19869_), .B(new_n19633_), .ZN(new_n19871_));
  AOI21_X1   g19679(.A1(new_n19870_), .A2(new_n19871_), .B(\asqrt[31] ), .ZN(new_n19872_));
  OAI21_X1   g19680(.A1(new_n19870_), .A2(new_n19871_), .B(new_n19639_), .ZN(new_n19873_));
  AOI21_X1   g19681(.A1(new_n19872_), .A2(new_n19873_), .B(\asqrt[32] ), .ZN(new_n19874_));
  OAI21_X1   g19682(.A1(new_n19872_), .A2(new_n19873_), .B(new_n19644_), .ZN(new_n19875_));
  AOI21_X1   g19683(.A1(new_n19874_), .A2(new_n19875_), .B(\asqrt[33] ), .ZN(new_n19876_));
  OAI21_X1   g19684(.A1(new_n19874_), .A2(new_n19875_), .B(new_n19650_), .ZN(new_n19877_));
  AOI21_X1   g19685(.A1(new_n19876_), .A2(new_n19877_), .B(\asqrt[34] ), .ZN(new_n19878_));
  OAI21_X1   g19686(.A1(new_n19876_), .A2(new_n19877_), .B(new_n19655_), .ZN(new_n19879_));
  AOI21_X1   g19687(.A1(new_n19878_), .A2(new_n19879_), .B(\asqrt[35] ), .ZN(new_n19880_));
  OAI21_X1   g19688(.A1(new_n19878_), .A2(new_n19879_), .B(new_n19661_), .ZN(new_n19881_));
  AOI21_X1   g19689(.A1(new_n19880_), .A2(new_n19881_), .B(\asqrt[36] ), .ZN(new_n19882_));
  OAI21_X1   g19690(.A1(new_n19880_), .A2(new_n19881_), .B(new_n19666_), .ZN(new_n19883_));
  AOI21_X1   g19691(.A1(new_n19882_), .A2(new_n19883_), .B(\asqrt[37] ), .ZN(new_n19884_));
  OAI21_X1   g19692(.A1(new_n19882_), .A2(new_n19883_), .B(new_n19672_), .ZN(new_n19885_));
  AOI21_X1   g19693(.A1(new_n19884_), .A2(new_n19885_), .B(\asqrt[38] ), .ZN(new_n19886_));
  OAI21_X1   g19694(.A1(new_n19884_), .A2(new_n19885_), .B(new_n19677_), .ZN(new_n19887_));
  AOI21_X1   g19695(.A1(new_n19886_), .A2(new_n19887_), .B(\asqrt[39] ), .ZN(new_n19888_));
  OAI21_X1   g19696(.A1(new_n19886_), .A2(new_n19887_), .B(new_n19683_), .ZN(new_n19889_));
  AOI21_X1   g19697(.A1(new_n19888_), .A2(new_n19889_), .B(\asqrt[40] ), .ZN(new_n19890_));
  OAI21_X1   g19698(.A1(new_n19888_), .A2(new_n19889_), .B(new_n19688_), .ZN(new_n19891_));
  AOI21_X1   g19699(.A1(new_n19890_), .A2(new_n19891_), .B(\asqrt[41] ), .ZN(new_n19892_));
  OAI21_X1   g19700(.A1(new_n19890_), .A2(new_n19891_), .B(new_n19694_), .ZN(new_n19893_));
  AOI21_X1   g19701(.A1(new_n19892_), .A2(new_n19893_), .B(\asqrt[42] ), .ZN(new_n19894_));
  OAI21_X1   g19702(.A1(new_n19892_), .A2(new_n19893_), .B(new_n19699_), .ZN(new_n19895_));
  AOI21_X1   g19703(.A1(new_n19894_), .A2(new_n19895_), .B(\asqrt[43] ), .ZN(new_n19896_));
  OAI21_X1   g19704(.A1(new_n19894_), .A2(new_n19895_), .B(new_n19705_), .ZN(new_n19897_));
  AOI21_X1   g19705(.A1(new_n19896_), .A2(new_n19897_), .B(\asqrt[44] ), .ZN(new_n19898_));
  OAI21_X1   g19706(.A1(new_n19896_), .A2(new_n19897_), .B(new_n19710_), .ZN(new_n19899_));
  AOI21_X1   g19707(.A1(new_n19898_), .A2(new_n19899_), .B(\asqrt[45] ), .ZN(new_n19900_));
  OAI21_X1   g19708(.A1(new_n19898_), .A2(new_n19899_), .B(new_n19716_), .ZN(new_n19901_));
  AOI21_X1   g19709(.A1(new_n19900_), .A2(new_n19901_), .B(\asqrt[46] ), .ZN(new_n19902_));
  OAI21_X1   g19710(.A1(new_n19900_), .A2(new_n19901_), .B(new_n19721_), .ZN(new_n19903_));
  AOI21_X1   g19711(.A1(new_n19902_), .A2(new_n19903_), .B(\asqrt[47] ), .ZN(new_n19904_));
  OAI21_X1   g19712(.A1(new_n19902_), .A2(new_n19903_), .B(new_n19727_), .ZN(new_n19905_));
  AOI21_X1   g19713(.A1(new_n19904_), .A2(new_n19905_), .B(\asqrt[48] ), .ZN(new_n19906_));
  OAI21_X1   g19714(.A1(new_n19904_), .A2(new_n19905_), .B(new_n19732_), .ZN(new_n19907_));
  AOI21_X1   g19715(.A1(new_n19906_), .A2(new_n19907_), .B(\asqrt[49] ), .ZN(new_n19908_));
  OAI21_X1   g19716(.A1(new_n19906_), .A2(new_n19907_), .B(new_n19738_), .ZN(new_n19909_));
  AOI21_X1   g19717(.A1(new_n19908_), .A2(new_n19909_), .B(\asqrt[50] ), .ZN(new_n19910_));
  OAI21_X1   g19718(.A1(new_n19908_), .A2(new_n19909_), .B(new_n19743_), .ZN(new_n19911_));
  AOI21_X1   g19719(.A1(new_n19910_), .A2(new_n19911_), .B(\asqrt[51] ), .ZN(new_n19912_));
  OAI21_X1   g19720(.A1(new_n19910_), .A2(new_n19911_), .B(new_n19749_), .ZN(new_n19913_));
  AOI21_X1   g19721(.A1(new_n19912_), .A2(new_n19913_), .B(\asqrt[52] ), .ZN(new_n19914_));
  OAI21_X1   g19722(.A1(new_n19912_), .A2(new_n19913_), .B(new_n19754_), .ZN(new_n19915_));
  AOI21_X1   g19723(.A1(new_n19914_), .A2(new_n19915_), .B(\asqrt[53] ), .ZN(new_n19916_));
  OAI21_X1   g19724(.A1(new_n19914_), .A2(new_n19915_), .B(new_n19760_), .ZN(new_n19917_));
  AOI21_X1   g19725(.A1(new_n19916_), .A2(new_n19917_), .B(\asqrt[54] ), .ZN(new_n19918_));
  OAI21_X1   g19726(.A1(new_n19916_), .A2(new_n19917_), .B(new_n19765_), .ZN(new_n19919_));
  AOI21_X1   g19727(.A1(new_n19918_), .A2(new_n19919_), .B(\asqrt[55] ), .ZN(new_n19920_));
  OAI21_X1   g19728(.A1(new_n19918_), .A2(new_n19919_), .B(new_n19771_), .ZN(new_n19921_));
  AOI21_X1   g19729(.A1(new_n19920_), .A2(new_n19921_), .B(\asqrt[56] ), .ZN(new_n19922_));
  OAI21_X1   g19730(.A1(new_n19920_), .A2(new_n19921_), .B(new_n19776_), .ZN(new_n19923_));
  AOI21_X1   g19731(.A1(new_n19922_), .A2(new_n19923_), .B(\asqrt[57] ), .ZN(new_n19924_));
  OAI21_X1   g19732(.A1(new_n19922_), .A2(new_n19923_), .B(new_n19782_), .ZN(new_n19925_));
  AOI21_X1   g19733(.A1(new_n19924_), .A2(new_n19925_), .B(\asqrt[58] ), .ZN(new_n19926_));
  OAI21_X1   g19734(.A1(new_n19924_), .A2(new_n19925_), .B(new_n19787_), .ZN(new_n19927_));
  AOI21_X1   g19735(.A1(new_n19926_), .A2(new_n19927_), .B(\asqrt[59] ), .ZN(new_n19928_));
  OAI21_X1   g19736(.A1(new_n19926_), .A2(new_n19927_), .B(new_n19793_), .ZN(new_n19929_));
  AOI21_X1   g19737(.A1(new_n19928_), .A2(new_n19929_), .B(\asqrt[60] ), .ZN(new_n19930_));
  OAI21_X1   g19738(.A1(new_n19928_), .A2(new_n19929_), .B(new_n19798_), .ZN(new_n19931_));
  AOI21_X1   g19739(.A1(new_n19930_), .A2(new_n19931_), .B(\asqrt[61] ), .ZN(new_n19932_));
  OAI21_X1   g19740(.A1(new_n19930_), .A2(new_n19931_), .B(new_n19804_), .ZN(new_n19933_));
  AOI21_X1   g19741(.A1(new_n19932_), .A2(new_n19933_), .B(\asqrt[62] ), .ZN(new_n19934_));
  AOI21_X1   g19742(.A1(new_n19445_), .A2(new_n19464_), .B(new_n19468_), .ZN(new_n19935_));
  NOR2_X1    g19743(.A1(new_n19809_), .A2(new_n19935_), .ZN(new_n19936_));
  OAI21_X1   g19744(.A1(new_n19932_), .A2(new_n19933_), .B(new_n19936_), .ZN(new_n19937_));
  OAI21_X1   g19745(.A1(new_n19934_), .A2(new_n19937_), .B(new_n193_), .ZN(new_n19938_));
  NOR2_X1    g19746(.A1(new_n19938_), .A2(new_n19811_), .ZN(\asqrt[0] ));
endmodule


