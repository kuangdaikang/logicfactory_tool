// Benchmark "sqrt" written by ABC on Mon Sep  4 17:10:25 2023

module sqrt ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] ,
    \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] , \asqrt[5] ,
    \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] , \asqrt[10] ,
    \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] , \asqrt[15] ,
    \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] , \asqrt[20] ,
    \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] , \asqrt[25] ,
    \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] , \asqrt[30] ,
    \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] , \asqrt[35] ,
    \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] , \asqrt[40] ,
    \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] , \asqrt[45] ,
    \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] , \asqrt[50] ,
    \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] , \asqrt[55] ,
    \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] , \asqrt[60] ,
    \asqrt[61] , \asqrt[62] , \asqrt[63]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] ;
  output \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] ,
    \asqrt[5] , \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] ,
    \asqrt[10] , \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] ,
    \asqrt[15] , \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] ,
    \asqrt[20] , \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] ,
    \asqrt[25] , \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] ,
    \asqrt[30] , \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] ,
    \asqrt[35] , \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] ,
    \asqrt[40] , \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] ,
    \asqrt[45] , \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] ,
    \asqrt[50] , \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] ,
    \asqrt[55] , \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] ,
    \asqrt[60] , \asqrt[61] , \asqrt[62] , \asqrt[63] ;
  wire new_n193_, new_n194_, new_n195_, new_n196_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_,
    new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_,
    new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_,
    new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_,
    new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3159_,
    new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_,
    new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_,
    new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_,
    new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_,
    new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_,
    new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_,
    new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_,
    new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_,
    new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_,
    new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_,
    new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_,
    new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_,
    new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_,
    new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_,
    new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_,
    new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_,
    new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_,
    new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_,
    new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4012_, new_n4013_, new_n4014_,
    new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_,
    new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_,
    new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_,
    new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_,
    new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_,
    new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_,
    new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_,
    new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_,
    new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_,
    new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_,
    new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_,
    new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_,
    new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_,
    new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_,
    new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_,
    new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_,
    new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_,
    new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_,
    new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_,
    new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_,
    new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_,
    new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_,
    new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_,
    new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_,
    new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_,
    new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_,
    new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_,
    new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_,
    new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_,
    new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_,
    new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_,
    new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_,
    new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_,
    new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_,
    new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_,
    new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_,
    new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_,
    new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_,
    new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_,
    new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_,
    new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_,
    new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_,
    new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_,
    new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_,
    new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_,
    new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_,
    new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_,
    new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_,
    new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_,
    new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_,
    new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_,
    new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_,
    new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_,
    new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_,
    new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_,
    new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_,
    new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_,
    new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_,
    new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_,
    new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_,
    new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_,
    new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_,
    new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_,
    new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_,
    new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_,
    new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_,
    new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_,
    new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_,
    new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_,
    new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_,
    new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_,
    new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_,
    new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_,
    new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_,
    new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_,
    new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_,
    new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_,
    new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_,
    new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_,
    new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_,
    new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_,
    new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_,
    new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_,
    new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_,
    new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_,
    new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_,
    new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_,
    new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_,
    new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_,
    new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_,
    new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_,
    new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_,
    new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_,
    new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_,
    new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_,
    new_n5627_, new_n5628_, new_n5629_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6018_,
    new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_,
    new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_,
    new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_,
    new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_,
    new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_,
    new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_,
    new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_,
    new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_,
    new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_,
    new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_,
    new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_,
    new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_,
    new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_,
    new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_,
    new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_,
    new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_,
    new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_,
    new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_,
    new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_,
    new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_,
    new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_,
    new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_,
    new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_,
    new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_,
    new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_,
    new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_,
    new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_,
    new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_,
    new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_,
    new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_,
    new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_,
    new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_,
    new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_,
    new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_,
    new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_,
    new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_,
    new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_,
    new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_,
    new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_,
    new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_,
    new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_,
    new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_,
    new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_,
    new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_,
    new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_,
    new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_,
    new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_,
    new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_,
    new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_,
    new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_,
    new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_,
    new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_,
    new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_,
    new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7170_, new_n7171_, new_n7172_, new_n7173_,
    new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_,
    new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_,
    new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_,
    new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_,
    new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_,
    new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_,
    new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_,
    new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_,
    new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_,
    new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_,
    new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_,
    new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_,
    new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_,
    new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_,
    new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_,
    new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_,
    new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_,
    new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_,
    new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_,
    new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_,
    new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_,
    new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_,
    new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7539_, new_n7540_,
    new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_,
    new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_,
    new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_,
    new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_,
    new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_,
    new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_,
    new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_,
    new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_,
    new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_,
    new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_,
    new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_,
    new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_,
    new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_,
    new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_,
    new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_,
    new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_,
    new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_,
    new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_,
    new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_,
    new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_,
    new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_,
    new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_,
    new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_,
    new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_,
    new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_,
    new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_,
    new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_,
    new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_,
    new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_,
    new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_,
    new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_,
    new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_,
    new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_,
    new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_,
    new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_,
    new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8424_,
    new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_,
    new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_,
    new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_,
    new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_,
    new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_,
    new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_,
    new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_,
    new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_,
    new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_,
    new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_,
    new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_,
    new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_,
    new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_,
    new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_,
    new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_,
    new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_,
    new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_,
    new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_,
    new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_,
    new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_,
    new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_,
    new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_,
    new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_,
    new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_,
    new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_,
    new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_,
    new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_,
    new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_,
    new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_,
    new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_,
    new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_,
    new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_,
    new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_,
    new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9272_,
    new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_,
    new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_,
    new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_,
    new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_,
    new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_,
    new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_,
    new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_,
    new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_,
    new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_,
    new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_,
    new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_,
    new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_,
    new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_,
    new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_,
    new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_,
    new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_,
    new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_,
    new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_,
    new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_,
    new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_,
    new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_,
    new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_,
    new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_,
    new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_,
    new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_,
    new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_,
    new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_,
    new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_,
    new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_,
    new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_,
    new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_,
    new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_,
    new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_,
    new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_,
    new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_,
    new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_,
    new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_,
    new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_,
    new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_,
    new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_,
    new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_,
    new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_,
    new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_,
    new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_,
    new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_,
    new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_,
    new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_,
    new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_,
    new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_,
    new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_,
    new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_,
    new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_,
    new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_,
    new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_,
    new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_,
    new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_,
    new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_,
    new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_,
    new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_,
    new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_,
    new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_,
    new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_,
    new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_,
    new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_,
    new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_,
    new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_,
    new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_,
    new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_,
    new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_,
    new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_,
    new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_,
    new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_,
    new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_,
    new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_,
    new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_,
    new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_,
    new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_,
    new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_,
    new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_,
    new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_,
    new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_,
    new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_,
    new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_,
    new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_,
    new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_,
    new_n9783_, new_n9784_, new_n9785_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_,
    new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_,
    new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_,
    new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10753_, new_n10754_, new_n10755_, new_n10756_,
    new_n10757_, new_n10758_, new_n10759_, new_n10760_, new_n10761_,
    new_n10762_, new_n10763_, new_n10764_, new_n10765_, new_n10766_,
    new_n10767_, new_n10768_, new_n10769_, new_n10770_, new_n10771_,
    new_n10772_, new_n10773_, new_n10774_, new_n10775_, new_n10776_,
    new_n10777_, new_n10778_, new_n10779_, new_n10780_, new_n10781_,
    new_n10782_, new_n10783_, new_n10784_, new_n10785_, new_n10786_,
    new_n10787_, new_n10788_, new_n10789_, new_n10790_, new_n10791_,
    new_n10792_, new_n10793_, new_n10794_, new_n10795_, new_n10796_,
    new_n10797_, new_n10798_, new_n10799_, new_n10800_, new_n10801_,
    new_n10802_, new_n10803_, new_n10804_, new_n10805_, new_n10806_,
    new_n10807_, new_n10808_, new_n10809_, new_n10810_, new_n10811_,
    new_n10812_, new_n10813_, new_n10814_, new_n10815_, new_n10816_,
    new_n10817_, new_n10818_, new_n10819_, new_n10820_, new_n10821_,
    new_n10822_, new_n10823_, new_n10824_, new_n10825_, new_n10826_,
    new_n10827_, new_n10828_, new_n10829_, new_n10830_, new_n10831_,
    new_n10832_, new_n10833_, new_n10834_, new_n10835_, new_n10836_,
    new_n10837_, new_n10838_, new_n10839_, new_n10840_, new_n10841_,
    new_n10842_, new_n10843_, new_n10844_, new_n10845_, new_n10846_,
    new_n10847_, new_n10848_, new_n10849_, new_n10850_, new_n10851_,
    new_n10852_, new_n10853_, new_n10854_, new_n10855_, new_n10856_,
    new_n10857_, new_n10858_, new_n10859_, new_n10860_, new_n10861_,
    new_n10862_, new_n10863_, new_n10864_, new_n10865_, new_n10866_,
    new_n10867_, new_n10868_, new_n10869_, new_n10870_, new_n10871_,
    new_n10872_, new_n10873_, new_n10874_, new_n10875_, new_n10876_,
    new_n10877_, new_n10878_, new_n10879_, new_n10880_, new_n10881_,
    new_n10882_, new_n10883_, new_n10884_, new_n10885_, new_n10886_,
    new_n10887_, new_n10888_, new_n10889_, new_n10890_, new_n10891_,
    new_n10892_, new_n10893_, new_n10894_, new_n10895_, new_n10896_,
    new_n10897_, new_n10898_, new_n10899_, new_n10900_, new_n10901_,
    new_n10902_, new_n10903_, new_n10904_, new_n10905_, new_n10906_,
    new_n10907_, new_n10908_, new_n10909_, new_n10910_, new_n10911_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10933_, new_n10934_, new_n10935_, new_n10936_,
    new_n10937_, new_n10938_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11025_, new_n11026_,
    new_n11027_, new_n11028_, new_n11029_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11093_, new_n11094_, new_n11095_, new_n11096_,
    new_n11097_, new_n11098_, new_n11099_, new_n11100_, new_n11101_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11126_,
    new_n11127_, new_n11128_, new_n11129_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11146_,
    new_n11147_, new_n11148_, new_n11149_, new_n11150_, new_n11151_,
    new_n11152_, new_n11153_, new_n11154_, new_n11155_, new_n11156_,
    new_n11157_, new_n11158_, new_n11159_, new_n11160_, new_n11161_,
    new_n11162_, new_n11163_, new_n11164_, new_n11165_, new_n11166_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11176_,
    new_n11177_, new_n11178_, new_n11179_, new_n11180_, new_n11181_,
    new_n11182_, new_n11183_, new_n11184_, new_n11185_, new_n11186_,
    new_n11187_, new_n11188_, new_n11189_, new_n11190_, new_n11191_,
    new_n11192_, new_n11193_, new_n11194_, new_n11195_, new_n11196_,
    new_n11197_, new_n11198_, new_n11199_, new_n11200_, new_n11201_,
    new_n11202_, new_n11203_, new_n11204_, new_n11205_, new_n11206_,
    new_n11207_, new_n11208_, new_n11209_, new_n11210_, new_n11211_,
    new_n11212_, new_n11213_, new_n11214_, new_n11215_, new_n11216_,
    new_n11217_, new_n11218_, new_n11219_, new_n11220_, new_n11221_,
    new_n11222_, new_n11223_, new_n11224_, new_n11225_, new_n11226_,
    new_n11227_, new_n11228_, new_n11229_, new_n11230_, new_n11231_,
    new_n11232_, new_n11233_, new_n11234_, new_n11235_, new_n11236_,
    new_n11237_, new_n11238_, new_n11239_, new_n11240_, new_n11241_,
    new_n11242_, new_n11243_, new_n11244_, new_n11245_, new_n11246_,
    new_n11247_, new_n11248_, new_n11249_, new_n11250_, new_n11251_,
    new_n11252_, new_n11253_, new_n11254_, new_n11255_, new_n11256_,
    new_n11257_, new_n11258_, new_n11259_, new_n11260_, new_n11261_,
    new_n11262_, new_n11263_, new_n11264_, new_n11265_, new_n11266_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11277_,
    new_n11278_, new_n11279_, new_n11280_, new_n11281_, new_n11282_,
    new_n11283_, new_n11284_, new_n11285_, new_n11286_, new_n11287_,
    new_n11288_, new_n11289_, new_n11290_, new_n11291_, new_n11292_,
    new_n11293_, new_n11294_, new_n11295_, new_n11296_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11308_, new_n11309_, new_n11310_, new_n11311_, new_n11312_,
    new_n11313_, new_n11314_, new_n11315_, new_n11316_, new_n11317_,
    new_n11318_, new_n11319_, new_n11320_, new_n11321_, new_n11322_,
    new_n11323_, new_n11324_, new_n11325_, new_n11326_, new_n11327_,
    new_n11328_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11398_, new_n11399_, new_n11400_, new_n11401_, new_n11402_,
    new_n11403_, new_n11404_, new_n11405_, new_n11406_, new_n11407_,
    new_n11408_, new_n11409_, new_n11410_, new_n11411_, new_n11412_,
    new_n11413_, new_n11414_, new_n11415_, new_n11416_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11423_, new_n11424_, new_n11425_, new_n11426_, new_n11427_,
    new_n11428_, new_n11429_, new_n11430_, new_n11431_, new_n11432_,
    new_n11433_, new_n11434_, new_n11435_, new_n11436_, new_n11437_,
    new_n11438_, new_n11439_, new_n11440_, new_n11441_, new_n11442_,
    new_n11443_, new_n11444_, new_n11445_, new_n11446_, new_n11447_,
    new_n11448_, new_n11449_, new_n11450_, new_n11451_, new_n11452_,
    new_n11453_, new_n11454_, new_n11455_, new_n11456_, new_n11457_,
    new_n11458_, new_n11459_, new_n11460_, new_n11461_, new_n11462_,
    new_n11463_, new_n11464_, new_n11465_, new_n11466_, new_n11467_,
    new_n11468_, new_n11469_, new_n11470_, new_n11471_, new_n11472_,
    new_n11473_, new_n11474_, new_n11475_, new_n11476_, new_n11477_,
    new_n11478_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11484_, new_n11485_, new_n11486_, new_n11487_,
    new_n11488_, new_n11489_, new_n11490_, new_n11491_, new_n11492_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11509_, new_n11510_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11554_, new_n11555_, new_n11556_, new_n11557_,
    new_n11558_, new_n11559_, new_n11560_, new_n11561_, new_n11562_,
    new_n11563_, new_n11564_, new_n11565_, new_n11566_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11575_, new_n11576_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11583_, new_n11584_, new_n11585_, new_n11586_, new_n11587_,
    new_n11588_, new_n11589_, new_n11590_, new_n11591_, new_n11592_,
    new_n11593_, new_n11594_, new_n11595_, new_n11596_, new_n11597_,
    new_n11598_, new_n11599_, new_n11600_, new_n11601_, new_n11602_,
    new_n11603_, new_n11604_, new_n11605_, new_n11606_, new_n11607_,
    new_n11608_, new_n11609_, new_n11610_, new_n11611_, new_n11612_,
    new_n11613_, new_n11614_, new_n11615_, new_n11616_, new_n11617_,
    new_n11618_, new_n11619_, new_n11620_, new_n11621_, new_n11622_,
    new_n11623_, new_n11624_, new_n11625_, new_n11626_, new_n11627_,
    new_n11628_, new_n11629_, new_n11630_, new_n11631_, new_n11632_,
    new_n11633_, new_n11634_, new_n11635_, new_n11636_, new_n11637_,
    new_n11638_, new_n11639_, new_n11640_, new_n11641_, new_n11642_,
    new_n11643_, new_n11644_, new_n11645_, new_n11646_, new_n11647_,
    new_n11648_, new_n11649_, new_n11650_, new_n11651_, new_n11652_,
    new_n11653_, new_n11654_, new_n11655_, new_n11656_, new_n11657_,
    new_n11658_, new_n11659_, new_n11660_, new_n11661_, new_n11662_,
    new_n11663_, new_n11664_, new_n11665_, new_n11666_, new_n11667_,
    new_n11668_, new_n11669_, new_n11670_, new_n11671_, new_n11672_,
    new_n11673_, new_n11674_, new_n11675_, new_n11676_, new_n11677_,
    new_n11678_, new_n11679_, new_n11680_, new_n11681_, new_n11682_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11689_, new_n11690_, new_n11691_, new_n11692_,
    new_n11693_, new_n11694_, new_n11695_, new_n11696_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11740_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11748_, new_n11749_, new_n11750_, new_n11751_, new_n11752_,
    new_n11753_, new_n11754_, new_n11755_, new_n11756_, new_n11757_,
    new_n11758_, new_n11759_, new_n11760_, new_n11761_, new_n11762_,
    new_n11763_, new_n11764_, new_n11765_, new_n11766_, new_n11767_,
    new_n11768_, new_n11769_, new_n11770_, new_n11771_, new_n11772_,
    new_n11773_, new_n11774_, new_n11775_, new_n11776_, new_n11777_,
    new_n11778_, new_n11779_, new_n11780_, new_n11781_, new_n11782_,
    new_n11783_, new_n11784_, new_n11785_, new_n11786_, new_n11787_,
    new_n11788_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11811_, new_n11812_, new_n11813_,
    new_n11814_, new_n11815_, new_n11816_, new_n11817_, new_n11818_,
    new_n11819_, new_n11820_, new_n11821_, new_n11822_, new_n11823_,
    new_n11824_, new_n11825_, new_n11826_, new_n11827_, new_n11828_,
    new_n11829_, new_n11830_, new_n11831_, new_n11832_, new_n11833_,
    new_n11834_, new_n11835_, new_n11836_, new_n11837_, new_n11838_,
    new_n11839_, new_n11840_, new_n11841_, new_n11842_, new_n11843_,
    new_n11844_, new_n11845_, new_n11846_, new_n11847_, new_n11848_,
    new_n11849_, new_n11850_, new_n11851_, new_n11852_, new_n11853_,
    new_n11854_, new_n11855_, new_n11856_, new_n11857_, new_n11858_,
    new_n11859_, new_n11860_, new_n11861_, new_n11862_, new_n11863_,
    new_n11864_, new_n11865_, new_n11866_, new_n11867_, new_n11868_,
    new_n11869_, new_n11870_, new_n11871_, new_n11872_, new_n11873_,
    new_n11874_, new_n11875_, new_n11876_, new_n11877_, new_n11878_,
    new_n11879_, new_n11880_, new_n11881_, new_n11882_, new_n11883_,
    new_n11884_, new_n11885_, new_n11886_, new_n11887_, new_n11888_,
    new_n11889_, new_n11890_, new_n11891_, new_n11892_, new_n11893_,
    new_n11894_, new_n11895_, new_n11896_, new_n11897_, new_n11898_,
    new_n11899_, new_n11900_, new_n11901_, new_n11902_, new_n11903_,
    new_n11904_, new_n11905_, new_n11906_, new_n11907_, new_n11908_,
    new_n11909_, new_n11910_, new_n11911_, new_n11912_, new_n11913_,
    new_n11914_, new_n11915_, new_n11916_, new_n11917_, new_n11918_,
    new_n11919_, new_n11920_, new_n11921_, new_n11922_, new_n11923_,
    new_n11924_, new_n11925_, new_n11926_, new_n11927_, new_n11928_,
    new_n11929_, new_n11930_, new_n11931_, new_n11932_, new_n11933_,
    new_n11934_, new_n11935_, new_n11936_, new_n11937_, new_n11938_,
    new_n11939_, new_n11940_, new_n11941_, new_n11942_, new_n11943_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11950_, new_n11951_, new_n11952_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11958_,
    new_n11959_, new_n11960_, new_n11961_, new_n11962_, new_n11963_,
    new_n11964_, new_n11965_, new_n11966_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12060_, new_n12061_, new_n12062_, new_n12063_,
    new_n12064_, new_n12065_, new_n12066_, new_n12067_, new_n12068_,
    new_n12069_, new_n12070_, new_n12071_, new_n12072_, new_n12073_,
    new_n12074_, new_n12075_, new_n12076_, new_n12077_, new_n12078_,
    new_n12079_, new_n12080_, new_n12081_, new_n12082_, new_n12083_,
    new_n12084_, new_n12085_, new_n12086_, new_n12087_, new_n12088_,
    new_n12089_, new_n12090_, new_n12091_, new_n12092_, new_n12093_,
    new_n12094_, new_n12095_, new_n12096_, new_n12097_, new_n12098_,
    new_n12099_, new_n12100_, new_n12101_, new_n12102_, new_n12103_,
    new_n12104_, new_n12105_, new_n12106_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12115_, new_n12116_, new_n12117_, new_n12118_,
    new_n12119_, new_n12120_, new_n12121_, new_n12122_, new_n12123_,
    new_n12124_, new_n12125_, new_n12126_, new_n12127_, new_n12128_,
    new_n12129_, new_n12130_, new_n12131_, new_n12132_, new_n12133_,
    new_n12134_, new_n12135_, new_n12136_, new_n12137_, new_n12138_,
    new_n12139_, new_n12140_, new_n12141_, new_n12142_, new_n12143_,
    new_n12144_, new_n12145_, new_n12146_, new_n12147_, new_n12148_,
    new_n12149_, new_n12150_, new_n12151_, new_n12152_, new_n12153_,
    new_n12154_, new_n12155_, new_n12156_, new_n12157_, new_n12158_,
    new_n12159_, new_n12160_, new_n12161_, new_n12162_, new_n12163_,
    new_n12164_, new_n12165_, new_n12166_, new_n12167_, new_n12168_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12173_,
    new_n12174_, new_n12175_, new_n12176_, new_n12177_, new_n12178_,
    new_n12179_, new_n12180_, new_n12181_, new_n12182_, new_n12183_,
    new_n12184_, new_n12185_, new_n12186_, new_n12187_, new_n12188_,
    new_n12189_, new_n12190_, new_n12191_, new_n12192_, new_n12193_,
    new_n12194_, new_n12195_, new_n12196_, new_n12197_, new_n12198_,
    new_n12199_, new_n12200_, new_n12201_, new_n12202_, new_n12203_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12254_, new_n12255_, new_n12256_, new_n12257_, new_n12258_,
    new_n12259_, new_n12260_, new_n12261_, new_n12262_, new_n12263_,
    new_n12264_, new_n12265_, new_n12266_, new_n12267_, new_n12268_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12280_, new_n12281_, new_n12282_, new_n12283_,
    new_n12284_, new_n12285_, new_n12286_, new_n12287_, new_n12288_,
    new_n12289_, new_n12290_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12296_, new_n12297_, new_n12298_,
    new_n12299_, new_n12300_, new_n12301_, new_n12302_, new_n12303_,
    new_n12305_, new_n12306_, new_n12307_, new_n12308_, new_n12309_,
    new_n12310_, new_n12311_, new_n12312_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12561_, new_n12562_, new_n12563_, new_n12564_,
    new_n12565_, new_n12566_, new_n12567_, new_n12568_, new_n12569_,
    new_n12570_, new_n12571_, new_n12572_, new_n12573_, new_n12574_,
    new_n12575_, new_n12576_, new_n12577_, new_n12578_, new_n12579_,
    new_n12580_, new_n12581_, new_n12582_, new_n12583_, new_n12584_,
    new_n12585_, new_n12586_, new_n12587_, new_n12588_, new_n12589_,
    new_n12590_, new_n12591_, new_n12592_, new_n12593_, new_n12594_,
    new_n12595_, new_n12596_, new_n12597_, new_n12598_, new_n12599_,
    new_n12600_, new_n12601_, new_n12602_, new_n12603_, new_n12604_,
    new_n12605_, new_n12606_, new_n12607_, new_n12608_, new_n12609_,
    new_n12610_, new_n12611_, new_n12612_, new_n12613_, new_n12614_,
    new_n12615_, new_n12616_, new_n12617_, new_n12618_, new_n12619_,
    new_n12620_, new_n12621_, new_n12622_, new_n12623_, new_n12624_,
    new_n12625_, new_n12626_, new_n12627_, new_n12628_, new_n12629_,
    new_n12630_, new_n12631_, new_n12632_, new_n12633_, new_n12634_,
    new_n12635_, new_n12636_, new_n12637_, new_n12638_, new_n12639_,
    new_n12640_, new_n12641_, new_n12642_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12649_,
    new_n12650_, new_n12651_, new_n12652_, new_n12653_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12663_, new_n12664_,
    new_n12665_, new_n12666_, new_n12667_, new_n12668_, new_n12669_,
    new_n12670_, new_n12671_, new_n12672_, new_n12673_, new_n12674_,
    new_n12675_, new_n12676_, new_n12677_, new_n12678_, new_n12679_,
    new_n12680_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12687_, new_n12688_, new_n12689_,
    new_n12690_, new_n12691_, new_n12692_, new_n12693_, new_n12694_,
    new_n12695_, new_n12696_, new_n12697_, new_n12698_, new_n12699_,
    new_n12700_, new_n12701_, new_n12702_, new_n12703_, new_n12704_,
    new_n12705_, new_n12706_, new_n12707_, new_n12708_, new_n12709_,
    new_n12710_, new_n12711_, new_n12712_, new_n12713_, new_n12714_,
    new_n12715_, new_n12716_, new_n12717_, new_n12718_, new_n12719_,
    new_n12720_, new_n12721_, new_n12722_, new_n12723_, new_n12724_,
    new_n12725_, new_n12726_, new_n12727_, new_n12728_, new_n12729_,
    new_n12730_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13428_, new_n13429_, new_n13430_, new_n13431_,
    new_n13432_, new_n13433_, new_n13434_, new_n13435_, new_n13436_,
    new_n13437_, new_n13438_, new_n13439_, new_n13440_, new_n13441_,
    new_n13442_, new_n13443_, new_n13444_, new_n13445_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13451_,
    new_n13452_, new_n13453_, new_n13454_, new_n13455_, new_n13456_,
    new_n13457_, new_n13458_, new_n13459_, new_n13460_, new_n13461_,
    new_n13462_, new_n13463_, new_n13464_, new_n13465_, new_n13466_,
    new_n13467_, new_n13468_, new_n13469_, new_n13470_, new_n13471_,
    new_n13472_, new_n13473_, new_n13474_, new_n13475_, new_n13476_,
    new_n13477_, new_n13478_, new_n13479_, new_n13480_, new_n13481_,
    new_n13482_, new_n13483_, new_n13484_, new_n13485_, new_n13486_,
    new_n13487_, new_n13488_, new_n13489_, new_n13490_, new_n13491_,
    new_n13492_, new_n13493_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13501_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13506_,
    new_n13507_, new_n13508_, new_n13509_, new_n13510_, new_n13511_,
    new_n13512_, new_n13513_, new_n13514_, new_n13515_, new_n13516_,
    new_n13517_, new_n13518_, new_n13519_, new_n13520_, new_n13521_,
    new_n13522_, new_n13523_, new_n13524_, new_n13525_, new_n13526_,
    new_n13527_, new_n13528_, new_n13529_, new_n13530_, new_n13531_,
    new_n13532_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13958_, new_n13959_, new_n13960_, new_n13961_, new_n13962_,
    new_n13963_, new_n13964_, new_n13965_, new_n13966_, new_n13967_,
    new_n13968_, new_n13969_, new_n13970_, new_n13971_, new_n13972_,
    new_n13973_, new_n13974_, new_n13975_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13998_, new_n13999_, new_n14000_, new_n14001_, new_n14002_,
    new_n14003_, new_n14004_, new_n14005_, new_n14006_, new_n14007_,
    new_n14008_, new_n14009_, new_n14010_, new_n14011_, new_n14012_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14019_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14031_, new_n14032_,
    new_n14033_, new_n14034_, new_n14035_, new_n14036_, new_n14037_,
    new_n14038_, new_n14039_, new_n14040_, new_n14041_, new_n14042_,
    new_n14043_, new_n14044_, new_n14045_, new_n14046_, new_n14047_,
    new_n14048_, new_n14049_, new_n14050_, new_n14051_, new_n14052_,
    new_n14053_, new_n14054_, new_n14055_, new_n14056_, new_n14057_,
    new_n14058_, new_n14059_, new_n14060_, new_n14061_, new_n14062_,
    new_n14063_, new_n14064_, new_n14065_, new_n14066_, new_n14067_,
    new_n14068_, new_n14069_, new_n14070_, new_n14071_, new_n14072_,
    new_n14073_, new_n14074_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14122_,
    new_n14123_, new_n14124_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14156_, new_n14157_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14170_, new_n14171_, new_n14172_,
    new_n14173_, new_n14174_, new_n14175_, new_n14176_, new_n14177_,
    new_n14178_, new_n14179_, new_n14180_, new_n14181_, new_n14182_,
    new_n14183_, new_n14184_, new_n14185_, new_n14186_, new_n14187_,
    new_n14188_, new_n14189_, new_n14190_, new_n14191_, new_n14192_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14206_, new_n14207_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14217_,
    new_n14218_, new_n14219_, new_n14220_, new_n14221_, new_n14222_,
    new_n14223_, new_n14224_, new_n14225_, new_n14226_, new_n14227_,
    new_n14228_, new_n14229_, new_n14230_, new_n14231_, new_n14232_,
    new_n14233_, new_n14234_, new_n14235_, new_n14236_, new_n14237_,
    new_n14238_, new_n14239_, new_n14240_, new_n14241_, new_n14242_,
    new_n14243_, new_n14244_, new_n14245_, new_n14246_, new_n14247_,
    new_n14248_, new_n14249_, new_n14250_, new_n14251_, new_n14252_,
    new_n14253_, new_n14254_, new_n14255_, new_n14256_, new_n14257_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14302_,
    new_n14303_, new_n14304_, new_n14305_, new_n14306_, new_n14307_,
    new_n14308_, new_n14309_, new_n14310_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14317_,
    new_n14318_, new_n14319_, new_n14320_, new_n14321_, new_n14322_,
    new_n14323_, new_n14324_, new_n14325_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14332_,
    new_n14333_, new_n14334_, new_n14335_, new_n14336_, new_n14337_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14344_, new_n14345_, new_n14346_, new_n14347_,
    new_n14348_, new_n14349_, new_n14350_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14355_, new_n14356_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14362_,
    new_n14363_, new_n14364_, new_n14365_, new_n14366_, new_n14367_,
    new_n14368_, new_n14369_, new_n14370_, new_n14371_, new_n14372_,
    new_n14373_, new_n14374_, new_n14375_, new_n14376_, new_n14377_,
    new_n14378_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14386_, new_n14387_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14393_, new_n14394_, new_n14395_, new_n14396_, new_n14397_,
    new_n14398_, new_n14399_, new_n14400_, new_n14401_, new_n14402_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14409_, new_n14410_, new_n14411_, new_n14412_,
    new_n14413_, new_n14414_, new_n14415_, new_n14416_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14422_,
    new_n14423_, new_n14424_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14545_, new_n14546_, new_n14547_,
    new_n14548_, new_n14549_, new_n14550_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14589_, new_n14590_, new_n14591_, new_n14592_, new_n14593_,
    new_n14594_, new_n14595_, new_n14596_, new_n14597_, new_n14598_,
    new_n14599_, new_n14600_, new_n14601_, new_n14602_, new_n14603_,
    new_n14604_, new_n14605_, new_n14606_, new_n14607_, new_n14608_,
    new_n14609_, new_n14610_, new_n14611_, new_n14612_, new_n14613_,
    new_n14614_, new_n14615_, new_n14616_, new_n14617_, new_n14618_,
    new_n14619_, new_n14620_, new_n14621_, new_n14622_, new_n14623_,
    new_n14624_, new_n14625_, new_n14626_, new_n14627_, new_n14628_,
    new_n14629_, new_n14630_, new_n14631_, new_n14632_, new_n14633_,
    new_n14634_, new_n14635_, new_n14636_, new_n14637_, new_n14638_,
    new_n14639_, new_n14640_, new_n14641_, new_n14642_, new_n14643_,
    new_n14644_, new_n14645_, new_n14646_, new_n14647_, new_n14648_,
    new_n14649_, new_n14650_, new_n14651_, new_n14652_, new_n14653_,
    new_n14654_, new_n14655_, new_n14656_, new_n14657_, new_n14658_,
    new_n14659_, new_n14660_, new_n14661_, new_n14662_, new_n14663_,
    new_n14664_, new_n14665_, new_n14666_, new_n14667_, new_n14668_,
    new_n14669_, new_n14670_, new_n14671_, new_n14672_, new_n14673_,
    new_n14674_, new_n14675_, new_n14676_, new_n14677_, new_n14678_,
    new_n14679_, new_n14680_, new_n14681_, new_n14682_, new_n14683_,
    new_n14684_, new_n14685_, new_n14686_, new_n14687_, new_n14688_,
    new_n14689_, new_n14690_, new_n14691_, new_n14692_, new_n14693_,
    new_n14694_, new_n14695_, new_n14696_, new_n14697_, new_n14698_,
    new_n14699_, new_n14700_, new_n14701_, new_n14702_, new_n14703_,
    new_n14704_, new_n14705_, new_n14706_, new_n14707_, new_n14708_,
    new_n14709_, new_n14710_, new_n14711_, new_n14712_, new_n14713_,
    new_n14714_, new_n14715_, new_n14716_, new_n14717_, new_n14718_,
    new_n14719_, new_n14720_, new_n14721_, new_n14722_, new_n14723_,
    new_n14724_, new_n14725_, new_n14726_, new_n14727_, new_n14728_,
    new_n14729_, new_n14730_, new_n14731_, new_n14732_, new_n14733_,
    new_n14734_, new_n14735_, new_n14736_, new_n14737_, new_n14738_,
    new_n14739_, new_n14740_, new_n14741_, new_n14742_, new_n14743_,
    new_n14744_, new_n14745_, new_n14746_, new_n14747_, new_n14748_,
    new_n14749_, new_n14750_, new_n14751_, new_n14752_, new_n14753_,
    new_n14754_, new_n14755_, new_n14756_, new_n14757_, new_n14758_,
    new_n14759_, new_n14760_, new_n14761_, new_n14762_, new_n14763_,
    new_n14764_, new_n14765_, new_n14766_, new_n14767_, new_n14768_,
    new_n14769_, new_n14770_, new_n14771_, new_n14772_, new_n14773_,
    new_n14774_, new_n14775_, new_n14776_, new_n14777_, new_n14778_,
    new_n14779_, new_n14780_, new_n14781_, new_n14782_, new_n14783_,
    new_n14784_, new_n14785_, new_n14786_, new_n14787_, new_n14788_,
    new_n14789_, new_n14790_, new_n14791_, new_n14792_, new_n14793_,
    new_n14794_, new_n14795_, new_n14796_, new_n14797_, new_n14798_,
    new_n14799_, new_n14800_, new_n14801_, new_n14802_, new_n14803_,
    new_n14804_, new_n14805_, new_n14806_, new_n14807_, new_n14808_,
    new_n14809_, new_n14810_, new_n14811_, new_n14812_, new_n14813_,
    new_n14814_, new_n14815_, new_n14816_, new_n14817_, new_n14818_,
    new_n14819_, new_n14820_, new_n14821_, new_n14822_, new_n14823_,
    new_n14824_, new_n14825_, new_n14826_, new_n14827_, new_n14828_,
    new_n14829_, new_n14830_, new_n14831_, new_n14832_, new_n14833_,
    new_n14834_, new_n14835_, new_n14836_, new_n14837_, new_n14838_,
    new_n14839_, new_n14840_, new_n14841_, new_n14842_, new_n14843_,
    new_n14844_, new_n14845_, new_n14846_, new_n14847_, new_n14848_,
    new_n14849_, new_n14850_, new_n14851_, new_n14852_, new_n14853_,
    new_n14854_, new_n14855_, new_n14856_, new_n14857_, new_n14858_,
    new_n14859_, new_n14860_, new_n14861_, new_n14862_, new_n14863_,
    new_n14864_, new_n14865_, new_n14866_, new_n14867_, new_n14868_,
    new_n14869_, new_n14870_, new_n14871_, new_n14872_, new_n14873_,
    new_n14874_, new_n14875_, new_n14876_, new_n14877_, new_n14878_,
    new_n14879_, new_n14880_, new_n14881_, new_n14882_, new_n14883_,
    new_n14884_, new_n14885_, new_n14886_, new_n14887_, new_n14888_,
    new_n14889_, new_n14890_, new_n14891_, new_n14892_, new_n14893_,
    new_n14894_, new_n14895_, new_n14896_, new_n14897_, new_n14898_,
    new_n14899_, new_n14900_, new_n14901_, new_n14902_, new_n14903_,
    new_n14904_, new_n14905_, new_n14906_, new_n14907_, new_n14908_,
    new_n14909_, new_n14910_, new_n14911_, new_n14912_, new_n14913_,
    new_n14914_, new_n14915_, new_n14916_, new_n14917_, new_n14918_,
    new_n14919_, new_n14920_, new_n14921_, new_n14922_, new_n14923_,
    new_n14924_, new_n14925_, new_n14926_, new_n14927_, new_n14928_,
    new_n14929_, new_n14930_, new_n14931_, new_n14932_, new_n14933_,
    new_n14934_, new_n14935_, new_n14936_, new_n14937_, new_n14938_,
    new_n14939_, new_n14940_, new_n14941_, new_n14942_, new_n14943_,
    new_n14944_, new_n14945_, new_n14946_, new_n14947_, new_n14948_,
    new_n14949_, new_n14950_, new_n14951_, new_n14952_, new_n14953_,
    new_n14954_, new_n14955_, new_n14956_, new_n14957_, new_n14958_,
    new_n14959_, new_n14960_, new_n14961_, new_n14962_, new_n14963_,
    new_n14964_, new_n14965_, new_n14966_, new_n14967_, new_n14968_,
    new_n14969_, new_n14970_, new_n14971_, new_n14972_, new_n14973_,
    new_n14974_, new_n14975_, new_n14976_, new_n14977_, new_n14978_,
    new_n14979_, new_n14980_, new_n14981_, new_n14982_, new_n14983_,
    new_n14984_, new_n14985_, new_n14986_, new_n14987_, new_n14988_,
    new_n14989_, new_n14990_, new_n14991_, new_n14992_, new_n14993_,
    new_n14994_, new_n14995_, new_n14996_, new_n14997_, new_n14998_,
    new_n14999_, new_n15000_, new_n15001_, new_n15002_, new_n15003_,
    new_n15004_, new_n15005_, new_n15006_, new_n15007_, new_n15008_,
    new_n15009_, new_n15010_, new_n15011_, new_n15012_, new_n15013_,
    new_n15014_, new_n15015_, new_n15016_, new_n15017_, new_n15018_,
    new_n15019_, new_n15020_, new_n15021_, new_n15022_, new_n15023_,
    new_n15024_, new_n15025_, new_n15026_, new_n15027_, new_n15028_,
    new_n15029_, new_n15030_, new_n15031_, new_n15032_, new_n15033_,
    new_n15034_, new_n15035_, new_n15036_, new_n15037_, new_n15038_,
    new_n15039_, new_n15040_, new_n15041_, new_n15042_, new_n15043_,
    new_n15044_, new_n15045_, new_n15046_, new_n15047_, new_n15048_,
    new_n15049_, new_n15050_, new_n15051_, new_n15052_, new_n15053_,
    new_n15054_, new_n15055_, new_n15056_, new_n15057_, new_n15058_,
    new_n15059_, new_n15060_, new_n15061_, new_n15062_, new_n15063_,
    new_n15064_, new_n15065_, new_n15066_, new_n15067_, new_n15068_,
    new_n15069_, new_n15070_, new_n15071_, new_n15072_, new_n15073_,
    new_n15074_, new_n15075_, new_n15076_, new_n15077_, new_n15078_,
    new_n15079_, new_n15080_, new_n15081_, new_n15082_, new_n15083_,
    new_n15084_, new_n15085_, new_n15086_, new_n15087_, new_n15088_,
    new_n15089_, new_n15090_, new_n15091_, new_n15092_, new_n15093_,
    new_n15094_, new_n15095_, new_n15096_, new_n15097_, new_n15098_,
    new_n15099_, new_n15100_, new_n15101_, new_n15102_, new_n15103_,
    new_n15104_, new_n15105_, new_n15106_, new_n15107_, new_n15108_,
    new_n15109_, new_n15110_, new_n15111_, new_n15112_, new_n15113_,
    new_n15114_, new_n15115_, new_n15116_, new_n15117_, new_n15118_,
    new_n15119_, new_n15120_, new_n15121_, new_n15122_, new_n15123_,
    new_n15124_, new_n15125_, new_n15126_, new_n15127_, new_n15128_,
    new_n15129_, new_n15130_, new_n15131_, new_n15132_, new_n15133_,
    new_n15134_, new_n15135_, new_n15136_, new_n15137_, new_n15138_,
    new_n15139_, new_n15140_, new_n15142_, new_n15143_, new_n15144_,
    new_n15145_, new_n15146_, new_n15147_, new_n15148_, new_n15149_,
    new_n15150_, new_n15151_, new_n15152_, new_n15153_, new_n15154_,
    new_n15155_, new_n15156_, new_n15157_, new_n15158_, new_n15159_,
    new_n15160_, new_n15161_, new_n15162_, new_n15163_, new_n15164_,
    new_n15165_, new_n15166_, new_n15167_, new_n15168_, new_n15169_,
    new_n15170_, new_n15171_, new_n15172_, new_n15173_, new_n15174_,
    new_n15175_, new_n15176_, new_n15177_, new_n15178_, new_n15179_,
    new_n15180_, new_n15181_, new_n15182_, new_n15183_, new_n15184_,
    new_n15185_, new_n15186_, new_n15187_, new_n15188_, new_n15189_,
    new_n15190_, new_n15191_, new_n15192_, new_n15193_, new_n15194_,
    new_n15195_, new_n15196_, new_n15197_, new_n15198_, new_n15199_,
    new_n15200_, new_n15201_, new_n15202_, new_n15203_, new_n15204_,
    new_n15205_, new_n15206_, new_n15207_, new_n15208_, new_n15209_,
    new_n15210_, new_n15211_, new_n15212_, new_n15213_, new_n15214_,
    new_n15215_, new_n15216_, new_n15217_, new_n15218_, new_n15219_,
    new_n15220_, new_n15221_, new_n15222_, new_n15223_, new_n15224_,
    new_n15225_, new_n15226_, new_n15227_, new_n15228_, new_n15229_,
    new_n15230_, new_n15231_, new_n15232_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15369_,
    new_n15370_, new_n15371_, new_n15372_, new_n15373_, new_n15374_,
    new_n15375_, new_n15376_, new_n15377_, new_n15378_, new_n15379_,
    new_n15380_, new_n15381_, new_n15382_, new_n15383_, new_n15384_,
    new_n15385_, new_n15386_, new_n15387_, new_n15388_, new_n15389_,
    new_n15390_, new_n15391_, new_n15392_, new_n15393_, new_n15394_,
    new_n15395_, new_n15396_, new_n15397_, new_n15398_, new_n15399_,
    new_n15400_, new_n15401_, new_n15402_, new_n15403_, new_n15404_,
    new_n15405_, new_n15406_, new_n15407_, new_n15408_, new_n15409_,
    new_n15410_, new_n15411_, new_n15412_, new_n15413_, new_n15414_,
    new_n15415_, new_n15416_, new_n15417_, new_n15418_, new_n15419_,
    new_n15420_, new_n15421_, new_n15422_, new_n15423_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15428_, new_n15429_,
    new_n15430_, new_n15431_, new_n15432_, new_n15433_, new_n15434_,
    new_n15435_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15469_,
    new_n15470_, new_n15471_, new_n15472_, new_n15473_, new_n15474_,
    new_n15475_, new_n15476_, new_n15477_, new_n15478_, new_n15479_,
    new_n15480_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15488_, new_n15489_,
    new_n15490_, new_n15491_, new_n15492_, new_n15493_, new_n15494_,
    new_n15495_, new_n15496_, new_n15497_, new_n15498_, new_n15499_,
    new_n15500_, new_n15501_, new_n15502_, new_n15503_, new_n15504_,
    new_n15505_, new_n15506_, new_n15507_, new_n15508_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15575_, new_n15576_, new_n15577_, new_n15578_, new_n15579_,
    new_n15580_, new_n15581_, new_n15582_, new_n15583_, new_n15584_,
    new_n15585_, new_n15586_, new_n15587_, new_n15588_, new_n15589_,
    new_n15590_, new_n15591_, new_n15592_, new_n15593_, new_n15594_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15601_, new_n15602_, new_n15603_, new_n15604_,
    new_n15605_, new_n15606_, new_n15607_, new_n15608_, new_n15609_,
    new_n15610_, new_n15611_, new_n15612_, new_n15613_, new_n15614_,
    new_n15615_, new_n15616_, new_n15617_, new_n15618_, new_n15619_,
    new_n15620_, new_n15621_, new_n15622_, new_n15623_, new_n15624_,
    new_n15625_, new_n15626_, new_n15627_, new_n15628_, new_n15629_,
    new_n15630_, new_n15631_, new_n15632_, new_n15633_, new_n15634_,
    new_n15635_, new_n15636_, new_n15637_, new_n15638_, new_n15639_,
    new_n15640_, new_n15641_, new_n15642_, new_n15643_, new_n15644_,
    new_n15645_, new_n15646_, new_n15647_, new_n15648_, new_n15649_,
    new_n15650_, new_n15651_, new_n15652_, new_n15653_, new_n15654_,
    new_n15655_, new_n15656_, new_n15657_, new_n15658_, new_n15659_,
    new_n15660_, new_n15661_, new_n15662_, new_n15663_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15674_,
    new_n15675_, new_n15676_, new_n15677_, new_n15678_, new_n15679_,
    new_n15680_, new_n15681_, new_n15682_, new_n15683_, new_n15684_,
    new_n15685_, new_n15686_, new_n15687_, new_n15688_, new_n15689_,
    new_n15690_, new_n15691_, new_n15692_, new_n15693_, new_n15694_,
    new_n15695_, new_n15696_, new_n15697_, new_n15698_, new_n15699_,
    new_n15700_, new_n15701_, new_n15702_, new_n15703_, new_n15704_,
    new_n15705_, new_n15706_, new_n15707_, new_n15708_, new_n15709_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16181_, new_n16182_, new_n16183_, new_n16184_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16192_, new_n16193_, new_n16194_, new_n16195_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16340_, new_n16341_,
    new_n16342_, new_n16343_, new_n16344_, new_n16345_, new_n16346_,
    new_n16347_, new_n16348_, new_n16349_, new_n16350_, new_n16351_,
    new_n16352_, new_n16353_, new_n16354_, new_n16355_, new_n16356_,
    new_n16357_, new_n16358_, new_n16359_, new_n16360_, new_n16361_,
    new_n16362_, new_n16363_, new_n16364_, new_n16365_, new_n16366_,
    new_n16367_, new_n16368_, new_n16369_, new_n16370_, new_n16371_,
    new_n16372_, new_n16373_, new_n16374_, new_n16375_, new_n16376_,
    new_n16377_, new_n16378_, new_n16379_, new_n16380_, new_n16381_,
    new_n16382_, new_n16383_, new_n16384_, new_n16385_, new_n16386_,
    new_n16387_, new_n16388_, new_n16389_, new_n16390_, new_n16391_,
    new_n16392_, new_n16393_, new_n16394_, new_n16395_, new_n16396_,
    new_n16397_, new_n16398_, new_n16399_, new_n16400_, new_n16401_,
    new_n16402_, new_n16403_, new_n16404_, new_n16405_, new_n16406_,
    new_n16407_, new_n16408_, new_n16409_, new_n16410_, new_n16411_,
    new_n16412_, new_n16413_, new_n16414_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16426_,
    new_n16427_, new_n16428_, new_n16429_, new_n16430_, new_n16431_,
    new_n16432_, new_n16433_, new_n16434_, new_n16435_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16458_, new_n16459_, new_n16460_, new_n16461_,
    new_n16462_, new_n16463_, new_n16464_, new_n16465_, new_n16466_,
    new_n16467_, new_n16468_, new_n16469_, new_n16470_, new_n16471_,
    new_n16472_, new_n16473_, new_n16474_, new_n16475_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16490_, new_n16491_,
    new_n16492_, new_n16493_, new_n16494_, new_n16495_, new_n16496_,
    new_n16497_, new_n16498_, new_n16499_, new_n16500_, new_n16501_,
    new_n16502_, new_n16503_, new_n16504_, new_n16505_, new_n16506_,
    new_n16507_, new_n16508_, new_n16509_, new_n16510_, new_n16511_,
    new_n16512_, new_n16513_, new_n16514_, new_n16515_, new_n16516_,
    new_n16517_, new_n16518_, new_n16519_, new_n16520_, new_n16521_,
    new_n16522_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16530_, new_n16531_,
    new_n16532_, new_n16533_, new_n16534_, new_n16535_, new_n16536_,
    new_n16537_, new_n16538_, new_n16539_, new_n16540_, new_n16541_,
    new_n16542_, new_n16543_, new_n16544_, new_n16545_, new_n16546_,
    new_n16547_, new_n16548_, new_n16549_, new_n16550_, new_n16551_,
    new_n16552_, new_n16553_, new_n16554_, new_n16555_, new_n16556_,
    new_n16557_, new_n16558_, new_n16559_, new_n16560_, new_n16561_,
    new_n16562_, new_n16563_, new_n16564_, new_n16565_, new_n16566_,
    new_n16567_, new_n16568_, new_n16569_, new_n16570_, new_n16571_,
    new_n16572_, new_n16573_, new_n16574_, new_n16575_, new_n16576_,
    new_n16577_, new_n16578_, new_n16579_, new_n16580_, new_n16581_,
    new_n16582_, new_n16583_, new_n16584_, new_n16585_, new_n16586_,
    new_n16587_, new_n16588_, new_n16589_, new_n16590_, new_n16591_,
    new_n16592_, new_n16593_, new_n16594_, new_n16595_, new_n16596_,
    new_n16597_, new_n16598_, new_n16599_, new_n16600_, new_n16601_,
    new_n16602_, new_n16603_, new_n16604_, new_n16605_, new_n16606_,
    new_n16607_, new_n16608_, new_n16609_, new_n16610_, new_n16611_,
    new_n16612_, new_n16613_, new_n16614_, new_n16615_, new_n16616_,
    new_n16617_, new_n16618_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16623_, new_n16624_, new_n16625_, new_n16626_,
    new_n16627_, new_n16628_, new_n16629_, new_n16630_, new_n16631_,
    new_n16632_, new_n16633_, new_n16634_, new_n16635_, new_n16636_,
    new_n16637_, new_n16638_, new_n16639_, new_n16640_, new_n16641_,
    new_n16642_, new_n16643_, new_n16644_, new_n16645_, new_n16646_,
    new_n16647_, new_n16648_, new_n16649_, new_n16650_, new_n16651_,
    new_n16652_, new_n16653_, new_n16654_, new_n16655_, new_n16656_,
    new_n16657_, new_n16658_, new_n16659_, new_n16660_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16729_, new_n16730_, new_n16731_,
    new_n16732_, new_n16733_, new_n16734_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16905_, new_n16906_,
    new_n16907_, new_n16908_, new_n16909_, new_n16910_, new_n16911_,
    new_n16912_, new_n16913_, new_n16914_, new_n16915_, new_n16916_,
    new_n16917_, new_n16918_, new_n16919_, new_n16920_, new_n16921_,
    new_n16922_, new_n16923_, new_n16924_, new_n16925_, new_n16926_,
    new_n16927_, new_n16928_, new_n16929_, new_n16930_, new_n16931_,
    new_n16932_, new_n16933_, new_n16934_, new_n16935_, new_n16936_,
    new_n16937_, new_n16938_, new_n16939_, new_n16940_, new_n16941_,
    new_n16942_, new_n16943_, new_n16944_, new_n16945_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16952_, new_n16953_, new_n16954_, new_n16956_, new_n16957_,
    new_n16958_, new_n16959_, new_n16960_, new_n16961_, new_n16962_,
    new_n16963_, new_n16964_, new_n16965_, new_n16966_, new_n16967_,
    new_n16968_, new_n16969_, new_n16970_, new_n16971_, new_n16972_,
    new_n16973_, new_n16974_, new_n16975_, new_n16976_, new_n16977_,
    new_n16978_, new_n16979_, new_n16980_, new_n16981_, new_n16982_,
    new_n16983_, new_n16984_, new_n16985_, new_n16986_, new_n16987_,
    new_n16988_, new_n16989_, new_n16990_, new_n16991_, new_n16992_,
    new_n16993_, new_n16994_, new_n16995_, new_n16996_, new_n16997_,
    new_n16998_, new_n16999_, new_n17000_, new_n17001_, new_n17002_,
    new_n17003_, new_n17004_, new_n17005_, new_n17006_, new_n17007_,
    new_n17008_, new_n17009_, new_n17010_, new_n17011_, new_n17012_,
    new_n17013_, new_n17014_, new_n17015_, new_n17016_, new_n17017_,
    new_n17018_, new_n17019_, new_n17020_, new_n17021_, new_n17022_,
    new_n17023_, new_n17024_, new_n17025_, new_n17026_, new_n17027_,
    new_n17028_, new_n17029_, new_n17030_, new_n17031_, new_n17032_,
    new_n17033_, new_n17034_, new_n17035_, new_n17036_, new_n17037_,
    new_n17038_, new_n17039_, new_n17040_, new_n17041_, new_n17042_,
    new_n17043_, new_n17044_, new_n17045_, new_n17046_, new_n17047_,
    new_n17048_, new_n17049_, new_n17050_, new_n17051_, new_n17052_,
    new_n17053_, new_n17054_, new_n17055_, new_n17056_, new_n17057_,
    new_n17058_, new_n17059_, new_n17060_, new_n17061_, new_n17062_,
    new_n17063_, new_n17064_, new_n17065_, new_n17066_, new_n17067_,
    new_n17068_, new_n17069_, new_n17070_, new_n17071_, new_n17072_,
    new_n17073_, new_n17074_, new_n17075_, new_n17076_, new_n17077_,
    new_n17078_, new_n17079_, new_n17080_, new_n17081_, new_n17082_,
    new_n17083_, new_n17084_, new_n17085_, new_n17086_, new_n17087_,
    new_n17088_, new_n17089_, new_n17090_, new_n17091_, new_n17092_,
    new_n17093_, new_n17094_, new_n17095_, new_n17096_, new_n17097_,
    new_n17098_, new_n17099_, new_n17100_, new_n17101_, new_n17102_,
    new_n17103_, new_n17104_, new_n17105_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17124_, new_n17125_, new_n17126_, new_n17127_,
    new_n17128_, new_n17129_, new_n17130_, new_n17131_, new_n17132_,
    new_n17133_, new_n17134_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17147_,
    new_n17148_, new_n17149_, new_n17150_, new_n17151_, new_n17152_,
    new_n17153_, new_n17154_, new_n17155_, new_n17156_, new_n17157_,
    new_n17158_, new_n17159_, new_n17160_, new_n17161_, new_n17162_,
    new_n17163_, new_n17164_, new_n17165_, new_n17166_, new_n17167_,
    new_n17168_, new_n17169_, new_n17170_, new_n17171_, new_n17172_,
    new_n17173_, new_n17174_, new_n17175_, new_n17176_, new_n17177_,
    new_n17178_, new_n17179_, new_n17180_, new_n17181_, new_n17182_,
    new_n17183_, new_n17184_, new_n17185_, new_n17186_, new_n17187_,
    new_n17188_, new_n17189_, new_n17190_, new_n17191_, new_n17192_,
    new_n17193_, new_n17194_, new_n17195_, new_n17196_, new_n17197_,
    new_n17198_, new_n17199_, new_n17200_, new_n17201_, new_n17202_,
    new_n17203_, new_n17204_, new_n17205_, new_n17206_, new_n17207_,
    new_n17208_, new_n17209_, new_n17210_, new_n17211_, new_n17212_,
    new_n17213_, new_n17214_, new_n17215_, new_n17216_, new_n17217_,
    new_n17218_, new_n17219_, new_n17220_, new_n17221_, new_n17222_,
    new_n17223_, new_n17224_, new_n17225_, new_n17226_, new_n17227_,
    new_n17228_, new_n17229_, new_n17230_, new_n17231_, new_n17232_,
    new_n17233_, new_n17234_, new_n17235_, new_n17236_, new_n17237_,
    new_n17238_, new_n17239_, new_n17240_, new_n17241_, new_n17242_,
    new_n17243_, new_n17244_, new_n17245_, new_n17246_, new_n17247_,
    new_n17248_, new_n17249_, new_n17250_, new_n17251_, new_n17252_,
    new_n17253_, new_n17254_, new_n17255_, new_n17256_, new_n17257_,
    new_n17258_, new_n17259_, new_n17260_, new_n17261_, new_n17262_,
    new_n17263_, new_n17264_, new_n17265_, new_n17266_, new_n17267_,
    new_n17268_, new_n17269_, new_n17270_, new_n17271_, new_n17272_,
    new_n17273_, new_n17274_, new_n17275_, new_n17276_, new_n17277_,
    new_n17278_, new_n17279_, new_n17280_, new_n17281_, new_n17282_,
    new_n17283_, new_n17284_, new_n17285_, new_n17286_, new_n17287_,
    new_n17288_, new_n17289_, new_n17290_, new_n17291_, new_n17292_,
    new_n17293_, new_n17294_, new_n17295_, new_n17296_, new_n17297_,
    new_n17298_, new_n17299_, new_n17300_, new_n17301_, new_n17302_,
    new_n17303_, new_n17304_, new_n17305_, new_n17306_, new_n17307_,
    new_n17308_, new_n17309_, new_n17310_, new_n17311_, new_n17312_,
    new_n17313_, new_n17314_, new_n17315_, new_n17316_, new_n17317_,
    new_n17318_, new_n17319_, new_n17320_, new_n17321_, new_n17322_,
    new_n17323_, new_n17324_, new_n17325_, new_n17326_, new_n17327_,
    new_n17328_, new_n17329_, new_n17330_, new_n17331_, new_n17332_,
    new_n17333_, new_n17334_, new_n17335_, new_n17336_, new_n17337_,
    new_n17338_, new_n17339_, new_n17340_, new_n17341_, new_n17342_,
    new_n17343_, new_n17344_, new_n17345_, new_n17346_, new_n17347_,
    new_n17348_, new_n17349_, new_n17350_, new_n17351_, new_n17352_,
    new_n17353_, new_n17354_, new_n17355_, new_n17356_, new_n17357_,
    new_n17358_, new_n17359_, new_n17360_, new_n17361_, new_n17362_,
    new_n17363_, new_n17364_, new_n17365_, new_n17366_, new_n17367_,
    new_n17368_, new_n17369_, new_n17370_, new_n17371_, new_n17372_,
    new_n17373_, new_n17374_, new_n17375_, new_n17376_, new_n17377_,
    new_n17378_, new_n17379_, new_n17380_, new_n17381_, new_n17382_,
    new_n17383_, new_n17384_, new_n17385_, new_n17386_, new_n17387_,
    new_n17388_, new_n17389_, new_n17390_, new_n17391_, new_n17392_,
    new_n17393_, new_n17394_, new_n17395_, new_n17396_, new_n17397_,
    new_n17398_, new_n17399_, new_n17400_, new_n17401_, new_n17402_,
    new_n17403_, new_n17404_, new_n17405_, new_n17406_, new_n17407_,
    new_n17408_, new_n17409_, new_n17410_, new_n17411_, new_n17412_,
    new_n17413_, new_n17414_, new_n17415_, new_n17416_, new_n17417_,
    new_n17418_, new_n17419_, new_n17420_, new_n17421_, new_n17422_,
    new_n17423_, new_n17424_, new_n17425_, new_n17426_, new_n17427_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17441_, new_n17442_,
    new_n17443_, new_n17444_, new_n17445_, new_n17446_, new_n17447_,
    new_n17448_, new_n17449_, new_n17450_, new_n17451_, new_n17452_,
    new_n17453_, new_n17454_, new_n17455_, new_n17456_, new_n17457_,
    new_n17458_, new_n17459_, new_n17460_, new_n17461_, new_n17462_,
    new_n17463_, new_n17464_, new_n17465_, new_n17466_, new_n17467_,
    new_n17468_, new_n17469_, new_n17470_, new_n17471_, new_n17472_,
    new_n17473_, new_n17474_, new_n17475_, new_n17476_, new_n17477_,
    new_n17478_, new_n17479_, new_n17480_, new_n17481_, new_n17482_,
    new_n17483_, new_n17484_, new_n17485_, new_n17486_, new_n17487_,
    new_n17488_, new_n17489_, new_n17490_, new_n17491_, new_n17492_,
    new_n17493_, new_n17494_, new_n17495_, new_n17496_, new_n17497_,
    new_n17498_, new_n17499_, new_n17500_, new_n17501_, new_n17502_,
    new_n17503_, new_n17504_, new_n17505_, new_n17506_, new_n17507_,
    new_n17508_, new_n17509_, new_n17510_, new_n17511_, new_n17512_,
    new_n17513_, new_n17514_, new_n17515_, new_n17516_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17560_, new_n17561_, new_n17562_,
    new_n17564_, new_n17565_, new_n17566_, new_n17567_, new_n17568_,
    new_n17569_, new_n17570_, new_n17571_, new_n17572_, new_n17573_,
    new_n17574_, new_n17575_, new_n17576_, new_n17577_, new_n17578_,
    new_n17579_, new_n17580_, new_n17581_, new_n17582_, new_n17583_,
    new_n17584_, new_n17585_, new_n17586_, new_n17587_, new_n17588_,
    new_n17589_, new_n17590_, new_n17591_, new_n17592_, new_n17593_,
    new_n17594_, new_n17595_, new_n17596_, new_n17597_, new_n17598_,
    new_n17599_, new_n17600_, new_n17601_, new_n17602_, new_n17603_,
    new_n17604_, new_n17605_, new_n17606_, new_n17607_, new_n17608_,
    new_n17609_, new_n17610_, new_n17611_, new_n17612_, new_n17613_,
    new_n17614_, new_n17615_, new_n17616_, new_n17617_, new_n17618_,
    new_n17619_, new_n17620_, new_n17621_, new_n17622_, new_n17623_,
    new_n17624_, new_n17625_, new_n17626_, new_n17627_, new_n17628_,
    new_n17629_, new_n17630_, new_n17631_, new_n17632_, new_n17633_,
    new_n17634_, new_n17635_, new_n17636_, new_n17637_, new_n17638_,
    new_n17639_, new_n17640_, new_n17641_, new_n17642_, new_n17643_,
    new_n17644_, new_n17645_, new_n17646_, new_n17647_, new_n17648_,
    new_n17649_, new_n17650_, new_n17651_, new_n17652_, new_n17653_,
    new_n17654_, new_n17655_, new_n17656_, new_n17657_, new_n17658_,
    new_n17659_, new_n17660_, new_n17661_, new_n17662_, new_n17663_,
    new_n17664_, new_n17665_, new_n17666_, new_n17667_, new_n17668_,
    new_n17669_, new_n17670_, new_n17671_, new_n17672_, new_n17673_,
    new_n17674_, new_n17675_, new_n17676_, new_n17677_, new_n17678_,
    new_n17679_, new_n17680_, new_n17681_, new_n17682_, new_n17683_,
    new_n17684_, new_n17685_, new_n17686_, new_n17687_, new_n17688_,
    new_n17689_, new_n17690_, new_n17691_, new_n17692_, new_n17693_,
    new_n17694_, new_n17695_, new_n17696_, new_n17697_, new_n17698_,
    new_n17699_, new_n17700_, new_n17701_, new_n17702_, new_n17703_,
    new_n17704_, new_n17705_, new_n17706_, new_n17707_, new_n17708_,
    new_n17709_, new_n17710_, new_n17711_, new_n17712_, new_n17713_,
    new_n17714_, new_n17715_, new_n17716_, new_n17717_, new_n17718_,
    new_n17719_, new_n17720_, new_n17721_, new_n17722_, new_n17723_,
    new_n17724_, new_n17725_, new_n17726_, new_n17727_, new_n17728_,
    new_n17729_, new_n17730_, new_n17731_, new_n17732_, new_n17733_,
    new_n17734_, new_n17735_, new_n17736_, new_n17737_, new_n17738_,
    new_n17739_, new_n17740_, new_n17741_, new_n17742_, new_n17743_,
    new_n17744_, new_n17745_, new_n17746_, new_n17747_, new_n17748_,
    new_n17749_, new_n17750_, new_n17751_, new_n17752_, new_n17753_,
    new_n17754_, new_n17755_, new_n17756_, new_n17757_, new_n17758_,
    new_n17759_, new_n17760_, new_n17761_, new_n17762_, new_n17763_,
    new_n17764_, new_n17765_, new_n17766_, new_n17767_, new_n17768_,
    new_n17769_, new_n17770_, new_n17771_, new_n17772_, new_n17773_,
    new_n17774_, new_n17775_, new_n17776_, new_n17777_, new_n17778_,
    new_n17779_, new_n17780_, new_n17781_, new_n17782_, new_n17783_,
    new_n17784_, new_n17785_, new_n17786_, new_n17787_, new_n17788_,
    new_n17789_, new_n17790_, new_n17791_, new_n17792_, new_n17793_,
    new_n17794_, new_n17795_, new_n17796_, new_n17797_, new_n17798_,
    new_n17799_, new_n17800_, new_n17801_, new_n17802_, new_n17803_,
    new_n17804_, new_n17805_, new_n17806_, new_n17807_, new_n17808_,
    new_n17809_, new_n17810_, new_n17811_, new_n17812_, new_n17813_,
    new_n17814_, new_n17815_, new_n17816_, new_n17817_, new_n17818_,
    new_n17819_, new_n17820_, new_n17821_, new_n17822_, new_n17823_,
    new_n17824_, new_n17825_, new_n17826_, new_n17827_, new_n17828_,
    new_n17829_, new_n17830_, new_n17831_, new_n17832_, new_n17833_,
    new_n17834_, new_n17835_, new_n17836_, new_n17837_, new_n17838_,
    new_n17839_, new_n17840_, new_n17841_, new_n17842_, new_n17843_,
    new_n17844_, new_n17845_, new_n17846_, new_n17847_, new_n17848_,
    new_n17849_, new_n17850_, new_n17851_, new_n17852_, new_n17853_,
    new_n17854_, new_n17855_, new_n17856_, new_n17857_, new_n17858_,
    new_n17859_, new_n17860_, new_n17861_, new_n17862_, new_n17863_,
    new_n17864_, new_n17865_, new_n17866_, new_n17867_, new_n17868_,
    new_n17869_, new_n17870_, new_n17871_, new_n17872_, new_n17873_,
    new_n17874_, new_n17875_, new_n17876_, new_n17877_, new_n17878_,
    new_n17879_, new_n17880_, new_n17881_, new_n17882_, new_n17883_,
    new_n17884_, new_n17885_, new_n17886_, new_n17887_, new_n17888_,
    new_n17889_, new_n17890_, new_n17891_, new_n17892_, new_n17893_,
    new_n17894_, new_n17895_, new_n17896_, new_n17897_, new_n17898_,
    new_n17899_, new_n17900_, new_n17901_, new_n17902_, new_n17903_,
    new_n17904_, new_n17905_, new_n17906_, new_n17907_, new_n17908_,
    new_n17909_, new_n17910_, new_n17911_, new_n17912_, new_n17913_,
    new_n17914_, new_n17915_, new_n17916_, new_n17917_, new_n17918_,
    new_n17919_, new_n17920_, new_n17921_, new_n17922_, new_n17923_,
    new_n17924_, new_n17925_, new_n17926_, new_n17927_, new_n17928_,
    new_n17929_, new_n17930_, new_n17931_, new_n17932_, new_n17933_,
    new_n17934_, new_n17935_, new_n17936_, new_n17937_, new_n17938_,
    new_n17939_, new_n17940_, new_n17941_, new_n17942_, new_n17943_,
    new_n17944_, new_n17945_, new_n17946_, new_n17947_, new_n17948_,
    new_n17949_, new_n17950_, new_n17951_, new_n17952_, new_n17953_,
    new_n17954_, new_n17955_, new_n17956_, new_n17957_, new_n17958_,
    new_n17959_, new_n17960_, new_n17961_, new_n17962_, new_n17963_,
    new_n17964_, new_n17965_, new_n17966_, new_n17967_, new_n17968_,
    new_n17969_, new_n17970_, new_n17971_, new_n17972_, new_n17973_,
    new_n17974_, new_n17975_, new_n17976_, new_n17977_, new_n17978_,
    new_n17979_, new_n17980_, new_n17981_, new_n17982_, new_n17983_,
    new_n17984_, new_n17985_, new_n17986_, new_n17987_, new_n17988_,
    new_n17989_, new_n17990_, new_n17991_, new_n17992_, new_n17993_,
    new_n17994_, new_n17995_, new_n17996_, new_n17997_, new_n17998_,
    new_n17999_, new_n18000_, new_n18001_, new_n18002_, new_n18003_,
    new_n18004_, new_n18005_, new_n18006_, new_n18007_, new_n18008_,
    new_n18009_, new_n18010_, new_n18011_, new_n18012_, new_n18013_,
    new_n18014_, new_n18015_, new_n18016_, new_n18017_, new_n18018_,
    new_n18019_, new_n18020_, new_n18021_, new_n18022_, new_n18023_,
    new_n18024_, new_n18025_, new_n18026_, new_n18027_, new_n18028_,
    new_n18029_, new_n18030_, new_n18031_, new_n18032_, new_n18033_,
    new_n18034_, new_n18035_, new_n18036_, new_n18037_, new_n18038_,
    new_n18039_, new_n18040_, new_n18041_, new_n18042_, new_n18043_,
    new_n18044_, new_n18045_, new_n18046_, new_n18047_, new_n18048_,
    new_n18049_, new_n18050_, new_n18051_, new_n18052_, new_n18053_,
    new_n18054_, new_n18055_, new_n18056_, new_n18057_, new_n18058_,
    new_n18059_, new_n18060_, new_n18061_, new_n18062_, new_n18063_,
    new_n18064_, new_n18065_, new_n18066_, new_n18067_, new_n18068_,
    new_n18069_, new_n18070_, new_n18071_, new_n18072_, new_n18073_,
    new_n18074_, new_n18075_, new_n18076_, new_n18077_, new_n18078_,
    new_n18079_, new_n18080_, new_n18081_, new_n18082_, new_n18083_,
    new_n18084_, new_n18085_, new_n18086_, new_n18087_, new_n18088_,
    new_n18089_, new_n18090_, new_n18091_, new_n18092_, new_n18093_,
    new_n18094_, new_n18095_, new_n18096_, new_n18097_, new_n18098_,
    new_n18099_, new_n18100_, new_n18101_, new_n18102_, new_n18103_,
    new_n18104_, new_n18105_, new_n18106_, new_n18107_, new_n18108_,
    new_n18109_, new_n18110_, new_n18111_, new_n18112_, new_n18113_,
    new_n18114_, new_n18115_, new_n18116_, new_n18117_, new_n18118_,
    new_n18119_, new_n18120_, new_n18121_, new_n18122_, new_n18123_,
    new_n18124_, new_n18125_, new_n18126_, new_n18127_, new_n18128_,
    new_n18129_, new_n18130_, new_n18131_, new_n18132_, new_n18133_,
    new_n18134_, new_n18135_, new_n18136_, new_n18137_, new_n18138_,
    new_n18139_, new_n18140_, new_n18141_, new_n18142_, new_n18143_,
    new_n18144_, new_n18145_, new_n18146_, new_n18147_, new_n18148_,
    new_n18149_, new_n18150_, new_n18151_, new_n18152_, new_n18153_,
    new_n18154_, new_n18155_, new_n18156_, new_n18157_, new_n18158_,
    new_n18159_, new_n18160_, new_n18161_, new_n18162_, new_n18163_,
    new_n18164_, new_n18165_, new_n18166_, new_n18167_, new_n18168_,
    new_n18169_, new_n18170_, new_n18171_, new_n18172_, new_n18173_,
    new_n18174_, new_n18175_, new_n18176_, new_n18177_, new_n18178_,
    new_n18179_, new_n18180_, new_n18181_, new_n18182_, new_n18183_,
    new_n18184_, new_n18185_, new_n18186_, new_n18187_, new_n18188_,
    new_n18189_, new_n18190_, new_n18191_, new_n18192_, new_n18193_,
    new_n18194_, new_n18195_, new_n18196_, new_n18197_, new_n18198_,
    new_n18199_, new_n18200_, new_n18201_, new_n18202_, new_n18203_,
    new_n18204_, new_n18205_, new_n18206_, new_n18207_, new_n18208_,
    new_n18209_, new_n18210_, new_n18211_, new_n18212_, new_n18213_,
    new_n18214_, new_n18215_, new_n18216_, new_n18217_, new_n18218_,
    new_n18219_, new_n18220_, new_n18221_, new_n18222_, new_n18223_,
    new_n18224_, new_n18226_, new_n18227_, new_n18228_, new_n18229_,
    new_n18230_, new_n18231_, new_n18232_, new_n18233_, new_n18234_,
    new_n18235_, new_n18236_, new_n18237_, new_n18238_, new_n18239_,
    new_n18240_, new_n18241_, new_n18242_, new_n18243_, new_n18244_,
    new_n18245_, new_n18246_, new_n18247_, new_n18248_, new_n18249_,
    new_n18250_, new_n18251_, new_n18252_, new_n18253_, new_n18254_,
    new_n18255_, new_n18256_, new_n18257_, new_n18258_, new_n18259_,
    new_n18260_, new_n18261_, new_n18262_, new_n18263_, new_n18264_,
    new_n18265_, new_n18266_, new_n18267_, new_n18268_, new_n18269_,
    new_n18270_, new_n18271_, new_n18272_, new_n18273_, new_n18274_,
    new_n18275_, new_n18276_, new_n18277_, new_n18278_, new_n18279_,
    new_n18280_, new_n18281_, new_n18282_, new_n18283_, new_n18284_,
    new_n18285_, new_n18286_, new_n18287_, new_n18288_, new_n18289_,
    new_n18290_, new_n18291_, new_n18292_, new_n18293_, new_n18294_,
    new_n18295_, new_n18296_, new_n18297_, new_n18298_, new_n18299_,
    new_n18300_, new_n18301_, new_n18302_, new_n18303_, new_n18304_,
    new_n18305_, new_n18306_, new_n18307_, new_n18308_, new_n18309_,
    new_n18310_, new_n18311_, new_n18312_, new_n18313_, new_n18314_,
    new_n18315_, new_n18316_, new_n18317_, new_n18318_, new_n18319_,
    new_n18320_, new_n18321_, new_n18322_, new_n18323_, new_n18324_,
    new_n18325_, new_n18326_, new_n18327_, new_n18328_, new_n18329_,
    new_n18330_, new_n18331_, new_n18332_, new_n18333_, new_n18334_,
    new_n18335_, new_n18336_, new_n18337_, new_n18338_, new_n18339_,
    new_n18340_, new_n18341_, new_n18342_, new_n18343_, new_n18344_,
    new_n18345_, new_n18346_, new_n18347_, new_n18348_, new_n18349_,
    new_n18350_, new_n18351_, new_n18352_, new_n18353_, new_n18354_,
    new_n18355_, new_n18356_, new_n18357_, new_n18358_, new_n18359_,
    new_n18360_, new_n18361_, new_n18362_, new_n18363_, new_n18364_,
    new_n18365_, new_n18366_, new_n18367_, new_n18368_, new_n18369_,
    new_n18370_, new_n18371_, new_n18372_, new_n18373_, new_n18374_,
    new_n18375_, new_n18376_, new_n18377_, new_n18378_, new_n18379_,
    new_n18380_, new_n18381_, new_n18382_, new_n18383_, new_n18384_,
    new_n18385_, new_n18386_, new_n18387_, new_n18388_, new_n18389_,
    new_n18390_, new_n18391_, new_n18392_, new_n18393_, new_n18394_,
    new_n18395_, new_n18396_, new_n18397_, new_n18398_, new_n18399_,
    new_n18400_, new_n18401_, new_n18402_, new_n18403_, new_n18404_,
    new_n18405_, new_n18406_, new_n18407_, new_n18408_, new_n18409_,
    new_n18410_, new_n18411_, new_n18412_, new_n18413_, new_n18414_,
    new_n18415_, new_n18416_, new_n18417_, new_n18418_, new_n18419_,
    new_n18420_, new_n18421_, new_n18422_, new_n18423_, new_n18424_,
    new_n18425_, new_n18426_, new_n18427_, new_n18428_, new_n18429_,
    new_n18430_, new_n18431_, new_n18432_, new_n18433_, new_n18434_,
    new_n18435_, new_n18436_, new_n18437_, new_n18438_, new_n18439_,
    new_n18440_, new_n18441_, new_n18442_, new_n18443_, new_n18444_,
    new_n18445_, new_n18446_, new_n18447_, new_n18448_, new_n18449_,
    new_n18450_, new_n18451_, new_n18452_, new_n18453_, new_n18454_,
    new_n18455_, new_n18456_, new_n18457_, new_n18458_, new_n18459_,
    new_n18460_, new_n18461_, new_n18462_, new_n18463_, new_n18464_,
    new_n18465_, new_n18466_, new_n18467_, new_n18468_, new_n18469_,
    new_n18470_, new_n18471_, new_n18472_, new_n18473_, new_n18474_,
    new_n18475_, new_n18476_, new_n18477_, new_n18478_, new_n18479_,
    new_n18480_, new_n18481_, new_n18482_, new_n18483_, new_n18484_,
    new_n18485_, new_n18486_, new_n18487_, new_n18488_, new_n18489_,
    new_n18490_, new_n18491_, new_n18492_, new_n18493_, new_n18494_,
    new_n18495_, new_n18496_, new_n18497_, new_n18498_, new_n18499_,
    new_n18500_, new_n18501_, new_n18502_, new_n18503_, new_n18504_,
    new_n18505_, new_n18506_, new_n18507_, new_n18508_, new_n18509_,
    new_n18510_, new_n18511_, new_n18512_, new_n18513_, new_n18514_,
    new_n18515_, new_n18516_, new_n18517_, new_n18518_, new_n18519_,
    new_n18520_, new_n18521_, new_n18522_, new_n18523_, new_n18524_,
    new_n18525_, new_n18526_, new_n18527_, new_n18528_, new_n18529_,
    new_n18530_, new_n18531_, new_n18532_, new_n18533_, new_n18534_,
    new_n18535_, new_n18536_, new_n18537_, new_n18538_, new_n18539_,
    new_n18540_, new_n18541_, new_n18542_, new_n18543_, new_n18544_,
    new_n18545_, new_n18546_, new_n18547_, new_n18548_, new_n18549_,
    new_n18550_, new_n18551_, new_n18552_, new_n18553_, new_n18554_,
    new_n18555_, new_n18556_, new_n18557_, new_n18558_, new_n18559_,
    new_n18560_, new_n18561_, new_n18562_, new_n18563_, new_n18564_,
    new_n18565_, new_n18566_, new_n18567_, new_n18568_, new_n18569_,
    new_n18570_, new_n18571_, new_n18572_, new_n18573_, new_n18574_,
    new_n18575_, new_n18576_, new_n18577_, new_n18578_, new_n18579_,
    new_n18580_, new_n18581_, new_n18582_, new_n18583_, new_n18584_,
    new_n18585_, new_n18586_, new_n18587_, new_n18588_, new_n18589_,
    new_n18590_, new_n18591_, new_n18592_, new_n18593_, new_n18594_,
    new_n18595_, new_n18596_, new_n18597_, new_n18598_, new_n18599_,
    new_n18600_, new_n18601_, new_n18602_, new_n18603_, new_n18604_,
    new_n18605_, new_n18606_, new_n18607_, new_n18608_, new_n18609_,
    new_n18610_, new_n18611_, new_n18612_, new_n18613_, new_n18614_,
    new_n18615_, new_n18616_, new_n18617_, new_n18618_, new_n18619_,
    new_n18620_, new_n18621_, new_n18622_, new_n18623_, new_n18624_,
    new_n18625_, new_n18626_, new_n18627_, new_n18628_, new_n18629_,
    new_n18630_, new_n18631_, new_n18632_, new_n18633_, new_n18634_,
    new_n18635_, new_n18636_, new_n18637_, new_n18638_, new_n18639_,
    new_n18640_, new_n18641_, new_n18642_, new_n18643_, new_n18644_,
    new_n18645_, new_n18646_, new_n18647_, new_n18648_, new_n18649_,
    new_n18650_, new_n18651_, new_n18652_, new_n18653_, new_n18654_,
    new_n18655_, new_n18656_, new_n18657_, new_n18658_, new_n18659_,
    new_n18660_, new_n18661_, new_n18662_, new_n18663_, new_n18664_,
    new_n18665_, new_n18666_, new_n18667_, new_n18668_, new_n18669_,
    new_n18670_, new_n18671_, new_n18672_, new_n18673_, new_n18674_,
    new_n18675_, new_n18676_, new_n18677_, new_n18678_, new_n18679_,
    new_n18680_, new_n18681_, new_n18682_, new_n18683_, new_n18684_,
    new_n18685_, new_n18686_, new_n18687_, new_n18688_, new_n18689_,
    new_n18690_, new_n18691_, new_n18692_, new_n18693_, new_n18694_,
    new_n18695_, new_n18696_, new_n18697_, new_n18698_, new_n18699_,
    new_n18700_, new_n18701_, new_n18702_, new_n18703_, new_n18704_,
    new_n18705_, new_n18706_, new_n18707_, new_n18708_, new_n18709_,
    new_n18710_, new_n18711_, new_n18712_, new_n18713_, new_n18714_,
    new_n18715_, new_n18716_, new_n18717_, new_n18718_, new_n18719_,
    new_n18720_, new_n18721_, new_n18722_, new_n18723_, new_n18724_,
    new_n18725_, new_n18726_, new_n18727_, new_n18728_, new_n18729_,
    new_n18730_, new_n18731_, new_n18732_, new_n18733_, new_n18734_,
    new_n18735_, new_n18736_, new_n18737_, new_n18738_, new_n18739_,
    new_n18740_, new_n18741_, new_n18742_, new_n18743_, new_n18744_,
    new_n18745_, new_n18746_, new_n18747_, new_n18748_, new_n18749_,
    new_n18750_, new_n18751_, new_n18752_, new_n18753_, new_n18754_,
    new_n18755_, new_n18756_, new_n18757_, new_n18758_, new_n18759_,
    new_n18760_, new_n18761_, new_n18762_, new_n18763_, new_n18764_,
    new_n18765_, new_n18766_, new_n18767_, new_n18768_, new_n18769_,
    new_n18770_, new_n18771_, new_n18772_, new_n18773_, new_n18774_,
    new_n18775_, new_n18776_, new_n18777_, new_n18778_, new_n18779_,
    new_n18780_, new_n18781_, new_n18782_, new_n18783_, new_n18784_,
    new_n18785_, new_n18786_, new_n18787_, new_n18788_, new_n18789_,
    new_n18790_, new_n18791_, new_n18792_, new_n18793_, new_n18794_,
    new_n18795_, new_n18796_, new_n18797_, new_n18798_, new_n18799_,
    new_n18800_, new_n18801_, new_n18802_, new_n18803_, new_n18804_,
    new_n18805_, new_n18806_, new_n18807_, new_n18808_, new_n18809_,
    new_n18810_, new_n18811_, new_n18812_, new_n18813_, new_n18814_,
    new_n18815_, new_n18816_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18821_, new_n18822_, new_n18823_, new_n18824_,
    new_n18825_, new_n18826_, new_n18827_, new_n18828_, new_n18829_,
    new_n18830_, new_n18831_, new_n18832_, new_n18833_, new_n18834_,
    new_n18835_, new_n18836_, new_n18837_, new_n18838_, new_n18839_,
    new_n18840_, new_n18841_, new_n18842_, new_n18843_, new_n18844_,
    new_n18845_, new_n18846_, new_n18847_, new_n18848_, new_n18849_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18867_, new_n18868_, new_n18869_, new_n18870_,
    new_n18871_, new_n18872_, new_n18873_, new_n18874_, new_n18875_,
    new_n18876_, new_n18877_, new_n18878_, new_n18879_, new_n18880_,
    new_n18881_, new_n18882_, new_n18883_, new_n18884_, new_n18885_,
    new_n18886_, new_n18887_, new_n18888_, new_n18889_, new_n18890_,
    new_n18891_, new_n18892_, new_n18893_, new_n18894_, new_n18895_,
    new_n18896_, new_n18897_, new_n18898_, new_n18899_, new_n18900_,
    new_n18901_, new_n18902_, new_n18903_, new_n18904_, new_n18905_,
    new_n18906_, new_n18907_, new_n18908_, new_n18909_, new_n18910_,
    new_n18911_, new_n18912_, new_n18913_, new_n18914_, new_n18915_,
    new_n18916_, new_n18917_, new_n18918_, new_n18919_, new_n18920_,
    new_n18921_, new_n18922_, new_n18923_, new_n18924_, new_n18925_,
    new_n18926_, new_n18927_, new_n18928_, new_n18929_, new_n18930_,
    new_n18931_, new_n18932_, new_n18933_, new_n18934_, new_n18935_,
    new_n18936_, new_n18937_, new_n18938_, new_n18939_, new_n18940_,
    new_n18941_, new_n18942_, new_n18943_, new_n18944_, new_n18945_,
    new_n18946_, new_n18947_, new_n18948_, new_n18949_, new_n18950_,
    new_n18951_, new_n18952_, new_n18953_, new_n18954_, new_n18955_,
    new_n18956_, new_n18957_, new_n18958_, new_n18959_, new_n18960_,
    new_n18961_, new_n18962_, new_n18963_, new_n18964_, new_n18965_,
    new_n18966_, new_n18967_, new_n18968_, new_n18969_, new_n18970_,
    new_n18971_, new_n18972_, new_n18973_, new_n18974_, new_n18975_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19089_, new_n19090_,
    new_n19091_, new_n19092_, new_n19093_, new_n19094_, new_n19095_,
    new_n19096_, new_n19097_, new_n19098_, new_n19099_, new_n19100_,
    new_n19101_, new_n19102_, new_n19103_, new_n19104_, new_n19105_,
    new_n19106_, new_n19107_, new_n19108_, new_n19109_, new_n19110_,
    new_n19111_, new_n19112_, new_n19113_, new_n19114_, new_n19115_,
    new_n19116_, new_n19117_, new_n19118_, new_n19119_, new_n19120_,
    new_n19121_, new_n19122_, new_n19123_, new_n19124_, new_n19125_,
    new_n19126_, new_n19127_, new_n19128_, new_n19129_, new_n19130_,
    new_n19131_, new_n19132_, new_n19133_, new_n19134_, new_n19135_,
    new_n19136_, new_n19137_, new_n19138_, new_n19139_, new_n19140_,
    new_n19141_, new_n19142_, new_n19143_, new_n19144_, new_n19145_,
    new_n19146_, new_n19147_, new_n19148_, new_n19149_, new_n19150_,
    new_n19151_, new_n19152_, new_n19153_, new_n19154_, new_n19155_,
    new_n19156_, new_n19157_, new_n19158_, new_n19159_, new_n19160_,
    new_n19161_, new_n19162_, new_n19163_, new_n19164_, new_n19165_,
    new_n19166_, new_n19167_, new_n19168_, new_n19169_, new_n19170_,
    new_n19171_, new_n19172_, new_n19173_, new_n19174_, new_n19175_,
    new_n19176_, new_n19177_, new_n19178_, new_n19179_, new_n19180_,
    new_n19181_, new_n19182_, new_n19183_, new_n19184_, new_n19185_,
    new_n19186_, new_n19187_, new_n19188_, new_n19189_, new_n19190_,
    new_n19191_, new_n19192_, new_n19193_, new_n19194_, new_n19195_,
    new_n19196_, new_n19197_, new_n19198_, new_n19199_, new_n19200_,
    new_n19201_, new_n19202_, new_n19203_, new_n19204_, new_n19205_,
    new_n19206_, new_n19207_, new_n19208_, new_n19209_, new_n19210_,
    new_n19211_, new_n19212_, new_n19213_, new_n19214_, new_n19215_,
    new_n19216_, new_n19217_, new_n19218_, new_n19219_, new_n19220_,
    new_n19221_, new_n19222_, new_n19223_, new_n19224_, new_n19225_,
    new_n19226_, new_n19227_, new_n19228_, new_n19229_, new_n19230_,
    new_n19231_, new_n19232_, new_n19233_, new_n19234_, new_n19235_,
    new_n19236_, new_n19237_, new_n19238_, new_n19239_, new_n19240_,
    new_n19241_, new_n19242_, new_n19243_, new_n19244_, new_n19245_,
    new_n19246_, new_n19247_, new_n19248_, new_n19249_, new_n19250_,
    new_n19251_, new_n19252_, new_n19253_, new_n19254_, new_n19255_,
    new_n19256_, new_n19257_, new_n19258_, new_n19259_, new_n19260_,
    new_n19261_, new_n19262_, new_n19263_, new_n19264_, new_n19265_,
    new_n19266_, new_n19267_, new_n19268_, new_n19269_, new_n19270_,
    new_n19271_, new_n19272_, new_n19273_, new_n19274_, new_n19275_,
    new_n19276_, new_n19277_, new_n19278_, new_n19279_, new_n19280_,
    new_n19281_, new_n19282_, new_n19283_, new_n19284_, new_n19285_,
    new_n19286_, new_n19287_, new_n19288_, new_n19289_, new_n19290_,
    new_n19291_, new_n19292_, new_n19293_, new_n19294_, new_n19295_,
    new_n19296_, new_n19297_, new_n19298_, new_n19299_, new_n19300_,
    new_n19301_, new_n19302_, new_n19303_, new_n19304_, new_n19305_,
    new_n19306_, new_n19307_, new_n19308_, new_n19309_, new_n19310_,
    new_n19311_, new_n19312_, new_n19313_, new_n19314_, new_n19315_,
    new_n19316_, new_n19317_, new_n19318_, new_n19319_, new_n19320_,
    new_n19321_, new_n19322_, new_n19323_, new_n19324_, new_n19325_,
    new_n19326_, new_n19327_, new_n19328_, new_n19329_, new_n19330_,
    new_n19331_, new_n19332_, new_n19333_, new_n19334_, new_n19335_,
    new_n19336_, new_n19337_, new_n19338_, new_n19339_, new_n19340_,
    new_n19341_, new_n19342_, new_n19343_, new_n19344_, new_n19345_,
    new_n19346_, new_n19347_, new_n19348_, new_n19349_, new_n19350_,
    new_n19351_, new_n19352_, new_n19353_, new_n19354_, new_n19355_,
    new_n19356_, new_n19357_, new_n19358_, new_n19359_, new_n19360_,
    new_n19361_, new_n19362_, new_n19363_, new_n19364_, new_n19365_,
    new_n19366_, new_n19367_, new_n19368_, new_n19369_, new_n19370_,
    new_n19371_, new_n19372_, new_n19373_, new_n19374_, new_n19375_,
    new_n19376_, new_n19377_, new_n19378_, new_n19379_, new_n19380_,
    new_n19381_, new_n19382_, new_n19383_, new_n19384_, new_n19385_,
    new_n19386_, new_n19387_, new_n19388_, new_n19389_, new_n19390_,
    new_n19391_, new_n19392_, new_n19393_, new_n19394_, new_n19395_,
    new_n19396_, new_n19397_, new_n19398_, new_n19399_, new_n19400_,
    new_n19401_, new_n19402_, new_n19403_, new_n19404_, new_n19405_,
    new_n19406_, new_n19407_, new_n19408_, new_n19409_, new_n19410_,
    new_n19411_, new_n19412_, new_n19413_, new_n19414_, new_n19415_,
    new_n19416_, new_n19417_, new_n19418_, new_n19419_, new_n19420_,
    new_n19421_, new_n19422_, new_n19423_, new_n19424_, new_n19425_,
    new_n19426_, new_n19427_, new_n19428_, new_n19429_, new_n19430_,
    new_n19431_, new_n19432_, new_n19433_, new_n19434_, new_n19435_,
    new_n19436_, new_n19437_, new_n19438_, new_n19439_, new_n19440_,
    new_n19441_, new_n19442_, new_n19443_, new_n19444_, new_n19445_,
    new_n19446_, new_n19447_, new_n19448_, new_n19449_, new_n19450_,
    new_n19451_, new_n19452_, new_n19453_, new_n19454_, new_n19455_,
    new_n19456_, new_n19457_, new_n19458_, new_n19459_, new_n19460_,
    new_n19461_, new_n19462_, new_n19463_, new_n19464_, new_n19465_,
    new_n19466_, new_n19467_, new_n19468_, new_n19469_, new_n19470_,
    new_n19471_, new_n19472_, new_n19473_, new_n19474_, new_n19475_,
    new_n19476_, new_n19477_, new_n19478_, new_n19479_, new_n19480_,
    new_n19481_, new_n19482_, new_n19483_, new_n19484_, new_n19485_,
    new_n19486_, new_n19487_, new_n19488_, new_n19489_, new_n19490_,
    new_n19491_, new_n19492_, new_n19493_, new_n19494_, new_n19495_,
    new_n19496_, new_n19497_, new_n19498_, new_n19499_, new_n19500_,
    new_n19501_, new_n19502_, new_n19503_, new_n19504_, new_n19505_,
    new_n19506_, new_n19507_, new_n19508_, new_n19509_, new_n19510_,
    new_n19511_, new_n19512_, new_n19514_, new_n19515_, new_n19516_,
    new_n19517_, new_n19518_, new_n19519_, new_n19520_, new_n19521_,
    new_n19522_, new_n19523_, new_n19524_, new_n19525_, new_n19526_,
    new_n19527_, new_n19528_, new_n19529_, new_n19530_, new_n19531_,
    new_n19532_, new_n19533_, new_n19534_, new_n19535_, new_n19536_,
    new_n19537_, new_n19538_, new_n19539_, new_n19540_, new_n19541_,
    new_n19542_, new_n19543_, new_n19544_, new_n19545_, new_n19546_,
    new_n19547_, new_n19548_, new_n19549_, new_n19550_, new_n19551_,
    new_n19552_, new_n19553_, new_n19554_, new_n19555_, new_n19556_,
    new_n19557_, new_n19558_, new_n19559_, new_n19560_, new_n19561_,
    new_n19562_, new_n19563_, new_n19564_, new_n19565_, new_n19566_,
    new_n19567_, new_n19568_, new_n19569_, new_n19570_, new_n19571_,
    new_n19572_, new_n19573_, new_n19574_, new_n19575_, new_n19576_,
    new_n19577_, new_n19578_, new_n19579_, new_n19580_, new_n19581_,
    new_n19582_, new_n19583_, new_n19584_, new_n19585_, new_n19586_,
    new_n19587_, new_n19588_, new_n19589_, new_n19590_, new_n19591_,
    new_n19592_, new_n19593_, new_n19594_, new_n19595_, new_n19596_,
    new_n19597_, new_n19598_, new_n19599_, new_n19600_, new_n19601_,
    new_n19602_, new_n19603_, new_n19604_, new_n19605_, new_n19606_,
    new_n19607_, new_n19608_, new_n19609_, new_n19610_, new_n19611_,
    new_n19612_, new_n19613_, new_n19614_, new_n19615_, new_n19616_,
    new_n19617_, new_n19618_, new_n19619_, new_n19620_, new_n19621_,
    new_n19622_, new_n19623_, new_n19624_, new_n19625_, new_n19626_,
    new_n19627_, new_n19628_, new_n19629_, new_n19630_, new_n19631_,
    new_n19632_, new_n19633_, new_n19634_, new_n19635_, new_n19636_,
    new_n19637_, new_n19638_, new_n19639_, new_n19640_, new_n19641_,
    new_n19642_, new_n19643_, new_n19644_, new_n19645_, new_n19646_,
    new_n19647_, new_n19648_, new_n19649_, new_n19650_, new_n19651_,
    new_n19652_, new_n19653_, new_n19654_, new_n19655_, new_n19656_,
    new_n19657_, new_n19658_, new_n19659_, new_n19660_, new_n19661_,
    new_n19662_, new_n19663_, new_n19664_, new_n19665_, new_n19666_,
    new_n19667_, new_n19668_, new_n19669_, new_n19670_, new_n19671_,
    new_n19672_, new_n19673_, new_n19674_, new_n19675_, new_n19676_,
    new_n19677_, new_n19678_, new_n19679_, new_n19680_, new_n19681_,
    new_n19682_, new_n19683_, new_n19684_, new_n19685_, new_n19686_,
    new_n19687_, new_n19688_, new_n19689_, new_n19690_, new_n19691_,
    new_n19692_, new_n19693_, new_n19694_, new_n19695_, new_n19696_,
    new_n19697_, new_n19698_, new_n19699_, new_n19700_, new_n19701_,
    new_n19702_, new_n19703_, new_n19704_, new_n19705_, new_n19706_,
    new_n19707_, new_n19708_, new_n19709_, new_n19710_, new_n19711_,
    new_n19712_, new_n19713_, new_n19714_, new_n19715_, new_n19716_,
    new_n19717_, new_n19718_, new_n19719_, new_n19720_, new_n19721_,
    new_n19722_, new_n19723_, new_n19724_, new_n19725_, new_n19726_,
    new_n19727_, new_n19728_, new_n19729_, new_n19730_, new_n19731_,
    new_n19732_, new_n19733_, new_n19734_, new_n19735_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19804_, new_n19805_, new_n19806_,
    new_n19807_, new_n19808_, new_n19809_, new_n19810_, new_n19811_,
    new_n19812_, new_n19813_, new_n19814_, new_n19815_, new_n19816_,
    new_n19817_, new_n19818_, new_n19819_, new_n19820_, new_n19821_,
    new_n19822_, new_n19823_, new_n19824_, new_n19825_, new_n19826_,
    new_n19827_, new_n19828_, new_n19829_, new_n19830_, new_n19831_,
    new_n19832_, new_n19833_, new_n19834_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19840_, new_n19841_,
    new_n19842_, new_n19843_, new_n19844_, new_n19845_, new_n19846_,
    new_n19847_, new_n19848_, new_n19849_, new_n19850_, new_n19851_,
    new_n19852_, new_n19853_, new_n19854_, new_n19855_, new_n19856_,
    new_n19857_, new_n19858_, new_n19859_, new_n19860_, new_n19861_,
    new_n19862_, new_n19863_, new_n19864_, new_n19865_, new_n19866_,
    new_n19867_, new_n19868_, new_n19869_, new_n19870_, new_n19871_,
    new_n19872_, new_n19873_, new_n19874_, new_n19875_, new_n19876_,
    new_n19877_, new_n19878_, new_n19879_, new_n19880_, new_n19881_,
    new_n19882_, new_n19883_, new_n19884_, new_n19885_, new_n19886_,
    new_n19887_, new_n19888_, new_n19889_, new_n19890_, new_n19891_,
    new_n19892_, new_n19893_, new_n19894_, new_n19895_, new_n19896_,
    new_n19897_, new_n19898_, new_n19899_, new_n19900_, new_n19901_,
    new_n19902_, new_n19903_, new_n19904_, new_n19905_, new_n19906_,
    new_n19907_, new_n19908_, new_n19909_, new_n19910_, new_n19911_,
    new_n19912_, new_n19913_, new_n19914_, new_n19915_, new_n19916_,
    new_n19917_, new_n19918_, new_n19919_, new_n19920_, new_n19921_,
    new_n19922_, new_n19923_, new_n19924_, new_n19925_, new_n19926_,
    new_n19927_, new_n19928_, new_n19929_, new_n19930_, new_n19931_,
    new_n19932_, new_n19933_, new_n19934_, new_n19935_, new_n19936_,
    new_n19937_, new_n19938_, new_n19939_, new_n19940_, new_n19941_,
    new_n19942_, new_n19943_, new_n19944_, new_n19945_, new_n19946_,
    new_n19947_, new_n19948_, new_n19949_, new_n19950_, new_n19951_,
    new_n19952_, new_n19953_, new_n19954_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20127_, new_n20128_, new_n20129_, new_n20130_, new_n20131_,
    new_n20132_, new_n20133_, new_n20134_, new_n20135_, new_n20136_,
    new_n20137_, new_n20138_, new_n20139_, new_n20140_, new_n20141_,
    new_n20142_, new_n20143_, new_n20144_, new_n20145_, new_n20146_,
    new_n20147_, new_n20148_, new_n20149_, new_n20150_, new_n20151_,
    new_n20152_, new_n20153_, new_n20154_, new_n20155_, new_n20156_,
    new_n20157_, new_n20158_, new_n20159_, new_n20160_, new_n20161_,
    new_n20162_, new_n20163_, new_n20164_, new_n20165_, new_n20166_,
    new_n20167_, new_n20168_, new_n20169_, new_n20170_, new_n20171_,
    new_n20172_, new_n20173_, new_n20174_, new_n20175_, new_n20176_,
    new_n20177_, new_n20178_, new_n20179_, new_n20180_, new_n20181_,
    new_n20182_, new_n20183_, new_n20184_, new_n20185_, new_n20186_,
    new_n20187_, new_n20188_, new_n20189_, new_n20190_, new_n20191_,
    new_n20192_, new_n20193_, new_n20194_, new_n20195_, new_n20196_,
    new_n20197_, new_n20198_, new_n20199_, new_n20200_, new_n20201_,
    new_n20202_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20211_, new_n20212_,
    new_n20213_, new_n20214_, new_n20215_, new_n20216_, new_n20217_,
    new_n20218_, new_n20219_, new_n20220_, new_n20221_, new_n20222_,
    new_n20223_, new_n20224_, new_n20225_, new_n20226_, new_n20227_,
    new_n20228_, new_n20229_, new_n20230_, new_n20231_, new_n20232_,
    new_n20233_, new_n20234_, new_n20235_, new_n20236_, new_n20237_,
    new_n20238_, new_n20239_, new_n20240_, new_n20241_, new_n20242_,
    new_n20243_, new_n20244_, new_n20245_, new_n20246_, new_n20247_,
    new_n20248_, new_n20249_, new_n20250_, new_n20251_, new_n20252_,
    new_n20253_, new_n20254_, new_n20255_, new_n20256_, new_n20257_,
    new_n20258_, new_n20259_, new_n20260_, new_n20261_, new_n20262_,
    new_n20263_, new_n20264_, new_n20265_, new_n20266_, new_n20267_,
    new_n20268_, new_n20269_, new_n20270_, new_n20271_, new_n20272_,
    new_n20273_, new_n20274_, new_n20275_, new_n20276_, new_n20277_,
    new_n20278_, new_n20279_, new_n20280_, new_n20281_, new_n20282_,
    new_n20283_, new_n20284_, new_n20285_, new_n20286_, new_n20287_,
    new_n20288_, new_n20289_, new_n20290_, new_n20291_, new_n20292_,
    new_n20293_, new_n20294_, new_n20295_, new_n20296_, new_n20297_,
    new_n20298_, new_n20299_, new_n20300_, new_n20301_, new_n20302_,
    new_n20303_, new_n20304_, new_n20305_, new_n20306_, new_n20307_,
    new_n20308_, new_n20309_, new_n20310_, new_n20311_, new_n20312_,
    new_n20313_, new_n20314_, new_n20315_, new_n20316_, new_n20317_,
    new_n20318_, new_n20319_, new_n20320_, new_n20321_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20350_, new_n20351_, new_n20352_,
    new_n20353_, new_n20354_, new_n20355_, new_n20356_, new_n20357_,
    new_n20358_, new_n20359_, new_n20360_, new_n20361_, new_n20362_,
    new_n20363_, new_n20364_, new_n20365_, new_n20366_, new_n20367_,
    new_n20368_, new_n20369_, new_n20370_, new_n20371_, new_n20372_,
    new_n20373_, new_n20374_, new_n20375_, new_n20376_, new_n20377_,
    new_n20378_, new_n20379_, new_n20380_, new_n20381_, new_n20382_,
    new_n20383_, new_n20384_, new_n20385_, new_n20386_, new_n20387_,
    new_n20388_, new_n20389_, new_n20390_, new_n20391_, new_n20392_,
    new_n20393_, new_n20394_, new_n20395_, new_n20396_, new_n20397_,
    new_n20398_, new_n20399_, new_n20400_, new_n20401_, new_n20402_,
    new_n20403_, new_n20404_, new_n20405_, new_n20406_, new_n20407_,
    new_n20408_, new_n20409_, new_n20410_, new_n20411_, new_n20412_,
    new_n20413_, new_n20414_, new_n20415_, new_n20416_, new_n20417_,
    new_n20418_, new_n20419_, new_n20420_, new_n20421_, new_n20422_,
    new_n20423_, new_n20424_, new_n20425_, new_n20426_, new_n20427_,
    new_n20428_, new_n20429_, new_n20430_, new_n20431_, new_n20432_,
    new_n20433_, new_n20434_, new_n20435_, new_n20436_, new_n20437_,
    new_n20438_, new_n20439_, new_n20440_, new_n20441_, new_n20442_,
    new_n20443_, new_n20444_, new_n20445_, new_n20446_, new_n20447_,
    new_n20448_, new_n20449_, new_n20450_, new_n20451_, new_n20452_,
    new_n20453_, new_n20454_, new_n20455_, new_n20456_, new_n20457_,
    new_n20458_, new_n20459_, new_n20460_, new_n20461_, new_n20462_,
    new_n20463_, new_n20464_, new_n20465_, new_n20466_, new_n20467_,
    new_n20468_, new_n20469_, new_n20470_, new_n20471_, new_n20472_,
    new_n20473_, new_n20474_, new_n20475_, new_n20476_, new_n20477_,
    new_n20478_, new_n20479_, new_n20480_, new_n20481_, new_n20482_,
    new_n20483_, new_n20484_, new_n20485_, new_n20486_, new_n20487_,
    new_n20488_, new_n20489_, new_n20490_, new_n20491_, new_n20492_,
    new_n20493_, new_n20494_, new_n20495_, new_n20496_, new_n20497_,
    new_n20498_, new_n20499_, new_n20500_, new_n20501_, new_n20502_,
    new_n20503_, new_n20504_, new_n20505_, new_n20506_, new_n20507_,
    new_n20508_, new_n20509_, new_n20510_, new_n20511_, new_n20512_,
    new_n20513_, new_n20514_, new_n20515_, new_n20516_, new_n20517_,
    new_n20518_, new_n20519_, new_n20520_, new_n20521_, new_n20522_,
    new_n20523_, new_n20524_, new_n20525_, new_n20526_, new_n20527_,
    new_n20528_, new_n20529_, new_n20530_, new_n20531_, new_n20532_,
    new_n20533_, new_n20534_, new_n20535_, new_n20536_, new_n20537_,
    new_n20538_, new_n20539_, new_n20540_, new_n20541_, new_n20542_,
    new_n20543_, new_n20544_, new_n20545_, new_n20546_, new_n20547_,
    new_n20548_, new_n20549_, new_n20550_, new_n20551_, new_n20552_,
    new_n20553_, new_n20554_, new_n20555_, new_n20556_, new_n20557_,
    new_n20558_, new_n20559_, new_n20560_, new_n20561_, new_n20562_,
    new_n20563_, new_n20564_, new_n20565_, new_n20566_, new_n20567_,
    new_n20568_, new_n20569_, new_n20570_, new_n20571_, new_n20572_,
    new_n20573_, new_n20574_, new_n20575_, new_n20576_, new_n20577_,
    new_n20578_, new_n20579_, new_n20580_, new_n20581_, new_n20582_,
    new_n20583_, new_n20584_, new_n20585_, new_n20586_, new_n20587_,
    new_n20588_, new_n20589_, new_n20590_, new_n20591_, new_n20592_,
    new_n20593_, new_n20594_, new_n20595_, new_n20596_, new_n20597_,
    new_n20598_, new_n20599_, new_n20600_, new_n20601_, new_n20602_,
    new_n20603_, new_n20604_, new_n20605_, new_n20606_, new_n20607_,
    new_n20608_, new_n20609_, new_n20610_, new_n20611_, new_n20612_,
    new_n20613_, new_n20614_, new_n20615_, new_n20616_, new_n20617_,
    new_n20618_, new_n20619_, new_n20620_, new_n20621_, new_n20622_,
    new_n20623_, new_n20624_, new_n20625_, new_n20626_, new_n20627_,
    new_n20628_, new_n20629_, new_n20630_, new_n20631_, new_n20632_,
    new_n20633_, new_n20634_, new_n20635_, new_n20636_, new_n20637_,
    new_n20638_, new_n20639_, new_n20640_, new_n20641_, new_n20642_,
    new_n20643_, new_n20644_, new_n20645_, new_n20646_, new_n20647_,
    new_n20648_, new_n20649_, new_n20650_, new_n20651_, new_n20652_,
    new_n20653_, new_n20654_, new_n20655_, new_n20656_, new_n20657_,
    new_n20658_, new_n20659_, new_n20660_, new_n20661_, new_n20662_,
    new_n20663_, new_n20664_, new_n20665_, new_n20666_, new_n20667_,
    new_n20668_, new_n20669_, new_n20670_, new_n20671_, new_n20672_,
    new_n20673_, new_n20674_, new_n20675_, new_n20676_, new_n20677_,
    new_n20678_, new_n20679_, new_n20680_, new_n20681_, new_n20682_,
    new_n20683_, new_n20684_, new_n20685_, new_n20686_, new_n20687_,
    new_n20688_, new_n20689_, new_n20690_, new_n20691_, new_n20692_,
    new_n20693_, new_n20694_, new_n20695_, new_n20696_, new_n20697_,
    new_n20698_, new_n20699_, new_n20700_, new_n20701_, new_n20702_,
    new_n20703_, new_n20704_, new_n20705_, new_n20706_, new_n20707_,
    new_n20708_, new_n20709_, new_n20710_, new_n20711_, new_n20712_,
    new_n20713_, new_n20714_, new_n20715_, new_n20716_, new_n20717_,
    new_n20718_, new_n20719_, new_n20720_, new_n20721_, new_n20722_,
    new_n20723_, new_n20724_, new_n20725_, new_n20726_, new_n20727_,
    new_n20728_, new_n20729_, new_n20730_, new_n20731_, new_n20732_,
    new_n20733_, new_n20734_, new_n20735_, new_n20736_, new_n20737_,
    new_n20738_, new_n20739_, new_n20740_, new_n20741_, new_n20742_,
    new_n20743_, new_n20744_, new_n20745_, new_n20746_, new_n20747_,
    new_n20748_, new_n20749_, new_n20750_, new_n20751_, new_n20752_,
    new_n20753_, new_n20754_, new_n20755_, new_n20756_, new_n20757_,
    new_n20758_, new_n20759_, new_n20760_, new_n20761_, new_n20762_,
    new_n20763_, new_n20764_, new_n20765_, new_n20766_, new_n20767_,
    new_n20768_, new_n20769_, new_n20770_, new_n20771_, new_n20772_,
    new_n20773_, new_n20774_, new_n20775_, new_n20776_, new_n20777_,
    new_n20778_, new_n20779_, new_n20780_, new_n20781_, new_n20782_,
    new_n20783_, new_n20784_, new_n20785_, new_n20786_, new_n20787_,
    new_n20788_, new_n20789_, new_n20790_, new_n20791_, new_n20792_,
    new_n20793_, new_n20794_, new_n20795_, new_n20796_, new_n20797_,
    new_n20798_, new_n20799_, new_n20800_, new_n20801_, new_n20802_,
    new_n20803_, new_n20804_, new_n20805_, new_n20806_, new_n20807_,
    new_n20808_, new_n20809_, new_n20810_, new_n20811_, new_n20812_,
    new_n20813_, new_n20814_, new_n20815_, new_n20816_, new_n20817_,
    new_n20818_, new_n20819_, new_n20820_, new_n20821_, new_n20822_,
    new_n20823_, new_n20824_, new_n20825_, new_n20826_, new_n20827_,
    new_n20828_, new_n20829_, new_n20830_, new_n20831_, new_n20832_,
    new_n20833_, new_n20834_, new_n20835_, new_n20836_, new_n20837_,
    new_n20838_, new_n20839_, new_n20840_, new_n20841_, new_n20842_,
    new_n20843_, new_n20844_, new_n20845_, new_n20846_, new_n20847_,
    new_n20848_, new_n20849_, new_n20850_, new_n20851_, new_n20852_,
    new_n20853_, new_n20854_, new_n20855_, new_n20856_, new_n20857_,
    new_n20858_, new_n20859_, new_n20860_, new_n20861_, new_n20862_,
    new_n20863_, new_n20864_, new_n20865_, new_n20866_, new_n20867_,
    new_n20868_, new_n20869_, new_n20870_, new_n20871_, new_n20872_,
    new_n20873_, new_n20874_, new_n20875_, new_n20876_, new_n20877_,
    new_n20878_, new_n20880_, new_n20881_, new_n20882_, new_n20883_,
    new_n20884_, new_n20885_, new_n20886_, new_n20887_, new_n20888_,
    new_n20889_, new_n20890_, new_n20891_, new_n20892_, new_n20893_,
    new_n20894_, new_n20895_, new_n20896_, new_n20897_, new_n20898_,
    new_n20899_, new_n20900_, new_n20901_, new_n20902_, new_n20903_,
    new_n20904_, new_n20905_, new_n20906_, new_n20907_, new_n20908_,
    new_n20909_, new_n20910_, new_n20911_, new_n20912_, new_n20913_,
    new_n20914_, new_n20915_, new_n20916_, new_n20917_, new_n20918_,
    new_n20919_, new_n20920_, new_n20921_, new_n20922_, new_n20923_,
    new_n20924_, new_n20925_, new_n20926_, new_n20927_, new_n20928_,
    new_n20929_, new_n20930_, new_n20931_, new_n20932_, new_n20933_,
    new_n20934_, new_n20935_, new_n20936_, new_n20937_, new_n20938_,
    new_n20939_, new_n20940_, new_n20941_, new_n20942_, new_n20943_,
    new_n20944_, new_n20945_, new_n20946_, new_n20947_, new_n20948_,
    new_n20949_, new_n20950_, new_n20951_, new_n20952_, new_n20953_,
    new_n20954_, new_n20955_, new_n20956_, new_n20957_, new_n20958_,
    new_n20959_, new_n20960_, new_n20961_, new_n20962_, new_n20963_,
    new_n20964_, new_n20965_, new_n20966_, new_n20967_, new_n20968_,
    new_n20969_, new_n20970_, new_n20971_, new_n20972_, new_n20973_,
    new_n20974_, new_n20975_, new_n20976_, new_n20977_, new_n20978_,
    new_n20979_, new_n20980_, new_n20981_, new_n20982_, new_n20983_,
    new_n20984_, new_n20985_, new_n20986_, new_n20987_, new_n20988_,
    new_n20989_, new_n20990_, new_n20991_, new_n20992_, new_n20993_,
    new_n20994_, new_n20995_, new_n20996_, new_n20997_, new_n20998_,
    new_n20999_, new_n21000_, new_n21001_, new_n21002_, new_n21003_,
    new_n21004_, new_n21005_, new_n21006_, new_n21007_, new_n21008_,
    new_n21009_, new_n21010_, new_n21011_, new_n21012_, new_n21013_,
    new_n21014_, new_n21015_, new_n21016_, new_n21017_, new_n21018_,
    new_n21019_, new_n21020_, new_n21021_, new_n21022_, new_n21023_,
    new_n21024_, new_n21025_, new_n21026_, new_n21027_, new_n21028_,
    new_n21029_, new_n21030_, new_n21031_, new_n21032_, new_n21033_,
    new_n21034_, new_n21035_, new_n21036_, new_n21037_, new_n21038_,
    new_n21039_, new_n21040_, new_n21041_, new_n21042_, new_n21043_,
    new_n21044_, new_n21045_, new_n21046_, new_n21047_, new_n21048_,
    new_n21049_, new_n21050_, new_n21051_, new_n21052_, new_n21053_,
    new_n21054_, new_n21055_, new_n21056_, new_n21057_, new_n21058_,
    new_n21059_, new_n21060_, new_n21061_, new_n21062_, new_n21063_,
    new_n21064_, new_n21065_, new_n21066_, new_n21067_, new_n21068_,
    new_n21069_, new_n21070_, new_n21071_, new_n21072_, new_n21073_,
    new_n21074_, new_n21075_, new_n21076_, new_n21077_, new_n21078_,
    new_n21079_, new_n21080_, new_n21081_, new_n21082_, new_n21083_,
    new_n21084_, new_n21085_, new_n21086_, new_n21087_, new_n21088_,
    new_n21089_, new_n21090_, new_n21091_, new_n21092_, new_n21093_,
    new_n21094_, new_n21095_, new_n21096_, new_n21097_, new_n21098_,
    new_n21099_, new_n21100_, new_n21101_, new_n21102_, new_n21103_,
    new_n21104_, new_n21105_, new_n21106_, new_n21107_, new_n21108_,
    new_n21109_, new_n21110_, new_n21111_, new_n21112_, new_n21113_,
    new_n21114_, new_n21115_, new_n21116_, new_n21117_, new_n21118_,
    new_n21119_, new_n21120_, new_n21121_, new_n21122_, new_n21123_,
    new_n21124_, new_n21125_, new_n21126_, new_n21127_, new_n21128_,
    new_n21129_, new_n21130_, new_n21131_, new_n21132_, new_n21133_,
    new_n21134_, new_n21135_, new_n21136_, new_n21137_, new_n21138_,
    new_n21139_, new_n21140_, new_n21141_, new_n21142_, new_n21143_,
    new_n21144_, new_n21145_, new_n21146_, new_n21147_, new_n21148_,
    new_n21149_, new_n21150_, new_n21151_, new_n21152_, new_n21153_,
    new_n21154_, new_n21155_, new_n21156_, new_n21157_, new_n21158_,
    new_n21159_, new_n21160_, new_n21161_, new_n21162_, new_n21163_,
    new_n21164_, new_n21165_, new_n21166_, new_n21167_, new_n21168_,
    new_n21169_, new_n21170_, new_n21171_, new_n21172_, new_n21173_,
    new_n21174_, new_n21175_, new_n21176_, new_n21177_, new_n21178_,
    new_n21179_, new_n21180_, new_n21181_, new_n21182_, new_n21183_,
    new_n21184_, new_n21185_, new_n21186_, new_n21187_, new_n21188_,
    new_n21189_, new_n21190_, new_n21191_, new_n21192_, new_n21193_,
    new_n21194_, new_n21195_, new_n21196_, new_n21197_, new_n21198_,
    new_n21199_, new_n21200_, new_n21201_, new_n21202_, new_n21203_,
    new_n21204_, new_n21205_, new_n21206_, new_n21207_, new_n21208_,
    new_n21209_, new_n21210_, new_n21211_, new_n21212_, new_n21213_,
    new_n21214_, new_n21215_, new_n21216_, new_n21217_, new_n21218_,
    new_n21219_, new_n21220_, new_n21221_, new_n21222_, new_n21223_,
    new_n21224_, new_n21225_, new_n21226_, new_n21227_, new_n21228_,
    new_n21229_, new_n21230_, new_n21231_, new_n21232_, new_n21233_,
    new_n21234_, new_n21235_, new_n21236_, new_n21237_, new_n21238_,
    new_n21239_, new_n21240_, new_n21241_, new_n21242_, new_n21243_,
    new_n21244_, new_n21245_, new_n21246_, new_n21247_, new_n21248_,
    new_n21249_, new_n21250_, new_n21251_, new_n21252_, new_n21253_,
    new_n21254_, new_n21255_, new_n21256_, new_n21257_, new_n21258_,
    new_n21259_, new_n21260_, new_n21261_, new_n21262_, new_n21263_,
    new_n21264_, new_n21265_, new_n21266_, new_n21267_, new_n21268_,
    new_n21269_, new_n21270_, new_n21271_, new_n21272_, new_n21273_,
    new_n21274_, new_n21275_, new_n21276_, new_n21277_, new_n21278_,
    new_n21279_, new_n21280_, new_n21281_, new_n21282_, new_n21283_,
    new_n21284_, new_n21285_, new_n21286_, new_n21287_, new_n21288_,
    new_n21289_, new_n21290_, new_n21291_, new_n21292_, new_n21293_,
    new_n21294_, new_n21295_, new_n21296_, new_n21297_, new_n21298_,
    new_n21299_, new_n21300_, new_n21301_, new_n21302_, new_n21303_,
    new_n21304_, new_n21305_, new_n21306_, new_n21307_, new_n21308_,
    new_n21309_, new_n21310_, new_n21311_, new_n21312_, new_n21313_,
    new_n21314_, new_n21315_, new_n21316_, new_n21317_, new_n21318_,
    new_n21319_, new_n21320_, new_n21321_, new_n21322_, new_n21323_,
    new_n21324_, new_n21325_, new_n21326_, new_n21327_, new_n21328_,
    new_n21329_, new_n21330_, new_n21331_, new_n21332_, new_n21333_,
    new_n21334_, new_n21335_, new_n21336_, new_n21337_, new_n21338_,
    new_n21339_, new_n21340_, new_n21341_, new_n21342_, new_n21343_,
    new_n21344_, new_n21345_, new_n21346_, new_n21347_, new_n21348_,
    new_n21349_, new_n21350_, new_n21351_, new_n21352_, new_n21353_,
    new_n21354_, new_n21355_, new_n21356_, new_n21357_, new_n21358_,
    new_n21359_, new_n21360_, new_n21361_, new_n21362_, new_n21363_,
    new_n21364_, new_n21365_, new_n21366_, new_n21367_, new_n21368_,
    new_n21369_, new_n21370_, new_n21371_, new_n21372_, new_n21373_,
    new_n21374_, new_n21375_, new_n21376_, new_n21377_, new_n21378_,
    new_n21379_, new_n21380_, new_n21381_, new_n21382_, new_n21383_,
    new_n21384_, new_n21385_, new_n21386_, new_n21387_, new_n21388_,
    new_n21389_, new_n21390_, new_n21391_, new_n21392_, new_n21393_,
    new_n21394_, new_n21395_, new_n21396_, new_n21397_, new_n21398_,
    new_n21399_, new_n21400_, new_n21401_, new_n21402_, new_n21403_,
    new_n21404_, new_n21405_, new_n21406_, new_n21407_, new_n21408_,
    new_n21409_, new_n21410_, new_n21411_, new_n21412_, new_n21413_,
    new_n21414_, new_n21415_, new_n21416_, new_n21417_, new_n21418_,
    new_n21419_, new_n21420_, new_n21421_, new_n21422_, new_n21423_,
    new_n21424_, new_n21425_, new_n21426_, new_n21427_, new_n21428_,
    new_n21429_, new_n21430_, new_n21431_, new_n21432_, new_n21433_,
    new_n21434_, new_n21435_, new_n21436_, new_n21437_, new_n21438_,
    new_n21439_, new_n21440_, new_n21441_, new_n21442_, new_n21443_,
    new_n21444_, new_n21445_, new_n21446_, new_n21447_, new_n21448_,
    new_n21449_, new_n21450_, new_n21451_, new_n21452_, new_n21453_,
    new_n21454_, new_n21455_, new_n21456_, new_n21457_, new_n21458_,
    new_n21459_, new_n21460_, new_n21461_, new_n21462_, new_n21463_,
    new_n21464_, new_n21465_, new_n21466_, new_n21467_, new_n21468_,
    new_n21469_, new_n21470_, new_n21471_, new_n21472_, new_n21473_,
    new_n21474_, new_n21475_, new_n21476_, new_n21477_, new_n21478_,
    new_n21479_, new_n21480_, new_n21481_, new_n21482_, new_n21483_,
    new_n21484_, new_n21485_, new_n21486_, new_n21487_, new_n21488_,
    new_n21489_, new_n21490_, new_n21491_, new_n21492_, new_n21493_,
    new_n21494_, new_n21495_, new_n21496_, new_n21497_, new_n21498_,
    new_n21499_, new_n21500_, new_n21501_, new_n21502_, new_n21503_,
    new_n21504_, new_n21505_, new_n21506_, new_n21507_, new_n21508_,
    new_n21509_, new_n21510_, new_n21511_, new_n21512_, new_n21513_,
    new_n21514_, new_n21515_, new_n21516_, new_n21517_, new_n21518_,
    new_n21519_, new_n21520_, new_n21521_, new_n21522_, new_n21523_,
    new_n21524_, new_n21525_, new_n21526_, new_n21527_, new_n21528_,
    new_n21529_, new_n21530_, new_n21531_, new_n21532_, new_n21533_,
    new_n21534_, new_n21535_, new_n21536_, new_n21537_, new_n21538_,
    new_n21539_, new_n21540_, new_n21541_, new_n21542_, new_n21543_,
    new_n21544_, new_n21545_, new_n21546_, new_n21547_, new_n21548_,
    new_n21549_, new_n21550_, new_n21551_, new_n21552_, new_n21553_,
    new_n21554_, new_n21555_, new_n21556_, new_n21557_, new_n21558_,
    new_n21559_, new_n21560_, new_n21562_, new_n21563_, new_n21564_,
    new_n21565_, new_n21566_, new_n21567_, new_n21568_, new_n21569_,
    new_n21570_, new_n21571_, new_n21572_, new_n21573_, new_n21574_,
    new_n21575_, new_n21576_, new_n21577_, new_n21578_, new_n21579_,
    new_n21580_, new_n21581_, new_n21582_, new_n21583_, new_n21584_,
    new_n21585_, new_n21586_, new_n21587_, new_n21588_, new_n21589_,
    new_n21590_, new_n21591_, new_n21592_, new_n21593_, new_n21594_,
    new_n21595_, new_n21596_, new_n21597_, new_n21598_, new_n21599_,
    new_n21600_, new_n21601_, new_n21602_, new_n21603_, new_n21604_,
    new_n21605_, new_n21606_, new_n21607_, new_n21608_, new_n21609_,
    new_n21610_, new_n21611_, new_n21612_, new_n21613_, new_n21614_,
    new_n21615_, new_n21616_, new_n21617_, new_n21618_, new_n21619_,
    new_n21620_, new_n21621_, new_n21622_, new_n21623_, new_n21624_,
    new_n21625_, new_n21626_, new_n21627_, new_n21628_, new_n21629_,
    new_n21630_, new_n21631_, new_n21632_, new_n21633_, new_n21634_,
    new_n21635_, new_n21636_, new_n21637_, new_n21638_, new_n21639_,
    new_n21640_, new_n21641_, new_n21642_, new_n21643_, new_n21644_,
    new_n21645_, new_n21646_, new_n21647_, new_n21648_, new_n21649_,
    new_n21650_, new_n21651_, new_n21652_, new_n21653_, new_n21654_,
    new_n21655_, new_n21656_, new_n21657_, new_n21658_, new_n21659_,
    new_n21660_, new_n21661_, new_n21662_, new_n21663_, new_n21664_,
    new_n21665_, new_n21666_, new_n21667_, new_n21668_, new_n21669_,
    new_n21670_, new_n21671_, new_n21672_, new_n21673_, new_n21674_,
    new_n21675_, new_n21676_, new_n21677_, new_n21678_, new_n21679_,
    new_n21680_, new_n21681_, new_n21682_, new_n21683_, new_n21684_,
    new_n21685_, new_n21686_, new_n21687_, new_n21688_, new_n21689_,
    new_n21690_, new_n21691_, new_n21692_, new_n21693_, new_n21694_,
    new_n21695_, new_n21696_, new_n21697_, new_n21698_, new_n21699_,
    new_n21700_, new_n21701_, new_n21702_, new_n21703_, new_n21704_,
    new_n21705_, new_n21706_, new_n21707_, new_n21708_, new_n21709_,
    new_n21710_, new_n21711_, new_n21712_, new_n21713_, new_n21714_,
    new_n21715_, new_n21716_, new_n21717_, new_n21718_, new_n21719_,
    new_n21720_, new_n21721_, new_n21722_, new_n21723_, new_n21724_,
    new_n21725_, new_n21726_, new_n21727_, new_n21728_, new_n21729_,
    new_n21730_, new_n21731_, new_n21732_, new_n21733_, new_n21734_,
    new_n21735_, new_n21736_, new_n21737_, new_n21738_, new_n21739_,
    new_n21740_, new_n21741_, new_n21742_, new_n21743_, new_n21744_,
    new_n21745_, new_n21746_, new_n21747_, new_n21748_, new_n21749_,
    new_n21750_, new_n21751_, new_n21752_, new_n21753_, new_n21754_,
    new_n21755_, new_n21756_, new_n21757_, new_n21758_, new_n21759_,
    new_n21760_, new_n21761_, new_n21762_, new_n21763_, new_n21764_,
    new_n21765_, new_n21766_, new_n21767_, new_n21768_, new_n21769_,
    new_n21770_, new_n21771_, new_n21772_, new_n21773_, new_n21774_,
    new_n21775_, new_n21776_, new_n21777_, new_n21778_, new_n21779_,
    new_n21780_, new_n21781_, new_n21782_, new_n21783_, new_n21784_,
    new_n21785_, new_n21786_, new_n21787_, new_n21788_, new_n21789_,
    new_n21790_, new_n21791_, new_n21792_, new_n21793_, new_n21794_,
    new_n21795_, new_n21796_, new_n21797_, new_n21798_, new_n21799_,
    new_n21800_, new_n21801_, new_n21802_, new_n21803_, new_n21804_,
    new_n21805_, new_n21806_, new_n21807_, new_n21808_, new_n21809_,
    new_n21810_, new_n21811_, new_n21812_, new_n21813_, new_n21814_,
    new_n21815_, new_n21816_, new_n21817_, new_n21818_, new_n21819_,
    new_n21820_, new_n21821_, new_n21822_, new_n21823_, new_n21824_,
    new_n21825_, new_n21826_, new_n21827_, new_n21828_, new_n21829_,
    new_n21830_, new_n21831_, new_n21832_, new_n21833_, new_n21834_,
    new_n21835_, new_n21836_, new_n21837_, new_n21838_, new_n21839_,
    new_n21840_, new_n21841_, new_n21842_, new_n21843_, new_n21844_,
    new_n21845_, new_n21846_, new_n21847_, new_n21848_, new_n21849_,
    new_n21850_, new_n21851_, new_n21852_, new_n21853_, new_n21854_,
    new_n21855_, new_n21856_, new_n21857_, new_n21858_, new_n21859_,
    new_n21860_, new_n21861_, new_n21862_, new_n21863_, new_n21864_,
    new_n21865_, new_n21866_, new_n21867_, new_n21868_, new_n21869_,
    new_n21870_, new_n21871_, new_n21872_, new_n21873_, new_n21874_,
    new_n21875_, new_n21876_, new_n21877_, new_n21878_, new_n21879_,
    new_n21880_, new_n21881_, new_n21882_, new_n21883_, new_n21884_,
    new_n21885_, new_n21886_, new_n21887_, new_n21888_, new_n21889_,
    new_n21890_, new_n21891_, new_n21892_, new_n21893_, new_n21894_,
    new_n21895_, new_n21896_, new_n21897_, new_n21898_, new_n21899_,
    new_n21900_, new_n21901_, new_n21902_, new_n21903_, new_n21904_,
    new_n21905_, new_n21906_, new_n21907_, new_n21908_, new_n21909_,
    new_n21910_, new_n21911_, new_n21912_, new_n21913_, new_n21914_,
    new_n21915_, new_n21916_, new_n21917_, new_n21918_, new_n21919_,
    new_n21920_, new_n21921_, new_n21922_, new_n21923_, new_n21924_,
    new_n21925_, new_n21926_, new_n21927_, new_n21928_, new_n21929_,
    new_n21930_, new_n21931_, new_n21932_, new_n21933_, new_n21934_,
    new_n21935_, new_n21936_, new_n21937_, new_n21938_, new_n21939_,
    new_n21940_, new_n21941_, new_n21942_, new_n21943_, new_n21944_,
    new_n21945_, new_n21946_, new_n21947_, new_n21948_, new_n21949_,
    new_n21950_, new_n21951_, new_n21952_, new_n21953_, new_n21954_,
    new_n21955_, new_n21956_, new_n21957_, new_n21958_, new_n21959_,
    new_n21960_, new_n21961_, new_n21962_, new_n21963_, new_n21964_,
    new_n21965_, new_n21966_, new_n21967_, new_n21968_, new_n21969_,
    new_n21970_, new_n21971_, new_n21972_, new_n21973_, new_n21974_,
    new_n21975_, new_n21976_, new_n21977_, new_n21978_, new_n21979_,
    new_n21980_, new_n21981_, new_n21982_, new_n21983_, new_n21984_,
    new_n21985_, new_n21986_, new_n21987_, new_n21988_, new_n21989_,
    new_n21990_, new_n21991_, new_n21992_, new_n21993_, new_n21994_,
    new_n21995_, new_n21996_, new_n21997_, new_n21998_, new_n21999_,
    new_n22000_, new_n22001_, new_n22002_, new_n22003_, new_n22004_,
    new_n22005_, new_n22006_, new_n22007_, new_n22008_, new_n22009_,
    new_n22010_, new_n22011_, new_n22012_, new_n22013_, new_n22014_,
    new_n22015_, new_n22016_, new_n22017_, new_n22018_, new_n22019_,
    new_n22020_, new_n22021_, new_n22022_, new_n22023_, new_n22024_,
    new_n22025_, new_n22026_, new_n22027_, new_n22028_, new_n22029_,
    new_n22030_, new_n22031_, new_n22032_, new_n22033_, new_n22034_,
    new_n22035_, new_n22036_, new_n22037_, new_n22038_, new_n22039_,
    new_n22040_, new_n22041_, new_n22042_, new_n22043_, new_n22044_,
    new_n22045_, new_n22046_, new_n22047_, new_n22048_, new_n22049_,
    new_n22050_, new_n22051_, new_n22052_, new_n22053_, new_n22054_,
    new_n22055_, new_n22056_, new_n22057_, new_n22058_, new_n22059_,
    new_n22060_, new_n22061_, new_n22062_, new_n22063_, new_n22064_,
    new_n22065_, new_n22066_, new_n22067_, new_n22068_, new_n22069_,
    new_n22070_, new_n22071_, new_n22072_, new_n22073_, new_n22074_,
    new_n22075_, new_n22076_, new_n22077_, new_n22078_, new_n22079_,
    new_n22080_, new_n22081_, new_n22082_, new_n22083_, new_n22084_,
    new_n22085_, new_n22086_, new_n22087_, new_n22088_, new_n22089_,
    new_n22090_, new_n22091_, new_n22092_, new_n22093_, new_n22094_,
    new_n22095_, new_n22096_, new_n22097_, new_n22098_, new_n22099_,
    new_n22100_, new_n22101_, new_n22102_, new_n22103_, new_n22104_,
    new_n22105_, new_n22106_, new_n22107_, new_n22108_, new_n22109_,
    new_n22110_, new_n22111_, new_n22112_, new_n22113_, new_n22114_,
    new_n22115_, new_n22116_, new_n22117_, new_n22118_, new_n22119_,
    new_n22120_, new_n22121_, new_n22122_, new_n22123_, new_n22124_,
    new_n22125_, new_n22126_, new_n22127_, new_n22128_, new_n22129_,
    new_n22130_, new_n22131_, new_n22132_, new_n22133_, new_n22134_,
    new_n22135_, new_n22136_, new_n22137_, new_n22138_, new_n22139_,
    new_n22140_, new_n22141_, new_n22142_, new_n22143_, new_n22144_,
    new_n22145_, new_n22146_, new_n22147_, new_n22148_, new_n22149_,
    new_n22150_, new_n22151_, new_n22152_, new_n22153_, new_n22154_,
    new_n22155_, new_n22156_, new_n22157_, new_n22158_, new_n22159_,
    new_n22160_, new_n22161_, new_n22162_, new_n22163_, new_n22164_,
    new_n22165_, new_n22166_, new_n22167_, new_n22168_, new_n22169_,
    new_n22170_, new_n22171_, new_n22172_, new_n22173_, new_n22174_,
    new_n22175_, new_n22176_, new_n22177_, new_n22178_, new_n22179_,
    new_n22180_, new_n22181_, new_n22182_, new_n22183_, new_n22184_,
    new_n22185_, new_n22186_, new_n22187_, new_n22188_, new_n22189_,
    new_n22190_, new_n22191_, new_n22192_, new_n22193_, new_n22194_,
    new_n22195_, new_n22196_, new_n22197_, new_n22198_, new_n22199_,
    new_n22200_, new_n22201_, new_n22202_, new_n22203_, new_n22204_,
    new_n22205_, new_n22206_, new_n22207_, new_n22208_, new_n22209_,
    new_n22210_, new_n22211_, new_n22212_, new_n22213_, new_n22214_,
    new_n22215_, new_n22216_, new_n22217_, new_n22218_, new_n22219_,
    new_n22220_, new_n22221_, new_n22222_, new_n22223_, new_n22224_,
    new_n22225_, new_n22226_, new_n22227_, new_n22228_, new_n22229_,
    new_n22230_, new_n22231_, new_n22232_, new_n22233_, new_n22234_,
    new_n22235_, new_n22236_, new_n22237_, new_n22238_, new_n22239_,
    new_n22240_, new_n22241_, new_n22242_, new_n22243_, new_n22244_,
    new_n22245_, new_n22246_, new_n22247_, new_n22248_, new_n22249_,
    new_n22250_, new_n22251_, new_n22252_, new_n22253_, new_n22254_,
    new_n22255_, new_n22256_, new_n22257_, new_n22258_, new_n22259_,
    new_n22260_, new_n22261_, new_n22262_, new_n22263_, new_n22264_,
    new_n22265_, new_n22266_, new_n22267_, new_n22268_, new_n22269_,
    new_n22270_, new_n22271_, new_n22272_, new_n22273_, new_n22274_,
    new_n22275_, new_n22276_, new_n22277_, new_n22278_, new_n22279_,
    new_n22280_, new_n22281_, new_n22282_, new_n22283_, new_n22284_,
    new_n22285_, new_n22286_, new_n22287_, new_n22288_, new_n22290_,
    new_n22291_, new_n22292_, new_n22293_, new_n22294_, new_n22295_,
    new_n22296_, new_n22297_, new_n22298_, new_n22299_, new_n22300_,
    new_n22301_, new_n22302_, new_n22303_, new_n22304_, new_n22305_,
    new_n22306_, new_n22307_, new_n22308_, new_n22309_, new_n22310_,
    new_n22311_, new_n22312_, new_n22313_, new_n22314_, new_n22315_,
    new_n22316_, new_n22317_, new_n22318_, new_n22319_, new_n22320_,
    new_n22321_, new_n22322_, new_n22323_, new_n22324_, new_n22325_,
    new_n22326_, new_n22327_, new_n22328_, new_n22329_, new_n22330_,
    new_n22331_, new_n22332_, new_n22333_, new_n22334_, new_n22335_,
    new_n22336_, new_n22337_, new_n22338_, new_n22339_, new_n22340_,
    new_n22341_, new_n22342_, new_n22343_, new_n22344_, new_n22345_,
    new_n22346_, new_n22347_, new_n22348_, new_n22349_, new_n22350_,
    new_n22351_, new_n22352_, new_n22353_, new_n22354_, new_n22355_,
    new_n22356_, new_n22357_, new_n22358_, new_n22359_, new_n22360_,
    new_n22361_, new_n22362_, new_n22363_, new_n22364_, new_n22365_,
    new_n22366_, new_n22367_, new_n22368_, new_n22369_, new_n22370_,
    new_n22371_, new_n22372_, new_n22373_, new_n22374_, new_n22375_,
    new_n22376_, new_n22377_, new_n22378_, new_n22379_, new_n22380_,
    new_n22381_, new_n22382_, new_n22383_, new_n22384_, new_n22385_,
    new_n22386_, new_n22387_, new_n22388_, new_n22389_, new_n22390_,
    new_n22391_, new_n22392_, new_n22393_, new_n22394_, new_n22395_,
    new_n22396_, new_n22397_, new_n22398_, new_n22399_, new_n22400_,
    new_n22401_, new_n22402_, new_n22403_, new_n22404_, new_n22405_,
    new_n22406_, new_n22407_, new_n22408_, new_n22409_, new_n22410_,
    new_n22411_, new_n22412_, new_n22413_, new_n22414_, new_n22415_,
    new_n22416_, new_n22417_, new_n22418_, new_n22419_, new_n22420_,
    new_n22421_, new_n22422_, new_n22423_, new_n22424_, new_n22425_,
    new_n22426_, new_n22427_, new_n22428_, new_n22429_, new_n22430_,
    new_n22431_, new_n22432_, new_n22433_, new_n22434_, new_n22435_,
    new_n22436_, new_n22437_, new_n22438_, new_n22439_, new_n22440_,
    new_n22441_, new_n22442_, new_n22443_, new_n22444_, new_n22445_,
    new_n22446_, new_n22447_, new_n22448_, new_n22449_, new_n22450_,
    new_n22451_, new_n22452_, new_n22453_, new_n22454_, new_n22455_,
    new_n22456_, new_n22457_, new_n22458_, new_n22459_, new_n22460_,
    new_n22461_, new_n22462_, new_n22463_, new_n22464_, new_n22465_,
    new_n22466_, new_n22467_, new_n22468_, new_n22469_, new_n22470_,
    new_n22471_, new_n22472_, new_n22473_, new_n22474_, new_n22475_,
    new_n22476_, new_n22477_, new_n22478_, new_n22479_, new_n22480_,
    new_n22481_, new_n22482_, new_n22483_, new_n22484_, new_n22485_,
    new_n22486_, new_n22487_, new_n22488_, new_n22489_, new_n22490_,
    new_n22491_, new_n22492_, new_n22493_, new_n22494_, new_n22495_,
    new_n22496_, new_n22497_, new_n22498_, new_n22499_, new_n22500_,
    new_n22501_, new_n22502_, new_n22503_, new_n22504_, new_n22505_,
    new_n22506_, new_n22507_, new_n22508_, new_n22509_, new_n22510_,
    new_n22511_, new_n22512_, new_n22513_, new_n22514_, new_n22515_,
    new_n22516_, new_n22517_, new_n22518_, new_n22519_, new_n22520_,
    new_n22521_, new_n22522_, new_n22523_, new_n22524_, new_n22525_,
    new_n22526_, new_n22527_, new_n22528_, new_n22529_, new_n22530_,
    new_n22531_, new_n22532_, new_n22533_, new_n22534_, new_n22535_,
    new_n22536_, new_n22537_, new_n22538_, new_n22539_, new_n22540_,
    new_n22541_, new_n22542_, new_n22543_, new_n22544_, new_n22545_,
    new_n22546_, new_n22547_, new_n22548_, new_n22549_, new_n22550_,
    new_n22551_, new_n22552_, new_n22553_, new_n22554_, new_n22555_,
    new_n22556_, new_n22557_, new_n22558_, new_n22559_, new_n22560_,
    new_n22561_, new_n22562_, new_n22563_, new_n22564_, new_n22565_,
    new_n22566_, new_n22567_, new_n22568_, new_n22569_, new_n22570_,
    new_n22571_, new_n22572_, new_n22573_, new_n22574_, new_n22575_,
    new_n22576_, new_n22577_, new_n22578_, new_n22579_, new_n22580_,
    new_n22581_, new_n22582_, new_n22583_, new_n22584_, new_n22585_,
    new_n22586_, new_n22587_, new_n22588_, new_n22589_, new_n22590_,
    new_n22591_, new_n22592_, new_n22593_, new_n22594_, new_n22595_,
    new_n22596_, new_n22597_, new_n22598_, new_n22599_, new_n22600_,
    new_n22601_, new_n22602_, new_n22603_, new_n22604_, new_n22605_,
    new_n22606_, new_n22607_, new_n22608_, new_n22609_, new_n22610_,
    new_n22611_, new_n22612_, new_n22613_, new_n22614_, new_n22615_,
    new_n22616_, new_n22617_, new_n22618_, new_n22619_, new_n22620_,
    new_n22621_, new_n22622_, new_n22623_, new_n22624_, new_n22625_,
    new_n22626_, new_n22627_, new_n22628_, new_n22629_, new_n22630_,
    new_n22631_, new_n22632_, new_n22633_, new_n22634_, new_n22635_,
    new_n22636_, new_n22637_, new_n22638_, new_n22639_, new_n22640_,
    new_n22641_, new_n22642_, new_n22643_, new_n22644_, new_n22645_,
    new_n22646_, new_n22647_, new_n22648_, new_n22649_, new_n22650_,
    new_n22651_, new_n22652_, new_n22653_, new_n22654_, new_n22655_,
    new_n22656_, new_n22657_, new_n22658_, new_n22659_, new_n22660_,
    new_n22661_, new_n22662_, new_n22663_, new_n22664_, new_n22665_,
    new_n22666_, new_n22667_, new_n22668_, new_n22669_, new_n22670_,
    new_n22671_, new_n22672_, new_n22673_, new_n22674_, new_n22675_,
    new_n22676_, new_n22677_, new_n22678_, new_n22679_, new_n22680_,
    new_n22681_, new_n22682_, new_n22683_, new_n22684_, new_n22685_,
    new_n22686_, new_n22687_, new_n22688_, new_n22689_, new_n22690_,
    new_n22691_, new_n22692_, new_n22693_, new_n22694_, new_n22695_,
    new_n22696_, new_n22697_, new_n22698_, new_n22699_, new_n22700_,
    new_n22701_, new_n22702_, new_n22703_, new_n22704_, new_n22705_,
    new_n22706_, new_n22707_, new_n22708_, new_n22709_, new_n22710_,
    new_n22711_, new_n22712_, new_n22713_, new_n22714_, new_n22715_,
    new_n22716_, new_n22717_, new_n22718_, new_n22719_, new_n22720_,
    new_n22721_, new_n22722_, new_n22723_, new_n22724_, new_n22725_,
    new_n22726_, new_n22727_, new_n22728_, new_n22729_, new_n22730_,
    new_n22731_, new_n22732_, new_n22733_, new_n22734_, new_n22735_,
    new_n22736_, new_n22737_, new_n22738_, new_n22739_, new_n22740_,
    new_n22741_, new_n22742_, new_n22743_, new_n22744_, new_n22745_,
    new_n22746_, new_n22747_, new_n22748_, new_n22749_, new_n22750_,
    new_n22751_, new_n22752_, new_n22753_, new_n22754_, new_n22755_,
    new_n22756_, new_n22757_, new_n22758_, new_n22759_, new_n22760_,
    new_n22761_, new_n22762_, new_n22763_, new_n22764_, new_n22765_,
    new_n22766_, new_n22767_, new_n22768_, new_n22769_, new_n22770_,
    new_n22771_, new_n22772_, new_n22773_, new_n22774_, new_n22775_,
    new_n22776_, new_n22777_, new_n22778_, new_n22779_, new_n22780_,
    new_n22781_, new_n22782_, new_n22783_, new_n22784_, new_n22785_,
    new_n22786_, new_n22787_, new_n22788_, new_n22789_, new_n22790_,
    new_n22791_, new_n22792_, new_n22793_, new_n22794_, new_n22795_,
    new_n22796_, new_n22797_, new_n22798_, new_n22799_, new_n22800_,
    new_n22801_, new_n22802_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22876_, new_n22877_, new_n22878_, new_n22879_, new_n22880_,
    new_n22881_, new_n22882_, new_n22883_, new_n22884_, new_n22885_,
    new_n22886_, new_n22887_, new_n22888_, new_n22889_, new_n22890_,
    new_n22891_, new_n22892_, new_n22893_, new_n22894_, new_n22895_,
    new_n22896_, new_n22897_, new_n22898_, new_n22899_, new_n22900_,
    new_n22901_, new_n22902_, new_n22903_, new_n22904_, new_n22905_,
    new_n22906_, new_n22907_, new_n22908_, new_n22909_, new_n22910_,
    new_n22911_, new_n22912_, new_n22913_, new_n22914_, new_n22915_,
    new_n22916_, new_n22917_, new_n22918_, new_n22919_, new_n22920_,
    new_n22921_, new_n22922_, new_n22923_, new_n22924_, new_n22925_,
    new_n22926_, new_n22927_, new_n22928_, new_n22929_, new_n22930_,
    new_n22931_, new_n22932_, new_n22933_, new_n22934_, new_n22935_,
    new_n22936_, new_n22937_, new_n22938_, new_n22939_, new_n22940_,
    new_n22941_, new_n22942_, new_n22943_, new_n22944_, new_n22945_,
    new_n22946_, new_n22947_, new_n22948_, new_n22949_, new_n22950_,
    new_n22951_, new_n22952_, new_n22953_, new_n22954_, new_n22955_,
    new_n22956_, new_n22957_, new_n22958_, new_n22959_, new_n22960_,
    new_n22961_, new_n22962_, new_n22963_, new_n22964_, new_n22965_,
    new_n22966_, new_n22967_, new_n22968_, new_n22969_, new_n22970_,
    new_n22971_, new_n22972_, new_n22973_, new_n22974_, new_n22975_,
    new_n22976_, new_n22977_, new_n22978_, new_n22979_, new_n22980_,
    new_n22981_, new_n22982_, new_n22984_, new_n22985_, new_n22986_,
    new_n22987_, new_n22988_, new_n22989_, new_n22990_, new_n22991_,
    new_n22992_, new_n22993_, new_n22994_, new_n22995_, new_n22996_,
    new_n22997_, new_n22998_, new_n22999_, new_n23000_, new_n23001_,
    new_n23002_, new_n23003_, new_n23004_, new_n23005_, new_n23006_,
    new_n23007_, new_n23008_, new_n23009_, new_n23010_, new_n23011_,
    new_n23012_, new_n23013_, new_n23014_, new_n23015_, new_n23016_,
    new_n23017_, new_n23018_, new_n23019_, new_n23020_, new_n23021_,
    new_n23022_, new_n23023_, new_n23024_, new_n23025_, new_n23026_,
    new_n23027_, new_n23028_, new_n23029_, new_n23030_, new_n23031_,
    new_n23032_, new_n23033_, new_n23034_, new_n23035_, new_n23036_,
    new_n23037_, new_n23038_, new_n23039_, new_n23040_, new_n23041_,
    new_n23042_, new_n23043_, new_n23044_, new_n23045_, new_n23046_,
    new_n23047_, new_n23048_, new_n23049_, new_n23050_, new_n23051_,
    new_n23052_, new_n23053_, new_n23054_, new_n23055_, new_n23056_,
    new_n23057_, new_n23058_, new_n23059_, new_n23060_, new_n23061_,
    new_n23062_, new_n23063_, new_n23064_, new_n23065_, new_n23066_,
    new_n23067_, new_n23068_, new_n23069_, new_n23070_, new_n23071_,
    new_n23072_, new_n23073_, new_n23074_, new_n23075_, new_n23076_,
    new_n23077_, new_n23078_, new_n23079_, new_n23080_, new_n23081_,
    new_n23082_, new_n23083_, new_n23084_, new_n23085_, new_n23086_,
    new_n23087_, new_n23088_, new_n23089_, new_n23090_, new_n23091_,
    new_n23092_, new_n23093_, new_n23094_, new_n23095_, new_n23096_,
    new_n23097_, new_n23098_, new_n23099_, new_n23100_, new_n23101_,
    new_n23102_, new_n23103_, new_n23104_, new_n23105_, new_n23106_,
    new_n23107_, new_n23108_, new_n23109_, new_n23110_, new_n23111_,
    new_n23112_, new_n23113_, new_n23114_, new_n23115_, new_n23116_,
    new_n23117_, new_n23118_, new_n23119_, new_n23120_, new_n23121_,
    new_n23122_, new_n23123_, new_n23124_, new_n23125_, new_n23126_,
    new_n23127_, new_n23128_, new_n23129_, new_n23130_, new_n23131_,
    new_n23132_, new_n23133_, new_n23134_, new_n23135_, new_n23136_,
    new_n23137_, new_n23138_, new_n23139_, new_n23140_, new_n23141_,
    new_n23142_, new_n23143_, new_n23144_, new_n23145_, new_n23146_,
    new_n23147_, new_n23148_, new_n23149_, new_n23150_, new_n23151_,
    new_n23152_, new_n23153_, new_n23154_, new_n23155_, new_n23156_,
    new_n23157_, new_n23158_, new_n23159_, new_n23160_, new_n23161_,
    new_n23162_, new_n23163_, new_n23164_, new_n23165_, new_n23166_,
    new_n23167_, new_n23168_, new_n23169_, new_n23170_, new_n23171_,
    new_n23172_, new_n23173_, new_n23174_, new_n23175_, new_n23176_,
    new_n23177_, new_n23178_, new_n23179_, new_n23180_, new_n23181_,
    new_n23182_, new_n23183_, new_n23184_, new_n23185_, new_n23186_,
    new_n23187_, new_n23188_, new_n23189_, new_n23190_, new_n23191_,
    new_n23192_, new_n23193_, new_n23194_, new_n23195_, new_n23196_,
    new_n23197_, new_n23198_, new_n23199_, new_n23200_, new_n23201_,
    new_n23202_, new_n23203_, new_n23204_, new_n23205_, new_n23206_,
    new_n23207_, new_n23208_, new_n23209_, new_n23210_, new_n23211_,
    new_n23212_, new_n23213_, new_n23214_, new_n23215_, new_n23216_,
    new_n23217_, new_n23218_, new_n23219_, new_n23220_, new_n23221_,
    new_n23222_, new_n23223_, new_n23224_, new_n23225_, new_n23226_,
    new_n23227_, new_n23228_, new_n23229_, new_n23230_, new_n23231_,
    new_n23232_, new_n23233_, new_n23234_, new_n23235_, new_n23236_,
    new_n23237_, new_n23238_, new_n23239_, new_n23240_, new_n23241_,
    new_n23242_, new_n23243_, new_n23244_, new_n23245_, new_n23246_,
    new_n23247_, new_n23248_, new_n23249_, new_n23250_, new_n23251_,
    new_n23252_, new_n23253_, new_n23254_, new_n23255_, new_n23256_,
    new_n23257_, new_n23258_, new_n23259_, new_n23260_, new_n23261_,
    new_n23262_, new_n23263_, new_n23264_, new_n23265_, new_n23266_,
    new_n23267_, new_n23268_, new_n23269_, new_n23270_, new_n23271_,
    new_n23272_, new_n23273_, new_n23274_, new_n23275_, new_n23276_,
    new_n23277_, new_n23278_, new_n23279_, new_n23280_, new_n23281_,
    new_n23282_, new_n23283_, new_n23284_, new_n23285_, new_n23286_,
    new_n23287_, new_n23288_, new_n23289_, new_n23290_, new_n23291_,
    new_n23292_, new_n23293_, new_n23294_, new_n23295_, new_n23296_,
    new_n23297_, new_n23298_, new_n23299_, new_n23300_, new_n23301_,
    new_n23302_, new_n23303_, new_n23304_, new_n23305_, new_n23306_,
    new_n23307_, new_n23308_, new_n23309_, new_n23310_, new_n23311_,
    new_n23312_, new_n23313_, new_n23314_, new_n23315_, new_n23316_,
    new_n23317_, new_n23318_, new_n23319_, new_n23320_, new_n23321_,
    new_n23322_, new_n23323_, new_n23324_, new_n23325_, new_n23326_,
    new_n23327_, new_n23328_, new_n23329_, new_n23330_, new_n23331_,
    new_n23332_, new_n23333_, new_n23334_, new_n23335_, new_n23336_,
    new_n23337_, new_n23338_, new_n23339_, new_n23340_, new_n23341_,
    new_n23342_, new_n23343_, new_n23344_, new_n23345_, new_n23346_,
    new_n23347_, new_n23348_, new_n23349_, new_n23350_, new_n23351_,
    new_n23352_, new_n23353_, new_n23354_, new_n23355_, new_n23356_,
    new_n23357_, new_n23358_, new_n23359_, new_n23360_, new_n23361_,
    new_n23362_, new_n23363_, new_n23364_, new_n23365_, new_n23366_,
    new_n23367_, new_n23368_, new_n23369_, new_n23370_, new_n23371_,
    new_n23372_, new_n23373_, new_n23374_, new_n23375_, new_n23376_,
    new_n23377_, new_n23378_, new_n23379_, new_n23380_, new_n23381_,
    new_n23382_, new_n23383_, new_n23384_, new_n23385_, new_n23386_,
    new_n23387_, new_n23388_, new_n23389_, new_n23390_, new_n23391_,
    new_n23392_, new_n23393_, new_n23394_, new_n23395_, new_n23396_,
    new_n23397_, new_n23398_, new_n23399_, new_n23400_, new_n23401_,
    new_n23402_, new_n23403_, new_n23404_, new_n23405_, new_n23406_,
    new_n23407_, new_n23408_, new_n23409_, new_n23410_, new_n23411_,
    new_n23412_, new_n23413_, new_n23414_, new_n23415_, new_n23416_,
    new_n23417_, new_n23418_, new_n23419_, new_n23420_, new_n23421_,
    new_n23422_, new_n23423_, new_n23424_, new_n23425_, new_n23426_,
    new_n23427_, new_n23428_, new_n23429_, new_n23430_, new_n23431_,
    new_n23432_, new_n23433_, new_n23434_, new_n23435_, new_n23436_,
    new_n23437_, new_n23438_, new_n23439_, new_n23440_, new_n23441_,
    new_n23442_, new_n23443_, new_n23444_, new_n23445_, new_n23446_,
    new_n23447_, new_n23448_, new_n23449_, new_n23450_, new_n23451_,
    new_n23452_, new_n23453_, new_n23454_, new_n23455_, new_n23456_,
    new_n23457_, new_n23458_, new_n23459_, new_n23460_, new_n23461_,
    new_n23462_, new_n23463_, new_n23464_, new_n23465_, new_n23466_,
    new_n23467_, new_n23468_, new_n23469_, new_n23470_, new_n23471_,
    new_n23472_, new_n23473_, new_n23474_, new_n23475_, new_n23476_,
    new_n23477_, new_n23478_, new_n23479_, new_n23480_, new_n23481_,
    new_n23482_, new_n23483_, new_n23484_, new_n23485_, new_n23486_,
    new_n23487_, new_n23488_, new_n23489_, new_n23490_, new_n23491_,
    new_n23492_, new_n23493_, new_n23494_, new_n23495_, new_n23496_,
    new_n23497_, new_n23498_, new_n23499_, new_n23500_, new_n23501_,
    new_n23502_, new_n23503_, new_n23504_, new_n23505_, new_n23506_,
    new_n23507_, new_n23508_, new_n23509_, new_n23510_, new_n23511_,
    new_n23512_, new_n23513_, new_n23514_, new_n23515_, new_n23516_,
    new_n23517_, new_n23518_, new_n23519_, new_n23520_, new_n23521_,
    new_n23522_, new_n23523_, new_n23524_, new_n23525_, new_n23526_,
    new_n23527_, new_n23528_, new_n23529_, new_n23530_, new_n23531_,
    new_n23532_, new_n23533_, new_n23534_, new_n23535_, new_n23536_,
    new_n23537_, new_n23538_, new_n23539_, new_n23540_, new_n23541_,
    new_n23542_, new_n23543_, new_n23544_, new_n23545_, new_n23546_,
    new_n23547_, new_n23548_, new_n23549_, new_n23550_, new_n23551_,
    new_n23552_, new_n23553_, new_n23554_, new_n23555_, new_n23556_,
    new_n23557_, new_n23558_, new_n23559_, new_n23560_, new_n23561_,
    new_n23562_, new_n23563_, new_n23564_, new_n23565_, new_n23566_,
    new_n23567_, new_n23568_, new_n23569_, new_n23570_, new_n23571_,
    new_n23572_, new_n23573_, new_n23574_, new_n23575_, new_n23576_,
    new_n23577_, new_n23578_, new_n23579_, new_n23580_, new_n23581_,
    new_n23582_, new_n23583_, new_n23584_, new_n23585_, new_n23586_,
    new_n23587_, new_n23588_, new_n23589_, new_n23590_, new_n23591_,
    new_n23592_, new_n23593_, new_n23594_, new_n23595_, new_n23596_,
    new_n23597_, new_n23598_, new_n23599_, new_n23600_, new_n23601_,
    new_n23602_, new_n23603_, new_n23604_, new_n23605_, new_n23606_,
    new_n23607_, new_n23608_, new_n23609_, new_n23610_, new_n23611_,
    new_n23612_, new_n23613_, new_n23614_, new_n23615_, new_n23616_,
    new_n23617_, new_n23618_, new_n23619_, new_n23620_, new_n23621_,
    new_n23622_, new_n23623_, new_n23624_, new_n23625_, new_n23626_,
    new_n23627_, new_n23628_, new_n23629_, new_n23630_, new_n23631_,
    new_n23632_, new_n23633_, new_n23634_, new_n23635_, new_n23636_,
    new_n23637_, new_n23638_, new_n23639_, new_n23640_, new_n23641_,
    new_n23642_, new_n23643_, new_n23644_, new_n23645_, new_n23646_,
    new_n23647_, new_n23648_, new_n23649_, new_n23650_, new_n23651_,
    new_n23652_, new_n23653_, new_n23654_, new_n23655_, new_n23656_,
    new_n23657_, new_n23658_, new_n23659_, new_n23660_, new_n23661_,
    new_n23662_, new_n23663_, new_n23664_, new_n23665_, new_n23666_,
    new_n23667_, new_n23668_, new_n23669_, new_n23670_, new_n23671_,
    new_n23672_, new_n23673_, new_n23674_, new_n23675_, new_n23676_,
    new_n23677_, new_n23678_, new_n23679_, new_n23680_, new_n23681_,
    new_n23682_, new_n23683_, new_n23684_, new_n23685_, new_n23686_,
    new_n23687_, new_n23688_, new_n23689_, new_n23690_, new_n23691_,
    new_n23692_, new_n23693_, new_n23694_, new_n23695_, new_n23696_,
    new_n23697_, new_n23698_, new_n23699_, new_n23700_, new_n23701_,
    new_n23702_, new_n23703_, new_n23704_, new_n23705_, new_n23706_,
    new_n23707_, new_n23708_, new_n23709_, new_n23710_, new_n23711_,
    new_n23712_, new_n23713_, new_n23714_, new_n23715_, new_n23716_,
    new_n23717_, new_n23718_, new_n23719_, new_n23720_, new_n23721_,
    new_n23722_, new_n23723_, new_n23724_, new_n23725_, new_n23726_,
    new_n23727_, new_n23729_, new_n23730_, new_n23731_, new_n23732_,
    new_n23733_, new_n23734_, new_n23735_, new_n23736_, new_n23737_,
    new_n23738_, new_n23739_, new_n23740_, new_n23741_, new_n23742_,
    new_n23743_, new_n23744_, new_n23745_, new_n23746_, new_n23747_,
    new_n23748_, new_n23749_, new_n23750_, new_n23751_, new_n23752_,
    new_n23753_, new_n23754_, new_n23755_, new_n23756_, new_n23757_,
    new_n23758_, new_n23759_, new_n23760_, new_n23761_, new_n23762_,
    new_n23763_, new_n23764_, new_n23765_, new_n23766_, new_n23767_,
    new_n23768_, new_n23769_, new_n23770_, new_n23771_, new_n23772_,
    new_n23773_, new_n23774_, new_n23775_, new_n23776_, new_n23777_,
    new_n23778_, new_n23779_, new_n23780_, new_n23781_, new_n23782_,
    new_n23783_, new_n23784_, new_n23785_, new_n23786_, new_n23787_,
    new_n23788_, new_n23789_, new_n23790_, new_n23791_, new_n23792_,
    new_n23793_, new_n23794_, new_n23795_, new_n23796_, new_n23797_,
    new_n23798_, new_n23799_, new_n23800_, new_n23801_, new_n23802_,
    new_n23803_, new_n23804_, new_n23805_, new_n23806_, new_n23807_,
    new_n23808_, new_n23809_, new_n23810_, new_n23811_, new_n23812_,
    new_n23813_, new_n23814_, new_n23815_, new_n23816_, new_n23817_,
    new_n23818_, new_n23819_, new_n23820_, new_n23821_, new_n23822_,
    new_n23823_, new_n23824_, new_n23825_, new_n23826_, new_n23827_,
    new_n23828_, new_n23829_, new_n23830_, new_n23831_, new_n23832_,
    new_n23833_, new_n23834_, new_n23835_, new_n23836_, new_n23837_,
    new_n23838_, new_n23839_, new_n23840_, new_n23841_, new_n23842_,
    new_n23843_, new_n23844_, new_n23845_, new_n23846_, new_n23847_,
    new_n23848_, new_n23849_, new_n23850_, new_n23851_, new_n23852_,
    new_n23853_, new_n23854_, new_n23855_, new_n23856_, new_n23857_,
    new_n23858_, new_n23859_, new_n23860_, new_n23861_, new_n23862_,
    new_n23863_, new_n23864_, new_n23865_, new_n23866_, new_n23867_,
    new_n23868_, new_n23869_, new_n23870_, new_n23871_, new_n23872_,
    new_n23873_, new_n23874_, new_n23875_, new_n23876_, new_n23877_,
    new_n23878_, new_n23879_, new_n23880_, new_n23881_, new_n23882_,
    new_n23883_, new_n23884_, new_n23885_, new_n23886_, new_n23887_,
    new_n23888_, new_n23889_, new_n23890_, new_n23891_, new_n23892_,
    new_n23893_, new_n23894_, new_n23895_, new_n23896_, new_n23897_,
    new_n23898_, new_n23899_, new_n23900_, new_n23901_, new_n23902_,
    new_n23903_, new_n23904_, new_n23905_, new_n23906_, new_n23907_,
    new_n23908_, new_n23909_, new_n23910_, new_n23911_, new_n23912_,
    new_n23913_, new_n23914_, new_n23915_, new_n23916_, new_n23917_,
    new_n23918_, new_n23919_, new_n23920_, new_n23921_, new_n23922_,
    new_n23923_, new_n23924_, new_n23925_, new_n23926_, new_n23927_,
    new_n23928_, new_n23929_, new_n23930_, new_n23931_, new_n23932_,
    new_n23933_, new_n23934_, new_n23935_, new_n23936_, new_n23937_,
    new_n23938_, new_n23939_, new_n23940_, new_n23941_, new_n23942_,
    new_n23943_, new_n23944_, new_n23945_, new_n23946_, new_n23947_,
    new_n23948_, new_n23949_, new_n23950_, new_n23951_, new_n23952_,
    new_n23953_, new_n23954_, new_n23955_, new_n23956_, new_n23957_,
    new_n23958_, new_n23959_, new_n23960_, new_n23961_, new_n23962_,
    new_n23963_, new_n23964_, new_n23965_, new_n23966_, new_n23967_,
    new_n23968_, new_n23969_, new_n23970_, new_n23971_, new_n23972_,
    new_n23973_, new_n23974_, new_n23975_, new_n23976_, new_n23977_,
    new_n23978_, new_n23979_, new_n23980_, new_n23981_, new_n23982_,
    new_n23983_, new_n23984_, new_n23985_, new_n23986_, new_n23987_,
    new_n23988_, new_n23989_, new_n23990_, new_n23991_, new_n23992_,
    new_n23993_, new_n23994_, new_n23995_, new_n23996_, new_n23997_,
    new_n23998_, new_n23999_, new_n24000_, new_n24001_, new_n24002_,
    new_n24003_, new_n24004_, new_n24005_, new_n24006_, new_n24007_,
    new_n24008_, new_n24009_, new_n24010_, new_n24011_, new_n24012_,
    new_n24013_, new_n24014_, new_n24015_, new_n24016_, new_n24017_,
    new_n24018_, new_n24019_, new_n24020_, new_n24021_, new_n24022_,
    new_n24023_, new_n24024_, new_n24025_, new_n24026_, new_n24027_,
    new_n24028_, new_n24029_, new_n24030_, new_n24031_, new_n24032_,
    new_n24033_, new_n24034_, new_n24035_, new_n24036_, new_n24037_,
    new_n24038_, new_n24039_, new_n24040_, new_n24041_, new_n24042_,
    new_n24043_, new_n24044_, new_n24045_, new_n24046_, new_n24047_,
    new_n24048_, new_n24049_, new_n24050_, new_n24051_, new_n24052_,
    new_n24053_, new_n24054_, new_n24055_, new_n24056_, new_n24057_,
    new_n24058_, new_n24059_, new_n24060_, new_n24061_, new_n24062_,
    new_n24063_, new_n24064_, new_n24065_, new_n24066_, new_n24067_,
    new_n24068_, new_n24069_, new_n24070_, new_n24071_, new_n24072_,
    new_n24073_, new_n24074_, new_n24075_, new_n24076_, new_n24077_,
    new_n24078_, new_n24079_, new_n24080_, new_n24081_, new_n24082_,
    new_n24083_, new_n24084_, new_n24085_, new_n24086_, new_n24087_,
    new_n24088_, new_n24089_, new_n24090_, new_n24091_, new_n24092_,
    new_n24093_, new_n24094_, new_n24095_, new_n24096_, new_n24097_,
    new_n24098_, new_n24099_, new_n24100_, new_n24101_, new_n24102_,
    new_n24103_, new_n24104_, new_n24105_, new_n24106_, new_n24107_,
    new_n24108_, new_n24109_, new_n24110_, new_n24111_, new_n24112_,
    new_n24113_, new_n24114_, new_n24115_, new_n24116_, new_n24117_,
    new_n24118_, new_n24119_, new_n24120_, new_n24121_, new_n24122_,
    new_n24123_, new_n24124_, new_n24125_, new_n24126_, new_n24127_,
    new_n24128_, new_n24129_, new_n24130_, new_n24131_, new_n24132_,
    new_n24133_, new_n24134_, new_n24135_, new_n24136_, new_n24137_,
    new_n24138_, new_n24139_, new_n24140_, new_n24141_, new_n24142_,
    new_n24143_, new_n24144_, new_n24145_, new_n24146_, new_n24147_,
    new_n24148_, new_n24149_, new_n24150_, new_n24151_, new_n24152_,
    new_n24153_, new_n24154_, new_n24155_, new_n24156_, new_n24157_,
    new_n24158_, new_n24159_, new_n24160_, new_n24161_, new_n24162_,
    new_n24163_, new_n24164_, new_n24165_, new_n24166_, new_n24167_,
    new_n24168_, new_n24169_, new_n24170_, new_n24171_, new_n24172_,
    new_n24173_, new_n24174_, new_n24175_, new_n24176_, new_n24177_,
    new_n24178_, new_n24179_, new_n24180_, new_n24181_, new_n24182_,
    new_n24183_, new_n24184_, new_n24185_, new_n24186_, new_n24187_,
    new_n24188_, new_n24189_, new_n24190_, new_n24191_, new_n24192_,
    new_n24193_, new_n24194_, new_n24195_, new_n24196_, new_n24197_,
    new_n24198_, new_n24199_, new_n24200_, new_n24201_, new_n24202_,
    new_n24203_, new_n24204_, new_n24205_, new_n24206_, new_n24207_,
    new_n24208_, new_n24209_, new_n24210_, new_n24211_, new_n24212_,
    new_n24213_, new_n24214_, new_n24215_, new_n24216_, new_n24217_,
    new_n24218_, new_n24219_, new_n24220_, new_n24221_, new_n24222_,
    new_n24223_, new_n24224_, new_n24225_, new_n24226_, new_n24227_,
    new_n24228_, new_n24229_, new_n24230_, new_n24231_, new_n24232_,
    new_n24233_, new_n24234_, new_n24235_, new_n24236_, new_n24237_,
    new_n24238_, new_n24239_, new_n24240_, new_n24241_, new_n24242_,
    new_n24243_, new_n24244_, new_n24245_, new_n24246_, new_n24247_,
    new_n24248_, new_n24249_, new_n24250_, new_n24251_, new_n24252_,
    new_n24253_, new_n24254_, new_n24255_, new_n24256_, new_n24257_,
    new_n24258_, new_n24259_, new_n24260_, new_n24261_, new_n24262_,
    new_n24263_, new_n24264_, new_n24265_, new_n24266_, new_n24267_,
    new_n24268_, new_n24269_, new_n24270_, new_n24271_, new_n24272_,
    new_n24273_, new_n24274_, new_n24275_, new_n24276_, new_n24277_,
    new_n24278_, new_n24279_, new_n24280_, new_n24281_, new_n24282_,
    new_n24283_, new_n24284_, new_n24285_, new_n24286_, new_n24287_,
    new_n24288_, new_n24289_, new_n24290_, new_n24291_, new_n24292_,
    new_n24293_, new_n24294_, new_n24295_, new_n24296_, new_n24297_,
    new_n24298_, new_n24299_, new_n24300_, new_n24301_, new_n24302_,
    new_n24303_, new_n24304_, new_n24305_, new_n24306_, new_n24307_,
    new_n24308_, new_n24309_, new_n24310_, new_n24311_, new_n24312_,
    new_n24313_, new_n24314_, new_n24315_, new_n24316_, new_n24317_,
    new_n24318_, new_n24319_, new_n24320_, new_n24321_, new_n24322_,
    new_n24323_, new_n24324_, new_n24325_, new_n24326_, new_n24327_,
    new_n24328_, new_n24329_, new_n24330_, new_n24331_, new_n24332_,
    new_n24333_, new_n24334_, new_n24335_, new_n24336_, new_n24337_,
    new_n24338_, new_n24339_, new_n24340_, new_n24341_, new_n24342_,
    new_n24343_, new_n24344_, new_n24345_, new_n24346_, new_n24347_,
    new_n24348_, new_n24349_, new_n24350_, new_n24351_, new_n24352_,
    new_n24353_, new_n24354_, new_n24355_, new_n24356_, new_n24357_,
    new_n24358_, new_n24359_, new_n24360_, new_n24361_, new_n24362_,
    new_n24363_, new_n24364_, new_n24365_, new_n24366_, new_n24367_,
    new_n24368_, new_n24369_, new_n24370_, new_n24371_, new_n24372_,
    new_n24373_, new_n24374_, new_n24375_, new_n24376_, new_n24377_,
    new_n24378_, new_n24379_, new_n24380_, new_n24381_, new_n24382_,
    new_n24383_, new_n24384_, new_n24385_, new_n24386_, new_n24387_,
    new_n24388_, new_n24389_, new_n24390_, new_n24391_, new_n24392_,
    new_n24393_, new_n24394_, new_n24395_, new_n24396_, new_n24397_,
    new_n24398_, new_n24399_, new_n24400_, new_n24401_, new_n24402_,
    new_n24403_, new_n24404_, new_n24405_, new_n24406_, new_n24407_,
    new_n24408_, new_n24409_, new_n24410_, new_n24411_, new_n24412_,
    new_n24413_, new_n24414_, new_n24415_, new_n24416_, new_n24417_,
    new_n24418_, new_n24419_, new_n24420_, new_n24421_, new_n24422_,
    new_n24423_, new_n24424_, new_n24425_, new_n24426_, new_n24427_,
    new_n24428_, new_n24429_, new_n24430_, new_n24431_, new_n24432_,
    new_n24433_, new_n24434_, new_n24435_, new_n24436_, new_n24437_,
    new_n24438_, new_n24439_, new_n24440_, new_n24441_, new_n24442_,
    new_n24443_, new_n24444_, new_n24445_, new_n24446_, new_n24447_,
    new_n24448_, new_n24449_, new_n24450_, new_n24451_, new_n24452_,
    new_n24453_, new_n24454_, new_n24455_, new_n24456_, new_n24457_,
    new_n24458_, new_n24459_, new_n24460_, new_n24461_, new_n24462_,
    new_n24463_, new_n24464_, new_n24465_, new_n24466_, new_n24467_,
    new_n24468_, new_n24469_, new_n24470_, new_n24471_, new_n24472_,
    new_n24473_, new_n24474_, new_n24475_, new_n24476_, new_n24477_,
    new_n24478_, new_n24479_, new_n24480_, new_n24481_, new_n24483_,
    new_n24484_, new_n24485_, new_n24486_, new_n24487_, new_n24488_,
    new_n24489_, new_n24490_, new_n24491_, new_n24492_, new_n24493_,
    new_n24494_, new_n24495_, new_n24496_, new_n24497_, new_n24498_,
    new_n24499_, new_n24500_, new_n24501_, new_n24502_, new_n24503_,
    new_n24504_, new_n24505_, new_n24506_, new_n24507_, new_n24508_,
    new_n24509_, new_n24510_, new_n24511_, new_n24512_, new_n24513_,
    new_n24514_, new_n24515_, new_n24516_, new_n24517_, new_n24518_,
    new_n24519_, new_n24520_, new_n24521_, new_n24522_, new_n24523_,
    new_n24524_, new_n24525_, new_n24526_, new_n24527_, new_n24528_,
    new_n24529_, new_n24530_, new_n24531_, new_n24532_, new_n24533_,
    new_n24534_, new_n24535_, new_n24536_, new_n24537_, new_n24538_,
    new_n24539_, new_n24540_, new_n24541_, new_n24542_, new_n24543_,
    new_n24544_, new_n24545_, new_n24546_, new_n24547_, new_n24548_,
    new_n24549_, new_n24550_, new_n24551_, new_n24552_, new_n24553_,
    new_n24554_, new_n24555_, new_n24556_, new_n24557_, new_n24558_,
    new_n24559_, new_n24560_, new_n24561_, new_n24562_, new_n24563_,
    new_n24564_, new_n24565_, new_n24566_, new_n24567_, new_n24568_,
    new_n24569_, new_n24570_, new_n24571_, new_n24572_, new_n24573_,
    new_n24574_, new_n24575_, new_n24576_, new_n24577_, new_n24578_,
    new_n24579_, new_n24580_, new_n24581_, new_n24582_, new_n24583_,
    new_n24584_, new_n24585_, new_n24586_, new_n24587_, new_n24588_,
    new_n24589_, new_n24590_, new_n24591_, new_n24592_, new_n24593_,
    new_n24594_, new_n24595_, new_n24596_, new_n24597_, new_n24598_,
    new_n24599_, new_n24600_, new_n24601_, new_n24602_, new_n24603_,
    new_n24604_, new_n24605_, new_n24606_, new_n24607_, new_n24608_,
    new_n24609_, new_n24610_, new_n24611_, new_n24612_, new_n24613_,
    new_n24614_, new_n24615_, new_n24616_, new_n24617_, new_n24618_,
    new_n24619_, new_n24620_, new_n24621_, new_n24622_, new_n24623_,
    new_n24624_, new_n24625_, new_n24626_, new_n24627_, new_n24628_,
    new_n24629_, new_n24630_, new_n24631_, new_n24632_, new_n24633_,
    new_n24634_, new_n24635_, new_n24636_, new_n24637_, new_n24638_,
    new_n24639_, new_n24640_, new_n24641_, new_n24642_, new_n24643_,
    new_n24644_, new_n24645_, new_n24646_, new_n24647_, new_n24648_,
    new_n24649_, new_n24650_, new_n24651_, new_n24652_, new_n24653_,
    new_n24654_, new_n24655_, new_n24656_, new_n24657_, new_n24658_,
    new_n24659_, new_n24660_, new_n24661_, new_n24662_, new_n24663_,
    new_n24664_, new_n24665_, new_n24666_, new_n24667_, new_n24668_,
    new_n24669_, new_n24670_, new_n24671_, new_n24672_, new_n24673_,
    new_n24674_, new_n24675_, new_n24676_, new_n24677_, new_n24678_,
    new_n24679_, new_n24680_, new_n24681_, new_n24682_, new_n24683_,
    new_n24684_, new_n24685_, new_n24686_, new_n24687_, new_n24688_,
    new_n24689_, new_n24690_, new_n24691_, new_n24692_, new_n24693_,
    new_n24694_, new_n24695_, new_n24696_, new_n24697_, new_n24698_,
    new_n24699_, new_n24700_, new_n24701_, new_n24702_, new_n24703_,
    new_n24704_, new_n24705_, new_n24706_, new_n24707_, new_n24708_,
    new_n24709_, new_n24710_, new_n24711_, new_n24712_, new_n24713_,
    new_n24714_, new_n24715_, new_n24716_, new_n24717_, new_n24718_,
    new_n24719_, new_n24720_, new_n24721_, new_n24722_, new_n24723_,
    new_n24724_, new_n24725_, new_n24726_, new_n24727_, new_n24728_,
    new_n24729_, new_n24730_, new_n24731_, new_n24732_, new_n24733_,
    new_n24734_, new_n24735_, new_n24736_, new_n24737_, new_n24738_,
    new_n24739_, new_n24740_, new_n24741_, new_n24742_, new_n24743_,
    new_n24744_, new_n24745_, new_n24746_, new_n24747_, new_n24748_,
    new_n24749_, new_n24750_, new_n24751_, new_n24752_, new_n24753_,
    new_n24754_, new_n24755_, new_n24756_, new_n24757_, new_n24758_,
    new_n24759_, new_n24760_, new_n24761_, new_n24762_, new_n24763_,
    new_n24764_, new_n24765_, new_n24766_, new_n24767_, new_n24768_,
    new_n24769_, new_n24770_, new_n24771_, new_n24772_, new_n24773_,
    new_n24774_, new_n24775_, new_n24776_, new_n24777_, new_n24778_,
    new_n24779_, new_n24780_, new_n24781_, new_n24782_, new_n24783_,
    new_n24784_, new_n24785_, new_n24786_, new_n24787_, new_n24788_,
    new_n24789_, new_n24790_, new_n24791_, new_n24792_, new_n24793_,
    new_n24794_, new_n24795_, new_n24796_, new_n24797_, new_n24798_,
    new_n24799_, new_n24800_, new_n24801_, new_n24802_, new_n24803_,
    new_n24804_, new_n24805_, new_n24806_, new_n24807_, new_n24808_,
    new_n24809_, new_n24810_, new_n24811_, new_n24812_, new_n24813_,
    new_n24814_, new_n24815_, new_n24816_, new_n24817_, new_n24818_,
    new_n24819_, new_n24820_, new_n24821_, new_n24822_, new_n24823_,
    new_n24824_, new_n24825_, new_n24826_, new_n24827_, new_n24828_,
    new_n24829_, new_n24830_, new_n24831_, new_n24832_, new_n24833_,
    new_n24834_, new_n24835_, new_n24836_, new_n24837_, new_n24838_,
    new_n24839_, new_n24840_, new_n24841_, new_n24842_, new_n24843_,
    new_n24844_, new_n24845_, new_n24846_, new_n24847_, new_n24848_,
    new_n24849_, new_n24850_, new_n24851_, new_n24852_, new_n24853_,
    new_n24854_, new_n24855_, new_n24856_, new_n24857_, new_n24858_,
    new_n24859_, new_n24860_, new_n24861_, new_n24862_, new_n24863_,
    new_n24864_, new_n24865_, new_n24866_, new_n24867_, new_n24868_,
    new_n24869_, new_n24870_, new_n24871_, new_n24872_, new_n24873_,
    new_n24874_, new_n24875_, new_n24876_, new_n24877_, new_n24878_,
    new_n24879_, new_n24880_, new_n24881_, new_n24882_, new_n24883_,
    new_n24884_, new_n24885_, new_n24886_, new_n24887_, new_n24888_,
    new_n24889_, new_n24890_, new_n24891_, new_n24892_, new_n24893_,
    new_n24894_, new_n24895_, new_n24896_, new_n24897_, new_n24898_,
    new_n24899_, new_n24900_, new_n24901_, new_n24902_, new_n24903_,
    new_n24904_, new_n24905_, new_n24906_, new_n24907_, new_n24908_,
    new_n24909_, new_n24910_, new_n24911_, new_n24912_, new_n24913_,
    new_n24914_, new_n24915_, new_n24916_, new_n24917_, new_n24918_,
    new_n24919_, new_n24920_, new_n24921_, new_n24922_, new_n24923_,
    new_n24924_, new_n24925_, new_n24926_, new_n24927_, new_n24928_,
    new_n24929_, new_n24930_, new_n24931_, new_n24932_, new_n24933_,
    new_n24934_, new_n24935_, new_n24936_, new_n24937_, new_n24938_,
    new_n24939_, new_n24940_, new_n24941_, new_n24942_, new_n24943_,
    new_n24944_, new_n24945_, new_n24946_, new_n24947_, new_n24948_,
    new_n24949_, new_n24950_, new_n24951_, new_n24952_, new_n24953_,
    new_n24954_, new_n24955_, new_n24956_, new_n24957_, new_n24958_,
    new_n24959_, new_n24960_, new_n24961_, new_n24962_, new_n24963_,
    new_n24964_, new_n24965_, new_n24966_, new_n24967_, new_n24968_,
    new_n24969_, new_n24970_, new_n24971_, new_n24972_, new_n24973_,
    new_n24974_, new_n24975_, new_n24976_, new_n24977_, new_n24978_,
    new_n24979_, new_n24980_, new_n24981_, new_n24982_, new_n24983_,
    new_n24984_, new_n24985_, new_n24986_, new_n24987_, new_n24988_,
    new_n24989_, new_n24990_, new_n24991_, new_n24992_, new_n24993_,
    new_n24994_, new_n24995_, new_n24996_, new_n24997_, new_n24998_,
    new_n24999_, new_n25000_, new_n25001_, new_n25002_, new_n25003_,
    new_n25004_, new_n25005_, new_n25006_, new_n25007_, new_n25008_,
    new_n25009_, new_n25010_, new_n25011_, new_n25012_, new_n25013_,
    new_n25014_, new_n25015_, new_n25016_, new_n25017_, new_n25018_,
    new_n25019_, new_n25020_, new_n25021_, new_n25022_, new_n25023_,
    new_n25024_, new_n25025_, new_n25026_, new_n25027_, new_n25028_,
    new_n25029_, new_n25030_, new_n25031_, new_n25032_, new_n25033_,
    new_n25034_, new_n25035_, new_n25036_, new_n25037_, new_n25038_,
    new_n25039_, new_n25040_, new_n25041_, new_n25042_, new_n25043_,
    new_n25044_;
  NOR2_X1    g00000(.A1(\a[126] ), .A2(\a[127] ), .ZN(new_n193_));
  NAND2_X1   g00001(.A1(\a[126] ), .A2(\a[127] ), .ZN(new_n194_));
  INV_X1     g00002(.I(\a[126] ), .ZN(new_n195_));
  OAI21_X1   g00003(.A1(\a[124] ), .A2(\a[125] ), .B(new_n195_), .ZN(new_n196_));
  NAND2_X1   g00004(.A1(new_n196_), .A2(new_n194_), .ZN(\asqrt[62] ));
  INV_X1     g00005(.I(new_n193_), .ZN(\asqrt[63] ));
  INV_X1     g00006(.I(\a[124] ), .ZN(new_n199_));
  INV_X1     g00007(.I(new_n194_), .ZN(new_n200_));
  INV_X1     g00008(.I(\a[125] ), .ZN(new_n201_));
  AOI21_X1   g00009(.A1(new_n199_), .A2(new_n201_), .B(\a[126] ), .ZN(new_n202_));
  OAI21_X1   g00010(.A1(new_n202_), .A2(new_n200_), .B(new_n199_), .ZN(new_n203_));
  INV_X1     g00011(.I(\a[127] ), .ZN(new_n204_));
  NOR4_X1    g00012(.A1(new_n195_), .A2(new_n204_), .A3(\a[124] ), .A4(\a[125] ), .ZN(new_n205_));
  AOI21_X1   g00013(.A1(new_n203_), .A2(\a[125] ), .B(new_n205_), .ZN(new_n206_));
  NOR2_X1    g00014(.A1(new_n202_), .A2(new_n200_), .ZN(new_n207_));
  NOR2_X1    g00015(.A1(\a[122] ), .A2(\a[123] ), .ZN(new_n208_));
  NAND2_X1   g00016(.A1(new_n208_), .A2(new_n199_), .ZN(new_n209_));
  OAI21_X1   g00017(.A1(new_n207_), .A2(new_n199_), .B(new_n209_), .ZN(new_n210_));
  AOI21_X1   g00018(.A1(new_n206_), .A2(new_n210_), .B(\asqrt[63] ), .ZN(new_n211_));
  NOR3_X1    g00019(.A1(new_n195_), .A2(\a[124] ), .A3(\a[125] ), .ZN(new_n212_));
  NOR2_X1    g00020(.A1(\a[124] ), .A2(\a[125] ), .ZN(new_n213_));
  OAI21_X1   g00021(.A1(new_n213_), .A2(\a[126] ), .B(\a[127] ), .ZN(new_n214_));
  NOR2_X1    g00022(.A1(new_n214_), .A2(new_n212_), .ZN(new_n215_));
  INV_X1     g00023(.I(new_n215_), .ZN(new_n216_));
  OAI21_X1   g00024(.A1(new_n206_), .A2(new_n210_), .B(new_n216_), .ZN(new_n217_));
  NOR2_X1    g00025(.A1(new_n211_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1   g00026(.A1(new_n211_), .A2(new_n217_), .B(\a[122] ), .ZN(new_n219_));
  INV_X1     g00027(.I(\a[122] ), .ZN(new_n220_));
  NOR2_X1    g00028(.A1(\a[120] ), .A2(\a[121] ), .ZN(new_n221_));
  NAND2_X1   g00029(.A1(new_n221_), .A2(new_n220_), .ZN(new_n222_));
  NAND3_X1   g00030(.A1(new_n196_), .A2(new_n222_), .A3(new_n194_), .ZN(new_n223_));
  INV_X1     g00031(.I(new_n223_), .ZN(new_n224_));
  NAND2_X1   g00032(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  AOI21_X1   g00033(.A1(new_n196_), .A2(new_n194_), .B(\a[124] ), .ZN(new_n226_));
  INV_X1     g00034(.I(new_n205_), .ZN(new_n227_));
  OAI21_X1   g00035(.A1(new_n226_), .A2(new_n201_), .B(new_n227_), .ZN(new_n228_));
  INV_X1     g00036(.I(new_n209_), .ZN(new_n229_));
  AOI21_X1   g00037(.A1(\asqrt[62] ), .A2(\a[124] ), .B(new_n229_), .ZN(new_n230_));
  OAI21_X1   g00038(.A1(new_n228_), .A2(new_n230_), .B(new_n193_), .ZN(new_n231_));
  NAND2_X1   g00039(.A1(new_n228_), .A2(new_n230_), .ZN(new_n232_));
  NAND3_X1   g00040(.A1(new_n231_), .A2(new_n232_), .A3(new_n216_), .ZN(\asqrt[61] ));
  OAI21_X1   g00041(.A1(new_n211_), .A2(new_n217_), .B(new_n220_), .ZN(new_n234_));
  AOI22_X1   g00042(.A1(new_n234_), .A2(\a[123] ), .B1(\asqrt[61] ), .B2(new_n208_), .ZN(new_n235_));
  AOI21_X1   g00043(.A1(new_n219_), .A2(new_n222_), .B(new_n207_), .ZN(new_n236_));
  AOI21_X1   g00044(.A1(new_n235_), .A2(new_n225_), .B(new_n236_), .ZN(new_n237_));
  OAI21_X1   g00045(.A1(new_n211_), .A2(new_n217_), .B(new_n208_), .ZN(new_n238_));
  NOR2_X1    g00046(.A1(new_n215_), .A2(new_n207_), .ZN(new_n239_));
  NAND3_X1   g00047(.A1(new_n231_), .A2(new_n232_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1   g00048(.A1(new_n238_), .A2(new_n240_), .B(new_n199_), .ZN(new_n241_));
  INV_X1     g00049(.I(new_n208_), .ZN(new_n242_));
  AOI21_X1   g00050(.A1(new_n228_), .A2(new_n230_), .B(new_n215_), .ZN(new_n243_));
  AOI21_X1   g00051(.A1(new_n243_), .A2(new_n231_), .B(new_n242_), .ZN(new_n244_));
  OAI21_X1   g00052(.A1(new_n206_), .A2(new_n210_), .B(new_n239_), .ZN(new_n245_));
  OAI21_X1   g00053(.A1(new_n245_), .A2(new_n211_), .B(new_n199_), .ZN(new_n246_));
  NOR2_X1    g00054(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1    g00055(.A1(new_n228_), .A2(new_n230_), .ZN(new_n248_));
  INV_X1     g00056(.I(new_n232_), .ZN(new_n249_));
  AOI21_X1   g00057(.A1(\asqrt[61] ), .A2(new_n248_), .B(new_n249_), .ZN(new_n250_));
  OAI21_X1   g00058(.A1(new_n241_), .A2(new_n247_), .B(new_n250_), .ZN(new_n251_));
  OAI21_X1   g00059(.A1(new_n237_), .A2(new_n251_), .B(new_n193_), .ZN(new_n252_));
  NOR2_X1    g00060(.A1(new_n241_), .A2(new_n247_), .ZN(new_n253_));
  NAND2_X1   g00061(.A1(new_n237_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1   g00062(.A1(new_n218_), .A2(new_n228_), .B(new_n230_), .ZN(new_n255_));
  NOR2_X1    g00063(.A1(new_n248_), .A2(new_n193_), .ZN(new_n256_));
  NOR4_X1    g00064(.A1(new_n206_), .A2(new_n230_), .A3(new_n193_), .A4(new_n215_), .ZN(new_n257_));
  AOI21_X1   g00065(.A1(new_n255_), .A2(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND3_X1   g00066(.A1(new_n252_), .A2(new_n254_), .A3(new_n258_), .ZN(\asqrt[60] ));
  NOR2_X1    g00067(.A1(\a[118] ), .A2(\a[119] ), .ZN(new_n260_));
  INV_X1     g00068(.I(new_n260_), .ZN(new_n261_));
  NOR2_X1    g00069(.A1(new_n261_), .A2(\a[120] ), .ZN(new_n262_));
  INV_X1     g00070(.I(\a[120] ), .ZN(new_n263_));
  AOI21_X1   g00071(.A1(\asqrt[61] ), .A2(new_n206_), .B(new_n210_), .ZN(new_n264_));
  INV_X1     g00072(.I(new_n256_), .ZN(new_n265_));
  INV_X1     g00073(.I(new_n257_), .ZN(new_n266_));
  OAI21_X1   g00074(.A1(new_n264_), .A2(new_n265_), .B(new_n266_), .ZN(new_n267_));
  AOI21_X1   g00075(.A1(new_n237_), .A2(new_n253_), .B(new_n267_), .ZN(new_n268_));
  AOI21_X1   g00076(.A1(new_n268_), .A2(new_n252_), .B(new_n263_), .ZN(new_n269_));
  OAI21_X1   g00077(.A1(new_n269_), .A2(new_n262_), .B(\asqrt[61] ), .ZN(new_n270_));
  AOI21_X1   g00078(.A1(new_n243_), .A2(new_n231_), .B(new_n220_), .ZN(new_n271_));
  NOR2_X1    g00079(.A1(new_n271_), .A2(new_n223_), .ZN(new_n272_));
  INV_X1     g00080(.I(\a[123] ), .ZN(new_n273_));
  AOI21_X1   g00081(.A1(new_n243_), .A2(new_n231_), .B(\a[122] ), .ZN(new_n274_));
  OAI21_X1   g00082(.A1(new_n273_), .A2(new_n274_), .B(new_n238_), .ZN(new_n275_));
  INV_X1     g00083(.I(new_n222_), .ZN(new_n276_));
  OAI21_X1   g00084(.A1(new_n271_), .A2(new_n276_), .B(\asqrt[62] ), .ZN(new_n277_));
  OAI21_X1   g00085(.A1(new_n275_), .A2(new_n272_), .B(new_n277_), .ZN(new_n278_));
  NOR2_X1    g00086(.A1(new_n245_), .A2(new_n211_), .ZN(new_n279_));
  OAI21_X1   g00087(.A1(new_n244_), .A2(new_n279_), .B(\a[124] ), .ZN(new_n280_));
  NAND3_X1   g00088(.A1(new_n238_), .A2(new_n240_), .A3(new_n199_), .ZN(new_n281_));
  INV_X1     g00089(.I(new_n248_), .ZN(new_n282_));
  OAI21_X1   g00090(.A1(new_n218_), .A2(new_n282_), .B(new_n232_), .ZN(new_n283_));
  AOI21_X1   g00091(.A1(new_n280_), .A2(new_n281_), .B(new_n283_), .ZN(new_n284_));
  AOI21_X1   g00092(.A1(new_n278_), .A2(new_n284_), .B(\asqrt[63] ), .ZN(new_n285_));
  NAND2_X1   g00093(.A1(new_n280_), .A2(new_n281_), .ZN(new_n286_));
  OAI21_X1   g00094(.A1(new_n278_), .A2(new_n286_), .B(new_n258_), .ZN(new_n287_));
  OAI21_X1   g00095(.A1(new_n285_), .A2(new_n287_), .B(\a[120] ), .ZN(new_n288_));
  NOR4_X1    g00096(.A1(new_n249_), .A2(new_n211_), .A3(new_n215_), .A4(new_n262_), .ZN(new_n289_));
  NAND2_X1   g00097(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OAI21_X1   g00098(.A1(new_n285_), .A2(new_n287_), .B(new_n221_), .ZN(new_n291_));
  OAI21_X1   g00099(.A1(new_n285_), .A2(new_n287_), .B(new_n263_), .ZN(new_n292_));
  NAND2_X1   g00100(.A1(new_n292_), .A2(\a[121] ), .ZN(new_n293_));
  NAND3_X1   g00101(.A1(new_n290_), .A2(new_n293_), .A3(new_n291_), .ZN(new_n294_));
  AOI21_X1   g00102(.A1(new_n294_), .A2(new_n270_), .B(new_n207_), .ZN(new_n295_));
  NAND2_X1   g00103(.A1(new_n255_), .A2(new_n256_), .ZN(new_n296_));
  NOR2_X1    g00104(.A1(new_n218_), .A2(new_n257_), .ZN(new_n297_));
  NAND4_X1   g00105(.A1(new_n252_), .A2(new_n254_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  NAND2_X1   g00106(.A1(new_n291_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1   g00107(.A1(new_n299_), .A2(\a[122] ), .ZN(new_n300_));
  NAND3_X1   g00108(.A1(new_n291_), .A2(new_n298_), .A3(new_n220_), .ZN(new_n301_));
  INV_X1     g00109(.I(new_n262_), .ZN(new_n302_));
  AOI21_X1   g00110(.A1(new_n288_), .A2(new_n302_), .B(new_n218_), .ZN(new_n303_));
  NOR2_X1    g00111(.A1(new_n303_), .A2(\asqrt[62] ), .ZN(new_n304_));
  AOI22_X1   g00112(.A1(new_n294_), .A2(new_n304_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n305_));
  NOR2_X1    g00113(.A1(new_n285_), .A2(new_n287_), .ZN(new_n306_));
  NOR2_X1    g00114(.A1(new_n236_), .A2(new_n272_), .ZN(new_n307_));
  INV_X1     g00115(.I(new_n307_), .ZN(new_n308_));
  NOR3_X1    g00116(.A1(new_n306_), .A2(new_n235_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1   g00117(.A1(\asqrt[60] ), .A2(new_n307_), .B(new_n275_), .ZN(new_n310_));
  NOR2_X1    g00118(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1   g00119(.A1(\asqrt[60] ), .A2(new_n278_), .A3(new_n286_), .ZN(new_n312_));
  NAND2_X1   g00120(.A1(new_n312_), .A2(new_n254_), .ZN(new_n313_));
  NOR2_X1    g00121(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1   g00122(.A1(new_n305_), .A2(new_n295_), .B(new_n314_), .ZN(new_n315_));
  AOI22_X1   g00123(.A1(new_n292_), .A2(\a[121] ), .B1(\asqrt[60] ), .B2(new_n221_), .ZN(new_n316_));
  AOI21_X1   g00124(.A1(new_n316_), .A2(new_n290_), .B(new_n303_), .ZN(new_n317_));
  OAI21_X1   g00125(.A1(new_n317_), .A2(new_n207_), .B(new_n311_), .ZN(new_n318_));
  AOI21_X1   g00126(.A1(\asqrt[60] ), .A2(new_n237_), .B(new_n253_), .ZN(new_n319_));
  NAND2_X1   g00127(.A1(new_n254_), .A2(\asqrt[63] ), .ZN(new_n320_));
  NOR2_X1    g00128(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1    g00129(.A1(new_n247_), .A2(new_n257_), .ZN(new_n322_));
  NAND4_X1   g00130(.A1(new_n254_), .A2(new_n280_), .A3(new_n296_), .A4(new_n322_), .ZN(new_n323_));
  NOR2_X1    g00131(.A1(new_n323_), .A2(new_n285_), .ZN(new_n324_));
  NOR2_X1    g00132(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1   g00133(.A1(new_n318_), .A2(new_n305_), .B(new_n325_), .ZN(new_n326_));
  AOI21_X1   g00134(.A1(new_n193_), .A2(new_n315_), .B(new_n326_), .ZN(new_n327_));
  NOR2_X1    g00135(.A1(\a[116] ), .A2(\a[117] ), .ZN(new_n328_));
  INV_X1     g00136(.I(new_n328_), .ZN(new_n329_));
  NOR2_X1    g00137(.A1(new_n329_), .A2(\a[118] ), .ZN(new_n330_));
  INV_X1     g00138(.I(\a[118] ), .ZN(new_n331_));
  NAND2_X1   g00139(.A1(new_n315_), .A2(new_n193_), .ZN(new_n332_));
  INV_X1     g00140(.I(new_n289_), .ZN(new_n333_));
  NOR2_X1    g00141(.A1(new_n269_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1     g00142(.I(new_n291_), .ZN(new_n335_));
  INV_X1     g00143(.I(\a[121] ), .ZN(new_n336_));
  AOI21_X1   g00144(.A1(\asqrt[60] ), .A2(new_n263_), .B(new_n336_), .ZN(new_n337_));
  NOR3_X1    g00145(.A1(new_n334_), .A2(new_n337_), .A3(new_n335_), .ZN(new_n338_));
  AOI21_X1   g00146(.A1(new_n291_), .A2(new_n298_), .B(new_n220_), .ZN(new_n339_));
  AND3_X2    g00147(.A1(new_n291_), .A2(new_n298_), .A3(new_n220_), .Z(new_n340_));
  AOI21_X1   g00148(.A1(\asqrt[60] ), .A2(\a[120] ), .B(new_n262_), .ZN(new_n341_));
  OAI21_X1   g00149(.A1(new_n341_), .A2(new_n218_), .B(new_n207_), .ZN(new_n342_));
  OAI22_X1   g00150(.A1(new_n338_), .A2(new_n342_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n343_));
  AOI21_X1   g00151(.A1(new_n268_), .A2(new_n252_), .B(\a[120] ), .ZN(new_n344_));
  OAI21_X1   g00152(.A1(new_n336_), .A2(new_n344_), .B(new_n291_), .ZN(new_n345_));
  OAI21_X1   g00153(.A1(new_n345_), .A2(new_n334_), .B(new_n270_), .ZN(new_n346_));
  NAND3_X1   g00154(.A1(\asqrt[60] ), .A2(new_n275_), .A3(new_n307_), .ZN(new_n347_));
  NOR2_X1    g00155(.A1(new_n306_), .A2(new_n308_), .ZN(new_n348_));
  OAI21_X1   g00156(.A1(new_n275_), .A2(new_n348_), .B(new_n347_), .ZN(new_n349_));
  AOI21_X1   g00157(.A1(new_n346_), .A2(\asqrt[62] ), .B(new_n349_), .ZN(new_n350_));
  INV_X1     g00158(.I(new_n325_), .ZN(new_n351_));
  AOI21_X1   g00159(.A1(new_n350_), .A2(new_n343_), .B(new_n351_), .ZN(new_n352_));
  AOI21_X1   g00160(.A1(new_n332_), .A2(new_n352_), .B(new_n331_), .ZN(new_n353_));
  OAI21_X1   g00161(.A1(new_n353_), .A2(new_n330_), .B(\asqrt[60] ), .ZN(new_n354_));
  OAI21_X1   g00162(.A1(new_n338_), .A2(new_n303_), .B(\asqrt[62] ), .ZN(new_n355_));
  NAND2_X1   g00163(.A1(new_n343_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1   g00164(.A1(new_n356_), .A2(new_n314_), .B(\asqrt[63] ), .ZN(new_n357_));
  OAI21_X1   g00165(.A1(new_n357_), .A2(new_n326_), .B(\a[118] ), .ZN(new_n358_));
  INV_X1     g00166(.I(new_n330_), .ZN(new_n359_));
  AND3_X2    g00167(.A1(new_n296_), .A2(new_n266_), .A3(new_n359_), .Z(new_n360_));
  NAND3_X1   g00168(.A1(new_n252_), .A2(new_n360_), .A3(new_n254_), .ZN(new_n361_));
  INV_X1     g00169(.I(new_n361_), .ZN(new_n362_));
  NAND2_X1   g00170(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1   g00171(.A1(new_n349_), .A2(new_n254_), .A3(new_n312_), .ZN(new_n364_));
  AOI21_X1   g00172(.A1(new_n343_), .A2(new_n355_), .B(new_n364_), .ZN(new_n365_));
  OAI21_X1   g00173(.A1(\asqrt[63] ), .A2(new_n365_), .B(new_n352_), .ZN(\asqrt[59] ));
  NAND2_X1   g00174(.A1(\asqrt[59] ), .A2(new_n260_), .ZN(new_n367_));
  OAI21_X1   g00175(.A1(new_n327_), .A2(\a[118] ), .B(\a[119] ), .ZN(new_n368_));
  NAND3_X1   g00176(.A1(new_n363_), .A2(new_n368_), .A3(new_n367_), .ZN(new_n369_));
  AOI21_X1   g00177(.A1(new_n369_), .A2(new_n354_), .B(new_n218_), .ZN(new_n370_));
  NOR2_X1    g00178(.A1(new_n327_), .A2(new_n261_), .ZN(new_n371_));
  NAND2_X1   g00179(.A1(new_n350_), .A2(new_n343_), .ZN(new_n372_));
  INV_X1     g00180(.I(new_n321_), .ZN(new_n373_));
  NOR2_X1    g00181(.A1(new_n324_), .A2(new_n306_), .ZN(new_n374_));
  NAND3_X1   g00182(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NOR2_X1    g00183(.A1(new_n375_), .A2(new_n357_), .ZN(new_n376_));
  OAI21_X1   g00184(.A1(new_n371_), .A2(new_n376_), .B(\a[120] ), .ZN(new_n377_));
  NAND4_X1   g00185(.A1(new_n332_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n378_));
  NAND3_X1   g00186(.A1(new_n367_), .A2(new_n263_), .A3(new_n378_), .ZN(new_n379_));
  OAI21_X1   g00187(.A1(new_n327_), .A2(new_n331_), .B(new_n359_), .ZN(new_n380_));
  AOI21_X1   g00188(.A1(new_n380_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n381_));
  AOI22_X1   g00189(.A1(new_n369_), .A2(new_n381_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n382_));
  OAI21_X1   g00190(.A1(new_n382_), .A2(new_n370_), .B(\asqrt[62] ), .ZN(new_n383_));
  NOR3_X1    g00191(.A1(new_n316_), .A2(new_n303_), .A3(new_n334_), .ZN(new_n384_));
  NAND3_X1   g00192(.A1(\asqrt[59] ), .A2(new_n270_), .A3(new_n290_), .ZN(new_n385_));
  AOI22_X1   g00193(.A1(new_n385_), .A2(new_n316_), .B1(\asqrt[59] ), .B2(new_n384_), .ZN(new_n386_));
  INV_X1     g00194(.I(new_n386_), .ZN(new_n387_));
  AOI21_X1   g00195(.A1(new_n358_), .A2(new_n359_), .B(new_n306_), .ZN(new_n388_));
  OAI21_X1   g00196(.A1(new_n357_), .A2(new_n326_), .B(new_n331_), .ZN(new_n389_));
  AOI22_X1   g00197(.A1(new_n389_), .A2(\a[119] ), .B1(new_n260_), .B2(\asqrt[59] ), .ZN(new_n390_));
  AOI21_X1   g00198(.A1(new_n390_), .A2(new_n363_), .B(new_n388_), .ZN(new_n391_));
  OAI21_X1   g00199(.A1(new_n391_), .A2(new_n218_), .B(new_n207_), .ZN(new_n392_));
  OAI21_X1   g00200(.A1(new_n392_), .A2(new_n382_), .B(new_n387_), .ZN(new_n393_));
  NAND2_X1   g00201(.A1(new_n393_), .A2(new_n383_), .ZN(new_n394_));
  NOR2_X1    g00202(.A1(new_n340_), .A2(new_n339_), .ZN(new_n395_));
  INV_X1     g00203(.I(new_n395_), .ZN(new_n396_));
  NOR2_X1    g00204(.A1(new_n338_), .A2(new_n342_), .ZN(new_n397_));
  NOR3_X1    g00205(.A1(new_n396_), .A2(new_n295_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1   g00206(.A1(\asqrt[59] ), .A2(new_n398_), .ZN(new_n399_));
  OR3_X2     g00207(.A1(new_n327_), .A2(new_n295_), .A3(new_n397_), .Z(new_n400_));
  NAND2_X1   g00208(.A1(new_n400_), .A2(new_n396_), .ZN(new_n401_));
  NAND2_X1   g00209(.A1(new_n401_), .A2(new_n399_), .ZN(new_n402_));
  INV_X1     g00210(.I(new_n372_), .ZN(new_n403_));
  INV_X1     g00211(.I(new_n356_), .ZN(new_n404_));
  NOR2_X1    g00212(.A1(new_n404_), .A2(new_n311_), .ZN(new_n405_));
  AOI21_X1   g00213(.A1(\asqrt[59] ), .A2(new_n405_), .B(new_n403_), .ZN(new_n406_));
  NAND2_X1   g00214(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1     g00215(.I(new_n407_), .ZN(new_n408_));
  AOI21_X1   g00216(.A1(new_n394_), .A2(new_n408_), .B(\asqrt[63] ), .ZN(new_n409_));
  NOR2_X1    g00217(.A1(new_n353_), .A2(new_n361_), .ZN(new_n410_));
  INV_X1     g00218(.I(\a[119] ), .ZN(new_n411_));
  AOI21_X1   g00219(.A1(\asqrt[59] ), .A2(new_n331_), .B(new_n411_), .ZN(new_n412_));
  NOR3_X1    g00220(.A1(new_n410_), .A2(new_n412_), .A3(new_n371_), .ZN(new_n413_));
  AOI21_X1   g00221(.A1(new_n367_), .A2(new_n378_), .B(new_n263_), .ZN(new_n414_));
  NOR3_X1    g00222(.A1(new_n371_), .A2(\a[120] ), .A3(new_n376_), .ZN(new_n415_));
  AOI21_X1   g00223(.A1(\asqrt[59] ), .A2(\a[118] ), .B(new_n330_), .ZN(new_n416_));
  OAI21_X1   g00224(.A1(new_n416_), .A2(new_n306_), .B(new_n218_), .ZN(new_n417_));
  OAI22_X1   g00225(.A1(new_n413_), .A2(new_n417_), .B1(new_n415_), .B2(new_n414_), .ZN(new_n418_));
  AOI21_X1   g00226(.A1(new_n332_), .A2(new_n352_), .B(\a[118] ), .ZN(new_n419_));
  OAI22_X1   g00227(.A1(new_n419_), .A2(new_n411_), .B1(new_n261_), .B2(new_n327_), .ZN(new_n420_));
  OAI21_X1   g00228(.A1(new_n420_), .A2(new_n410_), .B(new_n354_), .ZN(new_n421_));
  AOI21_X1   g00229(.A1(new_n421_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n422_));
  AOI21_X1   g00230(.A1(new_n422_), .A2(new_n418_), .B(new_n386_), .ZN(new_n423_));
  INV_X1     g00231(.I(new_n402_), .ZN(new_n424_));
  NAND2_X1   g00232(.A1(new_n383_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1   g00233(.A1(\asqrt[59] ), .A2(new_n404_), .B(new_n311_), .ZN(new_n426_));
  NOR2_X1    g00234(.A1(new_n403_), .A2(new_n193_), .ZN(new_n427_));
  INV_X1     g00235(.I(new_n427_), .ZN(new_n428_));
  NOR2_X1    g00236(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1   g00237(.A1(new_n285_), .A2(new_n323_), .B(new_n347_), .ZN(new_n430_));
  NOR4_X1    g00238(.A1(new_n403_), .A2(new_n310_), .A3(new_n321_), .A4(new_n430_), .ZN(new_n431_));
  NAND2_X1   g00239(.A1(new_n431_), .A2(new_n332_), .ZN(new_n432_));
  INV_X1     g00240(.I(new_n432_), .ZN(new_n433_));
  NOR2_X1    g00241(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1   g00242(.A1(new_n425_), .A2(new_n423_), .B(new_n434_), .ZN(new_n435_));
  NOR2_X1    g00243(.A1(new_n409_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1    g00244(.A1(\a[114] ), .A2(\a[115] ), .ZN(new_n437_));
  INV_X1     g00245(.I(new_n437_), .ZN(new_n438_));
  NOR2_X1    g00246(.A1(new_n438_), .A2(\a[116] ), .ZN(new_n439_));
  INV_X1     g00247(.I(new_n439_), .ZN(new_n440_));
  OAI21_X1   g00248(.A1(new_n409_), .A2(new_n435_), .B(\a[116] ), .ZN(new_n441_));
  AOI21_X1   g00249(.A1(new_n441_), .A2(new_n440_), .B(new_n327_), .ZN(new_n442_));
  INV_X1     g00250(.I(\a[116] ), .ZN(new_n443_));
  OAI21_X1   g00251(.A1(new_n413_), .A2(new_n388_), .B(\asqrt[61] ), .ZN(new_n444_));
  AOI21_X1   g00252(.A1(new_n418_), .A2(new_n444_), .B(new_n207_), .ZN(new_n445_));
  NOR2_X1    g00253(.A1(new_n423_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1   g00254(.A1(new_n446_), .A2(new_n407_), .B(new_n193_), .ZN(new_n447_));
  NOR2_X1    g00255(.A1(new_n445_), .A2(new_n402_), .ZN(new_n448_));
  INV_X1     g00256(.I(new_n434_), .ZN(new_n449_));
  AOI21_X1   g00257(.A1(new_n448_), .A2(new_n393_), .B(new_n449_), .ZN(new_n450_));
  AOI21_X1   g00258(.A1(new_n447_), .A2(new_n450_), .B(new_n443_), .ZN(new_n451_));
  NOR2_X1    g00259(.A1(new_n324_), .A2(new_n439_), .ZN(new_n452_));
  NAND4_X1   g00260(.A1(new_n332_), .A2(new_n372_), .A3(new_n373_), .A4(new_n452_), .ZN(new_n453_));
  NOR2_X1    g00261(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1   g00262(.A1(new_n409_), .A2(new_n435_), .B(new_n328_), .ZN(new_n455_));
  INV_X1     g00263(.I(new_n455_), .ZN(new_n456_));
  INV_X1     g00264(.I(\a[117] ), .ZN(new_n457_));
  NAND2_X1   g00265(.A1(new_n447_), .A2(new_n450_), .ZN(\asqrt[58] ));
  AOI21_X1   g00266(.A1(\asqrt[58] ), .A2(new_n443_), .B(new_n457_), .ZN(new_n459_));
  NOR3_X1    g00267(.A1(new_n454_), .A2(new_n459_), .A3(new_n456_), .ZN(new_n460_));
  OAI21_X1   g00268(.A1(new_n460_), .A2(new_n442_), .B(\asqrt[60] ), .ZN(new_n461_));
  NAND2_X1   g00269(.A1(new_n448_), .A2(new_n393_), .ZN(new_n462_));
  INV_X1     g00270(.I(new_n429_), .ZN(new_n463_));
  NOR2_X1    g00271(.A1(new_n433_), .A2(new_n327_), .ZN(new_n464_));
  NAND4_X1   g00272(.A1(new_n447_), .A2(new_n462_), .A3(new_n463_), .A4(new_n464_), .ZN(new_n465_));
  AOI21_X1   g00273(.A1(new_n465_), .A2(new_n455_), .B(new_n331_), .ZN(new_n466_));
  NAND3_X1   g00274(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n467_));
  NOR2_X1    g00275(.A1(new_n467_), .A2(new_n409_), .ZN(new_n468_));
  NOR3_X1    g00276(.A1(new_n456_), .A2(new_n468_), .A3(\a[118] ), .ZN(new_n469_));
  OAI21_X1   g00277(.A1(new_n451_), .A2(new_n439_), .B(\asqrt[59] ), .ZN(new_n470_));
  NAND2_X1   g00278(.A1(new_n470_), .A2(new_n306_), .ZN(new_n471_));
  OAI22_X1   g00279(.A1(new_n460_), .A2(new_n471_), .B1(new_n469_), .B2(new_n466_), .ZN(new_n472_));
  AOI21_X1   g00280(.A1(new_n472_), .A2(new_n461_), .B(new_n218_), .ZN(new_n473_));
  NOR3_X1    g00281(.A1(new_n390_), .A2(new_n388_), .A3(new_n410_), .ZN(new_n474_));
  NAND3_X1   g00282(.A1(\asqrt[58] ), .A2(new_n354_), .A3(new_n363_), .ZN(new_n475_));
  AOI22_X1   g00283(.A1(new_n475_), .A2(new_n390_), .B1(\asqrt[58] ), .B2(new_n474_), .ZN(new_n476_));
  AOI21_X1   g00284(.A1(new_n447_), .A2(new_n450_), .B(\a[116] ), .ZN(new_n477_));
  OAI21_X1   g00285(.A1(new_n457_), .A2(new_n477_), .B(new_n455_), .ZN(new_n478_));
  OAI21_X1   g00286(.A1(new_n478_), .A2(new_n454_), .B(new_n470_), .ZN(new_n479_));
  AOI21_X1   g00287(.A1(new_n479_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n480_));
  AOI21_X1   g00288(.A1(new_n480_), .A2(new_n472_), .B(new_n476_), .ZN(new_n481_));
  OAI21_X1   g00289(.A1(new_n481_), .A2(new_n473_), .B(\asqrt[62] ), .ZN(new_n482_));
  NOR2_X1    g00290(.A1(new_n414_), .A2(new_n415_), .ZN(new_n483_));
  NOR2_X1    g00291(.A1(new_n413_), .A2(new_n417_), .ZN(new_n484_));
  INV_X1     g00292(.I(new_n484_), .ZN(new_n485_));
  NAND4_X1   g00293(.A1(\asqrt[58] ), .A2(new_n444_), .A3(new_n483_), .A4(new_n485_), .ZN(new_n486_));
  NOR3_X1    g00294(.A1(new_n436_), .A2(new_n370_), .A3(new_n484_), .ZN(new_n487_));
  OAI21_X1   g00295(.A1(new_n487_), .A2(new_n483_), .B(new_n486_), .ZN(new_n488_));
  INV_X1     g00296(.I(new_n453_), .ZN(new_n489_));
  NAND2_X1   g00297(.A1(new_n441_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1   g00298(.A1(new_n409_), .A2(new_n435_), .B(new_n443_), .ZN(new_n491_));
  NAND2_X1   g00299(.A1(new_n491_), .A2(\a[117] ), .ZN(new_n492_));
  NAND3_X1   g00300(.A1(new_n490_), .A2(new_n492_), .A3(new_n455_), .ZN(new_n493_));
  AOI21_X1   g00301(.A1(new_n493_), .A2(new_n470_), .B(new_n306_), .ZN(new_n494_));
  OAI21_X1   g00302(.A1(new_n456_), .A2(new_n468_), .B(\a[118] ), .ZN(new_n495_));
  NAND3_X1   g00303(.A1(new_n465_), .A2(new_n455_), .A3(new_n331_), .ZN(new_n496_));
  NAND2_X1   g00304(.A1(new_n441_), .A2(new_n440_), .ZN(new_n497_));
  AOI21_X1   g00305(.A1(new_n497_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n498_));
  AOI22_X1   g00306(.A1(new_n493_), .A2(new_n498_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n499_));
  OAI21_X1   g00307(.A1(new_n499_), .A2(new_n494_), .B(\asqrt[61] ), .ZN(new_n500_));
  NAND2_X1   g00308(.A1(new_n500_), .A2(new_n207_), .ZN(new_n501_));
  OAI21_X1   g00309(.A1(new_n501_), .A2(new_n481_), .B(new_n488_), .ZN(new_n502_));
  NOR2_X1    g00310(.A1(new_n392_), .A2(new_n382_), .ZN(new_n503_));
  NOR3_X1    g00311(.A1(new_n503_), .A2(new_n445_), .A3(new_n387_), .ZN(new_n504_));
  NAND2_X1   g00312(.A1(\asqrt[58] ), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1   g00313(.A1(new_n382_), .A2(new_n392_), .B(new_n383_), .ZN(new_n506_));
  OAI21_X1   g00314(.A1(new_n436_), .A2(new_n506_), .B(new_n387_), .ZN(new_n507_));
  NAND2_X1   g00315(.A1(new_n507_), .A2(new_n505_), .ZN(new_n508_));
  INV_X1     g00316(.I(new_n462_), .ZN(new_n509_));
  NOR2_X1    g00317(.A1(new_n446_), .A2(new_n424_), .ZN(new_n510_));
  AOI21_X1   g00318(.A1(\asqrt[58] ), .A2(new_n510_), .B(new_n509_), .ZN(new_n511_));
  NAND2_X1   g00319(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1   g00320(.A1(new_n502_), .A2(new_n482_), .B(new_n512_), .ZN(new_n513_));
  INV_X1     g00321(.I(new_n476_), .ZN(new_n514_));
  AOI22_X1   g00322(.A1(new_n491_), .A2(\a[117] ), .B1(\asqrt[58] ), .B2(new_n328_), .ZN(new_n515_));
  AOI21_X1   g00323(.A1(new_n515_), .A2(new_n490_), .B(new_n442_), .ZN(new_n516_));
  OAI21_X1   g00324(.A1(new_n516_), .A2(new_n306_), .B(new_n218_), .ZN(new_n517_));
  OAI21_X1   g00325(.A1(new_n517_), .A2(new_n499_), .B(new_n514_), .ZN(new_n518_));
  NAND2_X1   g00326(.A1(new_n518_), .A2(new_n500_), .ZN(new_n519_));
  AOI21_X1   g00327(.A1(new_n519_), .A2(\asqrt[62] ), .B(new_n508_), .ZN(new_n520_));
  OAI21_X1   g00328(.A1(new_n436_), .A2(new_n424_), .B(new_n446_), .ZN(new_n521_));
  NOR2_X1    g00329(.A1(new_n510_), .A2(new_n193_), .ZN(new_n522_));
  NAND2_X1   g00330(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1   g00331(.A1(\asqrt[59] ), .A2(new_n398_), .B(new_n433_), .ZN(new_n524_));
  NAND4_X1   g00332(.A1(new_n462_), .A2(new_n401_), .A3(new_n463_), .A4(new_n524_), .ZN(new_n525_));
  NOR2_X1    g00333(.A1(new_n525_), .A2(new_n409_), .ZN(new_n526_));
  INV_X1     g00334(.I(new_n526_), .ZN(new_n527_));
  NAND2_X1   g00335(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1   g00336(.A1(new_n520_), .A2(new_n502_), .B(new_n528_), .ZN(new_n529_));
  OAI21_X1   g00337(.A1(\asqrt[63] ), .A2(new_n513_), .B(new_n529_), .ZN(\asqrt[57] ));
  INV_X1     g00338(.I(\asqrt[57] ), .ZN(new_n531_));
  NOR2_X1    g00339(.A1(\a[112] ), .A2(\a[113] ), .ZN(new_n532_));
  INV_X1     g00340(.I(new_n532_), .ZN(new_n533_));
  NOR2_X1    g00341(.A1(new_n533_), .A2(\a[114] ), .ZN(new_n534_));
  INV_X1     g00342(.I(\a[114] ), .ZN(new_n535_));
  NAND3_X1   g00343(.A1(new_n518_), .A2(new_n500_), .A3(new_n207_), .ZN(new_n536_));
  AOI22_X1   g00344(.A1(new_n536_), .A2(new_n488_), .B1(new_n519_), .B2(\asqrt[62] ), .ZN(new_n537_));
  OAI21_X1   g00345(.A1(new_n537_), .A2(new_n512_), .B(new_n193_), .ZN(new_n538_));
  AOI21_X1   g00346(.A1(new_n538_), .A2(new_n529_), .B(new_n535_), .ZN(new_n539_));
  OAI21_X1   g00347(.A1(new_n539_), .A2(new_n534_), .B(\asqrt[58] ), .ZN(new_n540_));
  INV_X1     g00348(.I(new_n488_), .ZN(new_n541_));
  NOR3_X1    g00349(.A1(new_n481_), .A2(new_n473_), .A3(\asqrt[62] ), .ZN(new_n542_));
  OAI21_X1   g00350(.A1(new_n541_), .A2(new_n542_), .B(new_n482_), .ZN(new_n543_));
  INV_X1     g00351(.I(new_n512_), .ZN(new_n544_));
  AOI21_X1   g00352(.A1(new_n543_), .A2(new_n544_), .B(\asqrt[63] ), .ZN(new_n545_));
  NOR2_X1    g00353(.A1(new_n542_), .A2(new_n541_), .ZN(new_n546_));
  INV_X1     g00354(.I(new_n508_), .ZN(new_n547_));
  NAND2_X1   g00355(.A1(new_n482_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1     g00356(.I(new_n528_), .ZN(new_n549_));
  OAI21_X1   g00357(.A1(new_n546_), .A2(new_n548_), .B(new_n549_), .ZN(new_n550_));
  OAI21_X1   g00358(.A1(new_n545_), .A2(new_n550_), .B(\a[114] ), .ZN(new_n551_));
  INV_X1     g00359(.I(new_n534_), .ZN(new_n552_));
  NAND2_X1   g00360(.A1(new_n432_), .A2(new_n552_), .ZN(new_n553_));
  NOR4_X1    g00361(.A1(new_n509_), .A2(new_n409_), .A3(new_n429_), .A4(new_n553_), .ZN(new_n554_));
  NAND2_X1   g00362(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1   g00363(.A1(new_n545_), .A2(new_n550_), .B(new_n437_), .ZN(new_n556_));
  OAI21_X1   g00364(.A1(new_n545_), .A2(new_n550_), .B(new_n535_), .ZN(new_n557_));
  NAND2_X1   g00365(.A1(new_n557_), .A2(\a[115] ), .ZN(new_n558_));
  NAND3_X1   g00366(.A1(new_n555_), .A2(new_n558_), .A3(new_n556_), .ZN(new_n559_));
  AOI21_X1   g00367(.A1(new_n559_), .A2(new_n540_), .B(new_n327_), .ZN(new_n560_));
  AOI21_X1   g00368(.A1(new_n538_), .A2(new_n529_), .B(new_n438_), .ZN(new_n561_));
  NOR2_X1    g00369(.A1(new_n546_), .A2(new_n548_), .ZN(new_n562_));
  NOR2_X1    g00370(.A1(new_n526_), .A2(new_n436_), .ZN(new_n563_));
  NAND2_X1   g00371(.A1(new_n523_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1    g00372(.A1(new_n545_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  OAI21_X1   g00373(.A1(new_n565_), .A2(new_n561_), .B(\a[116] ), .ZN(new_n566_));
  INV_X1     g00374(.I(new_n565_), .ZN(new_n567_));
  NAND3_X1   g00375(.A1(new_n567_), .A2(new_n556_), .A3(new_n443_), .ZN(new_n568_));
  NAND2_X1   g00376(.A1(new_n551_), .A2(new_n552_), .ZN(new_n569_));
  AOI21_X1   g00377(.A1(new_n569_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n570_));
  AOI22_X1   g00378(.A1(new_n559_), .A2(new_n570_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n571_));
  OAI21_X1   g00379(.A1(new_n571_), .A2(new_n560_), .B(\asqrt[60] ), .ZN(new_n572_));
  NOR3_X1    g00380(.A1(new_n515_), .A2(new_n442_), .A3(new_n454_), .ZN(new_n573_));
  NAND3_X1   g00381(.A1(\asqrt[57] ), .A2(new_n470_), .A3(new_n490_), .ZN(new_n574_));
  AOI22_X1   g00382(.A1(new_n574_), .A2(new_n515_), .B1(\asqrt[57] ), .B2(new_n573_), .ZN(new_n575_));
  INV_X1     g00383(.I(new_n575_), .ZN(new_n576_));
  AOI21_X1   g00384(.A1(new_n551_), .A2(new_n552_), .B(new_n436_), .ZN(new_n577_));
  AOI21_X1   g00385(.A1(\a[115] ), .A2(new_n557_), .B(new_n561_), .ZN(new_n578_));
  AOI21_X1   g00386(.A1(new_n578_), .A2(new_n555_), .B(new_n577_), .ZN(new_n579_));
  OAI21_X1   g00387(.A1(new_n579_), .A2(new_n327_), .B(new_n306_), .ZN(new_n580_));
  OAI21_X1   g00388(.A1(new_n580_), .A2(new_n571_), .B(new_n576_), .ZN(new_n581_));
  AOI21_X1   g00389(.A1(new_n581_), .A2(new_n572_), .B(new_n218_), .ZN(new_n582_));
  NOR2_X1    g00390(.A1(new_n469_), .A2(new_n466_), .ZN(new_n583_));
  NOR2_X1    g00391(.A1(new_n460_), .A2(new_n471_), .ZN(new_n584_));
  INV_X1     g00392(.I(new_n584_), .ZN(new_n585_));
  NAND4_X1   g00393(.A1(\asqrt[57] ), .A2(new_n461_), .A3(new_n583_), .A4(new_n585_), .ZN(new_n586_));
  NOR3_X1    g00394(.A1(new_n531_), .A2(new_n494_), .A3(new_n584_), .ZN(new_n587_));
  OAI21_X1   g00395(.A1(new_n587_), .A2(new_n583_), .B(new_n586_), .ZN(new_n588_));
  INV_X1     g00396(.I(new_n588_), .ZN(new_n589_));
  INV_X1     g00397(.I(new_n554_), .ZN(new_n590_));
  NOR2_X1    g00398(.A1(new_n539_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1     g00399(.I(\a[115] ), .ZN(new_n592_));
  AOI21_X1   g00400(.A1(\asqrt[57] ), .A2(new_n535_), .B(new_n592_), .ZN(new_n593_));
  NOR3_X1    g00401(.A1(new_n591_), .A2(new_n593_), .A3(new_n561_), .ZN(new_n594_));
  OAI21_X1   g00402(.A1(new_n594_), .A2(new_n577_), .B(\asqrt[59] ), .ZN(new_n595_));
  AOI21_X1   g00403(.A1(new_n567_), .A2(new_n556_), .B(new_n443_), .ZN(new_n596_));
  NOR3_X1    g00404(.A1(new_n565_), .A2(new_n561_), .A3(\a[116] ), .ZN(new_n597_));
  AOI21_X1   g00405(.A1(\asqrt[57] ), .A2(\a[114] ), .B(new_n534_), .ZN(new_n598_));
  OAI21_X1   g00406(.A1(new_n598_), .A2(new_n436_), .B(new_n327_), .ZN(new_n599_));
  OAI22_X1   g00407(.A1(new_n594_), .A2(new_n599_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n600_));
  AOI21_X1   g00408(.A1(new_n600_), .A2(new_n595_), .B(new_n306_), .ZN(new_n601_));
  NOR2_X1    g00409(.A1(new_n601_), .A2(\asqrt[61] ), .ZN(new_n602_));
  AOI21_X1   g00410(.A1(new_n602_), .A2(new_n581_), .B(new_n589_), .ZN(new_n603_));
  OAI21_X1   g00411(.A1(new_n603_), .A2(new_n582_), .B(\asqrt[62] ), .ZN(new_n604_));
  NOR2_X1    g00412(.A1(new_n517_), .A2(new_n499_), .ZN(new_n605_));
  NOR3_X1    g00413(.A1(new_n531_), .A2(new_n473_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1     g00414(.I(new_n606_), .ZN(new_n607_));
  NOR3_X1    g00415(.A1(new_n473_), .A2(new_n605_), .A3(new_n514_), .ZN(new_n608_));
  AOI22_X1   g00416(.A1(new_n607_), .A2(new_n514_), .B1(\asqrt[57] ), .B2(new_n608_), .ZN(new_n609_));
  INV_X1     g00417(.I(new_n609_), .ZN(new_n610_));
  AOI21_X1   g00418(.A1(new_n538_), .A2(new_n529_), .B(\a[114] ), .ZN(new_n611_));
  OAI21_X1   g00419(.A1(new_n592_), .A2(new_n611_), .B(new_n556_), .ZN(new_n612_));
  OAI21_X1   g00420(.A1(new_n612_), .A2(new_n591_), .B(new_n540_), .ZN(new_n613_));
  AOI21_X1   g00421(.A1(new_n613_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n614_));
  AOI21_X1   g00422(.A1(new_n614_), .A2(new_n600_), .B(new_n575_), .ZN(new_n615_));
  OAI21_X1   g00423(.A1(new_n615_), .A2(new_n601_), .B(\asqrt[61] ), .ZN(new_n616_));
  NAND2_X1   g00424(.A1(new_n616_), .A2(new_n207_), .ZN(new_n617_));
  OAI21_X1   g00425(.A1(new_n617_), .A2(new_n603_), .B(new_n610_), .ZN(new_n618_));
  INV_X1     g00426(.I(new_n562_), .ZN(new_n619_));
  NAND4_X1   g00427(.A1(\asqrt[57] ), .A2(new_n482_), .A3(new_n541_), .A4(new_n536_), .ZN(new_n620_));
  NAND2_X1   g00428(.A1(new_n482_), .A2(new_n536_), .ZN(new_n621_));
  OAI21_X1   g00429(.A1(new_n531_), .A2(new_n621_), .B(new_n488_), .ZN(new_n622_));
  NAND2_X1   g00430(.A1(new_n622_), .A2(new_n620_), .ZN(new_n623_));
  NOR2_X1    g00431(.A1(new_n537_), .A2(new_n547_), .ZN(new_n624_));
  NAND2_X1   g00432(.A1(\asqrt[57] ), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1   g00433(.A1(new_n623_), .A2(new_n619_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1   g00434(.A1(new_n618_), .A2(new_n604_), .B(new_n626_), .ZN(new_n627_));
  NOR3_X1    g00435(.A1(new_n615_), .A2(new_n601_), .A3(\asqrt[61] ), .ZN(new_n628_));
  OAI21_X1   g00436(.A1(new_n589_), .A2(new_n628_), .B(new_n616_), .ZN(new_n629_));
  AOI21_X1   g00437(.A1(new_n629_), .A2(\asqrt[62] ), .B(new_n623_), .ZN(new_n630_));
  AOI21_X1   g00438(.A1(\asqrt[57] ), .A2(new_n508_), .B(new_n543_), .ZN(new_n631_));
  NOR2_X1    g00439(.A1(new_n624_), .A2(new_n193_), .ZN(new_n632_));
  INV_X1     g00440(.I(new_n632_), .ZN(new_n633_));
  NOR2_X1    g00441(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1   g00442(.A1(new_n523_), .A2(new_n505_), .A3(new_n507_), .A4(new_n527_), .ZN(new_n635_));
  NOR2_X1    g00443(.A1(new_n562_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1   g00444(.A1(new_n636_), .A2(new_n538_), .ZN(new_n637_));
  INV_X1     g00445(.I(new_n637_), .ZN(new_n638_));
  NOR2_X1    g00446(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1     g00447(.I(new_n639_), .ZN(new_n640_));
  AOI21_X1   g00448(.A1(new_n630_), .A2(new_n618_), .B(new_n640_), .ZN(new_n641_));
  OAI21_X1   g00449(.A1(\asqrt[63] ), .A2(new_n627_), .B(new_n641_), .ZN(\asqrt[56] ));
  NOR2_X1    g00450(.A1(\a[110] ), .A2(\a[111] ), .ZN(new_n643_));
  INV_X1     g00451(.I(new_n643_), .ZN(new_n644_));
  NOR2_X1    g00452(.A1(new_n644_), .A2(\a[112] ), .ZN(new_n645_));
  INV_X1     g00453(.I(new_n645_), .ZN(new_n646_));
  NAND2_X1   g00454(.A1(new_n618_), .A2(new_n604_), .ZN(new_n647_));
  INV_X1     g00455(.I(new_n626_), .ZN(new_n648_));
  AOI21_X1   g00456(.A1(new_n647_), .A2(new_n648_), .B(\asqrt[63] ), .ZN(new_n649_));
  NAND2_X1   g00457(.A1(new_n572_), .A2(new_n218_), .ZN(new_n650_));
  OAI21_X1   g00458(.A1(new_n650_), .A2(new_n615_), .B(new_n588_), .ZN(new_n651_));
  NAND2_X1   g00459(.A1(new_n581_), .A2(new_n572_), .ZN(new_n652_));
  AOI21_X1   g00460(.A1(new_n652_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n653_));
  AOI21_X1   g00461(.A1(new_n653_), .A2(new_n651_), .B(new_n609_), .ZN(new_n654_));
  INV_X1     g00462(.I(new_n623_), .ZN(new_n655_));
  NAND2_X1   g00463(.A1(new_n604_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1   g00464(.A1(new_n656_), .A2(new_n654_), .B(new_n639_), .ZN(new_n657_));
  OAI21_X1   g00465(.A1(new_n649_), .A2(new_n657_), .B(\a[112] ), .ZN(new_n658_));
  AOI21_X1   g00466(.A1(new_n658_), .A2(new_n646_), .B(new_n531_), .ZN(new_n659_));
  INV_X1     g00467(.I(\a[112] ), .ZN(new_n660_));
  AOI21_X1   g00468(.A1(new_n651_), .A2(new_n616_), .B(new_n207_), .ZN(new_n661_));
  OAI21_X1   g00469(.A1(new_n654_), .A2(new_n661_), .B(new_n648_), .ZN(new_n662_));
  NAND2_X1   g00470(.A1(new_n662_), .A2(new_n193_), .ZN(new_n663_));
  AOI21_X1   g00471(.A1(new_n663_), .A2(new_n641_), .B(new_n660_), .ZN(new_n664_));
  NAND4_X1   g00472(.A1(new_n619_), .A2(new_n523_), .A3(new_n527_), .A4(new_n646_), .ZN(new_n665_));
  NOR2_X1    g00473(.A1(new_n665_), .A2(new_n545_), .ZN(new_n666_));
  INV_X1     g00474(.I(new_n666_), .ZN(new_n667_));
  NOR2_X1    g00475(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1   g00476(.A1(new_n663_), .A2(new_n641_), .B(new_n533_), .ZN(new_n669_));
  INV_X1     g00477(.I(\a[113] ), .ZN(new_n670_));
  AOI21_X1   g00478(.A1(\asqrt[56] ), .A2(new_n660_), .B(new_n670_), .ZN(new_n671_));
  NOR3_X1    g00479(.A1(new_n668_), .A2(new_n671_), .A3(new_n669_), .ZN(new_n672_));
  OAI21_X1   g00480(.A1(new_n672_), .A2(new_n659_), .B(\asqrt[58] ), .ZN(new_n673_));
  OAI21_X1   g00481(.A1(new_n649_), .A2(new_n657_), .B(new_n532_), .ZN(new_n674_));
  NAND2_X1   g00482(.A1(new_n630_), .A2(new_n618_), .ZN(new_n675_));
  INV_X1     g00483(.I(new_n634_), .ZN(new_n676_));
  NOR2_X1    g00484(.A1(new_n638_), .A2(new_n531_), .ZN(new_n677_));
  NAND4_X1   g00485(.A1(new_n663_), .A2(new_n675_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n678_));
  AOI21_X1   g00486(.A1(new_n678_), .A2(new_n674_), .B(new_n535_), .ZN(new_n679_));
  INV_X1     g00487(.I(new_n675_), .ZN(new_n680_));
  NAND2_X1   g00488(.A1(new_n676_), .A2(new_n677_), .ZN(new_n681_));
  NOR3_X1    g00489(.A1(new_n680_), .A2(new_n649_), .A3(new_n681_), .ZN(new_n682_));
  NOR3_X1    g00490(.A1(new_n682_), .A2(new_n669_), .A3(\a[114] ), .ZN(new_n683_));
  AOI21_X1   g00491(.A1(\asqrt[56] ), .A2(\a[112] ), .B(new_n645_), .ZN(new_n684_));
  OAI21_X1   g00492(.A1(new_n684_), .A2(new_n531_), .B(new_n436_), .ZN(new_n685_));
  OAI22_X1   g00493(.A1(new_n672_), .A2(new_n685_), .B1(new_n679_), .B2(new_n683_), .ZN(new_n686_));
  AOI21_X1   g00494(.A1(new_n686_), .A2(new_n673_), .B(new_n327_), .ZN(new_n687_));
  NOR3_X1    g00495(.A1(new_n578_), .A2(new_n577_), .A3(new_n591_), .ZN(new_n688_));
  NAND3_X1   g00496(.A1(\asqrt[56] ), .A2(new_n540_), .A3(new_n555_), .ZN(new_n689_));
  AOI22_X1   g00497(.A1(new_n689_), .A2(new_n578_), .B1(\asqrt[56] ), .B2(new_n688_), .ZN(new_n690_));
  OAI21_X1   g00498(.A1(new_n664_), .A2(new_n645_), .B(\asqrt[57] ), .ZN(new_n691_));
  AOI21_X1   g00499(.A1(new_n663_), .A2(new_n641_), .B(\a[112] ), .ZN(new_n692_));
  OAI21_X1   g00500(.A1(new_n670_), .A2(new_n692_), .B(new_n674_), .ZN(new_n693_));
  OAI21_X1   g00501(.A1(new_n693_), .A2(new_n668_), .B(new_n691_), .ZN(new_n694_));
  AOI21_X1   g00502(.A1(new_n694_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n695_));
  AOI21_X1   g00503(.A1(new_n695_), .A2(new_n686_), .B(new_n690_), .ZN(new_n696_));
  OAI21_X1   g00504(.A1(new_n696_), .A2(new_n687_), .B(\asqrt[60] ), .ZN(new_n697_));
  INV_X1     g00505(.I(new_n697_), .ZN(new_n698_));
  NOR2_X1    g00506(.A1(new_n596_), .A2(new_n597_), .ZN(new_n699_));
  NOR2_X1    g00507(.A1(new_n594_), .A2(new_n599_), .ZN(new_n700_));
  INV_X1     g00508(.I(new_n700_), .ZN(new_n701_));
  NAND4_X1   g00509(.A1(\asqrt[56] ), .A2(new_n595_), .A3(new_n699_), .A4(new_n701_), .ZN(new_n702_));
  INV_X1     g00510(.I(\asqrt[56] ), .ZN(new_n703_));
  NOR3_X1    g00511(.A1(new_n703_), .A2(new_n560_), .A3(new_n700_), .ZN(new_n704_));
  OAI21_X1   g00512(.A1(new_n704_), .A2(new_n699_), .B(new_n702_), .ZN(new_n705_));
  INV_X1     g00513(.I(new_n705_), .ZN(new_n706_));
  NOR3_X1    g00514(.A1(new_n696_), .A2(new_n687_), .A3(\asqrt[60] ), .ZN(new_n707_));
  NOR2_X1    g00515(.A1(new_n707_), .A2(new_n706_), .ZN(new_n708_));
  OAI21_X1   g00516(.A1(new_n708_), .A2(new_n698_), .B(\asqrt[61] ), .ZN(new_n709_));
  NOR2_X1    g00517(.A1(new_n580_), .A2(new_n571_), .ZN(new_n710_));
  NOR3_X1    g00518(.A1(new_n703_), .A2(new_n601_), .A3(new_n710_), .ZN(new_n711_));
  INV_X1     g00519(.I(new_n711_), .ZN(new_n712_));
  NOR3_X1    g00520(.A1(new_n710_), .A2(new_n601_), .A3(new_n576_), .ZN(new_n713_));
  AOI22_X1   g00521(.A1(new_n712_), .A2(new_n576_), .B1(\asqrt[56] ), .B2(new_n713_), .ZN(new_n714_));
  INV_X1     g00522(.I(new_n714_), .ZN(new_n715_));
  NAND2_X1   g00523(.A1(new_n697_), .A2(new_n218_), .ZN(new_n716_));
  OAI21_X1   g00524(.A1(new_n708_), .A2(new_n716_), .B(new_n715_), .ZN(new_n717_));
  AOI21_X1   g00525(.A1(new_n717_), .A2(new_n709_), .B(new_n207_), .ZN(new_n718_));
  NOR3_X1    g00526(.A1(new_n582_), .A2(new_n628_), .A3(new_n588_), .ZN(new_n719_));
  NOR3_X1    g00527(.A1(new_n703_), .A2(new_n582_), .A3(new_n628_), .ZN(new_n720_));
  INV_X1     g00528(.I(new_n720_), .ZN(new_n721_));
  AOI22_X1   g00529(.A1(new_n721_), .A2(new_n588_), .B1(\asqrt[56] ), .B2(new_n719_), .ZN(new_n722_));
  OAI21_X1   g00530(.A1(new_n706_), .A2(new_n707_), .B(new_n697_), .ZN(new_n723_));
  AOI21_X1   g00531(.A1(new_n723_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n724_));
  AOI21_X1   g00532(.A1(new_n724_), .A2(new_n717_), .B(new_n722_), .ZN(new_n725_));
  NOR2_X1    g00533(.A1(new_n617_), .A2(new_n603_), .ZN(new_n726_));
  NOR3_X1    g00534(.A1(new_n661_), .A2(new_n726_), .A3(new_n610_), .ZN(new_n727_));
  NAND2_X1   g00535(.A1(\asqrt[56] ), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1   g00536(.A1(new_n603_), .A2(new_n617_), .B(new_n604_), .ZN(new_n729_));
  OAI21_X1   g00537(.A1(new_n703_), .A2(new_n729_), .B(new_n610_), .ZN(new_n730_));
  NAND2_X1   g00538(.A1(new_n730_), .A2(new_n728_), .ZN(new_n731_));
  INV_X1     g00539(.I(new_n731_), .ZN(new_n732_));
  INV_X1     g00540(.I(new_n647_), .ZN(new_n733_));
  NOR2_X1    g00541(.A1(new_n733_), .A2(new_n655_), .ZN(new_n734_));
  NAND2_X1   g00542(.A1(\asqrt[56] ), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1   g00543(.A1(new_n735_), .A2(new_n675_), .ZN(new_n736_));
  NOR2_X1    g00544(.A1(new_n732_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1   g00545(.A1(new_n725_), .A2(new_n718_), .B(new_n737_), .ZN(new_n738_));
  NAND2_X1   g00546(.A1(new_n738_), .A2(new_n193_), .ZN(new_n739_));
  NAND2_X1   g00547(.A1(new_n658_), .A2(new_n666_), .ZN(new_n740_));
  OAI21_X1   g00548(.A1(new_n649_), .A2(new_n657_), .B(new_n660_), .ZN(new_n741_));
  NAND2_X1   g00549(.A1(new_n741_), .A2(\a[113] ), .ZN(new_n742_));
  NAND3_X1   g00550(.A1(new_n740_), .A2(new_n742_), .A3(new_n674_), .ZN(new_n743_));
  AOI21_X1   g00551(.A1(new_n743_), .A2(new_n691_), .B(new_n436_), .ZN(new_n744_));
  OAI21_X1   g00552(.A1(new_n682_), .A2(new_n669_), .B(\a[114] ), .ZN(new_n745_));
  NAND3_X1   g00553(.A1(new_n678_), .A2(new_n674_), .A3(new_n535_), .ZN(new_n746_));
  NAND2_X1   g00554(.A1(new_n658_), .A2(new_n646_), .ZN(new_n747_));
  AOI21_X1   g00555(.A1(new_n747_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n748_));
  AOI22_X1   g00556(.A1(new_n743_), .A2(new_n748_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n749_));
  OAI21_X1   g00557(.A1(new_n749_), .A2(new_n744_), .B(\asqrt[59] ), .ZN(new_n750_));
  NAND2_X1   g00558(.A1(new_n750_), .A2(new_n306_), .ZN(new_n751_));
  OAI21_X1   g00559(.A1(new_n751_), .A2(new_n696_), .B(new_n705_), .ZN(new_n752_));
  INV_X1     g00560(.I(new_n690_), .ZN(new_n753_));
  AOI21_X1   g00561(.A1(\a[113] ), .A2(new_n741_), .B(new_n669_), .ZN(new_n754_));
  AOI21_X1   g00562(.A1(new_n754_), .A2(new_n740_), .B(new_n659_), .ZN(new_n755_));
  OAI21_X1   g00563(.A1(new_n755_), .A2(new_n436_), .B(new_n327_), .ZN(new_n756_));
  OAI21_X1   g00564(.A1(new_n756_), .A2(new_n749_), .B(new_n753_), .ZN(new_n757_));
  NAND2_X1   g00565(.A1(new_n757_), .A2(new_n750_), .ZN(new_n758_));
  AOI21_X1   g00566(.A1(new_n758_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n759_));
  AOI21_X1   g00567(.A1(new_n759_), .A2(new_n752_), .B(new_n714_), .ZN(new_n760_));
  INV_X1     g00568(.I(new_n722_), .ZN(new_n761_));
  NAND2_X1   g00569(.A1(new_n709_), .A2(new_n207_), .ZN(new_n762_));
  OAI21_X1   g00570(.A1(new_n762_), .A2(new_n760_), .B(new_n761_), .ZN(new_n763_));
  NOR2_X1    g00571(.A1(new_n718_), .A2(new_n731_), .ZN(new_n764_));
  AOI21_X1   g00572(.A1(\asqrt[56] ), .A2(new_n623_), .B(new_n647_), .ZN(new_n765_));
  NOR3_X1    g00573(.A1(new_n765_), .A2(new_n193_), .A3(new_n734_), .ZN(new_n766_));
  NAND4_X1   g00574(.A1(new_n676_), .A2(new_n620_), .A3(new_n622_), .A4(new_n637_), .ZN(new_n767_));
  NOR2_X1    g00575(.A1(new_n680_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1   g00576(.A1(new_n768_), .A2(new_n663_), .ZN(new_n769_));
  INV_X1     g00577(.I(new_n769_), .ZN(new_n770_));
  NOR2_X1    g00578(.A1(new_n766_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1     g00579(.I(new_n771_), .ZN(new_n772_));
  AOI21_X1   g00580(.A1(new_n764_), .A2(new_n763_), .B(new_n772_), .ZN(new_n773_));
  NAND2_X1   g00581(.A1(new_n739_), .A2(new_n773_), .ZN(\asqrt[55] ));
  NOR2_X1    g00582(.A1(\a[108] ), .A2(\a[109] ), .ZN(new_n775_));
  INV_X1     g00583(.I(new_n775_), .ZN(new_n776_));
  NOR2_X1    g00584(.A1(new_n776_), .A2(\a[110] ), .ZN(new_n777_));
  INV_X1     g00585(.I(new_n777_), .ZN(new_n778_));
  AOI21_X1   g00586(.A1(new_n752_), .A2(new_n697_), .B(new_n218_), .ZN(new_n779_));
  OAI21_X1   g00587(.A1(new_n760_), .A2(new_n779_), .B(\asqrt[62] ), .ZN(new_n780_));
  NOR3_X1    g00588(.A1(new_n760_), .A2(new_n779_), .A3(\asqrt[62] ), .ZN(new_n781_));
  OAI21_X1   g00589(.A1(new_n722_), .A2(new_n781_), .B(new_n780_), .ZN(new_n782_));
  AOI21_X1   g00590(.A1(new_n782_), .A2(new_n737_), .B(\asqrt[63] ), .ZN(new_n783_));
  NAND2_X1   g00591(.A1(new_n780_), .A2(new_n732_), .ZN(new_n784_));
  OAI21_X1   g00592(.A1(new_n784_), .A2(new_n725_), .B(new_n771_), .ZN(new_n785_));
  OAI21_X1   g00593(.A1(new_n783_), .A2(new_n785_), .B(\a[110] ), .ZN(new_n786_));
  AOI21_X1   g00594(.A1(new_n786_), .A2(new_n778_), .B(new_n703_), .ZN(new_n787_));
  NAND2_X1   g00595(.A1(new_n637_), .A2(new_n778_), .ZN(new_n788_));
  NOR4_X1    g00596(.A1(new_n680_), .A2(new_n649_), .A3(new_n634_), .A4(new_n788_), .ZN(new_n789_));
  NAND2_X1   g00597(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1   g00598(.A1(new_n739_), .A2(new_n773_), .B(new_n644_), .ZN(new_n791_));
  INV_X1     g00599(.I(\a[110] ), .ZN(new_n792_));
  OAI21_X1   g00600(.A1(new_n783_), .A2(new_n785_), .B(new_n792_), .ZN(new_n793_));
  AOI21_X1   g00601(.A1(\a[111] ), .A2(new_n793_), .B(new_n791_), .ZN(new_n794_));
  AOI21_X1   g00602(.A1(new_n794_), .A2(new_n790_), .B(new_n787_), .ZN(new_n795_));
  NOR2_X1    g00603(.A1(new_n795_), .A2(new_n531_), .ZN(new_n796_));
  NAND2_X1   g00604(.A1(new_n794_), .A2(new_n790_), .ZN(new_n797_));
  OAI21_X1   g00605(.A1(new_n783_), .A2(new_n785_), .B(new_n643_), .ZN(new_n798_));
  NAND2_X1   g00606(.A1(new_n764_), .A2(new_n763_), .ZN(new_n799_));
  INV_X1     g00607(.I(new_n766_), .ZN(new_n800_));
  NOR2_X1    g00608(.A1(new_n770_), .A2(new_n703_), .ZN(new_n801_));
  NAND4_X1   g00609(.A1(new_n739_), .A2(new_n799_), .A3(new_n800_), .A4(new_n801_), .ZN(new_n802_));
  AOI21_X1   g00610(.A1(new_n802_), .A2(new_n798_), .B(new_n660_), .ZN(new_n803_));
  INV_X1     g00611(.I(new_n799_), .ZN(new_n804_));
  NAND2_X1   g00612(.A1(new_n800_), .A2(new_n801_), .ZN(new_n805_));
  NOR3_X1    g00613(.A1(new_n804_), .A2(new_n783_), .A3(new_n805_), .ZN(new_n806_));
  NOR3_X1    g00614(.A1(new_n806_), .A2(\a[112] ), .A3(new_n791_), .ZN(new_n807_));
  NOR2_X1    g00615(.A1(new_n807_), .A2(new_n803_), .ZN(new_n808_));
  NOR2_X1    g00616(.A1(new_n787_), .A2(\asqrt[57] ), .ZN(new_n809_));
  AOI21_X1   g00617(.A1(new_n797_), .A2(new_n809_), .B(new_n808_), .ZN(new_n810_));
  OAI21_X1   g00618(.A1(new_n810_), .A2(new_n796_), .B(\asqrt[58] ), .ZN(new_n811_));
  NOR3_X1    g00619(.A1(new_n754_), .A2(new_n659_), .A3(new_n668_), .ZN(new_n812_));
  NAND3_X1   g00620(.A1(\asqrt[55] ), .A2(new_n691_), .A3(new_n740_), .ZN(new_n813_));
  AOI22_X1   g00621(.A1(new_n813_), .A2(new_n754_), .B1(\asqrt[55] ), .B2(new_n812_), .ZN(new_n814_));
  INV_X1     g00622(.I(new_n814_), .ZN(new_n815_));
  OAI21_X1   g00623(.A1(new_n795_), .A2(new_n531_), .B(new_n436_), .ZN(new_n816_));
  OAI21_X1   g00624(.A1(new_n810_), .A2(new_n816_), .B(new_n815_), .ZN(new_n817_));
  AOI21_X1   g00625(.A1(new_n817_), .A2(new_n811_), .B(new_n327_), .ZN(new_n818_));
  NOR2_X1    g00626(.A1(new_n679_), .A2(new_n683_), .ZN(new_n819_));
  INV_X1     g00627(.I(new_n819_), .ZN(new_n820_));
  NOR2_X1    g00628(.A1(new_n672_), .A2(new_n685_), .ZN(new_n821_));
  NOR3_X1    g00629(.A1(new_n744_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1     g00630(.I(\asqrt[55] ), .ZN(new_n823_));
  OR3_X2     g00631(.A1(new_n823_), .A2(new_n744_), .A3(new_n821_), .Z(new_n824_));
  AOI22_X1   g00632(.A1(new_n824_), .A2(new_n820_), .B1(\asqrt[55] ), .B2(new_n822_), .ZN(new_n825_));
  AOI21_X1   g00633(.A1(new_n739_), .A2(new_n773_), .B(new_n792_), .ZN(new_n826_));
  INV_X1     g00634(.I(new_n789_), .ZN(new_n827_));
  NOR2_X1    g00635(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1     g00636(.I(\a[111] ), .ZN(new_n829_));
  AOI21_X1   g00637(.A1(\asqrt[55] ), .A2(new_n792_), .B(new_n829_), .ZN(new_n830_));
  NOR3_X1    g00638(.A1(new_n828_), .A2(new_n830_), .A3(new_n791_), .ZN(new_n831_));
  OAI21_X1   g00639(.A1(new_n831_), .A2(new_n787_), .B(\asqrt[57] ), .ZN(new_n832_));
  OAI21_X1   g00640(.A1(new_n826_), .A2(new_n777_), .B(\asqrt[56] ), .ZN(new_n833_));
  NAND2_X1   g00641(.A1(new_n833_), .A2(new_n531_), .ZN(new_n834_));
  OAI22_X1   g00642(.A1(new_n831_), .A2(new_n834_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n835_));
  NAND2_X1   g00643(.A1(new_n835_), .A2(new_n832_), .ZN(new_n836_));
  AOI21_X1   g00644(.A1(new_n836_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n837_));
  AOI21_X1   g00645(.A1(new_n837_), .A2(new_n817_), .B(new_n825_), .ZN(new_n838_));
  OAI21_X1   g00646(.A1(new_n838_), .A2(new_n818_), .B(\asqrt[60] ), .ZN(new_n839_));
  NOR2_X1    g00647(.A1(new_n756_), .A2(new_n749_), .ZN(new_n840_));
  NOR3_X1    g00648(.A1(new_n823_), .A2(new_n687_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1     g00649(.I(new_n841_), .ZN(new_n842_));
  NOR3_X1    g00650(.A1(new_n840_), .A2(new_n687_), .A3(new_n753_), .ZN(new_n843_));
  AOI22_X1   g00651(.A1(new_n842_), .A2(new_n753_), .B1(\asqrt[55] ), .B2(new_n843_), .ZN(new_n844_));
  INV_X1     g00652(.I(new_n844_), .ZN(new_n845_));
  AOI21_X1   g00653(.A1(new_n835_), .A2(new_n832_), .B(new_n436_), .ZN(new_n846_));
  AOI21_X1   g00654(.A1(new_n739_), .A2(new_n773_), .B(\a[110] ), .ZN(new_n847_));
  OAI21_X1   g00655(.A1(new_n829_), .A2(new_n847_), .B(new_n798_), .ZN(new_n848_));
  OAI21_X1   g00656(.A1(new_n848_), .A2(new_n828_), .B(new_n833_), .ZN(new_n849_));
  AOI21_X1   g00657(.A1(new_n849_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n850_));
  AOI21_X1   g00658(.A1(new_n850_), .A2(new_n835_), .B(new_n814_), .ZN(new_n851_));
  OAI21_X1   g00659(.A1(new_n851_), .A2(new_n846_), .B(\asqrt[59] ), .ZN(new_n852_));
  NAND2_X1   g00660(.A1(new_n852_), .A2(new_n306_), .ZN(new_n853_));
  OAI21_X1   g00661(.A1(new_n853_), .A2(new_n838_), .B(new_n845_), .ZN(new_n854_));
  AOI21_X1   g00662(.A1(new_n854_), .A2(new_n839_), .B(new_n218_), .ZN(new_n855_));
  NOR3_X1    g00663(.A1(new_n698_), .A2(new_n707_), .A3(new_n705_), .ZN(new_n856_));
  NOR3_X1    g00664(.A1(new_n823_), .A2(new_n698_), .A3(new_n707_), .ZN(new_n857_));
  INV_X1     g00665(.I(new_n857_), .ZN(new_n858_));
  AOI22_X1   g00666(.A1(new_n858_), .A2(new_n705_), .B1(\asqrt[55] ), .B2(new_n856_), .ZN(new_n859_));
  NOR3_X1    g00667(.A1(new_n851_), .A2(new_n846_), .A3(\asqrt[59] ), .ZN(new_n860_));
  OAI21_X1   g00668(.A1(new_n825_), .A2(new_n860_), .B(new_n852_), .ZN(new_n861_));
  AOI21_X1   g00669(.A1(new_n861_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n862_));
  AOI21_X1   g00670(.A1(new_n862_), .A2(new_n854_), .B(new_n859_), .ZN(new_n863_));
  OAI21_X1   g00671(.A1(new_n863_), .A2(new_n855_), .B(\asqrt[62] ), .ZN(new_n864_));
  NOR2_X1    g00672(.A1(new_n708_), .A2(new_n716_), .ZN(new_n865_));
  NOR3_X1    g00673(.A1(new_n823_), .A2(new_n779_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1     g00674(.I(new_n866_), .ZN(new_n867_));
  NOR3_X1    g00675(.A1(new_n865_), .A2(new_n779_), .A3(new_n715_), .ZN(new_n868_));
  AOI22_X1   g00676(.A1(new_n867_), .A2(new_n715_), .B1(\asqrt[55] ), .B2(new_n868_), .ZN(new_n869_));
  NOR3_X1    g00677(.A1(new_n863_), .A2(\asqrt[62] ), .A3(new_n855_), .ZN(new_n870_));
  OAI21_X1   g00678(.A1(new_n869_), .A2(new_n870_), .B(new_n864_), .ZN(new_n871_));
  NOR3_X1    g00679(.A1(new_n718_), .A2(new_n781_), .A3(new_n761_), .ZN(new_n872_));
  NAND2_X1   g00680(.A1(\asqrt[55] ), .A2(new_n872_), .ZN(new_n873_));
  INV_X1     g00681(.I(new_n873_), .ZN(new_n874_));
  NOR2_X1    g00682(.A1(new_n718_), .A2(new_n781_), .ZN(new_n875_));
  AOI21_X1   g00683(.A1(\asqrt[55] ), .A2(new_n875_), .B(new_n722_), .ZN(new_n876_));
  NOR2_X1    g00684(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1     g00685(.I(new_n782_), .ZN(new_n878_));
  NOR3_X1    g00686(.A1(new_n823_), .A2(new_n878_), .A3(new_n732_), .ZN(new_n879_));
  NOR3_X1    g00687(.A1(new_n877_), .A2(new_n804_), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1   g00688(.A1(new_n871_), .A2(new_n880_), .B(\asqrt[63] ), .ZN(new_n881_));
  INV_X1     g00689(.I(new_n825_), .ZN(new_n882_));
  NAND2_X1   g00690(.A1(new_n811_), .A2(new_n327_), .ZN(new_n883_));
  OAI21_X1   g00691(.A1(new_n883_), .A2(new_n851_), .B(new_n882_), .ZN(new_n884_));
  NOR2_X1    g00692(.A1(new_n818_), .A2(\asqrt[60] ), .ZN(new_n885_));
  AOI21_X1   g00693(.A1(new_n885_), .A2(new_n884_), .B(new_n844_), .ZN(new_n886_));
  INV_X1     g00694(.I(new_n859_), .ZN(new_n887_));
  NAND2_X1   g00695(.A1(new_n839_), .A2(new_n218_), .ZN(new_n888_));
  OAI21_X1   g00696(.A1(new_n888_), .A2(new_n886_), .B(new_n887_), .ZN(new_n889_));
  NAND2_X1   g00697(.A1(new_n854_), .A2(new_n839_), .ZN(new_n890_));
  AOI21_X1   g00698(.A1(new_n890_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n891_));
  AOI21_X1   g00699(.A1(new_n891_), .A2(new_n889_), .B(new_n869_), .ZN(new_n892_));
  NAND2_X1   g00700(.A1(new_n864_), .A2(new_n877_), .ZN(new_n893_));
  OAI21_X1   g00701(.A1(new_n823_), .A2(new_n732_), .B(new_n878_), .ZN(new_n894_));
  AOI21_X1   g00702(.A1(new_n782_), .A2(new_n731_), .B(new_n193_), .ZN(new_n895_));
  NAND2_X1   g00703(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1     g00704(.I(new_n896_), .ZN(new_n897_));
  NAND4_X1   g00705(.A1(new_n800_), .A2(new_n730_), .A3(new_n728_), .A4(new_n769_), .ZN(new_n898_));
  NOR2_X1    g00706(.A1(new_n804_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1   g00707(.A1(new_n899_), .A2(new_n739_), .ZN(new_n900_));
  INV_X1     g00708(.I(new_n900_), .ZN(new_n901_));
  NOR2_X1    g00709(.A1(new_n897_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1   g00710(.A1(new_n893_), .A2(new_n892_), .B(new_n902_), .ZN(new_n903_));
  NOR2_X1    g00711(.A1(new_n881_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1    g00712(.A1(\a[106] ), .A2(\a[107] ), .ZN(new_n905_));
  INV_X1     g00713(.I(new_n905_), .ZN(new_n906_));
  NOR2_X1    g00714(.A1(new_n906_), .A2(\a[108] ), .ZN(new_n907_));
  INV_X1     g00715(.I(new_n907_), .ZN(new_n908_));
  OAI21_X1   g00716(.A1(new_n881_), .A2(new_n903_), .B(\a[108] ), .ZN(new_n909_));
  AOI21_X1   g00717(.A1(new_n909_), .A2(new_n908_), .B(new_n823_), .ZN(new_n910_));
  INV_X1     g00718(.I(\a[108] ), .ZN(new_n911_));
  AOI21_X1   g00719(.A1(new_n884_), .A2(new_n852_), .B(new_n306_), .ZN(new_n912_));
  OAI21_X1   g00720(.A1(new_n886_), .A2(new_n912_), .B(\asqrt[61] ), .ZN(new_n913_));
  AOI21_X1   g00721(.A1(new_n889_), .A2(new_n913_), .B(new_n207_), .ZN(new_n914_));
  OAI21_X1   g00722(.A1(new_n892_), .A2(new_n914_), .B(new_n880_), .ZN(new_n915_));
  NAND2_X1   g00723(.A1(new_n915_), .A2(new_n193_), .ZN(new_n916_));
  INV_X1     g00724(.I(new_n869_), .ZN(new_n917_));
  NAND2_X1   g00725(.A1(new_n913_), .A2(new_n207_), .ZN(new_n918_));
  OAI21_X1   g00726(.A1(new_n918_), .A2(new_n863_), .B(new_n917_), .ZN(new_n919_));
  NAND2_X1   g00727(.A1(new_n889_), .A2(new_n913_), .ZN(new_n920_));
  INV_X1     g00728(.I(new_n877_), .ZN(new_n921_));
  AOI21_X1   g00729(.A1(new_n920_), .A2(\asqrt[62] ), .B(new_n921_), .ZN(new_n922_));
  INV_X1     g00730(.I(new_n902_), .ZN(new_n923_));
  AOI21_X1   g00731(.A1(new_n922_), .A2(new_n919_), .B(new_n923_), .ZN(new_n924_));
  AOI21_X1   g00732(.A1(new_n916_), .A2(new_n924_), .B(new_n911_), .ZN(new_n925_));
  NOR3_X1    g00733(.A1(new_n766_), .A2(new_n770_), .A3(new_n907_), .ZN(new_n926_));
  NAND3_X1   g00734(.A1(new_n739_), .A2(new_n799_), .A3(new_n926_), .ZN(new_n927_));
  NOR2_X1    g00735(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  OAI21_X1   g00736(.A1(new_n881_), .A2(new_n903_), .B(new_n775_), .ZN(new_n929_));
  INV_X1     g00737(.I(new_n929_), .ZN(new_n930_));
  INV_X1     g00738(.I(\a[109] ), .ZN(new_n931_));
  NAND2_X1   g00739(.A1(new_n916_), .A2(new_n924_), .ZN(\asqrt[54] ));
  AOI21_X1   g00740(.A1(\asqrt[54] ), .A2(new_n911_), .B(new_n931_), .ZN(new_n933_));
  NOR3_X1    g00741(.A1(new_n928_), .A2(new_n933_), .A3(new_n930_), .ZN(new_n934_));
  OAI21_X1   g00742(.A1(new_n934_), .A2(new_n910_), .B(\asqrt[56] ), .ZN(new_n935_));
  NAND2_X1   g00743(.A1(new_n922_), .A2(new_n919_), .ZN(new_n936_));
  NAND3_X1   g00744(.A1(new_n896_), .A2(\asqrt[55] ), .A3(new_n900_), .ZN(new_n937_));
  INV_X1     g00745(.I(new_n937_), .ZN(new_n938_));
  NAND3_X1   g00746(.A1(new_n916_), .A2(new_n936_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1   g00747(.A1(new_n929_), .A2(new_n939_), .B(new_n792_), .ZN(new_n940_));
  AND3_X2    g00748(.A1(new_n929_), .A2(new_n939_), .A3(new_n792_), .Z(new_n941_));
  OAI21_X1   g00749(.A1(new_n925_), .A2(new_n907_), .B(\asqrt[55] ), .ZN(new_n942_));
  NAND2_X1   g00750(.A1(new_n942_), .A2(new_n703_), .ZN(new_n943_));
  OAI22_X1   g00751(.A1(new_n934_), .A2(new_n943_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n944_));
  AOI21_X1   g00752(.A1(new_n944_), .A2(new_n935_), .B(new_n531_), .ZN(new_n945_));
  NOR3_X1    g00753(.A1(new_n794_), .A2(new_n787_), .A3(new_n828_), .ZN(new_n946_));
  NAND3_X1   g00754(.A1(\asqrt[54] ), .A2(new_n833_), .A3(new_n790_), .ZN(new_n947_));
  AOI22_X1   g00755(.A1(new_n947_), .A2(new_n794_), .B1(\asqrt[54] ), .B2(new_n946_), .ZN(new_n948_));
  AOI21_X1   g00756(.A1(new_n916_), .A2(new_n924_), .B(\a[108] ), .ZN(new_n949_));
  OAI21_X1   g00757(.A1(new_n931_), .A2(new_n949_), .B(new_n929_), .ZN(new_n950_));
  OAI21_X1   g00758(.A1(new_n950_), .A2(new_n928_), .B(new_n942_), .ZN(new_n951_));
  AOI21_X1   g00759(.A1(new_n951_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n952_));
  AOI21_X1   g00760(.A1(new_n952_), .A2(new_n944_), .B(new_n948_), .ZN(new_n953_));
  OAI21_X1   g00761(.A1(new_n953_), .A2(new_n945_), .B(\asqrt[58] ), .ZN(new_n954_));
  NOR2_X1    g00762(.A1(new_n831_), .A2(new_n834_), .ZN(new_n955_));
  INV_X1     g00763(.I(new_n955_), .ZN(new_n956_));
  NAND4_X1   g00764(.A1(\asqrt[54] ), .A2(new_n832_), .A3(new_n808_), .A4(new_n956_), .ZN(new_n957_));
  NOR3_X1    g00765(.A1(new_n904_), .A2(new_n796_), .A3(new_n955_), .ZN(new_n958_));
  OAI21_X1   g00766(.A1(new_n958_), .A2(new_n808_), .B(new_n957_), .ZN(new_n959_));
  INV_X1     g00767(.I(new_n927_), .ZN(new_n960_));
  NAND2_X1   g00768(.A1(new_n909_), .A2(new_n960_), .ZN(new_n961_));
  OAI21_X1   g00769(.A1(new_n881_), .A2(new_n903_), .B(new_n911_), .ZN(new_n962_));
  AOI22_X1   g00770(.A1(new_n962_), .A2(\a[109] ), .B1(\asqrt[54] ), .B2(new_n775_), .ZN(new_n963_));
  AOI21_X1   g00771(.A1(new_n963_), .A2(new_n961_), .B(new_n910_), .ZN(new_n964_));
  NOR2_X1    g00772(.A1(new_n964_), .A2(new_n703_), .ZN(new_n965_));
  NAND2_X1   g00773(.A1(new_n963_), .A2(new_n961_), .ZN(new_n966_));
  INV_X1     g00774(.I(new_n940_), .ZN(new_n967_));
  NAND3_X1   g00775(.A1(new_n929_), .A2(new_n939_), .A3(new_n792_), .ZN(new_n968_));
  NOR2_X1    g00776(.A1(new_n910_), .A2(\asqrt[56] ), .ZN(new_n969_));
  AOI22_X1   g00777(.A1(new_n966_), .A2(new_n969_), .B1(new_n967_), .B2(new_n968_), .ZN(new_n970_));
  OAI21_X1   g00778(.A1(new_n970_), .A2(new_n965_), .B(\asqrt[57] ), .ZN(new_n971_));
  NAND2_X1   g00779(.A1(new_n971_), .A2(new_n436_), .ZN(new_n972_));
  OAI21_X1   g00780(.A1(new_n972_), .A2(new_n953_), .B(new_n959_), .ZN(new_n973_));
  AOI21_X1   g00781(.A1(new_n973_), .A2(new_n954_), .B(new_n327_), .ZN(new_n974_));
  NOR2_X1    g00782(.A1(new_n810_), .A2(new_n816_), .ZN(new_n975_));
  NOR3_X1    g00783(.A1(new_n904_), .A2(new_n846_), .A3(new_n975_), .ZN(new_n976_));
  INV_X1     g00784(.I(new_n976_), .ZN(new_n977_));
  NOR3_X1    g00785(.A1(new_n975_), .A2(new_n846_), .A3(new_n815_), .ZN(new_n978_));
  AOI22_X1   g00786(.A1(new_n977_), .A2(new_n815_), .B1(\asqrt[54] ), .B2(new_n978_), .ZN(new_n979_));
  INV_X1     g00787(.I(new_n948_), .ZN(new_n980_));
  OAI21_X1   g00788(.A1(new_n964_), .A2(new_n703_), .B(new_n531_), .ZN(new_n981_));
  OAI21_X1   g00789(.A1(new_n970_), .A2(new_n981_), .B(new_n980_), .ZN(new_n982_));
  NAND2_X1   g00790(.A1(new_n982_), .A2(new_n971_), .ZN(new_n983_));
  AOI21_X1   g00791(.A1(new_n983_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n984_));
  AOI21_X1   g00792(.A1(new_n984_), .A2(new_n973_), .B(new_n979_), .ZN(new_n985_));
  OAI21_X1   g00793(.A1(new_n985_), .A2(new_n974_), .B(\asqrt[60] ), .ZN(new_n986_));
  NOR3_X1    g00794(.A1(new_n818_), .A2(new_n860_), .A3(new_n882_), .ZN(new_n987_));
  NOR3_X1    g00795(.A1(new_n904_), .A2(new_n818_), .A3(new_n860_), .ZN(new_n988_));
  INV_X1     g00796(.I(new_n988_), .ZN(new_n989_));
  AOI22_X1   g00797(.A1(new_n989_), .A2(new_n882_), .B1(\asqrt[54] ), .B2(new_n987_), .ZN(new_n990_));
  INV_X1     g00798(.I(new_n990_), .ZN(new_n991_));
  INV_X1     g00799(.I(new_n954_), .ZN(new_n992_));
  INV_X1     g00800(.I(new_n959_), .ZN(new_n993_));
  NOR3_X1    g00801(.A1(new_n953_), .A2(new_n945_), .A3(\asqrt[58] ), .ZN(new_n994_));
  NOR2_X1    g00802(.A1(new_n994_), .A2(new_n993_), .ZN(new_n995_));
  OAI21_X1   g00803(.A1(new_n995_), .A2(new_n992_), .B(\asqrt[59] ), .ZN(new_n996_));
  NAND2_X1   g00804(.A1(new_n996_), .A2(new_n306_), .ZN(new_n997_));
  OAI21_X1   g00805(.A1(new_n997_), .A2(new_n985_), .B(new_n991_), .ZN(new_n998_));
  AOI21_X1   g00806(.A1(new_n998_), .A2(new_n986_), .B(new_n218_), .ZN(new_n999_));
  NOR2_X1    g00807(.A1(new_n853_), .A2(new_n838_), .ZN(new_n1000_));
  NOR3_X1    g00808(.A1(new_n904_), .A2(new_n912_), .A3(new_n1000_), .ZN(new_n1001_));
  INV_X1     g00809(.I(new_n1001_), .ZN(new_n1002_));
  NOR3_X1    g00810(.A1(new_n912_), .A2(new_n845_), .A3(new_n1000_), .ZN(new_n1003_));
  AOI22_X1   g00811(.A1(new_n1002_), .A2(new_n845_), .B1(\asqrt[54] ), .B2(new_n1003_), .ZN(new_n1004_));
  INV_X1     g00812(.I(new_n979_), .ZN(new_n1005_));
  NAND2_X1   g00813(.A1(new_n954_), .A2(new_n327_), .ZN(new_n1006_));
  OAI21_X1   g00814(.A1(new_n995_), .A2(new_n1006_), .B(new_n1005_), .ZN(new_n1007_));
  AOI21_X1   g00815(.A1(new_n1007_), .A2(new_n996_), .B(new_n306_), .ZN(new_n1008_));
  NOR2_X1    g00816(.A1(new_n1008_), .A2(\asqrt[61] ), .ZN(new_n1009_));
  AOI21_X1   g00817(.A1(new_n1009_), .A2(new_n998_), .B(new_n1004_), .ZN(new_n1010_));
  OAI21_X1   g00818(.A1(new_n1010_), .A2(new_n999_), .B(\asqrt[62] ), .ZN(new_n1011_));
  NOR2_X1    g00819(.A1(new_n888_), .A2(new_n886_), .ZN(new_n1012_));
  NOR3_X1    g00820(.A1(new_n1012_), .A2(new_n855_), .A3(new_n887_), .ZN(new_n1013_));
  NOR3_X1    g00821(.A1(new_n904_), .A2(new_n855_), .A3(new_n1012_), .ZN(new_n1014_));
  INV_X1     g00822(.I(new_n1014_), .ZN(new_n1015_));
  AOI22_X1   g00823(.A1(new_n1015_), .A2(new_n887_), .B1(\asqrt[54] ), .B2(new_n1013_), .ZN(new_n1016_));
  INV_X1     g00824(.I(new_n1016_), .ZN(new_n1017_));
  OAI21_X1   g00825(.A1(new_n993_), .A2(new_n994_), .B(new_n954_), .ZN(new_n1018_));
  AOI21_X1   g00826(.A1(new_n1018_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n1019_));
  AOI21_X1   g00827(.A1(new_n1019_), .A2(new_n1007_), .B(new_n990_), .ZN(new_n1020_));
  OAI21_X1   g00828(.A1(new_n1020_), .A2(new_n1008_), .B(\asqrt[61] ), .ZN(new_n1021_));
  NAND2_X1   g00829(.A1(new_n1021_), .A2(new_n207_), .ZN(new_n1022_));
  OAI21_X1   g00830(.A1(new_n1022_), .A2(new_n1010_), .B(new_n1017_), .ZN(new_n1023_));
  INV_X1     g00831(.I(new_n870_), .ZN(new_n1024_));
  NAND4_X1   g00832(.A1(\asqrt[54] ), .A2(new_n864_), .A3(new_n869_), .A4(new_n1024_), .ZN(new_n1025_));
  NAND2_X1   g00833(.A1(new_n1024_), .A2(new_n864_), .ZN(new_n1026_));
  OAI21_X1   g00834(.A1(new_n904_), .A2(new_n1026_), .B(new_n917_), .ZN(new_n1027_));
  NAND2_X1   g00835(.A1(new_n1025_), .A2(new_n1027_), .ZN(new_n1028_));
  AOI21_X1   g00836(.A1(new_n919_), .A2(new_n864_), .B(new_n877_), .ZN(new_n1029_));
  NAND2_X1   g00837(.A1(\asqrt[54] ), .A2(new_n1029_), .ZN(new_n1030_));
  NAND3_X1   g00838(.A1(new_n1028_), .A2(new_n936_), .A3(new_n1030_), .ZN(new_n1031_));
  AOI21_X1   g00839(.A1(new_n1023_), .A2(new_n1011_), .B(new_n1031_), .ZN(new_n1032_));
  NOR3_X1    g00840(.A1(new_n1020_), .A2(new_n1008_), .A3(\asqrt[61] ), .ZN(new_n1033_));
  OAI21_X1   g00841(.A1(new_n1004_), .A2(new_n1033_), .B(new_n1021_), .ZN(new_n1034_));
  AOI21_X1   g00842(.A1(new_n1034_), .A2(\asqrt[62] ), .B(new_n1028_), .ZN(new_n1035_));
  AOI21_X1   g00843(.A1(\asqrt[54] ), .A2(new_n921_), .B(new_n871_), .ZN(new_n1036_));
  OR3_X2     g00844(.A1(new_n1036_), .A2(new_n193_), .A3(new_n1029_), .Z(new_n1037_));
  INV_X1     g00845(.I(new_n936_), .ZN(new_n1038_));
  NAND2_X1   g00846(.A1(new_n900_), .A2(new_n873_), .ZN(new_n1039_));
  NOR4_X1    g00847(.A1(new_n1038_), .A2(new_n876_), .A3(new_n897_), .A4(new_n1039_), .ZN(new_n1040_));
  NAND2_X1   g00848(.A1(new_n1040_), .A2(new_n916_), .ZN(new_n1041_));
  NAND2_X1   g00849(.A1(new_n1037_), .A2(new_n1041_), .ZN(new_n1042_));
  AOI21_X1   g00850(.A1(new_n1035_), .A2(new_n1023_), .B(new_n1042_), .ZN(new_n1043_));
  OAI21_X1   g00851(.A1(\asqrt[63] ), .A2(new_n1032_), .B(new_n1043_), .ZN(\asqrt[53] ));
  NOR2_X1    g00852(.A1(\a[104] ), .A2(\a[105] ), .ZN(new_n1045_));
  INV_X1     g00853(.I(new_n1045_), .ZN(new_n1046_));
  NOR2_X1    g00854(.A1(new_n1046_), .A2(\a[106] ), .ZN(new_n1047_));
  INV_X1     g00855(.I(new_n1047_), .ZN(new_n1048_));
  NAND2_X1   g00856(.A1(new_n1023_), .A2(new_n1011_), .ZN(new_n1049_));
  INV_X1     g00857(.I(new_n1031_), .ZN(new_n1050_));
  AOI21_X1   g00858(.A1(new_n1049_), .A2(new_n1050_), .B(\asqrt[63] ), .ZN(new_n1051_));
  INV_X1     g00859(.I(new_n1004_), .ZN(new_n1052_));
  NAND2_X1   g00860(.A1(new_n986_), .A2(new_n218_), .ZN(new_n1053_));
  OAI21_X1   g00861(.A1(new_n1053_), .A2(new_n1020_), .B(new_n1052_), .ZN(new_n1054_));
  NOR2_X1    g00862(.A1(new_n999_), .A2(\asqrt[62] ), .ZN(new_n1055_));
  AOI21_X1   g00863(.A1(new_n1055_), .A2(new_n1054_), .B(new_n1016_), .ZN(new_n1056_));
  INV_X1     g00864(.I(new_n1028_), .ZN(new_n1057_));
  NAND2_X1   g00865(.A1(new_n1011_), .A2(new_n1057_), .ZN(new_n1058_));
  INV_X1     g00866(.I(new_n1042_), .ZN(new_n1059_));
  OAI21_X1   g00867(.A1(new_n1058_), .A2(new_n1056_), .B(new_n1059_), .ZN(new_n1060_));
  OAI21_X1   g00868(.A1(new_n1051_), .A2(new_n1060_), .B(\a[106] ), .ZN(new_n1061_));
  AOI21_X1   g00869(.A1(new_n1061_), .A2(new_n1048_), .B(new_n904_), .ZN(new_n1062_));
  INV_X1     g00870(.I(\a[106] ), .ZN(new_n1063_));
  NAND3_X1   g00871(.A1(new_n1054_), .A2(new_n207_), .A3(new_n1021_), .ZN(new_n1064_));
  AOI22_X1   g00872(.A1(new_n1064_), .A2(new_n1017_), .B1(new_n1034_), .B2(\asqrt[62] ), .ZN(new_n1065_));
  OAI21_X1   g00873(.A1(new_n1065_), .A2(new_n1031_), .B(new_n193_), .ZN(new_n1066_));
  AOI21_X1   g00874(.A1(new_n1066_), .A2(new_n1043_), .B(new_n1063_), .ZN(new_n1067_));
  NOR2_X1    g00875(.A1(new_n901_), .A2(new_n1047_), .ZN(new_n1068_));
  NAND4_X1   g00876(.A1(new_n916_), .A2(new_n936_), .A3(new_n896_), .A4(new_n1068_), .ZN(new_n1069_));
  NOR2_X1    g00877(.A1(new_n1067_), .A2(new_n1069_), .ZN(new_n1070_));
  AOI21_X1   g00878(.A1(new_n1066_), .A2(new_n1043_), .B(new_n906_), .ZN(new_n1071_));
  INV_X1     g00879(.I(\a[107] ), .ZN(new_n1072_));
  AOI21_X1   g00880(.A1(\asqrt[53] ), .A2(new_n1063_), .B(new_n1072_), .ZN(new_n1073_));
  NOR3_X1    g00881(.A1(new_n1070_), .A2(new_n1073_), .A3(new_n1071_), .ZN(new_n1074_));
  OAI21_X1   g00882(.A1(new_n1074_), .A2(new_n1062_), .B(\asqrt[55] ), .ZN(new_n1075_));
  OAI21_X1   g00883(.A1(new_n1051_), .A2(new_n1060_), .B(new_n905_), .ZN(new_n1076_));
  NOR2_X1    g00884(.A1(new_n1058_), .A2(new_n1056_), .ZN(new_n1077_));
  OAI21_X1   g00885(.A1(new_n1040_), .A2(new_n924_), .B(new_n916_), .ZN(new_n1078_));
  NAND2_X1   g00886(.A1(new_n1037_), .A2(new_n1078_), .ZN(new_n1079_));
  NOR3_X1    g00887(.A1(new_n1051_), .A2(new_n1077_), .A3(new_n1079_), .ZN(new_n1080_));
  INV_X1     g00888(.I(new_n1080_), .ZN(new_n1081_));
  AOI21_X1   g00889(.A1(new_n1081_), .A2(new_n1076_), .B(new_n911_), .ZN(new_n1082_));
  NOR3_X1    g00890(.A1(new_n1071_), .A2(new_n1080_), .A3(\a[108] ), .ZN(new_n1083_));
  AOI21_X1   g00891(.A1(\asqrt[53] ), .A2(\a[106] ), .B(new_n1047_), .ZN(new_n1084_));
  OAI21_X1   g00892(.A1(new_n1084_), .A2(new_n904_), .B(new_n823_), .ZN(new_n1085_));
  OAI22_X1   g00893(.A1(new_n1074_), .A2(new_n1085_), .B1(new_n1082_), .B2(new_n1083_), .ZN(new_n1086_));
  AOI21_X1   g00894(.A1(new_n1086_), .A2(new_n1075_), .B(new_n703_), .ZN(new_n1087_));
  NOR3_X1    g00895(.A1(new_n963_), .A2(new_n910_), .A3(new_n928_), .ZN(new_n1088_));
  NAND3_X1   g00896(.A1(\asqrt[53] ), .A2(new_n942_), .A3(new_n961_), .ZN(new_n1089_));
  AOI22_X1   g00897(.A1(new_n1089_), .A2(new_n963_), .B1(\asqrt[53] ), .B2(new_n1088_), .ZN(new_n1090_));
  OAI21_X1   g00898(.A1(new_n1067_), .A2(new_n1047_), .B(\asqrt[54] ), .ZN(new_n1091_));
  AOI21_X1   g00899(.A1(new_n1066_), .A2(new_n1043_), .B(\a[106] ), .ZN(new_n1092_));
  OAI21_X1   g00900(.A1(new_n1072_), .A2(new_n1092_), .B(new_n1076_), .ZN(new_n1093_));
  OAI21_X1   g00901(.A1(new_n1093_), .A2(new_n1070_), .B(new_n1091_), .ZN(new_n1094_));
  AOI21_X1   g00902(.A1(new_n1094_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n1095_));
  AOI21_X1   g00903(.A1(new_n1095_), .A2(new_n1086_), .B(new_n1090_), .ZN(new_n1096_));
  OAI21_X1   g00904(.A1(new_n1096_), .A2(new_n1087_), .B(\asqrt[57] ), .ZN(new_n1097_));
  INV_X1     g00905(.I(new_n1097_), .ZN(new_n1098_));
  NOR2_X1    g00906(.A1(new_n941_), .A2(new_n940_), .ZN(new_n1099_));
  NOR2_X1    g00907(.A1(new_n934_), .A2(new_n943_), .ZN(new_n1100_));
  INV_X1     g00908(.I(new_n1100_), .ZN(new_n1101_));
  NAND4_X1   g00909(.A1(\asqrt[53] ), .A2(new_n935_), .A3(new_n1099_), .A4(new_n1101_), .ZN(new_n1102_));
  INV_X1     g00910(.I(\asqrt[53] ), .ZN(new_n1103_));
  NOR3_X1    g00911(.A1(new_n1103_), .A2(new_n965_), .A3(new_n1100_), .ZN(new_n1104_));
  OAI21_X1   g00912(.A1(new_n1104_), .A2(new_n1099_), .B(new_n1102_), .ZN(new_n1105_));
  INV_X1     g00913(.I(new_n1105_), .ZN(new_n1106_));
  NOR3_X1    g00914(.A1(new_n1096_), .A2(new_n1087_), .A3(\asqrt[57] ), .ZN(new_n1107_));
  NOR2_X1    g00915(.A1(new_n1107_), .A2(new_n1106_), .ZN(new_n1108_));
  OAI21_X1   g00916(.A1(new_n1108_), .A2(new_n1098_), .B(\asqrt[58] ), .ZN(new_n1109_));
  NOR2_X1    g00917(.A1(new_n970_), .A2(new_n981_), .ZN(new_n1110_));
  NOR3_X1    g00918(.A1(new_n1103_), .A2(new_n945_), .A3(new_n1110_), .ZN(new_n1111_));
  INV_X1     g00919(.I(new_n1111_), .ZN(new_n1112_));
  NOR3_X1    g00920(.A1(new_n1110_), .A2(new_n945_), .A3(new_n980_), .ZN(new_n1113_));
  AOI22_X1   g00921(.A1(new_n1112_), .A2(new_n980_), .B1(\asqrt[53] ), .B2(new_n1113_), .ZN(new_n1114_));
  INV_X1     g00922(.I(new_n1114_), .ZN(new_n1115_));
  NAND2_X1   g00923(.A1(new_n1097_), .A2(new_n436_), .ZN(new_n1116_));
  OAI21_X1   g00924(.A1(new_n1108_), .A2(new_n1116_), .B(new_n1115_), .ZN(new_n1117_));
  AOI21_X1   g00925(.A1(new_n1117_), .A2(new_n1109_), .B(new_n327_), .ZN(new_n1118_));
  NOR3_X1    g00926(.A1(new_n992_), .A2(new_n994_), .A3(new_n959_), .ZN(new_n1119_));
  NOR3_X1    g00927(.A1(new_n1103_), .A2(new_n992_), .A3(new_n994_), .ZN(new_n1120_));
  INV_X1     g00928(.I(new_n1120_), .ZN(new_n1121_));
  AOI22_X1   g00929(.A1(new_n1121_), .A2(new_n959_), .B1(\asqrt[53] ), .B2(new_n1119_), .ZN(new_n1122_));
  OAI21_X1   g00930(.A1(new_n1106_), .A2(new_n1107_), .B(new_n1097_), .ZN(new_n1123_));
  AOI21_X1   g00931(.A1(new_n1123_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n1124_));
  AOI21_X1   g00932(.A1(new_n1124_), .A2(new_n1117_), .B(new_n1122_), .ZN(new_n1125_));
  OAI21_X1   g00933(.A1(new_n1125_), .A2(new_n1118_), .B(\asqrt[60] ), .ZN(new_n1126_));
  INV_X1     g00934(.I(new_n1126_), .ZN(new_n1127_));
  NOR2_X1    g00935(.A1(new_n995_), .A2(new_n1006_), .ZN(new_n1128_));
  NOR3_X1    g00936(.A1(new_n1103_), .A2(new_n974_), .A3(new_n1128_), .ZN(new_n1129_));
  INV_X1     g00937(.I(new_n1129_), .ZN(new_n1130_));
  NOR3_X1    g00938(.A1(new_n1128_), .A2(new_n974_), .A3(new_n1005_), .ZN(new_n1131_));
  AOI22_X1   g00939(.A1(new_n1130_), .A2(new_n1005_), .B1(\asqrt[53] ), .B2(new_n1131_), .ZN(new_n1132_));
  NOR3_X1    g00940(.A1(new_n1125_), .A2(new_n1118_), .A3(\asqrt[60] ), .ZN(new_n1133_));
  NOR2_X1    g00941(.A1(new_n1133_), .A2(new_n1132_), .ZN(new_n1134_));
  OAI21_X1   g00942(.A1(new_n1134_), .A2(new_n1127_), .B(\asqrt[61] ), .ZN(new_n1135_));
  NOR2_X1    g00943(.A1(new_n997_), .A2(new_n985_), .ZN(new_n1136_));
  NOR3_X1    g00944(.A1(new_n1136_), .A2(new_n1008_), .A3(new_n991_), .ZN(new_n1137_));
  NOR3_X1    g00945(.A1(new_n1103_), .A2(new_n1008_), .A3(new_n1136_), .ZN(new_n1138_));
  INV_X1     g00946(.I(new_n1138_), .ZN(new_n1139_));
  AOI22_X1   g00947(.A1(new_n1139_), .A2(new_n991_), .B1(\asqrt[53] ), .B2(new_n1137_), .ZN(new_n1140_));
  INV_X1     g00948(.I(new_n1140_), .ZN(new_n1141_));
  NAND2_X1   g00949(.A1(new_n1126_), .A2(new_n218_), .ZN(new_n1142_));
  OAI21_X1   g00950(.A1(new_n1134_), .A2(new_n1142_), .B(new_n1141_), .ZN(new_n1143_));
  AOI21_X1   g00951(.A1(new_n1143_), .A2(new_n1135_), .B(new_n207_), .ZN(new_n1144_));
  NOR3_X1    g00952(.A1(new_n1103_), .A2(new_n999_), .A3(new_n1033_), .ZN(new_n1145_));
  INV_X1     g00953(.I(new_n1145_), .ZN(new_n1146_));
  NOR3_X1    g00954(.A1(new_n999_), .A2(new_n1033_), .A3(new_n1052_), .ZN(new_n1147_));
  AOI22_X1   g00955(.A1(new_n1146_), .A2(new_n1052_), .B1(\asqrt[53] ), .B2(new_n1147_), .ZN(new_n1148_));
  OAI21_X1   g00956(.A1(new_n1132_), .A2(new_n1133_), .B(new_n1126_), .ZN(new_n1149_));
  AOI21_X1   g00957(.A1(new_n1149_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n1150_));
  AOI21_X1   g00958(.A1(new_n1150_), .A2(new_n1143_), .B(new_n1148_), .ZN(new_n1151_));
  AND3_X2    g00959(.A1(new_n1011_), .A2(new_n1016_), .A3(new_n1064_), .Z(new_n1152_));
  AND3_X2    g00960(.A1(\asqrt[53] ), .A2(new_n1011_), .A3(new_n1064_), .Z(new_n1153_));
  NOR2_X1    g00961(.A1(new_n1153_), .A2(new_n1016_), .ZN(new_n1154_));
  AOI21_X1   g00962(.A1(\asqrt[53] ), .A2(new_n1152_), .B(new_n1154_), .ZN(new_n1155_));
  NOR3_X1    g00963(.A1(new_n1103_), .A2(new_n1065_), .A3(new_n1057_), .ZN(new_n1156_));
  NOR3_X1    g00964(.A1(new_n1155_), .A2(new_n1077_), .A3(new_n1156_), .ZN(new_n1157_));
  OAI21_X1   g00965(.A1(new_n1151_), .A2(new_n1144_), .B(new_n1157_), .ZN(new_n1158_));
  NAND2_X1   g00966(.A1(new_n1158_), .A2(new_n193_), .ZN(new_n1159_));
  INV_X1     g00967(.I(new_n1132_), .ZN(new_n1160_));
  INV_X1     g00968(.I(new_n1069_), .ZN(new_n1161_));
  NAND2_X1   g00969(.A1(new_n1061_), .A2(new_n1161_), .ZN(new_n1162_));
  OAI21_X1   g00970(.A1(new_n1051_), .A2(new_n1060_), .B(new_n1063_), .ZN(new_n1163_));
  NAND2_X1   g00971(.A1(new_n1163_), .A2(\a[107] ), .ZN(new_n1164_));
  NAND3_X1   g00972(.A1(new_n1162_), .A2(new_n1164_), .A3(new_n1076_), .ZN(new_n1165_));
  AOI21_X1   g00973(.A1(new_n1165_), .A2(new_n1091_), .B(new_n823_), .ZN(new_n1166_));
  OAI21_X1   g00974(.A1(new_n1071_), .A2(new_n1080_), .B(\a[108] ), .ZN(new_n1167_));
  NAND3_X1   g00975(.A1(new_n1081_), .A2(new_n1076_), .A3(new_n911_), .ZN(new_n1168_));
  NAND2_X1   g00976(.A1(new_n1061_), .A2(new_n1048_), .ZN(new_n1169_));
  AOI21_X1   g00977(.A1(new_n1169_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1170_));
  AOI22_X1   g00978(.A1(new_n1165_), .A2(new_n1170_), .B1(new_n1167_), .B2(new_n1168_), .ZN(new_n1171_));
  OAI21_X1   g00979(.A1(new_n1171_), .A2(new_n1166_), .B(\asqrt[56] ), .ZN(new_n1172_));
  NAND2_X1   g00980(.A1(new_n1172_), .A2(new_n531_), .ZN(new_n1173_));
  OAI21_X1   g00981(.A1(new_n1173_), .A2(new_n1096_), .B(new_n1105_), .ZN(new_n1174_));
  AOI21_X1   g00982(.A1(new_n1174_), .A2(new_n1097_), .B(new_n436_), .ZN(new_n1175_));
  INV_X1     g00983(.I(new_n1090_), .ZN(new_n1176_));
  AOI21_X1   g00984(.A1(\a[107] ), .A2(new_n1163_), .B(new_n1071_), .ZN(new_n1177_));
  AOI21_X1   g00985(.A1(new_n1177_), .A2(new_n1162_), .B(new_n1062_), .ZN(new_n1178_));
  OAI21_X1   g00986(.A1(new_n1178_), .A2(new_n823_), .B(new_n703_), .ZN(new_n1179_));
  OAI21_X1   g00987(.A1(new_n1179_), .A2(new_n1171_), .B(new_n1176_), .ZN(new_n1180_));
  NAND2_X1   g00988(.A1(new_n1180_), .A2(new_n1172_), .ZN(new_n1181_));
  AOI21_X1   g00989(.A1(new_n1181_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n1182_));
  AOI21_X1   g00990(.A1(new_n1182_), .A2(new_n1174_), .B(new_n1114_), .ZN(new_n1183_));
  OAI21_X1   g00991(.A1(new_n1183_), .A2(new_n1175_), .B(\asqrt[59] ), .ZN(new_n1184_));
  NAND2_X1   g00992(.A1(new_n1184_), .A2(new_n306_), .ZN(new_n1185_));
  OAI21_X1   g00993(.A1(new_n1185_), .A2(new_n1125_), .B(new_n1160_), .ZN(new_n1186_));
  NOR3_X1    g00994(.A1(new_n1183_), .A2(new_n1175_), .A3(\asqrt[59] ), .ZN(new_n1187_));
  OAI21_X1   g00995(.A1(new_n1122_), .A2(new_n1187_), .B(new_n1184_), .ZN(new_n1188_));
  AOI21_X1   g00996(.A1(new_n1188_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n1189_));
  AOI21_X1   g00997(.A1(new_n1189_), .A2(new_n1186_), .B(new_n1140_), .ZN(new_n1190_));
  INV_X1     g00998(.I(new_n1148_), .ZN(new_n1191_));
  NAND2_X1   g00999(.A1(new_n1135_), .A2(new_n207_), .ZN(new_n1192_));
  OAI21_X1   g01000(.A1(new_n1192_), .A2(new_n1190_), .B(new_n1191_), .ZN(new_n1193_));
  INV_X1     g01001(.I(new_n1155_), .ZN(new_n1194_));
  NOR2_X1    g01002(.A1(new_n1144_), .A2(new_n1194_), .ZN(new_n1195_));
  NOR2_X1    g01003(.A1(new_n1065_), .A2(new_n1057_), .ZN(new_n1196_));
  AOI21_X1   g01004(.A1(\asqrt[53] ), .A2(new_n1028_), .B(new_n1049_), .ZN(new_n1197_));
  NOR3_X1    g01005(.A1(new_n1197_), .A2(new_n193_), .A3(new_n1196_), .ZN(new_n1198_));
  INV_X1     g01006(.I(new_n1077_), .ZN(new_n1199_));
  AND3_X2    g01007(.A1(new_n1041_), .A2(new_n1025_), .A3(new_n1027_), .Z(new_n1200_));
  NAND4_X1   g01008(.A1(new_n1199_), .A2(new_n1066_), .A3(new_n1037_), .A4(new_n1200_), .ZN(new_n1201_));
  INV_X1     g01009(.I(new_n1201_), .ZN(new_n1202_));
  NOR2_X1    g01010(.A1(new_n1198_), .A2(new_n1202_), .ZN(new_n1203_));
  INV_X1     g01011(.I(new_n1203_), .ZN(new_n1204_));
  AOI21_X1   g01012(.A1(new_n1195_), .A2(new_n1193_), .B(new_n1204_), .ZN(new_n1205_));
  NAND2_X1   g01013(.A1(new_n1159_), .A2(new_n1205_), .ZN(\asqrt[52] ));
  NOR2_X1    g01014(.A1(\a[102] ), .A2(\a[103] ), .ZN(new_n1207_));
  INV_X1     g01015(.I(new_n1207_), .ZN(new_n1208_));
  NOR2_X1    g01016(.A1(new_n1208_), .A2(\a[104] ), .ZN(new_n1209_));
  INV_X1     g01017(.I(new_n1209_), .ZN(new_n1210_));
  NAND3_X1   g01018(.A1(new_n1186_), .A2(new_n218_), .A3(new_n1126_), .ZN(new_n1211_));
  AOI22_X1   g01019(.A1(new_n1211_), .A2(new_n1141_), .B1(new_n1149_), .B2(\asqrt[61] ), .ZN(new_n1212_));
  AOI21_X1   g01020(.A1(new_n1186_), .A2(new_n1126_), .B(new_n218_), .ZN(new_n1213_));
  NOR3_X1    g01021(.A1(new_n1190_), .A2(\asqrt[62] ), .A3(new_n1213_), .ZN(new_n1214_));
  OAI22_X1   g01022(.A1(new_n1214_), .A2(new_n1148_), .B1(new_n1212_), .B2(new_n207_), .ZN(new_n1215_));
  AOI21_X1   g01023(.A1(new_n1215_), .A2(new_n1157_), .B(\asqrt[63] ), .ZN(new_n1216_));
  OAI21_X1   g01024(.A1(new_n1212_), .A2(new_n207_), .B(new_n1155_), .ZN(new_n1217_));
  OAI21_X1   g01025(.A1(new_n1217_), .A2(new_n1151_), .B(new_n1203_), .ZN(new_n1218_));
  OAI21_X1   g01026(.A1(new_n1216_), .A2(new_n1218_), .B(\a[104] ), .ZN(new_n1219_));
  AOI21_X1   g01027(.A1(new_n1219_), .A2(new_n1210_), .B(new_n1103_), .ZN(new_n1220_));
  INV_X1     g01028(.I(\a[104] ), .ZN(new_n1221_));
  AOI21_X1   g01029(.A1(new_n1159_), .A2(new_n1205_), .B(new_n1221_), .ZN(new_n1222_));
  NAND4_X1   g01030(.A1(new_n1199_), .A2(new_n1037_), .A3(new_n1041_), .A4(new_n1210_), .ZN(new_n1223_));
  NOR2_X1    g01031(.A1(new_n1223_), .A2(new_n1051_), .ZN(new_n1224_));
  INV_X1     g01032(.I(new_n1224_), .ZN(new_n1225_));
  NOR2_X1    g01033(.A1(new_n1222_), .A2(new_n1225_), .ZN(new_n1226_));
  AOI21_X1   g01034(.A1(new_n1159_), .A2(new_n1205_), .B(new_n1046_), .ZN(new_n1227_));
  INV_X1     g01035(.I(\a[105] ), .ZN(new_n1228_));
  AOI21_X1   g01036(.A1(\asqrt[52] ), .A2(new_n1221_), .B(new_n1228_), .ZN(new_n1229_));
  NOR3_X1    g01037(.A1(new_n1226_), .A2(new_n1229_), .A3(new_n1227_), .ZN(new_n1230_));
  OAI21_X1   g01038(.A1(new_n1230_), .A2(new_n1220_), .B(\asqrt[54] ), .ZN(new_n1231_));
  OAI21_X1   g01039(.A1(new_n1216_), .A2(new_n1218_), .B(new_n1045_), .ZN(new_n1232_));
  NAND2_X1   g01040(.A1(new_n1195_), .A2(new_n1193_), .ZN(new_n1233_));
  NOR3_X1    g01041(.A1(new_n1198_), .A2(new_n1103_), .A3(new_n1202_), .ZN(new_n1234_));
  NAND3_X1   g01042(.A1(new_n1159_), .A2(new_n1233_), .A3(new_n1234_), .ZN(new_n1235_));
  AOI21_X1   g01043(.A1(new_n1232_), .A2(new_n1235_), .B(new_n1063_), .ZN(new_n1236_));
  AND3_X2    g01044(.A1(new_n1159_), .A2(new_n1233_), .A3(new_n1234_), .Z(new_n1237_));
  NOR3_X1    g01045(.A1(new_n1237_), .A2(\a[106] ), .A3(new_n1227_), .ZN(new_n1238_));
  OAI21_X1   g01046(.A1(new_n1222_), .A2(new_n1209_), .B(\asqrt[53] ), .ZN(new_n1239_));
  NAND2_X1   g01047(.A1(new_n1239_), .A2(new_n904_), .ZN(new_n1240_));
  OAI22_X1   g01048(.A1(new_n1230_), .A2(new_n1240_), .B1(new_n1236_), .B2(new_n1238_), .ZN(new_n1241_));
  AOI21_X1   g01049(.A1(new_n1241_), .A2(new_n1231_), .B(new_n823_), .ZN(new_n1242_));
  NOR3_X1    g01050(.A1(new_n1177_), .A2(new_n1062_), .A3(new_n1070_), .ZN(new_n1243_));
  NAND3_X1   g01051(.A1(\asqrt[52] ), .A2(new_n1091_), .A3(new_n1162_), .ZN(new_n1244_));
  AOI22_X1   g01052(.A1(new_n1244_), .A2(new_n1177_), .B1(\asqrt[52] ), .B2(new_n1243_), .ZN(new_n1245_));
  AOI21_X1   g01053(.A1(new_n1159_), .A2(new_n1205_), .B(\a[104] ), .ZN(new_n1246_));
  OAI21_X1   g01054(.A1(new_n1228_), .A2(new_n1246_), .B(new_n1232_), .ZN(new_n1247_));
  OAI21_X1   g01055(.A1(new_n1247_), .A2(new_n1226_), .B(new_n1239_), .ZN(new_n1248_));
  AOI21_X1   g01056(.A1(new_n1248_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1249_));
  AOI21_X1   g01057(.A1(new_n1249_), .A2(new_n1241_), .B(new_n1245_), .ZN(new_n1250_));
  OAI21_X1   g01058(.A1(new_n1250_), .A2(new_n1242_), .B(\asqrt[56] ), .ZN(new_n1251_));
  NOR2_X1    g01059(.A1(new_n1082_), .A2(new_n1083_), .ZN(new_n1252_));
  NOR2_X1    g01060(.A1(new_n1074_), .A2(new_n1085_), .ZN(new_n1253_));
  INV_X1     g01061(.I(new_n1253_), .ZN(new_n1254_));
  NAND4_X1   g01062(.A1(\asqrt[52] ), .A2(new_n1075_), .A3(new_n1252_), .A4(new_n1254_), .ZN(new_n1255_));
  INV_X1     g01063(.I(\asqrt[52] ), .ZN(new_n1256_));
  NOR3_X1    g01064(.A1(new_n1256_), .A2(new_n1166_), .A3(new_n1253_), .ZN(new_n1257_));
  OAI21_X1   g01065(.A1(new_n1257_), .A2(new_n1252_), .B(new_n1255_), .ZN(new_n1258_));
  NAND2_X1   g01066(.A1(new_n1219_), .A2(new_n1224_), .ZN(new_n1259_));
  OAI21_X1   g01067(.A1(new_n1216_), .A2(new_n1218_), .B(new_n1221_), .ZN(new_n1260_));
  NAND2_X1   g01068(.A1(new_n1260_), .A2(\a[105] ), .ZN(new_n1261_));
  NAND3_X1   g01069(.A1(new_n1259_), .A2(new_n1261_), .A3(new_n1232_), .ZN(new_n1262_));
  AOI21_X1   g01070(.A1(new_n1262_), .A2(new_n1239_), .B(new_n904_), .ZN(new_n1263_));
  OAI21_X1   g01071(.A1(new_n1237_), .A2(new_n1227_), .B(\a[106] ), .ZN(new_n1264_));
  NAND3_X1   g01072(.A1(new_n1232_), .A2(new_n1235_), .A3(new_n1063_), .ZN(new_n1265_));
  NAND2_X1   g01073(.A1(new_n1219_), .A2(new_n1210_), .ZN(new_n1266_));
  AOI21_X1   g01074(.A1(new_n1266_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n1267_));
  AOI22_X1   g01075(.A1(new_n1262_), .A2(new_n1267_), .B1(new_n1264_), .B2(new_n1265_), .ZN(new_n1268_));
  OAI21_X1   g01076(.A1(new_n1268_), .A2(new_n1263_), .B(\asqrt[55] ), .ZN(new_n1269_));
  NAND2_X1   g01077(.A1(new_n1269_), .A2(new_n703_), .ZN(new_n1270_));
  OAI21_X1   g01078(.A1(new_n1270_), .A2(new_n1250_), .B(new_n1258_), .ZN(new_n1271_));
  AOI21_X1   g01079(.A1(new_n1271_), .A2(new_n1251_), .B(new_n531_), .ZN(new_n1272_));
  NOR2_X1    g01080(.A1(new_n1179_), .A2(new_n1171_), .ZN(new_n1273_));
  NOR3_X1    g01081(.A1(new_n1256_), .A2(new_n1087_), .A3(new_n1273_), .ZN(new_n1274_));
  INV_X1     g01082(.I(new_n1274_), .ZN(new_n1275_));
  NOR3_X1    g01083(.A1(new_n1273_), .A2(new_n1087_), .A3(new_n1176_), .ZN(new_n1276_));
  AOI22_X1   g01084(.A1(new_n1275_), .A2(new_n1176_), .B1(\asqrt[52] ), .B2(new_n1276_), .ZN(new_n1277_));
  INV_X1     g01085(.I(new_n1245_), .ZN(new_n1278_));
  AOI21_X1   g01086(.A1(\a[105] ), .A2(new_n1260_), .B(new_n1227_), .ZN(new_n1279_));
  AOI21_X1   g01087(.A1(new_n1279_), .A2(new_n1259_), .B(new_n1220_), .ZN(new_n1280_));
  OAI21_X1   g01088(.A1(new_n1280_), .A2(new_n904_), .B(new_n823_), .ZN(new_n1281_));
  OAI21_X1   g01089(.A1(new_n1281_), .A2(new_n1268_), .B(new_n1278_), .ZN(new_n1282_));
  NAND2_X1   g01090(.A1(new_n1282_), .A2(new_n1269_), .ZN(new_n1283_));
  AOI21_X1   g01091(.A1(new_n1283_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1284_));
  AOI21_X1   g01092(.A1(new_n1284_), .A2(new_n1271_), .B(new_n1277_), .ZN(new_n1285_));
  OAI21_X1   g01093(.A1(new_n1285_), .A2(new_n1272_), .B(\asqrt[58] ), .ZN(new_n1286_));
  NOR3_X1    g01094(.A1(new_n1098_), .A2(new_n1107_), .A3(new_n1105_), .ZN(new_n1287_));
  NOR3_X1    g01095(.A1(new_n1256_), .A2(new_n1098_), .A3(new_n1107_), .ZN(new_n1288_));
  INV_X1     g01096(.I(new_n1288_), .ZN(new_n1289_));
  AOI22_X1   g01097(.A1(new_n1289_), .A2(new_n1105_), .B1(\asqrt[52] ), .B2(new_n1287_), .ZN(new_n1290_));
  INV_X1     g01098(.I(new_n1290_), .ZN(new_n1291_));
  AOI21_X1   g01099(.A1(new_n1282_), .A2(new_n1269_), .B(new_n703_), .ZN(new_n1292_));
  INV_X1     g01100(.I(new_n1258_), .ZN(new_n1293_));
  NOR2_X1    g01101(.A1(new_n1242_), .A2(\asqrt[56] ), .ZN(new_n1294_));
  AOI21_X1   g01102(.A1(new_n1294_), .A2(new_n1282_), .B(new_n1293_), .ZN(new_n1295_));
  OAI21_X1   g01103(.A1(new_n1295_), .A2(new_n1292_), .B(\asqrt[57] ), .ZN(new_n1296_));
  NAND2_X1   g01104(.A1(new_n1296_), .A2(new_n436_), .ZN(new_n1297_));
  OAI21_X1   g01105(.A1(new_n1297_), .A2(new_n1285_), .B(new_n1291_), .ZN(new_n1298_));
  AOI21_X1   g01106(.A1(new_n1298_), .A2(new_n1286_), .B(new_n327_), .ZN(new_n1299_));
  NOR2_X1    g01107(.A1(new_n1108_), .A2(new_n1116_), .ZN(new_n1300_));
  NOR3_X1    g01108(.A1(new_n1256_), .A2(new_n1175_), .A3(new_n1300_), .ZN(new_n1301_));
  INV_X1     g01109(.I(new_n1301_), .ZN(new_n1302_));
  NOR3_X1    g01110(.A1(new_n1300_), .A2(new_n1175_), .A3(new_n1115_), .ZN(new_n1303_));
  AOI22_X1   g01111(.A1(new_n1302_), .A2(new_n1115_), .B1(\asqrt[52] ), .B2(new_n1303_), .ZN(new_n1304_));
  INV_X1     g01112(.I(new_n1277_), .ZN(new_n1305_));
  NAND2_X1   g01113(.A1(new_n1251_), .A2(new_n531_), .ZN(new_n1306_));
  OAI21_X1   g01114(.A1(new_n1306_), .A2(new_n1295_), .B(new_n1305_), .ZN(new_n1307_));
  AOI21_X1   g01115(.A1(new_n1307_), .A2(new_n1296_), .B(new_n436_), .ZN(new_n1308_));
  NOR2_X1    g01116(.A1(new_n1308_), .A2(\asqrt[59] ), .ZN(new_n1309_));
  AOI21_X1   g01117(.A1(new_n1309_), .A2(new_n1298_), .B(new_n1304_), .ZN(new_n1310_));
  OAI21_X1   g01118(.A1(new_n1310_), .A2(new_n1299_), .B(\asqrt[60] ), .ZN(new_n1311_));
  INV_X1     g01119(.I(new_n1122_), .ZN(new_n1312_));
  NOR3_X1    g01120(.A1(new_n1118_), .A2(new_n1187_), .A3(new_n1312_), .ZN(new_n1313_));
  NOR3_X1    g01121(.A1(new_n1256_), .A2(new_n1118_), .A3(new_n1187_), .ZN(new_n1314_));
  INV_X1     g01122(.I(new_n1314_), .ZN(new_n1315_));
  AOI22_X1   g01123(.A1(new_n1315_), .A2(new_n1312_), .B1(\asqrt[52] ), .B2(new_n1313_), .ZN(new_n1316_));
  INV_X1     g01124(.I(new_n1316_), .ZN(new_n1317_));
  NOR3_X1    g01125(.A1(new_n1250_), .A2(new_n1242_), .A3(\asqrt[56] ), .ZN(new_n1318_));
  OAI21_X1   g01126(.A1(new_n1293_), .A2(new_n1318_), .B(new_n1251_), .ZN(new_n1319_));
  AOI21_X1   g01127(.A1(new_n1319_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n1320_));
  AOI21_X1   g01128(.A1(new_n1320_), .A2(new_n1307_), .B(new_n1290_), .ZN(new_n1321_));
  OAI21_X1   g01129(.A1(new_n1321_), .A2(new_n1308_), .B(\asqrt[59] ), .ZN(new_n1322_));
  INV_X1     g01130(.I(new_n1304_), .ZN(new_n1323_));
  NAND2_X1   g01131(.A1(new_n1286_), .A2(new_n327_), .ZN(new_n1324_));
  OAI21_X1   g01132(.A1(new_n1324_), .A2(new_n1321_), .B(new_n1323_), .ZN(new_n1325_));
  NAND3_X1   g01133(.A1(new_n1325_), .A2(new_n306_), .A3(new_n1322_), .ZN(new_n1326_));
  NAND2_X1   g01134(.A1(new_n1326_), .A2(new_n1317_), .ZN(new_n1327_));
  AOI21_X1   g01135(.A1(new_n1327_), .A2(new_n1311_), .B(new_n218_), .ZN(new_n1328_));
  NOR3_X1    g01136(.A1(new_n1256_), .A2(new_n1127_), .A3(new_n1133_), .ZN(new_n1329_));
  INV_X1     g01137(.I(new_n1329_), .ZN(new_n1330_));
  NOR3_X1    g01138(.A1(new_n1127_), .A2(new_n1160_), .A3(new_n1133_), .ZN(new_n1331_));
  AOI22_X1   g01139(.A1(new_n1330_), .A2(new_n1160_), .B1(\asqrt[52] ), .B2(new_n1331_), .ZN(new_n1332_));
  AOI21_X1   g01140(.A1(new_n1325_), .A2(new_n1322_), .B(new_n306_), .ZN(new_n1333_));
  NOR2_X1    g01141(.A1(new_n1333_), .A2(\asqrt[61] ), .ZN(new_n1334_));
  AOI21_X1   g01142(.A1(new_n1334_), .A2(new_n1327_), .B(new_n1332_), .ZN(new_n1335_));
  OAI21_X1   g01143(.A1(new_n1335_), .A2(new_n1328_), .B(\asqrt[62] ), .ZN(new_n1336_));
  INV_X1     g01144(.I(new_n1211_), .ZN(new_n1337_));
  NOR3_X1    g01145(.A1(new_n1337_), .A2(new_n1213_), .A3(new_n1141_), .ZN(new_n1338_));
  NOR3_X1    g01146(.A1(new_n1256_), .A2(new_n1213_), .A3(new_n1337_), .ZN(new_n1339_));
  INV_X1     g01147(.I(new_n1339_), .ZN(new_n1340_));
  AOI22_X1   g01148(.A1(new_n1340_), .A2(new_n1141_), .B1(\asqrt[52] ), .B2(new_n1338_), .ZN(new_n1341_));
  INV_X1     g01149(.I(new_n1341_), .ZN(new_n1342_));
  NOR3_X1    g01150(.A1(new_n1285_), .A2(new_n1272_), .A3(\asqrt[58] ), .ZN(new_n1343_));
  OAI21_X1   g01151(.A1(new_n1290_), .A2(new_n1343_), .B(new_n1286_), .ZN(new_n1344_));
  AOI21_X1   g01152(.A1(new_n1344_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n1345_));
  AOI21_X1   g01153(.A1(new_n1345_), .A2(new_n1325_), .B(new_n1316_), .ZN(new_n1346_));
  OAI21_X1   g01154(.A1(new_n1346_), .A2(new_n1333_), .B(\asqrt[61] ), .ZN(new_n1347_));
  NAND2_X1   g01155(.A1(new_n1347_), .A2(new_n207_), .ZN(new_n1348_));
  OAI21_X1   g01156(.A1(new_n1348_), .A2(new_n1335_), .B(new_n1342_), .ZN(new_n1349_));
  INV_X1     g01157(.I(new_n1144_), .ZN(new_n1350_));
  INV_X1     g01158(.I(new_n1214_), .ZN(new_n1351_));
  NAND4_X1   g01159(.A1(\asqrt[52] ), .A2(new_n1350_), .A3(new_n1148_), .A4(new_n1351_), .ZN(new_n1352_));
  NAND2_X1   g01160(.A1(new_n1350_), .A2(new_n1351_), .ZN(new_n1353_));
  OAI21_X1   g01161(.A1(new_n1256_), .A2(new_n1353_), .B(new_n1191_), .ZN(new_n1354_));
  NAND2_X1   g01162(.A1(new_n1354_), .A2(new_n1352_), .ZN(new_n1355_));
  INV_X1     g01163(.I(new_n1233_), .ZN(new_n1356_));
  AOI21_X1   g01164(.A1(new_n1350_), .A2(new_n1193_), .B(new_n1155_), .ZN(new_n1357_));
  AOI21_X1   g01165(.A1(\asqrt[52] ), .A2(new_n1357_), .B(new_n1356_), .ZN(new_n1358_));
  NAND2_X1   g01166(.A1(new_n1355_), .A2(new_n1358_), .ZN(new_n1359_));
  AOI21_X1   g01167(.A1(new_n1349_), .A2(new_n1336_), .B(new_n1359_), .ZN(new_n1360_));
  NOR3_X1    g01168(.A1(new_n1321_), .A2(\asqrt[59] ), .A3(new_n1308_), .ZN(new_n1361_));
  OAI21_X1   g01169(.A1(new_n1304_), .A2(new_n1361_), .B(new_n1322_), .ZN(new_n1362_));
  AOI22_X1   g01170(.A1(new_n1326_), .A2(new_n1317_), .B1(new_n1362_), .B2(\asqrt[60] ), .ZN(new_n1363_));
  NOR3_X1    g01171(.A1(new_n1346_), .A2(\asqrt[61] ), .A3(new_n1333_), .ZN(new_n1364_));
  OAI22_X1   g01172(.A1(new_n1364_), .A2(new_n1332_), .B1(new_n1363_), .B2(new_n218_), .ZN(new_n1365_));
  AOI21_X1   g01173(.A1(new_n1365_), .A2(\asqrt[62] ), .B(new_n1355_), .ZN(new_n1366_));
  AOI21_X1   g01174(.A1(\asqrt[52] ), .A2(new_n1194_), .B(new_n1215_), .ZN(new_n1367_));
  OR3_X2     g01175(.A1(new_n1367_), .A2(new_n193_), .A3(new_n1357_), .Z(new_n1368_));
  NAND2_X1   g01176(.A1(\asqrt[53] ), .A2(new_n1152_), .ZN(new_n1369_));
  NAND2_X1   g01177(.A1(new_n1369_), .A2(new_n1201_), .ZN(new_n1370_));
  NOR4_X1    g01178(.A1(new_n1356_), .A2(new_n1154_), .A3(new_n1198_), .A4(new_n1370_), .ZN(new_n1371_));
  NAND2_X1   g01179(.A1(new_n1371_), .A2(new_n1159_), .ZN(new_n1372_));
  NAND2_X1   g01180(.A1(new_n1368_), .A2(new_n1372_), .ZN(new_n1373_));
  AOI21_X1   g01181(.A1(new_n1366_), .A2(new_n1349_), .B(new_n1373_), .ZN(new_n1374_));
  OAI21_X1   g01182(.A1(\asqrt[63] ), .A2(new_n1360_), .B(new_n1374_), .ZN(\asqrt[51] ));
  INV_X1     g01183(.I(\asqrt[51] ), .ZN(new_n1376_));
  NOR2_X1    g01184(.A1(\a[100] ), .A2(\a[101] ), .ZN(new_n1377_));
  INV_X1     g01185(.I(new_n1377_), .ZN(new_n1378_));
  NOR2_X1    g01186(.A1(new_n1378_), .A2(\a[102] ), .ZN(new_n1379_));
  INV_X1     g01187(.I(new_n1379_), .ZN(new_n1380_));
  NOR2_X1    g01188(.A1(new_n1360_), .A2(\asqrt[63] ), .ZN(new_n1381_));
  INV_X1     g01189(.I(new_n1349_), .ZN(new_n1382_));
  INV_X1     g01190(.I(new_n1355_), .ZN(new_n1383_));
  NAND2_X1   g01191(.A1(new_n1336_), .A2(new_n1383_), .ZN(new_n1384_));
  INV_X1     g01192(.I(new_n1373_), .ZN(new_n1385_));
  OAI21_X1   g01193(.A1(new_n1382_), .A2(new_n1384_), .B(new_n1385_), .ZN(new_n1386_));
  OAI21_X1   g01194(.A1(new_n1381_), .A2(new_n1386_), .B(\a[102] ), .ZN(new_n1387_));
  AOI21_X1   g01195(.A1(new_n1387_), .A2(new_n1380_), .B(new_n1256_), .ZN(new_n1388_));
  INV_X1     g01196(.I(\a[102] ), .ZN(new_n1389_));
  INV_X1     g01197(.I(new_n1332_), .ZN(new_n1390_));
  NAND2_X1   g01198(.A1(new_n1311_), .A2(new_n218_), .ZN(new_n1391_));
  OAI21_X1   g01199(.A1(new_n1391_), .A2(new_n1346_), .B(new_n1390_), .ZN(new_n1392_));
  NAND3_X1   g01200(.A1(new_n1392_), .A2(new_n207_), .A3(new_n1347_), .ZN(new_n1393_));
  AOI22_X1   g01201(.A1(new_n1393_), .A2(new_n1342_), .B1(new_n1365_), .B2(\asqrt[62] ), .ZN(new_n1394_));
  OAI21_X1   g01202(.A1(new_n1394_), .A2(new_n1359_), .B(new_n193_), .ZN(new_n1395_));
  AOI21_X1   g01203(.A1(new_n1395_), .A2(new_n1374_), .B(new_n1389_), .ZN(new_n1396_));
  NOR3_X1    g01204(.A1(new_n1198_), .A2(new_n1202_), .A3(new_n1379_), .ZN(new_n1397_));
  NAND3_X1   g01205(.A1(new_n1159_), .A2(new_n1233_), .A3(new_n1397_), .ZN(new_n1398_));
  NOR2_X1    g01206(.A1(new_n1396_), .A2(new_n1398_), .ZN(new_n1399_));
  AOI21_X1   g01207(.A1(new_n1395_), .A2(new_n1374_), .B(new_n1208_), .ZN(new_n1400_));
  INV_X1     g01208(.I(\a[103] ), .ZN(new_n1401_));
  AOI21_X1   g01209(.A1(\asqrt[51] ), .A2(new_n1389_), .B(new_n1401_), .ZN(new_n1402_));
  NOR3_X1    g01210(.A1(new_n1399_), .A2(new_n1402_), .A3(new_n1400_), .ZN(new_n1403_));
  OAI21_X1   g01211(.A1(new_n1403_), .A2(new_n1388_), .B(\asqrt[53] ), .ZN(new_n1404_));
  OAI21_X1   g01212(.A1(new_n1381_), .A2(new_n1386_), .B(new_n1207_), .ZN(new_n1405_));
  NOR2_X1    g01213(.A1(new_n1382_), .A2(new_n1384_), .ZN(new_n1406_));
  INV_X1     g01214(.I(new_n1406_), .ZN(new_n1407_));
  OAI21_X1   g01215(.A1(new_n1371_), .A2(new_n1205_), .B(new_n1159_), .ZN(new_n1408_));
  NAND4_X1   g01216(.A1(new_n1407_), .A2(new_n1395_), .A3(new_n1368_), .A4(new_n1408_), .ZN(new_n1409_));
  AOI21_X1   g01217(.A1(new_n1409_), .A2(new_n1405_), .B(new_n1221_), .ZN(new_n1410_));
  NAND2_X1   g01218(.A1(new_n1368_), .A2(new_n1408_), .ZN(new_n1411_));
  NOR3_X1    g01219(.A1(new_n1381_), .A2(new_n1406_), .A3(new_n1411_), .ZN(new_n1412_));
  NOR3_X1    g01220(.A1(new_n1412_), .A2(new_n1400_), .A3(\a[104] ), .ZN(new_n1413_));
  AOI21_X1   g01221(.A1(\asqrt[51] ), .A2(\a[102] ), .B(new_n1379_), .ZN(new_n1414_));
  OAI21_X1   g01222(.A1(new_n1414_), .A2(new_n1256_), .B(new_n1103_), .ZN(new_n1415_));
  OAI22_X1   g01223(.A1(new_n1403_), .A2(new_n1415_), .B1(new_n1410_), .B2(new_n1413_), .ZN(new_n1416_));
  AOI21_X1   g01224(.A1(new_n1416_), .A2(new_n1404_), .B(new_n904_), .ZN(new_n1417_));
  NOR3_X1    g01225(.A1(new_n1279_), .A2(new_n1220_), .A3(new_n1226_), .ZN(new_n1418_));
  NAND3_X1   g01226(.A1(\asqrt[51] ), .A2(new_n1239_), .A3(new_n1259_), .ZN(new_n1419_));
  AOI22_X1   g01227(.A1(new_n1419_), .A2(new_n1279_), .B1(\asqrt[51] ), .B2(new_n1418_), .ZN(new_n1420_));
  OAI21_X1   g01228(.A1(new_n1396_), .A2(new_n1379_), .B(\asqrt[52] ), .ZN(new_n1421_));
  AOI21_X1   g01229(.A1(new_n1395_), .A2(new_n1374_), .B(\a[102] ), .ZN(new_n1422_));
  OAI21_X1   g01230(.A1(new_n1401_), .A2(new_n1422_), .B(new_n1405_), .ZN(new_n1423_));
  OAI21_X1   g01231(.A1(new_n1423_), .A2(new_n1399_), .B(new_n1421_), .ZN(new_n1424_));
  AOI21_X1   g01232(.A1(new_n1424_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n1425_));
  AOI21_X1   g01233(.A1(new_n1425_), .A2(new_n1416_), .B(new_n1420_), .ZN(new_n1426_));
  OAI21_X1   g01234(.A1(new_n1426_), .A2(new_n1417_), .B(\asqrt[55] ), .ZN(new_n1427_));
  NOR2_X1    g01235(.A1(new_n1238_), .A2(new_n1236_), .ZN(new_n1428_));
  INV_X1     g01236(.I(new_n1428_), .ZN(new_n1429_));
  NAND2_X1   g01237(.A1(new_n1262_), .A2(new_n1267_), .ZN(new_n1430_));
  AND3_X2    g01238(.A1(new_n1231_), .A2(new_n1428_), .A3(new_n1430_), .Z(new_n1431_));
  NAND3_X1   g01239(.A1(\asqrt[51] ), .A2(new_n1231_), .A3(new_n1430_), .ZN(new_n1432_));
  AOI22_X1   g01240(.A1(new_n1432_), .A2(new_n1429_), .B1(\asqrt[51] ), .B2(new_n1431_), .ZN(new_n1433_));
  INV_X1     g01241(.I(new_n1433_), .ZN(new_n1434_));
  INV_X1     g01242(.I(new_n1398_), .ZN(new_n1435_));
  NAND2_X1   g01243(.A1(new_n1387_), .A2(new_n1435_), .ZN(new_n1436_));
  OAI21_X1   g01244(.A1(new_n1381_), .A2(new_n1386_), .B(new_n1389_), .ZN(new_n1437_));
  AOI21_X1   g01245(.A1(\a[103] ), .A2(new_n1437_), .B(new_n1400_), .ZN(new_n1438_));
  AOI21_X1   g01246(.A1(new_n1438_), .A2(new_n1436_), .B(new_n1388_), .ZN(new_n1439_));
  NOR2_X1    g01247(.A1(new_n1439_), .A2(new_n1103_), .ZN(new_n1440_));
  NAND2_X1   g01248(.A1(new_n1438_), .A2(new_n1436_), .ZN(new_n1441_));
  OAI21_X1   g01249(.A1(new_n1412_), .A2(new_n1400_), .B(\a[104] ), .ZN(new_n1442_));
  NAND3_X1   g01250(.A1(new_n1409_), .A2(new_n1405_), .A3(new_n1221_), .ZN(new_n1443_));
  NOR2_X1    g01251(.A1(new_n1388_), .A2(\asqrt[53] ), .ZN(new_n1444_));
  AOI22_X1   g01252(.A1(new_n1441_), .A2(new_n1444_), .B1(new_n1442_), .B2(new_n1443_), .ZN(new_n1445_));
  OAI21_X1   g01253(.A1(new_n1445_), .A2(new_n1440_), .B(\asqrt[54] ), .ZN(new_n1446_));
  NAND2_X1   g01254(.A1(new_n1446_), .A2(new_n823_), .ZN(new_n1447_));
  OAI21_X1   g01255(.A1(new_n1447_), .A2(new_n1426_), .B(new_n1434_), .ZN(new_n1448_));
  AOI21_X1   g01256(.A1(new_n1448_), .A2(new_n1427_), .B(new_n703_), .ZN(new_n1449_));
  NOR2_X1    g01257(.A1(new_n1281_), .A2(new_n1268_), .ZN(new_n1450_));
  NOR3_X1    g01258(.A1(new_n1376_), .A2(new_n1242_), .A3(new_n1450_), .ZN(new_n1451_));
  INV_X1     g01259(.I(new_n1451_), .ZN(new_n1452_));
  NOR3_X1    g01260(.A1(new_n1450_), .A2(new_n1242_), .A3(new_n1278_), .ZN(new_n1453_));
  AOI22_X1   g01261(.A1(new_n1452_), .A2(new_n1278_), .B1(\asqrt[51] ), .B2(new_n1453_), .ZN(new_n1454_));
  INV_X1     g01262(.I(new_n1420_), .ZN(new_n1455_));
  OAI21_X1   g01263(.A1(new_n1439_), .A2(new_n1103_), .B(new_n904_), .ZN(new_n1456_));
  OAI21_X1   g01264(.A1(new_n1456_), .A2(new_n1445_), .B(new_n1455_), .ZN(new_n1457_));
  AOI21_X1   g01265(.A1(new_n1457_), .A2(new_n1446_), .B(new_n823_), .ZN(new_n1458_));
  NOR2_X1    g01266(.A1(new_n1458_), .A2(\asqrt[56] ), .ZN(new_n1459_));
  AOI21_X1   g01267(.A1(new_n1459_), .A2(new_n1448_), .B(new_n1454_), .ZN(new_n1460_));
  OAI21_X1   g01268(.A1(new_n1460_), .A2(new_n1449_), .B(\asqrt[57] ), .ZN(new_n1461_));
  NOR3_X1    g01269(.A1(new_n1292_), .A2(new_n1318_), .A3(new_n1258_), .ZN(new_n1462_));
  NOR3_X1    g01270(.A1(new_n1376_), .A2(new_n1292_), .A3(new_n1318_), .ZN(new_n1463_));
  INV_X1     g01271(.I(new_n1463_), .ZN(new_n1464_));
  AOI22_X1   g01272(.A1(new_n1464_), .A2(new_n1258_), .B1(\asqrt[51] ), .B2(new_n1462_), .ZN(new_n1465_));
  INV_X1     g01273(.I(new_n1465_), .ZN(new_n1466_));
  NOR3_X1    g01274(.A1(new_n1426_), .A2(new_n1417_), .A3(\asqrt[55] ), .ZN(new_n1467_));
  NOR2_X1    g01275(.A1(new_n1467_), .A2(new_n1433_), .ZN(new_n1468_));
  OAI21_X1   g01276(.A1(new_n1468_), .A2(new_n1458_), .B(\asqrt[56] ), .ZN(new_n1469_));
  NAND2_X1   g01277(.A1(new_n1469_), .A2(new_n531_), .ZN(new_n1470_));
  OAI21_X1   g01278(.A1(new_n1470_), .A2(new_n1460_), .B(new_n1466_), .ZN(new_n1471_));
  AOI21_X1   g01279(.A1(new_n1471_), .A2(new_n1461_), .B(new_n436_), .ZN(new_n1472_));
  NOR2_X1    g01280(.A1(new_n1306_), .A2(new_n1295_), .ZN(new_n1473_));
  NOR3_X1    g01281(.A1(new_n1376_), .A2(new_n1272_), .A3(new_n1473_), .ZN(new_n1474_));
  INV_X1     g01282(.I(new_n1474_), .ZN(new_n1475_));
  NOR3_X1    g01283(.A1(new_n1272_), .A2(new_n1473_), .A3(new_n1305_), .ZN(new_n1476_));
  AOI22_X1   g01284(.A1(new_n1475_), .A2(new_n1305_), .B1(\asqrt[51] ), .B2(new_n1476_), .ZN(new_n1477_));
  INV_X1     g01285(.I(new_n1454_), .ZN(new_n1478_));
  NAND2_X1   g01286(.A1(new_n1427_), .A2(new_n703_), .ZN(new_n1479_));
  OAI21_X1   g01287(.A1(new_n1468_), .A2(new_n1479_), .B(new_n1478_), .ZN(new_n1480_));
  AOI21_X1   g01288(.A1(new_n1480_), .A2(new_n1469_), .B(new_n531_), .ZN(new_n1481_));
  NOR2_X1    g01289(.A1(new_n1481_), .A2(\asqrt[58] ), .ZN(new_n1482_));
  AOI21_X1   g01290(.A1(new_n1482_), .A2(new_n1471_), .B(new_n1477_), .ZN(new_n1483_));
  OAI21_X1   g01291(.A1(new_n1483_), .A2(new_n1472_), .B(\asqrt[59] ), .ZN(new_n1484_));
  INV_X1     g01292(.I(new_n1484_), .ZN(new_n1485_));
  OAI21_X1   g01293(.A1(new_n1433_), .A2(new_n1467_), .B(new_n1427_), .ZN(new_n1486_));
  AOI21_X1   g01294(.A1(new_n1486_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1487_));
  AOI21_X1   g01295(.A1(new_n1487_), .A2(new_n1480_), .B(new_n1465_), .ZN(new_n1488_));
  INV_X1     g01296(.I(new_n1477_), .ZN(new_n1489_));
  NAND2_X1   g01297(.A1(new_n1461_), .A2(new_n436_), .ZN(new_n1490_));
  OAI21_X1   g01298(.A1(new_n1490_), .A2(new_n1488_), .B(new_n1489_), .ZN(new_n1491_));
  NOR3_X1    g01299(.A1(new_n1343_), .A2(new_n1308_), .A3(new_n1291_), .ZN(new_n1492_));
  NOR3_X1    g01300(.A1(new_n1376_), .A2(new_n1308_), .A3(new_n1343_), .ZN(new_n1493_));
  INV_X1     g01301(.I(new_n1493_), .ZN(new_n1494_));
  AOI22_X1   g01302(.A1(new_n1494_), .A2(new_n1291_), .B1(\asqrt[51] ), .B2(new_n1492_), .ZN(new_n1495_));
  NOR2_X1    g01303(.A1(new_n1472_), .A2(\asqrt[59] ), .ZN(new_n1496_));
  AOI21_X1   g01304(.A1(new_n1496_), .A2(new_n1491_), .B(new_n1495_), .ZN(new_n1497_));
  OAI21_X1   g01305(.A1(new_n1485_), .A2(new_n1497_), .B(\asqrt[60] ), .ZN(new_n1498_));
  NOR3_X1    g01306(.A1(new_n1376_), .A2(new_n1299_), .A3(new_n1361_), .ZN(new_n1499_));
  INV_X1     g01307(.I(new_n1499_), .ZN(new_n1500_));
  NOR3_X1    g01308(.A1(new_n1299_), .A2(new_n1323_), .A3(new_n1361_), .ZN(new_n1501_));
  AOI22_X1   g01309(.A1(new_n1500_), .A2(new_n1323_), .B1(\asqrt[51] ), .B2(new_n1501_), .ZN(new_n1502_));
  INV_X1     g01310(.I(new_n1502_), .ZN(new_n1503_));
  NAND2_X1   g01311(.A1(new_n1484_), .A2(new_n306_), .ZN(new_n1504_));
  OAI21_X1   g01312(.A1(new_n1504_), .A2(new_n1497_), .B(new_n1503_), .ZN(new_n1505_));
  AOI21_X1   g01313(.A1(new_n1505_), .A2(new_n1498_), .B(new_n218_), .ZN(new_n1506_));
  AND3_X2    g01314(.A1(new_n1311_), .A2(new_n1326_), .A3(new_n1316_), .Z(new_n1507_));
  NAND3_X1   g01315(.A1(\asqrt[51] ), .A2(new_n1311_), .A3(new_n1326_), .ZN(new_n1508_));
  AOI22_X1   g01316(.A1(new_n1508_), .A2(new_n1317_), .B1(\asqrt[51] ), .B2(new_n1507_), .ZN(new_n1509_));
  INV_X1     g01317(.I(new_n1495_), .ZN(new_n1510_));
  OAI21_X1   g01318(.A1(new_n1488_), .A2(new_n1481_), .B(\asqrt[58] ), .ZN(new_n1511_));
  NAND2_X1   g01319(.A1(new_n1511_), .A2(new_n327_), .ZN(new_n1512_));
  OAI21_X1   g01320(.A1(new_n1512_), .A2(new_n1483_), .B(new_n1510_), .ZN(new_n1513_));
  AOI21_X1   g01321(.A1(new_n1513_), .A2(new_n1484_), .B(new_n306_), .ZN(new_n1514_));
  NOR2_X1    g01322(.A1(new_n1514_), .A2(\asqrt[61] ), .ZN(new_n1515_));
  AOI21_X1   g01323(.A1(new_n1515_), .A2(new_n1505_), .B(new_n1509_), .ZN(new_n1516_));
  OAI21_X1   g01324(.A1(new_n1516_), .A2(new_n1506_), .B(\asqrt[62] ), .ZN(new_n1517_));
  NOR3_X1    g01325(.A1(new_n1376_), .A2(new_n1328_), .A3(new_n1364_), .ZN(new_n1518_));
  INV_X1     g01326(.I(new_n1518_), .ZN(new_n1519_));
  NOR3_X1    g01327(.A1(new_n1328_), .A2(new_n1390_), .A3(new_n1364_), .ZN(new_n1520_));
  AOI22_X1   g01328(.A1(new_n1519_), .A2(new_n1390_), .B1(\asqrt[51] ), .B2(new_n1520_), .ZN(new_n1521_));
  INV_X1     g01329(.I(new_n1521_), .ZN(new_n1522_));
  NOR3_X1    g01330(.A1(new_n1488_), .A2(new_n1481_), .A3(\asqrt[58] ), .ZN(new_n1523_));
  OAI21_X1   g01331(.A1(new_n1477_), .A2(new_n1523_), .B(new_n1511_), .ZN(new_n1524_));
  AOI21_X1   g01332(.A1(new_n1524_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n1525_));
  AOI21_X1   g01333(.A1(new_n1525_), .A2(new_n1513_), .B(new_n1502_), .ZN(new_n1526_));
  OAI21_X1   g01334(.A1(new_n1526_), .A2(new_n1514_), .B(\asqrt[61] ), .ZN(new_n1527_));
  NAND2_X1   g01335(.A1(new_n1527_), .A2(new_n207_), .ZN(new_n1528_));
  OAI21_X1   g01336(.A1(new_n1528_), .A2(new_n1516_), .B(new_n1522_), .ZN(new_n1529_));
  NAND4_X1   g01337(.A1(\asqrt[51] ), .A2(new_n1336_), .A3(new_n1341_), .A4(new_n1393_), .ZN(new_n1530_));
  NAND2_X1   g01338(.A1(new_n1336_), .A2(new_n1393_), .ZN(new_n1531_));
  OAI21_X1   g01339(.A1(new_n1376_), .A2(new_n1531_), .B(new_n1342_), .ZN(new_n1532_));
  NAND2_X1   g01340(.A1(new_n1532_), .A2(new_n1530_), .ZN(new_n1533_));
  NOR2_X1    g01341(.A1(new_n1394_), .A2(new_n1383_), .ZN(new_n1534_));
  NAND2_X1   g01342(.A1(\asqrt[51] ), .A2(new_n1534_), .ZN(new_n1535_));
  NAND3_X1   g01343(.A1(new_n1533_), .A2(new_n1407_), .A3(new_n1535_), .ZN(new_n1536_));
  AOI21_X1   g01344(.A1(new_n1529_), .A2(new_n1517_), .B(new_n1536_), .ZN(new_n1537_));
  NOR3_X1    g01345(.A1(new_n1526_), .A2(\asqrt[61] ), .A3(new_n1514_), .ZN(new_n1538_));
  OAI21_X1   g01346(.A1(new_n1509_), .A2(new_n1538_), .B(new_n1527_), .ZN(new_n1539_));
  AOI21_X1   g01347(.A1(new_n1539_), .A2(\asqrt[62] ), .B(new_n1533_), .ZN(new_n1540_));
  OAI21_X1   g01348(.A1(new_n1376_), .A2(new_n1383_), .B(new_n1394_), .ZN(new_n1541_));
  NOR2_X1    g01349(.A1(new_n1534_), .A2(new_n193_), .ZN(new_n1542_));
  NAND2_X1   g01350(.A1(new_n1541_), .A2(new_n1542_), .ZN(new_n1543_));
  INV_X1     g01351(.I(new_n1543_), .ZN(new_n1544_));
  AND3_X2    g01352(.A1(new_n1354_), .A2(new_n1352_), .A3(new_n1372_), .Z(new_n1545_));
  NAND4_X1   g01353(.A1(new_n1407_), .A2(new_n1395_), .A3(new_n1368_), .A4(new_n1545_), .ZN(new_n1546_));
  INV_X1     g01354(.I(new_n1546_), .ZN(new_n1547_));
  NOR2_X1    g01355(.A1(new_n1544_), .A2(new_n1547_), .ZN(new_n1548_));
  INV_X1     g01356(.I(new_n1548_), .ZN(new_n1549_));
  AOI21_X1   g01357(.A1(new_n1540_), .A2(new_n1529_), .B(new_n1549_), .ZN(new_n1550_));
  OAI21_X1   g01358(.A1(\asqrt[63] ), .A2(new_n1537_), .B(new_n1550_), .ZN(\asqrt[50] ));
  NOR2_X1    g01359(.A1(\a[98] ), .A2(\a[99] ), .ZN(new_n1552_));
  INV_X1     g01360(.I(new_n1552_), .ZN(new_n1553_));
  NOR2_X1    g01361(.A1(new_n1553_), .A2(\a[100] ), .ZN(new_n1554_));
  INV_X1     g01362(.I(new_n1554_), .ZN(new_n1555_));
  NAND2_X1   g01363(.A1(new_n1529_), .A2(new_n1517_), .ZN(new_n1556_));
  INV_X1     g01364(.I(new_n1536_), .ZN(new_n1557_));
  AOI21_X1   g01365(.A1(new_n1556_), .A2(new_n1557_), .B(\asqrt[63] ), .ZN(new_n1558_));
  INV_X1     g01366(.I(new_n1529_), .ZN(new_n1559_));
  INV_X1     g01367(.I(new_n1533_), .ZN(new_n1560_));
  NAND2_X1   g01368(.A1(new_n1517_), .A2(new_n1560_), .ZN(new_n1561_));
  OAI21_X1   g01369(.A1(new_n1559_), .A2(new_n1561_), .B(new_n1548_), .ZN(new_n1562_));
  OAI21_X1   g01370(.A1(new_n1558_), .A2(new_n1562_), .B(\a[100] ), .ZN(new_n1563_));
  AOI21_X1   g01371(.A1(new_n1563_), .A2(new_n1555_), .B(new_n1376_), .ZN(new_n1564_));
  INV_X1     g01372(.I(\a[100] ), .ZN(new_n1565_));
  INV_X1     g01373(.I(new_n1509_), .ZN(new_n1566_));
  NAND3_X1   g01374(.A1(new_n1491_), .A2(new_n327_), .A3(new_n1511_), .ZN(new_n1567_));
  AOI22_X1   g01375(.A1(new_n1567_), .A2(new_n1510_), .B1(new_n1524_), .B2(\asqrt[59] ), .ZN(new_n1568_));
  OAI21_X1   g01376(.A1(new_n1568_), .A2(new_n306_), .B(new_n218_), .ZN(new_n1569_));
  OAI21_X1   g01377(.A1(new_n1569_), .A2(new_n1526_), .B(new_n1566_), .ZN(new_n1570_));
  NAND3_X1   g01378(.A1(new_n1570_), .A2(new_n207_), .A3(new_n1527_), .ZN(new_n1571_));
  AOI22_X1   g01379(.A1(new_n1571_), .A2(new_n1522_), .B1(new_n1539_), .B2(\asqrt[62] ), .ZN(new_n1572_));
  OAI21_X1   g01380(.A1(new_n1572_), .A2(new_n1536_), .B(new_n193_), .ZN(new_n1573_));
  AOI21_X1   g01381(.A1(new_n1573_), .A2(new_n1550_), .B(new_n1565_), .ZN(new_n1574_));
  NAND4_X1   g01382(.A1(new_n1407_), .A2(new_n1368_), .A3(new_n1372_), .A4(new_n1555_), .ZN(new_n1575_));
  NOR2_X1    g01383(.A1(new_n1575_), .A2(new_n1381_), .ZN(new_n1576_));
  INV_X1     g01384(.I(new_n1576_), .ZN(new_n1577_));
  NOR2_X1    g01385(.A1(new_n1574_), .A2(new_n1577_), .ZN(new_n1578_));
  AOI21_X1   g01386(.A1(new_n1573_), .A2(new_n1550_), .B(new_n1378_), .ZN(new_n1579_));
  INV_X1     g01387(.I(\a[101] ), .ZN(new_n1580_));
  AOI21_X1   g01388(.A1(\asqrt[50] ), .A2(new_n1565_), .B(new_n1580_), .ZN(new_n1581_));
  NOR3_X1    g01389(.A1(new_n1578_), .A2(new_n1581_), .A3(new_n1579_), .ZN(new_n1582_));
  OAI21_X1   g01390(.A1(new_n1582_), .A2(new_n1564_), .B(\asqrt[52] ), .ZN(new_n1583_));
  OAI21_X1   g01391(.A1(new_n1558_), .A2(new_n1562_), .B(new_n1377_), .ZN(new_n1584_));
  NOR2_X1    g01392(.A1(new_n1559_), .A2(new_n1561_), .ZN(new_n1585_));
  INV_X1     g01393(.I(new_n1585_), .ZN(new_n1586_));
  NOR2_X1    g01394(.A1(new_n1547_), .A2(new_n1376_), .ZN(new_n1587_));
  NAND4_X1   g01395(.A1(new_n1586_), .A2(new_n1573_), .A3(new_n1543_), .A4(new_n1587_), .ZN(new_n1588_));
  AOI21_X1   g01396(.A1(new_n1588_), .A2(new_n1584_), .B(new_n1389_), .ZN(new_n1589_));
  INV_X1     g01397(.I(new_n1587_), .ZN(new_n1590_));
  NOR4_X1    g01398(.A1(new_n1558_), .A2(new_n1585_), .A3(new_n1544_), .A4(new_n1590_), .ZN(new_n1591_));
  NOR3_X1    g01399(.A1(new_n1591_), .A2(new_n1579_), .A3(\a[102] ), .ZN(new_n1592_));
  AOI21_X1   g01400(.A1(\asqrt[50] ), .A2(\a[100] ), .B(new_n1554_), .ZN(new_n1593_));
  OAI21_X1   g01401(.A1(new_n1593_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n1594_));
  OAI22_X1   g01402(.A1(new_n1582_), .A2(new_n1594_), .B1(new_n1589_), .B2(new_n1592_), .ZN(new_n1595_));
  AOI21_X1   g01403(.A1(new_n1595_), .A2(new_n1583_), .B(new_n1103_), .ZN(new_n1596_));
  NOR3_X1    g01404(.A1(new_n1438_), .A2(new_n1388_), .A3(new_n1399_), .ZN(new_n1597_));
  NAND3_X1   g01405(.A1(\asqrt[50] ), .A2(new_n1421_), .A3(new_n1436_), .ZN(new_n1598_));
  AOI22_X1   g01406(.A1(new_n1598_), .A2(new_n1438_), .B1(\asqrt[50] ), .B2(new_n1597_), .ZN(new_n1599_));
  OAI21_X1   g01407(.A1(new_n1574_), .A2(new_n1554_), .B(\asqrt[51] ), .ZN(new_n1600_));
  AOI21_X1   g01408(.A1(new_n1573_), .A2(new_n1550_), .B(\a[100] ), .ZN(new_n1601_));
  OAI21_X1   g01409(.A1(new_n1580_), .A2(new_n1601_), .B(new_n1584_), .ZN(new_n1602_));
  OAI21_X1   g01410(.A1(new_n1602_), .A2(new_n1578_), .B(new_n1600_), .ZN(new_n1603_));
  AOI21_X1   g01411(.A1(new_n1603_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n1604_));
  AOI21_X1   g01412(.A1(new_n1604_), .A2(new_n1595_), .B(new_n1599_), .ZN(new_n1605_));
  OAI21_X1   g01413(.A1(new_n1605_), .A2(new_n1596_), .B(\asqrt[54] ), .ZN(new_n1606_));
  INV_X1     g01414(.I(new_n1606_), .ZN(new_n1607_));
  NOR2_X1    g01415(.A1(new_n1410_), .A2(new_n1413_), .ZN(new_n1608_));
  NOR2_X1    g01416(.A1(new_n1403_), .A2(new_n1415_), .ZN(new_n1609_));
  INV_X1     g01417(.I(new_n1609_), .ZN(new_n1610_));
  NAND4_X1   g01418(.A1(\asqrt[50] ), .A2(new_n1404_), .A3(new_n1608_), .A4(new_n1610_), .ZN(new_n1611_));
  INV_X1     g01419(.I(\asqrt[50] ), .ZN(new_n1612_));
  NOR3_X1    g01420(.A1(new_n1612_), .A2(new_n1440_), .A3(new_n1609_), .ZN(new_n1613_));
  OAI21_X1   g01421(.A1(new_n1613_), .A2(new_n1608_), .B(new_n1611_), .ZN(new_n1614_));
  INV_X1     g01422(.I(new_n1614_), .ZN(new_n1615_));
  NOR3_X1    g01423(.A1(new_n1605_), .A2(new_n1596_), .A3(\asqrt[54] ), .ZN(new_n1616_));
  NOR2_X1    g01424(.A1(new_n1616_), .A2(new_n1615_), .ZN(new_n1617_));
  OAI21_X1   g01425(.A1(new_n1617_), .A2(new_n1607_), .B(\asqrt[55] ), .ZN(new_n1618_));
  NOR2_X1    g01426(.A1(new_n1456_), .A2(new_n1445_), .ZN(new_n1619_));
  NOR3_X1    g01427(.A1(new_n1612_), .A2(new_n1417_), .A3(new_n1619_), .ZN(new_n1620_));
  INV_X1     g01428(.I(new_n1620_), .ZN(new_n1621_));
  NOR3_X1    g01429(.A1(new_n1619_), .A2(new_n1417_), .A3(new_n1455_), .ZN(new_n1622_));
  AOI22_X1   g01430(.A1(new_n1621_), .A2(new_n1455_), .B1(\asqrt[50] ), .B2(new_n1622_), .ZN(new_n1623_));
  INV_X1     g01431(.I(new_n1623_), .ZN(new_n1624_));
  NAND2_X1   g01432(.A1(new_n1606_), .A2(new_n823_), .ZN(new_n1625_));
  OAI21_X1   g01433(.A1(new_n1617_), .A2(new_n1625_), .B(new_n1624_), .ZN(new_n1626_));
  AOI21_X1   g01434(.A1(new_n1626_), .A2(new_n1618_), .B(new_n703_), .ZN(new_n1627_));
  NOR3_X1    g01435(.A1(new_n1458_), .A2(new_n1467_), .A3(new_n1434_), .ZN(new_n1628_));
  NOR3_X1    g01436(.A1(new_n1612_), .A2(new_n1458_), .A3(new_n1467_), .ZN(new_n1629_));
  INV_X1     g01437(.I(new_n1629_), .ZN(new_n1630_));
  AOI22_X1   g01438(.A1(new_n1630_), .A2(new_n1434_), .B1(\asqrt[50] ), .B2(new_n1628_), .ZN(new_n1631_));
  OAI21_X1   g01439(.A1(new_n1615_), .A2(new_n1616_), .B(new_n1606_), .ZN(new_n1632_));
  AOI21_X1   g01440(.A1(new_n1632_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n1633_));
  AOI21_X1   g01441(.A1(new_n1633_), .A2(new_n1626_), .B(new_n1631_), .ZN(new_n1634_));
  OAI21_X1   g01442(.A1(new_n1634_), .A2(new_n1627_), .B(\asqrt[57] ), .ZN(new_n1635_));
  INV_X1     g01443(.I(new_n1635_), .ZN(new_n1636_));
  NOR2_X1    g01444(.A1(new_n1468_), .A2(new_n1479_), .ZN(new_n1637_));
  NOR3_X1    g01445(.A1(new_n1612_), .A2(new_n1449_), .A3(new_n1637_), .ZN(new_n1638_));
  INV_X1     g01446(.I(new_n1638_), .ZN(new_n1639_));
  NOR3_X1    g01447(.A1(new_n1449_), .A2(new_n1637_), .A3(new_n1478_), .ZN(new_n1640_));
  AOI22_X1   g01448(.A1(new_n1639_), .A2(new_n1478_), .B1(\asqrt[50] ), .B2(new_n1640_), .ZN(new_n1641_));
  NOR3_X1    g01449(.A1(new_n1634_), .A2(new_n1627_), .A3(\asqrt[57] ), .ZN(new_n1642_));
  NOR2_X1    g01450(.A1(new_n1642_), .A2(new_n1641_), .ZN(new_n1643_));
  OAI21_X1   g01451(.A1(new_n1643_), .A2(new_n1636_), .B(\asqrt[58] ), .ZN(new_n1644_));
  NOR2_X1    g01452(.A1(new_n1470_), .A2(new_n1460_), .ZN(new_n1645_));
  NOR3_X1    g01453(.A1(new_n1645_), .A2(new_n1481_), .A3(new_n1466_), .ZN(new_n1646_));
  NOR3_X1    g01454(.A1(new_n1612_), .A2(new_n1481_), .A3(new_n1645_), .ZN(new_n1647_));
  INV_X1     g01455(.I(new_n1647_), .ZN(new_n1648_));
  AOI22_X1   g01456(.A1(new_n1648_), .A2(new_n1466_), .B1(\asqrt[50] ), .B2(new_n1646_), .ZN(new_n1649_));
  INV_X1     g01457(.I(new_n1649_), .ZN(new_n1650_));
  NAND2_X1   g01458(.A1(new_n1635_), .A2(new_n436_), .ZN(new_n1651_));
  OAI21_X1   g01459(.A1(new_n1643_), .A2(new_n1651_), .B(new_n1650_), .ZN(new_n1652_));
  AOI21_X1   g01460(.A1(new_n1652_), .A2(new_n1644_), .B(new_n327_), .ZN(new_n1653_));
  NOR3_X1    g01461(.A1(new_n1612_), .A2(new_n1472_), .A3(new_n1523_), .ZN(new_n1654_));
  INV_X1     g01462(.I(new_n1654_), .ZN(new_n1655_));
  NOR3_X1    g01463(.A1(new_n1472_), .A2(new_n1489_), .A3(new_n1523_), .ZN(new_n1656_));
  AOI22_X1   g01464(.A1(new_n1655_), .A2(new_n1489_), .B1(\asqrt[50] ), .B2(new_n1656_), .ZN(new_n1657_));
  OAI21_X1   g01465(.A1(new_n1641_), .A2(new_n1642_), .B(new_n1635_), .ZN(new_n1658_));
  AOI21_X1   g01466(.A1(new_n1658_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n1659_));
  AOI21_X1   g01467(.A1(new_n1659_), .A2(new_n1652_), .B(new_n1657_), .ZN(new_n1660_));
  OAI21_X1   g01468(.A1(new_n1660_), .A2(new_n1653_), .B(\asqrt[60] ), .ZN(new_n1661_));
  INV_X1     g01469(.I(new_n1661_), .ZN(new_n1662_));
  INV_X1     g01470(.I(new_n1660_), .ZN(new_n1663_));
  AND3_X2    g01471(.A1(new_n1484_), .A2(new_n1567_), .A3(new_n1495_), .Z(new_n1664_));
  NAND3_X1   g01472(.A1(\asqrt[50] ), .A2(new_n1484_), .A3(new_n1567_), .ZN(new_n1665_));
  AOI22_X1   g01473(.A1(new_n1665_), .A2(new_n1510_), .B1(\asqrt[50] ), .B2(new_n1664_), .ZN(new_n1666_));
  NOR2_X1    g01474(.A1(new_n1653_), .A2(\asqrt[60] ), .ZN(new_n1667_));
  AOI21_X1   g01475(.A1(new_n1663_), .A2(new_n1667_), .B(new_n1666_), .ZN(new_n1668_));
  OAI21_X1   g01476(.A1(new_n1668_), .A2(new_n1662_), .B(\asqrt[61] ), .ZN(new_n1669_));
  NOR2_X1    g01477(.A1(new_n1504_), .A2(new_n1497_), .ZN(new_n1670_));
  NOR3_X1    g01478(.A1(new_n1612_), .A2(new_n1514_), .A3(new_n1670_), .ZN(new_n1671_));
  INV_X1     g01479(.I(new_n1671_), .ZN(new_n1672_));
  NOR3_X1    g01480(.A1(new_n1670_), .A2(new_n1514_), .A3(new_n1503_), .ZN(new_n1673_));
  AOI22_X1   g01481(.A1(new_n1672_), .A2(new_n1503_), .B1(\asqrt[50] ), .B2(new_n1673_), .ZN(new_n1674_));
  INV_X1     g01482(.I(new_n1674_), .ZN(new_n1675_));
  NAND2_X1   g01483(.A1(new_n1661_), .A2(new_n218_), .ZN(new_n1676_));
  OAI21_X1   g01484(.A1(new_n1676_), .A2(new_n1668_), .B(new_n1675_), .ZN(new_n1677_));
  AOI21_X1   g01485(.A1(new_n1677_), .A2(new_n1669_), .B(new_n207_), .ZN(new_n1678_));
  NOR3_X1    g01486(.A1(new_n1506_), .A2(new_n1538_), .A3(new_n1566_), .ZN(new_n1679_));
  NOR3_X1    g01487(.A1(new_n1612_), .A2(new_n1506_), .A3(new_n1538_), .ZN(new_n1680_));
  INV_X1     g01488(.I(new_n1680_), .ZN(new_n1681_));
  AOI22_X1   g01489(.A1(new_n1681_), .A2(new_n1566_), .B1(\asqrt[50] ), .B2(new_n1679_), .ZN(new_n1682_));
  NOR3_X1    g01490(.A1(new_n1660_), .A2(new_n1653_), .A3(\asqrt[60] ), .ZN(new_n1683_));
  OAI21_X1   g01491(.A1(new_n1666_), .A2(new_n1683_), .B(new_n1661_), .ZN(new_n1684_));
  AOI21_X1   g01492(.A1(new_n1684_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n1685_));
  AOI21_X1   g01493(.A1(new_n1685_), .A2(new_n1677_), .B(new_n1682_), .ZN(new_n1686_));
  INV_X1     g01494(.I(new_n1517_), .ZN(new_n1687_));
  NOR2_X1    g01495(.A1(new_n1528_), .A2(new_n1516_), .ZN(new_n1688_));
  NOR3_X1    g01496(.A1(new_n1687_), .A2(new_n1522_), .A3(new_n1688_), .ZN(new_n1689_));
  NAND2_X1   g01497(.A1(\asqrt[50] ), .A2(new_n1689_), .ZN(new_n1690_));
  INV_X1     g01498(.I(new_n1690_), .ZN(new_n1691_));
  NOR2_X1    g01499(.A1(new_n1687_), .A2(new_n1688_), .ZN(new_n1692_));
  AOI21_X1   g01500(.A1(\asqrt[50] ), .A2(new_n1692_), .B(new_n1521_), .ZN(new_n1693_));
  NOR2_X1    g01501(.A1(new_n1691_), .A2(new_n1693_), .ZN(new_n1694_));
  NOR3_X1    g01502(.A1(new_n1612_), .A2(new_n1572_), .A3(new_n1560_), .ZN(new_n1695_));
  NOR3_X1    g01503(.A1(new_n1694_), .A2(new_n1585_), .A3(new_n1695_), .ZN(new_n1696_));
  OAI21_X1   g01504(.A1(new_n1686_), .A2(new_n1678_), .B(new_n1696_), .ZN(new_n1697_));
  NAND2_X1   g01505(.A1(new_n1697_), .A2(new_n193_), .ZN(new_n1698_));
  INV_X1     g01506(.I(new_n1682_), .ZN(new_n1699_));
  NAND3_X1   g01507(.A1(new_n1677_), .A2(new_n1669_), .A3(new_n207_), .ZN(new_n1700_));
  NAND2_X1   g01508(.A1(new_n1700_), .A2(new_n1699_), .ZN(new_n1701_));
  INV_X1     g01509(.I(new_n1694_), .ZN(new_n1702_));
  NOR2_X1    g01510(.A1(new_n1678_), .A2(new_n1702_), .ZN(new_n1703_));
  AOI21_X1   g01511(.A1(\asqrt[50] ), .A2(new_n1533_), .B(new_n1556_), .ZN(new_n1704_));
  AOI21_X1   g01512(.A1(new_n1556_), .A2(new_n1533_), .B(new_n193_), .ZN(new_n1705_));
  INV_X1     g01513(.I(new_n1705_), .ZN(new_n1706_));
  NOR2_X1    g01514(.A1(new_n1704_), .A2(new_n1706_), .ZN(new_n1707_));
  AND3_X2    g01515(.A1(new_n1532_), .A2(new_n1530_), .A3(new_n1546_), .Z(new_n1708_));
  NAND4_X1   g01516(.A1(new_n1586_), .A2(new_n1573_), .A3(new_n1543_), .A4(new_n1708_), .ZN(new_n1709_));
  INV_X1     g01517(.I(new_n1709_), .ZN(new_n1710_));
  NOR2_X1    g01518(.A1(new_n1707_), .A2(new_n1710_), .ZN(new_n1711_));
  INV_X1     g01519(.I(new_n1711_), .ZN(new_n1712_));
  AOI21_X1   g01520(.A1(new_n1703_), .A2(new_n1701_), .B(new_n1712_), .ZN(new_n1713_));
  NAND2_X1   g01521(.A1(new_n1698_), .A2(new_n1713_), .ZN(\asqrt[49] ));
  NOR2_X1    g01522(.A1(\a[96] ), .A2(\a[97] ), .ZN(new_n1715_));
  INV_X1     g01523(.I(new_n1715_), .ZN(new_n1716_));
  NOR2_X1    g01524(.A1(new_n1716_), .A2(\a[98] ), .ZN(new_n1717_));
  INV_X1     g01525(.I(new_n1717_), .ZN(new_n1718_));
  INV_X1     g01526(.I(new_n1666_), .ZN(new_n1719_));
  INV_X1     g01527(.I(new_n1641_), .ZN(new_n1720_));
  NAND2_X1   g01528(.A1(new_n1563_), .A2(new_n1576_), .ZN(new_n1721_));
  OAI21_X1   g01529(.A1(new_n1558_), .A2(new_n1562_), .B(new_n1565_), .ZN(new_n1722_));
  NAND2_X1   g01530(.A1(new_n1722_), .A2(\a[101] ), .ZN(new_n1723_));
  NAND3_X1   g01531(.A1(new_n1721_), .A2(new_n1723_), .A3(new_n1584_), .ZN(new_n1724_));
  AOI21_X1   g01532(.A1(new_n1724_), .A2(new_n1600_), .B(new_n1256_), .ZN(new_n1725_));
  OAI21_X1   g01533(.A1(new_n1591_), .A2(new_n1579_), .B(\a[102] ), .ZN(new_n1726_));
  NAND3_X1   g01534(.A1(new_n1588_), .A2(new_n1584_), .A3(new_n1389_), .ZN(new_n1727_));
  NAND2_X1   g01535(.A1(new_n1563_), .A2(new_n1555_), .ZN(new_n1728_));
  AOI21_X1   g01536(.A1(new_n1728_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n1729_));
  AOI22_X1   g01537(.A1(new_n1724_), .A2(new_n1729_), .B1(new_n1726_), .B2(new_n1727_), .ZN(new_n1730_));
  OAI21_X1   g01538(.A1(new_n1730_), .A2(new_n1725_), .B(\asqrt[53] ), .ZN(new_n1731_));
  NAND2_X1   g01539(.A1(new_n1731_), .A2(new_n904_), .ZN(new_n1732_));
  OAI21_X1   g01540(.A1(new_n1732_), .A2(new_n1605_), .B(new_n1614_), .ZN(new_n1733_));
  AOI21_X1   g01541(.A1(new_n1733_), .A2(new_n1606_), .B(new_n823_), .ZN(new_n1734_));
  INV_X1     g01542(.I(new_n1599_), .ZN(new_n1735_));
  AOI21_X1   g01543(.A1(\a[101] ), .A2(new_n1722_), .B(new_n1579_), .ZN(new_n1736_));
  AOI21_X1   g01544(.A1(new_n1736_), .A2(new_n1721_), .B(new_n1564_), .ZN(new_n1737_));
  OAI21_X1   g01545(.A1(new_n1737_), .A2(new_n1256_), .B(new_n1103_), .ZN(new_n1738_));
  OAI21_X1   g01546(.A1(new_n1738_), .A2(new_n1730_), .B(new_n1735_), .ZN(new_n1739_));
  NAND2_X1   g01547(.A1(new_n1739_), .A2(new_n1731_), .ZN(new_n1740_));
  AOI21_X1   g01548(.A1(new_n1740_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1741_));
  AOI21_X1   g01549(.A1(new_n1741_), .A2(new_n1733_), .B(new_n1623_), .ZN(new_n1742_));
  OAI21_X1   g01550(.A1(new_n1742_), .A2(new_n1734_), .B(\asqrt[56] ), .ZN(new_n1743_));
  NAND2_X1   g01551(.A1(new_n1743_), .A2(new_n531_), .ZN(new_n1744_));
  OAI21_X1   g01552(.A1(new_n1744_), .A2(new_n1634_), .B(new_n1720_), .ZN(new_n1745_));
  NAND3_X1   g01553(.A1(new_n1745_), .A2(new_n436_), .A3(new_n1635_), .ZN(new_n1746_));
  AOI22_X1   g01554(.A1(new_n1746_), .A2(new_n1650_), .B1(new_n1658_), .B2(\asqrt[58] ), .ZN(new_n1747_));
  OAI21_X1   g01555(.A1(new_n1747_), .A2(new_n327_), .B(new_n306_), .ZN(new_n1748_));
  OAI21_X1   g01556(.A1(new_n1748_), .A2(new_n1660_), .B(new_n1719_), .ZN(new_n1749_));
  AOI21_X1   g01557(.A1(new_n1749_), .A2(new_n1661_), .B(new_n218_), .ZN(new_n1750_));
  AOI21_X1   g01558(.A1(new_n1745_), .A2(new_n1635_), .B(new_n436_), .ZN(new_n1751_));
  NOR3_X1    g01559(.A1(new_n1742_), .A2(new_n1734_), .A3(\asqrt[56] ), .ZN(new_n1752_));
  OAI21_X1   g01560(.A1(new_n1631_), .A2(new_n1752_), .B(new_n1743_), .ZN(new_n1753_));
  AOI21_X1   g01561(.A1(new_n1753_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n1754_));
  AOI21_X1   g01562(.A1(new_n1754_), .A2(new_n1745_), .B(new_n1649_), .ZN(new_n1755_));
  NOR3_X1    g01563(.A1(new_n1755_), .A2(\asqrt[59] ), .A3(new_n1751_), .ZN(new_n1756_));
  OAI22_X1   g01564(.A1(new_n1756_), .A2(new_n1657_), .B1(new_n1747_), .B2(new_n327_), .ZN(new_n1757_));
  AOI21_X1   g01565(.A1(new_n1757_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n1758_));
  AOI21_X1   g01566(.A1(new_n1758_), .A2(new_n1749_), .B(new_n1674_), .ZN(new_n1759_));
  OAI21_X1   g01567(.A1(new_n1759_), .A2(new_n1750_), .B(\asqrt[62] ), .ZN(new_n1760_));
  NOR3_X1    g01568(.A1(new_n1759_), .A2(\asqrt[62] ), .A3(new_n1750_), .ZN(new_n1761_));
  OAI21_X1   g01569(.A1(new_n1682_), .A2(new_n1761_), .B(new_n1760_), .ZN(new_n1762_));
  AOI21_X1   g01570(.A1(new_n1762_), .A2(new_n1696_), .B(\asqrt[63] ), .ZN(new_n1763_));
  NAND2_X1   g01571(.A1(new_n1760_), .A2(new_n1694_), .ZN(new_n1764_));
  OAI21_X1   g01572(.A1(new_n1764_), .A2(new_n1686_), .B(new_n1711_), .ZN(new_n1765_));
  OAI21_X1   g01573(.A1(new_n1763_), .A2(new_n1765_), .B(\a[98] ), .ZN(new_n1766_));
  AOI21_X1   g01574(.A1(new_n1766_), .A2(new_n1718_), .B(new_n1612_), .ZN(new_n1767_));
  INV_X1     g01575(.I(\a[98] ), .ZN(new_n1768_));
  AOI21_X1   g01576(.A1(new_n1698_), .A2(new_n1713_), .B(new_n1768_), .ZN(new_n1769_));
  NAND2_X1   g01577(.A1(new_n1546_), .A2(new_n1718_), .ZN(new_n1770_));
  NOR4_X1    g01578(.A1(new_n1558_), .A2(new_n1585_), .A3(new_n1544_), .A4(new_n1770_), .ZN(new_n1771_));
  INV_X1     g01579(.I(new_n1771_), .ZN(new_n1772_));
  NOR2_X1    g01580(.A1(new_n1769_), .A2(new_n1772_), .ZN(new_n1773_));
  AOI21_X1   g01581(.A1(new_n1698_), .A2(new_n1713_), .B(new_n1553_), .ZN(new_n1774_));
  INV_X1     g01582(.I(\a[99] ), .ZN(new_n1775_));
  AOI21_X1   g01583(.A1(\asqrt[49] ), .A2(new_n1768_), .B(new_n1775_), .ZN(new_n1776_));
  NOR3_X1    g01584(.A1(new_n1773_), .A2(new_n1776_), .A3(new_n1774_), .ZN(new_n1777_));
  OAI21_X1   g01585(.A1(new_n1777_), .A2(new_n1767_), .B(\asqrt[51] ), .ZN(new_n1778_));
  OAI21_X1   g01586(.A1(new_n1763_), .A2(new_n1765_), .B(new_n1552_), .ZN(new_n1779_));
  NAND2_X1   g01587(.A1(new_n1703_), .A2(new_n1701_), .ZN(new_n1780_));
  INV_X1     g01588(.I(new_n1707_), .ZN(new_n1781_));
  NOR2_X1    g01589(.A1(new_n1710_), .A2(new_n1612_), .ZN(new_n1782_));
  NAND4_X1   g01590(.A1(new_n1698_), .A2(new_n1780_), .A3(new_n1781_), .A4(new_n1782_), .ZN(new_n1783_));
  AOI21_X1   g01591(.A1(new_n1783_), .A2(new_n1779_), .B(new_n1565_), .ZN(new_n1784_));
  INV_X1     g01592(.I(new_n1780_), .ZN(new_n1785_));
  NAND2_X1   g01593(.A1(new_n1781_), .A2(new_n1782_), .ZN(new_n1786_));
  NOR3_X1    g01594(.A1(new_n1785_), .A2(new_n1763_), .A3(new_n1786_), .ZN(new_n1787_));
  NOR3_X1    g01595(.A1(new_n1787_), .A2(new_n1774_), .A3(\a[100] ), .ZN(new_n1788_));
  OAI21_X1   g01596(.A1(new_n1769_), .A2(new_n1717_), .B(\asqrt[50] ), .ZN(new_n1789_));
  NAND2_X1   g01597(.A1(new_n1789_), .A2(new_n1376_), .ZN(new_n1790_));
  OAI22_X1   g01598(.A1(new_n1777_), .A2(new_n1790_), .B1(new_n1784_), .B2(new_n1788_), .ZN(new_n1791_));
  AOI21_X1   g01599(.A1(new_n1791_), .A2(new_n1778_), .B(new_n1256_), .ZN(new_n1792_));
  NOR3_X1    g01600(.A1(new_n1736_), .A2(new_n1564_), .A3(new_n1578_), .ZN(new_n1793_));
  NAND3_X1   g01601(.A1(\asqrt[49] ), .A2(new_n1600_), .A3(new_n1721_), .ZN(new_n1794_));
  AOI22_X1   g01602(.A1(new_n1794_), .A2(new_n1736_), .B1(\asqrt[49] ), .B2(new_n1793_), .ZN(new_n1795_));
  AOI21_X1   g01603(.A1(new_n1698_), .A2(new_n1713_), .B(\a[98] ), .ZN(new_n1796_));
  OAI21_X1   g01604(.A1(new_n1775_), .A2(new_n1796_), .B(new_n1779_), .ZN(new_n1797_));
  OAI21_X1   g01605(.A1(new_n1797_), .A2(new_n1773_), .B(new_n1789_), .ZN(new_n1798_));
  AOI21_X1   g01606(.A1(new_n1798_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n1799_));
  AOI21_X1   g01607(.A1(new_n1799_), .A2(new_n1791_), .B(new_n1795_), .ZN(new_n1800_));
  OAI21_X1   g01608(.A1(new_n1800_), .A2(new_n1792_), .B(\asqrt[53] ), .ZN(new_n1801_));
  NOR2_X1    g01609(.A1(new_n1589_), .A2(new_n1592_), .ZN(new_n1802_));
  NOR2_X1    g01610(.A1(new_n1582_), .A2(new_n1594_), .ZN(new_n1803_));
  INV_X1     g01611(.I(new_n1803_), .ZN(new_n1804_));
  NAND4_X1   g01612(.A1(\asqrt[49] ), .A2(new_n1583_), .A3(new_n1802_), .A4(new_n1804_), .ZN(new_n1805_));
  INV_X1     g01613(.I(\asqrt[49] ), .ZN(new_n1806_));
  NOR3_X1    g01614(.A1(new_n1806_), .A2(new_n1725_), .A3(new_n1803_), .ZN(new_n1807_));
  OAI21_X1   g01615(.A1(new_n1807_), .A2(new_n1802_), .B(new_n1805_), .ZN(new_n1808_));
  NAND2_X1   g01616(.A1(new_n1766_), .A2(new_n1771_), .ZN(new_n1809_));
  OAI21_X1   g01617(.A1(new_n1763_), .A2(new_n1765_), .B(new_n1768_), .ZN(new_n1810_));
  NAND2_X1   g01618(.A1(new_n1810_), .A2(\a[99] ), .ZN(new_n1811_));
  NAND3_X1   g01619(.A1(new_n1809_), .A2(new_n1811_), .A3(new_n1779_), .ZN(new_n1812_));
  AOI21_X1   g01620(.A1(new_n1812_), .A2(new_n1789_), .B(new_n1376_), .ZN(new_n1813_));
  OAI21_X1   g01621(.A1(new_n1787_), .A2(new_n1774_), .B(\a[100] ), .ZN(new_n1814_));
  NAND3_X1   g01622(.A1(new_n1783_), .A2(new_n1779_), .A3(new_n1565_), .ZN(new_n1815_));
  NAND2_X1   g01623(.A1(new_n1766_), .A2(new_n1718_), .ZN(new_n1816_));
  AOI21_X1   g01624(.A1(new_n1816_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n1817_));
  AOI22_X1   g01625(.A1(new_n1812_), .A2(new_n1817_), .B1(new_n1814_), .B2(new_n1815_), .ZN(new_n1818_));
  OAI21_X1   g01626(.A1(new_n1818_), .A2(new_n1813_), .B(\asqrt[52] ), .ZN(new_n1819_));
  NAND2_X1   g01627(.A1(new_n1819_), .A2(new_n1103_), .ZN(new_n1820_));
  OAI21_X1   g01628(.A1(new_n1820_), .A2(new_n1800_), .B(new_n1808_), .ZN(new_n1821_));
  AOI21_X1   g01629(.A1(new_n1821_), .A2(new_n1801_), .B(new_n904_), .ZN(new_n1822_));
  NOR2_X1    g01630(.A1(new_n1738_), .A2(new_n1730_), .ZN(new_n1823_));
  NOR3_X1    g01631(.A1(new_n1806_), .A2(new_n1596_), .A3(new_n1823_), .ZN(new_n1824_));
  INV_X1     g01632(.I(new_n1824_), .ZN(new_n1825_));
  NOR3_X1    g01633(.A1(new_n1823_), .A2(new_n1596_), .A3(new_n1735_), .ZN(new_n1826_));
  AOI22_X1   g01634(.A1(new_n1825_), .A2(new_n1735_), .B1(\asqrt[49] ), .B2(new_n1826_), .ZN(new_n1827_));
  INV_X1     g01635(.I(new_n1795_), .ZN(new_n1828_));
  AOI21_X1   g01636(.A1(\a[99] ), .A2(new_n1810_), .B(new_n1774_), .ZN(new_n1829_));
  AOI21_X1   g01637(.A1(new_n1829_), .A2(new_n1809_), .B(new_n1767_), .ZN(new_n1830_));
  OAI21_X1   g01638(.A1(new_n1830_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n1831_));
  OAI21_X1   g01639(.A1(new_n1831_), .A2(new_n1818_), .B(new_n1828_), .ZN(new_n1832_));
  NAND2_X1   g01640(.A1(new_n1832_), .A2(new_n1819_), .ZN(new_n1833_));
  AOI21_X1   g01641(.A1(new_n1833_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n1834_));
  AOI21_X1   g01642(.A1(new_n1834_), .A2(new_n1821_), .B(new_n1827_), .ZN(new_n1835_));
  OAI21_X1   g01643(.A1(new_n1835_), .A2(new_n1822_), .B(\asqrt[55] ), .ZN(new_n1836_));
  NOR3_X1    g01644(.A1(new_n1607_), .A2(new_n1616_), .A3(new_n1614_), .ZN(new_n1837_));
  NOR3_X1    g01645(.A1(new_n1806_), .A2(new_n1607_), .A3(new_n1616_), .ZN(new_n1838_));
  INV_X1     g01646(.I(new_n1838_), .ZN(new_n1839_));
  AOI22_X1   g01647(.A1(new_n1839_), .A2(new_n1614_), .B1(\asqrt[49] ), .B2(new_n1837_), .ZN(new_n1840_));
  INV_X1     g01648(.I(new_n1840_), .ZN(new_n1841_));
  INV_X1     g01649(.I(new_n1801_), .ZN(new_n1842_));
  INV_X1     g01650(.I(new_n1808_), .ZN(new_n1843_));
  NOR3_X1    g01651(.A1(new_n1800_), .A2(new_n1792_), .A3(\asqrt[53] ), .ZN(new_n1844_));
  NOR2_X1    g01652(.A1(new_n1844_), .A2(new_n1843_), .ZN(new_n1845_));
  OAI21_X1   g01653(.A1(new_n1845_), .A2(new_n1842_), .B(\asqrt[54] ), .ZN(new_n1846_));
  NAND2_X1   g01654(.A1(new_n1846_), .A2(new_n823_), .ZN(new_n1847_));
  OAI21_X1   g01655(.A1(new_n1847_), .A2(new_n1835_), .B(new_n1841_), .ZN(new_n1848_));
  AOI21_X1   g01656(.A1(new_n1848_), .A2(new_n1836_), .B(new_n703_), .ZN(new_n1849_));
  NOR2_X1    g01657(.A1(new_n1617_), .A2(new_n1625_), .ZN(new_n1850_));
  NOR3_X1    g01658(.A1(new_n1806_), .A2(new_n1734_), .A3(new_n1850_), .ZN(new_n1851_));
  INV_X1     g01659(.I(new_n1851_), .ZN(new_n1852_));
  NOR3_X1    g01660(.A1(new_n1850_), .A2(new_n1734_), .A3(new_n1624_), .ZN(new_n1853_));
  AOI22_X1   g01661(.A1(new_n1852_), .A2(new_n1624_), .B1(\asqrt[49] ), .B2(new_n1853_), .ZN(new_n1854_));
  INV_X1     g01662(.I(new_n1827_), .ZN(new_n1855_));
  NAND2_X1   g01663(.A1(new_n1801_), .A2(new_n904_), .ZN(new_n1856_));
  OAI21_X1   g01664(.A1(new_n1845_), .A2(new_n1856_), .B(new_n1855_), .ZN(new_n1857_));
  NAND2_X1   g01665(.A1(new_n1857_), .A2(new_n1846_), .ZN(new_n1858_));
  AOI21_X1   g01666(.A1(new_n1858_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n1859_));
  AOI21_X1   g01667(.A1(new_n1859_), .A2(new_n1848_), .B(new_n1854_), .ZN(new_n1860_));
  OAI21_X1   g01668(.A1(new_n1860_), .A2(new_n1849_), .B(\asqrt[57] ), .ZN(new_n1861_));
  INV_X1     g01669(.I(new_n1631_), .ZN(new_n1862_));
  NOR3_X1    g01670(.A1(new_n1627_), .A2(new_n1752_), .A3(new_n1862_), .ZN(new_n1863_));
  NOR3_X1    g01671(.A1(new_n1806_), .A2(new_n1627_), .A3(new_n1752_), .ZN(new_n1864_));
  INV_X1     g01672(.I(new_n1864_), .ZN(new_n1865_));
  AOI22_X1   g01673(.A1(new_n1865_), .A2(new_n1862_), .B1(\asqrt[49] ), .B2(new_n1863_), .ZN(new_n1866_));
  INV_X1     g01674(.I(new_n1866_), .ZN(new_n1867_));
  AOI21_X1   g01675(.A1(new_n1857_), .A2(new_n1846_), .B(new_n823_), .ZN(new_n1868_));
  OAI21_X1   g01676(.A1(new_n1843_), .A2(new_n1844_), .B(new_n1801_), .ZN(new_n1869_));
  AOI21_X1   g01677(.A1(new_n1869_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n1870_));
  AOI21_X1   g01678(.A1(new_n1870_), .A2(new_n1857_), .B(new_n1840_), .ZN(new_n1871_));
  OAI21_X1   g01679(.A1(new_n1871_), .A2(new_n1868_), .B(\asqrt[56] ), .ZN(new_n1872_));
  INV_X1     g01680(.I(new_n1854_), .ZN(new_n1873_));
  NAND2_X1   g01681(.A1(new_n1836_), .A2(new_n703_), .ZN(new_n1874_));
  OAI21_X1   g01682(.A1(new_n1874_), .A2(new_n1871_), .B(new_n1873_), .ZN(new_n1875_));
  NAND3_X1   g01683(.A1(new_n1875_), .A2(new_n531_), .A3(new_n1872_), .ZN(new_n1876_));
  NAND2_X1   g01684(.A1(new_n1876_), .A2(new_n1867_), .ZN(new_n1877_));
  AOI21_X1   g01685(.A1(new_n1877_), .A2(new_n1861_), .B(new_n436_), .ZN(new_n1878_));
  NOR3_X1    g01686(.A1(new_n1806_), .A2(new_n1636_), .A3(new_n1642_), .ZN(new_n1879_));
  INV_X1     g01687(.I(new_n1879_), .ZN(new_n1880_));
  NOR3_X1    g01688(.A1(new_n1636_), .A2(new_n1720_), .A3(new_n1642_), .ZN(new_n1881_));
  AOI22_X1   g01689(.A1(new_n1880_), .A2(new_n1720_), .B1(\asqrt[49] ), .B2(new_n1881_), .ZN(new_n1882_));
  AOI21_X1   g01690(.A1(new_n1875_), .A2(new_n1872_), .B(new_n531_), .ZN(new_n1883_));
  NOR2_X1    g01691(.A1(new_n1883_), .A2(\asqrt[58] ), .ZN(new_n1884_));
  AOI21_X1   g01692(.A1(new_n1884_), .A2(new_n1877_), .B(new_n1882_), .ZN(new_n1885_));
  OAI21_X1   g01693(.A1(new_n1885_), .A2(new_n1878_), .B(\asqrt[59] ), .ZN(new_n1886_));
  INV_X1     g01694(.I(new_n1886_), .ZN(new_n1887_));
  INV_X1     g01695(.I(new_n1746_), .ZN(new_n1888_));
  NOR3_X1    g01696(.A1(new_n1888_), .A2(new_n1751_), .A3(new_n1650_), .ZN(new_n1889_));
  NOR3_X1    g01697(.A1(new_n1806_), .A2(new_n1751_), .A3(new_n1888_), .ZN(new_n1890_));
  INV_X1     g01698(.I(new_n1890_), .ZN(new_n1891_));
  AOI22_X1   g01699(.A1(new_n1891_), .A2(new_n1650_), .B1(\asqrt[49] ), .B2(new_n1889_), .ZN(new_n1892_));
  NOR3_X1    g01700(.A1(new_n1885_), .A2(new_n1878_), .A3(\asqrt[59] ), .ZN(new_n1893_));
  NOR2_X1    g01701(.A1(new_n1893_), .A2(new_n1892_), .ZN(new_n1894_));
  OAI21_X1   g01702(.A1(new_n1894_), .A2(new_n1887_), .B(\asqrt[60] ), .ZN(new_n1895_));
  INV_X1     g01703(.I(new_n1657_), .ZN(new_n1896_));
  NOR3_X1    g01704(.A1(new_n1806_), .A2(new_n1653_), .A3(new_n1756_), .ZN(new_n1897_));
  INV_X1     g01705(.I(new_n1897_), .ZN(new_n1898_));
  NOR3_X1    g01706(.A1(new_n1653_), .A2(new_n1756_), .A3(new_n1896_), .ZN(new_n1899_));
  AOI22_X1   g01707(.A1(new_n1898_), .A2(new_n1896_), .B1(\asqrt[49] ), .B2(new_n1899_), .ZN(new_n1900_));
  INV_X1     g01708(.I(new_n1900_), .ZN(new_n1901_));
  NAND2_X1   g01709(.A1(new_n1886_), .A2(new_n306_), .ZN(new_n1902_));
  OAI21_X1   g01710(.A1(new_n1894_), .A2(new_n1902_), .B(new_n1901_), .ZN(new_n1903_));
  AOI21_X1   g01711(.A1(new_n1903_), .A2(new_n1895_), .B(new_n218_), .ZN(new_n1904_));
  NOR3_X1    g01712(.A1(new_n1662_), .A2(new_n1719_), .A3(new_n1683_), .ZN(new_n1905_));
  NOR3_X1    g01713(.A1(new_n1806_), .A2(new_n1662_), .A3(new_n1683_), .ZN(new_n1906_));
  INV_X1     g01714(.I(new_n1906_), .ZN(new_n1907_));
  AOI22_X1   g01715(.A1(new_n1907_), .A2(new_n1719_), .B1(\asqrt[49] ), .B2(new_n1905_), .ZN(new_n1908_));
  INV_X1     g01716(.I(new_n1892_), .ZN(new_n1909_));
  NOR3_X1    g01717(.A1(new_n1835_), .A2(new_n1822_), .A3(\asqrt[55] ), .ZN(new_n1910_));
  OAI21_X1   g01718(.A1(new_n1840_), .A2(new_n1910_), .B(new_n1836_), .ZN(new_n1911_));
  AOI21_X1   g01719(.A1(new_n1911_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n1912_));
  AOI21_X1   g01720(.A1(new_n1912_), .A2(new_n1875_), .B(new_n1866_), .ZN(new_n1913_));
  OAI21_X1   g01721(.A1(new_n1913_), .A2(new_n1883_), .B(\asqrt[58] ), .ZN(new_n1914_));
  NAND2_X1   g01722(.A1(new_n1914_), .A2(new_n327_), .ZN(new_n1915_));
  OAI21_X1   g01723(.A1(new_n1915_), .A2(new_n1885_), .B(new_n1909_), .ZN(new_n1916_));
  AOI21_X1   g01724(.A1(new_n1916_), .A2(new_n1886_), .B(new_n306_), .ZN(new_n1917_));
  NOR2_X1    g01725(.A1(new_n1917_), .A2(\asqrt[61] ), .ZN(new_n1918_));
  AOI21_X1   g01726(.A1(new_n1918_), .A2(new_n1903_), .B(new_n1908_), .ZN(new_n1919_));
  OAI21_X1   g01727(.A1(new_n1919_), .A2(new_n1904_), .B(\asqrt[62] ), .ZN(new_n1920_));
  NOR2_X1    g01728(.A1(new_n1676_), .A2(new_n1668_), .ZN(new_n1921_));
  NOR3_X1    g01729(.A1(new_n1806_), .A2(new_n1750_), .A3(new_n1921_), .ZN(new_n1922_));
  INV_X1     g01730(.I(new_n1922_), .ZN(new_n1923_));
  NOR3_X1    g01731(.A1(new_n1921_), .A2(new_n1750_), .A3(new_n1675_), .ZN(new_n1924_));
  AOI22_X1   g01732(.A1(new_n1923_), .A2(new_n1675_), .B1(\asqrt[49] ), .B2(new_n1924_), .ZN(new_n1925_));
  INV_X1     g01733(.I(new_n1925_), .ZN(new_n1926_));
  NOR3_X1    g01734(.A1(new_n1871_), .A2(new_n1868_), .A3(\asqrt[56] ), .ZN(new_n1927_));
  OAI21_X1   g01735(.A1(new_n1854_), .A2(new_n1927_), .B(new_n1872_), .ZN(new_n1928_));
  AOI22_X1   g01736(.A1(new_n1876_), .A2(new_n1867_), .B1(new_n1928_), .B2(\asqrt[57] ), .ZN(new_n1929_));
  NOR3_X1    g01737(.A1(new_n1913_), .A2(\asqrt[58] ), .A3(new_n1883_), .ZN(new_n1930_));
  OAI22_X1   g01738(.A1(new_n1930_), .A2(new_n1882_), .B1(new_n1929_), .B2(new_n436_), .ZN(new_n1931_));
  AOI21_X1   g01739(.A1(new_n1931_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n1932_));
  AOI21_X1   g01740(.A1(new_n1932_), .A2(new_n1916_), .B(new_n1900_), .ZN(new_n1933_));
  OAI21_X1   g01741(.A1(new_n1933_), .A2(new_n1917_), .B(\asqrt[61] ), .ZN(new_n1934_));
  NAND2_X1   g01742(.A1(new_n1934_), .A2(new_n207_), .ZN(new_n1935_));
  OAI21_X1   g01743(.A1(new_n1935_), .A2(new_n1919_), .B(new_n1926_), .ZN(new_n1936_));
  NAND4_X1   g01744(.A1(\asqrt[49] ), .A2(new_n1760_), .A3(new_n1682_), .A4(new_n1700_), .ZN(new_n1937_));
  NAND2_X1   g01745(.A1(new_n1700_), .A2(new_n1760_), .ZN(new_n1938_));
  OAI21_X1   g01746(.A1(new_n1806_), .A2(new_n1938_), .B(new_n1699_), .ZN(new_n1939_));
  NAND2_X1   g01747(.A1(new_n1939_), .A2(new_n1937_), .ZN(new_n1940_));
  AOI21_X1   g01748(.A1(new_n1701_), .A2(new_n1760_), .B(new_n1694_), .ZN(new_n1941_));
  AOI21_X1   g01749(.A1(\asqrt[49] ), .A2(new_n1941_), .B(new_n1785_), .ZN(new_n1942_));
  NAND2_X1   g01750(.A1(new_n1940_), .A2(new_n1942_), .ZN(new_n1943_));
  AOI21_X1   g01751(.A1(new_n1936_), .A2(new_n1920_), .B(new_n1943_), .ZN(new_n1944_));
  NOR3_X1    g01752(.A1(new_n1933_), .A2(\asqrt[61] ), .A3(new_n1917_), .ZN(new_n1945_));
  OAI21_X1   g01753(.A1(new_n1908_), .A2(new_n1945_), .B(new_n1934_), .ZN(new_n1946_));
  AOI21_X1   g01754(.A1(new_n1946_), .A2(\asqrt[62] ), .B(new_n1940_), .ZN(new_n1947_));
  AOI21_X1   g01755(.A1(\asqrt[49] ), .A2(new_n1702_), .B(new_n1762_), .ZN(new_n1948_));
  OR3_X2     g01756(.A1(new_n1948_), .A2(new_n193_), .A3(new_n1941_), .Z(new_n1949_));
  NAND2_X1   g01757(.A1(new_n1690_), .A2(new_n1709_), .ZN(new_n1950_));
  NOR4_X1    g01758(.A1(new_n1785_), .A2(new_n1693_), .A3(new_n1707_), .A4(new_n1950_), .ZN(new_n1951_));
  NAND2_X1   g01759(.A1(new_n1951_), .A2(new_n1698_), .ZN(new_n1952_));
  NAND2_X1   g01760(.A1(new_n1949_), .A2(new_n1952_), .ZN(new_n1953_));
  AOI21_X1   g01761(.A1(new_n1947_), .A2(new_n1936_), .B(new_n1953_), .ZN(new_n1954_));
  OAI21_X1   g01762(.A1(\asqrt[63] ), .A2(new_n1944_), .B(new_n1954_), .ZN(\asqrt[48] ));
  INV_X1     g01763(.I(\asqrt[48] ), .ZN(new_n1956_));
  NOR2_X1    g01764(.A1(\a[94] ), .A2(\a[95] ), .ZN(new_n1957_));
  INV_X1     g01765(.I(new_n1957_), .ZN(new_n1958_));
  NOR2_X1    g01766(.A1(new_n1958_), .A2(\a[96] ), .ZN(new_n1959_));
  INV_X1     g01767(.I(new_n1959_), .ZN(new_n1960_));
  NOR2_X1    g01768(.A1(new_n1944_), .A2(\asqrt[63] ), .ZN(new_n1961_));
  INV_X1     g01769(.I(new_n1936_), .ZN(new_n1962_));
  INV_X1     g01770(.I(new_n1940_), .ZN(new_n1963_));
  NAND2_X1   g01771(.A1(new_n1920_), .A2(new_n1963_), .ZN(new_n1964_));
  INV_X1     g01772(.I(new_n1953_), .ZN(new_n1965_));
  OAI21_X1   g01773(.A1(new_n1962_), .A2(new_n1964_), .B(new_n1965_), .ZN(new_n1966_));
  OAI21_X1   g01774(.A1(new_n1961_), .A2(new_n1966_), .B(\a[96] ), .ZN(new_n1967_));
  AOI21_X1   g01775(.A1(new_n1967_), .A2(new_n1960_), .B(new_n1806_), .ZN(new_n1968_));
  NOR3_X1    g01776(.A1(new_n1707_), .A2(new_n1710_), .A3(new_n1959_), .ZN(new_n1969_));
  NAND3_X1   g01777(.A1(new_n1698_), .A2(new_n1780_), .A3(new_n1969_), .ZN(new_n1970_));
  INV_X1     g01778(.I(new_n1970_), .ZN(new_n1971_));
  NAND2_X1   g01779(.A1(new_n1967_), .A2(new_n1971_), .ZN(new_n1972_));
  INV_X1     g01780(.I(\a[96] ), .ZN(new_n1973_));
  OAI21_X1   g01781(.A1(new_n1961_), .A2(new_n1966_), .B(new_n1973_), .ZN(new_n1974_));
  AOI22_X1   g01782(.A1(new_n1974_), .A2(\a[97] ), .B1(\asqrt[48] ), .B2(new_n1715_), .ZN(new_n1975_));
  AOI21_X1   g01783(.A1(new_n1975_), .A2(new_n1972_), .B(new_n1968_), .ZN(new_n1976_));
  NOR2_X1    g01784(.A1(new_n1976_), .A2(new_n1612_), .ZN(new_n1977_));
  NAND2_X1   g01785(.A1(new_n1975_), .A2(new_n1972_), .ZN(new_n1978_));
  INV_X1     g01786(.I(new_n1908_), .ZN(new_n1979_));
  INV_X1     g01787(.I(new_n1882_), .ZN(new_n1980_));
  NAND2_X1   g01788(.A1(new_n1861_), .A2(new_n436_), .ZN(new_n1981_));
  OAI21_X1   g01789(.A1(new_n1981_), .A2(new_n1913_), .B(new_n1980_), .ZN(new_n1982_));
  NAND3_X1   g01790(.A1(new_n1982_), .A2(new_n327_), .A3(new_n1914_), .ZN(new_n1983_));
  AOI22_X1   g01791(.A1(new_n1983_), .A2(new_n1909_), .B1(\asqrt[59] ), .B2(new_n1931_), .ZN(new_n1984_));
  OAI21_X1   g01792(.A1(new_n1984_), .A2(new_n306_), .B(new_n218_), .ZN(new_n1985_));
  OAI21_X1   g01793(.A1(new_n1985_), .A2(new_n1933_), .B(new_n1979_), .ZN(new_n1986_));
  NAND3_X1   g01794(.A1(new_n1986_), .A2(new_n207_), .A3(new_n1934_), .ZN(new_n1987_));
  AOI22_X1   g01795(.A1(new_n1987_), .A2(new_n1926_), .B1(new_n1946_), .B2(\asqrt[62] ), .ZN(new_n1988_));
  OAI21_X1   g01796(.A1(new_n1988_), .A2(new_n1943_), .B(new_n193_), .ZN(new_n1989_));
  AOI21_X1   g01797(.A1(new_n1989_), .A2(new_n1954_), .B(new_n1716_), .ZN(new_n1990_));
  NOR2_X1    g01798(.A1(new_n1962_), .A2(new_n1964_), .ZN(new_n1991_));
  OAI21_X1   g01799(.A1(new_n1951_), .A2(new_n1713_), .B(new_n1698_), .ZN(new_n1992_));
  NAND2_X1   g01800(.A1(new_n1949_), .A2(new_n1992_), .ZN(new_n1993_));
  NOR3_X1    g01801(.A1(new_n1961_), .A2(new_n1991_), .A3(new_n1993_), .ZN(new_n1994_));
  OAI21_X1   g01802(.A1(new_n1990_), .A2(new_n1994_), .B(\a[98] ), .ZN(new_n1995_));
  OAI21_X1   g01803(.A1(new_n1961_), .A2(new_n1966_), .B(new_n1715_), .ZN(new_n1996_));
  INV_X1     g01804(.I(new_n1994_), .ZN(new_n1997_));
  NAND3_X1   g01805(.A1(new_n1997_), .A2(new_n1996_), .A3(new_n1768_), .ZN(new_n1998_));
  NOR2_X1    g01806(.A1(new_n1968_), .A2(\asqrt[50] ), .ZN(new_n1999_));
  AOI22_X1   g01807(.A1(new_n1978_), .A2(new_n1999_), .B1(new_n1995_), .B2(new_n1998_), .ZN(new_n2000_));
  OAI21_X1   g01808(.A1(new_n2000_), .A2(new_n1977_), .B(\asqrt[51] ), .ZN(new_n2001_));
  NOR3_X1    g01809(.A1(new_n1829_), .A2(new_n1767_), .A3(new_n1773_), .ZN(new_n2002_));
  NAND3_X1   g01810(.A1(\asqrt[48] ), .A2(new_n1789_), .A3(new_n1809_), .ZN(new_n2003_));
  AOI22_X1   g01811(.A1(new_n2003_), .A2(new_n1829_), .B1(\asqrt[48] ), .B2(new_n2002_), .ZN(new_n2004_));
  INV_X1     g01812(.I(new_n2004_), .ZN(new_n2005_));
  OAI21_X1   g01813(.A1(new_n1976_), .A2(new_n1612_), .B(new_n1376_), .ZN(new_n2006_));
  OAI21_X1   g01814(.A1(new_n2006_), .A2(new_n2000_), .B(new_n2005_), .ZN(new_n2007_));
  AOI21_X1   g01815(.A1(new_n2007_), .A2(new_n2001_), .B(new_n1256_), .ZN(new_n2008_));
  NOR2_X1    g01816(.A1(new_n1788_), .A2(new_n1784_), .ZN(new_n2009_));
  NOR2_X1    g01817(.A1(new_n1777_), .A2(new_n1790_), .ZN(new_n2010_));
  INV_X1     g01818(.I(new_n2010_), .ZN(new_n2011_));
  NAND4_X1   g01819(.A1(\asqrt[48] ), .A2(new_n1778_), .A3(new_n2009_), .A4(new_n2011_), .ZN(new_n2012_));
  NOR3_X1    g01820(.A1(new_n1956_), .A2(new_n1813_), .A3(new_n2010_), .ZN(new_n2013_));
  OAI21_X1   g01821(.A1(new_n2013_), .A2(new_n2009_), .B(new_n2012_), .ZN(new_n2014_));
  INV_X1     g01822(.I(new_n2014_), .ZN(new_n2015_));
  AOI21_X1   g01823(.A1(new_n1989_), .A2(new_n1954_), .B(new_n1973_), .ZN(new_n2016_));
  NOR2_X1    g01824(.A1(new_n2016_), .A2(new_n1970_), .ZN(new_n2017_));
  INV_X1     g01825(.I(\a[97] ), .ZN(new_n2018_));
  AOI21_X1   g01826(.A1(\asqrt[48] ), .A2(new_n1973_), .B(new_n2018_), .ZN(new_n2019_));
  NOR3_X1    g01827(.A1(new_n2017_), .A2(new_n2019_), .A3(new_n1990_), .ZN(new_n2020_));
  OAI21_X1   g01828(.A1(new_n2020_), .A2(new_n1968_), .B(\asqrt[50] ), .ZN(new_n2021_));
  AOI21_X1   g01829(.A1(new_n1997_), .A2(new_n1996_), .B(new_n1768_), .ZN(new_n2022_));
  NOR3_X1    g01830(.A1(new_n1990_), .A2(new_n1994_), .A3(\a[98] ), .ZN(new_n2023_));
  AOI21_X1   g01831(.A1(\asqrt[48] ), .A2(\a[96] ), .B(new_n1959_), .ZN(new_n2024_));
  OAI21_X1   g01832(.A1(new_n2024_), .A2(new_n1806_), .B(new_n1612_), .ZN(new_n2025_));
  OAI22_X1   g01833(.A1(new_n2020_), .A2(new_n2025_), .B1(new_n2022_), .B2(new_n2023_), .ZN(new_n2026_));
  AOI21_X1   g01834(.A1(new_n2026_), .A2(new_n2021_), .B(new_n1376_), .ZN(new_n2027_));
  OAI21_X1   g01835(.A1(new_n2016_), .A2(new_n1959_), .B(\asqrt[49] ), .ZN(new_n2028_));
  AOI21_X1   g01836(.A1(new_n1989_), .A2(new_n1954_), .B(\a[96] ), .ZN(new_n2029_));
  OAI21_X1   g01837(.A1(new_n2018_), .A2(new_n2029_), .B(new_n1996_), .ZN(new_n2030_));
  OAI21_X1   g01838(.A1(new_n2030_), .A2(new_n2017_), .B(new_n2028_), .ZN(new_n2031_));
  AOI21_X1   g01839(.A1(new_n2031_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n2032_));
  AOI21_X1   g01840(.A1(new_n2032_), .A2(new_n2026_), .B(new_n2004_), .ZN(new_n2033_));
  NOR3_X1    g01841(.A1(new_n2033_), .A2(new_n2027_), .A3(\asqrt[52] ), .ZN(new_n2034_));
  NOR2_X1    g01842(.A1(new_n2034_), .A2(new_n2015_), .ZN(new_n2035_));
  OAI21_X1   g01843(.A1(new_n2035_), .A2(new_n2008_), .B(\asqrt[53] ), .ZN(new_n2036_));
  NOR2_X1    g01844(.A1(new_n1831_), .A2(new_n1818_), .ZN(new_n2037_));
  NOR3_X1    g01845(.A1(new_n1956_), .A2(new_n1792_), .A3(new_n2037_), .ZN(new_n2038_));
  INV_X1     g01846(.I(new_n2038_), .ZN(new_n2039_));
  NOR3_X1    g01847(.A1(new_n2037_), .A2(new_n1792_), .A3(new_n1828_), .ZN(new_n2040_));
  AOI22_X1   g01848(.A1(new_n2039_), .A2(new_n1828_), .B1(\asqrt[48] ), .B2(new_n2040_), .ZN(new_n2041_));
  INV_X1     g01849(.I(new_n2041_), .ZN(new_n2042_));
  OAI21_X1   g01850(.A1(new_n2033_), .A2(new_n2027_), .B(\asqrt[52] ), .ZN(new_n2043_));
  NAND2_X1   g01851(.A1(new_n2043_), .A2(new_n1103_), .ZN(new_n2044_));
  OAI21_X1   g01852(.A1(new_n2035_), .A2(new_n2044_), .B(new_n2042_), .ZN(new_n2045_));
  AOI21_X1   g01853(.A1(new_n2045_), .A2(new_n2036_), .B(new_n904_), .ZN(new_n2046_));
  NOR3_X1    g01854(.A1(new_n1842_), .A2(new_n1844_), .A3(new_n1808_), .ZN(new_n2047_));
  NOR3_X1    g01855(.A1(new_n1956_), .A2(new_n1842_), .A3(new_n1844_), .ZN(new_n2048_));
  INV_X1     g01856(.I(new_n2048_), .ZN(new_n2049_));
  AOI22_X1   g01857(.A1(new_n2049_), .A2(new_n1808_), .B1(\asqrt[48] ), .B2(new_n2047_), .ZN(new_n2050_));
  OAI21_X1   g01858(.A1(new_n2015_), .A2(new_n2034_), .B(new_n2043_), .ZN(new_n2051_));
  AOI21_X1   g01859(.A1(new_n2051_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n2052_));
  AOI21_X1   g01860(.A1(new_n2052_), .A2(new_n2045_), .B(new_n2050_), .ZN(new_n2053_));
  OAI21_X1   g01861(.A1(new_n2053_), .A2(new_n2046_), .B(\asqrt[55] ), .ZN(new_n2054_));
  INV_X1     g01862(.I(new_n2054_), .ZN(new_n2055_));
  NOR2_X1    g01863(.A1(new_n1845_), .A2(new_n1856_), .ZN(new_n2056_));
  NOR3_X1    g01864(.A1(new_n1956_), .A2(new_n1822_), .A3(new_n2056_), .ZN(new_n2057_));
  INV_X1     g01865(.I(new_n2057_), .ZN(new_n2058_));
  NOR3_X1    g01866(.A1(new_n2056_), .A2(new_n1822_), .A3(new_n1855_), .ZN(new_n2059_));
  AOI22_X1   g01867(.A1(new_n2058_), .A2(new_n1855_), .B1(\asqrt[48] ), .B2(new_n2059_), .ZN(new_n2060_));
  NOR3_X1    g01868(.A1(new_n2053_), .A2(new_n2046_), .A3(\asqrt[55] ), .ZN(new_n2061_));
  NOR2_X1    g01869(.A1(new_n2061_), .A2(new_n2060_), .ZN(new_n2062_));
  OAI21_X1   g01870(.A1(new_n2062_), .A2(new_n2055_), .B(\asqrt[56] ), .ZN(new_n2063_));
  NOR3_X1    g01871(.A1(new_n1868_), .A2(new_n1910_), .A3(new_n1841_), .ZN(new_n2064_));
  NOR3_X1    g01872(.A1(new_n1956_), .A2(new_n1868_), .A3(new_n1910_), .ZN(new_n2065_));
  INV_X1     g01873(.I(new_n2065_), .ZN(new_n2066_));
  AOI22_X1   g01874(.A1(new_n2066_), .A2(new_n1841_), .B1(\asqrt[48] ), .B2(new_n2064_), .ZN(new_n2067_));
  INV_X1     g01875(.I(new_n2067_), .ZN(new_n2068_));
  NAND2_X1   g01876(.A1(new_n2054_), .A2(new_n703_), .ZN(new_n2069_));
  OAI21_X1   g01877(.A1(new_n2062_), .A2(new_n2069_), .B(new_n2068_), .ZN(new_n2070_));
  AOI21_X1   g01878(.A1(new_n2070_), .A2(new_n2063_), .B(new_n531_), .ZN(new_n2071_));
  NOR3_X1    g01879(.A1(new_n1956_), .A2(new_n1849_), .A3(new_n1927_), .ZN(new_n2072_));
  INV_X1     g01880(.I(new_n2072_), .ZN(new_n2073_));
  NOR3_X1    g01881(.A1(new_n1849_), .A2(new_n1873_), .A3(new_n1927_), .ZN(new_n2074_));
  AOI22_X1   g01882(.A1(new_n2073_), .A2(new_n1873_), .B1(\asqrt[48] ), .B2(new_n2074_), .ZN(new_n2075_));
  OAI21_X1   g01883(.A1(new_n2060_), .A2(new_n2061_), .B(new_n2054_), .ZN(new_n2076_));
  AOI21_X1   g01884(.A1(new_n2076_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n2077_));
  AOI21_X1   g01885(.A1(new_n2077_), .A2(new_n2070_), .B(new_n2075_), .ZN(new_n2078_));
  OAI21_X1   g01886(.A1(new_n2078_), .A2(new_n2071_), .B(\asqrt[58] ), .ZN(new_n2079_));
  AND3_X2    g01887(.A1(new_n1861_), .A2(new_n1866_), .A3(new_n1876_), .Z(new_n2080_));
  NAND3_X1   g01888(.A1(\asqrt[48] ), .A2(new_n1861_), .A3(new_n1876_), .ZN(new_n2081_));
  AOI22_X1   g01889(.A1(new_n2081_), .A2(new_n1867_), .B1(\asqrt[48] ), .B2(new_n2080_), .ZN(new_n2082_));
  INV_X1     g01890(.I(new_n2082_), .ZN(new_n2083_));
  INV_X1     g01891(.I(new_n2060_), .ZN(new_n2084_));
  NAND2_X1   g01892(.A1(new_n2001_), .A2(new_n1256_), .ZN(new_n2085_));
  OAI21_X1   g01893(.A1(new_n2085_), .A2(new_n2033_), .B(new_n2014_), .ZN(new_n2086_));
  AOI21_X1   g01894(.A1(new_n2086_), .A2(new_n2043_), .B(new_n1103_), .ZN(new_n2087_));
  NOR2_X1    g01895(.A1(new_n2008_), .A2(\asqrt[53] ), .ZN(new_n2088_));
  AOI21_X1   g01896(.A1(new_n2088_), .A2(new_n2086_), .B(new_n2041_), .ZN(new_n2089_));
  OAI21_X1   g01897(.A1(new_n2089_), .A2(new_n2087_), .B(\asqrt[54] ), .ZN(new_n2090_));
  NAND2_X1   g01898(.A1(new_n2090_), .A2(new_n823_), .ZN(new_n2091_));
  OAI21_X1   g01899(.A1(new_n2091_), .A2(new_n2053_), .B(new_n2084_), .ZN(new_n2092_));
  NAND3_X1   g01900(.A1(new_n2092_), .A2(new_n703_), .A3(new_n2054_), .ZN(new_n2093_));
  AOI22_X1   g01901(.A1(new_n2093_), .A2(new_n2068_), .B1(new_n2076_), .B2(\asqrt[56] ), .ZN(new_n2094_));
  OAI21_X1   g01902(.A1(new_n2094_), .A2(new_n531_), .B(new_n436_), .ZN(new_n2095_));
  OAI21_X1   g01903(.A1(new_n2095_), .A2(new_n2078_), .B(new_n2083_), .ZN(new_n2096_));
  AOI21_X1   g01904(.A1(new_n2096_), .A2(new_n2079_), .B(new_n327_), .ZN(new_n2097_));
  NOR3_X1    g01905(.A1(new_n1956_), .A2(new_n1878_), .A3(new_n1930_), .ZN(new_n2098_));
  INV_X1     g01906(.I(new_n2098_), .ZN(new_n2099_));
  NOR3_X1    g01907(.A1(new_n1878_), .A2(new_n1980_), .A3(new_n1930_), .ZN(new_n2100_));
  AOI22_X1   g01908(.A1(new_n2099_), .A2(new_n1980_), .B1(\asqrt[48] ), .B2(new_n2100_), .ZN(new_n2101_));
  INV_X1     g01909(.I(new_n2071_), .ZN(new_n2102_));
  INV_X1     g01910(.I(new_n2070_), .ZN(new_n2103_));
  INV_X1     g01911(.I(new_n2075_), .ZN(new_n2104_));
  NAND2_X1   g01912(.A1(new_n2063_), .A2(new_n531_), .ZN(new_n2105_));
  OAI21_X1   g01913(.A1(new_n2105_), .A2(new_n2103_), .B(new_n2104_), .ZN(new_n2106_));
  AOI21_X1   g01914(.A1(new_n2106_), .A2(new_n2102_), .B(new_n436_), .ZN(new_n2107_));
  NOR2_X1    g01915(.A1(new_n2107_), .A2(\asqrt[59] ), .ZN(new_n2108_));
  AOI21_X1   g01916(.A1(new_n2108_), .A2(new_n2096_), .B(new_n2101_), .ZN(new_n2109_));
  OAI21_X1   g01917(.A1(new_n2109_), .A2(new_n2097_), .B(\asqrt[60] ), .ZN(new_n2110_));
  NOR3_X1    g01918(.A1(new_n1887_), .A2(new_n1893_), .A3(new_n1909_), .ZN(new_n2111_));
  NOR3_X1    g01919(.A1(new_n1956_), .A2(new_n1887_), .A3(new_n1893_), .ZN(new_n2112_));
  INV_X1     g01920(.I(new_n2112_), .ZN(new_n2113_));
  AOI22_X1   g01921(.A1(new_n2113_), .A2(new_n1909_), .B1(\asqrt[48] ), .B2(new_n2111_), .ZN(new_n2114_));
  INV_X1     g01922(.I(new_n2114_), .ZN(new_n2115_));
  NOR2_X1    g01923(.A1(new_n2071_), .A2(\asqrt[58] ), .ZN(new_n2116_));
  AOI21_X1   g01924(.A1(new_n2116_), .A2(new_n2106_), .B(new_n2082_), .ZN(new_n2117_));
  OAI21_X1   g01925(.A1(new_n2117_), .A2(new_n2107_), .B(\asqrt[59] ), .ZN(new_n2118_));
  NAND2_X1   g01926(.A1(new_n2118_), .A2(new_n306_), .ZN(new_n2119_));
  OAI21_X1   g01927(.A1(new_n2119_), .A2(new_n2109_), .B(new_n2115_), .ZN(new_n2120_));
  AOI21_X1   g01928(.A1(new_n2120_), .A2(new_n2110_), .B(new_n218_), .ZN(new_n2121_));
  NOR2_X1    g01929(.A1(new_n1894_), .A2(new_n1902_), .ZN(new_n2122_));
  NOR3_X1    g01930(.A1(new_n1956_), .A2(new_n1917_), .A3(new_n2122_), .ZN(new_n2123_));
  INV_X1     g01931(.I(new_n2123_), .ZN(new_n2124_));
  NOR3_X1    g01932(.A1(new_n2122_), .A2(new_n1917_), .A3(new_n1901_), .ZN(new_n2125_));
  AOI22_X1   g01933(.A1(new_n2124_), .A2(new_n1901_), .B1(\asqrt[48] ), .B2(new_n2125_), .ZN(new_n2126_));
  INV_X1     g01934(.I(new_n2101_), .ZN(new_n2127_));
  NAND2_X1   g01935(.A1(new_n2079_), .A2(new_n327_), .ZN(new_n2128_));
  OAI21_X1   g01936(.A1(new_n2128_), .A2(new_n2117_), .B(new_n2127_), .ZN(new_n2129_));
  AOI21_X1   g01937(.A1(new_n2129_), .A2(new_n2118_), .B(new_n306_), .ZN(new_n2130_));
  NOR2_X1    g01938(.A1(new_n2130_), .A2(\asqrt[61] ), .ZN(new_n2131_));
  AOI21_X1   g01939(.A1(new_n2131_), .A2(new_n2120_), .B(new_n2126_), .ZN(new_n2132_));
  OAI21_X1   g01940(.A1(new_n2132_), .A2(new_n2121_), .B(\asqrt[62] ), .ZN(new_n2133_));
  NOR3_X1    g01941(.A1(new_n1904_), .A2(new_n1979_), .A3(new_n1945_), .ZN(new_n2134_));
  NOR3_X1    g01942(.A1(new_n1956_), .A2(new_n1904_), .A3(new_n1945_), .ZN(new_n2135_));
  INV_X1     g01943(.I(new_n2135_), .ZN(new_n2136_));
  AOI22_X1   g01944(.A1(new_n2136_), .A2(new_n1979_), .B1(\asqrt[48] ), .B2(new_n2134_), .ZN(new_n2137_));
  INV_X1     g01945(.I(new_n2137_), .ZN(new_n2138_));
  NOR3_X1    g01946(.A1(new_n2078_), .A2(new_n2071_), .A3(\asqrt[58] ), .ZN(new_n2139_));
  OAI21_X1   g01947(.A1(new_n2082_), .A2(new_n2139_), .B(new_n2079_), .ZN(new_n2140_));
  AOI21_X1   g01948(.A1(new_n2140_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n2141_));
  AOI21_X1   g01949(.A1(new_n2141_), .A2(new_n2129_), .B(new_n2114_), .ZN(new_n2142_));
  OAI21_X1   g01950(.A1(new_n2142_), .A2(new_n2130_), .B(\asqrt[61] ), .ZN(new_n2143_));
  NAND2_X1   g01951(.A1(new_n2143_), .A2(new_n207_), .ZN(new_n2144_));
  OAI21_X1   g01952(.A1(new_n2144_), .A2(new_n2132_), .B(new_n2138_), .ZN(new_n2145_));
  INV_X1     g01953(.I(new_n1991_), .ZN(new_n2146_));
  NAND4_X1   g01954(.A1(\asqrt[48] ), .A2(new_n1920_), .A3(new_n1925_), .A4(new_n1987_), .ZN(new_n2147_));
  NAND2_X1   g01955(.A1(new_n1987_), .A2(new_n1920_), .ZN(new_n2148_));
  OAI21_X1   g01956(.A1(new_n1956_), .A2(new_n2148_), .B(new_n1926_), .ZN(new_n2149_));
  NAND2_X1   g01957(.A1(new_n2149_), .A2(new_n2147_), .ZN(new_n2150_));
  NOR2_X1    g01958(.A1(new_n1988_), .A2(new_n1963_), .ZN(new_n2151_));
  NAND2_X1   g01959(.A1(\asqrt[48] ), .A2(new_n2151_), .ZN(new_n2152_));
  NAND3_X1   g01960(.A1(new_n2150_), .A2(new_n2146_), .A3(new_n2152_), .ZN(new_n2153_));
  AOI21_X1   g01961(.A1(new_n2145_), .A2(new_n2133_), .B(new_n2153_), .ZN(new_n2154_));
  NOR3_X1    g01962(.A1(new_n2142_), .A2(\asqrt[61] ), .A3(new_n2130_), .ZN(new_n2155_));
  OAI21_X1   g01963(.A1(new_n2126_), .A2(new_n2155_), .B(new_n2143_), .ZN(new_n2156_));
  AOI21_X1   g01964(.A1(new_n2156_), .A2(\asqrt[62] ), .B(new_n2150_), .ZN(new_n2157_));
  OAI21_X1   g01965(.A1(new_n1956_), .A2(new_n1963_), .B(new_n1988_), .ZN(new_n2158_));
  NOR2_X1    g01966(.A1(new_n2151_), .A2(new_n193_), .ZN(new_n2159_));
  NAND2_X1   g01967(.A1(new_n2158_), .A2(new_n2159_), .ZN(new_n2160_));
  INV_X1     g01968(.I(new_n2160_), .ZN(new_n2161_));
  AND3_X2    g01969(.A1(new_n1939_), .A2(new_n1937_), .A3(new_n1952_), .Z(new_n2162_));
  NAND4_X1   g01970(.A1(new_n2146_), .A2(new_n1989_), .A3(new_n1949_), .A4(new_n2162_), .ZN(new_n2163_));
  INV_X1     g01971(.I(new_n2163_), .ZN(new_n2164_));
  NOR2_X1    g01972(.A1(new_n2161_), .A2(new_n2164_), .ZN(new_n2165_));
  INV_X1     g01973(.I(new_n2165_), .ZN(new_n2166_));
  AOI21_X1   g01974(.A1(new_n2157_), .A2(new_n2145_), .B(new_n2166_), .ZN(new_n2167_));
  OAI21_X1   g01975(.A1(\asqrt[63] ), .A2(new_n2154_), .B(new_n2167_), .ZN(\asqrt[47] ));
  NOR2_X1    g01976(.A1(\a[92] ), .A2(\a[93] ), .ZN(new_n2169_));
  INV_X1     g01977(.I(new_n2169_), .ZN(new_n2170_));
  NOR2_X1    g01978(.A1(new_n2170_), .A2(\a[94] ), .ZN(new_n2171_));
  INV_X1     g01979(.I(new_n2171_), .ZN(new_n2172_));
  NAND2_X1   g01980(.A1(new_n2145_), .A2(new_n2133_), .ZN(new_n2173_));
  INV_X1     g01981(.I(new_n2153_), .ZN(new_n2174_));
  AOI21_X1   g01982(.A1(new_n2173_), .A2(new_n2174_), .B(\asqrt[63] ), .ZN(new_n2175_));
  INV_X1     g01983(.I(new_n2145_), .ZN(new_n2176_));
  INV_X1     g01984(.I(new_n2150_), .ZN(new_n2177_));
  NAND2_X1   g01985(.A1(new_n2133_), .A2(new_n2177_), .ZN(new_n2178_));
  OAI21_X1   g01986(.A1(new_n2176_), .A2(new_n2178_), .B(new_n2165_), .ZN(new_n2179_));
  OAI21_X1   g01987(.A1(new_n2175_), .A2(new_n2179_), .B(\a[94] ), .ZN(new_n2180_));
  AOI21_X1   g01988(.A1(new_n2180_), .A2(new_n2172_), .B(new_n1956_), .ZN(new_n2181_));
  INV_X1     g01989(.I(\a[94] ), .ZN(new_n2182_));
  INV_X1     g01990(.I(new_n2126_), .ZN(new_n2183_));
  NAND3_X1   g01991(.A1(new_n2096_), .A2(new_n327_), .A3(new_n2079_), .ZN(new_n2184_));
  AOI21_X1   g01992(.A1(new_n2127_), .A2(new_n2184_), .B(new_n2097_), .ZN(new_n2185_));
  OAI21_X1   g01993(.A1(new_n2185_), .A2(new_n306_), .B(new_n218_), .ZN(new_n2186_));
  OAI21_X1   g01994(.A1(new_n2186_), .A2(new_n2142_), .B(new_n2183_), .ZN(new_n2187_));
  NAND3_X1   g01995(.A1(new_n2187_), .A2(new_n207_), .A3(new_n2143_), .ZN(new_n2188_));
  AOI22_X1   g01996(.A1(new_n2188_), .A2(new_n2138_), .B1(new_n2156_), .B2(\asqrt[62] ), .ZN(new_n2189_));
  OAI21_X1   g01997(.A1(new_n2189_), .A2(new_n2153_), .B(new_n193_), .ZN(new_n2190_));
  AOI21_X1   g01998(.A1(new_n2190_), .A2(new_n2167_), .B(new_n2182_), .ZN(new_n2191_));
  NAND4_X1   g01999(.A1(new_n2146_), .A2(new_n1949_), .A3(new_n1952_), .A4(new_n2172_), .ZN(new_n2192_));
  NOR2_X1    g02000(.A1(new_n2192_), .A2(new_n1961_), .ZN(new_n2193_));
  INV_X1     g02001(.I(new_n2193_), .ZN(new_n2194_));
  NOR2_X1    g02002(.A1(new_n2191_), .A2(new_n2194_), .ZN(new_n2195_));
  AOI21_X1   g02003(.A1(new_n2190_), .A2(new_n2167_), .B(new_n1958_), .ZN(new_n2196_));
  INV_X1     g02004(.I(\a[95] ), .ZN(new_n2197_));
  AOI21_X1   g02005(.A1(\asqrt[47] ), .A2(new_n2182_), .B(new_n2197_), .ZN(new_n2198_));
  NOR3_X1    g02006(.A1(new_n2195_), .A2(new_n2198_), .A3(new_n2196_), .ZN(new_n2199_));
  OAI21_X1   g02007(.A1(new_n2199_), .A2(new_n2181_), .B(\asqrt[49] ), .ZN(new_n2200_));
  OAI21_X1   g02008(.A1(new_n2175_), .A2(new_n2179_), .B(new_n1957_), .ZN(new_n2201_));
  NOR2_X1    g02009(.A1(new_n2176_), .A2(new_n2178_), .ZN(new_n2202_));
  INV_X1     g02010(.I(new_n2202_), .ZN(new_n2203_));
  NOR2_X1    g02011(.A1(new_n2164_), .A2(new_n1956_), .ZN(new_n2204_));
  NAND4_X1   g02012(.A1(new_n2203_), .A2(new_n2190_), .A3(new_n2160_), .A4(new_n2204_), .ZN(new_n2205_));
  AOI21_X1   g02013(.A1(new_n2205_), .A2(new_n2201_), .B(new_n1973_), .ZN(new_n2206_));
  INV_X1     g02014(.I(new_n2204_), .ZN(new_n2207_));
  NOR4_X1    g02015(.A1(new_n2175_), .A2(new_n2202_), .A3(new_n2161_), .A4(new_n2207_), .ZN(new_n2208_));
  NOR3_X1    g02016(.A1(new_n2208_), .A2(new_n2196_), .A3(\a[96] ), .ZN(new_n2209_));
  AOI21_X1   g02017(.A1(\asqrt[47] ), .A2(\a[94] ), .B(new_n2171_), .ZN(new_n2210_));
  OAI21_X1   g02018(.A1(new_n2210_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n2211_));
  OAI22_X1   g02019(.A1(new_n2199_), .A2(new_n2211_), .B1(new_n2206_), .B2(new_n2209_), .ZN(new_n2212_));
  AOI21_X1   g02020(.A1(new_n2212_), .A2(new_n2200_), .B(new_n1612_), .ZN(new_n2213_));
  NOR3_X1    g02021(.A1(new_n1975_), .A2(new_n1968_), .A3(new_n2017_), .ZN(new_n2214_));
  NAND3_X1   g02022(.A1(\asqrt[47] ), .A2(new_n2028_), .A3(new_n1972_), .ZN(new_n2215_));
  AOI22_X1   g02023(.A1(new_n2215_), .A2(new_n1975_), .B1(\asqrt[47] ), .B2(new_n2214_), .ZN(new_n2216_));
  OAI21_X1   g02024(.A1(new_n2191_), .A2(new_n2171_), .B(\asqrt[48] ), .ZN(new_n2217_));
  AOI21_X1   g02025(.A1(new_n2190_), .A2(new_n2167_), .B(\a[94] ), .ZN(new_n2218_));
  OAI21_X1   g02026(.A1(new_n2197_), .A2(new_n2218_), .B(new_n2201_), .ZN(new_n2219_));
  OAI21_X1   g02027(.A1(new_n2219_), .A2(new_n2195_), .B(new_n2217_), .ZN(new_n2220_));
  AOI21_X1   g02028(.A1(new_n2220_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n2221_));
  AOI21_X1   g02029(.A1(new_n2221_), .A2(new_n2212_), .B(new_n2216_), .ZN(new_n2222_));
  OAI21_X1   g02030(.A1(new_n2222_), .A2(new_n2213_), .B(\asqrt[51] ), .ZN(new_n2223_));
  INV_X1     g02031(.I(new_n2223_), .ZN(new_n2224_));
  NOR2_X1    g02032(.A1(new_n2022_), .A2(new_n2023_), .ZN(new_n2225_));
  NOR2_X1    g02033(.A1(new_n2020_), .A2(new_n2025_), .ZN(new_n2226_));
  INV_X1     g02034(.I(new_n2226_), .ZN(new_n2227_));
  NAND4_X1   g02035(.A1(\asqrt[47] ), .A2(new_n2021_), .A3(new_n2225_), .A4(new_n2227_), .ZN(new_n2228_));
  INV_X1     g02036(.I(\asqrt[47] ), .ZN(new_n2229_));
  NOR3_X1    g02037(.A1(new_n2229_), .A2(new_n1977_), .A3(new_n2226_), .ZN(new_n2230_));
  OAI21_X1   g02038(.A1(new_n2230_), .A2(new_n2225_), .B(new_n2228_), .ZN(new_n2231_));
  INV_X1     g02039(.I(new_n2231_), .ZN(new_n2232_));
  NOR3_X1    g02040(.A1(new_n2222_), .A2(new_n2213_), .A3(\asqrt[51] ), .ZN(new_n2233_));
  NOR2_X1    g02041(.A1(new_n2233_), .A2(new_n2232_), .ZN(new_n2234_));
  OAI21_X1   g02042(.A1(new_n2234_), .A2(new_n2224_), .B(\asqrt[52] ), .ZN(new_n2235_));
  NOR2_X1    g02043(.A1(new_n2006_), .A2(new_n2000_), .ZN(new_n2236_));
  NOR3_X1    g02044(.A1(new_n2229_), .A2(new_n2027_), .A3(new_n2236_), .ZN(new_n2237_));
  INV_X1     g02045(.I(new_n2237_), .ZN(new_n2238_));
  NOR3_X1    g02046(.A1(new_n2236_), .A2(new_n2027_), .A3(new_n2005_), .ZN(new_n2239_));
  AOI22_X1   g02047(.A1(new_n2238_), .A2(new_n2005_), .B1(\asqrt[47] ), .B2(new_n2239_), .ZN(new_n2240_));
  INV_X1     g02048(.I(new_n2240_), .ZN(new_n2241_));
  NAND2_X1   g02049(.A1(new_n2223_), .A2(new_n1256_), .ZN(new_n2242_));
  OAI21_X1   g02050(.A1(new_n2234_), .A2(new_n2242_), .B(new_n2241_), .ZN(new_n2243_));
  AOI21_X1   g02051(.A1(new_n2243_), .A2(new_n2235_), .B(new_n1103_), .ZN(new_n2244_));
  NOR3_X1    g02052(.A1(new_n2008_), .A2(new_n2034_), .A3(new_n2014_), .ZN(new_n2245_));
  NOR3_X1    g02053(.A1(new_n2229_), .A2(new_n2008_), .A3(new_n2034_), .ZN(new_n2246_));
  INV_X1     g02054(.I(new_n2246_), .ZN(new_n2247_));
  AOI22_X1   g02055(.A1(new_n2247_), .A2(new_n2014_), .B1(\asqrt[47] ), .B2(new_n2245_), .ZN(new_n2248_));
  OAI21_X1   g02056(.A1(new_n2232_), .A2(new_n2233_), .B(new_n2223_), .ZN(new_n2249_));
  AOI21_X1   g02057(.A1(new_n2249_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n2250_));
  AOI21_X1   g02058(.A1(new_n2250_), .A2(new_n2243_), .B(new_n2248_), .ZN(new_n2251_));
  OAI21_X1   g02059(.A1(new_n2251_), .A2(new_n2244_), .B(\asqrt[54] ), .ZN(new_n2252_));
  INV_X1     g02060(.I(new_n2252_), .ZN(new_n2253_));
  NOR2_X1    g02061(.A1(new_n2035_), .A2(new_n2044_), .ZN(new_n2254_));
  NOR3_X1    g02062(.A1(new_n2229_), .A2(new_n2087_), .A3(new_n2254_), .ZN(new_n2255_));
  INV_X1     g02063(.I(new_n2255_), .ZN(new_n2256_));
  NOR3_X1    g02064(.A1(new_n2254_), .A2(new_n2087_), .A3(new_n2042_), .ZN(new_n2257_));
  AOI22_X1   g02065(.A1(new_n2256_), .A2(new_n2042_), .B1(\asqrt[47] ), .B2(new_n2257_), .ZN(new_n2258_));
  NOR3_X1    g02066(.A1(new_n2251_), .A2(new_n2244_), .A3(\asqrt[54] ), .ZN(new_n2259_));
  NOR2_X1    g02067(.A1(new_n2259_), .A2(new_n2258_), .ZN(new_n2260_));
  OAI21_X1   g02068(.A1(new_n2260_), .A2(new_n2253_), .B(\asqrt[55] ), .ZN(new_n2261_));
  INV_X1     g02069(.I(new_n2050_), .ZN(new_n2262_));
  INV_X1     g02070(.I(new_n2052_), .ZN(new_n2263_));
  NOR2_X1    g02071(.A1(new_n2263_), .A2(new_n2089_), .ZN(new_n2264_));
  NOR3_X1    g02072(.A1(new_n2264_), .A2(new_n2046_), .A3(new_n2262_), .ZN(new_n2265_));
  NOR3_X1    g02073(.A1(new_n2229_), .A2(new_n2046_), .A3(new_n2264_), .ZN(new_n2266_));
  INV_X1     g02074(.I(new_n2266_), .ZN(new_n2267_));
  AOI22_X1   g02075(.A1(new_n2267_), .A2(new_n2262_), .B1(\asqrt[47] ), .B2(new_n2265_), .ZN(new_n2268_));
  INV_X1     g02076(.I(new_n2268_), .ZN(new_n2269_));
  NAND2_X1   g02077(.A1(new_n2252_), .A2(new_n823_), .ZN(new_n2270_));
  OAI21_X1   g02078(.A1(new_n2260_), .A2(new_n2270_), .B(new_n2269_), .ZN(new_n2271_));
  AOI21_X1   g02079(.A1(new_n2271_), .A2(new_n2261_), .B(new_n703_), .ZN(new_n2272_));
  NOR3_X1    g02080(.A1(new_n2229_), .A2(new_n2055_), .A3(new_n2061_), .ZN(new_n2273_));
  INV_X1     g02081(.I(new_n2273_), .ZN(new_n2274_));
  NOR3_X1    g02082(.A1(new_n2055_), .A2(new_n2084_), .A3(new_n2061_), .ZN(new_n2275_));
  AOI22_X1   g02083(.A1(new_n2274_), .A2(new_n2084_), .B1(\asqrt[47] ), .B2(new_n2275_), .ZN(new_n2276_));
  OAI21_X1   g02084(.A1(new_n2258_), .A2(new_n2259_), .B(new_n2252_), .ZN(new_n2277_));
  AOI21_X1   g02085(.A1(new_n2277_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n2278_));
  AOI21_X1   g02086(.A1(new_n2278_), .A2(new_n2271_), .B(new_n2276_), .ZN(new_n2279_));
  OAI21_X1   g02087(.A1(new_n2279_), .A2(new_n2272_), .B(\asqrt[57] ), .ZN(new_n2280_));
  AND3_X2    g02088(.A1(new_n2063_), .A2(new_n2067_), .A3(new_n2093_), .Z(new_n2281_));
  NAND3_X1   g02089(.A1(\asqrt[47] ), .A2(new_n2063_), .A3(new_n2093_), .ZN(new_n2282_));
  AOI22_X1   g02090(.A1(new_n2282_), .A2(new_n2068_), .B1(\asqrt[47] ), .B2(new_n2281_), .ZN(new_n2283_));
  INV_X1     g02091(.I(new_n2283_), .ZN(new_n2284_));
  INV_X1     g02092(.I(new_n2258_), .ZN(new_n2285_));
  NAND2_X1   g02093(.A1(new_n2180_), .A2(new_n2193_), .ZN(new_n2286_));
  OAI21_X1   g02094(.A1(new_n2175_), .A2(new_n2179_), .B(new_n2182_), .ZN(new_n2287_));
  NAND2_X1   g02095(.A1(new_n2287_), .A2(\a[95] ), .ZN(new_n2288_));
  NAND3_X1   g02096(.A1(new_n2286_), .A2(new_n2288_), .A3(new_n2201_), .ZN(new_n2289_));
  AOI21_X1   g02097(.A1(new_n2289_), .A2(new_n2217_), .B(new_n1806_), .ZN(new_n2290_));
  OAI21_X1   g02098(.A1(new_n2208_), .A2(new_n2196_), .B(\a[96] ), .ZN(new_n2291_));
  NAND3_X1   g02099(.A1(new_n2205_), .A2(new_n2201_), .A3(new_n1973_), .ZN(new_n2292_));
  NAND2_X1   g02100(.A1(new_n2180_), .A2(new_n2172_), .ZN(new_n2293_));
  AOI21_X1   g02101(.A1(new_n2293_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n2294_));
  AOI22_X1   g02102(.A1(new_n2289_), .A2(new_n2294_), .B1(new_n2291_), .B2(new_n2292_), .ZN(new_n2295_));
  OAI21_X1   g02103(.A1(new_n2295_), .A2(new_n2290_), .B(\asqrt[50] ), .ZN(new_n2296_));
  NAND2_X1   g02104(.A1(new_n2296_), .A2(new_n1376_), .ZN(new_n2297_));
  OAI21_X1   g02105(.A1(new_n2297_), .A2(new_n2222_), .B(new_n2231_), .ZN(new_n2298_));
  AOI21_X1   g02106(.A1(new_n2298_), .A2(new_n2223_), .B(new_n1256_), .ZN(new_n2299_));
  INV_X1     g02107(.I(new_n2216_), .ZN(new_n2300_));
  AOI21_X1   g02108(.A1(\a[95] ), .A2(new_n2287_), .B(new_n2196_), .ZN(new_n2301_));
  AOI21_X1   g02109(.A1(new_n2301_), .A2(new_n2286_), .B(new_n2181_), .ZN(new_n2302_));
  OAI21_X1   g02110(.A1(new_n2302_), .A2(new_n1806_), .B(new_n1612_), .ZN(new_n2303_));
  OAI21_X1   g02111(.A1(new_n2303_), .A2(new_n2295_), .B(new_n2300_), .ZN(new_n2304_));
  NAND2_X1   g02112(.A1(new_n2304_), .A2(new_n2296_), .ZN(new_n2305_));
  AOI21_X1   g02113(.A1(new_n2305_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n2306_));
  AOI21_X1   g02114(.A1(new_n2306_), .A2(new_n2298_), .B(new_n2240_), .ZN(new_n2307_));
  OAI21_X1   g02115(.A1(new_n2307_), .A2(new_n2299_), .B(\asqrt[53] ), .ZN(new_n2308_));
  NAND2_X1   g02116(.A1(new_n2308_), .A2(new_n904_), .ZN(new_n2309_));
  OAI21_X1   g02117(.A1(new_n2309_), .A2(new_n2251_), .B(new_n2285_), .ZN(new_n2310_));
  NAND3_X1   g02118(.A1(new_n2310_), .A2(new_n823_), .A3(new_n2252_), .ZN(new_n2311_));
  AOI22_X1   g02119(.A1(new_n2311_), .A2(new_n2269_), .B1(new_n2277_), .B2(\asqrt[55] ), .ZN(new_n2312_));
  OAI21_X1   g02120(.A1(new_n2312_), .A2(new_n703_), .B(new_n531_), .ZN(new_n2313_));
  OAI21_X1   g02121(.A1(new_n2313_), .A2(new_n2279_), .B(new_n2284_), .ZN(new_n2314_));
  AOI21_X1   g02122(.A1(new_n2314_), .A2(new_n2280_), .B(new_n436_), .ZN(new_n2315_));
  NOR2_X1    g02123(.A1(new_n2105_), .A2(new_n2103_), .ZN(new_n2316_));
  NOR3_X1    g02124(.A1(new_n2229_), .A2(new_n2071_), .A3(new_n2316_), .ZN(new_n2317_));
  INV_X1     g02125(.I(new_n2317_), .ZN(new_n2318_));
  NOR3_X1    g02126(.A1(new_n2316_), .A2(new_n2071_), .A3(new_n2104_), .ZN(new_n2319_));
  AOI22_X1   g02127(.A1(new_n2318_), .A2(new_n2104_), .B1(\asqrt[47] ), .B2(new_n2319_), .ZN(new_n2320_));
  AOI21_X1   g02128(.A1(new_n2310_), .A2(new_n2252_), .B(new_n823_), .ZN(new_n2321_));
  NOR3_X1    g02129(.A1(new_n2307_), .A2(new_n2299_), .A3(\asqrt[53] ), .ZN(new_n2322_));
  OAI21_X1   g02130(.A1(new_n2248_), .A2(new_n2322_), .B(new_n2308_), .ZN(new_n2323_));
  AOI21_X1   g02131(.A1(new_n2323_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n2324_));
  AOI21_X1   g02132(.A1(new_n2324_), .A2(new_n2310_), .B(new_n2268_), .ZN(new_n2325_));
  NOR3_X1    g02133(.A1(new_n2325_), .A2(\asqrt[56] ), .A3(new_n2321_), .ZN(new_n2326_));
  OAI22_X1   g02134(.A1(new_n2326_), .A2(new_n2276_), .B1(new_n2312_), .B2(new_n703_), .ZN(new_n2327_));
  AOI21_X1   g02135(.A1(new_n2327_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n2328_));
  AOI21_X1   g02136(.A1(new_n2328_), .A2(new_n2314_), .B(new_n2320_), .ZN(new_n2329_));
  OAI21_X1   g02137(.A1(new_n2329_), .A2(new_n2315_), .B(\asqrt[59] ), .ZN(new_n2330_));
  NOR3_X1    g02138(.A1(new_n2107_), .A2(new_n2139_), .A3(new_n2083_), .ZN(new_n2331_));
  NOR3_X1    g02139(.A1(new_n2229_), .A2(new_n2107_), .A3(new_n2139_), .ZN(new_n2332_));
  INV_X1     g02140(.I(new_n2332_), .ZN(new_n2333_));
  AOI22_X1   g02141(.A1(new_n2333_), .A2(new_n2083_), .B1(\asqrt[47] ), .B2(new_n2331_), .ZN(new_n2334_));
  INV_X1     g02142(.I(new_n2334_), .ZN(new_n2335_));
  INV_X1     g02143(.I(new_n2280_), .ZN(new_n2336_));
  INV_X1     g02144(.I(new_n2276_), .ZN(new_n2337_));
  NAND2_X1   g02145(.A1(new_n2261_), .A2(new_n703_), .ZN(new_n2338_));
  OAI21_X1   g02146(.A1(new_n2338_), .A2(new_n2325_), .B(new_n2337_), .ZN(new_n2339_));
  NOR2_X1    g02147(.A1(new_n2272_), .A2(\asqrt[57] ), .ZN(new_n2340_));
  AOI21_X1   g02148(.A1(new_n2340_), .A2(new_n2339_), .B(new_n2283_), .ZN(new_n2341_));
  OAI21_X1   g02149(.A1(new_n2336_), .A2(new_n2341_), .B(\asqrt[58] ), .ZN(new_n2342_));
  NAND2_X1   g02150(.A1(new_n2342_), .A2(new_n327_), .ZN(new_n2343_));
  OAI21_X1   g02151(.A1(new_n2343_), .A2(new_n2329_), .B(new_n2335_), .ZN(new_n2344_));
  AOI21_X1   g02152(.A1(new_n2344_), .A2(new_n2330_), .B(new_n306_), .ZN(new_n2345_));
  INV_X1     g02153(.I(new_n2184_), .ZN(new_n2346_));
  NOR3_X1    g02154(.A1(new_n2229_), .A2(new_n2097_), .A3(new_n2346_), .ZN(new_n2347_));
  INV_X1     g02155(.I(new_n2347_), .ZN(new_n2348_));
  NOR3_X1    g02156(.A1(new_n2346_), .A2(new_n2097_), .A3(new_n2127_), .ZN(new_n2349_));
  AOI22_X1   g02157(.A1(new_n2348_), .A2(new_n2127_), .B1(\asqrt[47] ), .B2(new_n2349_), .ZN(new_n2350_));
  INV_X1     g02158(.I(new_n2320_), .ZN(new_n2351_));
  NAND2_X1   g02159(.A1(new_n2280_), .A2(new_n436_), .ZN(new_n2352_));
  OAI21_X1   g02160(.A1(new_n2352_), .A2(new_n2341_), .B(new_n2351_), .ZN(new_n2353_));
  AOI21_X1   g02161(.A1(new_n2353_), .A2(new_n2342_), .B(new_n327_), .ZN(new_n2354_));
  NOR2_X1    g02162(.A1(new_n2354_), .A2(\asqrt[60] ), .ZN(new_n2355_));
  AOI21_X1   g02163(.A1(new_n2355_), .A2(new_n2344_), .B(new_n2350_), .ZN(new_n2356_));
  OAI21_X1   g02164(.A1(new_n2356_), .A2(new_n2345_), .B(\asqrt[61] ), .ZN(new_n2357_));
  NOR2_X1    g02165(.A1(new_n2119_), .A2(new_n2109_), .ZN(new_n2358_));
  NOR3_X1    g02166(.A1(new_n2358_), .A2(new_n2130_), .A3(new_n2115_), .ZN(new_n2359_));
  NOR3_X1    g02167(.A1(new_n2229_), .A2(new_n2130_), .A3(new_n2358_), .ZN(new_n2360_));
  INV_X1     g02168(.I(new_n2360_), .ZN(new_n2361_));
  AOI22_X1   g02169(.A1(new_n2361_), .A2(new_n2115_), .B1(\asqrt[47] ), .B2(new_n2359_), .ZN(new_n2362_));
  INV_X1     g02170(.I(new_n2362_), .ZN(new_n2363_));
  NOR3_X1    g02171(.A1(new_n2279_), .A2(new_n2272_), .A3(\asqrt[57] ), .ZN(new_n2364_));
  OAI21_X1   g02172(.A1(new_n2283_), .A2(new_n2364_), .B(new_n2280_), .ZN(new_n2365_));
  AOI21_X1   g02173(.A1(new_n2365_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n2366_));
  AOI21_X1   g02174(.A1(new_n2366_), .A2(new_n2353_), .B(new_n2334_), .ZN(new_n2367_));
  OAI21_X1   g02175(.A1(new_n2367_), .A2(new_n2354_), .B(\asqrt[60] ), .ZN(new_n2368_));
  NAND2_X1   g02176(.A1(new_n2368_), .A2(new_n218_), .ZN(new_n2369_));
  OAI21_X1   g02177(.A1(new_n2369_), .A2(new_n2356_), .B(new_n2363_), .ZN(new_n2370_));
  AOI21_X1   g02178(.A1(new_n2370_), .A2(new_n2357_), .B(new_n207_), .ZN(new_n2371_));
  NOR3_X1    g02179(.A1(new_n2229_), .A2(new_n2121_), .A3(new_n2155_), .ZN(new_n2372_));
  INV_X1     g02180(.I(new_n2372_), .ZN(new_n2373_));
  NOR3_X1    g02181(.A1(new_n2121_), .A2(new_n2155_), .A3(new_n2183_), .ZN(new_n2374_));
  AOI22_X1   g02182(.A1(new_n2373_), .A2(new_n2183_), .B1(\asqrt[47] ), .B2(new_n2374_), .ZN(new_n2375_));
  NOR3_X1    g02183(.A1(new_n2367_), .A2(\asqrt[60] ), .A3(new_n2354_), .ZN(new_n2376_));
  OAI21_X1   g02184(.A1(new_n2350_), .A2(new_n2376_), .B(new_n2368_), .ZN(new_n2377_));
  AOI21_X1   g02185(.A1(new_n2377_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n2378_));
  AOI21_X1   g02186(.A1(new_n2378_), .A2(new_n2370_), .B(new_n2375_), .ZN(new_n2379_));
  INV_X1     g02187(.I(new_n2133_), .ZN(new_n2380_));
  NOR2_X1    g02188(.A1(new_n2144_), .A2(new_n2132_), .ZN(new_n2381_));
  NOR3_X1    g02189(.A1(new_n2380_), .A2(new_n2138_), .A3(new_n2381_), .ZN(new_n2382_));
  NAND2_X1   g02190(.A1(\asqrt[47] ), .A2(new_n2382_), .ZN(new_n2383_));
  INV_X1     g02191(.I(new_n2383_), .ZN(new_n2384_));
  NOR2_X1    g02192(.A1(new_n2380_), .A2(new_n2381_), .ZN(new_n2385_));
  AOI21_X1   g02193(.A1(\asqrt[47] ), .A2(new_n2385_), .B(new_n2137_), .ZN(new_n2386_));
  NOR2_X1    g02194(.A1(new_n2384_), .A2(new_n2386_), .ZN(new_n2387_));
  NOR3_X1    g02195(.A1(new_n2229_), .A2(new_n2189_), .A3(new_n2177_), .ZN(new_n2388_));
  NOR3_X1    g02196(.A1(new_n2387_), .A2(new_n2202_), .A3(new_n2388_), .ZN(new_n2389_));
  OAI21_X1   g02197(.A1(new_n2379_), .A2(new_n2371_), .B(new_n2389_), .ZN(new_n2390_));
  NAND2_X1   g02198(.A1(new_n2390_), .A2(new_n193_), .ZN(new_n2391_));
  INV_X1     g02199(.I(new_n2375_), .ZN(new_n2392_));
  NAND3_X1   g02200(.A1(new_n2370_), .A2(new_n207_), .A3(new_n2357_), .ZN(new_n2393_));
  NAND2_X1   g02201(.A1(new_n2393_), .A2(new_n2392_), .ZN(new_n2394_));
  INV_X1     g02202(.I(new_n2387_), .ZN(new_n2395_));
  NOR2_X1    g02203(.A1(new_n2371_), .A2(new_n2395_), .ZN(new_n2396_));
  AOI21_X1   g02204(.A1(\asqrt[47] ), .A2(new_n2150_), .B(new_n2173_), .ZN(new_n2397_));
  OAI21_X1   g02205(.A1(new_n2189_), .A2(new_n2177_), .B(\asqrt[63] ), .ZN(new_n2398_));
  NOR2_X1    g02206(.A1(new_n2397_), .A2(new_n2398_), .ZN(new_n2399_));
  AND3_X2    g02207(.A1(new_n2149_), .A2(new_n2147_), .A3(new_n2163_), .Z(new_n2400_));
  NAND4_X1   g02208(.A1(new_n2203_), .A2(new_n2190_), .A3(new_n2160_), .A4(new_n2400_), .ZN(new_n2401_));
  INV_X1     g02209(.I(new_n2401_), .ZN(new_n2402_));
  NOR2_X1    g02210(.A1(new_n2399_), .A2(new_n2402_), .ZN(new_n2403_));
  INV_X1     g02211(.I(new_n2403_), .ZN(new_n2404_));
  AOI21_X1   g02212(.A1(new_n2396_), .A2(new_n2394_), .B(new_n2404_), .ZN(new_n2405_));
  NAND2_X1   g02213(.A1(new_n2391_), .A2(new_n2405_), .ZN(\asqrt[46] ));
  NOR2_X1    g02214(.A1(\a[90] ), .A2(\a[91] ), .ZN(new_n2407_));
  INV_X1     g02215(.I(new_n2407_), .ZN(new_n2408_));
  NOR2_X1    g02216(.A1(new_n2408_), .A2(\a[92] ), .ZN(new_n2409_));
  INV_X1     g02217(.I(new_n2409_), .ZN(new_n2410_));
  INV_X1     g02218(.I(new_n2350_), .ZN(new_n2411_));
  NAND2_X1   g02219(.A1(new_n2330_), .A2(new_n306_), .ZN(new_n2412_));
  OAI21_X1   g02220(.A1(new_n2412_), .A2(new_n2367_), .B(new_n2411_), .ZN(new_n2413_));
  AOI21_X1   g02221(.A1(new_n2413_), .A2(new_n2368_), .B(new_n218_), .ZN(new_n2414_));
  NOR3_X1    g02222(.A1(new_n2329_), .A2(\asqrt[59] ), .A3(new_n2315_), .ZN(new_n2415_));
  OAI21_X1   g02223(.A1(new_n2334_), .A2(new_n2415_), .B(new_n2330_), .ZN(new_n2416_));
  AOI21_X1   g02224(.A1(new_n2416_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n2417_));
  AOI21_X1   g02225(.A1(new_n2417_), .A2(new_n2413_), .B(new_n2362_), .ZN(new_n2418_));
  OAI21_X1   g02226(.A1(new_n2418_), .A2(new_n2414_), .B(\asqrt[62] ), .ZN(new_n2419_));
  NOR3_X1    g02227(.A1(new_n2418_), .A2(\asqrt[62] ), .A3(new_n2414_), .ZN(new_n2420_));
  OAI21_X1   g02228(.A1(new_n2375_), .A2(new_n2420_), .B(new_n2419_), .ZN(new_n2421_));
  AOI21_X1   g02229(.A1(new_n2421_), .A2(new_n2389_), .B(\asqrt[63] ), .ZN(new_n2422_));
  NAND2_X1   g02230(.A1(new_n2419_), .A2(new_n2387_), .ZN(new_n2423_));
  OAI21_X1   g02231(.A1(new_n2423_), .A2(new_n2379_), .B(new_n2403_), .ZN(new_n2424_));
  OAI21_X1   g02232(.A1(new_n2422_), .A2(new_n2424_), .B(\a[92] ), .ZN(new_n2425_));
  AOI21_X1   g02233(.A1(new_n2425_), .A2(new_n2410_), .B(new_n2229_), .ZN(new_n2426_));
  INV_X1     g02234(.I(\a[92] ), .ZN(new_n2427_));
  AOI21_X1   g02235(.A1(new_n2391_), .A2(new_n2405_), .B(new_n2427_), .ZN(new_n2428_));
  NAND2_X1   g02236(.A1(new_n2163_), .A2(new_n2410_), .ZN(new_n2429_));
  NOR4_X1    g02237(.A1(new_n2175_), .A2(new_n2202_), .A3(new_n2161_), .A4(new_n2429_), .ZN(new_n2430_));
  INV_X1     g02238(.I(new_n2430_), .ZN(new_n2431_));
  NOR2_X1    g02239(.A1(new_n2428_), .A2(new_n2431_), .ZN(new_n2432_));
  AOI21_X1   g02240(.A1(new_n2391_), .A2(new_n2405_), .B(new_n2170_), .ZN(new_n2433_));
  INV_X1     g02241(.I(\a[93] ), .ZN(new_n2434_));
  AOI21_X1   g02242(.A1(\asqrt[46] ), .A2(new_n2427_), .B(new_n2434_), .ZN(new_n2435_));
  NOR3_X1    g02243(.A1(new_n2432_), .A2(new_n2435_), .A3(new_n2433_), .ZN(new_n2436_));
  OAI21_X1   g02244(.A1(new_n2436_), .A2(new_n2426_), .B(\asqrt[48] ), .ZN(new_n2437_));
  OAI21_X1   g02245(.A1(new_n2422_), .A2(new_n2424_), .B(new_n2169_), .ZN(new_n2438_));
  NAND2_X1   g02246(.A1(new_n2396_), .A2(new_n2394_), .ZN(new_n2439_));
  INV_X1     g02247(.I(new_n2399_), .ZN(new_n2440_));
  NOR2_X1    g02248(.A1(new_n2402_), .A2(new_n2229_), .ZN(new_n2441_));
  NAND4_X1   g02249(.A1(new_n2391_), .A2(new_n2439_), .A3(new_n2440_), .A4(new_n2441_), .ZN(new_n2442_));
  AOI21_X1   g02250(.A1(new_n2442_), .A2(new_n2438_), .B(new_n2182_), .ZN(new_n2443_));
  INV_X1     g02251(.I(new_n2439_), .ZN(new_n2444_));
  NAND2_X1   g02252(.A1(new_n2440_), .A2(new_n2441_), .ZN(new_n2445_));
  NOR3_X1    g02253(.A1(new_n2444_), .A2(new_n2422_), .A3(new_n2445_), .ZN(new_n2446_));
  NOR3_X1    g02254(.A1(new_n2446_), .A2(new_n2433_), .A3(\a[94] ), .ZN(new_n2447_));
  OAI21_X1   g02255(.A1(new_n2428_), .A2(new_n2409_), .B(\asqrt[47] ), .ZN(new_n2448_));
  NAND2_X1   g02256(.A1(new_n2448_), .A2(new_n1956_), .ZN(new_n2449_));
  OAI22_X1   g02257(.A1(new_n2436_), .A2(new_n2449_), .B1(new_n2443_), .B2(new_n2447_), .ZN(new_n2450_));
  AOI21_X1   g02258(.A1(new_n2450_), .A2(new_n2437_), .B(new_n1806_), .ZN(new_n2451_));
  NOR3_X1    g02259(.A1(new_n2301_), .A2(new_n2181_), .A3(new_n2195_), .ZN(new_n2452_));
  NAND3_X1   g02260(.A1(\asqrt[46] ), .A2(new_n2217_), .A3(new_n2286_), .ZN(new_n2453_));
  AOI22_X1   g02261(.A1(new_n2453_), .A2(new_n2301_), .B1(\asqrt[46] ), .B2(new_n2452_), .ZN(new_n2454_));
  AOI21_X1   g02262(.A1(new_n2391_), .A2(new_n2405_), .B(\a[92] ), .ZN(new_n2455_));
  OAI21_X1   g02263(.A1(new_n2434_), .A2(new_n2455_), .B(new_n2438_), .ZN(new_n2456_));
  OAI21_X1   g02264(.A1(new_n2456_), .A2(new_n2432_), .B(new_n2448_), .ZN(new_n2457_));
  AOI21_X1   g02265(.A1(new_n2457_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n2458_));
  AOI21_X1   g02266(.A1(new_n2458_), .A2(new_n2450_), .B(new_n2454_), .ZN(new_n2459_));
  OAI21_X1   g02267(.A1(new_n2459_), .A2(new_n2451_), .B(\asqrt[50] ), .ZN(new_n2460_));
  NOR2_X1    g02268(.A1(new_n2206_), .A2(new_n2209_), .ZN(new_n2461_));
  NOR2_X1    g02269(.A1(new_n2199_), .A2(new_n2211_), .ZN(new_n2462_));
  INV_X1     g02270(.I(new_n2462_), .ZN(new_n2463_));
  NAND4_X1   g02271(.A1(\asqrt[46] ), .A2(new_n2200_), .A3(new_n2461_), .A4(new_n2463_), .ZN(new_n2464_));
  INV_X1     g02272(.I(\asqrt[46] ), .ZN(new_n2465_));
  NOR3_X1    g02273(.A1(new_n2465_), .A2(new_n2290_), .A3(new_n2462_), .ZN(new_n2466_));
  OAI21_X1   g02274(.A1(new_n2466_), .A2(new_n2461_), .B(new_n2464_), .ZN(new_n2467_));
  NAND2_X1   g02275(.A1(new_n2425_), .A2(new_n2430_), .ZN(new_n2468_));
  OAI21_X1   g02276(.A1(new_n2422_), .A2(new_n2424_), .B(new_n2427_), .ZN(new_n2469_));
  NAND2_X1   g02277(.A1(new_n2469_), .A2(\a[93] ), .ZN(new_n2470_));
  NAND3_X1   g02278(.A1(new_n2468_), .A2(new_n2470_), .A3(new_n2438_), .ZN(new_n2471_));
  AOI21_X1   g02279(.A1(new_n2471_), .A2(new_n2448_), .B(new_n1956_), .ZN(new_n2472_));
  OAI21_X1   g02280(.A1(new_n2446_), .A2(new_n2433_), .B(\a[94] ), .ZN(new_n2473_));
  NAND3_X1   g02281(.A1(new_n2442_), .A2(new_n2438_), .A3(new_n2182_), .ZN(new_n2474_));
  NAND2_X1   g02282(.A1(new_n2425_), .A2(new_n2410_), .ZN(new_n2475_));
  AOI21_X1   g02283(.A1(new_n2475_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n2476_));
  AOI22_X1   g02284(.A1(new_n2471_), .A2(new_n2476_), .B1(new_n2473_), .B2(new_n2474_), .ZN(new_n2477_));
  OAI21_X1   g02285(.A1(new_n2477_), .A2(new_n2472_), .B(\asqrt[49] ), .ZN(new_n2478_));
  NAND2_X1   g02286(.A1(new_n2478_), .A2(new_n1612_), .ZN(new_n2479_));
  OAI21_X1   g02287(.A1(new_n2479_), .A2(new_n2459_), .B(new_n2467_), .ZN(new_n2480_));
  AOI21_X1   g02288(.A1(new_n2480_), .A2(new_n2460_), .B(new_n1376_), .ZN(new_n2481_));
  NOR2_X1    g02289(.A1(new_n2303_), .A2(new_n2295_), .ZN(new_n2482_));
  NOR3_X1    g02290(.A1(new_n2465_), .A2(new_n2213_), .A3(new_n2482_), .ZN(new_n2483_));
  INV_X1     g02291(.I(new_n2483_), .ZN(new_n2484_));
  NOR3_X1    g02292(.A1(new_n2482_), .A2(new_n2213_), .A3(new_n2300_), .ZN(new_n2485_));
  AOI22_X1   g02293(.A1(new_n2484_), .A2(new_n2300_), .B1(\asqrt[46] ), .B2(new_n2485_), .ZN(new_n2486_));
  INV_X1     g02294(.I(new_n2454_), .ZN(new_n2487_));
  AOI21_X1   g02295(.A1(\a[93] ), .A2(new_n2469_), .B(new_n2433_), .ZN(new_n2488_));
  AOI21_X1   g02296(.A1(new_n2488_), .A2(new_n2468_), .B(new_n2426_), .ZN(new_n2489_));
  OAI21_X1   g02297(.A1(new_n2489_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n2490_));
  OAI21_X1   g02298(.A1(new_n2490_), .A2(new_n2477_), .B(new_n2487_), .ZN(new_n2491_));
  NAND2_X1   g02299(.A1(new_n2491_), .A2(new_n2478_), .ZN(new_n2492_));
  AOI21_X1   g02300(.A1(new_n2492_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n2493_));
  AOI21_X1   g02301(.A1(new_n2493_), .A2(new_n2480_), .B(new_n2486_), .ZN(new_n2494_));
  OAI21_X1   g02302(.A1(new_n2494_), .A2(new_n2481_), .B(\asqrt[52] ), .ZN(new_n2495_));
  NOR3_X1    g02303(.A1(new_n2224_), .A2(new_n2233_), .A3(new_n2231_), .ZN(new_n2496_));
  NOR3_X1    g02304(.A1(new_n2465_), .A2(new_n2224_), .A3(new_n2233_), .ZN(new_n2497_));
  INV_X1     g02305(.I(new_n2497_), .ZN(new_n2498_));
  AOI22_X1   g02306(.A1(new_n2498_), .A2(new_n2231_), .B1(\asqrt[46] ), .B2(new_n2496_), .ZN(new_n2499_));
  INV_X1     g02307(.I(new_n2499_), .ZN(new_n2500_));
  INV_X1     g02308(.I(new_n2460_), .ZN(new_n2501_));
  INV_X1     g02309(.I(new_n2467_), .ZN(new_n2502_));
  NOR3_X1    g02310(.A1(new_n2459_), .A2(new_n2451_), .A3(\asqrt[50] ), .ZN(new_n2503_));
  NOR2_X1    g02311(.A1(new_n2503_), .A2(new_n2502_), .ZN(new_n2504_));
  OAI21_X1   g02312(.A1(new_n2504_), .A2(new_n2501_), .B(\asqrt[51] ), .ZN(new_n2505_));
  NAND2_X1   g02313(.A1(new_n2505_), .A2(new_n1256_), .ZN(new_n2506_));
  OAI21_X1   g02314(.A1(new_n2506_), .A2(new_n2494_), .B(new_n2500_), .ZN(new_n2507_));
  AOI21_X1   g02315(.A1(new_n2507_), .A2(new_n2495_), .B(new_n1103_), .ZN(new_n2508_));
  NAND2_X1   g02316(.A1(new_n2306_), .A2(new_n2298_), .ZN(new_n2509_));
  NAND3_X1   g02317(.A1(\asqrt[46] ), .A2(new_n2235_), .A3(new_n2509_), .ZN(new_n2510_));
  AND3_X2    g02318(.A1(new_n2235_), .A2(new_n2240_), .A3(new_n2509_), .Z(new_n2511_));
  AOI22_X1   g02319(.A1(new_n2510_), .A2(new_n2241_), .B1(\asqrt[46] ), .B2(new_n2511_), .ZN(new_n2512_));
  INV_X1     g02320(.I(new_n2486_), .ZN(new_n2513_));
  NAND2_X1   g02321(.A1(new_n2460_), .A2(new_n1376_), .ZN(new_n2514_));
  OAI21_X1   g02322(.A1(new_n2504_), .A2(new_n2514_), .B(new_n2513_), .ZN(new_n2515_));
  AOI21_X1   g02323(.A1(new_n2515_), .A2(new_n2505_), .B(new_n1256_), .ZN(new_n2516_));
  NOR2_X1    g02324(.A1(new_n2516_), .A2(\asqrt[53] ), .ZN(new_n2517_));
  AOI21_X1   g02325(.A1(new_n2517_), .A2(new_n2507_), .B(new_n2512_), .ZN(new_n2518_));
  OAI21_X1   g02326(.A1(new_n2518_), .A2(new_n2508_), .B(\asqrt[54] ), .ZN(new_n2519_));
  INV_X1     g02327(.I(new_n2248_), .ZN(new_n2520_));
  NOR3_X1    g02328(.A1(new_n2244_), .A2(new_n2322_), .A3(new_n2520_), .ZN(new_n2521_));
  NOR3_X1    g02329(.A1(new_n2465_), .A2(new_n2244_), .A3(new_n2322_), .ZN(new_n2522_));
  INV_X1     g02330(.I(new_n2522_), .ZN(new_n2523_));
  AOI22_X1   g02331(.A1(new_n2523_), .A2(new_n2520_), .B1(\asqrt[46] ), .B2(new_n2521_), .ZN(new_n2524_));
  INV_X1     g02332(.I(new_n2524_), .ZN(new_n2525_));
  OAI21_X1   g02333(.A1(new_n2502_), .A2(new_n2503_), .B(new_n2460_), .ZN(new_n2526_));
  AOI21_X1   g02334(.A1(new_n2526_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n2527_));
  AOI21_X1   g02335(.A1(new_n2527_), .A2(new_n2515_), .B(new_n2499_), .ZN(new_n2528_));
  OAI21_X1   g02336(.A1(new_n2528_), .A2(new_n2516_), .B(\asqrt[53] ), .ZN(new_n2529_));
  INV_X1     g02337(.I(new_n2512_), .ZN(new_n2530_));
  NAND2_X1   g02338(.A1(new_n2495_), .A2(new_n1103_), .ZN(new_n2531_));
  OAI21_X1   g02339(.A1(new_n2531_), .A2(new_n2528_), .B(new_n2530_), .ZN(new_n2532_));
  NAND3_X1   g02340(.A1(new_n2532_), .A2(new_n904_), .A3(new_n2529_), .ZN(new_n2533_));
  NAND2_X1   g02341(.A1(new_n2533_), .A2(new_n2525_), .ZN(new_n2534_));
  AOI21_X1   g02342(.A1(new_n2534_), .A2(new_n2519_), .B(new_n823_), .ZN(new_n2535_));
  NOR3_X1    g02343(.A1(new_n2465_), .A2(new_n2253_), .A3(new_n2259_), .ZN(new_n2536_));
  INV_X1     g02344(.I(new_n2536_), .ZN(new_n2537_));
  NOR3_X1    g02345(.A1(new_n2253_), .A2(new_n2285_), .A3(new_n2259_), .ZN(new_n2538_));
  AOI22_X1   g02346(.A1(new_n2537_), .A2(new_n2285_), .B1(\asqrt[46] ), .B2(new_n2538_), .ZN(new_n2539_));
  AOI21_X1   g02347(.A1(new_n2532_), .A2(new_n2529_), .B(new_n904_), .ZN(new_n2540_));
  NOR2_X1    g02348(.A1(new_n2540_), .A2(\asqrt[55] ), .ZN(new_n2541_));
  AOI21_X1   g02349(.A1(new_n2541_), .A2(new_n2534_), .B(new_n2539_), .ZN(new_n2542_));
  OAI21_X1   g02350(.A1(new_n2542_), .A2(new_n2535_), .B(\asqrt[56] ), .ZN(new_n2543_));
  INV_X1     g02351(.I(new_n2311_), .ZN(new_n2544_));
  NOR3_X1    g02352(.A1(new_n2544_), .A2(new_n2321_), .A3(new_n2269_), .ZN(new_n2545_));
  NOR3_X1    g02353(.A1(new_n2465_), .A2(new_n2321_), .A3(new_n2544_), .ZN(new_n2546_));
  INV_X1     g02354(.I(new_n2546_), .ZN(new_n2547_));
  AOI22_X1   g02355(.A1(new_n2547_), .A2(new_n2269_), .B1(\asqrt[46] ), .B2(new_n2545_), .ZN(new_n2548_));
  INV_X1     g02356(.I(new_n2548_), .ZN(new_n2549_));
  NOR3_X1    g02357(.A1(new_n2494_), .A2(new_n2481_), .A3(\asqrt[52] ), .ZN(new_n2550_));
  OAI21_X1   g02358(.A1(new_n2499_), .A2(new_n2550_), .B(new_n2495_), .ZN(new_n2551_));
  AOI21_X1   g02359(.A1(new_n2551_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n2552_));
  AOI21_X1   g02360(.A1(new_n2552_), .A2(new_n2532_), .B(new_n2524_), .ZN(new_n2553_));
  OAI21_X1   g02361(.A1(new_n2553_), .A2(new_n2540_), .B(\asqrt[55] ), .ZN(new_n2554_));
  NAND2_X1   g02362(.A1(new_n2554_), .A2(new_n703_), .ZN(new_n2555_));
  OAI21_X1   g02363(.A1(new_n2555_), .A2(new_n2542_), .B(new_n2549_), .ZN(new_n2556_));
  AOI21_X1   g02364(.A1(new_n2556_), .A2(new_n2543_), .B(new_n531_), .ZN(new_n2557_));
  INV_X1     g02365(.I(new_n2557_), .ZN(new_n2558_));
  INV_X1     g02366(.I(new_n2556_), .ZN(new_n2559_));
  NOR3_X1    g02367(.A1(new_n2465_), .A2(new_n2272_), .A3(new_n2326_), .ZN(new_n2560_));
  INV_X1     g02368(.I(new_n2560_), .ZN(new_n2561_));
  NOR3_X1    g02369(.A1(new_n2272_), .A2(new_n2326_), .A3(new_n2337_), .ZN(new_n2562_));
  AOI22_X1   g02370(.A1(new_n2561_), .A2(new_n2337_), .B1(\asqrt[46] ), .B2(new_n2562_), .ZN(new_n2563_));
  INV_X1     g02371(.I(new_n2563_), .ZN(new_n2564_));
  NAND2_X1   g02372(.A1(new_n2543_), .A2(new_n531_), .ZN(new_n2565_));
  OAI21_X1   g02373(.A1(new_n2559_), .A2(new_n2565_), .B(new_n2564_), .ZN(new_n2566_));
  AOI21_X1   g02374(.A1(new_n2566_), .A2(new_n2558_), .B(new_n436_), .ZN(new_n2567_));
  NOR3_X1    g02375(.A1(new_n2336_), .A2(new_n2284_), .A3(new_n2364_), .ZN(new_n2568_));
  NOR3_X1    g02376(.A1(new_n2465_), .A2(new_n2336_), .A3(new_n2364_), .ZN(new_n2569_));
  INV_X1     g02377(.I(new_n2569_), .ZN(new_n2570_));
  AOI22_X1   g02378(.A1(new_n2570_), .A2(new_n2284_), .B1(\asqrt[46] ), .B2(new_n2568_), .ZN(new_n2571_));
  NOR2_X1    g02379(.A1(new_n2557_), .A2(\asqrt[58] ), .ZN(new_n2572_));
  AOI21_X1   g02380(.A1(new_n2572_), .A2(new_n2566_), .B(new_n2571_), .ZN(new_n2573_));
  OAI21_X1   g02381(.A1(new_n2573_), .A2(new_n2567_), .B(\asqrt[59] ), .ZN(new_n2574_));
  NOR2_X1    g02382(.A1(new_n2352_), .A2(new_n2341_), .ZN(new_n2575_));
  NOR3_X1    g02383(.A1(new_n2465_), .A2(new_n2315_), .A3(new_n2575_), .ZN(new_n2576_));
  INV_X1     g02384(.I(new_n2576_), .ZN(new_n2577_));
  NOR3_X1    g02385(.A1(new_n2575_), .A2(new_n2315_), .A3(new_n2351_), .ZN(new_n2578_));
  AOI22_X1   g02386(.A1(new_n2577_), .A2(new_n2351_), .B1(\asqrt[46] ), .B2(new_n2578_), .ZN(new_n2579_));
  INV_X1     g02387(.I(new_n2579_), .ZN(new_n2580_));
  NOR3_X1    g02388(.A1(new_n2528_), .A2(new_n2516_), .A3(\asqrt[53] ), .ZN(new_n2581_));
  OAI21_X1   g02389(.A1(new_n2512_), .A2(new_n2581_), .B(new_n2529_), .ZN(new_n2582_));
  AOI22_X1   g02390(.A1(new_n2533_), .A2(new_n2525_), .B1(new_n2582_), .B2(\asqrt[54] ), .ZN(new_n2583_));
  NOR3_X1    g02391(.A1(new_n2553_), .A2(\asqrt[55] ), .A3(new_n2540_), .ZN(new_n2584_));
  OAI22_X1   g02392(.A1(new_n2584_), .A2(new_n2539_), .B1(new_n2583_), .B2(new_n823_), .ZN(new_n2585_));
  AOI21_X1   g02393(.A1(new_n2585_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n2586_));
  AOI21_X1   g02394(.A1(new_n2586_), .A2(new_n2556_), .B(new_n2563_), .ZN(new_n2587_));
  OAI21_X1   g02395(.A1(new_n2587_), .A2(new_n2557_), .B(\asqrt[58] ), .ZN(new_n2588_));
  NAND2_X1   g02396(.A1(new_n2588_), .A2(new_n327_), .ZN(new_n2589_));
  OAI21_X1   g02397(.A1(new_n2589_), .A2(new_n2573_), .B(new_n2580_), .ZN(new_n2590_));
  AOI21_X1   g02398(.A1(new_n2590_), .A2(new_n2574_), .B(new_n306_), .ZN(new_n2591_));
  INV_X1     g02399(.I(new_n2591_), .ZN(new_n2592_));
  INV_X1     g02400(.I(new_n2590_), .ZN(new_n2593_));
  NOR3_X1    g02401(.A1(new_n2354_), .A2(new_n2415_), .A3(new_n2335_), .ZN(new_n2594_));
  NOR3_X1    g02402(.A1(new_n2465_), .A2(new_n2354_), .A3(new_n2415_), .ZN(new_n2595_));
  INV_X1     g02403(.I(new_n2595_), .ZN(new_n2596_));
  AOI22_X1   g02404(.A1(new_n2596_), .A2(new_n2335_), .B1(\asqrt[46] ), .B2(new_n2594_), .ZN(new_n2597_));
  INV_X1     g02405(.I(new_n2597_), .ZN(new_n2598_));
  NAND2_X1   g02406(.A1(new_n2574_), .A2(new_n306_), .ZN(new_n2599_));
  OAI21_X1   g02407(.A1(new_n2593_), .A2(new_n2599_), .B(new_n2598_), .ZN(new_n2600_));
  AOI21_X1   g02408(.A1(new_n2600_), .A2(new_n2592_), .B(new_n218_), .ZN(new_n2601_));
  NOR3_X1    g02409(.A1(new_n2465_), .A2(new_n2345_), .A3(new_n2376_), .ZN(new_n2602_));
  INV_X1     g02410(.I(new_n2602_), .ZN(new_n2603_));
  NOR3_X1    g02411(.A1(new_n2345_), .A2(new_n2411_), .A3(new_n2376_), .ZN(new_n2604_));
  AOI22_X1   g02412(.A1(new_n2603_), .A2(new_n2411_), .B1(\asqrt[46] ), .B2(new_n2604_), .ZN(new_n2605_));
  NOR2_X1    g02413(.A1(new_n2591_), .A2(\asqrt[61] ), .ZN(new_n2606_));
  AOI21_X1   g02414(.A1(new_n2606_), .A2(new_n2600_), .B(new_n2605_), .ZN(new_n2607_));
  OAI21_X1   g02415(.A1(new_n2607_), .A2(new_n2601_), .B(\asqrt[62] ), .ZN(new_n2608_));
  NOR2_X1    g02416(.A1(new_n2369_), .A2(new_n2356_), .ZN(new_n2609_));
  NOR3_X1    g02417(.A1(new_n2609_), .A2(new_n2414_), .A3(new_n2363_), .ZN(new_n2610_));
  NOR3_X1    g02418(.A1(new_n2465_), .A2(new_n2414_), .A3(new_n2609_), .ZN(new_n2611_));
  INV_X1     g02419(.I(new_n2611_), .ZN(new_n2612_));
  AOI22_X1   g02420(.A1(new_n2612_), .A2(new_n2363_), .B1(\asqrt[46] ), .B2(new_n2610_), .ZN(new_n2613_));
  INV_X1     g02421(.I(new_n2613_), .ZN(new_n2614_));
  NOR3_X1    g02422(.A1(new_n2587_), .A2(\asqrt[58] ), .A3(new_n2557_), .ZN(new_n2615_));
  OAI21_X1   g02423(.A1(new_n2571_), .A2(new_n2615_), .B(new_n2588_), .ZN(new_n2616_));
  AOI21_X1   g02424(.A1(new_n2616_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n2617_));
  AOI21_X1   g02425(.A1(new_n2617_), .A2(new_n2590_), .B(new_n2597_), .ZN(new_n2618_));
  OAI21_X1   g02426(.A1(new_n2618_), .A2(new_n2591_), .B(\asqrt[61] ), .ZN(new_n2619_));
  NAND2_X1   g02427(.A1(new_n2619_), .A2(new_n207_), .ZN(new_n2620_));
  OAI21_X1   g02428(.A1(new_n2620_), .A2(new_n2607_), .B(new_n2614_), .ZN(new_n2621_));
  NAND4_X1   g02429(.A1(\asqrt[46] ), .A2(new_n2419_), .A3(new_n2375_), .A4(new_n2393_), .ZN(new_n2622_));
  NAND2_X1   g02430(.A1(new_n2419_), .A2(new_n2393_), .ZN(new_n2623_));
  OAI21_X1   g02431(.A1(new_n2465_), .A2(new_n2623_), .B(new_n2392_), .ZN(new_n2624_));
  NAND2_X1   g02432(.A1(new_n2624_), .A2(new_n2622_), .ZN(new_n2625_));
  AOI21_X1   g02433(.A1(new_n2394_), .A2(new_n2419_), .B(new_n2387_), .ZN(new_n2626_));
  AOI21_X1   g02434(.A1(\asqrt[46] ), .A2(new_n2626_), .B(new_n2444_), .ZN(new_n2627_));
  NAND2_X1   g02435(.A1(new_n2625_), .A2(new_n2627_), .ZN(new_n2628_));
  AOI21_X1   g02436(.A1(new_n2621_), .A2(new_n2608_), .B(new_n2628_), .ZN(new_n2629_));
  NOR3_X1    g02437(.A1(new_n2618_), .A2(\asqrt[61] ), .A3(new_n2591_), .ZN(new_n2630_));
  OAI21_X1   g02438(.A1(new_n2605_), .A2(new_n2630_), .B(new_n2619_), .ZN(new_n2631_));
  AOI21_X1   g02439(.A1(new_n2631_), .A2(\asqrt[62] ), .B(new_n2625_), .ZN(new_n2632_));
  AOI21_X1   g02440(.A1(\asqrt[46] ), .A2(new_n2395_), .B(new_n2421_), .ZN(new_n2633_));
  OR3_X2     g02441(.A1(new_n2633_), .A2(new_n193_), .A3(new_n2626_), .Z(new_n2634_));
  NAND2_X1   g02442(.A1(new_n2383_), .A2(new_n2401_), .ZN(new_n2635_));
  NOR4_X1    g02443(.A1(new_n2444_), .A2(new_n2386_), .A3(new_n2399_), .A4(new_n2635_), .ZN(new_n2636_));
  NAND2_X1   g02444(.A1(new_n2636_), .A2(new_n2391_), .ZN(new_n2637_));
  NAND2_X1   g02445(.A1(new_n2634_), .A2(new_n2637_), .ZN(new_n2638_));
  AOI21_X1   g02446(.A1(new_n2632_), .A2(new_n2621_), .B(new_n2638_), .ZN(new_n2639_));
  OAI21_X1   g02447(.A1(\asqrt[63] ), .A2(new_n2629_), .B(new_n2639_), .ZN(\asqrt[45] ));
  INV_X1     g02448(.I(\asqrt[45] ), .ZN(new_n2641_));
  NOR2_X1    g02449(.A1(\a[88] ), .A2(\a[89] ), .ZN(new_n2642_));
  INV_X1     g02450(.I(new_n2642_), .ZN(new_n2643_));
  NOR2_X1    g02451(.A1(new_n2643_), .A2(\a[90] ), .ZN(new_n2644_));
  INV_X1     g02452(.I(new_n2644_), .ZN(new_n2645_));
  NOR2_X1    g02453(.A1(new_n2629_), .A2(\asqrt[63] ), .ZN(new_n2646_));
  INV_X1     g02454(.I(new_n2621_), .ZN(new_n2647_));
  INV_X1     g02455(.I(new_n2625_), .ZN(new_n2648_));
  NAND2_X1   g02456(.A1(new_n2608_), .A2(new_n2648_), .ZN(new_n2649_));
  INV_X1     g02457(.I(new_n2638_), .ZN(new_n2650_));
  OAI21_X1   g02458(.A1(new_n2647_), .A2(new_n2649_), .B(new_n2650_), .ZN(new_n2651_));
  OAI21_X1   g02459(.A1(new_n2646_), .A2(new_n2651_), .B(\a[90] ), .ZN(new_n2652_));
  AOI21_X1   g02460(.A1(new_n2652_), .A2(new_n2645_), .B(new_n2465_), .ZN(new_n2653_));
  INV_X1     g02461(.I(\a[90] ), .ZN(new_n2654_));
  INV_X1     g02462(.I(new_n2605_), .ZN(new_n2655_));
  INV_X1     g02463(.I(new_n2571_), .ZN(new_n2656_));
  INV_X1     g02464(.I(new_n2539_), .ZN(new_n2657_));
  NAND2_X1   g02465(.A1(new_n2519_), .A2(new_n823_), .ZN(new_n2658_));
  OAI21_X1   g02466(.A1(new_n2658_), .A2(new_n2553_), .B(new_n2657_), .ZN(new_n2659_));
  NAND3_X1   g02467(.A1(new_n2659_), .A2(new_n703_), .A3(new_n2554_), .ZN(new_n2660_));
  AOI22_X1   g02468(.A1(new_n2660_), .A2(new_n2549_), .B1(\asqrt[56] ), .B2(new_n2585_), .ZN(new_n2661_));
  OAI21_X1   g02469(.A1(new_n2661_), .A2(new_n531_), .B(new_n436_), .ZN(new_n2662_));
  OAI21_X1   g02470(.A1(new_n2662_), .A2(new_n2587_), .B(new_n2656_), .ZN(new_n2663_));
  NAND3_X1   g02471(.A1(new_n2663_), .A2(new_n327_), .A3(new_n2588_), .ZN(new_n2664_));
  AOI22_X1   g02472(.A1(new_n2664_), .A2(new_n2580_), .B1(new_n2616_), .B2(\asqrt[59] ), .ZN(new_n2665_));
  OAI21_X1   g02473(.A1(new_n2665_), .A2(new_n306_), .B(new_n218_), .ZN(new_n2666_));
  OAI21_X1   g02474(.A1(new_n2666_), .A2(new_n2618_), .B(new_n2655_), .ZN(new_n2667_));
  NAND3_X1   g02475(.A1(new_n2667_), .A2(new_n207_), .A3(new_n2619_), .ZN(new_n2668_));
  AOI22_X1   g02476(.A1(new_n2668_), .A2(new_n2614_), .B1(new_n2631_), .B2(\asqrt[62] ), .ZN(new_n2669_));
  OAI21_X1   g02477(.A1(new_n2669_), .A2(new_n2628_), .B(new_n193_), .ZN(new_n2670_));
  AOI21_X1   g02478(.A1(new_n2670_), .A2(new_n2639_), .B(new_n2654_), .ZN(new_n2671_));
  NOR3_X1    g02479(.A1(new_n2399_), .A2(new_n2402_), .A3(new_n2644_), .ZN(new_n2672_));
  NAND3_X1   g02480(.A1(new_n2391_), .A2(new_n2439_), .A3(new_n2672_), .ZN(new_n2673_));
  NOR2_X1    g02481(.A1(new_n2671_), .A2(new_n2673_), .ZN(new_n2674_));
  INV_X1     g02482(.I(new_n2674_), .ZN(new_n2675_));
  AOI21_X1   g02483(.A1(new_n2670_), .A2(new_n2639_), .B(new_n2408_), .ZN(new_n2676_));
  INV_X1     g02484(.I(\a[91] ), .ZN(new_n2677_));
  AOI21_X1   g02485(.A1(\asqrt[45] ), .A2(new_n2654_), .B(new_n2677_), .ZN(new_n2678_));
  NOR2_X1    g02486(.A1(new_n2678_), .A2(new_n2676_), .ZN(new_n2679_));
  AOI21_X1   g02487(.A1(new_n2679_), .A2(new_n2675_), .B(new_n2653_), .ZN(new_n2680_));
  NOR2_X1    g02488(.A1(new_n2680_), .A2(new_n2229_), .ZN(new_n2681_));
  OAI21_X1   g02489(.A1(new_n2646_), .A2(new_n2651_), .B(new_n2407_), .ZN(new_n2682_));
  NAND2_X1   g02490(.A1(new_n2632_), .A2(new_n2621_), .ZN(new_n2683_));
  OAI21_X1   g02491(.A1(new_n2636_), .A2(new_n2405_), .B(new_n2391_), .ZN(new_n2684_));
  NAND4_X1   g02492(.A1(new_n2670_), .A2(new_n2683_), .A3(new_n2634_), .A4(new_n2684_), .ZN(new_n2685_));
  AOI21_X1   g02493(.A1(new_n2685_), .A2(new_n2682_), .B(new_n2427_), .ZN(new_n2686_));
  NAND3_X1   g02494(.A1(new_n2683_), .A2(new_n2634_), .A3(new_n2684_), .ZN(new_n2687_));
  NOR2_X1    g02495(.A1(new_n2687_), .A2(new_n2646_), .ZN(new_n2688_));
  NOR3_X1    g02496(.A1(new_n2688_), .A2(new_n2676_), .A3(\a[92] ), .ZN(new_n2689_));
  NOR2_X1    g02497(.A1(new_n2689_), .A2(new_n2686_), .ZN(new_n2690_));
  NOR3_X1    g02498(.A1(new_n2674_), .A2(new_n2678_), .A3(new_n2676_), .ZN(new_n2691_));
  AOI21_X1   g02499(.A1(\asqrt[45] ), .A2(\a[90] ), .B(new_n2644_), .ZN(new_n2692_));
  OAI21_X1   g02500(.A1(new_n2692_), .A2(new_n2465_), .B(new_n2229_), .ZN(new_n2693_));
  NOR2_X1    g02501(.A1(new_n2691_), .A2(new_n2693_), .ZN(new_n2694_));
  NOR2_X1    g02502(.A1(new_n2694_), .A2(new_n2690_), .ZN(new_n2695_));
  OAI21_X1   g02503(.A1(new_n2695_), .A2(new_n2681_), .B(\asqrt[48] ), .ZN(new_n2696_));
  NOR3_X1    g02504(.A1(new_n2488_), .A2(new_n2426_), .A3(new_n2432_), .ZN(new_n2697_));
  NAND3_X1   g02505(.A1(\asqrt[45] ), .A2(new_n2448_), .A3(new_n2468_), .ZN(new_n2698_));
  AOI22_X1   g02506(.A1(new_n2698_), .A2(new_n2488_), .B1(\asqrt[45] ), .B2(new_n2697_), .ZN(new_n2699_));
  INV_X1     g02507(.I(new_n2699_), .ZN(new_n2700_));
  OAI21_X1   g02508(.A1(new_n2680_), .A2(new_n2229_), .B(new_n1956_), .ZN(new_n2701_));
  OAI21_X1   g02509(.A1(new_n2701_), .A2(new_n2695_), .B(new_n2700_), .ZN(new_n2702_));
  AOI21_X1   g02510(.A1(new_n2702_), .A2(new_n2696_), .B(new_n1806_), .ZN(new_n2703_));
  NOR2_X1    g02511(.A1(new_n2447_), .A2(new_n2443_), .ZN(new_n2704_));
  NOR2_X1    g02512(.A1(new_n2436_), .A2(new_n2449_), .ZN(new_n2705_));
  INV_X1     g02513(.I(new_n2705_), .ZN(new_n2706_));
  NAND4_X1   g02514(.A1(\asqrt[45] ), .A2(new_n2437_), .A3(new_n2704_), .A4(new_n2706_), .ZN(new_n2707_));
  NOR3_X1    g02515(.A1(new_n2641_), .A2(new_n2472_), .A3(new_n2705_), .ZN(new_n2708_));
  OAI21_X1   g02516(.A1(new_n2708_), .A2(new_n2704_), .B(new_n2707_), .ZN(new_n2709_));
  INV_X1     g02517(.I(new_n2709_), .ZN(new_n2710_));
  OAI21_X1   g02518(.A1(new_n2691_), .A2(new_n2653_), .B(\asqrt[47] ), .ZN(new_n2711_));
  OAI22_X1   g02519(.A1(new_n2691_), .A2(new_n2693_), .B1(new_n2686_), .B2(new_n2689_), .ZN(new_n2712_));
  AOI21_X1   g02520(.A1(new_n2712_), .A2(new_n2711_), .B(new_n1956_), .ZN(new_n2713_));
  OAI21_X1   g02521(.A1(new_n2671_), .A2(new_n2644_), .B(\asqrt[46] ), .ZN(new_n2714_));
  AOI21_X1   g02522(.A1(new_n2670_), .A2(new_n2639_), .B(\a[90] ), .ZN(new_n2715_));
  OAI21_X1   g02523(.A1(new_n2677_), .A2(new_n2715_), .B(new_n2682_), .ZN(new_n2716_));
  OAI21_X1   g02524(.A1(new_n2716_), .A2(new_n2674_), .B(new_n2714_), .ZN(new_n2717_));
  AOI21_X1   g02525(.A1(new_n2717_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n2718_));
  AOI21_X1   g02526(.A1(new_n2718_), .A2(new_n2712_), .B(new_n2699_), .ZN(new_n2719_));
  NOR3_X1    g02527(.A1(new_n2719_), .A2(new_n2713_), .A3(\asqrt[49] ), .ZN(new_n2720_));
  NOR2_X1    g02528(.A1(new_n2720_), .A2(new_n2710_), .ZN(new_n2721_));
  OAI21_X1   g02529(.A1(new_n2721_), .A2(new_n2703_), .B(\asqrt[50] ), .ZN(new_n2722_));
  NOR2_X1    g02530(.A1(new_n2490_), .A2(new_n2477_), .ZN(new_n2723_));
  NOR3_X1    g02531(.A1(new_n2641_), .A2(new_n2451_), .A3(new_n2723_), .ZN(new_n2724_));
  INV_X1     g02532(.I(new_n2724_), .ZN(new_n2725_));
  NOR3_X1    g02533(.A1(new_n2723_), .A2(new_n2451_), .A3(new_n2487_), .ZN(new_n2726_));
  AOI22_X1   g02534(.A1(new_n2725_), .A2(new_n2487_), .B1(\asqrt[45] ), .B2(new_n2726_), .ZN(new_n2727_));
  INV_X1     g02535(.I(new_n2727_), .ZN(new_n2728_));
  OAI21_X1   g02536(.A1(new_n2719_), .A2(new_n2713_), .B(\asqrt[49] ), .ZN(new_n2729_));
  NAND2_X1   g02537(.A1(new_n2729_), .A2(new_n1612_), .ZN(new_n2730_));
  OAI21_X1   g02538(.A1(new_n2721_), .A2(new_n2730_), .B(new_n2728_), .ZN(new_n2731_));
  AOI21_X1   g02539(.A1(new_n2731_), .A2(new_n2722_), .B(new_n1376_), .ZN(new_n2732_));
  NOR3_X1    g02540(.A1(new_n2501_), .A2(new_n2503_), .A3(new_n2467_), .ZN(new_n2733_));
  NOR3_X1    g02541(.A1(new_n2641_), .A2(new_n2501_), .A3(new_n2503_), .ZN(new_n2734_));
  INV_X1     g02542(.I(new_n2734_), .ZN(new_n2735_));
  AOI22_X1   g02543(.A1(new_n2735_), .A2(new_n2467_), .B1(\asqrt[45] ), .B2(new_n2733_), .ZN(new_n2736_));
  OAI21_X1   g02544(.A1(new_n2710_), .A2(new_n2720_), .B(new_n2729_), .ZN(new_n2737_));
  AOI21_X1   g02545(.A1(new_n2737_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n2738_));
  AOI21_X1   g02546(.A1(new_n2738_), .A2(new_n2731_), .B(new_n2736_), .ZN(new_n2739_));
  OAI21_X1   g02547(.A1(new_n2739_), .A2(new_n2732_), .B(\asqrt[52] ), .ZN(new_n2740_));
  NOR2_X1    g02548(.A1(new_n2504_), .A2(new_n2514_), .ZN(new_n2741_));
  NOR3_X1    g02549(.A1(new_n2641_), .A2(new_n2481_), .A3(new_n2741_), .ZN(new_n2742_));
  INV_X1     g02550(.I(new_n2742_), .ZN(new_n2743_));
  NOR3_X1    g02551(.A1(new_n2741_), .A2(new_n2481_), .A3(new_n2513_), .ZN(new_n2744_));
  AOI22_X1   g02552(.A1(new_n2743_), .A2(new_n2513_), .B1(\asqrt[45] ), .B2(new_n2744_), .ZN(new_n2745_));
  INV_X1     g02553(.I(new_n2745_), .ZN(new_n2746_));
  NAND2_X1   g02554(.A1(new_n2696_), .A2(new_n1806_), .ZN(new_n2747_));
  OAI21_X1   g02555(.A1(new_n2747_), .A2(new_n2719_), .B(new_n2709_), .ZN(new_n2748_));
  AOI21_X1   g02556(.A1(new_n2748_), .A2(new_n2729_), .B(new_n1612_), .ZN(new_n2749_));
  NOR2_X1    g02557(.A1(new_n2703_), .A2(\asqrt[50] ), .ZN(new_n2750_));
  AOI21_X1   g02558(.A1(new_n2750_), .A2(new_n2748_), .B(new_n2727_), .ZN(new_n2751_));
  OAI21_X1   g02559(.A1(new_n2751_), .A2(new_n2749_), .B(\asqrt[51] ), .ZN(new_n2752_));
  NAND2_X1   g02560(.A1(new_n2752_), .A2(new_n1256_), .ZN(new_n2753_));
  OAI21_X1   g02561(.A1(new_n2753_), .A2(new_n2739_), .B(new_n2746_), .ZN(new_n2754_));
  AOI21_X1   g02562(.A1(new_n2754_), .A2(new_n2740_), .B(new_n1103_), .ZN(new_n2755_));
  NOR3_X1    g02563(.A1(new_n2516_), .A2(new_n2550_), .A3(new_n2500_), .ZN(new_n2756_));
  NOR3_X1    g02564(.A1(new_n2641_), .A2(new_n2516_), .A3(new_n2550_), .ZN(new_n2757_));
  INV_X1     g02565(.I(new_n2757_), .ZN(new_n2758_));
  AOI22_X1   g02566(.A1(new_n2758_), .A2(new_n2500_), .B1(\asqrt[45] ), .B2(new_n2756_), .ZN(new_n2759_));
  INV_X1     g02567(.I(new_n2736_), .ZN(new_n2760_));
  NAND2_X1   g02568(.A1(new_n2722_), .A2(new_n1376_), .ZN(new_n2761_));
  OAI21_X1   g02569(.A1(new_n2761_), .A2(new_n2751_), .B(new_n2760_), .ZN(new_n2762_));
  AOI21_X1   g02570(.A1(new_n2762_), .A2(new_n2752_), .B(new_n1256_), .ZN(new_n2763_));
  NOR2_X1    g02571(.A1(new_n2763_), .A2(\asqrt[53] ), .ZN(new_n2764_));
  AOI21_X1   g02572(.A1(new_n2764_), .A2(new_n2754_), .B(new_n2759_), .ZN(new_n2765_));
  OAI21_X1   g02573(.A1(new_n2765_), .A2(new_n2755_), .B(\asqrt[54] ), .ZN(new_n2766_));
  NOR3_X1    g02574(.A1(new_n2641_), .A2(new_n2508_), .A3(new_n2581_), .ZN(new_n2767_));
  INV_X1     g02575(.I(new_n2767_), .ZN(new_n2768_));
  NOR3_X1    g02576(.A1(new_n2508_), .A2(new_n2530_), .A3(new_n2581_), .ZN(new_n2769_));
  AOI22_X1   g02577(.A1(new_n2768_), .A2(new_n2530_), .B1(\asqrt[45] ), .B2(new_n2769_), .ZN(new_n2770_));
  INV_X1     g02578(.I(new_n2770_), .ZN(new_n2771_));
  NOR2_X1    g02579(.A1(new_n2732_), .A2(\asqrt[52] ), .ZN(new_n2772_));
  AOI21_X1   g02580(.A1(new_n2772_), .A2(new_n2762_), .B(new_n2745_), .ZN(new_n2773_));
  OAI21_X1   g02581(.A1(new_n2773_), .A2(new_n2763_), .B(\asqrt[53] ), .ZN(new_n2774_));
  NAND2_X1   g02582(.A1(new_n2774_), .A2(new_n904_), .ZN(new_n2775_));
  OAI21_X1   g02583(.A1(new_n2775_), .A2(new_n2765_), .B(new_n2771_), .ZN(new_n2776_));
  AOI21_X1   g02584(.A1(new_n2776_), .A2(new_n2766_), .B(new_n823_), .ZN(new_n2777_));
  AND3_X2    g02585(.A1(new_n2519_), .A2(new_n2524_), .A3(new_n2533_), .Z(new_n2778_));
  NAND3_X1   g02586(.A1(\asqrt[45] ), .A2(new_n2519_), .A3(new_n2533_), .ZN(new_n2779_));
  AOI22_X1   g02587(.A1(new_n2779_), .A2(new_n2525_), .B1(\asqrt[45] ), .B2(new_n2778_), .ZN(new_n2780_));
  INV_X1     g02588(.I(new_n2759_), .ZN(new_n2781_));
  NAND2_X1   g02589(.A1(new_n2740_), .A2(new_n1103_), .ZN(new_n2782_));
  OAI21_X1   g02590(.A1(new_n2782_), .A2(new_n2773_), .B(new_n2781_), .ZN(new_n2783_));
  AOI21_X1   g02591(.A1(new_n2783_), .A2(new_n2774_), .B(new_n904_), .ZN(new_n2784_));
  NOR2_X1    g02592(.A1(new_n2784_), .A2(\asqrt[55] ), .ZN(new_n2785_));
  AOI21_X1   g02593(.A1(new_n2785_), .A2(new_n2776_), .B(new_n2780_), .ZN(new_n2786_));
  OAI21_X1   g02594(.A1(new_n2786_), .A2(new_n2777_), .B(\asqrt[56] ), .ZN(new_n2787_));
  NOR3_X1    g02595(.A1(new_n2641_), .A2(new_n2535_), .A3(new_n2584_), .ZN(new_n2788_));
  INV_X1     g02596(.I(new_n2788_), .ZN(new_n2789_));
  NOR3_X1    g02597(.A1(new_n2535_), .A2(new_n2657_), .A3(new_n2584_), .ZN(new_n2790_));
  AOI22_X1   g02598(.A1(new_n2789_), .A2(new_n2657_), .B1(\asqrt[45] ), .B2(new_n2790_), .ZN(new_n2791_));
  INV_X1     g02599(.I(new_n2791_), .ZN(new_n2792_));
  NOR3_X1    g02600(.A1(new_n2739_), .A2(new_n2732_), .A3(\asqrt[52] ), .ZN(new_n2793_));
  OAI21_X1   g02601(.A1(new_n2745_), .A2(new_n2793_), .B(new_n2740_), .ZN(new_n2794_));
  AOI21_X1   g02602(.A1(new_n2794_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n2795_));
  AOI21_X1   g02603(.A1(new_n2795_), .A2(new_n2783_), .B(new_n2770_), .ZN(new_n2796_));
  OAI21_X1   g02604(.A1(new_n2796_), .A2(new_n2784_), .B(\asqrt[55] ), .ZN(new_n2797_));
  NAND2_X1   g02605(.A1(new_n2797_), .A2(new_n703_), .ZN(new_n2798_));
  OAI21_X1   g02606(.A1(new_n2798_), .A2(new_n2786_), .B(new_n2792_), .ZN(new_n2799_));
  AOI21_X1   g02607(.A1(new_n2799_), .A2(new_n2787_), .B(new_n531_), .ZN(new_n2800_));
  INV_X1     g02608(.I(new_n2543_), .ZN(new_n2801_));
  NOR2_X1    g02609(.A1(new_n2555_), .A2(new_n2542_), .ZN(new_n2802_));
  NOR3_X1    g02610(.A1(new_n2801_), .A2(new_n2549_), .A3(new_n2802_), .ZN(new_n2803_));
  NOR3_X1    g02611(.A1(new_n2641_), .A2(new_n2801_), .A3(new_n2802_), .ZN(new_n2804_));
  INV_X1     g02612(.I(new_n2804_), .ZN(new_n2805_));
  AOI22_X1   g02613(.A1(new_n2805_), .A2(new_n2549_), .B1(\asqrt[45] ), .B2(new_n2803_), .ZN(new_n2806_));
  NOR3_X1    g02614(.A1(new_n2796_), .A2(\asqrt[55] ), .A3(new_n2784_), .ZN(new_n2807_));
  OAI21_X1   g02615(.A1(new_n2780_), .A2(new_n2807_), .B(new_n2797_), .ZN(new_n2808_));
  AOI21_X1   g02616(.A1(new_n2808_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n2809_));
  AOI21_X1   g02617(.A1(new_n2809_), .A2(new_n2799_), .B(new_n2806_), .ZN(new_n2810_));
  OAI21_X1   g02618(.A1(new_n2810_), .A2(new_n2800_), .B(\asqrt[58] ), .ZN(new_n2811_));
  NOR2_X1    g02619(.A1(new_n2559_), .A2(new_n2565_), .ZN(new_n2812_));
  NOR3_X1    g02620(.A1(new_n2641_), .A2(new_n2557_), .A3(new_n2812_), .ZN(new_n2813_));
  INV_X1     g02621(.I(new_n2813_), .ZN(new_n2814_));
  NOR3_X1    g02622(.A1(new_n2812_), .A2(new_n2557_), .A3(new_n2564_), .ZN(new_n2815_));
  AOI22_X1   g02623(.A1(new_n2814_), .A2(new_n2564_), .B1(\asqrt[45] ), .B2(new_n2815_), .ZN(new_n2816_));
  INV_X1     g02624(.I(new_n2816_), .ZN(new_n2817_));
  INV_X1     g02625(.I(new_n2780_), .ZN(new_n2818_));
  NAND2_X1   g02626(.A1(new_n2766_), .A2(new_n823_), .ZN(new_n2819_));
  OAI21_X1   g02627(.A1(new_n2819_), .A2(new_n2796_), .B(new_n2818_), .ZN(new_n2820_));
  AOI21_X1   g02628(.A1(new_n2820_), .A2(new_n2797_), .B(new_n703_), .ZN(new_n2821_));
  NOR2_X1    g02629(.A1(new_n2777_), .A2(\asqrt[56] ), .ZN(new_n2822_));
  AOI21_X1   g02630(.A1(new_n2822_), .A2(new_n2820_), .B(new_n2791_), .ZN(new_n2823_));
  OAI21_X1   g02631(.A1(new_n2823_), .A2(new_n2821_), .B(\asqrt[57] ), .ZN(new_n2824_));
  NAND2_X1   g02632(.A1(new_n2824_), .A2(new_n436_), .ZN(new_n2825_));
  OAI21_X1   g02633(.A1(new_n2825_), .A2(new_n2810_), .B(new_n2817_), .ZN(new_n2826_));
  AOI21_X1   g02634(.A1(new_n2826_), .A2(new_n2811_), .B(new_n327_), .ZN(new_n2827_));
  NOR3_X1    g02635(.A1(new_n2567_), .A2(new_n2656_), .A3(new_n2615_), .ZN(new_n2828_));
  NOR3_X1    g02636(.A1(new_n2641_), .A2(new_n2567_), .A3(new_n2615_), .ZN(new_n2829_));
  INV_X1     g02637(.I(new_n2829_), .ZN(new_n2830_));
  AOI22_X1   g02638(.A1(new_n2830_), .A2(new_n2656_), .B1(\asqrt[45] ), .B2(new_n2828_), .ZN(new_n2831_));
  INV_X1     g02639(.I(new_n2806_), .ZN(new_n2832_));
  NAND2_X1   g02640(.A1(new_n2787_), .A2(new_n531_), .ZN(new_n2833_));
  OAI21_X1   g02641(.A1(new_n2833_), .A2(new_n2823_), .B(new_n2832_), .ZN(new_n2834_));
  AOI21_X1   g02642(.A1(new_n2834_), .A2(new_n2824_), .B(new_n436_), .ZN(new_n2835_));
  NOR2_X1    g02643(.A1(new_n2835_), .A2(\asqrt[59] ), .ZN(new_n2836_));
  AOI21_X1   g02644(.A1(new_n2836_), .A2(new_n2826_), .B(new_n2831_), .ZN(new_n2837_));
  OAI21_X1   g02645(.A1(new_n2837_), .A2(new_n2827_), .B(\asqrt[60] ), .ZN(new_n2838_));
  INV_X1     g02646(.I(new_n2574_), .ZN(new_n2839_));
  NOR2_X1    g02647(.A1(new_n2589_), .A2(new_n2573_), .ZN(new_n2840_));
  NOR3_X1    g02648(.A1(new_n2641_), .A2(new_n2839_), .A3(new_n2840_), .ZN(new_n2841_));
  INV_X1     g02649(.I(new_n2841_), .ZN(new_n2842_));
  NOR3_X1    g02650(.A1(new_n2839_), .A2(new_n2580_), .A3(new_n2840_), .ZN(new_n2843_));
  AOI22_X1   g02651(.A1(new_n2842_), .A2(new_n2580_), .B1(\asqrt[45] ), .B2(new_n2843_), .ZN(new_n2844_));
  INV_X1     g02652(.I(new_n2844_), .ZN(new_n2845_));
  NOR2_X1    g02653(.A1(new_n2800_), .A2(\asqrt[58] ), .ZN(new_n2846_));
  AOI21_X1   g02654(.A1(new_n2846_), .A2(new_n2834_), .B(new_n2816_), .ZN(new_n2847_));
  OAI21_X1   g02655(.A1(new_n2847_), .A2(new_n2835_), .B(\asqrt[59] ), .ZN(new_n2848_));
  NAND2_X1   g02656(.A1(new_n2848_), .A2(new_n306_), .ZN(new_n2849_));
  OAI21_X1   g02657(.A1(new_n2849_), .A2(new_n2837_), .B(new_n2845_), .ZN(new_n2850_));
  AOI21_X1   g02658(.A1(new_n2850_), .A2(new_n2838_), .B(new_n218_), .ZN(new_n2851_));
  NOR2_X1    g02659(.A1(new_n2593_), .A2(new_n2599_), .ZN(new_n2852_));
  NOR3_X1    g02660(.A1(new_n2852_), .A2(new_n2591_), .A3(new_n2598_), .ZN(new_n2853_));
  NOR3_X1    g02661(.A1(new_n2641_), .A2(new_n2591_), .A3(new_n2852_), .ZN(new_n2854_));
  INV_X1     g02662(.I(new_n2854_), .ZN(new_n2855_));
  AOI22_X1   g02663(.A1(new_n2855_), .A2(new_n2598_), .B1(\asqrt[45] ), .B2(new_n2853_), .ZN(new_n2856_));
  INV_X1     g02664(.I(new_n2831_), .ZN(new_n2857_));
  NAND2_X1   g02665(.A1(new_n2811_), .A2(new_n327_), .ZN(new_n2858_));
  OAI21_X1   g02666(.A1(new_n2858_), .A2(new_n2847_), .B(new_n2857_), .ZN(new_n2859_));
  AOI21_X1   g02667(.A1(new_n2859_), .A2(new_n2848_), .B(new_n306_), .ZN(new_n2860_));
  NOR2_X1    g02668(.A1(new_n2860_), .A2(\asqrt[61] ), .ZN(new_n2861_));
  AOI21_X1   g02669(.A1(new_n2861_), .A2(new_n2850_), .B(new_n2856_), .ZN(new_n2862_));
  OAI21_X1   g02670(.A1(new_n2862_), .A2(new_n2851_), .B(\asqrt[62] ), .ZN(new_n2863_));
  NOR3_X1    g02671(.A1(new_n2641_), .A2(new_n2601_), .A3(new_n2630_), .ZN(new_n2864_));
  INV_X1     g02672(.I(new_n2864_), .ZN(new_n2865_));
  NOR3_X1    g02673(.A1(new_n2601_), .A2(new_n2655_), .A3(new_n2630_), .ZN(new_n2866_));
  AOI22_X1   g02674(.A1(new_n2865_), .A2(new_n2655_), .B1(\asqrt[45] ), .B2(new_n2866_), .ZN(new_n2867_));
  INV_X1     g02675(.I(new_n2867_), .ZN(new_n2868_));
  NOR3_X1    g02676(.A1(new_n2810_), .A2(\asqrt[58] ), .A3(new_n2800_), .ZN(new_n2869_));
  OAI21_X1   g02677(.A1(new_n2816_), .A2(new_n2869_), .B(new_n2811_), .ZN(new_n2870_));
  AOI21_X1   g02678(.A1(new_n2870_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n2871_));
  AOI21_X1   g02679(.A1(new_n2871_), .A2(new_n2859_), .B(new_n2844_), .ZN(new_n2872_));
  OAI21_X1   g02680(.A1(new_n2872_), .A2(new_n2860_), .B(\asqrt[61] ), .ZN(new_n2873_));
  NAND2_X1   g02681(.A1(new_n2873_), .A2(new_n207_), .ZN(new_n2874_));
  OAI21_X1   g02682(.A1(new_n2874_), .A2(new_n2862_), .B(new_n2868_), .ZN(new_n2875_));
  NAND4_X1   g02683(.A1(\asqrt[45] ), .A2(new_n2608_), .A3(new_n2613_), .A4(new_n2668_), .ZN(new_n2876_));
  NAND2_X1   g02684(.A1(new_n2608_), .A2(new_n2668_), .ZN(new_n2877_));
  OAI21_X1   g02685(.A1(new_n2641_), .A2(new_n2877_), .B(new_n2614_), .ZN(new_n2878_));
  NAND2_X1   g02686(.A1(new_n2878_), .A2(new_n2876_), .ZN(new_n2879_));
  NOR2_X1    g02687(.A1(new_n2669_), .A2(new_n2648_), .ZN(new_n2880_));
  NAND2_X1   g02688(.A1(\asqrt[45] ), .A2(new_n2880_), .ZN(new_n2881_));
  NAND3_X1   g02689(.A1(new_n2879_), .A2(new_n2683_), .A3(new_n2881_), .ZN(new_n2882_));
  AOI21_X1   g02690(.A1(new_n2875_), .A2(new_n2863_), .B(new_n2882_), .ZN(new_n2883_));
  NOR3_X1    g02691(.A1(new_n2872_), .A2(\asqrt[61] ), .A3(new_n2860_), .ZN(new_n2884_));
  OAI21_X1   g02692(.A1(new_n2856_), .A2(new_n2884_), .B(new_n2873_), .ZN(new_n2885_));
  AOI21_X1   g02693(.A1(new_n2885_), .A2(\asqrt[62] ), .B(new_n2879_), .ZN(new_n2886_));
  OAI21_X1   g02694(.A1(new_n2641_), .A2(new_n2648_), .B(new_n2669_), .ZN(new_n2887_));
  NOR2_X1    g02695(.A1(new_n2880_), .A2(new_n193_), .ZN(new_n2888_));
  NAND2_X1   g02696(.A1(new_n2887_), .A2(new_n2888_), .ZN(new_n2889_));
  INV_X1     g02697(.I(new_n2889_), .ZN(new_n2890_));
  AND3_X2    g02698(.A1(new_n2624_), .A2(new_n2622_), .A3(new_n2637_), .Z(new_n2891_));
  NAND4_X1   g02699(.A1(new_n2670_), .A2(new_n2683_), .A3(new_n2634_), .A4(new_n2891_), .ZN(new_n2892_));
  INV_X1     g02700(.I(new_n2892_), .ZN(new_n2893_));
  NOR2_X1    g02701(.A1(new_n2890_), .A2(new_n2893_), .ZN(new_n2894_));
  INV_X1     g02702(.I(new_n2894_), .ZN(new_n2895_));
  AOI21_X1   g02703(.A1(new_n2886_), .A2(new_n2875_), .B(new_n2895_), .ZN(new_n2896_));
  OAI21_X1   g02704(.A1(\asqrt[63] ), .A2(new_n2883_), .B(new_n2896_), .ZN(\asqrt[44] ));
  NOR2_X1    g02705(.A1(\a[86] ), .A2(\a[87] ), .ZN(new_n2898_));
  INV_X1     g02706(.I(new_n2898_), .ZN(new_n2899_));
  NOR2_X1    g02707(.A1(new_n2899_), .A2(\a[88] ), .ZN(new_n2900_));
  INV_X1     g02708(.I(new_n2900_), .ZN(new_n2901_));
  NAND2_X1   g02709(.A1(new_n2875_), .A2(new_n2863_), .ZN(new_n2902_));
  INV_X1     g02710(.I(new_n2882_), .ZN(new_n2903_));
  AOI21_X1   g02711(.A1(new_n2902_), .A2(new_n2903_), .B(\asqrt[63] ), .ZN(new_n2904_));
  INV_X1     g02712(.I(new_n2875_), .ZN(new_n2905_));
  INV_X1     g02713(.I(new_n2879_), .ZN(new_n2906_));
  NAND2_X1   g02714(.A1(new_n2863_), .A2(new_n2906_), .ZN(new_n2907_));
  OAI21_X1   g02715(.A1(new_n2905_), .A2(new_n2907_), .B(new_n2894_), .ZN(new_n2908_));
  OAI21_X1   g02716(.A1(new_n2904_), .A2(new_n2908_), .B(\a[88] ), .ZN(new_n2909_));
  AOI21_X1   g02717(.A1(new_n2909_), .A2(new_n2901_), .B(new_n2641_), .ZN(new_n2910_));
  INV_X1     g02718(.I(\a[88] ), .ZN(new_n2911_));
  INV_X1     g02719(.I(new_n2856_), .ZN(new_n2912_));
  NAND2_X1   g02720(.A1(new_n2838_), .A2(new_n218_), .ZN(new_n2913_));
  OAI21_X1   g02721(.A1(new_n2913_), .A2(new_n2872_), .B(new_n2912_), .ZN(new_n2914_));
  NAND3_X1   g02722(.A1(new_n2914_), .A2(new_n207_), .A3(new_n2873_), .ZN(new_n2915_));
  AOI22_X1   g02723(.A1(new_n2915_), .A2(new_n2868_), .B1(new_n2885_), .B2(\asqrt[62] ), .ZN(new_n2916_));
  OAI21_X1   g02724(.A1(new_n2916_), .A2(new_n2882_), .B(new_n193_), .ZN(new_n2917_));
  AOI21_X1   g02725(.A1(new_n2917_), .A2(new_n2896_), .B(new_n2911_), .ZN(new_n2918_));
  NAND4_X1   g02726(.A1(new_n2683_), .A2(new_n2634_), .A3(new_n2637_), .A4(new_n2901_), .ZN(new_n2919_));
  NOR2_X1    g02727(.A1(new_n2919_), .A2(new_n2646_), .ZN(new_n2920_));
  INV_X1     g02728(.I(new_n2920_), .ZN(new_n2921_));
  NOR2_X1    g02729(.A1(new_n2918_), .A2(new_n2921_), .ZN(new_n2922_));
  AOI21_X1   g02730(.A1(new_n2917_), .A2(new_n2896_), .B(new_n2643_), .ZN(new_n2923_));
  INV_X1     g02731(.I(\a[89] ), .ZN(new_n2924_));
  AOI21_X1   g02732(.A1(\asqrt[44] ), .A2(new_n2911_), .B(new_n2924_), .ZN(new_n2925_));
  NOR3_X1    g02733(.A1(new_n2922_), .A2(new_n2925_), .A3(new_n2923_), .ZN(new_n2926_));
  OAI21_X1   g02734(.A1(new_n2926_), .A2(new_n2910_), .B(\asqrt[46] ), .ZN(new_n2927_));
  OAI21_X1   g02735(.A1(new_n2904_), .A2(new_n2908_), .B(new_n2642_), .ZN(new_n2928_));
  NOR2_X1    g02736(.A1(new_n2905_), .A2(new_n2907_), .ZN(new_n2929_));
  INV_X1     g02737(.I(new_n2929_), .ZN(new_n2930_));
  NOR2_X1    g02738(.A1(new_n2893_), .A2(new_n2641_), .ZN(new_n2931_));
  NAND4_X1   g02739(.A1(new_n2930_), .A2(new_n2917_), .A3(new_n2889_), .A4(new_n2931_), .ZN(new_n2932_));
  AOI21_X1   g02740(.A1(new_n2932_), .A2(new_n2928_), .B(new_n2654_), .ZN(new_n2933_));
  INV_X1     g02741(.I(new_n2931_), .ZN(new_n2934_));
  NOR4_X1    g02742(.A1(new_n2904_), .A2(new_n2929_), .A3(new_n2890_), .A4(new_n2934_), .ZN(new_n2935_));
  NOR3_X1    g02743(.A1(new_n2935_), .A2(new_n2923_), .A3(\a[90] ), .ZN(new_n2936_));
  AOI21_X1   g02744(.A1(\asqrt[44] ), .A2(\a[88] ), .B(new_n2900_), .ZN(new_n2937_));
  OAI21_X1   g02745(.A1(new_n2937_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n2938_));
  OAI22_X1   g02746(.A1(new_n2926_), .A2(new_n2938_), .B1(new_n2933_), .B2(new_n2936_), .ZN(new_n2939_));
  AOI21_X1   g02747(.A1(new_n2939_), .A2(new_n2927_), .B(new_n2229_), .ZN(new_n2940_));
  NOR3_X1    g02748(.A1(new_n2679_), .A2(new_n2653_), .A3(new_n2674_), .ZN(new_n2941_));
  NAND3_X1   g02749(.A1(\asqrt[44] ), .A2(new_n2714_), .A3(new_n2675_), .ZN(new_n2942_));
  AOI22_X1   g02750(.A1(new_n2942_), .A2(new_n2679_), .B1(\asqrt[44] ), .B2(new_n2941_), .ZN(new_n2943_));
  OAI21_X1   g02751(.A1(new_n2918_), .A2(new_n2900_), .B(\asqrt[45] ), .ZN(new_n2944_));
  AOI21_X1   g02752(.A1(new_n2917_), .A2(new_n2896_), .B(\a[88] ), .ZN(new_n2945_));
  OAI21_X1   g02753(.A1(new_n2924_), .A2(new_n2945_), .B(new_n2928_), .ZN(new_n2946_));
  OAI21_X1   g02754(.A1(new_n2946_), .A2(new_n2922_), .B(new_n2944_), .ZN(new_n2947_));
  AOI21_X1   g02755(.A1(new_n2947_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n2948_));
  AOI21_X1   g02756(.A1(new_n2948_), .A2(new_n2939_), .B(new_n2943_), .ZN(new_n2949_));
  OAI21_X1   g02757(.A1(new_n2949_), .A2(new_n2940_), .B(\asqrt[48] ), .ZN(new_n2950_));
  INV_X1     g02758(.I(new_n2950_), .ZN(new_n2951_));
  INV_X1     g02759(.I(new_n2694_), .ZN(new_n2952_));
  NAND4_X1   g02760(.A1(\asqrt[44] ), .A2(new_n2711_), .A3(new_n2690_), .A4(new_n2952_), .ZN(new_n2953_));
  INV_X1     g02761(.I(\asqrt[44] ), .ZN(new_n2954_));
  NOR3_X1    g02762(.A1(new_n2954_), .A2(new_n2681_), .A3(new_n2694_), .ZN(new_n2955_));
  OAI21_X1   g02763(.A1(new_n2955_), .A2(new_n2690_), .B(new_n2953_), .ZN(new_n2956_));
  INV_X1     g02764(.I(new_n2956_), .ZN(new_n2957_));
  NOR3_X1    g02765(.A1(new_n2949_), .A2(new_n2940_), .A3(\asqrt[48] ), .ZN(new_n2958_));
  NOR2_X1    g02766(.A1(new_n2958_), .A2(new_n2957_), .ZN(new_n2959_));
  OAI21_X1   g02767(.A1(new_n2959_), .A2(new_n2951_), .B(\asqrt[49] ), .ZN(new_n2960_));
  NAND2_X1   g02768(.A1(new_n2718_), .A2(new_n2712_), .ZN(new_n2961_));
  NAND3_X1   g02769(.A1(\asqrt[44] ), .A2(new_n2696_), .A3(new_n2961_), .ZN(new_n2962_));
  AND3_X2    g02770(.A1(new_n2696_), .A2(new_n2699_), .A3(new_n2961_), .Z(new_n2963_));
  AOI22_X1   g02771(.A1(new_n2962_), .A2(new_n2700_), .B1(\asqrt[44] ), .B2(new_n2963_), .ZN(new_n2964_));
  INV_X1     g02772(.I(new_n2964_), .ZN(new_n2965_));
  NAND2_X1   g02773(.A1(new_n2950_), .A2(new_n1806_), .ZN(new_n2966_));
  OAI21_X1   g02774(.A1(new_n2959_), .A2(new_n2966_), .B(new_n2965_), .ZN(new_n2967_));
  AOI21_X1   g02775(.A1(new_n2967_), .A2(new_n2960_), .B(new_n1612_), .ZN(new_n2968_));
  NOR3_X1    g02776(.A1(new_n2703_), .A2(new_n2709_), .A3(new_n2720_), .ZN(new_n2969_));
  NOR3_X1    g02777(.A1(new_n2954_), .A2(new_n2703_), .A3(new_n2720_), .ZN(new_n2970_));
  INV_X1     g02778(.I(new_n2970_), .ZN(new_n2971_));
  AOI22_X1   g02779(.A1(new_n2971_), .A2(new_n2709_), .B1(\asqrt[44] ), .B2(new_n2969_), .ZN(new_n2972_));
  OAI21_X1   g02780(.A1(new_n2957_), .A2(new_n2958_), .B(new_n2950_), .ZN(new_n2973_));
  AOI21_X1   g02781(.A1(new_n2973_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n2974_));
  AOI21_X1   g02782(.A1(new_n2974_), .A2(new_n2967_), .B(new_n2972_), .ZN(new_n2975_));
  OAI21_X1   g02783(.A1(new_n2975_), .A2(new_n2968_), .B(\asqrt[51] ), .ZN(new_n2976_));
  INV_X1     g02784(.I(new_n2976_), .ZN(new_n2977_));
  NAND2_X1   g02785(.A1(new_n2750_), .A2(new_n2748_), .ZN(new_n2978_));
  NAND3_X1   g02786(.A1(\asqrt[44] ), .A2(new_n2722_), .A3(new_n2978_), .ZN(new_n2979_));
  AND3_X2    g02787(.A1(new_n2978_), .A2(new_n2722_), .A3(new_n2727_), .Z(new_n2980_));
  AOI22_X1   g02788(.A1(new_n2979_), .A2(new_n2728_), .B1(\asqrt[44] ), .B2(new_n2980_), .ZN(new_n2981_));
  NOR3_X1    g02789(.A1(new_n2975_), .A2(new_n2968_), .A3(\asqrt[51] ), .ZN(new_n2982_));
  NOR2_X1    g02790(.A1(new_n2982_), .A2(new_n2981_), .ZN(new_n2983_));
  OAI21_X1   g02791(.A1(new_n2983_), .A2(new_n2977_), .B(\asqrt[52] ), .ZN(new_n2984_));
  NOR2_X1    g02792(.A1(new_n2761_), .A2(new_n2751_), .ZN(new_n2985_));
  NOR3_X1    g02793(.A1(new_n2985_), .A2(new_n2732_), .A3(new_n2760_), .ZN(new_n2986_));
  NOR3_X1    g02794(.A1(new_n2954_), .A2(new_n2732_), .A3(new_n2985_), .ZN(new_n2987_));
  INV_X1     g02795(.I(new_n2987_), .ZN(new_n2988_));
  AOI22_X1   g02796(.A1(new_n2988_), .A2(new_n2760_), .B1(\asqrt[44] ), .B2(new_n2986_), .ZN(new_n2989_));
  INV_X1     g02797(.I(new_n2989_), .ZN(new_n2990_));
  NAND2_X1   g02798(.A1(new_n2976_), .A2(new_n1256_), .ZN(new_n2991_));
  OAI21_X1   g02799(.A1(new_n2983_), .A2(new_n2991_), .B(new_n2990_), .ZN(new_n2992_));
  AOI21_X1   g02800(.A1(new_n2992_), .A2(new_n2984_), .B(new_n1103_), .ZN(new_n2993_));
  NOR3_X1    g02801(.A1(new_n2954_), .A2(new_n2763_), .A3(new_n2793_), .ZN(new_n2994_));
  INV_X1     g02802(.I(new_n2994_), .ZN(new_n2995_));
  NOR3_X1    g02803(.A1(new_n2763_), .A2(new_n2746_), .A3(new_n2793_), .ZN(new_n2996_));
  AOI22_X1   g02804(.A1(new_n2995_), .A2(new_n2746_), .B1(\asqrt[44] ), .B2(new_n2996_), .ZN(new_n2997_));
  OAI21_X1   g02805(.A1(new_n2981_), .A2(new_n2982_), .B(new_n2976_), .ZN(new_n2998_));
  AOI21_X1   g02806(.A1(new_n2998_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n2999_));
  AOI21_X1   g02807(.A1(new_n2999_), .A2(new_n2992_), .B(new_n2997_), .ZN(new_n3000_));
  OAI21_X1   g02808(.A1(new_n3000_), .A2(new_n2993_), .B(\asqrt[54] ), .ZN(new_n3001_));
  INV_X1     g02809(.I(new_n3001_), .ZN(new_n3002_));
  NAND3_X1   g02810(.A1(new_n2754_), .A2(new_n1103_), .A3(new_n2740_), .ZN(new_n3003_));
  AND3_X2    g02811(.A1(new_n3003_), .A2(new_n2774_), .A3(new_n2759_), .Z(new_n3004_));
  NAND3_X1   g02812(.A1(\asqrt[44] ), .A2(new_n2774_), .A3(new_n3003_), .ZN(new_n3005_));
  AOI22_X1   g02813(.A1(new_n3005_), .A2(new_n2781_), .B1(\asqrt[44] ), .B2(new_n3004_), .ZN(new_n3006_));
  NOR3_X1    g02814(.A1(new_n3000_), .A2(new_n2993_), .A3(\asqrt[54] ), .ZN(new_n3007_));
  NOR2_X1    g02815(.A1(new_n3007_), .A2(new_n3006_), .ZN(new_n3008_));
  OAI21_X1   g02816(.A1(new_n3008_), .A2(new_n3002_), .B(\asqrt[55] ), .ZN(new_n3009_));
  NOR2_X1    g02817(.A1(new_n2775_), .A2(new_n2765_), .ZN(new_n3010_));
  NOR3_X1    g02818(.A1(new_n2954_), .A2(new_n2784_), .A3(new_n3010_), .ZN(new_n3011_));
  INV_X1     g02819(.I(new_n3011_), .ZN(new_n3012_));
  NOR3_X1    g02820(.A1(new_n3010_), .A2(new_n2784_), .A3(new_n2771_), .ZN(new_n3013_));
  AOI22_X1   g02821(.A1(new_n3012_), .A2(new_n2771_), .B1(\asqrt[44] ), .B2(new_n3013_), .ZN(new_n3014_));
  INV_X1     g02822(.I(new_n3014_), .ZN(new_n3015_));
  NAND2_X1   g02823(.A1(new_n3001_), .A2(new_n823_), .ZN(new_n3016_));
  OAI21_X1   g02824(.A1(new_n3008_), .A2(new_n3016_), .B(new_n3015_), .ZN(new_n3017_));
  AOI21_X1   g02825(.A1(new_n3017_), .A2(new_n3009_), .B(new_n703_), .ZN(new_n3018_));
  NOR3_X1    g02826(.A1(new_n2777_), .A2(new_n2807_), .A3(new_n2818_), .ZN(new_n3019_));
  NOR3_X1    g02827(.A1(new_n2954_), .A2(new_n2777_), .A3(new_n2807_), .ZN(new_n3020_));
  INV_X1     g02828(.I(new_n3020_), .ZN(new_n3021_));
  AOI22_X1   g02829(.A1(new_n3021_), .A2(new_n2818_), .B1(\asqrt[44] ), .B2(new_n3019_), .ZN(new_n3022_));
  OAI21_X1   g02830(.A1(new_n3006_), .A2(new_n3007_), .B(new_n3001_), .ZN(new_n3023_));
  AOI21_X1   g02831(.A1(new_n3023_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n3024_));
  AOI21_X1   g02832(.A1(new_n3024_), .A2(new_n3017_), .B(new_n3022_), .ZN(new_n3025_));
  OAI21_X1   g02833(.A1(new_n3025_), .A2(new_n3018_), .B(\asqrt[57] ), .ZN(new_n3026_));
  NAND2_X1   g02834(.A1(new_n2822_), .A2(new_n2820_), .ZN(new_n3027_));
  INV_X1     g02835(.I(new_n3027_), .ZN(new_n3028_));
  NOR3_X1    g02836(.A1(new_n2954_), .A2(new_n2821_), .A3(new_n3028_), .ZN(new_n3029_));
  INV_X1     g02837(.I(new_n3029_), .ZN(new_n3030_));
  NOR3_X1    g02838(.A1(new_n3028_), .A2(new_n2821_), .A3(new_n2792_), .ZN(new_n3031_));
  AOI22_X1   g02839(.A1(new_n3030_), .A2(new_n2792_), .B1(\asqrt[44] ), .B2(new_n3031_), .ZN(new_n3032_));
  INV_X1     g02840(.I(new_n3032_), .ZN(new_n3033_));
  INV_X1     g02841(.I(new_n3006_), .ZN(new_n3034_));
  INV_X1     g02842(.I(new_n2981_), .ZN(new_n3035_));
  NAND2_X1   g02843(.A1(new_n2909_), .A2(new_n2920_), .ZN(new_n3036_));
  OAI21_X1   g02844(.A1(new_n2904_), .A2(new_n2908_), .B(new_n2911_), .ZN(new_n3037_));
  NAND2_X1   g02845(.A1(new_n3037_), .A2(\a[89] ), .ZN(new_n3038_));
  NAND3_X1   g02846(.A1(new_n3036_), .A2(new_n3038_), .A3(new_n2928_), .ZN(new_n3039_));
  AOI21_X1   g02847(.A1(new_n3039_), .A2(new_n2944_), .B(new_n2465_), .ZN(new_n3040_));
  OAI21_X1   g02848(.A1(new_n2935_), .A2(new_n2923_), .B(\a[90] ), .ZN(new_n3041_));
  NAND3_X1   g02849(.A1(new_n2932_), .A2(new_n2928_), .A3(new_n2654_), .ZN(new_n3042_));
  NAND2_X1   g02850(.A1(new_n2909_), .A2(new_n2901_), .ZN(new_n3043_));
  AOI21_X1   g02851(.A1(new_n3043_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n3044_));
  AOI22_X1   g02852(.A1(new_n3039_), .A2(new_n3044_), .B1(new_n3041_), .B2(new_n3042_), .ZN(new_n3045_));
  OAI21_X1   g02853(.A1(new_n3045_), .A2(new_n3040_), .B(\asqrt[47] ), .ZN(new_n3046_));
  NAND2_X1   g02854(.A1(new_n3046_), .A2(new_n1956_), .ZN(new_n3047_));
  OAI21_X1   g02855(.A1(new_n3047_), .A2(new_n2949_), .B(new_n2956_), .ZN(new_n3048_));
  AOI21_X1   g02856(.A1(new_n3048_), .A2(new_n2950_), .B(new_n1806_), .ZN(new_n3049_));
  INV_X1     g02857(.I(new_n2943_), .ZN(new_n3050_));
  AOI21_X1   g02858(.A1(\a[89] ), .A2(new_n3037_), .B(new_n2923_), .ZN(new_n3051_));
  AOI21_X1   g02859(.A1(new_n3051_), .A2(new_n3036_), .B(new_n2910_), .ZN(new_n3052_));
  OAI21_X1   g02860(.A1(new_n3052_), .A2(new_n2465_), .B(new_n2229_), .ZN(new_n3053_));
  OAI21_X1   g02861(.A1(new_n3053_), .A2(new_n3045_), .B(new_n3050_), .ZN(new_n3054_));
  NAND2_X1   g02862(.A1(new_n3054_), .A2(new_n3046_), .ZN(new_n3055_));
  AOI21_X1   g02863(.A1(new_n3055_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n3056_));
  AOI21_X1   g02864(.A1(new_n3056_), .A2(new_n3048_), .B(new_n2964_), .ZN(new_n3057_));
  OAI21_X1   g02865(.A1(new_n3057_), .A2(new_n3049_), .B(\asqrt[50] ), .ZN(new_n3058_));
  NAND2_X1   g02866(.A1(new_n3058_), .A2(new_n1376_), .ZN(new_n3059_));
  OAI21_X1   g02867(.A1(new_n3059_), .A2(new_n2975_), .B(new_n3035_), .ZN(new_n3060_));
  NAND3_X1   g02868(.A1(new_n3060_), .A2(new_n1256_), .A3(new_n2976_), .ZN(new_n3061_));
  AOI22_X1   g02869(.A1(new_n3061_), .A2(new_n2990_), .B1(new_n2998_), .B2(\asqrt[52] ), .ZN(new_n3062_));
  OAI21_X1   g02870(.A1(new_n3062_), .A2(new_n1103_), .B(new_n904_), .ZN(new_n3063_));
  OAI21_X1   g02871(.A1(new_n3063_), .A2(new_n3000_), .B(new_n3034_), .ZN(new_n3064_));
  AOI21_X1   g02872(.A1(new_n3064_), .A2(new_n3001_), .B(new_n823_), .ZN(new_n3065_));
  AOI21_X1   g02873(.A1(new_n3060_), .A2(new_n2976_), .B(new_n1256_), .ZN(new_n3066_));
  NOR3_X1    g02874(.A1(new_n3057_), .A2(new_n3049_), .A3(\asqrt[50] ), .ZN(new_n3067_));
  OAI21_X1   g02875(.A1(new_n2972_), .A2(new_n3067_), .B(new_n3058_), .ZN(new_n3068_));
  AOI21_X1   g02876(.A1(new_n3068_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n3069_));
  AOI21_X1   g02877(.A1(new_n3069_), .A2(new_n3060_), .B(new_n2989_), .ZN(new_n3070_));
  NOR3_X1    g02878(.A1(new_n3070_), .A2(\asqrt[53] ), .A3(new_n3066_), .ZN(new_n3071_));
  OAI22_X1   g02879(.A1(new_n3071_), .A2(new_n2997_), .B1(new_n3062_), .B2(new_n1103_), .ZN(new_n3072_));
  AOI21_X1   g02880(.A1(new_n3072_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n3073_));
  AOI21_X1   g02881(.A1(new_n3073_), .A2(new_n3064_), .B(new_n3014_), .ZN(new_n3074_));
  OAI21_X1   g02882(.A1(new_n3074_), .A2(new_n3065_), .B(\asqrt[56] ), .ZN(new_n3075_));
  NAND2_X1   g02883(.A1(new_n3075_), .A2(new_n531_), .ZN(new_n3076_));
  OAI21_X1   g02884(.A1(new_n3076_), .A2(new_n3025_), .B(new_n3033_), .ZN(new_n3077_));
  AOI21_X1   g02885(.A1(new_n3077_), .A2(new_n3026_), .B(new_n436_), .ZN(new_n3078_));
  NOR2_X1    g02886(.A1(new_n2833_), .A2(new_n2823_), .ZN(new_n3079_));
  NOR3_X1    g02887(.A1(new_n3079_), .A2(new_n2800_), .A3(new_n2832_), .ZN(new_n3080_));
  NOR3_X1    g02888(.A1(new_n2954_), .A2(new_n2800_), .A3(new_n3079_), .ZN(new_n3081_));
  INV_X1     g02889(.I(new_n3081_), .ZN(new_n3082_));
  AOI22_X1   g02890(.A1(new_n3082_), .A2(new_n2832_), .B1(\asqrt[44] ), .B2(new_n3080_), .ZN(new_n3083_));
  NOR3_X1    g02891(.A1(new_n3074_), .A2(\asqrt[56] ), .A3(new_n3065_), .ZN(new_n3084_));
  OAI21_X1   g02892(.A1(new_n3022_), .A2(new_n3084_), .B(new_n3075_), .ZN(new_n3085_));
  AOI21_X1   g02893(.A1(new_n3085_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n3086_));
  AOI21_X1   g02894(.A1(new_n3086_), .A2(new_n3077_), .B(new_n3083_), .ZN(new_n3087_));
  OAI21_X1   g02895(.A1(new_n3087_), .A2(new_n3078_), .B(\asqrt[59] ), .ZN(new_n3088_));
  NOR3_X1    g02896(.A1(new_n2954_), .A2(new_n2835_), .A3(new_n2869_), .ZN(new_n3089_));
  INV_X1     g02897(.I(new_n3089_), .ZN(new_n3090_));
  NOR3_X1    g02898(.A1(new_n2835_), .A2(new_n2869_), .A3(new_n2817_), .ZN(new_n3091_));
  AOI22_X1   g02899(.A1(new_n3090_), .A2(new_n2817_), .B1(\asqrt[44] ), .B2(new_n3091_), .ZN(new_n3092_));
  INV_X1     g02900(.I(new_n3092_), .ZN(new_n3093_));
  INV_X1     g02901(.I(new_n3026_), .ZN(new_n3094_));
  NOR3_X1    g02902(.A1(new_n3025_), .A2(new_n3018_), .A3(\asqrt[57] ), .ZN(new_n3095_));
  NOR2_X1    g02903(.A1(new_n3095_), .A2(new_n3032_), .ZN(new_n3096_));
  OAI21_X1   g02904(.A1(new_n3096_), .A2(new_n3094_), .B(\asqrt[58] ), .ZN(new_n3097_));
  NAND2_X1   g02905(.A1(new_n3097_), .A2(new_n327_), .ZN(new_n3098_));
  OAI21_X1   g02906(.A1(new_n3098_), .A2(new_n3087_), .B(new_n3093_), .ZN(new_n3099_));
  AOI21_X1   g02907(.A1(new_n3099_), .A2(new_n3088_), .B(new_n306_), .ZN(new_n3100_));
  NOR2_X1    g02908(.A1(new_n2858_), .A2(new_n2847_), .ZN(new_n3101_));
  NOR3_X1    g02909(.A1(new_n2827_), .A2(new_n3101_), .A3(new_n2857_), .ZN(new_n3102_));
  NOR3_X1    g02910(.A1(new_n2954_), .A2(new_n2827_), .A3(new_n3101_), .ZN(new_n3103_));
  INV_X1     g02911(.I(new_n3103_), .ZN(new_n3104_));
  AOI22_X1   g02912(.A1(new_n3104_), .A2(new_n2857_), .B1(\asqrt[44] ), .B2(new_n3102_), .ZN(new_n3105_));
  INV_X1     g02913(.I(new_n3083_), .ZN(new_n3106_));
  NAND2_X1   g02914(.A1(new_n3026_), .A2(new_n436_), .ZN(new_n3107_));
  OAI21_X1   g02915(.A1(new_n3096_), .A2(new_n3107_), .B(new_n3106_), .ZN(new_n3108_));
  AOI21_X1   g02916(.A1(new_n3108_), .A2(new_n3097_), .B(new_n327_), .ZN(new_n3109_));
  NOR2_X1    g02917(.A1(new_n3109_), .A2(\asqrt[60] ), .ZN(new_n3110_));
  AOI21_X1   g02918(.A1(new_n3110_), .A2(new_n3099_), .B(new_n3105_), .ZN(new_n3111_));
  OAI21_X1   g02919(.A1(new_n3111_), .A2(new_n3100_), .B(\asqrt[61] ), .ZN(new_n3112_));
  NOR2_X1    g02920(.A1(new_n2849_), .A2(new_n2837_), .ZN(new_n3113_));
  NOR3_X1    g02921(.A1(new_n2954_), .A2(new_n2860_), .A3(new_n3113_), .ZN(new_n3114_));
  INV_X1     g02922(.I(new_n3114_), .ZN(new_n3115_));
  NOR3_X1    g02923(.A1(new_n3113_), .A2(new_n2860_), .A3(new_n2845_), .ZN(new_n3116_));
  AOI22_X1   g02924(.A1(new_n3115_), .A2(new_n2845_), .B1(\asqrt[44] ), .B2(new_n3116_), .ZN(new_n3117_));
  INV_X1     g02925(.I(new_n3117_), .ZN(new_n3118_));
  OAI21_X1   g02926(.A1(new_n3032_), .A2(new_n3095_), .B(new_n3026_), .ZN(new_n3119_));
  AOI21_X1   g02927(.A1(new_n3119_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n3120_));
  AOI21_X1   g02928(.A1(new_n3120_), .A2(new_n3108_), .B(new_n3092_), .ZN(new_n3121_));
  OAI21_X1   g02929(.A1(new_n3121_), .A2(new_n3109_), .B(\asqrt[60] ), .ZN(new_n3122_));
  NAND2_X1   g02930(.A1(new_n3122_), .A2(new_n218_), .ZN(new_n3123_));
  OAI21_X1   g02931(.A1(new_n3123_), .A2(new_n3111_), .B(new_n3118_), .ZN(new_n3124_));
  AOI21_X1   g02932(.A1(new_n3124_), .A2(new_n3112_), .B(new_n207_), .ZN(new_n3125_));
  NOR3_X1    g02933(.A1(new_n2851_), .A2(new_n2884_), .A3(new_n2912_), .ZN(new_n3126_));
  NOR3_X1    g02934(.A1(new_n2954_), .A2(new_n2851_), .A3(new_n2884_), .ZN(new_n3127_));
  INV_X1     g02935(.I(new_n3127_), .ZN(new_n3128_));
  AOI22_X1   g02936(.A1(new_n3128_), .A2(new_n2912_), .B1(\asqrt[44] ), .B2(new_n3126_), .ZN(new_n3129_));
  NOR3_X1    g02937(.A1(new_n3121_), .A2(new_n3109_), .A3(\asqrt[60] ), .ZN(new_n3130_));
  OAI21_X1   g02938(.A1(new_n3105_), .A2(new_n3130_), .B(new_n3122_), .ZN(new_n3131_));
  AOI21_X1   g02939(.A1(new_n3131_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n3132_));
  AOI21_X1   g02940(.A1(new_n3132_), .A2(new_n3124_), .B(new_n3129_), .ZN(new_n3133_));
  AND3_X2    g02941(.A1(new_n2863_), .A2(new_n2915_), .A3(new_n2867_), .Z(new_n3134_));
  NAND2_X1   g02942(.A1(\asqrt[44] ), .A2(new_n3134_), .ZN(new_n3135_));
  INV_X1     g02943(.I(new_n3135_), .ZN(new_n3136_));
  AND2_X2    g02944(.A1(new_n2863_), .A2(new_n2915_), .Z(new_n3137_));
  AOI21_X1   g02945(.A1(\asqrt[44] ), .A2(new_n3137_), .B(new_n2867_), .ZN(new_n3138_));
  NOR2_X1    g02946(.A1(new_n3136_), .A2(new_n3138_), .ZN(new_n3139_));
  NOR3_X1    g02947(.A1(new_n2954_), .A2(new_n2916_), .A3(new_n2906_), .ZN(new_n3140_));
  NOR3_X1    g02948(.A1(new_n3139_), .A2(new_n2929_), .A3(new_n3140_), .ZN(new_n3141_));
  OAI21_X1   g02949(.A1(new_n3133_), .A2(new_n3125_), .B(new_n3141_), .ZN(new_n3142_));
  NAND2_X1   g02950(.A1(new_n3142_), .A2(new_n193_), .ZN(new_n3143_));
  INV_X1     g02951(.I(new_n3129_), .ZN(new_n3144_));
  NAND3_X1   g02952(.A1(new_n3124_), .A2(new_n3112_), .A3(new_n207_), .ZN(new_n3145_));
  NAND2_X1   g02953(.A1(new_n3145_), .A2(new_n3144_), .ZN(new_n3146_));
  INV_X1     g02954(.I(new_n3139_), .ZN(new_n3147_));
  NOR2_X1    g02955(.A1(new_n3125_), .A2(new_n3147_), .ZN(new_n3148_));
  AOI21_X1   g02956(.A1(\asqrt[44] ), .A2(new_n2879_), .B(new_n2902_), .ZN(new_n3149_));
  OAI21_X1   g02957(.A1(new_n2916_), .A2(new_n2906_), .B(\asqrt[63] ), .ZN(new_n3150_));
  NOR2_X1    g02958(.A1(new_n3149_), .A2(new_n3150_), .ZN(new_n3151_));
  AND3_X2    g02959(.A1(new_n2878_), .A2(new_n2876_), .A3(new_n2892_), .Z(new_n3152_));
  NAND4_X1   g02960(.A1(new_n2930_), .A2(new_n2917_), .A3(new_n2889_), .A4(new_n3152_), .ZN(new_n3153_));
  INV_X1     g02961(.I(new_n3153_), .ZN(new_n3154_));
  NOR2_X1    g02962(.A1(new_n3151_), .A2(new_n3154_), .ZN(new_n3155_));
  INV_X1     g02963(.I(new_n3155_), .ZN(new_n3156_));
  AOI21_X1   g02964(.A1(new_n3148_), .A2(new_n3146_), .B(new_n3156_), .ZN(new_n3157_));
  NAND2_X1   g02965(.A1(new_n3143_), .A2(new_n3157_), .ZN(\asqrt[43] ));
  NOR2_X1    g02966(.A1(\a[84] ), .A2(\a[85] ), .ZN(new_n3159_));
  INV_X1     g02967(.I(new_n3159_), .ZN(new_n3160_));
  NOR2_X1    g02968(.A1(new_n3160_), .A2(\a[86] ), .ZN(new_n3161_));
  INV_X1     g02969(.I(new_n3161_), .ZN(new_n3162_));
  INV_X1     g02970(.I(new_n3105_), .ZN(new_n3163_));
  NAND2_X1   g02971(.A1(new_n3088_), .A2(new_n306_), .ZN(new_n3164_));
  OAI21_X1   g02972(.A1(new_n3164_), .A2(new_n3121_), .B(new_n3163_), .ZN(new_n3165_));
  AOI21_X1   g02973(.A1(new_n3165_), .A2(new_n3122_), .B(new_n218_), .ZN(new_n3166_));
  NOR3_X1    g02974(.A1(new_n3087_), .A2(\asqrt[59] ), .A3(new_n3078_), .ZN(new_n3167_));
  OAI21_X1   g02975(.A1(new_n3092_), .A2(new_n3167_), .B(new_n3088_), .ZN(new_n3168_));
  AOI21_X1   g02976(.A1(new_n3168_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n3169_));
  AOI21_X1   g02977(.A1(new_n3169_), .A2(new_n3165_), .B(new_n3117_), .ZN(new_n3170_));
  OAI21_X1   g02978(.A1(new_n3170_), .A2(new_n3166_), .B(\asqrt[62] ), .ZN(new_n3171_));
  NOR3_X1    g02979(.A1(new_n3170_), .A2(\asqrt[62] ), .A3(new_n3166_), .ZN(new_n3172_));
  OAI21_X1   g02980(.A1(new_n3129_), .A2(new_n3172_), .B(new_n3171_), .ZN(new_n3173_));
  AOI21_X1   g02981(.A1(new_n3173_), .A2(new_n3141_), .B(\asqrt[63] ), .ZN(new_n3174_));
  NAND2_X1   g02982(.A1(new_n3171_), .A2(new_n3139_), .ZN(new_n3175_));
  OAI21_X1   g02983(.A1(new_n3175_), .A2(new_n3133_), .B(new_n3155_), .ZN(new_n3176_));
  OAI21_X1   g02984(.A1(new_n3174_), .A2(new_n3176_), .B(\a[86] ), .ZN(new_n3177_));
  AOI21_X1   g02985(.A1(new_n3177_), .A2(new_n3162_), .B(new_n2954_), .ZN(new_n3178_));
  INV_X1     g02986(.I(\a[86] ), .ZN(new_n3179_));
  AOI21_X1   g02987(.A1(new_n3143_), .A2(new_n3157_), .B(new_n3179_), .ZN(new_n3180_));
  NAND2_X1   g02988(.A1(new_n2892_), .A2(new_n3162_), .ZN(new_n3181_));
  NOR4_X1    g02989(.A1(new_n2904_), .A2(new_n2929_), .A3(new_n2890_), .A4(new_n3181_), .ZN(new_n3182_));
  INV_X1     g02990(.I(new_n3182_), .ZN(new_n3183_));
  NOR2_X1    g02991(.A1(new_n3180_), .A2(new_n3183_), .ZN(new_n3184_));
  AOI21_X1   g02992(.A1(new_n3143_), .A2(new_n3157_), .B(new_n2899_), .ZN(new_n3185_));
  INV_X1     g02993(.I(\a[87] ), .ZN(new_n3186_));
  AOI21_X1   g02994(.A1(\asqrt[43] ), .A2(new_n3179_), .B(new_n3186_), .ZN(new_n3187_));
  NOR3_X1    g02995(.A1(new_n3184_), .A2(new_n3187_), .A3(new_n3185_), .ZN(new_n3188_));
  OAI21_X1   g02996(.A1(new_n3188_), .A2(new_n3178_), .B(\asqrt[45] ), .ZN(new_n3189_));
  OAI21_X1   g02997(.A1(new_n3174_), .A2(new_n3176_), .B(new_n2898_), .ZN(new_n3190_));
  NAND2_X1   g02998(.A1(new_n3148_), .A2(new_n3146_), .ZN(new_n3191_));
  INV_X1     g02999(.I(new_n3151_), .ZN(new_n3192_));
  NOR2_X1    g03000(.A1(new_n3154_), .A2(new_n2954_), .ZN(new_n3193_));
  NAND4_X1   g03001(.A1(new_n3143_), .A2(new_n3191_), .A3(new_n3192_), .A4(new_n3193_), .ZN(new_n3194_));
  AOI21_X1   g03002(.A1(new_n3194_), .A2(new_n3190_), .B(new_n2911_), .ZN(new_n3195_));
  INV_X1     g03003(.I(new_n3191_), .ZN(new_n3196_));
  NAND2_X1   g03004(.A1(new_n3192_), .A2(new_n3193_), .ZN(new_n3197_));
  NOR3_X1    g03005(.A1(new_n3196_), .A2(new_n3174_), .A3(new_n3197_), .ZN(new_n3198_));
  NOR3_X1    g03006(.A1(new_n3198_), .A2(new_n3185_), .A3(\a[88] ), .ZN(new_n3199_));
  OAI21_X1   g03007(.A1(new_n3180_), .A2(new_n3161_), .B(\asqrt[44] ), .ZN(new_n3200_));
  NAND2_X1   g03008(.A1(new_n3200_), .A2(new_n2641_), .ZN(new_n3201_));
  OAI22_X1   g03009(.A1(new_n3188_), .A2(new_n3201_), .B1(new_n3195_), .B2(new_n3199_), .ZN(new_n3202_));
  AOI21_X1   g03010(.A1(new_n3202_), .A2(new_n3189_), .B(new_n2465_), .ZN(new_n3203_));
  NOR3_X1    g03011(.A1(new_n3051_), .A2(new_n2910_), .A3(new_n2922_), .ZN(new_n3204_));
  NAND3_X1   g03012(.A1(\asqrt[43] ), .A2(new_n2944_), .A3(new_n3036_), .ZN(new_n3205_));
  AOI22_X1   g03013(.A1(new_n3205_), .A2(new_n3051_), .B1(\asqrt[43] ), .B2(new_n3204_), .ZN(new_n3206_));
  AOI21_X1   g03014(.A1(new_n3143_), .A2(new_n3157_), .B(\a[86] ), .ZN(new_n3207_));
  OAI21_X1   g03015(.A1(new_n3186_), .A2(new_n3207_), .B(new_n3190_), .ZN(new_n3208_));
  OAI21_X1   g03016(.A1(new_n3208_), .A2(new_n3184_), .B(new_n3200_), .ZN(new_n3209_));
  AOI21_X1   g03017(.A1(new_n3209_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n3210_));
  AOI21_X1   g03018(.A1(new_n3210_), .A2(new_n3202_), .B(new_n3206_), .ZN(new_n3211_));
  OAI21_X1   g03019(.A1(new_n3211_), .A2(new_n3203_), .B(\asqrt[47] ), .ZN(new_n3212_));
  INV_X1     g03020(.I(new_n3212_), .ZN(new_n3213_));
  NOR2_X1    g03021(.A1(new_n2933_), .A2(new_n2936_), .ZN(new_n3214_));
  NOR2_X1    g03022(.A1(new_n2926_), .A2(new_n2938_), .ZN(new_n3215_));
  INV_X1     g03023(.I(new_n3215_), .ZN(new_n3216_));
  NAND4_X1   g03024(.A1(\asqrt[43] ), .A2(new_n2927_), .A3(new_n3214_), .A4(new_n3216_), .ZN(new_n3217_));
  INV_X1     g03025(.I(\asqrt[43] ), .ZN(new_n3218_));
  NOR3_X1    g03026(.A1(new_n3218_), .A2(new_n3040_), .A3(new_n3215_), .ZN(new_n3219_));
  OAI21_X1   g03027(.A1(new_n3219_), .A2(new_n3214_), .B(new_n3217_), .ZN(new_n3220_));
  INV_X1     g03028(.I(new_n3220_), .ZN(new_n3221_));
  NOR3_X1    g03029(.A1(new_n3211_), .A2(new_n3203_), .A3(\asqrt[47] ), .ZN(new_n3222_));
  NOR2_X1    g03030(.A1(new_n3222_), .A2(new_n3221_), .ZN(new_n3223_));
  OAI21_X1   g03031(.A1(new_n3223_), .A2(new_n3213_), .B(\asqrt[48] ), .ZN(new_n3224_));
  NOR2_X1    g03032(.A1(new_n3053_), .A2(new_n3045_), .ZN(new_n3225_));
  NOR3_X1    g03033(.A1(new_n3218_), .A2(new_n2940_), .A3(new_n3225_), .ZN(new_n3226_));
  INV_X1     g03034(.I(new_n3226_), .ZN(new_n3227_));
  NOR3_X1    g03035(.A1(new_n3225_), .A2(new_n2940_), .A3(new_n3050_), .ZN(new_n3228_));
  AOI22_X1   g03036(.A1(new_n3227_), .A2(new_n3050_), .B1(\asqrt[43] ), .B2(new_n3228_), .ZN(new_n3229_));
  INV_X1     g03037(.I(new_n3229_), .ZN(new_n3230_));
  NAND2_X1   g03038(.A1(new_n3212_), .A2(new_n1956_), .ZN(new_n3231_));
  OAI21_X1   g03039(.A1(new_n3223_), .A2(new_n3231_), .B(new_n3230_), .ZN(new_n3232_));
  AOI21_X1   g03040(.A1(new_n3232_), .A2(new_n3224_), .B(new_n1806_), .ZN(new_n3233_));
  NOR3_X1    g03041(.A1(new_n2951_), .A2(new_n2958_), .A3(new_n2956_), .ZN(new_n3234_));
  NOR3_X1    g03042(.A1(new_n3218_), .A2(new_n2951_), .A3(new_n2958_), .ZN(new_n3235_));
  INV_X1     g03043(.I(new_n3235_), .ZN(new_n3236_));
  AOI22_X1   g03044(.A1(new_n3236_), .A2(new_n2956_), .B1(\asqrt[43] ), .B2(new_n3234_), .ZN(new_n3237_));
  OAI21_X1   g03045(.A1(new_n3221_), .A2(new_n3222_), .B(new_n3212_), .ZN(new_n3238_));
  AOI21_X1   g03046(.A1(new_n3238_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n3239_));
  AOI21_X1   g03047(.A1(new_n3239_), .A2(new_n3232_), .B(new_n3237_), .ZN(new_n3240_));
  OAI21_X1   g03048(.A1(new_n3240_), .A2(new_n3233_), .B(\asqrt[50] ), .ZN(new_n3241_));
  NAND2_X1   g03049(.A1(new_n3056_), .A2(new_n3048_), .ZN(new_n3242_));
  NAND3_X1   g03050(.A1(\asqrt[43] ), .A2(new_n2960_), .A3(new_n3242_), .ZN(new_n3243_));
  AND3_X2    g03051(.A1(new_n2960_), .A2(new_n2964_), .A3(new_n3242_), .Z(new_n3244_));
  AOI22_X1   g03052(.A1(new_n3243_), .A2(new_n2965_), .B1(\asqrt[43] ), .B2(new_n3244_), .ZN(new_n3245_));
  INV_X1     g03053(.I(new_n3245_), .ZN(new_n3246_));
  NAND2_X1   g03054(.A1(new_n3177_), .A2(new_n3182_), .ZN(new_n3247_));
  OAI21_X1   g03055(.A1(new_n3174_), .A2(new_n3176_), .B(new_n3179_), .ZN(new_n3248_));
  NAND2_X1   g03056(.A1(new_n3248_), .A2(\a[87] ), .ZN(new_n3249_));
  NAND3_X1   g03057(.A1(new_n3247_), .A2(new_n3249_), .A3(new_n3190_), .ZN(new_n3250_));
  AOI21_X1   g03058(.A1(new_n3250_), .A2(new_n3200_), .B(new_n2641_), .ZN(new_n3251_));
  OAI21_X1   g03059(.A1(new_n3198_), .A2(new_n3185_), .B(\a[88] ), .ZN(new_n3252_));
  NAND3_X1   g03060(.A1(new_n3194_), .A2(new_n3190_), .A3(new_n2911_), .ZN(new_n3253_));
  NAND2_X1   g03061(.A1(new_n3177_), .A2(new_n3162_), .ZN(new_n3254_));
  AOI21_X1   g03062(.A1(new_n3254_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n3255_));
  AOI22_X1   g03063(.A1(new_n3250_), .A2(new_n3255_), .B1(new_n3252_), .B2(new_n3253_), .ZN(new_n3256_));
  OAI21_X1   g03064(.A1(new_n3256_), .A2(new_n3251_), .B(\asqrt[46] ), .ZN(new_n3257_));
  NAND2_X1   g03065(.A1(new_n3257_), .A2(new_n2229_), .ZN(new_n3258_));
  OAI21_X1   g03066(.A1(new_n3258_), .A2(new_n3211_), .B(new_n3220_), .ZN(new_n3259_));
  AOI21_X1   g03067(.A1(new_n3259_), .A2(new_n3212_), .B(new_n1956_), .ZN(new_n3260_));
  INV_X1     g03068(.I(new_n3206_), .ZN(new_n3261_));
  AOI21_X1   g03069(.A1(\a[87] ), .A2(new_n3248_), .B(new_n3185_), .ZN(new_n3262_));
  AOI21_X1   g03070(.A1(new_n3262_), .A2(new_n3247_), .B(new_n3178_), .ZN(new_n3263_));
  OAI21_X1   g03071(.A1(new_n3263_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n3264_));
  OAI21_X1   g03072(.A1(new_n3264_), .A2(new_n3256_), .B(new_n3261_), .ZN(new_n3265_));
  NAND2_X1   g03073(.A1(new_n3265_), .A2(new_n3257_), .ZN(new_n3266_));
  AOI21_X1   g03074(.A1(new_n3266_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n3267_));
  AOI21_X1   g03075(.A1(new_n3267_), .A2(new_n3259_), .B(new_n3229_), .ZN(new_n3268_));
  OAI21_X1   g03076(.A1(new_n3268_), .A2(new_n3260_), .B(\asqrt[49] ), .ZN(new_n3269_));
  NAND2_X1   g03077(.A1(new_n3269_), .A2(new_n1612_), .ZN(new_n3270_));
  OAI21_X1   g03078(.A1(new_n3270_), .A2(new_n3240_), .B(new_n3246_), .ZN(new_n3271_));
  AOI21_X1   g03079(.A1(new_n3271_), .A2(new_n3241_), .B(new_n1376_), .ZN(new_n3272_));
  INV_X1     g03080(.I(new_n2972_), .ZN(new_n3273_));
  NOR3_X1    g03081(.A1(new_n2968_), .A2(new_n3067_), .A3(new_n3273_), .ZN(new_n3274_));
  NOR3_X1    g03082(.A1(new_n3218_), .A2(new_n2968_), .A3(new_n3067_), .ZN(new_n3275_));
  INV_X1     g03083(.I(new_n3275_), .ZN(new_n3276_));
  AOI22_X1   g03084(.A1(new_n3276_), .A2(new_n3273_), .B1(\asqrt[43] ), .B2(new_n3274_), .ZN(new_n3277_));
  NOR3_X1    g03085(.A1(new_n3268_), .A2(new_n3260_), .A3(\asqrt[49] ), .ZN(new_n3278_));
  OAI21_X1   g03086(.A1(new_n3237_), .A2(new_n3278_), .B(new_n3269_), .ZN(new_n3279_));
  AOI21_X1   g03087(.A1(new_n3279_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n3280_));
  AOI21_X1   g03088(.A1(new_n3280_), .A2(new_n3271_), .B(new_n3277_), .ZN(new_n3281_));
  OAI21_X1   g03089(.A1(new_n3281_), .A2(new_n3272_), .B(\asqrt[52] ), .ZN(new_n3282_));
  INV_X1     g03090(.I(new_n3282_), .ZN(new_n3283_));
  INV_X1     g03091(.I(new_n3277_), .ZN(new_n3284_));
  NAND3_X1   g03092(.A1(new_n3271_), .A2(new_n1376_), .A3(new_n3241_), .ZN(new_n3285_));
  NAND2_X1   g03093(.A1(new_n3285_), .A2(new_n3284_), .ZN(new_n3286_));
  NOR3_X1    g03094(.A1(new_n3218_), .A2(new_n2977_), .A3(new_n2982_), .ZN(new_n3287_));
  INV_X1     g03095(.I(new_n3287_), .ZN(new_n3288_));
  NOR3_X1    g03096(.A1(new_n2977_), .A2(new_n3035_), .A3(new_n2982_), .ZN(new_n3289_));
  AOI22_X1   g03097(.A1(new_n3288_), .A2(new_n3035_), .B1(\asqrt[43] ), .B2(new_n3289_), .ZN(new_n3290_));
  NOR2_X1    g03098(.A1(new_n3272_), .A2(\asqrt[52] ), .ZN(new_n3291_));
  AOI21_X1   g03099(.A1(new_n3291_), .A2(new_n3286_), .B(new_n3290_), .ZN(new_n3292_));
  OAI21_X1   g03100(.A1(new_n3283_), .A2(new_n3292_), .B(\asqrt[53] ), .ZN(new_n3293_));
  INV_X1     g03101(.I(new_n3061_), .ZN(new_n3294_));
  NOR3_X1    g03102(.A1(new_n3294_), .A2(new_n3066_), .A3(new_n2990_), .ZN(new_n3295_));
  NOR3_X1    g03103(.A1(new_n3218_), .A2(new_n3066_), .A3(new_n3294_), .ZN(new_n3296_));
  INV_X1     g03104(.I(new_n3296_), .ZN(new_n3297_));
  AOI22_X1   g03105(.A1(new_n3297_), .A2(new_n2990_), .B1(\asqrt[43] ), .B2(new_n3295_), .ZN(new_n3298_));
  INV_X1     g03106(.I(new_n3298_), .ZN(new_n3299_));
  NAND2_X1   g03107(.A1(new_n3282_), .A2(new_n1103_), .ZN(new_n3300_));
  OAI21_X1   g03108(.A1(new_n3300_), .A2(new_n3292_), .B(new_n3299_), .ZN(new_n3301_));
  AOI21_X1   g03109(.A1(new_n3301_), .A2(new_n3293_), .B(new_n904_), .ZN(new_n3302_));
  INV_X1     g03110(.I(new_n3302_), .ZN(new_n3303_));
  INV_X1     g03111(.I(new_n3301_), .ZN(new_n3304_));
  INV_X1     g03112(.I(new_n2997_), .ZN(new_n3305_));
  NOR3_X1    g03113(.A1(new_n3218_), .A2(new_n2993_), .A3(new_n3071_), .ZN(new_n3306_));
  INV_X1     g03114(.I(new_n3306_), .ZN(new_n3307_));
  NOR3_X1    g03115(.A1(new_n2993_), .A2(new_n3071_), .A3(new_n3305_), .ZN(new_n3308_));
  AOI22_X1   g03116(.A1(new_n3307_), .A2(new_n3305_), .B1(\asqrt[43] ), .B2(new_n3308_), .ZN(new_n3309_));
  INV_X1     g03117(.I(new_n3309_), .ZN(new_n3310_));
  NAND2_X1   g03118(.A1(new_n3293_), .A2(new_n904_), .ZN(new_n3311_));
  OAI21_X1   g03119(.A1(new_n3311_), .A2(new_n3304_), .B(new_n3310_), .ZN(new_n3312_));
  AOI21_X1   g03120(.A1(new_n3312_), .A2(new_n3303_), .B(new_n823_), .ZN(new_n3313_));
  NOR3_X1    g03121(.A1(new_n3002_), .A2(new_n3034_), .A3(new_n3007_), .ZN(new_n3314_));
  NOR3_X1    g03122(.A1(new_n3218_), .A2(new_n3002_), .A3(new_n3007_), .ZN(new_n3315_));
  INV_X1     g03123(.I(new_n3315_), .ZN(new_n3316_));
  AOI22_X1   g03124(.A1(new_n3316_), .A2(new_n3034_), .B1(\asqrt[43] ), .B2(new_n3314_), .ZN(new_n3317_));
  NOR2_X1    g03125(.A1(new_n3302_), .A2(\asqrt[55] ), .ZN(new_n3318_));
  AOI21_X1   g03126(.A1(new_n3318_), .A2(new_n3312_), .B(new_n3317_), .ZN(new_n3319_));
  OAI21_X1   g03127(.A1(new_n3319_), .A2(new_n3313_), .B(\asqrt[56] ), .ZN(new_n3320_));
  NOR2_X1    g03128(.A1(new_n3008_), .A2(new_n3016_), .ZN(new_n3321_));
  NOR3_X1    g03129(.A1(new_n3218_), .A2(new_n3065_), .A3(new_n3321_), .ZN(new_n3322_));
  INV_X1     g03130(.I(new_n3322_), .ZN(new_n3323_));
  NOR3_X1    g03131(.A1(new_n3321_), .A2(new_n3065_), .A3(new_n3015_), .ZN(new_n3324_));
  AOI22_X1   g03132(.A1(new_n3323_), .A2(new_n3015_), .B1(\asqrt[43] ), .B2(new_n3324_), .ZN(new_n3325_));
  INV_X1     g03133(.I(new_n3325_), .ZN(new_n3326_));
  NOR3_X1    g03134(.A1(new_n3240_), .A2(new_n3233_), .A3(\asqrt[50] ), .ZN(new_n3327_));
  OAI21_X1   g03135(.A1(new_n3245_), .A2(new_n3327_), .B(new_n3241_), .ZN(new_n3328_));
  AOI22_X1   g03136(.A1(new_n3285_), .A2(new_n3284_), .B1(new_n3328_), .B2(\asqrt[51] ), .ZN(new_n3329_));
  NOR3_X1    g03137(.A1(new_n3281_), .A2(\asqrt[52] ), .A3(new_n3272_), .ZN(new_n3330_));
  OAI22_X1   g03138(.A1(new_n3330_), .A2(new_n3290_), .B1(new_n3329_), .B2(new_n1256_), .ZN(new_n3331_));
  AOI21_X1   g03139(.A1(new_n3331_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n3332_));
  AOI21_X1   g03140(.A1(new_n3332_), .A2(new_n3301_), .B(new_n3309_), .ZN(new_n3333_));
  OAI21_X1   g03141(.A1(new_n3333_), .A2(new_n3302_), .B(\asqrt[55] ), .ZN(new_n3334_));
  NAND2_X1   g03142(.A1(new_n3334_), .A2(new_n703_), .ZN(new_n3335_));
  OAI21_X1   g03143(.A1(new_n3335_), .A2(new_n3319_), .B(new_n3326_), .ZN(new_n3336_));
  AOI21_X1   g03144(.A1(new_n3336_), .A2(new_n3320_), .B(new_n531_), .ZN(new_n3337_));
  INV_X1     g03145(.I(new_n3337_), .ZN(new_n3338_));
  INV_X1     g03146(.I(new_n3336_), .ZN(new_n3339_));
  INV_X1     g03147(.I(new_n3022_), .ZN(new_n3340_));
  NOR3_X1    g03148(.A1(new_n3018_), .A2(new_n3084_), .A3(new_n3340_), .ZN(new_n3341_));
  NOR3_X1    g03149(.A1(new_n3218_), .A2(new_n3018_), .A3(new_n3084_), .ZN(new_n3342_));
  INV_X1     g03150(.I(new_n3342_), .ZN(new_n3343_));
  AOI22_X1   g03151(.A1(new_n3343_), .A2(new_n3340_), .B1(\asqrt[43] ), .B2(new_n3341_), .ZN(new_n3344_));
  INV_X1     g03152(.I(new_n3344_), .ZN(new_n3345_));
  NAND2_X1   g03153(.A1(new_n3320_), .A2(new_n531_), .ZN(new_n3346_));
  OAI21_X1   g03154(.A1(new_n3339_), .A2(new_n3346_), .B(new_n3345_), .ZN(new_n3347_));
  AOI21_X1   g03155(.A1(new_n3347_), .A2(new_n3338_), .B(new_n436_), .ZN(new_n3348_));
  NOR3_X1    g03156(.A1(new_n3218_), .A2(new_n3094_), .A3(new_n3095_), .ZN(new_n3349_));
  INV_X1     g03157(.I(new_n3349_), .ZN(new_n3350_));
  NOR3_X1    g03158(.A1(new_n3094_), .A2(new_n3033_), .A3(new_n3095_), .ZN(new_n3351_));
  AOI22_X1   g03159(.A1(new_n3350_), .A2(new_n3033_), .B1(\asqrt[43] ), .B2(new_n3351_), .ZN(new_n3352_));
  NOR2_X1    g03160(.A1(new_n3337_), .A2(\asqrt[58] ), .ZN(new_n3353_));
  AOI21_X1   g03161(.A1(new_n3353_), .A2(new_n3347_), .B(new_n3352_), .ZN(new_n3354_));
  OAI21_X1   g03162(.A1(new_n3354_), .A2(new_n3348_), .B(\asqrt[59] ), .ZN(new_n3355_));
  NOR2_X1    g03163(.A1(new_n3096_), .A2(new_n3107_), .ZN(new_n3356_));
  NOR3_X1    g03164(.A1(new_n3356_), .A2(new_n3078_), .A3(new_n3106_), .ZN(new_n3357_));
  NOR3_X1    g03165(.A1(new_n3218_), .A2(new_n3078_), .A3(new_n3356_), .ZN(new_n3358_));
  INV_X1     g03166(.I(new_n3358_), .ZN(new_n3359_));
  AOI22_X1   g03167(.A1(new_n3359_), .A2(new_n3106_), .B1(\asqrt[43] ), .B2(new_n3357_), .ZN(new_n3360_));
  INV_X1     g03168(.I(new_n3360_), .ZN(new_n3361_));
  NOR3_X1    g03169(.A1(new_n3333_), .A2(\asqrt[55] ), .A3(new_n3302_), .ZN(new_n3362_));
  OAI21_X1   g03170(.A1(new_n3317_), .A2(new_n3362_), .B(new_n3334_), .ZN(new_n3363_));
  AOI21_X1   g03171(.A1(new_n3363_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n3364_));
  AOI21_X1   g03172(.A1(new_n3364_), .A2(new_n3336_), .B(new_n3344_), .ZN(new_n3365_));
  OAI21_X1   g03173(.A1(new_n3365_), .A2(new_n3337_), .B(\asqrt[58] ), .ZN(new_n3366_));
  NAND2_X1   g03174(.A1(new_n3366_), .A2(new_n327_), .ZN(new_n3367_));
  OAI21_X1   g03175(.A1(new_n3367_), .A2(new_n3354_), .B(new_n3361_), .ZN(new_n3368_));
  AOI21_X1   g03176(.A1(new_n3368_), .A2(new_n3355_), .B(new_n306_), .ZN(new_n3369_));
  INV_X1     g03177(.I(new_n3369_), .ZN(new_n3370_));
  INV_X1     g03178(.I(new_n3368_), .ZN(new_n3371_));
  NOR3_X1    g03179(.A1(new_n3218_), .A2(new_n3109_), .A3(new_n3167_), .ZN(new_n3372_));
  INV_X1     g03180(.I(new_n3372_), .ZN(new_n3373_));
  NOR3_X1    g03181(.A1(new_n3109_), .A2(new_n3167_), .A3(new_n3093_), .ZN(new_n3374_));
  AOI22_X1   g03182(.A1(new_n3373_), .A2(new_n3093_), .B1(\asqrt[43] ), .B2(new_n3374_), .ZN(new_n3375_));
  INV_X1     g03183(.I(new_n3375_), .ZN(new_n3376_));
  NAND2_X1   g03184(.A1(new_n3355_), .A2(new_n306_), .ZN(new_n3377_));
  OAI21_X1   g03185(.A1(new_n3371_), .A2(new_n3377_), .B(new_n3376_), .ZN(new_n3378_));
  AOI21_X1   g03186(.A1(new_n3378_), .A2(new_n3370_), .B(new_n218_), .ZN(new_n3379_));
  NOR3_X1    g03187(.A1(new_n3100_), .A2(new_n3130_), .A3(new_n3163_), .ZN(new_n3380_));
  NOR3_X1    g03188(.A1(new_n3218_), .A2(new_n3100_), .A3(new_n3130_), .ZN(new_n3381_));
  INV_X1     g03189(.I(new_n3381_), .ZN(new_n3382_));
  AOI22_X1   g03190(.A1(new_n3382_), .A2(new_n3163_), .B1(\asqrt[43] ), .B2(new_n3380_), .ZN(new_n3383_));
  NOR2_X1    g03191(.A1(new_n3369_), .A2(\asqrt[61] ), .ZN(new_n3384_));
  AOI21_X1   g03192(.A1(new_n3384_), .A2(new_n3378_), .B(new_n3383_), .ZN(new_n3385_));
  OAI21_X1   g03193(.A1(new_n3385_), .A2(new_n3379_), .B(\asqrt[62] ), .ZN(new_n3386_));
  NOR2_X1    g03194(.A1(new_n3123_), .A2(new_n3111_), .ZN(new_n3387_));
  NOR3_X1    g03195(.A1(new_n3218_), .A2(new_n3166_), .A3(new_n3387_), .ZN(new_n3388_));
  INV_X1     g03196(.I(new_n3388_), .ZN(new_n3389_));
  NOR3_X1    g03197(.A1(new_n3387_), .A2(new_n3166_), .A3(new_n3118_), .ZN(new_n3390_));
  AOI22_X1   g03198(.A1(new_n3389_), .A2(new_n3118_), .B1(\asqrt[43] ), .B2(new_n3390_), .ZN(new_n3391_));
  INV_X1     g03199(.I(new_n3391_), .ZN(new_n3392_));
  NOR3_X1    g03200(.A1(new_n3365_), .A2(\asqrt[58] ), .A3(new_n3337_), .ZN(new_n3393_));
  OAI21_X1   g03201(.A1(new_n3352_), .A2(new_n3393_), .B(new_n3366_), .ZN(new_n3394_));
  AOI21_X1   g03202(.A1(new_n3394_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n3395_));
  AOI21_X1   g03203(.A1(new_n3395_), .A2(new_n3368_), .B(new_n3375_), .ZN(new_n3396_));
  OAI21_X1   g03204(.A1(new_n3396_), .A2(new_n3369_), .B(\asqrt[61] ), .ZN(new_n3397_));
  NAND2_X1   g03205(.A1(new_n3397_), .A2(new_n207_), .ZN(new_n3398_));
  OAI21_X1   g03206(.A1(new_n3398_), .A2(new_n3385_), .B(new_n3392_), .ZN(new_n3399_));
  NAND4_X1   g03207(.A1(\asqrt[43] ), .A2(new_n3171_), .A3(new_n3129_), .A4(new_n3145_), .ZN(new_n3400_));
  NAND2_X1   g03208(.A1(new_n3171_), .A2(new_n3145_), .ZN(new_n3401_));
  OAI21_X1   g03209(.A1(new_n3218_), .A2(new_n3401_), .B(new_n3144_), .ZN(new_n3402_));
  NAND2_X1   g03210(.A1(new_n3402_), .A2(new_n3400_), .ZN(new_n3403_));
  AOI21_X1   g03211(.A1(new_n3146_), .A2(new_n3171_), .B(new_n3139_), .ZN(new_n3404_));
  AOI21_X1   g03212(.A1(\asqrt[43] ), .A2(new_n3404_), .B(new_n3196_), .ZN(new_n3405_));
  NAND2_X1   g03213(.A1(new_n3403_), .A2(new_n3405_), .ZN(new_n3406_));
  AOI21_X1   g03214(.A1(new_n3399_), .A2(new_n3386_), .B(new_n3406_), .ZN(new_n3407_));
  NOR3_X1    g03215(.A1(new_n3396_), .A2(\asqrt[61] ), .A3(new_n3369_), .ZN(new_n3408_));
  OAI21_X1   g03216(.A1(new_n3383_), .A2(new_n3408_), .B(new_n3397_), .ZN(new_n3409_));
  AOI21_X1   g03217(.A1(new_n3409_), .A2(\asqrt[62] ), .B(new_n3403_), .ZN(new_n3410_));
  AOI21_X1   g03218(.A1(\asqrt[43] ), .A2(new_n3147_), .B(new_n3173_), .ZN(new_n3411_));
  OR3_X2     g03219(.A1(new_n3411_), .A2(new_n193_), .A3(new_n3404_), .Z(new_n3412_));
  NAND2_X1   g03220(.A1(new_n3135_), .A2(new_n3153_), .ZN(new_n3413_));
  NOR4_X1    g03221(.A1(new_n3196_), .A2(new_n3138_), .A3(new_n3151_), .A4(new_n3413_), .ZN(new_n3414_));
  NAND2_X1   g03222(.A1(new_n3414_), .A2(new_n3143_), .ZN(new_n3415_));
  NAND2_X1   g03223(.A1(new_n3412_), .A2(new_n3415_), .ZN(new_n3416_));
  AOI21_X1   g03224(.A1(new_n3410_), .A2(new_n3399_), .B(new_n3416_), .ZN(new_n3417_));
  OAI21_X1   g03225(.A1(\asqrt[63] ), .A2(new_n3407_), .B(new_n3417_), .ZN(\asqrt[42] ));
  INV_X1     g03226(.I(\asqrt[42] ), .ZN(new_n3419_));
  NOR2_X1    g03227(.A1(\a[82] ), .A2(\a[83] ), .ZN(new_n3420_));
  INV_X1     g03228(.I(new_n3420_), .ZN(new_n3421_));
  NOR2_X1    g03229(.A1(new_n3421_), .A2(\a[84] ), .ZN(new_n3422_));
  INV_X1     g03230(.I(\a[84] ), .ZN(new_n3423_));
  INV_X1     g03231(.I(new_n3383_), .ZN(new_n3424_));
  INV_X1     g03232(.I(new_n3352_), .ZN(new_n3425_));
  INV_X1     g03233(.I(new_n3317_), .ZN(new_n3426_));
  INV_X1     g03234(.I(new_n3290_), .ZN(new_n3427_));
  INV_X1     g03235(.I(new_n3237_), .ZN(new_n3428_));
  NAND2_X1   g03236(.A1(new_n3224_), .A2(new_n1806_), .ZN(new_n3429_));
  OAI21_X1   g03237(.A1(new_n3429_), .A2(new_n3268_), .B(new_n3428_), .ZN(new_n3430_));
  AOI21_X1   g03238(.A1(new_n3430_), .A2(new_n3269_), .B(new_n1612_), .ZN(new_n3431_));
  NOR2_X1    g03239(.A1(new_n3233_), .A2(\asqrt[50] ), .ZN(new_n3432_));
  AOI21_X1   g03240(.A1(new_n3432_), .A2(new_n3430_), .B(new_n3245_), .ZN(new_n3433_));
  OAI21_X1   g03241(.A1(new_n3433_), .A2(new_n3431_), .B(\asqrt[51] ), .ZN(new_n3434_));
  NAND2_X1   g03242(.A1(new_n3434_), .A2(new_n1256_), .ZN(new_n3435_));
  OAI21_X1   g03243(.A1(new_n3435_), .A2(new_n3281_), .B(new_n3427_), .ZN(new_n3436_));
  NAND3_X1   g03244(.A1(new_n3436_), .A2(new_n1103_), .A3(new_n3282_), .ZN(new_n3437_));
  AOI22_X1   g03245(.A1(new_n3437_), .A2(new_n3299_), .B1(\asqrt[53] ), .B2(new_n3331_), .ZN(new_n3438_));
  OAI21_X1   g03246(.A1(new_n3438_), .A2(new_n904_), .B(new_n823_), .ZN(new_n3439_));
  OAI21_X1   g03247(.A1(new_n3439_), .A2(new_n3333_), .B(new_n3426_), .ZN(new_n3440_));
  NAND3_X1   g03248(.A1(new_n3440_), .A2(new_n703_), .A3(new_n3334_), .ZN(new_n3441_));
  AOI22_X1   g03249(.A1(new_n3441_), .A2(new_n3326_), .B1(new_n3363_), .B2(\asqrt[56] ), .ZN(new_n3442_));
  OAI21_X1   g03250(.A1(new_n3442_), .A2(new_n531_), .B(new_n436_), .ZN(new_n3443_));
  OAI21_X1   g03251(.A1(new_n3443_), .A2(new_n3365_), .B(new_n3425_), .ZN(new_n3444_));
  NAND3_X1   g03252(.A1(new_n3444_), .A2(new_n327_), .A3(new_n3366_), .ZN(new_n3445_));
  AOI22_X1   g03253(.A1(new_n3445_), .A2(new_n3361_), .B1(new_n3394_), .B2(\asqrt[59] ), .ZN(new_n3446_));
  OAI21_X1   g03254(.A1(new_n3446_), .A2(new_n306_), .B(new_n218_), .ZN(new_n3447_));
  OAI21_X1   g03255(.A1(new_n3447_), .A2(new_n3396_), .B(new_n3424_), .ZN(new_n3448_));
  NAND3_X1   g03256(.A1(new_n3448_), .A2(new_n207_), .A3(new_n3397_), .ZN(new_n3449_));
  AOI22_X1   g03257(.A1(new_n3449_), .A2(new_n3392_), .B1(new_n3409_), .B2(\asqrt[62] ), .ZN(new_n3450_));
  OAI21_X1   g03258(.A1(new_n3450_), .A2(new_n3406_), .B(new_n193_), .ZN(new_n3451_));
  AOI21_X1   g03259(.A1(new_n3451_), .A2(new_n3417_), .B(new_n3423_), .ZN(new_n3452_));
  OAI21_X1   g03260(.A1(new_n3452_), .A2(new_n3422_), .B(\asqrt[43] ), .ZN(new_n3453_));
  INV_X1     g03261(.I(new_n3453_), .ZN(new_n3454_));
  NOR2_X1    g03262(.A1(new_n3154_), .A2(new_n3422_), .ZN(new_n3455_));
  NAND4_X1   g03263(.A1(new_n3143_), .A2(new_n3191_), .A3(new_n3192_), .A4(new_n3455_), .ZN(new_n3456_));
  NOR2_X1    g03264(.A1(new_n3452_), .A2(new_n3456_), .ZN(new_n3457_));
  AOI21_X1   g03265(.A1(new_n3451_), .A2(new_n3417_), .B(new_n3160_), .ZN(new_n3458_));
  INV_X1     g03266(.I(\a[85] ), .ZN(new_n3459_));
  AOI21_X1   g03267(.A1(\asqrt[42] ), .A2(new_n3423_), .B(new_n3459_), .ZN(new_n3460_));
  NOR3_X1    g03268(.A1(new_n3457_), .A2(new_n3460_), .A3(new_n3458_), .ZN(new_n3461_));
  OAI21_X1   g03269(.A1(new_n3461_), .A2(new_n3454_), .B(\asqrt[44] ), .ZN(new_n3462_));
  NOR2_X1    g03270(.A1(new_n3407_), .A2(\asqrt[63] ), .ZN(new_n3463_));
  INV_X1     g03271(.I(new_n3399_), .ZN(new_n3464_));
  INV_X1     g03272(.I(new_n3403_), .ZN(new_n3465_));
  NAND2_X1   g03273(.A1(new_n3386_), .A2(new_n3465_), .ZN(new_n3466_));
  INV_X1     g03274(.I(new_n3416_), .ZN(new_n3467_));
  OAI21_X1   g03275(.A1(new_n3464_), .A2(new_n3466_), .B(new_n3467_), .ZN(new_n3468_));
  OAI21_X1   g03276(.A1(new_n3463_), .A2(new_n3468_), .B(new_n3159_), .ZN(new_n3469_));
  NOR2_X1    g03277(.A1(new_n3464_), .A2(new_n3466_), .ZN(new_n3470_));
  OAI21_X1   g03278(.A1(new_n3414_), .A2(new_n3157_), .B(new_n3143_), .ZN(new_n3471_));
  NAND2_X1   g03279(.A1(new_n3412_), .A2(new_n3471_), .ZN(new_n3472_));
  NOR3_X1    g03280(.A1(new_n3463_), .A2(new_n3470_), .A3(new_n3472_), .ZN(new_n3473_));
  INV_X1     g03281(.I(new_n3473_), .ZN(new_n3474_));
  AOI21_X1   g03282(.A1(new_n3474_), .A2(new_n3469_), .B(new_n3179_), .ZN(new_n3475_));
  NOR3_X1    g03283(.A1(new_n3473_), .A2(new_n3458_), .A3(\a[86] ), .ZN(new_n3476_));
  AOI21_X1   g03284(.A1(\asqrt[42] ), .A2(\a[84] ), .B(new_n3422_), .ZN(new_n3477_));
  OAI21_X1   g03285(.A1(new_n3477_), .A2(new_n3218_), .B(new_n2954_), .ZN(new_n3478_));
  OAI22_X1   g03286(.A1(new_n3461_), .A2(new_n3478_), .B1(new_n3475_), .B2(new_n3476_), .ZN(new_n3479_));
  AOI21_X1   g03287(.A1(new_n3479_), .A2(new_n3462_), .B(new_n2641_), .ZN(new_n3480_));
  NOR3_X1    g03288(.A1(new_n3262_), .A2(new_n3178_), .A3(new_n3184_), .ZN(new_n3481_));
  NAND3_X1   g03289(.A1(\asqrt[42] ), .A2(new_n3200_), .A3(new_n3247_), .ZN(new_n3482_));
  AOI22_X1   g03290(.A1(new_n3482_), .A2(new_n3262_), .B1(\asqrt[42] ), .B2(new_n3481_), .ZN(new_n3483_));
  AOI21_X1   g03291(.A1(new_n3451_), .A2(new_n3417_), .B(\a[84] ), .ZN(new_n3484_));
  OAI21_X1   g03292(.A1(new_n3459_), .A2(new_n3484_), .B(new_n3469_), .ZN(new_n3485_));
  OAI21_X1   g03293(.A1(new_n3485_), .A2(new_n3457_), .B(new_n3453_), .ZN(new_n3486_));
  AOI21_X1   g03294(.A1(new_n3486_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n3487_));
  AOI21_X1   g03295(.A1(new_n3487_), .A2(new_n3479_), .B(new_n3483_), .ZN(new_n3488_));
  OAI21_X1   g03296(.A1(new_n3488_), .A2(new_n3480_), .B(\asqrt[46] ), .ZN(new_n3489_));
  INV_X1     g03297(.I(new_n3489_), .ZN(new_n3490_));
  NOR2_X1    g03298(.A1(new_n3199_), .A2(new_n3195_), .ZN(new_n3491_));
  INV_X1     g03299(.I(new_n3491_), .ZN(new_n3492_));
  NOR2_X1    g03300(.A1(new_n3188_), .A2(new_n3201_), .ZN(new_n3493_));
  NOR3_X1    g03301(.A1(new_n3251_), .A2(new_n3492_), .A3(new_n3493_), .ZN(new_n3494_));
  NOR3_X1    g03302(.A1(new_n3419_), .A2(new_n3251_), .A3(new_n3493_), .ZN(new_n3495_));
  INV_X1     g03303(.I(new_n3495_), .ZN(new_n3496_));
  AOI22_X1   g03304(.A1(new_n3496_), .A2(new_n3492_), .B1(\asqrt[42] ), .B2(new_n3494_), .ZN(new_n3497_));
  NOR3_X1    g03305(.A1(new_n3488_), .A2(new_n3480_), .A3(\asqrt[46] ), .ZN(new_n3498_));
  NOR2_X1    g03306(.A1(new_n3498_), .A2(new_n3497_), .ZN(new_n3499_));
  OAI21_X1   g03307(.A1(new_n3499_), .A2(new_n3490_), .B(\asqrt[47] ), .ZN(new_n3500_));
  NOR2_X1    g03308(.A1(new_n3264_), .A2(new_n3256_), .ZN(new_n3501_));
  NOR3_X1    g03309(.A1(new_n3419_), .A2(new_n3203_), .A3(new_n3501_), .ZN(new_n3502_));
  INV_X1     g03310(.I(new_n3502_), .ZN(new_n3503_));
  NOR3_X1    g03311(.A1(new_n3501_), .A2(new_n3203_), .A3(new_n3261_), .ZN(new_n3504_));
  AOI22_X1   g03312(.A1(new_n3503_), .A2(new_n3261_), .B1(\asqrt[42] ), .B2(new_n3504_), .ZN(new_n3505_));
  INV_X1     g03313(.I(new_n3505_), .ZN(new_n3506_));
  NAND2_X1   g03314(.A1(new_n3489_), .A2(new_n2229_), .ZN(new_n3507_));
  OAI21_X1   g03315(.A1(new_n3499_), .A2(new_n3507_), .B(new_n3506_), .ZN(new_n3508_));
  AOI21_X1   g03316(.A1(new_n3508_), .A2(new_n3500_), .B(new_n1956_), .ZN(new_n3509_));
  NOR3_X1    g03317(.A1(new_n3213_), .A2(new_n3222_), .A3(new_n3220_), .ZN(new_n3510_));
  NOR3_X1    g03318(.A1(new_n3419_), .A2(new_n3213_), .A3(new_n3222_), .ZN(new_n3511_));
  INV_X1     g03319(.I(new_n3511_), .ZN(new_n3512_));
  AOI22_X1   g03320(.A1(new_n3512_), .A2(new_n3220_), .B1(\asqrt[42] ), .B2(new_n3510_), .ZN(new_n3513_));
  OAI21_X1   g03321(.A1(new_n3497_), .A2(new_n3498_), .B(new_n3489_), .ZN(new_n3514_));
  AOI21_X1   g03322(.A1(new_n3514_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n3515_));
  AOI21_X1   g03323(.A1(new_n3515_), .A2(new_n3508_), .B(new_n3513_), .ZN(new_n3516_));
  OAI21_X1   g03324(.A1(new_n3516_), .A2(new_n3509_), .B(\asqrt[49] ), .ZN(new_n3517_));
  INV_X1     g03325(.I(new_n3517_), .ZN(new_n3518_));
  NOR2_X1    g03326(.A1(new_n3223_), .A2(new_n3231_), .ZN(new_n3519_));
  NOR3_X1    g03327(.A1(new_n3419_), .A2(new_n3260_), .A3(new_n3519_), .ZN(new_n3520_));
  INV_X1     g03328(.I(new_n3520_), .ZN(new_n3521_));
  NOR3_X1    g03329(.A1(new_n3519_), .A2(new_n3260_), .A3(new_n3230_), .ZN(new_n3522_));
  AOI22_X1   g03330(.A1(new_n3521_), .A2(new_n3230_), .B1(\asqrt[42] ), .B2(new_n3522_), .ZN(new_n3523_));
  NOR3_X1    g03331(.A1(new_n3516_), .A2(new_n3509_), .A3(\asqrt[49] ), .ZN(new_n3524_));
  NOR2_X1    g03332(.A1(new_n3524_), .A2(new_n3523_), .ZN(new_n3525_));
  OAI21_X1   g03333(.A1(new_n3525_), .A2(new_n3518_), .B(\asqrt[50] ), .ZN(new_n3526_));
  NOR3_X1    g03334(.A1(new_n3233_), .A2(new_n3278_), .A3(new_n3428_), .ZN(new_n3527_));
  NOR3_X1    g03335(.A1(new_n3419_), .A2(new_n3233_), .A3(new_n3278_), .ZN(new_n3528_));
  INV_X1     g03336(.I(new_n3528_), .ZN(new_n3529_));
  AOI22_X1   g03337(.A1(new_n3529_), .A2(new_n3428_), .B1(\asqrt[42] ), .B2(new_n3527_), .ZN(new_n3530_));
  INV_X1     g03338(.I(new_n3530_), .ZN(new_n3531_));
  NAND2_X1   g03339(.A1(new_n3517_), .A2(new_n1612_), .ZN(new_n3532_));
  OAI21_X1   g03340(.A1(new_n3525_), .A2(new_n3532_), .B(new_n3531_), .ZN(new_n3533_));
  AOI21_X1   g03341(.A1(new_n3533_), .A2(new_n3526_), .B(new_n1376_), .ZN(new_n3534_));
  NOR3_X1    g03342(.A1(new_n3419_), .A2(new_n3431_), .A3(new_n3327_), .ZN(new_n3535_));
  INV_X1     g03343(.I(new_n3535_), .ZN(new_n3536_));
  NOR3_X1    g03344(.A1(new_n3431_), .A2(new_n3246_), .A3(new_n3327_), .ZN(new_n3537_));
  AOI22_X1   g03345(.A1(new_n3536_), .A2(new_n3246_), .B1(\asqrt[42] ), .B2(new_n3537_), .ZN(new_n3538_));
  OAI21_X1   g03346(.A1(new_n3523_), .A2(new_n3524_), .B(new_n3517_), .ZN(new_n3539_));
  AOI21_X1   g03347(.A1(new_n3539_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n3540_));
  AOI21_X1   g03348(.A1(new_n3540_), .A2(new_n3533_), .B(new_n3538_), .ZN(new_n3541_));
  OAI21_X1   g03349(.A1(new_n3541_), .A2(new_n3534_), .B(\asqrt[52] ), .ZN(new_n3542_));
  AND3_X2    g03350(.A1(new_n3434_), .A2(new_n3277_), .A3(new_n3285_), .Z(new_n3543_));
  NAND3_X1   g03351(.A1(\asqrt[42] ), .A2(new_n3434_), .A3(new_n3285_), .ZN(new_n3544_));
  AOI22_X1   g03352(.A1(new_n3544_), .A2(new_n3284_), .B1(\asqrt[42] ), .B2(new_n3543_), .ZN(new_n3545_));
  INV_X1     g03353(.I(new_n3545_), .ZN(new_n3546_));
  INV_X1     g03354(.I(new_n3523_), .ZN(new_n3547_));
  OR2_X2     g03355(.A1(new_n3509_), .A2(\asqrt[49] ), .Z(new_n3548_));
  OAI21_X1   g03356(.A1(new_n3548_), .A2(new_n3516_), .B(new_n3547_), .ZN(new_n3549_));
  AOI21_X1   g03357(.A1(new_n3549_), .A2(new_n3517_), .B(new_n1612_), .ZN(new_n3550_));
  INV_X1     g03358(.I(new_n3532_), .ZN(new_n3551_));
  AOI21_X1   g03359(.A1(new_n3551_), .A2(new_n3549_), .B(new_n3530_), .ZN(new_n3552_));
  OAI21_X1   g03360(.A1(new_n3552_), .A2(new_n3550_), .B(\asqrt[51] ), .ZN(new_n3553_));
  NAND2_X1   g03361(.A1(new_n3553_), .A2(new_n1256_), .ZN(new_n3554_));
  OAI21_X1   g03362(.A1(new_n3554_), .A2(new_n3541_), .B(new_n3546_), .ZN(new_n3555_));
  AOI21_X1   g03363(.A1(new_n3555_), .A2(new_n3542_), .B(new_n1103_), .ZN(new_n3556_));
  NOR3_X1    g03364(.A1(new_n3419_), .A2(new_n3283_), .A3(new_n3330_), .ZN(new_n3557_));
  INV_X1     g03365(.I(new_n3557_), .ZN(new_n3558_));
  NOR3_X1    g03366(.A1(new_n3283_), .A2(new_n3427_), .A3(new_n3330_), .ZN(new_n3559_));
  AOI22_X1   g03367(.A1(new_n3558_), .A2(new_n3427_), .B1(\asqrt[42] ), .B2(new_n3559_), .ZN(new_n3560_));
  INV_X1     g03368(.I(new_n3538_), .ZN(new_n3561_));
  NAND2_X1   g03369(.A1(new_n3526_), .A2(new_n1376_), .ZN(new_n3562_));
  OAI21_X1   g03370(.A1(new_n3562_), .A2(new_n3552_), .B(new_n3561_), .ZN(new_n3563_));
  AOI21_X1   g03371(.A1(new_n3563_), .A2(new_n3553_), .B(new_n1256_), .ZN(new_n3564_));
  NOR2_X1    g03372(.A1(new_n3564_), .A2(\asqrt[53] ), .ZN(new_n3565_));
  AOI21_X1   g03373(.A1(new_n3565_), .A2(new_n3555_), .B(new_n3560_), .ZN(new_n3566_));
  OAI21_X1   g03374(.A1(new_n3566_), .A2(new_n3556_), .B(\asqrt[54] ), .ZN(new_n3567_));
  INV_X1     g03375(.I(new_n3293_), .ZN(new_n3568_));
  NOR2_X1    g03376(.A1(new_n3300_), .A2(new_n3292_), .ZN(new_n3569_));
  NOR3_X1    g03377(.A1(new_n3568_), .A2(new_n3299_), .A3(new_n3569_), .ZN(new_n3570_));
  NOR3_X1    g03378(.A1(new_n3419_), .A2(new_n3568_), .A3(new_n3569_), .ZN(new_n3571_));
  INV_X1     g03379(.I(new_n3571_), .ZN(new_n3572_));
  AOI22_X1   g03380(.A1(new_n3572_), .A2(new_n3299_), .B1(\asqrt[42] ), .B2(new_n3570_), .ZN(new_n3573_));
  INV_X1     g03381(.I(new_n3573_), .ZN(new_n3574_));
  NOR2_X1    g03382(.A1(new_n3534_), .A2(\asqrt[52] ), .ZN(new_n3575_));
  AOI21_X1   g03383(.A1(new_n3575_), .A2(new_n3563_), .B(new_n3545_), .ZN(new_n3576_));
  OAI21_X1   g03384(.A1(new_n3576_), .A2(new_n3564_), .B(\asqrt[53] ), .ZN(new_n3577_));
  NAND2_X1   g03385(.A1(new_n3577_), .A2(new_n904_), .ZN(new_n3578_));
  OAI21_X1   g03386(.A1(new_n3578_), .A2(new_n3566_), .B(new_n3574_), .ZN(new_n3579_));
  AOI21_X1   g03387(.A1(new_n3579_), .A2(new_n3567_), .B(new_n823_), .ZN(new_n3580_));
  NOR2_X1    g03388(.A1(new_n3311_), .A2(new_n3304_), .ZN(new_n3581_));
  NOR3_X1    g03389(.A1(new_n3419_), .A2(new_n3302_), .A3(new_n3581_), .ZN(new_n3582_));
  INV_X1     g03390(.I(new_n3582_), .ZN(new_n3583_));
  NOR3_X1    g03391(.A1(new_n3581_), .A2(new_n3302_), .A3(new_n3310_), .ZN(new_n3584_));
  AOI22_X1   g03392(.A1(new_n3583_), .A2(new_n3310_), .B1(\asqrt[42] ), .B2(new_n3584_), .ZN(new_n3585_));
  INV_X1     g03393(.I(new_n3560_), .ZN(new_n3586_));
  NAND2_X1   g03394(.A1(new_n3542_), .A2(new_n1103_), .ZN(new_n3587_));
  OAI21_X1   g03395(.A1(new_n3587_), .A2(new_n3576_), .B(new_n3586_), .ZN(new_n3588_));
  AOI21_X1   g03396(.A1(new_n3588_), .A2(new_n3577_), .B(new_n904_), .ZN(new_n3589_));
  NOR2_X1    g03397(.A1(new_n3589_), .A2(\asqrt[55] ), .ZN(new_n3590_));
  AOI21_X1   g03398(.A1(new_n3590_), .A2(new_n3579_), .B(new_n3585_), .ZN(new_n3591_));
  OAI21_X1   g03399(.A1(new_n3591_), .A2(new_n3580_), .B(\asqrt[56] ), .ZN(new_n3592_));
  NOR3_X1    g03400(.A1(new_n3313_), .A2(new_n3426_), .A3(new_n3362_), .ZN(new_n3593_));
  NOR3_X1    g03401(.A1(new_n3419_), .A2(new_n3313_), .A3(new_n3362_), .ZN(new_n3594_));
  INV_X1     g03402(.I(new_n3594_), .ZN(new_n3595_));
  AOI22_X1   g03403(.A1(new_n3595_), .A2(new_n3426_), .B1(\asqrt[42] ), .B2(new_n3593_), .ZN(new_n3596_));
  INV_X1     g03404(.I(new_n3596_), .ZN(new_n3597_));
  NOR3_X1    g03405(.A1(new_n3541_), .A2(new_n3534_), .A3(\asqrt[52] ), .ZN(new_n3598_));
  OAI21_X1   g03406(.A1(new_n3545_), .A2(new_n3598_), .B(new_n3542_), .ZN(new_n3599_));
  AOI21_X1   g03407(.A1(new_n3599_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n3600_));
  AOI21_X1   g03408(.A1(new_n3600_), .A2(new_n3588_), .B(new_n3573_), .ZN(new_n3601_));
  OAI21_X1   g03409(.A1(new_n3601_), .A2(new_n3589_), .B(\asqrt[55] ), .ZN(new_n3602_));
  NAND2_X1   g03410(.A1(new_n3602_), .A2(new_n703_), .ZN(new_n3603_));
  OAI21_X1   g03411(.A1(new_n3603_), .A2(new_n3591_), .B(new_n3597_), .ZN(new_n3604_));
  AOI21_X1   g03412(.A1(new_n3604_), .A2(new_n3592_), .B(new_n531_), .ZN(new_n3605_));
  INV_X1     g03413(.I(new_n3320_), .ZN(new_n3606_));
  NOR2_X1    g03414(.A1(new_n3335_), .A2(new_n3319_), .ZN(new_n3607_));
  NOR3_X1    g03415(.A1(new_n3419_), .A2(new_n3606_), .A3(new_n3607_), .ZN(new_n3608_));
  INV_X1     g03416(.I(new_n3608_), .ZN(new_n3609_));
  NOR3_X1    g03417(.A1(new_n3606_), .A2(new_n3326_), .A3(new_n3607_), .ZN(new_n3610_));
  AOI22_X1   g03418(.A1(new_n3609_), .A2(new_n3326_), .B1(\asqrt[42] ), .B2(new_n3610_), .ZN(new_n3611_));
  NOR3_X1    g03419(.A1(new_n3601_), .A2(\asqrt[55] ), .A3(new_n3589_), .ZN(new_n3612_));
  OAI21_X1   g03420(.A1(new_n3585_), .A2(new_n3612_), .B(new_n3602_), .ZN(new_n3613_));
  AOI21_X1   g03421(.A1(new_n3613_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n3614_));
  AOI21_X1   g03422(.A1(new_n3614_), .A2(new_n3604_), .B(new_n3611_), .ZN(new_n3615_));
  OAI21_X1   g03423(.A1(new_n3615_), .A2(new_n3605_), .B(\asqrt[58] ), .ZN(new_n3616_));
  NOR2_X1    g03424(.A1(new_n3339_), .A2(new_n3346_), .ZN(new_n3617_));
  NOR3_X1    g03425(.A1(new_n3617_), .A2(new_n3337_), .A3(new_n3345_), .ZN(new_n3618_));
  NOR3_X1    g03426(.A1(new_n3419_), .A2(new_n3337_), .A3(new_n3617_), .ZN(new_n3619_));
  INV_X1     g03427(.I(new_n3619_), .ZN(new_n3620_));
  AOI22_X1   g03428(.A1(new_n3620_), .A2(new_n3345_), .B1(\asqrt[42] ), .B2(new_n3618_), .ZN(new_n3621_));
  INV_X1     g03429(.I(new_n3621_), .ZN(new_n3622_));
  INV_X1     g03430(.I(new_n3585_), .ZN(new_n3623_));
  NAND2_X1   g03431(.A1(new_n3567_), .A2(new_n823_), .ZN(new_n3624_));
  OAI21_X1   g03432(.A1(new_n3624_), .A2(new_n3601_), .B(new_n3623_), .ZN(new_n3625_));
  AOI21_X1   g03433(.A1(new_n3625_), .A2(new_n3602_), .B(new_n703_), .ZN(new_n3626_));
  NOR2_X1    g03434(.A1(new_n3580_), .A2(\asqrt[56] ), .ZN(new_n3627_));
  AOI21_X1   g03435(.A1(new_n3627_), .A2(new_n3625_), .B(new_n3596_), .ZN(new_n3628_));
  OAI21_X1   g03436(.A1(new_n3628_), .A2(new_n3626_), .B(\asqrt[57] ), .ZN(new_n3629_));
  NAND2_X1   g03437(.A1(new_n3629_), .A2(new_n436_), .ZN(new_n3630_));
  OAI21_X1   g03438(.A1(new_n3630_), .A2(new_n3615_), .B(new_n3622_), .ZN(new_n3631_));
  AOI21_X1   g03439(.A1(new_n3631_), .A2(new_n3616_), .B(new_n327_), .ZN(new_n3632_));
  NOR3_X1    g03440(.A1(new_n3419_), .A2(new_n3348_), .A3(new_n3393_), .ZN(new_n3633_));
  INV_X1     g03441(.I(new_n3633_), .ZN(new_n3634_));
  NOR3_X1    g03442(.A1(new_n3348_), .A2(new_n3425_), .A3(new_n3393_), .ZN(new_n3635_));
  AOI22_X1   g03443(.A1(new_n3634_), .A2(new_n3425_), .B1(\asqrt[42] ), .B2(new_n3635_), .ZN(new_n3636_));
  INV_X1     g03444(.I(new_n3611_), .ZN(new_n3637_));
  NAND2_X1   g03445(.A1(new_n3592_), .A2(new_n531_), .ZN(new_n3638_));
  OAI21_X1   g03446(.A1(new_n3638_), .A2(new_n3628_), .B(new_n3637_), .ZN(new_n3639_));
  AOI21_X1   g03447(.A1(new_n3639_), .A2(new_n3629_), .B(new_n436_), .ZN(new_n3640_));
  NOR2_X1    g03448(.A1(new_n3640_), .A2(\asqrt[59] ), .ZN(new_n3641_));
  AOI21_X1   g03449(.A1(new_n3641_), .A2(new_n3631_), .B(new_n3636_), .ZN(new_n3642_));
  OAI21_X1   g03450(.A1(new_n3642_), .A2(new_n3632_), .B(\asqrt[60] ), .ZN(new_n3643_));
  INV_X1     g03451(.I(new_n3355_), .ZN(new_n3644_));
  NOR2_X1    g03452(.A1(new_n3367_), .A2(new_n3354_), .ZN(new_n3645_));
  NOR3_X1    g03453(.A1(new_n3644_), .A2(new_n3361_), .A3(new_n3645_), .ZN(new_n3646_));
  NOR3_X1    g03454(.A1(new_n3419_), .A2(new_n3644_), .A3(new_n3645_), .ZN(new_n3647_));
  INV_X1     g03455(.I(new_n3647_), .ZN(new_n3648_));
  AOI22_X1   g03456(.A1(new_n3648_), .A2(new_n3361_), .B1(\asqrt[42] ), .B2(new_n3646_), .ZN(new_n3649_));
  INV_X1     g03457(.I(new_n3649_), .ZN(new_n3650_));
  NOR2_X1    g03458(.A1(new_n3605_), .A2(\asqrt[58] ), .ZN(new_n3651_));
  AOI21_X1   g03459(.A1(new_n3651_), .A2(new_n3639_), .B(new_n3621_), .ZN(new_n3652_));
  OAI21_X1   g03460(.A1(new_n3652_), .A2(new_n3640_), .B(\asqrt[59] ), .ZN(new_n3653_));
  NAND2_X1   g03461(.A1(new_n3653_), .A2(new_n306_), .ZN(new_n3654_));
  OAI21_X1   g03462(.A1(new_n3654_), .A2(new_n3642_), .B(new_n3650_), .ZN(new_n3655_));
  AOI21_X1   g03463(.A1(new_n3655_), .A2(new_n3643_), .B(new_n218_), .ZN(new_n3656_));
  NOR2_X1    g03464(.A1(new_n3371_), .A2(new_n3377_), .ZN(new_n3657_));
  NOR3_X1    g03465(.A1(new_n3419_), .A2(new_n3369_), .A3(new_n3657_), .ZN(new_n3658_));
  INV_X1     g03466(.I(new_n3658_), .ZN(new_n3659_));
  NOR3_X1    g03467(.A1(new_n3657_), .A2(new_n3369_), .A3(new_n3376_), .ZN(new_n3660_));
  AOI22_X1   g03468(.A1(new_n3659_), .A2(new_n3376_), .B1(\asqrt[42] ), .B2(new_n3660_), .ZN(new_n3661_));
  INV_X1     g03469(.I(new_n3636_), .ZN(new_n3662_));
  NAND2_X1   g03470(.A1(new_n3616_), .A2(new_n327_), .ZN(new_n3663_));
  OAI21_X1   g03471(.A1(new_n3663_), .A2(new_n3652_), .B(new_n3662_), .ZN(new_n3664_));
  AOI21_X1   g03472(.A1(new_n3664_), .A2(new_n3653_), .B(new_n306_), .ZN(new_n3665_));
  NOR2_X1    g03473(.A1(new_n3665_), .A2(\asqrt[61] ), .ZN(new_n3666_));
  AOI21_X1   g03474(.A1(new_n3666_), .A2(new_n3655_), .B(new_n3661_), .ZN(new_n3667_));
  OAI21_X1   g03475(.A1(new_n3667_), .A2(new_n3656_), .B(\asqrt[62] ), .ZN(new_n3668_));
  NOR3_X1    g03476(.A1(new_n3379_), .A2(new_n3424_), .A3(new_n3408_), .ZN(new_n3669_));
  NOR3_X1    g03477(.A1(new_n3419_), .A2(new_n3379_), .A3(new_n3408_), .ZN(new_n3670_));
  INV_X1     g03478(.I(new_n3670_), .ZN(new_n3671_));
  AOI22_X1   g03479(.A1(new_n3671_), .A2(new_n3424_), .B1(\asqrt[42] ), .B2(new_n3669_), .ZN(new_n3672_));
  INV_X1     g03480(.I(new_n3672_), .ZN(new_n3673_));
  NOR3_X1    g03481(.A1(new_n3615_), .A2(\asqrt[58] ), .A3(new_n3605_), .ZN(new_n3674_));
  OAI21_X1   g03482(.A1(new_n3621_), .A2(new_n3674_), .B(new_n3616_), .ZN(new_n3675_));
  AOI21_X1   g03483(.A1(new_n3675_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n3676_));
  AOI21_X1   g03484(.A1(new_n3676_), .A2(new_n3664_), .B(new_n3649_), .ZN(new_n3677_));
  OAI21_X1   g03485(.A1(new_n3677_), .A2(new_n3665_), .B(\asqrt[61] ), .ZN(new_n3678_));
  NAND2_X1   g03486(.A1(new_n3678_), .A2(new_n207_), .ZN(new_n3679_));
  OAI21_X1   g03487(.A1(new_n3679_), .A2(new_n3667_), .B(new_n3673_), .ZN(new_n3680_));
  INV_X1     g03488(.I(new_n3470_), .ZN(new_n3681_));
  NAND4_X1   g03489(.A1(\asqrt[42] ), .A2(new_n3386_), .A3(new_n3391_), .A4(new_n3449_), .ZN(new_n3682_));
  NAND2_X1   g03490(.A1(new_n3386_), .A2(new_n3449_), .ZN(new_n3683_));
  OAI21_X1   g03491(.A1(new_n3419_), .A2(new_n3683_), .B(new_n3392_), .ZN(new_n3684_));
  NAND2_X1   g03492(.A1(new_n3684_), .A2(new_n3682_), .ZN(new_n3685_));
  NOR2_X1    g03493(.A1(new_n3450_), .A2(new_n3465_), .ZN(new_n3686_));
  NAND2_X1   g03494(.A1(\asqrt[42] ), .A2(new_n3686_), .ZN(new_n3687_));
  NAND3_X1   g03495(.A1(new_n3685_), .A2(new_n3681_), .A3(new_n3687_), .ZN(new_n3688_));
  AOI21_X1   g03496(.A1(new_n3680_), .A2(new_n3668_), .B(new_n3688_), .ZN(new_n3689_));
  NOR3_X1    g03497(.A1(new_n3677_), .A2(\asqrt[61] ), .A3(new_n3665_), .ZN(new_n3690_));
  OAI21_X1   g03498(.A1(new_n3661_), .A2(new_n3690_), .B(new_n3678_), .ZN(new_n3691_));
  AOI21_X1   g03499(.A1(new_n3691_), .A2(\asqrt[62] ), .B(new_n3685_), .ZN(new_n3692_));
  OAI21_X1   g03500(.A1(new_n3419_), .A2(new_n3465_), .B(new_n3450_), .ZN(new_n3693_));
  NOR2_X1    g03501(.A1(new_n3686_), .A2(new_n193_), .ZN(new_n3694_));
  NAND2_X1   g03502(.A1(new_n3693_), .A2(new_n3694_), .ZN(new_n3695_));
  INV_X1     g03503(.I(new_n3695_), .ZN(new_n3696_));
  AND3_X2    g03504(.A1(new_n3402_), .A2(new_n3400_), .A3(new_n3415_), .Z(new_n3697_));
  NAND4_X1   g03505(.A1(new_n3681_), .A2(new_n3451_), .A3(new_n3412_), .A4(new_n3697_), .ZN(new_n3698_));
  INV_X1     g03506(.I(new_n3698_), .ZN(new_n3699_));
  NOR2_X1    g03507(.A1(new_n3696_), .A2(new_n3699_), .ZN(new_n3700_));
  INV_X1     g03508(.I(new_n3700_), .ZN(new_n3701_));
  AOI21_X1   g03509(.A1(new_n3692_), .A2(new_n3680_), .B(new_n3701_), .ZN(new_n3702_));
  OAI21_X1   g03510(.A1(\asqrt[63] ), .A2(new_n3689_), .B(new_n3702_), .ZN(\asqrt[41] ));
  NOR2_X1    g03511(.A1(\a[80] ), .A2(\a[81] ), .ZN(new_n3704_));
  INV_X1     g03512(.I(new_n3704_), .ZN(new_n3705_));
  NOR2_X1    g03513(.A1(new_n3705_), .A2(\a[82] ), .ZN(new_n3706_));
  INV_X1     g03514(.I(new_n3706_), .ZN(new_n3707_));
  NAND2_X1   g03515(.A1(new_n3680_), .A2(new_n3668_), .ZN(new_n3708_));
  INV_X1     g03516(.I(new_n3688_), .ZN(new_n3709_));
  AOI21_X1   g03517(.A1(new_n3708_), .A2(new_n3709_), .B(\asqrt[63] ), .ZN(new_n3710_));
  INV_X1     g03518(.I(new_n3680_), .ZN(new_n3711_));
  INV_X1     g03519(.I(new_n3685_), .ZN(new_n3712_));
  NAND2_X1   g03520(.A1(new_n3668_), .A2(new_n3712_), .ZN(new_n3713_));
  OAI21_X1   g03521(.A1(new_n3711_), .A2(new_n3713_), .B(new_n3700_), .ZN(new_n3714_));
  OAI21_X1   g03522(.A1(new_n3710_), .A2(new_n3714_), .B(\a[82] ), .ZN(new_n3715_));
  AOI21_X1   g03523(.A1(new_n3715_), .A2(new_n3707_), .B(new_n3419_), .ZN(new_n3716_));
  INV_X1     g03524(.I(\a[82] ), .ZN(new_n3717_));
  INV_X1     g03525(.I(new_n3661_), .ZN(new_n3718_));
  NAND2_X1   g03526(.A1(new_n3643_), .A2(new_n218_), .ZN(new_n3719_));
  OAI21_X1   g03527(.A1(new_n3719_), .A2(new_n3677_), .B(new_n3718_), .ZN(new_n3720_));
  NAND3_X1   g03528(.A1(new_n3720_), .A2(new_n207_), .A3(new_n3678_), .ZN(new_n3721_));
  AOI22_X1   g03529(.A1(new_n3721_), .A2(new_n3673_), .B1(new_n3691_), .B2(\asqrt[62] ), .ZN(new_n3722_));
  OAI21_X1   g03530(.A1(new_n3722_), .A2(new_n3688_), .B(new_n193_), .ZN(new_n3723_));
  AOI21_X1   g03531(.A1(new_n3723_), .A2(new_n3702_), .B(new_n3717_), .ZN(new_n3724_));
  NAND4_X1   g03532(.A1(new_n3681_), .A2(new_n3412_), .A3(new_n3415_), .A4(new_n3707_), .ZN(new_n3725_));
  NOR2_X1    g03533(.A1(new_n3725_), .A2(new_n3463_), .ZN(new_n3726_));
  INV_X1     g03534(.I(new_n3726_), .ZN(new_n3727_));
  NOR2_X1    g03535(.A1(new_n3724_), .A2(new_n3727_), .ZN(new_n3728_));
  AOI21_X1   g03536(.A1(new_n3723_), .A2(new_n3702_), .B(new_n3421_), .ZN(new_n3729_));
  INV_X1     g03537(.I(\a[83] ), .ZN(new_n3730_));
  AOI21_X1   g03538(.A1(\asqrt[41] ), .A2(new_n3717_), .B(new_n3730_), .ZN(new_n3731_));
  NOR3_X1    g03539(.A1(new_n3728_), .A2(new_n3731_), .A3(new_n3729_), .ZN(new_n3732_));
  OAI21_X1   g03540(.A1(new_n3732_), .A2(new_n3716_), .B(\asqrt[43] ), .ZN(new_n3733_));
  OAI21_X1   g03541(.A1(new_n3710_), .A2(new_n3714_), .B(new_n3420_), .ZN(new_n3734_));
  NOR2_X1    g03542(.A1(new_n3711_), .A2(new_n3713_), .ZN(new_n3735_));
  INV_X1     g03543(.I(new_n3735_), .ZN(new_n3736_));
  NOR2_X1    g03544(.A1(new_n3699_), .A2(new_n3419_), .ZN(new_n3737_));
  NAND4_X1   g03545(.A1(new_n3736_), .A2(new_n3723_), .A3(new_n3695_), .A4(new_n3737_), .ZN(new_n3738_));
  AOI21_X1   g03546(.A1(new_n3738_), .A2(new_n3734_), .B(new_n3423_), .ZN(new_n3739_));
  INV_X1     g03547(.I(new_n3737_), .ZN(new_n3740_));
  NOR4_X1    g03548(.A1(new_n3710_), .A2(new_n3735_), .A3(new_n3696_), .A4(new_n3740_), .ZN(new_n3741_));
  NOR3_X1    g03549(.A1(new_n3741_), .A2(new_n3729_), .A3(\a[84] ), .ZN(new_n3742_));
  AOI21_X1   g03550(.A1(\asqrt[41] ), .A2(\a[82] ), .B(new_n3706_), .ZN(new_n3743_));
  OAI21_X1   g03551(.A1(new_n3743_), .A2(new_n3419_), .B(new_n3218_), .ZN(new_n3744_));
  OAI22_X1   g03552(.A1(new_n3732_), .A2(new_n3744_), .B1(new_n3739_), .B2(new_n3742_), .ZN(new_n3745_));
  AOI21_X1   g03553(.A1(new_n3745_), .A2(new_n3733_), .B(new_n2954_), .ZN(new_n3746_));
  INV_X1     g03554(.I(new_n3485_), .ZN(new_n3747_));
  NOR3_X1    g03555(.A1(new_n3454_), .A2(new_n3747_), .A3(new_n3457_), .ZN(new_n3748_));
  NOR2_X1    g03556(.A1(new_n3454_), .A2(new_n3457_), .ZN(new_n3749_));
  NAND2_X1   g03557(.A1(\asqrt[41] ), .A2(new_n3749_), .ZN(new_n3750_));
  AOI22_X1   g03558(.A1(new_n3750_), .A2(new_n3747_), .B1(\asqrt[41] ), .B2(new_n3748_), .ZN(new_n3751_));
  OAI21_X1   g03559(.A1(new_n3724_), .A2(new_n3706_), .B(\asqrt[42] ), .ZN(new_n3752_));
  AOI21_X1   g03560(.A1(new_n3723_), .A2(new_n3702_), .B(\a[82] ), .ZN(new_n3753_));
  OAI21_X1   g03561(.A1(new_n3730_), .A2(new_n3753_), .B(new_n3734_), .ZN(new_n3754_));
  OAI21_X1   g03562(.A1(new_n3754_), .A2(new_n3728_), .B(new_n3752_), .ZN(new_n3755_));
  AOI21_X1   g03563(.A1(new_n3755_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n3756_));
  AOI21_X1   g03564(.A1(new_n3756_), .A2(new_n3745_), .B(new_n3751_), .ZN(new_n3757_));
  OAI21_X1   g03565(.A1(new_n3757_), .A2(new_n3746_), .B(\asqrt[45] ), .ZN(new_n3758_));
  INV_X1     g03566(.I(new_n3758_), .ZN(new_n3759_));
  NOR2_X1    g03567(.A1(new_n3475_), .A2(new_n3476_), .ZN(new_n3760_));
  NOR2_X1    g03568(.A1(new_n3461_), .A2(new_n3478_), .ZN(new_n3761_));
  INV_X1     g03569(.I(new_n3761_), .ZN(new_n3762_));
  NAND4_X1   g03570(.A1(\asqrt[41] ), .A2(new_n3462_), .A3(new_n3760_), .A4(new_n3762_), .ZN(new_n3763_));
  AND3_X2    g03571(.A1(\asqrt[41] ), .A2(new_n3462_), .A3(new_n3762_), .Z(new_n3764_));
  OAI21_X1   g03572(.A1(new_n3764_), .A2(new_n3760_), .B(new_n3763_), .ZN(new_n3765_));
  INV_X1     g03573(.I(new_n3765_), .ZN(new_n3766_));
  NOR3_X1    g03574(.A1(new_n3757_), .A2(new_n3746_), .A3(\asqrt[45] ), .ZN(new_n3767_));
  NOR2_X1    g03575(.A1(new_n3767_), .A2(new_n3766_), .ZN(new_n3768_));
  OAI21_X1   g03576(.A1(new_n3768_), .A2(new_n3759_), .B(\asqrt[46] ), .ZN(new_n3769_));
  INV_X1     g03577(.I(new_n3483_), .ZN(new_n3770_));
  INV_X1     g03578(.I(new_n3480_), .ZN(new_n3771_));
  NAND2_X1   g03579(.A1(new_n3487_), .A2(new_n3479_), .ZN(new_n3772_));
  NAND3_X1   g03580(.A1(\asqrt[41] ), .A2(new_n3771_), .A3(new_n3772_), .ZN(new_n3773_));
  AND3_X2    g03581(.A1(new_n3771_), .A2(new_n3483_), .A3(new_n3772_), .Z(new_n3774_));
  AOI22_X1   g03582(.A1(new_n3773_), .A2(new_n3770_), .B1(\asqrt[41] ), .B2(new_n3774_), .ZN(new_n3775_));
  INV_X1     g03583(.I(new_n3775_), .ZN(new_n3776_));
  NAND2_X1   g03584(.A1(new_n3758_), .A2(new_n2465_), .ZN(new_n3777_));
  OAI21_X1   g03585(.A1(new_n3768_), .A2(new_n3777_), .B(new_n3776_), .ZN(new_n3778_));
  AOI21_X1   g03586(.A1(new_n3778_), .A2(new_n3769_), .B(new_n2229_), .ZN(new_n3779_));
  INV_X1     g03587(.I(new_n3497_), .ZN(new_n3780_));
  NOR3_X1    g03588(.A1(new_n3490_), .A2(new_n3780_), .A3(new_n3498_), .ZN(new_n3781_));
  INV_X1     g03589(.I(\asqrt[41] ), .ZN(new_n3782_));
  NOR3_X1    g03590(.A1(new_n3782_), .A2(new_n3490_), .A3(new_n3498_), .ZN(new_n3783_));
  INV_X1     g03591(.I(new_n3783_), .ZN(new_n3784_));
  AOI22_X1   g03592(.A1(new_n3784_), .A2(new_n3780_), .B1(\asqrt[41] ), .B2(new_n3781_), .ZN(new_n3785_));
  OAI21_X1   g03593(.A1(new_n3766_), .A2(new_n3767_), .B(new_n3758_), .ZN(new_n3786_));
  AOI21_X1   g03594(.A1(new_n3786_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n3787_));
  AOI21_X1   g03595(.A1(new_n3787_), .A2(new_n3778_), .B(new_n3785_), .ZN(new_n3788_));
  OAI21_X1   g03596(.A1(new_n3788_), .A2(new_n3779_), .B(\asqrt[48] ), .ZN(new_n3789_));
  INV_X1     g03597(.I(new_n3789_), .ZN(new_n3790_));
  INV_X1     g03598(.I(new_n3499_), .ZN(new_n3791_));
  INV_X1     g03599(.I(new_n3507_), .ZN(new_n3792_));
  NAND2_X1   g03600(.A1(new_n3791_), .A2(new_n3792_), .ZN(new_n3793_));
  NAND3_X1   g03601(.A1(\asqrt[41] ), .A2(new_n3500_), .A3(new_n3793_), .ZN(new_n3794_));
  AND3_X2    g03602(.A1(new_n3793_), .A2(new_n3500_), .A3(new_n3505_), .Z(new_n3795_));
  AOI22_X1   g03603(.A1(new_n3794_), .A2(new_n3506_), .B1(\asqrt[41] ), .B2(new_n3795_), .ZN(new_n3796_));
  NOR3_X1    g03604(.A1(new_n3788_), .A2(new_n3779_), .A3(\asqrt[48] ), .ZN(new_n3797_));
  NOR2_X1    g03605(.A1(new_n3797_), .A2(new_n3796_), .ZN(new_n3798_));
  OAI21_X1   g03606(.A1(new_n3798_), .A2(new_n3790_), .B(\asqrt[49] ), .ZN(new_n3799_));
  INV_X1     g03607(.I(new_n3513_), .ZN(new_n3800_));
  INV_X1     g03608(.I(new_n3508_), .ZN(new_n3801_));
  INV_X1     g03609(.I(new_n3515_), .ZN(new_n3802_));
  NOR2_X1    g03610(.A1(new_n3802_), .A2(new_n3801_), .ZN(new_n3803_));
  NOR3_X1    g03611(.A1(new_n3803_), .A2(new_n3509_), .A3(new_n3800_), .ZN(new_n3804_));
  NOR3_X1    g03612(.A1(new_n3782_), .A2(new_n3509_), .A3(new_n3803_), .ZN(new_n3805_));
  INV_X1     g03613(.I(new_n3805_), .ZN(new_n3806_));
  AOI22_X1   g03614(.A1(new_n3806_), .A2(new_n3800_), .B1(\asqrt[41] ), .B2(new_n3804_), .ZN(new_n3807_));
  INV_X1     g03615(.I(new_n3807_), .ZN(new_n3808_));
  NAND2_X1   g03616(.A1(new_n3789_), .A2(new_n1806_), .ZN(new_n3809_));
  OAI21_X1   g03617(.A1(new_n3798_), .A2(new_n3809_), .B(new_n3808_), .ZN(new_n3810_));
  AOI21_X1   g03618(.A1(new_n3810_), .A2(new_n3799_), .B(new_n1612_), .ZN(new_n3811_));
  NOR3_X1    g03619(.A1(new_n3782_), .A2(new_n3518_), .A3(new_n3524_), .ZN(new_n3812_));
  INV_X1     g03620(.I(new_n3812_), .ZN(new_n3813_));
  NOR3_X1    g03621(.A1(new_n3518_), .A2(new_n3547_), .A3(new_n3524_), .ZN(new_n3814_));
  AOI22_X1   g03622(.A1(new_n3813_), .A2(new_n3547_), .B1(\asqrt[41] ), .B2(new_n3814_), .ZN(new_n3815_));
  OAI21_X1   g03623(.A1(new_n3796_), .A2(new_n3797_), .B(new_n3789_), .ZN(new_n3816_));
  AOI21_X1   g03624(.A1(new_n3816_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n3817_));
  AOI21_X1   g03625(.A1(new_n3817_), .A2(new_n3810_), .B(new_n3815_), .ZN(new_n3818_));
  OAI21_X1   g03626(.A1(new_n3818_), .A2(new_n3811_), .B(\asqrt[51] ), .ZN(new_n3819_));
  INV_X1     g03627(.I(new_n3819_), .ZN(new_n3820_));
  NOR2_X1    g03628(.A1(new_n3525_), .A2(new_n3532_), .ZN(new_n3821_));
  NOR3_X1    g03629(.A1(new_n3550_), .A2(new_n3821_), .A3(new_n3531_), .ZN(new_n3822_));
  NOR3_X1    g03630(.A1(new_n3782_), .A2(new_n3550_), .A3(new_n3821_), .ZN(new_n3823_));
  INV_X1     g03631(.I(new_n3823_), .ZN(new_n3824_));
  AOI22_X1   g03632(.A1(new_n3824_), .A2(new_n3531_), .B1(\asqrt[41] ), .B2(new_n3822_), .ZN(new_n3825_));
  NOR3_X1    g03633(.A1(new_n3818_), .A2(new_n3811_), .A3(\asqrt[51] ), .ZN(new_n3826_));
  NOR2_X1    g03634(.A1(new_n3826_), .A2(new_n3825_), .ZN(new_n3827_));
  OAI21_X1   g03635(.A1(new_n3827_), .A2(new_n3820_), .B(\asqrt[52] ), .ZN(new_n3828_));
  NOR2_X1    g03636(.A1(new_n3562_), .A2(new_n3552_), .ZN(new_n3829_));
  NOR3_X1    g03637(.A1(new_n3782_), .A2(new_n3534_), .A3(new_n3829_), .ZN(new_n3830_));
  INV_X1     g03638(.I(new_n3830_), .ZN(new_n3831_));
  NOR3_X1    g03639(.A1(new_n3829_), .A2(new_n3534_), .A3(new_n3561_), .ZN(new_n3832_));
  AOI22_X1   g03640(.A1(new_n3831_), .A2(new_n3561_), .B1(\asqrt[41] ), .B2(new_n3832_), .ZN(new_n3833_));
  INV_X1     g03641(.I(new_n3833_), .ZN(new_n3834_));
  NAND2_X1   g03642(.A1(new_n3819_), .A2(new_n1256_), .ZN(new_n3835_));
  OAI21_X1   g03643(.A1(new_n3827_), .A2(new_n3835_), .B(new_n3834_), .ZN(new_n3836_));
  AOI21_X1   g03644(.A1(new_n3836_), .A2(new_n3828_), .B(new_n1103_), .ZN(new_n3837_));
  NOR3_X1    g03645(.A1(new_n3564_), .A2(new_n3598_), .A3(new_n3546_), .ZN(new_n3838_));
  NOR3_X1    g03646(.A1(new_n3782_), .A2(new_n3564_), .A3(new_n3598_), .ZN(new_n3839_));
  INV_X1     g03647(.I(new_n3839_), .ZN(new_n3840_));
  AOI22_X1   g03648(.A1(new_n3840_), .A2(new_n3546_), .B1(\asqrt[41] ), .B2(new_n3838_), .ZN(new_n3841_));
  OAI21_X1   g03649(.A1(new_n3825_), .A2(new_n3826_), .B(new_n3819_), .ZN(new_n3842_));
  AOI21_X1   g03650(.A1(new_n3842_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n3843_));
  AOI21_X1   g03651(.A1(new_n3843_), .A2(new_n3836_), .B(new_n3841_), .ZN(new_n3844_));
  OAI21_X1   g03652(.A1(new_n3844_), .A2(new_n3837_), .B(\asqrt[54] ), .ZN(new_n3845_));
  INV_X1     g03653(.I(new_n3845_), .ZN(new_n3846_));
  NOR2_X1    g03654(.A1(new_n3587_), .A2(new_n3576_), .ZN(new_n3847_));
  NOR3_X1    g03655(.A1(new_n3782_), .A2(new_n3556_), .A3(new_n3847_), .ZN(new_n3848_));
  INV_X1     g03656(.I(new_n3848_), .ZN(new_n3849_));
  NOR3_X1    g03657(.A1(new_n3556_), .A2(new_n3847_), .A3(new_n3586_), .ZN(new_n3850_));
  AOI22_X1   g03658(.A1(new_n3849_), .A2(new_n3586_), .B1(\asqrt[41] ), .B2(new_n3850_), .ZN(new_n3851_));
  NOR3_X1    g03659(.A1(new_n3844_), .A2(new_n3837_), .A3(\asqrt[54] ), .ZN(new_n3852_));
  NOR2_X1    g03660(.A1(new_n3852_), .A2(new_n3851_), .ZN(new_n3853_));
  OAI21_X1   g03661(.A1(new_n3853_), .A2(new_n3846_), .B(\asqrt[55] ), .ZN(new_n3854_));
  NOR2_X1    g03662(.A1(new_n3578_), .A2(new_n3566_), .ZN(new_n3855_));
  NOR3_X1    g03663(.A1(new_n3855_), .A2(new_n3589_), .A3(new_n3574_), .ZN(new_n3856_));
  NOR3_X1    g03664(.A1(new_n3782_), .A2(new_n3589_), .A3(new_n3855_), .ZN(new_n3857_));
  INV_X1     g03665(.I(new_n3857_), .ZN(new_n3858_));
  AOI22_X1   g03666(.A1(new_n3858_), .A2(new_n3574_), .B1(\asqrt[41] ), .B2(new_n3856_), .ZN(new_n3859_));
  INV_X1     g03667(.I(new_n3859_), .ZN(new_n3860_));
  NAND2_X1   g03668(.A1(new_n3845_), .A2(new_n823_), .ZN(new_n3861_));
  OAI21_X1   g03669(.A1(new_n3853_), .A2(new_n3861_), .B(new_n3860_), .ZN(new_n3862_));
  AOI21_X1   g03670(.A1(new_n3862_), .A2(new_n3854_), .B(new_n703_), .ZN(new_n3863_));
  NOR3_X1    g03671(.A1(new_n3782_), .A2(new_n3580_), .A3(new_n3612_), .ZN(new_n3864_));
  INV_X1     g03672(.I(new_n3864_), .ZN(new_n3865_));
  NOR3_X1    g03673(.A1(new_n3580_), .A2(new_n3612_), .A3(new_n3623_), .ZN(new_n3866_));
  AOI22_X1   g03674(.A1(new_n3865_), .A2(new_n3623_), .B1(\asqrt[41] ), .B2(new_n3866_), .ZN(new_n3867_));
  OAI21_X1   g03675(.A1(new_n3851_), .A2(new_n3852_), .B(new_n3845_), .ZN(new_n3868_));
  AOI21_X1   g03676(.A1(new_n3868_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n3869_));
  AOI21_X1   g03677(.A1(new_n3869_), .A2(new_n3862_), .B(new_n3867_), .ZN(new_n3870_));
  OAI21_X1   g03678(.A1(new_n3870_), .A2(new_n3863_), .B(\asqrt[57] ), .ZN(new_n3871_));
  NOR2_X1    g03679(.A1(new_n3603_), .A2(new_n3591_), .ZN(new_n3872_));
  NOR3_X1    g03680(.A1(new_n3626_), .A2(new_n3872_), .A3(new_n3597_), .ZN(new_n3873_));
  NOR3_X1    g03681(.A1(new_n3782_), .A2(new_n3626_), .A3(new_n3872_), .ZN(new_n3874_));
  INV_X1     g03682(.I(new_n3874_), .ZN(new_n3875_));
  AOI22_X1   g03683(.A1(new_n3875_), .A2(new_n3597_), .B1(\asqrt[41] ), .B2(new_n3873_), .ZN(new_n3876_));
  INV_X1     g03684(.I(new_n3876_), .ZN(new_n3877_));
  INV_X1     g03685(.I(new_n3851_), .ZN(new_n3878_));
  INV_X1     g03686(.I(new_n3825_), .ZN(new_n3879_));
  INV_X1     g03687(.I(new_n3796_), .ZN(new_n3880_));
  NAND2_X1   g03688(.A1(new_n3715_), .A2(new_n3726_), .ZN(new_n3881_));
  OAI21_X1   g03689(.A1(new_n3710_), .A2(new_n3714_), .B(new_n3717_), .ZN(new_n3882_));
  NAND2_X1   g03690(.A1(new_n3882_), .A2(\a[83] ), .ZN(new_n3883_));
  NAND3_X1   g03691(.A1(new_n3881_), .A2(new_n3883_), .A3(new_n3734_), .ZN(new_n3884_));
  AOI21_X1   g03692(.A1(new_n3884_), .A2(new_n3752_), .B(new_n3218_), .ZN(new_n3885_));
  OAI21_X1   g03693(.A1(new_n3741_), .A2(new_n3729_), .B(\a[84] ), .ZN(new_n3886_));
  NAND3_X1   g03694(.A1(new_n3738_), .A2(new_n3734_), .A3(new_n3423_), .ZN(new_n3887_));
  NAND2_X1   g03695(.A1(new_n3715_), .A2(new_n3707_), .ZN(new_n3888_));
  AOI21_X1   g03696(.A1(new_n3888_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n3889_));
  AOI22_X1   g03697(.A1(new_n3884_), .A2(new_n3889_), .B1(new_n3886_), .B2(new_n3887_), .ZN(new_n3890_));
  OAI21_X1   g03698(.A1(new_n3890_), .A2(new_n3885_), .B(\asqrt[44] ), .ZN(new_n3891_));
  NAND2_X1   g03699(.A1(new_n3891_), .A2(new_n2641_), .ZN(new_n3892_));
  OAI21_X1   g03700(.A1(new_n3892_), .A2(new_n3757_), .B(new_n3765_), .ZN(new_n3893_));
  AOI21_X1   g03701(.A1(new_n3893_), .A2(new_n3758_), .B(new_n2465_), .ZN(new_n3894_));
  INV_X1     g03702(.I(new_n3751_), .ZN(new_n3895_));
  AOI21_X1   g03703(.A1(\a[83] ), .A2(new_n3882_), .B(new_n3729_), .ZN(new_n3896_));
  AOI21_X1   g03704(.A1(new_n3896_), .A2(new_n3881_), .B(new_n3716_), .ZN(new_n3897_));
  OAI21_X1   g03705(.A1(new_n3897_), .A2(new_n3218_), .B(new_n2954_), .ZN(new_n3898_));
  OAI21_X1   g03706(.A1(new_n3898_), .A2(new_n3890_), .B(new_n3895_), .ZN(new_n3899_));
  NAND2_X1   g03707(.A1(new_n3899_), .A2(new_n3891_), .ZN(new_n3900_));
  AOI21_X1   g03708(.A1(new_n3900_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n3901_));
  AOI21_X1   g03709(.A1(new_n3901_), .A2(new_n3893_), .B(new_n3775_), .ZN(new_n3902_));
  OAI21_X1   g03710(.A1(new_n3902_), .A2(new_n3894_), .B(\asqrt[47] ), .ZN(new_n3903_));
  NAND2_X1   g03711(.A1(new_n3903_), .A2(new_n1956_), .ZN(new_n3904_));
  OAI21_X1   g03712(.A1(new_n3904_), .A2(new_n3788_), .B(new_n3880_), .ZN(new_n3905_));
  NAND3_X1   g03713(.A1(new_n3905_), .A2(new_n1806_), .A3(new_n3789_), .ZN(new_n3906_));
  AOI22_X1   g03714(.A1(new_n3906_), .A2(new_n3808_), .B1(new_n3816_), .B2(\asqrt[49] ), .ZN(new_n3907_));
  OAI21_X1   g03715(.A1(new_n3907_), .A2(new_n1612_), .B(new_n1376_), .ZN(new_n3908_));
  OAI21_X1   g03716(.A1(new_n3908_), .A2(new_n3818_), .B(new_n3879_), .ZN(new_n3909_));
  AOI21_X1   g03717(.A1(new_n3909_), .A2(new_n3819_), .B(new_n1256_), .ZN(new_n3910_));
  AOI21_X1   g03718(.A1(new_n3905_), .A2(new_n3789_), .B(new_n1806_), .ZN(new_n3911_));
  NOR3_X1    g03719(.A1(new_n3902_), .A2(new_n3894_), .A3(\asqrt[47] ), .ZN(new_n3912_));
  OAI21_X1   g03720(.A1(new_n3785_), .A2(new_n3912_), .B(new_n3903_), .ZN(new_n3913_));
  AOI21_X1   g03721(.A1(new_n3913_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n3914_));
  AOI21_X1   g03722(.A1(new_n3914_), .A2(new_n3905_), .B(new_n3807_), .ZN(new_n3915_));
  NOR3_X1    g03723(.A1(new_n3915_), .A2(\asqrt[50] ), .A3(new_n3911_), .ZN(new_n3916_));
  OAI22_X1   g03724(.A1(new_n3916_), .A2(new_n3815_), .B1(new_n3907_), .B2(new_n1612_), .ZN(new_n3917_));
  AOI21_X1   g03725(.A1(new_n3917_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n3918_));
  AOI21_X1   g03726(.A1(new_n3918_), .A2(new_n3909_), .B(new_n3833_), .ZN(new_n3919_));
  OAI21_X1   g03727(.A1(new_n3919_), .A2(new_n3910_), .B(\asqrt[53] ), .ZN(new_n3920_));
  NAND2_X1   g03728(.A1(new_n3920_), .A2(new_n904_), .ZN(new_n3921_));
  OAI21_X1   g03729(.A1(new_n3921_), .A2(new_n3844_), .B(new_n3878_), .ZN(new_n3922_));
  AOI21_X1   g03730(.A1(new_n3922_), .A2(new_n3845_), .B(new_n823_), .ZN(new_n3923_));
  NOR3_X1    g03731(.A1(new_n3919_), .A2(\asqrt[53] ), .A3(new_n3910_), .ZN(new_n3924_));
  OAI21_X1   g03732(.A1(new_n3841_), .A2(new_n3924_), .B(new_n3920_), .ZN(new_n3925_));
  AOI21_X1   g03733(.A1(new_n3925_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n3926_));
  AOI21_X1   g03734(.A1(new_n3926_), .A2(new_n3922_), .B(new_n3859_), .ZN(new_n3927_));
  OAI21_X1   g03735(.A1(new_n3927_), .A2(new_n3923_), .B(\asqrt[56] ), .ZN(new_n3928_));
  NAND2_X1   g03736(.A1(new_n3928_), .A2(new_n531_), .ZN(new_n3929_));
  OAI21_X1   g03737(.A1(new_n3929_), .A2(new_n3870_), .B(new_n3877_), .ZN(new_n3930_));
  AOI21_X1   g03738(.A1(new_n3930_), .A2(new_n3871_), .B(new_n436_), .ZN(new_n3931_));
  NOR2_X1    g03739(.A1(new_n3638_), .A2(new_n3628_), .ZN(new_n3932_));
  NOR3_X1    g03740(.A1(new_n3782_), .A2(new_n3605_), .A3(new_n3932_), .ZN(new_n3933_));
  INV_X1     g03741(.I(new_n3933_), .ZN(new_n3934_));
  NOR3_X1    g03742(.A1(new_n3932_), .A2(new_n3605_), .A3(new_n3637_), .ZN(new_n3935_));
  AOI22_X1   g03743(.A1(new_n3934_), .A2(new_n3637_), .B1(\asqrt[41] ), .B2(new_n3935_), .ZN(new_n3936_));
  NOR3_X1    g03744(.A1(new_n3927_), .A2(\asqrt[56] ), .A3(new_n3923_), .ZN(new_n3937_));
  OAI21_X1   g03745(.A1(new_n3867_), .A2(new_n3937_), .B(new_n3928_), .ZN(new_n3938_));
  AOI21_X1   g03746(.A1(new_n3938_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n3939_));
  AOI21_X1   g03747(.A1(new_n3939_), .A2(new_n3930_), .B(new_n3936_), .ZN(new_n3940_));
  OAI21_X1   g03748(.A1(new_n3940_), .A2(new_n3931_), .B(\asqrt[59] ), .ZN(new_n3941_));
  NOR3_X1    g03749(.A1(new_n3640_), .A2(new_n3674_), .A3(new_n3622_), .ZN(new_n3942_));
  NOR3_X1    g03750(.A1(new_n3782_), .A2(new_n3640_), .A3(new_n3674_), .ZN(new_n3943_));
  INV_X1     g03751(.I(new_n3943_), .ZN(new_n3944_));
  AOI22_X1   g03752(.A1(new_n3944_), .A2(new_n3622_), .B1(\asqrt[41] ), .B2(new_n3942_), .ZN(new_n3945_));
  INV_X1     g03753(.I(new_n3945_), .ZN(new_n3946_));
  INV_X1     g03754(.I(new_n3871_), .ZN(new_n3947_));
  NOR3_X1    g03755(.A1(new_n3870_), .A2(new_n3863_), .A3(\asqrt[57] ), .ZN(new_n3948_));
  NOR2_X1    g03756(.A1(new_n3948_), .A2(new_n3876_), .ZN(new_n3949_));
  OAI21_X1   g03757(.A1(new_n3949_), .A2(new_n3947_), .B(\asqrt[58] ), .ZN(new_n3950_));
  NAND2_X1   g03758(.A1(new_n3950_), .A2(new_n327_), .ZN(new_n3951_));
  OAI21_X1   g03759(.A1(new_n3951_), .A2(new_n3940_), .B(new_n3946_), .ZN(new_n3952_));
  AOI21_X1   g03760(.A1(new_n3952_), .A2(new_n3941_), .B(new_n306_), .ZN(new_n3953_));
  NOR2_X1    g03761(.A1(new_n3663_), .A2(new_n3652_), .ZN(new_n3954_));
  NOR3_X1    g03762(.A1(new_n3782_), .A2(new_n3632_), .A3(new_n3954_), .ZN(new_n3955_));
  INV_X1     g03763(.I(new_n3955_), .ZN(new_n3956_));
  NOR3_X1    g03764(.A1(new_n3632_), .A2(new_n3954_), .A3(new_n3662_), .ZN(new_n3957_));
  AOI22_X1   g03765(.A1(new_n3956_), .A2(new_n3662_), .B1(\asqrt[41] ), .B2(new_n3957_), .ZN(new_n3958_));
  INV_X1     g03766(.I(new_n3936_), .ZN(new_n3959_));
  NAND2_X1   g03767(.A1(new_n3871_), .A2(new_n436_), .ZN(new_n3960_));
  OAI21_X1   g03768(.A1(new_n3949_), .A2(new_n3960_), .B(new_n3959_), .ZN(new_n3961_));
  AOI21_X1   g03769(.A1(new_n3961_), .A2(new_n3950_), .B(new_n327_), .ZN(new_n3962_));
  NOR2_X1    g03770(.A1(new_n3962_), .A2(\asqrt[60] ), .ZN(new_n3963_));
  AOI21_X1   g03771(.A1(new_n3963_), .A2(new_n3952_), .B(new_n3958_), .ZN(new_n3964_));
  OAI21_X1   g03772(.A1(new_n3964_), .A2(new_n3953_), .B(\asqrt[61] ), .ZN(new_n3965_));
  NOR2_X1    g03773(.A1(new_n3654_), .A2(new_n3642_), .ZN(new_n3966_));
  NOR3_X1    g03774(.A1(new_n3966_), .A2(new_n3665_), .A3(new_n3650_), .ZN(new_n3967_));
  NOR3_X1    g03775(.A1(new_n3782_), .A2(new_n3665_), .A3(new_n3966_), .ZN(new_n3968_));
  INV_X1     g03776(.I(new_n3968_), .ZN(new_n3969_));
  AOI22_X1   g03777(.A1(new_n3969_), .A2(new_n3650_), .B1(\asqrt[41] ), .B2(new_n3967_), .ZN(new_n3970_));
  INV_X1     g03778(.I(new_n3970_), .ZN(new_n3971_));
  OAI21_X1   g03779(.A1(new_n3876_), .A2(new_n3948_), .B(new_n3871_), .ZN(new_n3972_));
  AOI21_X1   g03780(.A1(new_n3972_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n3973_));
  AOI21_X1   g03781(.A1(new_n3973_), .A2(new_n3961_), .B(new_n3945_), .ZN(new_n3974_));
  OAI21_X1   g03782(.A1(new_n3974_), .A2(new_n3962_), .B(\asqrt[60] ), .ZN(new_n3975_));
  NAND2_X1   g03783(.A1(new_n3975_), .A2(new_n218_), .ZN(new_n3976_));
  OAI21_X1   g03784(.A1(new_n3976_), .A2(new_n3964_), .B(new_n3971_), .ZN(new_n3977_));
  AOI21_X1   g03785(.A1(new_n3977_), .A2(new_n3965_), .B(new_n207_), .ZN(new_n3978_));
  NOR3_X1    g03786(.A1(new_n3782_), .A2(new_n3656_), .A3(new_n3690_), .ZN(new_n3979_));
  INV_X1     g03787(.I(new_n3979_), .ZN(new_n3980_));
  NOR3_X1    g03788(.A1(new_n3656_), .A2(new_n3690_), .A3(new_n3718_), .ZN(new_n3981_));
  AOI22_X1   g03789(.A1(new_n3980_), .A2(new_n3718_), .B1(\asqrt[41] ), .B2(new_n3981_), .ZN(new_n3982_));
  NOR3_X1    g03790(.A1(new_n3974_), .A2(new_n3962_), .A3(\asqrt[60] ), .ZN(new_n3983_));
  OAI21_X1   g03791(.A1(new_n3958_), .A2(new_n3983_), .B(new_n3975_), .ZN(new_n3984_));
  AOI21_X1   g03792(.A1(new_n3984_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n3985_));
  AOI21_X1   g03793(.A1(new_n3985_), .A2(new_n3977_), .B(new_n3982_), .ZN(new_n3986_));
  AND3_X2    g03794(.A1(new_n3668_), .A2(new_n3721_), .A3(new_n3672_), .Z(new_n3987_));
  NAND2_X1   g03795(.A1(\asqrt[41] ), .A2(new_n3987_), .ZN(new_n3988_));
  INV_X1     g03796(.I(new_n3988_), .ZN(new_n3989_));
  AND2_X2    g03797(.A1(new_n3668_), .A2(new_n3721_), .Z(new_n3990_));
  AOI21_X1   g03798(.A1(\asqrt[41] ), .A2(new_n3990_), .B(new_n3672_), .ZN(new_n3991_));
  NOR2_X1    g03799(.A1(new_n3989_), .A2(new_n3991_), .ZN(new_n3992_));
  NOR3_X1    g03800(.A1(new_n3782_), .A2(new_n3722_), .A3(new_n3712_), .ZN(new_n3993_));
  NOR3_X1    g03801(.A1(new_n3992_), .A2(new_n3735_), .A3(new_n3993_), .ZN(new_n3994_));
  OAI21_X1   g03802(.A1(new_n3986_), .A2(new_n3978_), .B(new_n3994_), .ZN(new_n3995_));
  NAND2_X1   g03803(.A1(new_n3995_), .A2(new_n193_), .ZN(new_n3996_));
  INV_X1     g03804(.I(new_n3982_), .ZN(new_n3997_));
  NAND3_X1   g03805(.A1(new_n3977_), .A2(new_n3965_), .A3(new_n207_), .ZN(new_n3998_));
  NAND2_X1   g03806(.A1(new_n3998_), .A2(new_n3997_), .ZN(new_n3999_));
  INV_X1     g03807(.I(new_n3992_), .ZN(new_n4000_));
  NOR2_X1    g03808(.A1(new_n3978_), .A2(new_n4000_), .ZN(new_n4001_));
  AOI21_X1   g03809(.A1(\asqrt[41] ), .A2(new_n3685_), .B(new_n3708_), .ZN(new_n4002_));
  OAI21_X1   g03810(.A1(new_n3722_), .A2(new_n3712_), .B(\asqrt[63] ), .ZN(new_n4003_));
  NOR2_X1    g03811(.A1(new_n4002_), .A2(new_n4003_), .ZN(new_n4004_));
  AND3_X2    g03812(.A1(new_n3684_), .A2(new_n3682_), .A3(new_n3698_), .Z(new_n4005_));
  NAND4_X1   g03813(.A1(new_n3736_), .A2(new_n3723_), .A3(new_n3695_), .A4(new_n4005_), .ZN(new_n4006_));
  INV_X1     g03814(.I(new_n4006_), .ZN(new_n4007_));
  NOR2_X1    g03815(.A1(new_n4004_), .A2(new_n4007_), .ZN(new_n4008_));
  INV_X1     g03816(.I(new_n4008_), .ZN(new_n4009_));
  AOI21_X1   g03817(.A1(new_n4001_), .A2(new_n3999_), .B(new_n4009_), .ZN(new_n4010_));
  NAND2_X1   g03818(.A1(new_n3996_), .A2(new_n4010_), .ZN(\asqrt[40] ));
  NOR2_X1    g03819(.A1(\a[78] ), .A2(\a[79] ), .ZN(new_n4012_));
  INV_X1     g03820(.I(new_n4012_), .ZN(new_n4013_));
  NOR2_X1    g03821(.A1(new_n4013_), .A2(\a[80] ), .ZN(new_n4014_));
  INV_X1     g03822(.I(new_n4014_), .ZN(new_n4015_));
  INV_X1     g03823(.I(new_n3958_), .ZN(new_n4016_));
  NAND2_X1   g03824(.A1(new_n3941_), .A2(new_n306_), .ZN(new_n4017_));
  OAI21_X1   g03825(.A1(new_n4017_), .A2(new_n3974_), .B(new_n4016_), .ZN(new_n4018_));
  AOI21_X1   g03826(.A1(new_n4018_), .A2(new_n3975_), .B(new_n218_), .ZN(new_n4019_));
  NOR3_X1    g03827(.A1(new_n3940_), .A2(\asqrt[59] ), .A3(new_n3931_), .ZN(new_n4020_));
  OAI21_X1   g03828(.A1(new_n3945_), .A2(new_n4020_), .B(new_n3941_), .ZN(new_n4021_));
  AOI21_X1   g03829(.A1(new_n4021_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n4022_));
  AOI21_X1   g03830(.A1(new_n4022_), .A2(new_n4018_), .B(new_n3970_), .ZN(new_n4023_));
  OAI21_X1   g03831(.A1(new_n4023_), .A2(new_n4019_), .B(\asqrt[62] ), .ZN(new_n4024_));
  NOR3_X1    g03832(.A1(new_n4023_), .A2(\asqrt[62] ), .A3(new_n4019_), .ZN(new_n4025_));
  OAI21_X1   g03833(.A1(new_n3982_), .A2(new_n4025_), .B(new_n4024_), .ZN(new_n4026_));
  AOI21_X1   g03834(.A1(new_n4026_), .A2(new_n3994_), .B(\asqrt[63] ), .ZN(new_n4027_));
  NAND2_X1   g03835(.A1(new_n4024_), .A2(new_n3992_), .ZN(new_n4028_));
  OAI21_X1   g03836(.A1(new_n4028_), .A2(new_n3986_), .B(new_n4008_), .ZN(new_n4029_));
  OAI21_X1   g03837(.A1(new_n4027_), .A2(new_n4029_), .B(\a[80] ), .ZN(new_n4030_));
  AOI21_X1   g03838(.A1(new_n4030_), .A2(new_n4015_), .B(new_n3782_), .ZN(new_n4031_));
  INV_X1     g03839(.I(\a[80] ), .ZN(new_n4032_));
  AOI21_X1   g03840(.A1(new_n3996_), .A2(new_n4010_), .B(new_n4032_), .ZN(new_n4033_));
  NAND2_X1   g03841(.A1(new_n3698_), .A2(new_n4015_), .ZN(new_n4034_));
  NOR4_X1    g03842(.A1(new_n3710_), .A2(new_n3735_), .A3(new_n3696_), .A4(new_n4034_), .ZN(new_n4035_));
  INV_X1     g03843(.I(new_n4035_), .ZN(new_n4036_));
  NOR2_X1    g03844(.A1(new_n4033_), .A2(new_n4036_), .ZN(new_n4037_));
  AOI21_X1   g03845(.A1(new_n3996_), .A2(new_n4010_), .B(new_n3705_), .ZN(new_n4038_));
  INV_X1     g03846(.I(\a[81] ), .ZN(new_n4039_));
  AOI21_X1   g03847(.A1(\asqrt[40] ), .A2(new_n4032_), .B(new_n4039_), .ZN(new_n4040_));
  NOR3_X1    g03848(.A1(new_n4037_), .A2(new_n4040_), .A3(new_n4038_), .ZN(new_n4041_));
  OAI21_X1   g03849(.A1(new_n4041_), .A2(new_n4031_), .B(\asqrt[42] ), .ZN(new_n4042_));
  OAI21_X1   g03850(.A1(new_n4027_), .A2(new_n4029_), .B(new_n3704_), .ZN(new_n4043_));
  NAND2_X1   g03851(.A1(new_n4001_), .A2(new_n3999_), .ZN(new_n4044_));
  INV_X1     g03852(.I(new_n4004_), .ZN(new_n4045_));
  NOR2_X1    g03853(.A1(new_n4007_), .A2(new_n3782_), .ZN(new_n4046_));
  NAND4_X1   g03854(.A1(new_n3996_), .A2(new_n4044_), .A3(new_n4045_), .A4(new_n4046_), .ZN(new_n4047_));
  AOI21_X1   g03855(.A1(new_n4047_), .A2(new_n4043_), .B(new_n3717_), .ZN(new_n4048_));
  INV_X1     g03856(.I(new_n4044_), .ZN(new_n4049_));
  NAND2_X1   g03857(.A1(new_n4045_), .A2(new_n4046_), .ZN(new_n4050_));
  NOR3_X1    g03858(.A1(new_n4049_), .A2(new_n4027_), .A3(new_n4050_), .ZN(new_n4051_));
  NOR3_X1    g03859(.A1(new_n4051_), .A2(new_n4038_), .A3(\a[82] ), .ZN(new_n4052_));
  OAI21_X1   g03860(.A1(new_n4033_), .A2(new_n4014_), .B(\asqrt[41] ), .ZN(new_n4053_));
  NAND2_X1   g03861(.A1(new_n4053_), .A2(new_n3419_), .ZN(new_n4054_));
  OAI22_X1   g03862(.A1(new_n4041_), .A2(new_n4054_), .B1(new_n4048_), .B2(new_n4052_), .ZN(new_n4055_));
  AOI21_X1   g03863(.A1(new_n4055_), .A2(new_n4042_), .B(new_n3218_), .ZN(new_n4056_));
  NOR3_X1    g03864(.A1(new_n3896_), .A2(new_n3716_), .A3(new_n3728_), .ZN(new_n4057_));
  NAND3_X1   g03865(.A1(\asqrt[40] ), .A2(new_n3752_), .A3(new_n3881_), .ZN(new_n4058_));
  AOI22_X1   g03866(.A1(new_n4058_), .A2(new_n3896_), .B1(\asqrt[40] ), .B2(new_n4057_), .ZN(new_n4059_));
  AOI21_X1   g03867(.A1(new_n3996_), .A2(new_n4010_), .B(\a[80] ), .ZN(new_n4060_));
  OAI21_X1   g03868(.A1(new_n4039_), .A2(new_n4060_), .B(new_n4043_), .ZN(new_n4061_));
  OAI21_X1   g03869(.A1(new_n4061_), .A2(new_n4037_), .B(new_n4053_), .ZN(new_n4062_));
  AOI21_X1   g03870(.A1(new_n4062_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n4063_));
  AOI21_X1   g03871(.A1(new_n4063_), .A2(new_n4055_), .B(new_n4059_), .ZN(new_n4064_));
  OAI21_X1   g03872(.A1(new_n4064_), .A2(new_n4056_), .B(\asqrt[44] ), .ZN(new_n4065_));
  INV_X1     g03873(.I(new_n4065_), .ZN(new_n4066_));
  NOR2_X1    g03874(.A1(new_n3739_), .A2(new_n3742_), .ZN(new_n4067_));
  NOR2_X1    g03875(.A1(new_n3732_), .A2(new_n3744_), .ZN(new_n4068_));
  INV_X1     g03876(.I(new_n4068_), .ZN(new_n4069_));
  NAND4_X1   g03877(.A1(\asqrt[40] ), .A2(new_n3733_), .A3(new_n4067_), .A4(new_n4069_), .ZN(new_n4070_));
  INV_X1     g03878(.I(\asqrt[40] ), .ZN(new_n4071_));
  NOR3_X1    g03879(.A1(new_n4071_), .A2(new_n3885_), .A3(new_n4068_), .ZN(new_n4072_));
  OAI21_X1   g03880(.A1(new_n4072_), .A2(new_n4067_), .B(new_n4070_), .ZN(new_n4073_));
  INV_X1     g03881(.I(new_n4073_), .ZN(new_n4074_));
  NOR3_X1    g03882(.A1(new_n4064_), .A2(new_n4056_), .A3(\asqrt[44] ), .ZN(new_n4075_));
  NOR2_X1    g03883(.A1(new_n4075_), .A2(new_n4074_), .ZN(new_n4076_));
  OAI21_X1   g03884(.A1(new_n4076_), .A2(new_n4066_), .B(\asqrt[45] ), .ZN(new_n4077_));
  NOR2_X1    g03885(.A1(new_n3898_), .A2(new_n3890_), .ZN(new_n4078_));
  NOR3_X1    g03886(.A1(new_n4071_), .A2(new_n3746_), .A3(new_n4078_), .ZN(new_n4079_));
  INV_X1     g03887(.I(new_n4079_), .ZN(new_n4080_));
  NOR3_X1    g03888(.A1(new_n4078_), .A2(new_n3746_), .A3(new_n3895_), .ZN(new_n4081_));
  AOI22_X1   g03889(.A1(new_n4080_), .A2(new_n3895_), .B1(\asqrt[40] ), .B2(new_n4081_), .ZN(new_n4082_));
  INV_X1     g03890(.I(new_n4082_), .ZN(new_n4083_));
  NAND2_X1   g03891(.A1(new_n4065_), .A2(new_n2641_), .ZN(new_n4084_));
  OAI21_X1   g03892(.A1(new_n4076_), .A2(new_n4084_), .B(new_n4083_), .ZN(new_n4085_));
  AOI21_X1   g03893(.A1(new_n4085_), .A2(new_n4077_), .B(new_n2465_), .ZN(new_n4086_));
  NOR3_X1    g03894(.A1(new_n3759_), .A2(new_n3767_), .A3(new_n3765_), .ZN(new_n4087_));
  NOR3_X1    g03895(.A1(new_n4071_), .A2(new_n3759_), .A3(new_n3767_), .ZN(new_n4088_));
  INV_X1     g03896(.I(new_n4088_), .ZN(new_n4089_));
  AOI22_X1   g03897(.A1(new_n4089_), .A2(new_n3765_), .B1(\asqrt[40] ), .B2(new_n4087_), .ZN(new_n4090_));
  OAI21_X1   g03898(.A1(new_n4074_), .A2(new_n4075_), .B(new_n4065_), .ZN(new_n4091_));
  AOI21_X1   g03899(.A1(new_n4091_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n4092_));
  AOI21_X1   g03900(.A1(new_n4092_), .A2(new_n4085_), .B(new_n4090_), .ZN(new_n4093_));
  OAI21_X1   g03901(.A1(new_n4093_), .A2(new_n4086_), .B(\asqrt[47] ), .ZN(new_n4094_));
  NAND2_X1   g03902(.A1(new_n3901_), .A2(new_n3893_), .ZN(new_n4095_));
  NAND3_X1   g03903(.A1(\asqrt[40] ), .A2(new_n3769_), .A3(new_n4095_), .ZN(new_n4096_));
  AND3_X2    g03904(.A1(new_n3769_), .A2(new_n3775_), .A3(new_n4095_), .Z(new_n4097_));
  AOI22_X1   g03905(.A1(new_n4096_), .A2(new_n3776_), .B1(\asqrt[40] ), .B2(new_n4097_), .ZN(new_n4098_));
  INV_X1     g03906(.I(new_n4098_), .ZN(new_n4099_));
  NAND2_X1   g03907(.A1(new_n4030_), .A2(new_n4035_), .ZN(new_n4100_));
  OAI21_X1   g03908(.A1(new_n4027_), .A2(new_n4029_), .B(new_n4032_), .ZN(new_n4101_));
  NAND2_X1   g03909(.A1(new_n4101_), .A2(\a[81] ), .ZN(new_n4102_));
  NAND3_X1   g03910(.A1(new_n4100_), .A2(new_n4102_), .A3(new_n4043_), .ZN(new_n4103_));
  AOI21_X1   g03911(.A1(new_n4103_), .A2(new_n4053_), .B(new_n3419_), .ZN(new_n4104_));
  OAI21_X1   g03912(.A1(new_n4051_), .A2(new_n4038_), .B(\a[82] ), .ZN(new_n4105_));
  NAND3_X1   g03913(.A1(new_n4047_), .A2(new_n4043_), .A3(new_n3717_), .ZN(new_n4106_));
  NAND2_X1   g03914(.A1(new_n4030_), .A2(new_n4015_), .ZN(new_n4107_));
  AOI21_X1   g03915(.A1(new_n4107_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n4108_));
  AOI22_X1   g03916(.A1(new_n4103_), .A2(new_n4108_), .B1(new_n4105_), .B2(new_n4106_), .ZN(new_n4109_));
  OAI21_X1   g03917(.A1(new_n4109_), .A2(new_n4104_), .B(\asqrt[43] ), .ZN(new_n4110_));
  NAND2_X1   g03918(.A1(new_n4110_), .A2(new_n2954_), .ZN(new_n4111_));
  OAI21_X1   g03919(.A1(new_n4111_), .A2(new_n4064_), .B(new_n4073_), .ZN(new_n4112_));
  AOI21_X1   g03920(.A1(new_n4112_), .A2(new_n4065_), .B(new_n2641_), .ZN(new_n4113_));
  INV_X1     g03921(.I(new_n4059_), .ZN(new_n4114_));
  AOI21_X1   g03922(.A1(\a[81] ), .A2(new_n4101_), .B(new_n4038_), .ZN(new_n4115_));
  AOI21_X1   g03923(.A1(new_n4115_), .A2(new_n4100_), .B(new_n4031_), .ZN(new_n4116_));
  OAI21_X1   g03924(.A1(new_n4116_), .A2(new_n3419_), .B(new_n3218_), .ZN(new_n4117_));
  OAI21_X1   g03925(.A1(new_n4117_), .A2(new_n4109_), .B(new_n4114_), .ZN(new_n4118_));
  NAND2_X1   g03926(.A1(new_n4118_), .A2(new_n4110_), .ZN(new_n4119_));
  AOI21_X1   g03927(.A1(new_n4119_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n4120_));
  AOI21_X1   g03928(.A1(new_n4120_), .A2(new_n4112_), .B(new_n4082_), .ZN(new_n4121_));
  OAI21_X1   g03929(.A1(new_n4121_), .A2(new_n4113_), .B(\asqrt[46] ), .ZN(new_n4122_));
  NAND2_X1   g03930(.A1(new_n4122_), .A2(new_n2229_), .ZN(new_n4123_));
  OAI21_X1   g03931(.A1(new_n4123_), .A2(new_n4093_), .B(new_n4099_), .ZN(new_n4124_));
  AOI21_X1   g03932(.A1(new_n4124_), .A2(new_n4094_), .B(new_n1956_), .ZN(new_n4125_));
  INV_X1     g03933(.I(new_n3785_), .ZN(new_n4126_));
  NOR3_X1    g03934(.A1(new_n3779_), .A2(new_n3912_), .A3(new_n4126_), .ZN(new_n4127_));
  NOR3_X1    g03935(.A1(new_n4071_), .A2(new_n3779_), .A3(new_n3912_), .ZN(new_n4128_));
  INV_X1     g03936(.I(new_n4128_), .ZN(new_n4129_));
  AOI22_X1   g03937(.A1(new_n4129_), .A2(new_n4126_), .B1(\asqrt[40] ), .B2(new_n4127_), .ZN(new_n4130_));
  NOR3_X1    g03938(.A1(new_n4121_), .A2(new_n4113_), .A3(\asqrt[46] ), .ZN(new_n4131_));
  OAI21_X1   g03939(.A1(new_n4090_), .A2(new_n4131_), .B(new_n4122_), .ZN(new_n4132_));
  AOI21_X1   g03940(.A1(new_n4132_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n4133_));
  AOI21_X1   g03941(.A1(new_n4133_), .A2(new_n4124_), .B(new_n4130_), .ZN(new_n4134_));
  OAI21_X1   g03942(.A1(new_n4134_), .A2(new_n4125_), .B(\asqrt[49] ), .ZN(new_n4135_));
  INV_X1     g03943(.I(new_n4135_), .ZN(new_n4136_));
  NOR3_X1    g03944(.A1(new_n4071_), .A2(new_n3790_), .A3(new_n3797_), .ZN(new_n4137_));
  INV_X1     g03945(.I(new_n4137_), .ZN(new_n4138_));
  NOR3_X1    g03946(.A1(new_n3790_), .A2(new_n3880_), .A3(new_n3797_), .ZN(new_n4139_));
  AOI22_X1   g03947(.A1(new_n4138_), .A2(new_n3880_), .B1(\asqrt[40] ), .B2(new_n4139_), .ZN(new_n4140_));
  NOR3_X1    g03948(.A1(new_n4134_), .A2(\asqrt[49] ), .A3(new_n4125_), .ZN(new_n4141_));
  NOR2_X1    g03949(.A1(new_n4141_), .A2(new_n4140_), .ZN(new_n4142_));
  OAI21_X1   g03950(.A1(new_n4142_), .A2(new_n4136_), .B(\asqrt[50] ), .ZN(new_n4143_));
  INV_X1     g03951(.I(new_n3906_), .ZN(new_n4144_));
  NOR3_X1    g03952(.A1(new_n4144_), .A2(new_n3911_), .A3(new_n3808_), .ZN(new_n4145_));
  NOR3_X1    g03953(.A1(new_n4071_), .A2(new_n3911_), .A3(new_n4144_), .ZN(new_n4146_));
  INV_X1     g03954(.I(new_n4146_), .ZN(new_n4147_));
  AOI22_X1   g03955(.A1(new_n4147_), .A2(new_n3808_), .B1(\asqrt[40] ), .B2(new_n4145_), .ZN(new_n4148_));
  INV_X1     g03956(.I(new_n4148_), .ZN(new_n4149_));
  NAND2_X1   g03957(.A1(new_n4135_), .A2(new_n1612_), .ZN(new_n4150_));
  OAI21_X1   g03958(.A1(new_n4142_), .A2(new_n4150_), .B(new_n4149_), .ZN(new_n4151_));
  AOI21_X1   g03959(.A1(new_n4151_), .A2(new_n4143_), .B(new_n1376_), .ZN(new_n4152_));
  INV_X1     g03960(.I(new_n3815_), .ZN(new_n4153_));
  NOR3_X1    g03961(.A1(new_n4071_), .A2(new_n3811_), .A3(new_n3916_), .ZN(new_n4154_));
  INV_X1     g03962(.I(new_n4154_), .ZN(new_n4155_));
  NOR3_X1    g03963(.A1(new_n3811_), .A2(new_n3916_), .A3(new_n4153_), .ZN(new_n4156_));
  AOI22_X1   g03964(.A1(new_n4155_), .A2(new_n4153_), .B1(\asqrt[40] ), .B2(new_n4156_), .ZN(new_n4157_));
  NOR3_X1    g03965(.A1(new_n4093_), .A2(new_n4086_), .A3(\asqrt[47] ), .ZN(new_n4158_));
  OAI21_X1   g03966(.A1(new_n4098_), .A2(new_n4158_), .B(new_n4094_), .ZN(new_n4159_));
  INV_X1     g03967(.I(new_n4130_), .ZN(new_n4160_));
  NAND3_X1   g03968(.A1(new_n4124_), .A2(new_n1956_), .A3(new_n4094_), .ZN(new_n4161_));
  AOI22_X1   g03969(.A1(new_n4161_), .A2(new_n4160_), .B1(new_n4159_), .B2(\asqrt[48] ), .ZN(new_n4162_));
  OAI22_X1   g03970(.A1(new_n4141_), .A2(new_n4140_), .B1(new_n4162_), .B2(new_n1806_), .ZN(new_n4163_));
  AOI21_X1   g03971(.A1(new_n4163_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n4164_));
  AOI21_X1   g03972(.A1(new_n4164_), .A2(new_n4151_), .B(new_n4157_), .ZN(new_n4165_));
  OAI21_X1   g03973(.A1(new_n4165_), .A2(new_n4152_), .B(\asqrt[52] ), .ZN(new_n4166_));
  INV_X1     g03974(.I(new_n4166_), .ZN(new_n4167_));
  INV_X1     g03975(.I(new_n4165_), .ZN(new_n4168_));
  NOR3_X1    g03976(.A1(new_n3820_), .A2(new_n3879_), .A3(new_n3826_), .ZN(new_n4169_));
  NOR3_X1    g03977(.A1(new_n4071_), .A2(new_n3820_), .A3(new_n3826_), .ZN(new_n4170_));
  INV_X1     g03978(.I(new_n4170_), .ZN(new_n4171_));
  AOI22_X1   g03979(.A1(new_n4171_), .A2(new_n3879_), .B1(\asqrt[40] ), .B2(new_n4169_), .ZN(new_n4172_));
  NOR2_X1    g03980(.A1(new_n4152_), .A2(\asqrt[52] ), .ZN(new_n4173_));
  AOI21_X1   g03981(.A1(new_n4168_), .A2(new_n4173_), .B(new_n4172_), .ZN(new_n4174_));
  OAI21_X1   g03982(.A1(new_n4174_), .A2(new_n4167_), .B(\asqrt[53] ), .ZN(new_n4175_));
  NOR2_X1    g03983(.A1(new_n3827_), .A2(new_n3835_), .ZN(new_n4176_));
  NOR3_X1    g03984(.A1(new_n4071_), .A2(new_n3910_), .A3(new_n4176_), .ZN(new_n4177_));
  INV_X1     g03985(.I(new_n4177_), .ZN(new_n4178_));
  NOR3_X1    g03986(.A1(new_n4176_), .A2(new_n3910_), .A3(new_n3834_), .ZN(new_n4179_));
  AOI22_X1   g03987(.A1(new_n4178_), .A2(new_n3834_), .B1(\asqrt[40] ), .B2(new_n4179_), .ZN(new_n4180_));
  INV_X1     g03988(.I(new_n4180_), .ZN(new_n4181_));
  NAND2_X1   g03989(.A1(new_n4166_), .A2(new_n1103_), .ZN(new_n4182_));
  OAI21_X1   g03990(.A1(new_n4182_), .A2(new_n4174_), .B(new_n4181_), .ZN(new_n4183_));
  AOI21_X1   g03991(.A1(new_n4183_), .A2(new_n4175_), .B(new_n904_), .ZN(new_n4184_));
  INV_X1     g03992(.I(new_n4184_), .ZN(new_n4185_));
  INV_X1     g03993(.I(new_n4183_), .ZN(new_n4186_));
  INV_X1     g03994(.I(new_n3841_), .ZN(new_n4187_));
  NOR3_X1    g03995(.A1(new_n3837_), .A2(new_n3924_), .A3(new_n4187_), .ZN(new_n4188_));
  NOR3_X1    g03996(.A1(new_n4071_), .A2(new_n3837_), .A3(new_n3924_), .ZN(new_n4189_));
  INV_X1     g03997(.I(new_n4189_), .ZN(new_n4190_));
  AOI22_X1   g03998(.A1(new_n4190_), .A2(new_n4187_), .B1(\asqrt[40] ), .B2(new_n4188_), .ZN(new_n4191_));
  INV_X1     g03999(.I(new_n4191_), .ZN(new_n4192_));
  NAND2_X1   g04000(.A1(new_n4175_), .A2(new_n904_), .ZN(new_n4193_));
  OAI21_X1   g04001(.A1(new_n4193_), .A2(new_n4186_), .B(new_n4192_), .ZN(new_n4194_));
  AOI21_X1   g04002(.A1(new_n4194_), .A2(new_n4185_), .B(new_n823_), .ZN(new_n4195_));
  NOR3_X1    g04003(.A1(new_n4071_), .A2(new_n3846_), .A3(new_n3852_), .ZN(new_n4196_));
  INV_X1     g04004(.I(new_n4196_), .ZN(new_n4197_));
  NOR3_X1    g04005(.A1(new_n3846_), .A2(new_n3878_), .A3(new_n3852_), .ZN(new_n4198_));
  AOI22_X1   g04006(.A1(new_n4197_), .A2(new_n3878_), .B1(\asqrt[40] ), .B2(new_n4198_), .ZN(new_n4199_));
  NOR2_X1    g04007(.A1(new_n4184_), .A2(\asqrt[55] ), .ZN(new_n4200_));
  AOI21_X1   g04008(.A1(new_n4200_), .A2(new_n4194_), .B(new_n4199_), .ZN(new_n4201_));
  OAI21_X1   g04009(.A1(new_n4201_), .A2(new_n4195_), .B(\asqrt[56] ), .ZN(new_n4202_));
  NOR2_X1    g04010(.A1(new_n3853_), .A2(new_n3861_), .ZN(new_n4203_));
  NOR3_X1    g04011(.A1(new_n4203_), .A2(new_n3923_), .A3(new_n3860_), .ZN(new_n4204_));
  NOR3_X1    g04012(.A1(new_n4071_), .A2(new_n3923_), .A3(new_n4203_), .ZN(new_n4205_));
  INV_X1     g04013(.I(new_n4205_), .ZN(new_n4206_));
  AOI22_X1   g04014(.A1(new_n4206_), .A2(new_n3860_), .B1(\asqrt[40] ), .B2(new_n4204_), .ZN(new_n4207_));
  INV_X1     g04015(.I(new_n4207_), .ZN(new_n4208_));
  NOR3_X1    g04016(.A1(new_n4165_), .A2(new_n4152_), .A3(\asqrt[52] ), .ZN(new_n4209_));
  OAI21_X1   g04017(.A1(new_n4172_), .A2(new_n4209_), .B(new_n4166_), .ZN(new_n4210_));
  AOI21_X1   g04018(.A1(new_n4210_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n4211_));
  AOI21_X1   g04019(.A1(new_n4211_), .A2(new_n4183_), .B(new_n4191_), .ZN(new_n4212_));
  OAI21_X1   g04020(.A1(new_n4212_), .A2(new_n4184_), .B(\asqrt[55] ), .ZN(new_n4213_));
  NAND2_X1   g04021(.A1(new_n4213_), .A2(new_n703_), .ZN(new_n4214_));
  OAI21_X1   g04022(.A1(new_n4214_), .A2(new_n4201_), .B(new_n4208_), .ZN(new_n4215_));
  AOI21_X1   g04023(.A1(new_n4215_), .A2(new_n4202_), .B(new_n531_), .ZN(new_n4216_));
  INV_X1     g04024(.I(new_n4216_), .ZN(new_n4217_));
  INV_X1     g04025(.I(new_n4215_), .ZN(new_n4218_));
  INV_X1     g04026(.I(new_n3867_), .ZN(new_n4219_));
  NOR3_X1    g04027(.A1(new_n4071_), .A2(new_n3863_), .A3(new_n3937_), .ZN(new_n4220_));
  INV_X1     g04028(.I(new_n4220_), .ZN(new_n4221_));
  NOR3_X1    g04029(.A1(new_n3863_), .A2(new_n3937_), .A3(new_n4219_), .ZN(new_n4222_));
  AOI22_X1   g04030(.A1(new_n4221_), .A2(new_n4219_), .B1(\asqrt[40] ), .B2(new_n4222_), .ZN(new_n4223_));
  INV_X1     g04031(.I(new_n4223_), .ZN(new_n4224_));
  NAND2_X1   g04032(.A1(new_n4202_), .A2(new_n531_), .ZN(new_n4225_));
  OAI21_X1   g04033(.A1(new_n4225_), .A2(new_n4218_), .B(new_n4224_), .ZN(new_n4226_));
  AOI21_X1   g04034(.A1(new_n4226_), .A2(new_n4217_), .B(new_n436_), .ZN(new_n4227_));
  NOR3_X1    g04035(.A1(new_n3947_), .A2(new_n3877_), .A3(new_n3948_), .ZN(new_n4228_));
  NOR3_X1    g04036(.A1(new_n4071_), .A2(new_n3947_), .A3(new_n3948_), .ZN(new_n4229_));
  INV_X1     g04037(.I(new_n4229_), .ZN(new_n4230_));
  AOI22_X1   g04038(.A1(new_n4230_), .A2(new_n3877_), .B1(\asqrt[40] ), .B2(new_n4228_), .ZN(new_n4231_));
  NOR2_X1    g04039(.A1(new_n4216_), .A2(\asqrt[58] ), .ZN(new_n4232_));
  AOI21_X1   g04040(.A1(new_n4232_), .A2(new_n4226_), .B(new_n4231_), .ZN(new_n4233_));
  OAI21_X1   g04041(.A1(new_n4233_), .A2(new_n4227_), .B(\asqrt[59] ), .ZN(new_n4234_));
  NOR2_X1    g04042(.A1(new_n3949_), .A2(new_n3960_), .ZN(new_n4235_));
  NOR3_X1    g04043(.A1(new_n4071_), .A2(new_n3931_), .A3(new_n4235_), .ZN(new_n4236_));
  INV_X1     g04044(.I(new_n4236_), .ZN(new_n4237_));
  NOR3_X1    g04045(.A1(new_n4235_), .A2(new_n3931_), .A3(new_n3959_), .ZN(new_n4238_));
  AOI22_X1   g04046(.A1(new_n4237_), .A2(new_n3959_), .B1(\asqrt[40] ), .B2(new_n4238_), .ZN(new_n4239_));
  INV_X1     g04047(.I(new_n4239_), .ZN(new_n4240_));
  NOR3_X1    g04048(.A1(new_n4212_), .A2(\asqrt[55] ), .A3(new_n4184_), .ZN(new_n4241_));
  OAI21_X1   g04049(.A1(new_n4199_), .A2(new_n4241_), .B(new_n4213_), .ZN(new_n4242_));
  AOI21_X1   g04050(.A1(new_n4242_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n4243_));
  AOI21_X1   g04051(.A1(new_n4243_), .A2(new_n4215_), .B(new_n4223_), .ZN(new_n4244_));
  OAI21_X1   g04052(.A1(new_n4244_), .A2(new_n4216_), .B(\asqrt[58] ), .ZN(new_n4245_));
  NAND2_X1   g04053(.A1(new_n4245_), .A2(new_n327_), .ZN(new_n4246_));
  OAI21_X1   g04054(.A1(new_n4246_), .A2(new_n4233_), .B(new_n4240_), .ZN(new_n4247_));
  AOI21_X1   g04055(.A1(new_n4247_), .A2(new_n4234_), .B(new_n306_), .ZN(new_n4248_));
  INV_X1     g04056(.I(new_n4248_), .ZN(new_n4249_));
  INV_X1     g04057(.I(new_n4247_), .ZN(new_n4250_));
  NOR3_X1    g04058(.A1(new_n3962_), .A2(new_n4020_), .A3(new_n3946_), .ZN(new_n4251_));
  NOR3_X1    g04059(.A1(new_n4071_), .A2(new_n3962_), .A3(new_n4020_), .ZN(new_n4252_));
  INV_X1     g04060(.I(new_n4252_), .ZN(new_n4253_));
  AOI22_X1   g04061(.A1(new_n4253_), .A2(new_n3946_), .B1(\asqrt[40] ), .B2(new_n4251_), .ZN(new_n4254_));
  INV_X1     g04062(.I(new_n4254_), .ZN(new_n4255_));
  NAND2_X1   g04063(.A1(new_n4234_), .A2(new_n306_), .ZN(new_n4256_));
  OAI21_X1   g04064(.A1(new_n4250_), .A2(new_n4256_), .B(new_n4255_), .ZN(new_n4257_));
  AOI21_X1   g04065(.A1(new_n4257_), .A2(new_n4249_), .B(new_n218_), .ZN(new_n4258_));
  NOR3_X1    g04066(.A1(new_n4071_), .A2(new_n3953_), .A3(new_n3983_), .ZN(new_n4259_));
  INV_X1     g04067(.I(new_n4259_), .ZN(new_n4260_));
  NOR3_X1    g04068(.A1(new_n3953_), .A2(new_n3983_), .A3(new_n4016_), .ZN(new_n4261_));
  AOI22_X1   g04069(.A1(new_n4260_), .A2(new_n4016_), .B1(\asqrt[40] ), .B2(new_n4261_), .ZN(new_n4262_));
  NOR2_X1    g04070(.A1(new_n4248_), .A2(\asqrt[61] ), .ZN(new_n4263_));
  AOI21_X1   g04071(.A1(new_n4263_), .A2(new_n4257_), .B(new_n4262_), .ZN(new_n4264_));
  OAI21_X1   g04072(.A1(new_n4264_), .A2(new_n4258_), .B(\asqrt[62] ), .ZN(new_n4265_));
  NOR2_X1    g04073(.A1(new_n3976_), .A2(new_n3964_), .ZN(new_n4266_));
  NOR3_X1    g04074(.A1(new_n4266_), .A2(new_n4019_), .A3(new_n3971_), .ZN(new_n4267_));
  NOR3_X1    g04075(.A1(new_n4071_), .A2(new_n4019_), .A3(new_n4266_), .ZN(new_n4268_));
  INV_X1     g04076(.I(new_n4268_), .ZN(new_n4269_));
  AOI22_X1   g04077(.A1(new_n4269_), .A2(new_n3971_), .B1(\asqrt[40] ), .B2(new_n4267_), .ZN(new_n4270_));
  INV_X1     g04078(.I(new_n4270_), .ZN(new_n4271_));
  NOR3_X1    g04079(.A1(new_n4244_), .A2(\asqrt[58] ), .A3(new_n4216_), .ZN(new_n4272_));
  OAI21_X1   g04080(.A1(new_n4231_), .A2(new_n4272_), .B(new_n4245_), .ZN(new_n4273_));
  AOI21_X1   g04081(.A1(new_n4273_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n4274_));
  AOI21_X1   g04082(.A1(new_n4274_), .A2(new_n4247_), .B(new_n4254_), .ZN(new_n4275_));
  OAI21_X1   g04083(.A1(new_n4275_), .A2(new_n4248_), .B(\asqrt[61] ), .ZN(new_n4276_));
  NAND2_X1   g04084(.A1(new_n4276_), .A2(new_n207_), .ZN(new_n4277_));
  OAI21_X1   g04085(.A1(new_n4277_), .A2(new_n4264_), .B(new_n4271_), .ZN(new_n4278_));
  NAND4_X1   g04086(.A1(\asqrt[40] ), .A2(new_n4024_), .A3(new_n3982_), .A4(new_n3998_), .ZN(new_n4279_));
  NAND2_X1   g04087(.A1(new_n4024_), .A2(new_n3998_), .ZN(new_n4280_));
  OAI21_X1   g04088(.A1(new_n4071_), .A2(new_n4280_), .B(new_n3997_), .ZN(new_n4281_));
  NAND2_X1   g04089(.A1(new_n4281_), .A2(new_n4279_), .ZN(new_n4282_));
  AOI21_X1   g04090(.A1(new_n3999_), .A2(new_n4024_), .B(new_n3992_), .ZN(new_n4283_));
  AOI21_X1   g04091(.A1(\asqrt[40] ), .A2(new_n4283_), .B(new_n4049_), .ZN(new_n4284_));
  NAND2_X1   g04092(.A1(new_n4282_), .A2(new_n4284_), .ZN(new_n4285_));
  AOI21_X1   g04093(.A1(new_n4278_), .A2(new_n4265_), .B(new_n4285_), .ZN(new_n4286_));
  NOR3_X1    g04094(.A1(new_n4275_), .A2(\asqrt[61] ), .A3(new_n4248_), .ZN(new_n4287_));
  OAI21_X1   g04095(.A1(new_n4262_), .A2(new_n4287_), .B(new_n4276_), .ZN(new_n4288_));
  AOI21_X1   g04096(.A1(new_n4288_), .A2(\asqrt[62] ), .B(new_n4282_), .ZN(new_n4289_));
  AOI21_X1   g04097(.A1(\asqrt[40] ), .A2(new_n4000_), .B(new_n4026_), .ZN(new_n4290_));
  OR3_X2     g04098(.A1(new_n4290_), .A2(new_n193_), .A3(new_n4283_), .Z(new_n4291_));
  NAND2_X1   g04099(.A1(new_n3988_), .A2(new_n4006_), .ZN(new_n4292_));
  NOR4_X1    g04100(.A1(new_n4049_), .A2(new_n3991_), .A3(new_n4004_), .A4(new_n4292_), .ZN(new_n4293_));
  NAND2_X1   g04101(.A1(new_n4293_), .A2(new_n3996_), .ZN(new_n4294_));
  NAND2_X1   g04102(.A1(new_n4291_), .A2(new_n4294_), .ZN(new_n4295_));
  AOI21_X1   g04103(.A1(new_n4289_), .A2(new_n4278_), .B(new_n4295_), .ZN(new_n4296_));
  OAI21_X1   g04104(.A1(\asqrt[63] ), .A2(new_n4286_), .B(new_n4296_), .ZN(\asqrt[39] ));
  INV_X1     g04105(.I(\asqrt[39] ), .ZN(new_n4298_));
  NOR2_X1    g04106(.A1(\a[76] ), .A2(\a[77] ), .ZN(new_n4299_));
  INV_X1     g04107(.I(new_n4299_), .ZN(new_n4300_));
  NOR2_X1    g04108(.A1(new_n4300_), .A2(\a[78] ), .ZN(new_n4301_));
  INV_X1     g04109(.I(\a[78] ), .ZN(new_n4302_));
  INV_X1     g04110(.I(new_n4262_), .ZN(new_n4303_));
  INV_X1     g04111(.I(new_n4231_), .ZN(new_n4304_));
  INV_X1     g04112(.I(new_n4199_), .ZN(new_n4305_));
  INV_X1     g04113(.I(new_n4172_), .ZN(new_n4306_));
  INV_X1     g04114(.I(new_n4140_), .ZN(new_n4307_));
  INV_X1     g04115(.I(new_n4090_), .ZN(new_n4308_));
  NAND2_X1   g04116(.A1(new_n4077_), .A2(new_n2465_), .ZN(new_n4309_));
  OAI21_X1   g04117(.A1(new_n4309_), .A2(new_n4121_), .B(new_n4308_), .ZN(new_n4310_));
  AOI21_X1   g04118(.A1(new_n4310_), .A2(new_n4122_), .B(new_n2229_), .ZN(new_n4311_));
  NOR2_X1    g04119(.A1(new_n4086_), .A2(\asqrt[47] ), .ZN(new_n4312_));
  AOI21_X1   g04120(.A1(new_n4312_), .A2(new_n4310_), .B(new_n4098_), .ZN(new_n4313_));
  OAI21_X1   g04121(.A1(new_n4313_), .A2(new_n4311_), .B(\asqrt[48] ), .ZN(new_n4314_));
  NAND2_X1   g04122(.A1(new_n4314_), .A2(new_n1806_), .ZN(new_n4315_));
  OAI21_X1   g04123(.A1(new_n4315_), .A2(new_n4134_), .B(new_n4307_), .ZN(new_n4316_));
  AOI21_X1   g04124(.A1(new_n4316_), .A2(new_n4135_), .B(new_n1612_), .ZN(new_n4317_));
  NAND3_X1   g04125(.A1(new_n4316_), .A2(new_n1612_), .A3(new_n4135_), .ZN(new_n4318_));
  AOI21_X1   g04126(.A1(new_n4149_), .A2(new_n4318_), .B(new_n4317_), .ZN(new_n4319_));
  OAI21_X1   g04127(.A1(new_n4319_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n4320_));
  OAI21_X1   g04128(.A1(new_n4320_), .A2(new_n4165_), .B(new_n4306_), .ZN(new_n4321_));
  NAND3_X1   g04129(.A1(new_n4321_), .A2(new_n1103_), .A3(new_n4166_), .ZN(new_n4322_));
  AOI22_X1   g04130(.A1(new_n4322_), .A2(new_n4181_), .B1(\asqrt[53] ), .B2(new_n4210_), .ZN(new_n4323_));
  OAI21_X1   g04131(.A1(new_n4323_), .A2(new_n904_), .B(new_n823_), .ZN(new_n4324_));
  OAI21_X1   g04132(.A1(new_n4324_), .A2(new_n4212_), .B(new_n4305_), .ZN(new_n4325_));
  NAND3_X1   g04133(.A1(new_n4325_), .A2(new_n703_), .A3(new_n4213_), .ZN(new_n4326_));
  AOI22_X1   g04134(.A1(new_n4326_), .A2(new_n4208_), .B1(new_n4242_), .B2(\asqrt[56] ), .ZN(new_n4327_));
  OAI21_X1   g04135(.A1(new_n4327_), .A2(new_n531_), .B(new_n436_), .ZN(new_n4328_));
  OAI21_X1   g04136(.A1(new_n4328_), .A2(new_n4244_), .B(new_n4304_), .ZN(new_n4329_));
  NAND3_X1   g04137(.A1(new_n4329_), .A2(new_n327_), .A3(new_n4245_), .ZN(new_n4330_));
  AOI22_X1   g04138(.A1(new_n4330_), .A2(new_n4240_), .B1(new_n4273_), .B2(\asqrt[59] ), .ZN(new_n4331_));
  OAI21_X1   g04139(.A1(new_n4331_), .A2(new_n306_), .B(new_n218_), .ZN(new_n4332_));
  OAI21_X1   g04140(.A1(new_n4332_), .A2(new_n4275_), .B(new_n4303_), .ZN(new_n4333_));
  NAND3_X1   g04141(.A1(new_n4333_), .A2(new_n207_), .A3(new_n4276_), .ZN(new_n4334_));
  AOI22_X1   g04142(.A1(new_n4334_), .A2(new_n4271_), .B1(new_n4288_), .B2(\asqrt[62] ), .ZN(new_n4335_));
  OAI21_X1   g04143(.A1(new_n4335_), .A2(new_n4285_), .B(new_n193_), .ZN(new_n4336_));
  AOI21_X1   g04144(.A1(new_n4336_), .A2(new_n4296_), .B(new_n4302_), .ZN(new_n4337_));
  OAI21_X1   g04145(.A1(new_n4337_), .A2(new_n4301_), .B(\asqrt[40] ), .ZN(new_n4338_));
  INV_X1     g04146(.I(new_n4338_), .ZN(new_n4339_));
  NOR2_X1    g04147(.A1(new_n4007_), .A2(new_n4301_), .ZN(new_n4340_));
  NAND4_X1   g04148(.A1(new_n3996_), .A2(new_n4044_), .A3(new_n4045_), .A4(new_n4340_), .ZN(new_n4341_));
  NOR2_X1    g04149(.A1(new_n4337_), .A2(new_n4341_), .ZN(new_n4342_));
  AOI21_X1   g04150(.A1(new_n4336_), .A2(new_n4296_), .B(new_n4013_), .ZN(new_n4343_));
  INV_X1     g04151(.I(\a[79] ), .ZN(new_n4344_));
  AOI21_X1   g04152(.A1(\asqrt[39] ), .A2(new_n4302_), .B(new_n4344_), .ZN(new_n4345_));
  NOR3_X1    g04153(.A1(new_n4342_), .A2(new_n4345_), .A3(new_n4343_), .ZN(new_n4346_));
  OAI21_X1   g04154(.A1(new_n4346_), .A2(new_n4339_), .B(\asqrt[41] ), .ZN(new_n4347_));
  NOR2_X1    g04155(.A1(new_n4286_), .A2(\asqrt[63] ), .ZN(new_n4348_));
  INV_X1     g04156(.I(new_n4278_), .ZN(new_n4349_));
  INV_X1     g04157(.I(new_n4282_), .ZN(new_n4350_));
  NAND2_X1   g04158(.A1(new_n4265_), .A2(new_n4350_), .ZN(new_n4351_));
  INV_X1     g04159(.I(new_n4295_), .ZN(new_n4352_));
  OAI21_X1   g04160(.A1(new_n4349_), .A2(new_n4351_), .B(new_n4352_), .ZN(new_n4353_));
  OAI21_X1   g04161(.A1(new_n4348_), .A2(new_n4353_), .B(new_n4012_), .ZN(new_n4354_));
  NOR2_X1    g04162(.A1(new_n4349_), .A2(new_n4351_), .ZN(new_n4355_));
  OAI21_X1   g04163(.A1(new_n4293_), .A2(new_n4010_), .B(new_n3996_), .ZN(new_n4356_));
  NAND2_X1   g04164(.A1(new_n4291_), .A2(new_n4356_), .ZN(new_n4357_));
  NOR3_X1    g04165(.A1(new_n4348_), .A2(new_n4355_), .A3(new_n4357_), .ZN(new_n4358_));
  INV_X1     g04166(.I(new_n4358_), .ZN(new_n4359_));
  AOI21_X1   g04167(.A1(new_n4359_), .A2(new_n4354_), .B(new_n4032_), .ZN(new_n4360_));
  NOR3_X1    g04168(.A1(new_n4358_), .A2(new_n4343_), .A3(\a[80] ), .ZN(new_n4361_));
  AOI21_X1   g04169(.A1(\asqrt[39] ), .A2(\a[78] ), .B(new_n4301_), .ZN(new_n4362_));
  OAI21_X1   g04170(.A1(new_n4362_), .A2(new_n4071_), .B(new_n3782_), .ZN(new_n4363_));
  OAI22_X1   g04171(.A1(new_n4346_), .A2(new_n4363_), .B1(new_n4360_), .B2(new_n4361_), .ZN(new_n4364_));
  AOI21_X1   g04172(.A1(new_n4364_), .A2(new_n4347_), .B(new_n3419_), .ZN(new_n4365_));
  NOR3_X1    g04173(.A1(new_n4115_), .A2(new_n4031_), .A3(new_n4037_), .ZN(new_n4366_));
  NAND3_X1   g04174(.A1(\asqrt[39] ), .A2(new_n4053_), .A3(new_n4100_), .ZN(new_n4367_));
  AOI22_X1   g04175(.A1(new_n4367_), .A2(new_n4115_), .B1(\asqrt[39] ), .B2(new_n4366_), .ZN(new_n4368_));
  AOI21_X1   g04176(.A1(new_n4336_), .A2(new_n4296_), .B(\a[78] ), .ZN(new_n4369_));
  OAI21_X1   g04177(.A1(new_n4344_), .A2(new_n4369_), .B(new_n4354_), .ZN(new_n4370_));
  OAI21_X1   g04178(.A1(new_n4370_), .A2(new_n4342_), .B(new_n4338_), .ZN(new_n4371_));
  AOI21_X1   g04179(.A1(new_n4371_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n4372_));
  AOI21_X1   g04180(.A1(new_n4372_), .A2(new_n4364_), .B(new_n4368_), .ZN(new_n4373_));
  OAI21_X1   g04181(.A1(new_n4373_), .A2(new_n4365_), .B(\asqrt[43] ), .ZN(new_n4374_));
  INV_X1     g04182(.I(new_n4374_), .ZN(new_n4375_));
  NOR2_X1    g04183(.A1(new_n4052_), .A2(new_n4048_), .ZN(new_n4376_));
  INV_X1     g04184(.I(new_n4376_), .ZN(new_n4377_));
  NOR2_X1    g04185(.A1(new_n4041_), .A2(new_n4054_), .ZN(new_n4378_));
  NOR3_X1    g04186(.A1(new_n4104_), .A2(new_n4377_), .A3(new_n4378_), .ZN(new_n4379_));
  NOR3_X1    g04187(.A1(new_n4298_), .A2(new_n4104_), .A3(new_n4378_), .ZN(new_n4380_));
  INV_X1     g04188(.I(new_n4380_), .ZN(new_n4381_));
  AOI22_X1   g04189(.A1(new_n4381_), .A2(new_n4377_), .B1(\asqrt[39] ), .B2(new_n4379_), .ZN(new_n4382_));
  NOR3_X1    g04190(.A1(new_n4373_), .A2(new_n4365_), .A3(\asqrt[43] ), .ZN(new_n4383_));
  NOR2_X1    g04191(.A1(new_n4383_), .A2(new_n4382_), .ZN(new_n4384_));
  OAI21_X1   g04192(.A1(new_n4384_), .A2(new_n4375_), .B(\asqrt[44] ), .ZN(new_n4385_));
  NOR2_X1    g04193(.A1(new_n4117_), .A2(new_n4109_), .ZN(new_n4386_));
  NOR3_X1    g04194(.A1(new_n4298_), .A2(new_n4056_), .A3(new_n4386_), .ZN(new_n4387_));
  INV_X1     g04195(.I(new_n4387_), .ZN(new_n4388_));
  NOR3_X1    g04196(.A1(new_n4386_), .A2(new_n4056_), .A3(new_n4114_), .ZN(new_n4389_));
  AOI22_X1   g04197(.A1(new_n4388_), .A2(new_n4114_), .B1(\asqrt[39] ), .B2(new_n4389_), .ZN(new_n4390_));
  INV_X1     g04198(.I(new_n4390_), .ZN(new_n4391_));
  NAND2_X1   g04199(.A1(new_n4374_), .A2(new_n2954_), .ZN(new_n4392_));
  OAI21_X1   g04200(.A1(new_n4384_), .A2(new_n4392_), .B(new_n4391_), .ZN(new_n4393_));
  AOI21_X1   g04201(.A1(new_n4393_), .A2(new_n4385_), .B(new_n2641_), .ZN(new_n4394_));
  NOR3_X1    g04202(.A1(new_n4066_), .A2(new_n4075_), .A3(new_n4073_), .ZN(new_n4395_));
  NOR3_X1    g04203(.A1(new_n4298_), .A2(new_n4066_), .A3(new_n4075_), .ZN(new_n4396_));
  INV_X1     g04204(.I(new_n4396_), .ZN(new_n4397_));
  AOI22_X1   g04205(.A1(new_n4397_), .A2(new_n4073_), .B1(\asqrt[39] ), .B2(new_n4395_), .ZN(new_n4398_));
  OAI21_X1   g04206(.A1(new_n4382_), .A2(new_n4383_), .B(new_n4374_), .ZN(new_n4399_));
  AOI21_X1   g04207(.A1(new_n4399_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n4400_));
  AOI21_X1   g04208(.A1(new_n4400_), .A2(new_n4393_), .B(new_n4398_), .ZN(new_n4401_));
  OAI21_X1   g04209(.A1(new_n4401_), .A2(new_n4394_), .B(\asqrt[46] ), .ZN(new_n4402_));
  INV_X1     g04210(.I(new_n4402_), .ZN(new_n4403_));
  NOR2_X1    g04211(.A1(new_n4076_), .A2(new_n4084_), .ZN(new_n4404_));
  NOR3_X1    g04212(.A1(new_n4298_), .A2(new_n4113_), .A3(new_n4404_), .ZN(new_n4405_));
  INV_X1     g04213(.I(new_n4405_), .ZN(new_n4406_));
  NOR3_X1    g04214(.A1(new_n4404_), .A2(new_n4113_), .A3(new_n4083_), .ZN(new_n4407_));
  AOI22_X1   g04215(.A1(new_n4406_), .A2(new_n4083_), .B1(\asqrt[39] ), .B2(new_n4407_), .ZN(new_n4408_));
  NOR3_X1    g04216(.A1(new_n4401_), .A2(new_n4394_), .A3(\asqrt[46] ), .ZN(new_n4409_));
  NOR2_X1    g04217(.A1(new_n4409_), .A2(new_n4408_), .ZN(new_n4410_));
  OAI21_X1   g04218(.A1(new_n4410_), .A2(new_n4403_), .B(\asqrt[47] ), .ZN(new_n4411_));
  NOR3_X1    g04219(.A1(new_n4086_), .A2(new_n4131_), .A3(new_n4308_), .ZN(new_n4412_));
  NOR3_X1    g04220(.A1(new_n4298_), .A2(new_n4086_), .A3(new_n4131_), .ZN(new_n4413_));
  INV_X1     g04221(.I(new_n4413_), .ZN(new_n4414_));
  AOI22_X1   g04222(.A1(new_n4414_), .A2(new_n4308_), .B1(\asqrt[39] ), .B2(new_n4412_), .ZN(new_n4415_));
  INV_X1     g04223(.I(new_n4415_), .ZN(new_n4416_));
  NAND2_X1   g04224(.A1(new_n4402_), .A2(new_n2229_), .ZN(new_n4417_));
  OAI21_X1   g04225(.A1(new_n4410_), .A2(new_n4417_), .B(new_n4416_), .ZN(new_n4418_));
  AOI21_X1   g04226(.A1(new_n4418_), .A2(new_n4411_), .B(new_n1956_), .ZN(new_n4419_));
  NOR3_X1    g04227(.A1(new_n4298_), .A2(new_n4311_), .A3(new_n4158_), .ZN(new_n4420_));
  INV_X1     g04228(.I(new_n4420_), .ZN(new_n4421_));
  NOR3_X1    g04229(.A1(new_n4311_), .A2(new_n4099_), .A3(new_n4158_), .ZN(new_n4422_));
  AOI22_X1   g04230(.A1(new_n4421_), .A2(new_n4099_), .B1(\asqrt[39] ), .B2(new_n4422_), .ZN(new_n4423_));
  OAI21_X1   g04231(.A1(new_n4408_), .A2(new_n4409_), .B(new_n4402_), .ZN(new_n4424_));
  AOI21_X1   g04232(.A1(new_n4424_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n4425_));
  AOI21_X1   g04233(.A1(new_n4425_), .A2(new_n4418_), .B(new_n4423_), .ZN(new_n4426_));
  OAI21_X1   g04234(.A1(new_n4426_), .A2(new_n4419_), .B(\asqrt[49] ), .ZN(new_n4427_));
  INV_X1     g04235(.I(new_n4427_), .ZN(new_n4428_));
  AND3_X2    g04236(.A1(new_n4314_), .A2(new_n4130_), .A3(new_n4161_), .Z(new_n4429_));
  NAND3_X1   g04237(.A1(\asqrt[39] ), .A2(new_n4314_), .A3(new_n4161_), .ZN(new_n4430_));
  AOI22_X1   g04238(.A1(new_n4430_), .A2(new_n4160_), .B1(\asqrt[39] ), .B2(new_n4429_), .ZN(new_n4431_));
  NOR3_X1    g04239(.A1(new_n4426_), .A2(new_n4419_), .A3(\asqrt[49] ), .ZN(new_n4432_));
  NOR2_X1    g04240(.A1(new_n4432_), .A2(new_n4431_), .ZN(new_n4433_));
  OAI21_X1   g04241(.A1(new_n4433_), .A2(new_n4428_), .B(\asqrt[50] ), .ZN(new_n4434_));
  NOR3_X1    g04242(.A1(new_n4298_), .A2(new_n4136_), .A3(new_n4141_), .ZN(new_n4435_));
  INV_X1     g04243(.I(new_n4435_), .ZN(new_n4436_));
  NOR3_X1    g04244(.A1(new_n4136_), .A2(new_n4307_), .A3(new_n4141_), .ZN(new_n4437_));
  AOI22_X1   g04245(.A1(new_n4436_), .A2(new_n4307_), .B1(\asqrt[39] ), .B2(new_n4437_), .ZN(new_n4438_));
  INV_X1     g04246(.I(new_n4438_), .ZN(new_n4439_));
  NAND2_X1   g04247(.A1(new_n4427_), .A2(new_n1612_), .ZN(new_n4440_));
  OAI21_X1   g04248(.A1(new_n4433_), .A2(new_n4440_), .B(new_n4439_), .ZN(new_n4441_));
  AOI21_X1   g04249(.A1(new_n4441_), .A2(new_n4434_), .B(new_n1376_), .ZN(new_n4442_));
  NOR2_X1    g04250(.A1(new_n4142_), .A2(new_n4150_), .ZN(new_n4443_));
  NOR3_X1    g04251(.A1(new_n4443_), .A2(new_n4317_), .A3(new_n4149_), .ZN(new_n4444_));
  NOR3_X1    g04252(.A1(new_n4298_), .A2(new_n4317_), .A3(new_n4443_), .ZN(new_n4445_));
  INV_X1     g04253(.I(new_n4445_), .ZN(new_n4446_));
  AOI22_X1   g04254(.A1(new_n4446_), .A2(new_n4149_), .B1(\asqrt[39] ), .B2(new_n4444_), .ZN(new_n4447_));
  OAI21_X1   g04255(.A1(new_n4431_), .A2(new_n4432_), .B(new_n4427_), .ZN(new_n4448_));
  AOI21_X1   g04256(.A1(new_n4448_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n4449_));
  AOI21_X1   g04257(.A1(new_n4449_), .A2(new_n4441_), .B(new_n4447_), .ZN(new_n4450_));
  OAI21_X1   g04258(.A1(new_n4450_), .A2(new_n4442_), .B(\asqrt[52] ), .ZN(new_n4451_));
  INV_X1     g04259(.I(new_n4157_), .ZN(new_n4452_));
  INV_X1     g04260(.I(new_n4151_), .ZN(new_n4453_));
  INV_X1     g04261(.I(new_n4164_), .ZN(new_n4454_));
  NOR2_X1    g04262(.A1(new_n4454_), .A2(new_n4453_), .ZN(new_n4455_));
  NOR3_X1    g04263(.A1(new_n4298_), .A2(new_n4152_), .A3(new_n4455_), .ZN(new_n4456_));
  INV_X1     g04264(.I(new_n4456_), .ZN(new_n4457_));
  NOR3_X1    g04265(.A1(new_n4455_), .A2(new_n4152_), .A3(new_n4452_), .ZN(new_n4458_));
  AOI22_X1   g04266(.A1(new_n4457_), .A2(new_n4452_), .B1(\asqrt[39] ), .B2(new_n4458_), .ZN(new_n4459_));
  INV_X1     g04267(.I(new_n4459_), .ZN(new_n4460_));
  INV_X1     g04268(.I(new_n4431_), .ZN(new_n4461_));
  OR2_X2     g04269(.A1(new_n4419_), .A2(\asqrt[49] ), .Z(new_n4462_));
  OAI21_X1   g04270(.A1(new_n4462_), .A2(new_n4426_), .B(new_n4461_), .ZN(new_n4463_));
  AOI21_X1   g04271(.A1(new_n4463_), .A2(new_n4427_), .B(new_n1612_), .ZN(new_n4464_));
  INV_X1     g04272(.I(new_n4440_), .ZN(new_n4465_));
  AOI21_X1   g04273(.A1(new_n4465_), .A2(new_n4463_), .B(new_n4438_), .ZN(new_n4466_));
  OAI21_X1   g04274(.A1(new_n4466_), .A2(new_n4464_), .B(\asqrt[51] ), .ZN(new_n4467_));
  NAND2_X1   g04275(.A1(new_n4467_), .A2(new_n1256_), .ZN(new_n4468_));
  OAI21_X1   g04276(.A1(new_n4468_), .A2(new_n4450_), .B(new_n4460_), .ZN(new_n4469_));
  AOI21_X1   g04277(.A1(new_n4469_), .A2(new_n4451_), .B(new_n1103_), .ZN(new_n4470_));
  NOR3_X1    g04278(.A1(new_n4167_), .A2(new_n4306_), .A3(new_n4209_), .ZN(new_n4471_));
  NOR3_X1    g04279(.A1(new_n4298_), .A2(new_n4167_), .A3(new_n4209_), .ZN(new_n4472_));
  INV_X1     g04280(.I(new_n4472_), .ZN(new_n4473_));
  AOI22_X1   g04281(.A1(new_n4473_), .A2(new_n4306_), .B1(\asqrt[39] ), .B2(new_n4471_), .ZN(new_n4474_));
  INV_X1     g04282(.I(new_n4447_), .ZN(new_n4475_));
  NAND2_X1   g04283(.A1(new_n4434_), .A2(new_n1376_), .ZN(new_n4476_));
  OAI21_X1   g04284(.A1(new_n4476_), .A2(new_n4466_), .B(new_n4475_), .ZN(new_n4477_));
  AOI21_X1   g04285(.A1(new_n4477_), .A2(new_n4467_), .B(new_n1256_), .ZN(new_n4478_));
  NOR2_X1    g04286(.A1(new_n4478_), .A2(\asqrt[53] ), .ZN(new_n4479_));
  AOI21_X1   g04287(.A1(new_n4479_), .A2(new_n4469_), .B(new_n4474_), .ZN(new_n4480_));
  OAI21_X1   g04288(.A1(new_n4480_), .A2(new_n4470_), .B(\asqrt[54] ), .ZN(new_n4481_));
  INV_X1     g04289(.I(new_n4175_), .ZN(new_n4482_));
  NOR2_X1    g04290(.A1(new_n4182_), .A2(new_n4174_), .ZN(new_n4483_));
  NOR3_X1    g04291(.A1(new_n4298_), .A2(new_n4482_), .A3(new_n4483_), .ZN(new_n4484_));
  INV_X1     g04292(.I(new_n4484_), .ZN(new_n4485_));
  NOR3_X1    g04293(.A1(new_n4482_), .A2(new_n4181_), .A3(new_n4483_), .ZN(new_n4486_));
  AOI22_X1   g04294(.A1(new_n4485_), .A2(new_n4181_), .B1(\asqrt[39] ), .B2(new_n4486_), .ZN(new_n4487_));
  INV_X1     g04295(.I(new_n4487_), .ZN(new_n4488_));
  NOR2_X1    g04296(.A1(new_n4442_), .A2(\asqrt[52] ), .ZN(new_n4489_));
  AOI21_X1   g04297(.A1(new_n4489_), .A2(new_n4477_), .B(new_n4459_), .ZN(new_n4490_));
  OAI21_X1   g04298(.A1(new_n4490_), .A2(new_n4478_), .B(\asqrt[53] ), .ZN(new_n4491_));
  NAND2_X1   g04299(.A1(new_n4491_), .A2(new_n904_), .ZN(new_n4492_));
  OAI21_X1   g04300(.A1(new_n4492_), .A2(new_n4480_), .B(new_n4488_), .ZN(new_n4493_));
  AOI21_X1   g04301(.A1(new_n4493_), .A2(new_n4481_), .B(new_n823_), .ZN(new_n4494_));
  NOR2_X1    g04302(.A1(new_n4193_), .A2(new_n4186_), .ZN(new_n4495_));
  NOR3_X1    g04303(.A1(new_n4495_), .A2(new_n4184_), .A3(new_n4192_), .ZN(new_n4496_));
  NOR3_X1    g04304(.A1(new_n4298_), .A2(new_n4184_), .A3(new_n4495_), .ZN(new_n4497_));
  INV_X1     g04305(.I(new_n4497_), .ZN(new_n4498_));
  AOI22_X1   g04306(.A1(new_n4498_), .A2(new_n4192_), .B1(\asqrt[39] ), .B2(new_n4496_), .ZN(new_n4499_));
  INV_X1     g04307(.I(new_n4474_), .ZN(new_n4500_));
  NAND2_X1   g04308(.A1(new_n4451_), .A2(new_n1103_), .ZN(new_n4501_));
  OAI21_X1   g04309(.A1(new_n4501_), .A2(new_n4490_), .B(new_n4500_), .ZN(new_n4502_));
  AOI21_X1   g04310(.A1(new_n4502_), .A2(new_n4491_), .B(new_n904_), .ZN(new_n4503_));
  NOR2_X1    g04311(.A1(new_n4503_), .A2(\asqrt[55] ), .ZN(new_n4504_));
  AOI21_X1   g04312(.A1(new_n4504_), .A2(new_n4493_), .B(new_n4499_), .ZN(new_n4505_));
  OAI21_X1   g04313(.A1(new_n4505_), .A2(new_n4494_), .B(\asqrt[56] ), .ZN(new_n4506_));
  NOR3_X1    g04314(.A1(new_n4298_), .A2(new_n4195_), .A3(new_n4241_), .ZN(new_n4507_));
  INV_X1     g04315(.I(new_n4507_), .ZN(new_n4508_));
  NOR3_X1    g04316(.A1(new_n4195_), .A2(new_n4305_), .A3(new_n4241_), .ZN(new_n4509_));
  AOI22_X1   g04317(.A1(new_n4508_), .A2(new_n4305_), .B1(\asqrt[39] ), .B2(new_n4509_), .ZN(new_n4510_));
  INV_X1     g04318(.I(new_n4510_), .ZN(new_n4511_));
  NOR3_X1    g04319(.A1(new_n4450_), .A2(new_n4442_), .A3(\asqrt[52] ), .ZN(new_n4512_));
  OAI21_X1   g04320(.A1(new_n4459_), .A2(new_n4512_), .B(new_n4451_), .ZN(new_n4513_));
  AOI21_X1   g04321(.A1(new_n4513_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n4514_));
  AOI21_X1   g04322(.A1(new_n4514_), .A2(new_n4502_), .B(new_n4487_), .ZN(new_n4515_));
  OAI21_X1   g04323(.A1(new_n4515_), .A2(new_n4503_), .B(\asqrt[55] ), .ZN(new_n4516_));
  NAND2_X1   g04324(.A1(new_n4516_), .A2(new_n703_), .ZN(new_n4517_));
  OAI21_X1   g04325(.A1(new_n4517_), .A2(new_n4505_), .B(new_n4511_), .ZN(new_n4518_));
  AOI21_X1   g04326(.A1(new_n4518_), .A2(new_n4506_), .B(new_n531_), .ZN(new_n4519_));
  INV_X1     g04327(.I(new_n4202_), .ZN(new_n4520_));
  NOR2_X1    g04328(.A1(new_n4214_), .A2(new_n4201_), .ZN(new_n4521_));
  NOR3_X1    g04329(.A1(new_n4520_), .A2(new_n4208_), .A3(new_n4521_), .ZN(new_n4522_));
  NOR3_X1    g04330(.A1(new_n4298_), .A2(new_n4520_), .A3(new_n4521_), .ZN(new_n4523_));
  INV_X1     g04331(.I(new_n4523_), .ZN(new_n4524_));
  AOI22_X1   g04332(.A1(new_n4524_), .A2(new_n4208_), .B1(\asqrt[39] ), .B2(new_n4522_), .ZN(new_n4525_));
  NOR3_X1    g04333(.A1(new_n4515_), .A2(\asqrt[55] ), .A3(new_n4503_), .ZN(new_n4526_));
  OAI21_X1   g04334(.A1(new_n4499_), .A2(new_n4526_), .B(new_n4516_), .ZN(new_n4527_));
  AOI21_X1   g04335(.A1(new_n4527_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n4528_));
  AOI21_X1   g04336(.A1(new_n4528_), .A2(new_n4518_), .B(new_n4525_), .ZN(new_n4529_));
  OAI21_X1   g04337(.A1(new_n4529_), .A2(new_n4519_), .B(\asqrt[58] ), .ZN(new_n4530_));
  NOR2_X1    g04338(.A1(new_n4225_), .A2(new_n4218_), .ZN(new_n4531_));
  NOR3_X1    g04339(.A1(new_n4298_), .A2(new_n4216_), .A3(new_n4531_), .ZN(new_n4532_));
  INV_X1     g04340(.I(new_n4532_), .ZN(new_n4533_));
  NOR3_X1    g04341(.A1(new_n4531_), .A2(new_n4216_), .A3(new_n4224_), .ZN(new_n4534_));
  AOI22_X1   g04342(.A1(new_n4533_), .A2(new_n4224_), .B1(\asqrt[39] ), .B2(new_n4534_), .ZN(new_n4535_));
  INV_X1     g04343(.I(new_n4535_), .ZN(new_n4536_));
  INV_X1     g04344(.I(new_n4499_), .ZN(new_n4537_));
  NAND2_X1   g04345(.A1(new_n4481_), .A2(new_n823_), .ZN(new_n4538_));
  OAI21_X1   g04346(.A1(new_n4538_), .A2(new_n4515_), .B(new_n4537_), .ZN(new_n4539_));
  AOI21_X1   g04347(.A1(new_n4539_), .A2(new_n4516_), .B(new_n703_), .ZN(new_n4540_));
  NOR2_X1    g04348(.A1(new_n4494_), .A2(\asqrt[56] ), .ZN(new_n4541_));
  AOI21_X1   g04349(.A1(new_n4541_), .A2(new_n4539_), .B(new_n4510_), .ZN(new_n4542_));
  OAI21_X1   g04350(.A1(new_n4542_), .A2(new_n4540_), .B(\asqrt[57] ), .ZN(new_n4543_));
  NAND2_X1   g04351(.A1(new_n4543_), .A2(new_n436_), .ZN(new_n4544_));
  OAI21_X1   g04352(.A1(new_n4544_), .A2(new_n4529_), .B(new_n4536_), .ZN(new_n4545_));
  AOI21_X1   g04353(.A1(new_n4545_), .A2(new_n4530_), .B(new_n327_), .ZN(new_n4546_));
  NOR3_X1    g04354(.A1(new_n4227_), .A2(new_n4304_), .A3(new_n4272_), .ZN(new_n4547_));
  NOR3_X1    g04355(.A1(new_n4298_), .A2(new_n4227_), .A3(new_n4272_), .ZN(new_n4548_));
  INV_X1     g04356(.I(new_n4548_), .ZN(new_n4549_));
  AOI22_X1   g04357(.A1(new_n4549_), .A2(new_n4304_), .B1(\asqrt[39] ), .B2(new_n4547_), .ZN(new_n4550_));
  INV_X1     g04358(.I(new_n4525_), .ZN(new_n4551_));
  NAND2_X1   g04359(.A1(new_n4506_), .A2(new_n531_), .ZN(new_n4552_));
  OAI21_X1   g04360(.A1(new_n4552_), .A2(new_n4542_), .B(new_n4551_), .ZN(new_n4553_));
  AOI21_X1   g04361(.A1(new_n4553_), .A2(new_n4543_), .B(new_n436_), .ZN(new_n4554_));
  NOR2_X1    g04362(.A1(new_n4554_), .A2(\asqrt[59] ), .ZN(new_n4555_));
  AOI21_X1   g04363(.A1(new_n4555_), .A2(new_n4545_), .B(new_n4550_), .ZN(new_n4556_));
  OAI21_X1   g04364(.A1(new_n4556_), .A2(new_n4546_), .B(\asqrt[60] ), .ZN(new_n4557_));
  INV_X1     g04365(.I(new_n4234_), .ZN(new_n4558_));
  NOR2_X1    g04366(.A1(new_n4246_), .A2(new_n4233_), .ZN(new_n4559_));
  NOR3_X1    g04367(.A1(new_n4298_), .A2(new_n4558_), .A3(new_n4559_), .ZN(new_n4560_));
  INV_X1     g04368(.I(new_n4560_), .ZN(new_n4561_));
  NOR3_X1    g04369(.A1(new_n4558_), .A2(new_n4240_), .A3(new_n4559_), .ZN(new_n4562_));
  AOI22_X1   g04370(.A1(new_n4561_), .A2(new_n4240_), .B1(\asqrt[39] ), .B2(new_n4562_), .ZN(new_n4563_));
  INV_X1     g04371(.I(new_n4563_), .ZN(new_n4564_));
  NOR2_X1    g04372(.A1(new_n4519_), .A2(\asqrt[58] ), .ZN(new_n4565_));
  AOI21_X1   g04373(.A1(new_n4565_), .A2(new_n4553_), .B(new_n4535_), .ZN(new_n4566_));
  OAI21_X1   g04374(.A1(new_n4566_), .A2(new_n4554_), .B(\asqrt[59] ), .ZN(new_n4567_));
  NAND2_X1   g04375(.A1(new_n4567_), .A2(new_n306_), .ZN(new_n4568_));
  OAI21_X1   g04376(.A1(new_n4568_), .A2(new_n4556_), .B(new_n4564_), .ZN(new_n4569_));
  AOI21_X1   g04377(.A1(new_n4569_), .A2(new_n4557_), .B(new_n218_), .ZN(new_n4570_));
  NOR2_X1    g04378(.A1(new_n4250_), .A2(new_n4256_), .ZN(new_n4571_));
  NOR3_X1    g04379(.A1(new_n4571_), .A2(new_n4248_), .A3(new_n4255_), .ZN(new_n4572_));
  NOR3_X1    g04380(.A1(new_n4298_), .A2(new_n4248_), .A3(new_n4571_), .ZN(new_n4573_));
  INV_X1     g04381(.I(new_n4573_), .ZN(new_n4574_));
  AOI22_X1   g04382(.A1(new_n4574_), .A2(new_n4255_), .B1(\asqrt[39] ), .B2(new_n4572_), .ZN(new_n4575_));
  INV_X1     g04383(.I(new_n4550_), .ZN(new_n4576_));
  NAND2_X1   g04384(.A1(new_n4530_), .A2(new_n327_), .ZN(new_n4577_));
  OAI21_X1   g04385(.A1(new_n4577_), .A2(new_n4566_), .B(new_n4576_), .ZN(new_n4578_));
  AOI21_X1   g04386(.A1(new_n4578_), .A2(new_n4567_), .B(new_n306_), .ZN(new_n4579_));
  NOR2_X1    g04387(.A1(new_n4579_), .A2(\asqrt[61] ), .ZN(new_n4580_));
  AOI21_X1   g04388(.A1(new_n4580_), .A2(new_n4569_), .B(new_n4575_), .ZN(new_n4581_));
  OAI21_X1   g04389(.A1(new_n4581_), .A2(new_n4570_), .B(\asqrt[62] ), .ZN(new_n4582_));
  NOR3_X1    g04390(.A1(new_n4298_), .A2(new_n4258_), .A3(new_n4287_), .ZN(new_n4583_));
  INV_X1     g04391(.I(new_n4583_), .ZN(new_n4584_));
  NOR3_X1    g04392(.A1(new_n4258_), .A2(new_n4303_), .A3(new_n4287_), .ZN(new_n4585_));
  AOI22_X1   g04393(.A1(new_n4584_), .A2(new_n4303_), .B1(\asqrt[39] ), .B2(new_n4585_), .ZN(new_n4586_));
  INV_X1     g04394(.I(new_n4586_), .ZN(new_n4587_));
  NOR3_X1    g04395(.A1(new_n4529_), .A2(\asqrt[58] ), .A3(new_n4519_), .ZN(new_n4588_));
  OAI21_X1   g04396(.A1(new_n4535_), .A2(new_n4588_), .B(new_n4530_), .ZN(new_n4589_));
  AOI21_X1   g04397(.A1(new_n4589_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n4590_));
  AOI21_X1   g04398(.A1(new_n4590_), .A2(new_n4578_), .B(new_n4563_), .ZN(new_n4591_));
  OAI21_X1   g04399(.A1(new_n4591_), .A2(new_n4579_), .B(\asqrt[61] ), .ZN(new_n4592_));
  NAND2_X1   g04400(.A1(new_n4592_), .A2(new_n207_), .ZN(new_n4593_));
  OAI21_X1   g04401(.A1(new_n4593_), .A2(new_n4581_), .B(new_n4587_), .ZN(new_n4594_));
  INV_X1     g04402(.I(new_n4355_), .ZN(new_n4595_));
  NAND4_X1   g04403(.A1(\asqrt[39] ), .A2(new_n4265_), .A3(new_n4270_), .A4(new_n4334_), .ZN(new_n4596_));
  NAND2_X1   g04404(.A1(new_n4265_), .A2(new_n4334_), .ZN(new_n4597_));
  OAI21_X1   g04405(.A1(new_n4298_), .A2(new_n4597_), .B(new_n4271_), .ZN(new_n4598_));
  NAND2_X1   g04406(.A1(new_n4598_), .A2(new_n4596_), .ZN(new_n4599_));
  NOR2_X1    g04407(.A1(new_n4335_), .A2(new_n4350_), .ZN(new_n4600_));
  NAND2_X1   g04408(.A1(\asqrt[39] ), .A2(new_n4600_), .ZN(new_n4601_));
  NAND3_X1   g04409(.A1(new_n4599_), .A2(new_n4595_), .A3(new_n4601_), .ZN(new_n4602_));
  AOI21_X1   g04410(.A1(new_n4594_), .A2(new_n4582_), .B(new_n4602_), .ZN(new_n4603_));
  NOR3_X1    g04411(.A1(new_n4591_), .A2(\asqrt[61] ), .A3(new_n4579_), .ZN(new_n4604_));
  OAI21_X1   g04412(.A1(new_n4575_), .A2(new_n4604_), .B(new_n4592_), .ZN(new_n4605_));
  AOI21_X1   g04413(.A1(new_n4605_), .A2(\asqrt[62] ), .B(new_n4599_), .ZN(new_n4606_));
  OAI21_X1   g04414(.A1(new_n4298_), .A2(new_n4350_), .B(new_n4335_), .ZN(new_n4607_));
  NOR2_X1    g04415(.A1(new_n4600_), .A2(new_n193_), .ZN(new_n4608_));
  NAND2_X1   g04416(.A1(new_n4607_), .A2(new_n4608_), .ZN(new_n4609_));
  INV_X1     g04417(.I(new_n4609_), .ZN(new_n4610_));
  AND3_X2    g04418(.A1(new_n4281_), .A2(new_n4279_), .A3(new_n4294_), .Z(new_n4611_));
  NAND4_X1   g04419(.A1(new_n4595_), .A2(new_n4336_), .A3(new_n4291_), .A4(new_n4611_), .ZN(new_n4612_));
  INV_X1     g04420(.I(new_n4612_), .ZN(new_n4613_));
  NOR2_X1    g04421(.A1(new_n4610_), .A2(new_n4613_), .ZN(new_n4614_));
  INV_X1     g04422(.I(new_n4614_), .ZN(new_n4615_));
  AOI21_X1   g04423(.A1(new_n4606_), .A2(new_n4594_), .B(new_n4615_), .ZN(new_n4616_));
  OAI21_X1   g04424(.A1(\asqrt[63] ), .A2(new_n4603_), .B(new_n4616_), .ZN(\asqrt[38] ));
  NOR2_X1    g04425(.A1(\a[74] ), .A2(\a[75] ), .ZN(new_n4618_));
  INV_X1     g04426(.I(new_n4618_), .ZN(new_n4619_));
  NOR2_X1    g04427(.A1(new_n4619_), .A2(\a[76] ), .ZN(new_n4620_));
  INV_X1     g04428(.I(new_n4620_), .ZN(new_n4621_));
  NAND2_X1   g04429(.A1(new_n4594_), .A2(new_n4582_), .ZN(new_n4622_));
  INV_X1     g04430(.I(new_n4602_), .ZN(new_n4623_));
  AOI21_X1   g04431(.A1(new_n4622_), .A2(new_n4623_), .B(\asqrt[63] ), .ZN(new_n4624_));
  INV_X1     g04432(.I(new_n4594_), .ZN(new_n4625_));
  INV_X1     g04433(.I(new_n4599_), .ZN(new_n4626_));
  NAND2_X1   g04434(.A1(new_n4582_), .A2(new_n4626_), .ZN(new_n4627_));
  OAI21_X1   g04435(.A1(new_n4625_), .A2(new_n4627_), .B(new_n4614_), .ZN(new_n4628_));
  OAI21_X1   g04436(.A1(new_n4624_), .A2(new_n4628_), .B(\a[76] ), .ZN(new_n4629_));
  AOI21_X1   g04437(.A1(new_n4629_), .A2(new_n4621_), .B(new_n4298_), .ZN(new_n4630_));
  INV_X1     g04438(.I(\a[76] ), .ZN(new_n4631_));
  INV_X1     g04439(.I(new_n4575_), .ZN(new_n4632_));
  NAND2_X1   g04440(.A1(new_n4557_), .A2(new_n218_), .ZN(new_n4633_));
  OAI21_X1   g04441(.A1(new_n4633_), .A2(new_n4591_), .B(new_n4632_), .ZN(new_n4634_));
  NAND3_X1   g04442(.A1(new_n4634_), .A2(new_n207_), .A3(new_n4592_), .ZN(new_n4635_));
  AOI22_X1   g04443(.A1(new_n4635_), .A2(new_n4587_), .B1(new_n4605_), .B2(\asqrt[62] ), .ZN(new_n4636_));
  OAI21_X1   g04444(.A1(new_n4636_), .A2(new_n4602_), .B(new_n193_), .ZN(new_n4637_));
  AOI21_X1   g04445(.A1(new_n4637_), .A2(new_n4616_), .B(new_n4631_), .ZN(new_n4638_));
  NAND4_X1   g04446(.A1(new_n4595_), .A2(new_n4291_), .A3(new_n4294_), .A4(new_n4621_), .ZN(new_n4639_));
  NOR2_X1    g04447(.A1(new_n4639_), .A2(new_n4348_), .ZN(new_n4640_));
  INV_X1     g04448(.I(new_n4640_), .ZN(new_n4641_));
  NOR2_X1    g04449(.A1(new_n4638_), .A2(new_n4641_), .ZN(new_n4642_));
  AOI21_X1   g04450(.A1(new_n4637_), .A2(new_n4616_), .B(new_n4300_), .ZN(new_n4643_));
  INV_X1     g04451(.I(\a[77] ), .ZN(new_n4644_));
  AOI21_X1   g04452(.A1(\asqrt[38] ), .A2(new_n4631_), .B(new_n4644_), .ZN(new_n4645_));
  NOR3_X1    g04453(.A1(new_n4642_), .A2(new_n4645_), .A3(new_n4643_), .ZN(new_n4646_));
  OAI21_X1   g04454(.A1(new_n4646_), .A2(new_n4630_), .B(\asqrt[40] ), .ZN(new_n4647_));
  OAI21_X1   g04455(.A1(new_n4624_), .A2(new_n4628_), .B(new_n4299_), .ZN(new_n4648_));
  NOR2_X1    g04456(.A1(new_n4625_), .A2(new_n4627_), .ZN(new_n4649_));
  INV_X1     g04457(.I(new_n4649_), .ZN(new_n4650_));
  NOR2_X1    g04458(.A1(new_n4613_), .A2(new_n4298_), .ZN(new_n4651_));
  NAND4_X1   g04459(.A1(new_n4650_), .A2(new_n4637_), .A3(new_n4609_), .A4(new_n4651_), .ZN(new_n4652_));
  AOI21_X1   g04460(.A1(new_n4652_), .A2(new_n4648_), .B(new_n4302_), .ZN(new_n4653_));
  INV_X1     g04461(.I(new_n4651_), .ZN(new_n4654_));
  NOR4_X1    g04462(.A1(new_n4624_), .A2(new_n4649_), .A3(new_n4610_), .A4(new_n4654_), .ZN(new_n4655_));
  NOR3_X1    g04463(.A1(new_n4655_), .A2(new_n4643_), .A3(\a[78] ), .ZN(new_n4656_));
  AOI21_X1   g04464(.A1(\asqrt[38] ), .A2(\a[76] ), .B(new_n4620_), .ZN(new_n4657_));
  OAI21_X1   g04465(.A1(new_n4657_), .A2(new_n4298_), .B(new_n4071_), .ZN(new_n4658_));
  OAI22_X1   g04466(.A1(new_n4646_), .A2(new_n4658_), .B1(new_n4653_), .B2(new_n4656_), .ZN(new_n4659_));
  AOI21_X1   g04467(.A1(new_n4659_), .A2(new_n4647_), .B(new_n3782_), .ZN(new_n4660_));
  INV_X1     g04468(.I(new_n4370_), .ZN(new_n4661_));
  NOR3_X1    g04469(.A1(new_n4339_), .A2(new_n4661_), .A3(new_n4342_), .ZN(new_n4662_));
  NOR2_X1    g04470(.A1(new_n4339_), .A2(new_n4342_), .ZN(new_n4663_));
  NAND2_X1   g04471(.A1(\asqrt[38] ), .A2(new_n4663_), .ZN(new_n4664_));
  AOI22_X1   g04472(.A1(new_n4664_), .A2(new_n4661_), .B1(\asqrt[38] ), .B2(new_n4662_), .ZN(new_n4665_));
  OAI21_X1   g04473(.A1(new_n4638_), .A2(new_n4620_), .B(\asqrt[39] ), .ZN(new_n4666_));
  AOI21_X1   g04474(.A1(new_n4637_), .A2(new_n4616_), .B(\a[76] ), .ZN(new_n4667_));
  OAI21_X1   g04475(.A1(new_n4644_), .A2(new_n4667_), .B(new_n4648_), .ZN(new_n4668_));
  OAI21_X1   g04476(.A1(new_n4668_), .A2(new_n4642_), .B(new_n4666_), .ZN(new_n4669_));
  AOI21_X1   g04477(.A1(new_n4669_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n4670_));
  AOI21_X1   g04478(.A1(new_n4670_), .A2(new_n4659_), .B(new_n4665_), .ZN(new_n4671_));
  OAI21_X1   g04479(.A1(new_n4671_), .A2(new_n4660_), .B(\asqrt[42] ), .ZN(new_n4672_));
  INV_X1     g04480(.I(new_n4672_), .ZN(new_n4673_));
  NOR2_X1    g04481(.A1(new_n4360_), .A2(new_n4361_), .ZN(new_n4674_));
  NOR2_X1    g04482(.A1(new_n4346_), .A2(new_n4363_), .ZN(new_n4675_));
  INV_X1     g04483(.I(new_n4675_), .ZN(new_n4676_));
  NAND4_X1   g04484(.A1(\asqrt[38] ), .A2(new_n4347_), .A3(new_n4674_), .A4(new_n4676_), .ZN(new_n4677_));
  AND3_X2    g04485(.A1(\asqrt[38] ), .A2(new_n4347_), .A3(new_n4676_), .Z(new_n4678_));
  OAI21_X1   g04486(.A1(new_n4678_), .A2(new_n4674_), .B(new_n4677_), .ZN(new_n4679_));
  INV_X1     g04487(.I(new_n4679_), .ZN(new_n4680_));
  NOR3_X1    g04488(.A1(new_n4671_), .A2(new_n4660_), .A3(\asqrt[42] ), .ZN(new_n4681_));
  NOR2_X1    g04489(.A1(new_n4681_), .A2(new_n4680_), .ZN(new_n4682_));
  OAI21_X1   g04490(.A1(new_n4682_), .A2(new_n4673_), .B(\asqrt[43] ), .ZN(new_n4683_));
  INV_X1     g04491(.I(new_n4368_), .ZN(new_n4684_));
  INV_X1     g04492(.I(new_n4365_), .ZN(new_n4685_));
  NAND2_X1   g04493(.A1(new_n4372_), .A2(new_n4364_), .ZN(new_n4686_));
  NAND3_X1   g04494(.A1(\asqrt[38] ), .A2(new_n4685_), .A3(new_n4686_), .ZN(new_n4687_));
  AND3_X2    g04495(.A1(new_n4685_), .A2(new_n4368_), .A3(new_n4686_), .Z(new_n4688_));
  AOI22_X1   g04496(.A1(new_n4687_), .A2(new_n4684_), .B1(\asqrt[38] ), .B2(new_n4688_), .ZN(new_n4689_));
  INV_X1     g04497(.I(new_n4689_), .ZN(new_n4690_));
  NAND2_X1   g04498(.A1(new_n4672_), .A2(new_n3218_), .ZN(new_n4691_));
  OAI21_X1   g04499(.A1(new_n4682_), .A2(new_n4691_), .B(new_n4690_), .ZN(new_n4692_));
  AOI21_X1   g04500(.A1(new_n4692_), .A2(new_n4683_), .B(new_n2954_), .ZN(new_n4693_));
  INV_X1     g04501(.I(new_n4382_), .ZN(new_n4694_));
  NOR3_X1    g04502(.A1(new_n4375_), .A2(new_n4383_), .A3(new_n4694_), .ZN(new_n4695_));
  INV_X1     g04503(.I(\asqrt[38] ), .ZN(new_n4696_));
  NOR3_X1    g04504(.A1(new_n4696_), .A2(new_n4375_), .A3(new_n4383_), .ZN(new_n4697_));
  INV_X1     g04505(.I(new_n4697_), .ZN(new_n4698_));
  AOI22_X1   g04506(.A1(new_n4698_), .A2(new_n4694_), .B1(\asqrt[38] ), .B2(new_n4695_), .ZN(new_n4699_));
  OAI21_X1   g04507(.A1(new_n4680_), .A2(new_n4681_), .B(new_n4672_), .ZN(new_n4700_));
  AOI21_X1   g04508(.A1(new_n4700_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n4701_));
  AOI21_X1   g04509(.A1(new_n4701_), .A2(new_n4692_), .B(new_n4699_), .ZN(new_n4702_));
  OAI21_X1   g04510(.A1(new_n4702_), .A2(new_n4693_), .B(\asqrt[45] ), .ZN(new_n4703_));
  INV_X1     g04511(.I(new_n4703_), .ZN(new_n4704_));
  INV_X1     g04512(.I(new_n4384_), .ZN(new_n4705_));
  INV_X1     g04513(.I(new_n4392_), .ZN(new_n4706_));
  NAND2_X1   g04514(.A1(new_n4705_), .A2(new_n4706_), .ZN(new_n4707_));
  NAND3_X1   g04515(.A1(\asqrt[38] ), .A2(new_n4385_), .A3(new_n4707_), .ZN(new_n4708_));
  AND3_X2    g04516(.A1(new_n4707_), .A2(new_n4385_), .A3(new_n4390_), .Z(new_n4709_));
  AOI22_X1   g04517(.A1(new_n4708_), .A2(new_n4391_), .B1(\asqrt[38] ), .B2(new_n4709_), .ZN(new_n4710_));
  NOR3_X1    g04518(.A1(new_n4702_), .A2(new_n4693_), .A3(\asqrt[45] ), .ZN(new_n4711_));
  NOR2_X1    g04519(.A1(new_n4711_), .A2(new_n4710_), .ZN(new_n4712_));
  OAI21_X1   g04520(.A1(new_n4712_), .A2(new_n4704_), .B(\asqrt[46] ), .ZN(new_n4713_));
  INV_X1     g04521(.I(new_n4398_), .ZN(new_n4714_));
  INV_X1     g04522(.I(new_n4393_), .ZN(new_n4715_));
  INV_X1     g04523(.I(new_n4400_), .ZN(new_n4716_));
  NOR2_X1    g04524(.A1(new_n4716_), .A2(new_n4715_), .ZN(new_n4717_));
  NOR3_X1    g04525(.A1(new_n4717_), .A2(new_n4394_), .A3(new_n4714_), .ZN(new_n4718_));
  NOR3_X1    g04526(.A1(new_n4696_), .A2(new_n4394_), .A3(new_n4717_), .ZN(new_n4719_));
  INV_X1     g04527(.I(new_n4719_), .ZN(new_n4720_));
  AOI22_X1   g04528(.A1(new_n4720_), .A2(new_n4714_), .B1(\asqrt[38] ), .B2(new_n4718_), .ZN(new_n4721_));
  INV_X1     g04529(.I(new_n4721_), .ZN(new_n4722_));
  NAND2_X1   g04530(.A1(new_n4703_), .A2(new_n2465_), .ZN(new_n4723_));
  OAI21_X1   g04531(.A1(new_n4712_), .A2(new_n4723_), .B(new_n4722_), .ZN(new_n4724_));
  AOI21_X1   g04532(.A1(new_n4724_), .A2(new_n4713_), .B(new_n2229_), .ZN(new_n4725_));
  INV_X1     g04533(.I(new_n4408_), .ZN(new_n4726_));
  NOR3_X1    g04534(.A1(new_n4696_), .A2(new_n4403_), .A3(new_n4409_), .ZN(new_n4727_));
  INV_X1     g04535(.I(new_n4727_), .ZN(new_n4728_));
  NOR3_X1    g04536(.A1(new_n4403_), .A2(new_n4726_), .A3(new_n4409_), .ZN(new_n4729_));
  AOI22_X1   g04537(.A1(new_n4728_), .A2(new_n4726_), .B1(\asqrt[38] ), .B2(new_n4729_), .ZN(new_n4730_));
  OAI21_X1   g04538(.A1(new_n4710_), .A2(new_n4711_), .B(new_n4703_), .ZN(new_n4731_));
  AOI21_X1   g04539(.A1(new_n4731_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n4732_));
  AOI21_X1   g04540(.A1(new_n4732_), .A2(new_n4724_), .B(new_n4730_), .ZN(new_n4733_));
  OAI21_X1   g04541(.A1(new_n4733_), .A2(new_n4725_), .B(\asqrt[48] ), .ZN(new_n4734_));
  INV_X1     g04542(.I(new_n4734_), .ZN(new_n4735_));
  NOR2_X1    g04543(.A1(new_n4410_), .A2(new_n4417_), .ZN(new_n4736_));
  INV_X1     g04544(.I(new_n4736_), .ZN(new_n4737_));
  AND3_X2    g04545(.A1(new_n4737_), .A2(new_n4411_), .A3(new_n4415_), .Z(new_n4738_));
  NAND3_X1   g04546(.A1(\asqrt[38] ), .A2(new_n4411_), .A3(new_n4737_), .ZN(new_n4739_));
  AOI22_X1   g04547(.A1(new_n4739_), .A2(new_n4416_), .B1(\asqrt[38] ), .B2(new_n4738_), .ZN(new_n4740_));
  NOR3_X1    g04548(.A1(new_n4733_), .A2(new_n4725_), .A3(\asqrt[48] ), .ZN(new_n4741_));
  NOR2_X1    g04549(.A1(new_n4741_), .A2(new_n4740_), .ZN(new_n4742_));
  OAI21_X1   g04550(.A1(new_n4742_), .A2(new_n4735_), .B(\asqrt[49] ), .ZN(new_n4743_));
  INV_X1     g04551(.I(new_n4423_), .ZN(new_n4744_));
  INV_X1     g04552(.I(new_n4418_), .ZN(new_n4745_));
  NAND2_X1   g04553(.A1(new_n4411_), .A2(new_n1956_), .ZN(new_n4746_));
  NOR2_X1    g04554(.A1(new_n4746_), .A2(new_n4745_), .ZN(new_n4747_));
  NOR3_X1    g04555(.A1(new_n4696_), .A2(new_n4419_), .A3(new_n4747_), .ZN(new_n4748_));
  INV_X1     g04556(.I(new_n4748_), .ZN(new_n4749_));
  NOR3_X1    g04557(.A1(new_n4747_), .A2(new_n4419_), .A3(new_n4744_), .ZN(new_n4750_));
  AOI22_X1   g04558(.A1(new_n4749_), .A2(new_n4744_), .B1(\asqrt[38] ), .B2(new_n4750_), .ZN(new_n4751_));
  INV_X1     g04559(.I(new_n4751_), .ZN(new_n4752_));
  NAND2_X1   g04560(.A1(new_n4734_), .A2(new_n1806_), .ZN(new_n4753_));
  OAI21_X1   g04561(.A1(new_n4742_), .A2(new_n4753_), .B(new_n4752_), .ZN(new_n4754_));
  AOI21_X1   g04562(.A1(new_n4754_), .A2(new_n4743_), .B(new_n1612_), .ZN(new_n4755_));
  NOR3_X1    g04563(.A1(new_n4428_), .A2(new_n4432_), .A3(new_n4461_), .ZN(new_n4756_));
  NOR3_X1    g04564(.A1(new_n4696_), .A2(new_n4428_), .A3(new_n4432_), .ZN(new_n4757_));
  INV_X1     g04565(.I(new_n4757_), .ZN(new_n4758_));
  AOI22_X1   g04566(.A1(new_n4758_), .A2(new_n4461_), .B1(\asqrt[38] ), .B2(new_n4756_), .ZN(new_n4759_));
  OAI21_X1   g04567(.A1(new_n4740_), .A2(new_n4741_), .B(new_n4734_), .ZN(new_n4760_));
  AOI21_X1   g04568(.A1(new_n4760_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n4761_));
  AOI21_X1   g04569(.A1(new_n4761_), .A2(new_n4754_), .B(new_n4759_), .ZN(new_n4762_));
  OAI21_X1   g04570(.A1(new_n4762_), .A2(new_n4755_), .B(\asqrt[51] ), .ZN(new_n4763_));
  INV_X1     g04571(.I(new_n4763_), .ZN(new_n4764_));
  NOR2_X1    g04572(.A1(new_n4433_), .A2(new_n4440_), .ZN(new_n4765_));
  NOR3_X1    g04573(.A1(new_n4696_), .A2(new_n4464_), .A3(new_n4765_), .ZN(new_n4766_));
  INV_X1     g04574(.I(new_n4766_), .ZN(new_n4767_));
  NOR3_X1    g04575(.A1(new_n4464_), .A2(new_n4439_), .A3(new_n4765_), .ZN(new_n4768_));
  AOI22_X1   g04576(.A1(new_n4767_), .A2(new_n4439_), .B1(\asqrt[38] ), .B2(new_n4768_), .ZN(new_n4769_));
  NOR3_X1    g04577(.A1(new_n4762_), .A2(new_n4755_), .A3(\asqrt[51] ), .ZN(new_n4770_));
  NOR2_X1    g04578(.A1(new_n4770_), .A2(new_n4769_), .ZN(new_n4771_));
  OAI21_X1   g04579(.A1(new_n4771_), .A2(new_n4764_), .B(\asqrt[52] ), .ZN(new_n4772_));
  NOR2_X1    g04580(.A1(new_n4476_), .A2(new_n4466_), .ZN(new_n4773_));
  NOR3_X1    g04581(.A1(new_n4773_), .A2(new_n4442_), .A3(new_n4475_), .ZN(new_n4774_));
  NOR3_X1    g04582(.A1(new_n4696_), .A2(new_n4442_), .A3(new_n4773_), .ZN(new_n4775_));
  INV_X1     g04583(.I(new_n4775_), .ZN(new_n4776_));
  AOI22_X1   g04584(.A1(new_n4776_), .A2(new_n4475_), .B1(\asqrt[38] ), .B2(new_n4774_), .ZN(new_n4777_));
  INV_X1     g04585(.I(new_n4777_), .ZN(new_n4778_));
  NAND2_X1   g04586(.A1(new_n4763_), .A2(new_n1256_), .ZN(new_n4779_));
  OAI21_X1   g04587(.A1(new_n4771_), .A2(new_n4779_), .B(new_n4778_), .ZN(new_n4780_));
  AOI21_X1   g04588(.A1(new_n4780_), .A2(new_n4772_), .B(new_n1103_), .ZN(new_n4781_));
  NOR3_X1    g04589(.A1(new_n4696_), .A2(new_n4478_), .A3(new_n4512_), .ZN(new_n4782_));
  INV_X1     g04590(.I(new_n4782_), .ZN(new_n4783_));
  NOR3_X1    g04591(.A1(new_n4478_), .A2(new_n4512_), .A3(new_n4460_), .ZN(new_n4784_));
  AOI22_X1   g04592(.A1(new_n4783_), .A2(new_n4460_), .B1(\asqrt[38] ), .B2(new_n4784_), .ZN(new_n4785_));
  OAI21_X1   g04593(.A1(new_n4769_), .A2(new_n4770_), .B(new_n4763_), .ZN(new_n4786_));
  AOI21_X1   g04594(.A1(new_n4786_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n4787_));
  AOI21_X1   g04595(.A1(new_n4787_), .A2(new_n4780_), .B(new_n4785_), .ZN(new_n4788_));
  OAI21_X1   g04596(.A1(new_n4788_), .A2(new_n4781_), .B(\asqrt[54] ), .ZN(new_n4789_));
  INV_X1     g04597(.I(new_n4789_), .ZN(new_n4790_));
  NOR2_X1    g04598(.A1(new_n4501_), .A2(new_n4490_), .ZN(new_n4791_));
  NOR3_X1    g04599(.A1(new_n4470_), .A2(new_n4791_), .A3(new_n4500_), .ZN(new_n4792_));
  NOR3_X1    g04600(.A1(new_n4696_), .A2(new_n4470_), .A3(new_n4791_), .ZN(new_n4793_));
  INV_X1     g04601(.I(new_n4793_), .ZN(new_n4794_));
  AOI22_X1   g04602(.A1(new_n4794_), .A2(new_n4500_), .B1(\asqrt[38] ), .B2(new_n4792_), .ZN(new_n4795_));
  NOR3_X1    g04603(.A1(new_n4788_), .A2(new_n4781_), .A3(\asqrt[54] ), .ZN(new_n4796_));
  NOR2_X1    g04604(.A1(new_n4796_), .A2(new_n4795_), .ZN(new_n4797_));
  OAI21_X1   g04605(.A1(new_n4797_), .A2(new_n4790_), .B(\asqrt[55] ), .ZN(new_n4798_));
  NOR2_X1    g04606(.A1(new_n4492_), .A2(new_n4480_), .ZN(new_n4799_));
  NOR3_X1    g04607(.A1(new_n4696_), .A2(new_n4503_), .A3(new_n4799_), .ZN(new_n4800_));
  INV_X1     g04608(.I(new_n4800_), .ZN(new_n4801_));
  NOR3_X1    g04609(.A1(new_n4799_), .A2(new_n4503_), .A3(new_n4488_), .ZN(new_n4802_));
  AOI22_X1   g04610(.A1(new_n4801_), .A2(new_n4488_), .B1(\asqrt[38] ), .B2(new_n4802_), .ZN(new_n4803_));
  INV_X1     g04611(.I(new_n4803_), .ZN(new_n4804_));
  NAND2_X1   g04612(.A1(new_n4789_), .A2(new_n823_), .ZN(new_n4805_));
  OAI21_X1   g04613(.A1(new_n4797_), .A2(new_n4805_), .B(new_n4804_), .ZN(new_n4806_));
  AOI21_X1   g04614(.A1(new_n4806_), .A2(new_n4798_), .B(new_n703_), .ZN(new_n4807_));
  NOR3_X1    g04615(.A1(new_n4494_), .A2(new_n4526_), .A3(new_n4537_), .ZN(new_n4808_));
  NOR3_X1    g04616(.A1(new_n4696_), .A2(new_n4494_), .A3(new_n4526_), .ZN(new_n4809_));
  INV_X1     g04617(.I(new_n4809_), .ZN(new_n4810_));
  AOI22_X1   g04618(.A1(new_n4810_), .A2(new_n4537_), .B1(\asqrt[38] ), .B2(new_n4808_), .ZN(new_n4811_));
  OAI21_X1   g04619(.A1(new_n4795_), .A2(new_n4796_), .B(new_n4789_), .ZN(new_n4812_));
  AOI21_X1   g04620(.A1(new_n4812_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n4813_));
  AOI21_X1   g04621(.A1(new_n4813_), .A2(new_n4806_), .B(new_n4811_), .ZN(new_n4814_));
  OAI21_X1   g04622(.A1(new_n4814_), .A2(new_n4807_), .B(\asqrt[57] ), .ZN(new_n4815_));
  NOR2_X1    g04623(.A1(new_n4517_), .A2(new_n4505_), .ZN(new_n4816_));
  NOR3_X1    g04624(.A1(new_n4696_), .A2(new_n4540_), .A3(new_n4816_), .ZN(new_n4817_));
  INV_X1     g04625(.I(new_n4817_), .ZN(new_n4818_));
  NOR3_X1    g04626(.A1(new_n4540_), .A2(new_n4816_), .A3(new_n4511_), .ZN(new_n4819_));
  AOI22_X1   g04627(.A1(new_n4818_), .A2(new_n4511_), .B1(\asqrt[38] ), .B2(new_n4819_), .ZN(new_n4820_));
  INV_X1     g04628(.I(new_n4820_), .ZN(new_n4821_));
  INV_X1     g04629(.I(new_n4795_), .ZN(new_n4822_));
  INV_X1     g04630(.I(new_n4769_), .ZN(new_n4823_));
  INV_X1     g04631(.I(new_n4740_), .ZN(new_n4824_));
  INV_X1     g04632(.I(new_n4710_), .ZN(new_n4825_));
  NAND2_X1   g04633(.A1(new_n4629_), .A2(new_n4640_), .ZN(new_n4826_));
  OAI21_X1   g04634(.A1(new_n4624_), .A2(new_n4628_), .B(new_n4631_), .ZN(new_n4827_));
  NAND2_X1   g04635(.A1(new_n4827_), .A2(\a[77] ), .ZN(new_n4828_));
  NAND3_X1   g04636(.A1(new_n4826_), .A2(new_n4828_), .A3(new_n4648_), .ZN(new_n4829_));
  AOI21_X1   g04637(.A1(new_n4829_), .A2(new_n4666_), .B(new_n4071_), .ZN(new_n4830_));
  OAI21_X1   g04638(.A1(new_n4655_), .A2(new_n4643_), .B(\a[78] ), .ZN(new_n4831_));
  NAND3_X1   g04639(.A1(new_n4652_), .A2(new_n4648_), .A3(new_n4302_), .ZN(new_n4832_));
  NAND2_X1   g04640(.A1(new_n4629_), .A2(new_n4621_), .ZN(new_n4833_));
  AOI21_X1   g04641(.A1(new_n4833_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n4834_));
  AOI22_X1   g04642(.A1(new_n4829_), .A2(new_n4834_), .B1(new_n4831_), .B2(new_n4832_), .ZN(new_n4835_));
  OAI21_X1   g04643(.A1(new_n4835_), .A2(new_n4830_), .B(\asqrt[41] ), .ZN(new_n4836_));
  NAND2_X1   g04644(.A1(new_n4836_), .A2(new_n3419_), .ZN(new_n4837_));
  OAI21_X1   g04645(.A1(new_n4837_), .A2(new_n4671_), .B(new_n4679_), .ZN(new_n4838_));
  AOI21_X1   g04646(.A1(new_n4838_), .A2(new_n4672_), .B(new_n3218_), .ZN(new_n4839_));
  INV_X1     g04647(.I(new_n4665_), .ZN(new_n4840_));
  AOI21_X1   g04648(.A1(\a[77] ), .A2(new_n4827_), .B(new_n4643_), .ZN(new_n4841_));
  AOI21_X1   g04649(.A1(new_n4841_), .A2(new_n4826_), .B(new_n4630_), .ZN(new_n4842_));
  OAI21_X1   g04650(.A1(new_n4842_), .A2(new_n4071_), .B(new_n3782_), .ZN(new_n4843_));
  OAI21_X1   g04651(.A1(new_n4843_), .A2(new_n4835_), .B(new_n4840_), .ZN(new_n4844_));
  NAND2_X1   g04652(.A1(new_n4844_), .A2(new_n4836_), .ZN(new_n4845_));
  AOI21_X1   g04653(.A1(new_n4845_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n4846_));
  AOI21_X1   g04654(.A1(new_n4846_), .A2(new_n4838_), .B(new_n4689_), .ZN(new_n4847_));
  OAI21_X1   g04655(.A1(new_n4847_), .A2(new_n4839_), .B(\asqrt[44] ), .ZN(new_n4848_));
  NAND2_X1   g04656(.A1(new_n4848_), .A2(new_n2641_), .ZN(new_n4849_));
  OAI21_X1   g04657(.A1(new_n4849_), .A2(new_n4702_), .B(new_n4825_), .ZN(new_n4850_));
  NAND3_X1   g04658(.A1(new_n4850_), .A2(new_n2465_), .A3(new_n4703_), .ZN(new_n4851_));
  AOI22_X1   g04659(.A1(new_n4851_), .A2(new_n4722_), .B1(new_n4731_), .B2(\asqrt[46] ), .ZN(new_n4852_));
  OAI21_X1   g04660(.A1(new_n4852_), .A2(new_n2229_), .B(new_n1956_), .ZN(new_n4853_));
  OAI21_X1   g04661(.A1(new_n4853_), .A2(new_n4733_), .B(new_n4824_), .ZN(new_n4854_));
  AOI21_X1   g04662(.A1(new_n4854_), .A2(new_n4734_), .B(new_n1806_), .ZN(new_n4855_));
  AOI21_X1   g04663(.A1(new_n4850_), .A2(new_n4703_), .B(new_n2465_), .ZN(new_n4856_));
  NOR3_X1    g04664(.A1(new_n4847_), .A2(new_n4839_), .A3(\asqrt[44] ), .ZN(new_n4857_));
  OAI21_X1   g04665(.A1(new_n4699_), .A2(new_n4857_), .B(new_n4848_), .ZN(new_n4858_));
  AOI21_X1   g04666(.A1(new_n4858_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n4859_));
  AOI21_X1   g04667(.A1(new_n4859_), .A2(new_n4850_), .B(new_n4721_), .ZN(new_n4860_));
  NOR3_X1    g04668(.A1(new_n4860_), .A2(\asqrt[47] ), .A3(new_n4856_), .ZN(new_n4861_));
  OAI22_X1   g04669(.A1(new_n4861_), .A2(new_n4730_), .B1(new_n4852_), .B2(new_n2229_), .ZN(new_n4862_));
  AOI21_X1   g04670(.A1(new_n4862_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n4863_));
  AOI21_X1   g04671(.A1(new_n4863_), .A2(new_n4854_), .B(new_n4751_), .ZN(new_n4864_));
  OAI21_X1   g04672(.A1(new_n4864_), .A2(new_n4855_), .B(\asqrt[50] ), .ZN(new_n4865_));
  NAND2_X1   g04673(.A1(new_n4865_), .A2(new_n1376_), .ZN(new_n4866_));
  OAI21_X1   g04674(.A1(new_n4866_), .A2(new_n4762_), .B(new_n4823_), .ZN(new_n4867_));
  AOI21_X1   g04675(.A1(new_n4867_), .A2(new_n4763_), .B(new_n1256_), .ZN(new_n4868_));
  NOR3_X1    g04676(.A1(new_n4864_), .A2(\asqrt[50] ), .A3(new_n4855_), .ZN(new_n4869_));
  OAI21_X1   g04677(.A1(new_n4759_), .A2(new_n4869_), .B(new_n4865_), .ZN(new_n4870_));
  AOI21_X1   g04678(.A1(new_n4870_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n4871_));
  AOI21_X1   g04679(.A1(new_n4871_), .A2(new_n4867_), .B(new_n4777_), .ZN(new_n4872_));
  OAI21_X1   g04680(.A1(new_n4872_), .A2(new_n4868_), .B(\asqrt[53] ), .ZN(new_n4873_));
  NAND2_X1   g04681(.A1(new_n4873_), .A2(new_n904_), .ZN(new_n4874_));
  OAI21_X1   g04682(.A1(new_n4874_), .A2(new_n4788_), .B(new_n4822_), .ZN(new_n4875_));
  AOI21_X1   g04683(.A1(new_n4875_), .A2(new_n4789_), .B(new_n823_), .ZN(new_n4876_));
  NOR3_X1    g04684(.A1(new_n4872_), .A2(\asqrt[53] ), .A3(new_n4868_), .ZN(new_n4877_));
  OAI21_X1   g04685(.A1(new_n4785_), .A2(new_n4877_), .B(new_n4873_), .ZN(new_n4878_));
  AOI21_X1   g04686(.A1(new_n4878_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n4879_));
  AOI21_X1   g04687(.A1(new_n4879_), .A2(new_n4875_), .B(new_n4803_), .ZN(new_n4880_));
  OAI21_X1   g04688(.A1(new_n4880_), .A2(new_n4876_), .B(\asqrt[56] ), .ZN(new_n4881_));
  NAND2_X1   g04689(.A1(new_n4881_), .A2(new_n531_), .ZN(new_n4882_));
  OAI21_X1   g04690(.A1(new_n4882_), .A2(new_n4814_), .B(new_n4821_), .ZN(new_n4883_));
  AOI21_X1   g04691(.A1(new_n4883_), .A2(new_n4815_), .B(new_n436_), .ZN(new_n4884_));
  NOR2_X1    g04692(.A1(new_n4552_), .A2(new_n4542_), .ZN(new_n4885_));
  NOR3_X1    g04693(.A1(new_n4885_), .A2(new_n4519_), .A3(new_n4551_), .ZN(new_n4886_));
  NOR3_X1    g04694(.A1(new_n4696_), .A2(new_n4519_), .A3(new_n4885_), .ZN(new_n4887_));
  INV_X1     g04695(.I(new_n4887_), .ZN(new_n4888_));
  AOI22_X1   g04696(.A1(new_n4888_), .A2(new_n4551_), .B1(\asqrt[38] ), .B2(new_n4886_), .ZN(new_n4889_));
  NOR3_X1    g04697(.A1(new_n4880_), .A2(\asqrt[56] ), .A3(new_n4876_), .ZN(new_n4890_));
  OAI21_X1   g04698(.A1(new_n4811_), .A2(new_n4890_), .B(new_n4881_), .ZN(new_n4891_));
  AOI21_X1   g04699(.A1(new_n4891_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n4892_));
  AOI21_X1   g04700(.A1(new_n4892_), .A2(new_n4883_), .B(new_n4889_), .ZN(new_n4893_));
  OAI21_X1   g04701(.A1(new_n4893_), .A2(new_n4884_), .B(\asqrt[59] ), .ZN(new_n4894_));
  NOR3_X1    g04702(.A1(new_n4696_), .A2(new_n4554_), .A3(new_n4588_), .ZN(new_n4895_));
  INV_X1     g04703(.I(new_n4895_), .ZN(new_n4896_));
  NOR3_X1    g04704(.A1(new_n4554_), .A2(new_n4588_), .A3(new_n4536_), .ZN(new_n4897_));
  AOI22_X1   g04705(.A1(new_n4896_), .A2(new_n4536_), .B1(\asqrt[38] ), .B2(new_n4897_), .ZN(new_n4898_));
  INV_X1     g04706(.I(new_n4898_), .ZN(new_n4899_));
  INV_X1     g04707(.I(new_n4815_), .ZN(new_n4900_));
  NOR3_X1    g04708(.A1(new_n4814_), .A2(new_n4807_), .A3(\asqrt[57] ), .ZN(new_n4901_));
  NOR2_X1    g04709(.A1(new_n4901_), .A2(new_n4820_), .ZN(new_n4902_));
  OAI21_X1   g04710(.A1(new_n4902_), .A2(new_n4900_), .B(\asqrt[58] ), .ZN(new_n4903_));
  NAND2_X1   g04711(.A1(new_n4903_), .A2(new_n327_), .ZN(new_n4904_));
  OAI21_X1   g04712(.A1(new_n4904_), .A2(new_n4893_), .B(new_n4899_), .ZN(new_n4905_));
  AOI21_X1   g04713(.A1(new_n4905_), .A2(new_n4894_), .B(new_n306_), .ZN(new_n4906_));
  NOR2_X1    g04714(.A1(new_n4577_), .A2(new_n4566_), .ZN(new_n4907_));
  NOR3_X1    g04715(.A1(new_n4546_), .A2(new_n4907_), .A3(new_n4576_), .ZN(new_n4908_));
  NOR3_X1    g04716(.A1(new_n4696_), .A2(new_n4546_), .A3(new_n4907_), .ZN(new_n4909_));
  INV_X1     g04717(.I(new_n4909_), .ZN(new_n4910_));
  AOI22_X1   g04718(.A1(new_n4910_), .A2(new_n4576_), .B1(\asqrt[38] ), .B2(new_n4908_), .ZN(new_n4911_));
  INV_X1     g04719(.I(new_n4889_), .ZN(new_n4912_));
  NAND2_X1   g04720(.A1(new_n4815_), .A2(new_n436_), .ZN(new_n4913_));
  OAI21_X1   g04721(.A1(new_n4902_), .A2(new_n4913_), .B(new_n4912_), .ZN(new_n4914_));
  AOI21_X1   g04722(.A1(new_n4914_), .A2(new_n4903_), .B(new_n327_), .ZN(new_n4915_));
  NOR2_X1    g04723(.A1(new_n4915_), .A2(\asqrt[60] ), .ZN(new_n4916_));
  AOI21_X1   g04724(.A1(new_n4916_), .A2(new_n4905_), .B(new_n4911_), .ZN(new_n4917_));
  OAI21_X1   g04725(.A1(new_n4917_), .A2(new_n4906_), .B(\asqrt[61] ), .ZN(new_n4918_));
  NOR2_X1    g04726(.A1(new_n4568_), .A2(new_n4556_), .ZN(new_n4919_));
  NOR3_X1    g04727(.A1(new_n4696_), .A2(new_n4579_), .A3(new_n4919_), .ZN(new_n4920_));
  INV_X1     g04728(.I(new_n4920_), .ZN(new_n4921_));
  NOR3_X1    g04729(.A1(new_n4919_), .A2(new_n4579_), .A3(new_n4564_), .ZN(new_n4922_));
  AOI22_X1   g04730(.A1(new_n4921_), .A2(new_n4564_), .B1(\asqrt[38] ), .B2(new_n4922_), .ZN(new_n4923_));
  INV_X1     g04731(.I(new_n4923_), .ZN(new_n4924_));
  OAI21_X1   g04732(.A1(new_n4820_), .A2(new_n4901_), .B(new_n4815_), .ZN(new_n4925_));
  AOI21_X1   g04733(.A1(new_n4925_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n4926_));
  AOI21_X1   g04734(.A1(new_n4926_), .A2(new_n4914_), .B(new_n4898_), .ZN(new_n4927_));
  OAI21_X1   g04735(.A1(new_n4927_), .A2(new_n4915_), .B(\asqrt[60] ), .ZN(new_n4928_));
  NAND2_X1   g04736(.A1(new_n4928_), .A2(new_n218_), .ZN(new_n4929_));
  OAI21_X1   g04737(.A1(new_n4929_), .A2(new_n4917_), .B(new_n4924_), .ZN(new_n4930_));
  AOI21_X1   g04738(.A1(new_n4930_), .A2(new_n4918_), .B(new_n207_), .ZN(new_n4931_));
  NOR3_X1    g04739(.A1(new_n4570_), .A2(new_n4604_), .A3(new_n4632_), .ZN(new_n4932_));
  NOR3_X1    g04740(.A1(new_n4696_), .A2(new_n4570_), .A3(new_n4604_), .ZN(new_n4933_));
  INV_X1     g04741(.I(new_n4933_), .ZN(new_n4934_));
  AOI22_X1   g04742(.A1(new_n4934_), .A2(new_n4632_), .B1(\asqrt[38] ), .B2(new_n4932_), .ZN(new_n4935_));
  NOR3_X1    g04743(.A1(new_n4927_), .A2(new_n4915_), .A3(\asqrt[60] ), .ZN(new_n4936_));
  OAI21_X1   g04744(.A1(new_n4911_), .A2(new_n4936_), .B(new_n4928_), .ZN(new_n4937_));
  AOI21_X1   g04745(.A1(new_n4937_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n4938_));
  AOI21_X1   g04746(.A1(new_n4938_), .A2(new_n4930_), .B(new_n4935_), .ZN(new_n4939_));
  AND3_X2    g04747(.A1(new_n4582_), .A2(new_n4635_), .A3(new_n4586_), .Z(new_n4940_));
  NAND2_X1   g04748(.A1(\asqrt[38] ), .A2(new_n4940_), .ZN(new_n4941_));
  INV_X1     g04749(.I(new_n4941_), .ZN(new_n4942_));
  AND2_X2    g04750(.A1(new_n4582_), .A2(new_n4635_), .Z(new_n4943_));
  AOI21_X1   g04751(.A1(\asqrt[38] ), .A2(new_n4943_), .B(new_n4586_), .ZN(new_n4944_));
  NOR2_X1    g04752(.A1(new_n4942_), .A2(new_n4944_), .ZN(new_n4945_));
  NOR3_X1    g04753(.A1(new_n4696_), .A2(new_n4636_), .A3(new_n4626_), .ZN(new_n4946_));
  NOR3_X1    g04754(.A1(new_n4945_), .A2(new_n4649_), .A3(new_n4946_), .ZN(new_n4947_));
  OAI21_X1   g04755(.A1(new_n4939_), .A2(new_n4931_), .B(new_n4947_), .ZN(new_n4948_));
  NAND2_X1   g04756(.A1(new_n4948_), .A2(new_n193_), .ZN(new_n4949_));
  INV_X1     g04757(.I(new_n4935_), .ZN(new_n4950_));
  NAND3_X1   g04758(.A1(new_n4930_), .A2(new_n4918_), .A3(new_n207_), .ZN(new_n4951_));
  NAND2_X1   g04759(.A1(new_n4951_), .A2(new_n4950_), .ZN(new_n4952_));
  INV_X1     g04760(.I(new_n4945_), .ZN(new_n4953_));
  NOR2_X1    g04761(.A1(new_n4931_), .A2(new_n4953_), .ZN(new_n4954_));
  AOI21_X1   g04762(.A1(\asqrt[38] ), .A2(new_n4599_), .B(new_n4622_), .ZN(new_n4955_));
  OAI21_X1   g04763(.A1(new_n4636_), .A2(new_n4626_), .B(\asqrt[63] ), .ZN(new_n4956_));
  NOR2_X1    g04764(.A1(new_n4955_), .A2(new_n4956_), .ZN(new_n4957_));
  AND3_X2    g04765(.A1(new_n4598_), .A2(new_n4596_), .A3(new_n4612_), .Z(new_n4958_));
  NAND4_X1   g04766(.A1(new_n4650_), .A2(new_n4637_), .A3(new_n4609_), .A4(new_n4958_), .ZN(new_n4959_));
  INV_X1     g04767(.I(new_n4959_), .ZN(new_n4960_));
  NOR2_X1    g04768(.A1(new_n4957_), .A2(new_n4960_), .ZN(new_n4961_));
  INV_X1     g04769(.I(new_n4961_), .ZN(new_n4962_));
  AOI21_X1   g04770(.A1(new_n4954_), .A2(new_n4952_), .B(new_n4962_), .ZN(new_n4963_));
  NAND2_X1   g04771(.A1(new_n4949_), .A2(new_n4963_), .ZN(\asqrt[37] ));
  NOR2_X1    g04772(.A1(\a[72] ), .A2(\a[73] ), .ZN(new_n4965_));
  INV_X1     g04773(.I(new_n4965_), .ZN(new_n4966_));
  NOR2_X1    g04774(.A1(new_n4966_), .A2(\a[74] ), .ZN(new_n4967_));
  INV_X1     g04775(.I(new_n4967_), .ZN(new_n4968_));
  INV_X1     g04776(.I(new_n4911_), .ZN(new_n4969_));
  NAND2_X1   g04777(.A1(new_n4894_), .A2(new_n306_), .ZN(new_n4970_));
  OAI21_X1   g04778(.A1(new_n4970_), .A2(new_n4927_), .B(new_n4969_), .ZN(new_n4971_));
  AOI21_X1   g04779(.A1(new_n4971_), .A2(new_n4928_), .B(new_n218_), .ZN(new_n4972_));
  NOR3_X1    g04780(.A1(new_n4893_), .A2(\asqrt[59] ), .A3(new_n4884_), .ZN(new_n4973_));
  OAI21_X1   g04781(.A1(new_n4898_), .A2(new_n4973_), .B(new_n4894_), .ZN(new_n4974_));
  AOI21_X1   g04782(.A1(new_n4974_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n4975_));
  AOI21_X1   g04783(.A1(new_n4975_), .A2(new_n4971_), .B(new_n4923_), .ZN(new_n4976_));
  OAI21_X1   g04784(.A1(new_n4976_), .A2(new_n4972_), .B(\asqrt[62] ), .ZN(new_n4977_));
  NOR3_X1    g04785(.A1(new_n4976_), .A2(\asqrt[62] ), .A3(new_n4972_), .ZN(new_n4978_));
  OAI21_X1   g04786(.A1(new_n4935_), .A2(new_n4978_), .B(new_n4977_), .ZN(new_n4979_));
  AOI21_X1   g04787(.A1(new_n4979_), .A2(new_n4947_), .B(\asqrt[63] ), .ZN(new_n4980_));
  NAND2_X1   g04788(.A1(new_n4977_), .A2(new_n4945_), .ZN(new_n4981_));
  OAI21_X1   g04789(.A1(new_n4981_), .A2(new_n4939_), .B(new_n4961_), .ZN(new_n4982_));
  OAI21_X1   g04790(.A1(new_n4980_), .A2(new_n4982_), .B(\a[74] ), .ZN(new_n4983_));
  AOI21_X1   g04791(.A1(new_n4983_), .A2(new_n4968_), .B(new_n4696_), .ZN(new_n4984_));
  INV_X1     g04792(.I(\a[74] ), .ZN(new_n4985_));
  AOI21_X1   g04793(.A1(new_n4949_), .A2(new_n4963_), .B(new_n4985_), .ZN(new_n4986_));
  NAND2_X1   g04794(.A1(new_n4612_), .A2(new_n4968_), .ZN(new_n4987_));
  NOR4_X1    g04795(.A1(new_n4624_), .A2(new_n4649_), .A3(new_n4610_), .A4(new_n4987_), .ZN(new_n4988_));
  INV_X1     g04796(.I(new_n4988_), .ZN(new_n4989_));
  NOR2_X1    g04797(.A1(new_n4986_), .A2(new_n4989_), .ZN(new_n4990_));
  AOI21_X1   g04798(.A1(new_n4949_), .A2(new_n4963_), .B(new_n4619_), .ZN(new_n4991_));
  INV_X1     g04799(.I(\a[75] ), .ZN(new_n4992_));
  AOI21_X1   g04800(.A1(\asqrt[37] ), .A2(new_n4985_), .B(new_n4992_), .ZN(new_n4993_));
  NOR3_X1    g04801(.A1(new_n4990_), .A2(new_n4993_), .A3(new_n4991_), .ZN(new_n4994_));
  OAI21_X1   g04802(.A1(new_n4994_), .A2(new_n4984_), .B(\asqrt[39] ), .ZN(new_n4995_));
  OAI21_X1   g04803(.A1(new_n4980_), .A2(new_n4982_), .B(new_n4618_), .ZN(new_n4996_));
  NAND2_X1   g04804(.A1(new_n4954_), .A2(new_n4952_), .ZN(new_n4997_));
  INV_X1     g04805(.I(new_n4957_), .ZN(new_n4998_));
  NOR2_X1    g04806(.A1(new_n4960_), .A2(new_n4696_), .ZN(new_n4999_));
  NAND4_X1   g04807(.A1(new_n4949_), .A2(new_n4997_), .A3(new_n4998_), .A4(new_n4999_), .ZN(new_n5000_));
  AOI21_X1   g04808(.A1(new_n5000_), .A2(new_n4996_), .B(new_n4631_), .ZN(new_n5001_));
  INV_X1     g04809(.I(new_n4997_), .ZN(new_n5002_));
  NAND2_X1   g04810(.A1(new_n4998_), .A2(new_n4999_), .ZN(new_n5003_));
  NOR3_X1    g04811(.A1(new_n5002_), .A2(new_n4980_), .A3(new_n5003_), .ZN(new_n5004_));
  NOR3_X1    g04812(.A1(new_n5004_), .A2(new_n4991_), .A3(\a[76] ), .ZN(new_n5005_));
  OAI21_X1   g04813(.A1(new_n4986_), .A2(new_n4967_), .B(\asqrt[38] ), .ZN(new_n5006_));
  NAND2_X1   g04814(.A1(new_n5006_), .A2(new_n4298_), .ZN(new_n5007_));
  OAI22_X1   g04815(.A1(new_n4994_), .A2(new_n5007_), .B1(new_n5001_), .B2(new_n5005_), .ZN(new_n5008_));
  AOI21_X1   g04816(.A1(new_n5008_), .A2(new_n4995_), .B(new_n4071_), .ZN(new_n5009_));
  NOR3_X1    g04817(.A1(new_n4841_), .A2(new_n4630_), .A3(new_n4642_), .ZN(new_n5010_));
  NAND3_X1   g04818(.A1(\asqrt[37] ), .A2(new_n4666_), .A3(new_n4826_), .ZN(new_n5011_));
  AOI22_X1   g04819(.A1(new_n5011_), .A2(new_n4841_), .B1(\asqrt[37] ), .B2(new_n5010_), .ZN(new_n5012_));
  AOI21_X1   g04820(.A1(new_n4949_), .A2(new_n4963_), .B(\a[74] ), .ZN(new_n5013_));
  OAI21_X1   g04821(.A1(new_n4992_), .A2(new_n5013_), .B(new_n4996_), .ZN(new_n5014_));
  OAI21_X1   g04822(.A1(new_n5014_), .A2(new_n4990_), .B(new_n5006_), .ZN(new_n5015_));
  AOI21_X1   g04823(.A1(new_n5015_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n5016_));
  AOI21_X1   g04824(.A1(new_n5016_), .A2(new_n5008_), .B(new_n5012_), .ZN(new_n5017_));
  OAI21_X1   g04825(.A1(new_n5017_), .A2(new_n5009_), .B(\asqrt[41] ), .ZN(new_n5018_));
  INV_X1     g04826(.I(new_n5018_), .ZN(new_n5019_));
  NOR2_X1    g04827(.A1(new_n4653_), .A2(new_n4656_), .ZN(new_n5020_));
  NOR2_X1    g04828(.A1(new_n4646_), .A2(new_n4658_), .ZN(new_n5021_));
  INV_X1     g04829(.I(new_n5021_), .ZN(new_n5022_));
  NAND4_X1   g04830(.A1(\asqrt[37] ), .A2(new_n4647_), .A3(new_n5020_), .A4(new_n5022_), .ZN(new_n5023_));
  INV_X1     g04831(.I(\asqrt[37] ), .ZN(new_n5024_));
  NOR3_X1    g04832(.A1(new_n5024_), .A2(new_n4830_), .A3(new_n5021_), .ZN(new_n5025_));
  OAI21_X1   g04833(.A1(new_n5025_), .A2(new_n5020_), .B(new_n5023_), .ZN(new_n5026_));
  INV_X1     g04834(.I(new_n5026_), .ZN(new_n5027_));
  NOR3_X1    g04835(.A1(new_n5017_), .A2(new_n5009_), .A3(\asqrt[41] ), .ZN(new_n5028_));
  NOR2_X1    g04836(.A1(new_n5028_), .A2(new_n5027_), .ZN(new_n5029_));
  OAI21_X1   g04837(.A1(new_n5029_), .A2(new_n5019_), .B(\asqrt[42] ), .ZN(new_n5030_));
  NOR2_X1    g04838(.A1(new_n4843_), .A2(new_n4835_), .ZN(new_n5031_));
  NOR3_X1    g04839(.A1(new_n5024_), .A2(new_n4660_), .A3(new_n5031_), .ZN(new_n5032_));
  INV_X1     g04840(.I(new_n5032_), .ZN(new_n5033_));
  NOR3_X1    g04841(.A1(new_n5031_), .A2(new_n4660_), .A3(new_n4840_), .ZN(new_n5034_));
  AOI22_X1   g04842(.A1(new_n5033_), .A2(new_n4840_), .B1(\asqrt[37] ), .B2(new_n5034_), .ZN(new_n5035_));
  INV_X1     g04843(.I(new_n5035_), .ZN(new_n5036_));
  NAND2_X1   g04844(.A1(new_n5018_), .A2(new_n3419_), .ZN(new_n5037_));
  OAI21_X1   g04845(.A1(new_n5029_), .A2(new_n5037_), .B(new_n5036_), .ZN(new_n5038_));
  AOI21_X1   g04846(.A1(new_n5038_), .A2(new_n5030_), .B(new_n3218_), .ZN(new_n5039_));
  NOR3_X1    g04847(.A1(new_n4673_), .A2(new_n4681_), .A3(new_n4679_), .ZN(new_n5040_));
  NOR3_X1    g04848(.A1(new_n5024_), .A2(new_n4673_), .A3(new_n4681_), .ZN(new_n5041_));
  INV_X1     g04849(.I(new_n5041_), .ZN(new_n5042_));
  AOI22_X1   g04850(.A1(new_n5042_), .A2(new_n4679_), .B1(\asqrt[37] ), .B2(new_n5040_), .ZN(new_n5043_));
  OAI21_X1   g04851(.A1(new_n5027_), .A2(new_n5028_), .B(new_n5018_), .ZN(new_n5044_));
  AOI21_X1   g04852(.A1(new_n5044_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n5045_));
  AOI21_X1   g04853(.A1(new_n5045_), .A2(new_n5038_), .B(new_n5043_), .ZN(new_n5046_));
  OAI21_X1   g04854(.A1(new_n5046_), .A2(new_n5039_), .B(\asqrt[44] ), .ZN(new_n5047_));
  NAND2_X1   g04855(.A1(new_n4846_), .A2(new_n4838_), .ZN(new_n5048_));
  NAND3_X1   g04856(.A1(\asqrt[37] ), .A2(new_n4683_), .A3(new_n5048_), .ZN(new_n5049_));
  AND3_X2    g04857(.A1(new_n4683_), .A2(new_n4689_), .A3(new_n5048_), .Z(new_n5050_));
  AOI22_X1   g04858(.A1(new_n5049_), .A2(new_n4690_), .B1(\asqrt[37] ), .B2(new_n5050_), .ZN(new_n5051_));
  INV_X1     g04859(.I(new_n5051_), .ZN(new_n5052_));
  NAND2_X1   g04860(.A1(new_n4983_), .A2(new_n4988_), .ZN(new_n5053_));
  OAI21_X1   g04861(.A1(new_n4980_), .A2(new_n4982_), .B(new_n4985_), .ZN(new_n5054_));
  NAND2_X1   g04862(.A1(new_n5054_), .A2(\a[75] ), .ZN(new_n5055_));
  NAND3_X1   g04863(.A1(new_n5053_), .A2(new_n5055_), .A3(new_n4996_), .ZN(new_n5056_));
  AOI21_X1   g04864(.A1(new_n5056_), .A2(new_n5006_), .B(new_n4298_), .ZN(new_n5057_));
  OAI21_X1   g04865(.A1(new_n5004_), .A2(new_n4991_), .B(\a[76] ), .ZN(new_n5058_));
  NAND3_X1   g04866(.A1(new_n5000_), .A2(new_n4996_), .A3(new_n4631_), .ZN(new_n5059_));
  NAND2_X1   g04867(.A1(new_n4983_), .A2(new_n4968_), .ZN(new_n5060_));
  AOI21_X1   g04868(.A1(new_n5060_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n5061_));
  AOI22_X1   g04869(.A1(new_n5056_), .A2(new_n5061_), .B1(new_n5058_), .B2(new_n5059_), .ZN(new_n5062_));
  OAI21_X1   g04870(.A1(new_n5062_), .A2(new_n5057_), .B(\asqrt[40] ), .ZN(new_n5063_));
  NAND2_X1   g04871(.A1(new_n5063_), .A2(new_n3782_), .ZN(new_n5064_));
  OAI21_X1   g04872(.A1(new_n5064_), .A2(new_n5017_), .B(new_n5026_), .ZN(new_n5065_));
  AOI21_X1   g04873(.A1(new_n5065_), .A2(new_n5018_), .B(new_n3419_), .ZN(new_n5066_));
  INV_X1     g04874(.I(new_n5012_), .ZN(new_n5067_));
  AOI21_X1   g04875(.A1(\a[75] ), .A2(new_n5054_), .B(new_n4991_), .ZN(new_n5068_));
  AOI21_X1   g04876(.A1(new_n5068_), .A2(new_n5053_), .B(new_n4984_), .ZN(new_n5069_));
  OAI21_X1   g04877(.A1(new_n5069_), .A2(new_n4298_), .B(new_n4071_), .ZN(new_n5070_));
  OAI21_X1   g04878(.A1(new_n5070_), .A2(new_n5062_), .B(new_n5067_), .ZN(new_n5071_));
  NAND2_X1   g04879(.A1(new_n5071_), .A2(new_n5063_), .ZN(new_n5072_));
  AOI21_X1   g04880(.A1(new_n5072_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n5073_));
  AOI21_X1   g04881(.A1(new_n5073_), .A2(new_n5065_), .B(new_n5035_), .ZN(new_n5074_));
  OAI21_X1   g04882(.A1(new_n5074_), .A2(new_n5066_), .B(\asqrt[43] ), .ZN(new_n5075_));
  NAND2_X1   g04883(.A1(new_n5075_), .A2(new_n2954_), .ZN(new_n5076_));
  OAI21_X1   g04884(.A1(new_n5076_), .A2(new_n5046_), .B(new_n5052_), .ZN(new_n5077_));
  AOI21_X1   g04885(.A1(new_n5077_), .A2(new_n5047_), .B(new_n2641_), .ZN(new_n5078_));
  INV_X1     g04886(.I(new_n4699_), .ZN(new_n5079_));
  NOR3_X1    g04887(.A1(new_n4693_), .A2(new_n4857_), .A3(new_n5079_), .ZN(new_n5080_));
  NOR3_X1    g04888(.A1(new_n5024_), .A2(new_n4693_), .A3(new_n4857_), .ZN(new_n5081_));
  INV_X1     g04889(.I(new_n5081_), .ZN(new_n5082_));
  AOI22_X1   g04890(.A1(new_n5082_), .A2(new_n5079_), .B1(\asqrt[37] ), .B2(new_n5080_), .ZN(new_n5083_));
  NOR3_X1    g04891(.A1(new_n5074_), .A2(new_n5066_), .A3(\asqrt[43] ), .ZN(new_n5084_));
  OAI21_X1   g04892(.A1(new_n5043_), .A2(new_n5084_), .B(new_n5075_), .ZN(new_n5085_));
  AOI21_X1   g04893(.A1(new_n5085_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n5086_));
  AOI21_X1   g04894(.A1(new_n5086_), .A2(new_n5077_), .B(new_n5083_), .ZN(new_n5087_));
  OAI21_X1   g04895(.A1(new_n5087_), .A2(new_n5078_), .B(\asqrt[46] ), .ZN(new_n5088_));
  INV_X1     g04896(.I(new_n5088_), .ZN(new_n5089_));
  NOR3_X1    g04897(.A1(new_n5024_), .A2(new_n4704_), .A3(new_n4711_), .ZN(new_n5090_));
  INV_X1     g04898(.I(new_n5090_), .ZN(new_n5091_));
  NOR3_X1    g04899(.A1(new_n4704_), .A2(new_n4825_), .A3(new_n4711_), .ZN(new_n5092_));
  AOI22_X1   g04900(.A1(new_n5091_), .A2(new_n4825_), .B1(\asqrt[37] ), .B2(new_n5092_), .ZN(new_n5093_));
  NOR3_X1    g04901(.A1(new_n5087_), .A2(\asqrt[46] ), .A3(new_n5078_), .ZN(new_n5094_));
  NOR2_X1    g04902(.A1(new_n5094_), .A2(new_n5093_), .ZN(new_n5095_));
  OAI21_X1   g04903(.A1(new_n5095_), .A2(new_n5089_), .B(\asqrt[47] ), .ZN(new_n5096_));
  INV_X1     g04904(.I(new_n4851_), .ZN(new_n5097_));
  NOR3_X1    g04905(.A1(new_n5097_), .A2(new_n4856_), .A3(new_n4722_), .ZN(new_n5098_));
  NOR3_X1    g04906(.A1(new_n5024_), .A2(new_n4856_), .A3(new_n5097_), .ZN(new_n5099_));
  INV_X1     g04907(.I(new_n5099_), .ZN(new_n5100_));
  AOI22_X1   g04908(.A1(new_n5100_), .A2(new_n4722_), .B1(\asqrt[37] ), .B2(new_n5098_), .ZN(new_n5101_));
  INV_X1     g04909(.I(new_n5101_), .ZN(new_n5102_));
  NAND2_X1   g04910(.A1(new_n5088_), .A2(new_n2229_), .ZN(new_n5103_));
  OAI21_X1   g04911(.A1(new_n5095_), .A2(new_n5103_), .B(new_n5102_), .ZN(new_n5104_));
  AOI21_X1   g04912(.A1(new_n5104_), .A2(new_n5096_), .B(new_n1956_), .ZN(new_n5105_));
  INV_X1     g04913(.I(new_n4730_), .ZN(new_n5106_));
  NOR3_X1    g04914(.A1(new_n5024_), .A2(new_n4725_), .A3(new_n4861_), .ZN(new_n5107_));
  INV_X1     g04915(.I(new_n5107_), .ZN(new_n5108_));
  NOR3_X1    g04916(.A1(new_n4725_), .A2(new_n4861_), .A3(new_n5106_), .ZN(new_n5109_));
  AOI22_X1   g04917(.A1(new_n5108_), .A2(new_n5106_), .B1(\asqrt[37] ), .B2(new_n5109_), .ZN(new_n5110_));
  NOR3_X1    g04918(.A1(new_n5046_), .A2(new_n5039_), .A3(\asqrt[44] ), .ZN(new_n5111_));
  OAI21_X1   g04919(.A1(new_n5051_), .A2(new_n5111_), .B(new_n5047_), .ZN(new_n5112_));
  INV_X1     g04920(.I(new_n5083_), .ZN(new_n5113_));
  NAND3_X1   g04921(.A1(new_n5077_), .A2(new_n2641_), .A3(new_n5047_), .ZN(new_n5114_));
  AOI22_X1   g04922(.A1(new_n5114_), .A2(new_n5113_), .B1(new_n5112_), .B2(\asqrt[45] ), .ZN(new_n5115_));
  OAI22_X1   g04923(.A1(new_n5094_), .A2(new_n5093_), .B1(new_n5115_), .B2(new_n2465_), .ZN(new_n5116_));
  AOI21_X1   g04924(.A1(new_n5116_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n5117_));
  AOI21_X1   g04925(.A1(new_n5117_), .A2(new_n5104_), .B(new_n5110_), .ZN(new_n5118_));
  OAI21_X1   g04926(.A1(new_n5118_), .A2(new_n5105_), .B(\asqrt[49] ), .ZN(new_n5119_));
  INV_X1     g04927(.I(new_n5119_), .ZN(new_n5120_));
  NOR3_X1    g04928(.A1(new_n4735_), .A2(new_n4824_), .A3(new_n4741_), .ZN(new_n5121_));
  NOR3_X1    g04929(.A1(new_n5024_), .A2(new_n4735_), .A3(new_n4741_), .ZN(new_n5122_));
  INV_X1     g04930(.I(new_n5122_), .ZN(new_n5123_));
  AOI22_X1   g04931(.A1(new_n5123_), .A2(new_n4824_), .B1(\asqrt[37] ), .B2(new_n5121_), .ZN(new_n5124_));
  NOR3_X1    g04932(.A1(new_n5118_), .A2(new_n5105_), .A3(\asqrt[49] ), .ZN(new_n5125_));
  NOR2_X1    g04933(.A1(new_n5125_), .A2(new_n5124_), .ZN(new_n5126_));
  OAI21_X1   g04934(.A1(new_n5126_), .A2(new_n5120_), .B(\asqrt[50] ), .ZN(new_n5127_));
  NOR2_X1    g04935(.A1(new_n4742_), .A2(new_n4753_), .ZN(new_n5128_));
  NOR3_X1    g04936(.A1(new_n5024_), .A2(new_n4855_), .A3(new_n5128_), .ZN(new_n5129_));
  INV_X1     g04937(.I(new_n5129_), .ZN(new_n5130_));
  NOR3_X1    g04938(.A1(new_n5128_), .A2(new_n4855_), .A3(new_n4752_), .ZN(new_n5131_));
  AOI22_X1   g04939(.A1(new_n5130_), .A2(new_n4752_), .B1(\asqrt[37] ), .B2(new_n5131_), .ZN(new_n5132_));
  INV_X1     g04940(.I(new_n5132_), .ZN(new_n5133_));
  NAND2_X1   g04941(.A1(new_n5119_), .A2(new_n1612_), .ZN(new_n5134_));
  OAI21_X1   g04942(.A1(new_n5126_), .A2(new_n5134_), .B(new_n5133_), .ZN(new_n5135_));
  AOI21_X1   g04943(.A1(new_n5135_), .A2(new_n5127_), .B(new_n1376_), .ZN(new_n5136_));
  INV_X1     g04944(.I(new_n4759_), .ZN(new_n5137_));
  NOR3_X1    g04945(.A1(new_n4755_), .A2(new_n4869_), .A3(new_n5137_), .ZN(new_n5138_));
  NOR3_X1    g04946(.A1(new_n5024_), .A2(new_n4755_), .A3(new_n4869_), .ZN(new_n5139_));
  INV_X1     g04947(.I(new_n5139_), .ZN(new_n5140_));
  AOI22_X1   g04948(.A1(new_n5140_), .A2(new_n5137_), .B1(\asqrt[37] ), .B2(new_n5138_), .ZN(new_n5141_));
  OAI21_X1   g04949(.A1(new_n5124_), .A2(new_n5125_), .B(new_n5119_), .ZN(new_n5142_));
  AOI21_X1   g04950(.A1(new_n5142_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n5143_));
  AOI21_X1   g04951(.A1(new_n5143_), .A2(new_n5135_), .B(new_n5141_), .ZN(new_n5144_));
  OAI21_X1   g04952(.A1(new_n5144_), .A2(new_n5136_), .B(\asqrt[52] ), .ZN(new_n5145_));
  INV_X1     g04953(.I(new_n5145_), .ZN(new_n5146_));
  INV_X1     g04954(.I(new_n5144_), .ZN(new_n5147_));
  NOR3_X1    g04955(.A1(new_n5024_), .A2(new_n4764_), .A3(new_n4770_), .ZN(new_n5148_));
  INV_X1     g04956(.I(new_n5148_), .ZN(new_n5149_));
  NOR3_X1    g04957(.A1(new_n4764_), .A2(new_n4823_), .A3(new_n4770_), .ZN(new_n5150_));
  AOI22_X1   g04958(.A1(new_n5149_), .A2(new_n4823_), .B1(\asqrt[37] ), .B2(new_n5150_), .ZN(new_n5151_));
  NOR2_X1    g04959(.A1(new_n5136_), .A2(\asqrt[52] ), .ZN(new_n5152_));
  AOI21_X1   g04960(.A1(new_n5147_), .A2(new_n5152_), .B(new_n5151_), .ZN(new_n5153_));
  OAI21_X1   g04961(.A1(new_n5153_), .A2(new_n5146_), .B(\asqrt[53] ), .ZN(new_n5154_));
  NOR2_X1    g04962(.A1(new_n4771_), .A2(new_n4779_), .ZN(new_n5155_));
  NOR3_X1    g04963(.A1(new_n5155_), .A2(new_n4868_), .A3(new_n4778_), .ZN(new_n5156_));
  NOR3_X1    g04964(.A1(new_n5024_), .A2(new_n4868_), .A3(new_n5155_), .ZN(new_n5157_));
  INV_X1     g04965(.I(new_n5157_), .ZN(new_n5158_));
  AOI22_X1   g04966(.A1(new_n5158_), .A2(new_n4778_), .B1(\asqrt[37] ), .B2(new_n5156_), .ZN(new_n5159_));
  INV_X1     g04967(.I(new_n5159_), .ZN(new_n5160_));
  NAND2_X1   g04968(.A1(new_n5145_), .A2(new_n1103_), .ZN(new_n5161_));
  OAI21_X1   g04969(.A1(new_n5161_), .A2(new_n5153_), .B(new_n5160_), .ZN(new_n5162_));
  AOI21_X1   g04970(.A1(new_n5162_), .A2(new_n5154_), .B(new_n904_), .ZN(new_n5163_));
  INV_X1     g04971(.I(new_n5163_), .ZN(new_n5164_));
  INV_X1     g04972(.I(new_n5162_), .ZN(new_n5165_));
  INV_X1     g04973(.I(new_n4785_), .ZN(new_n5166_));
  NOR3_X1    g04974(.A1(new_n5024_), .A2(new_n4781_), .A3(new_n4877_), .ZN(new_n5167_));
  INV_X1     g04975(.I(new_n5167_), .ZN(new_n5168_));
  NOR3_X1    g04976(.A1(new_n4781_), .A2(new_n4877_), .A3(new_n5166_), .ZN(new_n5169_));
  AOI22_X1   g04977(.A1(new_n5168_), .A2(new_n5166_), .B1(\asqrt[37] ), .B2(new_n5169_), .ZN(new_n5170_));
  INV_X1     g04978(.I(new_n5170_), .ZN(new_n5171_));
  NAND2_X1   g04979(.A1(new_n5154_), .A2(new_n904_), .ZN(new_n5172_));
  OAI21_X1   g04980(.A1(new_n5172_), .A2(new_n5165_), .B(new_n5171_), .ZN(new_n5173_));
  AOI21_X1   g04981(.A1(new_n5173_), .A2(new_n5164_), .B(new_n823_), .ZN(new_n5174_));
  NOR3_X1    g04982(.A1(new_n4790_), .A2(new_n4822_), .A3(new_n4796_), .ZN(new_n5175_));
  NOR3_X1    g04983(.A1(new_n5024_), .A2(new_n4790_), .A3(new_n4796_), .ZN(new_n5176_));
  INV_X1     g04984(.I(new_n5176_), .ZN(new_n5177_));
  AOI22_X1   g04985(.A1(new_n5177_), .A2(new_n4822_), .B1(\asqrt[37] ), .B2(new_n5175_), .ZN(new_n5178_));
  NOR2_X1    g04986(.A1(new_n5163_), .A2(\asqrt[55] ), .ZN(new_n5179_));
  AOI21_X1   g04987(.A1(new_n5179_), .A2(new_n5173_), .B(new_n5178_), .ZN(new_n5180_));
  OAI21_X1   g04988(.A1(new_n5180_), .A2(new_n5174_), .B(\asqrt[56] ), .ZN(new_n5181_));
  NOR2_X1    g04989(.A1(new_n4797_), .A2(new_n4805_), .ZN(new_n5182_));
  NOR3_X1    g04990(.A1(new_n5024_), .A2(new_n4876_), .A3(new_n5182_), .ZN(new_n5183_));
  INV_X1     g04991(.I(new_n5183_), .ZN(new_n5184_));
  NOR3_X1    g04992(.A1(new_n5182_), .A2(new_n4876_), .A3(new_n4804_), .ZN(new_n5185_));
  AOI22_X1   g04993(.A1(new_n5184_), .A2(new_n4804_), .B1(\asqrt[37] ), .B2(new_n5185_), .ZN(new_n5186_));
  INV_X1     g04994(.I(new_n5186_), .ZN(new_n5187_));
  NOR3_X1    g04995(.A1(new_n5144_), .A2(new_n5136_), .A3(\asqrt[52] ), .ZN(new_n5188_));
  OAI21_X1   g04996(.A1(new_n5151_), .A2(new_n5188_), .B(new_n5145_), .ZN(new_n5189_));
  AOI21_X1   g04997(.A1(new_n5189_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n5190_));
  AOI21_X1   g04998(.A1(new_n5190_), .A2(new_n5162_), .B(new_n5170_), .ZN(new_n5191_));
  OAI21_X1   g04999(.A1(new_n5191_), .A2(new_n5163_), .B(\asqrt[55] ), .ZN(new_n5192_));
  NAND2_X1   g05000(.A1(new_n5192_), .A2(new_n703_), .ZN(new_n5193_));
  OAI21_X1   g05001(.A1(new_n5193_), .A2(new_n5180_), .B(new_n5187_), .ZN(new_n5194_));
  AOI21_X1   g05002(.A1(new_n5194_), .A2(new_n5181_), .B(new_n531_), .ZN(new_n5195_));
  INV_X1     g05003(.I(new_n5195_), .ZN(new_n5196_));
  INV_X1     g05004(.I(new_n5194_), .ZN(new_n5197_));
  INV_X1     g05005(.I(new_n4811_), .ZN(new_n5198_));
  NOR3_X1    g05006(.A1(new_n4807_), .A2(new_n4890_), .A3(new_n5198_), .ZN(new_n5199_));
  NOR3_X1    g05007(.A1(new_n5024_), .A2(new_n4807_), .A3(new_n4890_), .ZN(new_n5200_));
  INV_X1     g05008(.I(new_n5200_), .ZN(new_n5201_));
  AOI22_X1   g05009(.A1(new_n5201_), .A2(new_n5198_), .B1(\asqrt[37] ), .B2(new_n5199_), .ZN(new_n5202_));
  INV_X1     g05010(.I(new_n5202_), .ZN(new_n5203_));
  NAND2_X1   g05011(.A1(new_n5181_), .A2(new_n531_), .ZN(new_n5204_));
  OAI21_X1   g05012(.A1(new_n5204_), .A2(new_n5197_), .B(new_n5203_), .ZN(new_n5205_));
  AOI21_X1   g05013(.A1(new_n5205_), .A2(new_n5196_), .B(new_n436_), .ZN(new_n5206_));
  NOR3_X1    g05014(.A1(new_n5024_), .A2(new_n4900_), .A3(new_n4901_), .ZN(new_n5207_));
  INV_X1     g05015(.I(new_n5207_), .ZN(new_n5208_));
  NOR3_X1    g05016(.A1(new_n4900_), .A2(new_n4901_), .A3(new_n4821_), .ZN(new_n5209_));
  AOI22_X1   g05017(.A1(new_n5208_), .A2(new_n4821_), .B1(\asqrt[37] ), .B2(new_n5209_), .ZN(new_n5210_));
  NOR2_X1    g05018(.A1(new_n5195_), .A2(\asqrt[58] ), .ZN(new_n5211_));
  AOI21_X1   g05019(.A1(new_n5211_), .A2(new_n5205_), .B(new_n5210_), .ZN(new_n5212_));
  OAI21_X1   g05020(.A1(new_n5212_), .A2(new_n5206_), .B(\asqrt[59] ), .ZN(new_n5213_));
  NOR2_X1    g05021(.A1(new_n4902_), .A2(new_n4913_), .ZN(new_n5214_));
  NOR3_X1    g05022(.A1(new_n5214_), .A2(new_n4884_), .A3(new_n4912_), .ZN(new_n5215_));
  NOR3_X1    g05023(.A1(new_n5024_), .A2(new_n4884_), .A3(new_n5214_), .ZN(new_n5216_));
  INV_X1     g05024(.I(new_n5216_), .ZN(new_n5217_));
  AOI22_X1   g05025(.A1(new_n5217_), .A2(new_n4912_), .B1(\asqrt[37] ), .B2(new_n5215_), .ZN(new_n5218_));
  INV_X1     g05026(.I(new_n5218_), .ZN(new_n5219_));
  NOR3_X1    g05027(.A1(new_n5191_), .A2(\asqrt[55] ), .A3(new_n5163_), .ZN(new_n5220_));
  OAI21_X1   g05028(.A1(new_n5178_), .A2(new_n5220_), .B(new_n5192_), .ZN(new_n5221_));
  AOI21_X1   g05029(.A1(new_n5221_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n5222_));
  AOI21_X1   g05030(.A1(new_n5222_), .A2(new_n5194_), .B(new_n5202_), .ZN(new_n5223_));
  OAI21_X1   g05031(.A1(new_n5223_), .A2(new_n5195_), .B(\asqrt[58] ), .ZN(new_n5224_));
  NAND2_X1   g05032(.A1(new_n5224_), .A2(new_n327_), .ZN(new_n5225_));
  OAI21_X1   g05033(.A1(new_n5225_), .A2(new_n5212_), .B(new_n5219_), .ZN(new_n5226_));
  AOI21_X1   g05034(.A1(new_n5226_), .A2(new_n5213_), .B(new_n306_), .ZN(new_n5227_));
  INV_X1     g05035(.I(new_n5227_), .ZN(new_n5228_));
  INV_X1     g05036(.I(new_n5226_), .ZN(new_n5229_));
  NOR3_X1    g05037(.A1(new_n5024_), .A2(new_n4915_), .A3(new_n4973_), .ZN(new_n5230_));
  INV_X1     g05038(.I(new_n5230_), .ZN(new_n5231_));
  NOR3_X1    g05039(.A1(new_n4915_), .A2(new_n4973_), .A3(new_n4899_), .ZN(new_n5232_));
  AOI22_X1   g05040(.A1(new_n5231_), .A2(new_n4899_), .B1(\asqrt[37] ), .B2(new_n5232_), .ZN(new_n5233_));
  INV_X1     g05041(.I(new_n5233_), .ZN(new_n5234_));
  NAND2_X1   g05042(.A1(new_n5213_), .A2(new_n306_), .ZN(new_n5235_));
  OAI21_X1   g05043(.A1(new_n5229_), .A2(new_n5235_), .B(new_n5234_), .ZN(new_n5236_));
  AOI21_X1   g05044(.A1(new_n5236_), .A2(new_n5228_), .B(new_n218_), .ZN(new_n5237_));
  NOR3_X1    g05045(.A1(new_n4906_), .A2(new_n4936_), .A3(new_n4969_), .ZN(new_n5238_));
  NOR3_X1    g05046(.A1(new_n5024_), .A2(new_n4906_), .A3(new_n4936_), .ZN(new_n5239_));
  INV_X1     g05047(.I(new_n5239_), .ZN(new_n5240_));
  AOI22_X1   g05048(.A1(new_n5240_), .A2(new_n4969_), .B1(\asqrt[37] ), .B2(new_n5238_), .ZN(new_n5241_));
  NOR2_X1    g05049(.A1(new_n5227_), .A2(\asqrt[61] ), .ZN(new_n5242_));
  AOI21_X1   g05050(.A1(new_n5242_), .A2(new_n5236_), .B(new_n5241_), .ZN(new_n5243_));
  OAI21_X1   g05051(.A1(new_n5243_), .A2(new_n5237_), .B(\asqrt[62] ), .ZN(new_n5244_));
  NOR2_X1    g05052(.A1(new_n4929_), .A2(new_n4917_), .ZN(new_n5245_));
  NOR3_X1    g05053(.A1(new_n5024_), .A2(new_n4972_), .A3(new_n5245_), .ZN(new_n5246_));
  INV_X1     g05054(.I(new_n5246_), .ZN(new_n5247_));
  NOR3_X1    g05055(.A1(new_n5245_), .A2(new_n4972_), .A3(new_n4924_), .ZN(new_n5248_));
  AOI22_X1   g05056(.A1(new_n5247_), .A2(new_n4924_), .B1(\asqrt[37] ), .B2(new_n5248_), .ZN(new_n5249_));
  INV_X1     g05057(.I(new_n5249_), .ZN(new_n5250_));
  NOR3_X1    g05058(.A1(new_n5223_), .A2(\asqrt[58] ), .A3(new_n5195_), .ZN(new_n5251_));
  OAI21_X1   g05059(.A1(new_n5210_), .A2(new_n5251_), .B(new_n5224_), .ZN(new_n5252_));
  AOI21_X1   g05060(.A1(new_n5252_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n5253_));
  AOI21_X1   g05061(.A1(new_n5253_), .A2(new_n5226_), .B(new_n5233_), .ZN(new_n5254_));
  OAI21_X1   g05062(.A1(new_n5254_), .A2(new_n5227_), .B(\asqrt[61] ), .ZN(new_n5255_));
  NAND2_X1   g05063(.A1(new_n5255_), .A2(new_n207_), .ZN(new_n5256_));
  OAI21_X1   g05064(.A1(new_n5256_), .A2(new_n5243_), .B(new_n5250_), .ZN(new_n5257_));
  NAND4_X1   g05065(.A1(\asqrt[37] ), .A2(new_n4977_), .A3(new_n4935_), .A4(new_n4951_), .ZN(new_n5258_));
  NAND2_X1   g05066(.A1(new_n4977_), .A2(new_n4951_), .ZN(new_n5259_));
  OAI21_X1   g05067(.A1(new_n5024_), .A2(new_n5259_), .B(new_n4950_), .ZN(new_n5260_));
  NAND2_X1   g05068(.A1(new_n5260_), .A2(new_n5258_), .ZN(new_n5261_));
  AOI21_X1   g05069(.A1(new_n4952_), .A2(new_n4977_), .B(new_n4945_), .ZN(new_n5262_));
  AOI21_X1   g05070(.A1(\asqrt[37] ), .A2(new_n5262_), .B(new_n5002_), .ZN(new_n5263_));
  NAND2_X1   g05071(.A1(new_n5261_), .A2(new_n5263_), .ZN(new_n5264_));
  AOI21_X1   g05072(.A1(new_n5257_), .A2(new_n5244_), .B(new_n5264_), .ZN(new_n5265_));
  NOR3_X1    g05073(.A1(new_n5254_), .A2(\asqrt[61] ), .A3(new_n5227_), .ZN(new_n5266_));
  OAI21_X1   g05074(.A1(new_n5241_), .A2(new_n5266_), .B(new_n5255_), .ZN(new_n5267_));
  AOI21_X1   g05075(.A1(new_n5267_), .A2(\asqrt[62] ), .B(new_n5261_), .ZN(new_n5268_));
  AOI21_X1   g05076(.A1(\asqrt[37] ), .A2(new_n4953_), .B(new_n4979_), .ZN(new_n5269_));
  OR3_X2     g05077(.A1(new_n5269_), .A2(new_n193_), .A3(new_n5262_), .Z(new_n5270_));
  NAND2_X1   g05078(.A1(new_n4941_), .A2(new_n4959_), .ZN(new_n5271_));
  NOR4_X1    g05079(.A1(new_n5002_), .A2(new_n4944_), .A3(new_n4957_), .A4(new_n5271_), .ZN(new_n5272_));
  NAND2_X1   g05080(.A1(new_n5272_), .A2(new_n4949_), .ZN(new_n5273_));
  NAND2_X1   g05081(.A1(new_n5270_), .A2(new_n5273_), .ZN(new_n5274_));
  AOI21_X1   g05082(.A1(new_n5268_), .A2(new_n5257_), .B(new_n5274_), .ZN(new_n5275_));
  OAI21_X1   g05083(.A1(\asqrt[63] ), .A2(new_n5265_), .B(new_n5275_), .ZN(\asqrt[36] ));
  INV_X1     g05084(.I(\asqrt[36] ), .ZN(new_n5277_));
  NOR2_X1    g05085(.A1(\a[70] ), .A2(\a[71] ), .ZN(new_n5278_));
  INV_X1     g05086(.I(new_n5278_), .ZN(new_n5279_));
  NOR2_X1    g05087(.A1(new_n5279_), .A2(\a[72] ), .ZN(new_n5280_));
  INV_X1     g05088(.I(\a[72] ), .ZN(new_n5281_));
  INV_X1     g05089(.I(new_n5241_), .ZN(new_n5282_));
  INV_X1     g05090(.I(new_n5210_), .ZN(new_n5283_));
  INV_X1     g05091(.I(new_n5178_), .ZN(new_n5284_));
  INV_X1     g05092(.I(new_n5151_), .ZN(new_n5285_));
  INV_X1     g05093(.I(new_n5124_), .ZN(new_n5286_));
  INV_X1     g05094(.I(new_n5093_), .ZN(new_n5287_));
  INV_X1     g05095(.I(new_n5047_), .ZN(new_n5288_));
  NOR2_X1    g05096(.A1(new_n5111_), .A2(new_n5051_), .ZN(new_n5289_));
  OAI21_X1   g05097(.A1(new_n5289_), .A2(new_n5288_), .B(\asqrt[45] ), .ZN(new_n5290_));
  NAND2_X1   g05098(.A1(new_n5290_), .A2(new_n2465_), .ZN(new_n5291_));
  OAI21_X1   g05099(.A1(new_n5291_), .A2(new_n5087_), .B(new_n5287_), .ZN(new_n5292_));
  NAND3_X1   g05100(.A1(new_n5292_), .A2(new_n2229_), .A3(new_n5088_), .ZN(new_n5293_));
  AOI22_X1   g05101(.A1(new_n5293_), .A2(new_n5102_), .B1(\asqrt[47] ), .B2(new_n5116_), .ZN(new_n5294_));
  OAI21_X1   g05102(.A1(new_n5294_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n5295_));
  OAI21_X1   g05103(.A1(new_n5295_), .A2(new_n5118_), .B(new_n5286_), .ZN(new_n5296_));
  NAND3_X1   g05104(.A1(new_n5296_), .A2(new_n1612_), .A3(new_n5119_), .ZN(new_n5297_));
  AOI22_X1   g05105(.A1(new_n5297_), .A2(new_n5133_), .B1(\asqrt[50] ), .B2(new_n5142_), .ZN(new_n5298_));
  OAI21_X1   g05106(.A1(new_n5298_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n5299_));
  OAI21_X1   g05107(.A1(new_n5299_), .A2(new_n5144_), .B(new_n5285_), .ZN(new_n5300_));
  NAND3_X1   g05108(.A1(new_n5300_), .A2(new_n1103_), .A3(new_n5145_), .ZN(new_n5301_));
  AOI22_X1   g05109(.A1(new_n5301_), .A2(new_n5160_), .B1(\asqrt[53] ), .B2(new_n5189_), .ZN(new_n5302_));
  OAI21_X1   g05110(.A1(new_n5302_), .A2(new_n904_), .B(new_n823_), .ZN(new_n5303_));
  OAI21_X1   g05111(.A1(new_n5303_), .A2(new_n5191_), .B(new_n5284_), .ZN(new_n5304_));
  NAND3_X1   g05112(.A1(new_n5304_), .A2(new_n703_), .A3(new_n5192_), .ZN(new_n5305_));
  AOI22_X1   g05113(.A1(new_n5305_), .A2(new_n5187_), .B1(\asqrt[56] ), .B2(new_n5221_), .ZN(new_n5306_));
  OAI21_X1   g05114(.A1(new_n5306_), .A2(new_n531_), .B(new_n436_), .ZN(new_n5307_));
  OAI21_X1   g05115(.A1(new_n5307_), .A2(new_n5223_), .B(new_n5283_), .ZN(new_n5308_));
  NAND3_X1   g05116(.A1(new_n5308_), .A2(new_n327_), .A3(new_n5224_), .ZN(new_n5309_));
  AOI22_X1   g05117(.A1(new_n5309_), .A2(new_n5219_), .B1(\asqrt[59] ), .B2(new_n5252_), .ZN(new_n5310_));
  OAI21_X1   g05118(.A1(new_n5310_), .A2(new_n306_), .B(new_n218_), .ZN(new_n5311_));
  OAI21_X1   g05119(.A1(new_n5311_), .A2(new_n5254_), .B(new_n5282_), .ZN(new_n5312_));
  NAND3_X1   g05120(.A1(new_n5312_), .A2(new_n207_), .A3(new_n5255_), .ZN(new_n5313_));
  AOI22_X1   g05121(.A1(new_n5313_), .A2(new_n5250_), .B1(new_n5267_), .B2(\asqrt[62] ), .ZN(new_n5314_));
  OAI21_X1   g05122(.A1(new_n5314_), .A2(new_n5264_), .B(new_n193_), .ZN(new_n5315_));
  AOI21_X1   g05123(.A1(new_n5315_), .A2(new_n5275_), .B(new_n5281_), .ZN(new_n5316_));
  OAI21_X1   g05124(.A1(new_n5316_), .A2(new_n5280_), .B(\asqrt[37] ), .ZN(new_n5317_));
  INV_X1     g05125(.I(new_n5317_), .ZN(new_n5318_));
  NOR2_X1    g05126(.A1(new_n4960_), .A2(new_n5280_), .ZN(new_n5319_));
  NAND4_X1   g05127(.A1(new_n4949_), .A2(new_n4997_), .A3(new_n4998_), .A4(new_n5319_), .ZN(new_n5320_));
  NOR2_X1    g05128(.A1(new_n5316_), .A2(new_n5320_), .ZN(new_n5321_));
  AOI21_X1   g05129(.A1(new_n5315_), .A2(new_n5275_), .B(new_n4966_), .ZN(new_n5322_));
  INV_X1     g05130(.I(\a[73] ), .ZN(new_n5323_));
  AOI21_X1   g05131(.A1(\asqrt[36] ), .A2(new_n5281_), .B(new_n5323_), .ZN(new_n5324_));
  NOR3_X1    g05132(.A1(new_n5321_), .A2(new_n5324_), .A3(new_n5322_), .ZN(new_n5325_));
  OAI21_X1   g05133(.A1(new_n5325_), .A2(new_n5318_), .B(\asqrt[38] ), .ZN(new_n5326_));
  NOR2_X1    g05134(.A1(new_n5265_), .A2(\asqrt[63] ), .ZN(new_n5327_));
  INV_X1     g05135(.I(new_n5257_), .ZN(new_n5328_));
  INV_X1     g05136(.I(new_n5261_), .ZN(new_n5329_));
  NAND2_X1   g05137(.A1(new_n5244_), .A2(new_n5329_), .ZN(new_n5330_));
  INV_X1     g05138(.I(new_n5274_), .ZN(new_n5331_));
  OAI21_X1   g05139(.A1(new_n5328_), .A2(new_n5330_), .B(new_n5331_), .ZN(new_n5332_));
  OAI21_X1   g05140(.A1(new_n5327_), .A2(new_n5332_), .B(new_n4965_), .ZN(new_n5333_));
  NOR2_X1    g05141(.A1(new_n5328_), .A2(new_n5330_), .ZN(new_n5334_));
  OAI21_X1   g05142(.A1(new_n5272_), .A2(new_n4963_), .B(new_n4949_), .ZN(new_n5335_));
  NAND2_X1   g05143(.A1(new_n5270_), .A2(new_n5335_), .ZN(new_n5336_));
  NOR3_X1    g05144(.A1(new_n5327_), .A2(new_n5334_), .A3(new_n5336_), .ZN(new_n5337_));
  INV_X1     g05145(.I(new_n5337_), .ZN(new_n5338_));
  AOI21_X1   g05146(.A1(new_n5338_), .A2(new_n5333_), .B(new_n4985_), .ZN(new_n5339_));
  NOR3_X1    g05147(.A1(new_n5322_), .A2(new_n5337_), .A3(\a[74] ), .ZN(new_n5340_));
  AOI21_X1   g05148(.A1(\asqrt[36] ), .A2(\a[72] ), .B(new_n5280_), .ZN(new_n5341_));
  OAI21_X1   g05149(.A1(new_n5341_), .A2(new_n5024_), .B(new_n4696_), .ZN(new_n5342_));
  OAI22_X1   g05150(.A1(new_n5325_), .A2(new_n5342_), .B1(new_n5339_), .B2(new_n5340_), .ZN(new_n5343_));
  AOI21_X1   g05151(.A1(new_n5343_), .A2(new_n5326_), .B(new_n4298_), .ZN(new_n5344_));
  NOR3_X1    g05152(.A1(new_n5068_), .A2(new_n4984_), .A3(new_n4990_), .ZN(new_n5345_));
  NAND3_X1   g05153(.A1(\asqrt[36] ), .A2(new_n5006_), .A3(new_n5053_), .ZN(new_n5346_));
  AOI22_X1   g05154(.A1(new_n5346_), .A2(new_n5068_), .B1(\asqrt[36] ), .B2(new_n5345_), .ZN(new_n5347_));
  AOI21_X1   g05155(.A1(new_n5315_), .A2(new_n5275_), .B(\a[72] ), .ZN(new_n5348_));
  OAI21_X1   g05156(.A1(new_n5323_), .A2(new_n5348_), .B(new_n5333_), .ZN(new_n5349_));
  OAI21_X1   g05157(.A1(new_n5349_), .A2(new_n5321_), .B(new_n5317_), .ZN(new_n5350_));
  AOI21_X1   g05158(.A1(new_n5350_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n5351_));
  AOI21_X1   g05159(.A1(new_n5351_), .A2(new_n5343_), .B(new_n5347_), .ZN(new_n5352_));
  OAI21_X1   g05160(.A1(new_n5352_), .A2(new_n5344_), .B(\asqrt[40] ), .ZN(new_n5353_));
  INV_X1     g05161(.I(new_n5353_), .ZN(new_n5354_));
  NOR2_X1    g05162(.A1(new_n5005_), .A2(new_n5001_), .ZN(new_n5355_));
  INV_X1     g05163(.I(new_n5355_), .ZN(new_n5356_));
  NOR2_X1    g05164(.A1(new_n4994_), .A2(new_n5007_), .ZN(new_n5357_));
  NOR3_X1    g05165(.A1(new_n5057_), .A2(new_n5356_), .A3(new_n5357_), .ZN(new_n5358_));
  NOR3_X1    g05166(.A1(new_n5277_), .A2(new_n5057_), .A3(new_n5357_), .ZN(new_n5359_));
  INV_X1     g05167(.I(new_n5359_), .ZN(new_n5360_));
  AOI22_X1   g05168(.A1(new_n5360_), .A2(new_n5356_), .B1(\asqrt[36] ), .B2(new_n5358_), .ZN(new_n5361_));
  NOR3_X1    g05169(.A1(new_n5352_), .A2(new_n5344_), .A3(\asqrt[40] ), .ZN(new_n5362_));
  NOR2_X1    g05170(.A1(new_n5362_), .A2(new_n5361_), .ZN(new_n5363_));
  OAI21_X1   g05171(.A1(new_n5363_), .A2(new_n5354_), .B(\asqrt[41] ), .ZN(new_n5364_));
  NOR2_X1    g05172(.A1(new_n5070_), .A2(new_n5062_), .ZN(new_n5365_));
  NOR3_X1    g05173(.A1(new_n5277_), .A2(new_n5009_), .A3(new_n5365_), .ZN(new_n5366_));
  INV_X1     g05174(.I(new_n5366_), .ZN(new_n5367_));
  NOR3_X1    g05175(.A1(new_n5365_), .A2(new_n5009_), .A3(new_n5067_), .ZN(new_n5368_));
  AOI22_X1   g05176(.A1(new_n5367_), .A2(new_n5067_), .B1(\asqrt[36] ), .B2(new_n5368_), .ZN(new_n5369_));
  INV_X1     g05177(.I(new_n5369_), .ZN(new_n5370_));
  NAND2_X1   g05178(.A1(new_n5353_), .A2(new_n3782_), .ZN(new_n5371_));
  OAI21_X1   g05179(.A1(new_n5363_), .A2(new_n5371_), .B(new_n5370_), .ZN(new_n5372_));
  AOI21_X1   g05180(.A1(new_n5372_), .A2(new_n5364_), .B(new_n3419_), .ZN(new_n5373_));
  NOR3_X1    g05181(.A1(new_n5019_), .A2(new_n5028_), .A3(new_n5026_), .ZN(new_n5374_));
  NOR3_X1    g05182(.A1(new_n5277_), .A2(new_n5019_), .A3(new_n5028_), .ZN(new_n5375_));
  INV_X1     g05183(.I(new_n5375_), .ZN(new_n5376_));
  AOI22_X1   g05184(.A1(new_n5376_), .A2(new_n5026_), .B1(\asqrt[36] ), .B2(new_n5374_), .ZN(new_n5377_));
  OAI21_X1   g05185(.A1(new_n5361_), .A2(new_n5362_), .B(new_n5353_), .ZN(new_n5378_));
  AOI21_X1   g05186(.A1(new_n5378_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n5379_));
  AOI21_X1   g05187(.A1(new_n5379_), .A2(new_n5372_), .B(new_n5377_), .ZN(new_n5380_));
  OAI21_X1   g05188(.A1(new_n5380_), .A2(new_n5373_), .B(\asqrt[43] ), .ZN(new_n5381_));
  INV_X1     g05189(.I(new_n5381_), .ZN(new_n5382_));
  NOR2_X1    g05190(.A1(new_n5029_), .A2(new_n5037_), .ZN(new_n5383_));
  NOR3_X1    g05191(.A1(new_n5277_), .A2(new_n5066_), .A3(new_n5383_), .ZN(new_n5384_));
  INV_X1     g05192(.I(new_n5384_), .ZN(new_n5385_));
  NOR3_X1    g05193(.A1(new_n5383_), .A2(new_n5066_), .A3(new_n5036_), .ZN(new_n5386_));
  AOI22_X1   g05194(.A1(new_n5385_), .A2(new_n5036_), .B1(\asqrt[36] ), .B2(new_n5386_), .ZN(new_n5387_));
  NOR3_X1    g05195(.A1(new_n5380_), .A2(new_n5373_), .A3(\asqrt[43] ), .ZN(new_n5388_));
  NOR2_X1    g05196(.A1(new_n5388_), .A2(new_n5387_), .ZN(new_n5389_));
  OAI21_X1   g05197(.A1(new_n5389_), .A2(new_n5382_), .B(\asqrt[44] ), .ZN(new_n5390_));
  INV_X1     g05198(.I(new_n5043_), .ZN(new_n5391_));
  NOR3_X1    g05199(.A1(new_n5039_), .A2(new_n5084_), .A3(new_n5391_), .ZN(new_n5392_));
  NOR3_X1    g05200(.A1(new_n5277_), .A2(new_n5039_), .A3(new_n5084_), .ZN(new_n5393_));
  INV_X1     g05201(.I(new_n5393_), .ZN(new_n5394_));
  AOI22_X1   g05202(.A1(new_n5394_), .A2(new_n5391_), .B1(\asqrt[36] ), .B2(new_n5392_), .ZN(new_n5395_));
  INV_X1     g05203(.I(new_n5395_), .ZN(new_n5396_));
  NAND2_X1   g05204(.A1(new_n5381_), .A2(new_n2954_), .ZN(new_n5397_));
  OAI21_X1   g05205(.A1(new_n5389_), .A2(new_n5397_), .B(new_n5396_), .ZN(new_n5398_));
  AOI21_X1   g05206(.A1(new_n5398_), .A2(new_n5390_), .B(new_n2641_), .ZN(new_n5399_));
  NOR3_X1    g05207(.A1(new_n5277_), .A2(new_n5288_), .A3(new_n5111_), .ZN(new_n5400_));
  INV_X1     g05208(.I(new_n5400_), .ZN(new_n5401_));
  NOR3_X1    g05209(.A1(new_n5288_), .A2(new_n5052_), .A3(new_n5111_), .ZN(new_n5402_));
  AOI22_X1   g05210(.A1(new_n5401_), .A2(new_n5052_), .B1(\asqrt[36] ), .B2(new_n5402_), .ZN(new_n5403_));
  OAI21_X1   g05211(.A1(new_n5387_), .A2(new_n5388_), .B(new_n5381_), .ZN(new_n5404_));
  AOI21_X1   g05212(.A1(new_n5404_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n5405_));
  AOI21_X1   g05213(.A1(new_n5405_), .A2(new_n5398_), .B(new_n5403_), .ZN(new_n5406_));
  OAI21_X1   g05214(.A1(new_n5406_), .A2(new_n5399_), .B(\asqrt[46] ), .ZN(new_n5407_));
  INV_X1     g05215(.I(new_n5407_), .ZN(new_n5408_));
  INV_X1     g05216(.I(new_n5114_), .ZN(new_n5409_));
  NOR3_X1    g05217(.A1(new_n5409_), .A2(new_n5078_), .A3(new_n5113_), .ZN(new_n5410_));
  NOR3_X1    g05218(.A1(new_n5277_), .A2(new_n5078_), .A3(new_n5409_), .ZN(new_n5411_));
  INV_X1     g05219(.I(new_n5411_), .ZN(new_n5412_));
  AOI22_X1   g05220(.A1(new_n5412_), .A2(new_n5113_), .B1(\asqrt[36] ), .B2(new_n5410_), .ZN(new_n5413_));
  NOR3_X1    g05221(.A1(new_n5406_), .A2(new_n5399_), .A3(\asqrt[46] ), .ZN(new_n5414_));
  NOR2_X1    g05222(.A1(new_n5414_), .A2(new_n5413_), .ZN(new_n5415_));
  OAI21_X1   g05223(.A1(new_n5415_), .A2(new_n5408_), .B(\asqrt[47] ), .ZN(new_n5416_));
  NOR3_X1    g05224(.A1(new_n5277_), .A2(new_n5089_), .A3(new_n5094_), .ZN(new_n5417_));
  INV_X1     g05225(.I(new_n5417_), .ZN(new_n5418_));
  NOR3_X1    g05226(.A1(new_n5089_), .A2(new_n5094_), .A3(new_n5287_), .ZN(new_n5419_));
  AOI22_X1   g05227(.A1(new_n5418_), .A2(new_n5287_), .B1(\asqrt[36] ), .B2(new_n5419_), .ZN(new_n5420_));
  INV_X1     g05228(.I(new_n5420_), .ZN(new_n5421_));
  NAND2_X1   g05229(.A1(new_n5407_), .A2(new_n2229_), .ZN(new_n5422_));
  OAI21_X1   g05230(.A1(new_n5415_), .A2(new_n5422_), .B(new_n5421_), .ZN(new_n5423_));
  AOI21_X1   g05231(.A1(new_n5423_), .A2(new_n5416_), .B(new_n1956_), .ZN(new_n5424_));
  INV_X1     g05232(.I(new_n5096_), .ZN(new_n5425_));
  NOR2_X1    g05233(.A1(new_n5095_), .A2(new_n5103_), .ZN(new_n5426_));
  NOR3_X1    g05234(.A1(new_n5425_), .A2(new_n5102_), .A3(new_n5426_), .ZN(new_n5427_));
  NOR3_X1    g05235(.A1(new_n5277_), .A2(new_n5425_), .A3(new_n5426_), .ZN(new_n5428_));
  INV_X1     g05236(.I(new_n5428_), .ZN(new_n5429_));
  AOI22_X1   g05237(.A1(new_n5429_), .A2(new_n5102_), .B1(\asqrt[36] ), .B2(new_n5427_), .ZN(new_n5430_));
  OAI21_X1   g05238(.A1(new_n5413_), .A2(new_n5414_), .B(new_n5407_), .ZN(new_n5431_));
  AOI21_X1   g05239(.A1(new_n5431_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n5432_));
  AOI21_X1   g05240(.A1(new_n5432_), .A2(new_n5423_), .B(new_n5430_), .ZN(new_n5433_));
  OAI21_X1   g05241(.A1(new_n5433_), .A2(new_n5424_), .B(\asqrt[49] ), .ZN(new_n5434_));
  INV_X1     g05242(.I(new_n5434_), .ZN(new_n5435_));
  INV_X1     g05243(.I(new_n5110_), .ZN(new_n5436_));
  INV_X1     g05244(.I(new_n5104_), .ZN(new_n5437_));
  INV_X1     g05245(.I(new_n5117_), .ZN(new_n5438_));
  NOR2_X1    g05246(.A1(new_n5438_), .A2(new_n5437_), .ZN(new_n5439_));
  NOR3_X1    g05247(.A1(new_n5277_), .A2(new_n5105_), .A3(new_n5439_), .ZN(new_n5440_));
  INV_X1     g05248(.I(new_n5440_), .ZN(new_n5441_));
  NOR3_X1    g05249(.A1(new_n5439_), .A2(new_n5105_), .A3(new_n5436_), .ZN(new_n5442_));
  AOI22_X1   g05250(.A1(new_n5441_), .A2(new_n5436_), .B1(\asqrt[36] ), .B2(new_n5442_), .ZN(new_n5443_));
  NOR3_X1    g05251(.A1(new_n5433_), .A2(new_n5424_), .A3(\asqrt[49] ), .ZN(new_n5444_));
  NOR2_X1    g05252(.A1(new_n5444_), .A2(new_n5443_), .ZN(new_n5445_));
  OAI21_X1   g05253(.A1(new_n5445_), .A2(new_n5435_), .B(\asqrt[50] ), .ZN(new_n5446_));
  NOR3_X1    g05254(.A1(new_n5120_), .A2(new_n5286_), .A3(new_n5125_), .ZN(new_n5447_));
  NOR3_X1    g05255(.A1(new_n5277_), .A2(new_n5120_), .A3(new_n5125_), .ZN(new_n5448_));
  INV_X1     g05256(.I(new_n5448_), .ZN(new_n5449_));
  AOI22_X1   g05257(.A1(new_n5449_), .A2(new_n5286_), .B1(\asqrt[36] ), .B2(new_n5447_), .ZN(new_n5450_));
  INV_X1     g05258(.I(new_n5450_), .ZN(new_n5451_));
  NAND2_X1   g05259(.A1(new_n5434_), .A2(new_n1612_), .ZN(new_n5452_));
  OAI21_X1   g05260(.A1(new_n5445_), .A2(new_n5452_), .B(new_n5451_), .ZN(new_n5453_));
  AOI21_X1   g05261(.A1(new_n5453_), .A2(new_n5446_), .B(new_n1376_), .ZN(new_n5454_));
  INV_X1     g05262(.I(new_n5127_), .ZN(new_n5455_));
  NOR2_X1    g05263(.A1(new_n5126_), .A2(new_n5134_), .ZN(new_n5456_));
  NOR3_X1    g05264(.A1(new_n5277_), .A2(new_n5455_), .A3(new_n5456_), .ZN(new_n5457_));
  INV_X1     g05265(.I(new_n5457_), .ZN(new_n5458_));
  NOR3_X1    g05266(.A1(new_n5455_), .A2(new_n5133_), .A3(new_n5456_), .ZN(new_n5459_));
  AOI22_X1   g05267(.A1(new_n5458_), .A2(new_n5133_), .B1(\asqrt[36] ), .B2(new_n5459_), .ZN(new_n5460_));
  OAI21_X1   g05268(.A1(new_n5443_), .A2(new_n5444_), .B(new_n5434_), .ZN(new_n5461_));
  AOI21_X1   g05269(.A1(new_n5461_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n5462_));
  AOI21_X1   g05270(.A1(new_n5462_), .A2(new_n5453_), .B(new_n5460_), .ZN(new_n5463_));
  OAI21_X1   g05271(.A1(new_n5463_), .A2(new_n5454_), .B(\asqrt[52] ), .ZN(new_n5464_));
  INV_X1     g05272(.I(new_n5141_), .ZN(new_n5465_));
  INV_X1     g05273(.I(new_n5135_), .ZN(new_n5466_));
  INV_X1     g05274(.I(new_n5143_), .ZN(new_n5467_));
  NOR2_X1    g05275(.A1(new_n5467_), .A2(new_n5466_), .ZN(new_n5468_));
  NOR3_X1    g05276(.A1(new_n5468_), .A2(new_n5136_), .A3(new_n5465_), .ZN(new_n5469_));
  NOR3_X1    g05277(.A1(new_n5277_), .A2(new_n5136_), .A3(new_n5468_), .ZN(new_n5470_));
  INV_X1     g05278(.I(new_n5470_), .ZN(new_n5471_));
  AOI22_X1   g05279(.A1(new_n5471_), .A2(new_n5465_), .B1(\asqrt[36] ), .B2(new_n5469_), .ZN(new_n5472_));
  INV_X1     g05280(.I(new_n5472_), .ZN(new_n5473_));
  INV_X1     g05281(.I(new_n5443_), .ZN(new_n5474_));
  OR2_X2     g05282(.A1(new_n5424_), .A2(\asqrt[49] ), .Z(new_n5475_));
  OAI21_X1   g05283(.A1(new_n5475_), .A2(new_n5433_), .B(new_n5474_), .ZN(new_n5476_));
  AOI21_X1   g05284(.A1(new_n5476_), .A2(new_n5434_), .B(new_n1612_), .ZN(new_n5477_));
  INV_X1     g05285(.I(new_n5452_), .ZN(new_n5478_));
  AOI21_X1   g05286(.A1(new_n5478_), .A2(new_n5476_), .B(new_n5450_), .ZN(new_n5479_));
  OAI21_X1   g05287(.A1(new_n5479_), .A2(new_n5477_), .B(\asqrt[51] ), .ZN(new_n5480_));
  NAND2_X1   g05288(.A1(new_n5480_), .A2(new_n1256_), .ZN(new_n5481_));
  OAI21_X1   g05289(.A1(new_n5481_), .A2(new_n5463_), .B(new_n5473_), .ZN(new_n5482_));
  AOI21_X1   g05290(.A1(new_n5482_), .A2(new_n5464_), .B(new_n1103_), .ZN(new_n5483_));
  NOR3_X1    g05291(.A1(new_n5277_), .A2(new_n5146_), .A3(new_n5188_), .ZN(new_n5484_));
  INV_X1     g05292(.I(new_n5484_), .ZN(new_n5485_));
  NOR3_X1    g05293(.A1(new_n5146_), .A2(new_n5285_), .A3(new_n5188_), .ZN(new_n5486_));
  AOI22_X1   g05294(.A1(new_n5485_), .A2(new_n5285_), .B1(\asqrt[36] ), .B2(new_n5486_), .ZN(new_n5487_));
  INV_X1     g05295(.I(new_n5460_), .ZN(new_n5488_));
  NAND2_X1   g05296(.A1(new_n5446_), .A2(new_n1376_), .ZN(new_n5489_));
  OAI21_X1   g05297(.A1(new_n5489_), .A2(new_n5479_), .B(new_n5488_), .ZN(new_n5490_));
  AOI21_X1   g05298(.A1(new_n5490_), .A2(new_n5480_), .B(new_n1256_), .ZN(new_n5491_));
  NOR2_X1    g05299(.A1(new_n5491_), .A2(\asqrt[53] ), .ZN(new_n5492_));
  AOI21_X1   g05300(.A1(new_n5492_), .A2(new_n5482_), .B(new_n5487_), .ZN(new_n5493_));
  OAI21_X1   g05301(.A1(new_n5493_), .A2(new_n5483_), .B(\asqrt[54] ), .ZN(new_n5494_));
  INV_X1     g05302(.I(new_n5154_), .ZN(new_n5495_));
  NOR2_X1    g05303(.A1(new_n5161_), .A2(new_n5153_), .ZN(new_n5496_));
  NOR3_X1    g05304(.A1(new_n5495_), .A2(new_n5160_), .A3(new_n5496_), .ZN(new_n5497_));
  NOR3_X1    g05305(.A1(new_n5277_), .A2(new_n5495_), .A3(new_n5496_), .ZN(new_n5498_));
  INV_X1     g05306(.I(new_n5498_), .ZN(new_n5499_));
  AOI22_X1   g05307(.A1(new_n5499_), .A2(new_n5160_), .B1(\asqrt[36] ), .B2(new_n5497_), .ZN(new_n5500_));
  INV_X1     g05308(.I(new_n5500_), .ZN(new_n5501_));
  NOR2_X1    g05309(.A1(new_n5454_), .A2(\asqrt[52] ), .ZN(new_n5502_));
  AOI21_X1   g05310(.A1(new_n5502_), .A2(new_n5490_), .B(new_n5472_), .ZN(new_n5503_));
  OAI21_X1   g05311(.A1(new_n5503_), .A2(new_n5491_), .B(\asqrt[53] ), .ZN(new_n5504_));
  NAND2_X1   g05312(.A1(new_n5504_), .A2(new_n904_), .ZN(new_n5505_));
  OAI21_X1   g05313(.A1(new_n5505_), .A2(new_n5493_), .B(new_n5501_), .ZN(new_n5506_));
  AOI21_X1   g05314(.A1(new_n5506_), .A2(new_n5494_), .B(new_n823_), .ZN(new_n5507_));
  NOR2_X1    g05315(.A1(new_n5172_), .A2(new_n5165_), .ZN(new_n5508_));
  NOR3_X1    g05316(.A1(new_n5277_), .A2(new_n5163_), .A3(new_n5508_), .ZN(new_n5509_));
  INV_X1     g05317(.I(new_n5509_), .ZN(new_n5510_));
  NOR3_X1    g05318(.A1(new_n5508_), .A2(new_n5163_), .A3(new_n5171_), .ZN(new_n5511_));
  AOI22_X1   g05319(.A1(new_n5510_), .A2(new_n5171_), .B1(\asqrt[36] ), .B2(new_n5511_), .ZN(new_n5512_));
  INV_X1     g05320(.I(new_n5487_), .ZN(new_n5513_));
  NAND2_X1   g05321(.A1(new_n5464_), .A2(new_n1103_), .ZN(new_n5514_));
  OAI21_X1   g05322(.A1(new_n5514_), .A2(new_n5503_), .B(new_n5513_), .ZN(new_n5515_));
  AOI21_X1   g05323(.A1(new_n5515_), .A2(new_n5504_), .B(new_n904_), .ZN(new_n5516_));
  NOR2_X1    g05324(.A1(new_n5516_), .A2(\asqrt[55] ), .ZN(new_n5517_));
  AOI21_X1   g05325(.A1(new_n5517_), .A2(new_n5506_), .B(new_n5512_), .ZN(new_n5518_));
  OAI21_X1   g05326(.A1(new_n5518_), .A2(new_n5507_), .B(\asqrt[56] ), .ZN(new_n5519_));
  NOR3_X1    g05327(.A1(new_n5174_), .A2(new_n5284_), .A3(new_n5220_), .ZN(new_n5520_));
  NOR3_X1    g05328(.A1(new_n5277_), .A2(new_n5174_), .A3(new_n5220_), .ZN(new_n5521_));
  INV_X1     g05329(.I(new_n5521_), .ZN(new_n5522_));
  AOI22_X1   g05330(.A1(new_n5522_), .A2(new_n5284_), .B1(\asqrt[36] ), .B2(new_n5520_), .ZN(new_n5523_));
  INV_X1     g05331(.I(new_n5523_), .ZN(new_n5524_));
  NOR3_X1    g05332(.A1(new_n5463_), .A2(new_n5454_), .A3(\asqrt[52] ), .ZN(new_n5525_));
  OAI21_X1   g05333(.A1(new_n5472_), .A2(new_n5525_), .B(new_n5464_), .ZN(new_n5526_));
  AOI21_X1   g05334(.A1(new_n5526_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n5527_));
  AOI21_X1   g05335(.A1(new_n5527_), .A2(new_n5515_), .B(new_n5500_), .ZN(new_n5528_));
  OAI21_X1   g05336(.A1(new_n5528_), .A2(new_n5516_), .B(\asqrt[55] ), .ZN(new_n5529_));
  NAND2_X1   g05337(.A1(new_n5529_), .A2(new_n703_), .ZN(new_n5530_));
  OAI21_X1   g05338(.A1(new_n5530_), .A2(new_n5518_), .B(new_n5524_), .ZN(new_n5531_));
  AOI21_X1   g05339(.A1(new_n5531_), .A2(new_n5519_), .B(new_n531_), .ZN(new_n5532_));
  INV_X1     g05340(.I(new_n5181_), .ZN(new_n5533_));
  NOR2_X1    g05341(.A1(new_n5193_), .A2(new_n5180_), .ZN(new_n5534_));
  NOR3_X1    g05342(.A1(new_n5277_), .A2(new_n5533_), .A3(new_n5534_), .ZN(new_n5535_));
  INV_X1     g05343(.I(new_n5535_), .ZN(new_n5536_));
  NOR3_X1    g05344(.A1(new_n5533_), .A2(new_n5187_), .A3(new_n5534_), .ZN(new_n5537_));
  AOI22_X1   g05345(.A1(new_n5536_), .A2(new_n5187_), .B1(\asqrt[36] ), .B2(new_n5537_), .ZN(new_n5538_));
  NOR3_X1    g05346(.A1(new_n5528_), .A2(\asqrt[55] ), .A3(new_n5516_), .ZN(new_n5539_));
  OAI21_X1   g05347(.A1(new_n5512_), .A2(new_n5539_), .B(new_n5529_), .ZN(new_n5540_));
  AOI21_X1   g05348(.A1(new_n5540_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n5541_));
  AOI21_X1   g05349(.A1(new_n5541_), .A2(new_n5531_), .B(new_n5538_), .ZN(new_n5542_));
  OAI21_X1   g05350(.A1(new_n5542_), .A2(new_n5532_), .B(\asqrt[58] ), .ZN(new_n5543_));
  NOR2_X1    g05351(.A1(new_n5204_), .A2(new_n5197_), .ZN(new_n5544_));
  NOR3_X1    g05352(.A1(new_n5544_), .A2(new_n5195_), .A3(new_n5203_), .ZN(new_n5545_));
  NOR3_X1    g05353(.A1(new_n5277_), .A2(new_n5195_), .A3(new_n5544_), .ZN(new_n5546_));
  INV_X1     g05354(.I(new_n5546_), .ZN(new_n5547_));
  AOI22_X1   g05355(.A1(new_n5547_), .A2(new_n5203_), .B1(\asqrt[36] ), .B2(new_n5545_), .ZN(new_n5548_));
  INV_X1     g05356(.I(new_n5548_), .ZN(new_n5549_));
  INV_X1     g05357(.I(new_n5512_), .ZN(new_n5550_));
  NAND2_X1   g05358(.A1(new_n5494_), .A2(new_n823_), .ZN(new_n5551_));
  OAI21_X1   g05359(.A1(new_n5551_), .A2(new_n5528_), .B(new_n5550_), .ZN(new_n5552_));
  AOI21_X1   g05360(.A1(new_n5552_), .A2(new_n5529_), .B(new_n703_), .ZN(new_n5553_));
  NOR2_X1    g05361(.A1(new_n5507_), .A2(\asqrt[56] ), .ZN(new_n5554_));
  AOI21_X1   g05362(.A1(new_n5554_), .A2(new_n5552_), .B(new_n5523_), .ZN(new_n5555_));
  OAI21_X1   g05363(.A1(new_n5555_), .A2(new_n5553_), .B(\asqrt[57] ), .ZN(new_n5556_));
  NAND2_X1   g05364(.A1(new_n5556_), .A2(new_n436_), .ZN(new_n5557_));
  OAI21_X1   g05365(.A1(new_n5557_), .A2(new_n5542_), .B(new_n5549_), .ZN(new_n5558_));
  AOI21_X1   g05366(.A1(new_n5558_), .A2(new_n5543_), .B(new_n327_), .ZN(new_n5559_));
  NOR3_X1    g05367(.A1(new_n5277_), .A2(new_n5206_), .A3(new_n5251_), .ZN(new_n5560_));
  INV_X1     g05368(.I(new_n5560_), .ZN(new_n5561_));
  NOR3_X1    g05369(.A1(new_n5206_), .A2(new_n5283_), .A3(new_n5251_), .ZN(new_n5562_));
  AOI22_X1   g05370(.A1(new_n5561_), .A2(new_n5283_), .B1(\asqrt[36] ), .B2(new_n5562_), .ZN(new_n5563_));
  INV_X1     g05371(.I(new_n5538_), .ZN(new_n5564_));
  NAND2_X1   g05372(.A1(new_n5519_), .A2(new_n531_), .ZN(new_n5565_));
  OAI21_X1   g05373(.A1(new_n5565_), .A2(new_n5555_), .B(new_n5564_), .ZN(new_n5566_));
  AOI21_X1   g05374(.A1(new_n5566_), .A2(new_n5556_), .B(new_n436_), .ZN(new_n5567_));
  NOR2_X1    g05375(.A1(new_n5567_), .A2(\asqrt[59] ), .ZN(new_n5568_));
  AOI21_X1   g05376(.A1(new_n5568_), .A2(new_n5558_), .B(new_n5563_), .ZN(new_n5569_));
  OAI21_X1   g05377(.A1(new_n5569_), .A2(new_n5559_), .B(\asqrt[60] ), .ZN(new_n5570_));
  INV_X1     g05378(.I(new_n5213_), .ZN(new_n5571_));
  NOR2_X1    g05379(.A1(new_n5225_), .A2(new_n5212_), .ZN(new_n5572_));
  NOR3_X1    g05380(.A1(new_n5571_), .A2(new_n5219_), .A3(new_n5572_), .ZN(new_n5573_));
  NOR3_X1    g05381(.A1(new_n5277_), .A2(new_n5571_), .A3(new_n5572_), .ZN(new_n5574_));
  INV_X1     g05382(.I(new_n5574_), .ZN(new_n5575_));
  AOI22_X1   g05383(.A1(new_n5575_), .A2(new_n5219_), .B1(\asqrt[36] ), .B2(new_n5573_), .ZN(new_n5576_));
  INV_X1     g05384(.I(new_n5576_), .ZN(new_n5577_));
  NOR2_X1    g05385(.A1(new_n5532_), .A2(\asqrt[58] ), .ZN(new_n5578_));
  AOI21_X1   g05386(.A1(new_n5578_), .A2(new_n5566_), .B(new_n5548_), .ZN(new_n5579_));
  OAI21_X1   g05387(.A1(new_n5579_), .A2(new_n5567_), .B(\asqrt[59] ), .ZN(new_n5580_));
  NAND2_X1   g05388(.A1(new_n5580_), .A2(new_n306_), .ZN(new_n5581_));
  OAI21_X1   g05389(.A1(new_n5581_), .A2(new_n5569_), .B(new_n5577_), .ZN(new_n5582_));
  AOI21_X1   g05390(.A1(new_n5582_), .A2(new_n5570_), .B(new_n218_), .ZN(new_n5583_));
  NOR2_X1    g05391(.A1(new_n5229_), .A2(new_n5235_), .ZN(new_n5584_));
  NOR3_X1    g05392(.A1(new_n5277_), .A2(new_n5227_), .A3(new_n5584_), .ZN(new_n5585_));
  INV_X1     g05393(.I(new_n5585_), .ZN(new_n5586_));
  NOR3_X1    g05394(.A1(new_n5584_), .A2(new_n5227_), .A3(new_n5234_), .ZN(new_n5587_));
  AOI22_X1   g05395(.A1(new_n5586_), .A2(new_n5234_), .B1(\asqrt[36] ), .B2(new_n5587_), .ZN(new_n5588_));
  INV_X1     g05396(.I(new_n5563_), .ZN(new_n5589_));
  NAND2_X1   g05397(.A1(new_n5543_), .A2(new_n327_), .ZN(new_n5590_));
  OAI21_X1   g05398(.A1(new_n5590_), .A2(new_n5579_), .B(new_n5589_), .ZN(new_n5591_));
  AOI21_X1   g05399(.A1(new_n5591_), .A2(new_n5580_), .B(new_n306_), .ZN(new_n5592_));
  NOR2_X1    g05400(.A1(new_n5592_), .A2(\asqrt[61] ), .ZN(new_n5593_));
  AOI21_X1   g05401(.A1(new_n5593_), .A2(new_n5582_), .B(new_n5588_), .ZN(new_n5594_));
  OAI21_X1   g05402(.A1(new_n5594_), .A2(new_n5583_), .B(\asqrt[62] ), .ZN(new_n5595_));
  NOR3_X1    g05403(.A1(new_n5237_), .A2(new_n5282_), .A3(new_n5266_), .ZN(new_n5596_));
  NOR3_X1    g05404(.A1(new_n5277_), .A2(new_n5237_), .A3(new_n5266_), .ZN(new_n5597_));
  INV_X1     g05405(.I(new_n5597_), .ZN(new_n5598_));
  AOI22_X1   g05406(.A1(new_n5598_), .A2(new_n5282_), .B1(\asqrt[36] ), .B2(new_n5596_), .ZN(new_n5599_));
  INV_X1     g05407(.I(new_n5599_), .ZN(new_n5600_));
  NOR3_X1    g05408(.A1(new_n5542_), .A2(\asqrt[58] ), .A3(new_n5532_), .ZN(new_n5601_));
  OAI21_X1   g05409(.A1(new_n5548_), .A2(new_n5601_), .B(new_n5543_), .ZN(new_n5602_));
  AOI21_X1   g05410(.A1(new_n5602_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n5603_));
  AOI21_X1   g05411(.A1(new_n5603_), .A2(new_n5591_), .B(new_n5576_), .ZN(new_n5604_));
  OAI21_X1   g05412(.A1(new_n5604_), .A2(new_n5592_), .B(\asqrt[61] ), .ZN(new_n5605_));
  NAND2_X1   g05413(.A1(new_n5605_), .A2(new_n207_), .ZN(new_n5606_));
  OAI21_X1   g05414(.A1(new_n5606_), .A2(new_n5594_), .B(new_n5600_), .ZN(new_n5607_));
  INV_X1     g05415(.I(new_n5334_), .ZN(new_n5608_));
  NAND4_X1   g05416(.A1(\asqrt[36] ), .A2(new_n5244_), .A3(new_n5249_), .A4(new_n5313_), .ZN(new_n5609_));
  NAND2_X1   g05417(.A1(new_n5244_), .A2(new_n5313_), .ZN(new_n5610_));
  OAI21_X1   g05418(.A1(new_n5277_), .A2(new_n5610_), .B(new_n5250_), .ZN(new_n5611_));
  NAND2_X1   g05419(.A1(new_n5611_), .A2(new_n5609_), .ZN(new_n5612_));
  NOR2_X1    g05420(.A1(new_n5314_), .A2(new_n5329_), .ZN(new_n5613_));
  NAND2_X1   g05421(.A1(\asqrt[36] ), .A2(new_n5613_), .ZN(new_n5614_));
  NAND3_X1   g05422(.A1(new_n5612_), .A2(new_n5608_), .A3(new_n5614_), .ZN(new_n5615_));
  AOI21_X1   g05423(.A1(new_n5607_), .A2(new_n5595_), .B(new_n5615_), .ZN(new_n5616_));
  NOR3_X1    g05424(.A1(new_n5604_), .A2(\asqrt[61] ), .A3(new_n5592_), .ZN(new_n5617_));
  OAI21_X1   g05425(.A1(new_n5588_), .A2(new_n5617_), .B(new_n5605_), .ZN(new_n5618_));
  AOI21_X1   g05426(.A1(new_n5618_), .A2(\asqrt[62] ), .B(new_n5612_), .ZN(new_n5619_));
  OAI21_X1   g05427(.A1(new_n5277_), .A2(new_n5329_), .B(new_n5314_), .ZN(new_n5620_));
  NOR2_X1    g05428(.A1(new_n5613_), .A2(new_n193_), .ZN(new_n5621_));
  NAND2_X1   g05429(.A1(new_n5620_), .A2(new_n5621_), .ZN(new_n5622_));
  INV_X1     g05430(.I(new_n5622_), .ZN(new_n5623_));
  AND3_X2    g05431(.A1(new_n5260_), .A2(new_n5258_), .A3(new_n5273_), .Z(new_n5624_));
  NAND4_X1   g05432(.A1(new_n5608_), .A2(new_n5315_), .A3(new_n5270_), .A4(new_n5624_), .ZN(new_n5625_));
  INV_X1     g05433(.I(new_n5625_), .ZN(new_n5626_));
  NOR2_X1    g05434(.A1(new_n5623_), .A2(new_n5626_), .ZN(new_n5627_));
  INV_X1     g05435(.I(new_n5627_), .ZN(new_n5628_));
  AOI21_X1   g05436(.A1(new_n5619_), .A2(new_n5607_), .B(new_n5628_), .ZN(new_n5629_));
  OAI21_X1   g05437(.A1(\asqrt[63] ), .A2(new_n5616_), .B(new_n5629_), .ZN(\asqrt[35] ));
  NOR2_X1    g05438(.A1(\a[68] ), .A2(\a[69] ), .ZN(new_n5631_));
  INV_X1     g05439(.I(new_n5631_), .ZN(new_n5632_));
  NOR2_X1    g05440(.A1(new_n5632_), .A2(\a[70] ), .ZN(new_n5633_));
  INV_X1     g05441(.I(new_n5633_), .ZN(new_n5634_));
  NAND2_X1   g05442(.A1(new_n5607_), .A2(new_n5595_), .ZN(new_n5635_));
  INV_X1     g05443(.I(new_n5615_), .ZN(new_n5636_));
  AOI21_X1   g05444(.A1(new_n5635_), .A2(new_n5636_), .B(\asqrt[63] ), .ZN(new_n5637_));
  INV_X1     g05445(.I(new_n5607_), .ZN(new_n5638_));
  INV_X1     g05446(.I(new_n5612_), .ZN(new_n5639_));
  NAND2_X1   g05447(.A1(new_n5595_), .A2(new_n5639_), .ZN(new_n5640_));
  OAI21_X1   g05448(.A1(new_n5638_), .A2(new_n5640_), .B(new_n5627_), .ZN(new_n5641_));
  OAI21_X1   g05449(.A1(new_n5637_), .A2(new_n5641_), .B(\a[70] ), .ZN(new_n5642_));
  AOI21_X1   g05450(.A1(new_n5642_), .A2(new_n5634_), .B(new_n5277_), .ZN(new_n5643_));
  INV_X1     g05451(.I(\a[70] ), .ZN(new_n5644_));
  INV_X1     g05452(.I(new_n5588_), .ZN(new_n5645_));
  NAND2_X1   g05453(.A1(new_n5570_), .A2(new_n218_), .ZN(new_n5646_));
  OAI21_X1   g05454(.A1(new_n5646_), .A2(new_n5604_), .B(new_n5645_), .ZN(new_n5647_));
  NAND3_X1   g05455(.A1(new_n5647_), .A2(new_n207_), .A3(new_n5605_), .ZN(new_n5648_));
  AOI22_X1   g05456(.A1(new_n5648_), .A2(new_n5600_), .B1(new_n5618_), .B2(\asqrt[62] ), .ZN(new_n5649_));
  OAI21_X1   g05457(.A1(new_n5649_), .A2(new_n5615_), .B(new_n193_), .ZN(new_n5650_));
  AOI21_X1   g05458(.A1(new_n5650_), .A2(new_n5629_), .B(new_n5644_), .ZN(new_n5651_));
  NAND4_X1   g05459(.A1(new_n5608_), .A2(new_n5270_), .A3(new_n5273_), .A4(new_n5634_), .ZN(new_n5652_));
  NOR2_X1    g05460(.A1(new_n5652_), .A2(new_n5327_), .ZN(new_n5653_));
  INV_X1     g05461(.I(new_n5653_), .ZN(new_n5654_));
  NOR2_X1    g05462(.A1(new_n5651_), .A2(new_n5654_), .ZN(new_n5655_));
  AOI21_X1   g05463(.A1(new_n5650_), .A2(new_n5629_), .B(new_n5279_), .ZN(new_n5656_));
  INV_X1     g05464(.I(\a[71] ), .ZN(new_n5657_));
  AOI21_X1   g05465(.A1(\asqrt[35] ), .A2(new_n5644_), .B(new_n5657_), .ZN(new_n5658_));
  NOR3_X1    g05466(.A1(new_n5655_), .A2(new_n5658_), .A3(new_n5656_), .ZN(new_n5659_));
  OAI21_X1   g05467(.A1(new_n5659_), .A2(new_n5643_), .B(\asqrt[37] ), .ZN(new_n5660_));
  OAI21_X1   g05468(.A1(new_n5637_), .A2(new_n5641_), .B(new_n5278_), .ZN(new_n5661_));
  NOR2_X1    g05469(.A1(new_n5638_), .A2(new_n5640_), .ZN(new_n5662_));
  NOR2_X1    g05470(.A1(new_n5626_), .A2(new_n5277_), .ZN(new_n5663_));
  NAND2_X1   g05471(.A1(new_n5622_), .A2(new_n5663_), .ZN(new_n5664_));
  NOR3_X1    g05472(.A1(new_n5637_), .A2(new_n5662_), .A3(new_n5664_), .ZN(new_n5665_));
  INV_X1     g05473(.I(new_n5665_), .ZN(new_n5666_));
  AOI21_X1   g05474(.A1(new_n5666_), .A2(new_n5661_), .B(new_n5281_), .ZN(new_n5667_));
  NOR3_X1    g05475(.A1(new_n5665_), .A2(new_n5656_), .A3(\a[72] ), .ZN(new_n5668_));
  AOI21_X1   g05476(.A1(\asqrt[35] ), .A2(\a[70] ), .B(new_n5633_), .ZN(new_n5669_));
  OAI21_X1   g05477(.A1(new_n5669_), .A2(new_n5277_), .B(new_n5024_), .ZN(new_n5670_));
  OAI22_X1   g05478(.A1(new_n5659_), .A2(new_n5670_), .B1(new_n5667_), .B2(new_n5668_), .ZN(new_n5671_));
  AOI21_X1   g05479(.A1(new_n5671_), .A2(new_n5660_), .B(new_n4696_), .ZN(new_n5672_));
  INV_X1     g05480(.I(new_n5349_), .ZN(new_n5673_));
  NOR3_X1    g05481(.A1(new_n5318_), .A2(new_n5673_), .A3(new_n5321_), .ZN(new_n5674_));
  NOR2_X1    g05482(.A1(new_n5318_), .A2(new_n5321_), .ZN(new_n5675_));
  NAND2_X1   g05483(.A1(\asqrt[35] ), .A2(new_n5675_), .ZN(new_n5676_));
  AOI22_X1   g05484(.A1(new_n5676_), .A2(new_n5673_), .B1(\asqrt[35] ), .B2(new_n5674_), .ZN(new_n5677_));
  OAI21_X1   g05485(.A1(new_n5651_), .A2(new_n5633_), .B(\asqrt[36] ), .ZN(new_n5678_));
  AOI21_X1   g05486(.A1(new_n5650_), .A2(new_n5629_), .B(\a[70] ), .ZN(new_n5679_));
  OAI21_X1   g05487(.A1(new_n5657_), .A2(new_n5679_), .B(new_n5661_), .ZN(new_n5680_));
  OAI21_X1   g05488(.A1(new_n5680_), .A2(new_n5655_), .B(new_n5678_), .ZN(new_n5681_));
  AOI21_X1   g05489(.A1(new_n5681_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n5682_));
  AOI21_X1   g05490(.A1(new_n5682_), .A2(new_n5671_), .B(new_n5677_), .ZN(new_n5683_));
  OAI21_X1   g05491(.A1(new_n5683_), .A2(new_n5672_), .B(\asqrt[39] ), .ZN(new_n5684_));
  INV_X1     g05492(.I(new_n5684_), .ZN(new_n5685_));
  NOR2_X1    g05493(.A1(new_n5339_), .A2(new_n5340_), .ZN(new_n5686_));
  NOR2_X1    g05494(.A1(new_n5325_), .A2(new_n5342_), .ZN(new_n5687_));
  INV_X1     g05495(.I(new_n5687_), .ZN(new_n5688_));
  NAND4_X1   g05496(.A1(\asqrt[35] ), .A2(new_n5326_), .A3(new_n5686_), .A4(new_n5688_), .ZN(new_n5689_));
  AND3_X2    g05497(.A1(\asqrt[35] ), .A2(new_n5326_), .A3(new_n5688_), .Z(new_n5690_));
  OAI21_X1   g05498(.A1(new_n5690_), .A2(new_n5686_), .B(new_n5689_), .ZN(new_n5691_));
  INV_X1     g05499(.I(new_n5691_), .ZN(new_n5692_));
  NOR3_X1    g05500(.A1(new_n5683_), .A2(new_n5672_), .A3(\asqrt[39] ), .ZN(new_n5693_));
  NOR2_X1    g05501(.A1(new_n5693_), .A2(new_n5692_), .ZN(new_n5694_));
  OAI21_X1   g05502(.A1(new_n5694_), .A2(new_n5685_), .B(\asqrt[40] ), .ZN(new_n5695_));
  INV_X1     g05503(.I(new_n5347_), .ZN(new_n5696_));
  INV_X1     g05504(.I(new_n5344_), .ZN(new_n5697_));
  NAND2_X1   g05505(.A1(new_n5351_), .A2(new_n5343_), .ZN(new_n5698_));
  NAND3_X1   g05506(.A1(\asqrt[35] ), .A2(new_n5697_), .A3(new_n5698_), .ZN(new_n5699_));
  AND3_X2    g05507(.A1(new_n5697_), .A2(new_n5347_), .A3(new_n5698_), .Z(new_n5700_));
  AOI22_X1   g05508(.A1(new_n5699_), .A2(new_n5696_), .B1(\asqrt[35] ), .B2(new_n5700_), .ZN(new_n5701_));
  INV_X1     g05509(.I(new_n5701_), .ZN(new_n5702_));
  NAND2_X1   g05510(.A1(new_n5684_), .A2(new_n4071_), .ZN(new_n5703_));
  OAI21_X1   g05511(.A1(new_n5694_), .A2(new_n5703_), .B(new_n5702_), .ZN(new_n5704_));
  AOI21_X1   g05512(.A1(new_n5704_), .A2(new_n5695_), .B(new_n3782_), .ZN(new_n5705_));
  INV_X1     g05513(.I(new_n5361_), .ZN(new_n5706_));
  NOR3_X1    g05514(.A1(new_n5354_), .A2(new_n5706_), .A3(new_n5362_), .ZN(new_n5707_));
  INV_X1     g05515(.I(\asqrt[35] ), .ZN(new_n5708_));
  NOR3_X1    g05516(.A1(new_n5708_), .A2(new_n5354_), .A3(new_n5362_), .ZN(new_n5709_));
  INV_X1     g05517(.I(new_n5709_), .ZN(new_n5710_));
  AOI22_X1   g05518(.A1(new_n5710_), .A2(new_n5706_), .B1(\asqrt[35] ), .B2(new_n5707_), .ZN(new_n5711_));
  OAI21_X1   g05519(.A1(new_n5692_), .A2(new_n5693_), .B(new_n5684_), .ZN(new_n5712_));
  AOI21_X1   g05520(.A1(new_n5712_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n5713_));
  AOI21_X1   g05521(.A1(new_n5713_), .A2(new_n5704_), .B(new_n5711_), .ZN(new_n5714_));
  OAI21_X1   g05522(.A1(new_n5714_), .A2(new_n5705_), .B(\asqrt[42] ), .ZN(new_n5715_));
  INV_X1     g05523(.I(new_n5715_), .ZN(new_n5716_));
  INV_X1     g05524(.I(new_n5363_), .ZN(new_n5717_));
  INV_X1     g05525(.I(new_n5371_), .ZN(new_n5718_));
  NAND2_X1   g05526(.A1(new_n5717_), .A2(new_n5718_), .ZN(new_n5719_));
  NAND3_X1   g05527(.A1(\asqrt[35] ), .A2(new_n5364_), .A3(new_n5719_), .ZN(new_n5720_));
  AND3_X2    g05528(.A1(new_n5719_), .A2(new_n5364_), .A3(new_n5369_), .Z(new_n5721_));
  AOI22_X1   g05529(.A1(new_n5720_), .A2(new_n5370_), .B1(\asqrt[35] ), .B2(new_n5721_), .ZN(new_n5722_));
  NOR3_X1    g05530(.A1(new_n5714_), .A2(new_n5705_), .A3(\asqrt[42] ), .ZN(new_n5723_));
  NOR2_X1    g05531(.A1(new_n5723_), .A2(new_n5722_), .ZN(new_n5724_));
  OAI21_X1   g05532(.A1(new_n5724_), .A2(new_n5716_), .B(\asqrt[43] ), .ZN(new_n5725_));
  INV_X1     g05533(.I(new_n5377_), .ZN(new_n5726_));
  INV_X1     g05534(.I(new_n5372_), .ZN(new_n5727_));
  INV_X1     g05535(.I(new_n5379_), .ZN(new_n5728_));
  NOR2_X1    g05536(.A1(new_n5728_), .A2(new_n5727_), .ZN(new_n5729_));
  NOR3_X1    g05537(.A1(new_n5729_), .A2(new_n5373_), .A3(new_n5726_), .ZN(new_n5730_));
  NOR3_X1    g05538(.A1(new_n5708_), .A2(new_n5373_), .A3(new_n5729_), .ZN(new_n5731_));
  INV_X1     g05539(.I(new_n5731_), .ZN(new_n5732_));
  AOI22_X1   g05540(.A1(new_n5732_), .A2(new_n5726_), .B1(\asqrt[35] ), .B2(new_n5730_), .ZN(new_n5733_));
  INV_X1     g05541(.I(new_n5733_), .ZN(new_n5734_));
  NAND2_X1   g05542(.A1(new_n5715_), .A2(new_n3218_), .ZN(new_n5735_));
  OAI21_X1   g05543(.A1(new_n5724_), .A2(new_n5735_), .B(new_n5734_), .ZN(new_n5736_));
  AOI21_X1   g05544(.A1(new_n5736_), .A2(new_n5725_), .B(new_n2954_), .ZN(new_n5737_));
  INV_X1     g05545(.I(new_n5387_), .ZN(new_n5738_));
  NOR3_X1    g05546(.A1(new_n5708_), .A2(new_n5382_), .A3(new_n5388_), .ZN(new_n5739_));
  INV_X1     g05547(.I(new_n5739_), .ZN(new_n5740_));
  NOR3_X1    g05548(.A1(new_n5382_), .A2(new_n5738_), .A3(new_n5388_), .ZN(new_n5741_));
  AOI22_X1   g05549(.A1(new_n5740_), .A2(new_n5738_), .B1(\asqrt[35] ), .B2(new_n5741_), .ZN(new_n5742_));
  OAI21_X1   g05550(.A1(new_n5722_), .A2(new_n5723_), .B(new_n5715_), .ZN(new_n5743_));
  AOI21_X1   g05551(.A1(new_n5743_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n5744_));
  AOI21_X1   g05552(.A1(new_n5744_), .A2(new_n5736_), .B(new_n5742_), .ZN(new_n5745_));
  OAI21_X1   g05553(.A1(new_n5745_), .A2(new_n5737_), .B(\asqrt[45] ), .ZN(new_n5746_));
  INV_X1     g05554(.I(new_n5746_), .ZN(new_n5747_));
  NOR2_X1    g05555(.A1(new_n5389_), .A2(new_n5397_), .ZN(new_n5748_));
  INV_X1     g05556(.I(new_n5748_), .ZN(new_n5749_));
  AND3_X2    g05557(.A1(new_n5749_), .A2(new_n5390_), .A3(new_n5395_), .Z(new_n5750_));
  NAND3_X1   g05558(.A1(\asqrt[35] ), .A2(new_n5390_), .A3(new_n5749_), .ZN(new_n5751_));
  AOI22_X1   g05559(.A1(new_n5751_), .A2(new_n5396_), .B1(\asqrt[35] ), .B2(new_n5750_), .ZN(new_n5752_));
  NOR3_X1    g05560(.A1(new_n5745_), .A2(new_n5737_), .A3(\asqrt[45] ), .ZN(new_n5753_));
  NOR2_X1    g05561(.A1(new_n5753_), .A2(new_n5752_), .ZN(new_n5754_));
  OAI21_X1   g05562(.A1(new_n5754_), .A2(new_n5747_), .B(\asqrt[46] ), .ZN(new_n5755_));
  INV_X1     g05563(.I(new_n5403_), .ZN(new_n5756_));
  INV_X1     g05564(.I(new_n5398_), .ZN(new_n5757_));
  INV_X1     g05565(.I(new_n5405_), .ZN(new_n5758_));
  NOR2_X1    g05566(.A1(new_n5758_), .A2(new_n5757_), .ZN(new_n5759_));
  NOR3_X1    g05567(.A1(new_n5708_), .A2(new_n5399_), .A3(new_n5759_), .ZN(new_n5760_));
  INV_X1     g05568(.I(new_n5760_), .ZN(new_n5761_));
  NOR3_X1    g05569(.A1(new_n5759_), .A2(new_n5399_), .A3(new_n5756_), .ZN(new_n5762_));
  AOI22_X1   g05570(.A1(new_n5761_), .A2(new_n5756_), .B1(\asqrt[35] ), .B2(new_n5762_), .ZN(new_n5763_));
  INV_X1     g05571(.I(new_n5763_), .ZN(new_n5764_));
  NAND2_X1   g05572(.A1(new_n5746_), .A2(new_n2465_), .ZN(new_n5765_));
  OAI21_X1   g05573(.A1(new_n5754_), .A2(new_n5765_), .B(new_n5764_), .ZN(new_n5766_));
  AOI21_X1   g05574(.A1(new_n5766_), .A2(new_n5755_), .B(new_n2229_), .ZN(new_n5767_));
  INV_X1     g05575(.I(new_n5413_), .ZN(new_n5768_));
  NOR3_X1    g05576(.A1(new_n5408_), .A2(new_n5414_), .A3(new_n5768_), .ZN(new_n5769_));
  NOR3_X1    g05577(.A1(new_n5708_), .A2(new_n5408_), .A3(new_n5414_), .ZN(new_n5770_));
  INV_X1     g05578(.I(new_n5770_), .ZN(new_n5771_));
  AOI22_X1   g05579(.A1(new_n5771_), .A2(new_n5768_), .B1(\asqrt[35] ), .B2(new_n5769_), .ZN(new_n5772_));
  OAI21_X1   g05580(.A1(new_n5752_), .A2(new_n5753_), .B(new_n5746_), .ZN(new_n5773_));
  AOI21_X1   g05581(.A1(new_n5773_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n5774_));
  AOI21_X1   g05582(.A1(new_n5774_), .A2(new_n5766_), .B(new_n5772_), .ZN(new_n5775_));
  OAI21_X1   g05583(.A1(new_n5775_), .A2(new_n5767_), .B(\asqrt[48] ), .ZN(new_n5776_));
  INV_X1     g05584(.I(new_n5776_), .ZN(new_n5777_));
  INV_X1     g05585(.I(new_n5416_), .ZN(new_n5778_));
  NOR2_X1    g05586(.A1(new_n5415_), .A2(new_n5422_), .ZN(new_n5779_));
  NOR3_X1    g05587(.A1(new_n5708_), .A2(new_n5778_), .A3(new_n5779_), .ZN(new_n5780_));
  INV_X1     g05588(.I(new_n5780_), .ZN(new_n5781_));
  NOR3_X1    g05589(.A1(new_n5778_), .A2(new_n5421_), .A3(new_n5779_), .ZN(new_n5782_));
  AOI22_X1   g05590(.A1(new_n5781_), .A2(new_n5421_), .B1(\asqrt[35] ), .B2(new_n5782_), .ZN(new_n5783_));
  NOR3_X1    g05591(.A1(new_n5775_), .A2(new_n5767_), .A3(\asqrt[48] ), .ZN(new_n5784_));
  NOR2_X1    g05592(.A1(new_n5784_), .A2(new_n5783_), .ZN(new_n5785_));
  OAI21_X1   g05593(.A1(new_n5785_), .A2(new_n5777_), .B(\asqrt[49] ), .ZN(new_n5786_));
  INV_X1     g05594(.I(new_n5430_), .ZN(new_n5787_));
  INV_X1     g05595(.I(new_n5423_), .ZN(new_n5788_));
  INV_X1     g05596(.I(new_n5432_), .ZN(new_n5789_));
  NOR2_X1    g05597(.A1(new_n5789_), .A2(new_n5788_), .ZN(new_n5790_));
  NOR3_X1    g05598(.A1(new_n5790_), .A2(new_n5424_), .A3(new_n5787_), .ZN(new_n5791_));
  NOR3_X1    g05599(.A1(new_n5708_), .A2(new_n5424_), .A3(new_n5790_), .ZN(new_n5792_));
  INV_X1     g05600(.I(new_n5792_), .ZN(new_n5793_));
  AOI22_X1   g05601(.A1(new_n5793_), .A2(new_n5787_), .B1(\asqrt[35] ), .B2(new_n5791_), .ZN(new_n5794_));
  INV_X1     g05602(.I(new_n5794_), .ZN(new_n5795_));
  NAND2_X1   g05603(.A1(new_n5776_), .A2(new_n1806_), .ZN(new_n5796_));
  OAI21_X1   g05604(.A1(new_n5785_), .A2(new_n5796_), .B(new_n5795_), .ZN(new_n5797_));
  AOI21_X1   g05605(.A1(new_n5797_), .A2(new_n5786_), .B(new_n1612_), .ZN(new_n5798_));
  NOR3_X1    g05606(.A1(new_n5708_), .A2(new_n5435_), .A3(new_n5444_), .ZN(new_n5799_));
  INV_X1     g05607(.I(new_n5799_), .ZN(new_n5800_));
  NOR3_X1    g05608(.A1(new_n5435_), .A2(new_n5444_), .A3(new_n5474_), .ZN(new_n5801_));
  AOI22_X1   g05609(.A1(new_n5800_), .A2(new_n5474_), .B1(\asqrt[35] ), .B2(new_n5801_), .ZN(new_n5802_));
  OAI21_X1   g05610(.A1(new_n5783_), .A2(new_n5784_), .B(new_n5776_), .ZN(new_n5803_));
  AOI21_X1   g05611(.A1(new_n5803_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n5804_));
  AOI21_X1   g05612(.A1(new_n5804_), .A2(new_n5797_), .B(new_n5802_), .ZN(new_n5805_));
  OAI21_X1   g05613(.A1(new_n5805_), .A2(new_n5798_), .B(\asqrt[51] ), .ZN(new_n5806_));
  INV_X1     g05614(.I(new_n5806_), .ZN(new_n5807_));
  NOR2_X1    g05615(.A1(new_n5445_), .A2(new_n5452_), .ZN(new_n5808_));
  NOR3_X1    g05616(.A1(new_n5477_), .A2(new_n5808_), .A3(new_n5451_), .ZN(new_n5809_));
  NOR3_X1    g05617(.A1(new_n5708_), .A2(new_n5477_), .A3(new_n5808_), .ZN(new_n5810_));
  INV_X1     g05618(.I(new_n5810_), .ZN(new_n5811_));
  AOI22_X1   g05619(.A1(new_n5811_), .A2(new_n5451_), .B1(\asqrt[35] ), .B2(new_n5809_), .ZN(new_n5812_));
  NOR3_X1    g05620(.A1(new_n5805_), .A2(new_n5798_), .A3(\asqrt[51] ), .ZN(new_n5813_));
  NOR2_X1    g05621(.A1(new_n5813_), .A2(new_n5812_), .ZN(new_n5814_));
  OAI21_X1   g05622(.A1(new_n5814_), .A2(new_n5807_), .B(\asqrt[52] ), .ZN(new_n5815_));
  NOR2_X1    g05623(.A1(new_n5489_), .A2(new_n5479_), .ZN(new_n5816_));
  NOR3_X1    g05624(.A1(new_n5708_), .A2(new_n5454_), .A3(new_n5816_), .ZN(new_n5817_));
  INV_X1     g05625(.I(new_n5817_), .ZN(new_n5818_));
  NOR3_X1    g05626(.A1(new_n5816_), .A2(new_n5454_), .A3(new_n5488_), .ZN(new_n5819_));
  AOI22_X1   g05627(.A1(new_n5818_), .A2(new_n5488_), .B1(\asqrt[35] ), .B2(new_n5819_), .ZN(new_n5820_));
  INV_X1     g05628(.I(new_n5820_), .ZN(new_n5821_));
  NAND2_X1   g05629(.A1(new_n5806_), .A2(new_n1256_), .ZN(new_n5822_));
  OAI21_X1   g05630(.A1(new_n5814_), .A2(new_n5822_), .B(new_n5821_), .ZN(new_n5823_));
  AOI21_X1   g05631(.A1(new_n5823_), .A2(new_n5815_), .B(new_n1103_), .ZN(new_n5824_));
  NOR3_X1    g05632(.A1(new_n5491_), .A2(new_n5525_), .A3(new_n5473_), .ZN(new_n5825_));
  NOR3_X1    g05633(.A1(new_n5708_), .A2(new_n5491_), .A3(new_n5525_), .ZN(new_n5826_));
  INV_X1     g05634(.I(new_n5826_), .ZN(new_n5827_));
  AOI22_X1   g05635(.A1(new_n5827_), .A2(new_n5473_), .B1(\asqrt[35] ), .B2(new_n5825_), .ZN(new_n5828_));
  OAI21_X1   g05636(.A1(new_n5812_), .A2(new_n5813_), .B(new_n5806_), .ZN(new_n5829_));
  AOI21_X1   g05637(.A1(new_n5829_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n5830_));
  AOI21_X1   g05638(.A1(new_n5830_), .A2(new_n5823_), .B(new_n5828_), .ZN(new_n5831_));
  OAI21_X1   g05639(.A1(new_n5831_), .A2(new_n5824_), .B(\asqrt[54] ), .ZN(new_n5832_));
  INV_X1     g05640(.I(new_n5832_), .ZN(new_n5833_));
  NOR2_X1    g05641(.A1(new_n5514_), .A2(new_n5503_), .ZN(new_n5834_));
  NOR3_X1    g05642(.A1(new_n5708_), .A2(new_n5483_), .A3(new_n5834_), .ZN(new_n5835_));
  INV_X1     g05643(.I(new_n5835_), .ZN(new_n5836_));
  NOR3_X1    g05644(.A1(new_n5483_), .A2(new_n5834_), .A3(new_n5513_), .ZN(new_n5837_));
  AOI22_X1   g05645(.A1(new_n5836_), .A2(new_n5513_), .B1(\asqrt[35] ), .B2(new_n5837_), .ZN(new_n5838_));
  NOR3_X1    g05646(.A1(new_n5831_), .A2(new_n5824_), .A3(\asqrt[54] ), .ZN(new_n5839_));
  NOR2_X1    g05647(.A1(new_n5839_), .A2(new_n5838_), .ZN(new_n5840_));
  OAI21_X1   g05648(.A1(new_n5840_), .A2(new_n5833_), .B(\asqrt[55] ), .ZN(new_n5841_));
  NOR2_X1    g05649(.A1(new_n5505_), .A2(new_n5493_), .ZN(new_n5842_));
  NOR3_X1    g05650(.A1(new_n5842_), .A2(new_n5516_), .A3(new_n5501_), .ZN(new_n5843_));
  NOR3_X1    g05651(.A1(new_n5708_), .A2(new_n5516_), .A3(new_n5842_), .ZN(new_n5844_));
  INV_X1     g05652(.I(new_n5844_), .ZN(new_n5845_));
  AOI22_X1   g05653(.A1(new_n5845_), .A2(new_n5501_), .B1(\asqrt[35] ), .B2(new_n5843_), .ZN(new_n5846_));
  INV_X1     g05654(.I(new_n5846_), .ZN(new_n5847_));
  NAND2_X1   g05655(.A1(new_n5832_), .A2(new_n823_), .ZN(new_n5848_));
  OAI21_X1   g05656(.A1(new_n5840_), .A2(new_n5848_), .B(new_n5847_), .ZN(new_n5849_));
  AOI21_X1   g05657(.A1(new_n5849_), .A2(new_n5841_), .B(new_n703_), .ZN(new_n5850_));
  NOR3_X1    g05658(.A1(new_n5708_), .A2(new_n5507_), .A3(new_n5539_), .ZN(new_n5851_));
  INV_X1     g05659(.I(new_n5851_), .ZN(new_n5852_));
  NOR3_X1    g05660(.A1(new_n5507_), .A2(new_n5539_), .A3(new_n5550_), .ZN(new_n5853_));
  AOI22_X1   g05661(.A1(new_n5852_), .A2(new_n5550_), .B1(\asqrt[35] ), .B2(new_n5853_), .ZN(new_n5854_));
  OAI21_X1   g05662(.A1(new_n5838_), .A2(new_n5839_), .B(new_n5832_), .ZN(new_n5855_));
  AOI21_X1   g05663(.A1(new_n5855_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n5856_));
  AOI21_X1   g05664(.A1(new_n5856_), .A2(new_n5849_), .B(new_n5854_), .ZN(new_n5857_));
  OAI21_X1   g05665(.A1(new_n5857_), .A2(new_n5850_), .B(\asqrt[57] ), .ZN(new_n5858_));
  NOR2_X1    g05666(.A1(new_n5530_), .A2(new_n5518_), .ZN(new_n5859_));
  NOR3_X1    g05667(.A1(new_n5553_), .A2(new_n5859_), .A3(new_n5524_), .ZN(new_n5860_));
  NOR3_X1    g05668(.A1(new_n5708_), .A2(new_n5553_), .A3(new_n5859_), .ZN(new_n5861_));
  INV_X1     g05669(.I(new_n5861_), .ZN(new_n5862_));
  AOI22_X1   g05670(.A1(new_n5862_), .A2(new_n5524_), .B1(\asqrt[35] ), .B2(new_n5860_), .ZN(new_n5863_));
  INV_X1     g05671(.I(new_n5863_), .ZN(new_n5864_));
  INV_X1     g05672(.I(new_n5838_), .ZN(new_n5865_));
  INV_X1     g05673(.I(new_n5812_), .ZN(new_n5866_));
  INV_X1     g05674(.I(new_n5783_), .ZN(new_n5867_));
  INV_X1     g05675(.I(new_n5752_), .ZN(new_n5868_));
  INV_X1     g05676(.I(new_n5722_), .ZN(new_n5869_));
  NAND2_X1   g05677(.A1(new_n5642_), .A2(new_n5653_), .ZN(new_n5870_));
  OAI21_X1   g05678(.A1(new_n5637_), .A2(new_n5641_), .B(new_n5644_), .ZN(new_n5871_));
  NAND2_X1   g05679(.A1(new_n5871_), .A2(\a[71] ), .ZN(new_n5872_));
  NAND3_X1   g05680(.A1(new_n5870_), .A2(new_n5872_), .A3(new_n5661_), .ZN(new_n5873_));
  AOI21_X1   g05681(.A1(new_n5873_), .A2(new_n5678_), .B(new_n5024_), .ZN(new_n5874_));
  OAI21_X1   g05682(.A1(new_n5665_), .A2(new_n5656_), .B(\a[72] ), .ZN(new_n5875_));
  NAND3_X1   g05683(.A1(new_n5666_), .A2(new_n5661_), .A3(new_n5281_), .ZN(new_n5876_));
  NAND2_X1   g05684(.A1(new_n5642_), .A2(new_n5634_), .ZN(new_n5877_));
  AOI21_X1   g05685(.A1(new_n5877_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n5878_));
  AOI22_X1   g05686(.A1(new_n5873_), .A2(new_n5878_), .B1(new_n5875_), .B2(new_n5876_), .ZN(new_n5879_));
  OAI21_X1   g05687(.A1(new_n5879_), .A2(new_n5874_), .B(\asqrt[38] ), .ZN(new_n5880_));
  NAND2_X1   g05688(.A1(new_n5880_), .A2(new_n4298_), .ZN(new_n5881_));
  OAI21_X1   g05689(.A1(new_n5881_), .A2(new_n5683_), .B(new_n5691_), .ZN(new_n5882_));
  AOI21_X1   g05690(.A1(new_n5882_), .A2(new_n5684_), .B(new_n4071_), .ZN(new_n5883_));
  INV_X1     g05691(.I(new_n5677_), .ZN(new_n5884_));
  AOI21_X1   g05692(.A1(\a[71] ), .A2(new_n5871_), .B(new_n5656_), .ZN(new_n5885_));
  AOI21_X1   g05693(.A1(new_n5885_), .A2(new_n5870_), .B(new_n5643_), .ZN(new_n5886_));
  OAI21_X1   g05694(.A1(new_n5886_), .A2(new_n5024_), .B(new_n4696_), .ZN(new_n5887_));
  OAI21_X1   g05695(.A1(new_n5887_), .A2(new_n5879_), .B(new_n5884_), .ZN(new_n5888_));
  NAND2_X1   g05696(.A1(new_n5888_), .A2(new_n5880_), .ZN(new_n5889_));
  AOI21_X1   g05697(.A1(new_n5889_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n5890_));
  AOI21_X1   g05698(.A1(new_n5890_), .A2(new_n5882_), .B(new_n5701_), .ZN(new_n5891_));
  OAI21_X1   g05699(.A1(new_n5891_), .A2(new_n5883_), .B(\asqrt[41] ), .ZN(new_n5892_));
  NAND2_X1   g05700(.A1(new_n5892_), .A2(new_n3419_), .ZN(new_n5893_));
  OAI21_X1   g05701(.A1(new_n5893_), .A2(new_n5714_), .B(new_n5869_), .ZN(new_n5894_));
  NAND3_X1   g05702(.A1(new_n5894_), .A2(new_n3218_), .A3(new_n5715_), .ZN(new_n5895_));
  AOI22_X1   g05703(.A1(new_n5895_), .A2(new_n5734_), .B1(new_n5743_), .B2(\asqrt[43] ), .ZN(new_n5896_));
  OAI21_X1   g05704(.A1(new_n5896_), .A2(new_n2954_), .B(new_n2641_), .ZN(new_n5897_));
  OAI21_X1   g05705(.A1(new_n5897_), .A2(new_n5745_), .B(new_n5868_), .ZN(new_n5898_));
  AOI21_X1   g05706(.A1(new_n5898_), .A2(new_n5746_), .B(new_n2465_), .ZN(new_n5899_));
  AOI21_X1   g05707(.A1(new_n5894_), .A2(new_n5715_), .B(new_n3218_), .ZN(new_n5900_));
  NOR3_X1    g05708(.A1(new_n5891_), .A2(new_n5883_), .A3(\asqrt[41] ), .ZN(new_n5901_));
  OAI21_X1   g05709(.A1(new_n5711_), .A2(new_n5901_), .B(new_n5892_), .ZN(new_n5902_));
  AOI21_X1   g05710(.A1(new_n5902_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n5903_));
  AOI21_X1   g05711(.A1(new_n5903_), .A2(new_n5894_), .B(new_n5733_), .ZN(new_n5904_));
  NOR3_X1    g05712(.A1(new_n5904_), .A2(\asqrt[44] ), .A3(new_n5900_), .ZN(new_n5905_));
  OAI22_X1   g05713(.A1(new_n5905_), .A2(new_n5742_), .B1(new_n5896_), .B2(new_n2954_), .ZN(new_n5906_));
  AOI21_X1   g05714(.A1(new_n5906_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n5907_));
  AOI21_X1   g05715(.A1(new_n5907_), .A2(new_n5898_), .B(new_n5763_), .ZN(new_n5908_));
  OAI21_X1   g05716(.A1(new_n5908_), .A2(new_n5899_), .B(\asqrt[47] ), .ZN(new_n5909_));
  NAND2_X1   g05717(.A1(new_n5909_), .A2(new_n1956_), .ZN(new_n5910_));
  OAI21_X1   g05718(.A1(new_n5910_), .A2(new_n5775_), .B(new_n5867_), .ZN(new_n5911_));
  AOI21_X1   g05719(.A1(new_n5911_), .A2(new_n5776_), .B(new_n1806_), .ZN(new_n5912_));
  NOR3_X1    g05720(.A1(new_n5908_), .A2(\asqrt[47] ), .A3(new_n5899_), .ZN(new_n5913_));
  OAI21_X1   g05721(.A1(new_n5772_), .A2(new_n5913_), .B(new_n5909_), .ZN(new_n5914_));
  AOI21_X1   g05722(.A1(new_n5914_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n5915_));
  AOI21_X1   g05723(.A1(new_n5915_), .A2(new_n5911_), .B(new_n5794_), .ZN(new_n5916_));
  OAI21_X1   g05724(.A1(new_n5916_), .A2(new_n5912_), .B(\asqrt[50] ), .ZN(new_n5917_));
  NAND2_X1   g05725(.A1(new_n5917_), .A2(new_n1376_), .ZN(new_n5918_));
  OAI21_X1   g05726(.A1(new_n5918_), .A2(new_n5805_), .B(new_n5866_), .ZN(new_n5919_));
  AOI21_X1   g05727(.A1(new_n5919_), .A2(new_n5806_), .B(new_n1256_), .ZN(new_n5920_));
  NOR3_X1    g05728(.A1(new_n5916_), .A2(\asqrt[50] ), .A3(new_n5912_), .ZN(new_n5921_));
  OAI21_X1   g05729(.A1(new_n5802_), .A2(new_n5921_), .B(new_n5917_), .ZN(new_n5922_));
  AOI21_X1   g05730(.A1(new_n5922_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n5923_));
  AOI21_X1   g05731(.A1(new_n5923_), .A2(new_n5919_), .B(new_n5820_), .ZN(new_n5924_));
  OAI21_X1   g05732(.A1(new_n5924_), .A2(new_n5920_), .B(\asqrt[53] ), .ZN(new_n5925_));
  NAND2_X1   g05733(.A1(new_n5925_), .A2(new_n904_), .ZN(new_n5926_));
  OAI21_X1   g05734(.A1(new_n5926_), .A2(new_n5831_), .B(new_n5865_), .ZN(new_n5927_));
  AOI21_X1   g05735(.A1(new_n5927_), .A2(new_n5832_), .B(new_n823_), .ZN(new_n5928_));
  NOR3_X1    g05736(.A1(new_n5924_), .A2(\asqrt[53] ), .A3(new_n5920_), .ZN(new_n5929_));
  OAI21_X1   g05737(.A1(new_n5828_), .A2(new_n5929_), .B(new_n5925_), .ZN(new_n5930_));
  AOI21_X1   g05738(.A1(new_n5930_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n5931_));
  AOI21_X1   g05739(.A1(new_n5931_), .A2(new_n5927_), .B(new_n5846_), .ZN(new_n5932_));
  OAI21_X1   g05740(.A1(new_n5932_), .A2(new_n5928_), .B(\asqrt[56] ), .ZN(new_n5933_));
  NAND2_X1   g05741(.A1(new_n5933_), .A2(new_n531_), .ZN(new_n5934_));
  OAI21_X1   g05742(.A1(new_n5934_), .A2(new_n5857_), .B(new_n5864_), .ZN(new_n5935_));
  AOI21_X1   g05743(.A1(new_n5935_), .A2(new_n5858_), .B(new_n436_), .ZN(new_n5936_));
  NOR2_X1    g05744(.A1(new_n5565_), .A2(new_n5555_), .ZN(new_n5937_));
  NOR3_X1    g05745(.A1(new_n5708_), .A2(new_n5532_), .A3(new_n5937_), .ZN(new_n5938_));
  INV_X1     g05746(.I(new_n5938_), .ZN(new_n5939_));
  NOR3_X1    g05747(.A1(new_n5937_), .A2(new_n5532_), .A3(new_n5564_), .ZN(new_n5940_));
  AOI22_X1   g05748(.A1(new_n5939_), .A2(new_n5564_), .B1(\asqrt[35] ), .B2(new_n5940_), .ZN(new_n5941_));
  NOR3_X1    g05749(.A1(new_n5932_), .A2(\asqrt[56] ), .A3(new_n5928_), .ZN(new_n5942_));
  OAI21_X1   g05750(.A1(new_n5854_), .A2(new_n5942_), .B(new_n5933_), .ZN(new_n5943_));
  AOI21_X1   g05751(.A1(new_n5943_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n5944_));
  AOI21_X1   g05752(.A1(new_n5944_), .A2(new_n5935_), .B(new_n5941_), .ZN(new_n5945_));
  OAI21_X1   g05753(.A1(new_n5945_), .A2(new_n5936_), .B(\asqrt[59] ), .ZN(new_n5946_));
  NOR3_X1    g05754(.A1(new_n5567_), .A2(new_n5601_), .A3(new_n5549_), .ZN(new_n5947_));
  NOR3_X1    g05755(.A1(new_n5708_), .A2(new_n5567_), .A3(new_n5601_), .ZN(new_n5948_));
  INV_X1     g05756(.I(new_n5948_), .ZN(new_n5949_));
  AOI22_X1   g05757(.A1(new_n5949_), .A2(new_n5549_), .B1(\asqrt[35] ), .B2(new_n5947_), .ZN(new_n5950_));
  INV_X1     g05758(.I(new_n5950_), .ZN(new_n5951_));
  INV_X1     g05759(.I(new_n5858_), .ZN(new_n5952_));
  NOR3_X1    g05760(.A1(new_n5857_), .A2(new_n5850_), .A3(\asqrt[57] ), .ZN(new_n5953_));
  NOR2_X1    g05761(.A1(new_n5953_), .A2(new_n5863_), .ZN(new_n5954_));
  OAI21_X1   g05762(.A1(new_n5954_), .A2(new_n5952_), .B(\asqrt[58] ), .ZN(new_n5955_));
  NAND2_X1   g05763(.A1(new_n5955_), .A2(new_n327_), .ZN(new_n5956_));
  OAI21_X1   g05764(.A1(new_n5956_), .A2(new_n5945_), .B(new_n5951_), .ZN(new_n5957_));
  AOI21_X1   g05765(.A1(new_n5957_), .A2(new_n5946_), .B(new_n306_), .ZN(new_n5958_));
  NOR2_X1    g05766(.A1(new_n5590_), .A2(new_n5579_), .ZN(new_n5959_));
  NOR3_X1    g05767(.A1(new_n5708_), .A2(new_n5559_), .A3(new_n5959_), .ZN(new_n5960_));
  INV_X1     g05768(.I(new_n5960_), .ZN(new_n5961_));
  NOR3_X1    g05769(.A1(new_n5559_), .A2(new_n5959_), .A3(new_n5589_), .ZN(new_n5962_));
  AOI22_X1   g05770(.A1(new_n5961_), .A2(new_n5589_), .B1(\asqrt[35] ), .B2(new_n5962_), .ZN(new_n5963_));
  INV_X1     g05771(.I(new_n5941_), .ZN(new_n5964_));
  NAND2_X1   g05772(.A1(new_n5858_), .A2(new_n436_), .ZN(new_n5965_));
  OAI21_X1   g05773(.A1(new_n5954_), .A2(new_n5965_), .B(new_n5964_), .ZN(new_n5966_));
  AOI21_X1   g05774(.A1(new_n5966_), .A2(new_n5955_), .B(new_n327_), .ZN(new_n5967_));
  NOR2_X1    g05775(.A1(new_n5967_), .A2(\asqrt[60] ), .ZN(new_n5968_));
  AOI21_X1   g05776(.A1(new_n5968_), .A2(new_n5957_), .B(new_n5963_), .ZN(new_n5969_));
  OAI21_X1   g05777(.A1(new_n5969_), .A2(new_n5958_), .B(\asqrt[61] ), .ZN(new_n5970_));
  NOR2_X1    g05778(.A1(new_n5581_), .A2(new_n5569_), .ZN(new_n5971_));
  NOR3_X1    g05779(.A1(new_n5971_), .A2(new_n5592_), .A3(new_n5577_), .ZN(new_n5972_));
  NOR3_X1    g05780(.A1(new_n5708_), .A2(new_n5592_), .A3(new_n5971_), .ZN(new_n5973_));
  INV_X1     g05781(.I(new_n5973_), .ZN(new_n5974_));
  AOI22_X1   g05782(.A1(new_n5974_), .A2(new_n5577_), .B1(\asqrt[35] ), .B2(new_n5972_), .ZN(new_n5975_));
  INV_X1     g05783(.I(new_n5975_), .ZN(new_n5976_));
  OAI21_X1   g05784(.A1(new_n5863_), .A2(new_n5953_), .B(new_n5858_), .ZN(new_n5977_));
  AOI21_X1   g05785(.A1(new_n5977_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n5978_));
  AOI21_X1   g05786(.A1(new_n5978_), .A2(new_n5966_), .B(new_n5950_), .ZN(new_n5979_));
  OAI21_X1   g05787(.A1(new_n5979_), .A2(new_n5967_), .B(\asqrt[60] ), .ZN(new_n5980_));
  NAND2_X1   g05788(.A1(new_n5980_), .A2(new_n218_), .ZN(new_n5981_));
  OAI21_X1   g05789(.A1(new_n5981_), .A2(new_n5969_), .B(new_n5976_), .ZN(new_n5982_));
  AOI21_X1   g05790(.A1(new_n5982_), .A2(new_n5970_), .B(new_n207_), .ZN(new_n5983_));
  NOR3_X1    g05791(.A1(new_n5708_), .A2(new_n5583_), .A3(new_n5617_), .ZN(new_n5984_));
  INV_X1     g05792(.I(new_n5984_), .ZN(new_n5985_));
  NOR3_X1    g05793(.A1(new_n5583_), .A2(new_n5617_), .A3(new_n5645_), .ZN(new_n5986_));
  AOI22_X1   g05794(.A1(new_n5985_), .A2(new_n5645_), .B1(\asqrt[35] ), .B2(new_n5986_), .ZN(new_n5987_));
  NOR3_X1    g05795(.A1(new_n5979_), .A2(new_n5967_), .A3(\asqrt[60] ), .ZN(new_n5988_));
  OAI21_X1   g05796(.A1(new_n5963_), .A2(new_n5988_), .B(new_n5980_), .ZN(new_n5989_));
  AOI21_X1   g05797(.A1(new_n5989_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n5990_));
  AOI21_X1   g05798(.A1(new_n5990_), .A2(new_n5982_), .B(new_n5987_), .ZN(new_n5991_));
  AND3_X2    g05799(.A1(new_n5595_), .A2(new_n5648_), .A3(new_n5599_), .Z(new_n5992_));
  NAND2_X1   g05800(.A1(\asqrt[35] ), .A2(new_n5992_), .ZN(new_n5993_));
  INV_X1     g05801(.I(new_n5993_), .ZN(new_n5994_));
  AND2_X2    g05802(.A1(new_n5595_), .A2(new_n5648_), .Z(new_n5995_));
  AOI21_X1   g05803(.A1(\asqrt[35] ), .A2(new_n5995_), .B(new_n5599_), .ZN(new_n5996_));
  NOR2_X1    g05804(.A1(new_n5994_), .A2(new_n5996_), .ZN(new_n5997_));
  NOR3_X1    g05805(.A1(new_n5708_), .A2(new_n5649_), .A3(new_n5639_), .ZN(new_n5998_));
  NOR3_X1    g05806(.A1(new_n5997_), .A2(new_n5662_), .A3(new_n5998_), .ZN(new_n5999_));
  OAI21_X1   g05807(.A1(new_n5991_), .A2(new_n5983_), .B(new_n5999_), .ZN(new_n6000_));
  NAND2_X1   g05808(.A1(new_n6000_), .A2(new_n193_), .ZN(new_n6001_));
  INV_X1     g05809(.I(new_n5987_), .ZN(new_n6002_));
  NAND3_X1   g05810(.A1(new_n5982_), .A2(new_n5970_), .A3(new_n207_), .ZN(new_n6003_));
  NAND2_X1   g05811(.A1(new_n6003_), .A2(new_n6002_), .ZN(new_n6004_));
  INV_X1     g05812(.I(new_n5997_), .ZN(new_n6005_));
  NOR2_X1    g05813(.A1(new_n5983_), .A2(new_n6005_), .ZN(new_n6006_));
  AOI21_X1   g05814(.A1(\asqrt[35] ), .A2(new_n5612_), .B(new_n5635_), .ZN(new_n6007_));
  OAI21_X1   g05815(.A1(new_n5649_), .A2(new_n5639_), .B(\asqrt[63] ), .ZN(new_n6008_));
  NOR2_X1    g05816(.A1(new_n6007_), .A2(new_n6008_), .ZN(new_n6009_));
  INV_X1     g05817(.I(new_n5662_), .ZN(new_n6010_));
  AND3_X2    g05818(.A1(new_n5611_), .A2(new_n5609_), .A3(new_n5625_), .Z(new_n6011_));
  NAND4_X1   g05819(.A1(new_n6010_), .A2(new_n5650_), .A3(new_n5622_), .A4(new_n6011_), .ZN(new_n6012_));
  INV_X1     g05820(.I(new_n6012_), .ZN(new_n6013_));
  NOR2_X1    g05821(.A1(new_n6009_), .A2(new_n6013_), .ZN(new_n6014_));
  INV_X1     g05822(.I(new_n6014_), .ZN(new_n6015_));
  AOI21_X1   g05823(.A1(new_n6006_), .A2(new_n6004_), .B(new_n6015_), .ZN(new_n6016_));
  NAND2_X1   g05824(.A1(new_n6001_), .A2(new_n6016_), .ZN(\asqrt[34] ));
  NOR2_X1    g05825(.A1(\a[66] ), .A2(\a[67] ), .ZN(new_n6018_));
  INV_X1     g05826(.I(new_n6018_), .ZN(new_n6019_));
  NOR2_X1    g05827(.A1(new_n6019_), .A2(\a[68] ), .ZN(new_n6020_));
  INV_X1     g05828(.I(new_n6020_), .ZN(new_n6021_));
  INV_X1     g05829(.I(new_n5963_), .ZN(new_n6022_));
  NAND2_X1   g05830(.A1(new_n5946_), .A2(new_n306_), .ZN(new_n6023_));
  OAI21_X1   g05831(.A1(new_n6023_), .A2(new_n5979_), .B(new_n6022_), .ZN(new_n6024_));
  AOI21_X1   g05832(.A1(new_n6024_), .A2(new_n5980_), .B(new_n218_), .ZN(new_n6025_));
  NOR3_X1    g05833(.A1(new_n5945_), .A2(\asqrt[59] ), .A3(new_n5936_), .ZN(new_n6026_));
  OAI21_X1   g05834(.A1(new_n5950_), .A2(new_n6026_), .B(new_n5946_), .ZN(new_n6027_));
  AOI21_X1   g05835(.A1(new_n6027_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n6028_));
  AOI21_X1   g05836(.A1(new_n6028_), .A2(new_n6024_), .B(new_n5975_), .ZN(new_n6029_));
  OAI21_X1   g05837(.A1(new_n6029_), .A2(new_n6025_), .B(\asqrt[62] ), .ZN(new_n6030_));
  NOR3_X1    g05838(.A1(new_n6029_), .A2(\asqrt[62] ), .A3(new_n6025_), .ZN(new_n6031_));
  OAI21_X1   g05839(.A1(new_n5987_), .A2(new_n6031_), .B(new_n6030_), .ZN(new_n6032_));
  AOI21_X1   g05840(.A1(new_n6032_), .A2(new_n5999_), .B(\asqrt[63] ), .ZN(new_n6033_));
  NAND2_X1   g05841(.A1(new_n6030_), .A2(new_n5997_), .ZN(new_n6034_));
  OAI21_X1   g05842(.A1(new_n6034_), .A2(new_n5991_), .B(new_n6014_), .ZN(new_n6035_));
  OAI21_X1   g05843(.A1(new_n6033_), .A2(new_n6035_), .B(\a[68] ), .ZN(new_n6036_));
  AOI21_X1   g05844(.A1(new_n6036_), .A2(new_n6021_), .B(new_n5708_), .ZN(new_n6037_));
  INV_X1     g05845(.I(\a[68] ), .ZN(new_n6038_));
  AOI21_X1   g05846(.A1(new_n6001_), .A2(new_n6016_), .B(new_n6038_), .ZN(new_n6039_));
  NAND2_X1   g05847(.A1(new_n5625_), .A2(new_n6021_), .ZN(new_n6040_));
  NOR4_X1    g05848(.A1(new_n5637_), .A2(new_n5662_), .A3(new_n5623_), .A4(new_n6040_), .ZN(new_n6041_));
  INV_X1     g05849(.I(new_n6041_), .ZN(new_n6042_));
  NOR2_X1    g05850(.A1(new_n6039_), .A2(new_n6042_), .ZN(new_n6043_));
  AOI21_X1   g05851(.A1(new_n6001_), .A2(new_n6016_), .B(new_n5632_), .ZN(new_n6044_));
  INV_X1     g05852(.I(\a[69] ), .ZN(new_n6045_));
  AOI21_X1   g05853(.A1(\asqrt[34] ), .A2(new_n6038_), .B(new_n6045_), .ZN(new_n6046_));
  NOR3_X1    g05854(.A1(new_n6043_), .A2(new_n6046_), .A3(new_n6044_), .ZN(new_n6047_));
  OAI21_X1   g05855(.A1(new_n6047_), .A2(new_n6037_), .B(\asqrt[36] ), .ZN(new_n6048_));
  OAI21_X1   g05856(.A1(new_n6033_), .A2(new_n6035_), .B(new_n5631_), .ZN(new_n6049_));
  NAND2_X1   g05857(.A1(new_n6006_), .A2(new_n6004_), .ZN(new_n6050_));
  INV_X1     g05858(.I(new_n6009_), .ZN(new_n6051_));
  NOR2_X1    g05859(.A1(new_n6013_), .A2(new_n5708_), .ZN(new_n6052_));
  NAND4_X1   g05860(.A1(new_n6001_), .A2(new_n6050_), .A3(new_n6051_), .A4(new_n6052_), .ZN(new_n6053_));
  AOI21_X1   g05861(.A1(new_n6053_), .A2(new_n6049_), .B(new_n5644_), .ZN(new_n6054_));
  INV_X1     g05862(.I(new_n6050_), .ZN(new_n6055_));
  NAND2_X1   g05863(.A1(new_n6051_), .A2(new_n6052_), .ZN(new_n6056_));
  NOR3_X1    g05864(.A1(new_n6055_), .A2(new_n6033_), .A3(new_n6056_), .ZN(new_n6057_));
  NOR3_X1    g05865(.A1(new_n6057_), .A2(new_n6044_), .A3(\a[70] ), .ZN(new_n6058_));
  OAI21_X1   g05866(.A1(new_n6039_), .A2(new_n6020_), .B(\asqrt[35] ), .ZN(new_n6059_));
  NAND2_X1   g05867(.A1(new_n6059_), .A2(new_n5277_), .ZN(new_n6060_));
  OAI22_X1   g05868(.A1(new_n6047_), .A2(new_n6060_), .B1(new_n6054_), .B2(new_n6058_), .ZN(new_n6061_));
  AOI21_X1   g05869(.A1(new_n6061_), .A2(new_n6048_), .B(new_n5024_), .ZN(new_n6062_));
  NOR3_X1    g05870(.A1(new_n5885_), .A2(new_n5643_), .A3(new_n5655_), .ZN(new_n6063_));
  NAND3_X1   g05871(.A1(\asqrt[34] ), .A2(new_n5678_), .A3(new_n5870_), .ZN(new_n6064_));
  AOI22_X1   g05872(.A1(new_n6064_), .A2(new_n5885_), .B1(\asqrt[34] ), .B2(new_n6063_), .ZN(new_n6065_));
  AOI21_X1   g05873(.A1(new_n6001_), .A2(new_n6016_), .B(\a[68] ), .ZN(new_n6066_));
  OAI21_X1   g05874(.A1(new_n6045_), .A2(new_n6066_), .B(new_n6049_), .ZN(new_n6067_));
  OAI21_X1   g05875(.A1(new_n6067_), .A2(new_n6043_), .B(new_n6059_), .ZN(new_n6068_));
  AOI21_X1   g05876(.A1(new_n6068_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n6069_));
  AOI21_X1   g05877(.A1(new_n6069_), .A2(new_n6061_), .B(new_n6065_), .ZN(new_n6070_));
  OAI21_X1   g05878(.A1(new_n6070_), .A2(new_n6062_), .B(\asqrt[38] ), .ZN(new_n6071_));
  INV_X1     g05879(.I(new_n6071_), .ZN(new_n6072_));
  NOR2_X1    g05880(.A1(new_n5667_), .A2(new_n5668_), .ZN(new_n6073_));
  NOR2_X1    g05881(.A1(new_n5659_), .A2(new_n5670_), .ZN(new_n6074_));
  INV_X1     g05882(.I(new_n6074_), .ZN(new_n6075_));
  NAND4_X1   g05883(.A1(\asqrt[34] ), .A2(new_n5660_), .A3(new_n6073_), .A4(new_n6075_), .ZN(new_n6076_));
  INV_X1     g05884(.I(\asqrt[34] ), .ZN(new_n6077_));
  NOR3_X1    g05885(.A1(new_n6077_), .A2(new_n5874_), .A3(new_n6074_), .ZN(new_n6078_));
  OAI21_X1   g05886(.A1(new_n6078_), .A2(new_n6073_), .B(new_n6076_), .ZN(new_n6079_));
  INV_X1     g05887(.I(new_n6079_), .ZN(new_n6080_));
  NOR3_X1    g05888(.A1(new_n6070_), .A2(new_n6062_), .A3(\asqrt[38] ), .ZN(new_n6081_));
  NOR2_X1    g05889(.A1(new_n6081_), .A2(new_n6080_), .ZN(new_n6082_));
  OAI21_X1   g05890(.A1(new_n6082_), .A2(new_n6072_), .B(\asqrt[39] ), .ZN(new_n6083_));
  NOR2_X1    g05891(.A1(new_n5887_), .A2(new_n5879_), .ZN(new_n6084_));
  NOR3_X1    g05892(.A1(new_n6077_), .A2(new_n5672_), .A3(new_n6084_), .ZN(new_n6085_));
  INV_X1     g05893(.I(new_n6085_), .ZN(new_n6086_));
  NOR3_X1    g05894(.A1(new_n6084_), .A2(new_n5672_), .A3(new_n5884_), .ZN(new_n6087_));
  AOI22_X1   g05895(.A1(new_n6086_), .A2(new_n5884_), .B1(\asqrt[34] ), .B2(new_n6087_), .ZN(new_n6088_));
  INV_X1     g05896(.I(new_n6088_), .ZN(new_n6089_));
  NAND2_X1   g05897(.A1(new_n6071_), .A2(new_n4298_), .ZN(new_n6090_));
  OAI21_X1   g05898(.A1(new_n6082_), .A2(new_n6090_), .B(new_n6089_), .ZN(new_n6091_));
  AOI21_X1   g05899(.A1(new_n6091_), .A2(new_n6083_), .B(new_n4071_), .ZN(new_n6092_));
  NOR3_X1    g05900(.A1(new_n5685_), .A2(new_n5693_), .A3(new_n5691_), .ZN(new_n6093_));
  NOR3_X1    g05901(.A1(new_n6077_), .A2(new_n5685_), .A3(new_n5693_), .ZN(new_n6094_));
  INV_X1     g05902(.I(new_n6094_), .ZN(new_n6095_));
  AOI22_X1   g05903(.A1(new_n6095_), .A2(new_n5691_), .B1(\asqrt[34] ), .B2(new_n6093_), .ZN(new_n6096_));
  OAI21_X1   g05904(.A1(new_n6080_), .A2(new_n6081_), .B(new_n6071_), .ZN(new_n6097_));
  AOI21_X1   g05905(.A1(new_n6097_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n6098_));
  AOI21_X1   g05906(.A1(new_n6098_), .A2(new_n6091_), .B(new_n6096_), .ZN(new_n6099_));
  OAI21_X1   g05907(.A1(new_n6099_), .A2(new_n6092_), .B(\asqrt[41] ), .ZN(new_n6100_));
  NAND2_X1   g05908(.A1(new_n5890_), .A2(new_n5882_), .ZN(new_n6101_));
  NAND3_X1   g05909(.A1(\asqrt[34] ), .A2(new_n5695_), .A3(new_n6101_), .ZN(new_n6102_));
  AND3_X2    g05910(.A1(new_n5695_), .A2(new_n5701_), .A3(new_n6101_), .Z(new_n6103_));
  AOI22_X1   g05911(.A1(new_n6102_), .A2(new_n5702_), .B1(\asqrt[34] ), .B2(new_n6103_), .ZN(new_n6104_));
  INV_X1     g05912(.I(new_n6104_), .ZN(new_n6105_));
  NAND2_X1   g05913(.A1(new_n6036_), .A2(new_n6041_), .ZN(new_n6106_));
  OAI21_X1   g05914(.A1(new_n6033_), .A2(new_n6035_), .B(new_n6038_), .ZN(new_n6107_));
  NAND2_X1   g05915(.A1(new_n6107_), .A2(\a[69] ), .ZN(new_n6108_));
  NAND3_X1   g05916(.A1(new_n6106_), .A2(new_n6108_), .A3(new_n6049_), .ZN(new_n6109_));
  AOI21_X1   g05917(.A1(new_n6109_), .A2(new_n6059_), .B(new_n5277_), .ZN(new_n6110_));
  OAI21_X1   g05918(.A1(new_n6057_), .A2(new_n6044_), .B(\a[70] ), .ZN(new_n6111_));
  NAND3_X1   g05919(.A1(new_n6053_), .A2(new_n6049_), .A3(new_n5644_), .ZN(new_n6112_));
  NAND2_X1   g05920(.A1(new_n6036_), .A2(new_n6021_), .ZN(new_n6113_));
  AOI21_X1   g05921(.A1(new_n6113_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n6114_));
  AOI22_X1   g05922(.A1(new_n6109_), .A2(new_n6114_), .B1(new_n6111_), .B2(new_n6112_), .ZN(new_n6115_));
  OAI21_X1   g05923(.A1(new_n6115_), .A2(new_n6110_), .B(\asqrt[37] ), .ZN(new_n6116_));
  NAND2_X1   g05924(.A1(new_n6116_), .A2(new_n4696_), .ZN(new_n6117_));
  OAI21_X1   g05925(.A1(new_n6117_), .A2(new_n6070_), .B(new_n6079_), .ZN(new_n6118_));
  AOI21_X1   g05926(.A1(new_n6118_), .A2(new_n6071_), .B(new_n4298_), .ZN(new_n6119_));
  INV_X1     g05927(.I(new_n6065_), .ZN(new_n6120_));
  AOI21_X1   g05928(.A1(\a[69] ), .A2(new_n6107_), .B(new_n6044_), .ZN(new_n6121_));
  AOI21_X1   g05929(.A1(new_n6121_), .A2(new_n6106_), .B(new_n6037_), .ZN(new_n6122_));
  OAI21_X1   g05930(.A1(new_n6122_), .A2(new_n5277_), .B(new_n5024_), .ZN(new_n6123_));
  OAI21_X1   g05931(.A1(new_n6123_), .A2(new_n6115_), .B(new_n6120_), .ZN(new_n6124_));
  NAND2_X1   g05932(.A1(new_n6124_), .A2(new_n6116_), .ZN(new_n6125_));
  AOI21_X1   g05933(.A1(new_n6125_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n6126_));
  AOI21_X1   g05934(.A1(new_n6126_), .A2(new_n6118_), .B(new_n6088_), .ZN(new_n6127_));
  OAI21_X1   g05935(.A1(new_n6127_), .A2(new_n6119_), .B(\asqrt[40] ), .ZN(new_n6128_));
  NAND2_X1   g05936(.A1(new_n6128_), .A2(new_n3782_), .ZN(new_n6129_));
  OAI21_X1   g05937(.A1(new_n6129_), .A2(new_n6099_), .B(new_n6105_), .ZN(new_n6130_));
  AOI21_X1   g05938(.A1(new_n6130_), .A2(new_n6100_), .B(new_n3419_), .ZN(new_n6131_));
  INV_X1     g05939(.I(new_n5711_), .ZN(new_n6132_));
  NOR3_X1    g05940(.A1(new_n5705_), .A2(new_n5901_), .A3(new_n6132_), .ZN(new_n6133_));
  NOR3_X1    g05941(.A1(new_n6077_), .A2(new_n5705_), .A3(new_n5901_), .ZN(new_n6134_));
  INV_X1     g05942(.I(new_n6134_), .ZN(new_n6135_));
  AOI22_X1   g05943(.A1(new_n6135_), .A2(new_n6132_), .B1(\asqrt[34] ), .B2(new_n6133_), .ZN(new_n6136_));
  NOR3_X1    g05944(.A1(new_n6127_), .A2(new_n6119_), .A3(\asqrt[40] ), .ZN(new_n6137_));
  OAI21_X1   g05945(.A1(new_n6096_), .A2(new_n6137_), .B(new_n6128_), .ZN(new_n6138_));
  AOI21_X1   g05946(.A1(new_n6138_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n6139_));
  AOI21_X1   g05947(.A1(new_n6139_), .A2(new_n6130_), .B(new_n6136_), .ZN(new_n6140_));
  OAI21_X1   g05948(.A1(new_n6140_), .A2(new_n6131_), .B(\asqrt[43] ), .ZN(new_n6141_));
  INV_X1     g05949(.I(new_n6141_), .ZN(new_n6142_));
  NOR3_X1    g05950(.A1(new_n6077_), .A2(new_n5716_), .A3(new_n5723_), .ZN(new_n6143_));
  INV_X1     g05951(.I(new_n6143_), .ZN(new_n6144_));
  NOR3_X1    g05952(.A1(new_n5716_), .A2(new_n5869_), .A3(new_n5723_), .ZN(new_n6145_));
  AOI22_X1   g05953(.A1(new_n6144_), .A2(new_n5869_), .B1(\asqrt[34] ), .B2(new_n6145_), .ZN(new_n6146_));
  NOR3_X1    g05954(.A1(new_n6140_), .A2(\asqrt[43] ), .A3(new_n6131_), .ZN(new_n6147_));
  NOR2_X1    g05955(.A1(new_n6147_), .A2(new_n6146_), .ZN(new_n6148_));
  OAI21_X1   g05956(.A1(new_n6148_), .A2(new_n6142_), .B(\asqrt[44] ), .ZN(new_n6149_));
  INV_X1     g05957(.I(new_n5895_), .ZN(new_n6150_));
  NOR3_X1    g05958(.A1(new_n6150_), .A2(new_n5900_), .A3(new_n5734_), .ZN(new_n6151_));
  NOR3_X1    g05959(.A1(new_n6077_), .A2(new_n5900_), .A3(new_n6150_), .ZN(new_n6152_));
  INV_X1     g05960(.I(new_n6152_), .ZN(new_n6153_));
  AOI22_X1   g05961(.A1(new_n6153_), .A2(new_n5734_), .B1(\asqrt[34] ), .B2(new_n6151_), .ZN(new_n6154_));
  INV_X1     g05962(.I(new_n6154_), .ZN(new_n6155_));
  NAND2_X1   g05963(.A1(new_n6141_), .A2(new_n2954_), .ZN(new_n6156_));
  OAI21_X1   g05964(.A1(new_n6148_), .A2(new_n6156_), .B(new_n6155_), .ZN(new_n6157_));
  AOI21_X1   g05965(.A1(new_n6157_), .A2(new_n6149_), .B(new_n2641_), .ZN(new_n6158_));
  INV_X1     g05966(.I(new_n5742_), .ZN(new_n6159_));
  NOR3_X1    g05967(.A1(new_n6077_), .A2(new_n5737_), .A3(new_n5905_), .ZN(new_n6160_));
  INV_X1     g05968(.I(new_n6160_), .ZN(new_n6161_));
  NOR3_X1    g05969(.A1(new_n5737_), .A2(new_n5905_), .A3(new_n6159_), .ZN(new_n6162_));
  AOI22_X1   g05970(.A1(new_n6161_), .A2(new_n6159_), .B1(\asqrt[34] ), .B2(new_n6162_), .ZN(new_n6163_));
  NOR3_X1    g05971(.A1(new_n6099_), .A2(new_n6092_), .A3(\asqrt[41] ), .ZN(new_n6164_));
  OAI21_X1   g05972(.A1(new_n6104_), .A2(new_n6164_), .B(new_n6100_), .ZN(new_n6165_));
  INV_X1     g05973(.I(new_n6136_), .ZN(new_n6166_));
  NAND3_X1   g05974(.A1(new_n6130_), .A2(new_n3419_), .A3(new_n6100_), .ZN(new_n6167_));
  AOI22_X1   g05975(.A1(new_n6167_), .A2(new_n6166_), .B1(new_n6165_), .B2(\asqrt[42] ), .ZN(new_n6168_));
  OAI22_X1   g05976(.A1(new_n6147_), .A2(new_n6146_), .B1(new_n6168_), .B2(new_n3218_), .ZN(new_n6169_));
  AOI21_X1   g05977(.A1(new_n6169_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n6170_));
  AOI21_X1   g05978(.A1(new_n6170_), .A2(new_n6157_), .B(new_n6163_), .ZN(new_n6171_));
  OAI21_X1   g05979(.A1(new_n6171_), .A2(new_n6158_), .B(\asqrt[46] ), .ZN(new_n6172_));
  INV_X1     g05980(.I(new_n6172_), .ZN(new_n6173_));
  NOR3_X1    g05981(.A1(new_n5747_), .A2(new_n5868_), .A3(new_n5753_), .ZN(new_n6174_));
  NOR3_X1    g05982(.A1(new_n6077_), .A2(new_n5747_), .A3(new_n5753_), .ZN(new_n6175_));
  INV_X1     g05983(.I(new_n6175_), .ZN(new_n6176_));
  AOI22_X1   g05984(.A1(new_n6176_), .A2(new_n5868_), .B1(\asqrt[34] ), .B2(new_n6174_), .ZN(new_n6177_));
  NOR3_X1    g05985(.A1(new_n6171_), .A2(new_n6158_), .A3(\asqrt[46] ), .ZN(new_n6178_));
  NOR2_X1    g05986(.A1(new_n6178_), .A2(new_n6177_), .ZN(new_n6179_));
  OAI21_X1   g05987(.A1(new_n6179_), .A2(new_n6173_), .B(\asqrt[47] ), .ZN(new_n6180_));
  NOR2_X1    g05988(.A1(new_n5754_), .A2(new_n5765_), .ZN(new_n6181_));
  NOR3_X1    g05989(.A1(new_n6077_), .A2(new_n5899_), .A3(new_n6181_), .ZN(new_n6182_));
  INV_X1     g05990(.I(new_n6182_), .ZN(new_n6183_));
  NOR3_X1    g05991(.A1(new_n6181_), .A2(new_n5899_), .A3(new_n5764_), .ZN(new_n6184_));
  AOI22_X1   g05992(.A1(new_n6183_), .A2(new_n5764_), .B1(\asqrt[34] ), .B2(new_n6184_), .ZN(new_n6185_));
  INV_X1     g05993(.I(new_n6185_), .ZN(new_n6186_));
  NAND2_X1   g05994(.A1(new_n6172_), .A2(new_n2229_), .ZN(new_n6187_));
  OAI21_X1   g05995(.A1(new_n6179_), .A2(new_n6187_), .B(new_n6186_), .ZN(new_n6188_));
  AOI21_X1   g05996(.A1(new_n6188_), .A2(new_n6180_), .B(new_n1956_), .ZN(new_n6189_));
  INV_X1     g05997(.I(new_n5772_), .ZN(new_n6190_));
  NOR3_X1    g05998(.A1(new_n5767_), .A2(new_n5913_), .A3(new_n6190_), .ZN(new_n6191_));
  NOR3_X1    g05999(.A1(new_n6077_), .A2(new_n5767_), .A3(new_n5913_), .ZN(new_n6192_));
  INV_X1     g06000(.I(new_n6192_), .ZN(new_n6193_));
  AOI22_X1   g06001(.A1(new_n6193_), .A2(new_n6190_), .B1(\asqrt[34] ), .B2(new_n6191_), .ZN(new_n6194_));
  OAI21_X1   g06002(.A1(new_n6177_), .A2(new_n6178_), .B(new_n6172_), .ZN(new_n6195_));
  AOI21_X1   g06003(.A1(new_n6195_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n6196_));
  AOI21_X1   g06004(.A1(new_n6196_), .A2(new_n6188_), .B(new_n6194_), .ZN(new_n6197_));
  OAI21_X1   g06005(.A1(new_n6197_), .A2(new_n6189_), .B(\asqrt[49] ), .ZN(new_n6198_));
  INV_X1     g06006(.I(new_n6198_), .ZN(new_n6199_));
  NOR3_X1    g06007(.A1(new_n6077_), .A2(new_n5777_), .A3(new_n5784_), .ZN(new_n6200_));
  INV_X1     g06008(.I(new_n6200_), .ZN(new_n6201_));
  NOR3_X1    g06009(.A1(new_n5777_), .A2(new_n5867_), .A3(new_n5784_), .ZN(new_n6202_));
  AOI22_X1   g06010(.A1(new_n6201_), .A2(new_n5867_), .B1(\asqrt[34] ), .B2(new_n6202_), .ZN(new_n6203_));
  NOR3_X1    g06011(.A1(new_n6197_), .A2(new_n6189_), .A3(\asqrt[49] ), .ZN(new_n6204_));
  NOR2_X1    g06012(.A1(new_n6204_), .A2(new_n6203_), .ZN(new_n6205_));
  OAI21_X1   g06013(.A1(new_n6205_), .A2(new_n6199_), .B(\asqrt[50] ), .ZN(new_n6206_));
  NOR2_X1    g06014(.A1(new_n5785_), .A2(new_n5796_), .ZN(new_n6207_));
  NOR3_X1    g06015(.A1(new_n6207_), .A2(new_n5912_), .A3(new_n5795_), .ZN(new_n6208_));
  NOR3_X1    g06016(.A1(new_n6077_), .A2(new_n5912_), .A3(new_n6207_), .ZN(new_n6209_));
  INV_X1     g06017(.I(new_n6209_), .ZN(new_n6210_));
  AOI22_X1   g06018(.A1(new_n6210_), .A2(new_n5795_), .B1(\asqrt[34] ), .B2(new_n6208_), .ZN(new_n6211_));
  INV_X1     g06019(.I(new_n6211_), .ZN(new_n6212_));
  NAND2_X1   g06020(.A1(new_n6198_), .A2(new_n1612_), .ZN(new_n6213_));
  OAI21_X1   g06021(.A1(new_n6205_), .A2(new_n6213_), .B(new_n6212_), .ZN(new_n6214_));
  AOI21_X1   g06022(.A1(new_n6214_), .A2(new_n6206_), .B(new_n1376_), .ZN(new_n6215_));
  INV_X1     g06023(.I(new_n5802_), .ZN(new_n6216_));
  NOR3_X1    g06024(.A1(new_n6077_), .A2(new_n5798_), .A3(new_n5921_), .ZN(new_n6217_));
  INV_X1     g06025(.I(new_n6217_), .ZN(new_n6218_));
  NOR3_X1    g06026(.A1(new_n5798_), .A2(new_n5921_), .A3(new_n6216_), .ZN(new_n6219_));
  AOI22_X1   g06027(.A1(new_n6218_), .A2(new_n6216_), .B1(\asqrt[34] ), .B2(new_n6219_), .ZN(new_n6220_));
  OAI21_X1   g06028(.A1(new_n6203_), .A2(new_n6204_), .B(new_n6198_), .ZN(new_n6221_));
  AOI21_X1   g06029(.A1(new_n6221_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n6222_));
  AOI21_X1   g06030(.A1(new_n6222_), .A2(new_n6214_), .B(new_n6220_), .ZN(new_n6223_));
  OAI21_X1   g06031(.A1(new_n6223_), .A2(new_n6215_), .B(\asqrt[52] ), .ZN(new_n6224_));
  INV_X1     g06032(.I(new_n6224_), .ZN(new_n6225_));
  INV_X1     g06033(.I(new_n6223_), .ZN(new_n6226_));
  NOR3_X1    g06034(.A1(new_n5807_), .A2(new_n5866_), .A3(new_n5813_), .ZN(new_n6227_));
  NOR3_X1    g06035(.A1(new_n6077_), .A2(new_n5807_), .A3(new_n5813_), .ZN(new_n6228_));
  INV_X1     g06036(.I(new_n6228_), .ZN(new_n6229_));
  AOI22_X1   g06037(.A1(new_n6229_), .A2(new_n5866_), .B1(\asqrt[34] ), .B2(new_n6227_), .ZN(new_n6230_));
  NOR2_X1    g06038(.A1(new_n6215_), .A2(\asqrt[52] ), .ZN(new_n6231_));
  AOI21_X1   g06039(.A1(new_n6226_), .A2(new_n6231_), .B(new_n6230_), .ZN(new_n6232_));
  OAI21_X1   g06040(.A1(new_n6232_), .A2(new_n6225_), .B(\asqrt[53] ), .ZN(new_n6233_));
  NOR2_X1    g06041(.A1(new_n5814_), .A2(new_n5822_), .ZN(new_n6234_));
  NOR3_X1    g06042(.A1(new_n6077_), .A2(new_n5920_), .A3(new_n6234_), .ZN(new_n6235_));
  INV_X1     g06043(.I(new_n6235_), .ZN(new_n6236_));
  NOR3_X1    g06044(.A1(new_n6234_), .A2(new_n5920_), .A3(new_n5821_), .ZN(new_n6237_));
  AOI22_X1   g06045(.A1(new_n6236_), .A2(new_n5821_), .B1(\asqrt[34] ), .B2(new_n6237_), .ZN(new_n6238_));
  INV_X1     g06046(.I(new_n6238_), .ZN(new_n6239_));
  NAND2_X1   g06047(.A1(new_n6224_), .A2(new_n1103_), .ZN(new_n6240_));
  OAI21_X1   g06048(.A1(new_n6240_), .A2(new_n6232_), .B(new_n6239_), .ZN(new_n6241_));
  AOI21_X1   g06049(.A1(new_n6241_), .A2(new_n6233_), .B(new_n904_), .ZN(new_n6242_));
  INV_X1     g06050(.I(new_n6242_), .ZN(new_n6243_));
  INV_X1     g06051(.I(new_n6241_), .ZN(new_n6244_));
  INV_X1     g06052(.I(new_n5828_), .ZN(new_n6245_));
  NOR3_X1    g06053(.A1(new_n5824_), .A2(new_n5929_), .A3(new_n6245_), .ZN(new_n6246_));
  NOR3_X1    g06054(.A1(new_n6077_), .A2(new_n5824_), .A3(new_n5929_), .ZN(new_n6247_));
  INV_X1     g06055(.I(new_n6247_), .ZN(new_n6248_));
  AOI22_X1   g06056(.A1(new_n6248_), .A2(new_n6245_), .B1(\asqrt[34] ), .B2(new_n6246_), .ZN(new_n6249_));
  INV_X1     g06057(.I(new_n6249_), .ZN(new_n6250_));
  NAND2_X1   g06058(.A1(new_n6233_), .A2(new_n904_), .ZN(new_n6251_));
  OAI21_X1   g06059(.A1(new_n6251_), .A2(new_n6244_), .B(new_n6250_), .ZN(new_n6252_));
  AOI21_X1   g06060(.A1(new_n6252_), .A2(new_n6243_), .B(new_n823_), .ZN(new_n6253_));
  NOR3_X1    g06061(.A1(new_n6077_), .A2(new_n5833_), .A3(new_n5839_), .ZN(new_n6254_));
  INV_X1     g06062(.I(new_n6254_), .ZN(new_n6255_));
  NOR3_X1    g06063(.A1(new_n5833_), .A2(new_n5839_), .A3(new_n5865_), .ZN(new_n6256_));
  AOI22_X1   g06064(.A1(new_n6255_), .A2(new_n5865_), .B1(\asqrt[34] ), .B2(new_n6256_), .ZN(new_n6257_));
  NOR2_X1    g06065(.A1(new_n6242_), .A2(\asqrt[55] ), .ZN(new_n6258_));
  AOI21_X1   g06066(.A1(new_n6258_), .A2(new_n6252_), .B(new_n6257_), .ZN(new_n6259_));
  OAI21_X1   g06067(.A1(new_n6259_), .A2(new_n6253_), .B(\asqrt[56] ), .ZN(new_n6260_));
  NOR2_X1    g06068(.A1(new_n5840_), .A2(new_n5848_), .ZN(new_n6261_));
  NOR3_X1    g06069(.A1(new_n6261_), .A2(new_n5928_), .A3(new_n5847_), .ZN(new_n6262_));
  NOR3_X1    g06070(.A1(new_n6077_), .A2(new_n5928_), .A3(new_n6261_), .ZN(new_n6263_));
  INV_X1     g06071(.I(new_n6263_), .ZN(new_n6264_));
  AOI22_X1   g06072(.A1(new_n6264_), .A2(new_n5847_), .B1(\asqrt[34] ), .B2(new_n6262_), .ZN(new_n6265_));
  INV_X1     g06073(.I(new_n6265_), .ZN(new_n6266_));
  NOR3_X1    g06074(.A1(new_n6223_), .A2(new_n6215_), .A3(\asqrt[52] ), .ZN(new_n6267_));
  OAI21_X1   g06075(.A1(new_n6230_), .A2(new_n6267_), .B(new_n6224_), .ZN(new_n6268_));
  AOI21_X1   g06076(.A1(new_n6268_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n6269_));
  AOI21_X1   g06077(.A1(new_n6269_), .A2(new_n6241_), .B(new_n6249_), .ZN(new_n6270_));
  OAI21_X1   g06078(.A1(new_n6270_), .A2(new_n6242_), .B(\asqrt[55] ), .ZN(new_n6271_));
  NAND2_X1   g06079(.A1(new_n6271_), .A2(new_n703_), .ZN(new_n6272_));
  OAI21_X1   g06080(.A1(new_n6272_), .A2(new_n6259_), .B(new_n6266_), .ZN(new_n6273_));
  AOI21_X1   g06081(.A1(new_n6273_), .A2(new_n6260_), .B(new_n531_), .ZN(new_n6274_));
  INV_X1     g06082(.I(new_n6274_), .ZN(new_n6275_));
  INV_X1     g06083(.I(new_n6273_), .ZN(new_n6276_));
  INV_X1     g06084(.I(new_n5854_), .ZN(new_n6277_));
  NOR3_X1    g06085(.A1(new_n6077_), .A2(new_n5850_), .A3(new_n5942_), .ZN(new_n6278_));
  INV_X1     g06086(.I(new_n6278_), .ZN(new_n6279_));
  NOR3_X1    g06087(.A1(new_n5850_), .A2(new_n5942_), .A3(new_n6277_), .ZN(new_n6280_));
  AOI22_X1   g06088(.A1(new_n6279_), .A2(new_n6277_), .B1(\asqrt[34] ), .B2(new_n6280_), .ZN(new_n6281_));
  INV_X1     g06089(.I(new_n6281_), .ZN(new_n6282_));
  NAND2_X1   g06090(.A1(new_n6260_), .A2(new_n531_), .ZN(new_n6283_));
  OAI21_X1   g06091(.A1(new_n6283_), .A2(new_n6276_), .B(new_n6282_), .ZN(new_n6284_));
  AOI21_X1   g06092(.A1(new_n6284_), .A2(new_n6275_), .B(new_n436_), .ZN(new_n6285_));
  NOR3_X1    g06093(.A1(new_n5952_), .A2(new_n5953_), .A3(new_n5864_), .ZN(new_n6286_));
  NOR3_X1    g06094(.A1(new_n6077_), .A2(new_n5952_), .A3(new_n5953_), .ZN(new_n6287_));
  INV_X1     g06095(.I(new_n6287_), .ZN(new_n6288_));
  AOI22_X1   g06096(.A1(new_n6288_), .A2(new_n5864_), .B1(\asqrt[34] ), .B2(new_n6286_), .ZN(new_n6289_));
  NOR2_X1    g06097(.A1(new_n6274_), .A2(\asqrt[58] ), .ZN(new_n6290_));
  AOI21_X1   g06098(.A1(new_n6290_), .A2(new_n6284_), .B(new_n6289_), .ZN(new_n6291_));
  OAI21_X1   g06099(.A1(new_n6291_), .A2(new_n6285_), .B(\asqrt[59] ), .ZN(new_n6292_));
  NOR2_X1    g06100(.A1(new_n5954_), .A2(new_n5965_), .ZN(new_n6293_));
  NOR3_X1    g06101(.A1(new_n6077_), .A2(new_n5936_), .A3(new_n6293_), .ZN(new_n6294_));
  INV_X1     g06102(.I(new_n6294_), .ZN(new_n6295_));
  NOR3_X1    g06103(.A1(new_n6293_), .A2(new_n5936_), .A3(new_n5964_), .ZN(new_n6296_));
  AOI22_X1   g06104(.A1(new_n6295_), .A2(new_n5964_), .B1(\asqrt[34] ), .B2(new_n6296_), .ZN(new_n6297_));
  INV_X1     g06105(.I(new_n6297_), .ZN(new_n6298_));
  NOR3_X1    g06106(.A1(new_n6270_), .A2(\asqrt[55] ), .A3(new_n6242_), .ZN(new_n6299_));
  OAI21_X1   g06107(.A1(new_n6257_), .A2(new_n6299_), .B(new_n6271_), .ZN(new_n6300_));
  AOI21_X1   g06108(.A1(new_n6300_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n6301_));
  AOI21_X1   g06109(.A1(new_n6301_), .A2(new_n6273_), .B(new_n6281_), .ZN(new_n6302_));
  OAI21_X1   g06110(.A1(new_n6302_), .A2(new_n6274_), .B(\asqrt[58] ), .ZN(new_n6303_));
  NAND2_X1   g06111(.A1(new_n6303_), .A2(new_n327_), .ZN(new_n6304_));
  OAI21_X1   g06112(.A1(new_n6304_), .A2(new_n6291_), .B(new_n6298_), .ZN(new_n6305_));
  AOI21_X1   g06113(.A1(new_n6305_), .A2(new_n6292_), .B(new_n306_), .ZN(new_n6306_));
  INV_X1     g06114(.I(new_n6306_), .ZN(new_n6307_));
  INV_X1     g06115(.I(new_n6305_), .ZN(new_n6308_));
  NOR3_X1    g06116(.A1(new_n5967_), .A2(new_n6026_), .A3(new_n5951_), .ZN(new_n6309_));
  NOR3_X1    g06117(.A1(new_n6077_), .A2(new_n5967_), .A3(new_n6026_), .ZN(new_n6310_));
  INV_X1     g06118(.I(new_n6310_), .ZN(new_n6311_));
  AOI22_X1   g06119(.A1(new_n6311_), .A2(new_n5951_), .B1(\asqrt[34] ), .B2(new_n6309_), .ZN(new_n6312_));
  INV_X1     g06120(.I(new_n6312_), .ZN(new_n6313_));
  NAND2_X1   g06121(.A1(new_n6292_), .A2(new_n306_), .ZN(new_n6314_));
  OAI21_X1   g06122(.A1(new_n6308_), .A2(new_n6314_), .B(new_n6313_), .ZN(new_n6315_));
  AOI21_X1   g06123(.A1(new_n6315_), .A2(new_n6307_), .B(new_n218_), .ZN(new_n6316_));
  NOR3_X1    g06124(.A1(new_n6077_), .A2(new_n5958_), .A3(new_n5988_), .ZN(new_n6317_));
  INV_X1     g06125(.I(new_n6317_), .ZN(new_n6318_));
  NOR3_X1    g06126(.A1(new_n5958_), .A2(new_n5988_), .A3(new_n6022_), .ZN(new_n6319_));
  AOI22_X1   g06127(.A1(new_n6318_), .A2(new_n6022_), .B1(\asqrt[34] ), .B2(new_n6319_), .ZN(new_n6320_));
  NOR2_X1    g06128(.A1(new_n6306_), .A2(\asqrt[61] ), .ZN(new_n6321_));
  AOI21_X1   g06129(.A1(new_n6321_), .A2(new_n6315_), .B(new_n6320_), .ZN(new_n6322_));
  OAI21_X1   g06130(.A1(new_n6322_), .A2(new_n6316_), .B(\asqrt[62] ), .ZN(new_n6323_));
  NOR2_X1    g06131(.A1(new_n5981_), .A2(new_n5969_), .ZN(new_n6324_));
  NOR3_X1    g06132(.A1(new_n6324_), .A2(new_n6025_), .A3(new_n5976_), .ZN(new_n6325_));
  NOR3_X1    g06133(.A1(new_n6077_), .A2(new_n6025_), .A3(new_n6324_), .ZN(new_n6326_));
  INV_X1     g06134(.I(new_n6326_), .ZN(new_n6327_));
  AOI22_X1   g06135(.A1(new_n6327_), .A2(new_n5976_), .B1(\asqrt[34] ), .B2(new_n6325_), .ZN(new_n6328_));
  INV_X1     g06136(.I(new_n6328_), .ZN(new_n6329_));
  NOR3_X1    g06137(.A1(new_n6302_), .A2(\asqrt[58] ), .A3(new_n6274_), .ZN(new_n6330_));
  OAI21_X1   g06138(.A1(new_n6289_), .A2(new_n6330_), .B(new_n6303_), .ZN(new_n6331_));
  AOI21_X1   g06139(.A1(new_n6331_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n6332_));
  AOI21_X1   g06140(.A1(new_n6332_), .A2(new_n6305_), .B(new_n6312_), .ZN(new_n6333_));
  OAI21_X1   g06141(.A1(new_n6333_), .A2(new_n6306_), .B(\asqrt[61] ), .ZN(new_n6334_));
  NAND2_X1   g06142(.A1(new_n6334_), .A2(new_n207_), .ZN(new_n6335_));
  OAI21_X1   g06143(.A1(new_n6335_), .A2(new_n6322_), .B(new_n6329_), .ZN(new_n6336_));
  NAND4_X1   g06144(.A1(\asqrt[34] ), .A2(new_n6030_), .A3(new_n5987_), .A4(new_n6003_), .ZN(new_n6337_));
  NAND2_X1   g06145(.A1(new_n6030_), .A2(new_n6003_), .ZN(new_n6338_));
  OAI21_X1   g06146(.A1(new_n6077_), .A2(new_n6338_), .B(new_n6002_), .ZN(new_n6339_));
  NAND2_X1   g06147(.A1(new_n6339_), .A2(new_n6337_), .ZN(new_n6340_));
  AOI21_X1   g06148(.A1(new_n6004_), .A2(new_n6030_), .B(new_n5997_), .ZN(new_n6341_));
  AOI21_X1   g06149(.A1(\asqrt[34] ), .A2(new_n6341_), .B(new_n6055_), .ZN(new_n6342_));
  NAND2_X1   g06150(.A1(new_n6340_), .A2(new_n6342_), .ZN(new_n6343_));
  AOI21_X1   g06151(.A1(new_n6336_), .A2(new_n6323_), .B(new_n6343_), .ZN(new_n6344_));
  NOR3_X1    g06152(.A1(new_n6333_), .A2(\asqrt[61] ), .A3(new_n6306_), .ZN(new_n6345_));
  OAI21_X1   g06153(.A1(new_n6320_), .A2(new_n6345_), .B(new_n6334_), .ZN(new_n6346_));
  AOI21_X1   g06154(.A1(new_n6346_), .A2(\asqrt[62] ), .B(new_n6340_), .ZN(new_n6347_));
  AOI21_X1   g06155(.A1(\asqrt[34] ), .A2(new_n6005_), .B(new_n6032_), .ZN(new_n6348_));
  OR3_X2     g06156(.A1(new_n6348_), .A2(new_n193_), .A3(new_n6341_), .Z(new_n6349_));
  NAND2_X1   g06157(.A1(new_n5993_), .A2(new_n6012_), .ZN(new_n6350_));
  NOR4_X1    g06158(.A1(new_n6055_), .A2(new_n5996_), .A3(new_n6009_), .A4(new_n6350_), .ZN(new_n6351_));
  NAND2_X1   g06159(.A1(new_n6351_), .A2(new_n6001_), .ZN(new_n6352_));
  NAND2_X1   g06160(.A1(new_n6349_), .A2(new_n6352_), .ZN(new_n6353_));
  AOI21_X1   g06161(.A1(new_n6347_), .A2(new_n6336_), .B(new_n6353_), .ZN(new_n6354_));
  OAI21_X1   g06162(.A1(\asqrt[63] ), .A2(new_n6344_), .B(new_n6354_), .ZN(\asqrt[33] ));
  INV_X1     g06163(.I(\asqrt[33] ), .ZN(new_n6356_));
  NOR2_X1    g06164(.A1(\a[64] ), .A2(\a[65] ), .ZN(new_n6357_));
  INV_X1     g06165(.I(new_n6357_), .ZN(new_n6358_));
  NOR2_X1    g06166(.A1(new_n6358_), .A2(\a[66] ), .ZN(new_n6359_));
  INV_X1     g06167(.I(\a[66] ), .ZN(new_n6360_));
  INV_X1     g06168(.I(new_n6320_), .ZN(new_n6361_));
  INV_X1     g06169(.I(new_n6289_), .ZN(new_n6362_));
  INV_X1     g06170(.I(new_n6257_), .ZN(new_n6363_));
  INV_X1     g06171(.I(new_n6230_), .ZN(new_n6364_));
  INV_X1     g06172(.I(new_n6203_), .ZN(new_n6365_));
  INV_X1     g06173(.I(new_n6177_), .ZN(new_n6366_));
  INV_X1     g06174(.I(new_n6146_), .ZN(new_n6367_));
  INV_X1     g06175(.I(new_n6100_), .ZN(new_n6368_));
  NOR2_X1    g06176(.A1(new_n6164_), .A2(new_n6104_), .ZN(new_n6369_));
  OAI21_X1   g06177(.A1(new_n6369_), .A2(new_n6368_), .B(\asqrt[42] ), .ZN(new_n6370_));
  NAND2_X1   g06178(.A1(new_n6370_), .A2(new_n3218_), .ZN(new_n6371_));
  OAI21_X1   g06179(.A1(new_n6371_), .A2(new_n6140_), .B(new_n6367_), .ZN(new_n6372_));
  NAND3_X1   g06180(.A1(new_n6372_), .A2(new_n2954_), .A3(new_n6141_), .ZN(new_n6373_));
  AOI22_X1   g06181(.A1(new_n6373_), .A2(new_n6155_), .B1(\asqrt[44] ), .B2(new_n6169_), .ZN(new_n6374_));
  OAI21_X1   g06182(.A1(new_n6374_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n6375_));
  OAI21_X1   g06183(.A1(new_n6375_), .A2(new_n6171_), .B(new_n6366_), .ZN(new_n6376_));
  NAND3_X1   g06184(.A1(new_n6376_), .A2(new_n2229_), .A3(new_n6172_), .ZN(new_n6377_));
  AOI22_X1   g06185(.A1(new_n6377_), .A2(new_n6186_), .B1(\asqrt[47] ), .B2(new_n6195_), .ZN(new_n6378_));
  OAI21_X1   g06186(.A1(new_n6378_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n6379_));
  OAI21_X1   g06187(.A1(new_n6379_), .A2(new_n6197_), .B(new_n6365_), .ZN(new_n6380_));
  NAND3_X1   g06188(.A1(new_n6380_), .A2(new_n1612_), .A3(new_n6198_), .ZN(new_n6381_));
  AOI22_X1   g06189(.A1(new_n6381_), .A2(new_n6212_), .B1(\asqrt[50] ), .B2(new_n6221_), .ZN(new_n6382_));
  OAI21_X1   g06190(.A1(new_n6382_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n6383_));
  OAI21_X1   g06191(.A1(new_n6383_), .A2(new_n6223_), .B(new_n6364_), .ZN(new_n6384_));
  NAND3_X1   g06192(.A1(new_n6384_), .A2(new_n1103_), .A3(new_n6224_), .ZN(new_n6385_));
  AOI22_X1   g06193(.A1(new_n6385_), .A2(new_n6239_), .B1(\asqrt[53] ), .B2(new_n6268_), .ZN(new_n6386_));
  OAI21_X1   g06194(.A1(new_n6386_), .A2(new_n904_), .B(new_n823_), .ZN(new_n6387_));
  OAI21_X1   g06195(.A1(new_n6387_), .A2(new_n6270_), .B(new_n6363_), .ZN(new_n6388_));
  NAND3_X1   g06196(.A1(new_n6388_), .A2(new_n703_), .A3(new_n6271_), .ZN(new_n6389_));
  AOI22_X1   g06197(.A1(new_n6389_), .A2(new_n6266_), .B1(\asqrt[56] ), .B2(new_n6300_), .ZN(new_n6390_));
  OAI21_X1   g06198(.A1(new_n6390_), .A2(new_n531_), .B(new_n436_), .ZN(new_n6391_));
  OAI21_X1   g06199(.A1(new_n6391_), .A2(new_n6302_), .B(new_n6362_), .ZN(new_n6392_));
  NAND3_X1   g06200(.A1(new_n6392_), .A2(new_n327_), .A3(new_n6303_), .ZN(new_n6393_));
  AOI22_X1   g06201(.A1(new_n6393_), .A2(new_n6298_), .B1(new_n6331_), .B2(\asqrt[59] ), .ZN(new_n6394_));
  OAI21_X1   g06202(.A1(new_n6394_), .A2(new_n306_), .B(new_n218_), .ZN(new_n6395_));
  OAI21_X1   g06203(.A1(new_n6395_), .A2(new_n6333_), .B(new_n6361_), .ZN(new_n6396_));
  NAND3_X1   g06204(.A1(new_n6396_), .A2(new_n207_), .A3(new_n6334_), .ZN(new_n6397_));
  AOI22_X1   g06205(.A1(new_n6397_), .A2(new_n6329_), .B1(new_n6346_), .B2(\asqrt[62] ), .ZN(new_n6398_));
  OAI21_X1   g06206(.A1(new_n6398_), .A2(new_n6343_), .B(new_n193_), .ZN(new_n6399_));
  AOI21_X1   g06207(.A1(new_n6399_), .A2(new_n6354_), .B(new_n6360_), .ZN(new_n6400_));
  OAI21_X1   g06208(.A1(new_n6400_), .A2(new_n6359_), .B(\asqrt[34] ), .ZN(new_n6401_));
  INV_X1     g06209(.I(new_n6401_), .ZN(new_n6402_));
  OAI21_X1   g06210(.A1(\a[66] ), .A2(new_n6358_), .B(new_n6012_), .ZN(new_n6403_));
  NOR4_X1    g06211(.A1(new_n6055_), .A2(new_n6033_), .A3(new_n6009_), .A4(new_n6403_), .ZN(new_n6404_));
  INV_X1     g06212(.I(new_n6404_), .ZN(new_n6405_));
  NOR2_X1    g06213(.A1(new_n6400_), .A2(new_n6405_), .ZN(new_n6406_));
  AOI21_X1   g06214(.A1(new_n6399_), .A2(new_n6354_), .B(new_n6019_), .ZN(new_n6407_));
  INV_X1     g06215(.I(\a[67] ), .ZN(new_n6408_));
  AOI21_X1   g06216(.A1(\asqrt[33] ), .A2(new_n6360_), .B(new_n6408_), .ZN(new_n6409_));
  NOR3_X1    g06217(.A1(new_n6406_), .A2(new_n6409_), .A3(new_n6407_), .ZN(new_n6410_));
  OAI21_X1   g06218(.A1(new_n6410_), .A2(new_n6402_), .B(\asqrt[35] ), .ZN(new_n6411_));
  NOR2_X1    g06219(.A1(new_n6344_), .A2(\asqrt[63] ), .ZN(new_n6412_));
  INV_X1     g06220(.I(new_n6336_), .ZN(new_n6413_));
  INV_X1     g06221(.I(new_n6340_), .ZN(new_n6414_));
  NAND2_X1   g06222(.A1(new_n6323_), .A2(new_n6414_), .ZN(new_n6415_));
  INV_X1     g06223(.I(new_n6353_), .ZN(new_n6416_));
  OAI21_X1   g06224(.A1(new_n6413_), .A2(new_n6415_), .B(new_n6416_), .ZN(new_n6417_));
  OAI21_X1   g06225(.A1(new_n6412_), .A2(new_n6417_), .B(new_n6018_), .ZN(new_n6418_));
  NOR2_X1    g06226(.A1(new_n6413_), .A2(new_n6415_), .ZN(new_n6419_));
  OAI21_X1   g06227(.A1(new_n6351_), .A2(new_n6016_), .B(new_n6001_), .ZN(new_n6420_));
  NAND2_X1   g06228(.A1(new_n6349_), .A2(new_n6420_), .ZN(new_n6421_));
  NOR3_X1    g06229(.A1(new_n6412_), .A2(new_n6419_), .A3(new_n6421_), .ZN(new_n6422_));
  INV_X1     g06230(.I(new_n6422_), .ZN(new_n6423_));
  AOI21_X1   g06231(.A1(new_n6423_), .A2(new_n6418_), .B(new_n6038_), .ZN(new_n6424_));
  NOR3_X1    g06232(.A1(new_n6422_), .A2(new_n6407_), .A3(\a[68] ), .ZN(new_n6425_));
  AOI21_X1   g06233(.A1(\asqrt[33] ), .A2(\a[66] ), .B(new_n6359_), .ZN(new_n6426_));
  OAI21_X1   g06234(.A1(new_n6426_), .A2(new_n6077_), .B(new_n5708_), .ZN(new_n6427_));
  OAI22_X1   g06235(.A1(new_n6410_), .A2(new_n6427_), .B1(new_n6424_), .B2(new_n6425_), .ZN(new_n6428_));
  AOI21_X1   g06236(.A1(new_n6428_), .A2(new_n6411_), .B(new_n5277_), .ZN(new_n6429_));
  NOR3_X1    g06237(.A1(new_n6121_), .A2(new_n6037_), .A3(new_n6043_), .ZN(new_n6430_));
  NAND3_X1   g06238(.A1(\asqrt[33] ), .A2(new_n6059_), .A3(new_n6106_), .ZN(new_n6431_));
  AOI22_X1   g06239(.A1(new_n6431_), .A2(new_n6121_), .B1(\asqrt[33] ), .B2(new_n6430_), .ZN(new_n6432_));
  AOI21_X1   g06240(.A1(new_n6399_), .A2(new_n6354_), .B(\a[66] ), .ZN(new_n6433_));
  OAI21_X1   g06241(.A1(new_n6408_), .A2(new_n6433_), .B(new_n6418_), .ZN(new_n6434_));
  OAI21_X1   g06242(.A1(new_n6434_), .A2(new_n6406_), .B(new_n6401_), .ZN(new_n6435_));
  AOI21_X1   g06243(.A1(new_n6435_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n6436_));
  AOI21_X1   g06244(.A1(new_n6436_), .A2(new_n6428_), .B(new_n6432_), .ZN(new_n6437_));
  OAI21_X1   g06245(.A1(new_n6437_), .A2(new_n6429_), .B(\asqrt[37] ), .ZN(new_n6438_));
  INV_X1     g06246(.I(new_n6438_), .ZN(new_n6439_));
  NOR2_X1    g06247(.A1(new_n6058_), .A2(new_n6054_), .ZN(new_n6440_));
  INV_X1     g06248(.I(new_n6440_), .ZN(new_n6441_));
  NOR2_X1    g06249(.A1(new_n6047_), .A2(new_n6060_), .ZN(new_n6442_));
  NOR3_X1    g06250(.A1(new_n6110_), .A2(new_n6441_), .A3(new_n6442_), .ZN(new_n6443_));
  NOR3_X1    g06251(.A1(new_n6356_), .A2(new_n6110_), .A3(new_n6442_), .ZN(new_n6444_));
  INV_X1     g06252(.I(new_n6444_), .ZN(new_n6445_));
  AOI22_X1   g06253(.A1(new_n6445_), .A2(new_n6441_), .B1(\asqrt[33] ), .B2(new_n6443_), .ZN(new_n6446_));
  NOR3_X1    g06254(.A1(new_n6437_), .A2(new_n6429_), .A3(\asqrt[37] ), .ZN(new_n6447_));
  NOR2_X1    g06255(.A1(new_n6447_), .A2(new_n6446_), .ZN(new_n6448_));
  OAI21_X1   g06256(.A1(new_n6448_), .A2(new_n6439_), .B(\asqrt[38] ), .ZN(new_n6449_));
  NOR2_X1    g06257(.A1(new_n6123_), .A2(new_n6115_), .ZN(new_n6450_));
  NOR3_X1    g06258(.A1(new_n6356_), .A2(new_n6062_), .A3(new_n6450_), .ZN(new_n6451_));
  INV_X1     g06259(.I(new_n6451_), .ZN(new_n6452_));
  NOR3_X1    g06260(.A1(new_n6450_), .A2(new_n6062_), .A3(new_n6120_), .ZN(new_n6453_));
  AOI22_X1   g06261(.A1(new_n6452_), .A2(new_n6120_), .B1(\asqrt[33] ), .B2(new_n6453_), .ZN(new_n6454_));
  INV_X1     g06262(.I(new_n6454_), .ZN(new_n6455_));
  NAND2_X1   g06263(.A1(new_n6438_), .A2(new_n4696_), .ZN(new_n6456_));
  OAI21_X1   g06264(.A1(new_n6448_), .A2(new_n6456_), .B(new_n6455_), .ZN(new_n6457_));
  AOI21_X1   g06265(.A1(new_n6457_), .A2(new_n6449_), .B(new_n4298_), .ZN(new_n6458_));
  NOR3_X1    g06266(.A1(new_n6072_), .A2(new_n6081_), .A3(new_n6079_), .ZN(new_n6459_));
  NOR3_X1    g06267(.A1(new_n6356_), .A2(new_n6072_), .A3(new_n6081_), .ZN(new_n6460_));
  INV_X1     g06268(.I(new_n6460_), .ZN(new_n6461_));
  AOI22_X1   g06269(.A1(new_n6461_), .A2(new_n6079_), .B1(\asqrt[33] ), .B2(new_n6459_), .ZN(new_n6462_));
  OAI21_X1   g06270(.A1(new_n6446_), .A2(new_n6447_), .B(new_n6438_), .ZN(new_n6463_));
  AOI21_X1   g06271(.A1(new_n6463_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n6464_));
  AOI21_X1   g06272(.A1(new_n6464_), .A2(new_n6457_), .B(new_n6462_), .ZN(new_n6465_));
  OAI21_X1   g06273(.A1(new_n6465_), .A2(new_n6458_), .B(\asqrt[40] ), .ZN(new_n6466_));
  INV_X1     g06274(.I(new_n6466_), .ZN(new_n6467_));
  NOR2_X1    g06275(.A1(new_n6082_), .A2(new_n6090_), .ZN(new_n6468_));
  NOR3_X1    g06276(.A1(new_n6356_), .A2(new_n6119_), .A3(new_n6468_), .ZN(new_n6469_));
  INV_X1     g06277(.I(new_n6469_), .ZN(new_n6470_));
  NOR3_X1    g06278(.A1(new_n6468_), .A2(new_n6119_), .A3(new_n6089_), .ZN(new_n6471_));
  AOI22_X1   g06279(.A1(new_n6470_), .A2(new_n6089_), .B1(\asqrt[33] ), .B2(new_n6471_), .ZN(new_n6472_));
  NOR3_X1    g06280(.A1(new_n6465_), .A2(new_n6458_), .A3(\asqrt[40] ), .ZN(new_n6473_));
  NOR2_X1    g06281(.A1(new_n6473_), .A2(new_n6472_), .ZN(new_n6474_));
  OAI21_X1   g06282(.A1(new_n6474_), .A2(new_n6467_), .B(\asqrt[41] ), .ZN(new_n6475_));
  INV_X1     g06283(.I(new_n6096_), .ZN(new_n6476_));
  NOR3_X1    g06284(.A1(new_n6092_), .A2(new_n6137_), .A3(new_n6476_), .ZN(new_n6477_));
  NOR3_X1    g06285(.A1(new_n6356_), .A2(new_n6092_), .A3(new_n6137_), .ZN(new_n6478_));
  INV_X1     g06286(.I(new_n6478_), .ZN(new_n6479_));
  AOI22_X1   g06287(.A1(new_n6479_), .A2(new_n6476_), .B1(\asqrt[33] ), .B2(new_n6477_), .ZN(new_n6480_));
  INV_X1     g06288(.I(new_n6480_), .ZN(new_n6481_));
  NAND2_X1   g06289(.A1(new_n6466_), .A2(new_n3782_), .ZN(new_n6482_));
  OAI21_X1   g06290(.A1(new_n6474_), .A2(new_n6482_), .B(new_n6481_), .ZN(new_n6483_));
  AOI21_X1   g06291(.A1(new_n6483_), .A2(new_n6475_), .B(new_n3419_), .ZN(new_n6484_));
  NOR3_X1    g06292(.A1(new_n6356_), .A2(new_n6368_), .A3(new_n6164_), .ZN(new_n6485_));
  INV_X1     g06293(.I(new_n6485_), .ZN(new_n6486_));
  NOR3_X1    g06294(.A1(new_n6368_), .A2(new_n6105_), .A3(new_n6164_), .ZN(new_n6487_));
  AOI22_X1   g06295(.A1(new_n6486_), .A2(new_n6105_), .B1(\asqrt[33] ), .B2(new_n6487_), .ZN(new_n6488_));
  OAI21_X1   g06296(.A1(new_n6472_), .A2(new_n6473_), .B(new_n6466_), .ZN(new_n6489_));
  AOI21_X1   g06297(.A1(new_n6489_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n6490_));
  AOI21_X1   g06298(.A1(new_n6490_), .A2(new_n6483_), .B(new_n6488_), .ZN(new_n6491_));
  OAI21_X1   g06299(.A1(new_n6491_), .A2(new_n6484_), .B(\asqrt[43] ), .ZN(new_n6492_));
  INV_X1     g06300(.I(new_n6492_), .ZN(new_n6493_));
  INV_X1     g06301(.I(new_n6167_), .ZN(new_n6494_));
  NOR3_X1    g06302(.A1(new_n6494_), .A2(new_n6131_), .A3(new_n6166_), .ZN(new_n6495_));
  NOR3_X1    g06303(.A1(new_n6356_), .A2(new_n6131_), .A3(new_n6494_), .ZN(new_n6496_));
  INV_X1     g06304(.I(new_n6496_), .ZN(new_n6497_));
  AOI22_X1   g06305(.A1(new_n6497_), .A2(new_n6166_), .B1(\asqrt[33] ), .B2(new_n6495_), .ZN(new_n6498_));
  NOR3_X1    g06306(.A1(new_n6491_), .A2(new_n6484_), .A3(\asqrt[43] ), .ZN(new_n6499_));
  NOR2_X1    g06307(.A1(new_n6499_), .A2(new_n6498_), .ZN(new_n6500_));
  OAI21_X1   g06308(.A1(new_n6500_), .A2(new_n6493_), .B(\asqrt[44] ), .ZN(new_n6501_));
  NOR3_X1    g06309(.A1(new_n6356_), .A2(new_n6142_), .A3(new_n6147_), .ZN(new_n6502_));
  INV_X1     g06310(.I(new_n6502_), .ZN(new_n6503_));
  NOR3_X1    g06311(.A1(new_n6142_), .A2(new_n6147_), .A3(new_n6367_), .ZN(new_n6504_));
  AOI22_X1   g06312(.A1(new_n6503_), .A2(new_n6367_), .B1(\asqrt[33] ), .B2(new_n6504_), .ZN(new_n6505_));
  INV_X1     g06313(.I(new_n6505_), .ZN(new_n6506_));
  NAND2_X1   g06314(.A1(new_n6492_), .A2(new_n2954_), .ZN(new_n6507_));
  OAI21_X1   g06315(.A1(new_n6500_), .A2(new_n6507_), .B(new_n6506_), .ZN(new_n6508_));
  AOI21_X1   g06316(.A1(new_n6508_), .A2(new_n6501_), .B(new_n2641_), .ZN(new_n6509_));
  INV_X1     g06317(.I(new_n6149_), .ZN(new_n6510_));
  NOR2_X1    g06318(.A1(new_n6148_), .A2(new_n6156_), .ZN(new_n6511_));
  NOR3_X1    g06319(.A1(new_n6510_), .A2(new_n6155_), .A3(new_n6511_), .ZN(new_n6512_));
  NOR3_X1    g06320(.A1(new_n6356_), .A2(new_n6510_), .A3(new_n6511_), .ZN(new_n6513_));
  INV_X1     g06321(.I(new_n6513_), .ZN(new_n6514_));
  AOI22_X1   g06322(.A1(new_n6514_), .A2(new_n6155_), .B1(\asqrt[33] ), .B2(new_n6512_), .ZN(new_n6515_));
  OAI21_X1   g06323(.A1(new_n6498_), .A2(new_n6499_), .B(new_n6492_), .ZN(new_n6516_));
  AOI21_X1   g06324(.A1(new_n6516_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n6517_));
  AOI21_X1   g06325(.A1(new_n6517_), .A2(new_n6508_), .B(new_n6515_), .ZN(new_n6518_));
  OAI21_X1   g06326(.A1(new_n6518_), .A2(new_n6509_), .B(\asqrt[46] ), .ZN(new_n6519_));
  INV_X1     g06327(.I(new_n6519_), .ZN(new_n6520_));
  INV_X1     g06328(.I(new_n6163_), .ZN(new_n6521_));
  INV_X1     g06329(.I(new_n6157_), .ZN(new_n6522_));
  INV_X1     g06330(.I(new_n6170_), .ZN(new_n6523_));
  NOR2_X1    g06331(.A1(new_n6523_), .A2(new_n6522_), .ZN(new_n6524_));
  NOR3_X1    g06332(.A1(new_n6356_), .A2(new_n6158_), .A3(new_n6524_), .ZN(new_n6525_));
  INV_X1     g06333(.I(new_n6525_), .ZN(new_n6526_));
  NOR3_X1    g06334(.A1(new_n6524_), .A2(new_n6158_), .A3(new_n6521_), .ZN(new_n6527_));
  AOI22_X1   g06335(.A1(new_n6526_), .A2(new_n6521_), .B1(\asqrt[33] ), .B2(new_n6527_), .ZN(new_n6528_));
  NOR3_X1    g06336(.A1(new_n6518_), .A2(new_n6509_), .A3(\asqrt[46] ), .ZN(new_n6529_));
  NOR2_X1    g06337(.A1(new_n6529_), .A2(new_n6528_), .ZN(new_n6530_));
  OAI21_X1   g06338(.A1(new_n6530_), .A2(new_n6520_), .B(\asqrt[47] ), .ZN(new_n6531_));
  NOR3_X1    g06339(.A1(new_n6173_), .A2(new_n6366_), .A3(new_n6178_), .ZN(new_n6532_));
  NOR3_X1    g06340(.A1(new_n6356_), .A2(new_n6173_), .A3(new_n6178_), .ZN(new_n6533_));
  INV_X1     g06341(.I(new_n6533_), .ZN(new_n6534_));
  AOI22_X1   g06342(.A1(new_n6534_), .A2(new_n6366_), .B1(\asqrt[33] ), .B2(new_n6532_), .ZN(new_n6535_));
  INV_X1     g06343(.I(new_n6535_), .ZN(new_n6536_));
  NAND2_X1   g06344(.A1(new_n6519_), .A2(new_n2229_), .ZN(new_n6537_));
  OAI21_X1   g06345(.A1(new_n6530_), .A2(new_n6537_), .B(new_n6536_), .ZN(new_n6538_));
  AOI21_X1   g06346(.A1(new_n6538_), .A2(new_n6531_), .B(new_n1956_), .ZN(new_n6539_));
  INV_X1     g06347(.I(new_n6180_), .ZN(new_n6540_));
  NOR2_X1    g06348(.A1(new_n6179_), .A2(new_n6187_), .ZN(new_n6541_));
  NOR3_X1    g06349(.A1(new_n6356_), .A2(new_n6540_), .A3(new_n6541_), .ZN(new_n6542_));
  INV_X1     g06350(.I(new_n6542_), .ZN(new_n6543_));
  NOR3_X1    g06351(.A1(new_n6540_), .A2(new_n6186_), .A3(new_n6541_), .ZN(new_n6544_));
  AOI22_X1   g06352(.A1(new_n6543_), .A2(new_n6186_), .B1(\asqrt[33] ), .B2(new_n6544_), .ZN(new_n6545_));
  OAI21_X1   g06353(.A1(new_n6528_), .A2(new_n6529_), .B(new_n6519_), .ZN(new_n6546_));
  AOI21_X1   g06354(.A1(new_n6546_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n6547_));
  AOI21_X1   g06355(.A1(new_n6547_), .A2(new_n6538_), .B(new_n6545_), .ZN(new_n6548_));
  OAI21_X1   g06356(.A1(new_n6548_), .A2(new_n6539_), .B(\asqrt[49] ), .ZN(new_n6549_));
  INV_X1     g06357(.I(new_n6549_), .ZN(new_n6550_));
  INV_X1     g06358(.I(new_n6194_), .ZN(new_n6551_));
  INV_X1     g06359(.I(new_n6188_), .ZN(new_n6552_));
  INV_X1     g06360(.I(new_n6196_), .ZN(new_n6553_));
  NOR2_X1    g06361(.A1(new_n6553_), .A2(new_n6552_), .ZN(new_n6554_));
  NOR3_X1    g06362(.A1(new_n6554_), .A2(new_n6189_), .A3(new_n6551_), .ZN(new_n6555_));
  NOR3_X1    g06363(.A1(new_n6356_), .A2(new_n6189_), .A3(new_n6554_), .ZN(new_n6556_));
  INV_X1     g06364(.I(new_n6556_), .ZN(new_n6557_));
  AOI22_X1   g06365(.A1(new_n6557_), .A2(new_n6551_), .B1(\asqrt[33] ), .B2(new_n6555_), .ZN(new_n6558_));
  NOR3_X1    g06366(.A1(new_n6548_), .A2(new_n6539_), .A3(\asqrt[49] ), .ZN(new_n6559_));
  NOR2_X1    g06367(.A1(new_n6559_), .A2(new_n6558_), .ZN(new_n6560_));
  OAI21_X1   g06368(.A1(new_n6560_), .A2(new_n6550_), .B(\asqrt[50] ), .ZN(new_n6561_));
  NOR3_X1    g06369(.A1(new_n6356_), .A2(new_n6199_), .A3(new_n6204_), .ZN(new_n6562_));
  INV_X1     g06370(.I(new_n6562_), .ZN(new_n6563_));
  NOR3_X1    g06371(.A1(new_n6199_), .A2(new_n6365_), .A3(new_n6204_), .ZN(new_n6564_));
  AOI22_X1   g06372(.A1(new_n6563_), .A2(new_n6365_), .B1(\asqrt[33] ), .B2(new_n6564_), .ZN(new_n6565_));
  INV_X1     g06373(.I(new_n6565_), .ZN(new_n6566_));
  NAND2_X1   g06374(.A1(new_n6549_), .A2(new_n1612_), .ZN(new_n6567_));
  OAI21_X1   g06375(.A1(new_n6560_), .A2(new_n6567_), .B(new_n6566_), .ZN(new_n6568_));
  AOI21_X1   g06376(.A1(new_n6568_), .A2(new_n6561_), .B(new_n1376_), .ZN(new_n6569_));
  INV_X1     g06377(.I(new_n6206_), .ZN(new_n6570_));
  NOR2_X1    g06378(.A1(new_n6205_), .A2(new_n6213_), .ZN(new_n6571_));
  NOR3_X1    g06379(.A1(new_n6570_), .A2(new_n6212_), .A3(new_n6571_), .ZN(new_n6572_));
  NOR3_X1    g06380(.A1(new_n6356_), .A2(new_n6570_), .A3(new_n6571_), .ZN(new_n6573_));
  INV_X1     g06381(.I(new_n6573_), .ZN(new_n6574_));
  AOI22_X1   g06382(.A1(new_n6574_), .A2(new_n6212_), .B1(\asqrt[33] ), .B2(new_n6572_), .ZN(new_n6575_));
  OAI21_X1   g06383(.A1(new_n6558_), .A2(new_n6559_), .B(new_n6549_), .ZN(new_n6576_));
  AOI21_X1   g06384(.A1(new_n6576_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n6577_));
  AOI21_X1   g06385(.A1(new_n6577_), .A2(new_n6568_), .B(new_n6575_), .ZN(new_n6578_));
  OAI21_X1   g06386(.A1(new_n6578_), .A2(new_n6569_), .B(\asqrt[52] ), .ZN(new_n6579_));
  INV_X1     g06387(.I(new_n6220_), .ZN(new_n6580_));
  INV_X1     g06388(.I(new_n6214_), .ZN(new_n6581_));
  INV_X1     g06389(.I(new_n6222_), .ZN(new_n6582_));
  NOR2_X1    g06390(.A1(new_n6582_), .A2(new_n6581_), .ZN(new_n6583_));
  NOR3_X1    g06391(.A1(new_n6356_), .A2(new_n6215_), .A3(new_n6583_), .ZN(new_n6584_));
  INV_X1     g06392(.I(new_n6584_), .ZN(new_n6585_));
  NOR3_X1    g06393(.A1(new_n6583_), .A2(new_n6215_), .A3(new_n6580_), .ZN(new_n6586_));
  AOI22_X1   g06394(.A1(new_n6585_), .A2(new_n6580_), .B1(\asqrt[33] ), .B2(new_n6586_), .ZN(new_n6587_));
  INV_X1     g06395(.I(new_n6587_), .ZN(new_n6588_));
  INV_X1     g06396(.I(new_n6558_), .ZN(new_n6589_));
  INV_X1     g06397(.I(new_n6539_), .ZN(new_n6590_));
  NAND2_X1   g06398(.A1(new_n6590_), .A2(new_n1806_), .ZN(new_n6591_));
  OAI21_X1   g06399(.A1(new_n6591_), .A2(new_n6548_), .B(new_n6589_), .ZN(new_n6592_));
  AOI21_X1   g06400(.A1(new_n6592_), .A2(new_n6549_), .B(new_n1612_), .ZN(new_n6593_));
  INV_X1     g06401(.I(new_n6567_), .ZN(new_n6594_));
  AOI21_X1   g06402(.A1(new_n6594_), .A2(new_n6592_), .B(new_n6565_), .ZN(new_n6595_));
  OAI21_X1   g06403(.A1(new_n6595_), .A2(new_n6593_), .B(\asqrt[51] ), .ZN(new_n6596_));
  NAND2_X1   g06404(.A1(new_n6596_), .A2(new_n1256_), .ZN(new_n6597_));
  OAI21_X1   g06405(.A1(new_n6597_), .A2(new_n6578_), .B(new_n6588_), .ZN(new_n6598_));
  AOI21_X1   g06406(.A1(new_n6598_), .A2(new_n6579_), .B(new_n1103_), .ZN(new_n6599_));
  NOR3_X1    g06407(.A1(new_n6225_), .A2(new_n6364_), .A3(new_n6267_), .ZN(new_n6600_));
  NOR3_X1    g06408(.A1(new_n6356_), .A2(new_n6225_), .A3(new_n6267_), .ZN(new_n6601_));
  INV_X1     g06409(.I(new_n6601_), .ZN(new_n6602_));
  AOI22_X1   g06410(.A1(new_n6602_), .A2(new_n6364_), .B1(\asqrt[33] ), .B2(new_n6600_), .ZN(new_n6603_));
  INV_X1     g06411(.I(new_n6575_), .ZN(new_n6604_));
  NAND2_X1   g06412(.A1(new_n6561_), .A2(new_n1376_), .ZN(new_n6605_));
  OAI21_X1   g06413(.A1(new_n6605_), .A2(new_n6595_), .B(new_n6604_), .ZN(new_n6606_));
  AOI21_X1   g06414(.A1(new_n6606_), .A2(new_n6596_), .B(new_n1256_), .ZN(new_n6607_));
  NOR2_X1    g06415(.A1(new_n6607_), .A2(\asqrt[53] ), .ZN(new_n6608_));
  AOI21_X1   g06416(.A1(new_n6608_), .A2(new_n6598_), .B(new_n6603_), .ZN(new_n6609_));
  OAI21_X1   g06417(.A1(new_n6609_), .A2(new_n6599_), .B(\asqrt[54] ), .ZN(new_n6610_));
  INV_X1     g06418(.I(new_n6233_), .ZN(new_n6611_));
  NOR2_X1    g06419(.A1(new_n6240_), .A2(new_n6232_), .ZN(new_n6612_));
  NOR3_X1    g06420(.A1(new_n6356_), .A2(new_n6611_), .A3(new_n6612_), .ZN(new_n6613_));
  INV_X1     g06421(.I(new_n6613_), .ZN(new_n6614_));
  NOR3_X1    g06422(.A1(new_n6611_), .A2(new_n6239_), .A3(new_n6612_), .ZN(new_n6615_));
  AOI22_X1   g06423(.A1(new_n6614_), .A2(new_n6239_), .B1(\asqrt[33] ), .B2(new_n6615_), .ZN(new_n6616_));
  INV_X1     g06424(.I(new_n6616_), .ZN(new_n6617_));
  NOR2_X1    g06425(.A1(new_n6569_), .A2(\asqrt[52] ), .ZN(new_n6618_));
  AOI21_X1   g06426(.A1(new_n6618_), .A2(new_n6606_), .B(new_n6587_), .ZN(new_n6619_));
  OAI21_X1   g06427(.A1(new_n6619_), .A2(new_n6607_), .B(\asqrt[53] ), .ZN(new_n6620_));
  NAND2_X1   g06428(.A1(new_n6620_), .A2(new_n904_), .ZN(new_n6621_));
  OAI21_X1   g06429(.A1(new_n6621_), .A2(new_n6609_), .B(new_n6617_), .ZN(new_n6622_));
  AOI21_X1   g06430(.A1(new_n6622_), .A2(new_n6610_), .B(new_n823_), .ZN(new_n6623_));
  NOR2_X1    g06431(.A1(new_n6251_), .A2(new_n6244_), .ZN(new_n6624_));
  NOR3_X1    g06432(.A1(new_n6624_), .A2(new_n6242_), .A3(new_n6250_), .ZN(new_n6625_));
  NOR3_X1    g06433(.A1(new_n6356_), .A2(new_n6242_), .A3(new_n6624_), .ZN(new_n6626_));
  INV_X1     g06434(.I(new_n6626_), .ZN(new_n6627_));
  AOI22_X1   g06435(.A1(new_n6627_), .A2(new_n6250_), .B1(\asqrt[33] ), .B2(new_n6625_), .ZN(new_n6628_));
  INV_X1     g06436(.I(new_n6603_), .ZN(new_n6629_));
  NAND2_X1   g06437(.A1(new_n6579_), .A2(new_n1103_), .ZN(new_n6630_));
  OAI21_X1   g06438(.A1(new_n6630_), .A2(new_n6619_), .B(new_n6629_), .ZN(new_n6631_));
  AOI21_X1   g06439(.A1(new_n6631_), .A2(new_n6620_), .B(new_n904_), .ZN(new_n6632_));
  NOR2_X1    g06440(.A1(new_n6632_), .A2(\asqrt[55] ), .ZN(new_n6633_));
  AOI21_X1   g06441(.A1(new_n6633_), .A2(new_n6622_), .B(new_n6628_), .ZN(new_n6634_));
  OAI21_X1   g06442(.A1(new_n6634_), .A2(new_n6623_), .B(\asqrt[56] ), .ZN(new_n6635_));
  NOR3_X1    g06443(.A1(new_n6356_), .A2(new_n6253_), .A3(new_n6299_), .ZN(new_n6636_));
  INV_X1     g06444(.I(new_n6636_), .ZN(new_n6637_));
  NOR3_X1    g06445(.A1(new_n6253_), .A2(new_n6363_), .A3(new_n6299_), .ZN(new_n6638_));
  AOI22_X1   g06446(.A1(new_n6637_), .A2(new_n6363_), .B1(\asqrt[33] ), .B2(new_n6638_), .ZN(new_n6639_));
  INV_X1     g06447(.I(new_n6639_), .ZN(new_n6640_));
  NOR3_X1    g06448(.A1(new_n6578_), .A2(new_n6569_), .A3(\asqrt[52] ), .ZN(new_n6641_));
  OAI21_X1   g06449(.A1(new_n6587_), .A2(new_n6641_), .B(new_n6579_), .ZN(new_n6642_));
  AOI21_X1   g06450(.A1(new_n6642_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n6643_));
  AOI21_X1   g06451(.A1(new_n6643_), .A2(new_n6631_), .B(new_n6616_), .ZN(new_n6644_));
  OAI21_X1   g06452(.A1(new_n6644_), .A2(new_n6632_), .B(\asqrt[55] ), .ZN(new_n6645_));
  NAND2_X1   g06453(.A1(new_n6645_), .A2(new_n703_), .ZN(new_n6646_));
  OAI21_X1   g06454(.A1(new_n6646_), .A2(new_n6634_), .B(new_n6640_), .ZN(new_n6647_));
  AOI21_X1   g06455(.A1(new_n6647_), .A2(new_n6635_), .B(new_n531_), .ZN(new_n6648_));
  INV_X1     g06456(.I(new_n6260_), .ZN(new_n6649_));
  NOR2_X1    g06457(.A1(new_n6272_), .A2(new_n6259_), .ZN(new_n6650_));
  NOR3_X1    g06458(.A1(new_n6649_), .A2(new_n6266_), .A3(new_n6650_), .ZN(new_n6651_));
  NOR3_X1    g06459(.A1(new_n6356_), .A2(new_n6649_), .A3(new_n6650_), .ZN(new_n6652_));
  INV_X1     g06460(.I(new_n6652_), .ZN(new_n6653_));
  AOI22_X1   g06461(.A1(new_n6653_), .A2(new_n6266_), .B1(\asqrt[33] ), .B2(new_n6651_), .ZN(new_n6654_));
  NOR3_X1    g06462(.A1(new_n6644_), .A2(\asqrt[55] ), .A3(new_n6632_), .ZN(new_n6655_));
  OAI21_X1   g06463(.A1(new_n6628_), .A2(new_n6655_), .B(new_n6645_), .ZN(new_n6656_));
  AOI21_X1   g06464(.A1(new_n6656_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n6657_));
  AOI21_X1   g06465(.A1(new_n6657_), .A2(new_n6647_), .B(new_n6654_), .ZN(new_n6658_));
  OAI21_X1   g06466(.A1(new_n6658_), .A2(new_n6648_), .B(\asqrt[58] ), .ZN(new_n6659_));
  NOR2_X1    g06467(.A1(new_n6283_), .A2(new_n6276_), .ZN(new_n6660_));
  NOR3_X1    g06468(.A1(new_n6356_), .A2(new_n6274_), .A3(new_n6660_), .ZN(new_n6661_));
  INV_X1     g06469(.I(new_n6661_), .ZN(new_n6662_));
  NOR3_X1    g06470(.A1(new_n6660_), .A2(new_n6274_), .A3(new_n6282_), .ZN(new_n6663_));
  AOI22_X1   g06471(.A1(new_n6662_), .A2(new_n6282_), .B1(\asqrt[33] ), .B2(new_n6663_), .ZN(new_n6664_));
  INV_X1     g06472(.I(new_n6664_), .ZN(new_n6665_));
  INV_X1     g06473(.I(new_n6628_), .ZN(new_n6666_));
  NAND2_X1   g06474(.A1(new_n6610_), .A2(new_n823_), .ZN(new_n6667_));
  OAI21_X1   g06475(.A1(new_n6667_), .A2(new_n6644_), .B(new_n6666_), .ZN(new_n6668_));
  AOI21_X1   g06476(.A1(new_n6668_), .A2(new_n6645_), .B(new_n703_), .ZN(new_n6669_));
  NOR2_X1    g06477(.A1(new_n6623_), .A2(\asqrt[56] ), .ZN(new_n6670_));
  AOI21_X1   g06478(.A1(new_n6670_), .A2(new_n6668_), .B(new_n6639_), .ZN(new_n6671_));
  OAI21_X1   g06479(.A1(new_n6671_), .A2(new_n6669_), .B(\asqrt[57] ), .ZN(new_n6672_));
  NAND2_X1   g06480(.A1(new_n6672_), .A2(new_n436_), .ZN(new_n6673_));
  OAI21_X1   g06481(.A1(new_n6673_), .A2(new_n6658_), .B(new_n6665_), .ZN(new_n6674_));
  AOI21_X1   g06482(.A1(new_n6674_), .A2(new_n6659_), .B(new_n327_), .ZN(new_n6675_));
  NOR3_X1    g06483(.A1(new_n6285_), .A2(new_n6362_), .A3(new_n6330_), .ZN(new_n6676_));
  NOR3_X1    g06484(.A1(new_n6356_), .A2(new_n6285_), .A3(new_n6330_), .ZN(new_n6677_));
  INV_X1     g06485(.I(new_n6677_), .ZN(new_n6678_));
  AOI22_X1   g06486(.A1(new_n6678_), .A2(new_n6362_), .B1(\asqrt[33] ), .B2(new_n6676_), .ZN(new_n6679_));
  INV_X1     g06487(.I(new_n6654_), .ZN(new_n6680_));
  NAND2_X1   g06488(.A1(new_n6635_), .A2(new_n531_), .ZN(new_n6681_));
  OAI21_X1   g06489(.A1(new_n6681_), .A2(new_n6671_), .B(new_n6680_), .ZN(new_n6682_));
  AOI21_X1   g06490(.A1(new_n6682_), .A2(new_n6672_), .B(new_n436_), .ZN(new_n6683_));
  NOR2_X1    g06491(.A1(new_n6683_), .A2(\asqrt[59] ), .ZN(new_n6684_));
  AOI21_X1   g06492(.A1(new_n6684_), .A2(new_n6674_), .B(new_n6679_), .ZN(new_n6685_));
  OAI21_X1   g06493(.A1(new_n6685_), .A2(new_n6675_), .B(\asqrt[60] ), .ZN(new_n6686_));
  INV_X1     g06494(.I(new_n6292_), .ZN(new_n6687_));
  NOR2_X1    g06495(.A1(new_n6304_), .A2(new_n6291_), .ZN(new_n6688_));
  NOR3_X1    g06496(.A1(new_n6356_), .A2(new_n6687_), .A3(new_n6688_), .ZN(new_n6689_));
  INV_X1     g06497(.I(new_n6689_), .ZN(new_n6690_));
  NOR3_X1    g06498(.A1(new_n6687_), .A2(new_n6298_), .A3(new_n6688_), .ZN(new_n6691_));
  AOI22_X1   g06499(.A1(new_n6690_), .A2(new_n6298_), .B1(\asqrt[33] ), .B2(new_n6691_), .ZN(new_n6692_));
  INV_X1     g06500(.I(new_n6692_), .ZN(new_n6693_));
  NOR2_X1    g06501(.A1(new_n6648_), .A2(\asqrt[58] ), .ZN(new_n6694_));
  AOI21_X1   g06502(.A1(new_n6694_), .A2(new_n6682_), .B(new_n6664_), .ZN(new_n6695_));
  OAI21_X1   g06503(.A1(new_n6695_), .A2(new_n6683_), .B(\asqrt[59] ), .ZN(new_n6696_));
  NAND2_X1   g06504(.A1(new_n6696_), .A2(new_n306_), .ZN(new_n6697_));
  OAI21_X1   g06505(.A1(new_n6697_), .A2(new_n6685_), .B(new_n6693_), .ZN(new_n6698_));
  AOI21_X1   g06506(.A1(new_n6698_), .A2(new_n6686_), .B(new_n218_), .ZN(new_n6699_));
  NOR2_X1    g06507(.A1(new_n6308_), .A2(new_n6314_), .ZN(new_n6700_));
  NOR3_X1    g06508(.A1(new_n6700_), .A2(new_n6306_), .A3(new_n6313_), .ZN(new_n6701_));
  NOR3_X1    g06509(.A1(new_n6356_), .A2(new_n6306_), .A3(new_n6700_), .ZN(new_n6702_));
  INV_X1     g06510(.I(new_n6702_), .ZN(new_n6703_));
  AOI22_X1   g06511(.A1(new_n6703_), .A2(new_n6313_), .B1(\asqrt[33] ), .B2(new_n6701_), .ZN(new_n6704_));
  INV_X1     g06512(.I(new_n6679_), .ZN(new_n6705_));
  NAND2_X1   g06513(.A1(new_n6659_), .A2(new_n327_), .ZN(new_n6706_));
  OAI21_X1   g06514(.A1(new_n6706_), .A2(new_n6695_), .B(new_n6705_), .ZN(new_n6707_));
  AOI21_X1   g06515(.A1(new_n6707_), .A2(new_n6696_), .B(new_n306_), .ZN(new_n6708_));
  NOR2_X1    g06516(.A1(new_n6708_), .A2(\asqrt[61] ), .ZN(new_n6709_));
  AOI21_X1   g06517(.A1(new_n6709_), .A2(new_n6698_), .B(new_n6704_), .ZN(new_n6710_));
  OAI21_X1   g06518(.A1(new_n6710_), .A2(new_n6699_), .B(\asqrt[62] ), .ZN(new_n6711_));
  NOR3_X1    g06519(.A1(new_n6356_), .A2(new_n6316_), .A3(new_n6345_), .ZN(new_n6712_));
  INV_X1     g06520(.I(new_n6712_), .ZN(new_n6713_));
  NOR3_X1    g06521(.A1(new_n6316_), .A2(new_n6361_), .A3(new_n6345_), .ZN(new_n6714_));
  AOI22_X1   g06522(.A1(new_n6713_), .A2(new_n6361_), .B1(\asqrt[33] ), .B2(new_n6714_), .ZN(new_n6715_));
  INV_X1     g06523(.I(new_n6715_), .ZN(new_n6716_));
  NOR3_X1    g06524(.A1(new_n6658_), .A2(\asqrt[58] ), .A3(new_n6648_), .ZN(new_n6717_));
  OAI21_X1   g06525(.A1(new_n6664_), .A2(new_n6717_), .B(new_n6659_), .ZN(new_n6718_));
  AOI21_X1   g06526(.A1(new_n6718_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n6719_));
  AOI21_X1   g06527(.A1(new_n6719_), .A2(new_n6707_), .B(new_n6692_), .ZN(new_n6720_));
  OAI21_X1   g06528(.A1(new_n6720_), .A2(new_n6708_), .B(\asqrt[61] ), .ZN(new_n6721_));
  NAND2_X1   g06529(.A1(new_n6721_), .A2(new_n207_), .ZN(new_n6722_));
  OAI21_X1   g06530(.A1(new_n6722_), .A2(new_n6710_), .B(new_n6716_), .ZN(new_n6723_));
  INV_X1     g06531(.I(new_n6419_), .ZN(new_n6724_));
  NAND4_X1   g06532(.A1(\asqrt[33] ), .A2(new_n6323_), .A3(new_n6328_), .A4(new_n6397_), .ZN(new_n6725_));
  NAND2_X1   g06533(.A1(new_n6323_), .A2(new_n6397_), .ZN(new_n6726_));
  OAI21_X1   g06534(.A1(new_n6356_), .A2(new_n6726_), .B(new_n6329_), .ZN(new_n6727_));
  NAND2_X1   g06535(.A1(new_n6727_), .A2(new_n6725_), .ZN(new_n6728_));
  NOR2_X1    g06536(.A1(new_n6398_), .A2(new_n6414_), .ZN(new_n6729_));
  NAND2_X1   g06537(.A1(\asqrt[33] ), .A2(new_n6729_), .ZN(new_n6730_));
  NAND3_X1   g06538(.A1(new_n6728_), .A2(new_n6724_), .A3(new_n6730_), .ZN(new_n6731_));
  AOI21_X1   g06539(.A1(new_n6723_), .A2(new_n6711_), .B(new_n6731_), .ZN(new_n6732_));
  NOR3_X1    g06540(.A1(new_n6720_), .A2(\asqrt[61] ), .A3(new_n6708_), .ZN(new_n6733_));
  OAI21_X1   g06541(.A1(new_n6704_), .A2(new_n6733_), .B(new_n6721_), .ZN(new_n6734_));
  AOI21_X1   g06542(.A1(new_n6734_), .A2(\asqrt[62] ), .B(new_n6728_), .ZN(new_n6735_));
  OAI21_X1   g06543(.A1(new_n6356_), .A2(new_n6414_), .B(new_n6398_), .ZN(new_n6736_));
  NOR2_X1    g06544(.A1(new_n6729_), .A2(new_n193_), .ZN(new_n6737_));
  NAND2_X1   g06545(.A1(new_n6736_), .A2(new_n6737_), .ZN(new_n6738_));
  INV_X1     g06546(.I(new_n6738_), .ZN(new_n6739_));
  AND3_X2    g06547(.A1(new_n6339_), .A2(new_n6337_), .A3(new_n6352_), .Z(new_n6740_));
  NAND4_X1   g06548(.A1(new_n6724_), .A2(new_n6399_), .A3(new_n6349_), .A4(new_n6740_), .ZN(new_n6741_));
  INV_X1     g06549(.I(new_n6741_), .ZN(new_n6742_));
  NOR2_X1    g06550(.A1(new_n6739_), .A2(new_n6742_), .ZN(new_n6743_));
  INV_X1     g06551(.I(new_n6743_), .ZN(new_n6744_));
  AOI21_X1   g06552(.A1(new_n6735_), .A2(new_n6723_), .B(new_n6744_), .ZN(new_n6745_));
  OAI21_X1   g06553(.A1(\asqrt[63] ), .A2(new_n6732_), .B(new_n6745_), .ZN(\asqrt[32] ));
  NOR2_X1    g06554(.A1(\a[62] ), .A2(\a[63] ), .ZN(new_n6747_));
  INV_X1     g06555(.I(new_n6747_), .ZN(new_n6748_));
  NOR2_X1    g06556(.A1(new_n6748_), .A2(\a[64] ), .ZN(new_n6749_));
  INV_X1     g06557(.I(new_n6749_), .ZN(new_n6750_));
  NAND2_X1   g06558(.A1(new_n6723_), .A2(new_n6711_), .ZN(new_n6751_));
  INV_X1     g06559(.I(new_n6731_), .ZN(new_n6752_));
  AOI21_X1   g06560(.A1(new_n6751_), .A2(new_n6752_), .B(\asqrt[63] ), .ZN(new_n6753_));
  INV_X1     g06561(.I(new_n6723_), .ZN(new_n6754_));
  INV_X1     g06562(.I(new_n6728_), .ZN(new_n6755_));
  NAND2_X1   g06563(.A1(new_n6711_), .A2(new_n6755_), .ZN(new_n6756_));
  OAI21_X1   g06564(.A1(new_n6754_), .A2(new_n6756_), .B(new_n6743_), .ZN(new_n6757_));
  OAI21_X1   g06565(.A1(new_n6753_), .A2(new_n6757_), .B(\a[64] ), .ZN(new_n6758_));
  AOI21_X1   g06566(.A1(new_n6758_), .A2(new_n6750_), .B(new_n6356_), .ZN(new_n6759_));
  INV_X1     g06567(.I(\a[64] ), .ZN(new_n6760_));
  INV_X1     g06568(.I(new_n6704_), .ZN(new_n6761_));
  NAND2_X1   g06569(.A1(new_n6686_), .A2(new_n218_), .ZN(new_n6762_));
  OAI21_X1   g06570(.A1(new_n6762_), .A2(new_n6720_), .B(new_n6761_), .ZN(new_n6763_));
  NAND3_X1   g06571(.A1(new_n6763_), .A2(new_n207_), .A3(new_n6721_), .ZN(new_n6764_));
  AOI22_X1   g06572(.A1(new_n6764_), .A2(new_n6716_), .B1(new_n6734_), .B2(\asqrt[62] ), .ZN(new_n6765_));
  OAI21_X1   g06573(.A1(new_n6765_), .A2(new_n6731_), .B(new_n193_), .ZN(new_n6766_));
  AOI21_X1   g06574(.A1(new_n6766_), .A2(new_n6745_), .B(new_n6760_), .ZN(new_n6767_));
  NAND4_X1   g06575(.A1(new_n6724_), .A2(new_n6349_), .A3(new_n6352_), .A4(new_n6750_), .ZN(new_n6768_));
  NOR2_X1    g06576(.A1(new_n6768_), .A2(new_n6412_), .ZN(new_n6769_));
  INV_X1     g06577(.I(new_n6769_), .ZN(new_n6770_));
  NOR2_X1    g06578(.A1(new_n6767_), .A2(new_n6770_), .ZN(new_n6771_));
  AOI21_X1   g06579(.A1(new_n6766_), .A2(new_n6745_), .B(new_n6358_), .ZN(new_n6772_));
  INV_X1     g06580(.I(\a[65] ), .ZN(new_n6773_));
  AOI21_X1   g06581(.A1(\asqrt[32] ), .A2(new_n6760_), .B(new_n6773_), .ZN(new_n6774_));
  NOR3_X1    g06582(.A1(new_n6771_), .A2(new_n6774_), .A3(new_n6772_), .ZN(new_n6775_));
  OAI21_X1   g06583(.A1(new_n6775_), .A2(new_n6759_), .B(\asqrt[34] ), .ZN(new_n6776_));
  OAI21_X1   g06584(.A1(new_n6753_), .A2(new_n6757_), .B(new_n6357_), .ZN(new_n6777_));
  NOR2_X1    g06585(.A1(new_n6754_), .A2(new_n6756_), .ZN(new_n6778_));
  NOR2_X1    g06586(.A1(new_n6742_), .A2(new_n6356_), .ZN(new_n6779_));
  NAND2_X1   g06587(.A1(new_n6738_), .A2(new_n6779_), .ZN(new_n6780_));
  NOR3_X1    g06588(.A1(new_n6753_), .A2(new_n6778_), .A3(new_n6780_), .ZN(new_n6781_));
  INV_X1     g06589(.I(new_n6781_), .ZN(new_n6782_));
  AOI21_X1   g06590(.A1(new_n6782_), .A2(new_n6777_), .B(new_n6360_), .ZN(new_n6783_));
  NOR3_X1    g06591(.A1(new_n6781_), .A2(new_n6772_), .A3(\a[66] ), .ZN(new_n6784_));
  AOI21_X1   g06592(.A1(\asqrt[32] ), .A2(\a[64] ), .B(new_n6749_), .ZN(new_n6785_));
  OAI21_X1   g06593(.A1(new_n6785_), .A2(new_n6356_), .B(new_n6077_), .ZN(new_n6786_));
  OAI22_X1   g06594(.A1(new_n6775_), .A2(new_n6786_), .B1(new_n6783_), .B2(new_n6784_), .ZN(new_n6787_));
  AOI21_X1   g06595(.A1(new_n6787_), .A2(new_n6776_), .B(new_n5708_), .ZN(new_n6788_));
  INV_X1     g06596(.I(new_n6434_), .ZN(new_n6789_));
  NOR3_X1    g06597(.A1(new_n6402_), .A2(new_n6789_), .A3(new_n6406_), .ZN(new_n6790_));
  NOR2_X1    g06598(.A1(new_n6402_), .A2(new_n6406_), .ZN(new_n6791_));
  NAND2_X1   g06599(.A1(\asqrt[32] ), .A2(new_n6791_), .ZN(new_n6792_));
  AOI22_X1   g06600(.A1(new_n6792_), .A2(new_n6789_), .B1(\asqrt[32] ), .B2(new_n6790_), .ZN(new_n6793_));
  OAI21_X1   g06601(.A1(new_n6767_), .A2(new_n6749_), .B(\asqrt[33] ), .ZN(new_n6794_));
  AOI21_X1   g06602(.A1(new_n6766_), .A2(new_n6745_), .B(\a[64] ), .ZN(new_n6795_));
  OAI21_X1   g06603(.A1(new_n6773_), .A2(new_n6795_), .B(new_n6777_), .ZN(new_n6796_));
  OAI21_X1   g06604(.A1(new_n6796_), .A2(new_n6771_), .B(new_n6794_), .ZN(new_n6797_));
  AOI21_X1   g06605(.A1(new_n6797_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n6798_));
  AOI21_X1   g06606(.A1(new_n6798_), .A2(new_n6787_), .B(new_n6793_), .ZN(new_n6799_));
  OAI21_X1   g06607(.A1(new_n6799_), .A2(new_n6788_), .B(\asqrt[36] ), .ZN(new_n6800_));
  INV_X1     g06608(.I(new_n6800_), .ZN(new_n6801_));
  NOR2_X1    g06609(.A1(new_n6424_), .A2(new_n6425_), .ZN(new_n6802_));
  NOR2_X1    g06610(.A1(new_n6410_), .A2(new_n6427_), .ZN(new_n6803_));
  INV_X1     g06611(.I(new_n6803_), .ZN(new_n6804_));
  NAND4_X1   g06612(.A1(\asqrt[32] ), .A2(new_n6411_), .A3(new_n6802_), .A4(new_n6804_), .ZN(new_n6805_));
  AND3_X2    g06613(.A1(\asqrt[32] ), .A2(new_n6411_), .A3(new_n6804_), .Z(new_n6806_));
  OAI21_X1   g06614(.A1(new_n6806_), .A2(new_n6802_), .B(new_n6805_), .ZN(new_n6807_));
  INV_X1     g06615(.I(new_n6807_), .ZN(new_n6808_));
  NOR3_X1    g06616(.A1(new_n6799_), .A2(new_n6788_), .A3(\asqrt[36] ), .ZN(new_n6809_));
  NOR2_X1    g06617(.A1(new_n6809_), .A2(new_n6808_), .ZN(new_n6810_));
  OAI21_X1   g06618(.A1(new_n6810_), .A2(new_n6801_), .B(\asqrt[37] ), .ZN(new_n6811_));
  INV_X1     g06619(.I(new_n6432_), .ZN(new_n6812_));
  INV_X1     g06620(.I(new_n6429_), .ZN(new_n6813_));
  NAND2_X1   g06621(.A1(new_n6436_), .A2(new_n6428_), .ZN(new_n6814_));
  NAND3_X1   g06622(.A1(\asqrt[32] ), .A2(new_n6813_), .A3(new_n6814_), .ZN(new_n6815_));
  AND3_X2    g06623(.A1(new_n6813_), .A2(new_n6432_), .A3(new_n6814_), .Z(new_n6816_));
  AOI22_X1   g06624(.A1(new_n6815_), .A2(new_n6812_), .B1(\asqrt[32] ), .B2(new_n6816_), .ZN(new_n6817_));
  INV_X1     g06625(.I(new_n6817_), .ZN(new_n6818_));
  NAND2_X1   g06626(.A1(new_n6800_), .A2(new_n5024_), .ZN(new_n6819_));
  OAI21_X1   g06627(.A1(new_n6810_), .A2(new_n6819_), .B(new_n6818_), .ZN(new_n6820_));
  AOI21_X1   g06628(.A1(new_n6820_), .A2(new_n6811_), .B(new_n4696_), .ZN(new_n6821_));
  INV_X1     g06629(.I(new_n6446_), .ZN(new_n6822_));
  NOR3_X1    g06630(.A1(new_n6439_), .A2(new_n6822_), .A3(new_n6447_), .ZN(new_n6823_));
  INV_X1     g06631(.I(\asqrt[32] ), .ZN(new_n6824_));
  NOR3_X1    g06632(.A1(new_n6824_), .A2(new_n6439_), .A3(new_n6447_), .ZN(new_n6825_));
  INV_X1     g06633(.I(new_n6825_), .ZN(new_n6826_));
  AOI22_X1   g06634(.A1(new_n6826_), .A2(new_n6822_), .B1(\asqrt[32] ), .B2(new_n6823_), .ZN(new_n6827_));
  OAI21_X1   g06635(.A1(new_n6808_), .A2(new_n6809_), .B(new_n6800_), .ZN(new_n6828_));
  AOI21_X1   g06636(.A1(new_n6828_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n6829_));
  AOI21_X1   g06637(.A1(new_n6829_), .A2(new_n6820_), .B(new_n6827_), .ZN(new_n6830_));
  OAI21_X1   g06638(.A1(new_n6830_), .A2(new_n6821_), .B(\asqrt[39] ), .ZN(new_n6831_));
  INV_X1     g06639(.I(new_n6831_), .ZN(new_n6832_));
  INV_X1     g06640(.I(new_n6448_), .ZN(new_n6833_));
  INV_X1     g06641(.I(new_n6456_), .ZN(new_n6834_));
  NAND2_X1   g06642(.A1(new_n6833_), .A2(new_n6834_), .ZN(new_n6835_));
  NAND3_X1   g06643(.A1(\asqrt[32] ), .A2(new_n6449_), .A3(new_n6835_), .ZN(new_n6836_));
  AND3_X2    g06644(.A1(new_n6835_), .A2(new_n6449_), .A3(new_n6454_), .Z(new_n6837_));
  AOI22_X1   g06645(.A1(new_n6836_), .A2(new_n6455_), .B1(\asqrt[32] ), .B2(new_n6837_), .ZN(new_n6838_));
  NOR3_X1    g06646(.A1(new_n6830_), .A2(new_n6821_), .A3(\asqrt[39] ), .ZN(new_n6839_));
  NOR2_X1    g06647(.A1(new_n6839_), .A2(new_n6838_), .ZN(new_n6840_));
  OAI21_X1   g06648(.A1(new_n6840_), .A2(new_n6832_), .B(\asqrt[40] ), .ZN(new_n6841_));
  INV_X1     g06649(.I(new_n6462_), .ZN(new_n6842_));
  INV_X1     g06650(.I(new_n6457_), .ZN(new_n6843_));
  INV_X1     g06651(.I(new_n6464_), .ZN(new_n6844_));
  NOR2_X1    g06652(.A1(new_n6844_), .A2(new_n6843_), .ZN(new_n6845_));
  NOR3_X1    g06653(.A1(new_n6845_), .A2(new_n6458_), .A3(new_n6842_), .ZN(new_n6846_));
  NOR3_X1    g06654(.A1(new_n6824_), .A2(new_n6458_), .A3(new_n6845_), .ZN(new_n6847_));
  INV_X1     g06655(.I(new_n6847_), .ZN(new_n6848_));
  AOI22_X1   g06656(.A1(new_n6848_), .A2(new_n6842_), .B1(\asqrt[32] ), .B2(new_n6846_), .ZN(new_n6849_));
  INV_X1     g06657(.I(new_n6849_), .ZN(new_n6850_));
  NAND2_X1   g06658(.A1(new_n6831_), .A2(new_n4071_), .ZN(new_n6851_));
  OAI21_X1   g06659(.A1(new_n6840_), .A2(new_n6851_), .B(new_n6850_), .ZN(new_n6852_));
  AOI21_X1   g06660(.A1(new_n6852_), .A2(new_n6841_), .B(new_n3782_), .ZN(new_n6853_));
  INV_X1     g06661(.I(new_n6472_), .ZN(new_n6854_));
  NOR3_X1    g06662(.A1(new_n6824_), .A2(new_n6467_), .A3(new_n6473_), .ZN(new_n6855_));
  INV_X1     g06663(.I(new_n6855_), .ZN(new_n6856_));
  NOR3_X1    g06664(.A1(new_n6467_), .A2(new_n6854_), .A3(new_n6473_), .ZN(new_n6857_));
  AOI22_X1   g06665(.A1(new_n6856_), .A2(new_n6854_), .B1(\asqrt[32] ), .B2(new_n6857_), .ZN(new_n6858_));
  OAI21_X1   g06666(.A1(new_n6838_), .A2(new_n6839_), .B(new_n6831_), .ZN(new_n6859_));
  AOI21_X1   g06667(.A1(new_n6859_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n6860_));
  AOI21_X1   g06668(.A1(new_n6860_), .A2(new_n6852_), .B(new_n6858_), .ZN(new_n6861_));
  OAI21_X1   g06669(.A1(new_n6861_), .A2(new_n6853_), .B(\asqrt[42] ), .ZN(new_n6862_));
  INV_X1     g06670(.I(new_n6862_), .ZN(new_n6863_));
  NOR2_X1    g06671(.A1(new_n6474_), .A2(new_n6482_), .ZN(new_n6864_));
  INV_X1     g06672(.I(new_n6864_), .ZN(new_n6865_));
  AND3_X2    g06673(.A1(new_n6865_), .A2(new_n6475_), .A3(new_n6480_), .Z(new_n6866_));
  NAND3_X1   g06674(.A1(\asqrt[32] ), .A2(new_n6475_), .A3(new_n6865_), .ZN(new_n6867_));
  AOI22_X1   g06675(.A1(new_n6867_), .A2(new_n6481_), .B1(\asqrt[32] ), .B2(new_n6866_), .ZN(new_n6868_));
  NOR3_X1    g06676(.A1(new_n6861_), .A2(new_n6853_), .A3(\asqrt[42] ), .ZN(new_n6869_));
  NOR2_X1    g06677(.A1(new_n6869_), .A2(new_n6868_), .ZN(new_n6870_));
  OAI21_X1   g06678(.A1(new_n6870_), .A2(new_n6863_), .B(\asqrt[43] ), .ZN(new_n6871_));
  INV_X1     g06679(.I(new_n6488_), .ZN(new_n6872_));
  INV_X1     g06680(.I(new_n6483_), .ZN(new_n6873_));
  INV_X1     g06681(.I(new_n6490_), .ZN(new_n6874_));
  NOR2_X1    g06682(.A1(new_n6874_), .A2(new_n6873_), .ZN(new_n6875_));
  NOR3_X1    g06683(.A1(new_n6824_), .A2(new_n6484_), .A3(new_n6875_), .ZN(new_n6876_));
  INV_X1     g06684(.I(new_n6876_), .ZN(new_n6877_));
  NOR3_X1    g06685(.A1(new_n6875_), .A2(new_n6484_), .A3(new_n6872_), .ZN(new_n6878_));
  AOI22_X1   g06686(.A1(new_n6877_), .A2(new_n6872_), .B1(\asqrt[32] ), .B2(new_n6878_), .ZN(new_n6879_));
  INV_X1     g06687(.I(new_n6879_), .ZN(new_n6880_));
  NAND2_X1   g06688(.A1(new_n6862_), .A2(new_n3218_), .ZN(new_n6881_));
  OAI21_X1   g06689(.A1(new_n6870_), .A2(new_n6881_), .B(new_n6880_), .ZN(new_n6882_));
  AOI21_X1   g06690(.A1(new_n6882_), .A2(new_n6871_), .B(new_n2954_), .ZN(new_n6883_));
  INV_X1     g06691(.I(new_n6498_), .ZN(new_n6884_));
  NOR3_X1    g06692(.A1(new_n6493_), .A2(new_n6499_), .A3(new_n6884_), .ZN(new_n6885_));
  NOR3_X1    g06693(.A1(new_n6824_), .A2(new_n6493_), .A3(new_n6499_), .ZN(new_n6886_));
  INV_X1     g06694(.I(new_n6886_), .ZN(new_n6887_));
  AOI22_X1   g06695(.A1(new_n6887_), .A2(new_n6884_), .B1(\asqrt[32] ), .B2(new_n6885_), .ZN(new_n6888_));
  OAI21_X1   g06696(.A1(new_n6868_), .A2(new_n6869_), .B(new_n6862_), .ZN(new_n6889_));
  AOI21_X1   g06697(.A1(new_n6889_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n6890_));
  AOI21_X1   g06698(.A1(new_n6890_), .A2(new_n6882_), .B(new_n6888_), .ZN(new_n6891_));
  OAI21_X1   g06699(.A1(new_n6891_), .A2(new_n6883_), .B(\asqrt[45] ), .ZN(new_n6892_));
  INV_X1     g06700(.I(new_n6892_), .ZN(new_n6893_));
  INV_X1     g06701(.I(new_n6501_), .ZN(new_n6894_));
  NOR2_X1    g06702(.A1(new_n6500_), .A2(new_n6507_), .ZN(new_n6895_));
  NOR3_X1    g06703(.A1(new_n6824_), .A2(new_n6894_), .A3(new_n6895_), .ZN(new_n6896_));
  INV_X1     g06704(.I(new_n6896_), .ZN(new_n6897_));
  NOR3_X1    g06705(.A1(new_n6894_), .A2(new_n6506_), .A3(new_n6895_), .ZN(new_n6898_));
  AOI22_X1   g06706(.A1(new_n6897_), .A2(new_n6506_), .B1(\asqrt[32] ), .B2(new_n6898_), .ZN(new_n6899_));
  NOR3_X1    g06707(.A1(new_n6891_), .A2(new_n6883_), .A3(\asqrt[45] ), .ZN(new_n6900_));
  NOR2_X1    g06708(.A1(new_n6900_), .A2(new_n6899_), .ZN(new_n6901_));
  OAI21_X1   g06709(.A1(new_n6901_), .A2(new_n6893_), .B(\asqrt[46] ), .ZN(new_n6902_));
  INV_X1     g06710(.I(new_n6515_), .ZN(new_n6903_));
  INV_X1     g06711(.I(new_n6508_), .ZN(new_n6904_));
  INV_X1     g06712(.I(new_n6517_), .ZN(new_n6905_));
  NOR2_X1    g06713(.A1(new_n6905_), .A2(new_n6904_), .ZN(new_n6906_));
  NOR3_X1    g06714(.A1(new_n6906_), .A2(new_n6509_), .A3(new_n6903_), .ZN(new_n6907_));
  NOR3_X1    g06715(.A1(new_n6824_), .A2(new_n6509_), .A3(new_n6906_), .ZN(new_n6908_));
  INV_X1     g06716(.I(new_n6908_), .ZN(new_n6909_));
  AOI22_X1   g06717(.A1(new_n6909_), .A2(new_n6903_), .B1(\asqrt[32] ), .B2(new_n6907_), .ZN(new_n6910_));
  INV_X1     g06718(.I(new_n6910_), .ZN(new_n6911_));
  NAND2_X1   g06719(.A1(new_n6892_), .A2(new_n2465_), .ZN(new_n6912_));
  OAI21_X1   g06720(.A1(new_n6901_), .A2(new_n6912_), .B(new_n6911_), .ZN(new_n6913_));
  AOI21_X1   g06721(.A1(new_n6913_), .A2(new_n6902_), .B(new_n2229_), .ZN(new_n6914_));
  INV_X1     g06722(.I(new_n6528_), .ZN(new_n6915_));
  NOR3_X1    g06723(.A1(new_n6824_), .A2(new_n6520_), .A3(new_n6529_), .ZN(new_n6916_));
  INV_X1     g06724(.I(new_n6916_), .ZN(new_n6917_));
  NOR3_X1    g06725(.A1(new_n6520_), .A2(new_n6529_), .A3(new_n6915_), .ZN(new_n6918_));
  AOI22_X1   g06726(.A1(new_n6917_), .A2(new_n6915_), .B1(\asqrt[32] ), .B2(new_n6918_), .ZN(new_n6919_));
  OAI21_X1   g06727(.A1(new_n6899_), .A2(new_n6900_), .B(new_n6892_), .ZN(new_n6920_));
  AOI21_X1   g06728(.A1(new_n6920_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n6921_));
  AOI21_X1   g06729(.A1(new_n6921_), .A2(new_n6913_), .B(new_n6919_), .ZN(new_n6922_));
  OAI21_X1   g06730(.A1(new_n6922_), .A2(new_n6914_), .B(\asqrt[48] ), .ZN(new_n6923_));
  INV_X1     g06731(.I(new_n6923_), .ZN(new_n6924_));
  NOR2_X1    g06732(.A1(new_n6530_), .A2(new_n6537_), .ZN(new_n6925_));
  INV_X1     g06733(.I(new_n6925_), .ZN(new_n6926_));
  AND3_X2    g06734(.A1(new_n6926_), .A2(new_n6531_), .A3(new_n6535_), .Z(new_n6927_));
  NAND3_X1   g06735(.A1(\asqrt[32] ), .A2(new_n6531_), .A3(new_n6926_), .ZN(new_n6928_));
  AOI22_X1   g06736(.A1(new_n6928_), .A2(new_n6536_), .B1(\asqrt[32] ), .B2(new_n6927_), .ZN(new_n6929_));
  NOR3_X1    g06737(.A1(new_n6922_), .A2(new_n6914_), .A3(\asqrt[48] ), .ZN(new_n6930_));
  NOR2_X1    g06738(.A1(new_n6930_), .A2(new_n6929_), .ZN(new_n6931_));
  OAI21_X1   g06739(.A1(new_n6931_), .A2(new_n6924_), .B(\asqrt[49] ), .ZN(new_n6932_));
  INV_X1     g06740(.I(new_n6545_), .ZN(new_n6933_));
  NAND2_X1   g06741(.A1(new_n6547_), .A2(new_n6538_), .ZN(new_n6934_));
  NAND3_X1   g06742(.A1(\asqrt[32] ), .A2(new_n6590_), .A3(new_n6934_), .ZN(new_n6935_));
  AND3_X2    g06743(.A1(new_n6590_), .A2(new_n6545_), .A3(new_n6934_), .Z(new_n6936_));
  AOI22_X1   g06744(.A1(new_n6935_), .A2(new_n6933_), .B1(\asqrt[32] ), .B2(new_n6936_), .ZN(new_n6937_));
  INV_X1     g06745(.I(new_n6937_), .ZN(new_n6938_));
  NAND2_X1   g06746(.A1(new_n6923_), .A2(new_n1806_), .ZN(new_n6939_));
  OAI21_X1   g06747(.A1(new_n6931_), .A2(new_n6939_), .B(new_n6938_), .ZN(new_n6940_));
  AOI21_X1   g06748(.A1(new_n6940_), .A2(new_n6932_), .B(new_n1612_), .ZN(new_n6941_));
  NOR3_X1    g06749(.A1(new_n6550_), .A2(new_n6559_), .A3(new_n6589_), .ZN(new_n6942_));
  NOR3_X1    g06750(.A1(new_n6824_), .A2(new_n6550_), .A3(new_n6559_), .ZN(new_n6943_));
  INV_X1     g06751(.I(new_n6943_), .ZN(new_n6944_));
  AOI22_X1   g06752(.A1(new_n6944_), .A2(new_n6589_), .B1(\asqrt[32] ), .B2(new_n6942_), .ZN(new_n6945_));
  OAI21_X1   g06753(.A1(new_n6929_), .A2(new_n6930_), .B(new_n6923_), .ZN(new_n6946_));
  AOI21_X1   g06754(.A1(new_n6946_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n6947_));
  AOI21_X1   g06755(.A1(new_n6947_), .A2(new_n6940_), .B(new_n6945_), .ZN(new_n6948_));
  OAI21_X1   g06756(.A1(new_n6948_), .A2(new_n6941_), .B(\asqrt[51] ), .ZN(new_n6949_));
  INV_X1     g06757(.I(new_n6949_), .ZN(new_n6950_));
  NOR2_X1    g06758(.A1(new_n6560_), .A2(new_n6567_), .ZN(new_n6951_));
  NOR3_X1    g06759(.A1(new_n6824_), .A2(new_n6593_), .A3(new_n6951_), .ZN(new_n6952_));
  INV_X1     g06760(.I(new_n6952_), .ZN(new_n6953_));
  NOR3_X1    g06761(.A1(new_n6593_), .A2(new_n6951_), .A3(new_n6566_), .ZN(new_n6954_));
  AOI22_X1   g06762(.A1(new_n6953_), .A2(new_n6566_), .B1(\asqrt[32] ), .B2(new_n6954_), .ZN(new_n6955_));
  NOR3_X1    g06763(.A1(new_n6948_), .A2(new_n6941_), .A3(\asqrt[51] ), .ZN(new_n6956_));
  NOR2_X1    g06764(.A1(new_n6956_), .A2(new_n6955_), .ZN(new_n6957_));
  OAI21_X1   g06765(.A1(new_n6957_), .A2(new_n6950_), .B(\asqrt[52] ), .ZN(new_n6958_));
  NOR2_X1    g06766(.A1(new_n6605_), .A2(new_n6595_), .ZN(new_n6959_));
  NOR3_X1    g06767(.A1(new_n6959_), .A2(new_n6569_), .A3(new_n6604_), .ZN(new_n6960_));
  NOR3_X1    g06768(.A1(new_n6824_), .A2(new_n6569_), .A3(new_n6959_), .ZN(new_n6961_));
  INV_X1     g06769(.I(new_n6961_), .ZN(new_n6962_));
  AOI22_X1   g06770(.A1(new_n6962_), .A2(new_n6604_), .B1(\asqrt[32] ), .B2(new_n6960_), .ZN(new_n6963_));
  INV_X1     g06771(.I(new_n6963_), .ZN(new_n6964_));
  NAND2_X1   g06772(.A1(new_n6949_), .A2(new_n1256_), .ZN(new_n6965_));
  OAI21_X1   g06773(.A1(new_n6957_), .A2(new_n6965_), .B(new_n6964_), .ZN(new_n6966_));
  AOI21_X1   g06774(.A1(new_n6966_), .A2(new_n6958_), .B(new_n1103_), .ZN(new_n6967_));
  NOR3_X1    g06775(.A1(new_n6824_), .A2(new_n6607_), .A3(new_n6641_), .ZN(new_n6968_));
  INV_X1     g06776(.I(new_n6968_), .ZN(new_n6969_));
  NOR3_X1    g06777(.A1(new_n6607_), .A2(new_n6641_), .A3(new_n6588_), .ZN(new_n6970_));
  AOI22_X1   g06778(.A1(new_n6969_), .A2(new_n6588_), .B1(\asqrt[32] ), .B2(new_n6970_), .ZN(new_n6971_));
  OAI21_X1   g06779(.A1(new_n6955_), .A2(new_n6956_), .B(new_n6949_), .ZN(new_n6972_));
  AOI21_X1   g06780(.A1(new_n6972_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n6973_));
  AOI21_X1   g06781(.A1(new_n6973_), .A2(new_n6966_), .B(new_n6971_), .ZN(new_n6974_));
  OAI21_X1   g06782(.A1(new_n6974_), .A2(new_n6967_), .B(\asqrt[54] ), .ZN(new_n6975_));
  INV_X1     g06783(.I(new_n6975_), .ZN(new_n6976_));
  NOR2_X1    g06784(.A1(new_n6630_), .A2(new_n6619_), .ZN(new_n6977_));
  NOR3_X1    g06785(.A1(new_n6599_), .A2(new_n6977_), .A3(new_n6629_), .ZN(new_n6978_));
  NOR3_X1    g06786(.A1(new_n6824_), .A2(new_n6599_), .A3(new_n6977_), .ZN(new_n6979_));
  INV_X1     g06787(.I(new_n6979_), .ZN(new_n6980_));
  AOI22_X1   g06788(.A1(new_n6980_), .A2(new_n6629_), .B1(\asqrt[32] ), .B2(new_n6978_), .ZN(new_n6981_));
  NOR3_X1    g06789(.A1(new_n6974_), .A2(new_n6967_), .A3(\asqrt[54] ), .ZN(new_n6982_));
  NOR2_X1    g06790(.A1(new_n6982_), .A2(new_n6981_), .ZN(new_n6983_));
  OAI21_X1   g06791(.A1(new_n6983_), .A2(new_n6976_), .B(\asqrt[55] ), .ZN(new_n6984_));
  NOR2_X1    g06792(.A1(new_n6621_), .A2(new_n6609_), .ZN(new_n6985_));
  NOR3_X1    g06793(.A1(new_n6824_), .A2(new_n6632_), .A3(new_n6985_), .ZN(new_n6986_));
  INV_X1     g06794(.I(new_n6986_), .ZN(new_n6987_));
  NOR3_X1    g06795(.A1(new_n6985_), .A2(new_n6632_), .A3(new_n6617_), .ZN(new_n6988_));
  AOI22_X1   g06796(.A1(new_n6987_), .A2(new_n6617_), .B1(\asqrt[32] ), .B2(new_n6988_), .ZN(new_n6989_));
  INV_X1     g06797(.I(new_n6989_), .ZN(new_n6990_));
  NAND2_X1   g06798(.A1(new_n6975_), .A2(new_n823_), .ZN(new_n6991_));
  OAI21_X1   g06799(.A1(new_n6983_), .A2(new_n6991_), .B(new_n6990_), .ZN(new_n6992_));
  AOI21_X1   g06800(.A1(new_n6992_), .A2(new_n6984_), .B(new_n703_), .ZN(new_n6993_));
  NOR3_X1    g06801(.A1(new_n6623_), .A2(new_n6655_), .A3(new_n6666_), .ZN(new_n6994_));
  NOR3_X1    g06802(.A1(new_n6824_), .A2(new_n6623_), .A3(new_n6655_), .ZN(new_n6995_));
  INV_X1     g06803(.I(new_n6995_), .ZN(new_n6996_));
  AOI22_X1   g06804(.A1(new_n6996_), .A2(new_n6666_), .B1(\asqrt[32] ), .B2(new_n6994_), .ZN(new_n6997_));
  OAI21_X1   g06805(.A1(new_n6981_), .A2(new_n6982_), .B(new_n6975_), .ZN(new_n6998_));
  AOI21_X1   g06806(.A1(new_n6998_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n6999_));
  AOI21_X1   g06807(.A1(new_n6999_), .A2(new_n6992_), .B(new_n6997_), .ZN(new_n7000_));
  OAI21_X1   g06808(.A1(new_n7000_), .A2(new_n6993_), .B(\asqrt[57] ), .ZN(new_n7001_));
  NOR2_X1    g06809(.A1(new_n6646_), .A2(new_n6634_), .ZN(new_n7002_));
  NOR3_X1    g06810(.A1(new_n6824_), .A2(new_n6669_), .A3(new_n7002_), .ZN(new_n7003_));
  INV_X1     g06811(.I(new_n7003_), .ZN(new_n7004_));
  NOR3_X1    g06812(.A1(new_n6669_), .A2(new_n7002_), .A3(new_n6640_), .ZN(new_n7005_));
  AOI22_X1   g06813(.A1(new_n7004_), .A2(new_n6640_), .B1(\asqrt[32] ), .B2(new_n7005_), .ZN(new_n7006_));
  INV_X1     g06814(.I(new_n7006_), .ZN(new_n7007_));
  INV_X1     g06815(.I(new_n6981_), .ZN(new_n7008_));
  INV_X1     g06816(.I(new_n6955_), .ZN(new_n7009_));
  INV_X1     g06817(.I(new_n6929_), .ZN(new_n7010_));
  INV_X1     g06818(.I(new_n6899_), .ZN(new_n7011_));
  INV_X1     g06819(.I(new_n6868_), .ZN(new_n7012_));
  INV_X1     g06820(.I(new_n6838_), .ZN(new_n7013_));
  NAND2_X1   g06821(.A1(new_n6758_), .A2(new_n6769_), .ZN(new_n7014_));
  OAI21_X1   g06822(.A1(new_n6753_), .A2(new_n6757_), .B(new_n6760_), .ZN(new_n7015_));
  NAND2_X1   g06823(.A1(new_n7015_), .A2(\a[65] ), .ZN(new_n7016_));
  NAND3_X1   g06824(.A1(new_n7014_), .A2(new_n7016_), .A3(new_n6777_), .ZN(new_n7017_));
  AOI21_X1   g06825(.A1(new_n7017_), .A2(new_n6794_), .B(new_n6077_), .ZN(new_n7018_));
  OAI21_X1   g06826(.A1(new_n6781_), .A2(new_n6772_), .B(\a[66] ), .ZN(new_n7019_));
  NAND3_X1   g06827(.A1(new_n6782_), .A2(new_n6777_), .A3(new_n6360_), .ZN(new_n7020_));
  NAND2_X1   g06828(.A1(new_n6758_), .A2(new_n6750_), .ZN(new_n7021_));
  AOI21_X1   g06829(.A1(new_n7021_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n7022_));
  AOI22_X1   g06830(.A1(new_n7017_), .A2(new_n7022_), .B1(new_n7019_), .B2(new_n7020_), .ZN(new_n7023_));
  OAI21_X1   g06831(.A1(new_n7023_), .A2(new_n7018_), .B(\asqrt[35] ), .ZN(new_n7024_));
  NAND2_X1   g06832(.A1(new_n7024_), .A2(new_n5277_), .ZN(new_n7025_));
  OAI21_X1   g06833(.A1(new_n7025_), .A2(new_n6799_), .B(new_n6807_), .ZN(new_n7026_));
  AOI21_X1   g06834(.A1(new_n7026_), .A2(new_n6800_), .B(new_n5024_), .ZN(new_n7027_));
  INV_X1     g06835(.I(new_n6793_), .ZN(new_n7028_));
  AOI21_X1   g06836(.A1(\a[65] ), .A2(new_n7015_), .B(new_n6772_), .ZN(new_n7029_));
  AOI21_X1   g06837(.A1(new_n7029_), .A2(new_n7014_), .B(new_n6759_), .ZN(new_n7030_));
  OAI21_X1   g06838(.A1(new_n7030_), .A2(new_n6077_), .B(new_n5708_), .ZN(new_n7031_));
  OAI21_X1   g06839(.A1(new_n7031_), .A2(new_n7023_), .B(new_n7028_), .ZN(new_n7032_));
  NAND2_X1   g06840(.A1(new_n7032_), .A2(new_n7024_), .ZN(new_n7033_));
  AOI21_X1   g06841(.A1(new_n7033_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n7034_));
  AOI21_X1   g06842(.A1(new_n7034_), .A2(new_n7026_), .B(new_n6817_), .ZN(new_n7035_));
  OAI21_X1   g06843(.A1(new_n7035_), .A2(new_n7027_), .B(\asqrt[38] ), .ZN(new_n7036_));
  NAND2_X1   g06844(.A1(new_n7036_), .A2(new_n4298_), .ZN(new_n7037_));
  OAI21_X1   g06845(.A1(new_n7037_), .A2(new_n6830_), .B(new_n7013_), .ZN(new_n7038_));
  NAND3_X1   g06846(.A1(new_n7038_), .A2(new_n4071_), .A3(new_n6831_), .ZN(new_n7039_));
  AOI22_X1   g06847(.A1(new_n7039_), .A2(new_n6850_), .B1(new_n6859_), .B2(\asqrt[40] ), .ZN(new_n7040_));
  OAI21_X1   g06848(.A1(new_n7040_), .A2(new_n3782_), .B(new_n3419_), .ZN(new_n7041_));
  OAI21_X1   g06849(.A1(new_n7041_), .A2(new_n6861_), .B(new_n7012_), .ZN(new_n7042_));
  AOI21_X1   g06850(.A1(new_n7042_), .A2(new_n6862_), .B(new_n3218_), .ZN(new_n7043_));
  AOI21_X1   g06851(.A1(new_n7038_), .A2(new_n6831_), .B(new_n4071_), .ZN(new_n7044_));
  NOR3_X1    g06852(.A1(new_n7035_), .A2(new_n7027_), .A3(\asqrt[38] ), .ZN(new_n7045_));
  OAI21_X1   g06853(.A1(new_n6827_), .A2(new_n7045_), .B(new_n7036_), .ZN(new_n7046_));
  AOI21_X1   g06854(.A1(new_n7046_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n7047_));
  AOI21_X1   g06855(.A1(new_n7047_), .A2(new_n7038_), .B(new_n6849_), .ZN(new_n7048_));
  NOR3_X1    g06856(.A1(new_n7048_), .A2(\asqrt[41] ), .A3(new_n7044_), .ZN(new_n7049_));
  OAI22_X1   g06857(.A1(new_n7049_), .A2(new_n6858_), .B1(new_n7040_), .B2(new_n3782_), .ZN(new_n7050_));
  AOI21_X1   g06858(.A1(new_n7050_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n7051_));
  AOI21_X1   g06859(.A1(new_n7051_), .A2(new_n7042_), .B(new_n6879_), .ZN(new_n7052_));
  OAI21_X1   g06860(.A1(new_n7052_), .A2(new_n7043_), .B(\asqrt[44] ), .ZN(new_n7053_));
  NAND2_X1   g06861(.A1(new_n7053_), .A2(new_n2641_), .ZN(new_n7054_));
  OAI21_X1   g06862(.A1(new_n7054_), .A2(new_n6891_), .B(new_n7011_), .ZN(new_n7055_));
  AOI21_X1   g06863(.A1(new_n7055_), .A2(new_n6892_), .B(new_n2465_), .ZN(new_n7056_));
  NOR3_X1    g06864(.A1(new_n7052_), .A2(\asqrt[44] ), .A3(new_n7043_), .ZN(new_n7057_));
  OAI21_X1   g06865(.A1(new_n6888_), .A2(new_n7057_), .B(new_n7053_), .ZN(new_n7058_));
  AOI21_X1   g06866(.A1(new_n7058_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n7059_));
  AOI21_X1   g06867(.A1(new_n7059_), .A2(new_n7055_), .B(new_n6910_), .ZN(new_n7060_));
  OAI21_X1   g06868(.A1(new_n7060_), .A2(new_n7056_), .B(\asqrt[47] ), .ZN(new_n7061_));
  NAND2_X1   g06869(.A1(new_n7061_), .A2(new_n1956_), .ZN(new_n7062_));
  OAI21_X1   g06870(.A1(new_n7062_), .A2(new_n6922_), .B(new_n7010_), .ZN(new_n7063_));
  AOI21_X1   g06871(.A1(new_n7063_), .A2(new_n6923_), .B(new_n1806_), .ZN(new_n7064_));
  NOR3_X1    g06872(.A1(new_n7060_), .A2(\asqrt[47] ), .A3(new_n7056_), .ZN(new_n7065_));
  OAI21_X1   g06873(.A1(new_n6919_), .A2(new_n7065_), .B(new_n7061_), .ZN(new_n7066_));
  AOI21_X1   g06874(.A1(new_n7066_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n7067_));
  AOI21_X1   g06875(.A1(new_n7067_), .A2(new_n7063_), .B(new_n6937_), .ZN(new_n7068_));
  OAI21_X1   g06876(.A1(new_n7068_), .A2(new_n7064_), .B(\asqrt[50] ), .ZN(new_n7069_));
  NAND2_X1   g06877(.A1(new_n7069_), .A2(new_n1376_), .ZN(new_n7070_));
  OAI21_X1   g06878(.A1(new_n7070_), .A2(new_n6948_), .B(new_n7009_), .ZN(new_n7071_));
  AOI21_X1   g06879(.A1(new_n7071_), .A2(new_n6949_), .B(new_n1256_), .ZN(new_n7072_));
  NOR3_X1    g06880(.A1(new_n7068_), .A2(\asqrt[50] ), .A3(new_n7064_), .ZN(new_n7073_));
  OAI21_X1   g06881(.A1(new_n6945_), .A2(new_n7073_), .B(new_n7069_), .ZN(new_n7074_));
  AOI21_X1   g06882(.A1(new_n7074_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n7075_));
  AOI21_X1   g06883(.A1(new_n7075_), .A2(new_n7071_), .B(new_n6963_), .ZN(new_n7076_));
  OAI21_X1   g06884(.A1(new_n7076_), .A2(new_n7072_), .B(\asqrt[53] ), .ZN(new_n7077_));
  NAND2_X1   g06885(.A1(new_n7077_), .A2(new_n904_), .ZN(new_n7078_));
  OAI21_X1   g06886(.A1(new_n7078_), .A2(new_n6974_), .B(new_n7008_), .ZN(new_n7079_));
  AOI21_X1   g06887(.A1(new_n7079_), .A2(new_n6975_), .B(new_n823_), .ZN(new_n7080_));
  NOR3_X1    g06888(.A1(new_n7076_), .A2(\asqrt[53] ), .A3(new_n7072_), .ZN(new_n7081_));
  OAI21_X1   g06889(.A1(new_n6971_), .A2(new_n7081_), .B(new_n7077_), .ZN(new_n7082_));
  AOI21_X1   g06890(.A1(new_n7082_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n7083_));
  AOI21_X1   g06891(.A1(new_n7083_), .A2(new_n7079_), .B(new_n6989_), .ZN(new_n7084_));
  OAI21_X1   g06892(.A1(new_n7084_), .A2(new_n7080_), .B(\asqrt[56] ), .ZN(new_n7085_));
  NAND2_X1   g06893(.A1(new_n7085_), .A2(new_n531_), .ZN(new_n7086_));
  OAI21_X1   g06894(.A1(new_n7086_), .A2(new_n7000_), .B(new_n7007_), .ZN(new_n7087_));
  AOI21_X1   g06895(.A1(new_n7087_), .A2(new_n7001_), .B(new_n436_), .ZN(new_n7088_));
  NOR2_X1    g06896(.A1(new_n6681_), .A2(new_n6671_), .ZN(new_n7089_));
  NOR3_X1    g06897(.A1(new_n7089_), .A2(new_n6648_), .A3(new_n6680_), .ZN(new_n7090_));
  NOR3_X1    g06898(.A1(new_n6824_), .A2(new_n6648_), .A3(new_n7089_), .ZN(new_n7091_));
  INV_X1     g06899(.I(new_n7091_), .ZN(new_n7092_));
  AOI22_X1   g06900(.A1(new_n7092_), .A2(new_n6680_), .B1(\asqrt[32] ), .B2(new_n7090_), .ZN(new_n7093_));
  NOR3_X1    g06901(.A1(new_n7084_), .A2(\asqrt[56] ), .A3(new_n7080_), .ZN(new_n7094_));
  OAI21_X1   g06902(.A1(new_n6997_), .A2(new_n7094_), .B(new_n7085_), .ZN(new_n7095_));
  AOI21_X1   g06903(.A1(new_n7095_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n7096_));
  AOI21_X1   g06904(.A1(new_n7096_), .A2(new_n7087_), .B(new_n7093_), .ZN(new_n7097_));
  OAI21_X1   g06905(.A1(new_n7097_), .A2(new_n7088_), .B(\asqrt[59] ), .ZN(new_n7098_));
  NOR3_X1    g06906(.A1(new_n6824_), .A2(new_n6683_), .A3(new_n6717_), .ZN(new_n7099_));
  INV_X1     g06907(.I(new_n7099_), .ZN(new_n7100_));
  NOR3_X1    g06908(.A1(new_n6683_), .A2(new_n6717_), .A3(new_n6665_), .ZN(new_n7101_));
  AOI22_X1   g06909(.A1(new_n7100_), .A2(new_n6665_), .B1(\asqrt[32] ), .B2(new_n7101_), .ZN(new_n7102_));
  INV_X1     g06910(.I(new_n7102_), .ZN(new_n7103_));
  INV_X1     g06911(.I(new_n7001_), .ZN(new_n7104_));
  NOR3_X1    g06912(.A1(new_n7000_), .A2(new_n6993_), .A3(\asqrt[57] ), .ZN(new_n7105_));
  NOR2_X1    g06913(.A1(new_n7105_), .A2(new_n7006_), .ZN(new_n7106_));
  OAI21_X1   g06914(.A1(new_n7106_), .A2(new_n7104_), .B(\asqrt[58] ), .ZN(new_n7107_));
  NAND2_X1   g06915(.A1(new_n7107_), .A2(new_n327_), .ZN(new_n7108_));
  OAI21_X1   g06916(.A1(new_n7108_), .A2(new_n7097_), .B(new_n7103_), .ZN(new_n7109_));
  AOI21_X1   g06917(.A1(new_n7109_), .A2(new_n7098_), .B(new_n306_), .ZN(new_n7110_));
  NOR2_X1    g06918(.A1(new_n6706_), .A2(new_n6695_), .ZN(new_n7111_));
  NOR3_X1    g06919(.A1(new_n6675_), .A2(new_n7111_), .A3(new_n6705_), .ZN(new_n7112_));
  NOR3_X1    g06920(.A1(new_n6824_), .A2(new_n6675_), .A3(new_n7111_), .ZN(new_n7113_));
  INV_X1     g06921(.I(new_n7113_), .ZN(new_n7114_));
  AOI22_X1   g06922(.A1(new_n7114_), .A2(new_n6705_), .B1(\asqrt[32] ), .B2(new_n7112_), .ZN(new_n7115_));
  INV_X1     g06923(.I(new_n7093_), .ZN(new_n7116_));
  NAND2_X1   g06924(.A1(new_n7001_), .A2(new_n436_), .ZN(new_n7117_));
  OAI21_X1   g06925(.A1(new_n7106_), .A2(new_n7117_), .B(new_n7116_), .ZN(new_n7118_));
  AOI21_X1   g06926(.A1(new_n7118_), .A2(new_n7107_), .B(new_n327_), .ZN(new_n7119_));
  NOR2_X1    g06927(.A1(new_n7119_), .A2(\asqrt[60] ), .ZN(new_n7120_));
  AOI21_X1   g06928(.A1(new_n7120_), .A2(new_n7109_), .B(new_n7115_), .ZN(new_n7121_));
  OAI21_X1   g06929(.A1(new_n7121_), .A2(new_n7110_), .B(\asqrt[61] ), .ZN(new_n7122_));
  NOR2_X1    g06930(.A1(new_n6697_), .A2(new_n6685_), .ZN(new_n7123_));
  NOR3_X1    g06931(.A1(new_n6824_), .A2(new_n6708_), .A3(new_n7123_), .ZN(new_n7124_));
  INV_X1     g06932(.I(new_n7124_), .ZN(new_n7125_));
  NOR3_X1    g06933(.A1(new_n7123_), .A2(new_n6708_), .A3(new_n6693_), .ZN(new_n7126_));
  AOI22_X1   g06934(.A1(new_n7125_), .A2(new_n6693_), .B1(\asqrt[32] ), .B2(new_n7126_), .ZN(new_n7127_));
  INV_X1     g06935(.I(new_n7127_), .ZN(new_n7128_));
  OAI21_X1   g06936(.A1(new_n7006_), .A2(new_n7105_), .B(new_n7001_), .ZN(new_n7129_));
  AOI21_X1   g06937(.A1(new_n7129_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n7130_));
  AOI21_X1   g06938(.A1(new_n7130_), .A2(new_n7118_), .B(new_n7102_), .ZN(new_n7131_));
  OAI21_X1   g06939(.A1(new_n7131_), .A2(new_n7119_), .B(\asqrt[60] ), .ZN(new_n7132_));
  NAND2_X1   g06940(.A1(new_n7132_), .A2(new_n218_), .ZN(new_n7133_));
  OAI21_X1   g06941(.A1(new_n7133_), .A2(new_n7121_), .B(new_n7128_), .ZN(new_n7134_));
  AOI21_X1   g06942(.A1(new_n7134_), .A2(new_n7122_), .B(new_n207_), .ZN(new_n7135_));
  NOR3_X1    g06943(.A1(new_n6699_), .A2(new_n6733_), .A3(new_n6761_), .ZN(new_n7136_));
  NOR3_X1    g06944(.A1(new_n6824_), .A2(new_n6699_), .A3(new_n6733_), .ZN(new_n7137_));
  INV_X1     g06945(.I(new_n7137_), .ZN(new_n7138_));
  AOI22_X1   g06946(.A1(new_n7138_), .A2(new_n6761_), .B1(\asqrt[32] ), .B2(new_n7136_), .ZN(new_n7139_));
  NOR3_X1    g06947(.A1(new_n7131_), .A2(new_n7119_), .A3(\asqrt[60] ), .ZN(new_n7140_));
  OAI21_X1   g06948(.A1(new_n7115_), .A2(new_n7140_), .B(new_n7132_), .ZN(new_n7141_));
  AOI21_X1   g06949(.A1(new_n7141_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n7142_));
  AOI21_X1   g06950(.A1(new_n7142_), .A2(new_n7134_), .B(new_n7139_), .ZN(new_n7143_));
  AND3_X2    g06951(.A1(new_n6711_), .A2(new_n6764_), .A3(new_n6715_), .Z(new_n7144_));
  NAND2_X1   g06952(.A1(\asqrt[32] ), .A2(new_n7144_), .ZN(new_n7145_));
  INV_X1     g06953(.I(new_n7145_), .ZN(new_n7146_));
  AND2_X2    g06954(.A1(new_n6711_), .A2(new_n6764_), .Z(new_n7147_));
  AOI21_X1   g06955(.A1(\asqrt[32] ), .A2(new_n7147_), .B(new_n6715_), .ZN(new_n7148_));
  NOR2_X1    g06956(.A1(new_n7146_), .A2(new_n7148_), .ZN(new_n7149_));
  NOR3_X1    g06957(.A1(new_n6824_), .A2(new_n6765_), .A3(new_n6755_), .ZN(new_n7150_));
  NOR3_X1    g06958(.A1(new_n7149_), .A2(new_n6778_), .A3(new_n7150_), .ZN(new_n7151_));
  OAI21_X1   g06959(.A1(new_n7143_), .A2(new_n7135_), .B(new_n7151_), .ZN(new_n7152_));
  NAND2_X1   g06960(.A1(new_n7152_), .A2(new_n193_), .ZN(new_n7153_));
  INV_X1     g06961(.I(new_n7139_), .ZN(new_n7154_));
  NAND3_X1   g06962(.A1(new_n7134_), .A2(new_n7122_), .A3(new_n207_), .ZN(new_n7155_));
  NAND2_X1   g06963(.A1(new_n7155_), .A2(new_n7154_), .ZN(new_n7156_));
  INV_X1     g06964(.I(new_n7149_), .ZN(new_n7157_));
  NOR2_X1    g06965(.A1(new_n7135_), .A2(new_n7157_), .ZN(new_n7158_));
  AOI21_X1   g06966(.A1(\asqrt[32] ), .A2(new_n6728_), .B(new_n6751_), .ZN(new_n7159_));
  OAI21_X1   g06967(.A1(new_n6765_), .A2(new_n6755_), .B(\asqrt[63] ), .ZN(new_n7160_));
  NOR2_X1    g06968(.A1(new_n7159_), .A2(new_n7160_), .ZN(new_n7161_));
  INV_X1     g06969(.I(new_n6778_), .ZN(new_n7162_));
  AND3_X2    g06970(.A1(new_n6727_), .A2(new_n6725_), .A3(new_n6741_), .Z(new_n7163_));
  NAND4_X1   g06971(.A1(new_n7162_), .A2(new_n6766_), .A3(new_n6738_), .A4(new_n7163_), .ZN(new_n7164_));
  INV_X1     g06972(.I(new_n7164_), .ZN(new_n7165_));
  NOR2_X1    g06973(.A1(new_n7161_), .A2(new_n7165_), .ZN(new_n7166_));
  INV_X1     g06974(.I(new_n7166_), .ZN(new_n7167_));
  AOI21_X1   g06975(.A1(new_n7158_), .A2(new_n7156_), .B(new_n7167_), .ZN(new_n7168_));
  NAND2_X1   g06976(.A1(new_n7153_), .A2(new_n7168_), .ZN(\asqrt[31] ));
  NOR2_X1    g06977(.A1(\a[60] ), .A2(\a[61] ), .ZN(new_n7170_));
  INV_X1     g06978(.I(new_n7170_), .ZN(new_n7171_));
  NOR2_X1    g06979(.A1(new_n7171_), .A2(\a[62] ), .ZN(new_n7172_));
  INV_X1     g06980(.I(new_n7172_), .ZN(new_n7173_));
  INV_X1     g06981(.I(new_n7115_), .ZN(new_n7174_));
  NAND2_X1   g06982(.A1(new_n7098_), .A2(new_n306_), .ZN(new_n7175_));
  OAI21_X1   g06983(.A1(new_n7175_), .A2(new_n7131_), .B(new_n7174_), .ZN(new_n7176_));
  AOI21_X1   g06984(.A1(new_n7176_), .A2(new_n7132_), .B(new_n218_), .ZN(new_n7177_));
  NOR3_X1    g06985(.A1(new_n7097_), .A2(\asqrt[59] ), .A3(new_n7088_), .ZN(new_n7178_));
  OAI21_X1   g06986(.A1(new_n7102_), .A2(new_n7178_), .B(new_n7098_), .ZN(new_n7179_));
  AOI21_X1   g06987(.A1(new_n7179_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n7180_));
  AOI21_X1   g06988(.A1(new_n7180_), .A2(new_n7176_), .B(new_n7127_), .ZN(new_n7181_));
  OAI21_X1   g06989(.A1(new_n7181_), .A2(new_n7177_), .B(\asqrt[62] ), .ZN(new_n7182_));
  NOR3_X1    g06990(.A1(new_n7181_), .A2(\asqrt[62] ), .A3(new_n7177_), .ZN(new_n7183_));
  OAI21_X1   g06991(.A1(new_n7139_), .A2(new_n7183_), .B(new_n7182_), .ZN(new_n7184_));
  AOI21_X1   g06992(.A1(new_n7184_), .A2(new_n7151_), .B(\asqrt[63] ), .ZN(new_n7185_));
  NAND2_X1   g06993(.A1(new_n7182_), .A2(new_n7149_), .ZN(new_n7186_));
  OAI21_X1   g06994(.A1(new_n7186_), .A2(new_n7143_), .B(new_n7166_), .ZN(new_n7187_));
  OAI21_X1   g06995(.A1(new_n7185_), .A2(new_n7187_), .B(\a[62] ), .ZN(new_n7188_));
  AOI21_X1   g06996(.A1(new_n7188_), .A2(new_n7173_), .B(new_n6824_), .ZN(new_n7189_));
  INV_X1     g06997(.I(\a[62] ), .ZN(new_n7190_));
  AOI21_X1   g06998(.A1(new_n7153_), .A2(new_n7168_), .B(new_n7190_), .ZN(new_n7191_));
  NAND2_X1   g06999(.A1(new_n6741_), .A2(new_n7173_), .ZN(new_n7192_));
  NOR4_X1    g07000(.A1(new_n6753_), .A2(new_n6778_), .A3(new_n6739_), .A4(new_n7192_), .ZN(new_n7193_));
  INV_X1     g07001(.I(new_n7193_), .ZN(new_n7194_));
  NOR2_X1    g07002(.A1(new_n7191_), .A2(new_n7194_), .ZN(new_n7195_));
  AOI21_X1   g07003(.A1(new_n7153_), .A2(new_n7168_), .B(new_n6748_), .ZN(new_n7196_));
  INV_X1     g07004(.I(\a[63] ), .ZN(new_n7197_));
  AOI21_X1   g07005(.A1(\asqrt[31] ), .A2(new_n7190_), .B(new_n7197_), .ZN(new_n7198_));
  NOR3_X1    g07006(.A1(new_n7195_), .A2(new_n7198_), .A3(new_n7196_), .ZN(new_n7199_));
  OAI21_X1   g07007(.A1(new_n7199_), .A2(new_n7189_), .B(\asqrt[33] ), .ZN(new_n7200_));
  OAI21_X1   g07008(.A1(new_n7185_), .A2(new_n7187_), .B(new_n6747_), .ZN(new_n7201_));
  NAND2_X1   g07009(.A1(new_n7158_), .A2(new_n7156_), .ZN(new_n7202_));
  INV_X1     g07010(.I(new_n7161_), .ZN(new_n7203_));
  NOR2_X1    g07011(.A1(new_n7165_), .A2(new_n6824_), .ZN(new_n7204_));
  NAND4_X1   g07012(.A1(new_n7153_), .A2(new_n7202_), .A3(new_n7203_), .A4(new_n7204_), .ZN(new_n7205_));
  AOI21_X1   g07013(.A1(new_n7205_), .A2(new_n7201_), .B(new_n6760_), .ZN(new_n7206_));
  INV_X1     g07014(.I(new_n7202_), .ZN(new_n7207_));
  NAND2_X1   g07015(.A1(new_n7203_), .A2(new_n7204_), .ZN(new_n7208_));
  NOR3_X1    g07016(.A1(new_n7207_), .A2(new_n7185_), .A3(new_n7208_), .ZN(new_n7209_));
  NOR3_X1    g07017(.A1(new_n7209_), .A2(new_n7196_), .A3(\a[64] ), .ZN(new_n7210_));
  OAI21_X1   g07018(.A1(new_n7191_), .A2(new_n7172_), .B(\asqrt[32] ), .ZN(new_n7211_));
  NAND2_X1   g07019(.A1(new_n7211_), .A2(new_n6356_), .ZN(new_n7212_));
  OAI22_X1   g07020(.A1(new_n7199_), .A2(new_n7212_), .B1(new_n7206_), .B2(new_n7210_), .ZN(new_n7213_));
  AOI21_X1   g07021(.A1(new_n7213_), .A2(new_n7200_), .B(new_n6077_), .ZN(new_n7214_));
  NOR3_X1    g07022(.A1(new_n7029_), .A2(new_n6759_), .A3(new_n6771_), .ZN(new_n7215_));
  NAND3_X1   g07023(.A1(\asqrt[31] ), .A2(new_n6794_), .A3(new_n7014_), .ZN(new_n7216_));
  AOI22_X1   g07024(.A1(new_n7216_), .A2(new_n7029_), .B1(\asqrt[31] ), .B2(new_n7215_), .ZN(new_n7217_));
  AOI21_X1   g07025(.A1(new_n7153_), .A2(new_n7168_), .B(\a[62] ), .ZN(new_n7218_));
  OAI21_X1   g07026(.A1(new_n7197_), .A2(new_n7218_), .B(new_n7201_), .ZN(new_n7219_));
  OAI21_X1   g07027(.A1(new_n7219_), .A2(new_n7195_), .B(new_n7211_), .ZN(new_n7220_));
  AOI21_X1   g07028(.A1(new_n7220_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n7221_));
  AOI21_X1   g07029(.A1(new_n7221_), .A2(new_n7213_), .B(new_n7217_), .ZN(new_n7222_));
  OAI21_X1   g07030(.A1(new_n7222_), .A2(new_n7214_), .B(\asqrt[35] ), .ZN(new_n7223_));
  INV_X1     g07031(.I(new_n7223_), .ZN(new_n7224_));
  NOR2_X1    g07032(.A1(new_n6783_), .A2(new_n6784_), .ZN(new_n7225_));
  NOR2_X1    g07033(.A1(new_n6775_), .A2(new_n6786_), .ZN(new_n7226_));
  INV_X1     g07034(.I(new_n7226_), .ZN(new_n7227_));
  NAND4_X1   g07035(.A1(\asqrt[31] ), .A2(new_n6776_), .A3(new_n7225_), .A4(new_n7227_), .ZN(new_n7228_));
  INV_X1     g07036(.I(\asqrt[31] ), .ZN(new_n7229_));
  NOR3_X1    g07037(.A1(new_n7229_), .A2(new_n7018_), .A3(new_n7226_), .ZN(new_n7230_));
  OAI21_X1   g07038(.A1(new_n7230_), .A2(new_n7225_), .B(new_n7228_), .ZN(new_n7231_));
  INV_X1     g07039(.I(new_n7231_), .ZN(new_n7232_));
  NOR3_X1    g07040(.A1(new_n7222_), .A2(new_n7214_), .A3(\asqrt[35] ), .ZN(new_n7233_));
  NOR2_X1    g07041(.A1(new_n7233_), .A2(new_n7232_), .ZN(new_n7234_));
  OAI21_X1   g07042(.A1(new_n7234_), .A2(new_n7224_), .B(\asqrt[36] ), .ZN(new_n7235_));
  NOR2_X1    g07043(.A1(new_n7031_), .A2(new_n7023_), .ZN(new_n7236_));
  NOR3_X1    g07044(.A1(new_n7229_), .A2(new_n6788_), .A3(new_n7236_), .ZN(new_n7237_));
  INV_X1     g07045(.I(new_n7237_), .ZN(new_n7238_));
  NOR3_X1    g07046(.A1(new_n7236_), .A2(new_n6788_), .A3(new_n7028_), .ZN(new_n7239_));
  AOI22_X1   g07047(.A1(new_n7238_), .A2(new_n7028_), .B1(\asqrt[31] ), .B2(new_n7239_), .ZN(new_n7240_));
  INV_X1     g07048(.I(new_n7240_), .ZN(new_n7241_));
  NAND2_X1   g07049(.A1(new_n7223_), .A2(new_n5277_), .ZN(new_n7242_));
  OAI21_X1   g07050(.A1(new_n7234_), .A2(new_n7242_), .B(new_n7241_), .ZN(new_n7243_));
  AOI21_X1   g07051(.A1(new_n7243_), .A2(new_n7235_), .B(new_n5024_), .ZN(new_n7244_));
  NOR3_X1    g07052(.A1(new_n6801_), .A2(new_n6809_), .A3(new_n6807_), .ZN(new_n7245_));
  NOR3_X1    g07053(.A1(new_n7229_), .A2(new_n6801_), .A3(new_n6809_), .ZN(new_n7246_));
  INV_X1     g07054(.I(new_n7246_), .ZN(new_n7247_));
  AOI22_X1   g07055(.A1(new_n7247_), .A2(new_n6807_), .B1(\asqrt[31] ), .B2(new_n7245_), .ZN(new_n7248_));
  OAI21_X1   g07056(.A1(new_n7232_), .A2(new_n7233_), .B(new_n7223_), .ZN(new_n7249_));
  AOI21_X1   g07057(.A1(new_n7249_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n7250_));
  AOI21_X1   g07058(.A1(new_n7250_), .A2(new_n7243_), .B(new_n7248_), .ZN(new_n7251_));
  OAI21_X1   g07059(.A1(new_n7251_), .A2(new_n7244_), .B(\asqrt[38] ), .ZN(new_n7252_));
  INV_X1     g07060(.I(new_n7252_), .ZN(new_n7253_));
  NAND2_X1   g07061(.A1(new_n7034_), .A2(new_n7026_), .ZN(new_n7254_));
  NAND3_X1   g07062(.A1(\asqrt[31] ), .A2(new_n6811_), .A3(new_n7254_), .ZN(new_n7255_));
  AND3_X2    g07063(.A1(new_n6811_), .A2(new_n6817_), .A3(new_n7254_), .Z(new_n7256_));
  AOI22_X1   g07064(.A1(new_n7255_), .A2(new_n6818_), .B1(\asqrt[31] ), .B2(new_n7256_), .ZN(new_n7257_));
  NOR3_X1    g07065(.A1(new_n7251_), .A2(new_n7244_), .A3(\asqrt[38] ), .ZN(new_n7258_));
  NOR2_X1    g07066(.A1(new_n7258_), .A2(new_n7257_), .ZN(new_n7259_));
  OAI21_X1   g07067(.A1(new_n7259_), .A2(new_n7253_), .B(\asqrt[39] ), .ZN(new_n7260_));
  INV_X1     g07068(.I(new_n6827_), .ZN(new_n7261_));
  NOR3_X1    g07069(.A1(new_n6821_), .A2(new_n7045_), .A3(new_n7261_), .ZN(new_n7262_));
  NOR3_X1    g07070(.A1(new_n7229_), .A2(new_n6821_), .A3(new_n7045_), .ZN(new_n7263_));
  INV_X1     g07071(.I(new_n7263_), .ZN(new_n7264_));
  AOI22_X1   g07072(.A1(new_n7264_), .A2(new_n7261_), .B1(\asqrt[31] ), .B2(new_n7262_), .ZN(new_n7265_));
  INV_X1     g07073(.I(new_n7265_), .ZN(new_n7266_));
  NAND2_X1   g07074(.A1(new_n7252_), .A2(new_n4298_), .ZN(new_n7267_));
  OAI21_X1   g07075(.A1(new_n7259_), .A2(new_n7267_), .B(new_n7266_), .ZN(new_n7268_));
  AOI21_X1   g07076(.A1(new_n7268_), .A2(new_n7260_), .B(new_n4071_), .ZN(new_n7269_));
  NOR3_X1    g07077(.A1(new_n7229_), .A2(new_n6832_), .A3(new_n6839_), .ZN(new_n7270_));
  INV_X1     g07078(.I(new_n7270_), .ZN(new_n7271_));
  NOR3_X1    g07079(.A1(new_n6832_), .A2(new_n7013_), .A3(new_n6839_), .ZN(new_n7272_));
  AOI22_X1   g07080(.A1(new_n7271_), .A2(new_n7013_), .B1(\asqrt[31] ), .B2(new_n7272_), .ZN(new_n7273_));
  INV_X1     g07081(.I(new_n7257_), .ZN(new_n7274_));
  NAND2_X1   g07082(.A1(new_n7188_), .A2(new_n7193_), .ZN(new_n7275_));
  OAI21_X1   g07083(.A1(new_n7185_), .A2(new_n7187_), .B(new_n7190_), .ZN(new_n7276_));
  NAND2_X1   g07084(.A1(new_n7276_), .A2(\a[63] ), .ZN(new_n7277_));
  NAND3_X1   g07085(.A1(new_n7275_), .A2(new_n7277_), .A3(new_n7201_), .ZN(new_n7278_));
  AOI21_X1   g07086(.A1(new_n7278_), .A2(new_n7211_), .B(new_n6356_), .ZN(new_n7279_));
  OAI21_X1   g07087(.A1(new_n7209_), .A2(new_n7196_), .B(\a[64] ), .ZN(new_n7280_));
  NAND3_X1   g07088(.A1(new_n7205_), .A2(new_n7201_), .A3(new_n6760_), .ZN(new_n7281_));
  NAND2_X1   g07089(.A1(new_n7188_), .A2(new_n7173_), .ZN(new_n7282_));
  AOI21_X1   g07090(.A1(new_n7282_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n7283_));
  AOI22_X1   g07091(.A1(new_n7278_), .A2(new_n7283_), .B1(new_n7280_), .B2(new_n7281_), .ZN(new_n7284_));
  OAI21_X1   g07092(.A1(new_n7284_), .A2(new_n7279_), .B(\asqrt[34] ), .ZN(new_n7285_));
  NAND2_X1   g07093(.A1(new_n7285_), .A2(new_n5708_), .ZN(new_n7286_));
  OAI21_X1   g07094(.A1(new_n7286_), .A2(new_n7222_), .B(new_n7231_), .ZN(new_n7287_));
  AOI21_X1   g07095(.A1(new_n7287_), .A2(new_n7223_), .B(new_n5277_), .ZN(new_n7288_));
  INV_X1     g07096(.I(new_n7217_), .ZN(new_n7289_));
  AOI21_X1   g07097(.A1(\a[63] ), .A2(new_n7276_), .B(new_n7196_), .ZN(new_n7290_));
  AOI21_X1   g07098(.A1(new_n7290_), .A2(new_n7275_), .B(new_n7189_), .ZN(new_n7291_));
  OAI21_X1   g07099(.A1(new_n7291_), .A2(new_n6356_), .B(new_n6077_), .ZN(new_n7292_));
  OAI21_X1   g07100(.A1(new_n7292_), .A2(new_n7284_), .B(new_n7289_), .ZN(new_n7293_));
  NAND2_X1   g07101(.A1(new_n7293_), .A2(new_n7285_), .ZN(new_n7294_));
  AOI21_X1   g07102(.A1(new_n7294_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n7295_));
  AOI21_X1   g07103(.A1(new_n7295_), .A2(new_n7287_), .B(new_n7240_), .ZN(new_n7296_));
  OAI21_X1   g07104(.A1(new_n7296_), .A2(new_n7288_), .B(\asqrt[37] ), .ZN(new_n7297_));
  NAND2_X1   g07105(.A1(new_n7297_), .A2(new_n4696_), .ZN(new_n7298_));
  OAI21_X1   g07106(.A1(new_n7298_), .A2(new_n7251_), .B(new_n7274_), .ZN(new_n7299_));
  AOI21_X1   g07107(.A1(new_n7299_), .A2(new_n7252_), .B(new_n4298_), .ZN(new_n7300_));
  NOR2_X1    g07108(.A1(new_n7300_), .A2(\asqrt[40] ), .ZN(new_n7301_));
  AOI21_X1   g07109(.A1(new_n7301_), .A2(new_n7268_), .B(new_n7273_), .ZN(new_n7302_));
  OAI21_X1   g07110(.A1(new_n7302_), .A2(new_n7269_), .B(\asqrt[41] ), .ZN(new_n7303_));
  INV_X1     g07111(.I(new_n7039_), .ZN(new_n7304_));
  NOR3_X1    g07112(.A1(new_n7304_), .A2(new_n7044_), .A3(new_n6850_), .ZN(new_n7305_));
  NOR3_X1    g07113(.A1(new_n7229_), .A2(new_n7044_), .A3(new_n7304_), .ZN(new_n7306_));
  INV_X1     g07114(.I(new_n7306_), .ZN(new_n7307_));
  AOI22_X1   g07115(.A1(new_n7307_), .A2(new_n6850_), .B1(\asqrt[31] ), .B2(new_n7305_), .ZN(new_n7308_));
  INV_X1     g07116(.I(new_n7308_), .ZN(new_n7309_));
  OAI21_X1   g07117(.A1(new_n7257_), .A2(new_n7258_), .B(new_n7252_), .ZN(new_n7310_));
  NAND3_X1   g07118(.A1(new_n7299_), .A2(new_n4298_), .A3(new_n7252_), .ZN(new_n7311_));
  AOI22_X1   g07119(.A1(new_n7311_), .A2(new_n7266_), .B1(new_n7310_), .B2(\asqrt[39] ), .ZN(new_n7312_));
  OAI21_X1   g07120(.A1(new_n7312_), .A2(new_n4071_), .B(new_n3782_), .ZN(new_n7313_));
  OAI21_X1   g07121(.A1(new_n7313_), .A2(new_n7302_), .B(new_n7309_), .ZN(new_n7314_));
  AOI21_X1   g07122(.A1(new_n7314_), .A2(new_n7303_), .B(new_n3419_), .ZN(new_n7315_));
  INV_X1     g07123(.I(new_n6858_), .ZN(new_n7316_));
  NOR3_X1    g07124(.A1(new_n7229_), .A2(new_n6853_), .A3(new_n7049_), .ZN(new_n7317_));
  INV_X1     g07125(.I(new_n7317_), .ZN(new_n7318_));
  NOR3_X1    g07126(.A1(new_n6853_), .A2(new_n7049_), .A3(new_n7316_), .ZN(new_n7319_));
  AOI22_X1   g07127(.A1(new_n7318_), .A2(new_n7316_), .B1(\asqrt[31] ), .B2(new_n7319_), .ZN(new_n7320_));
  NOR3_X1    g07128(.A1(new_n7296_), .A2(new_n7288_), .A3(\asqrt[37] ), .ZN(new_n7321_));
  OAI21_X1   g07129(.A1(new_n7248_), .A2(new_n7321_), .B(new_n7297_), .ZN(new_n7322_));
  AOI21_X1   g07130(.A1(new_n7322_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n7323_));
  AOI21_X1   g07131(.A1(new_n7323_), .A2(new_n7299_), .B(new_n7265_), .ZN(new_n7324_));
  NOR3_X1    g07132(.A1(new_n7324_), .A2(\asqrt[40] ), .A3(new_n7300_), .ZN(new_n7325_));
  OAI22_X1   g07133(.A1(new_n7325_), .A2(new_n7273_), .B1(new_n7312_), .B2(new_n4071_), .ZN(new_n7326_));
  AOI21_X1   g07134(.A1(new_n7326_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n7327_));
  AOI21_X1   g07135(.A1(new_n7327_), .A2(new_n7314_), .B(new_n7320_), .ZN(new_n7328_));
  OAI21_X1   g07136(.A1(new_n7328_), .A2(new_n7315_), .B(\asqrt[43] ), .ZN(new_n7329_));
  INV_X1     g07137(.I(new_n7329_), .ZN(new_n7330_));
  NOR3_X1    g07138(.A1(new_n6863_), .A2(new_n7012_), .A3(new_n6869_), .ZN(new_n7331_));
  NOR3_X1    g07139(.A1(new_n7229_), .A2(new_n6863_), .A3(new_n6869_), .ZN(new_n7332_));
  INV_X1     g07140(.I(new_n7332_), .ZN(new_n7333_));
  AOI22_X1   g07141(.A1(new_n7333_), .A2(new_n7012_), .B1(\asqrt[31] ), .B2(new_n7331_), .ZN(new_n7334_));
  NOR3_X1    g07142(.A1(new_n7328_), .A2(\asqrt[43] ), .A3(new_n7315_), .ZN(new_n7335_));
  NOR2_X1    g07143(.A1(new_n7335_), .A2(new_n7334_), .ZN(new_n7336_));
  OAI21_X1   g07144(.A1(new_n7336_), .A2(new_n7330_), .B(\asqrt[44] ), .ZN(new_n7337_));
  NOR2_X1    g07145(.A1(new_n6870_), .A2(new_n6881_), .ZN(new_n7338_));
  NOR3_X1    g07146(.A1(new_n7229_), .A2(new_n7043_), .A3(new_n7338_), .ZN(new_n7339_));
  INV_X1     g07147(.I(new_n7339_), .ZN(new_n7340_));
  NOR3_X1    g07148(.A1(new_n7338_), .A2(new_n7043_), .A3(new_n6880_), .ZN(new_n7341_));
  AOI22_X1   g07149(.A1(new_n7340_), .A2(new_n6880_), .B1(\asqrt[31] ), .B2(new_n7341_), .ZN(new_n7342_));
  INV_X1     g07150(.I(new_n7342_), .ZN(new_n7343_));
  NAND2_X1   g07151(.A1(new_n7329_), .A2(new_n2954_), .ZN(new_n7344_));
  OAI21_X1   g07152(.A1(new_n7336_), .A2(new_n7344_), .B(new_n7343_), .ZN(new_n7345_));
  AOI21_X1   g07153(.A1(new_n7345_), .A2(new_n7337_), .B(new_n2641_), .ZN(new_n7346_));
  INV_X1     g07154(.I(new_n6888_), .ZN(new_n7347_));
  NOR3_X1    g07155(.A1(new_n6883_), .A2(new_n7057_), .A3(new_n7347_), .ZN(new_n7348_));
  NOR3_X1    g07156(.A1(new_n7229_), .A2(new_n6883_), .A3(new_n7057_), .ZN(new_n7349_));
  INV_X1     g07157(.I(new_n7349_), .ZN(new_n7350_));
  AOI22_X1   g07158(.A1(new_n7350_), .A2(new_n7347_), .B1(\asqrt[31] ), .B2(new_n7348_), .ZN(new_n7351_));
  OAI21_X1   g07159(.A1(new_n7334_), .A2(new_n7335_), .B(new_n7329_), .ZN(new_n7352_));
  AOI21_X1   g07160(.A1(new_n7352_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n7353_));
  AOI21_X1   g07161(.A1(new_n7353_), .A2(new_n7345_), .B(new_n7351_), .ZN(new_n7354_));
  OAI21_X1   g07162(.A1(new_n7354_), .A2(new_n7346_), .B(\asqrt[46] ), .ZN(new_n7355_));
  INV_X1     g07163(.I(new_n7355_), .ZN(new_n7356_));
  NOR3_X1    g07164(.A1(new_n7229_), .A2(new_n6893_), .A3(new_n6900_), .ZN(new_n7357_));
  INV_X1     g07165(.I(new_n7357_), .ZN(new_n7358_));
  NOR3_X1    g07166(.A1(new_n6893_), .A2(new_n7011_), .A3(new_n6900_), .ZN(new_n7359_));
  AOI22_X1   g07167(.A1(new_n7358_), .A2(new_n7011_), .B1(\asqrt[31] ), .B2(new_n7359_), .ZN(new_n7360_));
  NOR3_X1    g07168(.A1(new_n7354_), .A2(new_n7346_), .A3(\asqrt[46] ), .ZN(new_n7361_));
  NOR2_X1    g07169(.A1(new_n7361_), .A2(new_n7360_), .ZN(new_n7362_));
  OAI21_X1   g07170(.A1(new_n7362_), .A2(new_n7356_), .B(\asqrt[47] ), .ZN(new_n7363_));
  NOR2_X1    g07171(.A1(new_n6901_), .A2(new_n6912_), .ZN(new_n7364_));
  NOR3_X1    g07172(.A1(new_n7364_), .A2(new_n7056_), .A3(new_n6911_), .ZN(new_n7365_));
  NOR3_X1    g07173(.A1(new_n7229_), .A2(new_n7056_), .A3(new_n7364_), .ZN(new_n7366_));
  INV_X1     g07174(.I(new_n7366_), .ZN(new_n7367_));
  AOI22_X1   g07175(.A1(new_n7367_), .A2(new_n6911_), .B1(\asqrt[31] ), .B2(new_n7365_), .ZN(new_n7368_));
  INV_X1     g07176(.I(new_n7368_), .ZN(new_n7369_));
  NAND2_X1   g07177(.A1(new_n7355_), .A2(new_n2229_), .ZN(new_n7370_));
  OAI21_X1   g07178(.A1(new_n7362_), .A2(new_n7370_), .B(new_n7369_), .ZN(new_n7371_));
  AOI21_X1   g07179(.A1(new_n7371_), .A2(new_n7363_), .B(new_n1956_), .ZN(new_n7372_));
  INV_X1     g07180(.I(new_n6919_), .ZN(new_n7373_));
  NOR3_X1    g07181(.A1(new_n7229_), .A2(new_n6914_), .A3(new_n7065_), .ZN(new_n7374_));
  INV_X1     g07182(.I(new_n7374_), .ZN(new_n7375_));
  NOR3_X1    g07183(.A1(new_n6914_), .A2(new_n7065_), .A3(new_n7373_), .ZN(new_n7376_));
  AOI22_X1   g07184(.A1(new_n7375_), .A2(new_n7373_), .B1(\asqrt[31] ), .B2(new_n7376_), .ZN(new_n7377_));
  OAI21_X1   g07185(.A1(new_n7360_), .A2(new_n7361_), .B(new_n7355_), .ZN(new_n7378_));
  AOI21_X1   g07186(.A1(new_n7378_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n7379_));
  AOI21_X1   g07187(.A1(new_n7379_), .A2(new_n7371_), .B(new_n7377_), .ZN(new_n7380_));
  OAI21_X1   g07188(.A1(new_n7380_), .A2(new_n7372_), .B(\asqrt[49] ), .ZN(new_n7381_));
  INV_X1     g07189(.I(new_n7381_), .ZN(new_n7382_));
  NOR3_X1    g07190(.A1(new_n6924_), .A2(new_n7010_), .A3(new_n6930_), .ZN(new_n7383_));
  NOR3_X1    g07191(.A1(new_n7229_), .A2(new_n6924_), .A3(new_n6930_), .ZN(new_n7384_));
  INV_X1     g07192(.I(new_n7384_), .ZN(new_n7385_));
  AOI22_X1   g07193(.A1(new_n7385_), .A2(new_n7010_), .B1(\asqrt[31] ), .B2(new_n7383_), .ZN(new_n7386_));
  NOR3_X1    g07194(.A1(new_n7380_), .A2(new_n7372_), .A3(\asqrt[49] ), .ZN(new_n7387_));
  NOR2_X1    g07195(.A1(new_n7387_), .A2(new_n7386_), .ZN(new_n7388_));
  OAI21_X1   g07196(.A1(new_n7388_), .A2(new_n7382_), .B(\asqrt[50] ), .ZN(new_n7389_));
  NOR2_X1    g07197(.A1(new_n6931_), .A2(new_n6939_), .ZN(new_n7390_));
  NOR3_X1    g07198(.A1(new_n7229_), .A2(new_n7064_), .A3(new_n7390_), .ZN(new_n7391_));
  INV_X1     g07199(.I(new_n7391_), .ZN(new_n7392_));
  NOR3_X1    g07200(.A1(new_n7390_), .A2(new_n7064_), .A3(new_n6938_), .ZN(new_n7393_));
  AOI22_X1   g07201(.A1(new_n7392_), .A2(new_n6938_), .B1(\asqrt[31] ), .B2(new_n7393_), .ZN(new_n7394_));
  INV_X1     g07202(.I(new_n7394_), .ZN(new_n7395_));
  NAND2_X1   g07203(.A1(new_n7381_), .A2(new_n1612_), .ZN(new_n7396_));
  OAI21_X1   g07204(.A1(new_n7388_), .A2(new_n7396_), .B(new_n7395_), .ZN(new_n7397_));
  AOI21_X1   g07205(.A1(new_n7397_), .A2(new_n7389_), .B(new_n1376_), .ZN(new_n7398_));
  INV_X1     g07206(.I(new_n6945_), .ZN(new_n7399_));
  NOR3_X1    g07207(.A1(new_n6941_), .A2(new_n7073_), .A3(new_n7399_), .ZN(new_n7400_));
  NOR3_X1    g07208(.A1(new_n7229_), .A2(new_n6941_), .A3(new_n7073_), .ZN(new_n7401_));
  INV_X1     g07209(.I(new_n7401_), .ZN(new_n7402_));
  AOI22_X1   g07210(.A1(new_n7402_), .A2(new_n7399_), .B1(\asqrt[31] ), .B2(new_n7400_), .ZN(new_n7403_));
  OAI21_X1   g07211(.A1(new_n7386_), .A2(new_n7387_), .B(new_n7381_), .ZN(new_n7404_));
  AOI21_X1   g07212(.A1(new_n7404_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n7405_));
  AOI21_X1   g07213(.A1(new_n7405_), .A2(new_n7397_), .B(new_n7403_), .ZN(new_n7406_));
  OAI21_X1   g07214(.A1(new_n7406_), .A2(new_n7398_), .B(\asqrt[52] ), .ZN(new_n7407_));
  INV_X1     g07215(.I(new_n7407_), .ZN(new_n7408_));
  INV_X1     g07216(.I(new_n7406_), .ZN(new_n7409_));
  NOR3_X1    g07217(.A1(new_n7229_), .A2(new_n6950_), .A3(new_n6956_), .ZN(new_n7410_));
  INV_X1     g07218(.I(new_n7410_), .ZN(new_n7411_));
  NOR3_X1    g07219(.A1(new_n6950_), .A2(new_n7009_), .A3(new_n6956_), .ZN(new_n7412_));
  AOI22_X1   g07220(.A1(new_n7411_), .A2(new_n7009_), .B1(\asqrt[31] ), .B2(new_n7412_), .ZN(new_n7413_));
  NOR2_X1    g07221(.A1(new_n7398_), .A2(\asqrt[52] ), .ZN(new_n7414_));
  AOI21_X1   g07222(.A1(new_n7409_), .A2(new_n7414_), .B(new_n7413_), .ZN(new_n7415_));
  OAI21_X1   g07223(.A1(new_n7415_), .A2(new_n7408_), .B(\asqrt[53] ), .ZN(new_n7416_));
  NOR2_X1    g07224(.A1(new_n6957_), .A2(new_n6965_), .ZN(new_n7417_));
  NOR3_X1    g07225(.A1(new_n7417_), .A2(new_n7072_), .A3(new_n6964_), .ZN(new_n7418_));
  NOR3_X1    g07226(.A1(new_n7229_), .A2(new_n7072_), .A3(new_n7417_), .ZN(new_n7419_));
  INV_X1     g07227(.I(new_n7419_), .ZN(new_n7420_));
  AOI22_X1   g07228(.A1(new_n7420_), .A2(new_n6964_), .B1(\asqrt[31] ), .B2(new_n7418_), .ZN(new_n7421_));
  INV_X1     g07229(.I(new_n7421_), .ZN(new_n7422_));
  NAND2_X1   g07230(.A1(new_n7407_), .A2(new_n1103_), .ZN(new_n7423_));
  OAI21_X1   g07231(.A1(new_n7423_), .A2(new_n7415_), .B(new_n7422_), .ZN(new_n7424_));
  AOI21_X1   g07232(.A1(new_n7424_), .A2(new_n7416_), .B(new_n904_), .ZN(new_n7425_));
  INV_X1     g07233(.I(new_n7425_), .ZN(new_n7426_));
  INV_X1     g07234(.I(new_n7424_), .ZN(new_n7427_));
  INV_X1     g07235(.I(new_n6971_), .ZN(new_n7428_));
  NOR3_X1    g07236(.A1(new_n7229_), .A2(new_n6967_), .A3(new_n7081_), .ZN(new_n7429_));
  INV_X1     g07237(.I(new_n7429_), .ZN(new_n7430_));
  NOR3_X1    g07238(.A1(new_n6967_), .A2(new_n7081_), .A3(new_n7428_), .ZN(new_n7431_));
  AOI22_X1   g07239(.A1(new_n7430_), .A2(new_n7428_), .B1(\asqrt[31] ), .B2(new_n7431_), .ZN(new_n7432_));
  INV_X1     g07240(.I(new_n7432_), .ZN(new_n7433_));
  NAND2_X1   g07241(.A1(new_n7416_), .A2(new_n904_), .ZN(new_n7434_));
  OAI21_X1   g07242(.A1(new_n7434_), .A2(new_n7427_), .B(new_n7433_), .ZN(new_n7435_));
  AOI21_X1   g07243(.A1(new_n7435_), .A2(new_n7426_), .B(new_n823_), .ZN(new_n7436_));
  NOR3_X1    g07244(.A1(new_n6976_), .A2(new_n6982_), .A3(new_n7008_), .ZN(new_n7437_));
  NOR3_X1    g07245(.A1(new_n7229_), .A2(new_n6976_), .A3(new_n6982_), .ZN(new_n7438_));
  INV_X1     g07246(.I(new_n7438_), .ZN(new_n7439_));
  AOI22_X1   g07247(.A1(new_n7439_), .A2(new_n7008_), .B1(\asqrt[31] ), .B2(new_n7437_), .ZN(new_n7440_));
  NOR2_X1    g07248(.A1(new_n7425_), .A2(\asqrt[55] ), .ZN(new_n7441_));
  AOI21_X1   g07249(.A1(new_n7441_), .A2(new_n7435_), .B(new_n7440_), .ZN(new_n7442_));
  OAI21_X1   g07250(.A1(new_n7442_), .A2(new_n7436_), .B(\asqrt[56] ), .ZN(new_n7443_));
  NOR2_X1    g07251(.A1(new_n6983_), .A2(new_n6991_), .ZN(new_n7444_));
  NOR3_X1    g07252(.A1(new_n7229_), .A2(new_n7080_), .A3(new_n7444_), .ZN(new_n7445_));
  INV_X1     g07253(.I(new_n7445_), .ZN(new_n7446_));
  NOR3_X1    g07254(.A1(new_n7444_), .A2(new_n7080_), .A3(new_n6990_), .ZN(new_n7447_));
  AOI22_X1   g07255(.A1(new_n7446_), .A2(new_n6990_), .B1(\asqrt[31] ), .B2(new_n7447_), .ZN(new_n7448_));
  INV_X1     g07256(.I(new_n7448_), .ZN(new_n7449_));
  NOR3_X1    g07257(.A1(new_n7406_), .A2(new_n7398_), .A3(\asqrt[52] ), .ZN(new_n7450_));
  OAI21_X1   g07258(.A1(new_n7413_), .A2(new_n7450_), .B(new_n7407_), .ZN(new_n7451_));
  AOI21_X1   g07259(.A1(new_n7451_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n7452_));
  AOI21_X1   g07260(.A1(new_n7452_), .A2(new_n7424_), .B(new_n7432_), .ZN(new_n7453_));
  OAI21_X1   g07261(.A1(new_n7453_), .A2(new_n7425_), .B(\asqrt[55] ), .ZN(new_n7454_));
  NAND2_X1   g07262(.A1(new_n7454_), .A2(new_n703_), .ZN(new_n7455_));
  OAI21_X1   g07263(.A1(new_n7455_), .A2(new_n7442_), .B(new_n7449_), .ZN(new_n7456_));
  AOI21_X1   g07264(.A1(new_n7456_), .A2(new_n7443_), .B(new_n531_), .ZN(new_n7457_));
  INV_X1     g07265(.I(new_n7457_), .ZN(new_n7458_));
  INV_X1     g07266(.I(new_n7456_), .ZN(new_n7459_));
  INV_X1     g07267(.I(new_n6997_), .ZN(new_n7460_));
  NOR3_X1    g07268(.A1(new_n6993_), .A2(new_n7094_), .A3(new_n7460_), .ZN(new_n7461_));
  NOR3_X1    g07269(.A1(new_n7229_), .A2(new_n6993_), .A3(new_n7094_), .ZN(new_n7462_));
  INV_X1     g07270(.I(new_n7462_), .ZN(new_n7463_));
  AOI22_X1   g07271(.A1(new_n7463_), .A2(new_n7460_), .B1(\asqrt[31] ), .B2(new_n7461_), .ZN(new_n7464_));
  INV_X1     g07272(.I(new_n7464_), .ZN(new_n7465_));
  NAND2_X1   g07273(.A1(new_n7443_), .A2(new_n531_), .ZN(new_n7466_));
  OAI21_X1   g07274(.A1(new_n7466_), .A2(new_n7459_), .B(new_n7465_), .ZN(new_n7467_));
  AOI21_X1   g07275(.A1(new_n7467_), .A2(new_n7458_), .B(new_n436_), .ZN(new_n7468_));
  NOR3_X1    g07276(.A1(new_n7229_), .A2(new_n7104_), .A3(new_n7105_), .ZN(new_n7469_));
  INV_X1     g07277(.I(new_n7469_), .ZN(new_n7470_));
  NOR3_X1    g07278(.A1(new_n7104_), .A2(new_n7105_), .A3(new_n7007_), .ZN(new_n7471_));
  AOI22_X1   g07279(.A1(new_n7470_), .A2(new_n7007_), .B1(\asqrt[31] ), .B2(new_n7471_), .ZN(new_n7472_));
  NOR2_X1    g07280(.A1(new_n7457_), .A2(\asqrt[58] ), .ZN(new_n7473_));
  AOI21_X1   g07281(.A1(new_n7473_), .A2(new_n7467_), .B(new_n7472_), .ZN(new_n7474_));
  OAI21_X1   g07282(.A1(new_n7474_), .A2(new_n7468_), .B(\asqrt[59] ), .ZN(new_n7475_));
  NOR2_X1    g07283(.A1(new_n7106_), .A2(new_n7117_), .ZN(new_n7476_));
  NOR3_X1    g07284(.A1(new_n7476_), .A2(new_n7088_), .A3(new_n7116_), .ZN(new_n7477_));
  NOR3_X1    g07285(.A1(new_n7229_), .A2(new_n7088_), .A3(new_n7476_), .ZN(new_n7478_));
  INV_X1     g07286(.I(new_n7478_), .ZN(new_n7479_));
  AOI22_X1   g07287(.A1(new_n7479_), .A2(new_n7116_), .B1(\asqrt[31] ), .B2(new_n7477_), .ZN(new_n7480_));
  INV_X1     g07288(.I(new_n7480_), .ZN(new_n7481_));
  NOR3_X1    g07289(.A1(new_n7453_), .A2(\asqrt[55] ), .A3(new_n7425_), .ZN(new_n7482_));
  OAI21_X1   g07290(.A1(new_n7440_), .A2(new_n7482_), .B(new_n7454_), .ZN(new_n7483_));
  AOI21_X1   g07291(.A1(new_n7483_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n7484_));
  AOI21_X1   g07292(.A1(new_n7484_), .A2(new_n7456_), .B(new_n7464_), .ZN(new_n7485_));
  OAI21_X1   g07293(.A1(new_n7485_), .A2(new_n7457_), .B(\asqrt[58] ), .ZN(new_n7486_));
  NAND2_X1   g07294(.A1(new_n7486_), .A2(new_n327_), .ZN(new_n7487_));
  OAI21_X1   g07295(.A1(new_n7487_), .A2(new_n7474_), .B(new_n7481_), .ZN(new_n7488_));
  AOI21_X1   g07296(.A1(new_n7488_), .A2(new_n7475_), .B(new_n306_), .ZN(new_n7489_));
  INV_X1     g07297(.I(new_n7489_), .ZN(new_n7490_));
  INV_X1     g07298(.I(new_n7488_), .ZN(new_n7491_));
  NOR3_X1    g07299(.A1(new_n7229_), .A2(new_n7119_), .A3(new_n7178_), .ZN(new_n7492_));
  INV_X1     g07300(.I(new_n7492_), .ZN(new_n7493_));
  NOR3_X1    g07301(.A1(new_n7119_), .A2(new_n7178_), .A3(new_n7103_), .ZN(new_n7494_));
  AOI22_X1   g07302(.A1(new_n7493_), .A2(new_n7103_), .B1(\asqrt[31] ), .B2(new_n7494_), .ZN(new_n7495_));
  INV_X1     g07303(.I(new_n7495_), .ZN(new_n7496_));
  NAND2_X1   g07304(.A1(new_n7475_), .A2(new_n306_), .ZN(new_n7497_));
  OAI21_X1   g07305(.A1(new_n7491_), .A2(new_n7497_), .B(new_n7496_), .ZN(new_n7498_));
  AOI21_X1   g07306(.A1(new_n7498_), .A2(new_n7490_), .B(new_n218_), .ZN(new_n7499_));
  NOR3_X1    g07307(.A1(new_n7110_), .A2(new_n7140_), .A3(new_n7174_), .ZN(new_n7500_));
  NOR3_X1    g07308(.A1(new_n7229_), .A2(new_n7110_), .A3(new_n7140_), .ZN(new_n7501_));
  INV_X1     g07309(.I(new_n7501_), .ZN(new_n7502_));
  AOI22_X1   g07310(.A1(new_n7502_), .A2(new_n7174_), .B1(\asqrt[31] ), .B2(new_n7500_), .ZN(new_n7503_));
  NOR2_X1    g07311(.A1(new_n7489_), .A2(\asqrt[61] ), .ZN(new_n7504_));
  AOI21_X1   g07312(.A1(new_n7504_), .A2(new_n7498_), .B(new_n7503_), .ZN(new_n7505_));
  OAI21_X1   g07313(.A1(new_n7505_), .A2(new_n7499_), .B(\asqrt[62] ), .ZN(new_n7506_));
  NOR2_X1    g07314(.A1(new_n7133_), .A2(new_n7121_), .ZN(new_n7507_));
  NOR3_X1    g07315(.A1(new_n7229_), .A2(new_n7177_), .A3(new_n7507_), .ZN(new_n7508_));
  INV_X1     g07316(.I(new_n7508_), .ZN(new_n7509_));
  NOR3_X1    g07317(.A1(new_n7507_), .A2(new_n7177_), .A3(new_n7128_), .ZN(new_n7510_));
  AOI22_X1   g07318(.A1(new_n7509_), .A2(new_n7128_), .B1(\asqrt[31] ), .B2(new_n7510_), .ZN(new_n7511_));
  INV_X1     g07319(.I(new_n7511_), .ZN(new_n7512_));
  NOR3_X1    g07320(.A1(new_n7485_), .A2(\asqrt[58] ), .A3(new_n7457_), .ZN(new_n7513_));
  OAI21_X1   g07321(.A1(new_n7472_), .A2(new_n7513_), .B(new_n7486_), .ZN(new_n7514_));
  AOI21_X1   g07322(.A1(new_n7514_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n7515_));
  AOI21_X1   g07323(.A1(new_n7515_), .A2(new_n7488_), .B(new_n7495_), .ZN(new_n7516_));
  OAI21_X1   g07324(.A1(new_n7516_), .A2(new_n7489_), .B(\asqrt[61] ), .ZN(new_n7517_));
  NAND2_X1   g07325(.A1(new_n7517_), .A2(new_n207_), .ZN(new_n7518_));
  OAI21_X1   g07326(.A1(new_n7518_), .A2(new_n7505_), .B(new_n7512_), .ZN(new_n7519_));
  NAND4_X1   g07327(.A1(\asqrt[31] ), .A2(new_n7182_), .A3(new_n7139_), .A4(new_n7155_), .ZN(new_n7520_));
  NAND2_X1   g07328(.A1(new_n7182_), .A2(new_n7155_), .ZN(new_n7521_));
  OAI21_X1   g07329(.A1(new_n7229_), .A2(new_n7521_), .B(new_n7154_), .ZN(new_n7522_));
  NAND2_X1   g07330(.A1(new_n7522_), .A2(new_n7520_), .ZN(new_n7523_));
  AOI21_X1   g07331(.A1(new_n7156_), .A2(new_n7182_), .B(new_n7149_), .ZN(new_n7524_));
  AOI21_X1   g07332(.A1(\asqrt[31] ), .A2(new_n7524_), .B(new_n7207_), .ZN(new_n7525_));
  NAND2_X1   g07333(.A1(new_n7523_), .A2(new_n7525_), .ZN(new_n7526_));
  AOI21_X1   g07334(.A1(new_n7519_), .A2(new_n7506_), .B(new_n7526_), .ZN(new_n7527_));
  NOR3_X1    g07335(.A1(new_n7516_), .A2(\asqrt[61] ), .A3(new_n7489_), .ZN(new_n7528_));
  OAI21_X1   g07336(.A1(new_n7503_), .A2(new_n7528_), .B(new_n7517_), .ZN(new_n7529_));
  AOI21_X1   g07337(.A1(new_n7529_), .A2(\asqrt[62] ), .B(new_n7523_), .ZN(new_n7530_));
  AOI21_X1   g07338(.A1(\asqrt[31] ), .A2(new_n7157_), .B(new_n7184_), .ZN(new_n7531_));
  OR3_X2     g07339(.A1(new_n7531_), .A2(new_n193_), .A3(new_n7524_), .Z(new_n7532_));
  NAND2_X1   g07340(.A1(new_n7145_), .A2(new_n7164_), .ZN(new_n7533_));
  NOR4_X1    g07341(.A1(new_n7207_), .A2(new_n7148_), .A3(new_n7161_), .A4(new_n7533_), .ZN(new_n7534_));
  NAND2_X1   g07342(.A1(new_n7534_), .A2(new_n7153_), .ZN(new_n7535_));
  NAND2_X1   g07343(.A1(new_n7532_), .A2(new_n7535_), .ZN(new_n7536_));
  AOI21_X1   g07344(.A1(new_n7530_), .A2(new_n7519_), .B(new_n7536_), .ZN(new_n7537_));
  OAI21_X1   g07345(.A1(\asqrt[63] ), .A2(new_n7527_), .B(new_n7537_), .ZN(\asqrt[30] ));
  INV_X1     g07346(.I(\asqrt[30] ), .ZN(new_n7539_));
  NOR2_X1    g07347(.A1(\a[58] ), .A2(\a[59] ), .ZN(new_n7540_));
  INV_X1     g07348(.I(new_n7540_), .ZN(new_n7541_));
  NOR2_X1    g07349(.A1(new_n7541_), .A2(\a[60] ), .ZN(new_n7542_));
  INV_X1     g07350(.I(\a[60] ), .ZN(new_n7543_));
  INV_X1     g07351(.I(new_n7503_), .ZN(new_n7544_));
  INV_X1     g07352(.I(new_n7472_), .ZN(new_n7545_));
  INV_X1     g07353(.I(new_n7440_), .ZN(new_n7546_));
  INV_X1     g07354(.I(new_n7413_), .ZN(new_n7547_));
  INV_X1     g07355(.I(new_n7386_), .ZN(new_n7548_));
  INV_X1     g07356(.I(new_n7360_), .ZN(new_n7549_));
  INV_X1     g07357(.I(new_n7334_), .ZN(new_n7550_));
  INV_X1     g07358(.I(new_n7303_), .ZN(new_n7551_));
  NOR3_X1    g07359(.A1(new_n7302_), .A2(\asqrt[41] ), .A3(new_n7269_), .ZN(new_n7552_));
  NOR2_X1    g07360(.A1(new_n7552_), .A2(new_n7308_), .ZN(new_n7553_));
  OAI21_X1   g07361(.A1(new_n7553_), .A2(new_n7551_), .B(\asqrt[42] ), .ZN(new_n7554_));
  NAND2_X1   g07362(.A1(new_n7554_), .A2(new_n3218_), .ZN(new_n7555_));
  OAI21_X1   g07363(.A1(new_n7555_), .A2(new_n7328_), .B(new_n7550_), .ZN(new_n7556_));
  NAND3_X1   g07364(.A1(new_n7556_), .A2(new_n2954_), .A3(new_n7329_), .ZN(new_n7557_));
  AOI22_X1   g07365(.A1(new_n7557_), .A2(new_n7343_), .B1(\asqrt[44] ), .B2(new_n7352_), .ZN(new_n7558_));
  OAI21_X1   g07366(.A1(new_n7558_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n7559_));
  OAI21_X1   g07367(.A1(new_n7559_), .A2(new_n7354_), .B(new_n7549_), .ZN(new_n7560_));
  NAND3_X1   g07368(.A1(new_n7560_), .A2(new_n2229_), .A3(new_n7355_), .ZN(new_n7561_));
  AOI22_X1   g07369(.A1(new_n7561_), .A2(new_n7369_), .B1(\asqrt[47] ), .B2(new_n7378_), .ZN(new_n7562_));
  OAI21_X1   g07370(.A1(new_n7562_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n7563_));
  OAI21_X1   g07371(.A1(new_n7563_), .A2(new_n7380_), .B(new_n7548_), .ZN(new_n7564_));
  NAND3_X1   g07372(.A1(new_n7564_), .A2(new_n1612_), .A3(new_n7381_), .ZN(new_n7565_));
  AOI22_X1   g07373(.A1(new_n7565_), .A2(new_n7395_), .B1(\asqrt[50] ), .B2(new_n7404_), .ZN(new_n7566_));
  OAI21_X1   g07374(.A1(new_n7566_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n7567_));
  OAI21_X1   g07375(.A1(new_n7567_), .A2(new_n7406_), .B(new_n7547_), .ZN(new_n7568_));
  NAND3_X1   g07376(.A1(new_n7568_), .A2(new_n1103_), .A3(new_n7407_), .ZN(new_n7569_));
  AOI22_X1   g07377(.A1(new_n7569_), .A2(new_n7422_), .B1(\asqrt[53] ), .B2(new_n7451_), .ZN(new_n7570_));
  OAI21_X1   g07378(.A1(new_n7570_), .A2(new_n904_), .B(new_n823_), .ZN(new_n7571_));
  OAI21_X1   g07379(.A1(new_n7571_), .A2(new_n7453_), .B(new_n7546_), .ZN(new_n7572_));
  NAND3_X1   g07380(.A1(new_n7572_), .A2(new_n703_), .A3(new_n7454_), .ZN(new_n7573_));
  AOI22_X1   g07381(.A1(new_n7573_), .A2(new_n7449_), .B1(\asqrt[56] ), .B2(new_n7483_), .ZN(new_n7574_));
  OAI21_X1   g07382(.A1(new_n7574_), .A2(new_n531_), .B(new_n436_), .ZN(new_n7575_));
  OAI21_X1   g07383(.A1(new_n7575_), .A2(new_n7485_), .B(new_n7545_), .ZN(new_n7576_));
  NAND3_X1   g07384(.A1(new_n7576_), .A2(new_n327_), .A3(new_n7486_), .ZN(new_n7577_));
  AOI22_X1   g07385(.A1(new_n7577_), .A2(new_n7481_), .B1(\asqrt[59] ), .B2(new_n7514_), .ZN(new_n7578_));
  OAI21_X1   g07386(.A1(new_n7578_), .A2(new_n306_), .B(new_n218_), .ZN(new_n7579_));
  OAI21_X1   g07387(.A1(new_n7579_), .A2(new_n7516_), .B(new_n7544_), .ZN(new_n7580_));
  NAND3_X1   g07388(.A1(new_n7580_), .A2(new_n207_), .A3(new_n7517_), .ZN(new_n7581_));
  AOI22_X1   g07389(.A1(new_n7581_), .A2(new_n7512_), .B1(new_n7529_), .B2(\asqrt[62] ), .ZN(new_n7582_));
  OAI21_X1   g07390(.A1(new_n7582_), .A2(new_n7526_), .B(new_n193_), .ZN(new_n7583_));
  AOI21_X1   g07391(.A1(new_n7583_), .A2(new_n7537_), .B(new_n7543_), .ZN(new_n7584_));
  OAI21_X1   g07392(.A1(new_n7584_), .A2(new_n7542_), .B(\asqrt[31] ), .ZN(new_n7585_));
  INV_X1     g07393(.I(new_n7585_), .ZN(new_n7586_));
  OAI21_X1   g07394(.A1(\a[60] ), .A2(new_n7541_), .B(new_n7164_), .ZN(new_n7587_));
  NOR4_X1    g07395(.A1(new_n7207_), .A2(new_n7185_), .A3(new_n7161_), .A4(new_n7587_), .ZN(new_n7588_));
  INV_X1     g07396(.I(new_n7588_), .ZN(new_n7589_));
  NOR2_X1    g07397(.A1(new_n7584_), .A2(new_n7589_), .ZN(new_n7590_));
  AOI21_X1   g07398(.A1(new_n7583_), .A2(new_n7537_), .B(new_n7171_), .ZN(new_n7591_));
  INV_X1     g07399(.I(\a[61] ), .ZN(new_n7592_));
  AOI21_X1   g07400(.A1(\asqrt[30] ), .A2(new_n7543_), .B(new_n7592_), .ZN(new_n7593_));
  NOR3_X1    g07401(.A1(new_n7590_), .A2(new_n7593_), .A3(new_n7591_), .ZN(new_n7594_));
  OAI21_X1   g07402(.A1(new_n7594_), .A2(new_n7586_), .B(\asqrt[32] ), .ZN(new_n7595_));
  NOR2_X1    g07403(.A1(new_n7527_), .A2(\asqrt[63] ), .ZN(new_n7596_));
  INV_X1     g07404(.I(new_n7519_), .ZN(new_n7597_));
  INV_X1     g07405(.I(new_n7523_), .ZN(new_n7598_));
  NAND2_X1   g07406(.A1(new_n7506_), .A2(new_n7598_), .ZN(new_n7599_));
  INV_X1     g07407(.I(new_n7536_), .ZN(new_n7600_));
  OAI21_X1   g07408(.A1(new_n7597_), .A2(new_n7599_), .B(new_n7600_), .ZN(new_n7601_));
  OAI21_X1   g07409(.A1(new_n7596_), .A2(new_n7601_), .B(new_n7170_), .ZN(new_n7602_));
  NOR2_X1    g07410(.A1(new_n7597_), .A2(new_n7599_), .ZN(new_n7603_));
  OAI21_X1   g07411(.A1(new_n7534_), .A2(new_n7168_), .B(new_n7153_), .ZN(new_n7604_));
  NAND2_X1   g07412(.A1(new_n7532_), .A2(new_n7604_), .ZN(new_n7605_));
  NOR3_X1    g07413(.A1(new_n7596_), .A2(new_n7603_), .A3(new_n7605_), .ZN(new_n7606_));
  INV_X1     g07414(.I(new_n7606_), .ZN(new_n7607_));
  AOI21_X1   g07415(.A1(new_n7607_), .A2(new_n7602_), .B(new_n7190_), .ZN(new_n7608_));
  NOR3_X1    g07416(.A1(new_n7591_), .A2(new_n7606_), .A3(\a[62] ), .ZN(new_n7609_));
  AOI21_X1   g07417(.A1(\asqrt[30] ), .A2(\a[60] ), .B(new_n7542_), .ZN(new_n7610_));
  OAI21_X1   g07418(.A1(new_n7610_), .A2(new_n7229_), .B(new_n6824_), .ZN(new_n7611_));
  OAI22_X1   g07419(.A1(new_n7594_), .A2(new_n7611_), .B1(new_n7608_), .B2(new_n7609_), .ZN(new_n7612_));
  AOI21_X1   g07420(.A1(new_n7612_), .A2(new_n7595_), .B(new_n6356_), .ZN(new_n7613_));
  NOR3_X1    g07421(.A1(new_n7290_), .A2(new_n7189_), .A3(new_n7195_), .ZN(new_n7614_));
  NAND3_X1   g07422(.A1(\asqrt[30] ), .A2(new_n7211_), .A3(new_n7275_), .ZN(new_n7615_));
  AOI22_X1   g07423(.A1(new_n7615_), .A2(new_n7290_), .B1(\asqrt[30] ), .B2(new_n7614_), .ZN(new_n7616_));
  AOI21_X1   g07424(.A1(new_n7583_), .A2(new_n7537_), .B(\a[60] ), .ZN(new_n7617_));
  OAI21_X1   g07425(.A1(new_n7592_), .A2(new_n7617_), .B(new_n7602_), .ZN(new_n7618_));
  OAI21_X1   g07426(.A1(new_n7618_), .A2(new_n7590_), .B(new_n7585_), .ZN(new_n7619_));
  AOI21_X1   g07427(.A1(new_n7619_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n7620_));
  AOI21_X1   g07428(.A1(new_n7620_), .A2(new_n7612_), .B(new_n7616_), .ZN(new_n7621_));
  OAI21_X1   g07429(.A1(new_n7621_), .A2(new_n7613_), .B(\asqrt[34] ), .ZN(new_n7622_));
  INV_X1     g07430(.I(new_n7622_), .ZN(new_n7623_));
  NOR2_X1    g07431(.A1(new_n7210_), .A2(new_n7206_), .ZN(new_n7624_));
  INV_X1     g07432(.I(new_n7624_), .ZN(new_n7625_));
  NOR2_X1    g07433(.A1(new_n7199_), .A2(new_n7212_), .ZN(new_n7626_));
  NOR3_X1    g07434(.A1(new_n7279_), .A2(new_n7625_), .A3(new_n7626_), .ZN(new_n7627_));
  NOR3_X1    g07435(.A1(new_n7539_), .A2(new_n7279_), .A3(new_n7626_), .ZN(new_n7628_));
  INV_X1     g07436(.I(new_n7628_), .ZN(new_n7629_));
  AOI22_X1   g07437(.A1(new_n7629_), .A2(new_n7625_), .B1(\asqrt[30] ), .B2(new_n7627_), .ZN(new_n7630_));
  NOR3_X1    g07438(.A1(new_n7621_), .A2(new_n7613_), .A3(\asqrt[34] ), .ZN(new_n7631_));
  NOR2_X1    g07439(.A1(new_n7631_), .A2(new_n7630_), .ZN(new_n7632_));
  OAI21_X1   g07440(.A1(new_n7632_), .A2(new_n7623_), .B(\asqrt[35] ), .ZN(new_n7633_));
  NOR2_X1    g07441(.A1(new_n7292_), .A2(new_n7284_), .ZN(new_n7634_));
  NOR3_X1    g07442(.A1(new_n7539_), .A2(new_n7214_), .A3(new_n7634_), .ZN(new_n7635_));
  INV_X1     g07443(.I(new_n7635_), .ZN(new_n7636_));
  NOR3_X1    g07444(.A1(new_n7634_), .A2(new_n7214_), .A3(new_n7289_), .ZN(new_n7637_));
  AOI22_X1   g07445(.A1(new_n7636_), .A2(new_n7289_), .B1(\asqrt[30] ), .B2(new_n7637_), .ZN(new_n7638_));
  INV_X1     g07446(.I(new_n7638_), .ZN(new_n7639_));
  NAND2_X1   g07447(.A1(new_n7622_), .A2(new_n5708_), .ZN(new_n7640_));
  OAI21_X1   g07448(.A1(new_n7632_), .A2(new_n7640_), .B(new_n7639_), .ZN(new_n7641_));
  AOI21_X1   g07449(.A1(new_n7641_), .A2(new_n7633_), .B(new_n5277_), .ZN(new_n7642_));
  NOR3_X1    g07450(.A1(new_n7224_), .A2(new_n7233_), .A3(new_n7231_), .ZN(new_n7643_));
  NOR3_X1    g07451(.A1(new_n7539_), .A2(new_n7224_), .A3(new_n7233_), .ZN(new_n7644_));
  INV_X1     g07452(.I(new_n7644_), .ZN(new_n7645_));
  AOI22_X1   g07453(.A1(new_n7645_), .A2(new_n7231_), .B1(\asqrt[30] ), .B2(new_n7643_), .ZN(new_n7646_));
  OAI21_X1   g07454(.A1(new_n7630_), .A2(new_n7631_), .B(new_n7622_), .ZN(new_n7647_));
  AOI21_X1   g07455(.A1(new_n7647_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n7648_));
  AOI21_X1   g07456(.A1(new_n7648_), .A2(new_n7641_), .B(new_n7646_), .ZN(new_n7649_));
  OAI21_X1   g07457(.A1(new_n7649_), .A2(new_n7642_), .B(\asqrt[37] ), .ZN(new_n7650_));
  INV_X1     g07458(.I(new_n7650_), .ZN(new_n7651_));
  NOR2_X1    g07459(.A1(new_n7234_), .A2(new_n7242_), .ZN(new_n7652_));
  NOR3_X1    g07460(.A1(new_n7539_), .A2(new_n7288_), .A3(new_n7652_), .ZN(new_n7653_));
  INV_X1     g07461(.I(new_n7653_), .ZN(new_n7654_));
  NOR3_X1    g07462(.A1(new_n7652_), .A2(new_n7288_), .A3(new_n7241_), .ZN(new_n7655_));
  AOI22_X1   g07463(.A1(new_n7654_), .A2(new_n7241_), .B1(\asqrt[30] ), .B2(new_n7655_), .ZN(new_n7656_));
  NOR3_X1    g07464(.A1(new_n7649_), .A2(new_n7642_), .A3(\asqrt[37] ), .ZN(new_n7657_));
  NOR2_X1    g07465(.A1(new_n7657_), .A2(new_n7656_), .ZN(new_n7658_));
  OAI21_X1   g07466(.A1(new_n7658_), .A2(new_n7651_), .B(\asqrt[38] ), .ZN(new_n7659_));
  INV_X1     g07467(.I(new_n7248_), .ZN(new_n7660_));
  NOR3_X1    g07468(.A1(new_n7244_), .A2(new_n7321_), .A3(new_n7660_), .ZN(new_n7661_));
  NOR3_X1    g07469(.A1(new_n7539_), .A2(new_n7244_), .A3(new_n7321_), .ZN(new_n7662_));
  INV_X1     g07470(.I(new_n7662_), .ZN(new_n7663_));
  AOI22_X1   g07471(.A1(new_n7663_), .A2(new_n7660_), .B1(\asqrt[30] ), .B2(new_n7661_), .ZN(new_n7664_));
  INV_X1     g07472(.I(new_n7664_), .ZN(new_n7665_));
  NAND2_X1   g07473(.A1(new_n7650_), .A2(new_n4696_), .ZN(new_n7666_));
  OAI21_X1   g07474(.A1(new_n7658_), .A2(new_n7666_), .B(new_n7665_), .ZN(new_n7667_));
  AOI21_X1   g07475(.A1(new_n7667_), .A2(new_n7659_), .B(new_n4298_), .ZN(new_n7668_));
  NOR3_X1    g07476(.A1(new_n7539_), .A2(new_n7253_), .A3(new_n7258_), .ZN(new_n7669_));
  INV_X1     g07477(.I(new_n7669_), .ZN(new_n7670_));
  NOR3_X1    g07478(.A1(new_n7253_), .A2(new_n7274_), .A3(new_n7258_), .ZN(new_n7671_));
  AOI22_X1   g07479(.A1(new_n7670_), .A2(new_n7274_), .B1(\asqrt[30] ), .B2(new_n7671_), .ZN(new_n7672_));
  OAI21_X1   g07480(.A1(new_n7656_), .A2(new_n7657_), .B(new_n7650_), .ZN(new_n7673_));
  AOI21_X1   g07481(.A1(new_n7673_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n7674_));
  AOI21_X1   g07482(.A1(new_n7674_), .A2(new_n7667_), .B(new_n7672_), .ZN(new_n7675_));
  OAI21_X1   g07483(.A1(new_n7675_), .A2(new_n7668_), .B(\asqrt[40] ), .ZN(new_n7676_));
  INV_X1     g07484(.I(new_n7676_), .ZN(new_n7677_));
  INV_X1     g07485(.I(new_n7311_), .ZN(new_n7678_));
  NOR3_X1    g07486(.A1(new_n7678_), .A2(new_n7300_), .A3(new_n7266_), .ZN(new_n7679_));
  NOR3_X1    g07487(.A1(new_n7539_), .A2(new_n7300_), .A3(new_n7678_), .ZN(new_n7680_));
  INV_X1     g07488(.I(new_n7680_), .ZN(new_n7681_));
  AOI22_X1   g07489(.A1(new_n7681_), .A2(new_n7266_), .B1(\asqrt[30] ), .B2(new_n7679_), .ZN(new_n7682_));
  NOR3_X1    g07490(.A1(new_n7675_), .A2(new_n7668_), .A3(\asqrt[40] ), .ZN(new_n7683_));
  NOR2_X1    g07491(.A1(new_n7683_), .A2(new_n7682_), .ZN(new_n7684_));
  OAI21_X1   g07492(.A1(new_n7684_), .A2(new_n7677_), .B(\asqrt[41] ), .ZN(new_n7685_));
  INV_X1     g07493(.I(new_n7273_), .ZN(new_n7686_));
  NOR3_X1    g07494(.A1(new_n7539_), .A2(new_n7269_), .A3(new_n7325_), .ZN(new_n7687_));
  INV_X1     g07495(.I(new_n7687_), .ZN(new_n7688_));
  NOR3_X1    g07496(.A1(new_n7269_), .A2(new_n7325_), .A3(new_n7686_), .ZN(new_n7689_));
  AOI22_X1   g07497(.A1(new_n7688_), .A2(new_n7686_), .B1(\asqrt[30] ), .B2(new_n7689_), .ZN(new_n7690_));
  INV_X1     g07498(.I(new_n7690_), .ZN(new_n7691_));
  NAND2_X1   g07499(.A1(new_n7676_), .A2(new_n3782_), .ZN(new_n7692_));
  OAI21_X1   g07500(.A1(new_n7684_), .A2(new_n7692_), .B(new_n7691_), .ZN(new_n7693_));
  AOI21_X1   g07501(.A1(new_n7693_), .A2(new_n7685_), .B(new_n3419_), .ZN(new_n7694_));
  NOR3_X1    g07502(.A1(new_n7551_), .A2(new_n7309_), .A3(new_n7552_), .ZN(new_n7695_));
  NOR3_X1    g07503(.A1(new_n7539_), .A2(new_n7551_), .A3(new_n7552_), .ZN(new_n7696_));
  INV_X1     g07504(.I(new_n7696_), .ZN(new_n7697_));
  AOI22_X1   g07505(.A1(new_n7697_), .A2(new_n7309_), .B1(\asqrt[30] ), .B2(new_n7695_), .ZN(new_n7698_));
  OAI21_X1   g07506(.A1(new_n7682_), .A2(new_n7683_), .B(new_n7676_), .ZN(new_n7699_));
  AOI21_X1   g07507(.A1(new_n7699_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n7700_));
  AOI21_X1   g07508(.A1(new_n7700_), .A2(new_n7693_), .B(new_n7698_), .ZN(new_n7701_));
  OAI21_X1   g07509(.A1(new_n7701_), .A2(new_n7694_), .B(\asqrt[43] ), .ZN(new_n7702_));
  INV_X1     g07510(.I(new_n7702_), .ZN(new_n7703_));
  INV_X1     g07511(.I(new_n7320_), .ZN(new_n7704_));
  NAND2_X1   g07512(.A1(new_n7303_), .A2(new_n3419_), .ZN(new_n7705_));
  NOR2_X1    g07513(.A1(new_n7553_), .A2(new_n7705_), .ZN(new_n7706_));
  NOR3_X1    g07514(.A1(new_n7539_), .A2(new_n7315_), .A3(new_n7706_), .ZN(new_n7707_));
  INV_X1     g07515(.I(new_n7707_), .ZN(new_n7708_));
  NOR3_X1    g07516(.A1(new_n7706_), .A2(new_n7315_), .A3(new_n7704_), .ZN(new_n7709_));
  AOI22_X1   g07517(.A1(new_n7708_), .A2(new_n7704_), .B1(\asqrt[30] ), .B2(new_n7709_), .ZN(new_n7710_));
  NOR3_X1    g07518(.A1(new_n7701_), .A2(new_n7694_), .A3(\asqrt[43] ), .ZN(new_n7711_));
  NOR2_X1    g07519(.A1(new_n7711_), .A2(new_n7710_), .ZN(new_n7712_));
  OAI21_X1   g07520(.A1(new_n7712_), .A2(new_n7703_), .B(\asqrt[44] ), .ZN(new_n7713_));
  NOR3_X1    g07521(.A1(new_n7330_), .A2(new_n7550_), .A3(new_n7335_), .ZN(new_n7714_));
  NOR3_X1    g07522(.A1(new_n7539_), .A2(new_n7330_), .A3(new_n7335_), .ZN(new_n7715_));
  INV_X1     g07523(.I(new_n7715_), .ZN(new_n7716_));
  AOI22_X1   g07524(.A1(new_n7716_), .A2(new_n7550_), .B1(\asqrt[30] ), .B2(new_n7714_), .ZN(new_n7717_));
  INV_X1     g07525(.I(new_n7717_), .ZN(new_n7718_));
  NAND2_X1   g07526(.A1(new_n7702_), .A2(new_n2954_), .ZN(new_n7719_));
  OAI21_X1   g07527(.A1(new_n7712_), .A2(new_n7719_), .B(new_n7718_), .ZN(new_n7720_));
  AOI21_X1   g07528(.A1(new_n7720_), .A2(new_n7713_), .B(new_n2641_), .ZN(new_n7721_));
  INV_X1     g07529(.I(new_n7337_), .ZN(new_n7722_));
  NOR2_X1    g07530(.A1(new_n7336_), .A2(new_n7344_), .ZN(new_n7723_));
  NOR3_X1    g07531(.A1(new_n7539_), .A2(new_n7722_), .A3(new_n7723_), .ZN(new_n7724_));
  INV_X1     g07532(.I(new_n7724_), .ZN(new_n7725_));
  NOR3_X1    g07533(.A1(new_n7722_), .A2(new_n7723_), .A3(new_n7343_), .ZN(new_n7726_));
  AOI22_X1   g07534(.A1(new_n7725_), .A2(new_n7343_), .B1(\asqrt[30] ), .B2(new_n7726_), .ZN(new_n7727_));
  OAI21_X1   g07535(.A1(new_n7710_), .A2(new_n7711_), .B(new_n7702_), .ZN(new_n7728_));
  AOI21_X1   g07536(.A1(new_n7728_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n7729_));
  AOI21_X1   g07537(.A1(new_n7729_), .A2(new_n7720_), .B(new_n7727_), .ZN(new_n7730_));
  OAI21_X1   g07538(.A1(new_n7730_), .A2(new_n7721_), .B(\asqrt[46] ), .ZN(new_n7731_));
  INV_X1     g07539(.I(new_n7731_), .ZN(new_n7732_));
  INV_X1     g07540(.I(new_n7351_), .ZN(new_n7733_));
  INV_X1     g07541(.I(new_n7345_), .ZN(new_n7734_));
  INV_X1     g07542(.I(new_n7353_), .ZN(new_n7735_));
  NOR2_X1    g07543(.A1(new_n7735_), .A2(new_n7734_), .ZN(new_n7736_));
  NOR3_X1    g07544(.A1(new_n7736_), .A2(new_n7346_), .A3(new_n7733_), .ZN(new_n7737_));
  NOR3_X1    g07545(.A1(new_n7539_), .A2(new_n7346_), .A3(new_n7736_), .ZN(new_n7738_));
  INV_X1     g07546(.I(new_n7738_), .ZN(new_n7739_));
  AOI22_X1   g07547(.A1(new_n7739_), .A2(new_n7733_), .B1(\asqrt[30] ), .B2(new_n7737_), .ZN(new_n7740_));
  NOR3_X1    g07548(.A1(new_n7730_), .A2(new_n7721_), .A3(\asqrt[46] ), .ZN(new_n7741_));
  NOR2_X1    g07549(.A1(new_n7741_), .A2(new_n7740_), .ZN(new_n7742_));
  OAI21_X1   g07550(.A1(new_n7742_), .A2(new_n7732_), .B(\asqrt[47] ), .ZN(new_n7743_));
  NOR3_X1    g07551(.A1(new_n7539_), .A2(new_n7356_), .A3(new_n7361_), .ZN(new_n7744_));
  INV_X1     g07552(.I(new_n7744_), .ZN(new_n7745_));
  NOR3_X1    g07553(.A1(new_n7356_), .A2(new_n7549_), .A3(new_n7361_), .ZN(new_n7746_));
  AOI22_X1   g07554(.A1(new_n7745_), .A2(new_n7549_), .B1(\asqrt[30] ), .B2(new_n7746_), .ZN(new_n7747_));
  INV_X1     g07555(.I(new_n7747_), .ZN(new_n7748_));
  NAND2_X1   g07556(.A1(new_n7731_), .A2(new_n2229_), .ZN(new_n7749_));
  OAI21_X1   g07557(.A1(new_n7742_), .A2(new_n7749_), .B(new_n7748_), .ZN(new_n7750_));
  AOI21_X1   g07558(.A1(new_n7750_), .A2(new_n7743_), .B(new_n1956_), .ZN(new_n7751_));
  INV_X1     g07559(.I(new_n7363_), .ZN(new_n7752_));
  NOR2_X1    g07560(.A1(new_n7362_), .A2(new_n7370_), .ZN(new_n7753_));
  NOR3_X1    g07561(.A1(new_n7752_), .A2(new_n7753_), .A3(new_n7369_), .ZN(new_n7754_));
  NOR3_X1    g07562(.A1(new_n7539_), .A2(new_n7752_), .A3(new_n7753_), .ZN(new_n7755_));
  INV_X1     g07563(.I(new_n7755_), .ZN(new_n7756_));
  AOI22_X1   g07564(.A1(new_n7756_), .A2(new_n7369_), .B1(\asqrt[30] ), .B2(new_n7754_), .ZN(new_n7757_));
  OAI21_X1   g07565(.A1(new_n7740_), .A2(new_n7741_), .B(new_n7731_), .ZN(new_n7758_));
  AOI21_X1   g07566(.A1(new_n7758_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n7759_));
  AOI21_X1   g07567(.A1(new_n7759_), .A2(new_n7750_), .B(new_n7757_), .ZN(new_n7760_));
  OAI21_X1   g07568(.A1(new_n7760_), .A2(new_n7751_), .B(\asqrt[49] ), .ZN(new_n7761_));
  INV_X1     g07569(.I(new_n7761_), .ZN(new_n7762_));
  INV_X1     g07570(.I(new_n7377_), .ZN(new_n7763_));
  INV_X1     g07571(.I(new_n7371_), .ZN(new_n7764_));
  INV_X1     g07572(.I(new_n7379_), .ZN(new_n7765_));
  NOR2_X1    g07573(.A1(new_n7765_), .A2(new_n7764_), .ZN(new_n7766_));
  NOR3_X1    g07574(.A1(new_n7539_), .A2(new_n7372_), .A3(new_n7766_), .ZN(new_n7767_));
  INV_X1     g07575(.I(new_n7767_), .ZN(new_n7768_));
  NOR3_X1    g07576(.A1(new_n7766_), .A2(new_n7372_), .A3(new_n7763_), .ZN(new_n7769_));
  AOI22_X1   g07577(.A1(new_n7768_), .A2(new_n7763_), .B1(\asqrt[30] ), .B2(new_n7769_), .ZN(new_n7770_));
  NOR3_X1    g07578(.A1(new_n7760_), .A2(new_n7751_), .A3(\asqrt[49] ), .ZN(new_n7771_));
  NOR2_X1    g07579(.A1(new_n7771_), .A2(new_n7770_), .ZN(new_n7772_));
  OAI21_X1   g07580(.A1(new_n7772_), .A2(new_n7762_), .B(\asqrt[50] ), .ZN(new_n7773_));
  NOR3_X1    g07581(.A1(new_n7382_), .A2(new_n7548_), .A3(new_n7387_), .ZN(new_n7774_));
  NOR3_X1    g07582(.A1(new_n7539_), .A2(new_n7382_), .A3(new_n7387_), .ZN(new_n7775_));
  INV_X1     g07583(.I(new_n7775_), .ZN(new_n7776_));
  AOI22_X1   g07584(.A1(new_n7776_), .A2(new_n7548_), .B1(\asqrt[30] ), .B2(new_n7774_), .ZN(new_n7777_));
  INV_X1     g07585(.I(new_n7777_), .ZN(new_n7778_));
  NAND2_X1   g07586(.A1(new_n7761_), .A2(new_n1612_), .ZN(new_n7779_));
  OAI21_X1   g07587(.A1(new_n7772_), .A2(new_n7779_), .B(new_n7778_), .ZN(new_n7780_));
  AOI21_X1   g07588(.A1(new_n7780_), .A2(new_n7773_), .B(new_n1376_), .ZN(new_n7781_));
  INV_X1     g07589(.I(new_n7389_), .ZN(new_n7782_));
  NOR2_X1    g07590(.A1(new_n7388_), .A2(new_n7396_), .ZN(new_n7783_));
  NOR3_X1    g07591(.A1(new_n7539_), .A2(new_n7782_), .A3(new_n7783_), .ZN(new_n7784_));
  INV_X1     g07592(.I(new_n7784_), .ZN(new_n7785_));
  NOR3_X1    g07593(.A1(new_n7782_), .A2(new_n7395_), .A3(new_n7783_), .ZN(new_n7786_));
  AOI22_X1   g07594(.A1(new_n7785_), .A2(new_n7395_), .B1(\asqrt[30] ), .B2(new_n7786_), .ZN(new_n7787_));
  OAI21_X1   g07595(.A1(new_n7770_), .A2(new_n7771_), .B(new_n7761_), .ZN(new_n7788_));
  AOI21_X1   g07596(.A1(new_n7788_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n7789_));
  AOI21_X1   g07597(.A1(new_n7789_), .A2(new_n7780_), .B(new_n7787_), .ZN(new_n7790_));
  OAI21_X1   g07598(.A1(new_n7790_), .A2(new_n7781_), .B(\asqrt[52] ), .ZN(new_n7791_));
  INV_X1     g07599(.I(new_n7403_), .ZN(new_n7792_));
  INV_X1     g07600(.I(new_n7397_), .ZN(new_n7793_));
  INV_X1     g07601(.I(new_n7405_), .ZN(new_n7794_));
  NOR2_X1    g07602(.A1(new_n7794_), .A2(new_n7793_), .ZN(new_n7795_));
  NOR3_X1    g07603(.A1(new_n7795_), .A2(new_n7398_), .A3(new_n7792_), .ZN(new_n7796_));
  NOR3_X1    g07604(.A1(new_n7539_), .A2(new_n7398_), .A3(new_n7795_), .ZN(new_n7797_));
  INV_X1     g07605(.I(new_n7797_), .ZN(new_n7798_));
  AOI22_X1   g07606(.A1(new_n7798_), .A2(new_n7792_), .B1(\asqrt[30] ), .B2(new_n7796_), .ZN(new_n7799_));
  INV_X1     g07607(.I(new_n7799_), .ZN(new_n7800_));
  INV_X1     g07608(.I(new_n7770_), .ZN(new_n7801_));
  INV_X1     g07609(.I(new_n7751_), .ZN(new_n7802_));
  NAND2_X1   g07610(.A1(new_n7802_), .A2(new_n1806_), .ZN(new_n7803_));
  OAI21_X1   g07611(.A1(new_n7803_), .A2(new_n7760_), .B(new_n7801_), .ZN(new_n7804_));
  AOI21_X1   g07612(.A1(new_n7804_), .A2(new_n7761_), .B(new_n1612_), .ZN(new_n7805_));
  INV_X1     g07613(.I(new_n7779_), .ZN(new_n7806_));
  AOI21_X1   g07614(.A1(new_n7806_), .A2(new_n7804_), .B(new_n7777_), .ZN(new_n7807_));
  OAI21_X1   g07615(.A1(new_n7807_), .A2(new_n7805_), .B(\asqrt[51] ), .ZN(new_n7808_));
  NAND2_X1   g07616(.A1(new_n7808_), .A2(new_n1256_), .ZN(new_n7809_));
  OAI21_X1   g07617(.A1(new_n7809_), .A2(new_n7790_), .B(new_n7800_), .ZN(new_n7810_));
  AOI21_X1   g07618(.A1(new_n7810_), .A2(new_n7791_), .B(new_n1103_), .ZN(new_n7811_));
  NOR3_X1    g07619(.A1(new_n7539_), .A2(new_n7408_), .A3(new_n7450_), .ZN(new_n7812_));
  INV_X1     g07620(.I(new_n7812_), .ZN(new_n7813_));
  NOR3_X1    g07621(.A1(new_n7408_), .A2(new_n7547_), .A3(new_n7450_), .ZN(new_n7814_));
  AOI22_X1   g07622(.A1(new_n7813_), .A2(new_n7547_), .B1(\asqrt[30] ), .B2(new_n7814_), .ZN(new_n7815_));
  INV_X1     g07623(.I(new_n7787_), .ZN(new_n7816_));
  NAND2_X1   g07624(.A1(new_n7773_), .A2(new_n1376_), .ZN(new_n7817_));
  OAI21_X1   g07625(.A1(new_n7817_), .A2(new_n7807_), .B(new_n7816_), .ZN(new_n7818_));
  AOI21_X1   g07626(.A1(new_n7818_), .A2(new_n7808_), .B(new_n1256_), .ZN(new_n7819_));
  NOR2_X1    g07627(.A1(new_n7819_), .A2(\asqrt[53] ), .ZN(new_n7820_));
  AOI21_X1   g07628(.A1(new_n7820_), .A2(new_n7810_), .B(new_n7815_), .ZN(new_n7821_));
  OAI21_X1   g07629(.A1(new_n7821_), .A2(new_n7811_), .B(\asqrt[54] ), .ZN(new_n7822_));
  INV_X1     g07630(.I(new_n7416_), .ZN(new_n7823_));
  NOR2_X1    g07631(.A1(new_n7423_), .A2(new_n7415_), .ZN(new_n7824_));
  NOR3_X1    g07632(.A1(new_n7823_), .A2(new_n7422_), .A3(new_n7824_), .ZN(new_n7825_));
  NOR3_X1    g07633(.A1(new_n7539_), .A2(new_n7823_), .A3(new_n7824_), .ZN(new_n7826_));
  INV_X1     g07634(.I(new_n7826_), .ZN(new_n7827_));
  AOI22_X1   g07635(.A1(new_n7827_), .A2(new_n7422_), .B1(\asqrt[30] ), .B2(new_n7825_), .ZN(new_n7828_));
  INV_X1     g07636(.I(new_n7828_), .ZN(new_n7829_));
  NOR2_X1    g07637(.A1(new_n7781_), .A2(\asqrt[52] ), .ZN(new_n7830_));
  AOI21_X1   g07638(.A1(new_n7830_), .A2(new_n7818_), .B(new_n7799_), .ZN(new_n7831_));
  OAI21_X1   g07639(.A1(new_n7831_), .A2(new_n7819_), .B(\asqrt[53] ), .ZN(new_n7832_));
  NAND2_X1   g07640(.A1(new_n7832_), .A2(new_n904_), .ZN(new_n7833_));
  OAI21_X1   g07641(.A1(new_n7833_), .A2(new_n7821_), .B(new_n7829_), .ZN(new_n7834_));
  AOI21_X1   g07642(.A1(new_n7834_), .A2(new_n7822_), .B(new_n823_), .ZN(new_n7835_));
  NOR2_X1    g07643(.A1(new_n7434_), .A2(new_n7427_), .ZN(new_n7836_));
  NOR3_X1    g07644(.A1(new_n7539_), .A2(new_n7425_), .A3(new_n7836_), .ZN(new_n7837_));
  INV_X1     g07645(.I(new_n7837_), .ZN(new_n7838_));
  NOR3_X1    g07646(.A1(new_n7836_), .A2(new_n7425_), .A3(new_n7433_), .ZN(new_n7839_));
  AOI22_X1   g07647(.A1(new_n7838_), .A2(new_n7433_), .B1(\asqrt[30] ), .B2(new_n7839_), .ZN(new_n7840_));
  INV_X1     g07648(.I(new_n7815_), .ZN(new_n7841_));
  NAND2_X1   g07649(.A1(new_n7791_), .A2(new_n1103_), .ZN(new_n7842_));
  OAI21_X1   g07650(.A1(new_n7842_), .A2(new_n7831_), .B(new_n7841_), .ZN(new_n7843_));
  AOI21_X1   g07651(.A1(new_n7843_), .A2(new_n7832_), .B(new_n904_), .ZN(new_n7844_));
  NOR2_X1    g07652(.A1(new_n7844_), .A2(\asqrt[55] ), .ZN(new_n7845_));
  AOI21_X1   g07653(.A1(new_n7845_), .A2(new_n7834_), .B(new_n7840_), .ZN(new_n7846_));
  OAI21_X1   g07654(.A1(new_n7846_), .A2(new_n7835_), .B(\asqrt[56] ), .ZN(new_n7847_));
  NOR3_X1    g07655(.A1(new_n7436_), .A2(new_n7546_), .A3(new_n7482_), .ZN(new_n7848_));
  NOR3_X1    g07656(.A1(new_n7539_), .A2(new_n7436_), .A3(new_n7482_), .ZN(new_n7849_));
  INV_X1     g07657(.I(new_n7849_), .ZN(new_n7850_));
  AOI22_X1   g07658(.A1(new_n7850_), .A2(new_n7546_), .B1(\asqrt[30] ), .B2(new_n7848_), .ZN(new_n7851_));
  INV_X1     g07659(.I(new_n7851_), .ZN(new_n7852_));
  NOR3_X1    g07660(.A1(new_n7790_), .A2(new_n7781_), .A3(\asqrt[52] ), .ZN(new_n7853_));
  OAI21_X1   g07661(.A1(new_n7799_), .A2(new_n7853_), .B(new_n7791_), .ZN(new_n7854_));
  AOI21_X1   g07662(.A1(new_n7854_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n7855_));
  AOI21_X1   g07663(.A1(new_n7855_), .A2(new_n7843_), .B(new_n7828_), .ZN(new_n7856_));
  OAI21_X1   g07664(.A1(new_n7856_), .A2(new_n7844_), .B(\asqrt[55] ), .ZN(new_n7857_));
  NAND2_X1   g07665(.A1(new_n7857_), .A2(new_n703_), .ZN(new_n7858_));
  OAI21_X1   g07666(.A1(new_n7858_), .A2(new_n7846_), .B(new_n7852_), .ZN(new_n7859_));
  AOI21_X1   g07667(.A1(new_n7859_), .A2(new_n7847_), .B(new_n531_), .ZN(new_n7860_));
  INV_X1     g07668(.I(new_n7443_), .ZN(new_n7861_));
  NOR2_X1    g07669(.A1(new_n7455_), .A2(new_n7442_), .ZN(new_n7862_));
  NOR3_X1    g07670(.A1(new_n7539_), .A2(new_n7861_), .A3(new_n7862_), .ZN(new_n7863_));
  INV_X1     g07671(.I(new_n7863_), .ZN(new_n7864_));
  NOR3_X1    g07672(.A1(new_n7861_), .A2(new_n7449_), .A3(new_n7862_), .ZN(new_n7865_));
  AOI22_X1   g07673(.A1(new_n7864_), .A2(new_n7449_), .B1(\asqrt[30] ), .B2(new_n7865_), .ZN(new_n7866_));
  NOR3_X1    g07674(.A1(new_n7856_), .A2(\asqrt[55] ), .A3(new_n7844_), .ZN(new_n7867_));
  OAI21_X1   g07675(.A1(new_n7840_), .A2(new_n7867_), .B(new_n7857_), .ZN(new_n7868_));
  AOI21_X1   g07676(.A1(new_n7868_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n7869_));
  AOI21_X1   g07677(.A1(new_n7869_), .A2(new_n7859_), .B(new_n7866_), .ZN(new_n7870_));
  OAI21_X1   g07678(.A1(new_n7870_), .A2(new_n7860_), .B(\asqrt[58] ), .ZN(new_n7871_));
  NOR2_X1    g07679(.A1(new_n7466_), .A2(new_n7459_), .ZN(new_n7872_));
  NOR3_X1    g07680(.A1(new_n7872_), .A2(new_n7457_), .A3(new_n7465_), .ZN(new_n7873_));
  NOR3_X1    g07681(.A1(new_n7539_), .A2(new_n7457_), .A3(new_n7872_), .ZN(new_n7874_));
  INV_X1     g07682(.I(new_n7874_), .ZN(new_n7875_));
  AOI22_X1   g07683(.A1(new_n7875_), .A2(new_n7465_), .B1(\asqrt[30] ), .B2(new_n7873_), .ZN(new_n7876_));
  INV_X1     g07684(.I(new_n7876_), .ZN(new_n7877_));
  INV_X1     g07685(.I(new_n7840_), .ZN(new_n7878_));
  NAND2_X1   g07686(.A1(new_n7822_), .A2(new_n823_), .ZN(new_n7879_));
  OAI21_X1   g07687(.A1(new_n7879_), .A2(new_n7856_), .B(new_n7878_), .ZN(new_n7880_));
  AOI21_X1   g07688(.A1(new_n7880_), .A2(new_n7857_), .B(new_n703_), .ZN(new_n7881_));
  NOR2_X1    g07689(.A1(new_n7835_), .A2(\asqrt[56] ), .ZN(new_n7882_));
  AOI21_X1   g07690(.A1(new_n7882_), .A2(new_n7880_), .B(new_n7851_), .ZN(new_n7883_));
  OAI21_X1   g07691(.A1(new_n7883_), .A2(new_n7881_), .B(\asqrt[57] ), .ZN(new_n7884_));
  NAND2_X1   g07692(.A1(new_n7884_), .A2(new_n436_), .ZN(new_n7885_));
  OAI21_X1   g07693(.A1(new_n7885_), .A2(new_n7870_), .B(new_n7877_), .ZN(new_n7886_));
  AOI21_X1   g07694(.A1(new_n7886_), .A2(new_n7871_), .B(new_n327_), .ZN(new_n7887_));
  NOR3_X1    g07695(.A1(new_n7539_), .A2(new_n7468_), .A3(new_n7513_), .ZN(new_n7888_));
  INV_X1     g07696(.I(new_n7888_), .ZN(new_n7889_));
  NOR3_X1    g07697(.A1(new_n7468_), .A2(new_n7545_), .A3(new_n7513_), .ZN(new_n7890_));
  AOI22_X1   g07698(.A1(new_n7889_), .A2(new_n7545_), .B1(\asqrt[30] ), .B2(new_n7890_), .ZN(new_n7891_));
  INV_X1     g07699(.I(new_n7866_), .ZN(new_n7892_));
  NAND2_X1   g07700(.A1(new_n7847_), .A2(new_n531_), .ZN(new_n7893_));
  OAI21_X1   g07701(.A1(new_n7893_), .A2(new_n7883_), .B(new_n7892_), .ZN(new_n7894_));
  AOI21_X1   g07702(.A1(new_n7894_), .A2(new_n7884_), .B(new_n436_), .ZN(new_n7895_));
  NOR2_X1    g07703(.A1(new_n7895_), .A2(\asqrt[59] ), .ZN(new_n7896_));
  AOI21_X1   g07704(.A1(new_n7896_), .A2(new_n7886_), .B(new_n7891_), .ZN(new_n7897_));
  OAI21_X1   g07705(.A1(new_n7897_), .A2(new_n7887_), .B(\asqrt[60] ), .ZN(new_n7898_));
  INV_X1     g07706(.I(new_n7475_), .ZN(new_n7899_));
  NOR2_X1    g07707(.A1(new_n7487_), .A2(new_n7474_), .ZN(new_n7900_));
  NOR3_X1    g07708(.A1(new_n7899_), .A2(new_n7481_), .A3(new_n7900_), .ZN(new_n7901_));
  NOR3_X1    g07709(.A1(new_n7539_), .A2(new_n7899_), .A3(new_n7900_), .ZN(new_n7902_));
  INV_X1     g07710(.I(new_n7902_), .ZN(new_n7903_));
  AOI22_X1   g07711(.A1(new_n7903_), .A2(new_n7481_), .B1(\asqrt[30] ), .B2(new_n7901_), .ZN(new_n7904_));
  INV_X1     g07712(.I(new_n7904_), .ZN(new_n7905_));
  NOR2_X1    g07713(.A1(new_n7860_), .A2(\asqrt[58] ), .ZN(new_n7906_));
  AOI21_X1   g07714(.A1(new_n7906_), .A2(new_n7894_), .B(new_n7876_), .ZN(new_n7907_));
  OAI21_X1   g07715(.A1(new_n7907_), .A2(new_n7895_), .B(\asqrt[59] ), .ZN(new_n7908_));
  NAND2_X1   g07716(.A1(new_n7908_), .A2(new_n306_), .ZN(new_n7909_));
  OAI21_X1   g07717(.A1(new_n7909_), .A2(new_n7897_), .B(new_n7905_), .ZN(new_n7910_));
  AOI21_X1   g07718(.A1(new_n7910_), .A2(new_n7898_), .B(new_n218_), .ZN(new_n7911_));
  NOR2_X1    g07719(.A1(new_n7491_), .A2(new_n7497_), .ZN(new_n7912_));
  NOR3_X1    g07720(.A1(new_n7539_), .A2(new_n7489_), .A3(new_n7912_), .ZN(new_n7913_));
  INV_X1     g07721(.I(new_n7913_), .ZN(new_n7914_));
  NOR3_X1    g07722(.A1(new_n7912_), .A2(new_n7489_), .A3(new_n7496_), .ZN(new_n7915_));
  AOI22_X1   g07723(.A1(new_n7914_), .A2(new_n7496_), .B1(\asqrt[30] ), .B2(new_n7915_), .ZN(new_n7916_));
  INV_X1     g07724(.I(new_n7891_), .ZN(new_n7917_));
  NAND2_X1   g07725(.A1(new_n7871_), .A2(new_n327_), .ZN(new_n7918_));
  OAI21_X1   g07726(.A1(new_n7918_), .A2(new_n7907_), .B(new_n7917_), .ZN(new_n7919_));
  AOI21_X1   g07727(.A1(new_n7919_), .A2(new_n7908_), .B(new_n306_), .ZN(new_n7920_));
  NOR2_X1    g07728(.A1(new_n7920_), .A2(\asqrt[61] ), .ZN(new_n7921_));
  AOI21_X1   g07729(.A1(new_n7921_), .A2(new_n7910_), .B(new_n7916_), .ZN(new_n7922_));
  OAI21_X1   g07730(.A1(new_n7922_), .A2(new_n7911_), .B(\asqrt[62] ), .ZN(new_n7923_));
  NOR3_X1    g07731(.A1(new_n7499_), .A2(new_n7544_), .A3(new_n7528_), .ZN(new_n7924_));
  NOR3_X1    g07732(.A1(new_n7539_), .A2(new_n7499_), .A3(new_n7528_), .ZN(new_n7925_));
  INV_X1     g07733(.I(new_n7925_), .ZN(new_n7926_));
  AOI22_X1   g07734(.A1(new_n7926_), .A2(new_n7544_), .B1(\asqrt[30] ), .B2(new_n7924_), .ZN(new_n7927_));
  INV_X1     g07735(.I(new_n7927_), .ZN(new_n7928_));
  NOR3_X1    g07736(.A1(new_n7870_), .A2(\asqrt[58] ), .A3(new_n7860_), .ZN(new_n7929_));
  OAI21_X1   g07737(.A1(new_n7876_), .A2(new_n7929_), .B(new_n7871_), .ZN(new_n7930_));
  AOI21_X1   g07738(.A1(new_n7930_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n7931_));
  AOI21_X1   g07739(.A1(new_n7931_), .A2(new_n7919_), .B(new_n7904_), .ZN(new_n7932_));
  OAI21_X1   g07740(.A1(new_n7932_), .A2(new_n7920_), .B(\asqrt[61] ), .ZN(new_n7933_));
  NAND2_X1   g07741(.A1(new_n7933_), .A2(new_n207_), .ZN(new_n7934_));
  OAI21_X1   g07742(.A1(new_n7934_), .A2(new_n7922_), .B(new_n7928_), .ZN(new_n7935_));
  INV_X1     g07743(.I(new_n7603_), .ZN(new_n7936_));
  NAND4_X1   g07744(.A1(\asqrt[30] ), .A2(new_n7506_), .A3(new_n7511_), .A4(new_n7581_), .ZN(new_n7937_));
  NAND2_X1   g07745(.A1(new_n7506_), .A2(new_n7581_), .ZN(new_n7938_));
  OAI21_X1   g07746(.A1(new_n7539_), .A2(new_n7938_), .B(new_n7512_), .ZN(new_n7939_));
  NAND2_X1   g07747(.A1(new_n7939_), .A2(new_n7937_), .ZN(new_n7940_));
  NOR2_X1    g07748(.A1(new_n7582_), .A2(new_n7598_), .ZN(new_n7941_));
  NAND2_X1   g07749(.A1(\asqrt[30] ), .A2(new_n7941_), .ZN(new_n7942_));
  NAND3_X1   g07750(.A1(new_n7940_), .A2(new_n7936_), .A3(new_n7942_), .ZN(new_n7943_));
  AOI21_X1   g07751(.A1(new_n7935_), .A2(new_n7923_), .B(new_n7943_), .ZN(new_n7944_));
  NOR3_X1    g07752(.A1(new_n7932_), .A2(\asqrt[61] ), .A3(new_n7920_), .ZN(new_n7945_));
  OAI21_X1   g07753(.A1(new_n7916_), .A2(new_n7945_), .B(new_n7933_), .ZN(new_n7946_));
  AOI21_X1   g07754(.A1(new_n7946_), .A2(\asqrt[62] ), .B(new_n7940_), .ZN(new_n7947_));
  OAI21_X1   g07755(.A1(new_n7539_), .A2(new_n7598_), .B(new_n7582_), .ZN(new_n7948_));
  NOR2_X1    g07756(.A1(new_n7941_), .A2(new_n193_), .ZN(new_n7949_));
  NAND2_X1   g07757(.A1(new_n7948_), .A2(new_n7949_), .ZN(new_n7950_));
  INV_X1     g07758(.I(new_n7950_), .ZN(new_n7951_));
  AND3_X2    g07759(.A1(new_n7522_), .A2(new_n7520_), .A3(new_n7535_), .Z(new_n7952_));
  NAND4_X1   g07760(.A1(new_n7936_), .A2(new_n7583_), .A3(new_n7532_), .A4(new_n7952_), .ZN(new_n7953_));
  INV_X1     g07761(.I(new_n7953_), .ZN(new_n7954_));
  NOR2_X1    g07762(.A1(new_n7951_), .A2(new_n7954_), .ZN(new_n7955_));
  INV_X1     g07763(.I(new_n7955_), .ZN(new_n7956_));
  AOI21_X1   g07764(.A1(new_n7947_), .A2(new_n7935_), .B(new_n7956_), .ZN(new_n7957_));
  OAI21_X1   g07765(.A1(\asqrt[63] ), .A2(new_n7944_), .B(new_n7957_), .ZN(\asqrt[29] ));
  NOR2_X1    g07766(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n7959_));
  INV_X1     g07767(.I(new_n7959_), .ZN(new_n7960_));
  NOR2_X1    g07768(.A1(new_n7960_), .A2(\a[58] ), .ZN(new_n7961_));
  INV_X1     g07769(.I(new_n7961_), .ZN(new_n7962_));
  NAND2_X1   g07770(.A1(new_n7935_), .A2(new_n7923_), .ZN(new_n7963_));
  INV_X1     g07771(.I(new_n7943_), .ZN(new_n7964_));
  AOI21_X1   g07772(.A1(new_n7963_), .A2(new_n7964_), .B(\asqrt[63] ), .ZN(new_n7965_));
  INV_X1     g07773(.I(new_n7935_), .ZN(new_n7966_));
  INV_X1     g07774(.I(new_n7940_), .ZN(new_n7967_));
  NAND2_X1   g07775(.A1(new_n7923_), .A2(new_n7967_), .ZN(new_n7968_));
  OAI21_X1   g07776(.A1(new_n7966_), .A2(new_n7968_), .B(new_n7955_), .ZN(new_n7969_));
  OAI21_X1   g07777(.A1(new_n7965_), .A2(new_n7969_), .B(\a[58] ), .ZN(new_n7970_));
  AOI21_X1   g07778(.A1(new_n7970_), .A2(new_n7962_), .B(new_n7539_), .ZN(new_n7971_));
  INV_X1     g07779(.I(\a[58] ), .ZN(new_n7972_));
  INV_X1     g07780(.I(new_n7916_), .ZN(new_n7973_));
  NAND2_X1   g07781(.A1(new_n7898_), .A2(new_n218_), .ZN(new_n7974_));
  OAI21_X1   g07782(.A1(new_n7974_), .A2(new_n7932_), .B(new_n7973_), .ZN(new_n7975_));
  NAND3_X1   g07783(.A1(new_n7975_), .A2(new_n207_), .A3(new_n7933_), .ZN(new_n7976_));
  AOI22_X1   g07784(.A1(new_n7976_), .A2(new_n7928_), .B1(new_n7946_), .B2(\asqrt[62] ), .ZN(new_n7977_));
  OAI21_X1   g07785(.A1(new_n7977_), .A2(new_n7943_), .B(new_n193_), .ZN(new_n7978_));
  AOI21_X1   g07786(.A1(new_n7978_), .A2(new_n7957_), .B(new_n7972_), .ZN(new_n7979_));
  NAND4_X1   g07787(.A1(new_n7936_), .A2(new_n7532_), .A3(new_n7535_), .A4(new_n7962_), .ZN(new_n7980_));
  NOR2_X1    g07788(.A1(new_n7980_), .A2(new_n7596_), .ZN(new_n7981_));
  INV_X1     g07789(.I(new_n7981_), .ZN(new_n7982_));
  NOR2_X1    g07790(.A1(new_n7979_), .A2(new_n7982_), .ZN(new_n7983_));
  AOI21_X1   g07791(.A1(new_n7978_), .A2(new_n7957_), .B(new_n7541_), .ZN(new_n7984_));
  INV_X1     g07792(.I(\a[59] ), .ZN(new_n7985_));
  AOI21_X1   g07793(.A1(\asqrt[29] ), .A2(new_n7972_), .B(new_n7985_), .ZN(new_n7986_));
  NOR3_X1    g07794(.A1(new_n7983_), .A2(new_n7986_), .A3(new_n7984_), .ZN(new_n7987_));
  OAI21_X1   g07795(.A1(new_n7987_), .A2(new_n7971_), .B(\asqrt[31] ), .ZN(new_n7988_));
  OAI21_X1   g07796(.A1(new_n7965_), .A2(new_n7969_), .B(new_n7540_), .ZN(new_n7989_));
  NOR2_X1    g07797(.A1(new_n7966_), .A2(new_n7968_), .ZN(new_n7990_));
  NOR2_X1    g07798(.A1(new_n7954_), .A2(new_n7539_), .ZN(new_n7991_));
  NAND2_X1   g07799(.A1(new_n7950_), .A2(new_n7991_), .ZN(new_n7992_));
  NOR3_X1    g07800(.A1(new_n7965_), .A2(new_n7990_), .A3(new_n7992_), .ZN(new_n7993_));
  INV_X1     g07801(.I(new_n7993_), .ZN(new_n7994_));
  AOI21_X1   g07802(.A1(new_n7994_), .A2(new_n7989_), .B(new_n7543_), .ZN(new_n7995_));
  NOR3_X1    g07803(.A1(new_n7993_), .A2(new_n7984_), .A3(\a[60] ), .ZN(new_n7996_));
  AOI21_X1   g07804(.A1(\asqrt[29] ), .A2(\a[58] ), .B(new_n7961_), .ZN(new_n7997_));
  OAI21_X1   g07805(.A1(new_n7997_), .A2(new_n7539_), .B(new_n7229_), .ZN(new_n7998_));
  OAI22_X1   g07806(.A1(new_n7987_), .A2(new_n7998_), .B1(new_n7995_), .B2(new_n7996_), .ZN(new_n7999_));
  AOI21_X1   g07807(.A1(new_n7999_), .A2(new_n7988_), .B(new_n6824_), .ZN(new_n8000_));
  INV_X1     g07808(.I(new_n7618_), .ZN(new_n8001_));
  NOR3_X1    g07809(.A1(new_n7586_), .A2(new_n8001_), .A3(new_n7590_), .ZN(new_n8002_));
  NOR2_X1    g07810(.A1(new_n7586_), .A2(new_n7590_), .ZN(new_n8003_));
  NAND2_X1   g07811(.A1(\asqrt[29] ), .A2(new_n8003_), .ZN(new_n8004_));
  AOI22_X1   g07812(.A1(new_n8004_), .A2(new_n8001_), .B1(\asqrt[29] ), .B2(new_n8002_), .ZN(new_n8005_));
  OAI21_X1   g07813(.A1(new_n7979_), .A2(new_n7961_), .B(\asqrt[30] ), .ZN(new_n8006_));
  AOI21_X1   g07814(.A1(new_n7978_), .A2(new_n7957_), .B(\a[58] ), .ZN(new_n8007_));
  OAI21_X1   g07815(.A1(new_n7985_), .A2(new_n8007_), .B(new_n7989_), .ZN(new_n8008_));
  OAI21_X1   g07816(.A1(new_n8008_), .A2(new_n7983_), .B(new_n8006_), .ZN(new_n8009_));
  AOI21_X1   g07817(.A1(new_n8009_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n8010_));
  AOI21_X1   g07818(.A1(new_n8010_), .A2(new_n7999_), .B(new_n8005_), .ZN(new_n8011_));
  OAI21_X1   g07819(.A1(new_n8011_), .A2(new_n8000_), .B(\asqrt[33] ), .ZN(new_n8012_));
  INV_X1     g07820(.I(new_n8012_), .ZN(new_n8013_));
  NOR2_X1    g07821(.A1(new_n7608_), .A2(new_n7609_), .ZN(new_n8014_));
  NOR2_X1    g07822(.A1(new_n7594_), .A2(new_n7611_), .ZN(new_n8015_));
  INV_X1     g07823(.I(new_n8015_), .ZN(new_n8016_));
  NAND4_X1   g07824(.A1(\asqrt[29] ), .A2(new_n7595_), .A3(new_n8014_), .A4(new_n8016_), .ZN(new_n8017_));
  AND3_X2    g07825(.A1(\asqrt[29] ), .A2(new_n7595_), .A3(new_n8016_), .Z(new_n8018_));
  OAI21_X1   g07826(.A1(new_n8018_), .A2(new_n8014_), .B(new_n8017_), .ZN(new_n8019_));
  INV_X1     g07827(.I(new_n8019_), .ZN(new_n8020_));
  NOR3_X1    g07828(.A1(new_n8011_), .A2(new_n8000_), .A3(\asqrt[33] ), .ZN(new_n8021_));
  NOR2_X1    g07829(.A1(new_n8021_), .A2(new_n8020_), .ZN(new_n8022_));
  OAI21_X1   g07830(.A1(new_n8022_), .A2(new_n8013_), .B(\asqrt[34] ), .ZN(new_n8023_));
  INV_X1     g07831(.I(new_n7616_), .ZN(new_n8024_));
  INV_X1     g07832(.I(new_n7613_), .ZN(new_n8025_));
  NAND2_X1   g07833(.A1(new_n7620_), .A2(new_n7612_), .ZN(new_n8026_));
  NAND3_X1   g07834(.A1(\asqrt[29] ), .A2(new_n8025_), .A3(new_n8026_), .ZN(new_n8027_));
  AND3_X2    g07835(.A1(new_n8025_), .A2(new_n7616_), .A3(new_n8026_), .Z(new_n8028_));
  AOI22_X1   g07836(.A1(new_n8027_), .A2(new_n8024_), .B1(\asqrt[29] ), .B2(new_n8028_), .ZN(new_n8029_));
  INV_X1     g07837(.I(new_n8029_), .ZN(new_n8030_));
  NAND2_X1   g07838(.A1(new_n8012_), .A2(new_n6077_), .ZN(new_n8031_));
  OAI21_X1   g07839(.A1(new_n8022_), .A2(new_n8031_), .B(new_n8030_), .ZN(new_n8032_));
  AOI21_X1   g07840(.A1(new_n8032_), .A2(new_n8023_), .B(new_n5708_), .ZN(new_n8033_));
  INV_X1     g07841(.I(new_n7630_), .ZN(new_n8034_));
  NOR3_X1    g07842(.A1(new_n7623_), .A2(new_n8034_), .A3(new_n7631_), .ZN(new_n8035_));
  INV_X1     g07843(.I(\asqrt[29] ), .ZN(new_n8036_));
  NOR3_X1    g07844(.A1(new_n8036_), .A2(new_n7623_), .A3(new_n7631_), .ZN(new_n8037_));
  INV_X1     g07845(.I(new_n8037_), .ZN(new_n8038_));
  AOI22_X1   g07846(.A1(new_n8038_), .A2(new_n8034_), .B1(\asqrt[29] ), .B2(new_n8035_), .ZN(new_n8039_));
  OAI21_X1   g07847(.A1(new_n8020_), .A2(new_n8021_), .B(new_n8012_), .ZN(new_n8040_));
  AOI21_X1   g07848(.A1(new_n8040_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n8041_));
  AOI21_X1   g07849(.A1(new_n8041_), .A2(new_n8032_), .B(new_n8039_), .ZN(new_n8042_));
  OAI21_X1   g07850(.A1(new_n8042_), .A2(new_n8033_), .B(\asqrt[36] ), .ZN(new_n8043_));
  INV_X1     g07851(.I(new_n8043_), .ZN(new_n8044_));
  INV_X1     g07852(.I(new_n7632_), .ZN(new_n8045_));
  INV_X1     g07853(.I(new_n7640_), .ZN(new_n8046_));
  NAND2_X1   g07854(.A1(new_n8045_), .A2(new_n8046_), .ZN(new_n8047_));
  NAND3_X1   g07855(.A1(\asqrt[29] ), .A2(new_n7633_), .A3(new_n8047_), .ZN(new_n8048_));
  AND3_X2    g07856(.A1(new_n8047_), .A2(new_n7633_), .A3(new_n7638_), .Z(new_n8049_));
  AOI22_X1   g07857(.A1(new_n8048_), .A2(new_n7639_), .B1(\asqrt[29] ), .B2(new_n8049_), .ZN(new_n8050_));
  NOR3_X1    g07858(.A1(new_n8042_), .A2(new_n8033_), .A3(\asqrt[36] ), .ZN(new_n8051_));
  NOR2_X1    g07859(.A1(new_n8051_), .A2(new_n8050_), .ZN(new_n8052_));
  OAI21_X1   g07860(.A1(new_n8052_), .A2(new_n8044_), .B(\asqrt[37] ), .ZN(new_n8053_));
  INV_X1     g07861(.I(new_n7646_), .ZN(new_n8054_));
  INV_X1     g07862(.I(new_n7641_), .ZN(new_n8055_));
  INV_X1     g07863(.I(new_n7648_), .ZN(new_n8056_));
  NOR2_X1    g07864(.A1(new_n8056_), .A2(new_n8055_), .ZN(new_n8057_));
  NOR3_X1    g07865(.A1(new_n8057_), .A2(new_n7642_), .A3(new_n8054_), .ZN(new_n8058_));
  NOR3_X1    g07866(.A1(new_n8036_), .A2(new_n7642_), .A3(new_n8057_), .ZN(new_n8059_));
  INV_X1     g07867(.I(new_n8059_), .ZN(new_n8060_));
  AOI22_X1   g07868(.A1(new_n8060_), .A2(new_n8054_), .B1(\asqrt[29] ), .B2(new_n8058_), .ZN(new_n8061_));
  INV_X1     g07869(.I(new_n8061_), .ZN(new_n8062_));
  NAND2_X1   g07870(.A1(new_n8043_), .A2(new_n5024_), .ZN(new_n8063_));
  OAI21_X1   g07871(.A1(new_n8052_), .A2(new_n8063_), .B(new_n8062_), .ZN(new_n8064_));
  AOI21_X1   g07872(.A1(new_n8064_), .A2(new_n8053_), .B(new_n4696_), .ZN(new_n8065_));
  INV_X1     g07873(.I(new_n7656_), .ZN(new_n8066_));
  NOR3_X1    g07874(.A1(new_n8036_), .A2(new_n7651_), .A3(new_n7657_), .ZN(new_n8067_));
  INV_X1     g07875(.I(new_n8067_), .ZN(new_n8068_));
  NOR3_X1    g07876(.A1(new_n7651_), .A2(new_n8066_), .A3(new_n7657_), .ZN(new_n8069_));
  AOI22_X1   g07877(.A1(new_n8068_), .A2(new_n8066_), .B1(\asqrt[29] ), .B2(new_n8069_), .ZN(new_n8070_));
  OAI21_X1   g07878(.A1(new_n8050_), .A2(new_n8051_), .B(new_n8043_), .ZN(new_n8071_));
  AOI21_X1   g07879(.A1(new_n8071_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n8072_));
  AOI21_X1   g07880(.A1(new_n8072_), .A2(new_n8064_), .B(new_n8070_), .ZN(new_n8073_));
  OAI21_X1   g07881(.A1(new_n8073_), .A2(new_n8065_), .B(\asqrt[39] ), .ZN(new_n8074_));
  INV_X1     g07882(.I(new_n8074_), .ZN(new_n8075_));
  NOR2_X1    g07883(.A1(new_n7658_), .A2(new_n7666_), .ZN(new_n8076_));
  INV_X1     g07884(.I(new_n8076_), .ZN(new_n8077_));
  AND3_X2    g07885(.A1(new_n8077_), .A2(new_n7659_), .A3(new_n7664_), .Z(new_n8078_));
  NAND3_X1   g07886(.A1(\asqrt[29] ), .A2(new_n7659_), .A3(new_n8077_), .ZN(new_n8079_));
  AOI22_X1   g07887(.A1(new_n8079_), .A2(new_n7665_), .B1(\asqrt[29] ), .B2(new_n8078_), .ZN(new_n8080_));
  NOR3_X1    g07888(.A1(new_n8073_), .A2(new_n8065_), .A3(\asqrt[39] ), .ZN(new_n8081_));
  NOR2_X1    g07889(.A1(new_n8081_), .A2(new_n8080_), .ZN(new_n8082_));
  OAI21_X1   g07890(.A1(new_n8082_), .A2(new_n8075_), .B(\asqrt[40] ), .ZN(new_n8083_));
  INV_X1     g07891(.I(new_n7672_), .ZN(new_n8084_));
  INV_X1     g07892(.I(new_n7667_), .ZN(new_n8085_));
  INV_X1     g07893(.I(new_n7674_), .ZN(new_n8086_));
  NOR2_X1    g07894(.A1(new_n8086_), .A2(new_n8085_), .ZN(new_n8087_));
  NOR3_X1    g07895(.A1(new_n8036_), .A2(new_n7668_), .A3(new_n8087_), .ZN(new_n8088_));
  INV_X1     g07896(.I(new_n8088_), .ZN(new_n8089_));
  NOR3_X1    g07897(.A1(new_n8087_), .A2(new_n7668_), .A3(new_n8084_), .ZN(new_n8090_));
  AOI22_X1   g07898(.A1(new_n8089_), .A2(new_n8084_), .B1(\asqrt[29] ), .B2(new_n8090_), .ZN(new_n8091_));
  INV_X1     g07899(.I(new_n8091_), .ZN(new_n8092_));
  NAND2_X1   g07900(.A1(new_n8074_), .A2(new_n4071_), .ZN(new_n8093_));
  OAI21_X1   g07901(.A1(new_n8082_), .A2(new_n8093_), .B(new_n8092_), .ZN(new_n8094_));
  AOI21_X1   g07902(.A1(new_n8094_), .A2(new_n8083_), .B(new_n3782_), .ZN(new_n8095_));
  INV_X1     g07903(.I(new_n7682_), .ZN(new_n8096_));
  NOR3_X1    g07904(.A1(new_n7677_), .A2(new_n7683_), .A3(new_n8096_), .ZN(new_n8097_));
  NOR3_X1    g07905(.A1(new_n8036_), .A2(new_n7677_), .A3(new_n7683_), .ZN(new_n8098_));
  INV_X1     g07906(.I(new_n8098_), .ZN(new_n8099_));
  AOI22_X1   g07907(.A1(new_n8099_), .A2(new_n8096_), .B1(\asqrt[29] ), .B2(new_n8097_), .ZN(new_n8100_));
  OAI21_X1   g07908(.A1(new_n8080_), .A2(new_n8081_), .B(new_n8074_), .ZN(new_n8101_));
  AOI21_X1   g07909(.A1(new_n8101_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n8102_));
  AOI21_X1   g07910(.A1(new_n8102_), .A2(new_n8094_), .B(new_n8100_), .ZN(new_n8103_));
  OAI21_X1   g07911(.A1(new_n8103_), .A2(new_n8095_), .B(\asqrt[42] ), .ZN(new_n8104_));
  INV_X1     g07912(.I(new_n8104_), .ZN(new_n8105_));
  INV_X1     g07913(.I(new_n7685_), .ZN(new_n8106_));
  NOR2_X1    g07914(.A1(new_n7684_), .A2(new_n7692_), .ZN(new_n8107_));
  NOR3_X1    g07915(.A1(new_n8036_), .A2(new_n8106_), .A3(new_n8107_), .ZN(new_n8108_));
  INV_X1     g07916(.I(new_n8108_), .ZN(new_n8109_));
  NOR3_X1    g07917(.A1(new_n8106_), .A2(new_n7691_), .A3(new_n8107_), .ZN(new_n8110_));
  AOI22_X1   g07918(.A1(new_n8109_), .A2(new_n7691_), .B1(\asqrt[29] ), .B2(new_n8110_), .ZN(new_n8111_));
  NOR3_X1    g07919(.A1(new_n8103_), .A2(new_n8095_), .A3(\asqrt[42] ), .ZN(new_n8112_));
  NOR2_X1    g07920(.A1(new_n8112_), .A2(new_n8111_), .ZN(new_n8113_));
  OAI21_X1   g07921(.A1(new_n8113_), .A2(new_n8105_), .B(\asqrt[43] ), .ZN(new_n8114_));
  INV_X1     g07922(.I(new_n7698_), .ZN(new_n8115_));
  INV_X1     g07923(.I(new_n7693_), .ZN(new_n8116_));
  INV_X1     g07924(.I(new_n7700_), .ZN(new_n8117_));
  NOR2_X1    g07925(.A1(new_n8117_), .A2(new_n8116_), .ZN(new_n8118_));
  NOR3_X1    g07926(.A1(new_n8118_), .A2(new_n7694_), .A3(new_n8115_), .ZN(new_n8119_));
  NOR3_X1    g07927(.A1(new_n8036_), .A2(new_n7694_), .A3(new_n8118_), .ZN(new_n8120_));
  INV_X1     g07928(.I(new_n8120_), .ZN(new_n8121_));
  AOI22_X1   g07929(.A1(new_n8121_), .A2(new_n8115_), .B1(\asqrt[29] ), .B2(new_n8119_), .ZN(new_n8122_));
  INV_X1     g07930(.I(new_n8122_), .ZN(new_n8123_));
  NAND2_X1   g07931(.A1(new_n8104_), .A2(new_n3218_), .ZN(new_n8124_));
  OAI21_X1   g07932(.A1(new_n8113_), .A2(new_n8124_), .B(new_n8123_), .ZN(new_n8125_));
  AOI21_X1   g07933(.A1(new_n8125_), .A2(new_n8114_), .B(new_n2954_), .ZN(new_n8126_));
  INV_X1     g07934(.I(new_n7710_), .ZN(new_n8127_));
  NOR3_X1    g07935(.A1(new_n8036_), .A2(new_n7703_), .A3(new_n7711_), .ZN(new_n8128_));
  INV_X1     g07936(.I(new_n8128_), .ZN(new_n8129_));
  NOR3_X1    g07937(.A1(new_n7703_), .A2(new_n7711_), .A3(new_n8127_), .ZN(new_n8130_));
  AOI22_X1   g07938(.A1(new_n8129_), .A2(new_n8127_), .B1(\asqrt[29] ), .B2(new_n8130_), .ZN(new_n8131_));
  OAI21_X1   g07939(.A1(new_n8111_), .A2(new_n8112_), .B(new_n8104_), .ZN(new_n8132_));
  AOI21_X1   g07940(.A1(new_n8132_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n8133_));
  AOI21_X1   g07941(.A1(new_n8133_), .A2(new_n8125_), .B(new_n8131_), .ZN(new_n8134_));
  OAI21_X1   g07942(.A1(new_n8134_), .A2(new_n8126_), .B(\asqrt[45] ), .ZN(new_n8135_));
  INV_X1     g07943(.I(new_n8135_), .ZN(new_n8136_));
  NOR2_X1    g07944(.A1(new_n7712_), .A2(new_n7719_), .ZN(new_n8137_));
  INV_X1     g07945(.I(new_n8137_), .ZN(new_n8138_));
  AND3_X2    g07946(.A1(new_n8138_), .A2(new_n7713_), .A3(new_n7717_), .Z(new_n8139_));
  NAND3_X1   g07947(.A1(\asqrt[29] ), .A2(new_n7713_), .A3(new_n8138_), .ZN(new_n8140_));
  AOI22_X1   g07948(.A1(new_n8140_), .A2(new_n7718_), .B1(\asqrt[29] ), .B2(new_n8139_), .ZN(new_n8141_));
  NOR3_X1    g07949(.A1(new_n8134_), .A2(new_n8126_), .A3(\asqrt[45] ), .ZN(new_n8142_));
  NOR2_X1    g07950(.A1(new_n8142_), .A2(new_n8141_), .ZN(new_n8143_));
  OAI21_X1   g07951(.A1(new_n8143_), .A2(new_n8136_), .B(\asqrt[46] ), .ZN(new_n8144_));
  INV_X1     g07952(.I(new_n7727_), .ZN(new_n8145_));
  INV_X1     g07953(.I(new_n7721_), .ZN(new_n8146_));
  NAND2_X1   g07954(.A1(new_n7729_), .A2(new_n7720_), .ZN(new_n8147_));
  NAND3_X1   g07955(.A1(\asqrt[29] ), .A2(new_n8146_), .A3(new_n8147_), .ZN(new_n8148_));
  AND3_X2    g07956(.A1(new_n8146_), .A2(new_n7727_), .A3(new_n8147_), .Z(new_n8149_));
  AOI22_X1   g07957(.A1(new_n8148_), .A2(new_n8145_), .B1(\asqrt[29] ), .B2(new_n8149_), .ZN(new_n8150_));
  INV_X1     g07958(.I(new_n8150_), .ZN(new_n8151_));
  NAND2_X1   g07959(.A1(new_n8135_), .A2(new_n2465_), .ZN(new_n8152_));
  OAI21_X1   g07960(.A1(new_n8143_), .A2(new_n8152_), .B(new_n8151_), .ZN(new_n8153_));
  AOI21_X1   g07961(.A1(new_n8153_), .A2(new_n8144_), .B(new_n2229_), .ZN(new_n8154_));
  INV_X1     g07962(.I(new_n7740_), .ZN(new_n8155_));
  NOR3_X1    g07963(.A1(new_n7732_), .A2(new_n7741_), .A3(new_n8155_), .ZN(new_n8156_));
  NOR3_X1    g07964(.A1(new_n8036_), .A2(new_n7732_), .A3(new_n7741_), .ZN(new_n8157_));
  INV_X1     g07965(.I(new_n8157_), .ZN(new_n8158_));
  AOI22_X1   g07966(.A1(new_n8158_), .A2(new_n8155_), .B1(\asqrt[29] ), .B2(new_n8156_), .ZN(new_n8159_));
  OAI21_X1   g07967(.A1(new_n8141_), .A2(new_n8142_), .B(new_n8135_), .ZN(new_n8160_));
  AOI21_X1   g07968(.A1(new_n8160_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n8161_));
  AOI21_X1   g07969(.A1(new_n8161_), .A2(new_n8153_), .B(new_n8159_), .ZN(new_n8162_));
  OAI21_X1   g07970(.A1(new_n8162_), .A2(new_n8154_), .B(\asqrt[48] ), .ZN(new_n8163_));
  INV_X1     g07971(.I(new_n8163_), .ZN(new_n8164_));
  INV_X1     g07972(.I(new_n7743_), .ZN(new_n8165_));
  NOR2_X1    g07973(.A1(new_n7742_), .A2(new_n7749_), .ZN(new_n8166_));
  NOR3_X1    g07974(.A1(new_n8036_), .A2(new_n8165_), .A3(new_n8166_), .ZN(new_n8167_));
  INV_X1     g07975(.I(new_n8167_), .ZN(new_n8168_));
  NOR3_X1    g07976(.A1(new_n8165_), .A2(new_n7748_), .A3(new_n8166_), .ZN(new_n8169_));
  AOI22_X1   g07977(.A1(new_n8168_), .A2(new_n7748_), .B1(\asqrt[29] ), .B2(new_n8169_), .ZN(new_n8170_));
  NOR3_X1    g07978(.A1(new_n8162_), .A2(new_n8154_), .A3(\asqrt[48] ), .ZN(new_n8171_));
  NOR2_X1    g07979(.A1(new_n8171_), .A2(new_n8170_), .ZN(new_n8172_));
  OAI21_X1   g07980(.A1(new_n8172_), .A2(new_n8164_), .B(\asqrt[49] ), .ZN(new_n8173_));
  INV_X1     g07981(.I(new_n7757_), .ZN(new_n8174_));
  NAND2_X1   g07982(.A1(new_n7759_), .A2(new_n7750_), .ZN(new_n8175_));
  AND3_X2    g07983(.A1(new_n7802_), .A2(new_n7757_), .A3(new_n8175_), .Z(new_n8176_));
  NAND3_X1   g07984(.A1(\asqrt[29] ), .A2(new_n7802_), .A3(new_n8175_), .ZN(new_n8177_));
  AOI22_X1   g07985(.A1(new_n8177_), .A2(new_n8174_), .B1(\asqrt[29] ), .B2(new_n8176_), .ZN(new_n8178_));
  INV_X1     g07986(.I(new_n8178_), .ZN(new_n8179_));
  NAND2_X1   g07987(.A1(new_n8163_), .A2(new_n1806_), .ZN(new_n8180_));
  OAI21_X1   g07988(.A1(new_n8172_), .A2(new_n8180_), .B(new_n8179_), .ZN(new_n8181_));
  AOI21_X1   g07989(.A1(new_n8181_), .A2(new_n8173_), .B(new_n1612_), .ZN(new_n8182_));
  NOR3_X1    g07990(.A1(new_n8036_), .A2(new_n7762_), .A3(new_n7771_), .ZN(new_n8183_));
  INV_X1     g07991(.I(new_n8183_), .ZN(new_n8184_));
  NOR3_X1    g07992(.A1(new_n7762_), .A2(new_n7801_), .A3(new_n7771_), .ZN(new_n8185_));
  AOI22_X1   g07993(.A1(new_n8184_), .A2(new_n7801_), .B1(\asqrt[29] ), .B2(new_n8185_), .ZN(new_n8186_));
  OAI21_X1   g07994(.A1(new_n8170_), .A2(new_n8171_), .B(new_n8163_), .ZN(new_n8187_));
  AOI21_X1   g07995(.A1(new_n8187_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n8188_));
  AOI21_X1   g07996(.A1(new_n8188_), .A2(new_n8181_), .B(new_n8186_), .ZN(new_n8189_));
  OAI21_X1   g07997(.A1(new_n8189_), .A2(new_n8182_), .B(\asqrt[51] ), .ZN(new_n8190_));
  INV_X1     g07998(.I(new_n8190_), .ZN(new_n8191_));
  NOR2_X1    g07999(.A1(new_n7772_), .A2(new_n7779_), .ZN(new_n8192_));
  NOR3_X1    g08000(.A1(new_n7805_), .A2(new_n8192_), .A3(new_n7778_), .ZN(new_n8193_));
  NOR3_X1    g08001(.A1(new_n8036_), .A2(new_n7805_), .A3(new_n8192_), .ZN(new_n8194_));
  INV_X1     g08002(.I(new_n8194_), .ZN(new_n8195_));
  AOI22_X1   g08003(.A1(new_n8195_), .A2(new_n7778_), .B1(\asqrt[29] ), .B2(new_n8193_), .ZN(new_n8196_));
  NOR3_X1    g08004(.A1(new_n8189_), .A2(new_n8182_), .A3(\asqrt[51] ), .ZN(new_n8197_));
  NOR2_X1    g08005(.A1(new_n8197_), .A2(new_n8196_), .ZN(new_n8198_));
  OAI21_X1   g08006(.A1(new_n8198_), .A2(new_n8191_), .B(\asqrt[52] ), .ZN(new_n8199_));
  NOR2_X1    g08007(.A1(new_n7817_), .A2(new_n7807_), .ZN(new_n8200_));
  NOR3_X1    g08008(.A1(new_n8036_), .A2(new_n7781_), .A3(new_n8200_), .ZN(new_n8201_));
  INV_X1     g08009(.I(new_n8201_), .ZN(new_n8202_));
  NOR3_X1    g08010(.A1(new_n8200_), .A2(new_n7781_), .A3(new_n7816_), .ZN(new_n8203_));
  AOI22_X1   g08011(.A1(new_n8202_), .A2(new_n7816_), .B1(\asqrt[29] ), .B2(new_n8203_), .ZN(new_n8204_));
  INV_X1     g08012(.I(new_n8204_), .ZN(new_n8205_));
  NAND2_X1   g08013(.A1(new_n8190_), .A2(new_n1256_), .ZN(new_n8206_));
  OAI21_X1   g08014(.A1(new_n8198_), .A2(new_n8206_), .B(new_n8205_), .ZN(new_n8207_));
  AOI21_X1   g08015(.A1(new_n8207_), .A2(new_n8199_), .B(new_n1103_), .ZN(new_n8208_));
  NOR3_X1    g08016(.A1(new_n7819_), .A2(new_n7853_), .A3(new_n7800_), .ZN(new_n8209_));
  NOR3_X1    g08017(.A1(new_n8036_), .A2(new_n7819_), .A3(new_n7853_), .ZN(new_n8210_));
  INV_X1     g08018(.I(new_n8210_), .ZN(new_n8211_));
  AOI22_X1   g08019(.A1(new_n8211_), .A2(new_n7800_), .B1(\asqrt[29] ), .B2(new_n8209_), .ZN(new_n8212_));
  OAI21_X1   g08020(.A1(new_n8196_), .A2(new_n8197_), .B(new_n8190_), .ZN(new_n8213_));
  AOI21_X1   g08021(.A1(new_n8213_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n8214_));
  AOI21_X1   g08022(.A1(new_n8214_), .A2(new_n8207_), .B(new_n8212_), .ZN(new_n8215_));
  OAI21_X1   g08023(.A1(new_n8215_), .A2(new_n8208_), .B(\asqrt[54] ), .ZN(new_n8216_));
  INV_X1     g08024(.I(new_n8216_), .ZN(new_n8217_));
  NOR2_X1    g08025(.A1(new_n7842_), .A2(new_n7831_), .ZN(new_n8218_));
  NOR3_X1    g08026(.A1(new_n8036_), .A2(new_n7811_), .A3(new_n8218_), .ZN(new_n8219_));
  INV_X1     g08027(.I(new_n8219_), .ZN(new_n8220_));
  NOR3_X1    g08028(.A1(new_n7811_), .A2(new_n8218_), .A3(new_n7841_), .ZN(new_n8221_));
  AOI22_X1   g08029(.A1(new_n8220_), .A2(new_n7841_), .B1(\asqrt[29] ), .B2(new_n8221_), .ZN(new_n8222_));
  NOR3_X1    g08030(.A1(new_n8215_), .A2(new_n8208_), .A3(\asqrt[54] ), .ZN(new_n8223_));
  NOR2_X1    g08031(.A1(new_n8223_), .A2(new_n8222_), .ZN(new_n8224_));
  OAI21_X1   g08032(.A1(new_n8224_), .A2(new_n8217_), .B(\asqrt[55] ), .ZN(new_n8225_));
  NOR2_X1    g08033(.A1(new_n7833_), .A2(new_n7821_), .ZN(new_n8226_));
  NOR3_X1    g08034(.A1(new_n8226_), .A2(new_n7844_), .A3(new_n7829_), .ZN(new_n8227_));
  NOR3_X1    g08035(.A1(new_n8036_), .A2(new_n7844_), .A3(new_n8226_), .ZN(new_n8228_));
  INV_X1     g08036(.I(new_n8228_), .ZN(new_n8229_));
  AOI22_X1   g08037(.A1(new_n8229_), .A2(new_n7829_), .B1(\asqrt[29] ), .B2(new_n8227_), .ZN(new_n8230_));
  INV_X1     g08038(.I(new_n8230_), .ZN(new_n8231_));
  NAND2_X1   g08039(.A1(new_n8216_), .A2(new_n823_), .ZN(new_n8232_));
  OAI21_X1   g08040(.A1(new_n8224_), .A2(new_n8232_), .B(new_n8231_), .ZN(new_n8233_));
  AOI21_X1   g08041(.A1(new_n8233_), .A2(new_n8225_), .B(new_n703_), .ZN(new_n8234_));
  NOR3_X1    g08042(.A1(new_n8036_), .A2(new_n7835_), .A3(new_n7867_), .ZN(new_n8235_));
  INV_X1     g08043(.I(new_n8235_), .ZN(new_n8236_));
  NOR3_X1    g08044(.A1(new_n7835_), .A2(new_n7867_), .A3(new_n7878_), .ZN(new_n8237_));
  AOI22_X1   g08045(.A1(new_n8236_), .A2(new_n7878_), .B1(\asqrt[29] ), .B2(new_n8237_), .ZN(new_n8238_));
  OAI21_X1   g08046(.A1(new_n8222_), .A2(new_n8223_), .B(new_n8216_), .ZN(new_n8239_));
  AOI21_X1   g08047(.A1(new_n8239_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n8240_));
  AOI21_X1   g08048(.A1(new_n8240_), .A2(new_n8233_), .B(new_n8238_), .ZN(new_n8241_));
  OAI21_X1   g08049(.A1(new_n8241_), .A2(new_n8234_), .B(\asqrt[57] ), .ZN(new_n8242_));
  NOR2_X1    g08050(.A1(new_n7858_), .A2(new_n7846_), .ZN(new_n8243_));
  NOR3_X1    g08051(.A1(new_n7881_), .A2(new_n8243_), .A3(new_n7852_), .ZN(new_n8244_));
  NOR3_X1    g08052(.A1(new_n8036_), .A2(new_n7881_), .A3(new_n8243_), .ZN(new_n8245_));
  INV_X1     g08053(.I(new_n8245_), .ZN(new_n8246_));
  AOI22_X1   g08054(.A1(new_n8246_), .A2(new_n7852_), .B1(\asqrt[29] ), .B2(new_n8244_), .ZN(new_n8247_));
  INV_X1     g08055(.I(new_n8247_), .ZN(new_n8248_));
  INV_X1     g08056(.I(new_n8222_), .ZN(new_n8249_));
  INV_X1     g08057(.I(new_n8196_), .ZN(new_n8250_));
  INV_X1     g08058(.I(new_n8170_), .ZN(new_n8251_));
  INV_X1     g08059(.I(new_n8141_), .ZN(new_n8252_));
  INV_X1     g08060(.I(new_n8111_), .ZN(new_n8253_));
  INV_X1     g08061(.I(new_n8080_), .ZN(new_n8254_));
  INV_X1     g08062(.I(new_n8050_), .ZN(new_n8255_));
  NAND2_X1   g08063(.A1(new_n7970_), .A2(new_n7981_), .ZN(new_n8256_));
  OAI21_X1   g08064(.A1(new_n7965_), .A2(new_n7969_), .B(new_n7972_), .ZN(new_n8257_));
  NAND2_X1   g08065(.A1(new_n8257_), .A2(\a[59] ), .ZN(new_n8258_));
  NAND3_X1   g08066(.A1(new_n8256_), .A2(new_n8258_), .A3(new_n7989_), .ZN(new_n8259_));
  AOI21_X1   g08067(.A1(new_n8259_), .A2(new_n8006_), .B(new_n7229_), .ZN(new_n8260_));
  OAI21_X1   g08068(.A1(new_n7993_), .A2(new_n7984_), .B(\a[60] ), .ZN(new_n8261_));
  NAND3_X1   g08069(.A1(new_n7994_), .A2(new_n7989_), .A3(new_n7543_), .ZN(new_n8262_));
  NAND2_X1   g08070(.A1(new_n7970_), .A2(new_n7962_), .ZN(new_n8263_));
  AOI21_X1   g08071(.A1(new_n8263_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n8264_));
  AOI22_X1   g08072(.A1(new_n8259_), .A2(new_n8264_), .B1(new_n8261_), .B2(new_n8262_), .ZN(new_n8265_));
  OAI21_X1   g08073(.A1(new_n8265_), .A2(new_n8260_), .B(\asqrt[32] ), .ZN(new_n8266_));
  NAND2_X1   g08074(.A1(new_n8266_), .A2(new_n6356_), .ZN(new_n8267_));
  OAI21_X1   g08075(.A1(new_n8267_), .A2(new_n8011_), .B(new_n8019_), .ZN(new_n8268_));
  AOI21_X1   g08076(.A1(new_n8268_), .A2(new_n8012_), .B(new_n6077_), .ZN(new_n8269_));
  INV_X1     g08077(.I(new_n8005_), .ZN(new_n8270_));
  AOI21_X1   g08078(.A1(\a[59] ), .A2(new_n8257_), .B(new_n7984_), .ZN(new_n8271_));
  AOI21_X1   g08079(.A1(new_n8271_), .A2(new_n8256_), .B(new_n7971_), .ZN(new_n8272_));
  OAI21_X1   g08080(.A1(new_n8272_), .A2(new_n7229_), .B(new_n6824_), .ZN(new_n8273_));
  OAI21_X1   g08081(.A1(new_n8273_), .A2(new_n8265_), .B(new_n8270_), .ZN(new_n8274_));
  NAND2_X1   g08082(.A1(new_n8274_), .A2(new_n8266_), .ZN(new_n8275_));
  AOI21_X1   g08083(.A1(new_n8275_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n8276_));
  AOI21_X1   g08084(.A1(new_n8276_), .A2(new_n8268_), .B(new_n8029_), .ZN(new_n8277_));
  OAI21_X1   g08085(.A1(new_n8277_), .A2(new_n8269_), .B(\asqrt[35] ), .ZN(new_n8278_));
  NAND2_X1   g08086(.A1(new_n8278_), .A2(new_n5277_), .ZN(new_n8279_));
  OAI21_X1   g08087(.A1(new_n8279_), .A2(new_n8042_), .B(new_n8255_), .ZN(new_n8280_));
  NAND3_X1   g08088(.A1(new_n8280_), .A2(new_n5024_), .A3(new_n8043_), .ZN(new_n8281_));
  AOI22_X1   g08089(.A1(new_n8281_), .A2(new_n8062_), .B1(new_n8071_), .B2(\asqrt[37] ), .ZN(new_n8282_));
  OAI21_X1   g08090(.A1(new_n8282_), .A2(new_n4696_), .B(new_n4298_), .ZN(new_n8283_));
  OAI21_X1   g08091(.A1(new_n8283_), .A2(new_n8073_), .B(new_n8254_), .ZN(new_n8284_));
  AOI21_X1   g08092(.A1(new_n8284_), .A2(new_n8074_), .B(new_n4071_), .ZN(new_n8285_));
  AOI21_X1   g08093(.A1(new_n8280_), .A2(new_n8043_), .B(new_n5024_), .ZN(new_n8286_));
  NOR3_X1    g08094(.A1(new_n8277_), .A2(new_n8269_), .A3(\asqrt[35] ), .ZN(new_n8287_));
  OAI21_X1   g08095(.A1(new_n8039_), .A2(new_n8287_), .B(new_n8278_), .ZN(new_n8288_));
  AOI21_X1   g08096(.A1(new_n8288_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n8289_));
  AOI21_X1   g08097(.A1(new_n8289_), .A2(new_n8280_), .B(new_n8061_), .ZN(new_n8290_));
  NOR3_X1    g08098(.A1(new_n8290_), .A2(\asqrt[38] ), .A3(new_n8286_), .ZN(new_n8291_));
  OAI22_X1   g08099(.A1(new_n8291_), .A2(new_n8070_), .B1(new_n8282_), .B2(new_n4696_), .ZN(new_n8292_));
  AOI21_X1   g08100(.A1(new_n8292_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n8293_));
  AOI21_X1   g08101(.A1(new_n8293_), .A2(new_n8284_), .B(new_n8091_), .ZN(new_n8294_));
  OAI21_X1   g08102(.A1(new_n8294_), .A2(new_n8285_), .B(\asqrt[41] ), .ZN(new_n8295_));
  NAND2_X1   g08103(.A1(new_n8295_), .A2(new_n3419_), .ZN(new_n8296_));
  OAI21_X1   g08104(.A1(new_n8296_), .A2(new_n8103_), .B(new_n8253_), .ZN(new_n8297_));
  AOI21_X1   g08105(.A1(new_n8297_), .A2(new_n8104_), .B(new_n3218_), .ZN(new_n8298_));
  NOR3_X1    g08106(.A1(new_n8294_), .A2(\asqrt[41] ), .A3(new_n8285_), .ZN(new_n8299_));
  OAI21_X1   g08107(.A1(new_n8100_), .A2(new_n8299_), .B(new_n8295_), .ZN(new_n8300_));
  AOI21_X1   g08108(.A1(new_n8300_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n8301_));
  AOI21_X1   g08109(.A1(new_n8301_), .A2(new_n8297_), .B(new_n8122_), .ZN(new_n8302_));
  OAI21_X1   g08110(.A1(new_n8302_), .A2(new_n8298_), .B(\asqrt[44] ), .ZN(new_n8303_));
  NAND2_X1   g08111(.A1(new_n8303_), .A2(new_n2641_), .ZN(new_n8304_));
  OAI21_X1   g08112(.A1(new_n8304_), .A2(new_n8134_), .B(new_n8252_), .ZN(new_n8305_));
  AOI21_X1   g08113(.A1(new_n8305_), .A2(new_n8135_), .B(new_n2465_), .ZN(new_n8306_));
  NOR3_X1    g08114(.A1(new_n8302_), .A2(\asqrt[44] ), .A3(new_n8298_), .ZN(new_n8307_));
  OAI21_X1   g08115(.A1(new_n8131_), .A2(new_n8307_), .B(new_n8303_), .ZN(new_n8308_));
  AOI21_X1   g08116(.A1(new_n8308_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n8309_));
  AOI21_X1   g08117(.A1(new_n8309_), .A2(new_n8305_), .B(new_n8150_), .ZN(new_n8310_));
  OAI21_X1   g08118(.A1(new_n8310_), .A2(new_n8306_), .B(\asqrt[47] ), .ZN(new_n8311_));
  NAND2_X1   g08119(.A1(new_n8311_), .A2(new_n1956_), .ZN(new_n8312_));
  OAI21_X1   g08120(.A1(new_n8312_), .A2(new_n8162_), .B(new_n8251_), .ZN(new_n8313_));
  AOI21_X1   g08121(.A1(new_n8313_), .A2(new_n8163_), .B(new_n1806_), .ZN(new_n8314_));
  NOR3_X1    g08122(.A1(new_n8310_), .A2(\asqrt[47] ), .A3(new_n8306_), .ZN(new_n8315_));
  OAI21_X1   g08123(.A1(new_n8159_), .A2(new_n8315_), .B(new_n8311_), .ZN(new_n8316_));
  AOI21_X1   g08124(.A1(new_n8316_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n8317_));
  AOI21_X1   g08125(.A1(new_n8317_), .A2(new_n8313_), .B(new_n8178_), .ZN(new_n8318_));
  OAI21_X1   g08126(.A1(new_n8318_), .A2(new_n8314_), .B(\asqrt[50] ), .ZN(new_n8319_));
  NAND2_X1   g08127(.A1(new_n8319_), .A2(new_n1376_), .ZN(new_n8320_));
  OAI21_X1   g08128(.A1(new_n8320_), .A2(new_n8189_), .B(new_n8250_), .ZN(new_n8321_));
  AOI21_X1   g08129(.A1(new_n8321_), .A2(new_n8190_), .B(new_n1256_), .ZN(new_n8322_));
  NOR3_X1    g08130(.A1(new_n8318_), .A2(\asqrt[50] ), .A3(new_n8314_), .ZN(new_n8323_));
  OAI21_X1   g08131(.A1(new_n8186_), .A2(new_n8323_), .B(new_n8319_), .ZN(new_n8324_));
  AOI21_X1   g08132(.A1(new_n8324_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n8325_));
  AOI21_X1   g08133(.A1(new_n8325_), .A2(new_n8321_), .B(new_n8204_), .ZN(new_n8326_));
  OAI21_X1   g08134(.A1(new_n8326_), .A2(new_n8322_), .B(\asqrt[53] ), .ZN(new_n8327_));
  NAND2_X1   g08135(.A1(new_n8327_), .A2(new_n904_), .ZN(new_n8328_));
  OAI21_X1   g08136(.A1(new_n8328_), .A2(new_n8215_), .B(new_n8249_), .ZN(new_n8329_));
  AOI21_X1   g08137(.A1(new_n8329_), .A2(new_n8216_), .B(new_n823_), .ZN(new_n8330_));
  NOR3_X1    g08138(.A1(new_n8326_), .A2(\asqrt[53] ), .A3(new_n8322_), .ZN(new_n8331_));
  OAI21_X1   g08139(.A1(new_n8212_), .A2(new_n8331_), .B(new_n8327_), .ZN(new_n8332_));
  AOI21_X1   g08140(.A1(new_n8332_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n8333_));
  AOI21_X1   g08141(.A1(new_n8333_), .A2(new_n8329_), .B(new_n8230_), .ZN(new_n8334_));
  OAI21_X1   g08142(.A1(new_n8334_), .A2(new_n8330_), .B(\asqrt[56] ), .ZN(new_n8335_));
  NAND2_X1   g08143(.A1(new_n8335_), .A2(new_n531_), .ZN(new_n8336_));
  OAI21_X1   g08144(.A1(new_n8336_), .A2(new_n8241_), .B(new_n8248_), .ZN(new_n8337_));
  AOI21_X1   g08145(.A1(new_n8337_), .A2(new_n8242_), .B(new_n436_), .ZN(new_n8338_));
  NOR2_X1    g08146(.A1(new_n7893_), .A2(new_n7883_), .ZN(new_n8339_));
  NOR3_X1    g08147(.A1(new_n8036_), .A2(new_n7860_), .A3(new_n8339_), .ZN(new_n8340_));
  INV_X1     g08148(.I(new_n8340_), .ZN(new_n8341_));
  NOR3_X1    g08149(.A1(new_n8339_), .A2(new_n7860_), .A3(new_n7892_), .ZN(new_n8342_));
  AOI22_X1   g08150(.A1(new_n8341_), .A2(new_n7892_), .B1(\asqrt[29] ), .B2(new_n8342_), .ZN(new_n8343_));
  NOR3_X1    g08151(.A1(new_n8334_), .A2(\asqrt[56] ), .A3(new_n8330_), .ZN(new_n8344_));
  OAI21_X1   g08152(.A1(new_n8238_), .A2(new_n8344_), .B(new_n8335_), .ZN(new_n8345_));
  AOI21_X1   g08153(.A1(new_n8345_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n8346_));
  AOI21_X1   g08154(.A1(new_n8346_), .A2(new_n8337_), .B(new_n8343_), .ZN(new_n8347_));
  OAI21_X1   g08155(.A1(new_n8347_), .A2(new_n8338_), .B(\asqrt[59] ), .ZN(new_n8348_));
  NOR3_X1    g08156(.A1(new_n7895_), .A2(new_n7929_), .A3(new_n7877_), .ZN(new_n8349_));
  NOR3_X1    g08157(.A1(new_n8036_), .A2(new_n7895_), .A3(new_n7929_), .ZN(new_n8350_));
  INV_X1     g08158(.I(new_n8350_), .ZN(new_n8351_));
  AOI22_X1   g08159(.A1(new_n8351_), .A2(new_n7877_), .B1(\asqrt[29] ), .B2(new_n8349_), .ZN(new_n8352_));
  INV_X1     g08160(.I(new_n8352_), .ZN(new_n8353_));
  INV_X1     g08161(.I(new_n8238_), .ZN(new_n8354_));
  NAND2_X1   g08162(.A1(new_n8225_), .A2(new_n703_), .ZN(new_n8355_));
  OAI21_X1   g08163(.A1(new_n8355_), .A2(new_n8334_), .B(new_n8354_), .ZN(new_n8356_));
  AOI21_X1   g08164(.A1(new_n8356_), .A2(new_n8335_), .B(new_n531_), .ZN(new_n8357_));
  NOR2_X1    g08165(.A1(new_n8234_), .A2(\asqrt[57] ), .ZN(new_n8358_));
  AOI21_X1   g08166(.A1(new_n8358_), .A2(new_n8356_), .B(new_n8247_), .ZN(new_n8359_));
  OAI21_X1   g08167(.A1(new_n8359_), .A2(new_n8357_), .B(\asqrt[58] ), .ZN(new_n8360_));
  NAND2_X1   g08168(.A1(new_n8360_), .A2(new_n327_), .ZN(new_n8361_));
  OAI21_X1   g08169(.A1(new_n8361_), .A2(new_n8347_), .B(new_n8353_), .ZN(new_n8362_));
  AOI21_X1   g08170(.A1(new_n8362_), .A2(new_n8348_), .B(new_n306_), .ZN(new_n8363_));
  NOR2_X1    g08171(.A1(new_n7918_), .A2(new_n7907_), .ZN(new_n8364_));
  NOR3_X1    g08172(.A1(new_n8036_), .A2(new_n7887_), .A3(new_n8364_), .ZN(new_n8365_));
  INV_X1     g08173(.I(new_n8365_), .ZN(new_n8366_));
  NOR3_X1    g08174(.A1(new_n7887_), .A2(new_n8364_), .A3(new_n7917_), .ZN(new_n8367_));
  AOI22_X1   g08175(.A1(new_n8366_), .A2(new_n7917_), .B1(\asqrt[29] ), .B2(new_n8367_), .ZN(new_n8368_));
  INV_X1     g08176(.I(new_n8343_), .ZN(new_n8369_));
  NAND2_X1   g08177(.A1(new_n8242_), .A2(new_n436_), .ZN(new_n8370_));
  OAI21_X1   g08178(.A1(new_n8370_), .A2(new_n8359_), .B(new_n8369_), .ZN(new_n8371_));
  AOI21_X1   g08179(.A1(new_n8371_), .A2(new_n8360_), .B(new_n327_), .ZN(new_n8372_));
  NOR2_X1    g08180(.A1(new_n8372_), .A2(\asqrt[60] ), .ZN(new_n8373_));
  AOI21_X1   g08181(.A1(new_n8373_), .A2(new_n8362_), .B(new_n8368_), .ZN(new_n8374_));
  OAI21_X1   g08182(.A1(new_n8374_), .A2(new_n8363_), .B(\asqrt[61] ), .ZN(new_n8375_));
  NOR2_X1    g08183(.A1(new_n7909_), .A2(new_n7897_), .ZN(new_n8376_));
  NOR3_X1    g08184(.A1(new_n8376_), .A2(new_n7920_), .A3(new_n7905_), .ZN(new_n8377_));
  NOR3_X1    g08185(.A1(new_n8036_), .A2(new_n7920_), .A3(new_n8376_), .ZN(new_n8378_));
  INV_X1     g08186(.I(new_n8378_), .ZN(new_n8379_));
  AOI22_X1   g08187(.A1(new_n8379_), .A2(new_n7905_), .B1(\asqrt[29] ), .B2(new_n8377_), .ZN(new_n8380_));
  INV_X1     g08188(.I(new_n8380_), .ZN(new_n8381_));
  NOR3_X1    g08189(.A1(new_n8241_), .A2(new_n8234_), .A3(\asqrt[57] ), .ZN(new_n8382_));
  OAI21_X1   g08190(.A1(new_n8247_), .A2(new_n8382_), .B(new_n8242_), .ZN(new_n8383_));
  AOI21_X1   g08191(.A1(new_n8383_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n8384_));
  AOI21_X1   g08192(.A1(new_n8384_), .A2(new_n8371_), .B(new_n8352_), .ZN(new_n8385_));
  OAI21_X1   g08193(.A1(new_n8385_), .A2(new_n8372_), .B(\asqrt[60] ), .ZN(new_n8386_));
  NAND2_X1   g08194(.A1(new_n8386_), .A2(new_n218_), .ZN(new_n8387_));
  OAI21_X1   g08195(.A1(new_n8387_), .A2(new_n8374_), .B(new_n8381_), .ZN(new_n8388_));
  AOI21_X1   g08196(.A1(new_n8388_), .A2(new_n8375_), .B(new_n207_), .ZN(new_n8389_));
  NOR3_X1    g08197(.A1(new_n8036_), .A2(new_n7911_), .A3(new_n7945_), .ZN(new_n8390_));
  INV_X1     g08198(.I(new_n8390_), .ZN(new_n8391_));
  NOR3_X1    g08199(.A1(new_n7911_), .A2(new_n7945_), .A3(new_n7973_), .ZN(new_n8392_));
  AOI22_X1   g08200(.A1(new_n8391_), .A2(new_n7973_), .B1(\asqrt[29] ), .B2(new_n8392_), .ZN(new_n8393_));
  NOR3_X1    g08201(.A1(new_n8385_), .A2(\asqrt[60] ), .A3(new_n8372_), .ZN(new_n8394_));
  OAI21_X1   g08202(.A1(new_n8368_), .A2(new_n8394_), .B(new_n8386_), .ZN(new_n8395_));
  AOI21_X1   g08203(.A1(new_n8395_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n8396_));
  AOI21_X1   g08204(.A1(new_n8396_), .A2(new_n8388_), .B(new_n8393_), .ZN(new_n8397_));
  AND3_X2    g08205(.A1(new_n7923_), .A2(new_n7976_), .A3(new_n7927_), .Z(new_n8398_));
  NAND2_X1   g08206(.A1(\asqrt[29] ), .A2(new_n8398_), .ZN(new_n8399_));
  INV_X1     g08207(.I(new_n8399_), .ZN(new_n8400_));
  AND2_X2    g08208(.A1(new_n7923_), .A2(new_n7976_), .Z(new_n8401_));
  AOI21_X1   g08209(.A1(\asqrt[29] ), .A2(new_n8401_), .B(new_n7927_), .ZN(new_n8402_));
  NOR2_X1    g08210(.A1(new_n8400_), .A2(new_n8402_), .ZN(new_n8403_));
  NOR3_X1    g08211(.A1(new_n8036_), .A2(new_n7977_), .A3(new_n7967_), .ZN(new_n8404_));
  NOR3_X1    g08212(.A1(new_n8403_), .A2(new_n7990_), .A3(new_n8404_), .ZN(new_n8405_));
  OAI21_X1   g08213(.A1(new_n8397_), .A2(new_n8389_), .B(new_n8405_), .ZN(new_n8406_));
  NAND2_X1   g08214(.A1(new_n8406_), .A2(new_n193_), .ZN(new_n8407_));
  INV_X1     g08215(.I(new_n8393_), .ZN(new_n8408_));
  NAND3_X1   g08216(.A1(new_n8388_), .A2(new_n207_), .A3(new_n8375_), .ZN(new_n8409_));
  NAND2_X1   g08217(.A1(new_n8409_), .A2(new_n8408_), .ZN(new_n8410_));
  INV_X1     g08218(.I(new_n8403_), .ZN(new_n8411_));
  NOR2_X1    g08219(.A1(new_n8389_), .A2(new_n8411_), .ZN(new_n8412_));
  AOI21_X1   g08220(.A1(\asqrt[29] ), .A2(new_n7940_), .B(new_n7963_), .ZN(new_n8413_));
  OAI21_X1   g08221(.A1(new_n7977_), .A2(new_n7967_), .B(\asqrt[63] ), .ZN(new_n8414_));
  NOR2_X1    g08222(.A1(new_n8413_), .A2(new_n8414_), .ZN(new_n8415_));
  INV_X1     g08223(.I(new_n7990_), .ZN(new_n8416_));
  AND3_X2    g08224(.A1(new_n7939_), .A2(new_n7937_), .A3(new_n7953_), .Z(new_n8417_));
  NAND4_X1   g08225(.A1(new_n8416_), .A2(new_n7978_), .A3(new_n7950_), .A4(new_n8417_), .ZN(new_n8418_));
  INV_X1     g08226(.I(new_n8418_), .ZN(new_n8419_));
  NOR2_X1    g08227(.A1(new_n8415_), .A2(new_n8419_), .ZN(new_n8420_));
  INV_X1     g08228(.I(new_n8420_), .ZN(new_n8421_));
  AOI21_X1   g08229(.A1(new_n8412_), .A2(new_n8410_), .B(new_n8421_), .ZN(new_n8422_));
  NAND2_X1   g08230(.A1(new_n8407_), .A2(new_n8422_), .ZN(\asqrt[28] ));
  NOR2_X1    g08231(.A1(\a[54] ), .A2(\a[55] ), .ZN(new_n8424_));
  INV_X1     g08232(.I(new_n8424_), .ZN(new_n8425_));
  NOR2_X1    g08233(.A1(new_n8425_), .A2(\a[56] ), .ZN(new_n8426_));
  INV_X1     g08234(.I(new_n8426_), .ZN(new_n8427_));
  INV_X1     g08235(.I(new_n8368_), .ZN(new_n8428_));
  NAND2_X1   g08236(.A1(new_n8348_), .A2(new_n306_), .ZN(new_n8429_));
  OAI21_X1   g08237(.A1(new_n8429_), .A2(new_n8385_), .B(new_n8428_), .ZN(new_n8430_));
  AOI21_X1   g08238(.A1(new_n8430_), .A2(new_n8386_), .B(new_n218_), .ZN(new_n8431_));
  NOR3_X1    g08239(.A1(new_n8347_), .A2(\asqrt[59] ), .A3(new_n8338_), .ZN(new_n8432_));
  OAI21_X1   g08240(.A1(new_n8352_), .A2(new_n8432_), .B(new_n8348_), .ZN(new_n8433_));
  AOI21_X1   g08241(.A1(new_n8433_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n8434_));
  AOI21_X1   g08242(.A1(new_n8434_), .A2(new_n8430_), .B(new_n8380_), .ZN(new_n8435_));
  OAI21_X1   g08243(.A1(new_n8435_), .A2(new_n8431_), .B(\asqrt[62] ), .ZN(new_n8436_));
  NOR3_X1    g08244(.A1(new_n8435_), .A2(\asqrt[62] ), .A3(new_n8431_), .ZN(new_n8437_));
  OAI21_X1   g08245(.A1(new_n8393_), .A2(new_n8437_), .B(new_n8436_), .ZN(new_n8438_));
  AOI21_X1   g08246(.A1(new_n8438_), .A2(new_n8405_), .B(\asqrt[63] ), .ZN(new_n8439_));
  NAND2_X1   g08247(.A1(new_n8436_), .A2(new_n8403_), .ZN(new_n8440_));
  OAI21_X1   g08248(.A1(new_n8440_), .A2(new_n8397_), .B(new_n8420_), .ZN(new_n8441_));
  OAI21_X1   g08249(.A1(new_n8439_), .A2(new_n8441_), .B(\a[56] ), .ZN(new_n8442_));
  AOI21_X1   g08250(.A1(new_n8442_), .A2(new_n8427_), .B(new_n8036_), .ZN(new_n8443_));
  INV_X1     g08251(.I(\a[56] ), .ZN(new_n8444_));
  AOI21_X1   g08252(.A1(new_n8407_), .A2(new_n8422_), .B(new_n8444_), .ZN(new_n8445_));
  NAND2_X1   g08253(.A1(new_n7953_), .A2(new_n8427_), .ZN(new_n8446_));
  NOR4_X1    g08254(.A1(new_n7965_), .A2(new_n7990_), .A3(new_n7951_), .A4(new_n8446_), .ZN(new_n8447_));
  INV_X1     g08255(.I(new_n8447_), .ZN(new_n8448_));
  NOR2_X1    g08256(.A1(new_n8445_), .A2(new_n8448_), .ZN(new_n8449_));
  AOI21_X1   g08257(.A1(new_n8407_), .A2(new_n8422_), .B(new_n7960_), .ZN(new_n8450_));
  INV_X1     g08258(.I(\a[57] ), .ZN(new_n8451_));
  AOI21_X1   g08259(.A1(\asqrt[28] ), .A2(new_n8444_), .B(new_n8451_), .ZN(new_n8452_));
  NOR3_X1    g08260(.A1(new_n8449_), .A2(new_n8452_), .A3(new_n8450_), .ZN(new_n8453_));
  OAI21_X1   g08261(.A1(new_n8453_), .A2(new_n8443_), .B(\asqrt[30] ), .ZN(new_n8454_));
  OAI21_X1   g08262(.A1(new_n8439_), .A2(new_n8441_), .B(new_n7959_), .ZN(new_n8455_));
  NAND2_X1   g08263(.A1(new_n8412_), .A2(new_n8410_), .ZN(new_n8456_));
  INV_X1     g08264(.I(new_n8415_), .ZN(new_n8457_));
  NOR2_X1    g08265(.A1(new_n8419_), .A2(new_n8036_), .ZN(new_n8458_));
  NAND4_X1   g08266(.A1(new_n8407_), .A2(new_n8456_), .A3(new_n8457_), .A4(new_n8458_), .ZN(new_n8459_));
  AOI21_X1   g08267(.A1(new_n8459_), .A2(new_n8455_), .B(new_n7972_), .ZN(new_n8460_));
  INV_X1     g08268(.I(new_n8456_), .ZN(new_n8461_));
  NAND2_X1   g08269(.A1(new_n8457_), .A2(new_n8458_), .ZN(new_n8462_));
  NOR3_X1    g08270(.A1(new_n8461_), .A2(new_n8439_), .A3(new_n8462_), .ZN(new_n8463_));
  NOR3_X1    g08271(.A1(new_n8463_), .A2(new_n8450_), .A3(\a[58] ), .ZN(new_n8464_));
  OAI21_X1   g08272(.A1(new_n8445_), .A2(new_n8426_), .B(\asqrt[29] ), .ZN(new_n8465_));
  NAND2_X1   g08273(.A1(new_n8465_), .A2(new_n7539_), .ZN(new_n8466_));
  OAI22_X1   g08274(.A1(new_n8453_), .A2(new_n8466_), .B1(new_n8460_), .B2(new_n8464_), .ZN(new_n8467_));
  AOI21_X1   g08275(.A1(new_n8467_), .A2(new_n8454_), .B(new_n7229_), .ZN(new_n8468_));
  NOR3_X1    g08276(.A1(new_n8271_), .A2(new_n7971_), .A3(new_n7983_), .ZN(new_n8469_));
  NAND3_X1   g08277(.A1(\asqrt[28] ), .A2(new_n8006_), .A3(new_n8256_), .ZN(new_n8470_));
  AOI22_X1   g08278(.A1(new_n8470_), .A2(new_n8271_), .B1(\asqrt[28] ), .B2(new_n8469_), .ZN(new_n8471_));
  AOI21_X1   g08279(.A1(new_n8407_), .A2(new_n8422_), .B(\a[56] ), .ZN(new_n8472_));
  OAI21_X1   g08280(.A1(new_n8451_), .A2(new_n8472_), .B(new_n8455_), .ZN(new_n8473_));
  OAI21_X1   g08281(.A1(new_n8473_), .A2(new_n8449_), .B(new_n8465_), .ZN(new_n8474_));
  AOI21_X1   g08282(.A1(new_n8474_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n8475_));
  AOI21_X1   g08283(.A1(new_n8475_), .A2(new_n8467_), .B(new_n8471_), .ZN(new_n8476_));
  OAI21_X1   g08284(.A1(new_n8476_), .A2(new_n8468_), .B(\asqrt[32] ), .ZN(new_n8477_));
  INV_X1     g08285(.I(new_n8477_), .ZN(new_n8478_));
  NOR2_X1    g08286(.A1(new_n7995_), .A2(new_n7996_), .ZN(new_n8479_));
  NOR2_X1    g08287(.A1(new_n7987_), .A2(new_n7998_), .ZN(new_n8480_));
  INV_X1     g08288(.I(new_n8480_), .ZN(new_n8481_));
  NAND4_X1   g08289(.A1(\asqrt[28] ), .A2(new_n7988_), .A3(new_n8479_), .A4(new_n8481_), .ZN(new_n8482_));
  INV_X1     g08290(.I(\asqrt[28] ), .ZN(new_n8483_));
  NOR3_X1    g08291(.A1(new_n8483_), .A2(new_n8260_), .A3(new_n8480_), .ZN(new_n8484_));
  OAI21_X1   g08292(.A1(new_n8484_), .A2(new_n8479_), .B(new_n8482_), .ZN(new_n8485_));
  INV_X1     g08293(.I(new_n8485_), .ZN(new_n8486_));
  NOR3_X1    g08294(.A1(new_n8476_), .A2(new_n8468_), .A3(\asqrt[32] ), .ZN(new_n8487_));
  NOR2_X1    g08295(.A1(new_n8487_), .A2(new_n8486_), .ZN(new_n8488_));
  OAI21_X1   g08296(.A1(new_n8488_), .A2(new_n8478_), .B(\asqrt[33] ), .ZN(new_n8489_));
  NOR2_X1    g08297(.A1(new_n8273_), .A2(new_n8265_), .ZN(new_n8490_));
  NOR3_X1    g08298(.A1(new_n8483_), .A2(new_n8000_), .A3(new_n8490_), .ZN(new_n8491_));
  INV_X1     g08299(.I(new_n8491_), .ZN(new_n8492_));
  NOR3_X1    g08300(.A1(new_n8490_), .A2(new_n8000_), .A3(new_n8270_), .ZN(new_n8493_));
  AOI22_X1   g08301(.A1(new_n8492_), .A2(new_n8270_), .B1(\asqrt[28] ), .B2(new_n8493_), .ZN(new_n8494_));
  INV_X1     g08302(.I(new_n8494_), .ZN(new_n8495_));
  NAND2_X1   g08303(.A1(new_n8477_), .A2(new_n6356_), .ZN(new_n8496_));
  OAI21_X1   g08304(.A1(new_n8488_), .A2(new_n8496_), .B(new_n8495_), .ZN(new_n8497_));
  AOI21_X1   g08305(.A1(new_n8497_), .A2(new_n8489_), .B(new_n6077_), .ZN(new_n8498_));
  NOR3_X1    g08306(.A1(new_n8013_), .A2(new_n8021_), .A3(new_n8019_), .ZN(new_n8499_));
  NOR3_X1    g08307(.A1(new_n8483_), .A2(new_n8013_), .A3(new_n8021_), .ZN(new_n8500_));
  INV_X1     g08308(.I(new_n8500_), .ZN(new_n8501_));
  AOI22_X1   g08309(.A1(new_n8501_), .A2(new_n8019_), .B1(\asqrt[28] ), .B2(new_n8499_), .ZN(new_n8502_));
  OAI21_X1   g08310(.A1(new_n8486_), .A2(new_n8487_), .B(new_n8477_), .ZN(new_n8503_));
  AOI21_X1   g08311(.A1(new_n8503_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n8504_));
  AOI21_X1   g08312(.A1(new_n8504_), .A2(new_n8497_), .B(new_n8502_), .ZN(new_n8505_));
  OAI21_X1   g08313(.A1(new_n8505_), .A2(new_n8498_), .B(\asqrt[35] ), .ZN(new_n8506_));
  INV_X1     g08314(.I(new_n8506_), .ZN(new_n8507_));
  NAND2_X1   g08315(.A1(new_n8276_), .A2(new_n8268_), .ZN(new_n8508_));
  NAND3_X1   g08316(.A1(\asqrt[28] ), .A2(new_n8023_), .A3(new_n8508_), .ZN(new_n8509_));
  AND3_X2    g08317(.A1(new_n8023_), .A2(new_n8029_), .A3(new_n8508_), .Z(new_n8510_));
  AOI22_X1   g08318(.A1(new_n8509_), .A2(new_n8030_), .B1(\asqrt[28] ), .B2(new_n8510_), .ZN(new_n8511_));
  NOR3_X1    g08319(.A1(new_n8505_), .A2(new_n8498_), .A3(\asqrt[35] ), .ZN(new_n8512_));
  NOR2_X1    g08320(.A1(new_n8512_), .A2(new_n8511_), .ZN(new_n8513_));
  OAI21_X1   g08321(.A1(new_n8513_), .A2(new_n8507_), .B(\asqrt[36] ), .ZN(new_n8514_));
  INV_X1     g08322(.I(new_n8039_), .ZN(new_n8515_));
  NOR3_X1    g08323(.A1(new_n8033_), .A2(new_n8287_), .A3(new_n8515_), .ZN(new_n8516_));
  NOR3_X1    g08324(.A1(new_n8483_), .A2(new_n8033_), .A3(new_n8287_), .ZN(new_n8517_));
  INV_X1     g08325(.I(new_n8517_), .ZN(new_n8518_));
  AOI22_X1   g08326(.A1(new_n8518_), .A2(new_n8515_), .B1(\asqrt[28] ), .B2(new_n8516_), .ZN(new_n8519_));
  INV_X1     g08327(.I(new_n8519_), .ZN(new_n8520_));
  NAND2_X1   g08328(.A1(new_n8506_), .A2(new_n5277_), .ZN(new_n8521_));
  OAI21_X1   g08329(.A1(new_n8513_), .A2(new_n8521_), .B(new_n8520_), .ZN(new_n8522_));
  AOI21_X1   g08330(.A1(new_n8522_), .A2(new_n8514_), .B(new_n5024_), .ZN(new_n8523_));
  NOR3_X1    g08331(.A1(new_n8483_), .A2(new_n8044_), .A3(new_n8051_), .ZN(new_n8524_));
  INV_X1     g08332(.I(new_n8524_), .ZN(new_n8525_));
  NOR3_X1    g08333(.A1(new_n8044_), .A2(new_n8255_), .A3(new_n8051_), .ZN(new_n8526_));
  AOI22_X1   g08334(.A1(new_n8525_), .A2(new_n8255_), .B1(\asqrt[28] ), .B2(new_n8526_), .ZN(new_n8527_));
  INV_X1     g08335(.I(new_n8511_), .ZN(new_n8528_));
  NAND2_X1   g08336(.A1(new_n8442_), .A2(new_n8447_), .ZN(new_n8529_));
  OAI21_X1   g08337(.A1(new_n8439_), .A2(new_n8441_), .B(new_n8444_), .ZN(new_n8530_));
  NAND2_X1   g08338(.A1(new_n8530_), .A2(\a[57] ), .ZN(new_n8531_));
  NAND3_X1   g08339(.A1(new_n8529_), .A2(new_n8531_), .A3(new_n8455_), .ZN(new_n8532_));
  AOI21_X1   g08340(.A1(new_n8532_), .A2(new_n8465_), .B(new_n7539_), .ZN(new_n8533_));
  OAI21_X1   g08341(.A1(new_n8463_), .A2(new_n8450_), .B(\a[58] ), .ZN(new_n8534_));
  NAND3_X1   g08342(.A1(new_n8459_), .A2(new_n8455_), .A3(new_n7972_), .ZN(new_n8535_));
  NAND2_X1   g08343(.A1(new_n8442_), .A2(new_n8427_), .ZN(new_n8536_));
  AOI21_X1   g08344(.A1(new_n8536_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n8537_));
  AOI22_X1   g08345(.A1(new_n8532_), .A2(new_n8537_), .B1(new_n8534_), .B2(new_n8535_), .ZN(new_n8538_));
  OAI21_X1   g08346(.A1(new_n8538_), .A2(new_n8533_), .B(\asqrt[31] ), .ZN(new_n8539_));
  NAND2_X1   g08347(.A1(new_n8539_), .A2(new_n6824_), .ZN(new_n8540_));
  OAI21_X1   g08348(.A1(new_n8540_), .A2(new_n8476_), .B(new_n8485_), .ZN(new_n8541_));
  AOI21_X1   g08349(.A1(new_n8541_), .A2(new_n8477_), .B(new_n6356_), .ZN(new_n8542_));
  INV_X1     g08350(.I(new_n8471_), .ZN(new_n8543_));
  AOI21_X1   g08351(.A1(\a[57] ), .A2(new_n8530_), .B(new_n8450_), .ZN(new_n8544_));
  AOI21_X1   g08352(.A1(new_n8544_), .A2(new_n8529_), .B(new_n8443_), .ZN(new_n8545_));
  OAI21_X1   g08353(.A1(new_n8545_), .A2(new_n7539_), .B(new_n7229_), .ZN(new_n8546_));
  OAI21_X1   g08354(.A1(new_n8546_), .A2(new_n8538_), .B(new_n8543_), .ZN(new_n8547_));
  NAND2_X1   g08355(.A1(new_n8547_), .A2(new_n8539_), .ZN(new_n8548_));
  AOI21_X1   g08356(.A1(new_n8548_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n8549_));
  AOI21_X1   g08357(.A1(new_n8549_), .A2(new_n8541_), .B(new_n8494_), .ZN(new_n8550_));
  OAI21_X1   g08358(.A1(new_n8550_), .A2(new_n8542_), .B(\asqrt[34] ), .ZN(new_n8551_));
  NAND2_X1   g08359(.A1(new_n8551_), .A2(new_n5708_), .ZN(new_n8552_));
  OAI21_X1   g08360(.A1(new_n8552_), .A2(new_n8505_), .B(new_n8528_), .ZN(new_n8553_));
  AOI21_X1   g08361(.A1(new_n8553_), .A2(new_n8506_), .B(new_n5277_), .ZN(new_n8554_));
  NOR2_X1    g08362(.A1(new_n8554_), .A2(\asqrt[37] ), .ZN(new_n8555_));
  AOI21_X1   g08363(.A1(new_n8555_), .A2(new_n8522_), .B(new_n8527_), .ZN(new_n8556_));
  OAI21_X1   g08364(.A1(new_n8556_), .A2(new_n8523_), .B(\asqrt[38] ), .ZN(new_n8557_));
  INV_X1     g08365(.I(new_n8557_), .ZN(new_n8558_));
  INV_X1     g08366(.I(new_n8281_), .ZN(new_n8559_));
  NOR3_X1    g08367(.A1(new_n8559_), .A2(new_n8286_), .A3(new_n8062_), .ZN(new_n8560_));
  NOR3_X1    g08368(.A1(new_n8483_), .A2(new_n8286_), .A3(new_n8559_), .ZN(new_n8561_));
  INV_X1     g08369(.I(new_n8561_), .ZN(new_n8562_));
  AOI22_X1   g08370(.A1(new_n8562_), .A2(new_n8062_), .B1(\asqrt[28] ), .B2(new_n8560_), .ZN(new_n8563_));
  NOR3_X1    g08371(.A1(new_n8556_), .A2(\asqrt[38] ), .A3(new_n8523_), .ZN(new_n8564_));
  NOR2_X1    g08372(.A1(new_n8564_), .A2(new_n8563_), .ZN(new_n8565_));
  OAI21_X1   g08373(.A1(new_n8565_), .A2(new_n8558_), .B(\asqrt[39] ), .ZN(new_n8566_));
  INV_X1     g08374(.I(new_n8070_), .ZN(new_n8567_));
  NOR3_X1    g08375(.A1(new_n8483_), .A2(new_n8065_), .A3(new_n8291_), .ZN(new_n8568_));
  INV_X1     g08376(.I(new_n8568_), .ZN(new_n8569_));
  NOR3_X1    g08377(.A1(new_n8065_), .A2(new_n8291_), .A3(new_n8567_), .ZN(new_n8570_));
  AOI22_X1   g08378(.A1(new_n8569_), .A2(new_n8567_), .B1(\asqrt[28] ), .B2(new_n8570_), .ZN(new_n8571_));
  INV_X1     g08379(.I(new_n8571_), .ZN(new_n8572_));
  NAND2_X1   g08380(.A1(new_n8557_), .A2(new_n4298_), .ZN(new_n8573_));
  OAI21_X1   g08381(.A1(new_n8565_), .A2(new_n8573_), .B(new_n8572_), .ZN(new_n8574_));
  AOI21_X1   g08382(.A1(new_n8574_), .A2(new_n8566_), .B(new_n4071_), .ZN(new_n8575_));
  NOR3_X1    g08383(.A1(new_n8075_), .A2(new_n8254_), .A3(new_n8081_), .ZN(new_n8576_));
  NOR3_X1    g08384(.A1(new_n8483_), .A2(new_n8075_), .A3(new_n8081_), .ZN(new_n8577_));
  INV_X1     g08385(.I(new_n8577_), .ZN(new_n8578_));
  AOI22_X1   g08386(.A1(new_n8578_), .A2(new_n8254_), .B1(\asqrt[28] ), .B2(new_n8576_), .ZN(new_n8579_));
  INV_X1     g08387(.I(new_n8563_), .ZN(new_n8580_));
  OAI21_X1   g08388(.A1(new_n8511_), .A2(new_n8512_), .B(new_n8506_), .ZN(new_n8581_));
  NAND3_X1   g08389(.A1(new_n8553_), .A2(new_n5277_), .A3(new_n8506_), .ZN(new_n8582_));
  AOI22_X1   g08390(.A1(new_n8582_), .A2(new_n8520_), .B1(new_n8581_), .B2(\asqrt[36] ), .ZN(new_n8583_));
  OAI21_X1   g08391(.A1(new_n8583_), .A2(new_n5024_), .B(new_n4696_), .ZN(new_n8584_));
  OAI21_X1   g08392(.A1(new_n8584_), .A2(new_n8556_), .B(new_n8580_), .ZN(new_n8585_));
  AOI21_X1   g08393(.A1(new_n8585_), .A2(new_n8557_), .B(new_n4298_), .ZN(new_n8586_));
  NOR2_X1    g08394(.A1(new_n8586_), .A2(\asqrt[40] ), .ZN(new_n8587_));
  AOI21_X1   g08395(.A1(new_n8587_), .A2(new_n8574_), .B(new_n8579_), .ZN(new_n8588_));
  OAI21_X1   g08396(.A1(new_n8588_), .A2(new_n8575_), .B(\asqrt[41] ), .ZN(new_n8589_));
  NOR2_X1    g08397(.A1(new_n8082_), .A2(new_n8093_), .ZN(new_n8590_));
  NOR3_X1    g08398(.A1(new_n8483_), .A2(new_n8285_), .A3(new_n8590_), .ZN(new_n8591_));
  INV_X1     g08399(.I(new_n8591_), .ZN(new_n8592_));
  NOR3_X1    g08400(.A1(new_n8590_), .A2(new_n8285_), .A3(new_n8092_), .ZN(new_n8593_));
  AOI22_X1   g08401(.A1(new_n8592_), .A2(new_n8092_), .B1(\asqrt[28] ), .B2(new_n8593_), .ZN(new_n8594_));
  INV_X1     g08402(.I(new_n8594_), .ZN(new_n8595_));
  NOR3_X1    g08403(.A1(new_n8550_), .A2(new_n8542_), .A3(\asqrt[34] ), .ZN(new_n8596_));
  OAI21_X1   g08404(.A1(new_n8502_), .A2(new_n8596_), .B(new_n8551_), .ZN(new_n8597_));
  AOI21_X1   g08405(.A1(new_n8597_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n8598_));
  AOI21_X1   g08406(.A1(new_n8598_), .A2(new_n8553_), .B(new_n8519_), .ZN(new_n8599_));
  NOR3_X1    g08407(.A1(new_n8599_), .A2(\asqrt[37] ), .A3(new_n8554_), .ZN(new_n8600_));
  OAI22_X1   g08408(.A1(new_n8600_), .A2(new_n8527_), .B1(new_n8583_), .B2(new_n5024_), .ZN(new_n8601_));
  AOI21_X1   g08409(.A1(new_n8601_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n8602_));
  AOI21_X1   g08410(.A1(new_n8602_), .A2(new_n8585_), .B(new_n8571_), .ZN(new_n8603_));
  OAI21_X1   g08411(.A1(new_n8603_), .A2(new_n8586_), .B(\asqrt[40] ), .ZN(new_n8604_));
  NAND2_X1   g08412(.A1(new_n8604_), .A2(new_n3782_), .ZN(new_n8605_));
  OAI21_X1   g08413(.A1(new_n8605_), .A2(new_n8588_), .B(new_n8595_), .ZN(new_n8606_));
  AOI21_X1   g08414(.A1(new_n8606_), .A2(new_n8589_), .B(new_n3419_), .ZN(new_n8607_));
  INV_X1     g08415(.I(new_n8100_), .ZN(new_n8608_));
  NOR3_X1    g08416(.A1(new_n8095_), .A2(new_n8299_), .A3(new_n8608_), .ZN(new_n8609_));
  NOR3_X1    g08417(.A1(new_n8483_), .A2(new_n8095_), .A3(new_n8299_), .ZN(new_n8610_));
  INV_X1     g08418(.I(new_n8610_), .ZN(new_n8611_));
  AOI22_X1   g08419(.A1(new_n8611_), .A2(new_n8608_), .B1(\asqrt[28] ), .B2(new_n8609_), .ZN(new_n8612_));
  NOR3_X1    g08420(.A1(new_n8603_), .A2(\asqrt[40] ), .A3(new_n8586_), .ZN(new_n8613_));
  OAI21_X1   g08421(.A1(new_n8579_), .A2(new_n8613_), .B(new_n8604_), .ZN(new_n8614_));
  AOI21_X1   g08422(.A1(new_n8614_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n8615_));
  AOI21_X1   g08423(.A1(new_n8615_), .A2(new_n8606_), .B(new_n8612_), .ZN(new_n8616_));
  OAI21_X1   g08424(.A1(new_n8616_), .A2(new_n8607_), .B(\asqrt[43] ), .ZN(new_n8617_));
  INV_X1     g08425(.I(new_n8617_), .ZN(new_n8618_));
  NOR3_X1    g08426(.A1(new_n8483_), .A2(new_n8105_), .A3(new_n8112_), .ZN(new_n8619_));
  INV_X1     g08427(.I(new_n8619_), .ZN(new_n8620_));
  NOR3_X1    g08428(.A1(new_n8105_), .A2(new_n8253_), .A3(new_n8112_), .ZN(new_n8621_));
  AOI22_X1   g08429(.A1(new_n8620_), .A2(new_n8253_), .B1(\asqrt[28] ), .B2(new_n8621_), .ZN(new_n8622_));
  NOR3_X1    g08430(.A1(new_n8616_), .A2(\asqrt[43] ), .A3(new_n8607_), .ZN(new_n8623_));
  NOR2_X1    g08431(.A1(new_n8623_), .A2(new_n8622_), .ZN(new_n8624_));
  OAI21_X1   g08432(.A1(new_n8624_), .A2(new_n8618_), .B(\asqrt[44] ), .ZN(new_n8625_));
  NOR2_X1    g08433(.A1(new_n8113_), .A2(new_n8124_), .ZN(new_n8626_));
  NOR3_X1    g08434(.A1(new_n8626_), .A2(new_n8298_), .A3(new_n8123_), .ZN(new_n8627_));
  NOR3_X1    g08435(.A1(new_n8483_), .A2(new_n8298_), .A3(new_n8626_), .ZN(new_n8628_));
  INV_X1     g08436(.I(new_n8628_), .ZN(new_n8629_));
  AOI22_X1   g08437(.A1(new_n8629_), .A2(new_n8123_), .B1(\asqrt[28] ), .B2(new_n8627_), .ZN(new_n8630_));
  INV_X1     g08438(.I(new_n8630_), .ZN(new_n8631_));
  NAND2_X1   g08439(.A1(new_n8617_), .A2(new_n2954_), .ZN(new_n8632_));
  OAI21_X1   g08440(.A1(new_n8624_), .A2(new_n8632_), .B(new_n8631_), .ZN(new_n8633_));
  AOI21_X1   g08441(.A1(new_n8633_), .A2(new_n8625_), .B(new_n2641_), .ZN(new_n8634_));
  INV_X1     g08442(.I(new_n8131_), .ZN(new_n8635_));
  NOR3_X1    g08443(.A1(new_n8483_), .A2(new_n8126_), .A3(new_n8307_), .ZN(new_n8636_));
  INV_X1     g08444(.I(new_n8636_), .ZN(new_n8637_));
  NOR3_X1    g08445(.A1(new_n8126_), .A2(new_n8307_), .A3(new_n8635_), .ZN(new_n8638_));
  AOI22_X1   g08446(.A1(new_n8637_), .A2(new_n8635_), .B1(\asqrt[28] ), .B2(new_n8638_), .ZN(new_n8639_));
  OAI21_X1   g08447(.A1(new_n8622_), .A2(new_n8623_), .B(new_n8617_), .ZN(new_n8640_));
  AOI21_X1   g08448(.A1(new_n8640_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n8641_));
  AOI21_X1   g08449(.A1(new_n8641_), .A2(new_n8633_), .B(new_n8639_), .ZN(new_n8642_));
  OAI21_X1   g08450(.A1(new_n8642_), .A2(new_n8634_), .B(\asqrt[46] ), .ZN(new_n8643_));
  INV_X1     g08451(.I(new_n8643_), .ZN(new_n8644_));
  NOR3_X1    g08452(.A1(new_n8136_), .A2(new_n8252_), .A3(new_n8142_), .ZN(new_n8645_));
  NOR3_X1    g08453(.A1(new_n8483_), .A2(new_n8136_), .A3(new_n8142_), .ZN(new_n8646_));
  INV_X1     g08454(.I(new_n8646_), .ZN(new_n8647_));
  AOI22_X1   g08455(.A1(new_n8647_), .A2(new_n8252_), .B1(\asqrt[28] ), .B2(new_n8645_), .ZN(new_n8648_));
  NOR3_X1    g08456(.A1(new_n8642_), .A2(new_n8634_), .A3(\asqrt[46] ), .ZN(new_n8649_));
  NOR2_X1    g08457(.A1(new_n8649_), .A2(new_n8648_), .ZN(new_n8650_));
  OAI21_X1   g08458(.A1(new_n8650_), .A2(new_n8644_), .B(\asqrt[47] ), .ZN(new_n8651_));
  NOR2_X1    g08459(.A1(new_n8143_), .A2(new_n8152_), .ZN(new_n8652_));
  NOR3_X1    g08460(.A1(new_n8483_), .A2(new_n8306_), .A3(new_n8652_), .ZN(new_n8653_));
  INV_X1     g08461(.I(new_n8653_), .ZN(new_n8654_));
  NOR3_X1    g08462(.A1(new_n8652_), .A2(new_n8306_), .A3(new_n8151_), .ZN(new_n8655_));
  AOI22_X1   g08463(.A1(new_n8654_), .A2(new_n8151_), .B1(\asqrt[28] ), .B2(new_n8655_), .ZN(new_n8656_));
  INV_X1     g08464(.I(new_n8656_), .ZN(new_n8657_));
  NAND2_X1   g08465(.A1(new_n8643_), .A2(new_n2229_), .ZN(new_n8658_));
  OAI21_X1   g08466(.A1(new_n8650_), .A2(new_n8658_), .B(new_n8657_), .ZN(new_n8659_));
  AOI21_X1   g08467(.A1(new_n8659_), .A2(new_n8651_), .B(new_n1956_), .ZN(new_n8660_));
  INV_X1     g08468(.I(new_n8159_), .ZN(new_n8661_));
  NOR3_X1    g08469(.A1(new_n8154_), .A2(new_n8315_), .A3(new_n8661_), .ZN(new_n8662_));
  NOR3_X1    g08470(.A1(new_n8483_), .A2(new_n8154_), .A3(new_n8315_), .ZN(new_n8663_));
  INV_X1     g08471(.I(new_n8663_), .ZN(new_n8664_));
  AOI22_X1   g08472(.A1(new_n8664_), .A2(new_n8661_), .B1(\asqrt[28] ), .B2(new_n8662_), .ZN(new_n8665_));
  OAI21_X1   g08473(.A1(new_n8648_), .A2(new_n8649_), .B(new_n8643_), .ZN(new_n8666_));
  AOI21_X1   g08474(.A1(new_n8666_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n8667_));
  AOI21_X1   g08475(.A1(new_n8667_), .A2(new_n8659_), .B(new_n8665_), .ZN(new_n8668_));
  OAI21_X1   g08476(.A1(new_n8668_), .A2(new_n8660_), .B(\asqrt[49] ), .ZN(new_n8669_));
  INV_X1     g08477(.I(new_n8669_), .ZN(new_n8670_));
  NOR3_X1    g08478(.A1(new_n8483_), .A2(new_n8164_), .A3(new_n8171_), .ZN(new_n8671_));
  INV_X1     g08479(.I(new_n8671_), .ZN(new_n8672_));
  NOR3_X1    g08480(.A1(new_n8164_), .A2(new_n8251_), .A3(new_n8171_), .ZN(new_n8673_));
  AOI22_X1   g08481(.A1(new_n8672_), .A2(new_n8251_), .B1(\asqrt[28] ), .B2(new_n8673_), .ZN(new_n8674_));
  NOR3_X1    g08482(.A1(new_n8668_), .A2(new_n8660_), .A3(\asqrt[49] ), .ZN(new_n8675_));
  NOR2_X1    g08483(.A1(new_n8675_), .A2(new_n8674_), .ZN(new_n8676_));
  OAI21_X1   g08484(.A1(new_n8676_), .A2(new_n8670_), .B(\asqrt[50] ), .ZN(new_n8677_));
  NOR2_X1    g08485(.A1(new_n8172_), .A2(new_n8180_), .ZN(new_n8678_));
  NOR3_X1    g08486(.A1(new_n8678_), .A2(new_n8314_), .A3(new_n8179_), .ZN(new_n8679_));
  NOR3_X1    g08487(.A1(new_n8483_), .A2(new_n8314_), .A3(new_n8678_), .ZN(new_n8680_));
  INV_X1     g08488(.I(new_n8680_), .ZN(new_n8681_));
  AOI22_X1   g08489(.A1(new_n8681_), .A2(new_n8179_), .B1(\asqrt[28] ), .B2(new_n8679_), .ZN(new_n8682_));
  INV_X1     g08490(.I(new_n8682_), .ZN(new_n8683_));
  NAND2_X1   g08491(.A1(new_n8669_), .A2(new_n1612_), .ZN(new_n8684_));
  OAI21_X1   g08492(.A1(new_n8676_), .A2(new_n8684_), .B(new_n8683_), .ZN(new_n8685_));
  AOI21_X1   g08493(.A1(new_n8685_), .A2(new_n8677_), .B(new_n1376_), .ZN(new_n8686_));
  INV_X1     g08494(.I(new_n8186_), .ZN(new_n8687_));
  NOR3_X1    g08495(.A1(new_n8483_), .A2(new_n8182_), .A3(new_n8323_), .ZN(new_n8688_));
  INV_X1     g08496(.I(new_n8688_), .ZN(new_n8689_));
  NOR3_X1    g08497(.A1(new_n8182_), .A2(new_n8323_), .A3(new_n8687_), .ZN(new_n8690_));
  AOI22_X1   g08498(.A1(new_n8689_), .A2(new_n8687_), .B1(\asqrt[28] ), .B2(new_n8690_), .ZN(new_n8691_));
  OAI21_X1   g08499(.A1(new_n8674_), .A2(new_n8675_), .B(new_n8669_), .ZN(new_n8692_));
  AOI21_X1   g08500(.A1(new_n8692_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n8693_));
  AOI21_X1   g08501(.A1(new_n8693_), .A2(new_n8685_), .B(new_n8691_), .ZN(new_n8694_));
  OAI21_X1   g08502(.A1(new_n8694_), .A2(new_n8686_), .B(\asqrt[52] ), .ZN(new_n8695_));
  INV_X1     g08503(.I(new_n8695_), .ZN(new_n8696_));
  INV_X1     g08504(.I(new_n8694_), .ZN(new_n8697_));
  NOR3_X1    g08505(.A1(new_n8191_), .A2(new_n8250_), .A3(new_n8197_), .ZN(new_n8698_));
  NOR3_X1    g08506(.A1(new_n8483_), .A2(new_n8191_), .A3(new_n8197_), .ZN(new_n8699_));
  INV_X1     g08507(.I(new_n8699_), .ZN(new_n8700_));
  AOI22_X1   g08508(.A1(new_n8700_), .A2(new_n8250_), .B1(\asqrt[28] ), .B2(new_n8698_), .ZN(new_n8701_));
  NOR2_X1    g08509(.A1(new_n8686_), .A2(\asqrt[52] ), .ZN(new_n8702_));
  AOI21_X1   g08510(.A1(new_n8697_), .A2(new_n8702_), .B(new_n8701_), .ZN(new_n8703_));
  OAI21_X1   g08511(.A1(new_n8703_), .A2(new_n8696_), .B(\asqrt[53] ), .ZN(new_n8704_));
  NOR2_X1    g08512(.A1(new_n8198_), .A2(new_n8206_), .ZN(new_n8705_));
  NOR3_X1    g08513(.A1(new_n8483_), .A2(new_n8322_), .A3(new_n8705_), .ZN(new_n8706_));
  INV_X1     g08514(.I(new_n8706_), .ZN(new_n8707_));
  NOR3_X1    g08515(.A1(new_n8705_), .A2(new_n8322_), .A3(new_n8205_), .ZN(new_n8708_));
  AOI22_X1   g08516(.A1(new_n8707_), .A2(new_n8205_), .B1(\asqrt[28] ), .B2(new_n8708_), .ZN(new_n8709_));
  INV_X1     g08517(.I(new_n8709_), .ZN(new_n8710_));
  NAND2_X1   g08518(.A1(new_n8695_), .A2(new_n1103_), .ZN(new_n8711_));
  OAI21_X1   g08519(.A1(new_n8711_), .A2(new_n8703_), .B(new_n8710_), .ZN(new_n8712_));
  AOI21_X1   g08520(.A1(new_n8712_), .A2(new_n8704_), .B(new_n904_), .ZN(new_n8713_));
  INV_X1     g08521(.I(new_n8713_), .ZN(new_n8714_));
  INV_X1     g08522(.I(new_n8712_), .ZN(new_n8715_));
  INV_X1     g08523(.I(new_n8212_), .ZN(new_n8716_));
  NOR3_X1    g08524(.A1(new_n8208_), .A2(new_n8331_), .A3(new_n8716_), .ZN(new_n8717_));
  NOR3_X1    g08525(.A1(new_n8483_), .A2(new_n8208_), .A3(new_n8331_), .ZN(new_n8718_));
  INV_X1     g08526(.I(new_n8718_), .ZN(new_n8719_));
  AOI22_X1   g08527(.A1(new_n8719_), .A2(new_n8716_), .B1(\asqrt[28] ), .B2(new_n8717_), .ZN(new_n8720_));
  INV_X1     g08528(.I(new_n8720_), .ZN(new_n8721_));
  NAND2_X1   g08529(.A1(new_n8704_), .A2(new_n904_), .ZN(new_n8722_));
  OAI21_X1   g08530(.A1(new_n8722_), .A2(new_n8715_), .B(new_n8721_), .ZN(new_n8723_));
  AOI21_X1   g08531(.A1(new_n8723_), .A2(new_n8714_), .B(new_n823_), .ZN(new_n8724_));
  NOR3_X1    g08532(.A1(new_n8483_), .A2(new_n8217_), .A3(new_n8223_), .ZN(new_n8725_));
  INV_X1     g08533(.I(new_n8725_), .ZN(new_n8726_));
  NOR3_X1    g08534(.A1(new_n8217_), .A2(new_n8223_), .A3(new_n8249_), .ZN(new_n8727_));
  AOI22_X1   g08535(.A1(new_n8726_), .A2(new_n8249_), .B1(\asqrt[28] ), .B2(new_n8727_), .ZN(new_n8728_));
  NOR2_X1    g08536(.A1(new_n8713_), .A2(\asqrt[55] ), .ZN(new_n8729_));
  AOI21_X1   g08537(.A1(new_n8729_), .A2(new_n8723_), .B(new_n8728_), .ZN(new_n8730_));
  OAI21_X1   g08538(.A1(new_n8730_), .A2(new_n8724_), .B(\asqrt[56] ), .ZN(new_n8731_));
  NOR2_X1    g08539(.A1(new_n8224_), .A2(new_n8232_), .ZN(new_n8732_));
  NOR3_X1    g08540(.A1(new_n8732_), .A2(new_n8330_), .A3(new_n8231_), .ZN(new_n8733_));
  NOR3_X1    g08541(.A1(new_n8483_), .A2(new_n8330_), .A3(new_n8732_), .ZN(new_n8734_));
  INV_X1     g08542(.I(new_n8734_), .ZN(new_n8735_));
  AOI22_X1   g08543(.A1(new_n8735_), .A2(new_n8231_), .B1(\asqrt[28] ), .B2(new_n8733_), .ZN(new_n8736_));
  INV_X1     g08544(.I(new_n8736_), .ZN(new_n8737_));
  NOR3_X1    g08545(.A1(new_n8694_), .A2(new_n8686_), .A3(\asqrt[52] ), .ZN(new_n8738_));
  OAI21_X1   g08546(.A1(new_n8701_), .A2(new_n8738_), .B(new_n8695_), .ZN(new_n8739_));
  AOI21_X1   g08547(.A1(new_n8739_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n8740_));
  AOI21_X1   g08548(.A1(new_n8740_), .A2(new_n8712_), .B(new_n8720_), .ZN(new_n8741_));
  OAI21_X1   g08549(.A1(new_n8741_), .A2(new_n8713_), .B(\asqrt[55] ), .ZN(new_n8742_));
  NAND2_X1   g08550(.A1(new_n8742_), .A2(new_n703_), .ZN(new_n8743_));
  OAI21_X1   g08551(.A1(new_n8743_), .A2(new_n8730_), .B(new_n8737_), .ZN(new_n8744_));
  AOI21_X1   g08552(.A1(new_n8744_), .A2(new_n8731_), .B(new_n531_), .ZN(new_n8745_));
  INV_X1     g08553(.I(new_n8745_), .ZN(new_n8746_));
  INV_X1     g08554(.I(new_n8744_), .ZN(new_n8747_));
  NOR3_X1    g08555(.A1(new_n8483_), .A2(new_n8234_), .A3(new_n8344_), .ZN(new_n8748_));
  INV_X1     g08556(.I(new_n8748_), .ZN(new_n8749_));
  NOR3_X1    g08557(.A1(new_n8234_), .A2(new_n8344_), .A3(new_n8354_), .ZN(new_n8750_));
  AOI22_X1   g08558(.A1(new_n8749_), .A2(new_n8354_), .B1(\asqrt[28] ), .B2(new_n8750_), .ZN(new_n8751_));
  INV_X1     g08559(.I(new_n8751_), .ZN(new_n8752_));
  NAND2_X1   g08560(.A1(new_n8731_), .A2(new_n531_), .ZN(new_n8753_));
  OAI21_X1   g08561(.A1(new_n8753_), .A2(new_n8747_), .B(new_n8752_), .ZN(new_n8754_));
  AOI21_X1   g08562(.A1(new_n8754_), .A2(new_n8746_), .B(new_n436_), .ZN(new_n8755_));
  NOR3_X1    g08563(.A1(new_n8357_), .A2(new_n8382_), .A3(new_n8248_), .ZN(new_n8756_));
  NOR3_X1    g08564(.A1(new_n8483_), .A2(new_n8357_), .A3(new_n8382_), .ZN(new_n8757_));
  INV_X1     g08565(.I(new_n8757_), .ZN(new_n8758_));
  AOI22_X1   g08566(.A1(new_n8758_), .A2(new_n8248_), .B1(\asqrt[28] ), .B2(new_n8756_), .ZN(new_n8759_));
  NOR2_X1    g08567(.A1(new_n8745_), .A2(\asqrt[58] ), .ZN(new_n8760_));
  AOI21_X1   g08568(.A1(new_n8760_), .A2(new_n8754_), .B(new_n8759_), .ZN(new_n8761_));
  OAI21_X1   g08569(.A1(new_n8761_), .A2(new_n8755_), .B(\asqrt[59] ), .ZN(new_n8762_));
  NOR2_X1    g08570(.A1(new_n8370_), .A2(new_n8359_), .ZN(new_n8763_));
  NOR3_X1    g08571(.A1(new_n8483_), .A2(new_n8338_), .A3(new_n8763_), .ZN(new_n8764_));
  INV_X1     g08572(.I(new_n8764_), .ZN(new_n8765_));
  NOR3_X1    g08573(.A1(new_n8763_), .A2(new_n8338_), .A3(new_n8369_), .ZN(new_n8766_));
  AOI22_X1   g08574(.A1(new_n8765_), .A2(new_n8369_), .B1(\asqrt[28] ), .B2(new_n8766_), .ZN(new_n8767_));
  INV_X1     g08575(.I(new_n8767_), .ZN(new_n8768_));
  NOR3_X1    g08576(.A1(new_n8741_), .A2(\asqrt[55] ), .A3(new_n8713_), .ZN(new_n8769_));
  OAI21_X1   g08577(.A1(new_n8728_), .A2(new_n8769_), .B(new_n8742_), .ZN(new_n8770_));
  AOI21_X1   g08578(.A1(new_n8770_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n8771_));
  AOI21_X1   g08579(.A1(new_n8771_), .A2(new_n8744_), .B(new_n8751_), .ZN(new_n8772_));
  OAI21_X1   g08580(.A1(new_n8772_), .A2(new_n8745_), .B(\asqrt[58] ), .ZN(new_n8773_));
  NAND2_X1   g08581(.A1(new_n8773_), .A2(new_n327_), .ZN(new_n8774_));
  OAI21_X1   g08582(.A1(new_n8774_), .A2(new_n8761_), .B(new_n8768_), .ZN(new_n8775_));
  AOI21_X1   g08583(.A1(new_n8775_), .A2(new_n8762_), .B(new_n306_), .ZN(new_n8776_));
  INV_X1     g08584(.I(new_n8776_), .ZN(new_n8777_));
  INV_X1     g08585(.I(new_n8775_), .ZN(new_n8778_));
  NOR3_X1    g08586(.A1(new_n8432_), .A2(new_n8372_), .A3(new_n8353_), .ZN(new_n8779_));
  NOR3_X1    g08587(.A1(new_n8483_), .A2(new_n8372_), .A3(new_n8432_), .ZN(new_n8780_));
  INV_X1     g08588(.I(new_n8780_), .ZN(new_n8781_));
  AOI22_X1   g08589(.A1(new_n8781_), .A2(new_n8353_), .B1(\asqrt[28] ), .B2(new_n8779_), .ZN(new_n8782_));
  INV_X1     g08590(.I(new_n8782_), .ZN(new_n8783_));
  NAND2_X1   g08591(.A1(new_n8762_), .A2(new_n306_), .ZN(new_n8784_));
  OAI21_X1   g08592(.A1(new_n8778_), .A2(new_n8784_), .B(new_n8783_), .ZN(new_n8785_));
  AOI21_X1   g08593(.A1(new_n8785_), .A2(new_n8777_), .B(new_n218_), .ZN(new_n8786_));
  NOR3_X1    g08594(.A1(new_n8483_), .A2(new_n8363_), .A3(new_n8394_), .ZN(new_n8787_));
  INV_X1     g08595(.I(new_n8787_), .ZN(new_n8788_));
  NOR3_X1    g08596(.A1(new_n8363_), .A2(new_n8394_), .A3(new_n8428_), .ZN(new_n8789_));
  AOI22_X1   g08597(.A1(new_n8788_), .A2(new_n8428_), .B1(\asqrt[28] ), .B2(new_n8789_), .ZN(new_n8790_));
  NOR2_X1    g08598(.A1(new_n8776_), .A2(\asqrt[61] ), .ZN(new_n8791_));
  AOI21_X1   g08599(.A1(new_n8791_), .A2(new_n8785_), .B(new_n8790_), .ZN(new_n8792_));
  OAI21_X1   g08600(.A1(new_n8792_), .A2(new_n8786_), .B(\asqrt[62] ), .ZN(new_n8793_));
  NOR2_X1    g08601(.A1(new_n8387_), .A2(new_n8374_), .ZN(new_n8794_));
  NOR3_X1    g08602(.A1(new_n8794_), .A2(new_n8431_), .A3(new_n8381_), .ZN(new_n8795_));
  NOR3_X1    g08603(.A1(new_n8483_), .A2(new_n8431_), .A3(new_n8794_), .ZN(new_n8796_));
  INV_X1     g08604(.I(new_n8796_), .ZN(new_n8797_));
  AOI22_X1   g08605(.A1(new_n8797_), .A2(new_n8381_), .B1(\asqrt[28] ), .B2(new_n8795_), .ZN(new_n8798_));
  INV_X1     g08606(.I(new_n8798_), .ZN(new_n8799_));
  NOR3_X1    g08607(.A1(new_n8772_), .A2(\asqrt[58] ), .A3(new_n8745_), .ZN(new_n8800_));
  OAI21_X1   g08608(.A1(new_n8759_), .A2(new_n8800_), .B(new_n8773_), .ZN(new_n8801_));
  AOI21_X1   g08609(.A1(new_n8801_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n8802_));
  AOI21_X1   g08610(.A1(new_n8802_), .A2(new_n8775_), .B(new_n8782_), .ZN(new_n8803_));
  OAI21_X1   g08611(.A1(new_n8803_), .A2(new_n8776_), .B(\asqrt[61] ), .ZN(new_n8804_));
  NAND2_X1   g08612(.A1(new_n8804_), .A2(new_n207_), .ZN(new_n8805_));
  OAI21_X1   g08613(.A1(new_n8805_), .A2(new_n8792_), .B(new_n8799_), .ZN(new_n8806_));
  NAND4_X1   g08614(.A1(\asqrt[28] ), .A2(new_n8436_), .A3(new_n8393_), .A4(new_n8409_), .ZN(new_n8807_));
  NAND2_X1   g08615(.A1(new_n8436_), .A2(new_n8409_), .ZN(new_n8808_));
  OAI21_X1   g08616(.A1(new_n8483_), .A2(new_n8808_), .B(new_n8408_), .ZN(new_n8809_));
  NAND2_X1   g08617(.A1(new_n8809_), .A2(new_n8807_), .ZN(new_n8810_));
  AOI21_X1   g08618(.A1(new_n8410_), .A2(new_n8436_), .B(new_n8403_), .ZN(new_n8811_));
  AOI21_X1   g08619(.A1(\asqrt[28] ), .A2(new_n8811_), .B(new_n8461_), .ZN(new_n8812_));
  NAND2_X1   g08620(.A1(new_n8810_), .A2(new_n8812_), .ZN(new_n8813_));
  AOI21_X1   g08621(.A1(new_n8806_), .A2(new_n8793_), .B(new_n8813_), .ZN(new_n8814_));
  NOR3_X1    g08622(.A1(new_n8803_), .A2(\asqrt[61] ), .A3(new_n8776_), .ZN(new_n8815_));
  OAI21_X1   g08623(.A1(new_n8790_), .A2(new_n8815_), .B(new_n8804_), .ZN(new_n8816_));
  AOI21_X1   g08624(.A1(new_n8816_), .A2(\asqrt[62] ), .B(new_n8810_), .ZN(new_n8817_));
  AOI21_X1   g08625(.A1(\asqrt[28] ), .A2(new_n8411_), .B(new_n8438_), .ZN(new_n8818_));
  OR3_X2     g08626(.A1(new_n8818_), .A2(new_n193_), .A3(new_n8811_), .Z(new_n8819_));
  NAND2_X1   g08627(.A1(new_n8399_), .A2(new_n8418_), .ZN(new_n8820_));
  NOR4_X1    g08628(.A1(new_n8461_), .A2(new_n8402_), .A3(new_n8415_), .A4(new_n8820_), .ZN(new_n8821_));
  NAND2_X1   g08629(.A1(new_n8821_), .A2(new_n8407_), .ZN(new_n8822_));
  NAND2_X1   g08630(.A1(new_n8819_), .A2(new_n8822_), .ZN(new_n8823_));
  AOI21_X1   g08631(.A1(new_n8817_), .A2(new_n8806_), .B(new_n8823_), .ZN(new_n8824_));
  OAI21_X1   g08632(.A1(\asqrt[63] ), .A2(new_n8814_), .B(new_n8824_), .ZN(\asqrt[27] ));
  INV_X1     g08633(.I(\asqrt[27] ), .ZN(new_n8826_));
  NOR2_X1    g08634(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n8827_));
  INV_X1     g08635(.I(new_n8827_), .ZN(new_n8828_));
  NOR2_X1    g08636(.A1(new_n8828_), .A2(\a[54] ), .ZN(new_n8829_));
  INV_X1     g08637(.I(\a[54] ), .ZN(new_n8830_));
  INV_X1     g08638(.I(new_n8790_), .ZN(new_n8831_));
  INV_X1     g08639(.I(new_n8759_), .ZN(new_n8832_));
  INV_X1     g08640(.I(new_n8728_), .ZN(new_n8833_));
  INV_X1     g08641(.I(new_n8701_), .ZN(new_n8834_));
  INV_X1     g08642(.I(new_n8674_), .ZN(new_n8835_));
  INV_X1     g08643(.I(new_n8648_), .ZN(new_n8836_));
  INV_X1     g08644(.I(new_n8622_), .ZN(new_n8837_));
  INV_X1     g08645(.I(new_n8589_), .ZN(new_n8838_));
  NOR3_X1    g08646(.A1(new_n8588_), .A2(new_n8575_), .A3(\asqrt[41] ), .ZN(new_n8839_));
  NOR2_X1    g08647(.A1(new_n8839_), .A2(new_n8594_), .ZN(new_n8840_));
  OAI21_X1   g08648(.A1(new_n8840_), .A2(new_n8838_), .B(\asqrt[42] ), .ZN(new_n8841_));
  NAND2_X1   g08649(.A1(new_n8841_), .A2(new_n3218_), .ZN(new_n8842_));
  OAI21_X1   g08650(.A1(new_n8842_), .A2(new_n8616_), .B(new_n8837_), .ZN(new_n8843_));
  NAND3_X1   g08651(.A1(new_n8843_), .A2(new_n2954_), .A3(new_n8617_), .ZN(new_n8844_));
  AOI22_X1   g08652(.A1(new_n8844_), .A2(new_n8631_), .B1(\asqrt[44] ), .B2(new_n8640_), .ZN(new_n8845_));
  OAI21_X1   g08653(.A1(new_n8845_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n8846_));
  OAI21_X1   g08654(.A1(new_n8846_), .A2(new_n8642_), .B(new_n8836_), .ZN(new_n8847_));
  NAND3_X1   g08655(.A1(new_n8847_), .A2(new_n2229_), .A3(new_n8643_), .ZN(new_n8848_));
  AOI22_X1   g08656(.A1(new_n8848_), .A2(new_n8657_), .B1(\asqrt[47] ), .B2(new_n8666_), .ZN(new_n8849_));
  OAI21_X1   g08657(.A1(new_n8849_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n8850_));
  OAI21_X1   g08658(.A1(new_n8850_), .A2(new_n8668_), .B(new_n8835_), .ZN(new_n8851_));
  NAND3_X1   g08659(.A1(new_n8851_), .A2(new_n1612_), .A3(new_n8669_), .ZN(new_n8852_));
  AOI22_X1   g08660(.A1(new_n8852_), .A2(new_n8683_), .B1(\asqrt[50] ), .B2(new_n8692_), .ZN(new_n8853_));
  OAI21_X1   g08661(.A1(new_n8853_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n8854_));
  OAI21_X1   g08662(.A1(new_n8854_), .A2(new_n8694_), .B(new_n8834_), .ZN(new_n8855_));
  NAND3_X1   g08663(.A1(new_n8855_), .A2(new_n1103_), .A3(new_n8695_), .ZN(new_n8856_));
  AOI22_X1   g08664(.A1(new_n8856_), .A2(new_n8710_), .B1(\asqrt[53] ), .B2(new_n8739_), .ZN(new_n8857_));
  OAI21_X1   g08665(.A1(new_n8857_), .A2(new_n904_), .B(new_n823_), .ZN(new_n8858_));
  OAI21_X1   g08666(.A1(new_n8858_), .A2(new_n8741_), .B(new_n8833_), .ZN(new_n8859_));
  NAND3_X1   g08667(.A1(new_n8859_), .A2(new_n703_), .A3(new_n8742_), .ZN(new_n8860_));
  AOI22_X1   g08668(.A1(new_n8860_), .A2(new_n8737_), .B1(\asqrt[56] ), .B2(new_n8770_), .ZN(new_n8861_));
  OAI21_X1   g08669(.A1(new_n8861_), .A2(new_n531_), .B(new_n436_), .ZN(new_n8862_));
  OAI21_X1   g08670(.A1(new_n8862_), .A2(new_n8772_), .B(new_n8832_), .ZN(new_n8863_));
  NAND3_X1   g08671(.A1(new_n8863_), .A2(new_n327_), .A3(new_n8773_), .ZN(new_n8864_));
  AOI22_X1   g08672(.A1(new_n8864_), .A2(new_n8768_), .B1(new_n8801_), .B2(\asqrt[59] ), .ZN(new_n8865_));
  OAI21_X1   g08673(.A1(new_n8865_), .A2(new_n306_), .B(new_n218_), .ZN(new_n8866_));
  OAI21_X1   g08674(.A1(new_n8866_), .A2(new_n8803_), .B(new_n8831_), .ZN(new_n8867_));
  NAND3_X1   g08675(.A1(new_n8867_), .A2(new_n207_), .A3(new_n8804_), .ZN(new_n8868_));
  AOI22_X1   g08676(.A1(new_n8868_), .A2(new_n8799_), .B1(new_n8816_), .B2(\asqrt[62] ), .ZN(new_n8869_));
  OAI21_X1   g08677(.A1(new_n8869_), .A2(new_n8813_), .B(new_n193_), .ZN(new_n8870_));
  AOI21_X1   g08678(.A1(new_n8870_), .A2(new_n8824_), .B(new_n8830_), .ZN(new_n8871_));
  OAI21_X1   g08679(.A1(new_n8871_), .A2(new_n8829_), .B(\asqrt[28] ), .ZN(new_n8872_));
  INV_X1     g08680(.I(new_n8872_), .ZN(new_n8873_));
  OAI21_X1   g08681(.A1(\a[54] ), .A2(new_n8828_), .B(new_n8418_), .ZN(new_n8874_));
  NOR4_X1    g08682(.A1(new_n8461_), .A2(new_n8439_), .A3(new_n8415_), .A4(new_n8874_), .ZN(new_n8875_));
  INV_X1     g08683(.I(new_n8875_), .ZN(new_n8876_));
  NOR2_X1    g08684(.A1(new_n8871_), .A2(new_n8876_), .ZN(new_n8877_));
  AOI21_X1   g08685(.A1(new_n8870_), .A2(new_n8824_), .B(new_n8425_), .ZN(new_n8878_));
  INV_X1     g08686(.I(\a[55] ), .ZN(new_n8879_));
  AOI21_X1   g08687(.A1(\asqrt[27] ), .A2(new_n8830_), .B(new_n8879_), .ZN(new_n8880_));
  NOR3_X1    g08688(.A1(new_n8877_), .A2(new_n8880_), .A3(new_n8878_), .ZN(new_n8881_));
  OAI21_X1   g08689(.A1(new_n8881_), .A2(new_n8873_), .B(\asqrt[29] ), .ZN(new_n8882_));
  NOR2_X1    g08690(.A1(new_n8814_), .A2(\asqrt[63] ), .ZN(new_n8883_));
  INV_X1     g08691(.I(new_n8806_), .ZN(new_n8884_));
  INV_X1     g08692(.I(new_n8810_), .ZN(new_n8885_));
  NAND2_X1   g08693(.A1(new_n8793_), .A2(new_n8885_), .ZN(new_n8886_));
  INV_X1     g08694(.I(new_n8823_), .ZN(new_n8887_));
  OAI21_X1   g08695(.A1(new_n8884_), .A2(new_n8886_), .B(new_n8887_), .ZN(new_n8888_));
  OAI21_X1   g08696(.A1(new_n8883_), .A2(new_n8888_), .B(new_n8424_), .ZN(new_n8889_));
  NOR2_X1    g08697(.A1(new_n8884_), .A2(new_n8886_), .ZN(new_n8890_));
  OAI21_X1   g08698(.A1(new_n8821_), .A2(new_n8422_), .B(new_n8407_), .ZN(new_n8891_));
  NAND2_X1   g08699(.A1(new_n8819_), .A2(new_n8891_), .ZN(new_n8892_));
  NOR3_X1    g08700(.A1(new_n8883_), .A2(new_n8890_), .A3(new_n8892_), .ZN(new_n8893_));
  INV_X1     g08701(.I(new_n8893_), .ZN(new_n8894_));
  AOI21_X1   g08702(.A1(new_n8894_), .A2(new_n8889_), .B(new_n8444_), .ZN(new_n8895_));
  NOR3_X1    g08703(.A1(new_n8893_), .A2(new_n8878_), .A3(\a[56] ), .ZN(new_n8896_));
  AOI21_X1   g08704(.A1(\asqrt[27] ), .A2(\a[54] ), .B(new_n8829_), .ZN(new_n8897_));
  OAI21_X1   g08705(.A1(new_n8897_), .A2(new_n8483_), .B(new_n8036_), .ZN(new_n8898_));
  OAI22_X1   g08706(.A1(new_n8881_), .A2(new_n8898_), .B1(new_n8895_), .B2(new_n8896_), .ZN(new_n8899_));
  AOI21_X1   g08707(.A1(new_n8899_), .A2(new_n8882_), .B(new_n7539_), .ZN(new_n8900_));
  NOR3_X1    g08708(.A1(new_n8544_), .A2(new_n8443_), .A3(new_n8449_), .ZN(new_n8901_));
  NAND3_X1   g08709(.A1(\asqrt[27] ), .A2(new_n8465_), .A3(new_n8529_), .ZN(new_n8902_));
  AOI22_X1   g08710(.A1(new_n8902_), .A2(new_n8544_), .B1(\asqrt[27] ), .B2(new_n8901_), .ZN(new_n8903_));
  AOI21_X1   g08711(.A1(new_n8870_), .A2(new_n8824_), .B(\a[54] ), .ZN(new_n8904_));
  OAI21_X1   g08712(.A1(new_n8879_), .A2(new_n8904_), .B(new_n8889_), .ZN(new_n8905_));
  OAI21_X1   g08713(.A1(new_n8905_), .A2(new_n8877_), .B(new_n8872_), .ZN(new_n8906_));
  AOI21_X1   g08714(.A1(new_n8906_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n8907_));
  AOI21_X1   g08715(.A1(new_n8907_), .A2(new_n8899_), .B(new_n8903_), .ZN(new_n8908_));
  OAI21_X1   g08716(.A1(new_n8908_), .A2(new_n8900_), .B(\asqrt[31] ), .ZN(new_n8909_));
  INV_X1     g08717(.I(new_n8909_), .ZN(new_n8910_));
  NOR2_X1    g08718(.A1(new_n8464_), .A2(new_n8460_), .ZN(new_n8911_));
  INV_X1     g08719(.I(new_n8911_), .ZN(new_n8912_));
  NOR2_X1    g08720(.A1(new_n8453_), .A2(new_n8466_), .ZN(new_n8913_));
  NOR3_X1    g08721(.A1(new_n8533_), .A2(new_n8912_), .A3(new_n8913_), .ZN(new_n8914_));
  NOR3_X1    g08722(.A1(new_n8826_), .A2(new_n8533_), .A3(new_n8913_), .ZN(new_n8915_));
  INV_X1     g08723(.I(new_n8915_), .ZN(new_n8916_));
  AOI22_X1   g08724(.A1(new_n8916_), .A2(new_n8912_), .B1(\asqrt[27] ), .B2(new_n8914_), .ZN(new_n8917_));
  NOR3_X1    g08725(.A1(new_n8908_), .A2(new_n8900_), .A3(\asqrt[31] ), .ZN(new_n8918_));
  NOR2_X1    g08726(.A1(new_n8918_), .A2(new_n8917_), .ZN(new_n8919_));
  OAI21_X1   g08727(.A1(new_n8919_), .A2(new_n8910_), .B(\asqrt[32] ), .ZN(new_n8920_));
  NOR2_X1    g08728(.A1(new_n8546_), .A2(new_n8538_), .ZN(new_n8921_));
  NOR3_X1    g08729(.A1(new_n8826_), .A2(new_n8468_), .A3(new_n8921_), .ZN(new_n8922_));
  INV_X1     g08730(.I(new_n8922_), .ZN(new_n8923_));
  NOR3_X1    g08731(.A1(new_n8921_), .A2(new_n8468_), .A3(new_n8543_), .ZN(new_n8924_));
  AOI22_X1   g08732(.A1(new_n8923_), .A2(new_n8543_), .B1(\asqrt[27] ), .B2(new_n8924_), .ZN(new_n8925_));
  INV_X1     g08733(.I(new_n8925_), .ZN(new_n8926_));
  NAND2_X1   g08734(.A1(new_n8909_), .A2(new_n6824_), .ZN(new_n8927_));
  OAI21_X1   g08735(.A1(new_n8919_), .A2(new_n8927_), .B(new_n8926_), .ZN(new_n8928_));
  AOI21_X1   g08736(.A1(new_n8928_), .A2(new_n8920_), .B(new_n6356_), .ZN(new_n8929_));
  NOR3_X1    g08737(.A1(new_n8478_), .A2(new_n8487_), .A3(new_n8485_), .ZN(new_n8930_));
  NOR3_X1    g08738(.A1(new_n8826_), .A2(new_n8478_), .A3(new_n8487_), .ZN(new_n8931_));
  INV_X1     g08739(.I(new_n8931_), .ZN(new_n8932_));
  AOI22_X1   g08740(.A1(new_n8932_), .A2(new_n8485_), .B1(\asqrt[27] ), .B2(new_n8930_), .ZN(new_n8933_));
  OAI21_X1   g08741(.A1(new_n8917_), .A2(new_n8918_), .B(new_n8909_), .ZN(new_n8934_));
  AOI21_X1   g08742(.A1(new_n8934_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n8935_));
  AOI21_X1   g08743(.A1(new_n8935_), .A2(new_n8928_), .B(new_n8933_), .ZN(new_n8936_));
  OAI21_X1   g08744(.A1(new_n8936_), .A2(new_n8929_), .B(\asqrt[34] ), .ZN(new_n8937_));
  INV_X1     g08745(.I(new_n8937_), .ZN(new_n8938_));
  NOR2_X1    g08746(.A1(new_n8488_), .A2(new_n8496_), .ZN(new_n8939_));
  NOR3_X1    g08747(.A1(new_n8826_), .A2(new_n8542_), .A3(new_n8939_), .ZN(new_n8940_));
  INV_X1     g08748(.I(new_n8940_), .ZN(new_n8941_));
  NOR3_X1    g08749(.A1(new_n8939_), .A2(new_n8542_), .A3(new_n8495_), .ZN(new_n8942_));
  AOI22_X1   g08750(.A1(new_n8941_), .A2(new_n8495_), .B1(\asqrt[27] ), .B2(new_n8942_), .ZN(new_n8943_));
  NOR3_X1    g08751(.A1(new_n8936_), .A2(new_n8929_), .A3(\asqrt[34] ), .ZN(new_n8944_));
  NOR2_X1    g08752(.A1(new_n8944_), .A2(new_n8943_), .ZN(new_n8945_));
  OAI21_X1   g08753(.A1(new_n8945_), .A2(new_n8938_), .B(\asqrt[35] ), .ZN(new_n8946_));
  INV_X1     g08754(.I(new_n8502_), .ZN(new_n8947_));
  NOR3_X1    g08755(.A1(new_n8498_), .A2(new_n8596_), .A3(new_n8947_), .ZN(new_n8948_));
  NOR3_X1    g08756(.A1(new_n8826_), .A2(new_n8498_), .A3(new_n8596_), .ZN(new_n8949_));
  INV_X1     g08757(.I(new_n8949_), .ZN(new_n8950_));
  AOI22_X1   g08758(.A1(new_n8950_), .A2(new_n8947_), .B1(\asqrt[27] ), .B2(new_n8948_), .ZN(new_n8951_));
  INV_X1     g08759(.I(new_n8951_), .ZN(new_n8952_));
  NAND2_X1   g08760(.A1(new_n8937_), .A2(new_n5708_), .ZN(new_n8953_));
  OAI21_X1   g08761(.A1(new_n8945_), .A2(new_n8953_), .B(new_n8952_), .ZN(new_n8954_));
  AOI21_X1   g08762(.A1(new_n8954_), .A2(new_n8946_), .B(new_n5277_), .ZN(new_n8955_));
  NOR3_X1    g08763(.A1(new_n8826_), .A2(new_n8507_), .A3(new_n8512_), .ZN(new_n8956_));
  INV_X1     g08764(.I(new_n8956_), .ZN(new_n8957_));
  NOR3_X1    g08765(.A1(new_n8507_), .A2(new_n8528_), .A3(new_n8512_), .ZN(new_n8958_));
  AOI22_X1   g08766(.A1(new_n8957_), .A2(new_n8528_), .B1(\asqrt[27] ), .B2(new_n8958_), .ZN(new_n8959_));
  OAI21_X1   g08767(.A1(new_n8943_), .A2(new_n8944_), .B(new_n8937_), .ZN(new_n8960_));
  AOI21_X1   g08768(.A1(new_n8960_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n8961_));
  AOI21_X1   g08769(.A1(new_n8961_), .A2(new_n8954_), .B(new_n8959_), .ZN(new_n8962_));
  OAI21_X1   g08770(.A1(new_n8962_), .A2(new_n8955_), .B(\asqrt[37] ), .ZN(new_n8963_));
  INV_X1     g08771(.I(new_n8963_), .ZN(new_n8964_));
  INV_X1     g08772(.I(new_n8582_), .ZN(new_n8965_));
  NOR3_X1    g08773(.A1(new_n8965_), .A2(new_n8554_), .A3(new_n8520_), .ZN(new_n8966_));
  NOR3_X1    g08774(.A1(new_n8826_), .A2(new_n8554_), .A3(new_n8965_), .ZN(new_n8967_));
  INV_X1     g08775(.I(new_n8967_), .ZN(new_n8968_));
  AOI22_X1   g08776(.A1(new_n8968_), .A2(new_n8520_), .B1(\asqrt[27] ), .B2(new_n8966_), .ZN(new_n8969_));
  NOR3_X1    g08777(.A1(new_n8962_), .A2(new_n8955_), .A3(\asqrt[37] ), .ZN(new_n8970_));
  NOR2_X1    g08778(.A1(new_n8970_), .A2(new_n8969_), .ZN(new_n8971_));
  OAI21_X1   g08779(.A1(new_n8971_), .A2(new_n8964_), .B(\asqrt[38] ), .ZN(new_n8972_));
  INV_X1     g08780(.I(new_n8527_), .ZN(new_n8973_));
  NOR3_X1    g08781(.A1(new_n8826_), .A2(new_n8523_), .A3(new_n8600_), .ZN(new_n8974_));
  INV_X1     g08782(.I(new_n8974_), .ZN(new_n8975_));
  NOR3_X1    g08783(.A1(new_n8523_), .A2(new_n8600_), .A3(new_n8973_), .ZN(new_n8976_));
  AOI22_X1   g08784(.A1(new_n8975_), .A2(new_n8973_), .B1(\asqrt[27] ), .B2(new_n8976_), .ZN(new_n8977_));
  INV_X1     g08785(.I(new_n8977_), .ZN(new_n8978_));
  NAND2_X1   g08786(.A1(new_n8963_), .A2(new_n4696_), .ZN(new_n8979_));
  OAI21_X1   g08787(.A1(new_n8971_), .A2(new_n8979_), .B(new_n8978_), .ZN(new_n8980_));
  AOI21_X1   g08788(.A1(new_n8980_), .A2(new_n8972_), .B(new_n4298_), .ZN(new_n8981_));
  NOR3_X1    g08789(.A1(new_n8558_), .A2(new_n8580_), .A3(new_n8564_), .ZN(new_n8982_));
  NOR3_X1    g08790(.A1(new_n8826_), .A2(new_n8558_), .A3(new_n8564_), .ZN(new_n8983_));
  INV_X1     g08791(.I(new_n8983_), .ZN(new_n8984_));
  AOI22_X1   g08792(.A1(new_n8984_), .A2(new_n8580_), .B1(\asqrt[27] ), .B2(new_n8982_), .ZN(new_n8985_));
  OAI21_X1   g08793(.A1(new_n8969_), .A2(new_n8970_), .B(new_n8963_), .ZN(new_n8986_));
  AOI21_X1   g08794(.A1(new_n8986_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n8987_));
  AOI21_X1   g08795(.A1(new_n8987_), .A2(new_n8980_), .B(new_n8985_), .ZN(new_n8988_));
  OAI21_X1   g08796(.A1(new_n8988_), .A2(new_n8981_), .B(\asqrt[40] ), .ZN(new_n8989_));
  INV_X1     g08797(.I(new_n8989_), .ZN(new_n8990_));
  NOR2_X1    g08798(.A1(new_n8565_), .A2(new_n8573_), .ZN(new_n8991_));
  NOR3_X1    g08799(.A1(new_n8826_), .A2(new_n8586_), .A3(new_n8991_), .ZN(new_n8992_));
  INV_X1     g08800(.I(new_n8992_), .ZN(new_n8993_));
  NOR3_X1    g08801(.A1(new_n8991_), .A2(new_n8586_), .A3(new_n8572_), .ZN(new_n8994_));
  AOI22_X1   g08802(.A1(new_n8993_), .A2(new_n8572_), .B1(\asqrt[27] ), .B2(new_n8994_), .ZN(new_n8995_));
  NOR3_X1    g08803(.A1(new_n8988_), .A2(new_n8981_), .A3(\asqrt[40] ), .ZN(new_n8996_));
  NOR2_X1    g08804(.A1(new_n8996_), .A2(new_n8995_), .ZN(new_n8997_));
  OAI21_X1   g08805(.A1(new_n8997_), .A2(new_n8990_), .B(\asqrt[41] ), .ZN(new_n8998_));
  INV_X1     g08806(.I(new_n8579_), .ZN(new_n8999_));
  NOR3_X1    g08807(.A1(new_n8575_), .A2(new_n8613_), .A3(new_n8999_), .ZN(new_n9000_));
  NOR3_X1    g08808(.A1(new_n8826_), .A2(new_n8575_), .A3(new_n8613_), .ZN(new_n9001_));
  INV_X1     g08809(.I(new_n9001_), .ZN(new_n9002_));
  AOI22_X1   g08810(.A1(new_n9002_), .A2(new_n8999_), .B1(\asqrt[27] ), .B2(new_n9000_), .ZN(new_n9003_));
  INV_X1     g08811(.I(new_n9003_), .ZN(new_n9004_));
  NAND2_X1   g08812(.A1(new_n8989_), .A2(new_n3782_), .ZN(new_n9005_));
  OAI21_X1   g08813(.A1(new_n8997_), .A2(new_n9005_), .B(new_n9004_), .ZN(new_n9006_));
  AOI21_X1   g08814(.A1(new_n9006_), .A2(new_n8998_), .B(new_n3419_), .ZN(new_n9007_));
  NOR3_X1    g08815(.A1(new_n8826_), .A2(new_n8838_), .A3(new_n8839_), .ZN(new_n9008_));
  INV_X1     g08816(.I(new_n9008_), .ZN(new_n9009_));
  NOR3_X1    g08817(.A1(new_n8838_), .A2(new_n8595_), .A3(new_n8839_), .ZN(new_n9010_));
  AOI22_X1   g08818(.A1(new_n9009_), .A2(new_n8595_), .B1(\asqrt[27] ), .B2(new_n9010_), .ZN(new_n9011_));
  OAI21_X1   g08819(.A1(new_n8995_), .A2(new_n8996_), .B(new_n8989_), .ZN(new_n9012_));
  AOI21_X1   g08820(.A1(new_n9012_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n9013_));
  AOI21_X1   g08821(.A1(new_n9013_), .A2(new_n9006_), .B(new_n9011_), .ZN(new_n9014_));
  OAI21_X1   g08822(.A1(new_n9014_), .A2(new_n9007_), .B(\asqrt[43] ), .ZN(new_n9015_));
  INV_X1     g08823(.I(new_n9015_), .ZN(new_n9016_));
  INV_X1     g08824(.I(new_n8612_), .ZN(new_n9017_));
  NAND2_X1   g08825(.A1(new_n8589_), .A2(new_n3419_), .ZN(new_n9018_));
  NOR2_X1    g08826(.A1(new_n8840_), .A2(new_n9018_), .ZN(new_n9019_));
  NOR3_X1    g08827(.A1(new_n9019_), .A2(new_n8607_), .A3(new_n9017_), .ZN(new_n9020_));
  NOR3_X1    g08828(.A1(new_n8826_), .A2(new_n8607_), .A3(new_n9019_), .ZN(new_n9021_));
  INV_X1     g08829(.I(new_n9021_), .ZN(new_n9022_));
  AOI22_X1   g08830(.A1(new_n9022_), .A2(new_n9017_), .B1(\asqrt[27] ), .B2(new_n9020_), .ZN(new_n9023_));
  NOR3_X1    g08831(.A1(new_n9014_), .A2(new_n9007_), .A3(\asqrt[43] ), .ZN(new_n9024_));
  NOR2_X1    g08832(.A1(new_n9024_), .A2(new_n9023_), .ZN(new_n9025_));
  OAI21_X1   g08833(.A1(new_n9025_), .A2(new_n9016_), .B(\asqrt[44] ), .ZN(new_n9026_));
  NOR3_X1    g08834(.A1(new_n8826_), .A2(new_n8618_), .A3(new_n8623_), .ZN(new_n9027_));
  INV_X1     g08835(.I(new_n9027_), .ZN(new_n9028_));
  NOR3_X1    g08836(.A1(new_n8618_), .A2(new_n8837_), .A3(new_n8623_), .ZN(new_n9029_));
  AOI22_X1   g08837(.A1(new_n9028_), .A2(new_n8837_), .B1(\asqrt[27] ), .B2(new_n9029_), .ZN(new_n9030_));
  INV_X1     g08838(.I(new_n9030_), .ZN(new_n9031_));
  NAND2_X1   g08839(.A1(new_n9015_), .A2(new_n2954_), .ZN(new_n9032_));
  OAI21_X1   g08840(.A1(new_n9025_), .A2(new_n9032_), .B(new_n9031_), .ZN(new_n9033_));
  AOI21_X1   g08841(.A1(new_n9033_), .A2(new_n9026_), .B(new_n2641_), .ZN(new_n9034_));
  INV_X1     g08842(.I(new_n8625_), .ZN(new_n9035_));
  NOR2_X1    g08843(.A1(new_n8624_), .A2(new_n8632_), .ZN(new_n9036_));
  NOR3_X1    g08844(.A1(new_n9035_), .A2(new_n9036_), .A3(new_n8631_), .ZN(new_n9037_));
  NOR3_X1    g08845(.A1(new_n8826_), .A2(new_n9035_), .A3(new_n9036_), .ZN(new_n9038_));
  INV_X1     g08846(.I(new_n9038_), .ZN(new_n9039_));
  AOI22_X1   g08847(.A1(new_n9039_), .A2(new_n8631_), .B1(\asqrt[27] ), .B2(new_n9037_), .ZN(new_n9040_));
  OAI21_X1   g08848(.A1(new_n9023_), .A2(new_n9024_), .B(new_n9015_), .ZN(new_n9041_));
  AOI21_X1   g08849(.A1(new_n9041_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n9042_));
  AOI21_X1   g08850(.A1(new_n9042_), .A2(new_n9033_), .B(new_n9040_), .ZN(new_n9043_));
  OAI21_X1   g08851(.A1(new_n9043_), .A2(new_n9034_), .B(\asqrt[46] ), .ZN(new_n9044_));
  INV_X1     g08852(.I(new_n9044_), .ZN(new_n9045_));
  INV_X1     g08853(.I(new_n8639_), .ZN(new_n9046_));
  INV_X1     g08854(.I(new_n8633_), .ZN(new_n9047_));
  INV_X1     g08855(.I(new_n8641_), .ZN(new_n9048_));
  NOR2_X1    g08856(.A1(new_n9048_), .A2(new_n9047_), .ZN(new_n9049_));
  NOR3_X1    g08857(.A1(new_n8826_), .A2(new_n8634_), .A3(new_n9049_), .ZN(new_n9050_));
  INV_X1     g08858(.I(new_n9050_), .ZN(new_n9051_));
  NOR3_X1    g08859(.A1(new_n9049_), .A2(new_n8634_), .A3(new_n9046_), .ZN(new_n9052_));
  AOI22_X1   g08860(.A1(new_n9051_), .A2(new_n9046_), .B1(\asqrt[27] ), .B2(new_n9052_), .ZN(new_n9053_));
  NOR3_X1    g08861(.A1(new_n9043_), .A2(new_n9034_), .A3(\asqrt[46] ), .ZN(new_n9054_));
  NOR2_X1    g08862(.A1(new_n9054_), .A2(new_n9053_), .ZN(new_n9055_));
  OAI21_X1   g08863(.A1(new_n9055_), .A2(new_n9045_), .B(\asqrt[47] ), .ZN(new_n9056_));
  NOR3_X1    g08864(.A1(new_n8644_), .A2(new_n8836_), .A3(new_n8649_), .ZN(new_n9057_));
  NOR3_X1    g08865(.A1(new_n8826_), .A2(new_n8644_), .A3(new_n8649_), .ZN(new_n9058_));
  INV_X1     g08866(.I(new_n9058_), .ZN(new_n9059_));
  AOI22_X1   g08867(.A1(new_n9059_), .A2(new_n8836_), .B1(\asqrt[27] ), .B2(new_n9057_), .ZN(new_n9060_));
  INV_X1     g08868(.I(new_n9060_), .ZN(new_n9061_));
  NAND2_X1   g08869(.A1(new_n9044_), .A2(new_n2229_), .ZN(new_n9062_));
  OAI21_X1   g08870(.A1(new_n9055_), .A2(new_n9062_), .B(new_n9061_), .ZN(new_n9063_));
  AOI21_X1   g08871(.A1(new_n9063_), .A2(new_n9056_), .B(new_n1956_), .ZN(new_n9064_));
  INV_X1     g08872(.I(new_n8651_), .ZN(new_n9065_));
  NOR2_X1    g08873(.A1(new_n8650_), .A2(new_n8658_), .ZN(new_n9066_));
  NOR3_X1    g08874(.A1(new_n8826_), .A2(new_n9065_), .A3(new_n9066_), .ZN(new_n9067_));
  INV_X1     g08875(.I(new_n9067_), .ZN(new_n9068_));
  NOR3_X1    g08876(.A1(new_n9065_), .A2(new_n9066_), .A3(new_n8657_), .ZN(new_n9069_));
  AOI22_X1   g08877(.A1(new_n9068_), .A2(new_n8657_), .B1(\asqrt[27] ), .B2(new_n9069_), .ZN(new_n9070_));
  OAI21_X1   g08878(.A1(new_n9053_), .A2(new_n9054_), .B(new_n9044_), .ZN(new_n9071_));
  AOI21_X1   g08879(.A1(new_n9071_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n9072_));
  AOI21_X1   g08880(.A1(new_n9072_), .A2(new_n9063_), .B(new_n9070_), .ZN(new_n9073_));
  OAI21_X1   g08881(.A1(new_n9073_), .A2(new_n9064_), .B(\asqrt[49] ), .ZN(new_n9074_));
  INV_X1     g08882(.I(new_n9074_), .ZN(new_n9075_));
  INV_X1     g08883(.I(new_n8665_), .ZN(new_n9076_));
  INV_X1     g08884(.I(new_n8659_), .ZN(new_n9077_));
  INV_X1     g08885(.I(new_n8667_), .ZN(new_n9078_));
  NOR2_X1    g08886(.A1(new_n9078_), .A2(new_n9077_), .ZN(new_n9079_));
  NOR3_X1    g08887(.A1(new_n9079_), .A2(new_n8660_), .A3(new_n9076_), .ZN(new_n9080_));
  NOR3_X1    g08888(.A1(new_n8826_), .A2(new_n8660_), .A3(new_n9079_), .ZN(new_n9081_));
  INV_X1     g08889(.I(new_n9081_), .ZN(new_n9082_));
  AOI22_X1   g08890(.A1(new_n9082_), .A2(new_n9076_), .B1(\asqrt[27] ), .B2(new_n9080_), .ZN(new_n9083_));
  NOR3_X1    g08891(.A1(new_n9073_), .A2(new_n9064_), .A3(\asqrt[49] ), .ZN(new_n9084_));
  NOR2_X1    g08892(.A1(new_n9084_), .A2(new_n9083_), .ZN(new_n9085_));
  OAI21_X1   g08893(.A1(new_n9085_), .A2(new_n9075_), .B(\asqrt[50] ), .ZN(new_n9086_));
  NOR3_X1    g08894(.A1(new_n8826_), .A2(new_n8670_), .A3(new_n8675_), .ZN(new_n9087_));
  INV_X1     g08895(.I(new_n9087_), .ZN(new_n9088_));
  NOR3_X1    g08896(.A1(new_n8670_), .A2(new_n8835_), .A3(new_n8675_), .ZN(new_n9089_));
  AOI22_X1   g08897(.A1(new_n9088_), .A2(new_n8835_), .B1(\asqrt[27] ), .B2(new_n9089_), .ZN(new_n9090_));
  INV_X1     g08898(.I(new_n9090_), .ZN(new_n9091_));
  NAND2_X1   g08899(.A1(new_n9074_), .A2(new_n1612_), .ZN(new_n9092_));
  OAI21_X1   g08900(.A1(new_n9085_), .A2(new_n9092_), .B(new_n9091_), .ZN(new_n9093_));
  AOI21_X1   g08901(.A1(new_n9093_), .A2(new_n9086_), .B(new_n1376_), .ZN(new_n9094_));
  INV_X1     g08902(.I(new_n8677_), .ZN(new_n9095_));
  NOR2_X1    g08903(.A1(new_n8676_), .A2(new_n8684_), .ZN(new_n9096_));
  NOR3_X1    g08904(.A1(new_n9095_), .A2(new_n8683_), .A3(new_n9096_), .ZN(new_n9097_));
  NOR3_X1    g08905(.A1(new_n8826_), .A2(new_n9095_), .A3(new_n9096_), .ZN(new_n9098_));
  INV_X1     g08906(.I(new_n9098_), .ZN(new_n9099_));
  AOI22_X1   g08907(.A1(new_n9099_), .A2(new_n8683_), .B1(\asqrt[27] ), .B2(new_n9097_), .ZN(new_n9100_));
  OAI21_X1   g08908(.A1(new_n9083_), .A2(new_n9084_), .B(new_n9074_), .ZN(new_n9101_));
  AOI21_X1   g08909(.A1(new_n9101_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n9102_));
  AOI21_X1   g08910(.A1(new_n9102_), .A2(new_n9093_), .B(new_n9100_), .ZN(new_n9103_));
  OAI21_X1   g08911(.A1(new_n9103_), .A2(new_n9094_), .B(\asqrt[52] ), .ZN(new_n9104_));
  INV_X1     g08912(.I(new_n8691_), .ZN(new_n9105_));
  INV_X1     g08913(.I(new_n8685_), .ZN(new_n9106_));
  INV_X1     g08914(.I(new_n8693_), .ZN(new_n9107_));
  NOR2_X1    g08915(.A1(new_n9107_), .A2(new_n9106_), .ZN(new_n9108_));
  NOR3_X1    g08916(.A1(new_n8826_), .A2(new_n8686_), .A3(new_n9108_), .ZN(new_n9109_));
  INV_X1     g08917(.I(new_n9109_), .ZN(new_n9110_));
  NOR3_X1    g08918(.A1(new_n9108_), .A2(new_n8686_), .A3(new_n9105_), .ZN(new_n9111_));
  AOI22_X1   g08919(.A1(new_n9110_), .A2(new_n9105_), .B1(\asqrt[27] ), .B2(new_n9111_), .ZN(new_n9112_));
  INV_X1     g08920(.I(new_n9112_), .ZN(new_n9113_));
  INV_X1     g08921(.I(new_n9083_), .ZN(new_n9114_));
  INV_X1     g08922(.I(new_n9064_), .ZN(new_n9115_));
  NAND2_X1   g08923(.A1(new_n9115_), .A2(new_n1806_), .ZN(new_n9116_));
  OAI21_X1   g08924(.A1(new_n9116_), .A2(new_n9073_), .B(new_n9114_), .ZN(new_n9117_));
  AOI21_X1   g08925(.A1(new_n9117_), .A2(new_n9074_), .B(new_n1612_), .ZN(new_n9118_));
  INV_X1     g08926(.I(new_n9092_), .ZN(new_n9119_));
  AOI21_X1   g08927(.A1(new_n9119_), .A2(new_n9117_), .B(new_n9090_), .ZN(new_n9120_));
  OAI21_X1   g08928(.A1(new_n9120_), .A2(new_n9118_), .B(\asqrt[51] ), .ZN(new_n9121_));
  NAND2_X1   g08929(.A1(new_n9121_), .A2(new_n1256_), .ZN(new_n9122_));
  OAI21_X1   g08930(.A1(new_n9122_), .A2(new_n9103_), .B(new_n9113_), .ZN(new_n9123_));
  AOI21_X1   g08931(.A1(new_n9123_), .A2(new_n9104_), .B(new_n1103_), .ZN(new_n9124_));
  NOR3_X1    g08932(.A1(new_n8696_), .A2(new_n8834_), .A3(new_n8738_), .ZN(new_n9125_));
  NOR3_X1    g08933(.A1(new_n8826_), .A2(new_n8696_), .A3(new_n8738_), .ZN(new_n9126_));
  INV_X1     g08934(.I(new_n9126_), .ZN(new_n9127_));
  AOI22_X1   g08935(.A1(new_n9127_), .A2(new_n8834_), .B1(\asqrt[27] ), .B2(new_n9125_), .ZN(new_n9128_));
  INV_X1     g08936(.I(new_n9100_), .ZN(new_n9129_));
  NAND2_X1   g08937(.A1(new_n9086_), .A2(new_n1376_), .ZN(new_n9130_));
  OAI21_X1   g08938(.A1(new_n9130_), .A2(new_n9120_), .B(new_n9129_), .ZN(new_n9131_));
  AOI21_X1   g08939(.A1(new_n9131_), .A2(new_n9121_), .B(new_n1256_), .ZN(new_n9132_));
  NOR2_X1    g08940(.A1(new_n9132_), .A2(\asqrt[53] ), .ZN(new_n9133_));
  AOI21_X1   g08941(.A1(new_n9133_), .A2(new_n9123_), .B(new_n9128_), .ZN(new_n9134_));
  OAI21_X1   g08942(.A1(new_n9134_), .A2(new_n9124_), .B(\asqrt[54] ), .ZN(new_n9135_));
  INV_X1     g08943(.I(new_n8704_), .ZN(new_n9136_));
  NOR2_X1    g08944(.A1(new_n8711_), .A2(new_n8703_), .ZN(new_n9137_));
  NOR3_X1    g08945(.A1(new_n8826_), .A2(new_n9136_), .A3(new_n9137_), .ZN(new_n9138_));
  INV_X1     g08946(.I(new_n9138_), .ZN(new_n9139_));
  NOR3_X1    g08947(.A1(new_n9136_), .A2(new_n8710_), .A3(new_n9137_), .ZN(new_n9140_));
  AOI22_X1   g08948(.A1(new_n9139_), .A2(new_n8710_), .B1(\asqrt[27] ), .B2(new_n9140_), .ZN(new_n9141_));
  INV_X1     g08949(.I(new_n9141_), .ZN(new_n9142_));
  NOR2_X1    g08950(.A1(new_n9094_), .A2(\asqrt[52] ), .ZN(new_n9143_));
  AOI21_X1   g08951(.A1(new_n9143_), .A2(new_n9131_), .B(new_n9112_), .ZN(new_n9144_));
  OAI21_X1   g08952(.A1(new_n9144_), .A2(new_n9132_), .B(\asqrt[53] ), .ZN(new_n9145_));
  NAND2_X1   g08953(.A1(new_n9145_), .A2(new_n904_), .ZN(new_n9146_));
  OAI21_X1   g08954(.A1(new_n9146_), .A2(new_n9134_), .B(new_n9142_), .ZN(new_n9147_));
  AOI21_X1   g08955(.A1(new_n9147_), .A2(new_n9135_), .B(new_n823_), .ZN(new_n9148_));
  NOR2_X1    g08956(.A1(new_n8722_), .A2(new_n8715_), .ZN(new_n9149_));
  NOR3_X1    g08957(.A1(new_n9149_), .A2(new_n8713_), .A3(new_n8721_), .ZN(new_n9150_));
  NOR3_X1    g08958(.A1(new_n8826_), .A2(new_n8713_), .A3(new_n9149_), .ZN(new_n9151_));
  INV_X1     g08959(.I(new_n9151_), .ZN(new_n9152_));
  AOI22_X1   g08960(.A1(new_n9152_), .A2(new_n8721_), .B1(\asqrt[27] ), .B2(new_n9150_), .ZN(new_n9153_));
  INV_X1     g08961(.I(new_n9128_), .ZN(new_n9154_));
  NAND2_X1   g08962(.A1(new_n9104_), .A2(new_n1103_), .ZN(new_n9155_));
  OAI21_X1   g08963(.A1(new_n9155_), .A2(new_n9144_), .B(new_n9154_), .ZN(new_n9156_));
  AOI21_X1   g08964(.A1(new_n9156_), .A2(new_n9145_), .B(new_n904_), .ZN(new_n9157_));
  NOR2_X1    g08965(.A1(new_n9157_), .A2(\asqrt[55] ), .ZN(new_n9158_));
  AOI21_X1   g08966(.A1(new_n9158_), .A2(new_n9147_), .B(new_n9153_), .ZN(new_n9159_));
  OAI21_X1   g08967(.A1(new_n9159_), .A2(new_n9148_), .B(\asqrt[56] ), .ZN(new_n9160_));
  NOR3_X1    g08968(.A1(new_n8826_), .A2(new_n8724_), .A3(new_n8769_), .ZN(new_n9161_));
  INV_X1     g08969(.I(new_n9161_), .ZN(new_n9162_));
  NOR3_X1    g08970(.A1(new_n8724_), .A2(new_n8833_), .A3(new_n8769_), .ZN(new_n9163_));
  AOI22_X1   g08971(.A1(new_n9162_), .A2(new_n8833_), .B1(\asqrt[27] ), .B2(new_n9163_), .ZN(new_n9164_));
  INV_X1     g08972(.I(new_n9164_), .ZN(new_n9165_));
  NOR3_X1    g08973(.A1(new_n9103_), .A2(new_n9094_), .A3(\asqrt[52] ), .ZN(new_n9166_));
  OAI21_X1   g08974(.A1(new_n9112_), .A2(new_n9166_), .B(new_n9104_), .ZN(new_n9167_));
  AOI21_X1   g08975(.A1(new_n9167_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n9168_));
  AOI21_X1   g08976(.A1(new_n9168_), .A2(new_n9156_), .B(new_n9141_), .ZN(new_n9169_));
  OAI21_X1   g08977(.A1(new_n9169_), .A2(new_n9157_), .B(\asqrt[55] ), .ZN(new_n9170_));
  NAND2_X1   g08978(.A1(new_n9170_), .A2(new_n703_), .ZN(new_n9171_));
  OAI21_X1   g08979(.A1(new_n9171_), .A2(new_n9159_), .B(new_n9165_), .ZN(new_n9172_));
  AOI21_X1   g08980(.A1(new_n9172_), .A2(new_n9160_), .B(new_n531_), .ZN(new_n9173_));
  INV_X1     g08981(.I(new_n8731_), .ZN(new_n9174_));
  NOR2_X1    g08982(.A1(new_n8743_), .A2(new_n8730_), .ZN(new_n9175_));
  NOR3_X1    g08983(.A1(new_n9174_), .A2(new_n8737_), .A3(new_n9175_), .ZN(new_n9176_));
  NOR3_X1    g08984(.A1(new_n8826_), .A2(new_n9174_), .A3(new_n9175_), .ZN(new_n9177_));
  INV_X1     g08985(.I(new_n9177_), .ZN(new_n9178_));
  AOI22_X1   g08986(.A1(new_n9178_), .A2(new_n8737_), .B1(\asqrt[27] ), .B2(new_n9176_), .ZN(new_n9179_));
  NOR3_X1    g08987(.A1(new_n9169_), .A2(\asqrt[55] ), .A3(new_n9157_), .ZN(new_n9180_));
  OAI21_X1   g08988(.A1(new_n9153_), .A2(new_n9180_), .B(new_n9170_), .ZN(new_n9181_));
  AOI21_X1   g08989(.A1(new_n9181_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n9182_));
  AOI21_X1   g08990(.A1(new_n9182_), .A2(new_n9172_), .B(new_n9179_), .ZN(new_n9183_));
  OAI21_X1   g08991(.A1(new_n9183_), .A2(new_n9173_), .B(\asqrt[58] ), .ZN(new_n9184_));
  NOR2_X1    g08992(.A1(new_n8753_), .A2(new_n8747_), .ZN(new_n9185_));
  NOR3_X1    g08993(.A1(new_n8826_), .A2(new_n8745_), .A3(new_n9185_), .ZN(new_n9186_));
  INV_X1     g08994(.I(new_n9186_), .ZN(new_n9187_));
  NOR3_X1    g08995(.A1(new_n9185_), .A2(new_n8745_), .A3(new_n8752_), .ZN(new_n9188_));
  AOI22_X1   g08996(.A1(new_n9187_), .A2(new_n8752_), .B1(\asqrt[27] ), .B2(new_n9188_), .ZN(new_n9189_));
  INV_X1     g08997(.I(new_n9189_), .ZN(new_n9190_));
  INV_X1     g08998(.I(new_n9153_), .ZN(new_n9191_));
  NAND2_X1   g08999(.A1(new_n9135_), .A2(new_n823_), .ZN(new_n9192_));
  OAI21_X1   g09000(.A1(new_n9192_), .A2(new_n9169_), .B(new_n9191_), .ZN(new_n9193_));
  AOI21_X1   g09001(.A1(new_n9193_), .A2(new_n9170_), .B(new_n703_), .ZN(new_n9194_));
  NOR2_X1    g09002(.A1(new_n9148_), .A2(\asqrt[56] ), .ZN(new_n9195_));
  AOI21_X1   g09003(.A1(new_n9195_), .A2(new_n9193_), .B(new_n9164_), .ZN(new_n9196_));
  OAI21_X1   g09004(.A1(new_n9196_), .A2(new_n9194_), .B(\asqrt[57] ), .ZN(new_n9197_));
  NAND2_X1   g09005(.A1(new_n9197_), .A2(new_n436_), .ZN(new_n9198_));
  OAI21_X1   g09006(.A1(new_n9198_), .A2(new_n9183_), .B(new_n9190_), .ZN(new_n9199_));
  AOI21_X1   g09007(.A1(new_n9199_), .A2(new_n9184_), .B(new_n327_), .ZN(new_n9200_));
  NOR3_X1    g09008(.A1(new_n8755_), .A2(new_n8832_), .A3(new_n8800_), .ZN(new_n9201_));
  NOR3_X1    g09009(.A1(new_n8826_), .A2(new_n8755_), .A3(new_n8800_), .ZN(new_n9202_));
  INV_X1     g09010(.I(new_n9202_), .ZN(new_n9203_));
  AOI22_X1   g09011(.A1(new_n9203_), .A2(new_n8832_), .B1(\asqrt[27] ), .B2(new_n9201_), .ZN(new_n9204_));
  INV_X1     g09012(.I(new_n9179_), .ZN(new_n9205_));
  NAND2_X1   g09013(.A1(new_n9160_), .A2(new_n531_), .ZN(new_n9206_));
  OAI21_X1   g09014(.A1(new_n9206_), .A2(new_n9196_), .B(new_n9205_), .ZN(new_n9207_));
  AOI21_X1   g09015(.A1(new_n9207_), .A2(new_n9197_), .B(new_n436_), .ZN(new_n9208_));
  NOR2_X1    g09016(.A1(new_n9208_), .A2(\asqrt[59] ), .ZN(new_n9209_));
  AOI21_X1   g09017(.A1(new_n9209_), .A2(new_n9199_), .B(new_n9204_), .ZN(new_n9210_));
  OAI21_X1   g09018(.A1(new_n9210_), .A2(new_n9200_), .B(\asqrt[60] ), .ZN(new_n9211_));
  INV_X1     g09019(.I(new_n8762_), .ZN(new_n9212_));
  NOR2_X1    g09020(.A1(new_n8774_), .A2(new_n8761_), .ZN(new_n9213_));
  NOR3_X1    g09021(.A1(new_n8826_), .A2(new_n9212_), .A3(new_n9213_), .ZN(new_n9214_));
  INV_X1     g09022(.I(new_n9214_), .ZN(new_n9215_));
  NOR3_X1    g09023(.A1(new_n9212_), .A2(new_n8768_), .A3(new_n9213_), .ZN(new_n9216_));
  AOI22_X1   g09024(.A1(new_n9215_), .A2(new_n8768_), .B1(\asqrt[27] ), .B2(new_n9216_), .ZN(new_n9217_));
  INV_X1     g09025(.I(new_n9217_), .ZN(new_n9218_));
  NOR2_X1    g09026(.A1(new_n9173_), .A2(\asqrt[58] ), .ZN(new_n9219_));
  AOI21_X1   g09027(.A1(new_n9219_), .A2(new_n9207_), .B(new_n9189_), .ZN(new_n9220_));
  OAI21_X1   g09028(.A1(new_n9220_), .A2(new_n9208_), .B(\asqrt[59] ), .ZN(new_n9221_));
  NAND2_X1   g09029(.A1(new_n9221_), .A2(new_n306_), .ZN(new_n9222_));
  OAI21_X1   g09030(.A1(new_n9222_), .A2(new_n9210_), .B(new_n9218_), .ZN(new_n9223_));
  AOI21_X1   g09031(.A1(new_n9223_), .A2(new_n9211_), .B(new_n218_), .ZN(new_n9224_));
  NOR2_X1    g09032(.A1(new_n8778_), .A2(new_n8784_), .ZN(new_n9225_));
  NOR3_X1    g09033(.A1(new_n9225_), .A2(new_n8776_), .A3(new_n8783_), .ZN(new_n9226_));
  NOR3_X1    g09034(.A1(new_n8826_), .A2(new_n8776_), .A3(new_n9225_), .ZN(new_n9227_));
  INV_X1     g09035(.I(new_n9227_), .ZN(new_n9228_));
  AOI22_X1   g09036(.A1(new_n9228_), .A2(new_n8783_), .B1(\asqrt[27] ), .B2(new_n9226_), .ZN(new_n9229_));
  INV_X1     g09037(.I(new_n9204_), .ZN(new_n9230_));
  NAND2_X1   g09038(.A1(new_n9184_), .A2(new_n327_), .ZN(new_n9231_));
  OAI21_X1   g09039(.A1(new_n9231_), .A2(new_n9220_), .B(new_n9230_), .ZN(new_n9232_));
  AOI21_X1   g09040(.A1(new_n9232_), .A2(new_n9221_), .B(new_n306_), .ZN(new_n9233_));
  NOR2_X1    g09041(.A1(new_n9233_), .A2(\asqrt[61] ), .ZN(new_n9234_));
  AOI21_X1   g09042(.A1(new_n9234_), .A2(new_n9223_), .B(new_n9229_), .ZN(new_n9235_));
  OAI21_X1   g09043(.A1(new_n9235_), .A2(new_n9224_), .B(\asqrt[62] ), .ZN(new_n9236_));
  NOR3_X1    g09044(.A1(new_n8826_), .A2(new_n8786_), .A3(new_n8815_), .ZN(new_n9237_));
  INV_X1     g09045(.I(new_n9237_), .ZN(new_n9238_));
  NOR3_X1    g09046(.A1(new_n8786_), .A2(new_n8831_), .A3(new_n8815_), .ZN(new_n9239_));
  AOI22_X1   g09047(.A1(new_n9238_), .A2(new_n8831_), .B1(\asqrt[27] ), .B2(new_n9239_), .ZN(new_n9240_));
  INV_X1     g09048(.I(new_n9240_), .ZN(new_n9241_));
  NOR3_X1    g09049(.A1(new_n9183_), .A2(\asqrt[58] ), .A3(new_n9173_), .ZN(new_n9242_));
  OAI21_X1   g09050(.A1(new_n9189_), .A2(new_n9242_), .B(new_n9184_), .ZN(new_n9243_));
  AOI21_X1   g09051(.A1(new_n9243_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n9244_));
  AOI21_X1   g09052(.A1(new_n9244_), .A2(new_n9232_), .B(new_n9217_), .ZN(new_n9245_));
  OAI21_X1   g09053(.A1(new_n9245_), .A2(new_n9233_), .B(\asqrt[61] ), .ZN(new_n9246_));
  NAND2_X1   g09054(.A1(new_n9246_), .A2(new_n207_), .ZN(new_n9247_));
  OAI21_X1   g09055(.A1(new_n9247_), .A2(new_n9235_), .B(new_n9241_), .ZN(new_n9248_));
  INV_X1     g09056(.I(new_n8890_), .ZN(new_n9249_));
  NAND4_X1   g09057(.A1(\asqrt[27] ), .A2(new_n8793_), .A3(new_n8798_), .A4(new_n8868_), .ZN(new_n9250_));
  NAND2_X1   g09058(.A1(new_n8793_), .A2(new_n8868_), .ZN(new_n9251_));
  OAI21_X1   g09059(.A1(new_n8826_), .A2(new_n9251_), .B(new_n8799_), .ZN(new_n9252_));
  NAND2_X1   g09060(.A1(new_n9252_), .A2(new_n9250_), .ZN(new_n9253_));
  NOR2_X1    g09061(.A1(new_n8869_), .A2(new_n8885_), .ZN(new_n9254_));
  NAND2_X1   g09062(.A1(\asqrt[27] ), .A2(new_n9254_), .ZN(new_n9255_));
  NAND3_X1   g09063(.A1(new_n9253_), .A2(new_n9249_), .A3(new_n9255_), .ZN(new_n9256_));
  AOI21_X1   g09064(.A1(new_n9248_), .A2(new_n9236_), .B(new_n9256_), .ZN(new_n9257_));
  NOR3_X1    g09065(.A1(new_n9245_), .A2(\asqrt[61] ), .A3(new_n9233_), .ZN(new_n9258_));
  OAI21_X1   g09066(.A1(new_n9229_), .A2(new_n9258_), .B(new_n9246_), .ZN(new_n9259_));
  AOI21_X1   g09067(.A1(new_n9259_), .A2(\asqrt[62] ), .B(new_n9253_), .ZN(new_n9260_));
  OAI21_X1   g09068(.A1(new_n8826_), .A2(new_n8885_), .B(new_n8869_), .ZN(new_n9261_));
  NOR2_X1    g09069(.A1(new_n9254_), .A2(new_n193_), .ZN(new_n9262_));
  NAND2_X1   g09070(.A1(new_n9261_), .A2(new_n9262_), .ZN(new_n9263_));
  INV_X1     g09071(.I(new_n9263_), .ZN(new_n9264_));
  AND3_X2    g09072(.A1(new_n8809_), .A2(new_n8807_), .A3(new_n8822_), .Z(new_n9265_));
  NAND4_X1   g09073(.A1(new_n9249_), .A2(new_n8870_), .A3(new_n8819_), .A4(new_n9265_), .ZN(new_n9266_));
  INV_X1     g09074(.I(new_n9266_), .ZN(new_n9267_));
  NOR2_X1    g09075(.A1(new_n9264_), .A2(new_n9267_), .ZN(new_n9268_));
  INV_X1     g09076(.I(new_n9268_), .ZN(new_n9269_));
  AOI21_X1   g09077(.A1(new_n9260_), .A2(new_n9248_), .B(new_n9269_), .ZN(new_n9270_));
  OAI21_X1   g09078(.A1(\asqrt[63] ), .A2(new_n9257_), .B(new_n9270_), .ZN(\asqrt[26] ));
  NOR2_X1    g09079(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n9272_));
  INV_X1     g09080(.I(new_n9272_), .ZN(new_n9273_));
  NOR2_X1    g09081(.A1(new_n9273_), .A2(\a[52] ), .ZN(new_n9274_));
  INV_X1     g09082(.I(new_n9274_), .ZN(new_n9275_));
  NAND2_X1   g09083(.A1(new_n9248_), .A2(new_n9236_), .ZN(new_n9276_));
  INV_X1     g09084(.I(new_n9256_), .ZN(new_n9277_));
  AOI21_X1   g09085(.A1(new_n9276_), .A2(new_n9277_), .B(\asqrt[63] ), .ZN(new_n9278_));
  INV_X1     g09086(.I(new_n9248_), .ZN(new_n9279_));
  INV_X1     g09087(.I(new_n9253_), .ZN(new_n9280_));
  NAND2_X1   g09088(.A1(new_n9236_), .A2(new_n9280_), .ZN(new_n9281_));
  OAI21_X1   g09089(.A1(new_n9279_), .A2(new_n9281_), .B(new_n9268_), .ZN(new_n9282_));
  OAI21_X1   g09090(.A1(new_n9278_), .A2(new_n9282_), .B(\a[52] ), .ZN(new_n9283_));
  AOI21_X1   g09091(.A1(new_n9283_), .A2(new_n9275_), .B(new_n8826_), .ZN(new_n9284_));
  INV_X1     g09092(.I(\a[52] ), .ZN(new_n9285_));
  INV_X1     g09093(.I(new_n9229_), .ZN(new_n9286_));
  NAND2_X1   g09094(.A1(new_n9211_), .A2(new_n218_), .ZN(new_n9287_));
  OAI21_X1   g09095(.A1(new_n9287_), .A2(new_n9245_), .B(new_n9286_), .ZN(new_n9288_));
  NAND3_X1   g09096(.A1(new_n9288_), .A2(new_n207_), .A3(new_n9246_), .ZN(new_n9289_));
  AOI22_X1   g09097(.A1(new_n9289_), .A2(new_n9241_), .B1(new_n9259_), .B2(\asqrt[62] ), .ZN(new_n9290_));
  OAI21_X1   g09098(.A1(new_n9290_), .A2(new_n9256_), .B(new_n193_), .ZN(new_n9291_));
  AOI21_X1   g09099(.A1(new_n9291_), .A2(new_n9270_), .B(new_n9285_), .ZN(new_n9292_));
  NAND4_X1   g09100(.A1(new_n9249_), .A2(new_n8819_), .A3(new_n8822_), .A4(new_n9275_), .ZN(new_n9293_));
  NOR2_X1    g09101(.A1(new_n9293_), .A2(new_n8883_), .ZN(new_n9294_));
  INV_X1     g09102(.I(new_n9294_), .ZN(new_n9295_));
  NOR2_X1    g09103(.A1(new_n9292_), .A2(new_n9295_), .ZN(new_n9296_));
  AOI21_X1   g09104(.A1(new_n9291_), .A2(new_n9270_), .B(new_n8828_), .ZN(new_n9297_));
  INV_X1     g09105(.I(\a[53] ), .ZN(new_n9298_));
  AOI21_X1   g09106(.A1(\asqrt[26] ), .A2(new_n9285_), .B(new_n9298_), .ZN(new_n9299_));
  NOR3_X1    g09107(.A1(new_n9296_), .A2(new_n9299_), .A3(new_n9297_), .ZN(new_n9300_));
  OAI21_X1   g09108(.A1(new_n9300_), .A2(new_n9284_), .B(\asqrt[28] ), .ZN(new_n9301_));
  OAI21_X1   g09109(.A1(new_n9278_), .A2(new_n9282_), .B(new_n8827_), .ZN(new_n9302_));
  NOR2_X1    g09110(.A1(new_n9279_), .A2(new_n9281_), .ZN(new_n9303_));
  NOR2_X1    g09111(.A1(new_n9267_), .A2(new_n8826_), .ZN(new_n9304_));
  NAND2_X1   g09112(.A1(new_n9263_), .A2(new_n9304_), .ZN(new_n9305_));
  NOR3_X1    g09113(.A1(new_n9278_), .A2(new_n9303_), .A3(new_n9305_), .ZN(new_n9306_));
  INV_X1     g09114(.I(new_n9306_), .ZN(new_n9307_));
  AOI21_X1   g09115(.A1(new_n9307_), .A2(new_n9302_), .B(new_n8830_), .ZN(new_n9308_));
  NOR3_X1    g09116(.A1(new_n9306_), .A2(new_n9297_), .A3(\a[54] ), .ZN(new_n9309_));
  AOI21_X1   g09117(.A1(\asqrt[26] ), .A2(\a[52] ), .B(new_n9274_), .ZN(new_n9310_));
  OAI21_X1   g09118(.A1(new_n9310_), .A2(new_n8826_), .B(new_n8483_), .ZN(new_n9311_));
  OAI22_X1   g09119(.A1(new_n9300_), .A2(new_n9311_), .B1(new_n9308_), .B2(new_n9309_), .ZN(new_n9312_));
  AOI21_X1   g09120(.A1(new_n9312_), .A2(new_n9301_), .B(new_n8036_), .ZN(new_n9313_));
  INV_X1     g09121(.I(new_n8905_), .ZN(new_n9314_));
  OAI21_X1   g09122(.A1(new_n8871_), .A2(new_n8876_), .B(new_n8872_), .ZN(new_n9315_));
  NOR2_X1    g09123(.A1(new_n9315_), .A2(new_n9314_), .ZN(new_n9316_));
  NOR2_X1    g09124(.A1(new_n9278_), .A2(new_n9282_), .ZN(new_n9317_));
  OR2_X2     g09125(.A1(new_n9317_), .A2(new_n9315_), .Z(new_n9318_));
  AOI22_X1   g09126(.A1(new_n9318_), .A2(new_n9314_), .B1(\asqrt[26] ), .B2(new_n9316_), .ZN(new_n9319_));
  OAI21_X1   g09127(.A1(new_n9292_), .A2(new_n9274_), .B(\asqrt[27] ), .ZN(new_n9320_));
  AOI21_X1   g09128(.A1(new_n9291_), .A2(new_n9270_), .B(\a[52] ), .ZN(new_n9321_));
  OAI21_X1   g09129(.A1(new_n9298_), .A2(new_n9321_), .B(new_n9302_), .ZN(new_n9322_));
  OAI21_X1   g09130(.A1(new_n9322_), .A2(new_n9296_), .B(new_n9320_), .ZN(new_n9323_));
  AOI21_X1   g09131(.A1(new_n9323_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n9324_));
  AOI21_X1   g09132(.A1(new_n9324_), .A2(new_n9312_), .B(new_n9319_), .ZN(new_n9325_));
  OAI21_X1   g09133(.A1(new_n9325_), .A2(new_n9313_), .B(\asqrt[30] ), .ZN(new_n9326_));
  INV_X1     g09134(.I(new_n9326_), .ZN(new_n9327_));
  NOR2_X1    g09135(.A1(new_n8895_), .A2(new_n8896_), .ZN(new_n9328_));
  NOR2_X1    g09136(.A1(new_n8881_), .A2(new_n8898_), .ZN(new_n9329_));
  INV_X1     g09137(.I(new_n9329_), .ZN(new_n9330_));
  NAND4_X1   g09138(.A1(\asqrt[26] ), .A2(new_n8882_), .A3(new_n9328_), .A4(new_n9330_), .ZN(new_n9331_));
  NAND2_X1   g09139(.A1(new_n9330_), .A2(new_n8882_), .ZN(new_n9332_));
  NOR2_X1    g09140(.A1(new_n9317_), .A2(new_n9332_), .ZN(new_n9333_));
  OAI21_X1   g09141(.A1(new_n9328_), .A2(new_n9333_), .B(new_n9331_), .ZN(new_n9334_));
  INV_X1     g09142(.I(new_n9334_), .ZN(new_n9335_));
  NOR3_X1    g09143(.A1(new_n9325_), .A2(new_n9313_), .A3(\asqrt[30] ), .ZN(new_n9336_));
  NOR2_X1    g09144(.A1(new_n9336_), .A2(new_n9335_), .ZN(new_n9337_));
  OAI21_X1   g09145(.A1(new_n9337_), .A2(new_n9327_), .B(\asqrt[31] ), .ZN(new_n9338_));
  INV_X1     g09146(.I(new_n8903_), .ZN(new_n9339_));
  INV_X1     g09147(.I(new_n8900_), .ZN(new_n9340_));
  NAND2_X1   g09148(.A1(new_n8907_), .A2(new_n8899_), .ZN(new_n9341_));
  NAND3_X1   g09149(.A1(\asqrt[26] ), .A2(new_n9340_), .A3(new_n9341_), .ZN(new_n9342_));
  AND3_X2    g09150(.A1(new_n9340_), .A2(new_n8903_), .A3(new_n9341_), .Z(new_n9343_));
  AOI22_X1   g09151(.A1(new_n9342_), .A2(new_n9339_), .B1(\asqrt[26] ), .B2(new_n9343_), .ZN(new_n9344_));
  INV_X1     g09152(.I(new_n9344_), .ZN(new_n9345_));
  NAND2_X1   g09153(.A1(new_n9326_), .A2(new_n7229_), .ZN(new_n9346_));
  OAI21_X1   g09154(.A1(new_n9337_), .A2(new_n9346_), .B(new_n9345_), .ZN(new_n9347_));
  AOI21_X1   g09155(.A1(new_n9347_), .A2(new_n9338_), .B(new_n6824_), .ZN(new_n9348_));
  INV_X1     g09156(.I(new_n8917_), .ZN(new_n9349_));
  NOR3_X1    g09157(.A1(new_n8910_), .A2(new_n9349_), .A3(new_n8918_), .ZN(new_n9350_));
  NOR3_X1    g09158(.A1(new_n9317_), .A2(new_n8910_), .A3(new_n8918_), .ZN(new_n9351_));
  INV_X1     g09159(.I(new_n9351_), .ZN(new_n9352_));
  AOI22_X1   g09160(.A1(new_n9352_), .A2(new_n9349_), .B1(\asqrt[26] ), .B2(new_n9350_), .ZN(new_n9353_));
  OAI21_X1   g09161(.A1(new_n9335_), .A2(new_n9336_), .B(new_n9326_), .ZN(new_n9354_));
  AOI21_X1   g09162(.A1(new_n9354_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n9355_));
  AOI21_X1   g09163(.A1(new_n9355_), .A2(new_n9347_), .B(new_n9353_), .ZN(new_n9356_));
  OAI21_X1   g09164(.A1(new_n9356_), .A2(new_n9348_), .B(\asqrt[33] ), .ZN(new_n9357_));
  INV_X1     g09165(.I(new_n9357_), .ZN(new_n9358_));
  INV_X1     g09166(.I(new_n8919_), .ZN(new_n9359_));
  INV_X1     g09167(.I(new_n8927_), .ZN(new_n9360_));
  NAND2_X1   g09168(.A1(new_n9359_), .A2(new_n9360_), .ZN(new_n9361_));
  NAND3_X1   g09169(.A1(\asqrt[26] ), .A2(new_n8920_), .A3(new_n9361_), .ZN(new_n9362_));
  AND3_X2    g09170(.A1(new_n9361_), .A2(new_n8920_), .A3(new_n8925_), .Z(new_n9363_));
  AOI22_X1   g09171(.A1(new_n9362_), .A2(new_n8926_), .B1(\asqrt[26] ), .B2(new_n9363_), .ZN(new_n9364_));
  NOR3_X1    g09172(.A1(new_n9356_), .A2(new_n9348_), .A3(\asqrt[33] ), .ZN(new_n9365_));
  NOR2_X1    g09173(.A1(new_n9365_), .A2(new_n9364_), .ZN(new_n9366_));
  OAI21_X1   g09174(.A1(new_n9366_), .A2(new_n9358_), .B(\asqrt[34] ), .ZN(new_n9367_));
  INV_X1     g09175(.I(new_n8933_), .ZN(new_n9368_));
  INV_X1     g09176(.I(new_n8928_), .ZN(new_n9369_));
  INV_X1     g09177(.I(new_n8935_), .ZN(new_n9370_));
  OAI21_X1   g09178(.A1(new_n9370_), .A2(new_n9369_), .B(new_n8933_), .ZN(new_n9371_));
  NOR2_X1    g09179(.A1(new_n9371_), .A2(new_n8929_), .ZN(new_n9372_));
  NOR2_X1    g09180(.A1(new_n9370_), .A2(new_n9369_), .ZN(new_n9373_));
  NOR3_X1    g09181(.A1(new_n9317_), .A2(new_n8929_), .A3(new_n9373_), .ZN(new_n9374_));
  INV_X1     g09182(.I(new_n9374_), .ZN(new_n9375_));
  AOI22_X1   g09183(.A1(new_n9375_), .A2(new_n9368_), .B1(\asqrt[26] ), .B2(new_n9372_), .ZN(new_n9376_));
  INV_X1     g09184(.I(new_n9376_), .ZN(new_n9377_));
  NAND2_X1   g09185(.A1(new_n9357_), .A2(new_n6077_), .ZN(new_n9378_));
  OAI21_X1   g09186(.A1(new_n9366_), .A2(new_n9378_), .B(new_n9377_), .ZN(new_n9379_));
  AOI21_X1   g09187(.A1(new_n9379_), .A2(new_n9367_), .B(new_n5708_), .ZN(new_n9380_));
  INV_X1     g09188(.I(new_n8943_), .ZN(new_n9381_));
  NOR3_X1    g09189(.A1(new_n9317_), .A2(new_n8938_), .A3(new_n8944_), .ZN(new_n9382_));
  INV_X1     g09190(.I(new_n9382_), .ZN(new_n9383_));
  NOR3_X1    g09191(.A1(new_n8938_), .A2(new_n9381_), .A3(new_n8944_), .ZN(new_n9384_));
  AOI22_X1   g09192(.A1(new_n9383_), .A2(new_n9381_), .B1(\asqrt[26] ), .B2(new_n9384_), .ZN(new_n9385_));
  OAI21_X1   g09193(.A1(new_n9364_), .A2(new_n9365_), .B(new_n9357_), .ZN(new_n9386_));
  AOI21_X1   g09194(.A1(new_n9386_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n9387_));
  AOI21_X1   g09195(.A1(new_n9387_), .A2(new_n9379_), .B(new_n9385_), .ZN(new_n9388_));
  OAI21_X1   g09196(.A1(new_n9388_), .A2(new_n9380_), .B(\asqrt[36] ), .ZN(new_n9389_));
  INV_X1     g09197(.I(new_n9389_), .ZN(new_n9390_));
  NOR2_X1    g09198(.A1(new_n8945_), .A2(new_n8953_), .ZN(new_n9391_));
  INV_X1     g09199(.I(new_n9391_), .ZN(new_n9392_));
  AND3_X2    g09200(.A1(new_n9392_), .A2(new_n8946_), .A3(new_n8951_), .Z(new_n9393_));
  NAND3_X1   g09201(.A1(\asqrt[26] ), .A2(new_n8946_), .A3(new_n9392_), .ZN(new_n9394_));
  AOI22_X1   g09202(.A1(new_n9394_), .A2(new_n8952_), .B1(\asqrt[26] ), .B2(new_n9393_), .ZN(new_n9395_));
  NOR3_X1    g09203(.A1(new_n9388_), .A2(new_n9380_), .A3(\asqrt[36] ), .ZN(new_n9396_));
  NOR2_X1    g09204(.A1(new_n9396_), .A2(new_n9395_), .ZN(new_n9397_));
  OAI21_X1   g09205(.A1(new_n9397_), .A2(new_n9390_), .B(\asqrt[37] ), .ZN(new_n9398_));
  INV_X1     g09206(.I(new_n8959_), .ZN(new_n9399_));
  INV_X1     g09207(.I(new_n8954_), .ZN(new_n9400_));
  INV_X1     g09208(.I(new_n8961_), .ZN(new_n9401_));
  NOR2_X1    g09209(.A1(new_n9401_), .A2(new_n9400_), .ZN(new_n9402_));
  NOR3_X1    g09210(.A1(new_n9317_), .A2(new_n8955_), .A3(new_n9402_), .ZN(new_n9403_));
  INV_X1     g09211(.I(new_n9403_), .ZN(new_n9404_));
  NOR3_X1    g09212(.A1(new_n9402_), .A2(new_n8955_), .A3(new_n9399_), .ZN(new_n9405_));
  AOI22_X1   g09213(.A1(new_n9404_), .A2(new_n9399_), .B1(\asqrt[26] ), .B2(new_n9405_), .ZN(new_n9406_));
  INV_X1     g09214(.I(new_n9406_), .ZN(new_n9407_));
  NAND2_X1   g09215(.A1(new_n9389_), .A2(new_n5024_), .ZN(new_n9408_));
  OAI21_X1   g09216(.A1(new_n9397_), .A2(new_n9408_), .B(new_n9407_), .ZN(new_n9409_));
  AOI21_X1   g09217(.A1(new_n9409_), .A2(new_n9398_), .B(new_n4696_), .ZN(new_n9410_));
  INV_X1     g09218(.I(new_n8969_), .ZN(new_n9411_));
  NOR3_X1    g09219(.A1(new_n8964_), .A2(new_n8970_), .A3(new_n9411_), .ZN(new_n9412_));
  NOR3_X1    g09220(.A1(new_n9317_), .A2(new_n8964_), .A3(new_n8970_), .ZN(new_n9413_));
  INV_X1     g09221(.I(new_n9413_), .ZN(new_n9414_));
  AOI22_X1   g09222(.A1(new_n9414_), .A2(new_n9411_), .B1(\asqrt[26] ), .B2(new_n9412_), .ZN(new_n9415_));
  OAI21_X1   g09223(.A1(new_n9395_), .A2(new_n9396_), .B(new_n9389_), .ZN(new_n9416_));
  AOI21_X1   g09224(.A1(new_n9416_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n9417_));
  AOI21_X1   g09225(.A1(new_n9417_), .A2(new_n9409_), .B(new_n9415_), .ZN(new_n9418_));
  OAI21_X1   g09226(.A1(new_n9418_), .A2(new_n9410_), .B(\asqrt[39] ), .ZN(new_n9419_));
  INV_X1     g09227(.I(new_n9419_), .ZN(new_n9420_));
  INV_X1     g09228(.I(new_n8972_), .ZN(new_n9421_));
  NOR2_X1    g09229(.A1(new_n8971_), .A2(new_n8979_), .ZN(new_n9422_));
  NOR3_X1    g09230(.A1(new_n9317_), .A2(new_n9421_), .A3(new_n9422_), .ZN(new_n9423_));
  INV_X1     g09231(.I(new_n9423_), .ZN(new_n9424_));
  NOR3_X1    g09232(.A1(new_n9421_), .A2(new_n8978_), .A3(new_n9422_), .ZN(new_n9425_));
  AOI22_X1   g09233(.A1(new_n9424_), .A2(new_n8978_), .B1(\asqrt[26] ), .B2(new_n9425_), .ZN(new_n9426_));
  NOR3_X1    g09234(.A1(new_n9418_), .A2(new_n9410_), .A3(\asqrt[39] ), .ZN(new_n9427_));
  NOR2_X1    g09235(.A1(new_n9427_), .A2(new_n9426_), .ZN(new_n9428_));
  OAI21_X1   g09236(.A1(new_n9428_), .A2(new_n9420_), .B(\asqrt[40] ), .ZN(new_n9429_));
  INV_X1     g09237(.I(new_n8985_), .ZN(new_n9430_));
  INV_X1     g09238(.I(new_n8980_), .ZN(new_n9431_));
  INV_X1     g09239(.I(new_n8987_), .ZN(new_n9432_));
  NOR2_X1    g09240(.A1(new_n9432_), .A2(new_n9431_), .ZN(new_n9433_));
  NOR3_X1    g09241(.A1(new_n9433_), .A2(new_n8981_), .A3(new_n9430_), .ZN(new_n9434_));
  NOR3_X1    g09242(.A1(new_n9317_), .A2(new_n8981_), .A3(new_n9433_), .ZN(new_n9435_));
  INV_X1     g09243(.I(new_n9435_), .ZN(new_n9436_));
  AOI22_X1   g09244(.A1(new_n9436_), .A2(new_n9430_), .B1(\asqrt[26] ), .B2(new_n9434_), .ZN(new_n9437_));
  INV_X1     g09245(.I(new_n9437_), .ZN(new_n9438_));
  NAND2_X1   g09246(.A1(new_n9419_), .A2(new_n4071_), .ZN(new_n9439_));
  OAI21_X1   g09247(.A1(new_n9428_), .A2(new_n9439_), .B(new_n9438_), .ZN(new_n9440_));
  AOI21_X1   g09248(.A1(new_n9440_), .A2(new_n9429_), .B(new_n3782_), .ZN(new_n9441_));
  INV_X1     g09249(.I(new_n8995_), .ZN(new_n9442_));
  NOR3_X1    g09250(.A1(new_n9317_), .A2(new_n8990_), .A3(new_n8996_), .ZN(new_n9443_));
  INV_X1     g09251(.I(new_n9443_), .ZN(new_n9444_));
  NOR3_X1    g09252(.A1(new_n8990_), .A2(new_n8996_), .A3(new_n9442_), .ZN(new_n9445_));
  AOI22_X1   g09253(.A1(new_n9444_), .A2(new_n9442_), .B1(\asqrt[26] ), .B2(new_n9445_), .ZN(new_n9446_));
  OAI21_X1   g09254(.A1(new_n9426_), .A2(new_n9427_), .B(new_n9419_), .ZN(new_n9447_));
  AOI21_X1   g09255(.A1(new_n9447_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n9448_));
  AOI21_X1   g09256(.A1(new_n9448_), .A2(new_n9440_), .B(new_n9446_), .ZN(new_n9449_));
  OAI21_X1   g09257(.A1(new_n9449_), .A2(new_n9441_), .B(\asqrt[42] ), .ZN(new_n9450_));
  INV_X1     g09258(.I(new_n9450_), .ZN(new_n9451_));
  NOR2_X1    g09259(.A1(new_n8997_), .A2(new_n9005_), .ZN(new_n9452_));
  INV_X1     g09260(.I(new_n9452_), .ZN(new_n9453_));
  AND3_X2    g09261(.A1(new_n9453_), .A2(new_n8998_), .A3(new_n9003_), .Z(new_n9454_));
  NAND3_X1   g09262(.A1(\asqrt[26] ), .A2(new_n8998_), .A3(new_n9453_), .ZN(new_n9455_));
  AOI22_X1   g09263(.A1(new_n9455_), .A2(new_n9004_), .B1(\asqrt[26] ), .B2(new_n9454_), .ZN(new_n9456_));
  NOR3_X1    g09264(.A1(new_n9449_), .A2(new_n9441_), .A3(\asqrt[42] ), .ZN(new_n9457_));
  NOR2_X1    g09265(.A1(new_n9457_), .A2(new_n9456_), .ZN(new_n9458_));
  OAI21_X1   g09266(.A1(new_n9458_), .A2(new_n9451_), .B(\asqrt[43] ), .ZN(new_n9459_));
  INV_X1     g09267(.I(new_n9011_), .ZN(new_n9460_));
  INV_X1     g09268(.I(new_n9007_), .ZN(new_n9461_));
  NAND2_X1   g09269(.A1(new_n9013_), .A2(new_n9006_), .ZN(new_n9462_));
  NAND3_X1   g09270(.A1(\asqrt[26] ), .A2(new_n9461_), .A3(new_n9462_), .ZN(new_n9463_));
  AND3_X2    g09271(.A1(new_n9461_), .A2(new_n9011_), .A3(new_n9462_), .Z(new_n9464_));
  AOI22_X1   g09272(.A1(new_n9463_), .A2(new_n9460_), .B1(\asqrt[26] ), .B2(new_n9464_), .ZN(new_n9465_));
  INV_X1     g09273(.I(new_n9465_), .ZN(new_n9466_));
  NAND2_X1   g09274(.A1(new_n9450_), .A2(new_n3218_), .ZN(new_n9467_));
  OAI21_X1   g09275(.A1(new_n9458_), .A2(new_n9467_), .B(new_n9466_), .ZN(new_n9468_));
  AOI21_X1   g09276(.A1(new_n9468_), .A2(new_n9459_), .B(new_n2954_), .ZN(new_n9469_));
  INV_X1     g09277(.I(new_n9023_), .ZN(new_n9470_));
  NOR3_X1    g09278(.A1(new_n9016_), .A2(new_n9024_), .A3(new_n9470_), .ZN(new_n9471_));
  NOR3_X1    g09279(.A1(new_n9317_), .A2(new_n9016_), .A3(new_n9024_), .ZN(new_n9472_));
  INV_X1     g09280(.I(new_n9472_), .ZN(new_n9473_));
  AOI22_X1   g09281(.A1(new_n9473_), .A2(new_n9470_), .B1(\asqrt[26] ), .B2(new_n9471_), .ZN(new_n9474_));
  OAI21_X1   g09282(.A1(new_n9456_), .A2(new_n9457_), .B(new_n9450_), .ZN(new_n9475_));
  AOI21_X1   g09283(.A1(new_n9475_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n9476_));
  AOI21_X1   g09284(.A1(new_n9476_), .A2(new_n9468_), .B(new_n9474_), .ZN(new_n9477_));
  OAI21_X1   g09285(.A1(new_n9477_), .A2(new_n9469_), .B(\asqrt[45] ), .ZN(new_n9478_));
  INV_X1     g09286(.I(new_n9478_), .ZN(new_n9479_));
  OAI21_X1   g09287(.A1(new_n9025_), .A2(new_n9032_), .B(new_n9026_), .ZN(new_n9480_));
  NOR2_X1    g09288(.A1(new_n9317_), .A2(new_n9480_), .ZN(new_n9481_));
  INV_X1     g09289(.I(new_n9481_), .ZN(new_n9482_));
  NOR2_X1    g09290(.A1(new_n9025_), .A2(new_n9032_), .ZN(new_n9483_));
  NAND2_X1   g09291(.A1(new_n9026_), .A2(new_n9030_), .ZN(new_n9484_));
  NOR2_X1    g09292(.A1(new_n9484_), .A2(new_n9483_), .ZN(new_n9485_));
  AOI22_X1   g09293(.A1(new_n9482_), .A2(new_n9031_), .B1(\asqrt[26] ), .B2(new_n9485_), .ZN(new_n9486_));
  NOR3_X1    g09294(.A1(new_n9477_), .A2(new_n9469_), .A3(\asqrt[45] ), .ZN(new_n9487_));
  NOR2_X1    g09295(.A1(new_n9487_), .A2(new_n9486_), .ZN(new_n9488_));
  OAI21_X1   g09296(.A1(new_n9488_), .A2(new_n9479_), .B(\asqrt[46] ), .ZN(new_n9489_));
  INV_X1     g09297(.I(new_n9040_), .ZN(new_n9490_));
  INV_X1     g09298(.I(new_n9034_), .ZN(new_n9491_));
  NAND2_X1   g09299(.A1(new_n9042_), .A2(new_n9033_), .ZN(new_n9492_));
  AND3_X2    g09300(.A1(new_n9491_), .A2(new_n9040_), .A3(new_n9492_), .Z(new_n9493_));
  NAND3_X1   g09301(.A1(\asqrt[26] ), .A2(new_n9491_), .A3(new_n9492_), .ZN(new_n9494_));
  AOI22_X1   g09302(.A1(new_n9494_), .A2(new_n9490_), .B1(\asqrt[26] ), .B2(new_n9493_), .ZN(new_n9495_));
  INV_X1     g09303(.I(new_n9495_), .ZN(new_n9496_));
  NAND2_X1   g09304(.A1(new_n9478_), .A2(new_n2465_), .ZN(new_n9497_));
  OAI21_X1   g09305(.A1(new_n9488_), .A2(new_n9497_), .B(new_n9496_), .ZN(new_n9498_));
  AOI21_X1   g09306(.A1(new_n9498_), .A2(new_n9489_), .B(new_n2229_), .ZN(new_n9499_));
  INV_X1     g09307(.I(new_n9053_), .ZN(new_n9500_));
  NOR3_X1    g09308(.A1(new_n9317_), .A2(new_n9045_), .A3(new_n9054_), .ZN(new_n9501_));
  INV_X1     g09309(.I(new_n9501_), .ZN(new_n9502_));
  NOR3_X1    g09310(.A1(new_n9045_), .A2(new_n9500_), .A3(new_n9054_), .ZN(new_n9503_));
  AOI22_X1   g09311(.A1(new_n9502_), .A2(new_n9500_), .B1(\asqrt[26] ), .B2(new_n9503_), .ZN(new_n9504_));
  OAI21_X1   g09312(.A1(new_n9486_), .A2(new_n9487_), .B(new_n9478_), .ZN(new_n9505_));
  AOI21_X1   g09313(.A1(new_n9505_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n9506_));
  AOI21_X1   g09314(.A1(new_n9506_), .A2(new_n9498_), .B(new_n9504_), .ZN(new_n9507_));
  OAI21_X1   g09315(.A1(new_n9507_), .A2(new_n9499_), .B(\asqrt[48] ), .ZN(new_n9508_));
  INV_X1     g09316(.I(new_n9508_), .ZN(new_n9509_));
  OR2_X2     g09317(.A1(new_n9055_), .A2(new_n9062_), .Z(new_n9510_));
  AND3_X2    g09318(.A1(new_n9510_), .A2(new_n9056_), .A3(new_n9060_), .Z(new_n9511_));
  NAND3_X1   g09319(.A1(\asqrt[26] ), .A2(new_n9056_), .A3(new_n9510_), .ZN(new_n9512_));
  AOI22_X1   g09320(.A1(new_n9512_), .A2(new_n9061_), .B1(\asqrt[26] ), .B2(new_n9511_), .ZN(new_n9513_));
  NOR3_X1    g09321(.A1(new_n9507_), .A2(new_n9499_), .A3(\asqrt[48] ), .ZN(new_n9514_));
  NOR2_X1    g09322(.A1(new_n9514_), .A2(new_n9513_), .ZN(new_n9515_));
  OAI21_X1   g09323(.A1(new_n9515_), .A2(new_n9509_), .B(\asqrt[49] ), .ZN(new_n9516_));
  INV_X1     g09324(.I(new_n9070_), .ZN(new_n9517_));
  NAND2_X1   g09325(.A1(new_n9072_), .A2(new_n9063_), .ZN(new_n9518_));
  NAND3_X1   g09326(.A1(\asqrt[26] ), .A2(new_n9115_), .A3(new_n9518_), .ZN(new_n9519_));
  AND3_X2    g09327(.A1(new_n9115_), .A2(new_n9070_), .A3(new_n9518_), .Z(new_n9520_));
  AOI22_X1   g09328(.A1(new_n9519_), .A2(new_n9517_), .B1(\asqrt[26] ), .B2(new_n9520_), .ZN(new_n9521_));
  INV_X1     g09329(.I(new_n9521_), .ZN(new_n9522_));
  NAND2_X1   g09330(.A1(new_n9508_), .A2(new_n1806_), .ZN(new_n9523_));
  OAI21_X1   g09331(.A1(new_n9515_), .A2(new_n9523_), .B(new_n9522_), .ZN(new_n9524_));
  AOI21_X1   g09332(.A1(new_n9524_), .A2(new_n9516_), .B(new_n1612_), .ZN(new_n9525_));
  NOR3_X1    g09333(.A1(new_n9075_), .A2(new_n9114_), .A3(new_n9084_), .ZN(new_n9526_));
  NOR3_X1    g09334(.A1(new_n9317_), .A2(new_n9075_), .A3(new_n9084_), .ZN(new_n9527_));
  INV_X1     g09335(.I(new_n9527_), .ZN(new_n9528_));
  AOI22_X1   g09336(.A1(new_n9528_), .A2(new_n9114_), .B1(\asqrt[26] ), .B2(new_n9526_), .ZN(new_n9529_));
  OAI21_X1   g09337(.A1(new_n9513_), .A2(new_n9514_), .B(new_n9508_), .ZN(new_n9530_));
  AOI21_X1   g09338(.A1(new_n9530_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n9531_));
  AOI21_X1   g09339(.A1(new_n9531_), .A2(new_n9524_), .B(new_n9529_), .ZN(new_n9532_));
  OAI21_X1   g09340(.A1(new_n9532_), .A2(new_n9525_), .B(\asqrt[51] ), .ZN(new_n9533_));
  NOR2_X1    g09341(.A1(new_n9085_), .A2(new_n9092_), .ZN(new_n9534_));
  NOR3_X1    g09342(.A1(new_n9317_), .A2(new_n9118_), .A3(new_n9534_), .ZN(new_n9535_));
  INV_X1     g09343(.I(new_n9535_), .ZN(new_n9536_));
  NOR3_X1    g09344(.A1(new_n9118_), .A2(new_n9534_), .A3(new_n9091_), .ZN(new_n9537_));
  AOI22_X1   g09345(.A1(new_n9536_), .A2(new_n9091_), .B1(\asqrt[26] ), .B2(new_n9537_), .ZN(new_n9538_));
  INV_X1     g09346(.I(new_n9538_), .ZN(new_n9539_));
  INV_X1     g09347(.I(new_n9513_), .ZN(new_n9540_));
  INV_X1     g09348(.I(new_n9486_), .ZN(new_n9541_));
  INV_X1     g09349(.I(new_n9456_), .ZN(new_n9542_));
  INV_X1     g09350(.I(new_n9426_), .ZN(new_n9543_));
  INV_X1     g09351(.I(new_n9395_), .ZN(new_n9544_));
  INV_X1     g09352(.I(new_n9364_), .ZN(new_n9545_));
  NAND2_X1   g09353(.A1(new_n9283_), .A2(new_n9294_), .ZN(new_n9546_));
  OAI21_X1   g09354(.A1(new_n9278_), .A2(new_n9282_), .B(new_n9285_), .ZN(new_n9547_));
  NAND2_X1   g09355(.A1(new_n9547_), .A2(\a[53] ), .ZN(new_n9548_));
  NAND3_X1   g09356(.A1(new_n9546_), .A2(new_n9548_), .A3(new_n9302_), .ZN(new_n9549_));
  AOI21_X1   g09357(.A1(new_n9549_), .A2(new_n9320_), .B(new_n8483_), .ZN(new_n9550_));
  OAI21_X1   g09358(.A1(new_n9306_), .A2(new_n9297_), .B(\a[54] ), .ZN(new_n9551_));
  NAND3_X1   g09359(.A1(new_n9307_), .A2(new_n9302_), .A3(new_n8830_), .ZN(new_n9552_));
  NAND2_X1   g09360(.A1(new_n9283_), .A2(new_n9275_), .ZN(new_n9553_));
  AOI21_X1   g09361(.A1(new_n9553_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n9554_));
  AOI22_X1   g09362(.A1(new_n9549_), .A2(new_n9554_), .B1(new_n9551_), .B2(new_n9552_), .ZN(new_n9555_));
  OAI21_X1   g09363(.A1(new_n9555_), .A2(new_n9550_), .B(\asqrt[29] ), .ZN(new_n9556_));
  NAND2_X1   g09364(.A1(new_n9556_), .A2(new_n7539_), .ZN(new_n9557_));
  OAI21_X1   g09365(.A1(new_n9557_), .A2(new_n9325_), .B(new_n9334_), .ZN(new_n9558_));
  AOI21_X1   g09366(.A1(new_n9558_), .A2(new_n9326_), .B(new_n7229_), .ZN(new_n9559_));
  NAND2_X1   g09367(.A1(\asqrt[26] ), .A2(new_n9316_), .ZN(new_n9560_));
  NAND2_X1   g09368(.A1(new_n9318_), .A2(new_n9314_), .ZN(new_n9561_));
  NAND2_X1   g09369(.A1(new_n9561_), .A2(new_n9560_), .ZN(new_n9562_));
  AOI21_X1   g09370(.A1(\a[53] ), .A2(new_n9547_), .B(new_n9297_), .ZN(new_n9563_));
  AOI21_X1   g09371(.A1(new_n9563_), .A2(new_n9546_), .B(new_n9284_), .ZN(new_n9564_));
  OAI21_X1   g09372(.A1(new_n9564_), .A2(new_n8483_), .B(new_n8036_), .ZN(new_n9565_));
  OAI21_X1   g09373(.A1(new_n9565_), .A2(new_n9555_), .B(new_n9562_), .ZN(new_n9566_));
  NAND2_X1   g09374(.A1(new_n9566_), .A2(new_n9556_), .ZN(new_n9567_));
  AOI21_X1   g09375(.A1(new_n9567_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n9568_));
  AOI21_X1   g09376(.A1(new_n9568_), .A2(new_n9558_), .B(new_n9344_), .ZN(new_n9569_));
  OAI21_X1   g09377(.A1(new_n9569_), .A2(new_n9559_), .B(\asqrt[32] ), .ZN(new_n9570_));
  NAND2_X1   g09378(.A1(new_n9570_), .A2(new_n6356_), .ZN(new_n9571_));
  OAI21_X1   g09379(.A1(new_n9571_), .A2(new_n9356_), .B(new_n9545_), .ZN(new_n9572_));
  NAND3_X1   g09380(.A1(new_n9572_), .A2(new_n6077_), .A3(new_n9357_), .ZN(new_n9573_));
  AOI22_X1   g09381(.A1(new_n9573_), .A2(new_n9377_), .B1(new_n9386_), .B2(\asqrt[34] ), .ZN(new_n9574_));
  OAI21_X1   g09382(.A1(new_n9574_), .A2(new_n5708_), .B(new_n5277_), .ZN(new_n9575_));
  OAI21_X1   g09383(.A1(new_n9575_), .A2(new_n9388_), .B(new_n9544_), .ZN(new_n9576_));
  AOI21_X1   g09384(.A1(new_n9576_), .A2(new_n9389_), .B(new_n5024_), .ZN(new_n9577_));
  AOI21_X1   g09385(.A1(new_n9572_), .A2(new_n9357_), .B(new_n6077_), .ZN(new_n9578_));
  NOR3_X1    g09386(.A1(new_n9569_), .A2(new_n9559_), .A3(\asqrt[32] ), .ZN(new_n9579_));
  OAI21_X1   g09387(.A1(new_n9353_), .A2(new_n9579_), .B(new_n9570_), .ZN(new_n9580_));
  AOI21_X1   g09388(.A1(new_n9580_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n9581_));
  AOI21_X1   g09389(.A1(new_n9581_), .A2(new_n9572_), .B(new_n9376_), .ZN(new_n9582_));
  NOR3_X1    g09390(.A1(new_n9582_), .A2(\asqrt[35] ), .A3(new_n9578_), .ZN(new_n9583_));
  OAI22_X1   g09391(.A1(new_n9583_), .A2(new_n9385_), .B1(new_n9574_), .B2(new_n5708_), .ZN(new_n9584_));
  AOI21_X1   g09392(.A1(new_n9584_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n9585_));
  AOI21_X1   g09393(.A1(new_n9585_), .A2(new_n9576_), .B(new_n9406_), .ZN(new_n9586_));
  OAI21_X1   g09394(.A1(new_n9586_), .A2(new_n9577_), .B(\asqrt[38] ), .ZN(new_n9587_));
  NAND2_X1   g09395(.A1(new_n9587_), .A2(new_n4298_), .ZN(new_n9588_));
  OAI21_X1   g09396(.A1(new_n9588_), .A2(new_n9418_), .B(new_n9543_), .ZN(new_n9589_));
  AOI21_X1   g09397(.A1(new_n9589_), .A2(new_n9419_), .B(new_n4071_), .ZN(new_n9590_));
  NOR3_X1    g09398(.A1(new_n9586_), .A2(\asqrt[38] ), .A3(new_n9577_), .ZN(new_n9591_));
  OAI21_X1   g09399(.A1(new_n9415_), .A2(new_n9591_), .B(new_n9587_), .ZN(new_n9592_));
  AOI21_X1   g09400(.A1(new_n9592_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n9593_));
  AOI21_X1   g09401(.A1(new_n9593_), .A2(new_n9589_), .B(new_n9437_), .ZN(new_n9594_));
  OAI21_X1   g09402(.A1(new_n9594_), .A2(new_n9590_), .B(\asqrt[41] ), .ZN(new_n9595_));
  NAND2_X1   g09403(.A1(new_n9595_), .A2(new_n3419_), .ZN(new_n9596_));
  OAI21_X1   g09404(.A1(new_n9596_), .A2(new_n9449_), .B(new_n9542_), .ZN(new_n9597_));
  AOI21_X1   g09405(.A1(new_n9597_), .A2(new_n9450_), .B(new_n3218_), .ZN(new_n9598_));
  NOR3_X1    g09406(.A1(new_n9594_), .A2(\asqrt[41] ), .A3(new_n9590_), .ZN(new_n9599_));
  OAI21_X1   g09407(.A1(new_n9446_), .A2(new_n9599_), .B(new_n9595_), .ZN(new_n9600_));
  AOI21_X1   g09408(.A1(new_n9600_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n9601_));
  AOI21_X1   g09409(.A1(new_n9601_), .A2(new_n9597_), .B(new_n9465_), .ZN(new_n9602_));
  OAI21_X1   g09410(.A1(new_n9602_), .A2(new_n9598_), .B(\asqrt[44] ), .ZN(new_n9603_));
  NAND2_X1   g09411(.A1(new_n9603_), .A2(new_n2641_), .ZN(new_n9604_));
  OAI21_X1   g09412(.A1(new_n9604_), .A2(new_n9477_), .B(new_n9541_), .ZN(new_n9605_));
  AOI21_X1   g09413(.A1(new_n9605_), .A2(new_n9478_), .B(new_n2465_), .ZN(new_n9606_));
  NOR3_X1    g09414(.A1(new_n9602_), .A2(\asqrt[44] ), .A3(new_n9598_), .ZN(new_n9607_));
  OAI21_X1   g09415(.A1(new_n9474_), .A2(new_n9607_), .B(new_n9603_), .ZN(new_n9608_));
  AOI21_X1   g09416(.A1(new_n9608_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n9609_));
  AOI21_X1   g09417(.A1(new_n9609_), .A2(new_n9605_), .B(new_n9495_), .ZN(new_n9610_));
  OAI21_X1   g09418(.A1(new_n9610_), .A2(new_n9606_), .B(\asqrt[47] ), .ZN(new_n9611_));
  NAND2_X1   g09419(.A1(new_n9611_), .A2(new_n1956_), .ZN(new_n9612_));
  OAI21_X1   g09420(.A1(new_n9612_), .A2(new_n9507_), .B(new_n9540_), .ZN(new_n9613_));
  AOI21_X1   g09421(.A1(new_n9613_), .A2(new_n9508_), .B(new_n1806_), .ZN(new_n9614_));
  NOR3_X1    g09422(.A1(new_n9610_), .A2(\asqrt[47] ), .A3(new_n9606_), .ZN(new_n9615_));
  OAI21_X1   g09423(.A1(new_n9504_), .A2(new_n9615_), .B(new_n9611_), .ZN(new_n9616_));
  AOI21_X1   g09424(.A1(new_n9616_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n9617_));
  AOI21_X1   g09425(.A1(new_n9617_), .A2(new_n9613_), .B(new_n9521_), .ZN(new_n9618_));
  OAI21_X1   g09426(.A1(new_n9618_), .A2(new_n9614_), .B(\asqrt[50] ), .ZN(new_n9619_));
  NAND2_X1   g09427(.A1(new_n9619_), .A2(new_n1376_), .ZN(new_n9620_));
  OAI21_X1   g09428(.A1(new_n9620_), .A2(new_n9532_), .B(new_n9539_), .ZN(new_n9621_));
  AOI21_X1   g09429(.A1(new_n9621_), .A2(new_n9533_), .B(new_n1256_), .ZN(new_n9622_));
  NOR2_X1    g09430(.A1(new_n9130_), .A2(new_n9120_), .ZN(new_n9623_));
  NOR3_X1    g09431(.A1(new_n9623_), .A2(new_n9094_), .A3(new_n9129_), .ZN(new_n9624_));
  NOR3_X1    g09432(.A1(new_n9317_), .A2(new_n9094_), .A3(new_n9623_), .ZN(new_n9625_));
  INV_X1     g09433(.I(new_n9625_), .ZN(new_n9626_));
  AOI22_X1   g09434(.A1(new_n9626_), .A2(new_n9129_), .B1(\asqrt[26] ), .B2(new_n9624_), .ZN(new_n9627_));
  NOR3_X1    g09435(.A1(new_n9618_), .A2(\asqrt[50] ), .A3(new_n9614_), .ZN(new_n9628_));
  OAI21_X1   g09436(.A1(new_n9529_), .A2(new_n9628_), .B(new_n9619_), .ZN(new_n9629_));
  AOI21_X1   g09437(.A1(new_n9629_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n9630_));
  AOI21_X1   g09438(.A1(new_n9630_), .A2(new_n9621_), .B(new_n9627_), .ZN(new_n9631_));
  OAI21_X1   g09439(.A1(new_n9631_), .A2(new_n9622_), .B(\asqrt[53] ), .ZN(new_n9632_));
  NOR3_X1    g09440(.A1(new_n9317_), .A2(new_n9132_), .A3(new_n9166_), .ZN(new_n9633_));
  INV_X1     g09441(.I(new_n9633_), .ZN(new_n9634_));
  NOR3_X1    g09442(.A1(new_n9132_), .A2(new_n9166_), .A3(new_n9113_), .ZN(new_n9635_));
  AOI22_X1   g09443(.A1(new_n9634_), .A2(new_n9113_), .B1(\asqrt[26] ), .B2(new_n9635_), .ZN(new_n9636_));
  INV_X1     g09444(.I(new_n9636_), .ZN(new_n9637_));
  INV_X1     g09445(.I(new_n9529_), .ZN(new_n9638_));
  NAND2_X1   g09446(.A1(new_n9516_), .A2(new_n1612_), .ZN(new_n9639_));
  OAI21_X1   g09447(.A1(new_n9639_), .A2(new_n9618_), .B(new_n9638_), .ZN(new_n9640_));
  AOI21_X1   g09448(.A1(new_n9640_), .A2(new_n9619_), .B(new_n1376_), .ZN(new_n9641_));
  NOR2_X1    g09449(.A1(new_n9525_), .A2(\asqrt[51] ), .ZN(new_n9642_));
  AOI21_X1   g09450(.A1(new_n9642_), .A2(new_n9640_), .B(new_n9538_), .ZN(new_n9643_));
  OAI21_X1   g09451(.A1(new_n9643_), .A2(new_n9641_), .B(\asqrt[52] ), .ZN(new_n9644_));
  NAND2_X1   g09452(.A1(new_n9644_), .A2(new_n1103_), .ZN(new_n9645_));
  OAI21_X1   g09453(.A1(new_n9645_), .A2(new_n9631_), .B(new_n9637_), .ZN(new_n9646_));
  AOI21_X1   g09454(.A1(new_n9646_), .A2(new_n9632_), .B(new_n904_), .ZN(new_n9647_));
  OAI21_X1   g09455(.A1(new_n9155_), .A2(new_n9144_), .B(new_n9128_), .ZN(new_n9648_));
  NOR2_X1    g09456(.A1(new_n9648_), .A2(new_n9124_), .ZN(new_n9649_));
  OAI21_X1   g09457(.A1(new_n9144_), .A2(new_n9155_), .B(new_n9145_), .ZN(new_n9650_));
  NOR2_X1    g09458(.A1(new_n9317_), .A2(new_n9650_), .ZN(new_n9651_));
  INV_X1     g09459(.I(new_n9651_), .ZN(new_n9652_));
  AOI22_X1   g09460(.A1(new_n9652_), .A2(new_n9154_), .B1(\asqrt[26] ), .B2(new_n9649_), .ZN(new_n9653_));
  INV_X1     g09461(.I(new_n9627_), .ZN(new_n9654_));
  NAND2_X1   g09462(.A1(new_n9533_), .A2(new_n1256_), .ZN(new_n9655_));
  OAI21_X1   g09463(.A1(new_n9655_), .A2(new_n9643_), .B(new_n9654_), .ZN(new_n9656_));
  AOI21_X1   g09464(.A1(new_n9656_), .A2(new_n9644_), .B(new_n1103_), .ZN(new_n9657_));
  NOR2_X1    g09465(.A1(new_n9657_), .A2(\asqrt[54] ), .ZN(new_n9658_));
  AOI21_X1   g09466(.A1(new_n9658_), .A2(new_n9646_), .B(new_n9653_), .ZN(new_n9659_));
  OAI21_X1   g09467(.A1(new_n9659_), .A2(new_n9647_), .B(\asqrt[55] ), .ZN(new_n9660_));
  NOR2_X1    g09468(.A1(new_n9146_), .A2(new_n9134_), .ZN(new_n9661_));
  NOR3_X1    g09469(.A1(new_n9317_), .A2(new_n9157_), .A3(new_n9661_), .ZN(new_n9662_));
  INV_X1     g09470(.I(new_n9662_), .ZN(new_n9663_));
  NOR3_X1    g09471(.A1(new_n9661_), .A2(new_n9157_), .A3(new_n9142_), .ZN(new_n9664_));
  AOI22_X1   g09472(.A1(new_n9663_), .A2(new_n9142_), .B1(\asqrt[26] ), .B2(new_n9664_), .ZN(new_n9665_));
  INV_X1     g09473(.I(new_n9665_), .ZN(new_n9666_));
  NOR3_X1    g09474(.A1(new_n9532_), .A2(new_n9525_), .A3(\asqrt[51] ), .ZN(new_n9667_));
  OAI21_X1   g09475(.A1(new_n9538_), .A2(new_n9667_), .B(new_n9533_), .ZN(new_n9668_));
  AOI21_X1   g09476(.A1(new_n9668_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n9669_));
  AOI21_X1   g09477(.A1(new_n9669_), .A2(new_n9656_), .B(new_n9636_), .ZN(new_n9670_));
  OAI21_X1   g09478(.A1(new_n9670_), .A2(new_n9657_), .B(\asqrt[54] ), .ZN(new_n9671_));
  NAND2_X1   g09479(.A1(new_n9671_), .A2(new_n823_), .ZN(new_n9672_));
  OAI21_X1   g09480(.A1(new_n9672_), .A2(new_n9659_), .B(new_n9666_), .ZN(new_n9673_));
  AOI21_X1   g09481(.A1(new_n9673_), .A2(new_n9660_), .B(new_n703_), .ZN(new_n9674_));
  NOR3_X1    g09482(.A1(new_n9148_), .A2(new_n9180_), .A3(new_n9191_), .ZN(new_n9675_));
  NOR3_X1    g09483(.A1(new_n9317_), .A2(new_n9148_), .A3(new_n9180_), .ZN(new_n9676_));
  INV_X1     g09484(.I(new_n9676_), .ZN(new_n9677_));
  AOI22_X1   g09485(.A1(new_n9677_), .A2(new_n9191_), .B1(\asqrt[26] ), .B2(new_n9675_), .ZN(new_n9678_));
  NOR3_X1    g09486(.A1(new_n9670_), .A2(\asqrt[54] ), .A3(new_n9657_), .ZN(new_n9679_));
  OAI21_X1   g09487(.A1(new_n9653_), .A2(new_n9679_), .B(new_n9671_), .ZN(new_n9680_));
  AOI21_X1   g09488(.A1(new_n9680_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n9681_));
  AOI21_X1   g09489(.A1(new_n9681_), .A2(new_n9673_), .B(new_n9678_), .ZN(new_n9682_));
  OAI21_X1   g09490(.A1(new_n9682_), .A2(new_n9674_), .B(\asqrt[57] ), .ZN(new_n9683_));
  NOR2_X1    g09491(.A1(new_n9171_), .A2(new_n9159_), .ZN(new_n9684_));
  NOR3_X1    g09492(.A1(new_n9317_), .A2(new_n9194_), .A3(new_n9684_), .ZN(new_n9685_));
  INV_X1     g09493(.I(new_n9685_), .ZN(new_n9686_));
  NOR3_X1    g09494(.A1(new_n9194_), .A2(new_n9684_), .A3(new_n9165_), .ZN(new_n9687_));
  AOI22_X1   g09495(.A1(new_n9686_), .A2(new_n9165_), .B1(\asqrt[26] ), .B2(new_n9687_), .ZN(new_n9688_));
  INV_X1     g09496(.I(new_n9688_), .ZN(new_n9689_));
  INV_X1     g09497(.I(new_n9653_), .ZN(new_n9690_));
  NAND2_X1   g09498(.A1(new_n9632_), .A2(new_n904_), .ZN(new_n9691_));
  OAI21_X1   g09499(.A1(new_n9691_), .A2(new_n9670_), .B(new_n9690_), .ZN(new_n9692_));
  AOI21_X1   g09500(.A1(new_n9692_), .A2(new_n9671_), .B(new_n823_), .ZN(new_n9693_));
  NOR3_X1    g09501(.A1(new_n9631_), .A2(\asqrt[53] ), .A3(new_n9622_), .ZN(new_n9694_));
  OAI21_X1   g09502(.A1(new_n9636_), .A2(new_n9694_), .B(new_n9632_), .ZN(new_n9695_));
  AOI21_X1   g09503(.A1(new_n9695_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n9696_));
  AOI21_X1   g09504(.A1(new_n9696_), .A2(new_n9692_), .B(new_n9665_), .ZN(new_n9697_));
  OAI21_X1   g09505(.A1(new_n9697_), .A2(new_n9693_), .B(\asqrt[56] ), .ZN(new_n9698_));
  NAND2_X1   g09506(.A1(new_n9698_), .A2(new_n531_), .ZN(new_n9699_));
  OAI21_X1   g09507(.A1(new_n9699_), .A2(new_n9682_), .B(new_n9689_), .ZN(new_n9700_));
  AOI21_X1   g09508(.A1(new_n9700_), .A2(new_n9683_), .B(new_n436_), .ZN(new_n9701_));
  NOR2_X1    g09509(.A1(new_n9206_), .A2(new_n9196_), .ZN(new_n9702_));
  NOR3_X1    g09510(.A1(new_n9702_), .A2(new_n9173_), .A3(new_n9205_), .ZN(new_n9703_));
  NOR3_X1    g09511(.A1(new_n9317_), .A2(new_n9173_), .A3(new_n9702_), .ZN(new_n9704_));
  INV_X1     g09512(.I(new_n9704_), .ZN(new_n9705_));
  AOI22_X1   g09513(.A1(new_n9705_), .A2(new_n9205_), .B1(\asqrt[26] ), .B2(new_n9703_), .ZN(new_n9706_));
  NOR3_X1    g09514(.A1(new_n9697_), .A2(\asqrt[56] ), .A3(new_n9693_), .ZN(new_n9707_));
  OAI21_X1   g09515(.A1(new_n9678_), .A2(new_n9707_), .B(new_n9698_), .ZN(new_n9708_));
  AOI21_X1   g09516(.A1(new_n9708_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n9709_));
  AOI21_X1   g09517(.A1(new_n9709_), .A2(new_n9700_), .B(new_n9706_), .ZN(new_n9710_));
  OAI21_X1   g09518(.A1(new_n9710_), .A2(new_n9701_), .B(\asqrt[59] ), .ZN(new_n9711_));
  NOR3_X1    g09519(.A1(new_n9317_), .A2(new_n9208_), .A3(new_n9242_), .ZN(new_n9712_));
  INV_X1     g09520(.I(new_n9712_), .ZN(new_n9713_));
  NOR3_X1    g09521(.A1(new_n9208_), .A2(new_n9242_), .A3(new_n9190_), .ZN(new_n9714_));
  AOI22_X1   g09522(.A1(new_n9713_), .A2(new_n9190_), .B1(\asqrt[26] ), .B2(new_n9714_), .ZN(new_n9715_));
  INV_X1     g09523(.I(new_n9715_), .ZN(new_n9716_));
  INV_X1     g09524(.I(new_n9678_), .ZN(new_n9717_));
  NAND2_X1   g09525(.A1(new_n9660_), .A2(new_n703_), .ZN(new_n9718_));
  OAI21_X1   g09526(.A1(new_n9718_), .A2(new_n9697_), .B(new_n9717_), .ZN(new_n9719_));
  AOI21_X1   g09527(.A1(new_n9719_), .A2(new_n9698_), .B(new_n531_), .ZN(new_n9720_));
  NOR2_X1    g09528(.A1(new_n9674_), .A2(\asqrt[57] ), .ZN(new_n9721_));
  AOI21_X1   g09529(.A1(new_n9721_), .A2(new_n9719_), .B(new_n9688_), .ZN(new_n9722_));
  OAI21_X1   g09530(.A1(new_n9722_), .A2(new_n9720_), .B(\asqrt[58] ), .ZN(new_n9723_));
  NAND2_X1   g09531(.A1(new_n9723_), .A2(new_n327_), .ZN(new_n9724_));
  OAI21_X1   g09532(.A1(new_n9724_), .A2(new_n9710_), .B(new_n9716_), .ZN(new_n9725_));
  AOI21_X1   g09533(.A1(new_n9725_), .A2(new_n9711_), .B(new_n306_), .ZN(new_n9726_));
  NOR2_X1    g09534(.A1(new_n9231_), .A2(new_n9220_), .ZN(new_n9727_));
  NOR3_X1    g09535(.A1(new_n9200_), .A2(new_n9727_), .A3(new_n9230_), .ZN(new_n9728_));
  NOR3_X1    g09536(.A1(new_n9317_), .A2(new_n9200_), .A3(new_n9727_), .ZN(new_n9729_));
  INV_X1     g09537(.I(new_n9729_), .ZN(new_n9730_));
  AOI22_X1   g09538(.A1(new_n9730_), .A2(new_n9230_), .B1(\asqrt[26] ), .B2(new_n9728_), .ZN(new_n9731_));
  INV_X1     g09539(.I(new_n9706_), .ZN(new_n9732_));
  NAND2_X1   g09540(.A1(new_n9683_), .A2(new_n436_), .ZN(new_n9733_));
  OAI21_X1   g09541(.A1(new_n9733_), .A2(new_n9722_), .B(new_n9732_), .ZN(new_n9734_));
  AOI21_X1   g09542(.A1(new_n9734_), .A2(new_n9723_), .B(new_n327_), .ZN(new_n9735_));
  NOR2_X1    g09543(.A1(new_n9735_), .A2(\asqrt[60] ), .ZN(new_n9736_));
  AOI21_X1   g09544(.A1(new_n9736_), .A2(new_n9725_), .B(new_n9731_), .ZN(new_n9737_));
  OAI21_X1   g09545(.A1(new_n9737_), .A2(new_n9726_), .B(\asqrt[61] ), .ZN(new_n9738_));
  NOR2_X1    g09546(.A1(new_n9222_), .A2(new_n9210_), .ZN(new_n9739_));
  NOR3_X1    g09547(.A1(new_n9317_), .A2(new_n9233_), .A3(new_n9739_), .ZN(new_n9740_));
  INV_X1     g09548(.I(new_n9740_), .ZN(new_n9741_));
  NOR3_X1    g09549(.A1(new_n9739_), .A2(new_n9233_), .A3(new_n9218_), .ZN(new_n9742_));
  AOI22_X1   g09550(.A1(new_n9741_), .A2(new_n9218_), .B1(\asqrt[26] ), .B2(new_n9742_), .ZN(new_n9743_));
  INV_X1     g09551(.I(new_n9743_), .ZN(new_n9744_));
  NOR3_X1    g09552(.A1(new_n9682_), .A2(\asqrt[57] ), .A3(new_n9674_), .ZN(new_n9745_));
  OAI21_X1   g09553(.A1(new_n9688_), .A2(new_n9745_), .B(new_n9683_), .ZN(new_n9746_));
  AOI21_X1   g09554(.A1(new_n9746_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n9747_));
  AOI21_X1   g09555(.A1(new_n9747_), .A2(new_n9734_), .B(new_n9715_), .ZN(new_n9748_));
  OAI21_X1   g09556(.A1(new_n9748_), .A2(new_n9735_), .B(\asqrt[60] ), .ZN(new_n9749_));
  NAND2_X1   g09557(.A1(new_n9749_), .A2(new_n218_), .ZN(new_n9750_));
  OAI21_X1   g09558(.A1(new_n9750_), .A2(new_n9737_), .B(new_n9744_), .ZN(new_n9751_));
  AOI21_X1   g09559(.A1(new_n9751_), .A2(new_n9738_), .B(new_n207_), .ZN(new_n9752_));
  NOR3_X1    g09560(.A1(new_n9224_), .A2(new_n9258_), .A3(new_n9286_), .ZN(new_n9753_));
  NOR3_X1    g09561(.A1(new_n9317_), .A2(new_n9224_), .A3(new_n9258_), .ZN(new_n9754_));
  INV_X1     g09562(.I(new_n9754_), .ZN(new_n9755_));
  AOI22_X1   g09563(.A1(new_n9755_), .A2(new_n9286_), .B1(\asqrt[26] ), .B2(new_n9753_), .ZN(new_n9756_));
  NOR3_X1    g09564(.A1(new_n9748_), .A2(\asqrt[60] ), .A3(new_n9735_), .ZN(new_n9757_));
  OAI21_X1   g09565(.A1(new_n9731_), .A2(new_n9757_), .B(new_n9749_), .ZN(new_n9758_));
  AOI21_X1   g09566(.A1(new_n9758_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n9759_));
  AOI21_X1   g09567(.A1(new_n9759_), .A2(new_n9751_), .B(new_n9756_), .ZN(new_n9760_));
  AND3_X2    g09568(.A1(new_n9236_), .A2(new_n9289_), .A3(new_n9240_), .Z(new_n9761_));
  NAND2_X1   g09569(.A1(\asqrt[26] ), .A2(new_n9761_), .ZN(new_n9762_));
  INV_X1     g09570(.I(new_n9762_), .ZN(new_n9763_));
  AND2_X2    g09571(.A1(new_n9236_), .A2(new_n9289_), .Z(new_n9764_));
  AOI21_X1   g09572(.A1(\asqrt[26] ), .A2(new_n9764_), .B(new_n9240_), .ZN(new_n9765_));
  NOR2_X1    g09573(.A1(new_n9763_), .A2(new_n9765_), .ZN(new_n9766_));
  NOR3_X1    g09574(.A1(new_n9317_), .A2(new_n9290_), .A3(new_n9280_), .ZN(new_n9767_));
  NOR3_X1    g09575(.A1(new_n9766_), .A2(new_n9303_), .A3(new_n9767_), .ZN(new_n9768_));
  OAI21_X1   g09576(.A1(new_n9760_), .A2(new_n9752_), .B(new_n9768_), .ZN(new_n9769_));
  NAND2_X1   g09577(.A1(new_n9769_), .A2(new_n193_), .ZN(new_n9770_));
  INV_X1     g09578(.I(new_n9756_), .ZN(new_n9771_));
  NAND3_X1   g09579(.A1(new_n9751_), .A2(new_n207_), .A3(new_n9738_), .ZN(new_n9772_));
  NAND2_X1   g09580(.A1(new_n9772_), .A2(new_n9771_), .ZN(new_n9773_));
  INV_X1     g09581(.I(new_n9766_), .ZN(new_n9774_));
  NOR2_X1    g09582(.A1(new_n9752_), .A2(new_n9774_), .ZN(new_n9775_));
  AOI21_X1   g09583(.A1(\asqrt[26] ), .A2(new_n9253_), .B(new_n9276_), .ZN(new_n9776_));
  OAI21_X1   g09584(.A1(new_n9290_), .A2(new_n9280_), .B(\asqrt[63] ), .ZN(new_n9777_));
  NOR2_X1    g09585(.A1(new_n9776_), .A2(new_n9777_), .ZN(new_n9778_));
  INV_X1     g09586(.I(new_n9303_), .ZN(new_n9779_));
  AND3_X2    g09587(.A1(new_n9252_), .A2(new_n9250_), .A3(new_n9266_), .Z(new_n9780_));
  NAND4_X1   g09588(.A1(new_n9779_), .A2(new_n9291_), .A3(new_n9263_), .A4(new_n9780_), .ZN(new_n9781_));
  INV_X1     g09589(.I(new_n9781_), .ZN(new_n9782_));
  NOR2_X1    g09590(.A1(new_n9778_), .A2(new_n9782_), .ZN(new_n9783_));
  INV_X1     g09591(.I(new_n9783_), .ZN(new_n9784_));
  AOI21_X1   g09592(.A1(new_n9775_), .A2(new_n9773_), .B(new_n9784_), .ZN(new_n9785_));
  NAND2_X1   g09593(.A1(new_n9770_), .A2(new_n9785_), .ZN(\asqrt[25] ));
  NOR2_X1    g09594(.A1(\a[48] ), .A2(\a[49] ), .ZN(new_n9787_));
  INV_X1     g09595(.I(new_n9787_), .ZN(new_n9788_));
  NOR2_X1    g09596(.A1(new_n9788_), .A2(\a[50] ), .ZN(new_n9789_));
  INV_X1     g09597(.I(new_n9789_), .ZN(new_n9790_));
  INV_X1     g09598(.I(new_n9731_), .ZN(new_n9791_));
  NAND2_X1   g09599(.A1(new_n9711_), .A2(new_n306_), .ZN(new_n9792_));
  OAI21_X1   g09600(.A1(new_n9792_), .A2(new_n9748_), .B(new_n9791_), .ZN(new_n9793_));
  AOI21_X1   g09601(.A1(new_n9793_), .A2(new_n9749_), .B(new_n218_), .ZN(new_n9794_));
  NOR3_X1    g09602(.A1(new_n9710_), .A2(\asqrt[59] ), .A3(new_n9701_), .ZN(new_n9795_));
  OAI21_X1   g09603(.A1(new_n9715_), .A2(new_n9795_), .B(new_n9711_), .ZN(new_n9796_));
  AOI21_X1   g09604(.A1(new_n9796_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n9797_));
  AOI21_X1   g09605(.A1(new_n9797_), .A2(new_n9793_), .B(new_n9743_), .ZN(new_n9798_));
  OAI21_X1   g09606(.A1(new_n9798_), .A2(new_n9794_), .B(\asqrt[62] ), .ZN(new_n9799_));
  NOR3_X1    g09607(.A1(new_n9798_), .A2(\asqrt[62] ), .A3(new_n9794_), .ZN(new_n9800_));
  OAI21_X1   g09608(.A1(new_n9756_), .A2(new_n9800_), .B(new_n9799_), .ZN(new_n9801_));
  AOI21_X1   g09609(.A1(new_n9801_), .A2(new_n9768_), .B(\asqrt[63] ), .ZN(new_n9802_));
  NAND2_X1   g09610(.A1(new_n9799_), .A2(new_n9766_), .ZN(new_n9803_));
  OAI21_X1   g09611(.A1(new_n9803_), .A2(new_n9760_), .B(new_n9783_), .ZN(new_n9804_));
  OAI21_X1   g09612(.A1(new_n9802_), .A2(new_n9804_), .B(\a[50] ), .ZN(new_n9805_));
  AOI21_X1   g09613(.A1(new_n9805_), .A2(new_n9790_), .B(new_n9317_), .ZN(new_n9806_));
  INV_X1     g09614(.I(\a[50] ), .ZN(new_n9807_));
  AOI21_X1   g09615(.A1(new_n9770_), .A2(new_n9785_), .B(new_n9807_), .ZN(new_n9808_));
  NAND2_X1   g09616(.A1(new_n9266_), .A2(new_n9790_), .ZN(new_n9809_));
  NOR4_X1    g09617(.A1(new_n9278_), .A2(new_n9303_), .A3(new_n9264_), .A4(new_n9809_), .ZN(new_n9810_));
  INV_X1     g09618(.I(new_n9810_), .ZN(new_n9811_));
  NOR2_X1    g09619(.A1(new_n9808_), .A2(new_n9811_), .ZN(new_n9812_));
  AOI21_X1   g09620(.A1(new_n9770_), .A2(new_n9785_), .B(new_n9273_), .ZN(new_n9813_));
  INV_X1     g09621(.I(\a[51] ), .ZN(new_n9814_));
  AOI21_X1   g09622(.A1(\asqrt[25] ), .A2(new_n9807_), .B(new_n9814_), .ZN(new_n9815_));
  NOR3_X1    g09623(.A1(new_n9812_), .A2(new_n9815_), .A3(new_n9813_), .ZN(new_n9816_));
  OAI21_X1   g09624(.A1(new_n9816_), .A2(new_n9806_), .B(\asqrt[27] ), .ZN(new_n9817_));
  OAI21_X1   g09625(.A1(new_n9802_), .A2(new_n9804_), .B(new_n9272_), .ZN(new_n9818_));
  NAND2_X1   g09626(.A1(new_n9775_), .A2(new_n9773_), .ZN(new_n9819_));
  INV_X1     g09627(.I(new_n9778_), .ZN(new_n9820_));
  NOR2_X1    g09628(.A1(new_n9782_), .A2(new_n9317_), .ZN(new_n9821_));
  NAND4_X1   g09629(.A1(new_n9770_), .A2(new_n9819_), .A3(new_n9820_), .A4(new_n9821_), .ZN(new_n9822_));
  AOI21_X1   g09630(.A1(new_n9822_), .A2(new_n9818_), .B(new_n9285_), .ZN(new_n9823_));
  INV_X1     g09631(.I(new_n9819_), .ZN(new_n9824_));
  NAND2_X1   g09632(.A1(new_n9820_), .A2(new_n9821_), .ZN(new_n9825_));
  NOR3_X1    g09633(.A1(new_n9824_), .A2(new_n9802_), .A3(new_n9825_), .ZN(new_n9826_));
  NOR3_X1    g09634(.A1(new_n9826_), .A2(new_n9813_), .A3(\a[52] ), .ZN(new_n9827_));
  OAI21_X1   g09635(.A1(new_n9808_), .A2(new_n9789_), .B(\asqrt[26] ), .ZN(new_n9828_));
  NAND2_X1   g09636(.A1(new_n9828_), .A2(new_n8826_), .ZN(new_n9829_));
  OAI22_X1   g09637(.A1(new_n9816_), .A2(new_n9829_), .B1(new_n9823_), .B2(new_n9827_), .ZN(new_n9830_));
  AOI21_X1   g09638(.A1(new_n9830_), .A2(new_n9817_), .B(new_n8483_), .ZN(new_n9831_));
  NOR3_X1    g09639(.A1(new_n9563_), .A2(new_n9284_), .A3(new_n9296_), .ZN(new_n9832_));
  NAND3_X1   g09640(.A1(\asqrt[25] ), .A2(new_n9320_), .A3(new_n9546_), .ZN(new_n9833_));
  AOI22_X1   g09641(.A1(new_n9833_), .A2(new_n9563_), .B1(\asqrt[25] ), .B2(new_n9832_), .ZN(new_n9834_));
  AOI21_X1   g09642(.A1(new_n9770_), .A2(new_n9785_), .B(\a[50] ), .ZN(new_n9835_));
  OAI21_X1   g09643(.A1(new_n9814_), .A2(new_n9835_), .B(new_n9818_), .ZN(new_n9836_));
  OAI21_X1   g09644(.A1(new_n9836_), .A2(new_n9812_), .B(new_n9828_), .ZN(new_n9837_));
  AOI21_X1   g09645(.A1(new_n9837_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n9838_));
  AOI21_X1   g09646(.A1(new_n9838_), .A2(new_n9830_), .B(new_n9834_), .ZN(new_n9839_));
  OAI21_X1   g09647(.A1(new_n9839_), .A2(new_n9831_), .B(\asqrt[29] ), .ZN(new_n9840_));
  INV_X1     g09648(.I(new_n9840_), .ZN(new_n9841_));
  NOR2_X1    g09649(.A1(new_n9308_), .A2(new_n9309_), .ZN(new_n9842_));
  NOR2_X1    g09650(.A1(new_n9300_), .A2(new_n9311_), .ZN(new_n9843_));
  INV_X1     g09651(.I(new_n9843_), .ZN(new_n9844_));
  NAND4_X1   g09652(.A1(\asqrt[25] ), .A2(new_n9301_), .A3(new_n9842_), .A4(new_n9844_), .ZN(new_n9845_));
  INV_X1     g09653(.I(\asqrt[25] ), .ZN(new_n9846_));
  NOR3_X1    g09654(.A1(new_n9846_), .A2(new_n9550_), .A3(new_n9843_), .ZN(new_n9847_));
  OAI21_X1   g09655(.A1(new_n9847_), .A2(new_n9842_), .B(new_n9845_), .ZN(new_n9848_));
  INV_X1     g09656(.I(new_n9848_), .ZN(new_n9849_));
  NOR3_X1    g09657(.A1(new_n9839_), .A2(new_n9831_), .A3(\asqrt[29] ), .ZN(new_n9850_));
  NOR2_X1    g09658(.A1(new_n9850_), .A2(new_n9849_), .ZN(new_n9851_));
  OAI21_X1   g09659(.A1(new_n9851_), .A2(new_n9841_), .B(\asqrt[30] ), .ZN(new_n9852_));
  NOR2_X1    g09660(.A1(new_n9565_), .A2(new_n9555_), .ZN(new_n9853_));
  NOR3_X1    g09661(.A1(new_n9846_), .A2(new_n9313_), .A3(new_n9853_), .ZN(new_n9854_));
  INV_X1     g09662(.I(new_n9854_), .ZN(new_n9855_));
  NOR3_X1    g09663(.A1(new_n9853_), .A2(new_n9313_), .A3(new_n9562_), .ZN(new_n9856_));
  AOI22_X1   g09664(.A1(new_n9855_), .A2(new_n9562_), .B1(\asqrt[25] ), .B2(new_n9856_), .ZN(new_n9857_));
  INV_X1     g09665(.I(new_n9857_), .ZN(new_n9858_));
  NAND2_X1   g09666(.A1(new_n9840_), .A2(new_n7539_), .ZN(new_n9859_));
  OAI21_X1   g09667(.A1(new_n9851_), .A2(new_n9859_), .B(new_n9858_), .ZN(new_n9860_));
  AOI21_X1   g09668(.A1(new_n9860_), .A2(new_n9852_), .B(new_n7229_), .ZN(new_n9861_));
  NOR3_X1    g09669(.A1(new_n9327_), .A2(new_n9336_), .A3(new_n9334_), .ZN(new_n9862_));
  NOR3_X1    g09670(.A1(new_n9846_), .A2(new_n9327_), .A3(new_n9336_), .ZN(new_n9863_));
  INV_X1     g09671(.I(new_n9863_), .ZN(new_n9864_));
  AOI22_X1   g09672(.A1(new_n9864_), .A2(new_n9334_), .B1(\asqrt[25] ), .B2(new_n9862_), .ZN(new_n9865_));
  OAI21_X1   g09673(.A1(new_n9849_), .A2(new_n9850_), .B(new_n9840_), .ZN(new_n9866_));
  AOI21_X1   g09674(.A1(new_n9866_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n9867_));
  AOI21_X1   g09675(.A1(new_n9867_), .A2(new_n9860_), .B(new_n9865_), .ZN(new_n9868_));
  OAI21_X1   g09676(.A1(new_n9868_), .A2(new_n9861_), .B(\asqrt[32] ), .ZN(new_n9869_));
  NAND2_X1   g09677(.A1(new_n9568_), .A2(new_n9558_), .ZN(new_n9870_));
  NAND3_X1   g09678(.A1(\asqrt[25] ), .A2(new_n9338_), .A3(new_n9870_), .ZN(new_n9871_));
  AND3_X2    g09679(.A1(new_n9338_), .A2(new_n9344_), .A3(new_n9870_), .Z(new_n9872_));
  AOI22_X1   g09680(.A1(new_n9871_), .A2(new_n9345_), .B1(\asqrt[25] ), .B2(new_n9872_), .ZN(new_n9873_));
  INV_X1     g09681(.I(new_n9873_), .ZN(new_n9874_));
  NAND2_X1   g09682(.A1(new_n9805_), .A2(new_n9810_), .ZN(new_n9875_));
  OAI21_X1   g09683(.A1(new_n9802_), .A2(new_n9804_), .B(new_n9807_), .ZN(new_n9876_));
  NAND2_X1   g09684(.A1(new_n9876_), .A2(\a[51] ), .ZN(new_n9877_));
  NAND3_X1   g09685(.A1(new_n9875_), .A2(new_n9877_), .A3(new_n9818_), .ZN(new_n9878_));
  AOI21_X1   g09686(.A1(new_n9878_), .A2(new_n9828_), .B(new_n8826_), .ZN(new_n9879_));
  OAI21_X1   g09687(.A1(new_n9826_), .A2(new_n9813_), .B(\a[52] ), .ZN(new_n9880_));
  NAND3_X1   g09688(.A1(new_n9822_), .A2(new_n9818_), .A3(new_n9285_), .ZN(new_n9881_));
  NAND2_X1   g09689(.A1(new_n9805_), .A2(new_n9790_), .ZN(new_n9882_));
  AOI21_X1   g09690(.A1(new_n9882_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n9883_));
  AOI22_X1   g09691(.A1(new_n9878_), .A2(new_n9883_), .B1(new_n9880_), .B2(new_n9881_), .ZN(new_n9884_));
  OAI21_X1   g09692(.A1(new_n9884_), .A2(new_n9879_), .B(\asqrt[28] ), .ZN(new_n9885_));
  NAND2_X1   g09693(.A1(new_n9885_), .A2(new_n8036_), .ZN(new_n9886_));
  OAI21_X1   g09694(.A1(new_n9886_), .A2(new_n9839_), .B(new_n9848_), .ZN(new_n9887_));
  AOI21_X1   g09695(.A1(new_n9887_), .A2(new_n9840_), .B(new_n7539_), .ZN(new_n9888_));
  INV_X1     g09696(.I(new_n9834_), .ZN(new_n9889_));
  AOI21_X1   g09697(.A1(\a[51] ), .A2(new_n9876_), .B(new_n9813_), .ZN(new_n9890_));
  AOI21_X1   g09698(.A1(new_n9890_), .A2(new_n9875_), .B(new_n9806_), .ZN(new_n9891_));
  OAI21_X1   g09699(.A1(new_n9891_), .A2(new_n8826_), .B(new_n8483_), .ZN(new_n9892_));
  OAI21_X1   g09700(.A1(new_n9892_), .A2(new_n9884_), .B(new_n9889_), .ZN(new_n9893_));
  NAND2_X1   g09701(.A1(new_n9893_), .A2(new_n9885_), .ZN(new_n9894_));
  AOI21_X1   g09702(.A1(new_n9894_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n9895_));
  AOI21_X1   g09703(.A1(new_n9895_), .A2(new_n9887_), .B(new_n9857_), .ZN(new_n9896_));
  OAI21_X1   g09704(.A1(new_n9896_), .A2(new_n9888_), .B(\asqrt[31] ), .ZN(new_n9897_));
  NAND2_X1   g09705(.A1(new_n9897_), .A2(new_n6824_), .ZN(new_n9898_));
  OAI21_X1   g09706(.A1(new_n9898_), .A2(new_n9868_), .B(new_n9874_), .ZN(new_n9899_));
  AOI21_X1   g09707(.A1(new_n9899_), .A2(new_n9869_), .B(new_n6356_), .ZN(new_n9900_));
  INV_X1     g09708(.I(new_n9900_), .ZN(new_n9901_));
  INV_X1     g09709(.I(new_n9899_), .ZN(new_n9902_));
  INV_X1     g09710(.I(new_n9353_), .ZN(new_n9903_));
  NOR3_X1    g09711(.A1(new_n9348_), .A2(new_n9579_), .A3(new_n9903_), .ZN(new_n9904_));
  NOR3_X1    g09712(.A1(new_n9846_), .A2(new_n9348_), .A3(new_n9579_), .ZN(new_n9905_));
  INV_X1     g09713(.I(new_n9905_), .ZN(new_n9906_));
  AOI22_X1   g09714(.A1(new_n9906_), .A2(new_n9903_), .B1(\asqrt[25] ), .B2(new_n9904_), .ZN(new_n9907_));
  INV_X1     g09715(.I(new_n9907_), .ZN(new_n9908_));
  NAND2_X1   g09716(.A1(new_n9869_), .A2(new_n6356_), .ZN(new_n9909_));
  OAI21_X1   g09717(.A1(new_n9902_), .A2(new_n9909_), .B(new_n9908_), .ZN(new_n9910_));
  AOI21_X1   g09718(.A1(new_n9901_), .A2(new_n9910_), .B(new_n6077_), .ZN(new_n9911_));
  NOR3_X1    g09719(.A1(new_n9846_), .A2(new_n9358_), .A3(new_n9365_), .ZN(new_n9912_));
  INV_X1     g09720(.I(new_n9912_), .ZN(new_n9913_));
  NOR3_X1    g09721(.A1(new_n9358_), .A2(new_n9545_), .A3(new_n9365_), .ZN(new_n9914_));
  AOI22_X1   g09722(.A1(new_n9913_), .A2(new_n9545_), .B1(\asqrt[25] ), .B2(new_n9914_), .ZN(new_n9915_));
  NOR2_X1    g09723(.A1(new_n9900_), .A2(\asqrt[34] ), .ZN(new_n9916_));
  AOI21_X1   g09724(.A1(new_n9916_), .A2(new_n9910_), .B(new_n9915_), .ZN(new_n9917_));
  OAI21_X1   g09725(.A1(new_n9917_), .A2(new_n9911_), .B(\asqrt[35] ), .ZN(new_n9918_));
  INV_X1     g09726(.I(new_n9918_), .ZN(new_n9919_));
  INV_X1     g09727(.I(new_n9573_), .ZN(new_n9920_));
  NOR3_X1    g09728(.A1(new_n9920_), .A2(new_n9578_), .A3(new_n9377_), .ZN(new_n9921_));
  NOR3_X1    g09729(.A1(new_n9846_), .A2(new_n9578_), .A3(new_n9920_), .ZN(new_n9922_));
  INV_X1     g09730(.I(new_n9922_), .ZN(new_n9923_));
  AOI22_X1   g09731(.A1(new_n9923_), .A2(new_n9377_), .B1(\asqrt[25] ), .B2(new_n9921_), .ZN(new_n9924_));
  NOR3_X1    g09732(.A1(new_n9917_), .A2(new_n9911_), .A3(\asqrt[35] ), .ZN(new_n9925_));
  NOR2_X1    g09733(.A1(new_n9925_), .A2(new_n9924_), .ZN(new_n9926_));
  OAI21_X1   g09734(.A1(new_n9926_), .A2(new_n9919_), .B(\asqrt[36] ), .ZN(new_n9927_));
  INV_X1     g09735(.I(new_n9385_), .ZN(new_n9928_));
  NOR3_X1    g09736(.A1(new_n9846_), .A2(new_n9380_), .A3(new_n9583_), .ZN(new_n9929_));
  INV_X1     g09737(.I(new_n9929_), .ZN(new_n9930_));
  NOR3_X1    g09738(.A1(new_n9380_), .A2(new_n9583_), .A3(new_n9928_), .ZN(new_n9931_));
  AOI22_X1   g09739(.A1(new_n9930_), .A2(new_n9928_), .B1(\asqrt[25] ), .B2(new_n9931_), .ZN(new_n9932_));
  INV_X1     g09740(.I(new_n9932_), .ZN(new_n9933_));
  NAND2_X1   g09741(.A1(new_n9918_), .A2(new_n5277_), .ZN(new_n9934_));
  OAI21_X1   g09742(.A1(new_n9926_), .A2(new_n9934_), .B(new_n9933_), .ZN(new_n9935_));
  AOI21_X1   g09743(.A1(new_n9935_), .A2(new_n9927_), .B(new_n5024_), .ZN(new_n9936_));
  NOR3_X1    g09744(.A1(new_n9390_), .A2(new_n9544_), .A3(new_n9396_), .ZN(new_n9937_));
  NOR3_X1    g09745(.A1(new_n9846_), .A2(new_n9390_), .A3(new_n9396_), .ZN(new_n9938_));
  INV_X1     g09746(.I(new_n9938_), .ZN(new_n9939_));
  AOI22_X1   g09747(.A1(new_n9939_), .A2(new_n9544_), .B1(\asqrt[25] ), .B2(new_n9937_), .ZN(new_n9940_));
  INV_X1     g09748(.I(new_n9924_), .ZN(new_n9941_));
  NOR3_X1    g09749(.A1(new_n9868_), .A2(new_n9861_), .A3(\asqrt[32] ), .ZN(new_n9942_));
  OAI21_X1   g09750(.A1(new_n9873_), .A2(new_n9942_), .B(new_n9869_), .ZN(new_n9943_));
  NAND3_X1   g09751(.A1(new_n9899_), .A2(new_n6356_), .A3(new_n9869_), .ZN(new_n9944_));
  AOI22_X1   g09752(.A1(new_n9944_), .A2(new_n9908_), .B1(new_n9943_), .B2(\asqrt[33] ), .ZN(new_n9945_));
  OAI21_X1   g09753(.A1(new_n9945_), .A2(new_n6077_), .B(new_n5708_), .ZN(new_n9946_));
  OAI21_X1   g09754(.A1(new_n9946_), .A2(new_n9917_), .B(new_n9941_), .ZN(new_n9947_));
  AOI21_X1   g09755(.A1(new_n9947_), .A2(new_n9918_), .B(new_n5277_), .ZN(new_n9948_));
  NOR2_X1    g09756(.A1(new_n9948_), .A2(\asqrt[37] ), .ZN(new_n9949_));
  AOI21_X1   g09757(.A1(new_n9949_), .A2(new_n9935_), .B(new_n9940_), .ZN(new_n9950_));
  OAI21_X1   g09758(.A1(new_n9950_), .A2(new_n9936_), .B(\asqrt[38] ), .ZN(new_n9951_));
  INV_X1     g09759(.I(new_n9951_), .ZN(new_n9952_));
  NOR2_X1    g09760(.A1(new_n9397_), .A2(new_n9408_), .ZN(new_n9953_));
  NOR3_X1    g09761(.A1(new_n9846_), .A2(new_n9577_), .A3(new_n9953_), .ZN(new_n9954_));
  INV_X1     g09762(.I(new_n9954_), .ZN(new_n9955_));
  NOR3_X1    g09763(.A1(new_n9953_), .A2(new_n9577_), .A3(new_n9407_), .ZN(new_n9956_));
  AOI22_X1   g09764(.A1(new_n9955_), .A2(new_n9407_), .B1(\asqrt[25] ), .B2(new_n9956_), .ZN(new_n9957_));
  NOR3_X1    g09765(.A1(new_n9950_), .A2(new_n9936_), .A3(\asqrt[38] ), .ZN(new_n9958_));
  NOR2_X1    g09766(.A1(new_n9958_), .A2(new_n9957_), .ZN(new_n9959_));
  OAI21_X1   g09767(.A1(new_n9959_), .A2(new_n9952_), .B(\asqrt[39] ), .ZN(new_n9960_));
  INV_X1     g09768(.I(new_n9415_), .ZN(new_n9961_));
  NOR3_X1    g09769(.A1(new_n9410_), .A2(new_n9591_), .A3(new_n9961_), .ZN(new_n9962_));
  NOR3_X1    g09770(.A1(new_n9846_), .A2(new_n9410_), .A3(new_n9591_), .ZN(new_n9963_));
  INV_X1     g09771(.I(new_n9963_), .ZN(new_n9964_));
  AOI22_X1   g09772(.A1(new_n9964_), .A2(new_n9961_), .B1(\asqrt[25] ), .B2(new_n9962_), .ZN(new_n9965_));
  INV_X1     g09773(.I(new_n9965_), .ZN(new_n9966_));
  NAND2_X1   g09774(.A1(new_n9951_), .A2(new_n4298_), .ZN(new_n9967_));
  OAI21_X1   g09775(.A1(new_n9959_), .A2(new_n9967_), .B(new_n9966_), .ZN(new_n9968_));
  AOI21_X1   g09776(.A1(new_n9968_), .A2(new_n9960_), .B(new_n4071_), .ZN(new_n9969_));
  NOR3_X1    g09777(.A1(new_n9846_), .A2(new_n9420_), .A3(new_n9427_), .ZN(new_n9970_));
  INV_X1     g09778(.I(new_n9970_), .ZN(new_n9971_));
  NOR3_X1    g09779(.A1(new_n9420_), .A2(new_n9543_), .A3(new_n9427_), .ZN(new_n9972_));
  AOI22_X1   g09780(.A1(new_n9971_), .A2(new_n9543_), .B1(\asqrt[25] ), .B2(new_n9972_), .ZN(new_n9973_));
  INV_X1     g09781(.I(new_n9957_), .ZN(new_n9974_));
  NOR3_X1    g09782(.A1(new_n9896_), .A2(new_n9888_), .A3(\asqrt[31] ), .ZN(new_n9975_));
  OAI21_X1   g09783(.A1(new_n9865_), .A2(new_n9975_), .B(new_n9897_), .ZN(new_n9976_));
  AOI21_X1   g09784(.A1(new_n9976_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n9977_));
  AOI21_X1   g09785(.A1(new_n9977_), .A2(new_n9899_), .B(new_n9907_), .ZN(new_n9978_));
  NOR3_X1    g09786(.A1(new_n9978_), .A2(\asqrt[34] ), .A3(new_n9900_), .ZN(new_n9979_));
  OAI22_X1   g09787(.A1(new_n9979_), .A2(new_n9915_), .B1(new_n9945_), .B2(new_n6077_), .ZN(new_n9980_));
  AOI21_X1   g09788(.A1(new_n9980_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n9981_));
  AOI21_X1   g09789(.A1(new_n9981_), .A2(new_n9947_), .B(new_n9932_), .ZN(new_n9982_));
  OAI21_X1   g09790(.A1(new_n9982_), .A2(new_n9948_), .B(\asqrt[37] ), .ZN(new_n9983_));
  NAND2_X1   g09791(.A1(new_n9983_), .A2(new_n4696_), .ZN(new_n9984_));
  OAI21_X1   g09792(.A1(new_n9984_), .A2(new_n9950_), .B(new_n9974_), .ZN(new_n9985_));
  AOI21_X1   g09793(.A1(new_n9985_), .A2(new_n9951_), .B(new_n4298_), .ZN(new_n9986_));
  NOR2_X1    g09794(.A1(new_n9986_), .A2(\asqrt[40] ), .ZN(new_n9987_));
  AOI21_X1   g09795(.A1(new_n9987_), .A2(new_n9968_), .B(new_n9973_), .ZN(new_n9988_));
  OAI21_X1   g09796(.A1(new_n9988_), .A2(new_n9969_), .B(\asqrt[41] ), .ZN(new_n9989_));
  NOR2_X1    g09797(.A1(new_n9428_), .A2(new_n9439_), .ZN(new_n9990_));
  NOR3_X1    g09798(.A1(new_n9990_), .A2(new_n9590_), .A3(new_n9438_), .ZN(new_n9991_));
  NOR3_X1    g09799(.A1(new_n9846_), .A2(new_n9590_), .A3(new_n9990_), .ZN(new_n9992_));
  INV_X1     g09800(.I(new_n9992_), .ZN(new_n9993_));
  AOI22_X1   g09801(.A1(new_n9993_), .A2(new_n9438_), .B1(\asqrt[25] ), .B2(new_n9991_), .ZN(new_n9994_));
  INV_X1     g09802(.I(new_n9994_), .ZN(new_n9995_));
  NOR3_X1    g09803(.A1(new_n9982_), .A2(\asqrt[37] ), .A3(new_n9948_), .ZN(new_n9996_));
  OAI21_X1   g09804(.A1(new_n9940_), .A2(new_n9996_), .B(new_n9983_), .ZN(new_n9997_));
  AOI21_X1   g09805(.A1(new_n9997_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n9998_));
  AOI21_X1   g09806(.A1(new_n9998_), .A2(new_n9985_), .B(new_n9965_), .ZN(new_n9999_));
  OAI21_X1   g09807(.A1(new_n9999_), .A2(new_n9986_), .B(\asqrt[40] ), .ZN(new_n10000_));
  NAND2_X1   g09808(.A1(new_n10000_), .A2(new_n3782_), .ZN(new_n10001_));
  OAI21_X1   g09809(.A1(new_n10001_), .A2(new_n9988_), .B(new_n9995_), .ZN(new_n10002_));
  AOI21_X1   g09810(.A1(new_n10002_), .A2(new_n9989_), .B(new_n3419_), .ZN(new_n10003_));
  INV_X1     g09811(.I(new_n9446_), .ZN(new_n10004_));
  NOR3_X1    g09812(.A1(new_n9846_), .A2(new_n9441_), .A3(new_n9599_), .ZN(new_n10005_));
  INV_X1     g09813(.I(new_n10005_), .ZN(new_n10006_));
  NOR3_X1    g09814(.A1(new_n9441_), .A2(new_n9599_), .A3(new_n10004_), .ZN(new_n10007_));
  AOI22_X1   g09815(.A1(new_n10006_), .A2(new_n10004_), .B1(\asqrt[25] ), .B2(new_n10007_), .ZN(new_n10008_));
  NOR3_X1    g09816(.A1(new_n9999_), .A2(\asqrt[40] ), .A3(new_n9986_), .ZN(new_n10009_));
  OAI21_X1   g09817(.A1(new_n9973_), .A2(new_n10009_), .B(new_n10000_), .ZN(new_n10010_));
  AOI21_X1   g09818(.A1(new_n10010_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n10011_));
  AOI21_X1   g09819(.A1(new_n10011_), .A2(new_n10002_), .B(new_n10008_), .ZN(new_n10012_));
  OAI21_X1   g09820(.A1(new_n10012_), .A2(new_n10003_), .B(\asqrt[43] ), .ZN(new_n10013_));
  INV_X1     g09821(.I(new_n10013_), .ZN(new_n10014_));
  NOR3_X1    g09822(.A1(new_n9451_), .A2(new_n9542_), .A3(new_n9457_), .ZN(new_n10015_));
  NOR3_X1    g09823(.A1(new_n9846_), .A2(new_n9451_), .A3(new_n9457_), .ZN(new_n10016_));
  INV_X1     g09824(.I(new_n10016_), .ZN(new_n10017_));
  AOI22_X1   g09825(.A1(new_n10017_), .A2(new_n9542_), .B1(\asqrt[25] ), .B2(new_n10015_), .ZN(new_n10018_));
  NOR3_X1    g09826(.A1(new_n10012_), .A2(\asqrt[43] ), .A3(new_n10003_), .ZN(new_n10019_));
  NOR2_X1    g09827(.A1(new_n10019_), .A2(new_n10018_), .ZN(new_n10020_));
  OAI21_X1   g09828(.A1(new_n10020_), .A2(new_n10014_), .B(\asqrt[44] ), .ZN(new_n10021_));
  NOR2_X1    g09829(.A1(new_n9458_), .A2(new_n9467_), .ZN(new_n10022_));
  NOR3_X1    g09830(.A1(new_n9846_), .A2(new_n9598_), .A3(new_n10022_), .ZN(new_n10023_));
  INV_X1     g09831(.I(new_n10023_), .ZN(new_n10024_));
  NOR3_X1    g09832(.A1(new_n10022_), .A2(new_n9598_), .A3(new_n9466_), .ZN(new_n10025_));
  AOI22_X1   g09833(.A1(new_n10024_), .A2(new_n9466_), .B1(\asqrt[25] ), .B2(new_n10025_), .ZN(new_n10026_));
  INV_X1     g09834(.I(new_n10026_), .ZN(new_n10027_));
  NAND2_X1   g09835(.A1(new_n10013_), .A2(new_n2954_), .ZN(new_n10028_));
  OAI21_X1   g09836(.A1(new_n10020_), .A2(new_n10028_), .B(new_n10027_), .ZN(new_n10029_));
  AOI21_X1   g09837(.A1(new_n10029_), .A2(new_n10021_), .B(new_n2641_), .ZN(new_n10030_));
  INV_X1     g09838(.I(new_n9474_), .ZN(new_n10031_));
  NOR3_X1    g09839(.A1(new_n9469_), .A2(new_n9607_), .A3(new_n10031_), .ZN(new_n10032_));
  NOR3_X1    g09840(.A1(new_n9846_), .A2(new_n9469_), .A3(new_n9607_), .ZN(new_n10033_));
  INV_X1     g09841(.I(new_n10033_), .ZN(new_n10034_));
  AOI22_X1   g09842(.A1(new_n10034_), .A2(new_n10031_), .B1(\asqrt[25] ), .B2(new_n10032_), .ZN(new_n10035_));
  OAI21_X1   g09843(.A1(new_n10018_), .A2(new_n10019_), .B(new_n10013_), .ZN(new_n10036_));
  AOI21_X1   g09844(.A1(new_n10036_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n10037_));
  AOI21_X1   g09845(.A1(new_n10037_), .A2(new_n10029_), .B(new_n10035_), .ZN(new_n10038_));
  OAI21_X1   g09846(.A1(new_n10038_), .A2(new_n10030_), .B(\asqrt[46] ), .ZN(new_n10039_));
  INV_X1     g09847(.I(new_n10039_), .ZN(new_n10040_));
  NOR3_X1    g09848(.A1(new_n9846_), .A2(new_n9479_), .A3(new_n9487_), .ZN(new_n10041_));
  INV_X1     g09849(.I(new_n10041_), .ZN(new_n10042_));
  NOR3_X1    g09850(.A1(new_n9479_), .A2(new_n9541_), .A3(new_n9487_), .ZN(new_n10043_));
  AOI22_X1   g09851(.A1(new_n10042_), .A2(new_n9541_), .B1(\asqrt[25] ), .B2(new_n10043_), .ZN(new_n10044_));
  NOR3_X1    g09852(.A1(new_n10038_), .A2(new_n10030_), .A3(\asqrt[46] ), .ZN(new_n10045_));
  NOR2_X1    g09853(.A1(new_n10045_), .A2(new_n10044_), .ZN(new_n10046_));
  OAI21_X1   g09854(.A1(new_n10046_), .A2(new_n10040_), .B(\asqrt[47] ), .ZN(new_n10047_));
  NOR2_X1    g09855(.A1(new_n9488_), .A2(new_n9497_), .ZN(new_n10048_));
  NOR3_X1    g09856(.A1(new_n10048_), .A2(new_n9606_), .A3(new_n9496_), .ZN(new_n10049_));
  NOR3_X1    g09857(.A1(new_n9846_), .A2(new_n9606_), .A3(new_n10048_), .ZN(new_n10050_));
  INV_X1     g09858(.I(new_n10050_), .ZN(new_n10051_));
  AOI22_X1   g09859(.A1(new_n10051_), .A2(new_n9496_), .B1(\asqrt[25] ), .B2(new_n10049_), .ZN(new_n10052_));
  INV_X1     g09860(.I(new_n10052_), .ZN(new_n10053_));
  NAND2_X1   g09861(.A1(new_n10039_), .A2(new_n2229_), .ZN(new_n10054_));
  OAI21_X1   g09862(.A1(new_n10046_), .A2(new_n10054_), .B(new_n10053_), .ZN(new_n10055_));
  AOI21_X1   g09863(.A1(new_n10055_), .A2(new_n10047_), .B(new_n1956_), .ZN(new_n10056_));
  INV_X1     g09864(.I(new_n9504_), .ZN(new_n10057_));
  NOR3_X1    g09865(.A1(new_n9846_), .A2(new_n9499_), .A3(new_n9615_), .ZN(new_n10058_));
  INV_X1     g09866(.I(new_n10058_), .ZN(new_n10059_));
  NOR3_X1    g09867(.A1(new_n9499_), .A2(new_n9615_), .A3(new_n10057_), .ZN(new_n10060_));
  AOI22_X1   g09868(.A1(new_n10059_), .A2(new_n10057_), .B1(\asqrt[25] ), .B2(new_n10060_), .ZN(new_n10061_));
  OAI21_X1   g09869(.A1(new_n10044_), .A2(new_n10045_), .B(new_n10039_), .ZN(new_n10062_));
  AOI21_X1   g09870(.A1(new_n10062_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n10063_));
  AOI21_X1   g09871(.A1(new_n10063_), .A2(new_n10055_), .B(new_n10061_), .ZN(new_n10064_));
  OAI21_X1   g09872(.A1(new_n10064_), .A2(new_n10056_), .B(\asqrt[49] ), .ZN(new_n10065_));
  INV_X1     g09873(.I(new_n10065_), .ZN(new_n10066_));
  NOR3_X1    g09874(.A1(new_n9509_), .A2(new_n9540_), .A3(new_n9514_), .ZN(new_n10067_));
  NOR3_X1    g09875(.A1(new_n9846_), .A2(new_n9509_), .A3(new_n9514_), .ZN(new_n10068_));
  INV_X1     g09876(.I(new_n10068_), .ZN(new_n10069_));
  AOI22_X1   g09877(.A1(new_n10069_), .A2(new_n9540_), .B1(\asqrt[25] ), .B2(new_n10067_), .ZN(new_n10070_));
  NOR3_X1    g09878(.A1(new_n10064_), .A2(new_n10056_), .A3(\asqrt[49] ), .ZN(new_n10071_));
  NOR2_X1    g09879(.A1(new_n10071_), .A2(new_n10070_), .ZN(new_n10072_));
  OAI21_X1   g09880(.A1(new_n10072_), .A2(new_n10066_), .B(\asqrt[50] ), .ZN(new_n10073_));
  NOR2_X1    g09881(.A1(new_n9515_), .A2(new_n9523_), .ZN(new_n10074_));
  NOR3_X1    g09882(.A1(new_n9846_), .A2(new_n9614_), .A3(new_n10074_), .ZN(new_n10075_));
  INV_X1     g09883(.I(new_n10075_), .ZN(new_n10076_));
  NOR3_X1    g09884(.A1(new_n10074_), .A2(new_n9614_), .A3(new_n9522_), .ZN(new_n10077_));
  AOI22_X1   g09885(.A1(new_n10076_), .A2(new_n9522_), .B1(\asqrt[25] ), .B2(new_n10077_), .ZN(new_n10078_));
  INV_X1     g09886(.I(new_n10078_), .ZN(new_n10079_));
  NAND2_X1   g09887(.A1(new_n10065_), .A2(new_n1612_), .ZN(new_n10080_));
  OAI21_X1   g09888(.A1(new_n10072_), .A2(new_n10080_), .B(new_n10079_), .ZN(new_n10081_));
  AOI21_X1   g09889(.A1(new_n10081_), .A2(new_n10073_), .B(new_n1376_), .ZN(new_n10082_));
  NOR3_X1    g09890(.A1(new_n9525_), .A2(new_n9628_), .A3(new_n9638_), .ZN(new_n10083_));
  NOR3_X1    g09891(.A1(new_n9846_), .A2(new_n9525_), .A3(new_n9628_), .ZN(new_n10084_));
  INV_X1     g09892(.I(new_n10084_), .ZN(new_n10085_));
  AOI22_X1   g09893(.A1(new_n10085_), .A2(new_n9638_), .B1(\asqrt[25] ), .B2(new_n10083_), .ZN(new_n10086_));
  OAI21_X1   g09894(.A1(new_n10070_), .A2(new_n10071_), .B(new_n10065_), .ZN(new_n10087_));
  AOI21_X1   g09895(.A1(new_n10087_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n10088_));
  AOI21_X1   g09896(.A1(new_n10088_), .A2(new_n10081_), .B(new_n10086_), .ZN(new_n10089_));
  OAI21_X1   g09897(.A1(new_n10089_), .A2(new_n10082_), .B(\asqrt[52] ), .ZN(new_n10090_));
  INV_X1     g09898(.I(new_n10090_), .ZN(new_n10091_));
  INV_X1     g09899(.I(new_n10089_), .ZN(new_n10092_));
  NOR3_X1    g09900(.A1(new_n9846_), .A2(new_n9641_), .A3(new_n9667_), .ZN(new_n10093_));
  INV_X1     g09901(.I(new_n10093_), .ZN(new_n10094_));
  NOR3_X1    g09902(.A1(new_n9641_), .A2(new_n9539_), .A3(new_n9667_), .ZN(new_n10095_));
  AOI22_X1   g09903(.A1(new_n10094_), .A2(new_n9539_), .B1(\asqrt[25] ), .B2(new_n10095_), .ZN(new_n10096_));
  NOR2_X1    g09904(.A1(new_n10082_), .A2(\asqrt[52] ), .ZN(new_n10097_));
  AOI21_X1   g09905(.A1(new_n10092_), .A2(new_n10097_), .B(new_n10096_), .ZN(new_n10098_));
  OAI21_X1   g09906(.A1(new_n10098_), .A2(new_n10091_), .B(\asqrt[53] ), .ZN(new_n10099_));
  NOR2_X1    g09907(.A1(new_n9655_), .A2(new_n9643_), .ZN(new_n10100_));
  NOR3_X1    g09908(.A1(new_n10100_), .A2(new_n9622_), .A3(new_n9654_), .ZN(new_n10101_));
  NOR3_X1    g09909(.A1(new_n9846_), .A2(new_n9622_), .A3(new_n10100_), .ZN(new_n10102_));
  INV_X1     g09910(.I(new_n10102_), .ZN(new_n10103_));
  AOI22_X1   g09911(.A1(new_n10103_), .A2(new_n9654_), .B1(\asqrt[25] ), .B2(new_n10101_), .ZN(new_n10104_));
  INV_X1     g09912(.I(new_n10104_), .ZN(new_n10105_));
  NAND2_X1   g09913(.A1(new_n10090_), .A2(new_n1103_), .ZN(new_n10106_));
  OAI21_X1   g09914(.A1(new_n10106_), .A2(new_n10098_), .B(new_n10105_), .ZN(new_n10107_));
  AOI21_X1   g09915(.A1(new_n10107_), .A2(new_n10099_), .B(new_n904_), .ZN(new_n10108_));
  INV_X1     g09916(.I(new_n10108_), .ZN(new_n10109_));
  INV_X1     g09917(.I(new_n10107_), .ZN(new_n10110_));
  NOR3_X1    g09918(.A1(new_n9846_), .A2(new_n9657_), .A3(new_n9694_), .ZN(new_n10111_));
  INV_X1     g09919(.I(new_n10111_), .ZN(new_n10112_));
  NOR3_X1    g09920(.A1(new_n9694_), .A2(new_n9657_), .A3(new_n9637_), .ZN(new_n10113_));
  AOI22_X1   g09921(.A1(new_n10112_), .A2(new_n9637_), .B1(\asqrt[25] ), .B2(new_n10113_), .ZN(new_n10114_));
  INV_X1     g09922(.I(new_n10114_), .ZN(new_n10115_));
  NAND2_X1   g09923(.A1(new_n10099_), .A2(new_n904_), .ZN(new_n10116_));
  OAI21_X1   g09924(.A1(new_n10116_), .A2(new_n10110_), .B(new_n10115_), .ZN(new_n10117_));
  AOI21_X1   g09925(.A1(new_n10117_), .A2(new_n10109_), .B(new_n823_), .ZN(new_n10118_));
  NOR3_X1    g09926(.A1(new_n9647_), .A2(new_n9679_), .A3(new_n9690_), .ZN(new_n10119_));
  NOR3_X1    g09927(.A1(new_n9846_), .A2(new_n9647_), .A3(new_n9679_), .ZN(new_n10120_));
  INV_X1     g09928(.I(new_n10120_), .ZN(new_n10121_));
  AOI22_X1   g09929(.A1(new_n10121_), .A2(new_n9690_), .B1(\asqrt[25] ), .B2(new_n10119_), .ZN(new_n10122_));
  NOR2_X1    g09930(.A1(new_n10108_), .A2(\asqrt[55] ), .ZN(new_n10123_));
  AOI21_X1   g09931(.A1(new_n10123_), .A2(new_n10117_), .B(new_n10122_), .ZN(new_n10124_));
  OAI21_X1   g09932(.A1(new_n10124_), .A2(new_n10118_), .B(\asqrt[56] ), .ZN(new_n10125_));
  NOR2_X1    g09933(.A1(new_n9672_), .A2(new_n9659_), .ZN(new_n10126_));
  NOR3_X1    g09934(.A1(new_n9846_), .A2(new_n9693_), .A3(new_n10126_), .ZN(new_n10127_));
  INV_X1     g09935(.I(new_n10127_), .ZN(new_n10128_));
  NOR3_X1    g09936(.A1(new_n10126_), .A2(new_n9693_), .A3(new_n9666_), .ZN(new_n10129_));
  AOI22_X1   g09937(.A1(new_n10128_), .A2(new_n9666_), .B1(\asqrt[25] ), .B2(new_n10129_), .ZN(new_n10130_));
  INV_X1     g09938(.I(new_n10130_), .ZN(new_n10131_));
  NOR3_X1    g09939(.A1(new_n10089_), .A2(new_n10082_), .A3(\asqrt[52] ), .ZN(new_n10132_));
  OAI21_X1   g09940(.A1(new_n10096_), .A2(new_n10132_), .B(new_n10090_), .ZN(new_n10133_));
  AOI21_X1   g09941(.A1(new_n10133_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n10134_));
  AOI21_X1   g09942(.A1(new_n10134_), .A2(new_n10107_), .B(new_n10114_), .ZN(new_n10135_));
  OAI21_X1   g09943(.A1(new_n10135_), .A2(new_n10108_), .B(\asqrt[55] ), .ZN(new_n10136_));
  NAND2_X1   g09944(.A1(new_n10136_), .A2(new_n703_), .ZN(new_n10137_));
  OAI21_X1   g09945(.A1(new_n10137_), .A2(new_n10124_), .B(new_n10131_), .ZN(new_n10138_));
  AOI21_X1   g09946(.A1(new_n10138_), .A2(new_n10125_), .B(new_n531_), .ZN(new_n10139_));
  INV_X1     g09947(.I(new_n10139_), .ZN(new_n10140_));
  INV_X1     g09948(.I(new_n10138_), .ZN(new_n10141_));
  NOR3_X1    g09949(.A1(new_n9707_), .A2(new_n9674_), .A3(new_n9717_), .ZN(new_n10142_));
  NOR3_X1    g09950(.A1(new_n9846_), .A2(new_n9674_), .A3(new_n9707_), .ZN(new_n10143_));
  INV_X1     g09951(.I(new_n10143_), .ZN(new_n10144_));
  AOI22_X1   g09952(.A1(new_n10144_), .A2(new_n9717_), .B1(\asqrt[25] ), .B2(new_n10142_), .ZN(new_n10145_));
  INV_X1     g09953(.I(new_n10145_), .ZN(new_n10146_));
  NAND2_X1   g09954(.A1(new_n10125_), .A2(new_n531_), .ZN(new_n10147_));
  OAI21_X1   g09955(.A1(new_n10147_), .A2(new_n10141_), .B(new_n10146_), .ZN(new_n10148_));
  AOI21_X1   g09956(.A1(new_n10148_), .A2(new_n10140_), .B(new_n436_), .ZN(new_n10149_));
  NOR3_X1    g09957(.A1(new_n9846_), .A2(new_n9720_), .A3(new_n9745_), .ZN(new_n10150_));
  INV_X1     g09958(.I(new_n10150_), .ZN(new_n10151_));
  NOR3_X1    g09959(.A1(new_n9720_), .A2(new_n9745_), .A3(new_n9689_), .ZN(new_n10152_));
  AOI22_X1   g09960(.A1(new_n10151_), .A2(new_n9689_), .B1(\asqrt[25] ), .B2(new_n10152_), .ZN(new_n10153_));
  NOR2_X1    g09961(.A1(new_n10139_), .A2(\asqrt[58] ), .ZN(new_n10154_));
  AOI21_X1   g09962(.A1(new_n10154_), .A2(new_n10148_), .B(new_n10153_), .ZN(new_n10155_));
  OAI21_X1   g09963(.A1(new_n10155_), .A2(new_n10149_), .B(\asqrt[59] ), .ZN(new_n10156_));
  NOR2_X1    g09964(.A1(new_n9733_), .A2(new_n9722_), .ZN(new_n10157_));
  NOR3_X1    g09965(.A1(new_n10157_), .A2(new_n9701_), .A3(new_n9732_), .ZN(new_n10158_));
  NOR3_X1    g09966(.A1(new_n9846_), .A2(new_n9701_), .A3(new_n10157_), .ZN(new_n10159_));
  INV_X1     g09967(.I(new_n10159_), .ZN(new_n10160_));
  AOI22_X1   g09968(.A1(new_n10160_), .A2(new_n9732_), .B1(\asqrt[25] ), .B2(new_n10158_), .ZN(new_n10161_));
  INV_X1     g09969(.I(new_n10161_), .ZN(new_n10162_));
  NOR3_X1    g09970(.A1(new_n10135_), .A2(\asqrt[55] ), .A3(new_n10108_), .ZN(new_n10163_));
  OAI21_X1   g09971(.A1(new_n10122_), .A2(new_n10163_), .B(new_n10136_), .ZN(new_n10164_));
  AOI21_X1   g09972(.A1(new_n10164_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n10165_));
  AOI21_X1   g09973(.A1(new_n10165_), .A2(new_n10138_), .B(new_n10145_), .ZN(new_n10166_));
  OAI21_X1   g09974(.A1(new_n10166_), .A2(new_n10139_), .B(\asqrt[58] ), .ZN(new_n10167_));
  NAND2_X1   g09975(.A1(new_n10167_), .A2(new_n327_), .ZN(new_n10168_));
  OAI21_X1   g09976(.A1(new_n10168_), .A2(new_n10155_), .B(new_n10162_), .ZN(new_n10169_));
  AOI21_X1   g09977(.A1(new_n10169_), .A2(new_n10156_), .B(new_n306_), .ZN(new_n10170_));
  INV_X1     g09978(.I(new_n10170_), .ZN(new_n10171_));
  INV_X1     g09979(.I(new_n10169_), .ZN(new_n10172_));
  NOR3_X1    g09980(.A1(new_n9846_), .A2(new_n9735_), .A3(new_n9795_), .ZN(new_n10173_));
  INV_X1     g09981(.I(new_n10173_), .ZN(new_n10174_));
  NOR3_X1    g09982(.A1(new_n9795_), .A2(new_n9735_), .A3(new_n9716_), .ZN(new_n10175_));
  AOI22_X1   g09983(.A1(new_n10174_), .A2(new_n9716_), .B1(\asqrt[25] ), .B2(new_n10175_), .ZN(new_n10176_));
  INV_X1     g09984(.I(new_n10176_), .ZN(new_n10177_));
  NAND2_X1   g09985(.A1(new_n10156_), .A2(new_n306_), .ZN(new_n10178_));
  OAI21_X1   g09986(.A1(new_n10172_), .A2(new_n10178_), .B(new_n10177_), .ZN(new_n10179_));
  AOI21_X1   g09987(.A1(new_n10179_), .A2(new_n10171_), .B(new_n218_), .ZN(new_n10180_));
  NOR3_X1    g09988(.A1(new_n9726_), .A2(new_n9757_), .A3(new_n9791_), .ZN(new_n10181_));
  NOR3_X1    g09989(.A1(new_n9846_), .A2(new_n9726_), .A3(new_n9757_), .ZN(new_n10182_));
  INV_X1     g09990(.I(new_n10182_), .ZN(new_n10183_));
  AOI22_X1   g09991(.A1(new_n10183_), .A2(new_n9791_), .B1(\asqrt[25] ), .B2(new_n10181_), .ZN(new_n10184_));
  NOR2_X1    g09992(.A1(new_n10170_), .A2(\asqrt[61] ), .ZN(new_n10185_));
  AOI21_X1   g09993(.A1(new_n10185_), .A2(new_n10179_), .B(new_n10184_), .ZN(new_n10186_));
  OAI21_X1   g09994(.A1(new_n10186_), .A2(new_n10180_), .B(\asqrt[62] ), .ZN(new_n10187_));
  NOR2_X1    g09995(.A1(new_n9750_), .A2(new_n9737_), .ZN(new_n10188_));
  NOR3_X1    g09996(.A1(new_n9846_), .A2(new_n9794_), .A3(new_n10188_), .ZN(new_n10189_));
  INV_X1     g09997(.I(new_n10189_), .ZN(new_n10190_));
  NOR3_X1    g09998(.A1(new_n10188_), .A2(new_n9794_), .A3(new_n9744_), .ZN(new_n10191_));
  AOI22_X1   g09999(.A1(new_n10190_), .A2(new_n9744_), .B1(\asqrt[25] ), .B2(new_n10191_), .ZN(new_n10192_));
  INV_X1     g10000(.I(new_n10192_), .ZN(new_n10193_));
  NOR3_X1    g10001(.A1(new_n10166_), .A2(\asqrt[58] ), .A3(new_n10139_), .ZN(new_n10194_));
  OAI21_X1   g10002(.A1(new_n10153_), .A2(new_n10194_), .B(new_n10167_), .ZN(new_n10195_));
  AOI21_X1   g10003(.A1(new_n10195_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n10196_));
  AOI21_X1   g10004(.A1(new_n10196_), .A2(new_n10169_), .B(new_n10176_), .ZN(new_n10197_));
  OAI21_X1   g10005(.A1(new_n10197_), .A2(new_n10170_), .B(\asqrt[61] ), .ZN(new_n10198_));
  NAND2_X1   g10006(.A1(new_n10198_), .A2(new_n207_), .ZN(new_n10199_));
  OAI21_X1   g10007(.A1(new_n10199_), .A2(new_n10186_), .B(new_n10193_), .ZN(new_n10200_));
  NAND4_X1   g10008(.A1(\asqrt[25] ), .A2(new_n9799_), .A3(new_n9756_), .A4(new_n9772_), .ZN(new_n10201_));
  NAND2_X1   g10009(.A1(new_n9799_), .A2(new_n9772_), .ZN(new_n10202_));
  OAI21_X1   g10010(.A1(new_n9846_), .A2(new_n10202_), .B(new_n9771_), .ZN(new_n10203_));
  NAND2_X1   g10011(.A1(new_n10203_), .A2(new_n10201_), .ZN(new_n10204_));
  AOI21_X1   g10012(.A1(new_n9773_), .A2(new_n9799_), .B(new_n9766_), .ZN(new_n10205_));
  AOI21_X1   g10013(.A1(\asqrt[25] ), .A2(new_n10205_), .B(new_n9824_), .ZN(new_n10206_));
  NAND2_X1   g10014(.A1(new_n10204_), .A2(new_n10206_), .ZN(new_n10207_));
  AOI21_X1   g10015(.A1(new_n10200_), .A2(new_n10187_), .B(new_n10207_), .ZN(new_n10208_));
  NOR2_X1    g10016(.A1(new_n10208_), .A2(\asqrt[63] ), .ZN(new_n10209_));
  INV_X1     g10017(.I(new_n10200_), .ZN(new_n10210_));
  INV_X1     g10018(.I(new_n10204_), .ZN(new_n10211_));
  NAND2_X1   g10019(.A1(new_n10187_), .A2(new_n10211_), .ZN(new_n10212_));
  AOI21_X1   g10020(.A1(\asqrt[25] ), .A2(new_n9774_), .B(new_n9801_), .ZN(new_n10213_));
  OR3_X2     g10021(.A1(new_n10213_), .A2(new_n193_), .A3(new_n10205_), .Z(new_n10214_));
  NAND2_X1   g10022(.A1(new_n9762_), .A2(new_n9781_), .ZN(new_n10215_));
  NOR4_X1    g10023(.A1(new_n9824_), .A2(new_n9765_), .A3(new_n9778_), .A4(new_n10215_), .ZN(new_n10216_));
  NAND2_X1   g10024(.A1(new_n10216_), .A2(new_n9770_), .ZN(new_n10217_));
  NAND2_X1   g10025(.A1(new_n10214_), .A2(new_n10217_), .ZN(new_n10218_));
  INV_X1     g10026(.I(new_n10218_), .ZN(new_n10219_));
  OAI21_X1   g10027(.A1(new_n10210_), .A2(new_n10212_), .B(new_n10219_), .ZN(new_n10220_));
  NOR2_X1    g10028(.A1(new_n10209_), .A2(new_n10220_), .ZN(new_n10221_));
  INV_X1     g10029(.I(\a[48] ), .ZN(new_n10222_));
  NOR2_X1    g10030(.A1(\a[46] ), .A2(\a[47] ), .ZN(new_n10223_));
  INV_X1     g10031(.I(new_n10223_), .ZN(new_n10224_));
  NOR2_X1    g10032(.A1(new_n10224_), .A2(\a[48] ), .ZN(new_n10225_));
  INV_X1     g10033(.I(new_n10225_), .ZN(new_n10226_));
  OAI21_X1   g10034(.A1(new_n10221_), .A2(new_n10222_), .B(new_n10226_), .ZN(new_n10227_));
  NAND2_X1   g10035(.A1(new_n9781_), .A2(new_n10226_), .ZN(new_n10228_));
  NOR4_X1    g10036(.A1(new_n9824_), .A2(new_n9802_), .A3(new_n9778_), .A4(new_n10228_), .ZN(new_n10229_));
  OAI21_X1   g10037(.A1(new_n10221_), .A2(new_n10222_), .B(new_n10229_), .ZN(new_n10230_));
  NOR3_X1    g10038(.A1(new_n10197_), .A2(\asqrt[61] ), .A3(new_n10170_), .ZN(new_n10231_));
  OAI21_X1   g10039(.A1(new_n10184_), .A2(new_n10231_), .B(new_n10198_), .ZN(new_n10232_));
  INV_X1     g10040(.I(new_n10184_), .ZN(new_n10233_));
  INV_X1     g10041(.I(new_n10153_), .ZN(new_n10234_));
  INV_X1     g10042(.I(new_n10122_), .ZN(new_n10235_));
  INV_X1     g10043(.I(new_n10096_), .ZN(new_n10236_));
  INV_X1     g10044(.I(new_n10070_), .ZN(new_n10237_));
  INV_X1     g10045(.I(new_n10044_), .ZN(new_n10238_));
  INV_X1     g10046(.I(new_n10018_), .ZN(new_n10239_));
  INV_X1     g10047(.I(new_n9989_), .ZN(new_n10240_));
  NOR3_X1    g10048(.A1(new_n9988_), .A2(new_n9969_), .A3(\asqrt[41] ), .ZN(new_n10241_));
  NOR2_X1    g10049(.A1(new_n10241_), .A2(new_n9994_), .ZN(new_n10242_));
  OAI21_X1   g10050(.A1(new_n10242_), .A2(new_n10240_), .B(\asqrt[42] ), .ZN(new_n10243_));
  NAND2_X1   g10051(.A1(new_n10243_), .A2(new_n3218_), .ZN(new_n10244_));
  OAI21_X1   g10052(.A1(new_n10244_), .A2(new_n10012_), .B(new_n10239_), .ZN(new_n10245_));
  NAND3_X1   g10053(.A1(new_n10245_), .A2(new_n2954_), .A3(new_n10013_), .ZN(new_n10246_));
  AOI22_X1   g10054(.A1(new_n10246_), .A2(new_n10027_), .B1(\asqrt[44] ), .B2(new_n10036_), .ZN(new_n10247_));
  OAI21_X1   g10055(.A1(new_n10247_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n10248_));
  OAI21_X1   g10056(.A1(new_n10248_), .A2(new_n10038_), .B(new_n10238_), .ZN(new_n10249_));
  NAND3_X1   g10057(.A1(new_n10249_), .A2(new_n2229_), .A3(new_n10039_), .ZN(new_n10250_));
  AOI22_X1   g10058(.A1(new_n10250_), .A2(new_n10053_), .B1(\asqrt[47] ), .B2(new_n10062_), .ZN(new_n10251_));
  OAI21_X1   g10059(.A1(new_n10251_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n10252_));
  OAI21_X1   g10060(.A1(new_n10252_), .A2(new_n10064_), .B(new_n10237_), .ZN(new_n10253_));
  NAND3_X1   g10061(.A1(new_n10253_), .A2(new_n1612_), .A3(new_n10065_), .ZN(new_n10254_));
  AOI22_X1   g10062(.A1(new_n10254_), .A2(new_n10079_), .B1(\asqrt[50] ), .B2(new_n10087_), .ZN(new_n10255_));
  OAI21_X1   g10063(.A1(new_n10255_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n10256_));
  OAI21_X1   g10064(.A1(new_n10256_), .A2(new_n10089_), .B(new_n10236_), .ZN(new_n10257_));
  NAND3_X1   g10065(.A1(new_n10257_), .A2(new_n1103_), .A3(new_n10090_), .ZN(new_n10258_));
  AOI22_X1   g10066(.A1(new_n10258_), .A2(new_n10105_), .B1(\asqrt[53] ), .B2(new_n10133_), .ZN(new_n10259_));
  OAI21_X1   g10067(.A1(new_n10259_), .A2(new_n904_), .B(new_n823_), .ZN(new_n10260_));
  OAI21_X1   g10068(.A1(new_n10260_), .A2(new_n10135_), .B(new_n10235_), .ZN(new_n10261_));
  NAND3_X1   g10069(.A1(new_n10261_), .A2(new_n703_), .A3(new_n10136_), .ZN(new_n10262_));
  AOI22_X1   g10070(.A1(new_n10262_), .A2(new_n10131_), .B1(\asqrt[56] ), .B2(new_n10164_), .ZN(new_n10263_));
  OAI21_X1   g10071(.A1(new_n10263_), .A2(new_n531_), .B(new_n436_), .ZN(new_n10264_));
  OAI21_X1   g10072(.A1(new_n10264_), .A2(new_n10166_), .B(new_n10234_), .ZN(new_n10265_));
  NAND3_X1   g10073(.A1(new_n10265_), .A2(new_n327_), .A3(new_n10167_), .ZN(new_n10266_));
  AOI22_X1   g10074(.A1(new_n10266_), .A2(new_n10162_), .B1(new_n10195_), .B2(\asqrt[59] ), .ZN(new_n10267_));
  OAI21_X1   g10075(.A1(new_n10267_), .A2(new_n306_), .B(new_n218_), .ZN(new_n10268_));
  OAI21_X1   g10076(.A1(new_n10268_), .A2(new_n10197_), .B(new_n10233_), .ZN(new_n10269_));
  NAND3_X1   g10077(.A1(new_n10269_), .A2(new_n207_), .A3(new_n10198_), .ZN(new_n10270_));
  AOI22_X1   g10078(.A1(new_n10270_), .A2(new_n10193_), .B1(new_n10232_), .B2(\asqrt[62] ), .ZN(new_n10271_));
  OAI21_X1   g10079(.A1(new_n10271_), .A2(new_n10207_), .B(new_n193_), .ZN(new_n10272_));
  AOI21_X1   g10080(.A1(new_n10232_), .A2(\asqrt[62] ), .B(new_n10204_), .ZN(new_n10273_));
  AOI21_X1   g10081(.A1(new_n10273_), .A2(new_n10200_), .B(new_n10218_), .ZN(new_n10274_));
  AOI21_X1   g10082(.A1(new_n10272_), .A2(new_n10274_), .B(new_n9788_), .ZN(new_n10275_));
  OAI21_X1   g10083(.A1(new_n10209_), .A2(new_n10220_), .B(new_n10222_), .ZN(new_n10276_));
  AOI21_X1   g10084(.A1(\a[49] ), .A2(new_n10276_), .B(new_n10275_), .ZN(new_n10277_));
  AOI22_X1   g10085(.A1(new_n10277_), .A2(new_n10230_), .B1(\asqrt[25] ), .B2(new_n10227_), .ZN(new_n10278_));
  NOR2_X1    g10086(.A1(new_n10278_), .A2(new_n9317_), .ZN(new_n10279_));
  NAND2_X1   g10087(.A1(new_n10277_), .A2(new_n10230_), .ZN(new_n10280_));
  OAI21_X1   g10088(.A1(new_n10209_), .A2(new_n10220_), .B(new_n9787_), .ZN(new_n10281_));
  NAND2_X1   g10089(.A1(new_n10273_), .A2(new_n10200_), .ZN(new_n10282_));
  OAI21_X1   g10090(.A1(new_n10216_), .A2(new_n9785_), .B(new_n9770_), .ZN(new_n10283_));
  NAND4_X1   g10091(.A1(new_n10272_), .A2(new_n10282_), .A3(new_n10214_), .A4(new_n10283_), .ZN(new_n10284_));
  AOI21_X1   g10092(.A1(new_n10284_), .A2(new_n10281_), .B(new_n9807_), .ZN(new_n10285_));
  INV_X1     g10093(.I(new_n10282_), .ZN(new_n10286_));
  NAND2_X1   g10094(.A1(new_n10214_), .A2(new_n10283_), .ZN(new_n10287_));
  NOR3_X1    g10095(.A1(new_n10286_), .A2(new_n10209_), .A3(new_n10287_), .ZN(new_n10288_));
  NOR3_X1    g10096(.A1(new_n10288_), .A2(new_n10275_), .A3(\a[50] ), .ZN(new_n10289_));
  NOR2_X1    g10097(.A1(new_n10285_), .A2(new_n10289_), .ZN(new_n10290_));
  AOI21_X1   g10098(.A1(new_n10227_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n10291_));
  AOI21_X1   g10099(.A1(new_n10280_), .A2(new_n10291_), .B(new_n10290_), .ZN(new_n10292_));
  OAI21_X1   g10100(.A1(new_n10292_), .A2(new_n10279_), .B(\asqrt[27] ), .ZN(new_n10293_));
  OAI21_X1   g10101(.A1(\asqrt[63] ), .A2(new_n10208_), .B(new_n10274_), .ZN(\asqrt[24] ));
  NOR3_X1    g10102(.A1(new_n9890_), .A2(new_n9806_), .A3(new_n9812_), .ZN(new_n10295_));
  NAND3_X1   g10103(.A1(\asqrt[24] ), .A2(new_n9828_), .A3(new_n9875_), .ZN(new_n10296_));
  AOI22_X1   g10104(.A1(new_n10296_), .A2(new_n9890_), .B1(\asqrt[24] ), .B2(new_n10295_), .ZN(new_n10297_));
  INV_X1     g10105(.I(new_n10297_), .ZN(new_n10298_));
  OAI21_X1   g10106(.A1(new_n10278_), .A2(new_n9317_), .B(new_n8826_), .ZN(new_n10299_));
  OAI21_X1   g10107(.A1(new_n10299_), .A2(new_n10292_), .B(new_n10298_), .ZN(new_n10300_));
  AOI21_X1   g10108(.A1(new_n10300_), .A2(new_n10293_), .B(new_n8483_), .ZN(new_n10301_));
  NOR2_X1    g10109(.A1(new_n9827_), .A2(new_n9823_), .ZN(new_n10302_));
  NOR2_X1    g10110(.A1(new_n9816_), .A2(new_n9829_), .ZN(new_n10303_));
  INV_X1     g10111(.I(new_n10303_), .ZN(new_n10304_));
  NAND4_X1   g10112(.A1(\asqrt[24] ), .A2(new_n9817_), .A3(new_n10302_), .A4(new_n10304_), .ZN(new_n10305_));
  NOR3_X1    g10113(.A1(new_n10221_), .A2(new_n9879_), .A3(new_n10303_), .ZN(new_n10306_));
  OAI21_X1   g10114(.A1(new_n10306_), .A2(new_n10302_), .B(new_n10305_), .ZN(new_n10307_));
  INV_X1     g10115(.I(new_n10307_), .ZN(new_n10308_));
  AOI21_X1   g10116(.A1(new_n10272_), .A2(new_n10274_), .B(new_n10222_), .ZN(new_n10309_));
  OAI21_X1   g10117(.A1(new_n10309_), .A2(new_n10225_), .B(\asqrt[25] ), .ZN(new_n10310_));
  INV_X1     g10118(.I(new_n10310_), .ZN(new_n10311_));
  INV_X1     g10119(.I(new_n10229_), .ZN(new_n10312_));
  NOR2_X1    g10120(.A1(new_n10309_), .A2(new_n10312_), .ZN(new_n10313_));
  INV_X1     g10121(.I(\a[49] ), .ZN(new_n10314_));
  AOI21_X1   g10122(.A1(\asqrt[24] ), .A2(new_n10222_), .B(new_n10314_), .ZN(new_n10315_));
  NOR3_X1    g10123(.A1(new_n10313_), .A2(new_n10315_), .A3(new_n10275_), .ZN(new_n10316_));
  OAI21_X1   g10124(.A1(new_n10316_), .A2(new_n10311_), .B(\asqrt[26] ), .ZN(new_n10317_));
  AOI21_X1   g10125(.A1(\asqrt[24] ), .A2(\a[48] ), .B(new_n10225_), .ZN(new_n10318_));
  OAI21_X1   g10126(.A1(new_n10318_), .A2(new_n9846_), .B(new_n9317_), .ZN(new_n10319_));
  OAI22_X1   g10127(.A1(new_n10316_), .A2(new_n10319_), .B1(new_n10285_), .B2(new_n10289_), .ZN(new_n10320_));
  AOI21_X1   g10128(.A1(new_n10320_), .A2(new_n10317_), .B(new_n8826_), .ZN(new_n10321_));
  AOI21_X1   g10129(.A1(new_n10272_), .A2(new_n10274_), .B(\a[48] ), .ZN(new_n10322_));
  OAI21_X1   g10130(.A1(new_n10314_), .A2(new_n10322_), .B(new_n10281_), .ZN(new_n10323_));
  OAI21_X1   g10131(.A1(new_n10323_), .A2(new_n10313_), .B(new_n10310_), .ZN(new_n10324_));
  AOI21_X1   g10132(.A1(new_n10324_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n10325_));
  AOI21_X1   g10133(.A1(new_n10325_), .A2(new_n10320_), .B(new_n10297_), .ZN(new_n10326_));
  NOR3_X1    g10134(.A1(new_n10326_), .A2(new_n10321_), .A3(\asqrt[28] ), .ZN(new_n10327_));
  NOR2_X1    g10135(.A1(new_n10327_), .A2(new_n10308_), .ZN(new_n10328_));
  OAI21_X1   g10136(.A1(new_n10328_), .A2(new_n10301_), .B(\asqrt[29] ), .ZN(new_n10329_));
  NOR2_X1    g10137(.A1(new_n9892_), .A2(new_n9884_), .ZN(new_n10330_));
  NOR3_X1    g10138(.A1(new_n10221_), .A2(new_n9831_), .A3(new_n10330_), .ZN(new_n10331_));
  INV_X1     g10139(.I(new_n10331_), .ZN(new_n10332_));
  NOR3_X1    g10140(.A1(new_n10330_), .A2(new_n9831_), .A3(new_n9889_), .ZN(new_n10333_));
  AOI22_X1   g10141(.A1(new_n10332_), .A2(new_n9889_), .B1(\asqrt[24] ), .B2(new_n10333_), .ZN(new_n10334_));
  INV_X1     g10142(.I(new_n10334_), .ZN(new_n10335_));
  OAI21_X1   g10143(.A1(new_n10326_), .A2(new_n10321_), .B(\asqrt[28] ), .ZN(new_n10336_));
  NAND2_X1   g10144(.A1(new_n10336_), .A2(new_n8036_), .ZN(new_n10337_));
  OAI21_X1   g10145(.A1(new_n10328_), .A2(new_n10337_), .B(new_n10335_), .ZN(new_n10338_));
  AOI21_X1   g10146(.A1(new_n10338_), .A2(new_n10329_), .B(new_n7539_), .ZN(new_n10339_));
  NOR3_X1    g10147(.A1(new_n9841_), .A2(new_n9850_), .A3(new_n9848_), .ZN(new_n10340_));
  NOR3_X1    g10148(.A1(new_n10221_), .A2(new_n9841_), .A3(new_n9850_), .ZN(new_n10341_));
  INV_X1     g10149(.I(new_n10341_), .ZN(new_n10342_));
  AOI22_X1   g10150(.A1(new_n10342_), .A2(new_n9848_), .B1(\asqrt[24] ), .B2(new_n10340_), .ZN(new_n10343_));
  OAI21_X1   g10151(.A1(new_n10308_), .A2(new_n10327_), .B(new_n10336_), .ZN(new_n10344_));
  AOI21_X1   g10152(.A1(new_n10344_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n10345_));
  AOI21_X1   g10153(.A1(new_n10345_), .A2(new_n10338_), .B(new_n10343_), .ZN(new_n10346_));
  OAI21_X1   g10154(.A1(new_n10346_), .A2(new_n10339_), .B(\asqrt[31] ), .ZN(new_n10347_));
  INV_X1     g10155(.I(new_n10347_), .ZN(new_n10348_));
  NOR2_X1    g10156(.A1(new_n9851_), .A2(new_n9859_), .ZN(new_n10349_));
  NOR3_X1    g10157(.A1(new_n10221_), .A2(new_n9888_), .A3(new_n10349_), .ZN(new_n10350_));
  INV_X1     g10158(.I(new_n10350_), .ZN(new_n10351_));
  NOR3_X1    g10159(.A1(new_n10349_), .A2(new_n9888_), .A3(new_n9858_), .ZN(new_n10352_));
  AOI22_X1   g10160(.A1(new_n10351_), .A2(new_n9858_), .B1(\asqrt[24] ), .B2(new_n10352_), .ZN(new_n10353_));
  NOR3_X1    g10161(.A1(new_n10346_), .A2(new_n10339_), .A3(\asqrt[31] ), .ZN(new_n10354_));
  NOR2_X1    g10162(.A1(new_n10354_), .A2(new_n10353_), .ZN(new_n10355_));
  OAI21_X1   g10163(.A1(new_n10355_), .A2(new_n10348_), .B(\asqrt[32] ), .ZN(new_n10356_));
  INV_X1     g10164(.I(new_n9865_), .ZN(new_n10357_));
  NOR3_X1    g10165(.A1(new_n9861_), .A2(new_n9975_), .A3(new_n10357_), .ZN(new_n10358_));
  NOR3_X1    g10166(.A1(new_n10221_), .A2(new_n9861_), .A3(new_n9975_), .ZN(new_n10359_));
  INV_X1     g10167(.I(new_n10359_), .ZN(new_n10360_));
  AOI22_X1   g10168(.A1(new_n10360_), .A2(new_n10357_), .B1(\asqrt[24] ), .B2(new_n10358_), .ZN(new_n10361_));
  INV_X1     g10169(.I(new_n10361_), .ZN(new_n10362_));
  NAND2_X1   g10170(.A1(new_n10347_), .A2(new_n6824_), .ZN(new_n10363_));
  OAI21_X1   g10171(.A1(new_n10355_), .A2(new_n10363_), .B(new_n10362_), .ZN(new_n10364_));
  AOI21_X1   g10172(.A1(new_n10364_), .A2(new_n10356_), .B(new_n6356_), .ZN(new_n10365_));
  INV_X1     g10173(.I(new_n9942_), .ZN(new_n10366_));
  NAND3_X1   g10174(.A1(\asqrt[24] ), .A2(new_n9869_), .A3(new_n10366_), .ZN(new_n10367_));
  AND3_X2    g10175(.A1(new_n10366_), .A2(new_n9869_), .A3(new_n9873_), .Z(new_n10368_));
  AOI22_X1   g10176(.A1(new_n10367_), .A2(new_n9874_), .B1(\asqrt[24] ), .B2(new_n10368_), .ZN(new_n10369_));
  OAI21_X1   g10177(.A1(new_n10353_), .A2(new_n10354_), .B(new_n10347_), .ZN(new_n10370_));
  AOI21_X1   g10178(.A1(new_n10370_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n10371_));
  AOI21_X1   g10179(.A1(new_n10371_), .A2(new_n10364_), .B(new_n10369_), .ZN(new_n10372_));
  OAI21_X1   g10180(.A1(new_n10372_), .A2(new_n10365_), .B(\asqrt[34] ), .ZN(new_n10373_));
  INV_X1     g10181(.I(new_n10373_), .ZN(new_n10374_));
  INV_X1     g10182(.I(new_n9944_), .ZN(new_n10375_));
  NOR3_X1    g10183(.A1(new_n10375_), .A2(new_n9900_), .A3(new_n9908_), .ZN(new_n10376_));
  NOR3_X1    g10184(.A1(new_n10221_), .A2(new_n9900_), .A3(new_n10375_), .ZN(new_n10377_));
  INV_X1     g10185(.I(new_n10377_), .ZN(new_n10378_));
  AOI22_X1   g10186(.A1(new_n10378_), .A2(new_n9908_), .B1(\asqrt[24] ), .B2(new_n10376_), .ZN(new_n10379_));
  NOR3_X1    g10187(.A1(new_n10372_), .A2(new_n10365_), .A3(\asqrt[34] ), .ZN(new_n10380_));
  NOR2_X1    g10188(.A1(new_n10380_), .A2(new_n10379_), .ZN(new_n10381_));
  OAI21_X1   g10189(.A1(new_n10381_), .A2(new_n10374_), .B(\asqrt[35] ), .ZN(new_n10382_));
  INV_X1     g10190(.I(new_n9915_), .ZN(new_n10383_));
  NOR3_X1    g10191(.A1(new_n10221_), .A2(new_n9911_), .A3(new_n9979_), .ZN(new_n10384_));
  INV_X1     g10192(.I(new_n10384_), .ZN(new_n10385_));
  NOR3_X1    g10193(.A1(new_n9911_), .A2(new_n10383_), .A3(new_n9979_), .ZN(new_n10386_));
  AOI22_X1   g10194(.A1(new_n10385_), .A2(new_n10383_), .B1(\asqrt[24] ), .B2(new_n10386_), .ZN(new_n10387_));
  INV_X1     g10195(.I(new_n10387_), .ZN(new_n10388_));
  NAND2_X1   g10196(.A1(new_n10373_), .A2(new_n5708_), .ZN(new_n10389_));
  OAI21_X1   g10197(.A1(new_n10381_), .A2(new_n10389_), .B(new_n10388_), .ZN(new_n10390_));
  AOI21_X1   g10198(.A1(new_n10390_), .A2(new_n10382_), .B(new_n5277_), .ZN(new_n10391_));
  NOR3_X1    g10199(.A1(new_n9919_), .A2(new_n9941_), .A3(new_n9925_), .ZN(new_n10392_));
  NOR3_X1    g10200(.A1(new_n10221_), .A2(new_n9919_), .A3(new_n9925_), .ZN(new_n10393_));
  INV_X1     g10201(.I(new_n10393_), .ZN(new_n10394_));
  AOI22_X1   g10202(.A1(new_n10394_), .A2(new_n9941_), .B1(\asqrt[24] ), .B2(new_n10392_), .ZN(new_n10395_));
  OAI21_X1   g10203(.A1(new_n10379_), .A2(new_n10380_), .B(new_n10373_), .ZN(new_n10396_));
  AOI21_X1   g10204(.A1(new_n10396_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n10397_));
  AOI21_X1   g10205(.A1(new_n10397_), .A2(new_n10390_), .B(new_n10395_), .ZN(new_n10398_));
  OAI21_X1   g10206(.A1(new_n10398_), .A2(new_n10391_), .B(\asqrt[37] ), .ZN(new_n10399_));
  INV_X1     g10207(.I(new_n10399_), .ZN(new_n10400_));
  NOR2_X1    g10208(.A1(new_n9926_), .A2(new_n9934_), .ZN(new_n10401_));
  NOR3_X1    g10209(.A1(new_n10221_), .A2(new_n9948_), .A3(new_n10401_), .ZN(new_n10402_));
  INV_X1     g10210(.I(new_n10402_), .ZN(new_n10403_));
  NOR3_X1    g10211(.A1(new_n10401_), .A2(new_n9948_), .A3(new_n9933_), .ZN(new_n10404_));
  AOI22_X1   g10212(.A1(new_n10403_), .A2(new_n9933_), .B1(\asqrt[24] ), .B2(new_n10404_), .ZN(new_n10405_));
  NOR3_X1    g10213(.A1(new_n10398_), .A2(new_n10391_), .A3(\asqrt[37] ), .ZN(new_n10406_));
  NOR2_X1    g10214(.A1(new_n10406_), .A2(new_n10405_), .ZN(new_n10407_));
  OAI21_X1   g10215(.A1(new_n10407_), .A2(new_n10400_), .B(\asqrt[38] ), .ZN(new_n10408_));
  INV_X1     g10216(.I(new_n9940_), .ZN(new_n10409_));
  NOR3_X1    g10217(.A1(new_n9936_), .A2(new_n10409_), .A3(new_n9996_), .ZN(new_n10410_));
  NOR3_X1    g10218(.A1(new_n10221_), .A2(new_n9936_), .A3(new_n9996_), .ZN(new_n10411_));
  INV_X1     g10219(.I(new_n10411_), .ZN(new_n10412_));
  AOI22_X1   g10220(.A1(new_n10412_), .A2(new_n10409_), .B1(\asqrt[24] ), .B2(new_n10410_), .ZN(new_n10413_));
  INV_X1     g10221(.I(new_n10413_), .ZN(new_n10414_));
  NAND2_X1   g10222(.A1(new_n10399_), .A2(new_n4696_), .ZN(new_n10415_));
  OAI21_X1   g10223(.A1(new_n10407_), .A2(new_n10415_), .B(new_n10414_), .ZN(new_n10416_));
  AOI21_X1   g10224(.A1(new_n10416_), .A2(new_n10408_), .B(new_n4298_), .ZN(new_n10417_));
  NOR3_X1    g10225(.A1(new_n10221_), .A2(new_n9952_), .A3(new_n9958_), .ZN(new_n10418_));
  INV_X1     g10226(.I(new_n10418_), .ZN(new_n10419_));
  NOR3_X1    g10227(.A1(new_n9952_), .A2(new_n9974_), .A3(new_n9958_), .ZN(new_n10420_));
  AOI22_X1   g10228(.A1(new_n10419_), .A2(new_n9974_), .B1(\asqrt[24] ), .B2(new_n10420_), .ZN(new_n10421_));
  OAI21_X1   g10229(.A1(new_n10405_), .A2(new_n10406_), .B(new_n10399_), .ZN(new_n10422_));
  AOI21_X1   g10230(.A1(new_n10422_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n10423_));
  AOI21_X1   g10231(.A1(new_n10423_), .A2(new_n10416_), .B(new_n10421_), .ZN(new_n10424_));
  OAI21_X1   g10232(.A1(new_n10424_), .A2(new_n10417_), .B(\asqrt[40] ), .ZN(new_n10425_));
  INV_X1     g10233(.I(new_n10425_), .ZN(new_n10426_));
  NOR2_X1    g10234(.A1(new_n9959_), .A2(new_n9967_), .ZN(new_n10427_));
  NOR3_X1    g10235(.A1(new_n10427_), .A2(new_n9986_), .A3(new_n9966_), .ZN(new_n10428_));
  NOR3_X1    g10236(.A1(new_n10221_), .A2(new_n9986_), .A3(new_n10427_), .ZN(new_n10429_));
  INV_X1     g10237(.I(new_n10429_), .ZN(new_n10430_));
  AOI22_X1   g10238(.A1(new_n10430_), .A2(new_n9966_), .B1(\asqrt[24] ), .B2(new_n10428_), .ZN(new_n10431_));
  NOR3_X1    g10239(.A1(new_n10424_), .A2(new_n10417_), .A3(\asqrt[40] ), .ZN(new_n10432_));
  NOR2_X1    g10240(.A1(new_n10432_), .A2(new_n10431_), .ZN(new_n10433_));
  OAI21_X1   g10241(.A1(new_n10433_), .A2(new_n10426_), .B(\asqrt[41] ), .ZN(new_n10434_));
  INV_X1     g10242(.I(new_n9973_), .ZN(new_n10435_));
  NOR3_X1    g10243(.A1(new_n10221_), .A2(new_n9969_), .A3(new_n10009_), .ZN(new_n10436_));
  INV_X1     g10244(.I(new_n10436_), .ZN(new_n10437_));
  NOR3_X1    g10245(.A1(new_n9969_), .A2(new_n10435_), .A3(new_n10009_), .ZN(new_n10438_));
  AOI22_X1   g10246(.A1(new_n10437_), .A2(new_n10435_), .B1(\asqrt[24] ), .B2(new_n10438_), .ZN(new_n10439_));
  INV_X1     g10247(.I(new_n10439_), .ZN(new_n10440_));
  NAND2_X1   g10248(.A1(new_n10425_), .A2(new_n3782_), .ZN(new_n10441_));
  OAI21_X1   g10249(.A1(new_n10433_), .A2(new_n10441_), .B(new_n10440_), .ZN(new_n10442_));
  AOI21_X1   g10250(.A1(new_n10442_), .A2(new_n10434_), .B(new_n3419_), .ZN(new_n10443_));
  NOR3_X1    g10251(.A1(new_n10240_), .A2(new_n9995_), .A3(new_n10241_), .ZN(new_n10444_));
  NOR3_X1    g10252(.A1(new_n10221_), .A2(new_n10240_), .A3(new_n10241_), .ZN(new_n10445_));
  INV_X1     g10253(.I(new_n10445_), .ZN(new_n10446_));
  AOI22_X1   g10254(.A1(new_n10446_), .A2(new_n9995_), .B1(\asqrt[24] ), .B2(new_n10444_), .ZN(new_n10447_));
  OAI21_X1   g10255(.A1(new_n10431_), .A2(new_n10432_), .B(new_n10425_), .ZN(new_n10448_));
  AOI21_X1   g10256(.A1(new_n10448_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n10449_));
  AOI21_X1   g10257(.A1(new_n10449_), .A2(new_n10442_), .B(new_n10447_), .ZN(new_n10450_));
  OAI21_X1   g10258(.A1(new_n10450_), .A2(new_n10443_), .B(\asqrt[43] ), .ZN(new_n10451_));
  INV_X1     g10259(.I(new_n10451_), .ZN(new_n10452_));
  INV_X1     g10260(.I(new_n10008_), .ZN(new_n10453_));
  NAND2_X1   g10261(.A1(new_n9989_), .A2(new_n3419_), .ZN(new_n10454_));
  NOR2_X1    g10262(.A1(new_n10242_), .A2(new_n10454_), .ZN(new_n10455_));
  NOR3_X1    g10263(.A1(new_n10221_), .A2(new_n10003_), .A3(new_n10455_), .ZN(new_n10456_));
  INV_X1     g10264(.I(new_n10456_), .ZN(new_n10457_));
  NOR3_X1    g10265(.A1(new_n10455_), .A2(new_n10003_), .A3(new_n10453_), .ZN(new_n10458_));
  AOI22_X1   g10266(.A1(new_n10457_), .A2(new_n10453_), .B1(\asqrt[24] ), .B2(new_n10458_), .ZN(new_n10459_));
  NOR3_X1    g10267(.A1(new_n10450_), .A2(new_n10443_), .A3(\asqrt[43] ), .ZN(new_n10460_));
  NOR2_X1    g10268(.A1(new_n10460_), .A2(new_n10459_), .ZN(new_n10461_));
  OAI21_X1   g10269(.A1(new_n10461_), .A2(new_n10452_), .B(\asqrt[44] ), .ZN(new_n10462_));
  NOR3_X1    g10270(.A1(new_n10014_), .A2(new_n10019_), .A3(new_n10239_), .ZN(new_n10463_));
  NOR3_X1    g10271(.A1(new_n10221_), .A2(new_n10014_), .A3(new_n10019_), .ZN(new_n10464_));
  INV_X1     g10272(.I(new_n10464_), .ZN(new_n10465_));
  AOI22_X1   g10273(.A1(new_n10465_), .A2(new_n10239_), .B1(\asqrt[24] ), .B2(new_n10463_), .ZN(new_n10466_));
  INV_X1     g10274(.I(new_n10466_), .ZN(new_n10467_));
  NAND2_X1   g10275(.A1(new_n10451_), .A2(new_n2954_), .ZN(new_n10468_));
  OAI21_X1   g10276(.A1(new_n10461_), .A2(new_n10468_), .B(new_n10467_), .ZN(new_n10469_));
  AOI21_X1   g10277(.A1(new_n10469_), .A2(new_n10462_), .B(new_n2641_), .ZN(new_n10470_));
  INV_X1     g10278(.I(new_n10021_), .ZN(new_n10471_));
  NOR2_X1    g10279(.A1(new_n10020_), .A2(new_n10028_), .ZN(new_n10472_));
  NOR3_X1    g10280(.A1(new_n10221_), .A2(new_n10471_), .A3(new_n10472_), .ZN(new_n10473_));
  INV_X1     g10281(.I(new_n10473_), .ZN(new_n10474_));
  NOR3_X1    g10282(.A1(new_n10471_), .A2(new_n10472_), .A3(new_n10027_), .ZN(new_n10475_));
  AOI22_X1   g10283(.A1(new_n10474_), .A2(new_n10027_), .B1(\asqrt[24] ), .B2(new_n10475_), .ZN(new_n10476_));
  OAI21_X1   g10284(.A1(new_n10459_), .A2(new_n10460_), .B(new_n10451_), .ZN(new_n10477_));
  AOI21_X1   g10285(.A1(new_n10477_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n10478_));
  AOI21_X1   g10286(.A1(new_n10478_), .A2(new_n10469_), .B(new_n10476_), .ZN(new_n10479_));
  OAI21_X1   g10287(.A1(new_n10479_), .A2(new_n10470_), .B(\asqrt[46] ), .ZN(new_n10480_));
  INV_X1     g10288(.I(new_n10480_), .ZN(new_n10481_));
  INV_X1     g10289(.I(new_n10035_), .ZN(new_n10482_));
  INV_X1     g10290(.I(new_n10029_), .ZN(new_n10483_));
  INV_X1     g10291(.I(new_n10037_), .ZN(new_n10484_));
  NOR2_X1    g10292(.A1(new_n10484_), .A2(new_n10483_), .ZN(new_n10485_));
  NOR3_X1    g10293(.A1(new_n10485_), .A2(new_n10030_), .A3(new_n10482_), .ZN(new_n10486_));
  NOR3_X1    g10294(.A1(new_n10221_), .A2(new_n10030_), .A3(new_n10485_), .ZN(new_n10487_));
  INV_X1     g10295(.I(new_n10487_), .ZN(new_n10488_));
  AOI22_X1   g10296(.A1(new_n10488_), .A2(new_n10482_), .B1(\asqrt[24] ), .B2(new_n10486_), .ZN(new_n10489_));
  NOR3_X1    g10297(.A1(new_n10479_), .A2(new_n10470_), .A3(\asqrt[46] ), .ZN(new_n10490_));
  NOR2_X1    g10298(.A1(new_n10490_), .A2(new_n10489_), .ZN(new_n10491_));
  OAI21_X1   g10299(.A1(new_n10491_), .A2(new_n10481_), .B(\asqrt[47] ), .ZN(new_n10492_));
  NOR3_X1    g10300(.A1(new_n10221_), .A2(new_n10040_), .A3(new_n10045_), .ZN(new_n10493_));
  INV_X1     g10301(.I(new_n10493_), .ZN(new_n10494_));
  NOR3_X1    g10302(.A1(new_n10040_), .A2(new_n10238_), .A3(new_n10045_), .ZN(new_n10495_));
  AOI22_X1   g10303(.A1(new_n10494_), .A2(new_n10238_), .B1(\asqrt[24] ), .B2(new_n10495_), .ZN(new_n10496_));
  INV_X1     g10304(.I(new_n10496_), .ZN(new_n10497_));
  NAND2_X1   g10305(.A1(new_n10480_), .A2(new_n2229_), .ZN(new_n10498_));
  OAI21_X1   g10306(.A1(new_n10491_), .A2(new_n10498_), .B(new_n10497_), .ZN(new_n10499_));
  AOI21_X1   g10307(.A1(new_n10499_), .A2(new_n10492_), .B(new_n1956_), .ZN(new_n10500_));
  INV_X1     g10308(.I(new_n10047_), .ZN(new_n10501_));
  NOR2_X1    g10309(.A1(new_n10046_), .A2(new_n10054_), .ZN(new_n10502_));
  NOR3_X1    g10310(.A1(new_n10501_), .A2(new_n10502_), .A3(new_n10053_), .ZN(new_n10503_));
  NOR3_X1    g10311(.A1(new_n10221_), .A2(new_n10501_), .A3(new_n10502_), .ZN(new_n10504_));
  INV_X1     g10312(.I(new_n10504_), .ZN(new_n10505_));
  AOI22_X1   g10313(.A1(new_n10505_), .A2(new_n10053_), .B1(\asqrt[24] ), .B2(new_n10503_), .ZN(new_n10506_));
  OAI21_X1   g10314(.A1(new_n10489_), .A2(new_n10490_), .B(new_n10480_), .ZN(new_n10507_));
  AOI21_X1   g10315(.A1(new_n10507_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n10508_));
  AOI21_X1   g10316(.A1(new_n10508_), .A2(new_n10499_), .B(new_n10506_), .ZN(new_n10509_));
  OAI21_X1   g10317(.A1(new_n10509_), .A2(new_n10500_), .B(\asqrt[49] ), .ZN(new_n10510_));
  INV_X1     g10318(.I(new_n10510_), .ZN(new_n10511_));
  INV_X1     g10319(.I(new_n10061_), .ZN(new_n10512_));
  INV_X1     g10320(.I(new_n10055_), .ZN(new_n10513_));
  INV_X1     g10321(.I(new_n10063_), .ZN(new_n10514_));
  NOR2_X1    g10322(.A1(new_n10514_), .A2(new_n10513_), .ZN(new_n10515_));
  NOR3_X1    g10323(.A1(new_n10221_), .A2(new_n10056_), .A3(new_n10515_), .ZN(new_n10516_));
  INV_X1     g10324(.I(new_n10516_), .ZN(new_n10517_));
  NOR3_X1    g10325(.A1(new_n10515_), .A2(new_n10056_), .A3(new_n10512_), .ZN(new_n10518_));
  AOI22_X1   g10326(.A1(new_n10517_), .A2(new_n10512_), .B1(\asqrt[24] ), .B2(new_n10518_), .ZN(new_n10519_));
  NOR3_X1    g10327(.A1(new_n10509_), .A2(new_n10500_), .A3(\asqrt[49] ), .ZN(new_n10520_));
  NOR2_X1    g10328(.A1(new_n10520_), .A2(new_n10519_), .ZN(new_n10521_));
  OAI21_X1   g10329(.A1(new_n10521_), .A2(new_n10511_), .B(\asqrt[50] ), .ZN(new_n10522_));
  NOR3_X1    g10330(.A1(new_n10066_), .A2(new_n10237_), .A3(new_n10071_), .ZN(new_n10523_));
  NOR3_X1    g10331(.A1(new_n10221_), .A2(new_n10066_), .A3(new_n10071_), .ZN(new_n10524_));
  INV_X1     g10332(.I(new_n10524_), .ZN(new_n10525_));
  AOI22_X1   g10333(.A1(new_n10525_), .A2(new_n10237_), .B1(\asqrt[24] ), .B2(new_n10523_), .ZN(new_n10526_));
  INV_X1     g10334(.I(new_n10526_), .ZN(new_n10527_));
  NAND2_X1   g10335(.A1(new_n10510_), .A2(new_n1612_), .ZN(new_n10528_));
  OAI21_X1   g10336(.A1(new_n10521_), .A2(new_n10528_), .B(new_n10527_), .ZN(new_n10529_));
  AOI21_X1   g10337(.A1(new_n10529_), .A2(new_n10522_), .B(new_n1376_), .ZN(new_n10530_));
  INV_X1     g10338(.I(new_n10073_), .ZN(new_n10531_));
  NOR2_X1    g10339(.A1(new_n10072_), .A2(new_n10080_), .ZN(new_n10532_));
  NOR3_X1    g10340(.A1(new_n10221_), .A2(new_n10531_), .A3(new_n10532_), .ZN(new_n10533_));
  INV_X1     g10341(.I(new_n10533_), .ZN(new_n10534_));
  NOR3_X1    g10342(.A1(new_n10531_), .A2(new_n10079_), .A3(new_n10532_), .ZN(new_n10535_));
  AOI22_X1   g10343(.A1(new_n10534_), .A2(new_n10079_), .B1(\asqrt[24] ), .B2(new_n10535_), .ZN(new_n10536_));
  OAI21_X1   g10344(.A1(new_n10519_), .A2(new_n10520_), .B(new_n10510_), .ZN(new_n10537_));
  AOI21_X1   g10345(.A1(new_n10537_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n10538_));
  AOI21_X1   g10346(.A1(new_n10538_), .A2(new_n10529_), .B(new_n10536_), .ZN(new_n10539_));
  OAI21_X1   g10347(.A1(new_n10539_), .A2(new_n10530_), .B(\asqrt[52] ), .ZN(new_n10540_));
  INV_X1     g10348(.I(new_n10540_), .ZN(new_n10541_));
  INV_X1     g10349(.I(new_n10086_), .ZN(new_n10542_));
  INV_X1     g10350(.I(new_n10081_), .ZN(new_n10543_));
  INV_X1     g10351(.I(new_n10088_), .ZN(new_n10544_));
  NOR2_X1    g10352(.A1(new_n10544_), .A2(new_n10543_), .ZN(new_n10545_));
  NOR3_X1    g10353(.A1(new_n10545_), .A2(new_n10082_), .A3(new_n10542_), .ZN(new_n10546_));
  NOR3_X1    g10354(.A1(new_n10221_), .A2(new_n10082_), .A3(new_n10545_), .ZN(new_n10547_));
  INV_X1     g10355(.I(new_n10547_), .ZN(new_n10548_));
  AOI22_X1   g10356(.A1(new_n10548_), .A2(new_n10542_), .B1(\asqrt[24] ), .B2(new_n10546_), .ZN(new_n10549_));
  NOR3_X1    g10357(.A1(new_n10539_), .A2(new_n10530_), .A3(\asqrt[52] ), .ZN(new_n10550_));
  NOR2_X1    g10358(.A1(new_n10550_), .A2(new_n10549_), .ZN(new_n10551_));
  OAI21_X1   g10359(.A1(new_n10551_), .A2(new_n10541_), .B(\asqrt[53] ), .ZN(new_n10552_));
  NOR3_X1    g10360(.A1(new_n10221_), .A2(new_n10091_), .A3(new_n10132_), .ZN(new_n10553_));
  INV_X1     g10361(.I(new_n10553_), .ZN(new_n10554_));
  NOR3_X1    g10362(.A1(new_n10091_), .A2(new_n10236_), .A3(new_n10132_), .ZN(new_n10555_));
  AOI22_X1   g10363(.A1(new_n10554_), .A2(new_n10236_), .B1(\asqrt[24] ), .B2(new_n10555_), .ZN(new_n10556_));
  INV_X1     g10364(.I(new_n10556_), .ZN(new_n10557_));
  NAND2_X1   g10365(.A1(new_n10540_), .A2(new_n1103_), .ZN(new_n10558_));
  OAI21_X1   g10366(.A1(new_n10551_), .A2(new_n10558_), .B(new_n10557_), .ZN(new_n10559_));
  AOI21_X1   g10367(.A1(new_n10559_), .A2(new_n10552_), .B(new_n904_), .ZN(new_n10560_));
  INV_X1     g10368(.I(new_n10099_), .ZN(new_n10561_));
  NOR2_X1    g10369(.A1(new_n10106_), .A2(new_n10098_), .ZN(new_n10562_));
  NOR3_X1    g10370(.A1(new_n10561_), .A2(new_n10105_), .A3(new_n10562_), .ZN(new_n10563_));
  NOR3_X1    g10371(.A1(new_n10221_), .A2(new_n10561_), .A3(new_n10562_), .ZN(new_n10564_));
  INV_X1     g10372(.I(new_n10564_), .ZN(new_n10565_));
  AOI22_X1   g10373(.A1(new_n10565_), .A2(new_n10105_), .B1(\asqrt[24] ), .B2(new_n10563_), .ZN(new_n10566_));
  OAI21_X1   g10374(.A1(new_n10549_), .A2(new_n10550_), .B(new_n10540_), .ZN(new_n10567_));
  AOI21_X1   g10375(.A1(new_n10567_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n10568_));
  AOI21_X1   g10376(.A1(new_n10568_), .A2(new_n10559_), .B(new_n10566_), .ZN(new_n10569_));
  OAI21_X1   g10377(.A1(new_n10569_), .A2(new_n10560_), .B(\asqrt[55] ), .ZN(new_n10570_));
  INV_X1     g10378(.I(new_n10570_), .ZN(new_n10571_));
  NOR2_X1    g10379(.A1(new_n10116_), .A2(new_n10110_), .ZN(new_n10572_));
  NOR3_X1    g10380(.A1(new_n10221_), .A2(new_n10108_), .A3(new_n10572_), .ZN(new_n10573_));
  INV_X1     g10381(.I(new_n10573_), .ZN(new_n10574_));
  NOR3_X1    g10382(.A1(new_n10572_), .A2(new_n10108_), .A3(new_n10115_), .ZN(new_n10575_));
  AOI22_X1   g10383(.A1(new_n10574_), .A2(new_n10115_), .B1(\asqrt[24] ), .B2(new_n10575_), .ZN(new_n10576_));
  NOR3_X1    g10384(.A1(new_n10569_), .A2(new_n10560_), .A3(\asqrt[55] ), .ZN(new_n10577_));
  NOR2_X1    g10385(.A1(new_n10577_), .A2(new_n10576_), .ZN(new_n10578_));
  OAI21_X1   g10386(.A1(new_n10578_), .A2(new_n10571_), .B(\asqrt[56] ), .ZN(new_n10579_));
  NOR3_X1    g10387(.A1(new_n10118_), .A2(new_n10235_), .A3(new_n10163_), .ZN(new_n10580_));
  NOR3_X1    g10388(.A1(new_n10221_), .A2(new_n10118_), .A3(new_n10163_), .ZN(new_n10581_));
  INV_X1     g10389(.I(new_n10581_), .ZN(new_n10582_));
  AOI22_X1   g10390(.A1(new_n10582_), .A2(new_n10235_), .B1(\asqrt[24] ), .B2(new_n10580_), .ZN(new_n10583_));
  INV_X1     g10391(.I(new_n10583_), .ZN(new_n10584_));
  NAND2_X1   g10392(.A1(new_n10570_), .A2(new_n703_), .ZN(new_n10585_));
  OAI21_X1   g10393(.A1(new_n10578_), .A2(new_n10585_), .B(new_n10584_), .ZN(new_n10586_));
  AOI21_X1   g10394(.A1(new_n10586_), .A2(new_n10579_), .B(new_n531_), .ZN(new_n10587_));
  INV_X1     g10395(.I(new_n10125_), .ZN(new_n10588_));
  NOR2_X1    g10396(.A1(new_n10137_), .A2(new_n10124_), .ZN(new_n10589_));
  NOR3_X1    g10397(.A1(new_n10221_), .A2(new_n10588_), .A3(new_n10589_), .ZN(new_n10590_));
  INV_X1     g10398(.I(new_n10590_), .ZN(new_n10591_));
  NOR3_X1    g10399(.A1(new_n10588_), .A2(new_n10131_), .A3(new_n10589_), .ZN(new_n10592_));
  AOI22_X1   g10400(.A1(new_n10591_), .A2(new_n10131_), .B1(\asqrt[24] ), .B2(new_n10592_), .ZN(new_n10593_));
  OAI21_X1   g10401(.A1(new_n10576_), .A2(new_n10577_), .B(new_n10570_), .ZN(new_n10594_));
  AOI21_X1   g10402(.A1(new_n10594_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n10595_));
  AOI21_X1   g10403(.A1(new_n10595_), .A2(new_n10586_), .B(new_n10593_), .ZN(new_n10596_));
  OAI21_X1   g10404(.A1(new_n10596_), .A2(new_n10587_), .B(\asqrt[58] ), .ZN(new_n10597_));
  NOR2_X1    g10405(.A1(new_n10147_), .A2(new_n10141_), .ZN(new_n10598_));
  NOR3_X1    g10406(.A1(new_n10598_), .A2(new_n10139_), .A3(new_n10146_), .ZN(new_n10599_));
  NOR3_X1    g10407(.A1(new_n10221_), .A2(new_n10139_), .A3(new_n10598_), .ZN(new_n10600_));
  INV_X1     g10408(.I(new_n10600_), .ZN(new_n10601_));
  AOI22_X1   g10409(.A1(new_n10601_), .A2(new_n10146_), .B1(\asqrt[24] ), .B2(new_n10599_), .ZN(new_n10602_));
  INV_X1     g10410(.I(new_n10602_), .ZN(new_n10603_));
  INV_X1     g10411(.I(new_n10576_), .ZN(new_n10604_));
  INV_X1     g10412(.I(new_n10549_), .ZN(new_n10605_));
  INV_X1     g10413(.I(new_n10519_), .ZN(new_n10606_));
  INV_X1     g10414(.I(new_n10489_), .ZN(new_n10607_));
  INV_X1     g10415(.I(new_n10459_), .ZN(new_n10608_));
  INV_X1     g10416(.I(new_n10431_), .ZN(new_n10609_));
  INV_X1     g10417(.I(new_n10405_), .ZN(new_n10610_));
  INV_X1     g10418(.I(new_n10379_), .ZN(new_n10611_));
  INV_X1     g10419(.I(new_n10353_), .ZN(new_n10612_));
  NAND2_X1   g10420(.A1(new_n10293_), .A2(new_n8483_), .ZN(new_n10613_));
  OAI21_X1   g10421(.A1(new_n10613_), .A2(new_n10326_), .B(new_n10307_), .ZN(new_n10614_));
  AOI21_X1   g10422(.A1(new_n10614_), .A2(new_n10336_), .B(new_n8036_), .ZN(new_n10615_));
  NOR2_X1    g10423(.A1(new_n10301_), .A2(\asqrt[29] ), .ZN(new_n10616_));
  AOI21_X1   g10424(.A1(new_n10616_), .A2(new_n10614_), .B(new_n10334_), .ZN(new_n10617_));
  OAI21_X1   g10425(.A1(new_n10617_), .A2(new_n10615_), .B(\asqrt[30] ), .ZN(new_n10618_));
  NAND2_X1   g10426(.A1(new_n10618_), .A2(new_n7229_), .ZN(new_n10619_));
  OAI21_X1   g10427(.A1(new_n10619_), .A2(new_n10346_), .B(new_n10612_), .ZN(new_n10620_));
  NAND3_X1   g10428(.A1(new_n10620_), .A2(new_n6824_), .A3(new_n10347_), .ZN(new_n10621_));
  AOI22_X1   g10429(.A1(new_n10621_), .A2(new_n10362_), .B1(\asqrt[32] ), .B2(new_n10370_), .ZN(new_n10622_));
  OAI21_X1   g10430(.A1(new_n10622_), .A2(new_n6356_), .B(new_n6077_), .ZN(new_n10623_));
  OAI21_X1   g10431(.A1(new_n10623_), .A2(new_n10372_), .B(new_n10611_), .ZN(new_n10624_));
  AOI21_X1   g10432(.A1(new_n10624_), .A2(new_n10373_), .B(new_n5708_), .ZN(new_n10625_));
  AOI21_X1   g10433(.A1(new_n10620_), .A2(new_n10347_), .B(new_n6824_), .ZN(new_n10626_));
  NOR3_X1    g10434(.A1(new_n10617_), .A2(new_n10615_), .A3(\asqrt[30] ), .ZN(new_n10627_));
  OAI21_X1   g10435(.A1(new_n10343_), .A2(new_n10627_), .B(new_n10618_), .ZN(new_n10628_));
  AOI21_X1   g10436(.A1(new_n10628_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n10629_));
  AOI21_X1   g10437(.A1(new_n10629_), .A2(new_n10620_), .B(new_n10361_), .ZN(new_n10630_));
  NOR3_X1    g10438(.A1(new_n10630_), .A2(\asqrt[33] ), .A3(new_n10626_), .ZN(new_n10631_));
  OAI22_X1   g10439(.A1(new_n10631_), .A2(new_n10369_), .B1(new_n10622_), .B2(new_n6356_), .ZN(new_n10632_));
  AOI21_X1   g10440(.A1(new_n10632_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n10633_));
  AOI21_X1   g10441(.A1(new_n10633_), .A2(new_n10624_), .B(new_n10387_), .ZN(new_n10634_));
  OAI21_X1   g10442(.A1(new_n10634_), .A2(new_n10625_), .B(\asqrt[36] ), .ZN(new_n10635_));
  NAND2_X1   g10443(.A1(new_n10635_), .A2(new_n5024_), .ZN(new_n10636_));
  OAI21_X1   g10444(.A1(new_n10636_), .A2(new_n10398_), .B(new_n10610_), .ZN(new_n10637_));
  AOI21_X1   g10445(.A1(new_n10637_), .A2(new_n10399_), .B(new_n4696_), .ZN(new_n10638_));
  NOR3_X1    g10446(.A1(new_n10634_), .A2(\asqrt[36] ), .A3(new_n10625_), .ZN(new_n10639_));
  OAI21_X1   g10447(.A1(new_n10395_), .A2(new_n10639_), .B(new_n10635_), .ZN(new_n10640_));
  AOI21_X1   g10448(.A1(new_n10640_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n10641_));
  AOI21_X1   g10449(.A1(new_n10641_), .A2(new_n10637_), .B(new_n10413_), .ZN(new_n10642_));
  OAI21_X1   g10450(.A1(new_n10642_), .A2(new_n10638_), .B(\asqrt[39] ), .ZN(new_n10643_));
  NAND2_X1   g10451(.A1(new_n10643_), .A2(new_n4071_), .ZN(new_n10644_));
  OAI21_X1   g10452(.A1(new_n10644_), .A2(new_n10424_), .B(new_n10609_), .ZN(new_n10645_));
  AOI21_X1   g10453(.A1(new_n10645_), .A2(new_n10425_), .B(new_n3782_), .ZN(new_n10646_));
  NOR3_X1    g10454(.A1(new_n10642_), .A2(\asqrt[39] ), .A3(new_n10638_), .ZN(new_n10647_));
  OAI21_X1   g10455(.A1(new_n10421_), .A2(new_n10647_), .B(new_n10643_), .ZN(new_n10648_));
  AOI21_X1   g10456(.A1(new_n10648_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n10649_));
  AOI21_X1   g10457(.A1(new_n10649_), .A2(new_n10645_), .B(new_n10439_), .ZN(new_n10650_));
  OAI21_X1   g10458(.A1(new_n10650_), .A2(new_n10646_), .B(\asqrt[42] ), .ZN(new_n10651_));
  NAND2_X1   g10459(.A1(new_n10651_), .A2(new_n3218_), .ZN(new_n10652_));
  OAI21_X1   g10460(.A1(new_n10652_), .A2(new_n10450_), .B(new_n10608_), .ZN(new_n10653_));
  AOI21_X1   g10461(.A1(new_n10653_), .A2(new_n10451_), .B(new_n2954_), .ZN(new_n10654_));
  NOR3_X1    g10462(.A1(new_n10650_), .A2(\asqrt[42] ), .A3(new_n10646_), .ZN(new_n10655_));
  OAI21_X1   g10463(.A1(new_n10447_), .A2(new_n10655_), .B(new_n10651_), .ZN(new_n10656_));
  AOI21_X1   g10464(.A1(new_n10656_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n10657_));
  AOI21_X1   g10465(.A1(new_n10657_), .A2(new_n10653_), .B(new_n10466_), .ZN(new_n10658_));
  OAI21_X1   g10466(.A1(new_n10658_), .A2(new_n10654_), .B(\asqrt[45] ), .ZN(new_n10659_));
  NAND2_X1   g10467(.A1(new_n10659_), .A2(new_n2465_), .ZN(new_n10660_));
  OAI21_X1   g10468(.A1(new_n10660_), .A2(new_n10479_), .B(new_n10607_), .ZN(new_n10661_));
  AOI21_X1   g10469(.A1(new_n10661_), .A2(new_n10480_), .B(new_n2229_), .ZN(new_n10662_));
  NOR3_X1    g10470(.A1(new_n10658_), .A2(\asqrt[45] ), .A3(new_n10654_), .ZN(new_n10663_));
  OAI21_X1   g10471(.A1(new_n10476_), .A2(new_n10663_), .B(new_n10659_), .ZN(new_n10664_));
  AOI21_X1   g10472(.A1(new_n10664_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n10665_));
  AOI21_X1   g10473(.A1(new_n10665_), .A2(new_n10661_), .B(new_n10496_), .ZN(new_n10666_));
  OAI21_X1   g10474(.A1(new_n10666_), .A2(new_n10662_), .B(\asqrt[48] ), .ZN(new_n10667_));
  NAND2_X1   g10475(.A1(new_n10667_), .A2(new_n1806_), .ZN(new_n10668_));
  OAI21_X1   g10476(.A1(new_n10668_), .A2(new_n10509_), .B(new_n10606_), .ZN(new_n10669_));
  AOI21_X1   g10477(.A1(new_n10669_), .A2(new_n10510_), .B(new_n1612_), .ZN(new_n10670_));
  NOR3_X1    g10478(.A1(new_n10666_), .A2(\asqrt[48] ), .A3(new_n10662_), .ZN(new_n10671_));
  OAI21_X1   g10479(.A1(new_n10506_), .A2(new_n10671_), .B(new_n10667_), .ZN(new_n10672_));
  AOI21_X1   g10480(.A1(new_n10672_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n10673_));
  AOI21_X1   g10481(.A1(new_n10673_), .A2(new_n10669_), .B(new_n10526_), .ZN(new_n10674_));
  OAI21_X1   g10482(.A1(new_n10674_), .A2(new_n10670_), .B(\asqrt[51] ), .ZN(new_n10675_));
  NAND2_X1   g10483(.A1(new_n10675_), .A2(new_n1256_), .ZN(new_n10676_));
  OAI21_X1   g10484(.A1(new_n10676_), .A2(new_n10539_), .B(new_n10605_), .ZN(new_n10677_));
  NAND3_X1   g10485(.A1(new_n10677_), .A2(new_n1103_), .A3(new_n10540_), .ZN(new_n10678_));
  AOI22_X1   g10486(.A1(new_n10678_), .A2(new_n10557_), .B1(\asqrt[53] ), .B2(new_n10567_), .ZN(new_n10679_));
  OAI21_X1   g10487(.A1(new_n10679_), .A2(new_n904_), .B(new_n823_), .ZN(new_n10680_));
  OAI21_X1   g10488(.A1(new_n10680_), .A2(new_n10569_), .B(new_n10604_), .ZN(new_n10681_));
  NAND3_X1   g10489(.A1(new_n10681_), .A2(new_n703_), .A3(new_n10570_), .ZN(new_n10682_));
  AOI22_X1   g10490(.A1(new_n10682_), .A2(new_n10584_), .B1(\asqrt[56] ), .B2(new_n10594_), .ZN(new_n10683_));
  OAI21_X1   g10491(.A1(new_n10683_), .A2(new_n531_), .B(new_n436_), .ZN(new_n10684_));
  OAI21_X1   g10492(.A1(new_n10684_), .A2(new_n10596_), .B(new_n10603_), .ZN(new_n10685_));
  AOI21_X1   g10493(.A1(new_n10685_), .A2(new_n10597_), .B(new_n327_), .ZN(new_n10686_));
  NOR3_X1    g10494(.A1(new_n10221_), .A2(new_n10149_), .A3(new_n10194_), .ZN(new_n10687_));
  INV_X1     g10495(.I(new_n10687_), .ZN(new_n10688_));
  NOR3_X1    g10496(.A1(new_n10149_), .A2(new_n10234_), .A3(new_n10194_), .ZN(new_n10689_));
  AOI22_X1   g10497(.A1(new_n10688_), .A2(new_n10234_), .B1(\asqrt[24] ), .B2(new_n10689_), .ZN(new_n10690_));
  NAND2_X1   g10498(.A1(new_n10597_), .A2(new_n327_), .ZN(new_n10691_));
  INV_X1     g10499(.I(new_n10691_), .ZN(new_n10692_));
  AOI21_X1   g10500(.A1(new_n10692_), .A2(new_n10685_), .B(new_n10690_), .ZN(new_n10693_));
  OAI21_X1   g10501(.A1(new_n10693_), .A2(new_n10686_), .B(\asqrt[60] ), .ZN(new_n10694_));
  INV_X1     g10502(.I(new_n10156_), .ZN(new_n10695_));
  NOR2_X1    g10503(.A1(new_n10168_), .A2(new_n10155_), .ZN(new_n10696_));
  NOR3_X1    g10504(.A1(new_n10695_), .A2(new_n10162_), .A3(new_n10696_), .ZN(new_n10697_));
  NOR3_X1    g10505(.A1(new_n10221_), .A2(new_n10695_), .A3(new_n10696_), .ZN(new_n10698_));
  INV_X1     g10506(.I(new_n10698_), .ZN(new_n10699_));
  AOI22_X1   g10507(.A1(new_n10699_), .A2(new_n10162_), .B1(\asqrt[24] ), .B2(new_n10697_), .ZN(new_n10700_));
  INV_X1     g10508(.I(new_n10700_), .ZN(new_n10701_));
  INV_X1     g10509(.I(new_n10597_), .ZN(new_n10702_));
  NOR3_X1    g10510(.A1(new_n10596_), .A2(new_n10587_), .A3(\asqrt[58] ), .ZN(new_n10703_));
  NOR2_X1    g10511(.A1(new_n10703_), .A2(new_n10602_), .ZN(new_n10704_));
  OAI21_X1   g10512(.A1(new_n10704_), .A2(new_n10702_), .B(\asqrt[59] ), .ZN(new_n10705_));
  NAND2_X1   g10513(.A1(new_n10705_), .A2(new_n306_), .ZN(new_n10706_));
  OAI21_X1   g10514(.A1(new_n10706_), .A2(new_n10693_), .B(new_n10701_), .ZN(new_n10707_));
  AOI21_X1   g10515(.A1(new_n10707_), .A2(new_n10694_), .B(new_n218_), .ZN(new_n10708_));
  NOR2_X1    g10516(.A1(new_n10172_), .A2(new_n10178_), .ZN(new_n10709_));
  NOR3_X1    g10517(.A1(new_n10221_), .A2(new_n10170_), .A3(new_n10709_), .ZN(new_n10710_));
  INV_X1     g10518(.I(new_n10710_), .ZN(new_n10711_));
  NOR3_X1    g10519(.A1(new_n10709_), .A2(new_n10170_), .A3(new_n10177_), .ZN(new_n10712_));
  AOI22_X1   g10520(.A1(new_n10711_), .A2(new_n10177_), .B1(\asqrt[24] ), .B2(new_n10712_), .ZN(new_n10713_));
  INV_X1     g10521(.I(new_n10690_), .ZN(new_n10714_));
  OAI21_X1   g10522(.A1(new_n10704_), .A2(new_n10691_), .B(new_n10714_), .ZN(new_n10715_));
  AOI21_X1   g10523(.A1(new_n10715_), .A2(new_n10705_), .B(new_n306_), .ZN(new_n10716_));
  NOR2_X1    g10524(.A1(new_n10716_), .A2(\asqrt[61] ), .ZN(new_n10717_));
  AOI21_X1   g10525(.A1(new_n10717_), .A2(new_n10707_), .B(new_n10713_), .ZN(new_n10718_));
  OAI21_X1   g10526(.A1(new_n10718_), .A2(new_n10708_), .B(\asqrt[62] ), .ZN(new_n10719_));
  NOR3_X1    g10527(.A1(new_n10180_), .A2(new_n10233_), .A3(new_n10231_), .ZN(new_n10720_));
  NOR3_X1    g10528(.A1(new_n10221_), .A2(new_n10180_), .A3(new_n10231_), .ZN(new_n10721_));
  INV_X1     g10529(.I(new_n10721_), .ZN(new_n10722_));
  AOI22_X1   g10530(.A1(new_n10722_), .A2(new_n10233_), .B1(\asqrt[24] ), .B2(new_n10720_), .ZN(new_n10723_));
  INV_X1     g10531(.I(new_n10723_), .ZN(new_n10724_));
  OAI21_X1   g10532(.A1(new_n10602_), .A2(new_n10703_), .B(new_n10597_), .ZN(new_n10725_));
  AOI21_X1   g10533(.A1(new_n10725_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n10726_));
  AOI21_X1   g10534(.A1(new_n10726_), .A2(new_n10715_), .B(new_n10700_), .ZN(new_n10727_));
  OAI21_X1   g10535(.A1(new_n10727_), .A2(new_n10716_), .B(\asqrt[61] ), .ZN(new_n10728_));
  NAND2_X1   g10536(.A1(new_n10728_), .A2(new_n207_), .ZN(new_n10729_));
  OAI21_X1   g10537(.A1(new_n10729_), .A2(new_n10718_), .B(new_n10724_), .ZN(new_n10730_));
  NAND4_X1   g10538(.A1(\asqrt[24] ), .A2(new_n10187_), .A3(new_n10192_), .A4(new_n10270_), .ZN(new_n10731_));
  NAND2_X1   g10539(.A1(new_n10187_), .A2(new_n10270_), .ZN(new_n10732_));
  OAI21_X1   g10540(.A1(new_n10221_), .A2(new_n10732_), .B(new_n10193_), .ZN(new_n10733_));
  NAND2_X1   g10541(.A1(new_n10731_), .A2(new_n10733_), .ZN(new_n10734_));
  NOR2_X1    g10542(.A1(new_n10271_), .A2(new_n10211_), .ZN(new_n10735_));
  NAND2_X1   g10543(.A1(\asqrt[24] ), .A2(new_n10735_), .ZN(new_n10736_));
  NAND3_X1   g10544(.A1(new_n10734_), .A2(new_n10282_), .A3(new_n10736_), .ZN(new_n10737_));
  AOI21_X1   g10545(.A1(new_n10730_), .A2(new_n10719_), .B(new_n10737_), .ZN(new_n10738_));
  NOR3_X1    g10546(.A1(new_n10727_), .A2(new_n10716_), .A3(\asqrt[61] ), .ZN(new_n10739_));
  OAI21_X1   g10547(.A1(new_n10713_), .A2(new_n10739_), .B(new_n10728_), .ZN(new_n10740_));
  AOI21_X1   g10548(.A1(new_n10740_), .A2(\asqrt[62] ), .B(new_n10734_), .ZN(new_n10741_));
  OAI21_X1   g10549(.A1(new_n10221_), .A2(new_n10211_), .B(new_n10271_), .ZN(new_n10742_));
  NOR2_X1    g10550(.A1(new_n10735_), .A2(new_n193_), .ZN(new_n10743_));
  NAND2_X1   g10551(.A1(new_n10742_), .A2(new_n10743_), .ZN(new_n10744_));
  INV_X1     g10552(.I(new_n10744_), .ZN(new_n10745_));
  AND3_X2    g10553(.A1(new_n10203_), .A2(new_n10201_), .A3(new_n10217_), .Z(new_n10746_));
  NAND4_X1   g10554(.A1(new_n10272_), .A2(new_n10282_), .A3(new_n10214_), .A4(new_n10746_), .ZN(new_n10747_));
  INV_X1     g10555(.I(new_n10747_), .ZN(new_n10748_));
  NOR2_X1    g10556(.A1(new_n10745_), .A2(new_n10748_), .ZN(new_n10749_));
  INV_X1     g10557(.I(new_n10749_), .ZN(new_n10750_));
  AOI21_X1   g10558(.A1(new_n10741_), .A2(new_n10730_), .B(new_n10750_), .ZN(new_n10751_));
  OAI21_X1   g10559(.A1(\asqrt[63] ), .A2(new_n10738_), .B(new_n10751_), .ZN(\asqrt[23] ));
  NOR2_X1    g10560(.A1(\a[44] ), .A2(\a[45] ), .ZN(new_n10753_));
  INV_X1     g10561(.I(new_n10753_), .ZN(new_n10754_));
  NOR2_X1    g10562(.A1(new_n10754_), .A2(\a[46] ), .ZN(new_n10755_));
  INV_X1     g10563(.I(new_n10755_), .ZN(new_n10756_));
  NAND2_X1   g10564(.A1(new_n10730_), .A2(new_n10719_), .ZN(new_n10757_));
  INV_X1     g10565(.I(new_n10737_), .ZN(new_n10758_));
  AOI21_X1   g10566(.A1(new_n10757_), .A2(new_n10758_), .B(\asqrt[63] ), .ZN(new_n10759_));
  INV_X1     g10567(.I(new_n10713_), .ZN(new_n10760_));
  NAND3_X1   g10568(.A1(new_n10685_), .A2(new_n327_), .A3(new_n10597_), .ZN(new_n10761_));
  AOI22_X1   g10569(.A1(new_n10761_), .A2(new_n10714_), .B1(new_n10725_), .B2(\asqrt[59] ), .ZN(new_n10762_));
  OAI21_X1   g10570(.A1(new_n10762_), .A2(new_n306_), .B(new_n218_), .ZN(new_n10763_));
  OAI21_X1   g10571(.A1(new_n10763_), .A2(new_n10727_), .B(new_n10760_), .ZN(new_n10764_));
  NOR2_X1    g10572(.A1(new_n10708_), .A2(\asqrt[62] ), .ZN(new_n10765_));
  AOI21_X1   g10573(.A1(new_n10765_), .A2(new_n10764_), .B(new_n10723_), .ZN(new_n10766_));
  INV_X1     g10574(.I(new_n10734_), .ZN(new_n10767_));
  NAND2_X1   g10575(.A1(new_n10719_), .A2(new_n10767_), .ZN(new_n10768_));
  OAI21_X1   g10576(.A1(new_n10768_), .A2(new_n10766_), .B(new_n10749_), .ZN(new_n10769_));
  OAI21_X1   g10577(.A1(new_n10759_), .A2(new_n10769_), .B(\a[46] ), .ZN(new_n10770_));
  AOI21_X1   g10578(.A1(new_n10770_), .A2(new_n10756_), .B(new_n10221_), .ZN(new_n10771_));
  INV_X1     g10579(.I(\a[46] ), .ZN(new_n10772_));
  NAND3_X1   g10580(.A1(new_n10764_), .A2(new_n207_), .A3(new_n10728_), .ZN(new_n10773_));
  AOI22_X1   g10581(.A1(new_n10773_), .A2(new_n10724_), .B1(new_n10740_), .B2(\asqrt[62] ), .ZN(new_n10774_));
  OAI21_X1   g10582(.A1(new_n10774_), .A2(new_n10737_), .B(new_n193_), .ZN(new_n10775_));
  AOI21_X1   g10583(.A1(new_n10775_), .A2(new_n10751_), .B(new_n10772_), .ZN(new_n10776_));
  NAND4_X1   g10584(.A1(new_n10282_), .A2(new_n10214_), .A3(new_n10217_), .A4(new_n10756_), .ZN(new_n10777_));
  NOR2_X1    g10585(.A1(new_n10777_), .A2(new_n10209_), .ZN(new_n10778_));
  INV_X1     g10586(.I(new_n10778_), .ZN(new_n10779_));
  NOR2_X1    g10587(.A1(new_n10776_), .A2(new_n10779_), .ZN(new_n10780_));
  AOI21_X1   g10588(.A1(new_n10775_), .A2(new_n10751_), .B(new_n10224_), .ZN(new_n10781_));
  INV_X1     g10589(.I(\a[47] ), .ZN(new_n10782_));
  AOI21_X1   g10590(.A1(\asqrt[23] ), .A2(new_n10772_), .B(new_n10782_), .ZN(new_n10783_));
  NOR3_X1    g10591(.A1(new_n10780_), .A2(new_n10783_), .A3(new_n10781_), .ZN(new_n10784_));
  OAI21_X1   g10592(.A1(new_n10784_), .A2(new_n10771_), .B(\asqrt[25] ), .ZN(new_n10785_));
  OAI21_X1   g10593(.A1(new_n10759_), .A2(new_n10769_), .B(new_n10223_), .ZN(new_n10786_));
  NAND2_X1   g10594(.A1(new_n10741_), .A2(new_n10730_), .ZN(new_n10787_));
  NOR3_X1    g10595(.A1(new_n10745_), .A2(new_n10221_), .A3(new_n10748_), .ZN(new_n10788_));
  NAND3_X1   g10596(.A1(new_n10775_), .A2(new_n10787_), .A3(new_n10788_), .ZN(new_n10789_));
  AOI21_X1   g10597(.A1(new_n10789_), .A2(new_n10786_), .B(new_n10222_), .ZN(new_n10790_));
  NAND2_X1   g10598(.A1(new_n10787_), .A2(new_n10788_), .ZN(new_n10791_));
  NOR2_X1    g10599(.A1(new_n10791_), .A2(new_n10759_), .ZN(new_n10792_));
  NOR3_X1    g10600(.A1(new_n10792_), .A2(new_n10781_), .A3(\a[48] ), .ZN(new_n10793_));
  AOI21_X1   g10601(.A1(\asqrt[23] ), .A2(\a[46] ), .B(new_n10755_), .ZN(new_n10794_));
  OAI21_X1   g10602(.A1(new_n10794_), .A2(new_n10221_), .B(new_n9846_), .ZN(new_n10795_));
  OAI22_X1   g10603(.A1(new_n10784_), .A2(new_n10795_), .B1(new_n10790_), .B2(new_n10793_), .ZN(new_n10796_));
  AOI21_X1   g10604(.A1(new_n10796_), .A2(new_n10785_), .B(new_n9317_), .ZN(new_n10797_));
  NOR3_X1    g10605(.A1(new_n10311_), .A2(new_n10313_), .A3(new_n10277_), .ZN(new_n10798_));
  NAND3_X1   g10606(.A1(\asqrt[23] ), .A2(new_n10310_), .A3(new_n10230_), .ZN(new_n10799_));
  AOI22_X1   g10607(.A1(new_n10799_), .A2(new_n10277_), .B1(\asqrt[23] ), .B2(new_n10798_), .ZN(new_n10800_));
  OAI21_X1   g10608(.A1(new_n10776_), .A2(new_n10755_), .B(\asqrt[24] ), .ZN(new_n10801_));
  AOI21_X1   g10609(.A1(new_n10775_), .A2(new_n10751_), .B(\a[46] ), .ZN(new_n10802_));
  OAI21_X1   g10610(.A1(new_n10782_), .A2(new_n10802_), .B(new_n10786_), .ZN(new_n10803_));
  OAI21_X1   g10611(.A1(new_n10803_), .A2(new_n10780_), .B(new_n10801_), .ZN(new_n10804_));
  AOI21_X1   g10612(.A1(new_n10804_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n10805_));
  AOI21_X1   g10613(.A1(new_n10805_), .A2(new_n10796_), .B(new_n10800_), .ZN(new_n10806_));
  OAI21_X1   g10614(.A1(new_n10806_), .A2(new_n10797_), .B(\asqrt[27] ), .ZN(new_n10807_));
  INV_X1     g10615(.I(new_n10807_), .ZN(new_n10808_));
  NOR2_X1    g10616(.A1(new_n10316_), .A2(new_n10319_), .ZN(new_n10809_));
  INV_X1     g10617(.I(new_n10809_), .ZN(new_n10810_));
  NAND4_X1   g10618(.A1(\asqrt[23] ), .A2(new_n10317_), .A3(new_n10290_), .A4(new_n10810_), .ZN(new_n10811_));
  INV_X1     g10619(.I(\asqrt[23] ), .ZN(new_n10812_));
  NOR3_X1    g10620(.A1(new_n10812_), .A2(new_n10279_), .A3(new_n10809_), .ZN(new_n10813_));
  OAI21_X1   g10621(.A1(new_n10813_), .A2(new_n10290_), .B(new_n10811_), .ZN(new_n10814_));
  INV_X1     g10622(.I(new_n10814_), .ZN(new_n10815_));
  NOR3_X1    g10623(.A1(new_n10806_), .A2(new_n10797_), .A3(\asqrt[27] ), .ZN(new_n10816_));
  NOR2_X1    g10624(.A1(new_n10816_), .A2(new_n10815_), .ZN(new_n10817_));
  OAI21_X1   g10625(.A1(new_n10817_), .A2(new_n10808_), .B(\asqrt[28] ), .ZN(new_n10818_));
  NAND2_X1   g10626(.A1(new_n10325_), .A2(new_n10320_), .ZN(new_n10819_));
  NAND3_X1   g10627(.A1(\asqrt[23] ), .A2(new_n10293_), .A3(new_n10819_), .ZN(new_n10820_));
  AND3_X2    g10628(.A1(new_n10293_), .A2(new_n10297_), .A3(new_n10819_), .Z(new_n10821_));
  AOI22_X1   g10629(.A1(new_n10820_), .A2(new_n10298_), .B1(\asqrt[23] ), .B2(new_n10821_), .ZN(new_n10822_));
  INV_X1     g10630(.I(new_n10822_), .ZN(new_n10823_));
  NAND2_X1   g10631(.A1(new_n10807_), .A2(new_n8483_), .ZN(new_n10824_));
  OAI21_X1   g10632(.A1(new_n10817_), .A2(new_n10824_), .B(new_n10823_), .ZN(new_n10825_));
  AOI21_X1   g10633(.A1(new_n10825_), .A2(new_n10818_), .B(new_n8036_), .ZN(new_n10826_));
  NOR3_X1    g10634(.A1(new_n10301_), .A2(new_n10307_), .A3(new_n10327_), .ZN(new_n10827_));
  NOR3_X1    g10635(.A1(new_n10812_), .A2(new_n10301_), .A3(new_n10327_), .ZN(new_n10828_));
  INV_X1     g10636(.I(new_n10828_), .ZN(new_n10829_));
  AOI22_X1   g10637(.A1(new_n10829_), .A2(new_n10307_), .B1(\asqrt[23] ), .B2(new_n10827_), .ZN(new_n10830_));
  OAI21_X1   g10638(.A1(new_n10815_), .A2(new_n10816_), .B(new_n10807_), .ZN(new_n10831_));
  AOI21_X1   g10639(.A1(new_n10831_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n10832_));
  AOI21_X1   g10640(.A1(new_n10832_), .A2(new_n10825_), .B(new_n10830_), .ZN(new_n10833_));
  OAI21_X1   g10641(.A1(new_n10833_), .A2(new_n10826_), .B(\asqrt[30] ), .ZN(new_n10834_));
  INV_X1     g10642(.I(new_n10834_), .ZN(new_n10835_));
  NAND2_X1   g10643(.A1(new_n10616_), .A2(new_n10614_), .ZN(new_n10836_));
  NAND3_X1   g10644(.A1(\asqrt[23] ), .A2(new_n10329_), .A3(new_n10836_), .ZN(new_n10837_));
  AND3_X2    g10645(.A1(new_n10836_), .A2(new_n10329_), .A3(new_n10334_), .Z(new_n10838_));
  AOI22_X1   g10646(.A1(new_n10837_), .A2(new_n10335_), .B1(\asqrt[23] ), .B2(new_n10838_), .ZN(new_n10839_));
  NOR3_X1    g10647(.A1(new_n10833_), .A2(new_n10826_), .A3(\asqrt[30] ), .ZN(new_n10840_));
  NOR2_X1    g10648(.A1(new_n10840_), .A2(new_n10839_), .ZN(new_n10841_));
  OAI21_X1   g10649(.A1(new_n10841_), .A2(new_n10835_), .B(\asqrt[31] ), .ZN(new_n10842_));
  INV_X1     g10650(.I(new_n10343_), .ZN(new_n10843_));
  NOR3_X1    g10651(.A1(new_n10627_), .A2(new_n10339_), .A3(new_n10843_), .ZN(new_n10844_));
  NOR3_X1    g10652(.A1(new_n10812_), .A2(new_n10339_), .A3(new_n10627_), .ZN(new_n10845_));
  INV_X1     g10653(.I(new_n10845_), .ZN(new_n10846_));
  AOI22_X1   g10654(.A1(new_n10846_), .A2(new_n10843_), .B1(\asqrt[23] ), .B2(new_n10844_), .ZN(new_n10847_));
  INV_X1     g10655(.I(new_n10847_), .ZN(new_n10848_));
  NAND2_X1   g10656(.A1(new_n10834_), .A2(new_n7229_), .ZN(new_n10849_));
  OAI21_X1   g10657(.A1(new_n10841_), .A2(new_n10849_), .B(new_n10848_), .ZN(new_n10850_));
  AOI21_X1   g10658(.A1(new_n10850_), .A2(new_n10842_), .B(new_n6824_), .ZN(new_n10851_));
  NOR3_X1    g10659(.A1(new_n10812_), .A2(new_n10348_), .A3(new_n10354_), .ZN(new_n10852_));
  INV_X1     g10660(.I(new_n10852_), .ZN(new_n10853_));
  NOR3_X1    g10661(.A1(new_n10348_), .A2(new_n10612_), .A3(new_n10354_), .ZN(new_n10854_));
  AOI22_X1   g10662(.A1(new_n10853_), .A2(new_n10612_), .B1(\asqrt[23] ), .B2(new_n10854_), .ZN(new_n10855_));
  OAI21_X1   g10663(.A1(new_n10839_), .A2(new_n10840_), .B(new_n10834_), .ZN(new_n10856_));
  AOI21_X1   g10664(.A1(new_n10856_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n10857_));
  AOI21_X1   g10665(.A1(new_n10857_), .A2(new_n10850_), .B(new_n10855_), .ZN(new_n10858_));
  OAI21_X1   g10666(.A1(new_n10858_), .A2(new_n10851_), .B(\asqrt[33] ), .ZN(new_n10859_));
  INV_X1     g10667(.I(new_n10859_), .ZN(new_n10860_));
  INV_X1     g10668(.I(new_n10621_), .ZN(new_n10861_));
  NOR3_X1    g10669(.A1(new_n10861_), .A2(new_n10626_), .A3(new_n10362_), .ZN(new_n10862_));
  NOR3_X1    g10670(.A1(new_n10812_), .A2(new_n10626_), .A3(new_n10861_), .ZN(new_n10863_));
  INV_X1     g10671(.I(new_n10863_), .ZN(new_n10864_));
  AOI22_X1   g10672(.A1(new_n10864_), .A2(new_n10362_), .B1(\asqrt[23] ), .B2(new_n10862_), .ZN(new_n10865_));
  NOR3_X1    g10673(.A1(new_n10858_), .A2(new_n10851_), .A3(\asqrt[33] ), .ZN(new_n10866_));
  NOR2_X1    g10674(.A1(new_n10866_), .A2(new_n10865_), .ZN(new_n10867_));
  OAI21_X1   g10675(.A1(new_n10867_), .A2(new_n10860_), .B(\asqrt[34] ), .ZN(new_n10868_));
  INV_X1     g10676(.I(new_n10369_), .ZN(new_n10869_));
  NOR3_X1    g10677(.A1(new_n10812_), .A2(new_n10365_), .A3(new_n10631_), .ZN(new_n10870_));
  INV_X1     g10678(.I(new_n10870_), .ZN(new_n10871_));
  NOR3_X1    g10679(.A1(new_n10631_), .A2(new_n10365_), .A3(new_n10869_), .ZN(new_n10872_));
  AOI22_X1   g10680(.A1(new_n10871_), .A2(new_n10869_), .B1(\asqrt[23] ), .B2(new_n10872_), .ZN(new_n10873_));
  INV_X1     g10681(.I(new_n10873_), .ZN(new_n10874_));
  NAND2_X1   g10682(.A1(new_n10859_), .A2(new_n6077_), .ZN(new_n10875_));
  OAI21_X1   g10683(.A1(new_n10867_), .A2(new_n10875_), .B(new_n10874_), .ZN(new_n10876_));
  AOI21_X1   g10684(.A1(new_n10876_), .A2(new_n10868_), .B(new_n5708_), .ZN(new_n10877_));
  NOR3_X1    g10685(.A1(new_n10374_), .A2(new_n10611_), .A3(new_n10380_), .ZN(new_n10878_));
  NOR3_X1    g10686(.A1(new_n10812_), .A2(new_n10374_), .A3(new_n10380_), .ZN(new_n10879_));
  INV_X1     g10687(.I(new_n10879_), .ZN(new_n10880_));
  AOI22_X1   g10688(.A1(new_n10880_), .A2(new_n10611_), .B1(\asqrt[23] ), .B2(new_n10878_), .ZN(new_n10881_));
  OAI21_X1   g10689(.A1(new_n10865_), .A2(new_n10866_), .B(new_n10859_), .ZN(new_n10882_));
  AOI21_X1   g10690(.A1(new_n10882_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n10883_));
  AOI21_X1   g10691(.A1(new_n10883_), .A2(new_n10876_), .B(new_n10881_), .ZN(new_n10884_));
  OAI21_X1   g10692(.A1(new_n10884_), .A2(new_n10877_), .B(\asqrt[36] ), .ZN(new_n10885_));
  INV_X1     g10693(.I(new_n10885_), .ZN(new_n10886_));
  NOR2_X1    g10694(.A1(new_n10381_), .A2(new_n10389_), .ZN(new_n10887_));
  NOR3_X1    g10695(.A1(new_n10812_), .A2(new_n10625_), .A3(new_n10887_), .ZN(new_n10888_));
  INV_X1     g10696(.I(new_n10888_), .ZN(new_n10889_));
  NOR3_X1    g10697(.A1(new_n10887_), .A2(new_n10625_), .A3(new_n10388_), .ZN(new_n10890_));
  AOI22_X1   g10698(.A1(new_n10889_), .A2(new_n10388_), .B1(\asqrt[23] ), .B2(new_n10890_), .ZN(new_n10891_));
  NOR3_X1    g10699(.A1(new_n10884_), .A2(new_n10877_), .A3(\asqrt[36] ), .ZN(new_n10892_));
  NOR2_X1    g10700(.A1(new_n10892_), .A2(new_n10891_), .ZN(new_n10893_));
  OAI21_X1   g10701(.A1(new_n10893_), .A2(new_n10886_), .B(\asqrt[37] ), .ZN(new_n10894_));
  INV_X1     g10702(.I(new_n10395_), .ZN(new_n10895_));
  NOR3_X1    g10703(.A1(new_n10639_), .A2(new_n10391_), .A3(new_n10895_), .ZN(new_n10896_));
  NOR3_X1    g10704(.A1(new_n10812_), .A2(new_n10391_), .A3(new_n10639_), .ZN(new_n10897_));
  INV_X1     g10705(.I(new_n10897_), .ZN(new_n10898_));
  AOI22_X1   g10706(.A1(new_n10898_), .A2(new_n10895_), .B1(\asqrt[23] ), .B2(new_n10896_), .ZN(new_n10899_));
  INV_X1     g10707(.I(new_n10899_), .ZN(new_n10900_));
  NAND2_X1   g10708(.A1(new_n10885_), .A2(new_n5024_), .ZN(new_n10901_));
  OAI21_X1   g10709(.A1(new_n10893_), .A2(new_n10901_), .B(new_n10900_), .ZN(new_n10902_));
  AOI21_X1   g10710(.A1(new_n10902_), .A2(new_n10894_), .B(new_n4696_), .ZN(new_n10903_));
  NOR3_X1    g10711(.A1(new_n10812_), .A2(new_n10400_), .A3(new_n10406_), .ZN(new_n10904_));
  INV_X1     g10712(.I(new_n10904_), .ZN(new_n10905_));
  NOR3_X1    g10713(.A1(new_n10400_), .A2(new_n10610_), .A3(new_n10406_), .ZN(new_n10906_));
  AOI22_X1   g10714(.A1(new_n10905_), .A2(new_n10610_), .B1(\asqrt[23] ), .B2(new_n10906_), .ZN(new_n10907_));
  OAI21_X1   g10715(.A1(new_n10891_), .A2(new_n10892_), .B(new_n10885_), .ZN(new_n10908_));
  AOI21_X1   g10716(.A1(new_n10908_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n10909_));
  AOI21_X1   g10717(.A1(new_n10909_), .A2(new_n10902_), .B(new_n10907_), .ZN(new_n10910_));
  OAI21_X1   g10718(.A1(new_n10910_), .A2(new_n10903_), .B(\asqrt[39] ), .ZN(new_n10911_));
  INV_X1     g10719(.I(new_n10911_), .ZN(new_n10912_));
  NOR2_X1    g10720(.A1(new_n10407_), .A2(new_n10415_), .ZN(new_n10913_));
  NOR3_X1    g10721(.A1(new_n10913_), .A2(new_n10638_), .A3(new_n10414_), .ZN(new_n10914_));
  NOR3_X1    g10722(.A1(new_n10812_), .A2(new_n10638_), .A3(new_n10913_), .ZN(new_n10915_));
  INV_X1     g10723(.I(new_n10915_), .ZN(new_n10916_));
  AOI22_X1   g10724(.A1(new_n10916_), .A2(new_n10414_), .B1(\asqrt[23] ), .B2(new_n10914_), .ZN(new_n10917_));
  NOR3_X1    g10725(.A1(new_n10910_), .A2(new_n10903_), .A3(\asqrt[39] ), .ZN(new_n10918_));
  NOR2_X1    g10726(.A1(new_n10918_), .A2(new_n10917_), .ZN(new_n10919_));
  OAI21_X1   g10727(.A1(new_n10919_), .A2(new_n10912_), .B(\asqrt[40] ), .ZN(new_n10920_));
  INV_X1     g10728(.I(new_n10421_), .ZN(new_n10921_));
  NOR3_X1    g10729(.A1(new_n10812_), .A2(new_n10417_), .A3(new_n10647_), .ZN(new_n10922_));
  INV_X1     g10730(.I(new_n10922_), .ZN(new_n10923_));
  NOR3_X1    g10731(.A1(new_n10647_), .A2(new_n10417_), .A3(new_n10921_), .ZN(new_n10924_));
  AOI22_X1   g10732(.A1(new_n10923_), .A2(new_n10921_), .B1(\asqrt[23] ), .B2(new_n10924_), .ZN(new_n10925_));
  INV_X1     g10733(.I(new_n10925_), .ZN(new_n10926_));
  NAND2_X1   g10734(.A1(new_n10911_), .A2(new_n4071_), .ZN(new_n10927_));
  OAI21_X1   g10735(.A1(new_n10919_), .A2(new_n10927_), .B(new_n10926_), .ZN(new_n10928_));
  AOI21_X1   g10736(.A1(new_n10928_), .A2(new_n10920_), .B(new_n3782_), .ZN(new_n10929_));
  NOR3_X1    g10737(.A1(new_n10426_), .A2(new_n10609_), .A3(new_n10432_), .ZN(new_n10930_));
  NOR3_X1    g10738(.A1(new_n10812_), .A2(new_n10426_), .A3(new_n10432_), .ZN(new_n10931_));
  INV_X1     g10739(.I(new_n10931_), .ZN(new_n10932_));
  AOI22_X1   g10740(.A1(new_n10932_), .A2(new_n10609_), .B1(\asqrt[23] ), .B2(new_n10930_), .ZN(new_n10933_));
  OAI21_X1   g10741(.A1(new_n10917_), .A2(new_n10918_), .B(new_n10911_), .ZN(new_n10934_));
  AOI21_X1   g10742(.A1(new_n10934_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n10935_));
  AOI21_X1   g10743(.A1(new_n10935_), .A2(new_n10928_), .B(new_n10933_), .ZN(new_n10936_));
  OAI21_X1   g10744(.A1(new_n10936_), .A2(new_n10929_), .B(\asqrt[42] ), .ZN(new_n10937_));
  INV_X1     g10745(.I(new_n10937_), .ZN(new_n10938_));
  NOR2_X1    g10746(.A1(new_n10433_), .A2(new_n10441_), .ZN(new_n10939_));
  NOR3_X1    g10747(.A1(new_n10812_), .A2(new_n10646_), .A3(new_n10939_), .ZN(new_n10940_));
  INV_X1     g10748(.I(new_n10940_), .ZN(new_n10941_));
  NOR3_X1    g10749(.A1(new_n10939_), .A2(new_n10646_), .A3(new_n10440_), .ZN(new_n10942_));
  AOI22_X1   g10750(.A1(new_n10941_), .A2(new_n10440_), .B1(\asqrt[23] ), .B2(new_n10942_), .ZN(new_n10943_));
  NOR3_X1    g10751(.A1(new_n10936_), .A2(new_n10929_), .A3(\asqrt[42] ), .ZN(new_n10944_));
  NOR2_X1    g10752(.A1(new_n10944_), .A2(new_n10943_), .ZN(new_n10945_));
  OAI21_X1   g10753(.A1(new_n10945_), .A2(new_n10938_), .B(\asqrt[43] ), .ZN(new_n10946_));
  INV_X1     g10754(.I(new_n10447_), .ZN(new_n10947_));
  NOR3_X1    g10755(.A1(new_n10655_), .A2(new_n10443_), .A3(new_n10947_), .ZN(new_n10948_));
  NOR3_X1    g10756(.A1(new_n10812_), .A2(new_n10443_), .A3(new_n10655_), .ZN(new_n10949_));
  INV_X1     g10757(.I(new_n10949_), .ZN(new_n10950_));
  AOI22_X1   g10758(.A1(new_n10950_), .A2(new_n10947_), .B1(\asqrt[23] ), .B2(new_n10948_), .ZN(new_n10951_));
  INV_X1     g10759(.I(new_n10951_), .ZN(new_n10952_));
  NAND2_X1   g10760(.A1(new_n10937_), .A2(new_n3218_), .ZN(new_n10953_));
  OAI21_X1   g10761(.A1(new_n10945_), .A2(new_n10953_), .B(new_n10952_), .ZN(new_n10954_));
  AOI21_X1   g10762(.A1(new_n10954_), .A2(new_n10946_), .B(new_n2954_), .ZN(new_n10955_));
  NOR3_X1    g10763(.A1(new_n10812_), .A2(new_n10452_), .A3(new_n10460_), .ZN(new_n10956_));
  INV_X1     g10764(.I(new_n10956_), .ZN(new_n10957_));
  NOR3_X1    g10765(.A1(new_n10452_), .A2(new_n10608_), .A3(new_n10460_), .ZN(new_n10958_));
  AOI22_X1   g10766(.A1(new_n10957_), .A2(new_n10608_), .B1(\asqrt[23] ), .B2(new_n10958_), .ZN(new_n10959_));
  OAI21_X1   g10767(.A1(new_n10943_), .A2(new_n10944_), .B(new_n10937_), .ZN(new_n10960_));
  AOI21_X1   g10768(.A1(new_n10960_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n10961_));
  AOI21_X1   g10769(.A1(new_n10961_), .A2(new_n10954_), .B(new_n10959_), .ZN(new_n10962_));
  OAI21_X1   g10770(.A1(new_n10962_), .A2(new_n10955_), .B(\asqrt[45] ), .ZN(new_n10963_));
  INV_X1     g10771(.I(new_n10963_), .ZN(new_n10964_));
  NOR2_X1    g10772(.A1(new_n10461_), .A2(new_n10468_), .ZN(new_n10965_));
  NOR3_X1    g10773(.A1(new_n10965_), .A2(new_n10654_), .A3(new_n10467_), .ZN(new_n10966_));
  NOR3_X1    g10774(.A1(new_n10812_), .A2(new_n10654_), .A3(new_n10965_), .ZN(new_n10967_));
  INV_X1     g10775(.I(new_n10967_), .ZN(new_n10968_));
  AOI22_X1   g10776(.A1(new_n10968_), .A2(new_n10467_), .B1(\asqrt[23] ), .B2(new_n10966_), .ZN(new_n10969_));
  NOR3_X1    g10777(.A1(new_n10962_), .A2(new_n10955_), .A3(\asqrt[45] ), .ZN(new_n10970_));
  NOR2_X1    g10778(.A1(new_n10970_), .A2(new_n10969_), .ZN(new_n10971_));
  OAI21_X1   g10779(.A1(new_n10971_), .A2(new_n10964_), .B(\asqrt[46] ), .ZN(new_n10972_));
  INV_X1     g10780(.I(new_n10476_), .ZN(new_n10973_));
  NOR3_X1    g10781(.A1(new_n10812_), .A2(new_n10470_), .A3(new_n10663_), .ZN(new_n10974_));
  INV_X1     g10782(.I(new_n10974_), .ZN(new_n10975_));
  NOR3_X1    g10783(.A1(new_n10663_), .A2(new_n10470_), .A3(new_n10973_), .ZN(new_n10976_));
  AOI22_X1   g10784(.A1(new_n10975_), .A2(new_n10973_), .B1(\asqrt[23] ), .B2(new_n10976_), .ZN(new_n10977_));
  INV_X1     g10785(.I(new_n10977_), .ZN(new_n10978_));
  NAND2_X1   g10786(.A1(new_n10963_), .A2(new_n2465_), .ZN(new_n10979_));
  OAI21_X1   g10787(.A1(new_n10971_), .A2(new_n10979_), .B(new_n10978_), .ZN(new_n10980_));
  AOI21_X1   g10788(.A1(new_n10980_), .A2(new_n10972_), .B(new_n2229_), .ZN(new_n10981_));
  NOR3_X1    g10789(.A1(new_n10481_), .A2(new_n10607_), .A3(new_n10490_), .ZN(new_n10982_));
  NOR3_X1    g10790(.A1(new_n10812_), .A2(new_n10481_), .A3(new_n10490_), .ZN(new_n10983_));
  INV_X1     g10791(.I(new_n10983_), .ZN(new_n10984_));
  AOI22_X1   g10792(.A1(new_n10984_), .A2(new_n10607_), .B1(\asqrt[23] ), .B2(new_n10982_), .ZN(new_n10985_));
  OAI21_X1   g10793(.A1(new_n10969_), .A2(new_n10970_), .B(new_n10963_), .ZN(new_n10986_));
  AOI21_X1   g10794(.A1(new_n10986_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n10987_));
  AOI21_X1   g10795(.A1(new_n10987_), .A2(new_n10980_), .B(new_n10985_), .ZN(new_n10988_));
  OAI21_X1   g10796(.A1(new_n10988_), .A2(new_n10981_), .B(\asqrt[48] ), .ZN(new_n10989_));
  INV_X1     g10797(.I(new_n10989_), .ZN(new_n10990_));
  NOR2_X1    g10798(.A1(new_n10491_), .A2(new_n10498_), .ZN(new_n10991_));
  NOR3_X1    g10799(.A1(new_n10812_), .A2(new_n10662_), .A3(new_n10991_), .ZN(new_n10992_));
  INV_X1     g10800(.I(new_n10992_), .ZN(new_n10993_));
  NOR3_X1    g10801(.A1(new_n10991_), .A2(new_n10662_), .A3(new_n10497_), .ZN(new_n10994_));
  AOI22_X1   g10802(.A1(new_n10993_), .A2(new_n10497_), .B1(\asqrt[23] ), .B2(new_n10994_), .ZN(new_n10995_));
  NOR3_X1    g10803(.A1(new_n10988_), .A2(new_n10981_), .A3(\asqrt[48] ), .ZN(new_n10996_));
  NOR2_X1    g10804(.A1(new_n10996_), .A2(new_n10995_), .ZN(new_n10997_));
  OAI21_X1   g10805(.A1(new_n10997_), .A2(new_n10990_), .B(\asqrt[49] ), .ZN(new_n10998_));
  INV_X1     g10806(.I(new_n10506_), .ZN(new_n10999_));
  NOR3_X1    g10807(.A1(new_n10671_), .A2(new_n10500_), .A3(new_n10999_), .ZN(new_n11000_));
  NOR3_X1    g10808(.A1(new_n10812_), .A2(new_n10500_), .A3(new_n10671_), .ZN(new_n11001_));
  INV_X1     g10809(.I(new_n11001_), .ZN(new_n11002_));
  AOI22_X1   g10810(.A1(new_n11002_), .A2(new_n10999_), .B1(\asqrt[23] ), .B2(new_n11000_), .ZN(new_n11003_));
  INV_X1     g10811(.I(new_n11003_), .ZN(new_n11004_));
  NAND2_X1   g10812(.A1(new_n10989_), .A2(new_n1806_), .ZN(new_n11005_));
  OAI21_X1   g10813(.A1(new_n10997_), .A2(new_n11005_), .B(new_n11004_), .ZN(new_n11006_));
  AOI21_X1   g10814(.A1(new_n11006_), .A2(new_n10998_), .B(new_n1612_), .ZN(new_n11007_));
  NOR3_X1    g10815(.A1(new_n10812_), .A2(new_n10511_), .A3(new_n10520_), .ZN(new_n11008_));
  INV_X1     g10816(.I(new_n11008_), .ZN(new_n11009_));
  NOR3_X1    g10817(.A1(new_n10511_), .A2(new_n10606_), .A3(new_n10520_), .ZN(new_n11010_));
  AOI22_X1   g10818(.A1(new_n11009_), .A2(new_n10606_), .B1(\asqrt[23] ), .B2(new_n11010_), .ZN(new_n11011_));
  OAI21_X1   g10819(.A1(new_n10995_), .A2(new_n10996_), .B(new_n10989_), .ZN(new_n11012_));
  AOI21_X1   g10820(.A1(new_n11012_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n11013_));
  AOI21_X1   g10821(.A1(new_n11013_), .A2(new_n11006_), .B(new_n11011_), .ZN(new_n11014_));
  OAI21_X1   g10822(.A1(new_n11014_), .A2(new_n11007_), .B(\asqrt[51] ), .ZN(new_n11015_));
  INV_X1     g10823(.I(new_n11015_), .ZN(new_n11016_));
  NOR2_X1    g10824(.A1(new_n10521_), .A2(new_n10528_), .ZN(new_n11017_));
  NOR3_X1    g10825(.A1(new_n11017_), .A2(new_n10670_), .A3(new_n10527_), .ZN(new_n11018_));
  NOR3_X1    g10826(.A1(new_n10812_), .A2(new_n10670_), .A3(new_n11017_), .ZN(new_n11019_));
  INV_X1     g10827(.I(new_n11019_), .ZN(new_n11020_));
  AOI22_X1   g10828(.A1(new_n11020_), .A2(new_n10527_), .B1(\asqrt[23] ), .B2(new_n11018_), .ZN(new_n11021_));
  NOR3_X1    g10829(.A1(new_n11014_), .A2(new_n11007_), .A3(\asqrt[51] ), .ZN(new_n11022_));
  NOR2_X1    g10830(.A1(new_n11022_), .A2(new_n11021_), .ZN(new_n11023_));
  OAI21_X1   g10831(.A1(new_n11023_), .A2(new_n11016_), .B(\asqrt[52] ), .ZN(new_n11024_));
  INV_X1     g10832(.I(new_n10536_), .ZN(new_n11025_));
  NAND2_X1   g10833(.A1(new_n10538_), .A2(new_n10529_), .ZN(new_n11026_));
  INV_X1     g10834(.I(new_n11026_), .ZN(new_n11027_));
  NOR3_X1    g10835(.A1(new_n10812_), .A2(new_n10530_), .A3(new_n11027_), .ZN(new_n11028_));
  INV_X1     g10836(.I(new_n11028_), .ZN(new_n11029_));
  NOR3_X1    g10837(.A1(new_n11027_), .A2(new_n10530_), .A3(new_n11025_), .ZN(new_n11030_));
  AOI22_X1   g10838(.A1(new_n11029_), .A2(new_n11025_), .B1(\asqrt[23] ), .B2(new_n11030_), .ZN(new_n11031_));
  INV_X1     g10839(.I(new_n11031_), .ZN(new_n11032_));
  NAND2_X1   g10840(.A1(new_n11015_), .A2(new_n1256_), .ZN(new_n11033_));
  OAI21_X1   g10841(.A1(new_n11023_), .A2(new_n11033_), .B(new_n11032_), .ZN(new_n11034_));
  AOI21_X1   g10842(.A1(new_n11034_), .A2(new_n11024_), .B(new_n1103_), .ZN(new_n11035_));
  NOR3_X1    g10843(.A1(new_n10541_), .A2(new_n10605_), .A3(new_n10550_), .ZN(new_n11036_));
  NOR3_X1    g10844(.A1(new_n10812_), .A2(new_n10541_), .A3(new_n10550_), .ZN(new_n11037_));
  INV_X1     g10845(.I(new_n11037_), .ZN(new_n11038_));
  AOI22_X1   g10846(.A1(new_n11038_), .A2(new_n10605_), .B1(\asqrt[23] ), .B2(new_n11036_), .ZN(new_n11039_));
  OAI21_X1   g10847(.A1(new_n11021_), .A2(new_n11022_), .B(new_n11015_), .ZN(new_n11040_));
  AOI21_X1   g10848(.A1(new_n11040_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n11041_));
  AOI21_X1   g10849(.A1(new_n11041_), .A2(new_n11034_), .B(new_n11039_), .ZN(new_n11042_));
  OAI21_X1   g10850(.A1(new_n11042_), .A2(new_n11035_), .B(\asqrt[54] ), .ZN(new_n11043_));
  INV_X1     g10851(.I(new_n11043_), .ZN(new_n11044_));
  INV_X1     g10852(.I(new_n10552_), .ZN(new_n11045_));
  INV_X1     g10853(.I(new_n10678_), .ZN(new_n11046_));
  NOR3_X1    g10854(.A1(new_n10812_), .A2(new_n11045_), .A3(new_n11046_), .ZN(new_n11047_));
  INV_X1     g10855(.I(new_n11047_), .ZN(new_n11048_));
  NOR3_X1    g10856(.A1(new_n11045_), .A2(new_n11046_), .A3(new_n10557_), .ZN(new_n11049_));
  AOI22_X1   g10857(.A1(new_n11048_), .A2(new_n10557_), .B1(\asqrt[23] ), .B2(new_n11049_), .ZN(new_n11050_));
  NOR3_X1    g10858(.A1(new_n11042_), .A2(new_n11035_), .A3(\asqrt[54] ), .ZN(new_n11051_));
  NOR2_X1    g10859(.A1(new_n11051_), .A2(new_n11050_), .ZN(new_n11052_));
  OAI21_X1   g10860(.A1(new_n11052_), .A2(new_n11044_), .B(\asqrt[55] ), .ZN(new_n11053_));
  INV_X1     g10861(.I(new_n10566_), .ZN(new_n11054_));
  INV_X1     g10862(.I(new_n10559_), .ZN(new_n11055_));
  INV_X1     g10863(.I(new_n10568_), .ZN(new_n11056_));
  OAI21_X1   g10864(.A1(new_n11056_), .A2(new_n11055_), .B(new_n10566_), .ZN(new_n11057_));
  NOR2_X1    g10865(.A1(new_n11057_), .A2(new_n10560_), .ZN(new_n11058_));
  NOR2_X1    g10866(.A1(new_n11056_), .A2(new_n11055_), .ZN(new_n11059_));
  NOR3_X1    g10867(.A1(new_n10812_), .A2(new_n10560_), .A3(new_n11059_), .ZN(new_n11060_));
  INV_X1     g10868(.I(new_n11060_), .ZN(new_n11061_));
  AOI22_X1   g10869(.A1(new_n11061_), .A2(new_n11054_), .B1(\asqrt[23] ), .B2(new_n11058_), .ZN(new_n11062_));
  INV_X1     g10870(.I(new_n11062_), .ZN(new_n11063_));
  NAND2_X1   g10871(.A1(new_n11043_), .A2(new_n823_), .ZN(new_n11064_));
  OAI21_X1   g10872(.A1(new_n11052_), .A2(new_n11064_), .B(new_n11063_), .ZN(new_n11065_));
  AOI21_X1   g10873(.A1(new_n11065_), .A2(new_n11053_), .B(new_n703_), .ZN(new_n11066_));
  NOR3_X1    g10874(.A1(new_n10812_), .A2(new_n10571_), .A3(new_n10577_), .ZN(new_n11067_));
  INV_X1     g10875(.I(new_n11067_), .ZN(new_n11068_));
  NOR3_X1    g10876(.A1(new_n10571_), .A2(new_n10604_), .A3(new_n10577_), .ZN(new_n11069_));
  AOI22_X1   g10877(.A1(new_n11068_), .A2(new_n10604_), .B1(\asqrt[23] ), .B2(new_n11069_), .ZN(new_n11070_));
  OAI21_X1   g10878(.A1(new_n11050_), .A2(new_n11051_), .B(new_n11043_), .ZN(new_n11071_));
  AOI21_X1   g10879(.A1(new_n11071_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n11072_));
  AOI21_X1   g10880(.A1(new_n11072_), .A2(new_n11065_), .B(new_n11070_), .ZN(new_n11073_));
  OAI21_X1   g10881(.A1(new_n11073_), .A2(new_n11066_), .B(\asqrt[57] ), .ZN(new_n11074_));
  INV_X1     g10882(.I(new_n11074_), .ZN(new_n11075_));
  INV_X1     g10883(.I(new_n10579_), .ZN(new_n11076_));
  INV_X1     g10884(.I(new_n10682_), .ZN(new_n11077_));
  NOR3_X1    g10885(.A1(new_n11076_), .A2(new_n11077_), .A3(new_n10584_), .ZN(new_n11078_));
  NOR3_X1    g10886(.A1(new_n10812_), .A2(new_n11076_), .A3(new_n11077_), .ZN(new_n11079_));
  INV_X1     g10887(.I(new_n11079_), .ZN(new_n11080_));
  AOI22_X1   g10888(.A1(new_n11080_), .A2(new_n10584_), .B1(\asqrt[23] ), .B2(new_n11078_), .ZN(new_n11081_));
  NOR3_X1    g10889(.A1(new_n11073_), .A2(new_n11066_), .A3(\asqrt[57] ), .ZN(new_n11082_));
  NOR2_X1    g10890(.A1(new_n11082_), .A2(new_n11081_), .ZN(new_n11083_));
  OAI21_X1   g10891(.A1(new_n11083_), .A2(new_n11075_), .B(\asqrt[58] ), .ZN(new_n11084_));
  INV_X1     g10892(.I(new_n10593_), .ZN(new_n11085_));
  INV_X1     g10893(.I(new_n10586_), .ZN(new_n11086_));
  INV_X1     g10894(.I(new_n10595_), .ZN(new_n11087_));
  NOR2_X1    g10895(.A1(new_n11087_), .A2(new_n11086_), .ZN(new_n11088_));
  NOR3_X1    g10896(.A1(new_n10812_), .A2(new_n10587_), .A3(new_n11088_), .ZN(new_n11089_));
  INV_X1     g10897(.I(new_n11089_), .ZN(new_n11090_));
  NOR3_X1    g10898(.A1(new_n11088_), .A2(new_n10587_), .A3(new_n11085_), .ZN(new_n11091_));
  AOI22_X1   g10899(.A1(new_n11090_), .A2(new_n11085_), .B1(\asqrt[23] ), .B2(new_n11091_), .ZN(new_n11092_));
  INV_X1     g10900(.I(new_n11092_), .ZN(new_n11093_));
  NAND2_X1   g10901(.A1(new_n11074_), .A2(new_n436_), .ZN(new_n11094_));
  OAI21_X1   g10902(.A1(new_n11083_), .A2(new_n11094_), .B(new_n11093_), .ZN(new_n11095_));
  AOI21_X1   g10903(.A1(new_n11095_), .A2(new_n11084_), .B(new_n327_), .ZN(new_n11096_));
  NOR3_X1    g10904(.A1(new_n10702_), .A2(new_n10603_), .A3(new_n10703_), .ZN(new_n11097_));
  NOR3_X1    g10905(.A1(new_n10812_), .A2(new_n10702_), .A3(new_n10703_), .ZN(new_n11098_));
  INV_X1     g10906(.I(new_n11098_), .ZN(new_n11099_));
  AOI22_X1   g10907(.A1(new_n11099_), .A2(new_n10603_), .B1(\asqrt[23] ), .B2(new_n11097_), .ZN(new_n11100_));
  OAI21_X1   g10908(.A1(new_n11081_), .A2(new_n11082_), .B(new_n11074_), .ZN(new_n11101_));
  AOI21_X1   g10909(.A1(new_n11101_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n11102_));
  AOI21_X1   g10910(.A1(new_n11102_), .A2(new_n11095_), .B(new_n11100_), .ZN(new_n11103_));
  OAI21_X1   g10911(.A1(new_n11103_), .A2(new_n11096_), .B(\asqrt[60] ), .ZN(new_n11104_));
  INV_X1     g10912(.I(new_n11104_), .ZN(new_n11105_));
  INV_X1     g10913(.I(new_n10761_), .ZN(new_n11106_));
  NOR3_X1    g10914(.A1(new_n10812_), .A2(new_n10686_), .A3(new_n11106_), .ZN(new_n11107_));
  INV_X1     g10915(.I(new_n11107_), .ZN(new_n11108_));
  NOR3_X1    g10916(.A1(new_n11106_), .A2(new_n10686_), .A3(new_n10714_), .ZN(new_n11109_));
  AOI22_X1   g10917(.A1(new_n11108_), .A2(new_n10714_), .B1(\asqrt[23] ), .B2(new_n11109_), .ZN(new_n11110_));
  NOR3_X1    g10918(.A1(new_n11103_), .A2(new_n11096_), .A3(\asqrt[60] ), .ZN(new_n11111_));
  NOR2_X1    g10919(.A1(new_n11111_), .A2(new_n11110_), .ZN(new_n11112_));
  OAI21_X1   g10920(.A1(new_n11112_), .A2(new_n11105_), .B(\asqrt[61] ), .ZN(new_n11113_));
  NAND2_X1   g10921(.A1(new_n10726_), .A2(new_n10715_), .ZN(new_n11114_));
  AND3_X2    g10922(.A1(new_n10694_), .A2(new_n10700_), .A3(new_n11114_), .Z(new_n11115_));
  NAND3_X1   g10923(.A1(\asqrt[23] ), .A2(new_n10694_), .A3(new_n11114_), .ZN(new_n11116_));
  AOI22_X1   g10924(.A1(new_n11116_), .A2(new_n10701_), .B1(\asqrt[23] ), .B2(new_n11115_), .ZN(new_n11117_));
  INV_X1     g10925(.I(new_n11117_), .ZN(new_n11118_));
  NAND2_X1   g10926(.A1(new_n11104_), .A2(new_n218_), .ZN(new_n11119_));
  OAI21_X1   g10927(.A1(new_n11112_), .A2(new_n11119_), .B(new_n11118_), .ZN(new_n11120_));
  AOI21_X1   g10928(.A1(new_n11120_), .A2(new_n11113_), .B(new_n207_), .ZN(new_n11121_));
  NOR3_X1    g10929(.A1(new_n10812_), .A2(new_n10708_), .A3(new_n10739_), .ZN(new_n11122_));
  INV_X1     g10930(.I(new_n11122_), .ZN(new_n11123_));
  NOR3_X1    g10931(.A1(new_n10708_), .A2(new_n10760_), .A3(new_n10739_), .ZN(new_n11124_));
  AOI22_X1   g10932(.A1(new_n11123_), .A2(new_n10760_), .B1(\asqrt[23] ), .B2(new_n11124_), .ZN(new_n11125_));
  OAI21_X1   g10933(.A1(new_n11110_), .A2(new_n11111_), .B(new_n11104_), .ZN(new_n11126_));
  AOI21_X1   g10934(.A1(new_n11126_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n11127_));
  AOI21_X1   g10935(.A1(new_n11127_), .A2(new_n11120_), .B(new_n11125_), .ZN(new_n11128_));
  INV_X1     g10936(.I(new_n10719_), .ZN(new_n11129_));
  INV_X1     g10937(.I(new_n10773_), .ZN(new_n11130_));
  NOR3_X1    g10938(.A1(new_n11129_), .A2(new_n11130_), .A3(new_n10724_), .ZN(new_n11131_));
  NAND2_X1   g10939(.A1(\asqrt[23] ), .A2(new_n11131_), .ZN(new_n11132_));
  INV_X1     g10940(.I(new_n11132_), .ZN(new_n11133_));
  NOR2_X1    g10941(.A1(new_n11129_), .A2(new_n11130_), .ZN(new_n11134_));
  AOI21_X1   g10942(.A1(\asqrt[23] ), .A2(new_n11134_), .B(new_n10723_), .ZN(new_n11135_));
  NOR2_X1    g10943(.A1(new_n11133_), .A2(new_n11135_), .ZN(new_n11136_));
  INV_X1     g10944(.I(new_n11136_), .ZN(new_n11137_));
  NAND3_X1   g10945(.A1(\asqrt[23] ), .A2(new_n10757_), .A3(new_n10734_), .ZN(new_n11138_));
  AND3_X2    g10946(.A1(new_n11137_), .A2(new_n10787_), .A3(new_n11138_), .Z(new_n11139_));
  OAI21_X1   g10947(.A1(new_n11128_), .A2(new_n11121_), .B(new_n11139_), .ZN(new_n11140_));
  NAND2_X1   g10948(.A1(new_n11140_), .A2(new_n193_), .ZN(new_n11141_));
  INV_X1     g10949(.I(new_n11110_), .ZN(new_n11142_));
  INV_X1     g10950(.I(new_n11081_), .ZN(new_n11143_));
  INV_X1     g10951(.I(new_n11050_), .ZN(new_n11144_));
  INV_X1     g10952(.I(new_n11021_), .ZN(new_n11145_));
  INV_X1     g10953(.I(new_n10995_), .ZN(new_n11146_));
  INV_X1     g10954(.I(new_n10969_), .ZN(new_n11147_));
  INV_X1     g10955(.I(new_n10943_), .ZN(new_n11148_));
  INV_X1     g10956(.I(new_n10917_), .ZN(new_n11149_));
  INV_X1     g10957(.I(new_n10891_), .ZN(new_n11150_));
  INV_X1     g10958(.I(new_n10865_), .ZN(new_n11151_));
  INV_X1     g10959(.I(new_n10839_), .ZN(new_n11152_));
  NAND2_X1   g10960(.A1(new_n10770_), .A2(new_n10778_), .ZN(new_n11153_));
  OAI21_X1   g10961(.A1(new_n10759_), .A2(new_n10769_), .B(new_n10772_), .ZN(new_n11154_));
  NAND2_X1   g10962(.A1(new_n11154_), .A2(\a[47] ), .ZN(new_n11155_));
  NAND3_X1   g10963(.A1(new_n11153_), .A2(new_n11155_), .A3(new_n10786_), .ZN(new_n11156_));
  AOI21_X1   g10964(.A1(new_n11156_), .A2(new_n10801_), .B(new_n9846_), .ZN(new_n11157_));
  OAI21_X1   g10965(.A1(new_n10792_), .A2(new_n10781_), .B(\a[48] ), .ZN(new_n11158_));
  NAND3_X1   g10966(.A1(new_n10789_), .A2(new_n10786_), .A3(new_n10222_), .ZN(new_n11159_));
  NAND2_X1   g10967(.A1(new_n10770_), .A2(new_n10756_), .ZN(new_n11160_));
  AOI21_X1   g10968(.A1(new_n11160_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n11161_));
  AOI22_X1   g10969(.A1(new_n11156_), .A2(new_n11161_), .B1(new_n11158_), .B2(new_n11159_), .ZN(new_n11162_));
  OAI21_X1   g10970(.A1(new_n11162_), .A2(new_n11157_), .B(\asqrt[26] ), .ZN(new_n11163_));
  NAND2_X1   g10971(.A1(new_n11163_), .A2(new_n8826_), .ZN(new_n11164_));
  OAI21_X1   g10972(.A1(new_n11164_), .A2(new_n10806_), .B(new_n10814_), .ZN(new_n11165_));
  AOI21_X1   g10973(.A1(new_n11165_), .A2(new_n10807_), .B(new_n8483_), .ZN(new_n11166_));
  INV_X1     g10974(.I(new_n10800_), .ZN(new_n11167_));
  AOI21_X1   g10975(.A1(\a[47] ), .A2(new_n11154_), .B(new_n10781_), .ZN(new_n11168_));
  AOI21_X1   g10976(.A1(new_n11168_), .A2(new_n11153_), .B(new_n10771_), .ZN(new_n11169_));
  OAI21_X1   g10977(.A1(new_n11169_), .A2(new_n9846_), .B(new_n9317_), .ZN(new_n11170_));
  OAI21_X1   g10978(.A1(new_n11170_), .A2(new_n11162_), .B(new_n11167_), .ZN(new_n11171_));
  NAND2_X1   g10979(.A1(new_n11171_), .A2(new_n11163_), .ZN(new_n11172_));
  AOI21_X1   g10980(.A1(new_n11172_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n11173_));
  AOI21_X1   g10981(.A1(new_n11173_), .A2(new_n11165_), .B(new_n10822_), .ZN(new_n11174_));
  OAI21_X1   g10982(.A1(new_n11174_), .A2(new_n11166_), .B(\asqrt[29] ), .ZN(new_n11175_));
  NAND2_X1   g10983(.A1(new_n11175_), .A2(new_n7539_), .ZN(new_n11176_));
  OAI21_X1   g10984(.A1(new_n11176_), .A2(new_n10833_), .B(new_n11152_), .ZN(new_n11177_));
  NAND3_X1   g10985(.A1(new_n11177_), .A2(new_n7229_), .A3(new_n10834_), .ZN(new_n11178_));
  AOI22_X1   g10986(.A1(new_n11178_), .A2(new_n10848_), .B1(new_n10856_), .B2(\asqrt[31] ), .ZN(new_n11179_));
  OAI21_X1   g10987(.A1(new_n11179_), .A2(new_n6824_), .B(new_n6356_), .ZN(new_n11180_));
  OAI21_X1   g10988(.A1(new_n11180_), .A2(new_n10858_), .B(new_n11151_), .ZN(new_n11181_));
  AOI21_X1   g10989(.A1(new_n11181_), .A2(new_n10859_), .B(new_n6077_), .ZN(new_n11182_));
  AOI21_X1   g10990(.A1(new_n11177_), .A2(new_n10834_), .B(new_n7229_), .ZN(new_n11183_));
  NOR3_X1    g10991(.A1(new_n11174_), .A2(new_n11166_), .A3(\asqrt[29] ), .ZN(new_n11184_));
  OAI21_X1   g10992(.A1(new_n10830_), .A2(new_n11184_), .B(new_n11175_), .ZN(new_n11185_));
  AOI21_X1   g10993(.A1(new_n11185_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n11186_));
  AOI21_X1   g10994(.A1(new_n11186_), .A2(new_n11177_), .B(new_n10847_), .ZN(new_n11187_));
  NOR3_X1    g10995(.A1(new_n11187_), .A2(\asqrt[32] ), .A3(new_n11183_), .ZN(new_n11188_));
  OAI22_X1   g10996(.A1(new_n11188_), .A2(new_n10855_), .B1(new_n11179_), .B2(new_n6824_), .ZN(new_n11189_));
  AOI21_X1   g10997(.A1(new_n11189_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n11190_));
  AOI21_X1   g10998(.A1(new_n11190_), .A2(new_n11181_), .B(new_n10873_), .ZN(new_n11191_));
  OAI21_X1   g10999(.A1(new_n11191_), .A2(new_n11182_), .B(\asqrt[35] ), .ZN(new_n11192_));
  NAND2_X1   g11000(.A1(new_n11192_), .A2(new_n5277_), .ZN(new_n11193_));
  OAI21_X1   g11001(.A1(new_n11193_), .A2(new_n10884_), .B(new_n11150_), .ZN(new_n11194_));
  AOI21_X1   g11002(.A1(new_n11194_), .A2(new_n10885_), .B(new_n5024_), .ZN(new_n11195_));
  NOR3_X1    g11003(.A1(new_n11191_), .A2(\asqrt[35] ), .A3(new_n11182_), .ZN(new_n11196_));
  OAI21_X1   g11004(.A1(new_n10881_), .A2(new_n11196_), .B(new_n11192_), .ZN(new_n11197_));
  AOI21_X1   g11005(.A1(new_n11197_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n11198_));
  AOI21_X1   g11006(.A1(new_n11198_), .A2(new_n11194_), .B(new_n10899_), .ZN(new_n11199_));
  OAI21_X1   g11007(.A1(new_n11199_), .A2(new_n11195_), .B(\asqrt[38] ), .ZN(new_n11200_));
  NAND2_X1   g11008(.A1(new_n11200_), .A2(new_n4298_), .ZN(new_n11201_));
  OAI21_X1   g11009(.A1(new_n11201_), .A2(new_n10910_), .B(new_n11149_), .ZN(new_n11202_));
  AOI21_X1   g11010(.A1(new_n11202_), .A2(new_n10911_), .B(new_n4071_), .ZN(new_n11203_));
  NOR3_X1    g11011(.A1(new_n11199_), .A2(\asqrt[38] ), .A3(new_n11195_), .ZN(new_n11204_));
  OAI21_X1   g11012(.A1(new_n10907_), .A2(new_n11204_), .B(new_n11200_), .ZN(new_n11205_));
  AOI21_X1   g11013(.A1(new_n11205_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n11206_));
  AOI21_X1   g11014(.A1(new_n11206_), .A2(new_n11202_), .B(new_n10925_), .ZN(new_n11207_));
  OAI21_X1   g11015(.A1(new_n11207_), .A2(new_n11203_), .B(\asqrt[41] ), .ZN(new_n11208_));
  NAND2_X1   g11016(.A1(new_n11208_), .A2(new_n3419_), .ZN(new_n11209_));
  OAI21_X1   g11017(.A1(new_n11209_), .A2(new_n10936_), .B(new_n11148_), .ZN(new_n11210_));
  AOI21_X1   g11018(.A1(new_n11210_), .A2(new_n10937_), .B(new_n3218_), .ZN(new_n11211_));
  NOR3_X1    g11019(.A1(new_n11207_), .A2(\asqrt[41] ), .A3(new_n11203_), .ZN(new_n11212_));
  OAI21_X1   g11020(.A1(new_n10933_), .A2(new_n11212_), .B(new_n11208_), .ZN(new_n11213_));
  AOI21_X1   g11021(.A1(new_n11213_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n11214_));
  AOI21_X1   g11022(.A1(new_n11214_), .A2(new_n11210_), .B(new_n10951_), .ZN(new_n11215_));
  OAI21_X1   g11023(.A1(new_n11215_), .A2(new_n11211_), .B(\asqrt[44] ), .ZN(new_n11216_));
  NAND2_X1   g11024(.A1(new_n11216_), .A2(new_n2641_), .ZN(new_n11217_));
  OAI21_X1   g11025(.A1(new_n11217_), .A2(new_n10962_), .B(new_n11147_), .ZN(new_n11218_));
  AOI21_X1   g11026(.A1(new_n11218_), .A2(new_n10963_), .B(new_n2465_), .ZN(new_n11219_));
  NOR3_X1    g11027(.A1(new_n11215_), .A2(\asqrt[44] ), .A3(new_n11211_), .ZN(new_n11220_));
  OAI21_X1   g11028(.A1(new_n10959_), .A2(new_n11220_), .B(new_n11216_), .ZN(new_n11221_));
  AOI21_X1   g11029(.A1(new_n11221_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n11222_));
  AOI21_X1   g11030(.A1(new_n11222_), .A2(new_n11218_), .B(new_n10977_), .ZN(new_n11223_));
  OAI21_X1   g11031(.A1(new_n11223_), .A2(new_n11219_), .B(\asqrt[47] ), .ZN(new_n11224_));
  NAND2_X1   g11032(.A1(new_n11224_), .A2(new_n1956_), .ZN(new_n11225_));
  OAI21_X1   g11033(.A1(new_n11225_), .A2(new_n10988_), .B(new_n11146_), .ZN(new_n11226_));
  AOI21_X1   g11034(.A1(new_n11226_), .A2(new_n10989_), .B(new_n1806_), .ZN(new_n11227_));
  NOR3_X1    g11035(.A1(new_n11223_), .A2(\asqrt[47] ), .A3(new_n11219_), .ZN(new_n11228_));
  OAI21_X1   g11036(.A1(new_n10985_), .A2(new_n11228_), .B(new_n11224_), .ZN(new_n11229_));
  AOI21_X1   g11037(.A1(new_n11229_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n11230_));
  AOI21_X1   g11038(.A1(new_n11230_), .A2(new_n11226_), .B(new_n11003_), .ZN(new_n11231_));
  OAI21_X1   g11039(.A1(new_n11231_), .A2(new_n11227_), .B(\asqrt[50] ), .ZN(new_n11232_));
  NAND2_X1   g11040(.A1(new_n11232_), .A2(new_n1376_), .ZN(new_n11233_));
  OAI21_X1   g11041(.A1(new_n11233_), .A2(new_n11014_), .B(new_n11145_), .ZN(new_n11234_));
  AOI21_X1   g11042(.A1(new_n11234_), .A2(new_n11015_), .B(new_n1256_), .ZN(new_n11235_));
  NOR3_X1    g11043(.A1(new_n11231_), .A2(\asqrt[50] ), .A3(new_n11227_), .ZN(new_n11236_));
  OAI21_X1   g11044(.A1(new_n11011_), .A2(new_n11236_), .B(new_n11232_), .ZN(new_n11237_));
  AOI21_X1   g11045(.A1(new_n11237_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n11238_));
  AOI21_X1   g11046(.A1(new_n11238_), .A2(new_n11234_), .B(new_n11031_), .ZN(new_n11239_));
  OAI21_X1   g11047(.A1(new_n11239_), .A2(new_n11235_), .B(\asqrt[53] ), .ZN(new_n11240_));
  NAND2_X1   g11048(.A1(new_n11240_), .A2(new_n904_), .ZN(new_n11241_));
  OAI21_X1   g11049(.A1(new_n11241_), .A2(new_n11042_), .B(new_n11144_), .ZN(new_n11242_));
  AOI21_X1   g11050(.A1(new_n11242_), .A2(new_n11043_), .B(new_n823_), .ZN(new_n11243_));
  NOR3_X1    g11051(.A1(new_n11239_), .A2(\asqrt[53] ), .A3(new_n11235_), .ZN(new_n11244_));
  OAI21_X1   g11052(.A1(new_n11039_), .A2(new_n11244_), .B(new_n11240_), .ZN(new_n11245_));
  AOI21_X1   g11053(.A1(new_n11245_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n11246_));
  AOI21_X1   g11054(.A1(new_n11246_), .A2(new_n11242_), .B(new_n11062_), .ZN(new_n11247_));
  OAI21_X1   g11055(.A1(new_n11247_), .A2(new_n11243_), .B(\asqrt[56] ), .ZN(new_n11248_));
  NAND2_X1   g11056(.A1(new_n11248_), .A2(new_n531_), .ZN(new_n11249_));
  OAI21_X1   g11057(.A1(new_n11249_), .A2(new_n11073_), .B(new_n11143_), .ZN(new_n11250_));
  AOI21_X1   g11058(.A1(new_n11250_), .A2(new_n11074_), .B(new_n436_), .ZN(new_n11251_));
  NOR3_X1    g11059(.A1(new_n11247_), .A2(\asqrt[56] ), .A3(new_n11243_), .ZN(new_n11252_));
  OAI21_X1   g11060(.A1(new_n11070_), .A2(new_n11252_), .B(new_n11248_), .ZN(new_n11253_));
  AOI21_X1   g11061(.A1(new_n11253_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n11254_));
  AOI21_X1   g11062(.A1(new_n11254_), .A2(new_n11250_), .B(new_n11092_), .ZN(new_n11255_));
  OAI21_X1   g11063(.A1(new_n11255_), .A2(new_n11251_), .B(\asqrt[59] ), .ZN(new_n11256_));
  NAND2_X1   g11064(.A1(new_n11256_), .A2(new_n306_), .ZN(new_n11257_));
  OAI21_X1   g11065(.A1(new_n11257_), .A2(new_n11103_), .B(new_n11142_), .ZN(new_n11258_));
  NOR3_X1    g11066(.A1(new_n11255_), .A2(\asqrt[59] ), .A3(new_n11251_), .ZN(new_n11259_));
  OAI21_X1   g11067(.A1(new_n11100_), .A2(new_n11259_), .B(new_n11256_), .ZN(new_n11260_));
  AOI21_X1   g11068(.A1(new_n11260_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n11261_));
  AOI21_X1   g11069(.A1(new_n11261_), .A2(new_n11258_), .B(new_n11117_), .ZN(new_n11262_));
  INV_X1     g11070(.I(new_n11125_), .ZN(new_n11263_));
  NAND2_X1   g11071(.A1(new_n11113_), .A2(new_n207_), .ZN(new_n11264_));
  OAI21_X1   g11072(.A1(new_n11264_), .A2(new_n11262_), .B(new_n11263_), .ZN(new_n11265_));
  NOR2_X1    g11073(.A1(new_n11121_), .A2(new_n11137_), .ZN(new_n11266_));
  NAND2_X1   g11074(.A1(\asqrt[23] ), .A2(new_n10734_), .ZN(new_n11267_));
  OAI21_X1   g11075(.A1(new_n10774_), .A2(new_n10767_), .B(\asqrt[63] ), .ZN(new_n11268_));
  AOI21_X1   g11076(.A1(new_n11267_), .A2(new_n10774_), .B(new_n11268_), .ZN(new_n11269_));
  AND2_X2    g11077(.A1(new_n10731_), .A2(new_n10747_), .Z(new_n11270_));
  NAND4_X1   g11078(.A1(new_n10787_), .A2(new_n10733_), .A3(new_n10744_), .A4(new_n11270_), .ZN(new_n11271_));
  NOR2_X1    g11079(.A1(new_n11271_), .A2(new_n10759_), .ZN(new_n11272_));
  NOR2_X1    g11080(.A1(new_n11269_), .A2(new_n11272_), .ZN(new_n11273_));
  INV_X1     g11081(.I(new_n11273_), .ZN(new_n11274_));
  AOI21_X1   g11082(.A1(new_n11266_), .A2(new_n11265_), .B(new_n11274_), .ZN(new_n11275_));
  NAND2_X1   g11083(.A1(new_n11141_), .A2(new_n11275_), .ZN(\asqrt[22] ));
  NOR2_X1    g11084(.A1(\a[42] ), .A2(\a[43] ), .ZN(new_n11277_));
  INV_X1     g11085(.I(new_n11277_), .ZN(new_n11278_));
  NOR2_X1    g11086(.A1(new_n11278_), .A2(\a[44] ), .ZN(new_n11279_));
  INV_X1     g11087(.I(new_n11279_), .ZN(new_n11280_));
  AOI21_X1   g11088(.A1(new_n11258_), .A2(new_n11104_), .B(new_n218_), .ZN(new_n11281_));
  OAI21_X1   g11089(.A1(new_n11262_), .A2(new_n11281_), .B(\asqrt[62] ), .ZN(new_n11282_));
  NOR3_X1    g11090(.A1(new_n11262_), .A2(\asqrt[62] ), .A3(new_n11281_), .ZN(new_n11283_));
  OAI21_X1   g11091(.A1(new_n11125_), .A2(new_n11283_), .B(new_n11282_), .ZN(new_n11284_));
  AOI21_X1   g11092(.A1(new_n11284_), .A2(new_n11139_), .B(\asqrt[63] ), .ZN(new_n11285_));
  NAND2_X1   g11093(.A1(new_n11282_), .A2(new_n11136_), .ZN(new_n11286_));
  OAI21_X1   g11094(.A1(new_n11286_), .A2(new_n11128_), .B(new_n11273_), .ZN(new_n11287_));
  OAI21_X1   g11095(.A1(new_n11285_), .A2(new_n11287_), .B(\a[44] ), .ZN(new_n11288_));
  AOI21_X1   g11096(.A1(new_n11288_), .A2(new_n11280_), .B(new_n10812_), .ZN(new_n11289_));
  INV_X1     g11097(.I(\a[44] ), .ZN(new_n11290_));
  AOI21_X1   g11098(.A1(new_n11141_), .A2(new_n11275_), .B(new_n11290_), .ZN(new_n11291_));
  NAND4_X1   g11099(.A1(new_n10787_), .A2(new_n10744_), .A3(new_n10747_), .A4(new_n11280_), .ZN(new_n11292_));
  NOR2_X1    g11100(.A1(new_n11292_), .A2(new_n10759_), .ZN(new_n11293_));
  INV_X1     g11101(.I(new_n11293_), .ZN(new_n11294_));
  NOR2_X1    g11102(.A1(new_n11291_), .A2(new_n11294_), .ZN(new_n11295_));
  AOI21_X1   g11103(.A1(new_n11141_), .A2(new_n11275_), .B(new_n10754_), .ZN(new_n11296_));
  INV_X1     g11104(.I(\a[45] ), .ZN(new_n11297_));
  AOI21_X1   g11105(.A1(\asqrt[22] ), .A2(new_n11290_), .B(new_n11297_), .ZN(new_n11298_));
  NOR3_X1    g11106(.A1(new_n11295_), .A2(new_n11298_), .A3(new_n11296_), .ZN(new_n11299_));
  OAI21_X1   g11107(.A1(new_n11299_), .A2(new_n11289_), .B(\asqrt[24] ), .ZN(new_n11300_));
  OAI21_X1   g11108(.A1(new_n11285_), .A2(new_n11287_), .B(new_n10753_), .ZN(new_n11301_));
  NAND2_X1   g11109(.A1(new_n11266_), .A2(new_n11265_), .ZN(new_n11302_));
  NOR3_X1    g11110(.A1(new_n11269_), .A2(new_n10812_), .A3(new_n11272_), .ZN(new_n11303_));
  NAND3_X1   g11111(.A1(new_n11141_), .A2(new_n11302_), .A3(new_n11303_), .ZN(new_n11304_));
  AOI21_X1   g11112(.A1(new_n11301_), .A2(new_n11304_), .B(new_n10772_), .ZN(new_n11305_));
  AND3_X2    g11113(.A1(new_n11141_), .A2(new_n11302_), .A3(new_n11303_), .Z(new_n11306_));
  NOR3_X1    g11114(.A1(new_n11306_), .A2(\a[46] ), .A3(new_n11296_), .ZN(new_n11307_));
  OAI21_X1   g11115(.A1(new_n11291_), .A2(new_n11279_), .B(\asqrt[23] ), .ZN(new_n11308_));
  NAND2_X1   g11116(.A1(new_n11308_), .A2(new_n10221_), .ZN(new_n11309_));
  OAI22_X1   g11117(.A1(new_n11299_), .A2(new_n11309_), .B1(new_n11305_), .B2(new_n11307_), .ZN(new_n11310_));
  AOI21_X1   g11118(.A1(new_n11310_), .A2(new_n11300_), .B(new_n9846_), .ZN(new_n11311_));
  NOR3_X1    g11119(.A1(new_n11168_), .A2(new_n10771_), .A3(new_n10780_), .ZN(new_n11312_));
  NAND3_X1   g11120(.A1(\asqrt[22] ), .A2(new_n10801_), .A3(new_n11153_), .ZN(new_n11313_));
  AOI22_X1   g11121(.A1(new_n11313_), .A2(new_n11168_), .B1(\asqrt[22] ), .B2(new_n11312_), .ZN(new_n11314_));
  AOI21_X1   g11122(.A1(new_n11141_), .A2(new_n11275_), .B(\a[44] ), .ZN(new_n11315_));
  OAI21_X1   g11123(.A1(new_n11297_), .A2(new_n11315_), .B(new_n11301_), .ZN(new_n11316_));
  OAI21_X1   g11124(.A1(new_n11316_), .A2(new_n11295_), .B(new_n11308_), .ZN(new_n11317_));
  AOI21_X1   g11125(.A1(new_n11317_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n11318_));
  AOI21_X1   g11126(.A1(new_n11318_), .A2(new_n11310_), .B(new_n11314_), .ZN(new_n11319_));
  OAI21_X1   g11127(.A1(new_n11319_), .A2(new_n11311_), .B(\asqrt[26] ), .ZN(new_n11320_));
  INV_X1     g11128(.I(new_n11320_), .ZN(new_n11321_));
  NOR2_X1    g11129(.A1(new_n10793_), .A2(new_n10790_), .ZN(new_n11322_));
  NOR2_X1    g11130(.A1(new_n10784_), .A2(new_n10795_), .ZN(new_n11323_));
  INV_X1     g11131(.I(new_n11323_), .ZN(new_n11324_));
  NAND4_X1   g11132(.A1(\asqrt[22] ), .A2(new_n10785_), .A3(new_n11322_), .A4(new_n11324_), .ZN(new_n11325_));
  INV_X1     g11133(.I(\asqrt[22] ), .ZN(new_n11326_));
  NOR3_X1    g11134(.A1(new_n11326_), .A2(new_n11157_), .A3(new_n11323_), .ZN(new_n11327_));
  OAI21_X1   g11135(.A1(new_n11327_), .A2(new_n11322_), .B(new_n11325_), .ZN(new_n11328_));
  INV_X1     g11136(.I(new_n11328_), .ZN(new_n11329_));
  NOR3_X1    g11137(.A1(new_n11319_), .A2(new_n11311_), .A3(\asqrt[26] ), .ZN(new_n11330_));
  NOR2_X1    g11138(.A1(new_n11330_), .A2(new_n11329_), .ZN(new_n11331_));
  OAI21_X1   g11139(.A1(new_n11331_), .A2(new_n11321_), .B(\asqrt[27] ), .ZN(new_n11332_));
  NOR2_X1    g11140(.A1(new_n11170_), .A2(new_n11162_), .ZN(new_n11333_));
  NOR3_X1    g11141(.A1(new_n11326_), .A2(new_n10797_), .A3(new_n11333_), .ZN(new_n11334_));
  INV_X1     g11142(.I(new_n11334_), .ZN(new_n11335_));
  NOR3_X1    g11143(.A1(new_n11333_), .A2(new_n10797_), .A3(new_n11167_), .ZN(new_n11336_));
  AOI22_X1   g11144(.A1(new_n11335_), .A2(new_n11167_), .B1(\asqrt[22] ), .B2(new_n11336_), .ZN(new_n11337_));
  INV_X1     g11145(.I(new_n11337_), .ZN(new_n11338_));
  NAND2_X1   g11146(.A1(new_n11320_), .A2(new_n8826_), .ZN(new_n11339_));
  OAI21_X1   g11147(.A1(new_n11331_), .A2(new_n11339_), .B(new_n11338_), .ZN(new_n11340_));
  AOI21_X1   g11148(.A1(new_n11340_), .A2(new_n11332_), .B(new_n8483_), .ZN(new_n11341_));
  NOR3_X1    g11149(.A1(new_n10808_), .A2(new_n10816_), .A3(new_n10814_), .ZN(new_n11342_));
  NOR3_X1    g11150(.A1(new_n11326_), .A2(new_n10808_), .A3(new_n10816_), .ZN(new_n11343_));
  INV_X1     g11151(.I(new_n11343_), .ZN(new_n11344_));
  AOI22_X1   g11152(.A1(new_n11344_), .A2(new_n10814_), .B1(\asqrt[22] ), .B2(new_n11342_), .ZN(new_n11345_));
  OAI21_X1   g11153(.A1(new_n11329_), .A2(new_n11330_), .B(new_n11320_), .ZN(new_n11346_));
  AOI21_X1   g11154(.A1(new_n11346_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n11347_));
  AOI21_X1   g11155(.A1(new_n11347_), .A2(new_n11340_), .B(new_n11345_), .ZN(new_n11348_));
  OAI21_X1   g11156(.A1(new_n11348_), .A2(new_n11341_), .B(\asqrt[29] ), .ZN(new_n11349_));
  NAND2_X1   g11157(.A1(new_n11173_), .A2(new_n11165_), .ZN(new_n11350_));
  NAND3_X1   g11158(.A1(\asqrt[22] ), .A2(new_n10818_), .A3(new_n11350_), .ZN(new_n11351_));
  AND3_X2    g11159(.A1(new_n10818_), .A2(new_n10822_), .A3(new_n11350_), .Z(new_n11352_));
  AOI22_X1   g11160(.A1(new_n11351_), .A2(new_n10823_), .B1(\asqrt[22] ), .B2(new_n11352_), .ZN(new_n11353_));
  INV_X1     g11161(.I(new_n11353_), .ZN(new_n11354_));
  NAND2_X1   g11162(.A1(new_n11288_), .A2(new_n11293_), .ZN(new_n11355_));
  OAI21_X1   g11163(.A1(new_n11285_), .A2(new_n11287_), .B(new_n11290_), .ZN(new_n11356_));
  NAND2_X1   g11164(.A1(new_n11356_), .A2(\a[45] ), .ZN(new_n11357_));
  NAND3_X1   g11165(.A1(new_n11355_), .A2(new_n11357_), .A3(new_n11301_), .ZN(new_n11358_));
  AOI21_X1   g11166(.A1(new_n11358_), .A2(new_n11308_), .B(new_n10221_), .ZN(new_n11359_));
  OAI21_X1   g11167(.A1(new_n11306_), .A2(new_n11296_), .B(\a[46] ), .ZN(new_n11360_));
  NAND3_X1   g11168(.A1(new_n11301_), .A2(new_n11304_), .A3(new_n10772_), .ZN(new_n11361_));
  NAND2_X1   g11169(.A1(new_n11288_), .A2(new_n11280_), .ZN(new_n11362_));
  AOI21_X1   g11170(.A1(new_n11362_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n11363_));
  AOI22_X1   g11171(.A1(new_n11358_), .A2(new_n11363_), .B1(new_n11360_), .B2(new_n11361_), .ZN(new_n11364_));
  OAI21_X1   g11172(.A1(new_n11364_), .A2(new_n11359_), .B(\asqrt[25] ), .ZN(new_n11365_));
  NAND2_X1   g11173(.A1(new_n11365_), .A2(new_n9317_), .ZN(new_n11366_));
  OAI21_X1   g11174(.A1(new_n11366_), .A2(new_n11319_), .B(new_n11328_), .ZN(new_n11367_));
  AOI21_X1   g11175(.A1(new_n11367_), .A2(new_n11320_), .B(new_n8826_), .ZN(new_n11368_));
  INV_X1     g11176(.I(new_n11314_), .ZN(new_n11369_));
  AOI21_X1   g11177(.A1(\a[45] ), .A2(new_n11356_), .B(new_n11296_), .ZN(new_n11370_));
  AOI21_X1   g11178(.A1(new_n11370_), .A2(new_n11355_), .B(new_n11289_), .ZN(new_n11371_));
  OAI21_X1   g11179(.A1(new_n11371_), .A2(new_n10221_), .B(new_n9846_), .ZN(new_n11372_));
  OAI21_X1   g11180(.A1(new_n11372_), .A2(new_n11364_), .B(new_n11369_), .ZN(new_n11373_));
  NAND2_X1   g11181(.A1(new_n11373_), .A2(new_n11365_), .ZN(new_n11374_));
  AOI21_X1   g11182(.A1(new_n11374_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n11375_));
  AOI21_X1   g11183(.A1(new_n11375_), .A2(new_n11367_), .B(new_n11337_), .ZN(new_n11376_));
  OAI21_X1   g11184(.A1(new_n11376_), .A2(new_n11368_), .B(\asqrt[28] ), .ZN(new_n11377_));
  NAND2_X1   g11185(.A1(new_n11377_), .A2(new_n8036_), .ZN(new_n11378_));
  OAI21_X1   g11186(.A1(new_n11378_), .A2(new_n11348_), .B(new_n11354_), .ZN(new_n11379_));
  AOI21_X1   g11187(.A1(new_n11379_), .A2(new_n11349_), .B(new_n7539_), .ZN(new_n11380_));
  INV_X1     g11188(.I(new_n11380_), .ZN(new_n11381_));
  INV_X1     g11189(.I(new_n10830_), .ZN(new_n11382_));
  NOR3_X1    g11190(.A1(new_n10826_), .A2(new_n11184_), .A3(new_n11382_), .ZN(new_n11383_));
  NOR3_X1    g11191(.A1(new_n11326_), .A2(new_n10826_), .A3(new_n11184_), .ZN(new_n11384_));
  INV_X1     g11192(.I(new_n11384_), .ZN(new_n11385_));
  AOI22_X1   g11193(.A1(new_n11385_), .A2(new_n11382_), .B1(\asqrt[22] ), .B2(new_n11383_), .ZN(new_n11386_));
  INV_X1     g11194(.I(new_n11386_), .ZN(new_n11387_));
  NAND3_X1   g11195(.A1(new_n11379_), .A2(new_n7539_), .A3(new_n11349_), .ZN(new_n11388_));
  NAND2_X1   g11196(.A1(new_n11388_), .A2(new_n11387_), .ZN(new_n11389_));
  AOI21_X1   g11197(.A1(new_n11389_), .A2(new_n11381_), .B(new_n7229_), .ZN(new_n11390_));
  NOR3_X1    g11198(.A1(new_n11326_), .A2(new_n10835_), .A3(new_n10840_), .ZN(new_n11391_));
  INV_X1     g11199(.I(new_n11391_), .ZN(new_n11392_));
  NOR3_X1    g11200(.A1(new_n10835_), .A2(new_n11152_), .A3(new_n10840_), .ZN(new_n11393_));
  AOI22_X1   g11201(.A1(new_n11392_), .A2(new_n11152_), .B1(\asqrt[22] ), .B2(new_n11393_), .ZN(new_n11394_));
  NOR2_X1    g11202(.A1(new_n11380_), .A2(\asqrt[31] ), .ZN(new_n11395_));
  AOI21_X1   g11203(.A1(new_n11395_), .A2(new_n11389_), .B(new_n11394_), .ZN(new_n11396_));
  OAI21_X1   g11204(.A1(new_n11396_), .A2(new_n11390_), .B(\asqrt[32] ), .ZN(new_n11397_));
  INV_X1     g11205(.I(new_n11178_), .ZN(new_n11398_));
  NOR3_X1    g11206(.A1(new_n11398_), .A2(new_n11183_), .A3(new_n10848_), .ZN(new_n11399_));
  NOR3_X1    g11207(.A1(new_n11326_), .A2(new_n11183_), .A3(new_n11398_), .ZN(new_n11400_));
  INV_X1     g11208(.I(new_n11400_), .ZN(new_n11401_));
  AOI22_X1   g11209(.A1(new_n11401_), .A2(new_n10848_), .B1(\asqrt[22] ), .B2(new_n11399_), .ZN(new_n11402_));
  INV_X1     g11210(.I(new_n11402_), .ZN(new_n11403_));
  NOR3_X1    g11211(.A1(new_n11348_), .A2(new_n11341_), .A3(\asqrt[29] ), .ZN(new_n11404_));
  OAI21_X1   g11212(.A1(new_n11353_), .A2(new_n11404_), .B(new_n11349_), .ZN(new_n11405_));
  AOI22_X1   g11213(.A1(new_n11388_), .A2(new_n11387_), .B1(new_n11405_), .B2(\asqrt[30] ), .ZN(new_n11406_));
  OAI21_X1   g11214(.A1(new_n11406_), .A2(new_n7229_), .B(new_n6824_), .ZN(new_n11407_));
  OAI21_X1   g11215(.A1(new_n11407_), .A2(new_n11396_), .B(new_n11403_), .ZN(new_n11408_));
  AOI21_X1   g11216(.A1(new_n11408_), .A2(new_n11397_), .B(new_n6356_), .ZN(new_n11409_));
  INV_X1     g11217(.I(new_n11409_), .ZN(new_n11410_));
  INV_X1     g11218(.I(new_n11408_), .ZN(new_n11411_));
  INV_X1     g11219(.I(new_n10855_), .ZN(new_n11412_));
  NOR3_X1    g11220(.A1(new_n11326_), .A2(new_n10851_), .A3(new_n11188_), .ZN(new_n11413_));
  INV_X1     g11221(.I(new_n11413_), .ZN(new_n11414_));
  NOR3_X1    g11222(.A1(new_n10851_), .A2(new_n11188_), .A3(new_n11412_), .ZN(new_n11415_));
  AOI22_X1   g11223(.A1(new_n11414_), .A2(new_n11412_), .B1(\asqrt[22] ), .B2(new_n11415_), .ZN(new_n11416_));
  INV_X1     g11224(.I(new_n11416_), .ZN(new_n11417_));
  NAND2_X1   g11225(.A1(new_n11397_), .A2(new_n6356_), .ZN(new_n11418_));
  OAI21_X1   g11226(.A1(new_n11411_), .A2(new_n11418_), .B(new_n11417_), .ZN(new_n11419_));
  AOI21_X1   g11227(.A1(new_n11419_), .A2(new_n11410_), .B(new_n6077_), .ZN(new_n11420_));
  NOR3_X1    g11228(.A1(new_n10860_), .A2(new_n11151_), .A3(new_n10866_), .ZN(new_n11421_));
  NOR3_X1    g11229(.A1(new_n11326_), .A2(new_n10860_), .A3(new_n10866_), .ZN(new_n11422_));
  INV_X1     g11230(.I(new_n11422_), .ZN(new_n11423_));
  AOI22_X1   g11231(.A1(new_n11423_), .A2(new_n11151_), .B1(\asqrt[22] ), .B2(new_n11421_), .ZN(new_n11424_));
  NOR2_X1    g11232(.A1(new_n11409_), .A2(\asqrt[34] ), .ZN(new_n11425_));
  AOI21_X1   g11233(.A1(new_n11425_), .A2(new_n11419_), .B(new_n11424_), .ZN(new_n11426_));
  OAI21_X1   g11234(.A1(new_n11426_), .A2(new_n11420_), .B(\asqrt[35] ), .ZN(new_n11427_));
  NOR2_X1    g11235(.A1(new_n10867_), .A2(new_n10875_), .ZN(new_n11428_));
  NOR3_X1    g11236(.A1(new_n11326_), .A2(new_n11182_), .A3(new_n11428_), .ZN(new_n11429_));
  INV_X1     g11237(.I(new_n11429_), .ZN(new_n11430_));
  NOR3_X1    g11238(.A1(new_n11428_), .A2(new_n11182_), .A3(new_n10874_), .ZN(new_n11431_));
  AOI22_X1   g11239(.A1(new_n11430_), .A2(new_n10874_), .B1(\asqrt[22] ), .B2(new_n11431_), .ZN(new_n11432_));
  INV_X1     g11240(.I(new_n11432_), .ZN(new_n11433_));
  NOR3_X1    g11241(.A1(new_n11376_), .A2(new_n11368_), .A3(\asqrt[28] ), .ZN(new_n11434_));
  OAI21_X1   g11242(.A1(new_n11345_), .A2(new_n11434_), .B(new_n11377_), .ZN(new_n11435_));
  AOI21_X1   g11243(.A1(new_n11435_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n11436_));
  AOI21_X1   g11244(.A1(new_n11436_), .A2(new_n11379_), .B(new_n11386_), .ZN(new_n11437_));
  NOR3_X1    g11245(.A1(new_n11437_), .A2(\asqrt[31] ), .A3(new_n11380_), .ZN(new_n11438_));
  OAI22_X1   g11246(.A1(new_n11438_), .A2(new_n11394_), .B1(new_n11406_), .B2(new_n7229_), .ZN(new_n11439_));
  AOI21_X1   g11247(.A1(new_n11439_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n11440_));
  AOI21_X1   g11248(.A1(new_n11440_), .A2(new_n11408_), .B(new_n11416_), .ZN(new_n11441_));
  OAI21_X1   g11249(.A1(new_n11441_), .A2(new_n11409_), .B(\asqrt[34] ), .ZN(new_n11442_));
  NAND2_X1   g11250(.A1(new_n11442_), .A2(new_n5708_), .ZN(new_n11443_));
  OAI21_X1   g11251(.A1(new_n11443_), .A2(new_n11426_), .B(new_n11433_), .ZN(new_n11444_));
  NAND2_X1   g11252(.A1(new_n11444_), .A2(new_n11427_), .ZN(new_n11445_));
  NAND2_X1   g11253(.A1(new_n11445_), .A2(\asqrt[36] ), .ZN(new_n11446_));
  INV_X1     g11254(.I(new_n11444_), .ZN(new_n11447_));
  INV_X1     g11255(.I(new_n10881_), .ZN(new_n11448_));
  NOR3_X1    g11256(.A1(new_n10877_), .A2(new_n11196_), .A3(new_n11448_), .ZN(new_n11449_));
  NOR3_X1    g11257(.A1(new_n11326_), .A2(new_n10877_), .A3(new_n11196_), .ZN(new_n11450_));
  INV_X1     g11258(.I(new_n11450_), .ZN(new_n11451_));
  AOI22_X1   g11259(.A1(new_n11451_), .A2(new_n11448_), .B1(\asqrt[22] ), .B2(new_n11449_), .ZN(new_n11452_));
  INV_X1     g11260(.I(new_n11452_), .ZN(new_n11453_));
  NAND2_X1   g11261(.A1(new_n11427_), .A2(new_n5277_), .ZN(new_n11454_));
  OAI21_X1   g11262(.A1(new_n11447_), .A2(new_n11454_), .B(new_n11453_), .ZN(new_n11455_));
  AOI21_X1   g11263(.A1(new_n11455_), .A2(new_n11446_), .B(new_n5024_), .ZN(new_n11456_));
  NOR3_X1    g11264(.A1(new_n11326_), .A2(new_n10886_), .A3(new_n10892_), .ZN(new_n11457_));
  INV_X1     g11265(.I(new_n11457_), .ZN(new_n11458_));
  NOR3_X1    g11266(.A1(new_n10886_), .A2(new_n11150_), .A3(new_n10892_), .ZN(new_n11459_));
  AOI22_X1   g11267(.A1(new_n11458_), .A2(new_n11150_), .B1(\asqrt[22] ), .B2(new_n11459_), .ZN(new_n11460_));
  AOI21_X1   g11268(.A1(new_n11444_), .A2(new_n11427_), .B(new_n5277_), .ZN(new_n11461_));
  NOR2_X1    g11269(.A1(new_n11461_), .A2(\asqrt[37] ), .ZN(new_n11462_));
  AOI21_X1   g11270(.A1(new_n11462_), .A2(new_n11455_), .B(new_n11460_), .ZN(new_n11463_));
  OAI21_X1   g11271(.A1(new_n11463_), .A2(new_n11456_), .B(\asqrt[38] ), .ZN(new_n11464_));
  INV_X1     g11272(.I(new_n11464_), .ZN(new_n11465_));
  NOR2_X1    g11273(.A1(new_n10893_), .A2(new_n10901_), .ZN(new_n11466_));
  NOR3_X1    g11274(.A1(new_n11466_), .A2(new_n11195_), .A3(new_n10900_), .ZN(new_n11467_));
  NOR3_X1    g11275(.A1(new_n11326_), .A2(new_n11195_), .A3(new_n11466_), .ZN(new_n11468_));
  INV_X1     g11276(.I(new_n11468_), .ZN(new_n11469_));
  AOI22_X1   g11277(.A1(new_n11469_), .A2(new_n10900_), .B1(\asqrt[22] ), .B2(new_n11467_), .ZN(new_n11470_));
  NOR3_X1    g11278(.A1(new_n11463_), .A2(new_n11456_), .A3(\asqrt[38] ), .ZN(new_n11471_));
  NOR2_X1    g11279(.A1(new_n11471_), .A2(new_n11470_), .ZN(new_n11472_));
  OAI21_X1   g11280(.A1(new_n11472_), .A2(new_n11465_), .B(\asqrt[39] ), .ZN(new_n11473_));
  INV_X1     g11281(.I(new_n10907_), .ZN(new_n11474_));
  NOR3_X1    g11282(.A1(new_n11326_), .A2(new_n10903_), .A3(new_n11204_), .ZN(new_n11475_));
  INV_X1     g11283(.I(new_n11475_), .ZN(new_n11476_));
  NOR3_X1    g11284(.A1(new_n10903_), .A2(new_n11204_), .A3(new_n11474_), .ZN(new_n11477_));
  AOI22_X1   g11285(.A1(new_n11476_), .A2(new_n11474_), .B1(\asqrt[22] ), .B2(new_n11477_), .ZN(new_n11478_));
  INV_X1     g11286(.I(new_n11478_), .ZN(new_n11479_));
  NAND2_X1   g11287(.A1(new_n11464_), .A2(new_n4298_), .ZN(new_n11480_));
  OAI21_X1   g11288(.A1(new_n11472_), .A2(new_n11480_), .B(new_n11479_), .ZN(new_n11481_));
  AOI21_X1   g11289(.A1(new_n11481_), .A2(new_n11473_), .B(new_n4071_), .ZN(new_n11482_));
  NOR3_X1    g11290(.A1(new_n10912_), .A2(new_n11149_), .A3(new_n10918_), .ZN(new_n11483_));
  NOR3_X1    g11291(.A1(new_n11326_), .A2(new_n10912_), .A3(new_n10918_), .ZN(new_n11484_));
  INV_X1     g11292(.I(new_n11484_), .ZN(new_n11485_));
  AOI22_X1   g11293(.A1(new_n11485_), .A2(new_n11149_), .B1(\asqrt[22] ), .B2(new_n11483_), .ZN(new_n11486_));
  INV_X1     g11294(.I(new_n11470_), .ZN(new_n11487_));
  NOR3_X1    g11295(.A1(new_n11441_), .A2(\asqrt[34] ), .A3(new_n11409_), .ZN(new_n11488_));
  OAI21_X1   g11296(.A1(new_n11424_), .A2(new_n11488_), .B(new_n11442_), .ZN(new_n11489_));
  AOI21_X1   g11297(.A1(new_n11489_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n11490_));
  AOI21_X1   g11298(.A1(new_n11490_), .A2(new_n11444_), .B(new_n11452_), .ZN(new_n11491_));
  OAI21_X1   g11299(.A1(new_n11491_), .A2(new_n11461_), .B(\asqrt[37] ), .ZN(new_n11492_));
  NAND2_X1   g11300(.A1(new_n11492_), .A2(new_n4696_), .ZN(new_n11493_));
  OAI21_X1   g11301(.A1(new_n11493_), .A2(new_n11463_), .B(new_n11487_), .ZN(new_n11494_));
  AOI21_X1   g11302(.A1(new_n11494_), .A2(new_n11464_), .B(new_n4298_), .ZN(new_n11495_));
  NOR2_X1    g11303(.A1(new_n11495_), .A2(\asqrt[40] ), .ZN(new_n11496_));
  AOI21_X1   g11304(.A1(new_n11496_), .A2(new_n11481_), .B(new_n11486_), .ZN(new_n11497_));
  OAI21_X1   g11305(.A1(new_n11497_), .A2(new_n11482_), .B(\asqrt[41] ), .ZN(new_n11498_));
  NOR2_X1    g11306(.A1(new_n10919_), .A2(new_n10927_), .ZN(new_n11499_));
  NOR3_X1    g11307(.A1(new_n11326_), .A2(new_n11203_), .A3(new_n11499_), .ZN(new_n11500_));
  INV_X1     g11308(.I(new_n11500_), .ZN(new_n11501_));
  NOR3_X1    g11309(.A1(new_n11499_), .A2(new_n11203_), .A3(new_n10926_), .ZN(new_n11502_));
  AOI22_X1   g11310(.A1(new_n11501_), .A2(new_n10926_), .B1(\asqrt[22] ), .B2(new_n11502_), .ZN(new_n11503_));
  INV_X1     g11311(.I(new_n11503_), .ZN(new_n11504_));
  NOR3_X1    g11312(.A1(new_n11491_), .A2(\asqrt[37] ), .A3(new_n11461_), .ZN(new_n11505_));
  OAI21_X1   g11313(.A1(new_n11460_), .A2(new_n11505_), .B(new_n11492_), .ZN(new_n11506_));
  AOI21_X1   g11314(.A1(new_n11506_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n11507_));
  AOI21_X1   g11315(.A1(new_n11507_), .A2(new_n11494_), .B(new_n11478_), .ZN(new_n11508_));
  OAI21_X1   g11316(.A1(new_n11508_), .A2(new_n11495_), .B(\asqrt[40] ), .ZN(new_n11509_));
  NAND2_X1   g11317(.A1(new_n11509_), .A2(new_n3782_), .ZN(new_n11510_));
  OAI21_X1   g11318(.A1(new_n11510_), .A2(new_n11497_), .B(new_n11504_), .ZN(new_n11511_));
  AOI21_X1   g11319(.A1(new_n11511_), .A2(new_n11498_), .B(new_n3419_), .ZN(new_n11512_));
  INV_X1     g11320(.I(new_n10933_), .ZN(new_n11513_));
  NOR3_X1    g11321(.A1(new_n10929_), .A2(new_n11212_), .A3(new_n11513_), .ZN(new_n11514_));
  NOR3_X1    g11322(.A1(new_n11326_), .A2(new_n10929_), .A3(new_n11212_), .ZN(new_n11515_));
  INV_X1     g11323(.I(new_n11515_), .ZN(new_n11516_));
  AOI22_X1   g11324(.A1(new_n11516_), .A2(new_n11513_), .B1(\asqrt[22] ), .B2(new_n11514_), .ZN(new_n11517_));
  NOR3_X1    g11325(.A1(new_n11508_), .A2(\asqrt[40] ), .A3(new_n11495_), .ZN(new_n11518_));
  OAI21_X1   g11326(.A1(new_n11486_), .A2(new_n11518_), .B(new_n11509_), .ZN(new_n11519_));
  AOI21_X1   g11327(.A1(new_n11519_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n11520_));
  AOI21_X1   g11328(.A1(new_n11520_), .A2(new_n11511_), .B(new_n11517_), .ZN(new_n11521_));
  OAI21_X1   g11329(.A1(new_n11521_), .A2(new_n11512_), .B(\asqrt[43] ), .ZN(new_n11522_));
  INV_X1     g11330(.I(new_n11522_), .ZN(new_n11523_));
  NOR3_X1    g11331(.A1(new_n11326_), .A2(new_n10938_), .A3(new_n10944_), .ZN(new_n11524_));
  INV_X1     g11332(.I(new_n11524_), .ZN(new_n11525_));
  NOR3_X1    g11333(.A1(new_n10938_), .A2(new_n11148_), .A3(new_n10944_), .ZN(new_n11526_));
  AOI22_X1   g11334(.A1(new_n11525_), .A2(new_n11148_), .B1(\asqrt[22] ), .B2(new_n11526_), .ZN(new_n11527_));
  NOR3_X1    g11335(.A1(new_n11521_), .A2(\asqrt[43] ), .A3(new_n11512_), .ZN(new_n11528_));
  NOR2_X1    g11336(.A1(new_n11528_), .A2(new_n11527_), .ZN(new_n11529_));
  OAI21_X1   g11337(.A1(new_n11529_), .A2(new_n11523_), .B(\asqrt[44] ), .ZN(new_n11530_));
  NOR2_X1    g11338(.A1(new_n10945_), .A2(new_n10953_), .ZN(new_n11531_));
  NOR3_X1    g11339(.A1(new_n11531_), .A2(new_n11211_), .A3(new_n10952_), .ZN(new_n11532_));
  NOR3_X1    g11340(.A1(new_n11326_), .A2(new_n11211_), .A3(new_n11531_), .ZN(new_n11533_));
  INV_X1     g11341(.I(new_n11533_), .ZN(new_n11534_));
  AOI22_X1   g11342(.A1(new_n11534_), .A2(new_n10952_), .B1(\asqrt[22] ), .B2(new_n11532_), .ZN(new_n11535_));
  INV_X1     g11343(.I(new_n11535_), .ZN(new_n11536_));
  NAND2_X1   g11344(.A1(new_n11522_), .A2(new_n2954_), .ZN(new_n11537_));
  OAI21_X1   g11345(.A1(new_n11529_), .A2(new_n11537_), .B(new_n11536_), .ZN(new_n11538_));
  AOI21_X1   g11346(.A1(new_n11538_), .A2(new_n11530_), .B(new_n2641_), .ZN(new_n11539_));
  INV_X1     g11347(.I(new_n10959_), .ZN(new_n11540_));
  NOR3_X1    g11348(.A1(new_n11326_), .A2(new_n10955_), .A3(new_n11220_), .ZN(new_n11541_));
  INV_X1     g11349(.I(new_n11541_), .ZN(new_n11542_));
  NOR3_X1    g11350(.A1(new_n10955_), .A2(new_n11220_), .A3(new_n11540_), .ZN(new_n11543_));
  AOI22_X1   g11351(.A1(new_n11542_), .A2(new_n11540_), .B1(\asqrt[22] ), .B2(new_n11543_), .ZN(new_n11544_));
  OAI21_X1   g11352(.A1(new_n11527_), .A2(new_n11528_), .B(new_n11522_), .ZN(new_n11545_));
  AOI21_X1   g11353(.A1(new_n11545_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n11546_));
  AOI21_X1   g11354(.A1(new_n11546_), .A2(new_n11538_), .B(new_n11544_), .ZN(new_n11547_));
  OAI21_X1   g11355(.A1(new_n11547_), .A2(new_n11539_), .B(\asqrt[46] ), .ZN(new_n11548_));
  INV_X1     g11356(.I(new_n11548_), .ZN(new_n11549_));
  NOR3_X1    g11357(.A1(new_n10964_), .A2(new_n11147_), .A3(new_n10970_), .ZN(new_n11550_));
  NOR3_X1    g11358(.A1(new_n11326_), .A2(new_n10964_), .A3(new_n10970_), .ZN(new_n11551_));
  INV_X1     g11359(.I(new_n11551_), .ZN(new_n11552_));
  AOI22_X1   g11360(.A1(new_n11552_), .A2(new_n11147_), .B1(\asqrt[22] ), .B2(new_n11550_), .ZN(new_n11553_));
  NOR3_X1    g11361(.A1(new_n11547_), .A2(new_n11539_), .A3(\asqrt[46] ), .ZN(new_n11554_));
  NOR2_X1    g11362(.A1(new_n11554_), .A2(new_n11553_), .ZN(new_n11555_));
  OAI21_X1   g11363(.A1(new_n11555_), .A2(new_n11549_), .B(\asqrt[47] ), .ZN(new_n11556_));
  NOR2_X1    g11364(.A1(new_n10971_), .A2(new_n10979_), .ZN(new_n11557_));
  NOR3_X1    g11365(.A1(new_n11326_), .A2(new_n11219_), .A3(new_n11557_), .ZN(new_n11558_));
  INV_X1     g11366(.I(new_n11558_), .ZN(new_n11559_));
  NOR3_X1    g11367(.A1(new_n11557_), .A2(new_n11219_), .A3(new_n10978_), .ZN(new_n11560_));
  AOI22_X1   g11368(.A1(new_n11559_), .A2(new_n10978_), .B1(\asqrt[22] ), .B2(new_n11560_), .ZN(new_n11561_));
  INV_X1     g11369(.I(new_n11561_), .ZN(new_n11562_));
  NAND2_X1   g11370(.A1(new_n11548_), .A2(new_n2229_), .ZN(new_n11563_));
  OAI21_X1   g11371(.A1(new_n11555_), .A2(new_n11563_), .B(new_n11562_), .ZN(new_n11564_));
  AOI21_X1   g11372(.A1(new_n11564_), .A2(new_n11556_), .B(new_n1956_), .ZN(new_n11565_));
  INV_X1     g11373(.I(new_n10985_), .ZN(new_n11566_));
  NOR3_X1    g11374(.A1(new_n10981_), .A2(new_n11228_), .A3(new_n11566_), .ZN(new_n11567_));
  NOR3_X1    g11375(.A1(new_n11326_), .A2(new_n10981_), .A3(new_n11228_), .ZN(new_n11568_));
  INV_X1     g11376(.I(new_n11568_), .ZN(new_n11569_));
  AOI22_X1   g11377(.A1(new_n11569_), .A2(new_n11566_), .B1(\asqrt[22] ), .B2(new_n11567_), .ZN(new_n11570_));
  OAI21_X1   g11378(.A1(new_n11553_), .A2(new_n11554_), .B(new_n11548_), .ZN(new_n11571_));
  AOI21_X1   g11379(.A1(new_n11571_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n11572_));
  AOI21_X1   g11380(.A1(new_n11572_), .A2(new_n11564_), .B(new_n11570_), .ZN(new_n11573_));
  OAI21_X1   g11381(.A1(new_n11573_), .A2(new_n11565_), .B(\asqrt[49] ), .ZN(new_n11574_));
  INV_X1     g11382(.I(new_n11574_), .ZN(new_n11575_));
  NOR3_X1    g11383(.A1(new_n11326_), .A2(new_n10990_), .A3(new_n10996_), .ZN(new_n11576_));
  INV_X1     g11384(.I(new_n11576_), .ZN(new_n11577_));
  NOR3_X1    g11385(.A1(new_n10990_), .A2(new_n11146_), .A3(new_n10996_), .ZN(new_n11578_));
  AOI22_X1   g11386(.A1(new_n11577_), .A2(new_n11146_), .B1(\asqrt[22] ), .B2(new_n11578_), .ZN(new_n11579_));
  NOR3_X1    g11387(.A1(new_n11573_), .A2(new_n11565_), .A3(\asqrt[49] ), .ZN(new_n11580_));
  NOR2_X1    g11388(.A1(new_n11580_), .A2(new_n11579_), .ZN(new_n11581_));
  OAI21_X1   g11389(.A1(new_n11581_), .A2(new_n11575_), .B(\asqrt[50] ), .ZN(new_n11582_));
  NOR2_X1    g11390(.A1(new_n10997_), .A2(new_n11005_), .ZN(new_n11583_));
  NOR3_X1    g11391(.A1(new_n11583_), .A2(new_n11227_), .A3(new_n11004_), .ZN(new_n11584_));
  NOR3_X1    g11392(.A1(new_n11326_), .A2(new_n11227_), .A3(new_n11583_), .ZN(new_n11585_));
  INV_X1     g11393(.I(new_n11585_), .ZN(new_n11586_));
  AOI22_X1   g11394(.A1(new_n11586_), .A2(new_n11004_), .B1(\asqrt[22] ), .B2(new_n11584_), .ZN(new_n11587_));
  INV_X1     g11395(.I(new_n11587_), .ZN(new_n11588_));
  NAND2_X1   g11396(.A1(new_n11574_), .A2(new_n1612_), .ZN(new_n11589_));
  OAI21_X1   g11397(.A1(new_n11581_), .A2(new_n11589_), .B(new_n11588_), .ZN(new_n11590_));
  AOI21_X1   g11398(.A1(new_n11590_), .A2(new_n11582_), .B(new_n1376_), .ZN(new_n11591_));
  INV_X1     g11399(.I(new_n11011_), .ZN(new_n11592_));
  NOR3_X1    g11400(.A1(new_n11326_), .A2(new_n11007_), .A3(new_n11236_), .ZN(new_n11593_));
  INV_X1     g11401(.I(new_n11593_), .ZN(new_n11594_));
  NOR3_X1    g11402(.A1(new_n11007_), .A2(new_n11236_), .A3(new_n11592_), .ZN(new_n11595_));
  AOI22_X1   g11403(.A1(new_n11594_), .A2(new_n11592_), .B1(\asqrt[22] ), .B2(new_n11595_), .ZN(new_n11596_));
  OAI21_X1   g11404(.A1(new_n11579_), .A2(new_n11580_), .B(new_n11574_), .ZN(new_n11597_));
  AOI21_X1   g11405(.A1(new_n11597_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n11598_));
  AOI21_X1   g11406(.A1(new_n11598_), .A2(new_n11590_), .B(new_n11596_), .ZN(new_n11599_));
  OAI21_X1   g11407(.A1(new_n11599_), .A2(new_n11591_), .B(\asqrt[52] ), .ZN(new_n11600_));
  INV_X1     g11408(.I(new_n11600_), .ZN(new_n11601_));
  INV_X1     g11409(.I(new_n11599_), .ZN(new_n11602_));
  NOR3_X1    g11410(.A1(new_n11016_), .A2(new_n11145_), .A3(new_n11022_), .ZN(new_n11603_));
  NOR3_X1    g11411(.A1(new_n11326_), .A2(new_n11016_), .A3(new_n11022_), .ZN(new_n11604_));
  INV_X1     g11412(.I(new_n11604_), .ZN(new_n11605_));
  AOI22_X1   g11413(.A1(new_n11605_), .A2(new_n11145_), .B1(\asqrt[22] ), .B2(new_n11603_), .ZN(new_n11606_));
  NOR2_X1    g11414(.A1(new_n11591_), .A2(\asqrt[52] ), .ZN(new_n11607_));
  AOI21_X1   g11415(.A1(new_n11602_), .A2(new_n11607_), .B(new_n11606_), .ZN(new_n11608_));
  OAI21_X1   g11416(.A1(new_n11608_), .A2(new_n11601_), .B(\asqrt[53] ), .ZN(new_n11609_));
  NOR2_X1    g11417(.A1(new_n11023_), .A2(new_n11033_), .ZN(new_n11610_));
  NOR3_X1    g11418(.A1(new_n11326_), .A2(new_n11235_), .A3(new_n11610_), .ZN(new_n11611_));
  INV_X1     g11419(.I(new_n11611_), .ZN(new_n11612_));
  NOR3_X1    g11420(.A1(new_n11610_), .A2(new_n11235_), .A3(new_n11032_), .ZN(new_n11613_));
  AOI22_X1   g11421(.A1(new_n11612_), .A2(new_n11032_), .B1(\asqrt[22] ), .B2(new_n11613_), .ZN(new_n11614_));
  INV_X1     g11422(.I(new_n11614_), .ZN(new_n11615_));
  NAND2_X1   g11423(.A1(new_n11600_), .A2(new_n1103_), .ZN(new_n11616_));
  OAI21_X1   g11424(.A1(new_n11616_), .A2(new_n11608_), .B(new_n11615_), .ZN(new_n11617_));
  AOI21_X1   g11425(.A1(new_n11617_), .A2(new_n11609_), .B(new_n904_), .ZN(new_n11618_));
  INV_X1     g11426(.I(new_n11618_), .ZN(new_n11619_));
  INV_X1     g11427(.I(new_n11617_), .ZN(new_n11620_));
  INV_X1     g11428(.I(new_n11039_), .ZN(new_n11621_));
  NOR3_X1    g11429(.A1(new_n11035_), .A2(new_n11244_), .A3(new_n11621_), .ZN(new_n11622_));
  NOR3_X1    g11430(.A1(new_n11326_), .A2(new_n11035_), .A3(new_n11244_), .ZN(new_n11623_));
  INV_X1     g11431(.I(new_n11623_), .ZN(new_n11624_));
  AOI22_X1   g11432(.A1(new_n11624_), .A2(new_n11621_), .B1(\asqrt[22] ), .B2(new_n11622_), .ZN(new_n11625_));
  INV_X1     g11433(.I(new_n11625_), .ZN(new_n11626_));
  NAND2_X1   g11434(.A1(new_n11609_), .A2(new_n904_), .ZN(new_n11627_));
  OAI21_X1   g11435(.A1(new_n11627_), .A2(new_n11620_), .B(new_n11626_), .ZN(new_n11628_));
  AOI21_X1   g11436(.A1(new_n11628_), .A2(new_n11619_), .B(new_n823_), .ZN(new_n11629_));
  NOR3_X1    g11437(.A1(new_n11326_), .A2(new_n11044_), .A3(new_n11051_), .ZN(new_n11630_));
  INV_X1     g11438(.I(new_n11630_), .ZN(new_n11631_));
  NOR3_X1    g11439(.A1(new_n11044_), .A2(new_n11144_), .A3(new_n11051_), .ZN(new_n11632_));
  AOI22_X1   g11440(.A1(new_n11631_), .A2(new_n11144_), .B1(\asqrt[22] ), .B2(new_n11632_), .ZN(new_n11633_));
  NOR2_X1    g11441(.A1(new_n11618_), .A2(\asqrt[55] ), .ZN(new_n11634_));
  AOI21_X1   g11442(.A1(new_n11634_), .A2(new_n11628_), .B(new_n11633_), .ZN(new_n11635_));
  OAI21_X1   g11443(.A1(new_n11635_), .A2(new_n11629_), .B(\asqrt[56] ), .ZN(new_n11636_));
  NOR2_X1    g11444(.A1(new_n11052_), .A2(new_n11064_), .ZN(new_n11637_));
  NOR3_X1    g11445(.A1(new_n11637_), .A2(new_n11243_), .A3(new_n11063_), .ZN(new_n11638_));
  NOR3_X1    g11446(.A1(new_n11326_), .A2(new_n11243_), .A3(new_n11637_), .ZN(new_n11639_));
  INV_X1     g11447(.I(new_n11639_), .ZN(new_n11640_));
  AOI22_X1   g11448(.A1(new_n11640_), .A2(new_n11063_), .B1(\asqrt[22] ), .B2(new_n11638_), .ZN(new_n11641_));
  INV_X1     g11449(.I(new_n11641_), .ZN(new_n11642_));
  NOR3_X1    g11450(.A1(new_n11599_), .A2(new_n11591_), .A3(\asqrt[52] ), .ZN(new_n11643_));
  OAI21_X1   g11451(.A1(new_n11606_), .A2(new_n11643_), .B(new_n11600_), .ZN(new_n11644_));
  AOI21_X1   g11452(.A1(new_n11644_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n11645_));
  AOI21_X1   g11453(.A1(new_n11645_), .A2(new_n11617_), .B(new_n11625_), .ZN(new_n11646_));
  OAI21_X1   g11454(.A1(new_n11646_), .A2(new_n11618_), .B(\asqrt[55] ), .ZN(new_n11647_));
  NAND2_X1   g11455(.A1(new_n11647_), .A2(new_n703_), .ZN(new_n11648_));
  OAI21_X1   g11456(.A1(new_n11648_), .A2(new_n11635_), .B(new_n11642_), .ZN(new_n11649_));
  AOI21_X1   g11457(.A1(new_n11649_), .A2(new_n11636_), .B(new_n531_), .ZN(new_n11650_));
  INV_X1     g11458(.I(new_n11650_), .ZN(new_n11651_));
  INV_X1     g11459(.I(new_n11649_), .ZN(new_n11652_));
  INV_X1     g11460(.I(new_n11070_), .ZN(new_n11653_));
  NOR3_X1    g11461(.A1(new_n11326_), .A2(new_n11066_), .A3(new_n11252_), .ZN(new_n11654_));
  INV_X1     g11462(.I(new_n11654_), .ZN(new_n11655_));
  NOR3_X1    g11463(.A1(new_n11066_), .A2(new_n11252_), .A3(new_n11653_), .ZN(new_n11656_));
  AOI22_X1   g11464(.A1(new_n11655_), .A2(new_n11653_), .B1(\asqrt[22] ), .B2(new_n11656_), .ZN(new_n11657_));
  INV_X1     g11465(.I(new_n11657_), .ZN(new_n11658_));
  NAND2_X1   g11466(.A1(new_n11636_), .A2(new_n531_), .ZN(new_n11659_));
  OAI21_X1   g11467(.A1(new_n11659_), .A2(new_n11652_), .B(new_n11658_), .ZN(new_n11660_));
  AOI21_X1   g11468(.A1(new_n11660_), .A2(new_n11651_), .B(new_n436_), .ZN(new_n11661_));
  NOR3_X1    g11469(.A1(new_n11075_), .A2(new_n11143_), .A3(new_n11082_), .ZN(new_n11662_));
  NOR3_X1    g11470(.A1(new_n11326_), .A2(new_n11075_), .A3(new_n11082_), .ZN(new_n11663_));
  INV_X1     g11471(.I(new_n11663_), .ZN(new_n11664_));
  AOI22_X1   g11472(.A1(new_n11664_), .A2(new_n11143_), .B1(\asqrt[22] ), .B2(new_n11662_), .ZN(new_n11665_));
  NOR2_X1    g11473(.A1(new_n11650_), .A2(\asqrt[58] ), .ZN(new_n11666_));
  AOI21_X1   g11474(.A1(new_n11666_), .A2(new_n11660_), .B(new_n11665_), .ZN(new_n11667_));
  OAI21_X1   g11475(.A1(new_n11667_), .A2(new_n11661_), .B(\asqrt[59] ), .ZN(new_n11668_));
  NOR2_X1    g11476(.A1(new_n11083_), .A2(new_n11094_), .ZN(new_n11669_));
  NOR3_X1    g11477(.A1(new_n11326_), .A2(new_n11251_), .A3(new_n11669_), .ZN(new_n11670_));
  INV_X1     g11478(.I(new_n11670_), .ZN(new_n11671_));
  NOR3_X1    g11479(.A1(new_n11669_), .A2(new_n11251_), .A3(new_n11093_), .ZN(new_n11672_));
  AOI22_X1   g11480(.A1(new_n11671_), .A2(new_n11093_), .B1(\asqrt[22] ), .B2(new_n11672_), .ZN(new_n11673_));
  INV_X1     g11481(.I(new_n11673_), .ZN(new_n11674_));
  NOR3_X1    g11482(.A1(new_n11646_), .A2(\asqrt[55] ), .A3(new_n11618_), .ZN(new_n11675_));
  OAI21_X1   g11483(.A1(new_n11633_), .A2(new_n11675_), .B(new_n11647_), .ZN(new_n11676_));
  AOI21_X1   g11484(.A1(new_n11676_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n11677_));
  AOI21_X1   g11485(.A1(new_n11677_), .A2(new_n11649_), .B(new_n11657_), .ZN(new_n11678_));
  OAI21_X1   g11486(.A1(new_n11678_), .A2(new_n11650_), .B(\asqrt[58] ), .ZN(new_n11679_));
  NAND2_X1   g11487(.A1(new_n11679_), .A2(new_n327_), .ZN(new_n11680_));
  OAI21_X1   g11488(.A1(new_n11680_), .A2(new_n11667_), .B(new_n11674_), .ZN(new_n11681_));
  AOI21_X1   g11489(.A1(new_n11681_), .A2(new_n11668_), .B(new_n306_), .ZN(new_n11682_));
  INV_X1     g11490(.I(new_n11682_), .ZN(new_n11683_));
  INV_X1     g11491(.I(new_n11681_), .ZN(new_n11684_));
  INV_X1     g11492(.I(new_n11100_), .ZN(new_n11685_));
  NOR3_X1    g11493(.A1(new_n11096_), .A2(new_n11259_), .A3(new_n11685_), .ZN(new_n11686_));
  NOR3_X1    g11494(.A1(new_n11326_), .A2(new_n11096_), .A3(new_n11259_), .ZN(new_n11687_));
  INV_X1     g11495(.I(new_n11687_), .ZN(new_n11688_));
  AOI22_X1   g11496(.A1(new_n11688_), .A2(new_n11685_), .B1(\asqrt[22] ), .B2(new_n11686_), .ZN(new_n11689_));
  INV_X1     g11497(.I(new_n11689_), .ZN(new_n11690_));
  NAND2_X1   g11498(.A1(new_n11668_), .A2(new_n306_), .ZN(new_n11691_));
  OAI21_X1   g11499(.A1(new_n11684_), .A2(new_n11691_), .B(new_n11690_), .ZN(new_n11692_));
  AOI21_X1   g11500(.A1(new_n11692_), .A2(new_n11683_), .B(new_n218_), .ZN(new_n11693_));
  NOR3_X1    g11501(.A1(new_n11326_), .A2(new_n11105_), .A3(new_n11111_), .ZN(new_n11694_));
  INV_X1     g11502(.I(new_n11694_), .ZN(new_n11695_));
  NOR3_X1    g11503(.A1(new_n11105_), .A2(new_n11142_), .A3(new_n11111_), .ZN(new_n11696_));
  AOI22_X1   g11504(.A1(new_n11695_), .A2(new_n11142_), .B1(\asqrt[22] ), .B2(new_n11696_), .ZN(new_n11697_));
  NOR2_X1    g11505(.A1(new_n11682_), .A2(\asqrt[61] ), .ZN(new_n11698_));
  AOI21_X1   g11506(.A1(new_n11698_), .A2(new_n11692_), .B(new_n11697_), .ZN(new_n11699_));
  OAI21_X1   g11507(.A1(new_n11699_), .A2(new_n11693_), .B(\asqrt[62] ), .ZN(new_n11700_));
  NOR2_X1    g11508(.A1(new_n11112_), .A2(new_n11119_), .ZN(new_n11701_));
  NOR3_X1    g11509(.A1(new_n11701_), .A2(new_n11281_), .A3(new_n11118_), .ZN(new_n11702_));
  NOR3_X1    g11510(.A1(new_n11326_), .A2(new_n11281_), .A3(new_n11701_), .ZN(new_n11703_));
  INV_X1     g11511(.I(new_n11703_), .ZN(new_n11704_));
  AOI22_X1   g11512(.A1(new_n11704_), .A2(new_n11118_), .B1(\asqrt[22] ), .B2(new_n11702_), .ZN(new_n11705_));
  INV_X1     g11513(.I(new_n11705_), .ZN(new_n11706_));
  NOR3_X1    g11514(.A1(new_n11678_), .A2(\asqrt[58] ), .A3(new_n11650_), .ZN(new_n11707_));
  OAI21_X1   g11515(.A1(new_n11665_), .A2(new_n11707_), .B(new_n11679_), .ZN(new_n11708_));
  AOI21_X1   g11516(.A1(new_n11708_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n11709_));
  AOI21_X1   g11517(.A1(new_n11709_), .A2(new_n11681_), .B(new_n11689_), .ZN(new_n11710_));
  OAI21_X1   g11518(.A1(new_n11710_), .A2(new_n11682_), .B(\asqrt[61] ), .ZN(new_n11711_));
  NAND2_X1   g11519(.A1(new_n11711_), .A2(new_n207_), .ZN(new_n11712_));
  OAI21_X1   g11520(.A1(new_n11712_), .A2(new_n11699_), .B(new_n11706_), .ZN(new_n11713_));
  INV_X1     g11521(.I(new_n11283_), .ZN(new_n11714_));
  NAND4_X1   g11522(.A1(\asqrt[22] ), .A2(new_n11282_), .A3(new_n11125_), .A4(new_n11714_), .ZN(new_n11715_));
  NAND2_X1   g11523(.A1(new_n11714_), .A2(new_n11282_), .ZN(new_n11716_));
  OAI21_X1   g11524(.A1(new_n11326_), .A2(new_n11716_), .B(new_n11263_), .ZN(new_n11717_));
  NAND2_X1   g11525(.A1(new_n11717_), .A2(new_n11715_), .ZN(new_n11718_));
  INV_X1     g11526(.I(new_n11302_), .ZN(new_n11719_));
  AOI21_X1   g11527(.A1(new_n11265_), .A2(new_n11282_), .B(new_n11136_), .ZN(new_n11720_));
  AOI21_X1   g11528(.A1(\asqrt[22] ), .A2(new_n11720_), .B(new_n11719_), .ZN(new_n11721_));
  NAND2_X1   g11529(.A1(new_n11718_), .A2(new_n11721_), .ZN(new_n11722_));
  AOI21_X1   g11530(.A1(new_n11713_), .A2(new_n11700_), .B(new_n11722_), .ZN(new_n11723_));
  NOR2_X1    g11531(.A1(new_n11723_), .A2(\asqrt[63] ), .ZN(new_n11724_));
  INV_X1     g11532(.I(new_n11713_), .ZN(new_n11725_));
  INV_X1     g11533(.I(new_n11718_), .ZN(new_n11726_));
  NAND2_X1   g11534(.A1(new_n11700_), .A2(new_n11726_), .ZN(new_n11727_));
  AOI21_X1   g11535(.A1(\asqrt[22] ), .A2(new_n11137_), .B(new_n11284_), .ZN(new_n11728_));
  OR3_X2     g11536(.A1(new_n11728_), .A2(new_n193_), .A3(new_n11720_), .Z(new_n11729_));
  OAI21_X1   g11537(.A1(new_n10759_), .A2(new_n11271_), .B(new_n11132_), .ZN(new_n11730_));
  NOR4_X1    g11538(.A1(new_n11719_), .A2(new_n11135_), .A3(new_n11269_), .A4(new_n11730_), .ZN(new_n11731_));
  NAND2_X1   g11539(.A1(new_n11731_), .A2(new_n11141_), .ZN(new_n11732_));
  NAND2_X1   g11540(.A1(new_n11729_), .A2(new_n11732_), .ZN(new_n11733_));
  INV_X1     g11541(.I(new_n11733_), .ZN(new_n11734_));
  OAI21_X1   g11542(.A1(new_n11725_), .A2(new_n11727_), .B(new_n11734_), .ZN(new_n11735_));
  NOR2_X1    g11543(.A1(new_n11724_), .A2(new_n11735_), .ZN(new_n11736_));
  INV_X1     g11544(.I(\a[42] ), .ZN(new_n11737_));
  NOR2_X1    g11545(.A1(\a[40] ), .A2(\a[41] ), .ZN(new_n11738_));
  INV_X1     g11546(.I(new_n11738_), .ZN(new_n11739_));
  NOR2_X1    g11547(.A1(new_n11739_), .A2(\a[42] ), .ZN(new_n11740_));
  INV_X1     g11548(.I(new_n11740_), .ZN(new_n11741_));
  OAI21_X1   g11549(.A1(new_n11736_), .A2(new_n11737_), .B(new_n11741_), .ZN(new_n11742_));
  NOR3_X1    g11550(.A1(new_n11269_), .A2(new_n11272_), .A3(new_n11740_), .ZN(new_n11743_));
  NAND3_X1   g11551(.A1(new_n11141_), .A2(new_n11302_), .A3(new_n11743_), .ZN(new_n11744_));
  INV_X1     g11552(.I(new_n11744_), .ZN(new_n11745_));
  OAI21_X1   g11553(.A1(new_n11736_), .A2(new_n11737_), .B(new_n11745_), .ZN(new_n11746_));
  NOR3_X1    g11554(.A1(new_n11710_), .A2(\asqrt[61] ), .A3(new_n11682_), .ZN(new_n11747_));
  OAI21_X1   g11555(.A1(new_n11697_), .A2(new_n11747_), .B(new_n11711_), .ZN(new_n11748_));
  INV_X1     g11556(.I(new_n11697_), .ZN(new_n11749_));
  INV_X1     g11557(.I(new_n11665_), .ZN(new_n11750_));
  INV_X1     g11558(.I(new_n11633_), .ZN(new_n11751_));
  INV_X1     g11559(.I(new_n11606_), .ZN(new_n11752_));
  INV_X1     g11560(.I(new_n11579_), .ZN(new_n11753_));
  INV_X1     g11561(.I(new_n11553_), .ZN(new_n11754_));
  INV_X1     g11562(.I(new_n11527_), .ZN(new_n11755_));
  INV_X1     g11563(.I(new_n11498_), .ZN(new_n11756_));
  NOR3_X1    g11564(.A1(new_n11497_), .A2(new_n11482_), .A3(\asqrt[41] ), .ZN(new_n11757_));
  NOR2_X1    g11565(.A1(new_n11757_), .A2(new_n11503_), .ZN(new_n11758_));
  OAI21_X1   g11566(.A1(new_n11758_), .A2(new_n11756_), .B(\asqrt[42] ), .ZN(new_n11759_));
  NAND2_X1   g11567(.A1(new_n11759_), .A2(new_n3218_), .ZN(new_n11760_));
  OAI21_X1   g11568(.A1(new_n11760_), .A2(new_n11521_), .B(new_n11755_), .ZN(new_n11761_));
  NAND3_X1   g11569(.A1(new_n11761_), .A2(new_n2954_), .A3(new_n11522_), .ZN(new_n11762_));
  AOI22_X1   g11570(.A1(new_n11762_), .A2(new_n11536_), .B1(\asqrt[44] ), .B2(new_n11545_), .ZN(new_n11763_));
  OAI21_X1   g11571(.A1(new_n11763_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n11764_));
  OAI21_X1   g11572(.A1(new_n11764_), .A2(new_n11547_), .B(new_n11754_), .ZN(new_n11765_));
  NAND3_X1   g11573(.A1(new_n11765_), .A2(new_n2229_), .A3(new_n11548_), .ZN(new_n11766_));
  AOI22_X1   g11574(.A1(new_n11766_), .A2(new_n11562_), .B1(\asqrt[47] ), .B2(new_n11571_), .ZN(new_n11767_));
  OAI21_X1   g11575(.A1(new_n11767_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n11768_));
  OAI21_X1   g11576(.A1(new_n11768_), .A2(new_n11573_), .B(new_n11753_), .ZN(new_n11769_));
  NAND3_X1   g11577(.A1(new_n11769_), .A2(new_n1612_), .A3(new_n11574_), .ZN(new_n11770_));
  AOI22_X1   g11578(.A1(new_n11770_), .A2(new_n11588_), .B1(\asqrt[50] ), .B2(new_n11597_), .ZN(new_n11771_));
  OAI21_X1   g11579(.A1(new_n11771_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n11772_));
  OAI21_X1   g11580(.A1(new_n11772_), .A2(new_n11599_), .B(new_n11752_), .ZN(new_n11773_));
  NAND3_X1   g11581(.A1(new_n11773_), .A2(new_n1103_), .A3(new_n11600_), .ZN(new_n11774_));
  AOI22_X1   g11582(.A1(new_n11774_), .A2(new_n11615_), .B1(\asqrt[53] ), .B2(new_n11644_), .ZN(new_n11775_));
  OAI21_X1   g11583(.A1(new_n11775_), .A2(new_n904_), .B(new_n823_), .ZN(new_n11776_));
  OAI21_X1   g11584(.A1(new_n11776_), .A2(new_n11646_), .B(new_n11751_), .ZN(new_n11777_));
  NAND3_X1   g11585(.A1(new_n11777_), .A2(new_n703_), .A3(new_n11647_), .ZN(new_n11778_));
  AOI22_X1   g11586(.A1(new_n11778_), .A2(new_n11642_), .B1(\asqrt[56] ), .B2(new_n11676_), .ZN(new_n11779_));
  OAI21_X1   g11587(.A1(new_n11779_), .A2(new_n531_), .B(new_n436_), .ZN(new_n11780_));
  OAI21_X1   g11588(.A1(new_n11780_), .A2(new_n11678_), .B(new_n11750_), .ZN(new_n11781_));
  NAND3_X1   g11589(.A1(new_n11781_), .A2(new_n327_), .A3(new_n11679_), .ZN(new_n11782_));
  AOI22_X1   g11590(.A1(new_n11782_), .A2(new_n11674_), .B1(new_n11708_), .B2(\asqrt[59] ), .ZN(new_n11783_));
  OAI21_X1   g11591(.A1(new_n11783_), .A2(new_n306_), .B(new_n218_), .ZN(new_n11784_));
  OAI21_X1   g11592(.A1(new_n11784_), .A2(new_n11710_), .B(new_n11749_), .ZN(new_n11785_));
  NAND3_X1   g11593(.A1(new_n11785_), .A2(new_n207_), .A3(new_n11711_), .ZN(new_n11786_));
  AOI22_X1   g11594(.A1(new_n11786_), .A2(new_n11706_), .B1(new_n11748_), .B2(\asqrt[62] ), .ZN(new_n11787_));
  OAI21_X1   g11595(.A1(new_n11787_), .A2(new_n11722_), .B(new_n193_), .ZN(new_n11788_));
  AOI21_X1   g11596(.A1(new_n11748_), .A2(\asqrt[62] ), .B(new_n11718_), .ZN(new_n11789_));
  AOI21_X1   g11597(.A1(new_n11789_), .A2(new_n11713_), .B(new_n11733_), .ZN(new_n11790_));
  AOI21_X1   g11598(.A1(new_n11788_), .A2(new_n11790_), .B(new_n11278_), .ZN(new_n11791_));
  OAI21_X1   g11599(.A1(new_n11724_), .A2(new_n11735_), .B(new_n11737_), .ZN(new_n11792_));
  AOI21_X1   g11600(.A1(\a[43] ), .A2(new_n11792_), .B(new_n11791_), .ZN(new_n11793_));
  AOI22_X1   g11601(.A1(new_n11793_), .A2(new_n11746_), .B1(\asqrt[22] ), .B2(new_n11742_), .ZN(new_n11794_));
  NOR2_X1    g11602(.A1(new_n11794_), .A2(new_n10812_), .ZN(new_n11795_));
  NAND2_X1   g11603(.A1(new_n11793_), .A2(new_n11746_), .ZN(new_n11796_));
  OAI21_X1   g11604(.A1(new_n11724_), .A2(new_n11735_), .B(new_n11277_), .ZN(new_n11797_));
  NAND2_X1   g11605(.A1(new_n11789_), .A2(new_n11713_), .ZN(new_n11798_));
  OAI21_X1   g11606(.A1(new_n11731_), .A2(new_n11275_), .B(new_n11141_), .ZN(new_n11799_));
  NAND4_X1   g11607(.A1(new_n11788_), .A2(new_n11798_), .A3(new_n11729_), .A4(new_n11799_), .ZN(new_n11800_));
  AOI21_X1   g11608(.A1(new_n11800_), .A2(new_n11797_), .B(new_n11290_), .ZN(new_n11801_));
  INV_X1     g11609(.I(new_n11798_), .ZN(new_n11802_));
  NAND2_X1   g11610(.A1(new_n11729_), .A2(new_n11799_), .ZN(new_n11803_));
  NOR3_X1    g11611(.A1(new_n11802_), .A2(new_n11724_), .A3(new_n11803_), .ZN(new_n11804_));
  NOR3_X1    g11612(.A1(new_n11804_), .A2(new_n11791_), .A3(\a[44] ), .ZN(new_n11805_));
  NOR2_X1    g11613(.A1(new_n11801_), .A2(new_n11805_), .ZN(new_n11806_));
  AOI21_X1   g11614(.A1(new_n11742_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n11807_));
  AOI21_X1   g11615(.A1(new_n11796_), .A2(new_n11807_), .B(new_n11806_), .ZN(new_n11808_));
  OAI21_X1   g11616(.A1(new_n11808_), .A2(new_n11795_), .B(\asqrt[24] ), .ZN(new_n11809_));
  OAI21_X1   g11617(.A1(\asqrt[63] ), .A2(new_n11723_), .B(new_n11790_), .ZN(\asqrt[21] ));
  NOR3_X1    g11618(.A1(new_n11370_), .A2(new_n11289_), .A3(new_n11295_), .ZN(new_n11811_));
  NAND3_X1   g11619(.A1(\asqrt[21] ), .A2(new_n11308_), .A3(new_n11355_), .ZN(new_n11812_));
  AOI22_X1   g11620(.A1(new_n11812_), .A2(new_n11370_), .B1(\asqrt[21] ), .B2(new_n11811_), .ZN(new_n11813_));
  INV_X1     g11621(.I(new_n11813_), .ZN(new_n11814_));
  OAI21_X1   g11622(.A1(new_n11794_), .A2(new_n10812_), .B(new_n10221_), .ZN(new_n11815_));
  OAI21_X1   g11623(.A1(new_n11815_), .A2(new_n11808_), .B(new_n11814_), .ZN(new_n11816_));
  AOI21_X1   g11624(.A1(new_n11816_), .A2(new_n11809_), .B(new_n9846_), .ZN(new_n11817_));
  NOR2_X1    g11625(.A1(new_n11307_), .A2(new_n11305_), .ZN(new_n11818_));
  NOR2_X1    g11626(.A1(new_n11299_), .A2(new_n11309_), .ZN(new_n11819_));
  INV_X1     g11627(.I(new_n11819_), .ZN(new_n11820_));
  NAND4_X1   g11628(.A1(\asqrt[21] ), .A2(new_n11300_), .A3(new_n11818_), .A4(new_n11820_), .ZN(new_n11821_));
  NOR3_X1    g11629(.A1(new_n11736_), .A2(new_n11359_), .A3(new_n11819_), .ZN(new_n11822_));
  OAI21_X1   g11630(.A1(new_n11822_), .A2(new_n11818_), .B(new_n11821_), .ZN(new_n11823_));
  INV_X1     g11631(.I(new_n11823_), .ZN(new_n11824_));
  AOI21_X1   g11632(.A1(new_n11788_), .A2(new_n11790_), .B(new_n11737_), .ZN(new_n11825_));
  OAI21_X1   g11633(.A1(new_n11825_), .A2(new_n11740_), .B(\asqrt[22] ), .ZN(new_n11826_));
  INV_X1     g11634(.I(new_n11826_), .ZN(new_n11827_));
  NOR2_X1    g11635(.A1(new_n11825_), .A2(new_n11744_), .ZN(new_n11828_));
  INV_X1     g11636(.I(\a[43] ), .ZN(new_n11829_));
  AOI21_X1   g11637(.A1(\asqrt[21] ), .A2(new_n11737_), .B(new_n11829_), .ZN(new_n11830_));
  NOR3_X1    g11638(.A1(new_n11828_), .A2(new_n11830_), .A3(new_n11791_), .ZN(new_n11831_));
  OAI21_X1   g11639(.A1(new_n11831_), .A2(new_n11827_), .B(\asqrt[23] ), .ZN(new_n11832_));
  AOI21_X1   g11640(.A1(\asqrt[21] ), .A2(\a[42] ), .B(new_n11740_), .ZN(new_n11833_));
  OAI21_X1   g11641(.A1(new_n11833_), .A2(new_n11326_), .B(new_n10812_), .ZN(new_n11834_));
  OAI22_X1   g11642(.A1(new_n11831_), .A2(new_n11834_), .B1(new_n11801_), .B2(new_n11805_), .ZN(new_n11835_));
  AOI21_X1   g11643(.A1(new_n11835_), .A2(new_n11832_), .B(new_n10221_), .ZN(new_n11836_));
  AOI21_X1   g11644(.A1(new_n11788_), .A2(new_n11790_), .B(\a[42] ), .ZN(new_n11837_));
  OAI21_X1   g11645(.A1(new_n11829_), .A2(new_n11837_), .B(new_n11797_), .ZN(new_n11838_));
  OAI21_X1   g11646(.A1(new_n11838_), .A2(new_n11828_), .B(new_n11826_), .ZN(new_n11839_));
  AOI21_X1   g11647(.A1(new_n11839_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n11840_));
  AOI21_X1   g11648(.A1(new_n11840_), .A2(new_n11835_), .B(new_n11813_), .ZN(new_n11841_));
  NOR3_X1    g11649(.A1(new_n11841_), .A2(new_n11836_), .A3(\asqrt[25] ), .ZN(new_n11842_));
  NOR2_X1    g11650(.A1(new_n11842_), .A2(new_n11824_), .ZN(new_n11843_));
  OAI21_X1   g11651(.A1(new_n11843_), .A2(new_n11817_), .B(\asqrt[26] ), .ZN(new_n11844_));
  NOR2_X1    g11652(.A1(new_n11372_), .A2(new_n11364_), .ZN(new_n11845_));
  NOR3_X1    g11653(.A1(new_n11736_), .A2(new_n11311_), .A3(new_n11845_), .ZN(new_n11846_));
  INV_X1     g11654(.I(new_n11846_), .ZN(new_n11847_));
  NOR3_X1    g11655(.A1(new_n11845_), .A2(new_n11311_), .A3(new_n11369_), .ZN(new_n11848_));
  AOI22_X1   g11656(.A1(new_n11847_), .A2(new_n11369_), .B1(\asqrt[21] ), .B2(new_n11848_), .ZN(new_n11849_));
  INV_X1     g11657(.I(new_n11849_), .ZN(new_n11850_));
  OAI21_X1   g11658(.A1(new_n11841_), .A2(new_n11836_), .B(\asqrt[25] ), .ZN(new_n11851_));
  NAND2_X1   g11659(.A1(new_n11851_), .A2(new_n9317_), .ZN(new_n11852_));
  OAI21_X1   g11660(.A1(new_n11843_), .A2(new_n11852_), .B(new_n11850_), .ZN(new_n11853_));
  AOI21_X1   g11661(.A1(new_n11853_), .A2(new_n11844_), .B(new_n8826_), .ZN(new_n11854_));
  NOR3_X1    g11662(.A1(new_n11321_), .A2(new_n11330_), .A3(new_n11328_), .ZN(new_n11855_));
  NOR3_X1    g11663(.A1(new_n11736_), .A2(new_n11321_), .A3(new_n11330_), .ZN(new_n11856_));
  INV_X1     g11664(.I(new_n11856_), .ZN(new_n11857_));
  AOI22_X1   g11665(.A1(new_n11857_), .A2(new_n11328_), .B1(\asqrt[21] ), .B2(new_n11855_), .ZN(new_n11858_));
  OAI21_X1   g11666(.A1(new_n11824_), .A2(new_n11842_), .B(new_n11851_), .ZN(new_n11859_));
  AOI21_X1   g11667(.A1(new_n11859_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n11860_));
  AOI21_X1   g11668(.A1(new_n11860_), .A2(new_n11853_), .B(new_n11858_), .ZN(new_n11861_));
  OAI21_X1   g11669(.A1(new_n11861_), .A2(new_n11854_), .B(\asqrt[28] ), .ZN(new_n11862_));
  INV_X1     g11670(.I(new_n11862_), .ZN(new_n11863_));
  NAND2_X1   g11671(.A1(new_n11375_), .A2(new_n11367_), .ZN(new_n11864_));
  NAND3_X1   g11672(.A1(\asqrt[21] ), .A2(new_n11332_), .A3(new_n11864_), .ZN(new_n11865_));
  AND3_X2    g11673(.A1(new_n11332_), .A2(new_n11337_), .A3(new_n11864_), .Z(new_n11866_));
  AOI22_X1   g11674(.A1(new_n11865_), .A2(new_n11338_), .B1(\asqrt[21] ), .B2(new_n11866_), .ZN(new_n11867_));
  NOR3_X1    g11675(.A1(new_n11861_), .A2(new_n11854_), .A3(\asqrt[28] ), .ZN(new_n11868_));
  NOR2_X1    g11676(.A1(new_n11868_), .A2(new_n11867_), .ZN(new_n11869_));
  OAI21_X1   g11677(.A1(new_n11869_), .A2(new_n11863_), .B(\asqrt[29] ), .ZN(new_n11870_));
  INV_X1     g11678(.I(new_n11345_), .ZN(new_n11871_));
  NOR3_X1    g11679(.A1(new_n11341_), .A2(new_n11434_), .A3(new_n11871_), .ZN(new_n11872_));
  NOR3_X1    g11680(.A1(new_n11736_), .A2(new_n11341_), .A3(new_n11434_), .ZN(new_n11873_));
  INV_X1     g11681(.I(new_n11873_), .ZN(new_n11874_));
  AOI22_X1   g11682(.A1(new_n11874_), .A2(new_n11871_), .B1(\asqrt[21] ), .B2(new_n11872_), .ZN(new_n11875_));
  INV_X1     g11683(.I(new_n11875_), .ZN(new_n11876_));
  NAND2_X1   g11684(.A1(new_n11862_), .A2(new_n8036_), .ZN(new_n11877_));
  OAI21_X1   g11685(.A1(new_n11869_), .A2(new_n11877_), .B(new_n11876_), .ZN(new_n11878_));
  AOI21_X1   g11686(.A1(new_n11878_), .A2(new_n11870_), .B(new_n7539_), .ZN(new_n11879_));
  INV_X1     g11687(.I(new_n11404_), .ZN(new_n11880_));
  NAND3_X1   g11688(.A1(\asqrt[21] ), .A2(new_n11349_), .A3(new_n11880_), .ZN(new_n11881_));
  AND3_X2    g11689(.A1(new_n11880_), .A2(new_n11349_), .A3(new_n11353_), .Z(new_n11882_));
  AOI22_X1   g11690(.A1(new_n11881_), .A2(new_n11354_), .B1(\asqrt[21] ), .B2(new_n11882_), .ZN(new_n11883_));
  OAI21_X1   g11691(.A1(new_n11867_), .A2(new_n11868_), .B(new_n11862_), .ZN(new_n11884_));
  AOI21_X1   g11692(.A1(new_n11884_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n11885_));
  AOI21_X1   g11693(.A1(new_n11885_), .A2(new_n11878_), .B(new_n11883_), .ZN(new_n11886_));
  OAI21_X1   g11694(.A1(new_n11886_), .A2(new_n11879_), .B(\asqrt[31] ), .ZN(new_n11887_));
  INV_X1     g11695(.I(new_n11887_), .ZN(new_n11888_));
  INV_X1     g11696(.I(new_n11388_), .ZN(new_n11889_));
  NOR3_X1    g11697(.A1(new_n11889_), .A2(new_n11380_), .A3(new_n11387_), .ZN(new_n11890_));
  NOR3_X1    g11698(.A1(new_n11736_), .A2(new_n11380_), .A3(new_n11889_), .ZN(new_n11891_));
  INV_X1     g11699(.I(new_n11891_), .ZN(new_n11892_));
  AOI22_X1   g11700(.A1(new_n11892_), .A2(new_n11387_), .B1(\asqrt[21] ), .B2(new_n11890_), .ZN(new_n11893_));
  NOR3_X1    g11701(.A1(new_n11886_), .A2(new_n11879_), .A3(\asqrt[31] ), .ZN(new_n11894_));
  NOR2_X1    g11702(.A1(new_n11894_), .A2(new_n11893_), .ZN(new_n11895_));
  OAI21_X1   g11703(.A1(new_n11895_), .A2(new_n11888_), .B(\asqrt[32] ), .ZN(new_n11896_));
  INV_X1     g11704(.I(new_n11394_), .ZN(new_n11897_));
  NOR3_X1    g11705(.A1(new_n11736_), .A2(new_n11390_), .A3(new_n11438_), .ZN(new_n11898_));
  INV_X1     g11706(.I(new_n11898_), .ZN(new_n11899_));
  NOR3_X1    g11707(.A1(new_n11390_), .A2(new_n11897_), .A3(new_n11438_), .ZN(new_n11900_));
  AOI22_X1   g11708(.A1(new_n11899_), .A2(new_n11897_), .B1(\asqrt[21] ), .B2(new_n11900_), .ZN(new_n11901_));
  INV_X1     g11709(.I(new_n11901_), .ZN(new_n11902_));
  NAND2_X1   g11710(.A1(new_n11887_), .A2(new_n6824_), .ZN(new_n11903_));
  OAI21_X1   g11711(.A1(new_n11895_), .A2(new_n11903_), .B(new_n11902_), .ZN(new_n11904_));
  AOI21_X1   g11712(.A1(new_n11904_), .A2(new_n11896_), .B(new_n6356_), .ZN(new_n11905_));
  OAI21_X1   g11713(.A1(new_n11407_), .A2(new_n11396_), .B(new_n11402_), .ZN(new_n11906_));
  AOI21_X1   g11714(.A1(\asqrt[32] ), .A2(new_n11439_), .B(new_n11906_), .ZN(new_n11907_));
  OAI21_X1   g11715(.A1(new_n11396_), .A2(new_n11407_), .B(new_n11397_), .ZN(new_n11908_));
  NOR2_X1    g11716(.A1(new_n11736_), .A2(new_n11908_), .ZN(new_n11909_));
  INV_X1     g11717(.I(new_n11909_), .ZN(new_n11910_));
  AOI22_X1   g11718(.A1(new_n11910_), .A2(new_n11403_), .B1(\asqrt[21] ), .B2(new_n11907_), .ZN(new_n11911_));
  OAI21_X1   g11719(.A1(new_n11893_), .A2(new_n11894_), .B(new_n11887_), .ZN(new_n11912_));
  AOI21_X1   g11720(.A1(new_n11912_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n11913_));
  AOI21_X1   g11721(.A1(new_n11913_), .A2(new_n11904_), .B(new_n11911_), .ZN(new_n11914_));
  OAI21_X1   g11722(.A1(new_n11914_), .A2(new_n11905_), .B(\asqrt[34] ), .ZN(new_n11915_));
  INV_X1     g11723(.I(new_n11915_), .ZN(new_n11916_));
  NOR2_X1    g11724(.A1(new_n11411_), .A2(new_n11418_), .ZN(new_n11917_));
  NOR3_X1    g11725(.A1(new_n11736_), .A2(new_n11409_), .A3(new_n11917_), .ZN(new_n11918_));
  INV_X1     g11726(.I(new_n11918_), .ZN(new_n11919_));
  NOR3_X1    g11727(.A1(new_n11917_), .A2(new_n11409_), .A3(new_n11417_), .ZN(new_n11920_));
  AOI22_X1   g11728(.A1(new_n11919_), .A2(new_n11417_), .B1(\asqrt[21] ), .B2(new_n11920_), .ZN(new_n11921_));
  NOR3_X1    g11729(.A1(new_n11914_), .A2(new_n11905_), .A3(\asqrt[34] ), .ZN(new_n11922_));
  NOR2_X1    g11730(.A1(new_n11922_), .A2(new_n11921_), .ZN(new_n11923_));
  OAI21_X1   g11731(.A1(new_n11923_), .A2(new_n11916_), .B(\asqrt[35] ), .ZN(new_n11924_));
  INV_X1     g11732(.I(new_n11424_), .ZN(new_n11925_));
  NOR3_X1    g11733(.A1(new_n11420_), .A2(new_n11925_), .A3(new_n11488_), .ZN(new_n11926_));
  NOR3_X1    g11734(.A1(new_n11736_), .A2(new_n11420_), .A3(new_n11488_), .ZN(new_n11927_));
  INV_X1     g11735(.I(new_n11927_), .ZN(new_n11928_));
  AOI22_X1   g11736(.A1(new_n11928_), .A2(new_n11925_), .B1(\asqrt[21] ), .B2(new_n11926_), .ZN(new_n11929_));
  INV_X1     g11737(.I(new_n11929_), .ZN(new_n11930_));
  NAND2_X1   g11738(.A1(new_n11915_), .A2(new_n5708_), .ZN(new_n11931_));
  OAI21_X1   g11739(.A1(new_n11923_), .A2(new_n11931_), .B(new_n11930_), .ZN(new_n11932_));
  AOI21_X1   g11740(.A1(new_n11932_), .A2(new_n11924_), .B(new_n5277_), .ZN(new_n11933_));
  NOR2_X1    g11741(.A1(new_n11443_), .A2(new_n11426_), .ZN(new_n11934_));
  INV_X1     g11742(.I(new_n11934_), .ZN(new_n11935_));
  NAND3_X1   g11743(.A1(\asqrt[21] ), .A2(new_n11427_), .A3(new_n11935_), .ZN(new_n11936_));
  AND3_X2    g11744(.A1(new_n11935_), .A2(new_n11427_), .A3(new_n11432_), .Z(new_n11937_));
  AOI22_X1   g11745(.A1(new_n11936_), .A2(new_n11433_), .B1(\asqrt[21] ), .B2(new_n11937_), .ZN(new_n11938_));
  OAI21_X1   g11746(.A1(new_n11921_), .A2(new_n11922_), .B(new_n11915_), .ZN(new_n11939_));
  AOI21_X1   g11747(.A1(new_n11939_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n11940_));
  AOI21_X1   g11748(.A1(new_n11940_), .A2(new_n11932_), .B(new_n11938_), .ZN(new_n11941_));
  OAI21_X1   g11749(.A1(new_n11941_), .A2(new_n11933_), .B(\asqrt[37] ), .ZN(new_n11942_));
  INV_X1     g11750(.I(new_n11942_), .ZN(new_n11943_));
  NOR2_X1    g11751(.A1(new_n11447_), .A2(new_n11454_), .ZN(new_n11944_));
  NOR3_X1    g11752(.A1(new_n11944_), .A2(new_n11461_), .A3(new_n11453_), .ZN(new_n11945_));
  NOR3_X1    g11753(.A1(new_n11736_), .A2(new_n11461_), .A3(new_n11944_), .ZN(new_n11946_));
  INV_X1     g11754(.I(new_n11946_), .ZN(new_n11947_));
  AOI22_X1   g11755(.A1(new_n11947_), .A2(new_n11453_), .B1(\asqrt[21] ), .B2(new_n11945_), .ZN(new_n11948_));
  NOR3_X1    g11756(.A1(new_n11941_), .A2(new_n11933_), .A3(\asqrt[37] ), .ZN(new_n11949_));
  NOR2_X1    g11757(.A1(new_n11949_), .A2(new_n11948_), .ZN(new_n11950_));
  OAI21_X1   g11758(.A1(new_n11950_), .A2(new_n11943_), .B(\asqrt[38] ), .ZN(new_n11951_));
  INV_X1     g11759(.I(new_n11460_), .ZN(new_n11952_));
  NOR3_X1    g11760(.A1(new_n11736_), .A2(new_n11456_), .A3(new_n11505_), .ZN(new_n11953_));
  INV_X1     g11761(.I(new_n11953_), .ZN(new_n11954_));
  NOR3_X1    g11762(.A1(new_n11456_), .A2(new_n11952_), .A3(new_n11505_), .ZN(new_n11955_));
  AOI22_X1   g11763(.A1(new_n11954_), .A2(new_n11952_), .B1(\asqrt[21] ), .B2(new_n11955_), .ZN(new_n11956_));
  INV_X1     g11764(.I(new_n11956_), .ZN(new_n11957_));
  NAND2_X1   g11765(.A1(new_n11942_), .A2(new_n4696_), .ZN(new_n11958_));
  OAI21_X1   g11766(.A1(new_n11950_), .A2(new_n11958_), .B(new_n11957_), .ZN(new_n11959_));
  AOI21_X1   g11767(.A1(new_n11959_), .A2(new_n11951_), .B(new_n4298_), .ZN(new_n11960_));
  NOR3_X1    g11768(.A1(new_n11465_), .A2(new_n11487_), .A3(new_n11471_), .ZN(new_n11961_));
  NOR3_X1    g11769(.A1(new_n11736_), .A2(new_n11465_), .A3(new_n11471_), .ZN(new_n11962_));
  INV_X1     g11770(.I(new_n11962_), .ZN(new_n11963_));
  AOI22_X1   g11771(.A1(new_n11963_), .A2(new_n11487_), .B1(\asqrt[21] ), .B2(new_n11961_), .ZN(new_n11964_));
  OAI21_X1   g11772(.A1(new_n11948_), .A2(new_n11949_), .B(new_n11942_), .ZN(new_n11965_));
  AOI21_X1   g11773(.A1(new_n11965_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n11966_));
  AOI21_X1   g11774(.A1(new_n11966_), .A2(new_n11959_), .B(new_n11964_), .ZN(new_n11967_));
  OAI21_X1   g11775(.A1(new_n11967_), .A2(new_n11960_), .B(\asqrt[40] ), .ZN(new_n11968_));
  INV_X1     g11776(.I(new_n11968_), .ZN(new_n11969_));
  NOR2_X1    g11777(.A1(new_n11472_), .A2(new_n11480_), .ZN(new_n11970_));
  NOR3_X1    g11778(.A1(new_n11736_), .A2(new_n11495_), .A3(new_n11970_), .ZN(new_n11971_));
  INV_X1     g11779(.I(new_n11971_), .ZN(new_n11972_));
  NOR3_X1    g11780(.A1(new_n11970_), .A2(new_n11495_), .A3(new_n11479_), .ZN(new_n11973_));
  AOI22_X1   g11781(.A1(new_n11972_), .A2(new_n11479_), .B1(\asqrt[21] ), .B2(new_n11973_), .ZN(new_n11974_));
  NOR3_X1    g11782(.A1(new_n11967_), .A2(new_n11960_), .A3(\asqrt[40] ), .ZN(new_n11975_));
  NOR2_X1    g11783(.A1(new_n11975_), .A2(new_n11974_), .ZN(new_n11976_));
  OAI21_X1   g11784(.A1(new_n11976_), .A2(new_n11969_), .B(\asqrt[41] ), .ZN(new_n11977_));
  INV_X1     g11785(.I(new_n11486_), .ZN(new_n11978_));
  NOR3_X1    g11786(.A1(new_n11482_), .A2(new_n11978_), .A3(new_n11518_), .ZN(new_n11979_));
  NOR3_X1    g11787(.A1(new_n11736_), .A2(new_n11482_), .A3(new_n11518_), .ZN(new_n11980_));
  INV_X1     g11788(.I(new_n11980_), .ZN(new_n11981_));
  AOI22_X1   g11789(.A1(new_n11981_), .A2(new_n11978_), .B1(\asqrt[21] ), .B2(new_n11979_), .ZN(new_n11982_));
  INV_X1     g11790(.I(new_n11982_), .ZN(new_n11983_));
  NAND2_X1   g11791(.A1(new_n11968_), .A2(new_n3782_), .ZN(new_n11984_));
  OAI21_X1   g11792(.A1(new_n11976_), .A2(new_n11984_), .B(new_n11983_), .ZN(new_n11985_));
  AOI21_X1   g11793(.A1(new_n11985_), .A2(new_n11977_), .B(new_n3419_), .ZN(new_n11986_));
  NOR3_X1    g11794(.A1(new_n11736_), .A2(new_n11756_), .A3(new_n11757_), .ZN(new_n11987_));
  INV_X1     g11795(.I(new_n11987_), .ZN(new_n11988_));
  NOR3_X1    g11796(.A1(new_n11756_), .A2(new_n11504_), .A3(new_n11757_), .ZN(new_n11989_));
  AOI22_X1   g11797(.A1(new_n11988_), .A2(new_n11504_), .B1(\asqrt[21] ), .B2(new_n11989_), .ZN(new_n11990_));
  OAI21_X1   g11798(.A1(new_n11974_), .A2(new_n11975_), .B(new_n11968_), .ZN(new_n11991_));
  AOI21_X1   g11799(.A1(new_n11991_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n11992_));
  AOI21_X1   g11800(.A1(new_n11992_), .A2(new_n11985_), .B(new_n11990_), .ZN(new_n11993_));
  OAI21_X1   g11801(.A1(new_n11993_), .A2(new_n11986_), .B(\asqrt[43] ), .ZN(new_n11994_));
  INV_X1     g11802(.I(new_n11994_), .ZN(new_n11995_));
  INV_X1     g11803(.I(new_n11517_), .ZN(new_n11996_));
  NAND2_X1   g11804(.A1(new_n11498_), .A2(new_n3419_), .ZN(new_n11997_));
  NOR2_X1    g11805(.A1(new_n11758_), .A2(new_n11997_), .ZN(new_n11998_));
  NOR3_X1    g11806(.A1(new_n11998_), .A2(new_n11512_), .A3(new_n11996_), .ZN(new_n11999_));
  NOR3_X1    g11807(.A1(new_n11736_), .A2(new_n11512_), .A3(new_n11998_), .ZN(new_n12000_));
  INV_X1     g11808(.I(new_n12000_), .ZN(new_n12001_));
  AOI22_X1   g11809(.A1(new_n12001_), .A2(new_n11996_), .B1(\asqrt[21] ), .B2(new_n11999_), .ZN(new_n12002_));
  NOR3_X1    g11810(.A1(new_n11993_), .A2(new_n11986_), .A3(\asqrt[43] ), .ZN(new_n12003_));
  NOR2_X1    g11811(.A1(new_n12003_), .A2(new_n12002_), .ZN(new_n12004_));
  OAI21_X1   g11812(.A1(new_n12004_), .A2(new_n11995_), .B(\asqrt[44] ), .ZN(new_n12005_));
  NOR3_X1    g11813(.A1(new_n11736_), .A2(new_n11523_), .A3(new_n11528_), .ZN(new_n12006_));
  INV_X1     g11814(.I(new_n12006_), .ZN(new_n12007_));
  NOR3_X1    g11815(.A1(new_n11523_), .A2(new_n11528_), .A3(new_n11755_), .ZN(new_n12008_));
  AOI22_X1   g11816(.A1(new_n12007_), .A2(new_n11755_), .B1(\asqrt[21] ), .B2(new_n12008_), .ZN(new_n12009_));
  INV_X1     g11817(.I(new_n12009_), .ZN(new_n12010_));
  NAND2_X1   g11818(.A1(new_n11994_), .A2(new_n2954_), .ZN(new_n12011_));
  OAI21_X1   g11819(.A1(new_n12004_), .A2(new_n12011_), .B(new_n12010_), .ZN(new_n12012_));
  AOI21_X1   g11820(.A1(new_n12012_), .A2(new_n12005_), .B(new_n2641_), .ZN(new_n12013_));
  INV_X1     g11821(.I(new_n11530_), .ZN(new_n12014_));
  NOR2_X1    g11822(.A1(new_n11529_), .A2(new_n11537_), .ZN(new_n12015_));
  NOR3_X1    g11823(.A1(new_n12014_), .A2(new_n12015_), .A3(new_n11536_), .ZN(new_n12016_));
  NOR3_X1    g11824(.A1(new_n11736_), .A2(new_n12014_), .A3(new_n12015_), .ZN(new_n12017_));
  INV_X1     g11825(.I(new_n12017_), .ZN(new_n12018_));
  AOI22_X1   g11826(.A1(new_n12018_), .A2(new_n11536_), .B1(\asqrt[21] ), .B2(new_n12016_), .ZN(new_n12019_));
  OAI21_X1   g11827(.A1(new_n12002_), .A2(new_n12003_), .B(new_n11994_), .ZN(new_n12020_));
  AOI21_X1   g11828(.A1(new_n12020_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n12021_));
  AOI21_X1   g11829(.A1(new_n12021_), .A2(new_n12012_), .B(new_n12019_), .ZN(new_n12022_));
  OAI21_X1   g11830(.A1(new_n12022_), .A2(new_n12013_), .B(\asqrt[46] ), .ZN(new_n12023_));
  INV_X1     g11831(.I(new_n12023_), .ZN(new_n12024_));
  INV_X1     g11832(.I(new_n11544_), .ZN(new_n12025_));
  INV_X1     g11833(.I(new_n11538_), .ZN(new_n12026_));
  INV_X1     g11834(.I(new_n11546_), .ZN(new_n12027_));
  NOR2_X1    g11835(.A1(new_n12027_), .A2(new_n12026_), .ZN(new_n12028_));
  NOR3_X1    g11836(.A1(new_n11736_), .A2(new_n11539_), .A3(new_n12028_), .ZN(new_n12029_));
  INV_X1     g11837(.I(new_n12029_), .ZN(new_n12030_));
  NOR3_X1    g11838(.A1(new_n12028_), .A2(new_n11539_), .A3(new_n12025_), .ZN(new_n12031_));
  AOI22_X1   g11839(.A1(new_n12030_), .A2(new_n12025_), .B1(\asqrt[21] ), .B2(new_n12031_), .ZN(new_n12032_));
  NOR3_X1    g11840(.A1(new_n12022_), .A2(new_n12013_), .A3(\asqrt[46] ), .ZN(new_n12033_));
  NOR2_X1    g11841(.A1(new_n12033_), .A2(new_n12032_), .ZN(new_n12034_));
  OAI21_X1   g11842(.A1(new_n12034_), .A2(new_n12024_), .B(\asqrt[47] ), .ZN(new_n12035_));
  NOR3_X1    g11843(.A1(new_n11549_), .A2(new_n11754_), .A3(new_n11554_), .ZN(new_n12036_));
  NOR3_X1    g11844(.A1(new_n11736_), .A2(new_n11549_), .A3(new_n11554_), .ZN(new_n12037_));
  INV_X1     g11845(.I(new_n12037_), .ZN(new_n12038_));
  AOI22_X1   g11846(.A1(new_n12038_), .A2(new_n11754_), .B1(\asqrt[21] ), .B2(new_n12036_), .ZN(new_n12039_));
  INV_X1     g11847(.I(new_n12039_), .ZN(new_n12040_));
  NAND2_X1   g11848(.A1(new_n12023_), .A2(new_n2229_), .ZN(new_n12041_));
  OAI21_X1   g11849(.A1(new_n12034_), .A2(new_n12041_), .B(new_n12040_), .ZN(new_n12042_));
  AOI21_X1   g11850(.A1(new_n12042_), .A2(new_n12035_), .B(new_n1956_), .ZN(new_n12043_));
  INV_X1     g11851(.I(new_n11556_), .ZN(new_n12044_));
  NOR2_X1    g11852(.A1(new_n11555_), .A2(new_n11563_), .ZN(new_n12045_));
  NOR3_X1    g11853(.A1(new_n11736_), .A2(new_n12044_), .A3(new_n12045_), .ZN(new_n12046_));
  INV_X1     g11854(.I(new_n12046_), .ZN(new_n12047_));
  NOR3_X1    g11855(.A1(new_n12044_), .A2(new_n12045_), .A3(new_n11562_), .ZN(new_n12048_));
  AOI22_X1   g11856(.A1(new_n12047_), .A2(new_n11562_), .B1(\asqrt[21] ), .B2(new_n12048_), .ZN(new_n12049_));
  OAI21_X1   g11857(.A1(new_n12032_), .A2(new_n12033_), .B(new_n12023_), .ZN(new_n12050_));
  AOI21_X1   g11858(.A1(new_n12050_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n12051_));
  AOI21_X1   g11859(.A1(new_n12051_), .A2(new_n12042_), .B(new_n12049_), .ZN(new_n12052_));
  OAI21_X1   g11860(.A1(new_n12052_), .A2(new_n12043_), .B(\asqrt[49] ), .ZN(new_n12053_));
  INV_X1     g11861(.I(new_n12053_), .ZN(new_n12054_));
  INV_X1     g11862(.I(new_n11570_), .ZN(new_n12055_));
  INV_X1     g11863(.I(new_n11564_), .ZN(new_n12056_));
  INV_X1     g11864(.I(new_n11572_), .ZN(new_n12057_));
  NOR2_X1    g11865(.A1(new_n12057_), .A2(new_n12056_), .ZN(new_n12058_));
  NOR3_X1    g11866(.A1(new_n12058_), .A2(new_n11565_), .A3(new_n12055_), .ZN(new_n12059_));
  NOR3_X1    g11867(.A1(new_n11736_), .A2(new_n11565_), .A3(new_n12058_), .ZN(new_n12060_));
  INV_X1     g11868(.I(new_n12060_), .ZN(new_n12061_));
  AOI22_X1   g11869(.A1(new_n12061_), .A2(new_n12055_), .B1(\asqrt[21] ), .B2(new_n12059_), .ZN(new_n12062_));
  NOR3_X1    g11870(.A1(new_n12052_), .A2(new_n12043_), .A3(\asqrt[49] ), .ZN(new_n12063_));
  NOR2_X1    g11871(.A1(new_n12063_), .A2(new_n12062_), .ZN(new_n12064_));
  OAI21_X1   g11872(.A1(new_n12064_), .A2(new_n12054_), .B(\asqrt[50] ), .ZN(new_n12065_));
  NOR3_X1    g11873(.A1(new_n11736_), .A2(new_n11575_), .A3(new_n11580_), .ZN(new_n12066_));
  INV_X1     g11874(.I(new_n12066_), .ZN(new_n12067_));
  NOR3_X1    g11875(.A1(new_n11575_), .A2(new_n11753_), .A3(new_n11580_), .ZN(new_n12068_));
  AOI22_X1   g11876(.A1(new_n12067_), .A2(new_n11753_), .B1(\asqrt[21] ), .B2(new_n12068_), .ZN(new_n12069_));
  INV_X1     g11877(.I(new_n12069_), .ZN(new_n12070_));
  NAND2_X1   g11878(.A1(new_n12053_), .A2(new_n1612_), .ZN(new_n12071_));
  OAI21_X1   g11879(.A1(new_n12064_), .A2(new_n12071_), .B(new_n12070_), .ZN(new_n12072_));
  AOI21_X1   g11880(.A1(new_n12072_), .A2(new_n12065_), .B(new_n1376_), .ZN(new_n12073_));
  INV_X1     g11881(.I(new_n11582_), .ZN(new_n12074_));
  NOR2_X1    g11882(.A1(new_n11581_), .A2(new_n11589_), .ZN(new_n12075_));
  NOR3_X1    g11883(.A1(new_n12074_), .A2(new_n11588_), .A3(new_n12075_), .ZN(new_n12076_));
  NOR3_X1    g11884(.A1(new_n11736_), .A2(new_n12074_), .A3(new_n12075_), .ZN(new_n12077_));
  INV_X1     g11885(.I(new_n12077_), .ZN(new_n12078_));
  AOI22_X1   g11886(.A1(new_n12078_), .A2(new_n11588_), .B1(\asqrt[21] ), .B2(new_n12076_), .ZN(new_n12079_));
  OAI21_X1   g11887(.A1(new_n12062_), .A2(new_n12063_), .B(new_n12053_), .ZN(new_n12080_));
  AOI21_X1   g11888(.A1(new_n12080_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n12081_));
  AOI21_X1   g11889(.A1(new_n12081_), .A2(new_n12072_), .B(new_n12079_), .ZN(new_n12082_));
  OAI21_X1   g11890(.A1(new_n12082_), .A2(new_n12073_), .B(\asqrt[52] ), .ZN(new_n12083_));
  INV_X1     g11891(.I(new_n12083_), .ZN(new_n12084_));
  INV_X1     g11892(.I(new_n11596_), .ZN(new_n12085_));
  INV_X1     g11893(.I(new_n11590_), .ZN(new_n12086_));
  INV_X1     g11894(.I(new_n11598_), .ZN(new_n12087_));
  NOR2_X1    g11895(.A1(new_n12087_), .A2(new_n12086_), .ZN(new_n12088_));
  NOR3_X1    g11896(.A1(new_n11736_), .A2(new_n11591_), .A3(new_n12088_), .ZN(new_n12089_));
  INV_X1     g11897(.I(new_n12089_), .ZN(new_n12090_));
  NOR3_X1    g11898(.A1(new_n12088_), .A2(new_n11591_), .A3(new_n12085_), .ZN(new_n12091_));
  AOI22_X1   g11899(.A1(new_n12090_), .A2(new_n12085_), .B1(\asqrt[21] ), .B2(new_n12091_), .ZN(new_n12092_));
  NOR3_X1    g11900(.A1(new_n12082_), .A2(new_n12073_), .A3(\asqrt[52] ), .ZN(new_n12093_));
  NOR2_X1    g11901(.A1(new_n12093_), .A2(new_n12092_), .ZN(new_n12094_));
  OAI21_X1   g11902(.A1(new_n12094_), .A2(new_n12084_), .B(\asqrt[53] ), .ZN(new_n12095_));
  NOR3_X1    g11903(.A1(new_n11601_), .A2(new_n11752_), .A3(new_n11643_), .ZN(new_n12096_));
  NOR3_X1    g11904(.A1(new_n11736_), .A2(new_n11601_), .A3(new_n11643_), .ZN(new_n12097_));
  INV_X1     g11905(.I(new_n12097_), .ZN(new_n12098_));
  AOI22_X1   g11906(.A1(new_n12098_), .A2(new_n11752_), .B1(\asqrt[21] ), .B2(new_n12096_), .ZN(new_n12099_));
  INV_X1     g11907(.I(new_n12099_), .ZN(new_n12100_));
  NAND2_X1   g11908(.A1(new_n12083_), .A2(new_n1103_), .ZN(new_n12101_));
  OAI21_X1   g11909(.A1(new_n12094_), .A2(new_n12101_), .B(new_n12100_), .ZN(new_n12102_));
  AOI21_X1   g11910(.A1(new_n12102_), .A2(new_n12095_), .B(new_n904_), .ZN(new_n12103_));
  INV_X1     g11911(.I(new_n11609_), .ZN(new_n12104_));
  NOR2_X1    g11912(.A1(new_n11616_), .A2(new_n11608_), .ZN(new_n12105_));
  NOR3_X1    g11913(.A1(new_n11736_), .A2(new_n12104_), .A3(new_n12105_), .ZN(new_n12106_));
  INV_X1     g11914(.I(new_n12106_), .ZN(new_n12107_));
  NOR3_X1    g11915(.A1(new_n12104_), .A2(new_n11615_), .A3(new_n12105_), .ZN(new_n12108_));
  AOI22_X1   g11916(.A1(new_n12107_), .A2(new_n11615_), .B1(\asqrt[21] ), .B2(new_n12108_), .ZN(new_n12109_));
  OAI21_X1   g11917(.A1(new_n12092_), .A2(new_n12093_), .B(new_n12083_), .ZN(new_n12110_));
  AOI21_X1   g11918(.A1(new_n12110_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n12111_));
  AOI21_X1   g11919(.A1(new_n12111_), .A2(new_n12102_), .B(new_n12109_), .ZN(new_n12112_));
  OAI21_X1   g11920(.A1(new_n12112_), .A2(new_n12103_), .B(\asqrt[55] ), .ZN(new_n12113_));
  INV_X1     g11921(.I(new_n12113_), .ZN(new_n12114_));
  NOR2_X1    g11922(.A1(new_n11627_), .A2(new_n11620_), .ZN(new_n12115_));
  NOR3_X1    g11923(.A1(new_n12115_), .A2(new_n11618_), .A3(new_n11626_), .ZN(new_n12116_));
  NOR3_X1    g11924(.A1(new_n11736_), .A2(new_n11618_), .A3(new_n12115_), .ZN(new_n12117_));
  INV_X1     g11925(.I(new_n12117_), .ZN(new_n12118_));
  AOI22_X1   g11926(.A1(new_n12118_), .A2(new_n11626_), .B1(\asqrt[21] ), .B2(new_n12116_), .ZN(new_n12119_));
  NOR3_X1    g11927(.A1(new_n12112_), .A2(new_n12103_), .A3(\asqrt[55] ), .ZN(new_n12120_));
  NOR2_X1    g11928(.A1(new_n12120_), .A2(new_n12119_), .ZN(new_n12121_));
  OAI21_X1   g11929(.A1(new_n12121_), .A2(new_n12114_), .B(\asqrt[56] ), .ZN(new_n12122_));
  NOR3_X1    g11930(.A1(new_n11736_), .A2(new_n11629_), .A3(new_n11675_), .ZN(new_n12123_));
  INV_X1     g11931(.I(new_n12123_), .ZN(new_n12124_));
  NOR3_X1    g11932(.A1(new_n11629_), .A2(new_n11751_), .A3(new_n11675_), .ZN(new_n12125_));
  AOI22_X1   g11933(.A1(new_n12124_), .A2(new_n11751_), .B1(\asqrt[21] ), .B2(new_n12125_), .ZN(new_n12126_));
  INV_X1     g11934(.I(new_n12126_), .ZN(new_n12127_));
  NAND2_X1   g11935(.A1(new_n12113_), .A2(new_n703_), .ZN(new_n12128_));
  OAI21_X1   g11936(.A1(new_n12121_), .A2(new_n12128_), .B(new_n12127_), .ZN(new_n12129_));
  AOI21_X1   g11937(.A1(new_n12129_), .A2(new_n12122_), .B(new_n531_), .ZN(new_n12130_));
  INV_X1     g11938(.I(new_n11636_), .ZN(new_n12131_));
  NOR2_X1    g11939(.A1(new_n11648_), .A2(new_n11635_), .ZN(new_n12132_));
  NOR3_X1    g11940(.A1(new_n12131_), .A2(new_n11642_), .A3(new_n12132_), .ZN(new_n12133_));
  NOR3_X1    g11941(.A1(new_n11736_), .A2(new_n12131_), .A3(new_n12132_), .ZN(new_n12134_));
  INV_X1     g11942(.I(new_n12134_), .ZN(new_n12135_));
  AOI22_X1   g11943(.A1(new_n12135_), .A2(new_n11642_), .B1(\asqrt[21] ), .B2(new_n12133_), .ZN(new_n12136_));
  OAI21_X1   g11944(.A1(new_n12119_), .A2(new_n12120_), .B(new_n12113_), .ZN(new_n12137_));
  AOI21_X1   g11945(.A1(new_n12137_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n12138_));
  AOI21_X1   g11946(.A1(new_n12138_), .A2(new_n12129_), .B(new_n12136_), .ZN(new_n12139_));
  OAI21_X1   g11947(.A1(new_n12139_), .A2(new_n12130_), .B(\asqrt[58] ), .ZN(new_n12140_));
  NOR2_X1    g11948(.A1(new_n11659_), .A2(new_n11652_), .ZN(new_n12141_));
  NOR3_X1    g11949(.A1(new_n11736_), .A2(new_n11650_), .A3(new_n12141_), .ZN(new_n12142_));
  INV_X1     g11950(.I(new_n12142_), .ZN(new_n12143_));
  NOR3_X1    g11951(.A1(new_n12141_), .A2(new_n11650_), .A3(new_n11658_), .ZN(new_n12144_));
  AOI22_X1   g11952(.A1(new_n12143_), .A2(new_n11658_), .B1(\asqrt[21] ), .B2(new_n12144_), .ZN(new_n12145_));
  INV_X1     g11953(.I(new_n12145_), .ZN(new_n12146_));
  INV_X1     g11954(.I(new_n12119_), .ZN(new_n12147_));
  INV_X1     g11955(.I(new_n12092_), .ZN(new_n12148_));
  INV_X1     g11956(.I(new_n12062_), .ZN(new_n12149_));
  INV_X1     g11957(.I(new_n12032_), .ZN(new_n12150_));
  INV_X1     g11958(.I(new_n12002_), .ZN(new_n12151_));
  INV_X1     g11959(.I(new_n11974_), .ZN(new_n12152_));
  INV_X1     g11960(.I(new_n11948_), .ZN(new_n12153_));
  INV_X1     g11961(.I(new_n11921_), .ZN(new_n12154_));
  INV_X1     g11962(.I(new_n11893_), .ZN(new_n12155_));
  INV_X1     g11963(.I(new_n11867_), .ZN(new_n12156_));
  NAND2_X1   g11964(.A1(new_n11809_), .A2(new_n9846_), .ZN(new_n12157_));
  OAI21_X1   g11965(.A1(new_n12157_), .A2(new_n11841_), .B(new_n11823_), .ZN(new_n12158_));
  AOI21_X1   g11966(.A1(new_n12158_), .A2(new_n11851_), .B(new_n9317_), .ZN(new_n12159_));
  NOR2_X1    g11967(.A1(new_n11817_), .A2(\asqrt[26] ), .ZN(new_n12160_));
  AOI21_X1   g11968(.A1(new_n12160_), .A2(new_n12158_), .B(new_n11849_), .ZN(new_n12161_));
  OAI21_X1   g11969(.A1(new_n12161_), .A2(new_n12159_), .B(\asqrt[27] ), .ZN(new_n12162_));
  NAND2_X1   g11970(.A1(new_n12162_), .A2(new_n8483_), .ZN(new_n12163_));
  OAI21_X1   g11971(.A1(new_n12163_), .A2(new_n11861_), .B(new_n12156_), .ZN(new_n12164_));
  NAND3_X1   g11972(.A1(new_n12164_), .A2(new_n8036_), .A3(new_n11862_), .ZN(new_n12165_));
  AOI22_X1   g11973(.A1(new_n12165_), .A2(new_n11876_), .B1(\asqrt[29] ), .B2(new_n11884_), .ZN(new_n12166_));
  OAI21_X1   g11974(.A1(new_n12166_), .A2(new_n7539_), .B(new_n7229_), .ZN(new_n12167_));
  OAI21_X1   g11975(.A1(new_n12167_), .A2(new_n11886_), .B(new_n12155_), .ZN(new_n12168_));
  AOI21_X1   g11976(.A1(new_n12168_), .A2(new_n11887_), .B(new_n6824_), .ZN(new_n12169_));
  AOI21_X1   g11977(.A1(new_n12164_), .A2(new_n11862_), .B(new_n8036_), .ZN(new_n12170_));
  NOR3_X1    g11978(.A1(new_n12161_), .A2(new_n12159_), .A3(\asqrt[27] ), .ZN(new_n12171_));
  OAI21_X1   g11979(.A1(new_n11858_), .A2(new_n12171_), .B(new_n12162_), .ZN(new_n12172_));
  AOI21_X1   g11980(.A1(new_n12172_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n12173_));
  AOI21_X1   g11981(.A1(new_n12173_), .A2(new_n12164_), .B(new_n11875_), .ZN(new_n12174_));
  NOR3_X1    g11982(.A1(new_n12174_), .A2(\asqrt[30] ), .A3(new_n12170_), .ZN(new_n12175_));
  OAI22_X1   g11983(.A1(new_n12175_), .A2(new_n11883_), .B1(new_n12166_), .B2(new_n7539_), .ZN(new_n12176_));
  AOI21_X1   g11984(.A1(new_n12176_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n12177_));
  AOI21_X1   g11985(.A1(new_n12177_), .A2(new_n12168_), .B(new_n11901_), .ZN(new_n12178_));
  OAI21_X1   g11986(.A1(new_n12178_), .A2(new_n12169_), .B(\asqrt[33] ), .ZN(new_n12179_));
  NAND2_X1   g11987(.A1(new_n12179_), .A2(new_n6077_), .ZN(new_n12180_));
  OAI21_X1   g11988(.A1(new_n12180_), .A2(new_n11914_), .B(new_n12154_), .ZN(new_n12181_));
  AOI21_X1   g11989(.A1(new_n12181_), .A2(new_n11915_), .B(new_n5708_), .ZN(new_n12182_));
  NOR3_X1    g11990(.A1(new_n12178_), .A2(\asqrt[33] ), .A3(new_n12169_), .ZN(new_n12183_));
  OAI21_X1   g11991(.A1(new_n11911_), .A2(new_n12183_), .B(new_n12179_), .ZN(new_n12184_));
  AOI21_X1   g11992(.A1(new_n12184_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n12185_));
  AOI21_X1   g11993(.A1(new_n12185_), .A2(new_n12181_), .B(new_n11929_), .ZN(new_n12186_));
  OAI21_X1   g11994(.A1(new_n12186_), .A2(new_n12182_), .B(\asqrt[36] ), .ZN(new_n12187_));
  NAND2_X1   g11995(.A1(new_n12187_), .A2(new_n5024_), .ZN(new_n12188_));
  OAI21_X1   g11996(.A1(new_n12188_), .A2(new_n11941_), .B(new_n12153_), .ZN(new_n12189_));
  AOI21_X1   g11997(.A1(new_n12189_), .A2(new_n11942_), .B(new_n4696_), .ZN(new_n12190_));
  NOR3_X1    g11998(.A1(new_n12186_), .A2(\asqrt[36] ), .A3(new_n12182_), .ZN(new_n12191_));
  OAI21_X1   g11999(.A1(new_n11938_), .A2(new_n12191_), .B(new_n12187_), .ZN(new_n12192_));
  AOI21_X1   g12000(.A1(new_n12192_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n12193_));
  AOI21_X1   g12001(.A1(new_n12193_), .A2(new_n12189_), .B(new_n11956_), .ZN(new_n12194_));
  OAI21_X1   g12002(.A1(new_n12194_), .A2(new_n12190_), .B(\asqrt[39] ), .ZN(new_n12195_));
  NAND2_X1   g12003(.A1(new_n12195_), .A2(new_n4071_), .ZN(new_n12196_));
  OAI21_X1   g12004(.A1(new_n12196_), .A2(new_n11967_), .B(new_n12152_), .ZN(new_n12197_));
  AOI21_X1   g12005(.A1(new_n12197_), .A2(new_n11968_), .B(new_n3782_), .ZN(new_n12198_));
  NOR3_X1    g12006(.A1(new_n12194_), .A2(\asqrt[39] ), .A3(new_n12190_), .ZN(new_n12199_));
  OAI21_X1   g12007(.A1(new_n11964_), .A2(new_n12199_), .B(new_n12195_), .ZN(new_n12200_));
  AOI21_X1   g12008(.A1(new_n12200_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n12201_));
  AOI21_X1   g12009(.A1(new_n12201_), .A2(new_n12197_), .B(new_n11982_), .ZN(new_n12202_));
  OAI21_X1   g12010(.A1(new_n12202_), .A2(new_n12198_), .B(\asqrt[42] ), .ZN(new_n12203_));
  NAND2_X1   g12011(.A1(new_n12203_), .A2(new_n3218_), .ZN(new_n12204_));
  OAI21_X1   g12012(.A1(new_n12204_), .A2(new_n11993_), .B(new_n12151_), .ZN(new_n12205_));
  AOI21_X1   g12013(.A1(new_n12205_), .A2(new_n11994_), .B(new_n2954_), .ZN(new_n12206_));
  NOR3_X1    g12014(.A1(new_n12202_), .A2(\asqrt[42] ), .A3(new_n12198_), .ZN(new_n12207_));
  OAI21_X1   g12015(.A1(new_n11990_), .A2(new_n12207_), .B(new_n12203_), .ZN(new_n12208_));
  AOI21_X1   g12016(.A1(new_n12208_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n12209_));
  AOI21_X1   g12017(.A1(new_n12209_), .A2(new_n12205_), .B(new_n12009_), .ZN(new_n12210_));
  OAI21_X1   g12018(.A1(new_n12210_), .A2(new_n12206_), .B(\asqrt[45] ), .ZN(new_n12211_));
  NAND2_X1   g12019(.A1(new_n12211_), .A2(new_n2465_), .ZN(new_n12212_));
  OAI21_X1   g12020(.A1(new_n12212_), .A2(new_n12022_), .B(new_n12150_), .ZN(new_n12213_));
  AOI21_X1   g12021(.A1(new_n12213_), .A2(new_n12023_), .B(new_n2229_), .ZN(new_n12214_));
  NOR3_X1    g12022(.A1(new_n12210_), .A2(\asqrt[45] ), .A3(new_n12206_), .ZN(new_n12215_));
  OAI21_X1   g12023(.A1(new_n12019_), .A2(new_n12215_), .B(new_n12211_), .ZN(new_n12216_));
  AOI21_X1   g12024(.A1(new_n12216_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n12217_));
  AOI21_X1   g12025(.A1(new_n12217_), .A2(new_n12213_), .B(new_n12039_), .ZN(new_n12218_));
  OAI21_X1   g12026(.A1(new_n12218_), .A2(new_n12214_), .B(\asqrt[48] ), .ZN(new_n12219_));
  NAND2_X1   g12027(.A1(new_n12219_), .A2(new_n1806_), .ZN(new_n12220_));
  OAI21_X1   g12028(.A1(new_n12220_), .A2(new_n12052_), .B(new_n12149_), .ZN(new_n12221_));
  AOI21_X1   g12029(.A1(new_n12221_), .A2(new_n12053_), .B(new_n1612_), .ZN(new_n12222_));
  NOR3_X1    g12030(.A1(new_n12218_), .A2(\asqrt[48] ), .A3(new_n12214_), .ZN(new_n12223_));
  OAI21_X1   g12031(.A1(new_n12049_), .A2(new_n12223_), .B(new_n12219_), .ZN(new_n12224_));
  AOI21_X1   g12032(.A1(new_n12224_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n12225_));
  AOI21_X1   g12033(.A1(new_n12225_), .A2(new_n12221_), .B(new_n12069_), .ZN(new_n12226_));
  OAI21_X1   g12034(.A1(new_n12226_), .A2(new_n12222_), .B(\asqrt[51] ), .ZN(new_n12227_));
  NAND2_X1   g12035(.A1(new_n12227_), .A2(new_n1256_), .ZN(new_n12228_));
  OAI21_X1   g12036(.A1(new_n12228_), .A2(new_n12082_), .B(new_n12148_), .ZN(new_n12229_));
  NAND3_X1   g12037(.A1(new_n12229_), .A2(new_n1103_), .A3(new_n12083_), .ZN(new_n12230_));
  AOI22_X1   g12038(.A1(new_n12230_), .A2(new_n12100_), .B1(\asqrt[53] ), .B2(new_n12110_), .ZN(new_n12231_));
  OAI21_X1   g12039(.A1(new_n12231_), .A2(new_n904_), .B(new_n823_), .ZN(new_n12232_));
  OAI21_X1   g12040(.A1(new_n12232_), .A2(new_n12112_), .B(new_n12147_), .ZN(new_n12233_));
  NAND3_X1   g12041(.A1(new_n12233_), .A2(new_n703_), .A3(new_n12113_), .ZN(new_n12234_));
  AOI22_X1   g12042(.A1(new_n12234_), .A2(new_n12127_), .B1(\asqrt[56] ), .B2(new_n12137_), .ZN(new_n12235_));
  OAI21_X1   g12043(.A1(new_n12235_), .A2(new_n531_), .B(new_n436_), .ZN(new_n12236_));
  OAI21_X1   g12044(.A1(new_n12236_), .A2(new_n12139_), .B(new_n12146_), .ZN(new_n12237_));
  AOI21_X1   g12045(.A1(new_n12237_), .A2(new_n12140_), .B(new_n327_), .ZN(new_n12238_));
  NOR3_X1    g12046(.A1(new_n11661_), .A2(new_n11750_), .A3(new_n11707_), .ZN(new_n12239_));
  NOR3_X1    g12047(.A1(new_n11736_), .A2(new_n11661_), .A3(new_n11707_), .ZN(new_n12240_));
  INV_X1     g12048(.I(new_n12240_), .ZN(new_n12241_));
  AOI22_X1   g12049(.A1(new_n12241_), .A2(new_n11750_), .B1(\asqrt[21] ), .B2(new_n12239_), .ZN(new_n12242_));
  NAND2_X1   g12050(.A1(new_n12140_), .A2(new_n327_), .ZN(new_n12243_));
  INV_X1     g12051(.I(new_n12243_), .ZN(new_n12244_));
  AOI21_X1   g12052(.A1(new_n12244_), .A2(new_n12237_), .B(new_n12242_), .ZN(new_n12245_));
  OAI21_X1   g12053(.A1(new_n12245_), .A2(new_n12238_), .B(\asqrt[60] ), .ZN(new_n12246_));
  INV_X1     g12054(.I(new_n11668_), .ZN(new_n12247_));
  NOR2_X1    g12055(.A1(new_n11680_), .A2(new_n11667_), .ZN(new_n12248_));
  NOR3_X1    g12056(.A1(new_n11736_), .A2(new_n12247_), .A3(new_n12248_), .ZN(new_n12249_));
  INV_X1     g12057(.I(new_n12249_), .ZN(new_n12250_));
  NOR3_X1    g12058(.A1(new_n12247_), .A2(new_n11674_), .A3(new_n12248_), .ZN(new_n12251_));
  AOI22_X1   g12059(.A1(new_n12250_), .A2(new_n11674_), .B1(\asqrt[21] ), .B2(new_n12251_), .ZN(new_n12252_));
  INV_X1     g12060(.I(new_n12252_), .ZN(new_n12253_));
  INV_X1     g12061(.I(new_n12140_), .ZN(new_n12254_));
  NOR3_X1    g12062(.A1(new_n12139_), .A2(new_n12130_), .A3(\asqrt[58] ), .ZN(new_n12255_));
  NOR2_X1    g12063(.A1(new_n12255_), .A2(new_n12145_), .ZN(new_n12256_));
  OAI21_X1   g12064(.A1(new_n12256_), .A2(new_n12254_), .B(\asqrt[59] ), .ZN(new_n12257_));
  NAND2_X1   g12065(.A1(new_n12257_), .A2(new_n306_), .ZN(new_n12258_));
  OAI21_X1   g12066(.A1(new_n12258_), .A2(new_n12245_), .B(new_n12253_), .ZN(new_n12259_));
  AOI21_X1   g12067(.A1(new_n12259_), .A2(new_n12246_), .B(new_n218_), .ZN(new_n12260_));
  NOR2_X1    g12068(.A1(new_n11684_), .A2(new_n11691_), .ZN(new_n12261_));
  NOR3_X1    g12069(.A1(new_n12261_), .A2(new_n11682_), .A3(new_n11690_), .ZN(new_n12262_));
  NOR3_X1    g12070(.A1(new_n11736_), .A2(new_n11682_), .A3(new_n12261_), .ZN(new_n12263_));
  INV_X1     g12071(.I(new_n12263_), .ZN(new_n12264_));
  AOI22_X1   g12072(.A1(new_n12264_), .A2(new_n11690_), .B1(\asqrt[21] ), .B2(new_n12262_), .ZN(new_n12265_));
  INV_X1     g12073(.I(new_n12242_), .ZN(new_n12266_));
  OAI21_X1   g12074(.A1(new_n12256_), .A2(new_n12243_), .B(new_n12266_), .ZN(new_n12267_));
  AOI21_X1   g12075(.A1(new_n12267_), .A2(new_n12257_), .B(new_n306_), .ZN(new_n12268_));
  NOR2_X1    g12076(.A1(new_n12268_), .A2(\asqrt[61] ), .ZN(new_n12269_));
  AOI21_X1   g12077(.A1(new_n12269_), .A2(new_n12259_), .B(new_n12265_), .ZN(new_n12270_));
  OAI21_X1   g12078(.A1(new_n12270_), .A2(new_n12260_), .B(\asqrt[62] ), .ZN(new_n12271_));
  NOR3_X1    g12079(.A1(new_n11736_), .A2(new_n11693_), .A3(new_n11747_), .ZN(new_n12272_));
  INV_X1     g12080(.I(new_n12272_), .ZN(new_n12273_));
  NOR3_X1    g12081(.A1(new_n11693_), .A2(new_n11749_), .A3(new_n11747_), .ZN(new_n12274_));
  AOI22_X1   g12082(.A1(new_n12273_), .A2(new_n11749_), .B1(\asqrt[21] ), .B2(new_n12274_), .ZN(new_n12275_));
  INV_X1     g12083(.I(new_n12275_), .ZN(new_n12276_));
  OAI21_X1   g12084(.A1(new_n12145_), .A2(new_n12255_), .B(new_n12140_), .ZN(new_n12277_));
  AOI21_X1   g12085(.A1(new_n12277_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n12278_));
  AOI21_X1   g12086(.A1(new_n12278_), .A2(new_n12267_), .B(new_n12252_), .ZN(new_n12279_));
  OAI21_X1   g12087(.A1(new_n12279_), .A2(new_n12268_), .B(\asqrt[61] ), .ZN(new_n12280_));
  NAND2_X1   g12088(.A1(new_n12280_), .A2(new_n207_), .ZN(new_n12281_));
  OAI21_X1   g12089(.A1(new_n12281_), .A2(new_n12270_), .B(new_n12276_), .ZN(new_n12282_));
  NAND4_X1   g12090(.A1(\asqrt[21] ), .A2(new_n11700_), .A3(new_n11705_), .A4(new_n11786_), .ZN(new_n12283_));
  NAND2_X1   g12091(.A1(new_n11700_), .A2(new_n11786_), .ZN(new_n12284_));
  OAI21_X1   g12092(.A1(new_n11736_), .A2(new_n12284_), .B(new_n11706_), .ZN(new_n12285_));
  NAND2_X1   g12093(.A1(new_n12283_), .A2(new_n12285_), .ZN(new_n12286_));
  NOR2_X1    g12094(.A1(new_n11787_), .A2(new_n11726_), .ZN(new_n12287_));
  NAND2_X1   g12095(.A1(\asqrt[21] ), .A2(new_n12287_), .ZN(new_n12288_));
  NAND3_X1   g12096(.A1(new_n12286_), .A2(new_n11798_), .A3(new_n12288_), .ZN(new_n12289_));
  AOI21_X1   g12097(.A1(new_n12282_), .A2(new_n12271_), .B(new_n12289_), .ZN(new_n12290_));
  NOR3_X1    g12098(.A1(new_n12279_), .A2(new_n12268_), .A3(\asqrt[61] ), .ZN(new_n12291_));
  OAI21_X1   g12099(.A1(new_n12265_), .A2(new_n12291_), .B(new_n12280_), .ZN(new_n12292_));
  AOI21_X1   g12100(.A1(new_n12292_), .A2(\asqrt[62] ), .B(new_n12286_), .ZN(new_n12293_));
  OAI21_X1   g12101(.A1(new_n11736_), .A2(new_n11726_), .B(new_n11787_), .ZN(new_n12294_));
  NOR2_X1    g12102(.A1(new_n12287_), .A2(new_n193_), .ZN(new_n12295_));
  NAND2_X1   g12103(.A1(new_n12294_), .A2(new_n12295_), .ZN(new_n12296_));
  INV_X1     g12104(.I(new_n12296_), .ZN(new_n12297_));
  AND3_X2    g12105(.A1(new_n11717_), .A2(new_n11715_), .A3(new_n11732_), .Z(new_n12298_));
  NAND4_X1   g12106(.A1(new_n11788_), .A2(new_n11798_), .A3(new_n11729_), .A4(new_n12298_), .ZN(new_n12299_));
  INV_X1     g12107(.I(new_n12299_), .ZN(new_n12300_));
  NOR2_X1    g12108(.A1(new_n12297_), .A2(new_n12300_), .ZN(new_n12301_));
  INV_X1     g12109(.I(new_n12301_), .ZN(new_n12302_));
  AOI21_X1   g12110(.A1(new_n12293_), .A2(new_n12282_), .B(new_n12302_), .ZN(new_n12303_));
  OAI21_X1   g12111(.A1(\asqrt[63] ), .A2(new_n12290_), .B(new_n12303_), .ZN(\asqrt[20] ));
  NOR2_X1    g12112(.A1(\a[38] ), .A2(\a[39] ), .ZN(new_n12305_));
  INV_X1     g12113(.I(new_n12305_), .ZN(new_n12306_));
  NOR2_X1    g12114(.A1(new_n12306_), .A2(\a[40] ), .ZN(new_n12307_));
  INV_X1     g12115(.I(new_n12307_), .ZN(new_n12308_));
  NAND2_X1   g12116(.A1(new_n12282_), .A2(new_n12271_), .ZN(new_n12309_));
  INV_X1     g12117(.I(new_n12289_), .ZN(new_n12310_));
  AOI21_X1   g12118(.A1(new_n12309_), .A2(new_n12310_), .B(\asqrt[63] ), .ZN(new_n12311_));
  INV_X1     g12119(.I(new_n12265_), .ZN(new_n12312_));
  NAND3_X1   g12120(.A1(new_n12237_), .A2(new_n327_), .A3(new_n12140_), .ZN(new_n12313_));
  AOI22_X1   g12121(.A1(new_n12313_), .A2(new_n12266_), .B1(new_n12277_), .B2(\asqrt[59] ), .ZN(new_n12314_));
  OAI21_X1   g12122(.A1(new_n12314_), .A2(new_n306_), .B(new_n218_), .ZN(new_n12315_));
  OAI21_X1   g12123(.A1(new_n12315_), .A2(new_n12279_), .B(new_n12312_), .ZN(new_n12316_));
  NOR2_X1    g12124(.A1(new_n12260_), .A2(\asqrt[62] ), .ZN(new_n12317_));
  AOI21_X1   g12125(.A1(new_n12317_), .A2(new_n12316_), .B(new_n12275_), .ZN(new_n12318_));
  INV_X1     g12126(.I(new_n12286_), .ZN(new_n12319_));
  NAND2_X1   g12127(.A1(new_n12271_), .A2(new_n12319_), .ZN(new_n12320_));
  OAI21_X1   g12128(.A1(new_n12320_), .A2(new_n12318_), .B(new_n12301_), .ZN(new_n12321_));
  OAI21_X1   g12129(.A1(new_n12311_), .A2(new_n12321_), .B(\a[40] ), .ZN(new_n12322_));
  AOI21_X1   g12130(.A1(new_n12322_), .A2(new_n12308_), .B(new_n11736_), .ZN(new_n12323_));
  INV_X1     g12131(.I(\a[40] ), .ZN(new_n12324_));
  NAND3_X1   g12132(.A1(new_n12316_), .A2(new_n207_), .A3(new_n12280_), .ZN(new_n12325_));
  AOI22_X1   g12133(.A1(new_n12325_), .A2(new_n12276_), .B1(new_n12292_), .B2(\asqrt[62] ), .ZN(new_n12326_));
  OAI21_X1   g12134(.A1(new_n12326_), .A2(new_n12289_), .B(new_n193_), .ZN(new_n12327_));
  AOI21_X1   g12135(.A1(new_n12327_), .A2(new_n12303_), .B(new_n12324_), .ZN(new_n12328_));
  NAND4_X1   g12136(.A1(new_n11798_), .A2(new_n11729_), .A3(new_n11732_), .A4(new_n12308_), .ZN(new_n12329_));
  NOR2_X1    g12137(.A1(new_n12329_), .A2(new_n11724_), .ZN(new_n12330_));
  INV_X1     g12138(.I(new_n12330_), .ZN(new_n12331_));
  NOR2_X1    g12139(.A1(new_n12328_), .A2(new_n12331_), .ZN(new_n12332_));
  AOI21_X1   g12140(.A1(new_n12327_), .A2(new_n12303_), .B(new_n11739_), .ZN(new_n12333_));
  INV_X1     g12141(.I(\a[41] ), .ZN(new_n12334_));
  AOI21_X1   g12142(.A1(\asqrt[20] ), .A2(new_n12324_), .B(new_n12334_), .ZN(new_n12335_));
  NOR3_X1    g12143(.A1(new_n12332_), .A2(new_n12335_), .A3(new_n12333_), .ZN(new_n12336_));
  OAI21_X1   g12144(.A1(new_n12336_), .A2(new_n12323_), .B(\asqrt[22] ), .ZN(new_n12337_));
  OAI21_X1   g12145(.A1(new_n12311_), .A2(new_n12321_), .B(new_n11738_), .ZN(new_n12338_));
  NAND2_X1   g12146(.A1(new_n12293_), .A2(new_n12282_), .ZN(new_n12339_));
  NOR3_X1    g12147(.A1(new_n12297_), .A2(new_n11736_), .A3(new_n12300_), .ZN(new_n12340_));
  NAND3_X1   g12148(.A1(new_n12327_), .A2(new_n12339_), .A3(new_n12340_), .ZN(new_n12341_));
  AOI21_X1   g12149(.A1(new_n12341_), .A2(new_n12338_), .B(new_n11737_), .ZN(new_n12342_));
  NAND2_X1   g12150(.A1(new_n12339_), .A2(new_n12340_), .ZN(new_n12343_));
  NOR2_X1    g12151(.A1(new_n12343_), .A2(new_n12311_), .ZN(new_n12344_));
  NOR3_X1    g12152(.A1(new_n12344_), .A2(new_n12333_), .A3(\a[42] ), .ZN(new_n12345_));
  AOI21_X1   g12153(.A1(\asqrt[20] ), .A2(\a[40] ), .B(new_n12307_), .ZN(new_n12346_));
  OAI21_X1   g12154(.A1(new_n12346_), .A2(new_n11736_), .B(new_n11326_), .ZN(new_n12347_));
  OAI22_X1   g12155(.A1(new_n12336_), .A2(new_n12347_), .B1(new_n12342_), .B2(new_n12345_), .ZN(new_n12348_));
  AOI21_X1   g12156(.A1(new_n12348_), .A2(new_n12337_), .B(new_n10812_), .ZN(new_n12349_));
  NOR3_X1    g12157(.A1(new_n11827_), .A2(new_n11828_), .A3(new_n11793_), .ZN(new_n12350_));
  NAND3_X1   g12158(.A1(\asqrt[20] ), .A2(new_n11826_), .A3(new_n11746_), .ZN(new_n12351_));
  AOI22_X1   g12159(.A1(new_n12351_), .A2(new_n11793_), .B1(\asqrt[20] ), .B2(new_n12350_), .ZN(new_n12352_));
  OAI21_X1   g12160(.A1(new_n12328_), .A2(new_n12307_), .B(\asqrt[21] ), .ZN(new_n12353_));
  AOI21_X1   g12161(.A1(new_n12327_), .A2(new_n12303_), .B(\a[40] ), .ZN(new_n12354_));
  OAI21_X1   g12162(.A1(new_n12334_), .A2(new_n12354_), .B(new_n12338_), .ZN(new_n12355_));
  OAI21_X1   g12163(.A1(new_n12355_), .A2(new_n12332_), .B(new_n12353_), .ZN(new_n12356_));
  AOI21_X1   g12164(.A1(new_n12356_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n12357_));
  AOI21_X1   g12165(.A1(new_n12357_), .A2(new_n12348_), .B(new_n12352_), .ZN(new_n12358_));
  OAI21_X1   g12166(.A1(new_n12358_), .A2(new_n12349_), .B(\asqrt[24] ), .ZN(new_n12359_));
  INV_X1     g12167(.I(new_n12359_), .ZN(new_n12360_));
  NOR2_X1    g12168(.A1(new_n11831_), .A2(new_n11834_), .ZN(new_n12361_));
  INV_X1     g12169(.I(new_n12361_), .ZN(new_n12362_));
  NAND4_X1   g12170(.A1(\asqrt[20] ), .A2(new_n11832_), .A3(new_n11806_), .A4(new_n12362_), .ZN(new_n12363_));
  INV_X1     g12171(.I(\asqrt[20] ), .ZN(new_n12364_));
  NOR3_X1    g12172(.A1(new_n12364_), .A2(new_n11795_), .A3(new_n12361_), .ZN(new_n12365_));
  OAI21_X1   g12173(.A1(new_n12365_), .A2(new_n11806_), .B(new_n12363_), .ZN(new_n12366_));
  INV_X1     g12174(.I(new_n12366_), .ZN(new_n12367_));
  NOR3_X1    g12175(.A1(new_n12358_), .A2(new_n12349_), .A3(\asqrt[24] ), .ZN(new_n12368_));
  NOR2_X1    g12176(.A1(new_n12368_), .A2(new_n12367_), .ZN(new_n12369_));
  OAI21_X1   g12177(.A1(new_n12369_), .A2(new_n12360_), .B(\asqrt[25] ), .ZN(new_n12370_));
  NAND2_X1   g12178(.A1(new_n11840_), .A2(new_n11835_), .ZN(new_n12371_));
  NAND3_X1   g12179(.A1(\asqrt[20] ), .A2(new_n11809_), .A3(new_n12371_), .ZN(new_n12372_));
  AND3_X2    g12180(.A1(new_n11809_), .A2(new_n11813_), .A3(new_n12371_), .Z(new_n12373_));
  AOI22_X1   g12181(.A1(new_n12372_), .A2(new_n11814_), .B1(\asqrt[20] ), .B2(new_n12373_), .ZN(new_n12374_));
  INV_X1     g12182(.I(new_n12374_), .ZN(new_n12375_));
  NAND2_X1   g12183(.A1(new_n12359_), .A2(new_n9846_), .ZN(new_n12376_));
  OAI21_X1   g12184(.A1(new_n12369_), .A2(new_n12376_), .B(new_n12375_), .ZN(new_n12377_));
  AOI21_X1   g12185(.A1(new_n12377_), .A2(new_n12370_), .B(new_n9317_), .ZN(new_n12378_));
  NOR3_X1    g12186(.A1(new_n11817_), .A2(new_n11823_), .A3(new_n11842_), .ZN(new_n12379_));
  NOR3_X1    g12187(.A1(new_n12364_), .A2(new_n11817_), .A3(new_n11842_), .ZN(new_n12380_));
  INV_X1     g12188(.I(new_n12380_), .ZN(new_n12381_));
  AOI22_X1   g12189(.A1(new_n12381_), .A2(new_n11823_), .B1(\asqrt[20] ), .B2(new_n12379_), .ZN(new_n12382_));
  OAI21_X1   g12190(.A1(new_n12367_), .A2(new_n12368_), .B(new_n12359_), .ZN(new_n12383_));
  AOI21_X1   g12191(.A1(new_n12383_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n12384_));
  AOI21_X1   g12192(.A1(new_n12384_), .A2(new_n12377_), .B(new_n12382_), .ZN(new_n12385_));
  OAI21_X1   g12193(.A1(new_n12385_), .A2(new_n12378_), .B(\asqrt[27] ), .ZN(new_n12386_));
  INV_X1     g12194(.I(new_n12386_), .ZN(new_n12387_));
  NAND2_X1   g12195(.A1(new_n12160_), .A2(new_n12158_), .ZN(new_n12388_));
  NAND3_X1   g12196(.A1(\asqrt[20] ), .A2(new_n11844_), .A3(new_n12388_), .ZN(new_n12389_));
  AND3_X2    g12197(.A1(new_n12388_), .A2(new_n11844_), .A3(new_n11849_), .Z(new_n12390_));
  AOI22_X1   g12198(.A1(new_n12389_), .A2(new_n11850_), .B1(\asqrt[20] ), .B2(new_n12390_), .ZN(new_n12391_));
  NOR3_X1    g12199(.A1(new_n12385_), .A2(new_n12378_), .A3(\asqrt[27] ), .ZN(new_n12392_));
  NOR2_X1    g12200(.A1(new_n12392_), .A2(new_n12391_), .ZN(new_n12393_));
  OAI21_X1   g12201(.A1(new_n12393_), .A2(new_n12387_), .B(\asqrt[28] ), .ZN(new_n12394_));
  INV_X1     g12202(.I(new_n11858_), .ZN(new_n12395_));
  NOR3_X1    g12203(.A1(new_n12171_), .A2(new_n11854_), .A3(new_n12395_), .ZN(new_n12396_));
  NOR3_X1    g12204(.A1(new_n12364_), .A2(new_n11854_), .A3(new_n12171_), .ZN(new_n12397_));
  INV_X1     g12205(.I(new_n12397_), .ZN(new_n12398_));
  AOI22_X1   g12206(.A1(new_n12398_), .A2(new_n12395_), .B1(\asqrt[20] ), .B2(new_n12396_), .ZN(new_n12399_));
  INV_X1     g12207(.I(new_n12399_), .ZN(new_n12400_));
  NAND2_X1   g12208(.A1(new_n12386_), .A2(new_n8483_), .ZN(new_n12401_));
  OAI21_X1   g12209(.A1(new_n12393_), .A2(new_n12401_), .B(new_n12400_), .ZN(new_n12402_));
  AOI21_X1   g12210(.A1(new_n12402_), .A2(new_n12394_), .B(new_n8036_), .ZN(new_n12403_));
  NOR3_X1    g12211(.A1(new_n12364_), .A2(new_n11863_), .A3(new_n11868_), .ZN(new_n12404_));
  INV_X1     g12212(.I(new_n12404_), .ZN(new_n12405_));
  NOR3_X1    g12213(.A1(new_n11863_), .A2(new_n12156_), .A3(new_n11868_), .ZN(new_n12406_));
  AOI22_X1   g12214(.A1(new_n12405_), .A2(new_n12156_), .B1(\asqrt[20] ), .B2(new_n12406_), .ZN(new_n12407_));
  OAI21_X1   g12215(.A1(new_n12391_), .A2(new_n12392_), .B(new_n12386_), .ZN(new_n12408_));
  AOI21_X1   g12216(.A1(new_n12408_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n12409_));
  AOI21_X1   g12217(.A1(new_n12409_), .A2(new_n12402_), .B(new_n12407_), .ZN(new_n12410_));
  OAI21_X1   g12218(.A1(new_n12410_), .A2(new_n12403_), .B(\asqrt[30] ), .ZN(new_n12411_));
  INV_X1     g12219(.I(new_n12411_), .ZN(new_n12412_));
  INV_X1     g12220(.I(new_n12165_), .ZN(new_n12413_));
  NOR3_X1    g12221(.A1(new_n12413_), .A2(new_n12170_), .A3(new_n11876_), .ZN(new_n12414_));
  NOR3_X1    g12222(.A1(new_n12364_), .A2(new_n12170_), .A3(new_n12413_), .ZN(new_n12415_));
  INV_X1     g12223(.I(new_n12415_), .ZN(new_n12416_));
  AOI22_X1   g12224(.A1(new_n12416_), .A2(new_n11876_), .B1(\asqrt[20] ), .B2(new_n12414_), .ZN(new_n12417_));
  NOR3_X1    g12225(.A1(new_n12410_), .A2(new_n12403_), .A3(\asqrt[30] ), .ZN(new_n12418_));
  NOR2_X1    g12226(.A1(new_n12418_), .A2(new_n12417_), .ZN(new_n12419_));
  OAI21_X1   g12227(.A1(new_n12419_), .A2(new_n12412_), .B(\asqrt[31] ), .ZN(new_n12420_));
  INV_X1     g12228(.I(new_n11883_), .ZN(new_n12421_));
  NOR3_X1    g12229(.A1(new_n12364_), .A2(new_n11879_), .A3(new_n12175_), .ZN(new_n12422_));
  INV_X1     g12230(.I(new_n12422_), .ZN(new_n12423_));
  NOR3_X1    g12231(.A1(new_n12175_), .A2(new_n11879_), .A3(new_n12421_), .ZN(new_n12424_));
  AOI22_X1   g12232(.A1(new_n12423_), .A2(new_n12421_), .B1(\asqrt[20] ), .B2(new_n12424_), .ZN(new_n12425_));
  INV_X1     g12233(.I(new_n12425_), .ZN(new_n12426_));
  NAND2_X1   g12234(.A1(new_n12411_), .A2(new_n7229_), .ZN(new_n12427_));
  OAI21_X1   g12235(.A1(new_n12419_), .A2(new_n12427_), .B(new_n12426_), .ZN(new_n12428_));
  AOI21_X1   g12236(.A1(new_n12428_), .A2(new_n12420_), .B(new_n6824_), .ZN(new_n12429_));
  NOR3_X1    g12237(.A1(new_n11888_), .A2(new_n12155_), .A3(new_n11894_), .ZN(new_n12430_));
  NOR3_X1    g12238(.A1(new_n12364_), .A2(new_n11888_), .A3(new_n11894_), .ZN(new_n12431_));
  INV_X1     g12239(.I(new_n12431_), .ZN(new_n12432_));
  AOI22_X1   g12240(.A1(new_n12432_), .A2(new_n12155_), .B1(\asqrt[20] ), .B2(new_n12430_), .ZN(new_n12433_));
  OAI21_X1   g12241(.A1(new_n12417_), .A2(new_n12418_), .B(new_n12411_), .ZN(new_n12434_));
  AOI21_X1   g12242(.A1(new_n12434_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n12435_));
  AOI21_X1   g12243(.A1(new_n12435_), .A2(new_n12428_), .B(new_n12433_), .ZN(new_n12436_));
  OAI21_X1   g12244(.A1(new_n12436_), .A2(new_n12429_), .B(\asqrt[33] ), .ZN(new_n12437_));
  INV_X1     g12245(.I(new_n12437_), .ZN(new_n12438_));
  NOR2_X1    g12246(.A1(new_n11895_), .A2(new_n11903_), .ZN(new_n12439_));
  NOR3_X1    g12247(.A1(new_n12364_), .A2(new_n12169_), .A3(new_n12439_), .ZN(new_n12440_));
  INV_X1     g12248(.I(new_n12440_), .ZN(new_n12441_));
  NOR3_X1    g12249(.A1(new_n12439_), .A2(new_n12169_), .A3(new_n11902_), .ZN(new_n12442_));
  AOI22_X1   g12250(.A1(new_n12441_), .A2(new_n11902_), .B1(\asqrt[20] ), .B2(new_n12442_), .ZN(new_n12443_));
  NOR3_X1    g12251(.A1(new_n12436_), .A2(new_n12429_), .A3(\asqrt[33] ), .ZN(new_n12444_));
  NOR2_X1    g12252(.A1(new_n12444_), .A2(new_n12443_), .ZN(new_n12445_));
  OAI21_X1   g12253(.A1(new_n12445_), .A2(new_n12438_), .B(\asqrt[34] ), .ZN(new_n12446_));
  INV_X1     g12254(.I(new_n11911_), .ZN(new_n12447_));
  NOR3_X1    g12255(.A1(new_n12183_), .A2(new_n11905_), .A3(new_n12447_), .ZN(new_n12448_));
  NOR3_X1    g12256(.A1(new_n12364_), .A2(new_n11905_), .A3(new_n12183_), .ZN(new_n12449_));
  INV_X1     g12257(.I(new_n12449_), .ZN(new_n12450_));
  AOI22_X1   g12258(.A1(new_n12450_), .A2(new_n12447_), .B1(\asqrt[20] ), .B2(new_n12448_), .ZN(new_n12451_));
  INV_X1     g12259(.I(new_n12451_), .ZN(new_n12452_));
  NAND2_X1   g12260(.A1(new_n12437_), .A2(new_n6077_), .ZN(new_n12453_));
  OAI21_X1   g12261(.A1(new_n12445_), .A2(new_n12453_), .B(new_n12452_), .ZN(new_n12454_));
  AOI21_X1   g12262(.A1(new_n12454_), .A2(new_n12446_), .B(new_n5708_), .ZN(new_n12455_));
  NOR3_X1    g12263(.A1(new_n12364_), .A2(new_n11916_), .A3(new_n11922_), .ZN(new_n12456_));
  INV_X1     g12264(.I(new_n12456_), .ZN(new_n12457_));
  NOR3_X1    g12265(.A1(new_n11916_), .A2(new_n12154_), .A3(new_n11922_), .ZN(new_n12458_));
  AOI22_X1   g12266(.A1(new_n12457_), .A2(new_n12154_), .B1(\asqrt[20] ), .B2(new_n12458_), .ZN(new_n12459_));
  OAI21_X1   g12267(.A1(new_n12443_), .A2(new_n12444_), .B(new_n12437_), .ZN(new_n12460_));
  AOI21_X1   g12268(.A1(new_n12460_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n12461_));
  AOI21_X1   g12269(.A1(new_n12461_), .A2(new_n12454_), .B(new_n12459_), .ZN(new_n12462_));
  OAI21_X1   g12270(.A1(new_n12462_), .A2(new_n12455_), .B(\asqrt[36] ), .ZN(new_n12463_));
  INV_X1     g12271(.I(new_n12463_), .ZN(new_n12464_));
  NOR2_X1    g12272(.A1(new_n11923_), .A2(new_n11931_), .ZN(new_n12465_));
  NOR3_X1    g12273(.A1(new_n12465_), .A2(new_n12182_), .A3(new_n11930_), .ZN(new_n12466_));
  NOR3_X1    g12274(.A1(new_n12364_), .A2(new_n12182_), .A3(new_n12465_), .ZN(new_n12467_));
  INV_X1     g12275(.I(new_n12467_), .ZN(new_n12468_));
  AOI22_X1   g12276(.A1(new_n12468_), .A2(new_n11930_), .B1(\asqrt[20] ), .B2(new_n12466_), .ZN(new_n12469_));
  NOR3_X1    g12277(.A1(new_n12462_), .A2(new_n12455_), .A3(\asqrt[36] ), .ZN(new_n12470_));
  NOR2_X1    g12278(.A1(new_n12470_), .A2(new_n12469_), .ZN(new_n12471_));
  OAI21_X1   g12279(.A1(new_n12471_), .A2(new_n12464_), .B(\asqrt[37] ), .ZN(new_n12472_));
  INV_X1     g12280(.I(new_n11938_), .ZN(new_n12473_));
  NOR3_X1    g12281(.A1(new_n12364_), .A2(new_n11933_), .A3(new_n12191_), .ZN(new_n12474_));
  INV_X1     g12282(.I(new_n12474_), .ZN(new_n12475_));
  NOR3_X1    g12283(.A1(new_n12191_), .A2(new_n11933_), .A3(new_n12473_), .ZN(new_n12476_));
  AOI22_X1   g12284(.A1(new_n12475_), .A2(new_n12473_), .B1(\asqrt[20] ), .B2(new_n12476_), .ZN(new_n12477_));
  INV_X1     g12285(.I(new_n12477_), .ZN(new_n12478_));
  NAND2_X1   g12286(.A1(new_n12463_), .A2(new_n5024_), .ZN(new_n12479_));
  OAI21_X1   g12287(.A1(new_n12471_), .A2(new_n12479_), .B(new_n12478_), .ZN(new_n12480_));
  AOI21_X1   g12288(.A1(new_n12480_), .A2(new_n12472_), .B(new_n4696_), .ZN(new_n12481_));
  NOR3_X1    g12289(.A1(new_n11943_), .A2(new_n12153_), .A3(new_n11949_), .ZN(new_n12482_));
  NOR3_X1    g12290(.A1(new_n12364_), .A2(new_n11943_), .A3(new_n11949_), .ZN(new_n12483_));
  INV_X1     g12291(.I(new_n12483_), .ZN(new_n12484_));
  AOI22_X1   g12292(.A1(new_n12484_), .A2(new_n12153_), .B1(\asqrt[20] ), .B2(new_n12482_), .ZN(new_n12485_));
  OAI21_X1   g12293(.A1(new_n12469_), .A2(new_n12470_), .B(new_n12463_), .ZN(new_n12486_));
  AOI21_X1   g12294(.A1(new_n12486_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n12487_));
  AOI21_X1   g12295(.A1(new_n12487_), .A2(new_n12480_), .B(new_n12485_), .ZN(new_n12488_));
  OAI21_X1   g12296(.A1(new_n12488_), .A2(new_n12481_), .B(\asqrt[39] ), .ZN(new_n12489_));
  INV_X1     g12297(.I(new_n12489_), .ZN(new_n12490_));
  NOR2_X1    g12298(.A1(new_n11950_), .A2(new_n11958_), .ZN(new_n12491_));
  NOR3_X1    g12299(.A1(new_n12364_), .A2(new_n12190_), .A3(new_n12491_), .ZN(new_n12492_));
  INV_X1     g12300(.I(new_n12492_), .ZN(new_n12493_));
  NOR3_X1    g12301(.A1(new_n12491_), .A2(new_n12190_), .A3(new_n11957_), .ZN(new_n12494_));
  AOI22_X1   g12302(.A1(new_n12493_), .A2(new_n11957_), .B1(\asqrt[20] ), .B2(new_n12494_), .ZN(new_n12495_));
  NOR3_X1    g12303(.A1(new_n12488_), .A2(new_n12481_), .A3(\asqrt[39] ), .ZN(new_n12496_));
  NOR2_X1    g12304(.A1(new_n12496_), .A2(new_n12495_), .ZN(new_n12497_));
  OAI21_X1   g12305(.A1(new_n12497_), .A2(new_n12490_), .B(\asqrt[40] ), .ZN(new_n12498_));
  INV_X1     g12306(.I(new_n11964_), .ZN(new_n12499_));
  NOR3_X1    g12307(.A1(new_n12199_), .A2(new_n11960_), .A3(new_n12499_), .ZN(new_n12500_));
  NOR3_X1    g12308(.A1(new_n12364_), .A2(new_n11960_), .A3(new_n12199_), .ZN(new_n12501_));
  INV_X1     g12309(.I(new_n12501_), .ZN(new_n12502_));
  AOI22_X1   g12310(.A1(new_n12502_), .A2(new_n12499_), .B1(\asqrt[20] ), .B2(new_n12500_), .ZN(new_n12503_));
  INV_X1     g12311(.I(new_n12503_), .ZN(new_n12504_));
  NAND2_X1   g12312(.A1(new_n12489_), .A2(new_n4071_), .ZN(new_n12505_));
  OAI21_X1   g12313(.A1(new_n12497_), .A2(new_n12505_), .B(new_n12504_), .ZN(new_n12506_));
  AOI21_X1   g12314(.A1(new_n12506_), .A2(new_n12498_), .B(new_n3782_), .ZN(new_n12507_));
  NOR3_X1    g12315(.A1(new_n12364_), .A2(new_n11969_), .A3(new_n11975_), .ZN(new_n12508_));
  INV_X1     g12316(.I(new_n12508_), .ZN(new_n12509_));
  NOR3_X1    g12317(.A1(new_n11969_), .A2(new_n12152_), .A3(new_n11975_), .ZN(new_n12510_));
  AOI22_X1   g12318(.A1(new_n12509_), .A2(new_n12152_), .B1(\asqrt[20] ), .B2(new_n12510_), .ZN(new_n12511_));
  OAI21_X1   g12319(.A1(new_n12495_), .A2(new_n12496_), .B(new_n12489_), .ZN(new_n12512_));
  AOI21_X1   g12320(.A1(new_n12512_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n12513_));
  AOI21_X1   g12321(.A1(new_n12513_), .A2(new_n12506_), .B(new_n12511_), .ZN(new_n12514_));
  OAI21_X1   g12322(.A1(new_n12514_), .A2(new_n12507_), .B(\asqrt[42] ), .ZN(new_n12515_));
  INV_X1     g12323(.I(new_n12515_), .ZN(new_n12516_));
  NOR2_X1    g12324(.A1(new_n11976_), .A2(new_n11984_), .ZN(new_n12517_));
  NOR3_X1    g12325(.A1(new_n12517_), .A2(new_n12198_), .A3(new_n11983_), .ZN(new_n12518_));
  NOR3_X1    g12326(.A1(new_n12364_), .A2(new_n12198_), .A3(new_n12517_), .ZN(new_n12519_));
  INV_X1     g12327(.I(new_n12519_), .ZN(new_n12520_));
  AOI22_X1   g12328(.A1(new_n12520_), .A2(new_n11983_), .B1(\asqrt[20] ), .B2(new_n12518_), .ZN(new_n12521_));
  NOR3_X1    g12329(.A1(new_n12514_), .A2(new_n12507_), .A3(\asqrt[42] ), .ZN(new_n12522_));
  NOR2_X1    g12330(.A1(new_n12522_), .A2(new_n12521_), .ZN(new_n12523_));
  OAI21_X1   g12331(.A1(new_n12523_), .A2(new_n12516_), .B(\asqrt[43] ), .ZN(new_n12524_));
  INV_X1     g12332(.I(new_n11990_), .ZN(new_n12525_));
  NOR3_X1    g12333(.A1(new_n12364_), .A2(new_n11986_), .A3(new_n12207_), .ZN(new_n12526_));
  INV_X1     g12334(.I(new_n12526_), .ZN(new_n12527_));
  NOR3_X1    g12335(.A1(new_n12207_), .A2(new_n11986_), .A3(new_n12525_), .ZN(new_n12528_));
  AOI22_X1   g12336(.A1(new_n12527_), .A2(new_n12525_), .B1(\asqrt[20] ), .B2(new_n12528_), .ZN(new_n12529_));
  INV_X1     g12337(.I(new_n12529_), .ZN(new_n12530_));
  NAND2_X1   g12338(.A1(new_n12515_), .A2(new_n3218_), .ZN(new_n12531_));
  OAI21_X1   g12339(.A1(new_n12523_), .A2(new_n12531_), .B(new_n12530_), .ZN(new_n12532_));
  AOI21_X1   g12340(.A1(new_n12532_), .A2(new_n12524_), .B(new_n2954_), .ZN(new_n12533_));
  NOR3_X1    g12341(.A1(new_n11995_), .A2(new_n12151_), .A3(new_n12003_), .ZN(new_n12534_));
  NOR3_X1    g12342(.A1(new_n12364_), .A2(new_n11995_), .A3(new_n12003_), .ZN(new_n12535_));
  INV_X1     g12343(.I(new_n12535_), .ZN(new_n12536_));
  AOI22_X1   g12344(.A1(new_n12536_), .A2(new_n12151_), .B1(\asqrt[20] ), .B2(new_n12534_), .ZN(new_n12537_));
  OAI21_X1   g12345(.A1(new_n12521_), .A2(new_n12522_), .B(new_n12515_), .ZN(new_n12538_));
  AOI21_X1   g12346(.A1(new_n12538_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n12539_));
  AOI21_X1   g12347(.A1(new_n12539_), .A2(new_n12532_), .B(new_n12537_), .ZN(new_n12540_));
  OAI21_X1   g12348(.A1(new_n12540_), .A2(new_n12533_), .B(\asqrt[45] ), .ZN(new_n12541_));
  INV_X1     g12349(.I(new_n12541_), .ZN(new_n12542_));
  NOR2_X1    g12350(.A1(new_n12004_), .A2(new_n12011_), .ZN(new_n12543_));
  NOR3_X1    g12351(.A1(new_n12364_), .A2(new_n12206_), .A3(new_n12543_), .ZN(new_n12544_));
  INV_X1     g12352(.I(new_n12544_), .ZN(new_n12545_));
  NOR3_X1    g12353(.A1(new_n12543_), .A2(new_n12206_), .A3(new_n12010_), .ZN(new_n12546_));
  AOI22_X1   g12354(.A1(new_n12545_), .A2(new_n12010_), .B1(\asqrt[20] ), .B2(new_n12546_), .ZN(new_n12547_));
  NOR3_X1    g12355(.A1(new_n12540_), .A2(new_n12533_), .A3(\asqrt[45] ), .ZN(new_n12548_));
  NOR2_X1    g12356(.A1(new_n12548_), .A2(new_n12547_), .ZN(new_n12549_));
  OAI21_X1   g12357(.A1(new_n12549_), .A2(new_n12542_), .B(\asqrt[46] ), .ZN(new_n12550_));
  INV_X1     g12358(.I(new_n12019_), .ZN(new_n12551_));
  NOR3_X1    g12359(.A1(new_n12215_), .A2(new_n12013_), .A3(new_n12551_), .ZN(new_n12552_));
  NOR3_X1    g12360(.A1(new_n12364_), .A2(new_n12013_), .A3(new_n12215_), .ZN(new_n12553_));
  INV_X1     g12361(.I(new_n12553_), .ZN(new_n12554_));
  AOI22_X1   g12362(.A1(new_n12554_), .A2(new_n12551_), .B1(\asqrt[20] ), .B2(new_n12552_), .ZN(new_n12555_));
  INV_X1     g12363(.I(new_n12555_), .ZN(new_n12556_));
  NAND2_X1   g12364(.A1(new_n12541_), .A2(new_n2465_), .ZN(new_n12557_));
  OAI21_X1   g12365(.A1(new_n12549_), .A2(new_n12557_), .B(new_n12556_), .ZN(new_n12558_));
  AOI21_X1   g12366(.A1(new_n12558_), .A2(new_n12550_), .B(new_n2229_), .ZN(new_n12559_));
  NOR3_X1    g12367(.A1(new_n12364_), .A2(new_n12024_), .A3(new_n12033_), .ZN(new_n12560_));
  INV_X1     g12368(.I(new_n12560_), .ZN(new_n12561_));
  NOR3_X1    g12369(.A1(new_n12024_), .A2(new_n12150_), .A3(new_n12033_), .ZN(new_n12562_));
  AOI22_X1   g12370(.A1(new_n12561_), .A2(new_n12150_), .B1(\asqrt[20] ), .B2(new_n12562_), .ZN(new_n12563_));
  OAI21_X1   g12371(.A1(new_n12547_), .A2(new_n12548_), .B(new_n12541_), .ZN(new_n12564_));
  AOI21_X1   g12372(.A1(new_n12564_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n12565_));
  AOI21_X1   g12373(.A1(new_n12565_), .A2(new_n12558_), .B(new_n12563_), .ZN(new_n12566_));
  OAI21_X1   g12374(.A1(new_n12566_), .A2(new_n12559_), .B(\asqrt[48] ), .ZN(new_n12567_));
  INV_X1     g12375(.I(new_n12567_), .ZN(new_n12568_));
  NOR2_X1    g12376(.A1(new_n12034_), .A2(new_n12041_), .ZN(new_n12569_));
  NOR3_X1    g12377(.A1(new_n12569_), .A2(new_n12214_), .A3(new_n12040_), .ZN(new_n12570_));
  NOR3_X1    g12378(.A1(new_n12364_), .A2(new_n12214_), .A3(new_n12569_), .ZN(new_n12571_));
  INV_X1     g12379(.I(new_n12571_), .ZN(new_n12572_));
  AOI22_X1   g12380(.A1(new_n12572_), .A2(new_n12040_), .B1(\asqrt[20] ), .B2(new_n12570_), .ZN(new_n12573_));
  NOR3_X1    g12381(.A1(new_n12566_), .A2(new_n12559_), .A3(\asqrt[48] ), .ZN(new_n12574_));
  NOR2_X1    g12382(.A1(new_n12574_), .A2(new_n12573_), .ZN(new_n12575_));
  OAI21_X1   g12383(.A1(new_n12575_), .A2(new_n12568_), .B(\asqrt[49] ), .ZN(new_n12576_));
  INV_X1     g12384(.I(new_n12049_), .ZN(new_n12577_));
  NOR3_X1    g12385(.A1(new_n12364_), .A2(new_n12043_), .A3(new_n12223_), .ZN(new_n12578_));
  INV_X1     g12386(.I(new_n12578_), .ZN(new_n12579_));
  NOR3_X1    g12387(.A1(new_n12223_), .A2(new_n12043_), .A3(new_n12577_), .ZN(new_n12580_));
  AOI22_X1   g12388(.A1(new_n12579_), .A2(new_n12577_), .B1(\asqrt[20] ), .B2(new_n12580_), .ZN(new_n12581_));
  INV_X1     g12389(.I(new_n12581_), .ZN(new_n12582_));
  NAND2_X1   g12390(.A1(new_n12567_), .A2(new_n1806_), .ZN(new_n12583_));
  OAI21_X1   g12391(.A1(new_n12575_), .A2(new_n12583_), .B(new_n12582_), .ZN(new_n12584_));
  AOI21_X1   g12392(.A1(new_n12584_), .A2(new_n12576_), .B(new_n1612_), .ZN(new_n12585_));
  NOR3_X1    g12393(.A1(new_n12054_), .A2(new_n12149_), .A3(new_n12063_), .ZN(new_n12586_));
  NOR3_X1    g12394(.A1(new_n12364_), .A2(new_n12054_), .A3(new_n12063_), .ZN(new_n12587_));
  INV_X1     g12395(.I(new_n12587_), .ZN(new_n12588_));
  AOI22_X1   g12396(.A1(new_n12588_), .A2(new_n12149_), .B1(\asqrt[20] ), .B2(new_n12586_), .ZN(new_n12589_));
  OAI21_X1   g12397(.A1(new_n12573_), .A2(new_n12574_), .B(new_n12567_), .ZN(new_n12590_));
  AOI21_X1   g12398(.A1(new_n12590_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n12591_));
  AOI21_X1   g12399(.A1(new_n12591_), .A2(new_n12584_), .B(new_n12589_), .ZN(new_n12592_));
  OAI21_X1   g12400(.A1(new_n12592_), .A2(new_n12585_), .B(\asqrt[51] ), .ZN(new_n12593_));
  INV_X1     g12401(.I(new_n12593_), .ZN(new_n12594_));
  NOR2_X1    g12402(.A1(new_n12064_), .A2(new_n12071_), .ZN(new_n12595_));
  NOR3_X1    g12403(.A1(new_n12364_), .A2(new_n12222_), .A3(new_n12595_), .ZN(new_n12596_));
  INV_X1     g12404(.I(new_n12596_), .ZN(new_n12597_));
  NOR3_X1    g12405(.A1(new_n12595_), .A2(new_n12222_), .A3(new_n12070_), .ZN(new_n12598_));
  AOI22_X1   g12406(.A1(new_n12597_), .A2(new_n12070_), .B1(\asqrt[20] ), .B2(new_n12598_), .ZN(new_n12599_));
  NOR3_X1    g12407(.A1(new_n12592_), .A2(new_n12585_), .A3(\asqrt[51] ), .ZN(new_n12600_));
  NOR2_X1    g12408(.A1(new_n12600_), .A2(new_n12599_), .ZN(new_n12601_));
  OAI21_X1   g12409(.A1(new_n12601_), .A2(new_n12594_), .B(\asqrt[52] ), .ZN(new_n12602_));
  INV_X1     g12410(.I(new_n12079_), .ZN(new_n12603_));
  NAND2_X1   g12411(.A1(new_n12081_), .A2(new_n12072_), .ZN(new_n12604_));
  INV_X1     g12412(.I(new_n12604_), .ZN(new_n12605_));
  NOR3_X1    g12413(.A1(new_n12605_), .A2(new_n12073_), .A3(new_n12603_), .ZN(new_n12606_));
  NOR3_X1    g12414(.A1(new_n12364_), .A2(new_n12073_), .A3(new_n12605_), .ZN(new_n12607_));
  INV_X1     g12415(.I(new_n12607_), .ZN(new_n12608_));
  AOI22_X1   g12416(.A1(new_n12608_), .A2(new_n12603_), .B1(\asqrt[20] ), .B2(new_n12606_), .ZN(new_n12609_));
  INV_X1     g12417(.I(new_n12609_), .ZN(new_n12610_));
  NAND2_X1   g12418(.A1(new_n12593_), .A2(new_n1256_), .ZN(new_n12611_));
  OAI21_X1   g12419(.A1(new_n12601_), .A2(new_n12611_), .B(new_n12610_), .ZN(new_n12612_));
  AOI21_X1   g12420(.A1(new_n12612_), .A2(new_n12602_), .B(new_n1103_), .ZN(new_n12613_));
  NOR3_X1    g12421(.A1(new_n12364_), .A2(new_n12084_), .A3(new_n12093_), .ZN(new_n12614_));
  INV_X1     g12422(.I(new_n12614_), .ZN(new_n12615_));
  NOR3_X1    g12423(.A1(new_n12084_), .A2(new_n12148_), .A3(new_n12093_), .ZN(new_n12616_));
  AOI22_X1   g12424(.A1(new_n12615_), .A2(new_n12148_), .B1(\asqrt[20] ), .B2(new_n12616_), .ZN(new_n12617_));
  OAI21_X1   g12425(.A1(new_n12599_), .A2(new_n12600_), .B(new_n12593_), .ZN(new_n12618_));
  AOI21_X1   g12426(.A1(new_n12618_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n12619_));
  AOI21_X1   g12427(.A1(new_n12619_), .A2(new_n12612_), .B(new_n12617_), .ZN(new_n12620_));
  OAI21_X1   g12428(.A1(new_n12620_), .A2(new_n12613_), .B(\asqrt[54] ), .ZN(new_n12621_));
  INV_X1     g12429(.I(new_n12621_), .ZN(new_n12622_));
  INV_X1     g12430(.I(new_n12095_), .ZN(new_n12623_));
  INV_X1     g12431(.I(new_n12230_), .ZN(new_n12624_));
  NOR3_X1    g12432(.A1(new_n12623_), .A2(new_n12624_), .A3(new_n12100_), .ZN(new_n12625_));
  NOR3_X1    g12433(.A1(new_n12364_), .A2(new_n12623_), .A3(new_n12624_), .ZN(new_n12626_));
  INV_X1     g12434(.I(new_n12626_), .ZN(new_n12627_));
  AOI22_X1   g12435(.A1(new_n12627_), .A2(new_n12100_), .B1(\asqrt[20] ), .B2(new_n12625_), .ZN(new_n12628_));
  NOR3_X1    g12436(.A1(new_n12620_), .A2(new_n12613_), .A3(\asqrt[54] ), .ZN(new_n12629_));
  NOR2_X1    g12437(.A1(new_n12629_), .A2(new_n12628_), .ZN(new_n12630_));
  OAI21_X1   g12438(.A1(new_n12630_), .A2(new_n12622_), .B(\asqrt[55] ), .ZN(new_n12631_));
  INV_X1     g12439(.I(new_n12109_), .ZN(new_n12632_));
  INV_X1     g12440(.I(new_n12102_), .ZN(new_n12633_));
  INV_X1     g12441(.I(new_n12111_), .ZN(new_n12634_));
  NOR2_X1    g12442(.A1(new_n12634_), .A2(new_n12633_), .ZN(new_n12635_));
  NOR3_X1    g12443(.A1(new_n12364_), .A2(new_n12103_), .A3(new_n12635_), .ZN(new_n12636_));
  INV_X1     g12444(.I(new_n12636_), .ZN(new_n12637_));
  NOR3_X1    g12445(.A1(new_n12635_), .A2(new_n12103_), .A3(new_n12632_), .ZN(new_n12638_));
  AOI22_X1   g12446(.A1(new_n12637_), .A2(new_n12632_), .B1(\asqrt[20] ), .B2(new_n12638_), .ZN(new_n12639_));
  INV_X1     g12447(.I(new_n12639_), .ZN(new_n12640_));
  NAND2_X1   g12448(.A1(new_n12621_), .A2(new_n823_), .ZN(new_n12641_));
  OAI21_X1   g12449(.A1(new_n12630_), .A2(new_n12641_), .B(new_n12640_), .ZN(new_n12642_));
  AOI21_X1   g12450(.A1(new_n12642_), .A2(new_n12631_), .B(new_n703_), .ZN(new_n12643_));
  NOR3_X1    g12451(.A1(new_n12114_), .A2(new_n12147_), .A3(new_n12120_), .ZN(new_n12644_));
  NOR3_X1    g12452(.A1(new_n12364_), .A2(new_n12114_), .A3(new_n12120_), .ZN(new_n12645_));
  INV_X1     g12453(.I(new_n12645_), .ZN(new_n12646_));
  AOI22_X1   g12454(.A1(new_n12646_), .A2(new_n12147_), .B1(\asqrt[20] ), .B2(new_n12644_), .ZN(new_n12647_));
  OAI21_X1   g12455(.A1(new_n12628_), .A2(new_n12629_), .B(new_n12621_), .ZN(new_n12648_));
  AOI21_X1   g12456(.A1(new_n12648_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n12649_));
  AOI21_X1   g12457(.A1(new_n12649_), .A2(new_n12642_), .B(new_n12647_), .ZN(new_n12650_));
  OAI21_X1   g12458(.A1(new_n12650_), .A2(new_n12643_), .B(\asqrt[57] ), .ZN(new_n12651_));
  INV_X1     g12459(.I(new_n12651_), .ZN(new_n12652_));
  INV_X1     g12460(.I(new_n12122_), .ZN(new_n12653_));
  INV_X1     g12461(.I(new_n12234_), .ZN(new_n12654_));
  NOR3_X1    g12462(.A1(new_n12364_), .A2(new_n12653_), .A3(new_n12654_), .ZN(new_n12655_));
  INV_X1     g12463(.I(new_n12655_), .ZN(new_n12656_));
  NOR3_X1    g12464(.A1(new_n12653_), .A2(new_n12654_), .A3(new_n12127_), .ZN(new_n12657_));
  AOI22_X1   g12465(.A1(new_n12656_), .A2(new_n12127_), .B1(\asqrt[20] ), .B2(new_n12657_), .ZN(new_n12658_));
  NOR3_X1    g12466(.A1(new_n12650_), .A2(new_n12643_), .A3(\asqrt[57] ), .ZN(new_n12659_));
  NOR2_X1    g12467(.A1(new_n12659_), .A2(new_n12658_), .ZN(new_n12660_));
  OAI21_X1   g12468(.A1(new_n12660_), .A2(new_n12652_), .B(\asqrt[58] ), .ZN(new_n12661_));
  INV_X1     g12469(.I(new_n12136_), .ZN(new_n12662_));
  INV_X1     g12470(.I(new_n12129_), .ZN(new_n12663_));
  INV_X1     g12471(.I(new_n12138_), .ZN(new_n12664_));
  OAI21_X1   g12472(.A1(new_n12664_), .A2(new_n12663_), .B(new_n12136_), .ZN(new_n12665_));
  NOR2_X1    g12473(.A1(new_n12665_), .A2(new_n12130_), .ZN(new_n12666_));
  NOR2_X1    g12474(.A1(new_n12664_), .A2(new_n12663_), .ZN(new_n12667_));
  NOR3_X1    g12475(.A1(new_n12364_), .A2(new_n12130_), .A3(new_n12667_), .ZN(new_n12668_));
  INV_X1     g12476(.I(new_n12668_), .ZN(new_n12669_));
  AOI22_X1   g12477(.A1(new_n12669_), .A2(new_n12662_), .B1(\asqrt[20] ), .B2(new_n12666_), .ZN(new_n12670_));
  INV_X1     g12478(.I(new_n12670_), .ZN(new_n12671_));
  NAND2_X1   g12479(.A1(new_n12651_), .A2(new_n436_), .ZN(new_n12672_));
  OAI21_X1   g12480(.A1(new_n12660_), .A2(new_n12672_), .B(new_n12671_), .ZN(new_n12673_));
  AOI21_X1   g12481(.A1(new_n12673_), .A2(new_n12661_), .B(new_n327_), .ZN(new_n12674_));
  NOR3_X1    g12482(.A1(new_n12364_), .A2(new_n12254_), .A3(new_n12255_), .ZN(new_n12675_));
  INV_X1     g12483(.I(new_n12675_), .ZN(new_n12676_));
  NOR3_X1    g12484(.A1(new_n12254_), .A2(new_n12146_), .A3(new_n12255_), .ZN(new_n12677_));
  AOI22_X1   g12485(.A1(new_n12676_), .A2(new_n12146_), .B1(\asqrt[20] ), .B2(new_n12677_), .ZN(new_n12678_));
  OAI21_X1   g12486(.A1(new_n12658_), .A2(new_n12659_), .B(new_n12651_), .ZN(new_n12679_));
  AOI21_X1   g12487(.A1(new_n12679_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n12680_));
  AOI21_X1   g12488(.A1(new_n12680_), .A2(new_n12673_), .B(new_n12678_), .ZN(new_n12681_));
  OAI21_X1   g12489(.A1(new_n12681_), .A2(new_n12674_), .B(\asqrt[60] ), .ZN(new_n12682_));
  INV_X1     g12490(.I(new_n12682_), .ZN(new_n12683_));
  INV_X1     g12491(.I(new_n12313_), .ZN(new_n12684_));
  NOR3_X1    g12492(.A1(new_n12684_), .A2(new_n12238_), .A3(new_n12266_), .ZN(new_n12685_));
  NOR3_X1    g12493(.A1(new_n12364_), .A2(new_n12238_), .A3(new_n12684_), .ZN(new_n12686_));
  INV_X1     g12494(.I(new_n12686_), .ZN(new_n12687_));
  AOI22_X1   g12495(.A1(new_n12687_), .A2(new_n12266_), .B1(\asqrt[20] ), .B2(new_n12685_), .ZN(new_n12688_));
  NOR3_X1    g12496(.A1(new_n12681_), .A2(new_n12674_), .A3(\asqrt[60] ), .ZN(new_n12689_));
  NOR2_X1    g12497(.A1(new_n12689_), .A2(new_n12688_), .ZN(new_n12690_));
  OAI21_X1   g12498(.A1(new_n12690_), .A2(new_n12683_), .B(\asqrt[61] ), .ZN(new_n12691_));
  NAND2_X1   g12499(.A1(new_n12278_), .A2(new_n12267_), .ZN(new_n12692_));
  NAND3_X1   g12500(.A1(\asqrt[20] ), .A2(new_n12246_), .A3(new_n12692_), .ZN(new_n12693_));
  AND3_X2    g12501(.A1(new_n12246_), .A2(new_n12252_), .A3(new_n12692_), .Z(new_n12694_));
  AOI22_X1   g12502(.A1(new_n12693_), .A2(new_n12253_), .B1(\asqrt[20] ), .B2(new_n12694_), .ZN(new_n12695_));
  INV_X1     g12503(.I(new_n12695_), .ZN(new_n12696_));
  NAND2_X1   g12504(.A1(new_n12682_), .A2(new_n218_), .ZN(new_n12697_));
  OAI21_X1   g12505(.A1(new_n12690_), .A2(new_n12697_), .B(new_n12696_), .ZN(new_n12698_));
  AOI21_X1   g12506(.A1(new_n12698_), .A2(new_n12691_), .B(new_n207_), .ZN(new_n12699_));
  NOR3_X1    g12507(.A1(new_n12260_), .A2(new_n12312_), .A3(new_n12291_), .ZN(new_n12700_));
  NOR3_X1    g12508(.A1(new_n12364_), .A2(new_n12260_), .A3(new_n12291_), .ZN(new_n12701_));
  INV_X1     g12509(.I(new_n12701_), .ZN(new_n12702_));
  AOI22_X1   g12510(.A1(new_n12702_), .A2(new_n12312_), .B1(\asqrt[20] ), .B2(new_n12700_), .ZN(new_n12703_));
  OAI21_X1   g12511(.A1(new_n12688_), .A2(new_n12689_), .B(new_n12682_), .ZN(new_n12704_));
  AOI21_X1   g12512(.A1(new_n12704_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n12705_));
  AOI21_X1   g12513(.A1(new_n12705_), .A2(new_n12698_), .B(new_n12703_), .ZN(new_n12706_));
  INV_X1     g12514(.I(new_n12271_), .ZN(new_n12707_));
  INV_X1     g12515(.I(new_n12325_), .ZN(new_n12708_));
  NOR3_X1    g12516(.A1(new_n12707_), .A2(new_n12708_), .A3(new_n12276_), .ZN(new_n12709_));
  NAND2_X1   g12517(.A1(\asqrt[20] ), .A2(new_n12709_), .ZN(new_n12710_));
  INV_X1     g12518(.I(new_n12710_), .ZN(new_n12711_));
  NOR2_X1    g12519(.A1(new_n12707_), .A2(new_n12708_), .ZN(new_n12712_));
  AOI21_X1   g12520(.A1(\asqrt[20] ), .A2(new_n12712_), .B(new_n12275_), .ZN(new_n12713_));
  NOR2_X1    g12521(.A1(new_n12711_), .A2(new_n12713_), .ZN(new_n12714_));
  INV_X1     g12522(.I(new_n12714_), .ZN(new_n12715_));
  NAND3_X1   g12523(.A1(\asqrt[20] ), .A2(new_n12309_), .A3(new_n12286_), .ZN(new_n12716_));
  AND3_X2    g12524(.A1(new_n12715_), .A2(new_n12339_), .A3(new_n12716_), .Z(new_n12717_));
  OAI21_X1   g12525(.A1(new_n12706_), .A2(new_n12699_), .B(new_n12717_), .ZN(new_n12718_));
  NAND2_X1   g12526(.A1(new_n12718_), .A2(new_n193_), .ZN(new_n12719_));
  INV_X1     g12527(.I(new_n12688_), .ZN(new_n12720_));
  INV_X1     g12528(.I(new_n12658_), .ZN(new_n12721_));
  INV_X1     g12529(.I(new_n12628_), .ZN(new_n12722_));
  INV_X1     g12530(.I(new_n12599_), .ZN(new_n12723_));
  INV_X1     g12531(.I(new_n12573_), .ZN(new_n12724_));
  INV_X1     g12532(.I(new_n12547_), .ZN(new_n12725_));
  INV_X1     g12533(.I(new_n12521_), .ZN(new_n12726_));
  INV_X1     g12534(.I(new_n12495_), .ZN(new_n12727_));
  INV_X1     g12535(.I(new_n12469_), .ZN(new_n12728_));
  INV_X1     g12536(.I(new_n12443_), .ZN(new_n12729_));
  INV_X1     g12537(.I(new_n12417_), .ZN(new_n12730_));
  INV_X1     g12538(.I(new_n12391_), .ZN(new_n12731_));
  NAND2_X1   g12539(.A1(new_n12322_), .A2(new_n12330_), .ZN(new_n12732_));
  OAI21_X1   g12540(.A1(new_n12311_), .A2(new_n12321_), .B(new_n12324_), .ZN(new_n12733_));
  NAND2_X1   g12541(.A1(new_n12733_), .A2(\a[41] ), .ZN(new_n12734_));
  NAND3_X1   g12542(.A1(new_n12732_), .A2(new_n12734_), .A3(new_n12338_), .ZN(new_n12735_));
  AOI21_X1   g12543(.A1(new_n12735_), .A2(new_n12353_), .B(new_n11326_), .ZN(new_n12736_));
  OAI21_X1   g12544(.A1(new_n12344_), .A2(new_n12333_), .B(\a[42] ), .ZN(new_n12737_));
  NAND3_X1   g12545(.A1(new_n12341_), .A2(new_n12338_), .A3(new_n11737_), .ZN(new_n12738_));
  NAND2_X1   g12546(.A1(new_n12322_), .A2(new_n12308_), .ZN(new_n12739_));
  AOI21_X1   g12547(.A1(new_n12739_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n12740_));
  AOI22_X1   g12548(.A1(new_n12735_), .A2(new_n12740_), .B1(new_n12737_), .B2(new_n12738_), .ZN(new_n12741_));
  OAI21_X1   g12549(.A1(new_n12741_), .A2(new_n12736_), .B(\asqrt[23] ), .ZN(new_n12742_));
  NAND2_X1   g12550(.A1(new_n12742_), .A2(new_n10221_), .ZN(new_n12743_));
  OAI21_X1   g12551(.A1(new_n12743_), .A2(new_n12358_), .B(new_n12366_), .ZN(new_n12744_));
  AOI21_X1   g12552(.A1(new_n12744_), .A2(new_n12359_), .B(new_n9846_), .ZN(new_n12745_));
  INV_X1     g12553(.I(new_n12352_), .ZN(new_n12746_));
  AOI21_X1   g12554(.A1(\a[41] ), .A2(new_n12733_), .B(new_n12333_), .ZN(new_n12747_));
  AOI21_X1   g12555(.A1(new_n12747_), .A2(new_n12732_), .B(new_n12323_), .ZN(new_n12748_));
  OAI21_X1   g12556(.A1(new_n12748_), .A2(new_n11326_), .B(new_n10812_), .ZN(new_n12749_));
  OAI21_X1   g12557(.A1(new_n12749_), .A2(new_n12741_), .B(new_n12746_), .ZN(new_n12750_));
  NAND2_X1   g12558(.A1(new_n12750_), .A2(new_n12742_), .ZN(new_n12751_));
  AOI21_X1   g12559(.A1(new_n12751_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n12752_));
  AOI21_X1   g12560(.A1(new_n12752_), .A2(new_n12744_), .B(new_n12374_), .ZN(new_n12753_));
  OAI21_X1   g12561(.A1(new_n12753_), .A2(new_n12745_), .B(\asqrt[26] ), .ZN(new_n12754_));
  NAND2_X1   g12562(.A1(new_n12754_), .A2(new_n8826_), .ZN(new_n12755_));
  OAI21_X1   g12563(.A1(new_n12755_), .A2(new_n12385_), .B(new_n12731_), .ZN(new_n12756_));
  NAND3_X1   g12564(.A1(new_n12756_), .A2(new_n8483_), .A3(new_n12386_), .ZN(new_n12757_));
  AOI22_X1   g12565(.A1(new_n12757_), .A2(new_n12400_), .B1(new_n12408_), .B2(\asqrt[28] ), .ZN(new_n12758_));
  OAI21_X1   g12566(.A1(new_n12758_), .A2(new_n8036_), .B(new_n7539_), .ZN(new_n12759_));
  OAI21_X1   g12567(.A1(new_n12759_), .A2(new_n12410_), .B(new_n12730_), .ZN(new_n12760_));
  AOI21_X1   g12568(.A1(new_n12760_), .A2(new_n12411_), .B(new_n7229_), .ZN(new_n12761_));
  AOI21_X1   g12569(.A1(new_n12756_), .A2(new_n12386_), .B(new_n8483_), .ZN(new_n12762_));
  NOR3_X1    g12570(.A1(new_n12753_), .A2(new_n12745_), .A3(\asqrt[26] ), .ZN(new_n12763_));
  OAI21_X1   g12571(.A1(new_n12382_), .A2(new_n12763_), .B(new_n12754_), .ZN(new_n12764_));
  AOI21_X1   g12572(.A1(new_n12764_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n12765_));
  AOI21_X1   g12573(.A1(new_n12765_), .A2(new_n12756_), .B(new_n12399_), .ZN(new_n12766_));
  NOR3_X1    g12574(.A1(new_n12766_), .A2(\asqrt[29] ), .A3(new_n12762_), .ZN(new_n12767_));
  OAI22_X1   g12575(.A1(new_n12767_), .A2(new_n12407_), .B1(new_n12758_), .B2(new_n8036_), .ZN(new_n12768_));
  AOI21_X1   g12576(.A1(new_n12768_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n12769_));
  AOI21_X1   g12577(.A1(new_n12769_), .A2(new_n12760_), .B(new_n12425_), .ZN(new_n12770_));
  OAI21_X1   g12578(.A1(new_n12770_), .A2(new_n12761_), .B(\asqrt[32] ), .ZN(new_n12771_));
  NAND2_X1   g12579(.A1(new_n12771_), .A2(new_n6356_), .ZN(new_n12772_));
  OAI21_X1   g12580(.A1(new_n12772_), .A2(new_n12436_), .B(new_n12729_), .ZN(new_n12773_));
  AOI21_X1   g12581(.A1(new_n12773_), .A2(new_n12437_), .B(new_n6077_), .ZN(new_n12774_));
  NOR3_X1    g12582(.A1(new_n12770_), .A2(\asqrt[32] ), .A3(new_n12761_), .ZN(new_n12775_));
  OAI21_X1   g12583(.A1(new_n12433_), .A2(new_n12775_), .B(new_n12771_), .ZN(new_n12776_));
  AOI21_X1   g12584(.A1(new_n12776_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n12777_));
  AOI21_X1   g12585(.A1(new_n12777_), .A2(new_n12773_), .B(new_n12451_), .ZN(new_n12778_));
  OAI21_X1   g12586(.A1(new_n12778_), .A2(new_n12774_), .B(\asqrt[35] ), .ZN(new_n12779_));
  NAND2_X1   g12587(.A1(new_n12779_), .A2(new_n5277_), .ZN(new_n12780_));
  OAI21_X1   g12588(.A1(new_n12780_), .A2(new_n12462_), .B(new_n12728_), .ZN(new_n12781_));
  AOI21_X1   g12589(.A1(new_n12781_), .A2(new_n12463_), .B(new_n5024_), .ZN(new_n12782_));
  NOR3_X1    g12590(.A1(new_n12778_), .A2(\asqrt[35] ), .A3(new_n12774_), .ZN(new_n12783_));
  OAI21_X1   g12591(.A1(new_n12459_), .A2(new_n12783_), .B(new_n12779_), .ZN(new_n12784_));
  AOI21_X1   g12592(.A1(new_n12784_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n12785_));
  AOI21_X1   g12593(.A1(new_n12785_), .A2(new_n12781_), .B(new_n12477_), .ZN(new_n12786_));
  OAI21_X1   g12594(.A1(new_n12786_), .A2(new_n12782_), .B(\asqrt[38] ), .ZN(new_n12787_));
  NAND2_X1   g12595(.A1(new_n12787_), .A2(new_n4298_), .ZN(new_n12788_));
  OAI21_X1   g12596(.A1(new_n12788_), .A2(new_n12488_), .B(new_n12727_), .ZN(new_n12789_));
  AOI21_X1   g12597(.A1(new_n12789_), .A2(new_n12489_), .B(new_n4071_), .ZN(new_n12790_));
  NOR3_X1    g12598(.A1(new_n12786_), .A2(\asqrt[38] ), .A3(new_n12782_), .ZN(new_n12791_));
  OAI21_X1   g12599(.A1(new_n12485_), .A2(new_n12791_), .B(new_n12787_), .ZN(new_n12792_));
  AOI21_X1   g12600(.A1(new_n12792_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n12793_));
  AOI21_X1   g12601(.A1(new_n12793_), .A2(new_n12789_), .B(new_n12503_), .ZN(new_n12794_));
  OAI21_X1   g12602(.A1(new_n12794_), .A2(new_n12790_), .B(\asqrt[41] ), .ZN(new_n12795_));
  NAND2_X1   g12603(.A1(new_n12795_), .A2(new_n3419_), .ZN(new_n12796_));
  OAI21_X1   g12604(.A1(new_n12796_), .A2(new_n12514_), .B(new_n12726_), .ZN(new_n12797_));
  AOI21_X1   g12605(.A1(new_n12797_), .A2(new_n12515_), .B(new_n3218_), .ZN(new_n12798_));
  NOR3_X1    g12606(.A1(new_n12794_), .A2(\asqrt[41] ), .A3(new_n12790_), .ZN(new_n12799_));
  OAI21_X1   g12607(.A1(new_n12511_), .A2(new_n12799_), .B(new_n12795_), .ZN(new_n12800_));
  AOI21_X1   g12608(.A1(new_n12800_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n12801_));
  AOI21_X1   g12609(.A1(new_n12801_), .A2(new_n12797_), .B(new_n12529_), .ZN(new_n12802_));
  OAI21_X1   g12610(.A1(new_n12802_), .A2(new_n12798_), .B(\asqrt[44] ), .ZN(new_n12803_));
  NAND2_X1   g12611(.A1(new_n12803_), .A2(new_n2641_), .ZN(new_n12804_));
  OAI21_X1   g12612(.A1(new_n12804_), .A2(new_n12540_), .B(new_n12725_), .ZN(new_n12805_));
  AOI21_X1   g12613(.A1(new_n12805_), .A2(new_n12541_), .B(new_n2465_), .ZN(new_n12806_));
  NOR3_X1    g12614(.A1(new_n12802_), .A2(\asqrt[44] ), .A3(new_n12798_), .ZN(new_n12807_));
  OAI21_X1   g12615(.A1(new_n12537_), .A2(new_n12807_), .B(new_n12803_), .ZN(new_n12808_));
  AOI21_X1   g12616(.A1(new_n12808_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n12809_));
  AOI21_X1   g12617(.A1(new_n12809_), .A2(new_n12805_), .B(new_n12555_), .ZN(new_n12810_));
  OAI21_X1   g12618(.A1(new_n12810_), .A2(new_n12806_), .B(\asqrt[47] ), .ZN(new_n12811_));
  NAND2_X1   g12619(.A1(new_n12811_), .A2(new_n1956_), .ZN(new_n12812_));
  OAI21_X1   g12620(.A1(new_n12812_), .A2(new_n12566_), .B(new_n12724_), .ZN(new_n12813_));
  AOI21_X1   g12621(.A1(new_n12813_), .A2(new_n12567_), .B(new_n1806_), .ZN(new_n12814_));
  NOR3_X1    g12622(.A1(new_n12810_), .A2(\asqrt[47] ), .A3(new_n12806_), .ZN(new_n12815_));
  OAI21_X1   g12623(.A1(new_n12563_), .A2(new_n12815_), .B(new_n12811_), .ZN(new_n12816_));
  AOI21_X1   g12624(.A1(new_n12816_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n12817_));
  AOI21_X1   g12625(.A1(new_n12817_), .A2(new_n12813_), .B(new_n12581_), .ZN(new_n12818_));
  OAI21_X1   g12626(.A1(new_n12818_), .A2(new_n12814_), .B(\asqrt[50] ), .ZN(new_n12819_));
  NAND2_X1   g12627(.A1(new_n12819_), .A2(new_n1376_), .ZN(new_n12820_));
  OAI21_X1   g12628(.A1(new_n12820_), .A2(new_n12592_), .B(new_n12723_), .ZN(new_n12821_));
  AOI21_X1   g12629(.A1(new_n12821_), .A2(new_n12593_), .B(new_n1256_), .ZN(new_n12822_));
  NOR3_X1    g12630(.A1(new_n12818_), .A2(\asqrt[50] ), .A3(new_n12814_), .ZN(new_n12823_));
  OAI21_X1   g12631(.A1(new_n12589_), .A2(new_n12823_), .B(new_n12819_), .ZN(new_n12824_));
  AOI21_X1   g12632(.A1(new_n12824_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n12825_));
  AOI21_X1   g12633(.A1(new_n12825_), .A2(new_n12821_), .B(new_n12609_), .ZN(new_n12826_));
  OAI21_X1   g12634(.A1(new_n12826_), .A2(new_n12822_), .B(\asqrt[53] ), .ZN(new_n12827_));
  NAND2_X1   g12635(.A1(new_n12827_), .A2(new_n904_), .ZN(new_n12828_));
  OAI21_X1   g12636(.A1(new_n12828_), .A2(new_n12620_), .B(new_n12722_), .ZN(new_n12829_));
  AOI21_X1   g12637(.A1(new_n12829_), .A2(new_n12621_), .B(new_n823_), .ZN(new_n12830_));
  NOR3_X1    g12638(.A1(new_n12826_), .A2(\asqrt[53] ), .A3(new_n12822_), .ZN(new_n12831_));
  OAI21_X1   g12639(.A1(new_n12617_), .A2(new_n12831_), .B(new_n12827_), .ZN(new_n12832_));
  AOI21_X1   g12640(.A1(new_n12832_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n12833_));
  AOI21_X1   g12641(.A1(new_n12833_), .A2(new_n12829_), .B(new_n12639_), .ZN(new_n12834_));
  OAI21_X1   g12642(.A1(new_n12834_), .A2(new_n12830_), .B(\asqrt[56] ), .ZN(new_n12835_));
  NAND2_X1   g12643(.A1(new_n12835_), .A2(new_n531_), .ZN(new_n12836_));
  OAI21_X1   g12644(.A1(new_n12836_), .A2(new_n12650_), .B(new_n12721_), .ZN(new_n12837_));
  AOI21_X1   g12645(.A1(new_n12837_), .A2(new_n12651_), .B(new_n436_), .ZN(new_n12838_));
  NOR3_X1    g12646(.A1(new_n12834_), .A2(\asqrt[56] ), .A3(new_n12830_), .ZN(new_n12839_));
  OAI21_X1   g12647(.A1(new_n12647_), .A2(new_n12839_), .B(new_n12835_), .ZN(new_n12840_));
  AOI21_X1   g12648(.A1(new_n12840_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n12841_));
  AOI21_X1   g12649(.A1(new_n12841_), .A2(new_n12837_), .B(new_n12670_), .ZN(new_n12842_));
  OAI21_X1   g12650(.A1(new_n12842_), .A2(new_n12838_), .B(\asqrt[59] ), .ZN(new_n12843_));
  NAND2_X1   g12651(.A1(new_n12843_), .A2(new_n306_), .ZN(new_n12844_));
  OAI21_X1   g12652(.A1(new_n12844_), .A2(new_n12681_), .B(new_n12720_), .ZN(new_n12845_));
  NOR3_X1    g12653(.A1(new_n12842_), .A2(\asqrt[59] ), .A3(new_n12838_), .ZN(new_n12846_));
  OAI21_X1   g12654(.A1(new_n12678_), .A2(new_n12846_), .B(new_n12843_), .ZN(new_n12847_));
  AOI21_X1   g12655(.A1(new_n12847_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n12848_));
  AOI21_X1   g12656(.A1(new_n12848_), .A2(new_n12845_), .B(new_n12695_), .ZN(new_n12849_));
  INV_X1     g12657(.I(new_n12703_), .ZN(new_n12850_));
  NAND2_X1   g12658(.A1(new_n12691_), .A2(new_n207_), .ZN(new_n12851_));
  OAI21_X1   g12659(.A1(new_n12851_), .A2(new_n12849_), .B(new_n12850_), .ZN(new_n12852_));
  NOR2_X1    g12660(.A1(new_n12699_), .A2(new_n12715_), .ZN(new_n12853_));
  NAND2_X1   g12661(.A1(\asqrt[20] ), .A2(new_n12286_), .ZN(new_n12854_));
  OAI21_X1   g12662(.A1(new_n12326_), .A2(new_n12319_), .B(\asqrt[63] ), .ZN(new_n12855_));
  AOI21_X1   g12663(.A1(new_n12854_), .A2(new_n12326_), .B(new_n12855_), .ZN(new_n12856_));
  AND2_X2    g12664(.A1(new_n12283_), .A2(new_n12299_), .Z(new_n12857_));
  NAND4_X1   g12665(.A1(new_n12339_), .A2(new_n12285_), .A3(new_n12296_), .A4(new_n12857_), .ZN(new_n12858_));
  NOR2_X1    g12666(.A1(new_n12858_), .A2(new_n12311_), .ZN(new_n12859_));
  NOR2_X1    g12667(.A1(new_n12856_), .A2(new_n12859_), .ZN(new_n12860_));
  INV_X1     g12668(.I(new_n12860_), .ZN(new_n12861_));
  AOI21_X1   g12669(.A1(new_n12853_), .A2(new_n12852_), .B(new_n12861_), .ZN(new_n12862_));
  NAND2_X1   g12670(.A1(new_n12719_), .A2(new_n12862_), .ZN(\asqrt[19] ));
  NOR2_X1    g12671(.A1(\a[36] ), .A2(\a[37] ), .ZN(new_n12864_));
  INV_X1     g12672(.I(new_n12864_), .ZN(new_n12865_));
  NOR2_X1    g12673(.A1(new_n12865_), .A2(\a[38] ), .ZN(new_n12866_));
  INV_X1     g12674(.I(new_n12866_), .ZN(new_n12867_));
  AOI21_X1   g12675(.A1(new_n12845_), .A2(new_n12682_), .B(new_n218_), .ZN(new_n12868_));
  OAI21_X1   g12676(.A1(new_n12849_), .A2(new_n12868_), .B(\asqrt[62] ), .ZN(new_n12869_));
  NOR3_X1    g12677(.A1(new_n12849_), .A2(\asqrt[62] ), .A3(new_n12868_), .ZN(new_n12870_));
  OAI21_X1   g12678(.A1(new_n12703_), .A2(new_n12870_), .B(new_n12869_), .ZN(new_n12871_));
  AOI21_X1   g12679(.A1(new_n12871_), .A2(new_n12717_), .B(\asqrt[63] ), .ZN(new_n12872_));
  NAND2_X1   g12680(.A1(new_n12869_), .A2(new_n12714_), .ZN(new_n12873_));
  OAI21_X1   g12681(.A1(new_n12873_), .A2(new_n12706_), .B(new_n12860_), .ZN(new_n12874_));
  OAI21_X1   g12682(.A1(new_n12872_), .A2(new_n12874_), .B(\a[38] ), .ZN(new_n12875_));
  AOI21_X1   g12683(.A1(new_n12875_), .A2(new_n12867_), .B(new_n12364_), .ZN(new_n12876_));
  INV_X1     g12684(.I(\a[38] ), .ZN(new_n12877_));
  AOI21_X1   g12685(.A1(new_n12719_), .A2(new_n12862_), .B(new_n12877_), .ZN(new_n12878_));
  NAND4_X1   g12686(.A1(new_n12339_), .A2(new_n12296_), .A3(new_n12299_), .A4(new_n12867_), .ZN(new_n12879_));
  NOR2_X1    g12687(.A1(new_n12879_), .A2(new_n12311_), .ZN(new_n12880_));
  INV_X1     g12688(.I(new_n12880_), .ZN(new_n12881_));
  NOR2_X1    g12689(.A1(new_n12878_), .A2(new_n12881_), .ZN(new_n12882_));
  AOI21_X1   g12690(.A1(new_n12719_), .A2(new_n12862_), .B(new_n12306_), .ZN(new_n12883_));
  INV_X1     g12691(.I(\a[39] ), .ZN(new_n12884_));
  AOI21_X1   g12692(.A1(\asqrt[19] ), .A2(new_n12877_), .B(new_n12884_), .ZN(new_n12885_));
  NOR3_X1    g12693(.A1(new_n12882_), .A2(new_n12885_), .A3(new_n12883_), .ZN(new_n12886_));
  OAI21_X1   g12694(.A1(new_n12886_), .A2(new_n12876_), .B(\asqrt[21] ), .ZN(new_n12887_));
  OAI21_X1   g12695(.A1(new_n12872_), .A2(new_n12874_), .B(new_n12305_), .ZN(new_n12888_));
  NAND2_X1   g12696(.A1(new_n12853_), .A2(new_n12852_), .ZN(new_n12889_));
  NOR3_X1    g12697(.A1(new_n12856_), .A2(new_n12364_), .A3(new_n12859_), .ZN(new_n12890_));
  NAND3_X1   g12698(.A1(new_n12719_), .A2(new_n12889_), .A3(new_n12890_), .ZN(new_n12891_));
  AOI21_X1   g12699(.A1(new_n12888_), .A2(new_n12891_), .B(new_n12324_), .ZN(new_n12892_));
  AND3_X2    g12700(.A1(new_n12719_), .A2(new_n12889_), .A3(new_n12890_), .Z(new_n12893_));
  NOR3_X1    g12701(.A1(new_n12893_), .A2(\a[40] ), .A3(new_n12883_), .ZN(new_n12894_));
  OAI21_X1   g12702(.A1(new_n12878_), .A2(new_n12866_), .B(\asqrt[20] ), .ZN(new_n12895_));
  NAND2_X1   g12703(.A1(new_n12895_), .A2(new_n11736_), .ZN(new_n12896_));
  OAI22_X1   g12704(.A1(new_n12886_), .A2(new_n12896_), .B1(new_n12892_), .B2(new_n12894_), .ZN(new_n12897_));
  AOI21_X1   g12705(.A1(new_n12897_), .A2(new_n12887_), .B(new_n11326_), .ZN(new_n12898_));
  NOR3_X1    g12706(.A1(new_n12747_), .A2(new_n12323_), .A3(new_n12332_), .ZN(new_n12899_));
  NAND3_X1   g12707(.A1(\asqrt[19] ), .A2(new_n12353_), .A3(new_n12732_), .ZN(new_n12900_));
  AOI22_X1   g12708(.A1(new_n12900_), .A2(new_n12747_), .B1(\asqrt[19] ), .B2(new_n12899_), .ZN(new_n12901_));
  AOI21_X1   g12709(.A1(new_n12719_), .A2(new_n12862_), .B(\a[38] ), .ZN(new_n12902_));
  OAI21_X1   g12710(.A1(new_n12884_), .A2(new_n12902_), .B(new_n12888_), .ZN(new_n12903_));
  OAI21_X1   g12711(.A1(new_n12903_), .A2(new_n12882_), .B(new_n12895_), .ZN(new_n12904_));
  AOI21_X1   g12712(.A1(new_n12904_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n12905_));
  AOI21_X1   g12713(.A1(new_n12905_), .A2(new_n12897_), .B(new_n12901_), .ZN(new_n12906_));
  OAI21_X1   g12714(.A1(new_n12906_), .A2(new_n12898_), .B(\asqrt[23] ), .ZN(new_n12907_));
  INV_X1     g12715(.I(new_n12907_), .ZN(new_n12908_));
  NOR2_X1    g12716(.A1(new_n12345_), .A2(new_n12342_), .ZN(new_n12909_));
  NOR2_X1    g12717(.A1(new_n12336_), .A2(new_n12347_), .ZN(new_n12910_));
  INV_X1     g12718(.I(new_n12910_), .ZN(new_n12911_));
  NAND4_X1   g12719(.A1(\asqrt[19] ), .A2(new_n12337_), .A3(new_n12909_), .A4(new_n12911_), .ZN(new_n12912_));
  INV_X1     g12720(.I(\asqrt[19] ), .ZN(new_n12913_));
  NOR3_X1    g12721(.A1(new_n12913_), .A2(new_n12736_), .A3(new_n12910_), .ZN(new_n12914_));
  OAI21_X1   g12722(.A1(new_n12914_), .A2(new_n12909_), .B(new_n12912_), .ZN(new_n12915_));
  INV_X1     g12723(.I(new_n12915_), .ZN(new_n12916_));
  NOR3_X1    g12724(.A1(new_n12906_), .A2(new_n12898_), .A3(\asqrt[23] ), .ZN(new_n12917_));
  NOR2_X1    g12725(.A1(new_n12917_), .A2(new_n12916_), .ZN(new_n12918_));
  OAI21_X1   g12726(.A1(new_n12918_), .A2(new_n12908_), .B(\asqrt[24] ), .ZN(new_n12919_));
  NOR2_X1    g12727(.A1(new_n12749_), .A2(new_n12741_), .ZN(new_n12920_));
  NOR3_X1    g12728(.A1(new_n12913_), .A2(new_n12349_), .A3(new_n12920_), .ZN(new_n12921_));
  INV_X1     g12729(.I(new_n12921_), .ZN(new_n12922_));
  NOR3_X1    g12730(.A1(new_n12920_), .A2(new_n12349_), .A3(new_n12746_), .ZN(new_n12923_));
  AOI22_X1   g12731(.A1(new_n12922_), .A2(new_n12746_), .B1(\asqrt[19] ), .B2(new_n12923_), .ZN(new_n12924_));
  INV_X1     g12732(.I(new_n12924_), .ZN(new_n12925_));
  NAND2_X1   g12733(.A1(new_n12907_), .A2(new_n10221_), .ZN(new_n12926_));
  OAI21_X1   g12734(.A1(new_n12918_), .A2(new_n12926_), .B(new_n12925_), .ZN(new_n12927_));
  AOI21_X1   g12735(.A1(new_n12927_), .A2(new_n12919_), .B(new_n9846_), .ZN(new_n12928_));
  NOR3_X1    g12736(.A1(new_n12360_), .A2(new_n12368_), .A3(new_n12366_), .ZN(new_n12929_));
  NOR3_X1    g12737(.A1(new_n12913_), .A2(new_n12360_), .A3(new_n12368_), .ZN(new_n12930_));
  INV_X1     g12738(.I(new_n12930_), .ZN(new_n12931_));
  AOI22_X1   g12739(.A1(new_n12931_), .A2(new_n12366_), .B1(\asqrt[19] ), .B2(new_n12929_), .ZN(new_n12932_));
  OAI21_X1   g12740(.A1(new_n12916_), .A2(new_n12917_), .B(new_n12907_), .ZN(new_n12933_));
  AOI21_X1   g12741(.A1(new_n12933_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n12934_));
  AOI21_X1   g12742(.A1(new_n12934_), .A2(new_n12927_), .B(new_n12932_), .ZN(new_n12935_));
  OAI21_X1   g12743(.A1(new_n12935_), .A2(new_n12928_), .B(\asqrt[26] ), .ZN(new_n12936_));
  NAND2_X1   g12744(.A1(new_n12752_), .A2(new_n12744_), .ZN(new_n12937_));
  NAND3_X1   g12745(.A1(\asqrt[19] ), .A2(new_n12370_), .A3(new_n12937_), .ZN(new_n12938_));
  AND3_X2    g12746(.A1(new_n12370_), .A2(new_n12374_), .A3(new_n12937_), .Z(new_n12939_));
  AOI22_X1   g12747(.A1(new_n12938_), .A2(new_n12375_), .B1(\asqrt[19] ), .B2(new_n12939_), .ZN(new_n12940_));
  INV_X1     g12748(.I(new_n12940_), .ZN(new_n12941_));
  NAND2_X1   g12749(.A1(new_n12875_), .A2(new_n12880_), .ZN(new_n12942_));
  OAI21_X1   g12750(.A1(new_n12872_), .A2(new_n12874_), .B(new_n12877_), .ZN(new_n12943_));
  NAND2_X1   g12751(.A1(new_n12943_), .A2(\a[39] ), .ZN(new_n12944_));
  NAND3_X1   g12752(.A1(new_n12942_), .A2(new_n12944_), .A3(new_n12888_), .ZN(new_n12945_));
  AOI21_X1   g12753(.A1(new_n12945_), .A2(new_n12895_), .B(new_n11736_), .ZN(new_n12946_));
  OAI21_X1   g12754(.A1(new_n12893_), .A2(new_n12883_), .B(\a[40] ), .ZN(new_n12947_));
  NAND3_X1   g12755(.A1(new_n12888_), .A2(new_n12891_), .A3(new_n12324_), .ZN(new_n12948_));
  NAND2_X1   g12756(.A1(new_n12875_), .A2(new_n12867_), .ZN(new_n12949_));
  AOI21_X1   g12757(.A1(new_n12949_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n12950_));
  AOI22_X1   g12758(.A1(new_n12945_), .A2(new_n12950_), .B1(new_n12947_), .B2(new_n12948_), .ZN(new_n12951_));
  OAI21_X1   g12759(.A1(new_n12951_), .A2(new_n12946_), .B(\asqrt[22] ), .ZN(new_n12952_));
  NAND2_X1   g12760(.A1(new_n12952_), .A2(new_n10812_), .ZN(new_n12953_));
  OAI21_X1   g12761(.A1(new_n12953_), .A2(new_n12906_), .B(new_n12915_), .ZN(new_n12954_));
  AOI21_X1   g12762(.A1(new_n12954_), .A2(new_n12907_), .B(new_n10221_), .ZN(new_n12955_));
  INV_X1     g12763(.I(new_n12901_), .ZN(new_n12956_));
  AOI21_X1   g12764(.A1(\a[39] ), .A2(new_n12943_), .B(new_n12883_), .ZN(new_n12957_));
  AOI21_X1   g12765(.A1(new_n12957_), .A2(new_n12942_), .B(new_n12876_), .ZN(new_n12958_));
  OAI21_X1   g12766(.A1(new_n12958_), .A2(new_n11736_), .B(new_n11326_), .ZN(new_n12959_));
  OAI21_X1   g12767(.A1(new_n12959_), .A2(new_n12951_), .B(new_n12956_), .ZN(new_n12960_));
  NAND2_X1   g12768(.A1(new_n12960_), .A2(new_n12952_), .ZN(new_n12961_));
  AOI21_X1   g12769(.A1(new_n12961_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n12962_));
  AOI21_X1   g12770(.A1(new_n12962_), .A2(new_n12954_), .B(new_n12924_), .ZN(new_n12963_));
  OAI21_X1   g12771(.A1(new_n12963_), .A2(new_n12955_), .B(\asqrt[25] ), .ZN(new_n12964_));
  NAND2_X1   g12772(.A1(new_n12964_), .A2(new_n9317_), .ZN(new_n12965_));
  OAI21_X1   g12773(.A1(new_n12965_), .A2(new_n12935_), .B(new_n12941_), .ZN(new_n12966_));
  AOI21_X1   g12774(.A1(new_n12966_), .A2(new_n12936_), .B(new_n8826_), .ZN(new_n12967_));
  INV_X1     g12775(.I(new_n12382_), .ZN(new_n12968_));
  NOR3_X1    g12776(.A1(new_n12378_), .A2(new_n12763_), .A3(new_n12968_), .ZN(new_n12969_));
  NOR3_X1    g12777(.A1(new_n12913_), .A2(new_n12378_), .A3(new_n12763_), .ZN(new_n12970_));
  INV_X1     g12778(.I(new_n12970_), .ZN(new_n12971_));
  AOI22_X1   g12779(.A1(new_n12971_), .A2(new_n12968_), .B1(\asqrt[19] ), .B2(new_n12969_), .ZN(new_n12972_));
  NOR3_X1    g12780(.A1(new_n12963_), .A2(new_n12955_), .A3(\asqrt[25] ), .ZN(new_n12973_));
  OAI21_X1   g12781(.A1(new_n12932_), .A2(new_n12973_), .B(new_n12964_), .ZN(new_n12974_));
  AOI21_X1   g12782(.A1(new_n12974_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n12975_));
  AOI21_X1   g12783(.A1(new_n12975_), .A2(new_n12966_), .B(new_n12972_), .ZN(new_n12976_));
  OAI21_X1   g12784(.A1(new_n12976_), .A2(new_n12967_), .B(\asqrt[28] ), .ZN(new_n12977_));
  INV_X1     g12785(.I(new_n12977_), .ZN(new_n12978_));
  INV_X1     g12786(.I(new_n12972_), .ZN(new_n12979_));
  NAND3_X1   g12787(.A1(new_n12966_), .A2(new_n8826_), .A3(new_n12936_), .ZN(new_n12980_));
  NAND2_X1   g12788(.A1(new_n12980_), .A2(new_n12979_), .ZN(new_n12981_));
  NOR3_X1    g12789(.A1(new_n12913_), .A2(new_n12387_), .A3(new_n12392_), .ZN(new_n12982_));
  INV_X1     g12790(.I(new_n12982_), .ZN(new_n12983_));
  NOR3_X1    g12791(.A1(new_n12387_), .A2(new_n12731_), .A3(new_n12392_), .ZN(new_n12984_));
  AOI22_X1   g12792(.A1(new_n12983_), .A2(new_n12731_), .B1(\asqrt[19] ), .B2(new_n12984_), .ZN(new_n12985_));
  NOR2_X1    g12793(.A1(new_n12967_), .A2(\asqrt[28] ), .ZN(new_n12986_));
  AOI21_X1   g12794(.A1(new_n12986_), .A2(new_n12981_), .B(new_n12985_), .ZN(new_n12987_));
  OAI21_X1   g12795(.A1(new_n12978_), .A2(new_n12987_), .B(\asqrt[29] ), .ZN(new_n12988_));
  AND3_X2    g12796(.A1(new_n12394_), .A2(new_n12399_), .A3(new_n12757_), .Z(new_n12989_));
  NAND3_X1   g12797(.A1(\asqrt[19] ), .A2(new_n12394_), .A3(new_n12757_), .ZN(new_n12990_));
  AOI22_X1   g12798(.A1(new_n12990_), .A2(new_n12400_), .B1(\asqrt[19] ), .B2(new_n12989_), .ZN(new_n12991_));
  INV_X1     g12799(.I(new_n12991_), .ZN(new_n12992_));
  NAND2_X1   g12800(.A1(new_n12977_), .A2(new_n8036_), .ZN(new_n12993_));
  OAI21_X1   g12801(.A1(new_n12993_), .A2(new_n12987_), .B(new_n12992_), .ZN(new_n12994_));
  AOI21_X1   g12802(.A1(new_n12994_), .A2(new_n12988_), .B(new_n7539_), .ZN(new_n12995_));
  INV_X1     g12803(.I(new_n12995_), .ZN(new_n12996_));
  INV_X1     g12804(.I(new_n12994_), .ZN(new_n12997_));
  INV_X1     g12805(.I(new_n12407_), .ZN(new_n12998_));
  NOR3_X1    g12806(.A1(new_n12913_), .A2(new_n12403_), .A3(new_n12767_), .ZN(new_n12999_));
  INV_X1     g12807(.I(new_n12999_), .ZN(new_n13000_));
  NOR3_X1    g12808(.A1(new_n12403_), .A2(new_n12767_), .A3(new_n12998_), .ZN(new_n13001_));
  AOI22_X1   g12809(.A1(new_n13000_), .A2(new_n12998_), .B1(\asqrt[19] ), .B2(new_n13001_), .ZN(new_n13002_));
  INV_X1     g12810(.I(new_n13002_), .ZN(new_n13003_));
  NAND2_X1   g12811(.A1(new_n12988_), .A2(new_n7539_), .ZN(new_n13004_));
  OAI21_X1   g12812(.A1(new_n13004_), .A2(new_n12997_), .B(new_n13003_), .ZN(new_n13005_));
  AOI21_X1   g12813(.A1(new_n13005_), .A2(new_n12996_), .B(new_n7229_), .ZN(new_n13006_));
  NOR3_X1    g12814(.A1(new_n12412_), .A2(new_n12730_), .A3(new_n12418_), .ZN(new_n13007_));
  NOR3_X1    g12815(.A1(new_n12913_), .A2(new_n12412_), .A3(new_n12418_), .ZN(new_n13008_));
  INV_X1     g12816(.I(new_n13008_), .ZN(new_n13009_));
  AOI22_X1   g12817(.A1(new_n13009_), .A2(new_n12730_), .B1(\asqrt[19] ), .B2(new_n13007_), .ZN(new_n13010_));
  NOR2_X1    g12818(.A1(new_n12995_), .A2(\asqrt[31] ), .ZN(new_n13011_));
  AOI21_X1   g12819(.A1(new_n13011_), .A2(new_n13005_), .B(new_n13010_), .ZN(new_n13012_));
  OAI21_X1   g12820(.A1(new_n13012_), .A2(new_n13006_), .B(\asqrt[32] ), .ZN(new_n13013_));
  NOR2_X1    g12821(.A1(new_n12419_), .A2(new_n12427_), .ZN(new_n13014_));
  NOR3_X1    g12822(.A1(new_n12913_), .A2(new_n12761_), .A3(new_n13014_), .ZN(new_n13015_));
  INV_X1     g12823(.I(new_n13015_), .ZN(new_n13016_));
  NOR3_X1    g12824(.A1(new_n13014_), .A2(new_n12761_), .A3(new_n12426_), .ZN(new_n13017_));
  AOI22_X1   g12825(.A1(new_n13016_), .A2(new_n12426_), .B1(\asqrt[19] ), .B2(new_n13017_), .ZN(new_n13018_));
  INV_X1     g12826(.I(new_n13018_), .ZN(new_n13019_));
  NOR3_X1    g12827(.A1(new_n12935_), .A2(new_n12928_), .A3(\asqrt[26] ), .ZN(new_n13020_));
  OAI21_X1   g12828(.A1(new_n12940_), .A2(new_n13020_), .B(new_n12936_), .ZN(new_n13021_));
  AOI22_X1   g12829(.A1(new_n12980_), .A2(new_n12979_), .B1(new_n13021_), .B2(\asqrt[27] ), .ZN(new_n13022_));
  NOR3_X1    g12830(.A1(new_n12976_), .A2(\asqrt[28] ), .A3(new_n12967_), .ZN(new_n13023_));
  OAI22_X1   g12831(.A1(new_n13023_), .A2(new_n12985_), .B1(new_n13022_), .B2(new_n8483_), .ZN(new_n13024_));
  AOI21_X1   g12832(.A1(new_n13024_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n13025_));
  AOI21_X1   g12833(.A1(new_n13025_), .A2(new_n12994_), .B(new_n13002_), .ZN(new_n13026_));
  OAI21_X1   g12834(.A1(new_n13026_), .A2(new_n12995_), .B(\asqrt[31] ), .ZN(new_n13027_));
  NAND2_X1   g12835(.A1(new_n13027_), .A2(new_n6824_), .ZN(new_n13028_));
  OAI21_X1   g12836(.A1(new_n13028_), .A2(new_n13012_), .B(new_n13019_), .ZN(new_n13029_));
  AOI21_X1   g12837(.A1(new_n13029_), .A2(new_n13013_), .B(new_n6356_), .ZN(new_n13030_));
  INV_X1     g12838(.I(new_n13030_), .ZN(new_n13031_));
  INV_X1     g12839(.I(new_n13029_), .ZN(new_n13032_));
  INV_X1     g12840(.I(new_n12433_), .ZN(new_n13033_));
  NOR3_X1    g12841(.A1(new_n12429_), .A2(new_n12775_), .A3(new_n13033_), .ZN(new_n13034_));
  NOR3_X1    g12842(.A1(new_n12913_), .A2(new_n12429_), .A3(new_n12775_), .ZN(new_n13035_));
  INV_X1     g12843(.I(new_n13035_), .ZN(new_n13036_));
  AOI22_X1   g12844(.A1(new_n13036_), .A2(new_n13033_), .B1(\asqrt[19] ), .B2(new_n13034_), .ZN(new_n13037_));
  INV_X1     g12845(.I(new_n13037_), .ZN(new_n13038_));
  NAND2_X1   g12846(.A1(new_n13013_), .A2(new_n6356_), .ZN(new_n13039_));
  OAI21_X1   g12847(.A1(new_n13032_), .A2(new_n13039_), .B(new_n13038_), .ZN(new_n13040_));
  AOI21_X1   g12848(.A1(new_n13040_), .A2(new_n13031_), .B(new_n6077_), .ZN(new_n13041_));
  NOR3_X1    g12849(.A1(new_n12913_), .A2(new_n12438_), .A3(new_n12444_), .ZN(new_n13042_));
  INV_X1     g12850(.I(new_n13042_), .ZN(new_n13043_));
  NOR3_X1    g12851(.A1(new_n12438_), .A2(new_n12729_), .A3(new_n12444_), .ZN(new_n13044_));
  AOI22_X1   g12852(.A1(new_n13043_), .A2(new_n12729_), .B1(\asqrt[19] ), .B2(new_n13044_), .ZN(new_n13045_));
  NOR2_X1    g12853(.A1(new_n13030_), .A2(\asqrt[34] ), .ZN(new_n13046_));
  AOI21_X1   g12854(.A1(new_n13046_), .A2(new_n13040_), .B(new_n13045_), .ZN(new_n13047_));
  OAI21_X1   g12855(.A1(new_n13047_), .A2(new_n13041_), .B(\asqrt[35] ), .ZN(new_n13048_));
  NOR2_X1    g12856(.A1(new_n12445_), .A2(new_n12453_), .ZN(new_n13049_));
  NOR3_X1    g12857(.A1(new_n13049_), .A2(new_n12774_), .A3(new_n12452_), .ZN(new_n13050_));
  NOR3_X1    g12858(.A1(new_n12913_), .A2(new_n12774_), .A3(new_n13049_), .ZN(new_n13051_));
  INV_X1     g12859(.I(new_n13051_), .ZN(new_n13052_));
  AOI22_X1   g12860(.A1(new_n13052_), .A2(new_n12452_), .B1(\asqrt[19] ), .B2(new_n13050_), .ZN(new_n13053_));
  INV_X1     g12861(.I(new_n13053_), .ZN(new_n13054_));
  NOR3_X1    g12862(.A1(new_n13026_), .A2(\asqrt[31] ), .A3(new_n12995_), .ZN(new_n13055_));
  OAI21_X1   g12863(.A1(new_n13010_), .A2(new_n13055_), .B(new_n13027_), .ZN(new_n13056_));
  AOI21_X1   g12864(.A1(new_n13056_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n13057_));
  AOI21_X1   g12865(.A1(new_n13057_), .A2(new_n13029_), .B(new_n13037_), .ZN(new_n13058_));
  OAI21_X1   g12866(.A1(new_n13058_), .A2(new_n13030_), .B(\asqrt[34] ), .ZN(new_n13059_));
  NAND2_X1   g12867(.A1(new_n13059_), .A2(new_n5708_), .ZN(new_n13060_));
  OAI21_X1   g12868(.A1(new_n13060_), .A2(new_n13047_), .B(new_n13054_), .ZN(new_n13061_));
  NAND2_X1   g12869(.A1(new_n13061_), .A2(new_n13048_), .ZN(new_n13062_));
  NAND2_X1   g12870(.A1(new_n13062_), .A2(\asqrt[36] ), .ZN(new_n13063_));
  INV_X1     g12871(.I(new_n13061_), .ZN(new_n13064_));
  INV_X1     g12872(.I(new_n12459_), .ZN(new_n13065_));
  NOR3_X1    g12873(.A1(new_n12913_), .A2(new_n12455_), .A3(new_n12783_), .ZN(new_n13066_));
  INV_X1     g12874(.I(new_n13066_), .ZN(new_n13067_));
  NOR3_X1    g12875(.A1(new_n12455_), .A2(new_n12783_), .A3(new_n13065_), .ZN(new_n13068_));
  AOI22_X1   g12876(.A1(new_n13067_), .A2(new_n13065_), .B1(\asqrt[19] ), .B2(new_n13068_), .ZN(new_n13069_));
  INV_X1     g12877(.I(new_n13069_), .ZN(new_n13070_));
  NAND2_X1   g12878(.A1(new_n13048_), .A2(new_n5277_), .ZN(new_n13071_));
  OAI21_X1   g12879(.A1(new_n13064_), .A2(new_n13071_), .B(new_n13070_), .ZN(new_n13072_));
  AOI21_X1   g12880(.A1(new_n13072_), .A2(new_n13063_), .B(new_n5024_), .ZN(new_n13073_));
  NOR3_X1    g12881(.A1(new_n12464_), .A2(new_n12728_), .A3(new_n12470_), .ZN(new_n13074_));
  NOR3_X1    g12882(.A1(new_n12913_), .A2(new_n12464_), .A3(new_n12470_), .ZN(new_n13075_));
  INV_X1     g12883(.I(new_n13075_), .ZN(new_n13076_));
  AOI22_X1   g12884(.A1(new_n13076_), .A2(new_n12728_), .B1(\asqrt[19] ), .B2(new_n13074_), .ZN(new_n13077_));
  AOI21_X1   g12885(.A1(new_n13061_), .A2(new_n13048_), .B(new_n5277_), .ZN(new_n13078_));
  NOR2_X1    g12886(.A1(new_n13078_), .A2(\asqrt[37] ), .ZN(new_n13079_));
  AOI21_X1   g12887(.A1(new_n13079_), .A2(new_n13072_), .B(new_n13077_), .ZN(new_n13080_));
  OAI21_X1   g12888(.A1(new_n13080_), .A2(new_n13073_), .B(\asqrt[38] ), .ZN(new_n13081_));
  INV_X1     g12889(.I(new_n13081_), .ZN(new_n13082_));
  NOR2_X1    g12890(.A1(new_n12471_), .A2(new_n12479_), .ZN(new_n13083_));
  NOR3_X1    g12891(.A1(new_n12913_), .A2(new_n12782_), .A3(new_n13083_), .ZN(new_n13084_));
  INV_X1     g12892(.I(new_n13084_), .ZN(new_n13085_));
  NOR3_X1    g12893(.A1(new_n13083_), .A2(new_n12782_), .A3(new_n12478_), .ZN(new_n13086_));
  AOI22_X1   g12894(.A1(new_n13085_), .A2(new_n12478_), .B1(\asqrt[19] ), .B2(new_n13086_), .ZN(new_n13087_));
  NOR3_X1    g12895(.A1(new_n13080_), .A2(new_n13073_), .A3(\asqrt[38] ), .ZN(new_n13088_));
  NOR2_X1    g12896(.A1(new_n13088_), .A2(new_n13087_), .ZN(new_n13089_));
  OAI21_X1   g12897(.A1(new_n13089_), .A2(new_n13082_), .B(\asqrt[39] ), .ZN(new_n13090_));
  INV_X1     g12898(.I(new_n12485_), .ZN(new_n13091_));
  NOR3_X1    g12899(.A1(new_n12481_), .A2(new_n12791_), .A3(new_n13091_), .ZN(new_n13092_));
  NOR3_X1    g12900(.A1(new_n12913_), .A2(new_n12481_), .A3(new_n12791_), .ZN(new_n13093_));
  INV_X1     g12901(.I(new_n13093_), .ZN(new_n13094_));
  AOI22_X1   g12902(.A1(new_n13094_), .A2(new_n13091_), .B1(\asqrt[19] ), .B2(new_n13092_), .ZN(new_n13095_));
  INV_X1     g12903(.I(new_n13095_), .ZN(new_n13096_));
  NAND2_X1   g12904(.A1(new_n13081_), .A2(new_n4298_), .ZN(new_n13097_));
  OAI21_X1   g12905(.A1(new_n13089_), .A2(new_n13097_), .B(new_n13096_), .ZN(new_n13098_));
  AOI21_X1   g12906(.A1(new_n13098_), .A2(new_n13090_), .B(new_n4071_), .ZN(new_n13099_));
  NOR3_X1    g12907(.A1(new_n12913_), .A2(new_n12490_), .A3(new_n12496_), .ZN(new_n13100_));
  INV_X1     g12908(.I(new_n13100_), .ZN(new_n13101_));
  NOR3_X1    g12909(.A1(new_n12490_), .A2(new_n12727_), .A3(new_n12496_), .ZN(new_n13102_));
  AOI22_X1   g12910(.A1(new_n13101_), .A2(new_n12727_), .B1(\asqrt[19] ), .B2(new_n13102_), .ZN(new_n13103_));
  INV_X1     g12911(.I(new_n13087_), .ZN(new_n13104_));
  NOR3_X1    g12912(.A1(new_n13058_), .A2(\asqrt[34] ), .A3(new_n13030_), .ZN(new_n13105_));
  OAI21_X1   g12913(.A1(new_n13045_), .A2(new_n13105_), .B(new_n13059_), .ZN(new_n13106_));
  AOI21_X1   g12914(.A1(new_n13106_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n13107_));
  AOI21_X1   g12915(.A1(new_n13107_), .A2(new_n13061_), .B(new_n13069_), .ZN(new_n13108_));
  OAI21_X1   g12916(.A1(new_n13108_), .A2(new_n13078_), .B(\asqrt[37] ), .ZN(new_n13109_));
  NAND2_X1   g12917(.A1(new_n13109_), .A2(new_n4696_), .ZN(new_n13110_));
  OAI21_X1   g12918(.A1(new_n13110_), .A2(new_n13080_), .B(new_n13104_), .ZN(new_n13111_));
  AOI21_X1   g12919(.A1(new_n13111_), .A2(new_n13081_), .B(new_n4298_), .ZN(new_n13112_));
  NOR2_X1    g12920(.A1(new_n13112_), .A2(\asqrt[40] ), .ZN(new_n13113_));
  AOI21_X1   g12921(.A1(new_n13113_), .A2(new_n13098_), .B(new_n13103_), .ZN(new_n13114_));
  OAI21_X1   g12922(.A1(new_n13114_), .A2(new_n13099_), .B(\asqrt[41] ), .ZN(new_n13115_));
  NOR2_X1    g12923(.A1(new_n12497_), .A2(new_n12505_), .ZN(new_n13116_));
  NOR3_X1    g12924(.A1(new_n13116_), .A2(new_n12790_), .A3(new_n12504_), .ZN(new_n13117_));
  NOR3_X1    g12925(.A1(new_n12913_), .A2(new_n12790_), .A3(new_n13116_), .ZN(new_n13118_));
  INV_X1     g12926(.I(new_n13118_), .ZN(new_n13119_));
  AOI22_X1   g12927(.A1(new_n13119_), .A2(new_n12504_), .B1(\asqrt[19] ), .B2(new_n13117_), .ZN(new_n13120_));
  INV_X1     g12928(.I(new_n13120_), .ZN(new_n13121_));
  NOR3_X1    g12929(.A1(new_n13108_), .A2(\asqrt[37] ), .A3(new_n13078_), .ZN(new_n13122_));
  OAI21_X1   g12930(.A1(new_n13077_), .A2(new_n13122_), .B(new_n13109_), .ZN(new_n13123_));
  AOI21_X1   g12931(.A1(new_n13123_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n13124_));
  AOI21_X1   g12932(.A1(new_n13124_), .A2(new_n13111_), .B(new_n13095_), .ZN(new_n13125_));
  OAI21_X1   g12933(.A1(new_n13125_), .A2(new_n13112_), .B(\asqrt[40] ), .ZN(new_n13126_));
  NAND2_X1   g12934(.A1(new_n13126_), .A2(new_n3782_), .ZN(new_n13127_));
  OAI21_X1   g12935(.A1(new_n13127_), .A2(new_n13114_), .B(new_n13121_), .ZN(new_n13128_));
  AOI21_X1   g12936(.A1(new_n13128_), .A2(new_n13115_), .B(new_n3419_), .ZN(new_n13129_));
  INV_X1     g12937(.I(new_n12511_), .ZN(new_n13130_));
  NOR3_X1    g12938(.A1(new_n12913_), .A2(new_n12507_), .A3(new_n12799_), .ZN(new_n13131_));
  INV_X1     g12939(.I(new_n13131_), .ZN(new_n13132_));
  NOR3_X1    g12940(.A1(new_n12507_), .A2(new_n12799_), .A3(new_n13130_), .ZN(new_n13133_));
  AOI22_X1   g12941(.A1(new_n13132_), .A2(new_n13130_), .B1(\asqrt[19] ), .B2(new_n13133_), .ZN(new_n13134_));
  NOR3_X1    g12942(.A1(new_n13125_), .A2(\asqrt[40] ), .A3(new_n13112_), .ZN(new_n13135_));
  OAI21_X1   g12943(.A1(new_n13103_), .A2(new_n13135_), .B(new_n13126_), .ZN(new_n13136_));
  AOI21_X1   g12944(.A1(new_n13136_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n13137_));
  AOI21_X1   g12945(.A1(new_n13137_), .A2(new_n13128_), .B(new_n13134_), .ZN(new_n13138_));
  OAI21_X1   g12946(.A1(new_n13138_), .A2(new_n13129_), .B(\asqrt[43] ), .ZN(new_n13139_));
  INV_X1     g12947(.I(new_n13139_), .ZN(new_n13140_));
  NOR3_X1    g12948(.A1(new_n12516_), .A2(new_n12726_), .A3(new_n12522_), .ZN(new_n13141_));
  NOR3_X1    g12949(.A1(new_n12913_), .A2(new_n12516_), .A3(new_n12522_), .ZN(new_n13142_));
  INV_X1     g12950(.I(new_n13142_), .ZN(new_n13143_));
  AOI22_X1   g12951(.A1(new_n13143_), .A2(new_n12726_), .B1(\asqrt[19] ), .B2(new_n13141_), .ZN(new_n13144_));
  NOR3_X1    g12952(.A1(new_n13138_), .A2(\asqrt[43] ), .A3(new_n13129_), .ZN(new_n13145_));
  NOR2_X1    g12953(.A1(new_n13145_), .A2(new_n13144_), .ZN(new_n13146_));
  OAI21_X1   g12954(.A1(new_n13146_), .A2(new_n13140_), .B(\asqrt[44] ), .ZN(new_n13147_));
  NOR2_X1    g12955(.A1(new_n12523_), .A2(new_n12531_), .ZN(new_n13148_));
  NOR3_X1    g12956(.A1(new_n12913_), .A2(new_n12798_), .A3(new_n13148_), .ZN(new_n13149_));
  INV_X1     g12957(.I(new_n13149_), .ZN(new_n13150_));
  NOR3_X1    g12958(.A1(new_n13148_), .A2(new_n12798_), .A3(new_n12530_), .ZN(new_n13151_));
  AOI22_X1   g12959(.A1(new_n13150_), .A2(new_n12530_), .B1(\asqrt[19] ), .B2(new_n13151_), .ZN(new_n13152_));
  INV_X1     g12960(.I(new_n13152_), .ZN(new_n13153_));
  NAND2_X1   g12961(.A1(new_n13139_), .A2(new_n2954_), .ZN(new_n13154_));
  OAI21_X1   g12962(.A1(new_n13146_), .A2(new_n13154_), .B(new_n13153_), .ZN(new_n13155_));
  AOI21_X1   g12963(.A1(new_n13155_), .A2(new_n13147_), .B(new_n2641_), .ZN(new_n13156_));
  INV_X1     g12964(.I(new_n12537_), .ZN(new_n13157_));
  NOR3_X1    g12965(.A1(new_n12533_), .A2(new_n12807_), .A3(new_n13157_), .ZN(new_n13158_));
  NOR3_X1    g12966(.A1(new_n12913_), .A2(new_n12533_), .A3(new_n12807_), .ZN(new_n13159_));
  INV_X1     g12967(.I(new_n13159_), .ZN(new_n13160_));
  AOI22_X1   g12968(.A1(new_n13160_), .A2(new_n13157_), .B1(\asqrt[19] ), .B2(new_n13158_), .ZN(new_n13161_));
  OAI21_X1   g12969(.A1(new_n13144_), .A2(new_n13145_), .B(new_n13139_), .ZN(new_n13162_));
  AOI21_X1   g12970(.A1(new_n13162_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n13163_));
  AOI21_X1   g12971(.A1(new_n13163_), .A2(new_n13155_), .B(new_n13161_), .ZN(new_n13164_));
  OAI21_X1   g12972(.A1(new_n13164_), .A2(new_n13156_), .B(\asqrt[46] ), .ZN(new_n13165_));
  INV_X1     g12973(.I(new_n13165_), .ZN(new_n13166_));
  NOR3_X1    g12974(.A1(new_n12913_), .A2(new_n12542_), .A3(new_n12548_), .ZN(new_n13167_));
  INV_X1     g12975(.I(new_n13167_), .ZN(new_n13168_));
  NOR3_X1    g12976(.A1(new_n12542_), .A2(new_n12725_), .A3(new_n12548_), .ZN(new_n13169_));
  AOI22_X1   g12977(.A1(new_n13168_), .A2(new_n12725_), .B1(\asqrt[19] ), .B2(new_n13169_), .ZN(new_n13170_));
  NOR3_X1    g12978(.A1(new_n13164_), .A2(new_n13156_), .A3(\asqrt[46] ), .ZN(new_n13171_));
  NOR2_X1    g12979(.A1(new_n13171_), .A2(new_n13170_), .ZN(new_n13172_));
  OAI21_X1   g12980(.A1(new_n13172_), .A2(new_n13166_), .B(\asqrt[47] ), .ZN(new_n13173_));
  NOR2_X1    g12981(.A1(new_n12549_), .A2(new_n12557_), .ZN(new_n13174_));
  NOR3_X1    g12982(.A1(new_n13174_), .A2(new_n12806_), .A3(new_n12556_), .ZN(new_n13175_));
  NOR3_X1    g12983(.A1(new_n12913_), .A2(new_n12806_), .A3(new_n13174_), .ZN(new_n13176_));
  INV_X1     g12984(.I(new_n13176_), .ZN(new_n13177_));
  AOI22_X1   g12985(.A1(new_n13177_), .A2(new_n12556_), .B1(\asqrt[19] ), .B2(new_n13175_), .ZN(new_n13178_));
  INV_X1     g12986(.I(new_n13178_), .ZN(new_n13179_));
  NAND2_X1   g12987(.A1(new_n13165_), .A2(new_n2229_), .ZN(new_n13180_));
  OAI21_X1   g12988(.A1(new_n13172_), .A2(new_n13180_), .B(new_n13179_), .ZN(new_n13181_));
  AOI21_X1   g12989(.A1(new_n13181_), .A2(new_n13173_), .B(new_n1956_), .ZN(new_n13182_));
  INV_X1     g12990(.I(new_n12563_), .ZN(new_n13183_));
  NOR3_X1    g12991(.A1(new_n12913_), .A2(new_n12559_), .A3(new_n12815_), .ZN(new_n13184_));
  INV_X1     g12992(.I(new_n13184_), .ZN(new_n13185_));
  NOR3_X1    g12993(.A1(new_n12559_), .A2(new_n12815_), .A3(new_n13183_), .ZN(new_n13186_));
  AOI22_X1   g12994(.A1(new_n13185_), .A2(new_n13183_), .B1(\asqrt[19] ), .B2(new_n13186_), .ZN(new_n13187_));
  OAI21_X1   g12995(.A1(new_n13170_), .A2(new_n13171_), .B(new_n13165_), .ZN(new_n13188_));
  AOI21_X1   g12996(.A1(new_n13188_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n13189_));
  AOI21_X1   g12997(.A1(new_n13189_), .A2(new_n13181_), .B(new_n13187_), .ZN(new_n13190_));
  OAI21_X1   g12998(.A1(new_n13190_), .A2(new_n13182_), .B(\asqrt[49] ), .ZN(new_n13191_));
  INV_X1     g12999(.I(new_n13191_), .ZN(new_n13192_));
  NOR3_X1    g13000(.A1(new_n12568_), .A2(new_n12724_), .A3(new_n12574_), .ZN(new_n13193_));
  NOR3_X1    g13001(.A1(new_n12913_), .A2(new_n12568_), .A3(new_n12574_), .ZN(new_n13194_));
  INV_X1     g13002(.I(new_n13194_), .ZN(new_n13195_));
  AOI22_X1   g13003(.A1(new_n13195_), .A2(new_n12724_), .B1(\asqrt[19] ), .B2(new_n13193_), .ZN(new_n13196_));
  NOR3_X1    g13004(.A1(new_n13190_), .A2(new_n13182_), .A3(\asqrt[49] ), .ZN(new_n13197_));
  NOR2_X1    g13005(.A1(new_n13197_), .A2(new_n13196_), .ZN(new_n13198_));
  OAI21_X1   g13006(.A1(new_n13198_), .A2(new_n13192_), .B(\asqrt[50] ), .ZN(new_n13199_));
  NOR2_X1    g13007(.A1(new_n12575_), .A2(new_n12583_), .ZN(new_n13200_));
  NOR3_X1    g13008(.A1(new_n12913_), .A2(new_n12814_), .A3(new_n13200_), .ZN(new_n13201_));
  INV_X1     g13009(.I(new_n13201_), .ZN(new_n13202_));
  NOR3_X1    g13010(.A1(new_n13200_), .A2(new_n12814_), .A3(new_n12582_), .ZN(new_n13203_));
  AOI22_X1   g13011(.A1(new_n13202_), .A2(new_n12582_), .B1(\asqrt[19] ), .B2(new_n13203_), .ZN(new_n13204_));
  INV_X1     g13012(.I(new_n13204_), .ZN(new_n13205_));
  NAND2_X1   g13013(.A1(new_n13191_), .A2(new_n1612_), .ZN(new_n13206_));
  OAI21_X1   g13014(.A1(new_n13198_), .A2(new_n13206_), .B(new_n13205_), .ZN(new_n13207_));
  AOI21_X1   g13015(.A1(new_n13207_), .A2(new_n13199_), .B(new_n1376_), .ZN(new_n13208_));
  INV_X1     g13016(.I(new_n12589_), .ZN(new_n13209_));
  NOR3_X1    g13017(.A1(new_n12585_), .A2(new_n12823_), .A3(new_n13209_), .ZN(new_n13210_));
  NOR3_X1    g13018(.A1(new_n12913_), .A2(new_n12585_), .A3(new_n12823_), .ZN(new_n13211_));
  INV_X1     g13019(.I(new_n13211_), .ZN(new_n13212_));
  AOI22_X1   g13020(.A1(new_n13212_), .A2(new_n13209_), .B1(\asqrt[19] ), .B2(new_n13210_), .ZN(new_n13213_));
  OAI21_X1   g13021(.A1(new_n13196_), .A2(new_n13197_), .B(new_n13191_), .ZN(new_n13214_));
  AOI21_X1   g13022(.A1(new_n13214_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n13215_));
  AOI21_X1   g13023(.A1(new_n13215_), .A2(new_n13207_), .B(new_n13213_), .ZN(new_n13216_));
  OAI21_X1   g13024(.A1(new_n13216_), .A2(new_n13208_), .B(\asqrt[52] ), .ZN(new_n13217_));
  INV_X1     g13025(.I(new_n13217_), .ZN(new_n13218_));
  INV_X1     g13026(.I(new_n13216_), .ZN(new_n13219_));
  NOR3_X1    g13027(.A1(new_n12913_), .A2(new_n12594_), .A3(new_n12600_), .ZN(new_n13220_));
  INV_X1     g13028(.I(new_n13220_), .ZN(new_n13221_));
  NOR3_X1    g13029(.A1(new_n12594_), .A2(new_n12723_), .A3(new_n12600_), .ZN(new_n13222_));
  AOI22_X1   g13030(.A1(new_n13221_), .A2(new_n12723_), .B1(\asqrt[19] ), .B2(new_n13222_), .ZN(new_n13223_));
  NOR2_X1    g13031(.A1(new_n13208_), .A2(\asqrt[52] ), .ZN(new_n13224_));
  AOI21_X1   g13032(.A1(new_n13219_), .A2(new_n13224_), .B(new_n13223_), .ZN(new_n13225_));
  OAI21_X1   g13033(.A1(new_n13225_), .A2(new_n13218_), .B(\asqrt[53] ), .ZN(new_n13226_));
  NOR2_X1    g13034(.A1(new_n12601_), .A2(new_n12611_), .ZN(new_n13227_));
  NOR3_X1    g13035(.A1(new_n13227_), .A2(new_n12822_), .A3(new_n12610_), .ZN(new_n13228_));
  NOR3_X1    g13036(.A1(new_n12913_), .A2(new_n12822_), .A3(new_n13227_), .ZN(new_n13229_));
  INV_X1     g13037(.I(new_n13229_), .ZN(new_n13230_));
  AOI22_X1   g13038(.A1(new_n13230_), .A2(new_n12610_), .B1(\asqrt[19] ), .B2(new_n13228_), .ZN(new_n13231_));
  INV_X1     g13039(.I(new_n13231_), .ZN(new_n13232_));
  NAND2_X1   g13040(.A1(new_n13217_), .A2(new_n1103_), .ZN(new_n13233_));
  OAI21_X1   g13041(.A1(new_n13233_), .A2(new_n13225_), .B(new_n13232_), .ZN(new_n13234_));
  AOI21_X1   g13042(.A1(new_n13234_), .A2(new_n13226_), .B(new_n904_), .ZN(new_n13235_));
  INV_X1     g13043(.I(new_n13235_), .ZN(new_n13236_));
  INV_X1     g13044(.I(new_n13234_), .ZN(new_n13237_));
  INV_X1     g13045(.I(new_n12617_), .ZN(new_n13238_));
  NOR3_X1    g13046(.A1(new_n12913_), .A2(new_n12613_), .A3(new_n12831_), .ZN(new_n13239_));
  INV_X1     g13047(.I(new_n13239_), .ZN(new_n13240_));
  NOR3_X1    g13048(.A1(new_n12613_), .A2(new_n12831_), .A3(new_n13238_), .ZN(new_n13241_));
  AOI22_X1   g13049(.A1(new_n13240_), .A2(new_n13238_), .B1(\asqrt[19] ), .B2(new_n13241_), .ZN(new_n13242_));
  INV_X1     g13050(.I(new_n13242_), .ZN(new_n13243_));
  NAND2_X1   g13051(.A1(new_n13226_), .A2(new_n904_), .ZN(new_n13244_));
  OAI21_X1   g13052(.A1(new_n13244_), .A2(new_n13237_), .B(new_n13243_), .ZN(new_n13245_));
  AOI21_X1   g13053(.A1(new_n13245_), .A2(new_n13236_), .B(new_n823_), .ZN(new_n13246_));
  NOR3_X1    g13054(.A1(new_n12622_), .A2(new_n12722_), .A3(new_n12629_), .ZN(new_n13247_));
  NOR3_X1    g13055(.A1(new_n12913_), .A2(new_n12622_), .A3(new_n12629_), .ZN(new_n13248_));
  INV_X1     g13056(.I(new_n13248_), .ZN(new_n13249_));
  AOI22_X1   g13057(.A1(new_n13249_), .A2(new_n12722_), .B1(\asqrt[19] ), .B2(new_n13247_), .ZN(new_n13250_));
  NOR2_X1    g13058(.A1(new_n13235_), .A2(\asqrt[55] ), .ZN(new_n13251_));
  AOI21_X1   g13059(.A1(new_n13251_), .A2(new_n13245_), .B(new_n13250_), .ZN(new_n13252_));
  OAI21_X1   g13060(.A1(new_n13252_), .A2(new_n13246_), .B(\asqrt[56] ), .ZN(new_n13253_));
  NOR2_X1    g13061(.A1(new_n12630_), .A2(new_n12641_), .ZN(new_n13254_));
  NOR3_X1    g13062(.A1(new_n12913_), .A2(new_n12830_), .A3(new_n13254_), .ZN(new_n13255_));
  INV_X1     g13063(.I(new_n13255_), .ZN(new_n13256_));
  NOR3_X1    g13064(.A1(new_n13254_), .A2(new_n12830_), .A3(new_n12640_), .ZN(new_n13257_));
  AOI22_X1   g13065(.A1(new_n13256_), .A2(new_n12640_), .B1(\asqrt[19] ), .B2(new_n13257_), .ZN(new_n13258_));
  INV_X1     g13066(.I(new_n13258_), .ZN(new_n13259_));
  NOR3_X1    g13067(.A1(new_n13216_), .A2(new_n13208_), .A3(\asqrt[52] ), .ZN(new_n13260_));
  OAI21_X1   g13068(.A1(new_n13223_), .A2(new_n13260_), .B(new_n13217_), .ZN(new_n13261_));
  AOI21_X1   g13069(.A1(new_n13261_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n13262_));
  AOI21_X1   g13070(.A1(new_n13262_), .A2(new_n13234_), .B(new_n13242_), .ZN(new_n13263_));
  OAI21_X1   g13071(.A1(new_n13263_), .A2(new_n13235_), .B(\asqrt[55] ), .ZN(new_n13264_));
  NAND2_X1   g13072(.A1(new_n13264_), .A2(new_n703_), .ZN(new_n13265_));
  OAI21_X1   g13073(.A1(new_n13265_), .A2(new_n13252_), .B(new_n13259_), .ZN(new_n13266_));
  AOI21_X1   g13074(.A1(new_n13266_), .A2(new_n13253_), .B(new_n531_), .ZN(new_n13267_));
  INV_X1     g13075(.I(new_n13267_), .ZN(new_n13268_));
  INV_X1     g13076(.I(new_n13266_), .ZN(new_n13269_));
  INV_X1     g13077(.I(new_n12647_), .ZN(new_n13270_));
  NOR3_X1    g13078(.A1(new_n12643_), .A2(new_n12839_), .A3(new_n13270_), .ZN(new_n13271_));
  NOR3_X1    g13079(.A1(new_n12913_), .A2(new_n12643_), .A3(new_n12839_), .ZN(new_n13272_));
  INV_X1     g13080(.I(new_n13272_), .ZN(new_n13273_));
  AOI22_X1   g13081(.A1(new_n13273_), .A2(new_n13270_), .B1(\asqrt[19] ), .B2(new_n13271_), .ZN(new_n13274_));
  INV_X1     g13082(.I(new_n13274_), .ZN(new_n13275_));
  NAND2_X1   g13083(.A1(new_n13253_), .A2(new_n531_), .ZN(new_n13276_));
  OAI21_X1   g13084(.A1(new_n13276_), .A2(new_n13269_), .B(new_n13275_), .ZN(new_n13277_));
  AOI21_X1   g13085(.A1(new_n13277_), .A2(new_n13268_), .B(new_n436_), .ZN(new_n13278_));
  NOR3_X1    g13086(.A1(new_n12913_), .A2(new_n12652_), .A3(new_n12659_), .ZN(new_n13279_));
  INV_X1     g13087(.I(new_n13279_), .ZN(new_n13280_));
  NOR3_X1    g13088(.A1(new_n12652_), .A2(new_n12721_), .A3(new_n12659_), .ZN(new_n13281_));
  AOI22_X1   g13089(.A1(new_n13280_), .A2(new_n12721_), .B1(\asqrt[19] ), .B2(new_n13281_), .ZN(new_n13282_));
  NOR2_X1    g13090(.A1(new_n13267_), .A2(\asqrt[58] ), .ZN(new_n13283_));
  AOI21_X1   g13091(.A1(new_n13283_), .A2(new_n13277_), .B(new_n13282_), .ZN(new_n13284_));
  OAI21_X1   g13092(.A1(new_n13284_), .A2(new_n13278_), .B(\asqrt[59] ), .ZN(new_n13285_));
  NOR2_X1    g13093(.A1(new_n12660_), .A2(new_n12672_), .ZN(new_n13286_));
  NOR3_X1    g13094(.A1(new_n13286_), .A2(new_n12838_), .A3(new_n12671_), .ZN(new_n13287_));
  NOR3_X1    g13095(.A1(new_n12913_), .A2(new_n12838_), .A3(new_n13286_), .ZN(new_n13288_));
  INV_X1     g13096(.I(new_n13288_), .ZN(new_n13289_));
  AOI22_X1   g13097(.A1(new_n13289_), .A2(new_n12671_), .B1(\asqrt[19] ), .B2(new_n13287_), .ZN(new_n13290_));
  INV_X1     g13098(.I(new_n13290_), .ZN(new_n13291_));
  NOR3_X1    g13099(.A1(new_n13263_), .A2(\asqrt[55] ), .A3(new_n13235_), .ZN(new_n13292_));
  OAI21_X1   g13100(.A1(new_n13250_), .A2(new_n13292_), .B(new_n13264_), .ZN(new_n13293_));
  AOI21_X1   g13101(.A1(new_n13293_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n13294_));
  AOI21_X1   g13102(.A1(new_n13294_), .A2(new_n13266_), .B(new_n13274_), .ZN(new_n13295_));
  OAI21_X1   g13103(.A1(new_n13295_), .A2(new_n13267_), .B(\asqrt[58] ), .ZN(new_n13296_));
  NAND2_X1   g13104(.A1(new_n13296_), .A2(new_n327_), .ZN(new_n13297_));
  OAI21_X1   g13105(.A1(new_n13297_), .A2(new_n13284_), .B(new_n13291_), .ZN(new_n13298_));
  AOI21_X1   g13106(.A1(new_n13298_), .A2(new_n13285_), .B(new_n306_), .ZN(new_n13299_));
  INV_X1     g13107(.I(new_n13299_), .ZN(new_n13300_));
  INV_X1     g13108(.I(new_n13298_), .ZN(new_n13301_));
  INV_X1     g13109(.I(new_n12678_), .ZN(new_n13302_));
  NOR3_X1    g13110(.A1(new_n12913_), .A2(new_n12674_), .A3(new_n12846_), .ZN(new_n13303_));
  INV_X1     g13111(.I(new_n13303_), .ZN(new_n13304_));
  NOR3_X1    g13112(.A1(new_n12674_), .A2(new_n12846_), .A3(new_n13302_), .ZN(new_n13305_));
  AOI22_X1   g13113(.A1(new_n13304_), .A2(new_n13302_), .B1(\asqrt[19] ), .B2(new_n13305_), .ZN(new_n13306_));
  INV_X1     g13114(.I(new_n13306_), .ZN(new_n13307_));
  NAND2_X1   g13115(.A1(new_n13285_), .A2(new_n306_), .ZN(new_n13308_));
  OAI21_X1   g13116(.A1(new_n13301_), .A2(new_n13308_), .B(new_n13307_), .ZN(new_n13309_));
  AOI21_X1   g13117(.A1(new_n13309_), .A2(new_n13300_), .B(new_n218_), .ZN(new_n13310_));
  NOR3_X1    g13118(.A1(new_n12683_), .A2(new_n12720_), .A3(new_n12689_), .ZN(new_n13311_));
  NOR3_X1    g13119(.A1(new_n12913_), .A2(new_n12683_), .A3(new_n12689_), .ZN(new_n13312_));
  INV_X1     g13120(.I(new_n13312_), .ZN(new_n13313_));
  AOI22_X1   g13121(.A1(new_n13313_), .A2(new_n12720_), .B1(\asqrt[19] ), .B2(new_n13311_), .ZN(new_n13314_));
  NOR2_X1    g13122(.A1(new_n13299_), .A2(\asqrt[61] ), .ZN(new_n13315_));
  AOI21_X1   g13123(.A1(new_n13315_), .A2(new_n13309_), .B(new_n13314_), .ZN(new_n13316_));
  OAI21_X1   g13124(.A1(new_n13316_), .A2(new_n13310_), .B(\asqrt[62] ), .ZN(new_n13317_));
  NOR2_X1    g13125(.A1(new_n12690_), .A2(new_n12697_), .ZN(new_n13318_));
  NOR3_X1    g13126(.A1(new_n12913_), .A2(new_n12868_), .A3(new_n13318_), .ZN(new_n13319_));
  INV_X1     g13127(.I(new_n13319_), .ZN(new_n13320_));
  NOR3_X1    g13128(.A1(new_n13318_), .A2(new_n12868_), .A3(new_n12696_), .ZN(new_n13321_));
  AOI22_X1   g13129(.A1(new_n13320_), .A2(new_n12696_), .B1(\asqrt[19] ), .B2(new_n13321_), .ZN(new_n13322_));
  INV_X1     g13130(.I(new_n13322_), .ZN(new_n13323_));
  NOR3_X1    g13131(.A1(new_n13295_), .A2(\asqrt[58] ), .A3(new_n13267_), .ZN(new_n13324_));
  OAI21_X1   g13132(.A1(new_n13282_), .A2(new_n13324_), .B(new_n13296_), .ZN(new_n13325_));
  AOI21_X1   g13133(.A1(new_n13325_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n13326_));
  AOI21_X1   g13134(.A1(new_n13326_), .A2(new_n13298_), .B(new_n13306_), .ZN(new_n13327_));
  OAI21_X1   g13135(.A1(new_n13327_), .A2(new_n13299_), .B(\asqrt[61] ), .ZN(new_n13328_));
  NAND2_X1   g13136(.A1(new_n13328_), .A2(new_n207_), .ZN(new_n13329_));
  OAI21_X1   g13137(.A1(new_n13329_), .A2(new_n13316_), .B(new_n13323_), .ZN(new_n13330_));
  INV_X1     g13138(.I(new_n12870_), .ZN(new_n13331_));
  NAND4_X1   g13139(.A1(\asqrt[19] ), .A2(new_n12869_), .A3(new_n12703_), .A4(new_n13331_), .ZN(new_n13332_));
  NAND2_X1   g13140(.A1(new_n13331_), .A2(new_n12869_), .ZN(new_n13333_));
  OAI21_X1   g13141(.A1(new_n12913_), .A2(new_n13333_), .B(new_n12850_), .ZN(new_n13334_));
  NAND2_X1   g13142(.A1(new_n13334_), .A2(new_n13332_), .ZN(new_n13335_));
  INV_X1     g13143(.I(new_n12889_), .ZN(new_n13336_));
  AOI21_X1   g13144(.A1(new_n12852_), .A2(new_n12869_), .B(new_n12714_), .ZN(new_n13337_));
  AOI21_X1   g13145(.A1(\asqrt[19] ), .A2(new_n13337_), .B(new_n13336_), .ZN(new_n13338_));
  NAND2_X1   g13146(.A1(new_n13335_), .A2(new_n13338_), .ZN(new_n13339_));
  AOI21_X1   g13147(.A1(new_n13330_), .A2(new_n13317_), .B(new_n13339_), .ZN(new_n13340_));
  NOR2_X1    g13148(.A1(new_n13340_), .A2(\asqrt[63] ), .ZN(new_n13341_));
  INV_X1     g13149(.I(new_n13330_), .ZN(new_n13342_));
  INV_X1     g13150(.I(new_n13335_), .ZN(new_n13343_));
  NAND2_X1   g13151(.A1(new_n13317_), .A2(new_n13343_), .ZN(new_n13344_));
  AOI21_X1   g13152(.A1(\asqrt[19] ), .A2(new_n12715_), .B(new_n12871_), .ZN(new_n13345_));
  OR3_X2     g13153(.A1(new_n13345_), .A2(new_n193_), .A3(new_n13337_), .Z(new_n13346_));
  OAI21_X1   g13154(.A1(new_n12311_), .A2(new_n12858_), .B(new_n12710_), .ZN(new_n13347_));
  NOR4_X1    g13155(.A1(new_n13336_), .A2(new_n12713_), .A3(new_n12856_), .A4(new_n13347_), .ZN(new_n13348_));
  NAND2_X1   g13156(.A1(new_n13348_), .A2(new_n12719_), .ZN(new_n13349_));
  NAND2_X1   g13157(.A1(new_n13346_), .A2(new_n13349_), .ZN(new_n13350_));
  INV_X1     g13158(.I(new_n13350_), .ZN(new_n13351_));
  OAI21_X1   g13159(.A1(new_n13342_), .A2(new_n13344_), .B(new_n13351_), .ZN(new_n13352_));
  NOR2_X1    g13160(.A1(new_n13341_), .A2(new_n13352_), .ZN(new_n13353_));
  INV_X1     g13161(.I(\a[36] ), .ZN(new_n13354_));
  NOR2_X1    g13162(.A1(\a[34] ), .A2(\a[35] ), .ZN(new_n13355_));
  INV_X1     g13163(.I(new_n13355_), .ZN(new_n13356_));
  NOR2_X1    g13164(.A1(new_n13356_), .A2(\a[36] ), .ZN(new_n13357_));
  INV_X1     g13165(.I(new_n13357_), .ZN(new_n13358_));
  OAI21_X1   g13166(.A1(new_n13353_), .A2(new_n13354_), .B(new_n13358_), .ZN(new_n13359_));
  NOR3_X1    g13167(.A1(new_n12856_), .A2(new_n12859_), .A3(new_n13357_), .ZN(new_n13360_));
  NAND3_X1   g13168(.A1(new_n12719_), .A2(new_n12889_), .A3(new_n13360_), .ZN(new_n13361_));
  INV_X1     g13169(.I(new_n13361_), .ZN(new_n13362_));
  OAI21_X1   g13170(.A1(new_n13353_), .A2(new_n13354_), .B(new_n13362_), .ZN(new_n13363_));
  NOR3_X1    g13171(.A1(new_n13327_), .A2(\asqrt[61] ), .A3(new_n13299_), .ZN(new_n13364_));
  OAI21_X1   g13172(.A1(new_n13314_), .A2(new_n13364_), .B(new_n13328_), .ZN(new_n13365_));
  INV_X1     g13173(.I(new_n13314_), .ZN(new_n13366_));
  INV_X1     g13174(.I(new_n13282_), .ZN(new_n13367_));
  INV_X1     g13175(.I(new_n13250_), .ZN(new_n13368_));
  INV_X1     g13176(.I(new_n13223_), .ZN(new_n13369_));
  INV_X1     g13177(.I(new_n13196_), .ZN(new_n13370_));
  INV_X1     g13178(.I(new_n13170_), .ZN(new_n13371_));
  INV_X1     g13179(.I(new_n13144_), .ZN(new_n13372_));
  INV_X1     g13180(.I(new_n13115_), .ZN(new_n13373_));
  NOR3_X1    g13181(.A1(new_n13114_), .A2(new_n13099_), .A3(\asqrt[41] ), .ZN(new_n13374_));
  NOR2_X1    g13182(.A1(new_n13374_), .A2(new_n13120_), .ZN(new_n13375_));
  OAI21_X1   g13183(.A1(new_n13375_), .A2(new_n13373_), .B(\asqrt[42] ), .ZN(new_n13376_));
  NAND2_X1   g13184(.A1(new_n13376_), .A2(new_n3218_), .ZN(new_n13377_));
  OAI21_X1   g13185(.A1(new_n13377_), .A2(new_n13138_), .B(new_n13372_), .ZN(new_n13378_));
  NAND3_X1   g13186(.A1(new_n13378_), .A2(new_n2954_), .A3(new_n13139_), .ZN(new_n13379_));
  AOI22_X1   g13187(.A1(new_n13379_), .A2(new_n13153_), .B1(\asqrt[44] ), .B2(new_n13162_), .ZN(new_n13380_));
  OAI21_X1   g13188(.A1(new_n13380_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n13381_));
  OAI21_X1   g13189(.A1(new_n13381_), .A2(new_n13164_), .B(new_n13371_), .ZN(new_n13382_));
  NAND3_X1   g13190(.A1(new_n13382_), .A2(new_n2229_), .A3(new_n13165_), .ZN(new_n13383_));
  AOI22_X1   g13191(.A1(new_n13383_), .A2(new_n13179_), .B1(\asqrt[47] ), .B2(new_n13188_), .ZN(new_n13384_));
  OAI21_X1   g13192(.A1(new_n13384_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n13385_));
  OAI21_X1   g13193(.A1(new_n13385_), .A2(new_n13190_), .B(new_n13370_), .ZN(new_n13386_));
  NAND3_X1   g13194(.A1(new_n13386_), .A2(new_n1612_), .A3(new_n13191_), .ZN(new_n13387_));
  AOI22_X1   g13195(.A1(new_n13387_), .A2(new_n13205_), .B1(\asqrt[50] ), .B2(new_n13214_), .ZN(new_n13388_));
  OAI21_X1   g13196(.A1(new_n13388_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n13389_));
  OAI21_X1   g13197(.A1(new_n13389_), .A2(new_n13216_), .B(new_n13369_), .ZN(new_n13390_));
  NAND3_X1   g13198(.A1(new_n13390_), .A2(new_n1103_), .A3(new_n13217_), .ZN(new_n13391_));
  AOI22_X1   g13199(.A1(new_n13391_), .A2(new_n13232_), .B1(\asqrt[53] ), .B2(new_n13261_), .ZN(new_n13392_));
  OAI21_X1   g13200(.A1(new_n13392_), .A2(new_n904_), .B(new_n823_), .ZN(new_n13393_));
  OAI21_X1   g13201(.A1(new_n13393_), .A2(new_n13263_), .B(new_n13368_), .ZN(new_n13394_));
  NAND3_X1   g13202(.A1(new_n13394_), .A2(new_n703_), .A3(new_n13264_), .ZN(new_n13395_));
  AOI22_X1   g13203(.A1(new_n13395_), .A2(new_n13259_), .B1(\asqrt[56] ), .B2(new_n13293_), .ZN(new_n13396_));
  OAI21_X1   g13204(.A1(new_n13396_), .A2(new_n531_), .B(new_n436_), .ZN(new_n13397_));
  OAI21_X1   g13205(.A1(new_n13397_), .A2(new_n13295_), .B(new_n13367_), .ZN(new_n13398_));
  NAND3_X1   g13206(.A1(new_n13398_), .A2(new_n327_), .A3(new_n13296_), .ZN(new_n13399_));
  AOI22_X1   g13207(.A1(new_n13399_), .A2(new_n13291_), .B1(new_n13325_), .B2(\asqrt[59] ), .ZN(new_n13400_));
  OAI21_X1   g13208(.A1(new_n13400_), .A2(new_n306_), .B(new_n218_), .ZN(new_n13401_));
  OAI21_X1   g13209(.A1(new_n13401_), .A2(new_n13327_), .B(new_n13366_), .ZN(new_n13402_));
  NAND3_X1   g13210(.A1(new_n13402_), .A2(new_n207_), .A3(new_n13328_), .ZN(new_n13403_));
  AOI22_X1   g13211(.A1(new_n13403_), .A2(new_n13323_), .B1(new_n13365_), .B2(\asqrt[62] ), .ZN(new_n13404_));
  OAI21_X1   g13212(.A1(new_n13404_), .A2(new_n13339_), .B(new_n193_), .ZN(new_n13405_));
  AOI21_X1   g13213(.A1(new_n13365_), .A2(\asqrt[62] ), .B(new_n13335_), .ZN(new_n13406_));
  AOI21_X1   g13214(.A1(new_n13406_), .A2(new_n13330_), .B(new_n13350_), .ZN(new_n13407_));
  AOI21_X1   g13215(.A1(new_n13405_), .A2(new_n13407_), .B(new_n12865_), .ZN(new_n13408_));
  OAI21_X1   g13216(.A1(new_n13341_), .A2(new_n13352_), .B(new_n13354_), .ZN(new_n13409_));
  AOI21_X1   g13217(.A1(\a[37] ), .A2(new_n13409_), .B(new_n13408_), .ZN(new_n13410_));
  AOI22_X1   g13218(.A1(new_n13410_), .A2(new_n13363_), .B1(\asqrt[19] ), .B2(new_n13359_), .ZN(new_n13411_));
  NOR2_X1    g13219(.A1(new_n13411_), .A2(new_n12364_), .ZN(new_n13412_));
  NAND2_X1   g13220(.A1(new_n13410_), .A2(new_n13363_), .ZN(new_n13413_));
  OAI21_X1   g13221(.A1(new_n13341_), .A2(new_n13352_), .B(new_n12864_), .ZN(new_n13414_));
  NAND2_X1   g13222(.A1(new_n13406_), .A2(new_n13330_), .ZN(new_n13415_));
  OAI21_X1   g13223(.A1(new_n13348_), .A2(new_n12862_), .B(new_n12719_), .ZN(new_n13416_));
  NAND4_X1   g13224(.A1(new_n13405_), .A2(new_n13415_), .A3(new_n13346_), .A4(new_n13416_), .ZN(new_n13417_));
  AOI21_X1   g13225(.A1(new_n13417_), .A2(new_n13414_), .B(new_n12877_), .ZN(new_n13418_));
  INV_X1     g13226(.I(new_n13415_), .ZN(new_n13419_));
  NAND2_X1   g13227(.A1(new_n13346_), .A2(new_n13416_), .ZN(new_n13420_));
  NOR3_X1    g13228(.A1(new_n13419_), .A2(new_n13341_), .A3(new_n13420_), .ZN(new_n13421_));
  NOR3_X1    g13229(.A1(new_n13421_), .A2(new_n13408_), .A3(\a[38] ), .ZN(new_n13422_));
  NOR2_X1    g13230(.A1(new_n13418_), .A2(new_n13422_), .ZN(new_n13423_));
  AOI21_X1   g13231(.A1(new_n13359_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n13424_));
  AOI21_X1   g13232(.A1(new_n13413_), .A2(new_n13424_), .B(new_n13423_), .ZN(new_n13425_));
  OAI21_X1   g13233(.A1(new_n13425_), .A2(new_n13412_), .B(\asqrt[21] ), .ZN(new_n13426_));
  OAI21_X1   g13234(.A1(\asqrt[63] ), .A2(new_n13340_), .B(new_n13407_), .ZN(\asqrt[18] ));
  NOR3_X1    g13235(.A1(new_n12957_), .A2(new_n12876_), .A3(new_n12882_), .ZN(new_n13428_));
  NAND3_X1   g13236(.A1(\asqrt[18] ), .A2(new_n12895_), .A3(new_n12942_), .ZN(new_n13429_));
  AOI22_X1   g13237(.A1(new_n13429_), .A2(new_n12957_), .B1(\asqrt[18] ), .B2(new_n13428_), .ZN(new_n13430_));
  INV_X1     g13238(.I(new_n13430_), .ZN(new_n13431_));
  OAI21_X1   g13239(.A1(new_n13411_), .A2(new_n12364_), .B(new_n11736_), .ZN(new_n13432_));
  OAI21_X1   g13240(.A1(new_n13432_), .A2(new_n13425_), .B(new_n13431_), .ZN(new_n13433_));
  AOI21_X1   g13241(.A1(new_n13433_), .A2(new_n13426_), .B(new_n11326_), .ZN(new_n13434_));
  NOR2_X1    g13242(.A1(new_n12894_), .A2(new_n12892_), .ZN(new_n13435_));
  NOR2_X1    g13243(.A1(new_n12886_), .A2(new_n12896_), .ZN(new_n13436_));
  INV_X1     g13244(.I(new_n13436_), .ZN(new_n13437_));
  NAND4_X1   g13245(.A1(\asqrt[18] ), .A2(new_n12887_), .A3(new_n13435_), .A4(new_n13437_), .ZN(new_n13438_));
  NOR3_X1    g13246(.A1(new_n13353_), .A2(new_n12946_), .A3(new_n13436_), .ZN(new_n13439_));
  OAI21_X1   g13247(.A1(new_n13439_), .A2(new_n13435_), .B(new_n13438_), .ZN(new_n13440_));
  INV_X1     g13248(.I(new_n13440_), .ZN(new_n13441_));
  AOI21_X1   g13249(.A1(new_n13405_), .A2(new_n13407_), .B(new_n13354_), .ZN(new_n13442_));
  OAI21_X1   g13250(.A1(new_n13442_), .A2(new_n13357_), .B(\asqrt[19] ), .ZN(new_n13443_));
  INV_X1     g13251(.I(new_n13443_), .ZN(new_n13444_));
  NOR2_X1    g13252(.A1(new_n13442_), .A2(new_n13361_), .ZN(new_n13445_));
  INV_X1     g13253(.I(\a[37] ), .ZN(new_n13446_));
  AOI21_X1   g13254(.A1(\asqrt[18] ), .A2(new_n13354_), .B(new_n13446_), .ZN(new_n13447_));
  NOR3_X1    g13255(.A1(new_n13445_), .A2(new_n13447_), .A3(new_n13408_), .ZN(new_n13448_));
  OAI21_X1   g13256(.A1(new_n13448_), .A2(new_n13444_), .B(\asqrt[20] ), .ZN(new_n13449_));
  AOI21_X1   g13257(.A1(\asqrt[18] ), .A2(\a[36] ), .B(new_n13357_), .ZN(new_n13450_));
  OAI21_X1   g13258(.A1(new_n13450_), .A2(new_n12913_), .B(new_n12364_), .ZN(new_n13451_));
  OAI22_X1   g13259(.A1(new_n13448_), .A2(new_n13451_), .B1(new_n13418_), .B2(new_n13422_), .ZN(new_n13452_));
  AOI21_X1   g13260(.A1(new_n13452_), .A2(new_n13449_), .B(new_n11736_), .ZN(new_n13453_));
  AOI21_X1   g13261(.A1(new_n13405_), .A2(new_n13407_), .B(\a[36] ), .ZN(new_n13454_));
  OAI21_X1   g13262(.A1(new_n13446_), .A2(new_n13454_), .B(new_n13414_), .ZN(new_n13455_));
  OAI21_X1   g13263(.A1(new_n13455_), .A2(new_n13445_), .B(new_n13443_), .ZN(new_n13456_));
  AOI21_X1   g13264(.A1(new_n13456_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n13457_));
  AOI21_X1   g13265(.A1(new_n13457_), .A2(new_n13452_), .B(new_n13430_), .ZN(new_n13458_));
  NOR3_X1    g13266(.A1(new_n13458_), .A2(new_n13453_), .A3(\asqrt[22] ), .ZN(new_n13459_));
  NOR2_X1    g13267(.A1(new_n13459_), .A2(new_n13441_), .ZN(new_n13460_));
  OAI21_X1   g13268(.A1(new_n13460_), .A2(new_n13434_), .B(\asqrt[23] ), .ZN(new_n13461_));
  NOR2_X1    g13269(.A1(new_n12959_), .A2(new_n12951_), .ZN(new_n13462_));
  NOR3_X1    g13270(.A1(new_n13353_), .A2(new_n12898_), .A3(new_n13462_), .ZN(new_n13463_));
  INV_X1     g13271(.I(new_n13463_), .ZN(new_n13464_));
  NOR3_X1    g13272(.A1(new_n13462_), .A2(new_n12898_), .A3(new_n12956_), .ZN(new_n13465_));
  AOI22_X1   g13273(.A1(new_n13464_), .A2(new_n12956_), .B1(\asqrt[18] ), .B2(new_n13465_), .ZN(new_n13466_));
  INV_X1     g13274(.I(new_n13466_), .ZN(new_n13467_));
  OAI21_X1   g13275(.A1(new_n13458_), .A2(new_n13453_), .B(\asqrt[22] ), .ZN(new_n13468_));
  NAND2_X1   g13276(.A1(new_n13468_), .A2(new_n10812_), .ZN(new_n13469_));
  OAI21_X1   g13277(.A1(new_n13460_), .A2(new_n13469_), .B(new_n13467_), .ZN(new_n13470_));
  AOI21_X1   g13278(.A1(new_n13470_), .A2(new_n13461_), .B(new_n10221_), .ZN(new_n13471_));
  NOR3_X1    g13279(.A1(new_n12908_), .A2(new_n12917_), .A3(new_n12915_), .ZN(new_n13472_));
  NOR3_X1    g13280(.A1(new_n13353_), .A2(new_n12908_), .A3(new_n12917_), .ZN(new_n13473_));
  INV_X1     g13281(.I(new_n13473_), .ZN(new_n13474_));
  AOI22_X1   g13282(.A1(new_n13474_), .A2(new_n12915_), .B1(\asqrt[18] ), .B2(new_n13472_), .ZN(new_n13475_));
  OAI21_X1   g13283(.A1(new_n13441_), .A2(new_n13459_), .B(new_n13468_), .ZN(new_n13476_));
  AOI21_X1   g13284(.A1(new_n13476_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n13477_));
  AOI21_X1   g13285(.A1(new_n13477_), .A2(new_n13470_), .B(new_n13475_), .ZN(new_n13478_));
  OAI21_X1   g13286(.A1(new_n13478_), .A2(new_n13471_), .B(\asqrt[25] ), .ZN(new_n13479_));
  INV_X1     g13287(.I(new_n13479_), .ZN(new_n13480_));
  NAND2_X1   g13288(.A1(new_n12962_), .A2(new_n12954_), .ZN(new_n13481_));
  NAND3_X1   g13289(.A1(\asqrt[18] ), .A2(new_n12919_), .A3(new_n13481_), .ZN(new_n13482_));
  AND3_X2    g13290(.A1(new_n12919_), .A2(new_n12924_), .A3(new_n13481_), .Z(new_n13483_));
  AOI22_X1   g13291(.A1(new_n13482_), .A2(new_n12925_), .B1(\asqrt[18] ), .B2(new_n13483_), .ZN(new_n13484_));
  NOR3_X1    g13292(.A1(new_n13478_), .A2(new_n13471_), .A3(\asqrt[25] ), .ZN(new_n13485_));
  NOR2_X1    g13293(.A1(new_n13485_), .A2(new_n13484_), .ZN(new_n13486_));
  OAI21_X1   g13294(.A1(new_n13486_), .A2(new_n13480_), .B(\asqrt[26] ), .ZN(new_n13487_));
  INV_X1     g13295(.I(new_n12932_), .ZN(new_n13488_));
  NOR3_X1    g13296(.A1(new_n12928_), .A2(new_n12973_), .A3(new_n13488_), .ZN(new_n13489_));
  NOR3_X1    g13297(.A1(new_n13353_), .A2(new_n12928_), .A3(new_n12973_), .ZN(new_n13490_));
  INV_X1     g13298(.I(new_n13490_), .ZN(new_n13491_));
  AOI22_X1   g13299(.A1(new_n13491_), .A2(new_n13488_), .B1(\asqrt[18] ), .B2(new_n13489_), .ZN(new_n13492_));
  INV_X1     g13300(.I(new_n13492_), .ZN(new_n13493_));
  NAND2_X1   g13301(.A1(new_n13479_), .A2(new_n9317_), .ZN(new_n13494_));
  OAI21_X1   g13302(.A1(new_n13486_), .A2(new_n13494_), .B(new_n13493_), .ZN(new_n13495_));
  AOI21_X1   g13303(.A1(new_n13495_), .A2(new_n13487_), .B(new_n8826_), .ZN(new_n13496_));
  INV_X1     g13304(.I(new_n13020_), .ZN(new_n13497_));
  NAND3_X1   g13305(.A1(\asqrt[18] ), .A2(new_n12936_), .A3(new_n13497_), .ZN(new_n13498_));
  AND3_X2    g13306(.A1(new_n13497_), .A2(new_n12936_), .A3(new_n12940_), .Z(new_n13499_));
  AOI22_X1   g13307(.A1(new_n13498_), .A2(new_n12941_), .B1(\asqrt[18] ), .B2(new_n13499_), .ZN(new_n13500_));
  OAI21_X1   g13308(.A1(new_n13484_), .A2(new_n13485_), .B(new_n13479_), .ZN(new_n13501_));
  AOI21_X1   g13309(.A1(new_n13501_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n13502_));
  AOI21_X1   g13310(.A1(new_n13502_), .A2(new_n13495_), .B(new_n13500_), .ZN(new_n13503_));
  OAI21_X1   g13311(.A1(new_n13503_), .A2(new_n13496_), .B(\asqrt[28] ), .ZN(new_n13504_));
  INV_X1     g13312(.I(new_n13504_), .ZN(new_n13505_));
  INV_X1     g13313(.I(new_n12980_), .ZN(new_n13506_));
  NOR3_X1    g13314(.A1(new_n13506_), .A2(new_n12967_), .A3(new_n12979_), .ZN(new_n13507_));
  NOR3_X1    g13315(.A1(new_n13353_), .A2(new_n12967_), .A3(new_n13506_), .ZN(new_n13508_));
  INV_X1     g13316(.I(new_n13508_), .ZN(new_n13509_));
  AOI22_X1   g13317(.A1(new_n13509_), .A2(new_n12979_), .B1(\asqrt[18] ), .B2(new_n13507_), .ZN(new_n13510_));
  NOR3_X1    g13318(.A1(new_n13503_), .A2(new_n13496_), .A3(\asqrt[28] ), .ZN(new_n13511_));
  NOR2_X1    g13319(.A1(new_n13511_), .A2(new_n13510_), .ZN(new_n13512_));
  OAI21_X1   g13320(.A1(new_n13512_), .A2(new_n13505_), .B(\asqrt[29] ), .ZN(new_n13513_));
  INV_X1     g13321(.I(new_n12985_), .ZN(new_n13514_));
  NOR3_X1    g13322(.A1(new_n13353_), .A2(new_n12978_), .A3(new_n13023_), .ZN(new_n13515_));
  INV_X1     g13323(.I(new_n13515_), .ZN(new_n13516_));
  NOR3_X1    g13324(.A1(new_n12978_), .A2(new_n13514_), .A3(new_n13023_), .ZN(new_n13517_));
  AOI22_X1   g13325(.A1(new_n13516_), .A2(new_n13514_), .B1(\asqrt[18] ), .B2(new_n13517_), .ZN(new_n13518_));
  INV_X1     g13326(.I(new_n13518_), .ZN(new_n13519_));
  NAND2_X1   g13327(.A1(new_n13504_), .A2(new_n8036_), .ZN(new_n13520_));
  OAI21_X1   g13328(.A1(new_n13512_), .A2(new_n13520_), .B(new_n13519_), .ZN(new_n13521_));
  AOI21_X1   g13329(.A1(new_n13521_), .A2(new_n13513_), .B(new_n7539_), .ZN(new_n13522_));
  OAI21_X1   g13330(.A1(new_n12993_), .A2(new_n12987_), .B(new_n12991_), .ZN(new_n13523_));
  AOI21_X1   g13331(.A1(\asqrt[29] ), .A2(new_n13024_), .B(new_n13523_), .ZN(new_n13524_));
  OAI21_X1   g13332(.A1(new_n12987_), .A2(new_n12993_), .B(new_n12988_), .ZN(new_n13525_));
  NOR2_X1    g13333(.A1(new_n13353_), .A2(new_n13525_), .ZN(new_n13526_));
  INV_X1     g13334(.I(new_n13526_), .ZN(new_n13527_));
  AOI22_X1   g13335(.A1(new_n13527_), .A2(new_n12992_), .B1(\asqrt[18] ), .B2(new_n13524_), .ZN(new_n13528_));
  OAI21_X1   g13336(.A1(new_n13510_), .A2(new_n13511_), .B(new_n13504_), .ZN(new_n13529_));
  AOI21_X1   g13337(.A1(new_n13529_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n13530_));
  AOI21_X1   g13338(.A1(new_n13530_), .A2(new_n13521_), .B(new_n13528_), .ZN(new_n13531_));
  OAI21_X1   g13339(.A1(new_n13531_), .A2(new_n13522_), .B(\asqrt[31] ), .ZN(new_n13532_));
  INV_X1     g13340(.I(new_n13532_), .ZN(new_n13533_));
  NOR2_X1    g13341(.A1(new_n13004_), .A2(new_n12997_), .ZN(new_n13534_));
  NOR3_X1    g13342(.A1(new_n13353_), .A2(new_n12995_), .A3(new_n13534_), .ZN(new_n13535_));
  INV_X1     g13343(.I(new_n13535_), .ZN(new_n13536_));
  NOR3_X1    g13344(.A1(new_n13534_), .A2(new_n12995_), .A3(new_n13003_), .ZN(new_n13537_));
  AOI22_X1   g13345(.A1(new_n13536_), .A2(new_n13003_), .B1(\asqrt[18] ), .B2(new_n13537_), .ZN(new_n13538_));
  NOR3_X1    g13346(.A1(new_n13531_), .A2(new_n13522_), .A3(\asqrt[31] ), .ZN(new_n13539_));
  NOR2_X1    g13347(.A1(new_n13539_), .A2(new_n13538_), .ZN(new_n13540_));
  OAI21_X1   g13348(.A1(new_n13540_), .A2(new_n13533_), .B(\asqrt[32] ), .ZN(new_n13541_));
  INV_X1     g13349(.I(new_n13010_), .ZN(new_n13542_));
  NOR3_X1    g13350(.A1(new_n13006_), .A2(new_n13542_), .A3(new_n13055_), .ZN(new_n13543_));
  NOR3_X1    g13351(.A1(new_n13353_), .A2(new_n13006_), .A3(new_n13055_), .ZN(new_n13544_));
  INV_X1     g13352(.I(new_n13544_), .ZN(new_n13545_));
  AOI22_X1   g13353(.A1(new_n13545_), .A2(new_n13542_), .B1(\asqrt[18] ), .B2(new_n13543_), .ZN(new_n13546_));
  INV_X1     g13354(.I(new_n13546_), .ZN(new_n13547_));
  NAND2_X1   g13355(.A1(new_n13532_), .A2(new_n6824_), .ZN(new_n13548_));
  OAI21_X1   g13356(.A1(new_n13540_), .A2(new_n13548_), .B(new_n13547_), .ZN(new_n13549_));
  AOI21_X1   g13357(.A1(new_n13549_), .A2(new_n13541_), .B(new_n6356_), .ZN(new_n13550_));
  NOR2_X1    g13358(.A1(new_n13028_), .A2(new_n13012_), .ZN(new_n13551_));
  INV_X1     g13359(.I(new_n13551_), .ZN(new_n13552_));
  NAND3_X1   g13360(.A1(\asqrt[18] ), .A2(new_n13013_), .A3(new_n13552_), .ZN(new_n13553_));
  AND3_X2    g13361(.A1(new_n13552_), .A2(new_n13013_), .A3(new_n13018_), .Z(new_n13554_));
  AOI22_X1   g13362(.A1(new_n13553_), .A2(new_n13019_), .B1(\asqrt[18] ), .B2(new_n13554_), .ZN(new_n13555_));
  OAI21_X1   g13363(.A1(new_n13538_), .A2(new_n13539_), .B(new_n13532_), .ZN(new_n13556_));
  AOI21_X1   g13364(.A1(new_n13556_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n13557_));
  AOI21_X1   g13365(.A1(new_n13557_), .A2(new_n13549_), .B(new_n13555_), .ZN(new_n13558_));
  OAI21_X1   g13366(.A1(new_n13558_), .A2(new_n13550_), .B(\asqrt[34] ), .ZN(new_n13559_));
  INV_X1     g13367(.I(new_n13559_), .ZN(new_n13560_));
  NOR2_X1    g13368(.A1(new_n13032_), .A2(new_n13039_), .ZN(new_n13561_));
  NOR3_X1    g13369(.A1(new_n13561_), .A2(new_n13030_), .A3(new_n13038_), .ZN(new_n13562_));
  NOR3_X1    g13370(.A1(new_n13353_), .A2(new_n13030_), .A3(new_n13561_), .ZN(new_n13563_));
  INV_X1     g13371(.I(new_n13563_), .ZN(new_n13564_));
  AOI22_X1   g13372(.A1(new_n13564_), .A2(new_n13038_), .B1(\asqrt[18] ), .B2(new_n13562_), .ZN(new_n13565_));
  NOR3_X1    g13373(.A1(new_n13558_), .A2(new_n13550_), .A3(\asqrt[34] ), .ZN(new_n13566_));
  NOR2_X1    g13374(.A1(new_n13566_), .A2(new_n13565_), .ZN(new_n13567_));
  OAI21_X1   g13375(.A1(new_n13567_), .A2(new_n13560_), .B(\asqrt[35] ), .ZN(new_n13568_));
  INV_X1     g13376(.I(new_n13045_), .ZN(new_n13569_));
  NOR3_X1    g13377(.A1(new_n13353_), .A2(new_n13041_), .A3(new_n13105_), .ZN(new_n13570_));
  INV_X1     g13378(.I(new_n13570_), .ZN(new_n13571_));
  NOR3_X1    g13379(.A1(new_n13041_), .A2(new_n13569_), .A3(new_n13105_), .ZN(new_n13572_));
  AOI22_X1   g13380(.A1(new_n13571_), .A2(new_n13569_), .B1(\asqrt[18] ), .B2(new_n13572_), .ZN(new_n13573_));
  INV_X1     g13381(.I(new_n13573_), .ZN(new_n13574_));
  NAND2_X1   g13382(.A1(new_n13559_), .A2(new_n5708_), .ZN(new_n13575_));
  OAI21_X1   g13383(.A1(new_n13567_), .A2(new_n13575_), .B(new_n13574_), .ZN(new_n13576_));
  AOI21_X1   g13384(.A1(new_n13576_), .A2(new_n13568_), .B(new_n5277_), .ZN(new_n13577_));
  NOR2_X1    g13385(.A1(new_n13060_), .A2(new_n13047_), .ZN(new_n13578_));
  INV_X1     g13386(.I(new_n13578_), .ZN(new_n13579_));
  AND3_X2    g13387(.A1(new_n13579_), .A2(new_n13048_), .A3(new_n13053_), .Z(new_n13580_));
  NAND3_X1   g13388(.A1(\asqrt[18] ), .A2(new_n13048_), .A3(new_n13579_), .ZN(new_n13581_));
  AOI22_X1   g13389(.A1(new_n13581_), .A2(new_n13054_), .B1(\asqrt[18] ), .B2(new_n13580_), .ZN(new_n13582_));
  OAI21_X1   g13390(.A1(new_n13565_), .A2(new_n13566_), .B(new_n13559_), .ZN(new_n13583_));
  AOI21_X1   g13391(.A1(new_n13583_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n13584_));
  AOI21_X1   g13392(.A1(new_n13584_), .A2(new_n13576_), .B(new_n13582_), .ZN(new_n13585_));
  OAI21_X1   g13393(.A1(new_n13585_), .A2(new_n13577_), .B(\asqrt[37] ), .ZN(new_n13586_));
  INV_X1     g13394(.I(new_n13586_), .ZN(new_n13587_));
  NOR2_X1    g13395(.A1(new_n13064_), .A2(new_n13071_), .ZN(new_n13588_));
  NOR3_X1    g13396(.A1(new_n13353_), .A2(new_n13078_), .A3(new_n13588_), .ZN(new_n13589_));
  INV_X1     g13397(.I(new_n13589_), .ZN(new_n13590_));
  NOR3_X1    g13398(.A1(new_n13588_), .A2(new_n13078_), .A3(new_n13070_), .ZN(new_n13591_));
  AOI22_X1   g13399(.A1(new_n13590_), .A2(new_n13070_), .B1(\asqrt[18] ), .B2(new_n13591_), .ZN(new_n13592_));
  NOR3_X1    g13400(.A1(new_n13585_), .A2(new_n13577_), .A3(\asqrt[37] ), .ZN(new_n13593_));
  NOR2_X1    g13401(.A1(new_n13593_), .A2(new_n13592_), .ZN(new_n13594_));
  OAI21_X1   g13402(.A1(new_n13594_), .A2(new_n13587_), .B(\asqrt[38] ), .ZN(new_n13595_));
  INV_X1     g13403(.I(new_n13077_), .ZN(new_n13596_));
  NOR3_X1    g13404(.A1(new_n13073_), .A2(new_n13596_), .A3(new_n13122_), .ZN(new_n13597_));
  NOR3_X1    g13405(.A1(new_n13353_), .A2(new_n13073_), .A3(new_n13122_), .ZN(new_n13598_));
  INV_X1     g13406(.I(new_n13598_), .ZN(new_n13599_));
  AOI22_X1   g13407(.A1(new_n13599_), .A2(new_n13596_), .B1(\asqrt[18] ), .B2(new_n13597_), .ZN(new_n13600_));
  INV_X1     g13408(.I(new_n13600_), .ZN(new_n13601_));
  NAND2_X1   g13409(.A1(new_n13586_), .A2(new_n4696_), .ZN(new_n13602_));
  OAI21_X1   g13410(.A1(new_n13594_), .A2(new_n13602_), .B(new_n13601_), .ZN(new_n13603_));
  AOI21_X1   g13411(.A1(new_n13603_), .A2(new_n13595_), .B(new_n4298_), .ZN(new_n13604_));
  NOR3_X1    g13412(.A1(new_n13353_), .A2(new_n13082_), .A3(new_n13088_), .ZN(new_n13605_));
  INV_X1     g13413(.I(new_n13605_), .ZN(new_n13606_));
  NOR3_X1    g13414(.A1(new_n13082_), .A2(new_n13104_), .A3(new_n13088_), .ZN(new_n13607_));
  AOI22_X1   g13415(.A1(new_n13606_), .A2(new_n13104_), .B1(\asqrt[18] ), .B2(new_n13607_), .ZN(new_n13608_));
  OAI21_X1   g13416(.A1(new_n13592_), .A2(new_n13593_), .B(new_n13586_), .ZN(new_n13609_));
  AOI21_X1   g13417(.A1(new_n13609_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n13610_));
  AOI21_X1   g13418(.A1(new_n13610_), .A2(new_n13603_), .B(new_n13608_), .ZN(new_n13611_));
  OAI21_X1   g13419(.A1(new_n13611_), .A2(new_n13604_), .B(\asqrt[40] ), .ZN(new_n13612_));
  INV_X1     g13420(.I(new_n13612_), .ZN(new_n13613_));
  NOR2_X1    g13421(.A1(new_n13089_), .A2(new_n13097_), .ZN(new_n13614_));
  NOR3_X1    g13422(.A1(new_n13614_), .A2(new_n13112_), .A3(new_n13096_), .ZN(new_n13615_));
  NOR3_X1    g13423(.A1(new_n13353_), .A2(new_n13112_), .A3(new_n13614_), .ZN(new_n13616_));
  INV_X1     g13424(.I(new_n13616_), .ZN(new_n13617_));
  AOI22_X1   g13425(.A1(new_n13617_), .A2(new_n13096_), .B1(\asqrt[18] ), .B2(new_n13615_), .ZN(new_n13618_));
  NOR3_X1    g13426(.A1(new_n13611_), .A2(new_n13604_), .A3(\asqrt[40] ), .ZN(new_n13619_));
  NOR2_X1    g13427(.A1(new_n13619_), .A2(new_n13618_), .ZN(new_n13620_));
  OAI21_X1   g13428(.A1(new_n13620_), .A2(new_n13613_), .B(\asqrt[41] ), .ZN(new_n13621_));
  INV_X1     g13429(.I(new_n13103_), .ZN(new_n13622_));
  NOR3_X1    g13430(.A1(new_n13353_), .A2(new_n13099_), .A3(new_n13135_), .ZN(new_n13623_));
  INV_X1     g13431(.I(new_n13623_), .ZN(new_n13624_));
  NOR3_X1    g13432(.A1(new_n13099_), .A2(new_n13622_), .A3(new_n13135_), .ZN(new_n13625_));
  AOI22_X1   g13433(.A1(new_n13624_), .A2(new_n13622_), .B1(\asqrt[18] ), .B2(new_n13625_), .ZN(new_n13626_));
  INV_X1     g13434(.I(new_n13626_), .ZN(new_n13627_));
  NAND2_X1   g13435(.A1(new_n13612_), .A2(new_n3782_), .ZN(new_n13628_));
  OAI21_X1   g13436(.A1(new_n13620_), .A2(new_n13628_), .B(new_n13627_), .ZN(new_n13629_));
  AOI21_X1   g13437(.A1(new_n13629_), .A2(new_n13621_), .B(new_n3419_), .ZN(new_n13630_));
  NOR3_X1    g13438(.A1(new_n13373_), .A2(new_n13121_), .A3(new_n13374_), .ZN(new_n13631_));
  NOR3_X1    g13439(.A1(new_n13353_), .A2(new_n13373_), .A3(new_n13374_), .ZN(new_n13632_));
  INV_X1     g13440(.I(new_n13632_), .ZN(new_n13633_));
  AOI22_X1   g13441(.A1(new_n13633_), .A2(new_n13121_), .B1(\asqrt[18] ), .B2(new_n13631_), .ZN(new_n13634_));
  OAI21_X1   g13442(.A1(new_n13618_), .A2(new_n13619_), .B(new_n13612_), .ZN(new_n13635_));
  AOI21_X1   g13443(.A1(new_n13635_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n13636_));
  AOI21_X1   g13444(.A1(new_n13636_), .A2(new_n13629_), .B(new_n13634_), .ZN(new_n13637_));
  OAI21_X1   g13445(.A1(new_n13637_), .A2(new_n13630_), .B(\asqrt[43] ), .ZN(new_n13638_));
  INV_X1     g13446(.I(new_n13638_), .ZN(new_n13639_));
  INV_X1     g13447(.I(new_n13134_), .ZN(new_n13640_));
  NAND2_X1   g13448(.A1(new_n13115_), .A2(new_n3419_), .ZN(new_n13641_));
  NOR2_X1    g13449(.A1(new_n13375_), .A2(new_n13641_), .ZN(new_n13642_));
  NOR3_X1    g13450(.A1(new_n13353_), .A2(new_n13129_), .A3(new_n13642_), .ZN(new_n13643_));
  INV_X1     g13451(.I(new_n13643_), .ZN(new_n13644_));
  NOR3_X1    g13452(.A1(new_n13642_), .A2(new_n13129_), .A3(new_n13640_), .ZN(new_n13645_));
  AOI22_X1   g13453(.A1(new_n13644_), .A2(new_n13640_), .B1(\asqrt[18] ), .B2(new_n13645_), .ZN(new_n13646_));
  NOR3_X1    g13454(.A1(new_n13637_), .A2(new_n13630_), .A3(\asqrt[43] ), .ZN(new_n13647_));
  NOR2_X1    g13455(.A1(new_n13647_), .A2(new_n13646_), .ZN(new_n13648_));
  OAI21_X1   g13456(.A1(new_n13648_), .A2(new_n13639_), .B(\asqrt[44] ), .ZN(new_n13649_));
  NOR3_X1    g13457(.A1(new_n13140_), .A2(new_n13145_), .A3(new_n13372_), .ZN(new_n13650_));
  NOR3_X1    g13458(.A1(new_n13353_), .A2(new_n13140_), .A3(new_n13145_), .ZN(new_n13651_));
  INV_X1     g13459(.I(new_n13651_), .ZN(new_n13652_));
  AOI22_X1   g13460(.A1(new_n13652_), .A2(new_n13372_), .B1(\asqrt[18] ), .B2(new_n13650_), .ZN(new_n13653_));
  INV_X1     g13461(.I(new_n13653_), .ZN(new_n13654_));
  NAND2_X1   g13462(.A1(new_n13638_), .A2(new_n2954_), .ZN(new_n13655_));
  OAI21_X1   g13463(.A1(new_n13648_), .A2(new_n13655_), .B(new_n13654_), .ZN(new_n13656_));
  AOI21_X1   g13464(.A1(new_n13656_), .A2(new_n13649_), .B(new_n2641_), .ZN(new_n13657_));
  INV_X1     g13465(.I(new_n13147_), .ZN(new_n13658_));
  NOR2_X1    g13466(.A1(new_n13146_), .A2(new_n13154_), .ZN(new_n13659_));
  NOR3_X1    g13467(.A1(new_n13353_), .A2(new_n13658_), .A3(new_n13659_), .ZN(new_n13660_));
  INV_X1     g13468(.I(new_n13660_), .ZN(new_n13661_));
  NOR3_X1    g13469(.A1(new_n13658_), .A2(new_n13659_), .A3(new_n13153_), .ZN(new_n13662_));
  AOI22_X1   g13470(.A1(new_n13661_), .A2(new_n13153_), .B1(\asqrt[18] ), .B2(new_n13662_), .ZN(new_n13663_));
  OAI21_X1   g13471(.A1(new_n13646_), .A2(new_n13647_), .B(new_n13638_), .ZN(new_n13664_));
  AOI21_X1   g13472(.A1(new_n13664_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n13665_));
  AOI21_X1   g13473(.A1(new_n13665_), .A2(new_n13656_), .B(new_n13663_), .ZN(new_n13666_));
  OAI21_X1   g13474(.A1(new_n13666_), .A2(new_n13657_), .B(\asqrt[46] ), .ZN(new_n13667_));
  INV_X1     g13475(.I(new_n13667_), .ZN(new_n13668_));
  INV_X1     g13476(.I(new_n13161_), .ZN(new_n13669_));
  INV_X1     g13477(.I(new_n13155_), .ZN(new_n13670_));
  INV_X1     g13478(.I(new_n13163_), .ZN(new_n13671_));
  NOR2_X1    g13479(.A1(new_n13671_), .A2(new_n13670_), .ZN(new_n13672_));
  NOR3_X1    g13480(.A1(new_n13672_), .A2(new_n13156_), .A3(new_n13669_), .ZN(new_n13673_));
  NOR3_X1    g13481(.A1(new_n13353_), .A2(new_n13156_), .A3(new_n13672_), .ZN(new_n13674_));
  INV_X1     g13482(.I(new_n13674_), .ZN(new_n13675_));
  AOI22_X1   g13483(.A1(new_n13675_), .A2(new_n13669_), .B1(\asqrt[18] ), .B2(new_n13673_), .ZN(new_n13676_));
  NOR3_X1    g13484(.A1(new_n13666_), .A2(new_n13657_), .A3(\asqrt[46] ), .ZN(new_n13677_));
  NOR2_X1    g13485(.A1(new_n13677_), .A2(new_n13676_), .ZN(new_n13678_));
  OAI21_X1   g13486(.A1(new_n13678_), .A2(new_n13668_), .B(\asqrt[47] ), .ZN(new_n13679_));
  NOR3_X1    g13487(.A1(new_n13353_), .A2(new_n13166_), .A3(new_n13171_), .ZN(new_n13680_));
  INV_X1     g13488(.I(new_n13680_), .ZN(new_n13681_));
  NOR3_X1    g13489(.A1(new_n13166_), .A2(new_n13371_), .A3(new_n13171_), .ZN(new_n13682_));
  AOI22_X1   g13490(.A1(new_n13681_), .A2(new_n13371_), .B1(\asqrt[18] ), .B2(new_n13682_), .ZN(new_n13683_));
  INV_X1     g13491(.I(new_n13683_), .ZN(new_n13684_));
  NAND2_X1   g13492(.A1(new_n13667_), .A2(new_n2229_), .ZN(new_n13685_));
  OAI21_X1   g13493(.A1(new_n13678_), .A2(new_n13685_), .B(new_n13684_), .ZN(new_n13686_));
  AOI21_X1   g13494(.A1(new_n13686_), .A2(new_n13679_), .B(new_n1956_), .ZN(new_n13687_));
  INV_X1     g13495(.I(new_n13173_), .ZN(new_n13688_));
  NOR2_X1    g13496(.A1(new_n13172_), .A2(new_n13180_), .ZN(new_n13689_));
  NOR3_X1    g13497(.A1(new_n13688_), .A2(new_n13689_), .A3(new_n13179_), .ZN(new_n13690_));
  NOR3_X1    g13498(.A1(new_n13353_), .A2(new_n13688_), .A3(new_n13689_), .ZN(new_n13691_));
  INV_X1     g13499(.I(new_n13691_), .ZN(new_n13692_));
  AOI22_X1   g13500(.A1(new_n13692_), .A2(new_n13179_), .B1(\asqrt[18] ), .B2(new_n13690_), .ZN(new_n13693_));
  OAI21_X1   g13501(.A1(new_n13676_), .A2(new_n13677_), .B(new_n13667_), .ZN(new_n13694_));
  AOI21_X1   g13502(.A1(new_n13694_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n13695_));
  AOI21_X1   g13503(.A1(new_n13695_), .A2(new_n13686_), .B(new_n13693_), .ZN(new_n13696_));
  OAI21_X1   g13504(.A1(new_n13696_), .A2(new_n13687_), .B(\asqrt[49] ), .ZN(new_n13697_));
  INV_X1     g13505(.I(new_n13697_), .ZN(new_n13698_));
  INV_X1     g13506(.I(new_n13187_), .ZN(new_n13699_));
  INV_X1     g13507(.I(new_n13181_), .ZN(new_n13700_));
  INV_X1     g13508(.I(new_n13189_), .ZN(new_n13701_));
  NOR2_X1    g13509(.A1(new_n13701_), .A2(new_n13700_), .ZN(new_n13702_));
  NOR3_X1    g13510(.A1(new_n13353_), .A2(new_n13182_), .A3(new_n13702_), .ZN(new_n13703_));
  INV_X1     g13511(.I(new_n13703_), .ZN(new_n13704_));
  NOR3_X1    g13512(.A1(new_n13702_), .A2(new_n13182_), .A3(new_n13699_), .ZN(new_n13705_));
  AOI22_X1   g13513(.A1(new_n13704_), .A2(new_n13699_), .B1(\asqrt[18] ), .B2(new_n13705_), .ZN(new_n13706_));
  NOR3_X1    g13514(.A1(new_n13696_), .A2(new_n13687_), .A3(\asqrt[49] ), .ZN(new_n13707_));
  NOR2_X1    g13515(.A1(new_n13707_), .A2(new_n13706_), .ZN(new_n13708_));
  OAI21_X1   g13516(.A1(new_n13708_), .A2(new_n13698_), .B(\asqrt[50] ), .ZN(new_n13709_));
  NOR3_X1    g13517(.A1(new_n13192_), .A2(new_n13370_), .A3(new_n13197_), .ZN(new_n13710_));
  NOR3_X1    g13518(.A1(new_n13353_), .A2(new_n13192_), .A3(new_n13197_), .ZN(new_n13711_));
  INV_X1     g13519(.I(new_n13711_), .ZN(new_n13712_));
  AOI22_X1   g13520(.A1(new_n13712_), .A2(new_n13370_), .B1(\asqrt[18] ), .B2(new_n13710_), .ZN(new_n13713_));
  INV_X1     g13521(.I(new_n13713_), .ZN(new_n13714_));
  NAND2_X1   g13522(.A1(new_n13697_), .A2(new_n1612_), .ZN(new_n13715_));
  OAI21_X1   g13523(.A1(new_n13708_), .A2(new_n13715_), .B(new_n13714_), .ZN(new_n13716_));
  AOI21_X1   g13524(.A1(new_n13716_), .A2(new_n13709_), .B(new_n1376_), .ZN(new_n13717_));
  INV_X1     g13525(.I(new_n13199_), .ZN(new_n13718_));
  NOR2_X1    g13526(.A1(new_n13198_), .A2(new_n13206_), .ZN(new_n13719_));
  NOR3_X1    g13527(.A1(new_n13353_), .A2(new_n13718_), .A3(new_n13719_), .ZN(new_n13720_));
  INV_X1     g13528(.I(new_n13720_), .ZN(new_n13721_));
  NOR3_X1    g13529(.A1(new_n13718_), .A2(new_n13205_), .A3(new_n13719_), .ZN(new_n13722_));
  AOI22_X1   g13530(.A1(new_n13721_), .A2(new_n13205_), .B1(\asqrt[18] ), .B2(new_n13722_), .ZN(new_n13723_));
  OAI21_X1   g13531(.A1(new_n13706_), .A2(new_n13707_), .B(new_n13697_), .ZN(new_n13724_));
  AOI21_X1   g13532(.A1(new_n13724_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n13725_));
  AOI21_X1   g13533(.A1(new_n13725_), .A2(new_n13716_), .B(new_n13723_), .ZN(new_n13726_));
  OAI21_X1   g13534(.A1(new_n13726_), .A2(new_n13717_), .B(\asqrt[52] ), .ZN(new_n13727_));
  INV_X1     g13535(.I(new_n13727_), .ZN(new_n13728_));
  INV_X1     g13536(.I(new_n13213_), .ZN(new_n13729_));
  INV_X1     g13537(.I(new_n13207_), .ZN(new_n13730_));
  INV_X1     g13538(.I(new_n13215_), .ZN(new_n13731_));
  NOR2_X1    g13539(.A1(new_n13731_), .A2(new_n13730_), .ZN(new_n13732_));
  NOR3_X1    g13540(.A1(new_n13732_), .A2(new_n13208_), .A3(new_n13729_), .ZN(new_n13733_));
  NOR3_X1    g13541(.A1(new_n13353_), .A2(new_n13208_), .A3(new_n13732_), .ZN(new_n13734_));
  INV_X1     g13542(.I(new_n13734_), .ZN(new_n13735_));
  AOI22_X1   g13543(.A1(new_n13735_), .A2(new_n13729_), .B1(\asqrt[18] ), .B2(new_n13733_), .ZN(new_n13736_));
  NOR3_X1    g13544(.A1(new_n13726_), .A2(new_n13717_), .A3(\asqrt[52] ), .ZN(new_n13737_));
  NOR2_X1    g13545(.A1(new_n13737_), .A2(new_n13736_), .ZN(new_n13738_));
  OAI21_X1   g13546(.A1(new_n13738_), .A2(new_n13728_), .B(\asqrt[53] ), .ZN(new_n13739_));
  NOR3_X1    g13547(.A1(new_n13353_), .A2(new_n13218_), .A3(new_n13260_), .ZN(new_n13740_));
  INV_X1     g13548(.I(new_n13740_), .ZN(new_n13741_));
  NOR3_X1    g13549(.A1(new_n13218_), .A2(new_n13369_), .A3(new_n13260_), .ZN(new_n13742_));
  AOI22_X1   g13550(.A1(new_n13741_), .A2(new_n13369_), .B1(\asqrt[18] ), .B2(new_n13742_), .ZN(new_n13743_));
  INV_X1     g13551(.I(new_n13743_), .ZN(new_n13744_));
  NAND2_X1   g13552(.A1(new_n13727_), .A2(new_n1103_), .ZN(new_n13745_));
  OAI21_X1   g13553(.A1(new_n13738_), .A2(new_n13745_), .B(new_n13744_), .ZN(new_n13746_));
  AOI21_X1   g13554(.A1(new_n13746_), .A2(new_n13739_), .B(new_n904_), .ZN(new_n13747_));
  INV_X1     g13555(.I(new_n13226_), .ZN(new_n13748_));
  NOR2_X1    g13556(.A1(new_n13233_), .A2(new_n13225_), .ZN(new_n13749_));
  NOR3_X1    g13557(.A1(new_n13748_), .A2(new_n13232_), .A3(new_n13749_), .ZN(new_n13750_));
  NOR3_X1    g13558(.A1(new_n13353_), .A2(new_n13748_), .A3(new_n13749_), .ZN(new_n13751_));
  INV_X1     g13559(.I(new_n13751_), .ZN(new_n13752_));
  AOI22_X1   g13560(.A1(new_n13752_), .A2(new_n13232_), .B1(\asqrt[18] ), .B2(new_n13750_), .ZN(new_n13753_));
  OAI21_X1   g13561(.A1(new_n13736_), .A2(new_n13737_), .B(new_n13727_), .ZN(new_n13754_));
  AOI21_X1   g13562(.A1(new_n13754_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n13755_));
  AOI21_X1   g13563(.A1(new_n13755_), .A2(new_n13746_), .B(new_n13753_), .ZN(new_n13756_));
  OAI21_X1   g13564(.A1(new_n13756_), .A2(new_n13747_), .B(\asqrt[55] ), .ZN(new_n13757_));
  INV_X1     g13565(.I(new_n13757_), .ZN(new_n13758_));
  NOR2_X1    g13566(.A1(new_n13244_), .A2(new_n13237_), .ZN(new_n13759_));
  NOR3_X1    g13567(.A1(new_n13353_), .A2(new_n13235_), .A3(new_n13759_), .ZN(new_n13760_));
  INV_X1     g13568(.I(new_n13760_), .ZN(new_n13761_));
  NOR3_X1    g13569(.A1(new_n13759_), .A2(new_n13235_), .A3(new_n13243_), .ZN(new_n13762_));
  AOI22_X1   g13570(.A1(new_n13761_), .A2(new_n13243_), .B1(\asqrt[18] ), .B2(new_n13762_), .ZN(new_n13763_));
  NOR3_X1    g13571(.A1(new_n13756_), .A2(new_n13747_), .A3(\asqrt[55] ), .ZN(new_n13764_));
  NOR2_X1    g13572(.A1(new_n13764_), .A2(new_n13763_), .ZN(new_n13765_));
  OAI21_X1   g13573(.A1(new_n13765_), .A2(new_n13758_), .B(\asqrt[56] ), .ZN(new_n13766_));
  NOR3_X1    g13574(.A1(new_n13246_), .A2(new_n13368_), .A3(new_n13292_), .ZN(new_n13767_));
  NOR3_X1    g13575(.A1(new_n13353_), .A2(new_n13246_), .A3(new_n13292_), .ZN(new_n13768_));
  INV_X1     g13576(.I(new_n13768_), .ZN(new_n13769_));
  AOI22_X1   g13577(.A1(new_n13769_), .A2(new_n13368_), .B1(\asqrt[18] ), .B2(new_n13767_), .ZN(new_n13770_));
  INV_X1     g13578(.I(new_n13770_), .ZN(new_n13771_));
  NAND2_X1   g13579(.A1(new_n13757_), .A2(new_n703_), .ZN(new_n13772_));
  OAI21_X1   g13580(.A1(new_n13765_), .A2(new_n13772_), .B(new_n13771_), .ZN(new_n13773_));
  AOI21_X1   g13581(.A1(new_n13773_), .A2(new_n13766_), .B(new_n531_), .ZN(new_n13774_));
  INV_X1     g13582(.I(new_n13253_), .ZN(new_n13775_));
  NOR2_X1    g13583(.A1(new_n13265_), .A2(new_n13252_), .ZN(new_n13776_));
  NOR3_X1    g13584(.A1(new_n13353_), .A2(new_n13775_), .A3(new_n13776_), .ZN(new_n13777_));
  INV_X1     g13585(.I(new_n13777_), .ZN(new_n13778_));
  NOR3_X1    g13586(.A1(new_n13775_), .A2(new_n13259_), .A3(new_n13776_), .ZN(new_n13779_));
  AOI22_X1   g13587(.A1(new_n13778_), .A2(new_n13259_), .B1(\asqrt[18] ), .B2(new_n13779_), .ZN(new_n13780_));
  OAI21_X1   g13588(.A1(new_n13763_), .A2(new_n13764_), .B(new_n13757_), .ZN(new_n13781_));
  AOI21_X1   g13589(.A1(new_n13781_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n13782_));
  AOI21_X1   g13590(.A1(new_n13782_), .A2(new_n13773_), .B(new_n13780_), .ZN(new_n13783_));
  OAI21_X1   g13591(.A1(new_n13783_), .A2(new_n13774_), .B(\asqrt[58] ), .ZN(new_n13784_));
  NOR2_X1    g13592(.A1(new_n13276_), .A2(new_n13269_), .ZN(new_n13785_));
  NOR3_X1    g13593(.A1(new_n13785_), .A2(new_n13267_), .A3(new_n13275_), .ZN(new_n13786_));
  NOR3_X1    g13594(.A1(new_n13353_), .A2(new_n13267_), .A3(new_n13785_), .ZN(new_n13787_));
  INV_X1     g13595(.I(new_n13787_), .ZN(new_n13788_));
  AOI22_X1   g13596(.A1(new_n13788_), .A2(new_n13275_), .B1(\asqrt[18] ), .B2(new_n13786_), .ZN(new_n13789_));
  INV_X1     g13597(.I(new_n13789_), .ZN(new_n13790_));
  INV_X1     g13598(.I(new_n13763_), .ZN(new_n13791_));
  INV_X1     g13599(.I(new_n13736_), .ZN(new_n13792_));
  INV_X1     g13600(.I(new_n13706_), .ZN(new_n13793_));
  INV_X1     g13601(.I(new_n13676_), .ZN(new_n13794_));
  INV_X1     g13602(.I(new_n13646_), .ZN(new_n13795_));
  INV_X1     g13603(.I(new_n13618_), .ZN(new_n13796_));
  INV_X1     g13604(.I(new_n13592_), .ZN(new_n13797_));
  INV_X1     g13605(.I(new_n13565_), .ZN(new_n13798_));
  INV_X1     g13606(.I(new_n13538_), .ZN(new_n13799_));
  INV_X1     g13607(.I(new_n13510_), .ZN(new_n13800_));
  INV_X1     g13608(.I(new_n13484_), .ZN(new_n13801_));
  NAND2_X1   g13609(.A1(new_n13426_), .A2(new_n11326_), .ZN(new_n13802_));
  OAI21_X1   g13610(.A1(new_n13802_), .A2(new_n13458_), .B(new_n13440_), .ZN(new_n13803_));
  AOI21_X1   g13611(.A1(new_n13803_), .A2(new_n13468_), .B(new_n10812_), .ZN(new_n13804_));
  NOR2_X1    g13612(.A1(new_n13434_), .A2(\asqrt[23] ), .ZN(new_n13805_));
  AOI21_X1   g13613(.A1(new_n13805_), .A2(new_n13803_), .B(new_n13466_), .ZN(new_n13806_));
  OAI21_X1   g13614(.A1(new_n13806_), .A2(new_n13804_), .B(\asqrt[24] ), .ZN(new_n13807_));
  NAND2_X1   g13615(.A1(new_n13807_), .A2(new_n9846_), .ZN(new_n13808_));
  OAI21_X1   g13616(.A1(new_n13808_), .A2(new_n13478_), .B(new_n13801_), .ZN(new_n13809_));
  NAND3_X1   g13617(.A1(new_n13809_), .A2(new_n9317_), .A3(new_n13479_), .ZN(new_n13810_));
  AOI22_X1   g13618(.A1(new_n13810_), .A2(new_n13493_), .B1(\asqrt[26] ), .B2(new_n13501_), .ZN(new_n13811_));
  OAI21_X1   g13619(.A1(new_n13811_), .A2(new_n8826_), .B(new_n8483_), .ZN(new_n13812_));
  OAI21_X1   g13620(.A1(new_n13812_), .A2(new_n13503_), .B(new_n13800_), .ZN(new_n13813_));
  AOI21_X1   g13621(.A1(new_n13813_), .A2(new_n13504_), .B(new_n8036_), .ZN(new_n13814_));
  AOI21_X1   g13622(.A1(new_n13809_), .A2(new_n13479_), .B(new_n9317_), .ZN(new_n13815_));
  NOR3_X1    g13623(.A1(new_n13806_), .A2(new_n13804_), .A3(\asqrt[24] ), .ZN(new_n13816_));
  OAI21_X1   g13624(.A1(new_n13475_), .A2(new_n13816_), .B(new_n13807_), .ZN(new_n13817_));
  AOI21_X1   g13625(.A1(new_n13817_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n13818_));
  AOI21_X1   g13626(.A1(new_n13818_), .A2(new_n13809_), .B(new_n13492_), .ZN(new_n13819_));
  NOR3_X1    g13627(.A1(new_n13819_), .A2(\asqrt[27] ), .A3(new_n13815_), .ZN(new_n13820_));
  OAI22_X1   g13628(.A1(new_n13820_), .A2(new_n13500_), .B1(new_n13811_), .B2(new_n8826_), .ZN(new_n13821_));
  AOI21_X1   g13629(.A1(new_n13821_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n13822_));
  AOI21_X1   g13630(.A1(new_n13822_), .A2(new_n13813_), .B(new_n13518_), .ZN(new_n13823_));
  OAI21_X1   g13631(.A1(new_n13823_), .A2(new_n13814_), .B(\asqrt[30] ), .ZN(new_n13824_));
  NAND2_X1   g13632(.A1(new_n13824_), .A2(new_n7229_), .ZN(new_n13825_));
  OAI21_X1   g13633(.A1(new_n13825_), .A2(new_n13531_), .B(new_n13799_), .ZN(new_n13826_));
  AOI21_X1   g13634(.A1(new_n13826_), .A2(new_n13532_), .B(new_n6824_), .ZN(new_n13827_));
  NOR3_X1    g13635(.A1(new_n13823_), .A2(\asqrt[30] ), .A3(new_n13814_), .ZN(new_n13828_));
  OAI21_X1   g13636(.A1(new_n13528_), .A2(new_n13828_), .B(new_n13824_), .ZN(new_n13829_));
  AOI21_X1   g13637(.A1(new_n13829_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n13830_));
  AOI21_X1   g13638(.A1(new_n13830_), .A2(new_n13826_), .B(new_n13546_), .ZN(new_n13831_));
  OAI21_X1   g13639(.A1(new_n13831_), .A2(new_n13827_), .B(\asqrt[33] ), .ZN(new_n13832_));
  NAND2_X1   g13640(.A1(new_n13832_), .A2(new_n6077_), .ZN(new_n13833_));
  OAI21_X1   g13641(.A1(new_n13833_), .A2(new_n13558_), .B(new_n13798_), .ZN(new_n13834_));
  AOI21_X1   g13642(.A1(new_n13834_), .A2(new_n13559_), .B(new_n5708_), .ZN(new_n13835_));
  NOR3_X1    g13643(.A1(new_n13831_), .A2(\asqrt[33] ), .A3(new_n13827_), .ZN(new_n13836_));
  OAI21_X1   g13644(.A1(new_n13555_), .A2(new_n13836_), .B(new_n13832_), .ZN(new_n13837_));
  AOI21_X1   g13645(.A1(new_n13837_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n13838_));
  AOI21_X1   g13646(.A1(new_n13838_), .A2(new_n13834_), .B(new_n13573_), .ZN(new_n13839_));
  OAI21_X1   g13647(.A1(new_n13839_), .A2(new_n13835_), .B(\asqrt[36] ), .ZN(new_n13840_));
  NAND2_X1   g13648(.A1(new_n13840_), .A2(new_n5024_), .ZN(new_n13841_));
  OAI21_X1   g13649(.A1(new_n13841_), .A2(new_n13585_), .B(new_n13797_), .ZN(new_n13842_));
  AOI21_X1   g13650(.A1(new_n13842_), .A2(new_n13586_), .B(new_n4696_), .ZN(new_n13843_));
  NOR3_X1    g13651(.A1(new_n13839_), .A2(\asqrt[36] ), .A3(new_n13835_), .ZN(new_n13844_));
  OAI21_X1   g13652(.A1(new_n13582_), .A2(new_n13844_), .B(new_n13840_), .ZN(new_n13845_));
  AOI21_X1   g13653(.A1(new_n13845_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n13846_));
  AOI21_X1   g13654(.A1(new_n13846_), .A2(new_n13842_), .B(new_n13600_), .ZN(new_n13847_));
  OAI21_X1   g13655(.A1(new_n13847_), .A2(new_n13843_), .B(\asqrt[39] ), .ZN(new_n13848_));
  NAND2_X1   g13656(.A1(new_n13848_), .A2(new_n4071_), .ZN(new_n13849_));
  OAI21_X1   g13657(.A1(new_n13849_), .A2(new_n13611_), .B(new_n13796_), .ZN(new_n13850_));
  AOI21_X1   g13658(.A1(new_n13850_), .A2(new_n13612_), .B(new_n3782_), .ZN(new_n13851_));
  NOR3_X1    g13659(.A1(new_n13847_), .A2(\asqrt[39] ), .A3(new_n13843_), .ZN(new_n13852_));
  OAI21_X1   g13660(.A1(new_n13608_), .A2(new_n13852_), .B(new_n13848_), .ZN(new_n13853_));
  AOI21_X1   g13661(.A1(new_n13853_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n13854_));
  AOI21_X1   g13662(.A1(new_n13854_), .A2(new_n13850_), .B(new_n13626_), .ZN(new_n13855_));
  OAI21_X1   g13663(.A1(new_n13855_), .A2(new_n13851_), .B(\asqrt[42] ), .ZN(new_n13856_));
  NAND2_X1   g13664(.A1(new_n13856_), .A2(new_n3218_), .ZN(new_n13857_));
  OAI21_X1   g13665(.A1(new_n13857_), .A2(new_n13637_), .B(new_n13795_), .ZN(new_n13858_));
  AOI21_X1   g13666(.A1(new_n13858_), .A2(new_n13638_), .B(new_n2954_), .ZN(new_n13859_));
  NOR3_X1    g13667(.A1(new_n13855_), .A2(\asqrt[42] ), .A3(new_n13851_), .ZN(new_n13860_));
  OAI21_X1   g13668(.A1(new_n13634_), .A2(new_n13860_), .B(new_n13856_), .ZN(new_n13861_));
  AOI21_X1   g13669(.A1(new_n13861_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n13862_));
  AOI21_X1   g13670(.A1(new_n13862_), .A2(new_n13858_), .B(new_n13653_), .ZN(new_n13863_));
  OAI21_X1   g13671(.A1(new_n13863_), .A2(new_n13859_), .B(\asqrt[45] ), .ZN(new_n13864_));
  NAND2_X1   g13672(.A1(new_n13864_), .A2(new_n2465_), .ZN(new_n13865_));
  OAI21_X1   g13673(.A1(new_n13865_), .A2(new_n13666_), .B(new_n13794_), .ZN(new_n13866_));
  AOI21_X1   g13674(.A1(new_n13866_), .A2(new_n13667_), .B(new_n2229_), .ZN(new_n13867_));
  NOR3_X1    g13675(.A1(new_n13863_), .A2(\asqrt[45] ), .A3(new_n13859_), .ZN(new_n13868_));
  OAI21_X1   g13676(.A1(new_n13663_), .A2(new_n13868_), .B(new_n13864_), .ZN(new_n13869_));
  AOI21_X1   g13677(.A1(new_n13869_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n13870_));
  AOI21_X1   g13678(.A1(new_n13870_), .A2(new_n13866_), .B(new_n13683_), .ZN(new_n13871_));
  OAI21_X1   g13679(.A1(new_n13871_), .A2(new_n13867_), .B(\asqrt[48] ), .ZN(new_n13872_));
  NAND2_X1   g13680(.A1(new_n13872_), .A2(new_n1806_), .ZN(new_n13873_));
  OAI21_X1   g13681(.A1(new_n13873_), .A2(new_n13696_), .B(new_n13793_), .ZN(new_n13874_));
  AOI21_X1   g13682(.A1(new_n13874_), .A2(new_n13697_), .B(new_n1612_), .ZN(new_n13875_));
  NOR3_X1    g13683(.A1(new_n13871_), .A2(\asqrt[48] ), .A3(new_n13867_), .ZN(new_n13876_));
  OAI21_X1   g13684(.A1(new_n13693_), .A2(new_n13876_), .B(new_n13872_), .ZN(new_n13877_));
  AOI21_X1   g13685(.A1(new_n13877_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n13878_));
  AOI21_X1   g13686(.A1(new_n13878_), .A2(new_n13874_), .B(new_n13713_), .ZN(new_n13879_));
  OAI21_X1   g13687(.A1(new_n13879_), .A2(new_n13875_), .B(\asqrt[51] ), .ZN(new_n13880_));
  NAND2_X1   g13688(.A1(new_n13880_), .A2(new_n1256_), .ZN(new_n13881_));
  OAI21_X1   g13689(.A1(new_n13881_), .A2(new_n13726_), .B(new_n13792_), .ZN(new_n13882_));
  NAND3_X1   g13690(.A1(new_n13882_), .A2(new_n1103_), .A3(new_n13727_), .ZN(new_n13883_));
  AOI22_X1   g13691(.A1(new_n13883_), .A2(new_n13744_), .B1(\asqrt[53] ), .B2(new_n13754_), .ZN(new_n13884_));
  OAI21_X1   g13692(.A1(new_n13884_), .A2(new_n904_), .B(new_n823_), .ZN(new_n13885_));
  OAI21_X1   g13693(.A1(new_n13885_), .A2(new_n13756_), .B(new_n13791_), .ZN(new_n13886_));
  NAND3_X1   g13694(.A1(new_n13886_), .A2(new_n703_), .A3(new_n13757_), .ZN(new_n13887_));
  AOI22_X1   g13695(.A1(new_n13887_), .A2(new_n13771_), .B1(\asqrt[56] ), .B2(new_n13781_), .ZN(new_n13888_));
  OAI21_X1   g13696(.A1(new_n13888_), .A2(new_n531_), .B(new_n436_), .ZN(new_n13889_));
  OAI21_X1   g13697(.A1(new_n13889_), .A2(new_n13783_), .B(new_n13790_), .ZN(new_n13890_));
  AOI21_X1   g13698(.A1(new_n13890_), .A2(new_n13784_), .B(new_n327_), .ZN(new_n13891_));
  NOR3_X1    g13699(.A1(new_n13353_), .A2(new_n13278_), .A3(new_n13324_), .ZN(new_n13892_));
  INV_X1     g13700(.I(new_n13892_), .ZN(new_n13893_));
  NOR3_X1    g13701(.A1(new_n13278_), .A2(new_n13367_), .A3(new_n13324_), .ZN(new_n13894_));
  AOI22_X1   g13702(.A1(new_n13893_), .A2(new_n13367_), .B1(\asqrt[18] ), .B2(new_n13894_), .ZN(new_n13895_));
  NAND2_X1   g13703(.A1(new_n13784_), .A2(new_n327_), .ZN(new_n13896_));
  INV_X1     g13704(.I(new_n13896_), .ZN(new_n13897_));
  AOI21_X1   g13705(.A1(new_n13897_), .A2(new_n13890_), .B(new_n13895_), .ZN(new_n13898_));
  OAI21_X1   g13706(.A1(new_n13898_), .A2(new_n13891_), .B(\asqrt[60] ), .ZN(new_n13899_));
  INV_X1     g13707(.I(new_n13285_), .ZN(new_n13900_));
  NOR2_X1    g13708(.A1(new_n13297_), .A2(new_n13284_), .ZN(new_n13901_));
  NOR3_X1    g13709(.A1(new_n13900_), .A2(new_n13291_), .A3(new_n13901_), .ZN(new_n13902_));
  NOR3_X1    g13710(.A1(new_n13353_), .A2(new_n13900_), .A3(new_n13901_), .ZN(new_n13903_));
  INV_X1     g13711(.I(new_n13903_), .ZN(new_n13904_));
  AOI22_X1   g13712(.A1(new_n13904_), .A2(new_n13291_), .B1(\asqrt[18] ), .B2(new_n13902_), .ZN(new_n13905_));
  INV_X1     g13713(.I(new_n13905_), .ZN(new_n13906_));
  INV_X1     g13714(.I(new_n13784_), .ZN(new_n13907_));
  NOR3_X1    g13715(.A1(new_n13783_), .A2(new_n13774_), .A3(\asqrt[58] ), .ZN(new_n13908_));
  NOR2_X1    g13716(.A1(new_n13908_), .A2(new_n13789_), .ZN(new_n13909_));
  OAI21_X1   g13717(.A1(new_n13909_), .A2(new_n13907_), .B(\asqrt[59] ), .ZN(new_n13910_));
  NAND2_X1   g13718(.A1(new_n13910_), .A2(new_n306_), .ZN(new_n13911_));
  OAI21_X1   g13719(.A1(new_n13911_), .A2(new_n13898_), .B(new_n13906_), .ZN(new_n13912_));
  AOI21_X1   g13720(.A1(new_n13912_), .A2(new_n13899_), .B(new_n218_), .ZN(new_n13913_));
  NOR2_X1    g13721(.A1(new_n13301_), .A2(new_n13308_), .ZN(new_n13914_));
  NOR3_X1    g13722(.A1(new_n13353_), .A2(new_n13299_), .A3(new_n13914_), .ZN(new_n13915_));
  INV_X1     g13723(.I(new_n13915_), .ZN(new_n13916_));
  NOR3_X1    g13724(.A1(new_n13914_), .A2(new_n13299_), .A3(new_n13307_), .ZN(new_n13917_));
  AOI22_X1   g13725(.A1(new_n13916_), .A2(new_n13307_), .B1(\asqrt[18] ), .B2(new_n13917_), .ZN(new_n13918_));
  INV_X1     g13726(.I(new_n13895_), .ZN(new_n13919_));
  OAI21_X1   g13727(.A1(new_n13909_), .A2(new_n13896_), .B(new_n13919_), .ZN(new_n13920_));
  AOI21_X1   g13728(.A1(new_n13920_), .A2(new_n13910_), .B(new_n306_), .ZN(new_n13921_));
  NOR2_X1    g13729(.A1(new_n13921_), .A2(\asqrt[61] ), .ZN(new_n13922_));
  AOI21_X1   g13730(.A1(new_n13922_), .A2(new_n13912_), .B(new_n13918_), .ZN(new_n13923_));
  OAI21_X1   g13731(.A1(new_n13923_), .A2(new_n13913_), .B(\asqrt[62] ), .ZN(new_n13924_));
  NOR3_X1    g13732(.A1(new_n13310_), .A2(new_n13366_), .A3(new_n13364_), .ZN(new_n13925_));
  NOR3_X1    g13733(.A1(new_n13353_), .A2(new_n13310_), .A3(new_n13364_), .ZN(new_n13926_));
  INV_X1     g13734(.I(new_n13926_), .ZN(new_n13927_));
  AOI22_X1   g13735(.A1(new_n13927_), .A2(new_n13366_), .B1(\asqrt[18] ), .B2(new_n13925_), .ZN(new_n13928_));
  INV_X1     g13736(.I(new_n13928_), .ZN(new_n13929_));
  OAI21_X1   g13737(.A1(new_n13789_), .A2(new_n13908_), .B(new_n13784_), .ZN(new_n13930_));
  AOI21_X1   g13738(.A1(new_n13930_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n13931_));
  AOI21_X1   g13739(.A1(new_n13931_), .A2(new_n13920_), .B(new_n13905_), .ZN(new_n13932_));
  OAI21_X1   g13740(.A1(new_n13932_), .A2(new_n13921_), .B(\asqrt[61] ), .ZN(new_n13933_));
  NAND2_X1   g13741(.A1(new_n13933_), .A2(new_n207_), .ZN(new_n13934_));
  OAI21_X1   g13742(.A1(new_n13934_), .A2(new_n13923_), .B(new_n13929_), .ZN(new_n13935_));
  NAND4_X1   g13743(.A1(\asqrt[18] ), .A2(new_n13317_), .A3(new_n13322_), .A4(new_n13403_), .ZN(new_n13936_));
  NAND2_X1   g13744(.A1(new_n13317_), .A2(new_n13403_), .ZN(new_n13937_));
  OAI21_X1   g13745(.A1(new_n13353_), .A2(new_n13937_), .B(new_n13323_), .ZN(new_n13938_));
  NAND2_X1   g13746(.A1(new_n13936_), .A2(new_n13938_), .ZN(new_n13939_));
  NOR2_X1    g13747(.A1(new_n13404_), .A2(new_n13343_), .ZN(new_n13940_));
  NAND2_X1   g13748(.A1(\asqrt[18] ), .A2(new_n13940_), .ZN(new_n13941_));
  NAND3_X1   g13749(.A1(new_n13939_), .A2(new_n13415_), .A3(new_n13941_), .ZN(new_n13942_));
  AOI21_X1   g13750(.A1(new_n13935_), .A2(new_n13924_), .B(new_n13942_), .ZN(new_n13943_));
  NOR3_X1    g13751(.A1(new_n13932_), .A2(new_n13921_), .A3(\asqrt[61] ), .ZN(new_n13944_));
  OAI21_X1   g13752(.A1(new_n13918_), .A2(new_n13944_), .B(new_n13933_), .ZN(new_n13945_));
  AOI21_X1   g13753(.A1(new_n13945_), .A2(\asqrt[62] ), .B(new_n13939_), .ZN(new_n13946_));
  OAI21_X1   g13754(.A1(new_n13353_), .A2(new_n13343_), .B(new_n13404_), .ZN(new_n13947_));
  NOR2_X1    g13755(.A1(new_n13940_), .A2(new_n193_), .ZN(new_n13948_));
  NAND2_X1   g13756(.A1(new_n13947_), .A2(new_n13948_), .ZN(new_n13949_));
  INV_X1     g13757(.I(new_n13949_), .ZN(new_n13950_));
  AND3_X2    g13758(.A1(new_n13334_), .A2(new_n13332_), .A3(new_n13349_), .Z(new_n13951_));
  NAND4_X1   g13759(.A1(new_n13405_), .A2(new_n13415_), .A3(new_n13346_), .A4(new_n13951_), .ZN(new_n13952_));
  INV_X1     g13760(.I(new_n13952_), .ZN(new_n13953_));
  NOR2_X1    g13761(.A1(new_n13950_), .A2(new_n13953_), .ZN(new_n13954_));
  INV_X1     g13762(.I(new_n13954_), .ZN(new_n13955_));
  AOI21_X1   g13763(.A1(new_n13946_), .A2(new_n13935_), .B(new_n13955_), .ZN(new_n13956_));
  OAI21_X1   g13764(.A1(\asqrt[63] ), .A2(new_n13943_), .B(new_n13956_), .ZN(\asqrt[17] ));
  NOR2_X1    g13765(.A1(\a[32] ), .A2(\a[33] ), .ZN(new_n13958_));
  INV_X1     g13766(.I(new_n13958_), .ZN(new_n13959_));
  NOR2_X1    g13767(.A1(new_n13959_), .A2(\a[34] ), .ZN(new_n13960_));
  INV_X1     g13768(.I(new_n13960_), .ZN(new_n13961_));
  NAND2_X1   g13769(.A1(new_n13935_), .A2(new_n13924_), .ZN(new_n13962_));
  INV_X1     g13770(.I(new_n13942_), .ZN(new_n13963_));
  AOI21_X1   g13771(.A1(new_n13962_), .A2(new_n13963_), .B(\asqrt[63] ), .ZN(new_n13964_));
  INV_X1     g13772(.I(new_n13918_), .ZN(new_n13965_));
  NAND3_X1   g13773(.A1(new_n13890_), .A2(new_n327_), .A3(new_n13784_), .ZN(new_n13966_));
  AOI22_X1   g13774(.A1(new_n13966_), .A2(new_n13919_), .B1(new_n13930_), .B2(\asqrt[59] ), .ZN(new_n13967_));
  OAI21_X1   g13775(.A1(new_n13967_), .A2(new_n306_), .B(new_n218_), .ZN(new_n13968_));
  OAI21_X1   g13776(.A1(new_n13968_), .A2(new_n13932_), .B(new_n13965_), .ZN(new_n13969_));
  NOR2_X1    g13777(.A1(new_n13913_), .A2(\asqrt[62] ), .ZN(new_n13970_));
  AOI21_X1   g13778(.A1(new_n13970_), .A2(new_n13969_), .B(new_n13928_), .ZN(new_n13971_));
  INV_X1     g13779(.I(new_n13939_), .ZN(new_n13972_));
  NAND2_X1   g13780(.A1(new_n13924_), .A2(new_n13972_), .ZN(new_n13973_));
  OAI21_X1   g13781(.A1(new_n13973_), .A2(new_n13971_), .B(new_n13954_), .ZN(new_n13974_));
  OAI21_X1   g13782(.A1(new_n13964_), .A2(new_n13974_), .B(\a[34] ), .ZN(new_n13975_));
  AOI21_X1   g13783(.A1(new_n13975_), .A2(new_n13961_), .B(new_n13353_), .ZN(new_n13976_));
  INV_X1     g13784(.I(\a[34] ), .ZN(new_n13977_));
  NAND3_X1   g13785(.A1(new_n13969_), .A2(new_n207_), .A3(new_n13933_), .ZN(new_n13978_));
  AOI22_X1   g13786(.A1(new_n13978_), .A2(new_n13929_), .B1(new_n13945_), .B2(\asqrt[62] ), .ZN(new_n13979_));
  OAI21_X1   g13787(.A1(new_n13979_), .A2(new_n13942_), .B(new_n193_), .ZN(new_n13980_));
  AOI21_X1   g13788(.A1(new_n13980_), .A2(new_n13956_), .B(new_n13977_), .ZN(new_n13981_));
  NAND4_X1   g13789(.A1(new_n13415_), .A2(new_n13346_), .A3(new_n13349_), .A4(new_n13961_), .ZN(new_n13982_));
  NOR2_X1    g13790(.A1(new_n13982_), .A2(new_n13341_), .ZN(new_n13983_));
  INV_X1     g13791(.I(new_n13983_), .ZN(new_n13984_));
  NOR2_X1    g13792(.A1(new_n13981_), .A2(new_n13984_), .ZN(new_n13985_));
  AOI21_X1   g13793(.A1(new_n13980_), .A2(new_n13956_), .B(new_n13356_), .ZN(new_n13986_));
  INV_X1     g13794(.I(\a[35] ), .ZN(new_n13987_));
  AOI21_X1   g13795(.A1(\asqrt[17] ), .A2(new_n13977_), .B(new_n13987_), .ZN(new_n13988_));
  NOR3_X1    g13796(.A1(new_n13985_), .A2(new_n13988_), .A3(new_n13986_), .ZN(new_n13989_));
  OAI21_X1   g13797(.A1(new_n13989_), .A2(new_n13976_), .B(\asqrt[19] ), .ZN(new_n13990_));
  OAI21_X1   g13798(.A1(new_n13964_), .A2(new_n13974_), .B(new_n13355_), .ZN(new_n13991_));
  NAND2_X1   g13799(.A1(new_n13946_), .A2(new_n13935_), .ZN(new_n13992_));
  NOR3_X1    g13800(.A1(new_n13950_), .A2(new_n13353_), .A3(new_n13953_), .ZN(new_n13993_));
  NAND3_X1   g13801(.A1(new_n13980_), .A2(new_n13992_), .A3(new_n13993_), .ZN(new_n13994_));
  AOI21_X1   g13802(.A1(new_n13994_), .A2(new_n13991_), .B(new_n13354_), .ZN(new_n13995_));
  NAND2_X1   g13803(.A1(new_n13992_), .A2(new_n13993_), .ZN(new_n13996_));
  NOR2_X1    g13804(.A1(new_n13996_), .A2(new_n13964_), .ZN(new_n13997_));
  NOR3_X1    g13805(.A1(new_n13997_), .A2(new_n13986_), .A3(\a[36] ), .ZN(new_n13998_));
  AOI21_X1   g13806(.A1(\asqrt[17] ), .A2(\a[34] ), .B(new_n13960_), .ZN(new_n13999_));
  OAI21_X1   g13807(.A1(new_n13999_), .A2(new_n13353_), .B(new_n12913_), .ZN(new_n14000_));
  OAI22_X1   g13808(.A1(new_n13989_), .A2(new_n14000_), .B1(new_n13995_), .B2(new_n13998_), .ZN(new_n14001_));
  AOI21_X1   g13809(.A1(new_n14001_), .A2(new_n13990_), .B(new_n12364_), .ZN(new_n14002_));
  NOR3_X1    g13810(.A1(new_n13444_), .A2(new_n13445_), .A3(new_n13410_), .ZN(new_n14003_));
  NAND3_X1   g13811(.A1(\asqrt[17] ), .A2(new_n13443_), .A3(new_n13363_), .ZN(new_n14004_));
  AOI22_X1   g13812(.A1(new_n14004_), .A2(new_n13410_), .B1(\asqrt[17] ), .B2(new_n14003_), .ZN(new_n14005_));
  OAI21_X1   g13813(.A1(new_n13981_), .A2(new_n13960_), .B(\asqrt[18] ), .ZN(new_n14006_));
  AOI21_X1   g13814(.A1(new_n13980_), .A2(new_n13956_), .B(\a[34] ), .ZN(new_n14007_));
  OAI21_X1   g13815(.A1(new_n13987_), .A2(new_n14007_), .B(new_n13991_), .ZN(new_n14008_));
  OAI21_X1   g13816(.A1(new_n14008_), .A2(new_n13985_), .B(new_n14006_), .ZN(new_n14009_));
  AOI21_X1   g13817(.A1(new_n14009_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n14010_));
  AOI21_X1   g13818(.A1(new_n14010_), .A2(new_n14001_), .B(new_n14005_), .ZN(new_n14011_));
  OAI21_X1   g13819(.A1(new_n14011_), .A2(new_n14002_), .B(\asqrt[21] ), .ZN(new_n14012_));
  INV_X1     g13820(.I(new_n14012_), .ZN(new_n14013_));
  NOR2_X1    g13821(.A1(new_n13448_), .A2(new_n13451_), .ZN(new_n14014_));
  INV_X1     g13822(.I(new_n14014_), .ZN(new_n14015_));
  NAND4_X1   g13823(.A1(\asqrt[17] ), .A2(new_n13449_), .A3(new_n13423_), .A4(new_n14015_), .ZN(new_n14016_));
  INV_X1     g13824(.I(\asqrt[17] ), .ZN(new_n14017_));
  NOR3_X1    g13825(.A1(new_n14017_), .A2(new_n13412_), .A3(new_n14014_), .ZN(new_n14018_));
  OAI21_X1   g13826(.A1(new_n14018_), .A2(new_n13423_), .B(new_n14016_), .ZN(new_n14019_));
  INV_X1     g13827(.I(new_n14019_), .ZN(new_n14020_));
  NOR3_X1    g13828(.A1(new_n14011_), .A2(new_n14002_), .A3(\asqrt[21] ), .ZN(new_n14021_));
  NOR2_X1    g13829(.A1(new_n14021_), .A2(new_n14020_), .ZN(new_n14022_));
  OAI21_X1   g13830(.A1(new_n14022_), .A2(new_n14013_), .B(\asqrt[22] ), .ZN(new_n14023_));
  NAND2_X1   g13831(.A1(new_n13457_), .A2(new_n13452_), .ZN(new_n14024_));
  NAND3_X1   g13832(.A1(\asqrt[17] ), .A2(new_n13426_), .A3(new_n14024_), .ZN(new_n14025_));
  AND3_X2    g13833(.A1(new_n13426_), .A2(new_n13430_), .A3(new_n14024_), .Z(new_n14026_));
  AOI22_X1   g13834(.A1(new_n14025_), .A2(new_n13431_), .B1(\asqrt[17] ), .B2(new_n14026_), .ZN(new_n14027_));
  INV_X1     g13835(.I(new_n14027_), .ZN(new_n14028_));
  NAND2_X1   g13836(.A1(new_n14012_), .A2(new_n11326_), .ZN(new_n14029_));
  OAI21_X1   g13837(.A1(new_n14022_), .A2(new_n14029_), .B(new_n14028_), .ZN(new_n14030_));
  AOI21_X1   g13838(.A1(new_n14030_), .A2(new_n14023_), .B(new_n10812_), .ZN(new_n14031_));
  NOR3_X1    g13839(.A1(new_n13434_), .A2(new_n13440_), .A3(new_n13459_), .ZN(new_n14032_));
  NOR3_X1    g13840(.A1(new_n14017_), .A2(new_n13434_), .A3(new_n13459_), .ZN(new_n14033_));
  INV_X1     g13841(.I(new_n14033_), .ZN(new_n14034_));
  AOI22_X1   g13842(.A1(new_n14034_), .A2(new_n13440_), .B1(\asqrt[17] ), .B2(new_n14032_), .ZN(new_n14035_));
  OAI21_X1   g13843(.A1(new_n14020_), .A2(new_n14021_), .B(new_n14012_), .ZN(new_n14036_));
  AOI21_X1   g13844(.A1(new_n14036_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n14037_));
  AOI21_X1   g13845(.A1(new_n14037_), .A2(new_n14030_), .B(new_n14035_), .ZN(new_n14038_));
  OAI21_X1   g13846(.A1(new_n14038_), .A2(new_n14031_), .B(\asqrt[24] ), .ZN(new_n14039_));
  INV_X1     g13847(.I(new_n14039_), .ZN(new_n14040_));
  NAND2_X1   g13848(.A1(new_n13805_), .A2(new_n13803_), .ZN(new_n14041_));
  NAND3_X1   g13849(.A1(\asqrt[17] ), .A2(new_n13461_), .A3(new_n14041_), .ZN(new_n14042_));
  AND3_X2    g13850(.A1(new_n14041_), .A2(new_n13461_), .A3(new_n13466_), .Z(new_n14043_));
  AOI22_X1   g13851(.A1(new_n14042_), .A2(new_n13467_), .B1(\asqrt[17] ), .B2(new_n14043_), .ZN(new_n14044_));
  NOR3_X1    g13852(.A1(new_n14038_), .A2(new_n14031_), .A3(\asqrt[24] ), .ZN(new_n14045_));
  NOR2_X1    g13853(.A1(new_n14045_), .A2(new_n14044_), .ZN(new_n14046_));
  OAI21_X1   g13854(.A1(new_n14046_), .A2(new_n14040_), .B(\asqrt[25] ), .ZN(new_n14047_));
  INV_X1     g13855(.I(new_n13475_), .ZN(new_n14048_));
  NOR3_X1    g13856(.A1(new_n13816_), .A2(new_n13471_), .A3(new_n14048_), .ZN(new_n14049_));
  NOR3_X1    g13857(.A1(new_n14017_), .A2(new_n13471_), .A3(new_n13816_), .ZN(new_n14050_));
  INV_X1     g13858(.I(new_n14050_), .ZN(new_n14051_));
  AOI22_X1   g13859(.A1(new_n14051_), .A2(new_n14048_), .B1(\asqrt[17] ), .B2(new_n14049_), .ZN(new_n14052_));
  INV_X1     g13860(.I(new_n14052_), .ZN(new_n14053_));
  NAND2_X1   g13861(.A1(new_n14039_), .A2(new_n9846_), .ZN(new_n14054_));
  OAI21_X1   g13862(.A1(new_n14046_), .A2(new_n14054_), .B(new_n14053_), .ZN(new_n14055_));
  AOI21_X1   g13863(.A1(new_n14055_), .A2(new_n14047_), .B(new_n9317_), .ZN(new_n14056_));
  NOR3_X1    g13864(.A1(new_n14017_), .A2(new_n13480_), .A3(new_n13485_), .ZN(new_n14057_));
  INV_X1     g13865(.I(new_n14057_), .ZN(new_n14058_));
  NOR3_X1    g13866(.A1(new_n13480_), .A2(new_n13801_), .A3(new_n13485_), .ZN(new_n14059_));
  AOI22_X1   g13867(.A1(new_n14058_), .A2(new_n13801_), .B1(\asqrt[17] ), .B2(new_n14059_), .ZN(new_n14060_));
  OAI21_X1   g13868(.A1(new_n14044_), .A2(new_n14045_), .B(new_n14039_), .ZN(new_n14061_));
  AOI21_X1   g13869(.A1(new_n14061_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n14062_));
  AOI21_X1   g13870(.A1(new_n14062_), .A2(new_n14055_), .B(new_n14060_), .ZN(new_n14063_));
  OAI21_X1   g13871(.A1(new_n14063_), .A2(new_n14056_), .B(\asqrt[27] ), .ZN(new_n14064_));
  INV_X1     g13872(.I(new_n14064_), .ZN(new_n14065_));
  INV_X1     g13873(.I(new_n13810_), .ZN(new_n14066_));
  NOR3_X1    g13874(.A1(new_n14066_), .A2(new_n13815_), .A3(new_n13493_), .ZN(new_n14067_));
  NOR3_X1    g13875(.A1(new_n14017_), .A2(new_n13815_), .A3(new_n14066_), .ZN(new_n14068_));
  INV_X1     g13876(.I(new_n14068_), .ZN(new_n14069_));
  AOI22_X1   g13877(.A1(new_n14069_), .A2(new_n13493_), .B1(\asqrt[17] ), .B2(new_n14067_), .ZN(new_n14070_));
  NOR3_X1    g13878(.A1(new_n14063_), .A2(new_n14056_), .A3(\asqrt[27] ), .ZN(new_n14071_));
  NOR2_X1    g13879(.A1(new_n14071_), .A2(new_n14070_), .ZN(new_n14072_));
  OAI21_X1   g13880(.A1(new_n14072_), .A2(new_n14065_), .B(\asqrt[28] ), .ZN(new_n14073_));
  INV_X1     g13881(.I(new_n13500_), .ZN(new_n14074_));
  NOR3_X1    g13882(.A1(new_n14017_), .A2(new_n13496_), .A3(new_n13820_), .ZN(new_n14075_));
  INV_X1     g13883(.I(new_n14075_), .ZN(new_n14076_));
  NOR3_X1    g13884(.A1(new_n13820_), .A2(new_n13496_), .A3(new_n14074_), .ZN(new_n14077_));
  AOI22_X1   g13885(.A1(new_n14076_), .A2(new_n14074_), .B1(\asqrt[17] ), .B2(new_n14077_), .ZN(new_n14078_));
  INV_X1     g13886(.I(new_n14078_), .ZN(new_n14079_));
  NAND2_X1   g13887(.A1(new_n14064_), .A2(new_n8483_), .ZN(new_n14080_));
  OAI21_X1   g13888(.A1(new_n14072_), .A2(new_n14080_), .B(new_n14079_), .ZN(new_n14081_));
  AOI21_X1   g13889(.A1(new_n14081_), .A2(new_n14073_), .B(new_n8036_), .ZN(new_n14082_));
  NOR3_X1    g13890(.A1(new_n13505_), .A2(new_n13800_), .A3(new_n13511_), .ZN(new_n14083_));
  NOR3_X1    g13891(.A1(new_n14017_), .A2(new_n13505_), .A3(new_n13511_), .ZN(new_n14084_));
  INV_X1     g13892(.I(new_n14084_), .ZN(new_n14085_));
  AOI22_X1   g13893(.A1(new_n14085_), .A2(new_n13800_), .B1(\asqrt[17] ), .B2(new_n14083_), .ZN(new_n14086_));
  OAI21_X1   g13894(.A1(new_n14070_), .A2(new_n14071_), .B(new_n14064_), .ZN(new_n14087_));
  AOI21_X1   g13895(.A1(new_n14087_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n14088_));
  AOI21_X1   g13896(.A1(new_n14088_), .A2(new_n14081_), .B(new_n14086_), .ZN(new_n14089_));
  OAI21_X1   g13897(.A1(new_n14089_), .A2(new_n14082_), .B(\asqrt[30] ), .ZN(new_n14090_));
  INV_X1     g13898(.I(new_n14090_), .ZN(new_n14091_));
  NOR2_X1    g13899(.A1(new_n13512_), .A2(new_n13520_), .ZN(new_n14092_));
  NOR3_X1    g13900(.A1(new_n14017_), .A2(new_n13814_), .A3(new_n14092_), .ZN(new_n14093_));
  INV_X1     g13901(.I(new_n14093_), .ZN(new_n14094_));
  NOR3_X1    g13902(.A1(new_n14092_), .A2(new_n13814_), .A3(new_n13519_), .ZN(new_n14095_));
  AOI22_X1   g13903(.A1(new_n14094_), .A2(new_n13519_), .B1(\asqrt[17] ), .B2(new_n14095_), .ZN(new_n14096_));
  NOR3_X1    g13904(.A1(new_n14089_), .A2(new_n14082_), .A3(\asqrt[30] ), .ZN(new_n14097_));
  NOR2_X1    g13905(.A1(new_n14097_), .A2(new_n14096_), .ZN(new_n14098_));
  OAI21_X1   g13906(.A1(new_n14098_), .A2(new_n14091_), .B(\asqrt[31] ), .ZN(new_n14099_));
  INV_X1     g13907(.I(new_n13528_), .ZN(new_n14100_));
  NOR3_X1    g13908(.A1(new_n13828_), .A2(new_n13522_), .A3(new_n14100_), .ZN(new_n14101_));
  NOR3_X1    g13909(.A1(new_n14017_), .A2(new_n13522_), .A3(new_n13828_), .ZN(new_n14102_));
  INV_X1     g13910(.I(new_n14102_), .ZN(new_n14103_));
  AOI22_X1   g13911(.A1(new_n14103_), .A2(new_n14100_), .B1(\asqrt[17] ), .B2(new_n14101_), .ZN(new_n14104_));
  INV_X1     g13912(.I(new_n14104_), .ZN(new_n14105_));
  NAND2_X1   g13913(.A1(new_n14090_), .A2(new_n7229_), .ZN(new_n14106_));
  OAI21_X1   g13914(.A1(new_n14098_), .A2(new_n14106_), .B(new_n14105_), .ZN(new_n14107_));
  AOI21_X1   g13915(.A1(new_n14107_), .A2(new_n14099_), .B(new_n6824_), .ZN(new_n14108_));
  NOR3_X1    g13916(.A1(new_n14017_), .A2(new_n13533_), .A3(new_n13539_), .ZN(new_n14109_));
  INV_X1     g13917(.I(new_n14109_), .ZN(new_n14110_));
  NOR3_X1    g13918(.A1(new_n13533_), .A2(new_n13799_), .A3(new_n13539_), .ZN(new_n14111_));
  AOI22_X1   g13919(.A1(new_n14110_), .A2(new_n13799_), .B1(\asqrt[17] ), .B2(new_n14111_), .ZN(new_n14112_));
  OAI21_X1   g13920(.A1(new_n14096_), .A2(new_n14097_), .B(new_n14090_), .ZN(new_n14113_));
  AOI21_X1   g13921(.A1(new_n14113_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n14114_));
  AOI21_X1   g13922(.A1(new_n14114_), .A2(new_n14107_), .B(new_n14112_), .ZN(new_n14115_));
  OAI21_X1   g13923(.A1(new_n14115_), .A2(new_n14108_), .B(\asqrt[33] ), .ZN(new_n14116_));
  INV_X1     g13924(.I(new_n14116_), .ZN(new_n14117_));
  NOR2_X1    g13925(.A1(new_n13540_), .A2(new_n13548_), .ZN(new_n14118_));
  NOR3_X1    g13926(.A1(new_n14118_), .A2(new_n13827_), .A3(new_n13547_), .ZN(new_n14119_));
  NOR3_X1    g13927(.A1(new_n14017_), .A2(new_n13827_), .A3(new_n14118_), .ZN(new_n14120_));
  INV_X1     g13928(.I(new_n14120_), .ZN(new_n14121_));
  AOI22_X1   g13929(.A1(new_n14121_), .A2(new_n13547_), .B1(\asqrt[17] ), .B2(new_n14119_), .ZN(new_n14122_));
  NOR3_X1    g13930(.A1(new_n14115_), .A2(new_n14108_), .A3(\asqrt[33] ), .ZN(new_n14123_));
  NOR2_X1    g13931(.A1(new_n14123_), .A2(new_n14122_), .ZN(new_n14124_));
  OAI21_X1   g13932(.A1(new_n14124_), .A2(new_n14117_), .B(\asqrt[34] ), .ZN(new_n14125_));
  INV_X1     g13933(.I(new_n13555_), .ZN(new_n14126_));
  NOR3_X1    g13934(.A1(new_n14017_), .A2(new_n13550_), .A3(new_n13836_), .ZN(new_n14127_));
  INV_X1     g13935(.I(new_n14127_), .ZN(new_n14128_));
  NOR3_X1    g13936(.A1(new_n13836_), .A2(new_n13550_), .A3(new_n14126_), .ZN(new_n14129_));
  AOI22_X1   g13937(.A1(new_n14128_), .A2(new_n14126_), .B1(\asqrt[17] ), .B2(new_n14129_), .ZN(new_n14130_));
  INV_X1     g13938(.I(new_n14130_), .ZN(new_n14131_));
  NAND2_X1   g13939(.A1(new_n14116_), .A2(new_n6077_), .ZN(new_n14132_));
  OAI21_X1   g13940(.A1(new_n14124_), .A2(new_n14132_), .B(new_n14131_), .ZN(new_n14133_));
  AOI21_X1   g13941(.A1(new_n14133_), .A2(new_n14125_), .B(new_n5708_), .ZN(new_n14134_));
  NOR3_X1    g13942(.A1(new_n13560_), .A2(new_n13798_), .A3(new_n13566_), .ZN(new_n14135_));
  NOR3_X1    g13943(.A1(new_n14017_), .A2(new_n13560_), .A3(new_n13566_), .ZN(new_n14136_));
  INV_X1     g13944(.I(new_n14136_), .ZN(new_n14137_));
  AOI22_X1   g13945(.A1(new_n14137_), .A2(new_n13798_), .B1(\asqrt[17] ), .B2(new_n14135_), .ZN(new_n14138_));
  OAI21_X1   g13946(.A1(new_n14122_), .A2(new_n14123_), .B(new_n14116_), .ZN(new_n14139_));
  AOI21_X1   g13947(.A1(new_n14139_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n14140_));
  AOI21_X1   g13948(.A1(new_n14140_), .A2(new_n14133_), .B(new_n14138_), .ZN(new_n14141_));
  OAI21_X1   g13949(.A1(new_n14141_), .A2(new_n14134_), .B(\asqrt[36] ), .ZN(new_n14142_));
  INV_X1     g13950(.I(new_n14142_), .ZN(new_n14143_));
  NOR2_X1    g13951(.A1(new_n13567_), .A2(new_n13575_), .ZN(new_n14144_));
  NOR3_X1    g13952(.A1(new_n14017_), .A2(new_n13835_), .A3(new_n14144_), .ZN(new_n14145_));
  INV_X1     g13953(.I(new_n14145_), .ZN(new_n14146_));
  NOR3_X1    g13954(.A1(new_n14144_), .A2(new_n13835_), .A3(new_n13574_), .ZN(new_n14147_));
  AOI22_X1   g13955(.A1(new_n14146_), .A2(new_n13574_), .B1(\asqrt[17] ), .B2(new_n14147_), .ZN(new_n14148_));
  NOR3_X1    g13956(.A1(new_n14141_), .A2(new_n14134_), .A3(\asqrt[36] ), .ZN(new_n14149_));
  NOR2_X1    g13957(.A1(new_n14149_), .A2(new_n14148_), .ZN(new_n14150_));
  OAI21_X1   g13958(.A1(new_n14150_), .A2(new_n14143_), .B(\asqrt[37] ), .ZN(new_n14151_));
  INV_X1     g13959(.I(new_n13582_), .ZN(new_n14152_));
  NOR3_X1    g13960(.A1(new_n13844_), .A2(new_n13577_), .A3(new_n14152_), .ZN(new_n14153_));
  NOR3_X1    g13961(.A1(new_n14017_), .A2(new_n13577_), .A3(new_n13844_), .ZN(new_n14154_));
  INV_X1     g13962(.I(new_n14154_), .ZN(new_n14155_));
  AOI22_X1   g13963(.A1(new_n14155_), .A2(new_n14152_), .B1(\asqrt[17] ), .B2(new_n14153_), .ZN(new_n14156_));
  INV_X1     g13964(.I(new_n14156_), .ZN(new_n14157_));
  NAND2_X1   g13965(.A1(new_n14142_), .A2(new_n5024_), .ZN(new_n14158_));
  OAI21_X1   g13966(.A1(new_n14150_), .A2(new_n14158_), .B(new_n14157_), .ZN(new_n14159_));
  AOI21_X1   g13967(.A1(new_n14159_), .A2(new_n14151_), .B(new_n4696_), .ZN(new_n14160_));
  NOR3_X1    g13968(.A1(new_n14017_), .A2(new_n13587_), .A3(new_n13593_), .ZN(new_n14161_));
  INV_X1     g13969(.I(new_n14161_), .ZN(new_n14162_));
  NOR3_X1    g13970(.A1(new_n13587_), .A2(new_n13797_), .A3(new_n13593_), .ZN(new_n14163_));
  AOI22_X1   g13971(.A1(new_n14162_), .A2(new_n13797_), .B1(\asqrt[17] ), .B2(new_n14163_), .ZN(new_n14164_));
  OAI21_X1   g13972(.A1(new_n14148_), .A2(new_n14149_), .B(new_n14142_), .ZN(new_n14165_));
  AOI21_X1   g13973(.A1(new_n14165_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n14166_));
  AOI21_X1   g13974(.A1(new_n14166_), .A2(new_n14159_), .B(new_n14164_), .ZN(new_n14167_));
  OAI21_X1   g13975(.A1(new_n14167_), .A2(new_n14160_), .B(\asqrt[39] ), .ZN(new_n14168_));
  INV_X1     g13976(.I(new_n14168_), .ZN(new_n14169_));
  NOR2_X1    g13977(.A1(new_n13594_), .A2(new_n13602_), .ZN(new_n14170_));
  NOR3_X1    g13978(.A1(new_n14170_), .A2(new_n13843_), .A3(new_n13601_), .ZN(new_n14171_));
  NOR3_X1    g13979(.A1(new_n14017_), .A2(new_n13843_), .A3(new_n14170_), .ZN(new_n14172_));
  INV_X1     g13980(.I(new_n14172_), .ZN(new_n14173_));
  AOI22_X1   g13981(.A1(new_n14173_), .A2(new_n13601_), .B1(\asqrt[17] ), .B2(new_n14171_), .ZN(new_n14174_));
  NOR3_X1    g13982(.A1(new_n14167_), .A2(new_n14160_), .A3(\asqrt[39] ), .ZN(new_n14175_));
  NOR2_X1    g13983(.A1(new_n14175_), .A2(new_n14174_), .ZN(new_n14176_));
  OAI21_X1   g13984(.A1(new_n14176_), .A2(new_n14169_), .B(\asqrt[40] ), .ZN(new_n14177_));
  INV_X1     g13985(.I(new_n13608_), .ZN(new_n14178_));
  NOR3_X1    g13986(.A1(new_n14017_), .A2(new_n13604_), .A3(new_n13852_), .ZN(new_n14179_));
  INV_X1     g13987(.I(new_n14179_), .ZN(new_n14180_));
  NOR3_X1    g13988(.A1(new_n13852_), .A2(new_n13604_), .A3(new_n14178_), .ZN(new_n14181_));
  AOI22_X1   g13989(.A1(new_n14180_), .A2(new_n14178_), .B1(\asqrt[17] ), .B2(new_n14181_), .ZN(new_n14182_));
  INV_X1     g13990(.I(new_n14182_), .ZN(new_n14183_));
  NAND2_X1   g13991(.A1(new_n14168_), .A2(new_n4071_), .ZN(new_n14184_));
  OAI21_X1   g13992(.A1(new_n14176_), .A2(new_n14184_), .B(new_n14183_), .ZN(new_n14185_));
  AOI21_X1   g13993(.A1(new_n14185_), .A2(new_n14177_), .B(new_n3782_), .ZN(new_n14186_));
  NOR3_X1    g13994(.A1(new_n13613_), .A2(new_n13796_), .A3(new_n13619_), .ZN(new_n14187_));
  NOR3_X1    g13995(.A1(new_n14017_), .A2(new_n13613_), .A3(new_n13619_), .ZN(new_n14188_));
  INV_X1     g13996(.I(new_n14188_), .ZN(new_n14189_));
  AOI22_X1   g13997(.A1(new_n14189_), .A2(new_n13796_), .B1(\asqrt[17] ), .B2(new_n14187_), .ZN(new_n14190_));
  OAI21_X1   g13998(.A1(new_n14174_), .A2(new_n14175_), .B(new_n14168_), .ZN(new_n14191_));
  AOI21_X1   g13999(.A1(new_n14191_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n14192_));
  AOI21_X1   g14000(.A1(new_n14192_), .A2(new_n14185_), .B(new_n14190_), .ZN(new_n14193_));
  OAI21_X1   g14001(.A1(new_n14193_), .A2(new_n14186_), .B(\asqrt[42] ), .ZN(new_n14194_));
  INV_X1     g14002(.I(new_n14194_), .ZN(new_n14195_));
  NOR2_X1    g14003(.A1(new_n13620_), .A2(new_n13628_), .ZN(new_n14196_));
  NOR3_X1    g14004(.A1(new_n14017_), .A2(new_n13851_), .A3(new_n14196_), .ZN(new_n14197_));
  INV_X1     g14005(.I(new_n14197_), .ZN(new_n14198_));
  NOR3_X1    g14006(.A1(new_n14196_), .A2(new_n13851_), .A3(new_n13627_), .ZN(new_n14199_));
  AOI22_X1   g14007(.A1(new_n14198_), .A2(new_n13627_), .B1(\asqrt[17] ), .B2(new_n14199_), .ZN(new_n14200_));
  NOR3_X1    g14008(.A1(new_n14193_), .A2(new_n14186_), .A3(\asqrt[42] ), .ZN(new_n14201_));
  NOR2_X1    g14009(.A1(new_n14201_), .A2(new_n14200_), .ZN(new_n14202_));
  OAI21_X1   g14010(.A1(new_n14202_), .A2(new_n14195_), .B(\asqrt[43] ), .ZN(new_n14203_));
  INV_X1     g14011(.I(new_n13634_), .ZN(new_n14204_));
  NOR3_X1    g14012(.A1(new_n13860_), .A2(new_n13630_), .A3(new_n14204_), .ZN(new_n14205_));
  NOR3_X1    g14013(.A1(new_n14017_), .A2(new_n13630_), .A3(new_n13860_), .ZN(new_n14206_));
  INV_X1     g14014(.I(new_n14206_), .ZN(new_n14207_));
  AOI22_X1   g14015(.A1(new_n14207_), .A2(new_n14204_), .B1(\asqrt[17] ), .B2(new_n14205_), .ZN(new_n14208_));
  INV_X1     g14016(.I(new_n14208_), .ZN(new_n14209_));
  NAND2_X1   g14017(.A1(new_n14194_), .A2(new_n3218_), .ZN(new_n14210_));
  OAI21_X1   g14018(.A1(new_n14202_), .A2(new_n14210_), .B(new_n14209_), .ZN(new_n14211_));
  AOI21_X1   g14019(.A1(new_n14211_), .A2(new_n14203_), .B(new_n2954_), .ZN(new_n14212_));
  NOR3_X1    g14020(.A1(new_n14017_), .A2(new_n13639_), .A3(new_n13647_), .ZN(new_n14213_));
  INV_X1     g14021(.I(new_n14213_), .ZN(new_n14214_));
  NOR3_X1    g14022(.A1(new_n13639_), .A2(new_n13795_), .A3(new_n13647_), .ZN(new_n14215_));
  AOI22_X1   g14023(.A1(new_n14214_), .A2(new_n13795_), .B1(\asqrt[17] ), .B2(new_n14215_), .ZN(new_n14216_));
  OAI21_X1   g14024(.A1(new_n14200_), .A2(new_n14201_), .B(new_n14194_), .ZN(new_n14217_));
  AOI21_X1   g14025(.A1(new_n14217_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n14218_));
  AOI21_X1   g14026(.A1(new_n14218_), .A2(new_n14211_), .B(new_n14216_), .ZN(new_n14219_));
  OAI21_X1   g14027(.A1(new_n14219_), .A2(new_n14212_), .B(\asqrt[45] ), .ZN(new_n14220_));
  INV_X1     g14028(.I(new_n14220_), .ZN(new_n14221_));
  NOR2_X1    g14029(.A1(new_n13648_), .A2(new_n13655_), .ZN(new_n14222_));
  NOR3_X1    g14030(.A1(new_n14222_), .A2(new_n13859_), .A3(new_n13654_), .ZN(new_n14223_));
  NOR3_X1    g14031(.A1(new_n14017_), .A2(new_n13859_), .A3(new_n14222_), .ZN(new_n14224_));
  INV_X1     g14032(.I(new_n14224_), .ZN(new_n14225_));
  AOI22_X1   g14033(.A1(new_n14225_), .A2(new_n13654_), .B1(\asqrt[17] ), .B2(new_n14223_), .ZN(new_n14226_));
  NOR3_X1    g14034(.A1(new_n14219_), .A2(new_n14212_), .A3(\asqrt[45] ), .ZN(new_n14227_));
  NOR2_X1    g14035(.A1(new_n14227_), .A2(new_n14226_), .ZN(new_n14228_));
  OAI21_X1   g14036(.A1(new_n14228_), .A2(new_n14221_), .B(\asqrt[46] ), .ZN(new_n14229_));
  INV_X1     g14037(.I(new_n13663_), .ZN(new_n14230_));
  NOR3_X1    g14038(.A1(new_n14017_), .A2(new_n13657_), .A3(new_n13868_), .ZN(new_n14231_));
  INV_X1     g14039(.I(new_n14231_), .ZN(new_n14232_));
  NOR3_X1    g14040(.A1(new_n13868_), .A2(new_n13657_), .A3(new_n14230_), .ZN(new_n14233_));
  AOI22_X1   g14041(.A1(new_n14232_), .A2(new_n14230_), .B1(\asqrt[17] ), .B2(new_n14233_), .ZN(new_n14234_));
  INV_X1     g14042(.I(new_n14234_), .ZN(new_n14235_));
  NAND2_X1   g14043(.A1(new_n14220_), .A2(new_n2465_), .ZN(new_n14236_));
  OAI21_X1   g14044(.A1(new_n14228_), .A2(new_n14236_), .B(new_n14235_), .ZN(new_n14237_));
  AOI21_X1   g14045(.A1(new_n14237_), .A2(new_n14229_), .B(new_n2229_), .ZN(new_n14238_));
  NOR3_X1    g14046(.A1(new_n13668_), .A2(new_n13794_), .A3(new_n13677_), .ZN(new_n14239_));
  NOR3_X1    g14047(.A1(new_n14017_), .A2(new_n13668_), .A3(new_n13677_), .ZN(new_n14240_));
  INV_X1     g14048(.I(new_n14240_), .ZN(new_n14241_));
  AOI22_X1   g14049(.A1(new_n14241_), .A2(new_n13794_), .B1(\asqrt[17] ), .B2(new_n14239_), .ZN(new_n14242_));
  OAI21_X1   g14050(.A1(new_n14226_), .A2(new_n14227_), .B(new_n14220_), .ZN(new_n14243_));
  AOI21_X1   g14051(.A1(new_n14243_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n14244_));
  AOI21_X1   g14052(.A1(new_n14244_), .A2(new_n14237_), .B(new_n14242_), .ZN(new_n14245_));
  OAI21_X1   g14053(.A1(new_n14245_), .A2(new_n14238_), .B(\asqrt[48] ), .ZN(new_n14246_));
  INV_X1     g14054(.I(new_n14246_), .ZN(new_n14247_));
  NOR2_X1    g14055(.A1(new_n13678_), .A2(new_n13685_), .ZN(new_n14248_));
  NOR3_X1    g14056(.A1(new_n14017_), .A2(new_n13867_), .A3(new_n14248_), .ZN(new_n14249_));
  INV_X1     g14057(.I(new_n14249_), .ZN(new_n14250_));
  NOR3_X1    g14058(.A1(new_n14248_), .A2(new_n13867_), .A3(new_n13684_), .ZN(new_n14251_));
  AOI22_X1   g14059(.A1(new_n14250_), .A2(new_n13684_), .B1(\asqrt[17] ), .B2(new_n14251_), .ZN(new_n14252_));
  NOR3_X1    g14060(.A1(new_n14245_), .A2(new_n14238_), .A3(\asqrt[48] ), .ZN(new_n14253_));
  NOR2_X1    g14061(.A1(new_n14253_), .A2(new_n14252_), .ZN(new_n14254_));
  OAI21_X1   g14062(.A1(new_n14254_), .A2(new_n14247_), .B(\asqrt[49] ), .ZN(new_n14255_));
  INV_X1     g14063(.I(new_n13693_), .ZN(new_n14256_));
  NOR3_X1    g14064(.A1(new_n13876_), .A2(new_n13687_), .A3(new_n14256_), .ZN(new_n14257_));
  NOR3_X1    g14065(.A1(new_n14017_), .A2(new_n13687_), .A3(new_n13876_), .ZN(new_n14258_));
  INV_X1     g14066(.I(new_n14258_), .ZN(new_n14259_));
  AOI22_X1   g14067(.A1(new_n14259_), .A2(new_n14256_), .B1(\asqrt[17] ), .B2(new_n14257_), .ZN(new_n14260_));
  INV_X1     g14068(.I(new_n14260_), .ZN(new_n14261_));
  NAND2_X1   g14069(.A1(new_n14246_), .A2(new_n1806_), .ZN(new_n14262_));
  OAI21_X1   g14070(.A1(new_n14254_), .A2(new_n14262_), .B(new_n14261_), .ZN(new_n14263_));
  AOI21_X1   g14071(.A1(new_n14263_), .A2(new_n14255_), .B(new_n1612_), .ZN(new_n14264_));
  NOR3_X1    g14072(.A1(new_n14017_), .A2(new_n13698_), .A3(new_n13707_), .ZN(new_n14265_));
  INV_X1     g14073(.I(new_n14265_), .ZN(new_n14266_));
  NOR3_X1    g14074(.A1(new_n13698_), .A2(new_n13793_), .A3(new_n13707_), .ZN(new_n14267_));
  AOI22_X1   g14075(.A1(new_n14266_), .A2(new_n13793_), .B1(\asqrt[17] ), .B2(new_n14267_), .ZN(new_n14268_));
  OAI21_X1   g14076(.A1(new_n14252_), .A2(new_n14253_), .B(new_n14246_), .ZN(new_n14269_));
  AOI21_X1   g14077(.A1(new_n14269_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n14270_));
  AOI21_X1   g14078(.A1(new_n14270_), .A2(new_n14263_), .B(new_n14268_), .ZN(new_n14271_));
  OAI21_X1   g14079(.A1(new_n14271_), .A2(new_n14264_), .B(\asqrt[51] ), .ZN(new_n14272_));
  INV_X1     g14080(.I(new_n14272_), .ZN(new_n14273_));
  NOR2_X1    g14081(.A1(new_n13708_), .A2(new_n13715_), .ZN(new_n14274_));
  NOR3_X1    g14082(.A1(new_n14274_), .A2(new_n13875_), .A3(new_n13714_), .ZN(new_n14275_));
  NOR3_X1    g14083(.A1(new_n14017_), .A2(new_n13875_), .A3(new_n14274_), .ZN(new_n14276_));
  INV_X1     g14084(.I(new_n14276_), .ZN(new_n14277_));
  AOI22_X1   g14085(.A1(new_n14277_), .A2(new_n13714_), .B1(\asqrt[17] ), .B2(new_n14275_), .ZN(new_n14278_));
  NOR3_X1    g14086(.A1(new_n14271_), .A2(new_n14264_), .A3(\asqrt[51] ), .ZN(new_n14279_));
  NOR2_X1    g14087(.A1(new_n14279_), .A2(new_n14278_), .ZN(new_n14280_));
  OAI21_X1   g14088(.A1(new_n14280_), .A2(new_n14273_), .B(\asqrt[52] ), .ZN(new_n14281_));
  INV_X1     g14089(.I(new_n13723_), .ZN(new_n14282_));
  NAND2_X1   g14090(.A1(new_n13725_), .A2(new_n13716_), .ZN(new_n14283_));
  INV_X1     g14091(.I(new_n14283_), .ZN(new_n14284_));
  NOR3_X1    g14092(.A1(new_n14017_), .A2(new_n13717_), .A3(new_n14284_), .ZN(new_n14285_));
  INV_X1     g14093(.I(new_n14285_), .ZN(new_n14286_));
  NOR3_X1    g14094(.A1(new_n14284_), .A2(new_n13717_), .A3(new_n14282_), .ZN(new_n14287_));
  AOI22_X1   g14095(.A1(new_n14286_), .A2(new_n14282_), .B1(\asqrt[17] ), .B2(new_n14287_), .ZN(new_n14288_));
  INV_X1     g14096(.I(new_n14288_), .ZN(new_n14289_));
  NAND2_X1   g14097(.A1(new_n14272_), .A2(new_n1256_), .ZN(new_n14290_));
  OAI21_X1   g14098(.A1(new_n14280_), .A2(new_n14290_), .B(new_n14289_), .ZN(new_n14291_));
  AOI21_X1   g14099(.A1(new_n14291_), .A2(new_n14281_), .B(new_n1103_), .ZN(new_n14292_));
  NOR3_X1    g14100(.A1(new_n13728_), .A2(new_n13792_), .A3(new_n13737_), .ZN(new_n14293_));
  NOR3_X1    g14101(.A1(new_n14017_), .A2(new_n13728_), .A3(new_n13737_), .ZN(new_n14294_));
  INV_X1     g14102(.I(new_n14294_), .ZN(new_n14295_));
  AOI22_X1   g14103(.A1(new_n14295_), .A2(new_n13792_), .B1(\asqrt[17] ), .B2(new_n14293_), .ZN(new_n14296_));
  OAI21_X1   g14104(.A1(new_n14278_), .A2(new_n14279_), .B(new_n14272_), .ZN(new_n14297_));
  AOI21_X1   g14105(.A1(new_n14297_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n14298_));
  AOI21_X1   g14106(.A1(new_n14298_), .A2(new_n14291_), .B(new_n14296_), .ZN(new_n14299_));
  OAI21_X1   g14107(.A1(new_n14299_), .A2(new_n14292_), .B(\asqrt[54] ), .ZN(new_n14300_));
  INV_X1     g14108(.I(new_n14300_), .ZN(new_n14301_));
  INV_X1     g14109(.I(new_n13739_), .ZN(new_n14302_));
  INV_X1     g14110(.I(new_n13883_), .ZN(new_n14303_));
  NOR3_X1    g14111(.A1(new_n14017_), .A2(new_n14302_), .A3(new_n14303_), .ZN(new_n14304_));
  INV_X1     g14112(.I(new_n14304_), .ZN(new_n14305_));
  NOR3_X1    g14113(.A1(new_n14302_), .A2(new_n14303_), .A3(new_n13744_), .ZN(new_n14306_));
  AOI22_X1   g14114(.A1(new_n14305_), .A2(new_n13744_), .B1(\asqrt[17] ), .B2(new_n14306_), .ZN(new_n14307_));
  NOR3_X1    g14115(.A1(new_n14299_), .A2(new_n14292_), .A3(\asqrt[54] ), .ZN(new_n14308_));
  NOR2_X1    g14116(.A1(new_n14308_), .A2(new_n14307_), .ZN(new_n14309_));
  OAI21_X1   g14117(.A1(new_n14309_), .A2(new_n14301_), .B(\asqrt[55] ), .ZN(new_n14310_));
  INV_X1     g14118(.I(new_n13753_), .ZN(new_n14311_));
  INV_X1     g14119(.I(new_n13746_), .ZN(new_n14312_));
  INV_X1     g14120(.I(new_n13755_), .ZN(new_n14313_));
  OAI21_X1   g14121(.A1(new_n14313_), .A2(new_n14312_), .B(new_n13753_), .ZN(new_n14314_));
  NOR2_X1    g14122(.A1(new_n14314_), .A2(new_n13747_), .ZN(new_n14315_));
  NOR2_X1    g14123(.A1(new_n14313_), .A2(new_n14312_), .ZN(new_n14316_));
  NOR3_X1    g14124(.A1(new_n14017_), .A2(new_n13747_), .A3(new_n14316_), .ZN(new_n14317_));
  INV_X1     g14125(.I(new_n14317_), .ZN(new_n14318_));
  AOI22_X1   g14126(.A1(new_n14318_), .A2(new_n14311_), .B1(\asqrt[17] ), .B2(new_n14315_), .ZN(new_n14319_));
  INV_X1     g14127(.I(new_n14319_), .ZN(new_n14320_));
  NAND2_X1   g14128(.A1(new_n14300_), .A2(new_n823_), .ZN(new_n14321_));
  OAI21_X1   g14129(.A1(new_n14309_), .A2(new_n14321_), .B(new_n14320_), .ZN(new_n14322_));
  AOI21_X1   g14130(.A1(new_n14322_), .A2(new_n14310_), .B(new_n703_), .ZN(new_n14323_));
  NOR3_X1    g14131(.A1(new_n14017_), .A2(new_n13758_), .A3(new_n13764_), .ZN(new_n14324_));
  INV_X1     g14132(.I(new_n14324_), .ZN(new_n14325_));
  NOR3_X1    g14133(.A1(new_n13758_), .A2(new_n13791_), .A3(new_n13764_), .ZN(new_n14326_));
  AOI22_X1   g14134(.A1(new_n14325_), .A2(new_n13791_), .B1(\asqrt[17] ), .B2(new_n14326_), .ZN(new_n14327_));
  OAI21_X1   g14135(.A1(new_n14307_), .A2(new_n14308_), .B(new_n14300_), .ZN(new_n14328_));
  AOI21_X1   g14136(.A1(new_n14328_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n14329_));
  AOI21_X1   g14137(.A1(new_n14329_), .A2(new_n14322_), .B(new_n14327_), .ZN(new_n14330_));
  OAI21_X1   g14138(.A1(new_n14330_), .A2(new_n14323_), .B(\asqrt[57] ), .ZN(new_n14331_));
  INV_X1     g14139(.I(new_n14331_), .ZN(new_n14332_));
  INV_X1     g14140(.I(new_n13766_), .ZN(new_n14333_));
  INV_X1     g14141(.I(new_n13887_), .ZN(new_n14334_));
  NOR3_X1    g14142(.A1(new_n14333_), .A2(new_n14334_), .A3(new_n13771_), .ZN(new_n14335_));
  NOR3_X1    g14143(.A1(new_n14017_), .A2(new_n14333_), .A3(new_n14334_), .ZN(new_n14336_));
  INV_X1     g14144(.I(new_n14336_), .ZN(new_n14337_));
  AOI22_X1   g14145(.A1(new_n14337_), .A2(new_n13771_), .B1(\asqrt[17] ), .B2(new_n14335_), .ZN(new_n14338_));
  NOR3_X1    g14146(.A1(new_n14330_), .A2(new_n14323_), .A3(\asqrt[57] ), .ZN(new_n14339_));
  NOR2_X1    g14147(.A1(new_n14339_), .A2(new_n14338_), .ZN(new_n14340_));
  OAI21_X1   g14148(.A1(new_n14340_), .A2(new_n14332_), .B(\asqrt[58] ), .ZN(new_n14341_));
  INV_X1     g14149(.I(new_n13780_), .ZN(new_n14342_));
  INV_X1     g14150(.I(new_n13773_), .ZN(new_n14343_));
  INV_X1     g14151(.I(new_n13782_), .ZN(new_n14344_));
  NOR2_X1    g14152(.A1(new_n14344_), .A2(new_n14343_), .ZN(new_n14345_));
  NOR3_X1    g14153(.A1(new_n14017_), .A2(new_n13774_), .A3(new_n14345_), .ZN(new_n14346_));
  INV_X1     g14154(.I(new_n14346_), .ZN(new_n14347_));
  NOR3_X1    g14155(.A1(new_n14345_), .A2(new_n13774_), .A3(new_n14342_), .ZN(new_n14348_));
  AOI22_X1   g14156(.A1(new_n14347_), .A2(new_n14342_), .B1(\asqrt[17] ), .B2(new_n14348_), .ZN(new_n14349_));
  INV_X1     g14157(.I(new_n14349_), .ZN(new_n14350_));
  NAND2_X1   g14158(.A1(new_n14331_), .A2(new_n436_), .ZN(new_n14351_));
  OAI21_X1   g14159(.A1(new_n14340_), .A2(new_n14351_), .B(new_n14350_), .ZN(new_n14352_));
  AOI21_X1   g14160(.A1(new_n14352_), .A2(new_n14341_), .B(new_n327_), .ZN(new_n14353_));
  NOR3_X1    g14161(.A1(new_n13907_), .A2(new_n13790_), .A3(new_n13908_), .ZN(new_n14354_));
  NOR3_X1    g14162(.A1(new_n14017_), .A2(new_n13907_), .A3(new_n13908_), .ZN(new_n14355_));
  INV_X1     g14163(.I(new_n14355_), .ZN(new_n14356_));
  AOI22_X1   g14164(.A1(new_n14356_), .A2(new_n13790_), .B1(\asqrt[17] ), .B2(new_n14354_), .ZN(new_n14357_));
  OAI21_X1   g14165(.A1(new_n14338_), .A2(new_n14339_), .B(new_n14331_), .ZN(new_n14358_));
  AOI21_X1   g14166(.A1(new_n14358_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n14359_));
  AOI21_X1   g14167(.A1(new_n14359_), .A2(new_n14352_), .B(new_n14357_), .ZN(new_n14360_));
  OAI21_X1   g14168(.A1(new_n14360_), .A2(new_n14353_), .B(\asqrt[60] ), .ZN(new_n14361_));
  INV_X1     g14169(.I(new_n14361_), .ZN(new_n14362_));
  INV_X1     g14170(.I(new_n13966_), .ZN(new_n14363_));
  NOR3_X1    g14171(.A1(new_n14017_), .A2(new_n13891_), .A3(new_n14363_), .ZN(new_n14364_));
  INV_X1     g14172(.I(new_n14364_), .ZN(new_n14365_));
  NOR3_X1    g14173(.A1(new_n14363_), .A2(new_n13891_), .A3(new_n13919_), .ZN(new_n14366_));
  AOI22_X1   g14174(.A1(new_n14365_), .A2(new_n13919_), .B1(\asqrt[17] ), .B2(new_n14366_), .ZN(new_n14367_));
  NOR3_X1    g14175(.A1(new_n14360_), .A2(new_n14353_), .A3(\asqrt[60] ), .ZN(new_n14368_));
  NOR2_X1    g14176(.A1(new_n14368_), .A2(new_n14367_), .ZN(new_n14369_));
  OAI21_X1   g14177(.A1(new_n14369_), .A2(new_n14362_), .B(\asqrt[61] ), .ZN(new_n14370_));
  NAND2_X1   g14178(.A1(new_n13931_), .A2(new_n13920_), .ZN(new_n14371_));
  AND3_X2    g14179(.A1(new_n13899_), .A2(new_n13905_), .A3(new_n14371_), .Z(new_n14372_));
  NAND3_X1   g14180(.A1(\asqrt[17] ), .A2(new_n13899_), .A3(new_n14371_), .ZN(new_n14373_));
  AOI22_X1   g14181(.A1(new_n14373_), .A2(new_n13906_), .B1(\asqrt[17] ), .B2(new_n14372_), .ZN(new_n14374_));
  INV_X1     g14182(.I(new_n14374_), .ZN(new_n14375_));
  NAND2_X1   g14183(.A1(new_n14361_), .A2(new_n218_), .ZN(new_n14376_));
  OAI21_X1   g14184(.A1(new_n14369_), .A2(new_n14376_), .B(new_n14375_), .ZN(new_n14377_));
  AOI21_X1   g14185(.A1(new_n14377_), .A2(new_n14370_), .B(new_n207_), .ZN(new_n14378_));
  NOR3_X1    g14186(.A1(new_n14017_), .A2(new_n13913_), .A3(new_n13944_), .ZN(new_n14379_));
  INV_X1     g14187(.I(new_n14379_), .ZN(new_n14380_));
  NOR3_X1    g14188(.A1(new_n13913_), .A2(new_n13965_), .A3(new_n13944_), .ZN(new_n14381_));
  AOI22_X1   g14189(.A1(new_n14380_), .A2(new_n13965_), .B1(\asqrt[17] ), .B2(new_n14381_), .ZN(new_n14382_));
  OAI21_X1   g14190(.A1(new_n14367_), .A2(new_n14368_), .B(new_n14361_), .ZN(new_n14383_));
  AOI21_X1   g14191(.A1(new_n14383_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n14384_));
  AOI21_X1   g14192(.A1(new_n14384_), .A2(new_n14377_), .B(new_n14382_), .ZN(new_n14385_));
  INV_X1     g14193(.I(new_n13924_), .ZN(new_n14386_));
  INV_X1     g14194(.I(new_n13978_), .ZN(new_n14387_));
  NOR3_X1    g14195(.A1(new_n14386_), .A2(new_n14387_), .A3(new_n13929_), .ZN(new_n14388_));
  NAND2_X1   g14196(.A1(\asqrt[17] ), .A2(new_n14388_), .ZN(new_n14389_));
  INV_X1     g14197(.I(new_n14389_), .ZN(new_n14390_));
  NOR2_X1    g14198(.A1(new_n14386_), .A2(new_n14387_), .ZN(new_n14391_));
  AOI21_X1   g14199(.A1(\asqrt[17] ), .A2(new_n14391_), .B(new_n13928_), .ZN(new_n14392_));
  NOR2_X1    g14200(.A1(new_n14390_), .A2(new_n14392_), .ZN(new_n14393_));
  INV_X1     g14201(.I(new_n14393_), .ZN(new_n14394_));
  NAND3_X1   g14202(.A1(\asqrt[17] ), .A2(new_n13962_), .A3(new_n13939_), .ZN(new_n14395_));
  AND3_X2    g14203(.A1(new_n14394_), .A2(new_n13992_), .A3(new_n14395_), .Z(new_n14396_));
  OAI21_X1   g14204(.A1(new_n14385_), .A2(new_n14378_), .B(new_n14396_), .ZN(new_n14397_));
  NAND2_X1   g14205(.A1(new_n14397_), .A2(new_n193_), .ZN(new_n14398_));
  INV_X1     g14206(.I(new_n14367_), .ZN(new_n14399_));
  INV_X1     g14207(.I(new_n14338_), .ZN(new_n14400_));
  INV_X1     g14208(.I(new_n14307_), .ZN(new_n14401_));
  INV_X1     g14209(.I(new_n14278_), .ZN(new_n14402_));
  INV_X1     g14210(.I(new_n14252_), .ZN(new_n14403_));
  INV_X1     g14211(.I(new_n14226_), .ZN(new_n14404_));
  INV_X1     g14212(.I(new_n14200_), .ZN(new_n14405_));
  INV_X1     g14213(.I(new_n14174_), .ZN(new_n14406_));
  INV_X1     g14214(.I(new_n14148_), .ZN(new_n14407_));
  INV_X1     g14215(.I(new_n14122_), .ZN(new_n14408_));
  INV_X1     g14216(.I(new_n14096_), .ZN(new_n14409_));
  INV_X1     g14217(.I(new_n14070_), .ZN(new_n14410_));
  INV_X1     g14218(.I(new_n14044_), .ZN(new_n14411_));
  NAND2_X1   g14219(.A1(new_n13975_), .A2(new_n13983_), .ZN(new_n14412_));
  OAI21_X1   g14220(.A1(new_n13964_), .A2(new_n13974_), .B(new_n13977_), .ZN(new_n14413_));
  NAND2_X1   g14221(.A1(new_n14413_), .A2(\a[35] ), .ZN(new_n14414_));
  NAND3_X1   g14222(.A1(new_n14412_), .A2(new_n14414_), .A3(new_n13991_), .ZN(new_n14415_));
  AOI21_X1   g14223(.A1(new_n14415_), .A2(new_n14006_), .B(new_n12913_), .ZN(new_n14416_));
  OAI21_X1   g14224(.A1(new_n13997_), .A2(new_n13986_), .B(\a[36] ), .ZN(new_n14417_));
  NAND3_X1   g14225(.A1(new_n13994_), .A2(new_n13991_), .A3(new_n13354_), .ZN(new_n14418_));
  NAND2_X1   g14226(.A1(new_n13975_), .A2(new_n13961_), .ZN(new_n14419_));
  AOI21_X1   g14227(.A1(new_n14419_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n14420_));
  AOI22_X1   g14228(.A1(new_n14415_), .A2(new_n14420_), .B1(new_n14417_), .B2(new_n14418_), .ZN(new_n14421_));
  OAI21_X1   g14229(.A1(new_n14421_), .A2(new_n14416_), .B(\asqrt[20] ), .ZN(new_n14422_));
  NAND2_X1   g14230(.A1(new_n14422_), .A2(new_n11736_), .ZN(new_n14423_));
  OAI21_X1   g14231(.A1(new_n14423_), .A2(new_n14011_), .B(new_n14019_), .ZN(new_n14424_));
  AOI21_X1   g14232(.A1(new_n14424_), .A2(new_n14012_), .B(new_n11326_), .ZN(new_n14425_));
  INV_X1     g14233(.I(new_n14005_), .ZN(new_n14426_));
  AOI21_X1   g14234(.A1(\a[35] ), .A2(new_n14413_), .B(new_n13986_), .ZN(new_n14427_));
  AOI21_X1   g14235(.A1(new_n14427_), .A2(new_n14412_), .B(new_n13976_), .ZN(new_n14428_));
  OAI21_X1   g14236(.A1(new_n14428_), .A2(new_n12913_), .B(new_n12364_), .ZN(new_n14429_));
  OAI21_X1   g14237(.A1(new_n14429_), .A2(new_n14421_), .B(new_n14426_), .ZN(new_n14430_));
  NAND2_X1   g14238(.A1(new_n14430_), .A2(new_n14422_), .ZN(new_n14431_));
  AOI21_X1   g14239(.A1(new_n14431_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n14432_));
  AOI21_X1   g14240(.A1(new_n14432_), .A2(new_n14424_), .B(new_n14027_), .ZN(new_n14433_));
  OAI21_X1   g14241(.A1(new_n14433_), .A2(new_n14425_), .B(\asqrt[23] ), .ZN(new_n14434_));
  NAND2_X1   g14242(.A1(new_n14434_), .A2(new_n10221_), .ZN(new_n14435_));
  OAI21_X1   g14243(.A1(new_n14435_), .A2(new_n14038_), .B(new_n14411_), .ZN(new_n14436_));
  NAND3_X1   g14244(.A1(new_n14436_), .A2(new_n9846_), .A3(new_n14039_), .ZN(new_n14437_));
  AOI22_X1   g14245(.A1(new_n14437_), .A2(new_n14053_), .B1(new_n14061_), .B2(\asqrt[25] ), .ZN(new_n14438_));
  OAI21_X1   g14246(.A1(new_n14438_), .A2(new_n9317_), .B(new_n8826_), .ZN(new_n14439_));
  OAI21_X1   g14247(.A1(new_n14439_), .A2(new_n14063_), .B(new_n14410_), .ZN(new_n14440_));
  AOI21_X1   g14248(.A1(new_n14440_), .A2(new_n14064_), .B(new_n8483_), .ZN(new_n14441_));
  AOI21_X1   g14249(.A1(new_n14436_), .A2(new_n14039_), .B(new_n9846_), .ZN(new_n14442_));
  NOR3_X1    g14250(.A1(new_n14433_), .A2(new_n14425_), .A3(\asqrt[23] ), .ZN(new_n14443_));
  OAI21_X1   g14251(.A1(new_n14035_), .A2(new_n14443_), .B(new_n14434_), .ZN(new_n14444_));
  AOI21_X1   g14252(.A1(new_n14444_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n14445_));
  AOI21_X1   g14253(.A1(new_n14445_), .A2(new_n14436_), .B(new_n14052_), .ZN(new_n14446_));
  NOR3_X1    g14254(.A1(new_n14446_), .A2(\asqrt[26] ), .A3(new_n14442_), .ZN(new_n14447_));
  OAI22_X1   g14255(.A1(new_n14447_), .A2(new_n14060_), .B1(new_n14438_), .B2(new_n9317_), .ZN(new_n14448_));
  AOI21_X1   g14256(.A1(new_n14448_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n14449_));
  AOI21_X1   g14257(.A1(new_n14449_), .A2(new_n14440_), .B(new_n14078_), .ZN(new_n14450_));
  OAI21_X1   g14258(.A1(new_n14450_), .A2(new_n14441_), .B(\asqrt[29] ), .ZN(new_n14451_));
  NAND2_X1   g14259(.A1(new_n14451_), .A2(new_n7539_), .ZN(new_n14452_));
  OAI21_X1   g14260(.A1(new_n14452_), .A2(new_n14089_), .B(new_n14409_), .ZN(new_n14453_));
  AOI21_X1   g14261(.A1(new_n14453_), .A2(new_n14090_), .B(new_n7229_), .ZN(new_n14454_));
  NOR3_X1    g14262(.A1(new_n14450_), .A2(\asqrt[29] ), .A3(new_n14441_), .ZN(new_n14455_));
  OAI21_X1   g14263(.A1(new_n14086_), .A2(new_n14455_), .B(new_n14451_), .ZN(new_n14456_));
  AOI21_X1   g14264(.A1(new_n14456_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n14457_));
  AOI21_X1   g14265(.A1(new_n14457_), .A2(new_n14453_), .B(new_n14104_), .ZN(new_n14458_));
  OAI21_X1   g14266(.A1(new_n14458_), .A2(new_n14454_), .B(\asqrt[32] ), .ZN(new_n14459_));
  NAND2_X1   g14267(.A1(new_n14459_), .A2(new_n6356_), .ZN(new_n14460_));
  OAI21_X1   g14268(.A1(new_n14460_), .A2(new_n14115_), .B(new_n14408_), .ZN(new_n14461_));
  AOI21_X1   g14269(.A1(new_n14461_), .A2(new_n14116_), .B(new_n6077_), .ZN(new_n14462_));
  NOR3_X1    g14270(.A1(new_n14458_), .A2(\asqrt[32] ), .A3(new_n14454_), .ZN(new_n14463_));
  OAI21_X1   g14271(.A1(new_n14112_), .A2(new_n14463_), .B(new_n14459_), .ZN(new_n14464_));
  AOI21_X1   g14272(.A1(new_n14464_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n14465_));
  AOI21_X1   g14273(.A1(new_n14465_), .A2(new_n14461_), .B(new_n14130_), .ZN(new_n14466_));
  OAI21_X1   g14274(.A1(new_n14466_), .A2(new_n14462_), .B(\asqrt[35] ), .ZN(new_n14467_));
  NAND2_X1   g14275(.A1(new_n14467_), .A2(new_n5277_), .ZN(new_n14468_));
  OAI21_X1   g14276(.A1(new_n14468_), .A2(new_n14141_), .B(new_n14407_), .ZN(new_n14469_));
  AOI21_X1   g14277(.A1(new_n14469_), .A2(new_n14142_), .B(new_n5024_), .ZN(new_n14470_));
  NOR3_X1    g14278(.A1(new_n14466_), .A2(\asqrt[35] ), .A3(new_n14462_), .ZN(new_n14471_));
  OAI21_X1   g14279(.A1(new_n14138_), .A2(new_n14471_), .B(new_n14467_), .ZN(new_n14472_));
  AOI21_X1   g14280(.A1(new_n14472_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n14473_));
  AOI21_X1   g14281(.A1(new_n14473_), .A2(new_n14469_), .B(new_n14156_), .ZN(new_n14474_));
  OAI21_X1   g14282(.A1(new_n14474_), .A2(new_n14470_), .B(\asqrt[38] ), .ZN(new_n14475_));
  NAND2_X1   g14283(.A1(new_n14475_), .A2(new_n4298_), .ZN(new_n14476_));
  OAI21_X1   g14284(.A1(new_n14476_), .A2(new_n14167_), .B(new_n14406_), .ZN(new_n14477_));
  AOI21_X1   g14285(.A1(new_n14477_), .A2(new_n14168_), .B(new_n4071_), .ZN(new_n14478_));
  NOR3_X1    g14286(.A1(new_n14474_), .A2(\asqrt[38] ), .A3(new_n14470_), .ZN(new_n14479_));
  OAI21_X1   g14287(.A1(new_n14164_), .A2(new_n14479_), .B(new_n14475_), .ZN(new_n14480_));
  AOI21_X1   g14288(.A1(new_n14480_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n14481_));
  AOI21_X1   g14289(.A1(new_n14481_), .A2(new_n14477_), .B(new_n14182_), .ZN(new_n14482_));
  OAI21_X1   g14290(.A1(new_n14482_), .A2(new_n14478_), .B(\asqrt[41] ), .ZN(new_n14483_));
  NAND2_X1   g14291(.A1(new_n14483_), .A2(new_n3419_), .ZN(new_n14484_));
  OAI21_X1   g14292(.A1(new_n14484_), .A2(new_n14193_), .B(new_n14405_), .ZN(new_n14485_));
  AOI21_X1   g14293(.A1(new_n14485_), .A2(new_n14194_), .B(new_n3218_), .ZN(new_n14486_));
  NOR3_X1    g14294(.A1(new_n14482_), .A2(\asqrt[41] ), .A3(new_n14478_), .ZN(new_n14487_));
  OAI21_X1   g14295(.A1(new_n14190_), .A2(new_n14487_), .B(new_n14483_), .ZN(new_n14488_));
  AOI21_X1   g14296(.A1(new_n14488_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n14489_));
  AOI21_X1   g14297(.A1(new_n14489_), .A2(new_n14485_), .B(new_n14208_), .ZN(new_n14490_));
  OAI21_X1   g14298(.A1(new_n14490_), .A2(new_n14486_), .B(\asqrt[44] ), .ZN(new_n14491_));
  NAND2_X1   g14299(.A1(new_n14491_), .A2(new_n2641_), .ZN(new_n14492_));
  OAI21_X1   g14300(.A1(new_n14492_), .A2(new_n14219_), .B(new_n14404_), .ZN(new_n14493_));
  AOI21_X1   g14301(.A1(new_n14493_), .A2(new_n14220_), .B(new_n2465_), .ZN(new_n14494_));
  NOR3_X1    g14302(.A1(new_n14490_), .A2(\asqrt[44] ), .A3(new_n14486_), .ZN(new_n14495_));
  OAI21_X1   g14303(.A1(new_n14216_), .A2(new_n14495_), .B(new_n14491_), .ZN(new_n14496_));
  AOI21_X1   g14304(.A1(new_n14496_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n14497_));
  AOI21_X1   g14305(.A1(new_n14497_), .A2(new_n14493_), .B(new_n14234_), .ZN(new_n14498_));
  OAI21_X1   g14306(.A1(new_n14498_), .A2(new_n14494_), .B(\asqrt[47] ), .ZN(new_n14499_));
  NAND2_X1   g14307(.A1(new_n14499_), .A2(new_n1956_), .ZN(new_n14500_));
  OAI21_X1   g14308(.A1(new_n14500_), .A2(new_n14245_), .B(new_n14403_), .ZN(new_n14501_));
  AOI21_X1   g14309(.A1(new_n14501_), .A2(new_n14246_), .B(new_n1806_), .ZN(new_n14502_));
  NOR3_X1    g14310(.A1(new_n14498_), .A2(\asqrt[47] ), .A3(new_n14494_), .ZN(new_n14503_));
  OAI21_X1   g14311(.A1(new_n14242_), .A2(new_n14503_), .B(new_n14499_), .ZN(new_n14504_));
  AOI21_X1   g14312(.A1(new_n14504_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n14505_));
  AOI21_X1   g14313(.A1(new_n14505_), .A2(new_n14501_), .B(new_n14260_), .ZN(new_n14506_));
  OAI21_X1   g14314(.A1(new_n14506_), .A2(new_n14502_), .B(\asqrt[50] ), .ZN(new_n14507_));
  NAND2_X1   g14315(.A1(new_n14507_), .A2(new_n1376_), .ZN(new_n14508_));
  OAI21_X1   g14316(.A1(new_n14508_), .A2(new_n14271_), .B(new_n14402_), .ZN(new_n14509_));
  AOI21_X1   g14317(.A1(new_n14509_), .A2(new_n14272_), .B(new_n1256_), .ZN(new_n14510_));
  NOR3_X1    g14318(.A1(new_n14506_), .A2(\asqrt[50] ), .A3(new_n14502_), .ZN(new_n14511_));
  OAI21_X1   g14319(.A1(new_n14268_), .A2(new_n14511_), .B(new_n14507_), .ZN(new_n14512_));
  AOI21_X1   g14320(.A1(new_n14512_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n14513_));
  AOI21_X1   g14321(.A1(new_n14513_), .A2(new_n14509_), .B(new_n14288_), .ZN(new_n14514_));
  OAI21_X1   g14322(.A1(new_n14514_), .A2(new_n14510_), .B(\asqrt[53] ), .ZN(new_n14515_));
  NAND2_X1   g14323(.A1(new_n14515_), .A2(new_n904_), .ZN(new_n14516_));
  OAI21_X1   g14324(.A1(new_n14516_), .A2(new_n14299_), .B(new_n14401_), .ZN(new_n14517_));
  AOI21_X1   g14325(.A1(new_n14517_), .A2(new_n14300_), .B(new_n823_), .ZN(new_n14518_));
  NOR3_X1    g14326(.A1(new_n14514_), .A2(\asqrt[53] ), .A3(new_n14510_), .ZN(new_n14519_));
  OAI21_X1   g14327(.A1(new_n14296_), .A2(new_n14519_), .B(new_n14515_), .ZN(new_n14520_));
  AOI21_X1   g14328(.A1(new_n14520_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n14521_));
  AOI21_X1   g14329(.A1(new_n14521_), .A2(new_n14517_), .B(new_n14319_), .ZN(new_n14522_));
  OAI21_X1   g14330(.A1(new_n14522_), .A2(new_n14518_), .B(\asqrt[56] ), .ZN(new_n14523_));
  NAND2_X1   g14331(.A1(new_n14523_), .A2(new_n531_), .ZN(new_n14524_));
  OAI21_X1   g14332(.A1(new_n14524_), .A2(new_n14330_), .B(new_n14400_), .ZN(new_n14525_));
  AOI21_X1   g14333(.A1(new_n14525_), .A2(new_n14331_), .B(new_n436_), .ZN(new_n14526_));
  NOR3_X1    g14334(.A1(new_n14522_), .A2(\asqrt[56] ), .A3(new_n14518_), .ZN(new_n14527_));
  OAI21_X1   g14335(.A1(new_n14327_), .A2(new_n14527_), .B(new_n14523_), .ZN(new_n14528_));
  AOI21_X1   g14336(.A1(new_n14528_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n14529_));
  AOI21_X1   g14337(.A1(new_n14529_), .A2(new_n14525_), .B(new_n14349_), .ZN(new_n14530_));
  OAI21_X1   g14338(.A1(new_n14530_), .A2(new_n14526_), .B(\asqrt[59] ), .ZN(new_n14531_));
  NAND2_X1   g14339(.A1(new_n14531_), .A2(new_n306_), .ZN(new_n14532_));
  OAI21_X1   g14340(.A1(new_n14532_), .A2(new_n14360_), .B(new_n14399_), .ZN(new_n14533_));
  NOR3_X1    g14341(.A1(new_n14530_), .A2(\asqrt[59] ), .A3(new_n14526_), .ZN(new_n14534_));
  OAI21_X1   g14342(.A1(new_n14357_), .A2(new_n14534_), .B(new_n14531_), .ZN(new_n14535_));
  AOI21_X1   g14343(.A1(new_n14535_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n14536_));
  AOI21_X1   g14344(.A1(new_n14536_), .A2(new_n14533_), .B(new_n14374_), .ZN(new_n14537_));
  INV_X1     g14345(.I(new_n14382_), .ZN(new_n14538_));
  NAND2_X1   g14346(.A1(new_n14370_), .A2(new_n207_), .ZN(new_n14539_));
  OAI21_X1   g14347(.A1(new_n14539_), .A2(new_n14537_), .B(new_n14538_), .ZN(new_n14540_));
  NOR2_X1    g14348(.A1(new_n14378_), .A2(new_n14394_), .ZN(new_n14541_));
  NAND2_X1   g14349(.A1(\asqrt[17] ), .A2(new_n13939_), .ZN(new_n14542_));
  OAI21_X1   g14350(.A1(new_n13979_), .A2(new_n13972_), .B(\asqrt[63] ), .ZN(new_n14543_));
  AOI21_X1   g14351(.A1(new_n14542_), .A2(new_n13979_), .B(new_n14543_), .ZN(new_n14544_));
  AND2_X2    g14352(.A1(new_n13936_), .A2(new_n13952_), .Z(new_n14545_));
  NAND4_X1   g14353(.A1(new_n13992_), .A2(new_n13938_), .A3(new_n13949_), .A4(new_n14545_), .ZN(new_n14546_));
  NOR2_X1    g14354(.A1(new_n14546_), .A2(new_n13964_), .ZN(new_n14547_));
  NOR2_X1    g14355(.A1(new_n14544_), .A2(new_n14547_), .ZN(new_n14548_));
  INV_X1     g14356(.I(new_n14548_), .ZN(new_n14549_));
  AOI21_X1   g14357(.A1(new_n14541_), .A2(new_n14540_), .B(new_n14549_), .ZN(new_n14550_));
  NAND2_X1   g14358(.A1(new_n14398_), .A2(new_n14550_), .ZN(\asqrt[16] ));
  NOR2_X1    g14359(.A1(\a[30] ), .A2(\a[31] ), .ZN(new_n14552_));
  INV_X1     g14360(.I(new_n14552_), .ZN(new_n14553_));
  NOR2_X1    g14361(.A1(new_n14553_), .A2(\a[32] ), .ZN(new_n14554_));
  INV_X1     g14362(.I(new_n14554_), .ZN(new_n14555_));
  AOI21_X1   g14363(.A1(new_n14533_), .A2(new_n14361_), .B(new_n218_), .ZN(new_n14556_));
  OAI21_X1   g14364(.A1(new_n14537_), .A2(new_n14556_), .B(\asqrt[62] ), .ZN(new_n14557_));
  NOR3_X1    g14365(.A1(new_n14537_), .A2(\asqrt[62] ), .A3(new_n14556_), .ZN(new_n14558_));
  OAI21_X1   g14366(.A1(new_n14382_), .A2(new_n14558_), .B(new_n14557_), .ZN(new_n14559_));
  AOI21_X1   g14367(.A1(new_n14559_), .A2(new_n14396_), .B(\asqrt[63] ), .ZN(new_n14560_));
  NAND2_X1   g14368(.A1(new_n14557_), .A2(new_n14393_), .ZN(new_n14561_));
  OAI21_X1   g14369(.A1(new_n14561_), .A2(new_n14385_), .B(new_n14548_), .ZN(new_n14562_));
  OAI21_X1   g14370(.A1(new_n14560_), .A2(new_n14562_), .B(\a[32] ), .ZN(new_n14563_));
  AOI21_X1   g14371(.A1(new_n14563_), .A2(new_n14555_), .B(new_n14017_), .ZN(new_n14564_));
  INV_X1     g14372(.I(\a[32] ), .ZN(new_n14565_));
  AOI21_X1   g14373(.A1(new_n14398_), .A2(new_n14550_), .B(new_n14565_), .ZN(new_n14566_));
  NAND4_X1   g14374(.A1(new_n13992_), .A2(new_n13949_), .A3(new_n13952_), .A4(new_n14555_), .ZN(new_n14567_));
  NOR2_X1    g14375(.A1(new_n14567_), .A2(new_n13964_), .ZN(new_n14568_));
  INV_X1     g14376(.I(new_n14568_), .ZN(new_n14569_));
  NOR2_X1    g14377(.A1(new_n14566_), .A2(new_n14569_), .ZN(new_n14570_));
  AOI21_X1   g14378(.A1(new_n14398_), .A2(new_n14550_), .B(new_n13959_), .ZN(new_n14571_));
  INV_X1     g14379(.I(\a[33] ), .ZN(new_n14572_));
  AOI21_X1   g14380(.A1(\asqrt[16] ), .A2(new_n14565_), .B(new_n14572_), .ZN(new_n14573_));
  NOR3_X1    g14381(.A1(new_n14570_), .A2(new_n14573_), .A3(new_n14571_), .ZN(new_n14574_));
  OAI21_X1   g14382(.A1(new_n14574_), .A2(new_n14564_), .B(\asqrt[18] ), .ZN(new_n14575_));
  OAI21_X1   g14383(.A1(new_n14560_), .A2(new_n14562_), .B(new_n13958_), .ZN(new_n14576_));
  NAND2_X1   g14384(.A1(new_n14541_), .A2(new_n14540_), .ZN(new_n14577_));
  NOR3_X1    g14385(.A1(new_n14544_), .A2(new_n14017_), .A3(new_n14547_), .ZN(new_n14578_));
  NAND3_X1   g14386(.A1(new_n14398_), .A2(new_n14577_), .A3(new_n14578_), .ZN(new_n14579_));
  AOI21_X1   g14387(.A1(new_n14576_), .A2(new_n14579_), .B(new_n13977_), .ZN(new_n14580_));
  AND3_X2    g14388(.A1(new_n14398_), .A2(new_n14577_), .A3(new_n14578_), .Z(new_n14581_));
  NOR3_X1    g14389(.A1(new_n14581_), .A2(\a[34] ), .A3(new_n14571_), .ZN(new_n14582_));
  OAI21_X1   g14390(.A1(new_n14566_), .A2(new_n14554_), .B(\asqrt[17] ), .ZN(new_n14583_));
  NAND2_X1   g14391(.A1(new_n14583_), .A2(new_n13353_), .ZN(new_n14584_));
  OAI22_X1   g14392(.A1(new_n14574_), .A2(new_n14584_), .B1(new_n14580_), .B2(new_n14582_), .ZN(new_n14585_));
  AOI21_X1   g14393(.A1(new_n14585_), .A2(new_n14575_), .B(new_n12913_), .ZN(new_n14586_));
  NOR3_X1    g14394(.A1(new_n14427_), .A2(new_n13976_), .A3(new_n13985_), .ZN(new_n14587_));
  NAND3_X1   g14395(.A1(\asqrt[16] ), .A2(new_n14006_), .A3(new_n14412_), .ZN(new_n14588_));
  AOI22_X1   g14396(.A1(new_n14588_), .A2(new_n14427_), .B1(\asqrt[16] ), .B2(new_n14587_), .ZN(new_n14589_));
  AOI21_X1   g14397(.A1(new_n14398_), .A2(new_n14550_), .B(\a[32] ), .ZN(new_n14590_));
  OAI21_X1   g14398(.A1(new_n14572_), .A2(new_n14590_), .B(new_n14576_), .ZN(new_n14591_));
  OAI21_X1   g14399(.A1(new_n14591_), .A2(new_n14570_), .B(new_n14583_), .ZN(new_n14592_));
  AOI21_X1   g14400(.A1(new_n14592_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n14593_));
  AOI21_X1   g14401(.A1(new_n14593_), .A2(new_n14585_), .B(new_n14589_), .ZN(new_n14594_));
  OAI21_X1   g14402(.A1(new_n14594_), .A2(new_n14586_), .B(\asqrt[20] ), .ZN(new_n14595_));
  INV_X1     g14403(.I(new_n14595_), .ZN(new_n14596_));
  NOR2_X1    g14404(.A1(new_n13998_), .A2(new_n13995_), .ZN(new_n14597_));
  NOR2_X1    g14405(.A1(new_n13989_), .A2(new_n14000_), .ZN(new_n14598_));
  INV_X1     g14406(.I(new_n14598_), .ZN(new_n14599_));
  NAND4_X1   g14407(.A1(\asqrt[16] ), .A2(new_n13990_), .A3(new_n14597_), .A4(new_n14599_), .ZN(new_n14600_));
  INV_X1     g14408(.I(\asqrt[16] ), .ZN(new_n14601_));
  NOR3_X1    g14409(.A1(new_n14601_), .A2(new_n14416_), .A3(new_n14598_), .ZN(new_n14602_));
  OAI21_X1   g14410(.A1(new_n14602_), .A2(new_n14597_), .B(new_n14600_), .ZN(new_n14603_));
  INV_X1     g14411(.I(new_n14603_), .ZN(new_n14604_));
  NOR3_X1    g14412(.A1(new_n14594_), .A2(new_n14586_), .A3(\asqrt[20] ), .ZN(new_n14605_));
  NOR2_X1    g14413(.A1(new_n14605_), .A2(new_n14604_), .ZN(new_n14606_));
  OAI21_X1   g14414(.A1(new_n14606_), .A2(new_n14596_), .B(\asqrt[21] ), .ZN(new_n14607_));
  NOR2_X1    g14415(.A1(new_n14429_), .A2(new_n14421_), .ZN(new_n14608_));
  NOR3_X1    g14416(.A1(new_n14601_), .A2(new_n14002_), .A3(new_n14608_), .ZN(new_n14609_));
  INV_X1     g14417(.I(new_n14609_), .ZN(new_n14610_));
  NOR3_X1    g14418(.A1(new_n14608_), .A2(new_n14002_), .A3(new_n14426_), .ZN(new_n14611_));
  AOI22_X1   g14419(.A1(new_n14610_), .A2(new_n14426_), .B1(\asqrt[16] ), .B2(new_n14611_), .ZN(new_n14612_));
  INV_X1     g14420(.I(new_n14612_), .ZN(new_n14613_));
  NAND2_X1   g14421(.A1(new_n14595_), .A2(new_n11736_), .ZN(new_n14614_));
  OAI21_X1   g14422(.A1(new_n14606_), .A2(new_n14614_), .B(new_n14613_), .ZN(new_n14615_));
  AOI21_X1   g14423(.A1(new_n14615_), .A2(new_n14607_), .B(new_n11326_), .ZN(new_n14616_));
  NOR3_X1    g14424(.A1(new_n14013_), .A2(new_n14021_), .A3(new_n14019_), .ZN(new_n14617_));
  NOR3_X1    g14425(.A1(new_n14601_), .A2(new_n14013_), .A3(new_n14021_), .ZN(new_n14618_));
  INV_X1     g14426(.I(new_n14618_), .ZN(new_n14619_));
  AOI22_X1   g14427(.A1(new_n14619_), .A2(new_n14019_), .B1(\asqrt[16] ), .B2(new_n14617_), .ZN(new_n14620_));
  OAI21_X1   g14428(.A1(new_n14604_), .A2(new_n14605_), .B(new_n14595_), .ZN(new_n14621_));
  AOI21_X1   g14429(.A1(new_n14621_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n14622_));
  AOI21_X1   g14430(.A1(new_n14622_), .A2(new_n14615_), .B(new_n14620_), .ZN(new_n14623_));
  OAI21_X1   g14431(.A1(new_n14623_), .A2(new_n14616_), .B(\asqrt[23] ), .ZN(new_n14624_));
  NAND2_X1   g14432(.A1(new_n14432_), .A2(new_n14424_), .ZN(new_n14625_));
  NAND3_X1   g14433(.A1(\asqrt[16] ), .A2(new_n14023_), .A3(new_n14625_), .ZN(new_n14626_));
  AND3_X2    g14434(.A1(new_n14023_), .A2(new_n14027_), .A3(new_n14625_), .Z(new_n14627_));
  AOI22_X1   g14435(.A1(new_n14626_), .A2(new_n14028_), .B1(\asqrt[16] ), .B2(new_n14627_), .ZN(new_n14628_));
  INV_X1     g14436(.I(new_n14628_), .ZN(new_n14629_));
  NAND2_X1   g14437(.A1(new_n14563_), .A2(new_n14568_), .ZN(new_n14630_));
  OAI21_X1   g14438(.A1(new_n14560_), .A2(new_n14562_), .B(new_n14565_), .ZN(new_n14631_));
  NAND2_X1   g14439(.A1(new_n14631_), .A2(\a[33] ), .ZN(new_n14632_));
  NAND3_X1   g14440(.A1(new_n14630_), .A2(new_n14632_), .A3(new_n14576_), .ZN(new_n14633_));
  AOI21_X1   g14441(.A1(new_n14633_), .A2(new_n14583_), .B(new_n13353_), .ZN(new_n14634_));
  OAI21_X1   g14442(.A1(new_n14581_), .A2(new_n14571_), .B(\a[34] ), .ZN(new_n14635_));
  NAND3_X1   g14443(.A1(new_n14576_), .A2(new_n14579_), .A3(new_n13977_), .ZN(new_n14636_));
  NAND2_X1   g14444(.A1(new_n14563_), .A2(new_n14555_), .ZN(new_n14637_));
  AOI21_X1   g14445(.A1(new_n14637_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n14638_));
  AOI22_X1   g14446(.A1(new_n14633_), .A2(new_n14638_), .B1(new_n14635_), .B2(new_n14636_), .ZN(new_n14639_));
  OAI21_X1   g14447(.A1(new_n14639_), .A2(new_n14634_), .B(\asqrt[19] ), .ZN(new_n14640_));
  NAND2_X1   g14448(.A1(new_n14640_), .A2(new_n12364_), .ZN(new_n14641_));
  OAI21_X1   g14449(.A1(new_n14641_), .A2(new_n14594_), .B(new_n14603_), .ZN(new_n14642_));
  AOI21_X1   g14450(.A1(new_n14642_), .A2(new_n14595_), .B(new_n11736_), .ZN(new_n14643_));
  INV_X1     g14451(.I(new_n14589_), .ZN(new_n14644_));
  AOI21_X1   g14452(.A1(\a[33] ), .A2(new_n14631_), .B(new_n14571_), .ZN(new_n14645_));
  AOI21_X1   g14453(.A1(new_n14645_), .A2(new_n14630_), .B(new_n14564_), .ZN(new_n14646_));
  OAI21_X1   g14454(.A1(new_n14646_), .A2(new_n13353_), .B(new_n12913_), .ZN(new_n14647_));
  OAI21_X1   g14455(.A1(new_n14647_), .A2(new_n14639_), .B(new_n14644_), .ZN(new_n14648_));
  NAND2_X1   g14456(.A1(new_n14648_), .A2(new_n14640_), .ZN(new_n14649_));
  AOI21_X1   g14457(.A1(new_n14649_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n14650_));
  AOI21_X1   g14458(.A1(new_n14650_), .A2(new_n14642_), .B(new_n14612_), .ZN(new_n14651_));
  OAI21_X1   g14459(.A1(new_n14651_), .A2(new_n14643_), .B(\asqrt[22] ), .ZN(new_n14652_));
  NAND2_X1   g14460(.A1(new_n14652_), .A2(new_n10812_), .ZN(new_n14653_));
  OAI21_X1   g14461(.A1(new_n14653_), .A2(new_n14623_), .B(new_n14629_), .ZN(new_n14654_));
  AOI21_X1   g14462(.A1(new_n14654_), .A2(new_n14624_), .B(new_n10221_), .ZN(new_n14655_));
  INV_X1     g14463(.I(new_n14035_), .ZN(new_n14656_));
  NOR3_X1    g14464(.A1(new_n14031_), .A2(new_n14443_), .A3(new_n14656_), .ZN(new_n14657_));
  NOR3_X1    g14465(.A1(new_n14601_), .A2(new_n14031_), .A3(new_n14443_), .ZN(new_n14658_));
  INV_X1     g14466(.I(new_n14658_), .ZN(new_n14659_));
  AOI22_X1   g14467(.A1(new_n14659_), .A2(new_n14656_), .B1(\asqrt[16] ), .B2(new_n14657_), .ZN(new_n14660_));
  NOR3_X1    g14468(.A1(new_n14651_), .A2(new_n14643_), .A3(\asqrt[22] ), .ZN(new_n14661_));
  OAI21_X1   g14469(.A1(new_n14620_), .A2(new_n14661_), .B(new_n14652_), .ZN(new_n14662_));
  AOI21_X1   g14470(.A1(new_n14662_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n14663_));
  AOI21_X1   g14471(.A1(new_n14663_), .A2(new_n14654_), .B(new_n14660_), .ZN(new_n14664_));
  OAI21_X1   g14472(.A1(new_n14664_), .A2(new_n14655_), .B(\asqrt[25] ), .ZN(new_n14665_));
  INV_X1     g14473(.I(new_n14665_), .ZN(new_n14666_));
  NOR3_X1    g14474(.A1(new_n14601_), .A2(new_n14040_), .A3(new_n14045_), .ZN(new_n14667_));
  INV_X1     g14475(.I(new_n14667_), .ZN(new_n14668_));
  NOR3_X1    g14476(.A1(new_n14040_), .A2(new_n14411_), .A3(new_n14045_), .ZN(new_n14669_));
  AOI22_X1   g14477(.A1(new_n14668_), .A2(new_n14411_), .B1(\asqrt[16] ), .B2(new_n14669_), .ZN(new_n14670_));
  NOR3_X1    g14478(.A1(new_n14664_), .A2(\asqrt[25] ), .A3(new_n14655_), .ZN(new_n14671_));
  NOR2_X1    g14479(.A1(new_n14671_), .A2(new_n14670_), .ZN(new_n14672_));
  OAI21_X1   g14480(.A1(new_n14672_), .A2(new_n14666_), .B(\asqrt[26] ), .ZN(new_n14673_));
  AND3_X2    g14481(.A1(new_n14047_), .A2(new_n14052_), .A3(new_n14437_), .Z(new_n14674_));
  NAND3_X1   g14482(.A1(\asqrt[16] ), .A2(new_n14047_), .A3(new_n14437_), .ZN(new_n14675_));
  AOI22_X1   g14483(.A1(new_n14675_), .A2(new_n14053_), .B1(\asqrt[16] ), .B2(new_n14674_), .ZN(new_n14676_));
  INV_X1     g14484(.I(new_n14676_), .ZN(new_n14677_));
  NAND2_X1   g14485(.A1(new_n14665_), .A2(new_n9317_), .ZN(new_n14678_));
  OAI21_X1   g14486(.A1(new_n14672_), .A2(new_n14678_), .B(new_n14677_), .ZN(new_n14679_));
  AOI21_X1   g14487(.A1(new_n14679_), .A2(new_n14673_), .B(new_n8826_), .ZN(new_n14680_));
  INV_X1     g14488(.I(new_n14060_), .ZN(new_n14681_));
  NOR3_X1    g14489(.A1(new_n14601_), .A2(new_n14056_), .A3(new_n14447_), .ZN(new_n14682_));
  INV_X1     g14490(.I(new_n14682_), .ZN(new_n14683_));
  NOR3_X1    g14491(.A1(new_n14056_), .A2(new_n14447_), .A3(new_n14681_), .ZN(new_n14684_));
  AOI22_X1   g14492(.A1(new_n14683_), .A2(new_n14681_), .B1(\asqrt[16] ), .B2(new_n14684_), .ZN(new_n14685_));
  NOR3_X1    g14493(.A1(new_n14623_), .A2(new_n14616_), .A3(\asqrt[23] ), .ZN(new_n14686_));
  OAI21_X1   g14494(.A1(new_n14628_), .A2(new_n14686_), .B(new_n14624_), .ZN(new_n14687_));
  INV_X1     g14495(.I(new_n14660_), .ZN(new_n14688_));
  NAND3_X1   g14496(.A1(new_n14654_), .A2(new_n10221_), .A3(new_n14624_), .ZN(new_n14689_));
  AOI22_X1   g14497(.A1(new_n14689_), .A2(new_n14688_), .B1(new_n14687_), .B2(\asqrt[24] ), .ZN(new_n14690_));
  OAI22_X1   g14498(.A1(new_n14671_), .A2(new_n14670_), .B1(new_n14690_), .B2(new_n9846_), .ZN(new_n14691_));
  AOI21_X1   g14499(.A1(new_n14691_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n14692_));
  AOI21_X1   g14500(.A1(new_n14692_), .A2(new_n14679_), .B(new_n14685_), .ZN(new_n14693_));
  OAI21_X1   g14501(.A1(new_n14693_), .A2(new_n14680_), .B(\asqrt[28] ), .ZN(new_n14694_));
  INV_X1     g14502(.I(new_n14694_), .ZN(new_n14695_));
  INV_X1     g14503(.I(new_n14693_), .ZN(new_n14696_));
  NOR3_X1    g14504(.A1(new_n14065_), .A2(new_n14410_), .A3(new_n14071_), .ZN(new_n14697_));
  NOR3_X1    g14505(.A1(new_n14601_), .A2(new_n14065_), .A3(new_n14071_), .ZN(new_n14698_));
  INV_X1     g14506(.I(new_n14698_), .ZN(new_n14699_));
  AOI22_X1   g14507(.A1(new_n14699_), .A2(new_n14410_), .B1(\asqrt[16] ), .B2(new_n14697_), .ZN(new_n14700_));
  NOR2_X1    g14508(.A1(new_n14680_), .A2(\asqrt[28] ), .ZN(new_n14701_));
  AOI21_X1   g14509(.A1(new_n14696_), .A2(new_n14701_), .B(new_n14700_), .ZN(new_n14702_));
  OAI21_X1   g14510(.A1(new_n14702_), .A2(new_n14695_), .B(\asqrt[29] ), .ZN(new_n14703_));
  NOR2_X1    g14511(.A1(new_n14072_), .A2(new_n14080_), .ZN(new_n14704_));
  NOR3_X1    g14512(.A1(new_n14601_), .A2(new_n14441_), .A3(new_n14704_), .ZN(new_n14705_));
  INV_X1     g14513(.I(new_n14705_), .ZN(new_n14706_));
  NOR3_X1    g14514(.A1(new_n14704_), .A2(new_n14441_), .A3(new_n14079_), .ZN(new_n14707_));
  AOI22_X1   g14515(.A1(new_n14706_), .A2(new_n14079_), .B1(\asqrt[16] ), .B2(new_n14707_), .ZN(new_n14708_));
  INV_X1     g14516(.I(new_n14708_), .ZN(new_n14709_));
  NAND2_X1   g14517(.A1(new_n14694_), .A2(new_n8036_), .ZN(new_n14710_));
  OAI21_X1   g14518(.A1(new_n14710_), .A2(new_n14702_), .B(new_n14709_), .ZN(new_n14711_));
  AOI21_X1   g14519(.A1(new_n14711_), .A2(new_n14703_), .B(new_n7539_), .ZN(new_n14712_));
  INV_X1     g14520(.I(new_n14712_), .ZN(new_n14713_));
  INV_X1     g14521(.I(new_n14711_), .ZN(new_n14714_));
  INV_X1     g14522(.I(new_n14086_), .ZN(new_n14715_));
  NOR3_X1    g14523(.A1(new_n14082_), .A2(new_n14455_), .A3(new_n14715_), .ZN(new_n14716_));
  NOR3_X1    g14524(.A1(new_n14601_), .A2(new_n14082_), .A3(new_n14455_), .ZN(new_n14717_));
  INV_X1     g14525(.I(new_n14717_), .ZN(new_n14718_));
  AOI22_X1   g14526(.A1(new_n14718_), .A2(new_n14715_), .B1(\asqrt[16] ), .B2(new_n14716_), .ZN(new_n14719_));
  INV_X1     g14527(.I(new_n14719_), .ZN(new_n14720_));
  NAND2_X1   g14528(.A1(new_n14703_), .A2(new_n7539_), .ZN(new_n14721_));
  OAI21_X1   g14529(.A1(new_n14721_), .A2(new_n14714_), .B(new_n14720_), .ZN(new_n14722_));
  AOI21_X1   g14530(.A1(new_n14722_), .A2(new_n14713_), .B(new_n7229_), .ZN(new_n14723_));
  NOR3_X1    g14531(.A1(new_n14601_), .A2(new_n14091_), .A3(new_n14097_), .ZN(new_n14724_));
  INV_X1     g14532(.I(new_n14724_), .ZN(new_n14725_));
  NOR3_X1    g14533(.A1(new_n14091_), .A2(new_n14409_), .A3(new_n14097_), .ZN(new_n14726_));
  AOI22_X1   g14534(.A1(new_n14725_), .A2(new_n14409_), .B1(\asqrt[16] ), .B2(new_n14726_), .ZN(new_n14727_));
  NOR2_X1    g14535(.A1(new_n14712_), .A2(\asqrt[31] ), .ZN(new_n14728_));
  AOI21_X1   g14536(.A1(new_n14728_), .A2(new_n14722_), .B(new_n14727_), .ZN(new_n14729_));
  OAI21_X1   g14537(.A1(new_n14729_), .A2(new_n14723_), .B(\asqrt[32] ), .ZN(new_n14730_));
  NOR2_X1    g14538(.A1(new_n14098_), .A2(new_n14106_), .ZN(new_n14731_));
  NOR3_X1    g14539(.A1(new_n14731_), .A2(new_n14454_), .A3(new_n14105_), .ZN(new_n14732_));
  NOR3_X1    g14540(.A1(new_n14601_), .A2(new_n14454_), .A3(new_n14731_), .ZN(new_n14733_));
  INV_X1     g14541(.I(new_n14733_), .ZN(new_n14734_));
  AOI22_X1   g14542(.A1(new_n14734_), .A2(new_n14105_), .B1(\asqrt[16] ), .B2(new_n14732_), .ZN(new_n14735_));
  INV_X1     g14543(.I(new_n14735_), .ZN(new_n14736_));
  NOR3_X1    g14544(.A1(new_n14693_), .A2(new_n14680_), .A3(\asqrt[28] ), .ZN(new_n14737_));
  OAI21_X1   g14545(.A1(new_n14700_), .A2(new_n14737_), .B(new_n14694_), .ZN(new_n14738_));
  AOI21_X1   g14546(.A1(new_n14738_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n14739_));
  AOI21_X1   g14547(.A1(new_n14739_), .A2(new_n14711_), .B(new_n14719_), .ZN(new_n14740_));
  OAI21_X1   g14548(.A1(new_n14740_), .A2(new_n14712_), .B(\asqrt[31] ), .ZN(new_n14741_));
  NAND2_X1   g14549(.A1(new_n14741_), .A2(new_n6824_), .ZN(new_n14742_));
  OAI21_X1   g14550(.A1(new_n14742_), .A2(new_n14729_), .B(new_n14736_), .ZN(new_n14743_));
  AOI21_X1   g14551(.A1(new_n14743_), .A2(new_n14730_), .B(new_n6356_), .ZN(new_n14744_));
  INV_X1     g14552(.I(new_n14744_), .ZN(new_n14745_));
  INV_X1     g14553(.I(new_n14743_), .ZN(new_n14746_));
  INV_X1     g14554(.I(new_n14112_), .ZN(new_n14747_));
  NOR3_X1    g14555(.A1(new_n14601_), .A2(new_n14108_), .A3(new_n14463_), .ZN(new_n14748_));
  INV_X1     g14556(.I(new_n14748_), .ZN(new_n14749_));
  NOR3_X1    g14557(.A1(new_n14108_), .A2(new_n14463_), .A3(new_n14747_), .ZN(new_n14750_));
  AOI22_X1   g14558(.A1(new_n14749_), .A2(new_n14747_), .B1(\asqrt[16] ), .B2(new_n14750_), .ZN(new_n14751_));
  INV_X1     g14559(.I(new_n14751_), .ZN(new_n14752_));
  NAND2_X1   g14560(.A1(new_n14730_), .A2(new_n6356_), .ZN(new_n14753_));
  OAI21_X1   g14561(.A1(new_n14753_), .A2(new_n14746_), .B(new_n14752_), .ZN(new_n14754_));
  AOI21_X1   g14562(.A1(new_n14754_), .A2(new_n14745_), .B(new_n6077_), .ZN(new_n14755_));
  NOR3_X1    g14563(.A1(new_n14117_), .A2(new_n14408_), .A3(new_n14123_), .ZN(new_n14756_));
  NOR3_X1    g14564(.A1(new_n14601_), .A2(new_n14117_), .A3(new_n14123_), .ZN(new_n14757_));
  INV_X1     g14565(.I(new_n14757_), .ZN(new_n14758_));
  AOI22_X1   g14566(.A1(new_n14758_), .A2(new_n14408_), .B1(\asqrt[16] ), .B2(new_n14756_), .ZN(new_n14759_));
  NOR2_X1    g14567(.A1(new_n14744_), .A2(\asqrt[34] ), .ZN(new_n14760_));
  AOI21_X1   g14568(.A1(new_n14760_), .A2(new_n14754_), .B(new_n14759_), .ZN(new_n14761_));
  OAI21_X1   g14569(.A1(new_n14761_), .A2(new_n14755_), .B(\asqrt[35] ), .ZN(new_n14762_));
  NOR2_X1    g14570(.A1(new_n14124_), .A2(new_n14132_), .ZN(new_n14763_));
  NOR3_X1    g14571(.A1(new_n14601_), .A2(new_n14462_), .A3(new_n14763_), .ZN(new_n14764_));
  INV_X1     g14572(.I(new_n14764_), .ZN(new_n14765_));
  NOR3_X1    g14573(.A1(new_n14763_), .A2(new_n14462_), .A3(new_n14131_), .ZN(new_n14766_));
  AOI22_X1   g14574(.A1(new_n14765_), .A2(new_n14131_), .B1(\asqrt[16] ), .B2(new_n14766_), .ZN(new_n14767_));
  INV_X1     g14575(.I(new_n14767_), .ZN(new_n14768_));
  NOR3_X1    g14576(.A1(new_n14740_), .A2(\asqrt[31] ), .A3(new_n14712_), .ZN(new_n14769_));
  OAI21_X1   g14577(.A1(new_n14727_), .A2(new_n14769_), .B(new_n14741_), .ZN(new_n14770_));
  AOI21_X1   g14578(.A1(new_n14770_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n14771_));
  AOI21_X1   g14579(.A1(new_n14771_), .A2(new_n14743_), .B(new_n14751_), .ZN(new_n14772_));
  OAI21_X1   g14580(.A1(new_n14772_), .A2(new_n14744_), .B(\asqrt[34] ), .ZN(new_n14773_));
  NAND2_X1   g14581(.A1(new_n14773_), .A2(new_n5708_), .ZN(new_n14774_));
  OAI21_X1   g14582(.A1(new_n14774_), .A2(new_n14761_), .B(new_n14768_), .ZN(new_n14775_));
  NAND2_X1   g14583(.A1(new_n14775_), .A2(new_n14762_), .ZN(new_n14776_));
  NAND2_X1   g14584(.A1(new_n14776_), .A2(\asqrt[36] ), .ZN(new_n14777_));
  INV_X1     g14585(.I(new_n14775_), .ZN(new_n14778_));
  INV_X1     g14586(.I(new_n14138_), .ZN(new_n14779_));
  NOR3_X1    g14587(.A1(new_n14134_), .A2(new_n14471_), .A3(new_n14779_), .ZN(new_n14780_));
  NOR3_X1    g14588(.A1(new_n14601_), .A2(new_n14134_), .A3(new_n14471_), .ZN(new_n14781_));
  INV_X1     g14589(.I(new_n14781_), .ZN(new_n14782_));
  AOI22_X1   g14590(.A1(new_n14782_), .A2(new_n14779_), .B1(\asqrt[16] ), .B2(new_n14780_), .ZN(new_n14783_));
  INV_X1     g14591(.I(new_n14783_), .ZN(new_n14784_));
  NAND2_X1   g14592(.A1(new_n14762_), .A2(new_n5277_), .ZN(new_n14785_));
  OAI21_X1   g14593(.A1(new_n14778_), .A2(new_n14785_), .B(new_n14784_), .ZN(new_n14786_));
  AOI21_X1   g14594(.A1(new_n14786_), .A2(new_n14777_), .B(new_n5024_), .ZN(new_n14787_));
  NOR3_X1    g14595(.A1(new_n14601_), .A2(new_n14143_), .A3(new_n14149_), .ZN(new_n14788_));
  INV_X1     g14596(.I(new_n14788_), .ZN(new_n14789_));
  NOR3_X1    g14597(.A1(new_n14143_), .A2(new_n14407_), .A3(new_n14149_), .ZN(new_n14790_));
  AOI22_X1   g14598(.A1(new_n14789_), .A2(new_n14407_), .B1(\asqrt[16] ), .B2(new_n14790_), .ZN(new_n14791_));
  AOI21_X1   g14599(.A1(new_n14775_), .A2(new_n14762_), .B(new_n5277_), .ZN(new_n14792_));
  NOR2_X1    g14600(.A1(new_n14792_), .A2(\asqrt[37] ), .ZN(new_n14793_));
  AOI21_X1   g14601(.A1(new_n14793_), .A2(new_n14786_), .B(new_n14791_), .ZN(new_n14794_));
  OAI21_X1   g14602(.A1(new_n14794_), .A2(new_n14787_), .B(\asqrt[38] ), .ZN(new_n14795_));
  INV_X1     g14603(.I(new_n14795_), .ZN(new_n14796_));
  NOR2_X1    g14604(.A1(new_n14150_), .A2(new_n14158_), .ZN(new_n14797_));
  NOR3_X1    g14605(.A1(new_n14797_), .A2(new_n14470_), .A3(new_n14157_), .ZN(new_n14798_));
  NOR3_X1    g14606(.A1(new_n14601_), .A2(new_n14470_), .A3(new_n14797_), .ZN(new_n14799_));
  INV_X1     g14607(.I(new_n14799_), .ZN(new_n14800_));
  AOI22_X1   g14608(.A1(new_n14800_), .A2(new_n14157_), .B1(\asqrt[16] ), .B2(new_n14798_), .ZN(new_n14801_));
  NOR3_X1    g14609(.A1(new_n14794_), .A2(new_n14787_), .A3(\asqrt[38] ), .ZN(new_n14802_));
  NOR2_X1    g14610(.A1(new_n14802_), .A2(new_n14801_), .ZN(new_n14803_));
  OAI21_X1   g14611(.A1(new_n14803_), .A2(new_n14796_), .B(\asqrt[39] ), .ZN(new_n14804_));
  INV_X1     g14612(.I(new_n14164_), .ZN(new_n14805_));
  NOR3_X1    g14613(.A1(new_n14601_), .A2(new_n14160_), .A3(new_n14479_), .ZN(new_n14806_));
  INV_X1     g14614(.I(new_n14806_), .ZN(new_n14807_));
  NOR3_X1    g14615(.A1(new_n14160_), .A2(new_n14479_), .A3(new_n14805_), .ZN(new_n14808_));
  AOI22_X1   g14616(.A1(new_n14807_), .A2(new_n14805_), .B1(\asqrt[16] ), .B2(new_n14808_), .ZN(new_n14809_));
  INV_X1     g14617(.I(new_n14809_), .ZN(new_n14810_));
  NAND2_X1   g14618(.A1(new_n14795_), .A2(new_n4298_), .ZN(new_n14811_));
  OAI21_X1   g14619(.A1(new_n14803_), .A2(new_n14811_), .B(new_n14810_), .ZN(new_n14812_));
  AOI21_X1   g14620(.A1(new_n14812_), .A2(new_n14804_), .B(new_n4071_), .ZN(new_n14813_));
  NOR3_X1    g14621(.A1(new_n14169_), .A2(new_n14406_), .A3(new_n14175_), .ZN(new_n14814_));
  NOR3_X1    g14622(.A1(new_n14601_), .A2(new_n14169_), .A3(new_n14175_), .ZN(new_n14815_));
  INV_X1     g14623(.I(new_n14815_), .ZN(new_n14816_));
  AOI22_X1   g14624(.A1(new_n14816_), .A2(new_n14406_), .B1(\asqrt[16] ), .B2(new_n14814_), .ZN(new_n14817_));
  INV_X1     g14625(.I(new_n14801_), .ZN(new_n14818_));
  NOR3_X1    g14626(.A1(new_n14772_), .A2(\asqrt[34] ), .A3(new_n14744_), .ZN(new_n14819_));
  OAI21_X1   g14627(.A1(new_n14759_), .A2(new_n14819_), .B(new_n14773_), .ZN(new_n14820_));
  AOI21_X1   g14628(.A1(new_n14820_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n14821_));
  AOI21_X1   g14629(.A1(new_n14821_), .A2(new_n14775_), .B(new_n14783_), .ZN(new_n14822_));
  OAI21_X1   g14630(.A1(new_n14822_), .A2(new_n14792_), .B(\asqrt[37] ), .ZN(new_n14823_));
  NAND2_X1   g14631(.A1(new_n14823_), .A2(new_n4696_), .ZN(new_n14824_));
  OAI21_X1   g14632(.A1(new_n14824_), .A2(new_n14794_), .B(new_n14818_), .ZN(new_n14825_));
  AOI21_X1   g14633(.A1(new_n14825_), .A2(new_n14795_), .B(new_n4298_), .ZN(new_n14826_));
  NOR2_X1    g14634(.A1(new_n14826_), .A2(\asqrt[40] ), .ZN(new_n14827_));
  AOI21_X1   g14635(.A1(new_n14827_), .A2(new_n14812_), .B(new_n14817_), .ZN(new_n14828_));
  OAI21_X1   g14636(.A1(new_n14828_), .A2(new_n14813_), .B(\asqrt[41] ), .ZN(new_n14829_));
  NOR2_X1    g14637(.A1(new_n14176_), .A2(new_n14184_), .ZN(new_n14830_));
  NOR3_X1    g14638(.A1(new_n14601_), .A2(new_n14478_), .A3(new_n14830_), .ZN(new_n14831_));
  INV_X1     g14639(.I(new_n14831_), .ZN(new_n14832_));
  NOR3_X1    g14640(.A1(new_n14830_), .A2(new_n14478_), .A3(new_n14183_), .ZN(new_n14833_));
  AOI22_X1   g14641(.A1(new_n14832_), .A2(new_n14183_), .B1(\asqrt[16] ), .B2(new_n14833_), .ZN(new_n14834_));
  INV_X1     g14642(.I(new_n14834_), .ZN(new_n14835_));
  NOR3_X1    g14643(.A1(new_n14822_), .A2(\asqrt[37] ), .A3(new_n14792_), .ZN(new_n14836_));
  OAI21_X1   g14644(.A1(new_n14791_), .A2(new_n14836_), .B(new_n14823_), .ZN(new_n14837_));
  AOI21_X1   g14645(.A1(new_n14837_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n14838_));
  AOI21_X1   g14646(.A1(new_n14838_), .A2(new_n14825_), .B(new_n14809_), .ZN(new_n14839_));
  OAI21_X1   g14647(.A1(new_n14839_), .A2(new_n14826_), .B(\asqrt[40] ), .ZN(new_n14840_));
  NAND2_X1   g14648(.A1(new_n14840_), .A2(new_n3782_), .ZN(new_n14841_));
  OAI21_X1   g14649(.A1(new_n14841_), .A2(new_n14828_), .B(new_n14835_), .ZN(new_n14842_));
  AOI21_X1   g14650(.A1(new_n14842_), .A2(new_n14829_), .B(new_n3419_), .ZN(new_n14843_));
  INV_X1     g14651(.I(new_n14190_), .ZN(new_n14844_));
  NOR3_X1    g14652(.A1(new_n14186_), .A2(new_n14487_), .A3(new_n14844_), .ZN(new_n14845_));
  NOR3_X1    g14653(.A1(new_n14601_), .A2(new_n14186_), .A3(new_n14487_), .ZN(new_n14846_));
  INV_X1     g14654(.I(new_n14846_), .ZN(new_n14847_));
  AOI22_X1   g14655(.A1(new_n14847_), .A2(new_n14844_), .B1(\asqrt[16] ), .B2(new_n14845_), .ZN(new_n14848_));
  NOR3_X1    g14656(.A1(new_n14839_), .A2(\asqrt[40] ), .A3(new_n14826_), .ZN(new_n14849_));
  OAI21_X1   g14657(.A1(new_n14817_), .A2(new_n14849_), .B(new_n14840_), .ZN(new_n14850_));
  AOI21_X1   g14658(.A1(new_n14850_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n14851_));
  AOI21_X1   g14659(.A1(new_n14851_), .A2(new_n14842_), .B(new_n14848_), .ZN(new_n14852_));
  OAI21_X1   g14660(.A1(new_n14852_), .A2(new_n14843_), .B(\asqrt[43] ), .ZN(new_n14853_));
  INV_X1     g14661(.I(new_n14853_), .ZN(new_n14854_));
  NOR3_X1    g14662(.A1(new_n14601_), .A2(new_n14195_), .A3(new_n14201_), .ZN(new_n14855_));
  INV_X1     g14663(.I(new_n14855_), .ZN(new_n14856_));
  NOR3_X1    g14664(.A1(new_n14195_), .A2(new_n14405_), .A3(new_n14201_), .ZN(new_n14857_));
  AOI22_X1   g14665(.A1(new_n14856_), .A2(new_n14405_), .B1(\asqrt[16] ), .B2(new_n14857_), .ZN(new_n14858_));
  NOR3_X1    g14666(.A1(new_n14852_), .A2(\asqrt[43] ), .A3(new_n14843_), .ZN(new_n14859_));
  NOR2_X1    g14667(.A1(new_n14859_), .A2(new_n14858_), .ZN(new_n14860_));
  OAI21_X1   g14668(.A1(new_n14860_), .A2(new_n14854_), .B(\asqrt[44] ), .ZN(new_n14861_));
  NOR2_X1    g14669(.A1(new_n14202_), .A2(new_n14210_), .ZN(new_n14862_));
  NOR3_X1    g14670(.A1(new_n14862_), .A2(new_n14486_), .A3(new_n14209_), .ZN(new_n14863_));
  NOR3_X1    g14671(.A1(new_n14601_), .A2(new_n14486_), .A3(new_n14862_), .ZN(new_n14864_));
  INV_X1     g14672(.I(new_n14864_), .ZN(new_n14865_));
  AOI22_X1   g14673(.A1(new_n14865_), .A2(new_n14209_), .B1(\asqrt[16] ), .B2(new_n14863_), .ZN(new_n14866_));
  INV_X1     g14674(.I(new_n14866_), .ZN(new_n14867_));
  NAND2_X1   g14675(.A1(new_n14853_), .A2(new_n2954_), .ZN(new_n14868_));
  OAI21_X1   g14676(.A1(new_n14860_), .A2(new_n14868_), .B(new_n14867_), .ZN(new_n14869_));
  AOI21_X1   g14677(.A1(new_n14869_), .A2(new_n14861_), .B(new_n2641_), .ZN(new_n14870_));
  INV_X1     g14678(.I(new_n14216_), .ZN(new_n14871_));
  NOR3_X1    g14679(.A1(new_n14601_), .A2(new_n14212_), .A3(new_n14495_), .ZN(new_n14872_));
  INV_X1     g14680(.I(new_n14872_), .ZN(new_n14873_));
  NOR3_X1    g14681(.A1(new_n14212_), .A2(new_n14495_), .A3(new_n14871_), .ZN(new_n14874_));
  AOI22_X1   g14682(.A1(new_n14873_), .A2(new_n14871_), .B1(\asqrt[16] ), .B2(new_n14874_), .ZN(new_n14875_));
  OAI21_X1   g14683(.A1(new_n14858_), .A2(new_n14859_), .B(new_n14853_), .ZN(new_n14876_));
  AOI21_X1   g14684(.A1(new_n14876_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n14877_));
  AOI21_X1   g14685(.A1(new_n14877_), .A2(new_n14869_), .B(new_n14875_), .ZN(new_n14878_));
  OAI21_X1   g14686(.A1(new_n14878_), .A2(new_n14870_), .B(\asqrt[46] ), .ZN(new_n14879_));
  INV_X1     g14687(.I(new_n14879_), .ZN(new_n14880_));
  NOR3_X1    g14688(.A1(new_n14221_), .A2(new_n14404_), .A3(new_n14227_), .ZN(new_n14881_));
  NOR3_X1    g14689(.A1(new_n14601_), .A2(new_n14221_), .A3(new_n14227_), .ZN(new_n14882_));
  INV_X1     g14690(.I(new_n14882_), .ZN(new_n14883_));
  AOI22_X1   g14691(.A1(new_n14883_), .A2(new_n14404_), .B1(\asqrt[16] ), .B2(new_n14881_), .ZN(new_n14884_));
  NOR3_X1    g14692(.A1(new_n14878_), .A2(new_n14870_), .A3(\asqrt[46] ), .ZN(new_n14885_));
  NOR2_X1    g14693(.A1(new_n14885_), .A2(new_n14884_), .ZN(new_n14886_));
  OAI21_X1   g14694(.A1(new_n14886_), .A2(new_n14880_), .B(\asqrt[47] ), .ZN(new_n14887_));
  NOR2_X1    g14695(.A1(new_n14228_), .A2(new_n14236_), .ZN(new_n14888_));
  NOR3_X1    g14696(.A1(new_n14601_), .A2(new_n14494_), .A3(new_n14888_), .ZN(new_n14889_));
  INV_X1     g14697(.I(new_n14889_), .ZN(new_n14890_));
  NOR3_X1    g14698(.A1(new_n14888_), .A2(new_n14494_), .A3(new_n14235_), .ZN(new_n14891_));
  AOI22_X1   g14699(.A1(new_n14890_), .A2(new_n14235_), .B1(\asqrt[16] ), .B2(new_n14891_), .ZN(new_n14892_));
  INV_X1     g14700(.I(new_n14892_), .ZN(new_n14893_));
  NAND2_X1   g14701(.A1(new_n14879_), .A2(new_n2229_), .ZN(new_n14894_));
  OAI21_X1   g14702(.A1(new_n14886_), .A2(new_n14894_), .B(new_n14893_), .ZN(new_n14895_));
  AOI21_X1   g14703(.A1(new_n14895_), .A2(new_n14887_), .B(new_n1956_), .ZN(new_n14896_));
  INV_X1     g14704(.I(new_n14242_), .ZN(new_n14897_));
  NOR3_X1    g14705(.A1(new_n14238_), .A2(new_n14503_), .A3(new_n14897_), .ZN(new_n14898_));
  NOR3_X1    g14706(.A1(new_n14601_), .A2(new_n14238_), .A3(new_n14503_), .ZN(new_n14899_));
  INV_X1     g14707(.I(new_n14899_), .ZN(new_n14900_));
  AOI22_X1   g14708(.A1(new_n14900_), .A2(new_n14897_), .B1(\asqrt[16] ), .B2(new_n14898_), .ZN(new_n14901_));
  OAI21_X1   g14709(.A1(new_n14884_), .A2(new_n14885_), .B(new_n14879_), .ZN(new_n14902_));
  AOI21_X1   g14710(.A1(new_n14902_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n14903_));
  AOI21_X1   g14711(.A1(new_n14903_), .A2(new_n14895_), .B(new_n14901_), .ZN(new_n14904_));
  OAI21_X1   g14712(.A1(new_n14904_), .A2(new_n14896_), .B(\asqrt[49] ), .ZN(new_n14905_));
  INV_X1     g14713(.I(new_n14905_), .ZN(new_n14906_));
  NOR3_X1    g14714(.A1(new_n14601_), .A2(new_n14247_), .A3(new_n14253_), .ZN(new_n14907_));
  INV_X1     g14715(.I(new_n14907_), .ZN(new_n14908_));
  NOR3_X1    g14716(.A1(new_n14247_), .A2(new_n14403_), .A3(new_n14253_), .ZN(new_n14909_));
  AOI22_X1   g14717(.A1(new_n14908_), .A2(new_n14403_), .B1(\asqrt[16] ), .B2(new_n14909_), .ZN(new_n14910_));
  NOR3_X1    g14718(.A1(new_n14904_), .A2(new_n14896_), .A3(\asqrt[49] ), .ZN(new_n14911_));
  NOR2_X1    g14719(.A1(new_n14911_), .A2(new_n14910_), .ZN(new_n14912_));
  OAI21_X1   g14720(.A1(new_n14912_), .A2(new_n14906_), .B(\asqrt[50] ), .ZN(new_n14913_));
  NOR2_X1    g14721(.A1(new_n14254_), .A2(new_n14262_), .ZN(new_n14914_));
  NOR3_X1    g14722(.A1(new_n14914_), .A2(new_n14502_), .A3(new_n14261_), .ZN(new_n14915_));
  NOR3_X1    g14723(.A1(new_n14601_), .A2(new_n14502_), .A3(new_n14914_), .ZN(new_n14916_));
  INV_X1     g14724(.I(new_n14916_), .ZN(new_n14917_));
  AOI22_X1   g14725(.A1(new_n14917_), .A2(new_n14261_), .B1(\asqrt[16] ), .B2(new_n14915_), .ZN(new_n14918_));
  INV_X1     g14726(.I(new_n14918_), .ZN(new_n14919_));
  NAND2_X1   g14727(.A1(new_n14905_), .A2(new_n1612_), .ZN(new_n14920_));
  OAI21_X1   g14728(.A1(new_n14912_), .A2(new_n14920_), .B(new_n14919_), .ZN(new_n14921_));
  AOI21_X1   g14729(.A1(new_n14921_), .A2(new_n14913_), .B(new_n1376_), .ZN(new_n14922_));
  INV_X1     g14730(.I(new_n14268_), .ZN(new_n14923_));
  NOR3_X1    g14731(.A1(new_n14601_), .A2(new_n14264_), .A3(new_n14511_), .ZN(new_n14924_));
  INV_X1     g14732(.I(new_n14924_), .ZN(new_n14925_));
  NOR3_X1    g14733(.A1(new_n14264_), .A2(new_n14511_), .A3(new_n14923_), .ZN(new_n14926_));
  AOI22_X1   g14734(.A1(new_n14925_), .A2(new_n14923_), .B1(\asqrt[16] ), .B2(new_n14926_), .ZN(new_n14927_));
  OAI21_X1   g14735(.A1(new_n14910_), .A2(new_n14911_), .B(new_n14905_), .ZN(new_n14928_));
  AOI21_X1   g14736(.A1(new_n14928_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n14929_));
  AOI21_X1   g14737(.A1(new_n14929_), .A2(new_n14921_), .B(new_n14927_), .ZN(new_n14930_));
  OAI21_X1   g14738(.A1(new_n14930_), .A2(new_n14922_), .B(\asqrt[52] ), .ZN(new_n14931_));
  INV_X1     g14739(.I(new_n14931_), .ZN(new_n14932_));
  INV_X1     g14740(.I(new_n14930_), .ZN(new_n14933_));
  NOR3_X1    g14741(.A1(new_n14273_), .A2(new_n14402_), .A3(new_n14279_), .ZN(new_n14934_));
  NOR3_X1    g14742(.A1(new_n14601_), .A2(new_n14273_), .A3(new_n14279_), .ZN(new_n14935_));
  INV_X1     g14743(.I(new_n14935_), .ZN(new_n14936_));
  AOI22_X1   g14744(.A1(new_n14936_), .A2(new_n14402_), .B1(\asqrt[16] ), .B2(new_n14934_), .ZN(new_n14937_));
  NOR2_X1    g14745(.A1(new_n14922_), .A2(\asqrt[52] ), .ZN(new_n14938_));
  AOI21_X1   g14746(.A1(new_n14933_), .A2(new_n14938_), .B(new_n14937_), .ZN(new_n14939_));
  OAI21_X1   g14747(.A1(new_n14939_), .A2(new_n14932_), .B(\asqrt[53] ), .ZN(new_n14940_));
  NOR2_X1    g14748(.A1(new_n14280_), .A2(new_n14290_), .ZN(new_n14941_));
  NOR3_X1    g14749(.A1(new_n14601_), .A2(new_n14510_), .A3(new_n14941_), .ZN(new_n14942_));
  INV_X1     g14750(.I(new_n14942_), .ZN(new_n14943_));
  NOR3_X1    g14751(.A1(new_n14941_), .A2(new_n14510_), .A3(new_n14289_), .ZN(new_n14944_));
  AOI22_X1   g14752(.A1(new_n14943_), .A2(new_n14289_), .B1(\asqrt[16] ), .B2(new_n14944_), .ZN(new_n14945_));
  INV_X1     g14753(.I(new_n14945_), .ZN(new_n14946_));
  NAND2_X1   g14754(.A1(new_n14931_), .A2(new_n1103_), .ZN(new_n14947_));
  OAI21_X1   g14755(.A1(new_n14947_), .A2(new_n14939_), .B(new_n14946_), .ZN(new_n14948_));
  AOI21_X1   g14756(.A1(new_n14948_), .A2(new_n14940_), .B(new_n904_), .ZN(new_n14949_));
  INV_X1     g14757(.I(new_n14949_), .ZN(new_n14950_));
  INV_X1     g14758(.I(new_n14948_), .ZN(new_n14951_));
  INV_X1     g14759(.I(new_n14296_), .ZN(new_n14952_));
  NOR3_X1    g14760(.A1(new_n14292_), .A2(new_n14519_), .A3(new_n14952_), .ZN(new_n14953_));
  NOR3_X1    g14761(.A1(new_n14601_), .A2(new_n14292_), .A3(new_n14519_), .ZN(new_n14954_));
  INV_X1     g14762(.I(new_n14954_), .ZN(new_n14955_));
  AOI22_X1   g14763(.A1(new_n14955_), .A2(new_n14952_), .B1(\asqrt[16] ), .B2(new_n14953_), .ZN(new_n14956_));
  INV_X1     g14764(.I(new_n14956_), .ZN(new_n14957_));
  NAND2_X1   g14765(.A1(new_n14940_), .A2(new_n904_), .ZN(new_n14958_));
  OAI21_X1   g14766(.A1(new_n14958_), .A2(new_n14951_), .B(new_n14957_), .ZN(new_n14959_));
  AOI21_X1   g14767(.A1(new_n14959_), .A2(new_n14950_), .B(new_n823_), .ZN(new_n14960_));
  NOR3_X1    g14768(.A1(new_n14601_), .A2(new_n14301_), .A3(new_n14308_), .ZN(new_n14961_));
  INV_X1     g14769(.I(new_n14961_), .ZN(new_n14962_));
  NOR3_X1    g14770(.A1(new_n14301_), .A2(new_n14401_), .A3(new_n14308_), .ZN(new_n14963_));
  AOI22_X1   g14771(.A1(new_n14962_), .A2(new_n14401_), .B1(\asqrt[16] ), .B2(new_n14963_), .ZN(new_n14964_));
  NOR2_X1    g14772(.A1(new_n14949_), .A2(\asqrt[55] ), .ZN(new_n14965_));
  AOI21_X1   g14773(.A1(new_n14965_), .A2(new_n14959_), .B(new_n14964_), .ZN(new_n14966_));
  OAI21_X1   g14774(.A1(new_n14966_), .A2(new_n14960_), .B(\asqrt[56] ), .ZN(new_n14967_));
  NOR2_X1    g14775(.A1(new_n14309_), .A2(new_n14321_), .ZN(new_n14968_));
  NOR3_X1    g14776(.A1(new_n14968_), .A2(new_n14518_), .A3(new_n14320_), .ZN(new_n14969_));
  NOR3_X1    g14777(.A1(new_n14601_), .A2(new_n14518_), .A3(new_n14968_), .ZN(new_n14970_));
  INV_X1     g14778(.I(new_n14970_), .ZN(new_n14971_));
  AOI22_X1   g14779(.A1(new_n14971_), .A2(new_n14320_), .B1(\asqrt[16] ), .B2(new_n14969_), .ZN(new_n14972_));
  INV_X1     g14780(.I(new_n14972_), .ZN(new_n14973_));
  NOR3_X1    g14781(.A1(new_n14930_), .A2(new_n14922_), .A3(\asqrt[52] ), .ZN(new_n14974_));
  OAI21_X1   g14782(.A1(new_n14937_), .A2(new_n14974_), .B(new_n14931_), .ZN(new_n14975_));
  AOI21_X1   g14783(.A1(new_n14975_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n14976_));
  AOI21_X1   g14784(.A1(new_n14976_), .A2(new_n14948_), .B(new_n14956_), .ZN(new_n14977_));
  OAI21_X1   g14785(.A1(new_n14977_), .A2(new_n14949_), .B(\asqrt[55] ), .ZN(new_n14978_));
  NAND2_X1   g14786(.A1(new_n14978_), .A2(new_n703_), .ZN(new_n14979_));
  OAI21_X1   g14787(.A1(new_n14979_), .A2(new_n14966_), .B(new_n14973_), .ZN(new_n14980_));
  AOI21_X1   g14788(.A1(new_n14980_), .A2(new_n14967_), .B(new_n531_), .ZN(new_n14981_));
  INV_X1     g14789(.I(new_n14981_), .ZN(new_n14982_));
  INV_X1     g14790(.I(new_n14980_), .ZN(new_n14983_));
  INV_X1     g14791(.I(new_n14327_), .ZN(new_n14984_));
  NOR3_X1    g14792(.A1(new_n14601_), .A2(new_n14323_), .A3(new_n14527_), .ZN(new_n14985_));
  INV_X1     g14793(.I(new_n14985_), .ZN(new_n14986_));
  NOR3_X1    g14794(.A1(new_n14323_), .A2(new_n14527_), .A3(new_n14984_), .ZN(new_n14987_));
  AOI22_X1   g14795(.A1(new_n14986_), .A2(new_n14984_), .B1(\asqrt[16] ), .B2(new_n14987_), .ZN(new_n14988_));
  INV_X1     g14796(.I(new_n14988_), .ZN(new_n14989_));
  NAND2_X1   g14797(.A1(new_n14967_), .A2(new_n531_), .ZN(new_n14990_));
  OAI21_X1   g14798(.A1(new_n14990_), .A2(new_n14983_), .B(new_n14989_), .ZN(new_n14991_));
  AOI21_X1   g14799(.A1(new_n14991_), .A2(new_n14982_), .B(new_n436_), .ZN(new_n14992_));
  NOR3_X1    g14800(.A1(new_n14332_), .A2(new_n14400_), .A3(new_n14339_), .ZN(new_n14993_));
  NOR3_X1    g14801(.A1(new_n14601_), .A2(new_n14332_), .A3(new_n14339_), .ZN(new_n14994_));
  INV_X1     g14802(.I(new_n14994_), .ZN(new_n14995_));
  AOI22_X1   g14803(.A1(new_n14995_), .A2(new_n14400_), .B1(\asqrt[16] ), .B2(new_n14993_), .ZN(new_n14996_));
  NOR2_X1    g14804(.A1(new_n14981_), .A2(\asqrt[58] ), .ZN(new_n14997_));
  AOI21_X1   g14805(.A1(new_n14997_), .A2(new_n14991_), .B(new_n14996_), .ZN(new_n14998_));
  OAI21_X1   g14806(.A1(new_n14998_), .A2(new_n14992_), .B(\asqrt[59] ), .ZN(new_n14999_));
  NOR2_X1    g14807(.A1(new_n14340_), .A2(new_n14351_), .ZN(new_n15000_));
  NOR3_X1    g14808(.A1(new_n14601_), .A2(new_n14526_), .A3(new_n15000_), .ZN(new_n15001_));
  INV_X1     g14809(.I(new_n15001_), .ZN(new_n15002_));
  NOR3_X1    g14810(.A1(new_n15000_), .A2(new_n14526_), .A3(new_n14350_), .ZN(new_n15003_));
  AOI22_X1   g14811(.A1(new_n15002_), .A2(new_n14350_), .B1(\asqrt[16] ), .B2(new_n15003_), .ZN(new_n15004_));
  INV_X1     g14812(.I(new_n15004_), .ZN(new_n15005_));
  NOR3_X1    g14813(.A1(new_n14977_), .A2(\asqrt[55] ), .A3(new_n14949_), .ZN(new_n15006_));
  OAI21_X1   g14814(.A1(new_n14964_), .A2(new_n15006_), .B(new_n14978_), .ZN(new_n15007_));
  AOI21_X1   g14815(.A1(new_n15007_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n15008_));
  AOI21_X1   g14816(.A1(new_n15008_), .A2(new_n14980_), .B(new_n14988_), .ZN(new_n15009_));
  OAI21_X1   g14817(.A1(new_n15009_), .A2(new_n14981_), .B(\asqrt[58] ), .ZN(new_n15010_));
  NAND2_X1   g14818(.A1(new_n15010_), .A2(new_n327_), .ZN(new_n15011_));
  OAI21_X1   g14819(.A1(new_n15011_), .A2(new_n14998_), .B(new_n15005_), .ZN(new_n15012_));
  AOI21_X1   g14820(.A1(new_n15012_), .A2(new_n14999_), .B(new_n306_), .ZN(new_n15013_));
  INV_X1     g14821(.I(new_n15013_), .ZN(new_n15014_));
  INV_X1     g14822(.I(new_n15012_), .ZN(new_n15015_));
  INV_X1     g14823(.I(new_n14357_), .ZN(new_n15016_));
  NOR3_X1    g14824(.A1(new_n14353_), .A2(new_n14534_), .A3(new_n15016_), .ZN(new_n15017_));
  NOR3_X1    g14825(.A1(new_n14601_), .A2(new_n14353_), .A3(new_n14534_), .ZN(new_n15018_));
  INV_X1     g14826(.I(new_n15018_), .ZN(new_n15019_));
  AOI22_X1   g14827(.A1(new_n15019_), .A2(new_n15016_), .B1(\asqrt[16] ), .B2(new_n15017_), .ZN(new_n15020_));
  INV_X1     g14828(.I(new_n15020_), .ZN(new_n15021_));
  NAND2_X1   g14829(.A1(new_n14999_), .A2(new_n306_), .ZN(new_n15022_));
  OAI21_X1   g14830(.A1(new_n15015_), .A2(new_n15022_), .B(new_n15021_), .ZN(new_n15023_));
  AOI21_X1   g14831(.A1(new_n15023_), .A2(new_n15014_), .B(new_n218_), .ZN(new_n15024_));
  NOR3_X1    g14832(.A1(new_n14601_), .A2(new_n14362_), .A3(new_n14368_), .ZN(new_n15025_));
  INV_X1     g14833(.I(new_n15025_), .ZN(new_n15026_));
  NOR3_X1    g14834(.A1(new_n14362_), .A2(new_n14399_), .A3(new_n14368_), .ZN(new_n15027_));
  AOI22_X1   g14835(.A1(new_n15026_), .A2(new_n14399_), .B1(\asqrt[16] ), .B2(new_n15027_), .ZN(new_n15028_));
  NOR2_X1    g14836(.A1(new_n15013_), .A2(\asqrt[61] ), .ZN(new_n15029_));
  AOI21_X1   g14837(.A1(new_n15029_), .A2(new_n15023_), .B(new_n15028_), .ZN(new_n15030_));
  OAI21_X1   g14838(.A1(new_n15030_), .A2(new_n15024_), .B(\asqrt[62] ), .ZN(new_n15031_));
  NOR2_X1    g14839(.A1(new_n14369_), .A2(new_n14376_), .ZN(new_n15032_));
  NOR3_X1    g14840(.A1(new_n15032_), .A2(new_n14556_), .A3(new_n14375_), .ZN(new_n15033_));
  NOR3_X1    g14841(.A1(new_n14601_), .A2(new_n14556_), .A3(new_n15032_), .ZN(new_n15034_));
  INV_X1     g14842(.I(new_n15034_), .ZN(new_n15035_));
  AOI22_X1   g14843(.A1(new_n15035_), .A2(new_n14375_), .B1(\asqrt[16] ), .B2(new_n15033_), .ZN(new_n15036_));
  INV_X1     g14844(.I(new_n15036_), .ZN(new_n15037_));
  NOR3_X1    g14845(.A1(new_n15009_), .A2(\asqrt[58] ), .A3(new_n14981_), .ZN(new_n15038_));
  OAI21_X1   g14846(.A1(new_n14996_), .A2(new_n15038_), .B(new_n15010_), .ZN(new_n15039_));
  AOI21_X1   g14847(.A1(new_n15039_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n15040_));
  AOI21_X1   g14848(.A1(new_n15040_), .A2(new_n15012_), .B(new_n15020_), .ZN(new_n15041_));
  OAI21_X1   g14849(.A1(new_n15041_), .A2(new_n15013_), .B(\asqrt[61] ), .ZN(new_n15042_));
  NAND2_X1   g14850(.A1(new_n15042_), .A2(new_n207_), .ZN(new_n15043_));
  OAI21_X1   g14851(.A1(new_n15043_), .A2(new_n15030_), .B(new_n15037_), .ZN(new_n15044_));
  INV_X1     g14852(.I(new_n14558_), .ZN(new_n15045_));
  NAND4_X1   g14853(.A1(\asqrt[16] ), .A2(new_n14557_), .A3(new_n14382_), .A4(new_n15045_), .ZN(new_n15046_));
  NAND2_X1   g14854(.A1(new_n15045_), .A2(new_n14557_), .ZN(new_n15047_));
  OAI21_X1   g14855(.A1(new_n14601_), .A2(new_n15047_), .B(new_n14538_), .ZN(new_n15048_));
  NAND2_X1   g14856(.A1(new_n15048_), .A2(new_n15046_), .ZN(new_n15049_));
  INV_X1     g14857(.I(new_n14577_), .ZN(new_n15050_));
  AOI21_X1   g14858(.A1(new_n14540_), .A2(new_n14557_), .B(new_n14393_), .ZN(new_n15051_));
  AOI21_X1   g14859(.A1(\asqrt[16] ), .A2(new_n15051_), .B(new_n15050_), .ZN(new_n15052_));
  NAND2_X1   g14860(.A1(new_n15049_), .A2(new_n15052_), .ZN(new_n15053_));
  AOI21_X1   g14861(.A1(new_n15044_), .A2(new_n15031_), .B(new_n15053_), .ZN(new_n15054_));
  NOR2_X1    g14862(.A1(new_n15054_), .A2(\asqrt[63] ), .ZN(new_n15055_));
  INV_X1     g14863(.I(new_n15044_), .ZN(new_n15056_));
  INV_X1     g14864(.I(new_n15049_), .ZN(new_n15057_));
  NAND2_X1   g14865(.A1(new_n15031_), .A2(new_n15057_), .ZN(new_n15058_));
  AOI21_X1   g14866(.A1(\asqrt[16] ), .A2(new_n14394_), .B(new_n14559_), .ZN(new_n15059_));
  OR3_X2     g14867(.A1(new_n15059_), .A2(new_n193_), .A3(new_n15051_), .Z(new_n15060_));
  OAI21_X1   g14868(.A1(new_n13964_), .A2(new_n14546_), .B(new_n14389_), .ZN(new_n15061_));
  NOR4_X1    g14869(.A1(new_n15050_), .A2(new_n14392_), .A3(new_n14544_), .A4(new_n15061_), .ZN(new_n15062_));
  NAND2_X1   g14870(.A1(new_n15062_), .A2(new_n14398_), .ZN(new_n15063_));
  NAND2_X1   g14871(.A1(new_n15060_), .A2(new_n15063_), .ZN(new_n15064_));
  INV_X1     g14872(.I(new_n15064_), .ZN(new_n15065_));
  OAI21_X1   g14873(.A1(new_n15056_), .A2(new_n15058_), .B(new_n15065_), .ZN(new_n15066_));
  NOR2_X1    g14874(.A1(new_n15055_), .A2(new_n15066_), .ZN(new_n15067_));
  INV_X1     g14875(.I(\a[30] ), .ZN(new_n15068_));
  NOR2_X1    g14876(.A1(\a[28] ), .A2(\a[29] ), .ZN(new_n15069_));
  INV_X1     g14877(.I(new_n15069_), .ZN(new_n15070_));
  NOR2_X1    g14878(.A1(new_n15070_), .A2(\a[30] ), .ZN(new_n15071_));
  INV_X1     g14879(.I(new_n15071_), .ZN(new_n15072_));
  OAI21_X1   g14880(.A1(new_n15067_), .A2(new_n15068_), .B(new_n15072_), .ZN(new_n15073_));
  NOR3_X1    g14881(.A1(new_n14544_), .A2(new_n14547_), .A3(new_n15071_), .ZN(new_n15074_));
  NAND3_X1   g14882(.A1(new_n14398_), .A2(new_n14577_), .A3(new_n15074_), .ZN(new_n15075_));
  INV_X1     g14883(.I(new_n15075_), .ZN(new_n15076_));
  OAI21_X1   g14884(.A1(new_n15067_), .A2(new_n15068_), .B(new_n15076_), .ZN(new_n15077_));
  NOR3_X1    g14885(.A1(new_n15041_), .A2(\asqrt[61] ), .A3(new_n15013_), .ZN(new_n15078_));
  OAI21_X1   g14886(.A1(new_n15028_), .A2(new_n15078_), .B(new_n15042_), .ZN(new_n15079_));
  INV_X1     g14887(.I(new_n15028_), .ZN(new_n15080_));
  INV_X1     g14888(.I(new_n14996_), .ZN(new_n15081_));
  INV_X1     g14889(.I(new_n14964_), .ZN(new_n15082_));
  INV_X1     g14890(.I(new_n14937_), .ZN(new_n15083_));
  INV_X1     g14891(.I(new_n14910_), .ZN(new_n15084_));
  INV_X1     g14892(.I(new_n14884_), .ZN(new_n15085_));
  INV_X1     g14893(.I(new_n14858_), .ZN(new_n15086_));
  INV_X1     g14894(.I(new_n14829_), .ZN(new_n15087_));
  NOR3_X1    g14895(.A1(new_n14828_), .A2(new_n14813_), .A3(\asqrt[41] ), .ZN(new_n15088_));
  NOR2_X1    g14896(.A1(new_n15088_), .A2(new_n14834_), .ZN(new_n15089_));
  OAI21_X1   g14897(.A1(new_n15089_), .A2(new_n15087_), .B(\asqrt[42] ), .ZN(new_n15090_));
  NAND2_X1   g14898(.A1(new_n15090_), .A2(new_n3218_), .ZN(new_n15091_));
  OAI21_X1   g14899(.A1(new_n15091_), .A2(new_n14852_), .B(new_n15086_), .ZN(new_n15092_));
  NAND3_X1   g14900(.A1(new_n15092_), .A2(new_n2954_), .A3(new_n14853_), .ZN(new_n15093_));
  AOI22_X1   g14901(.A1(new_n15093_), .A2(new_n14867_), .B1(\asqrt[44] ), .B2(new_n14876_), .ZN(new_n15094_));
  OAI21_X1   g14902(.A1(new_n15094_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n15095_));
  OAI21_X1   g14903(.A1(new_n15095_), .A2(new_n14878_), .B(new_n15085_), .ZN(new_n15096_));
  NAND3_X1   g14904(.A1(new_n15096_), .A2(new_n2229_), .A3(new_n14879_), .ZN(new_n15097_));
  AOI22_X1   g14905(.A1(new_n15097_), .A2(new_n14893_), .B1(\asqrt[47] ), .B2(new_n14902_), .ZN(new_n15098_));
  OAI21_X1   g14906(.A1(new_n15098_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n15099_));
  OAI21_X1   g14907(.A1(new_n15099_), .A2(new_n14904_), .B(new_n15084_), .ZN(new_n15100_));
  NAND3_X1   g14908(.A1(new_n15100_), .A2(new_n1612_), .A3(new_n14905_), .ZN(new_n15101_));
  AOI22_X1   g14909(.A1(new_n15101_), .A2(new_n14919_), .B1(\asqrt[50] ), .B2(new_n14928_), .ZN(new_n15102_));
  OAI21_X1   g14910(.A1(new_n15102_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n15103_));
  OAI21_X1   g14911(.A1(new_n15103_), .A2(new_n14930_), .B(new_n15083_), .ZN(new_n15104_));
  NAND3_X1   g14912(.A1(new_n15104_), .A2(new_n1103_), .A3(new_n14931_), .ZN(new_n15105_));
  AOI22_X1   g14913(.A1(new_n15105_), .A2(new_n14946_), .B1(\asqrt[53] ), .B2(new_n14975_), .ZN(new_n15106_));
  OAI21_X1   g14914(.A1(new_n15106_), .A2(new_n904_), .B(new_n823_), .ZN(new_n15107_));
  OAI21_X1   g14915(.A1(new_n15107_), .A2(new_n14977_), .B(new_n15082_), .ZN(new_n15108_));
  NAND3_X1   g14916(.A1(new_n15108_), .A2(new_n703_), .A3(new_n14978_), .ZN(new_n15109_));
  AOI22_X1   g14917(.A1(new_n15109_), .A2(new_n14973_), .B1(\asqrt[56] ), .B2(new_n15007_), .ZN(new_n15110_));
  OAI21_X1   g14918(.A1(new_n15110_), .A2(new_n531_), .B(new_n436_), .ZN(new_n15111_));
  OAI21_X1   g14919(.A1(new_n15111_), .A2(new_n15009_), .B(new_n15081_), .ZN(new_n15112_));
  NAND3_X1   g14920(.A1(new_n15112_), .A2(new_n327_), .A3(new_n15010_), .ZN(new_n15113_));
  AOI22_X1   g14921(.A1(new_n15113_), .A2(new_n15005_), .B1(new_n15039_), .B2(\asqrt[59] ), .ZN(new_n15114_));
  OAI21_X1   g14922(.A1(new_n15114_), .A2(new_n306_), .B(new_n218_), .ZN(new_n15115_));
  OAI21_X1   g14923(.A1(new_n15115_), .A2(new_n15041_), .B(new_n15080_), .ZN(new_n15116_));
  NAND3_X1   g14924(.A1(new_n15116_), .A2(new_n207_), .A3(new_n15042_), .ZN(new_n15117_));
  AOI22_X1   g14925(.A1(new_n15117_), .A2(new_n15037_), .B1(new_n15079_), .B2(\asqrt[62] ), .ZN(new_n15118_));
  OAI21_X1   g14926(.A1(new_n15118_), .A2(new_n15053_), .B(new_n193_), .ZN(new_n15119_));
  AOI21_X1   g14927(.A1(new_n15079_), .A2(\asqrt[62] ), .B(new_n15049_), .ZN(new_n15120_));
  AOI21_X1   g14928(.A1(new_n15120_), .A2(new_n15044_), .B(new_n15064_), .ZN(new_n15121_));
  AOI21_X1   g14929(.A1(new_n15119_), .A2(new_n15121_), .B(new_n14553_), .ZN(new_n15122_));
  OAI21_X1   g14930(.A1(new_n15055_), .A2(new_n15066_), .B(new_n15068_), .ZN(new_n15123_));
  AOI21_X1   g14931(.A1(\a[31] ), .A2(new_n15123_), .B(new_n15122_), .ZN(new_n15124_));
  AOI22_X1   g14932(.A1(new_n15124_), .A2(new_n15077_), .B1(\asqrt[16] ), .B2(new_n15073_), .ZN(new_n15125_));
  NOR2_X1    g14933(.A1(new_n15125_), .A2(new_n14017_), .ZN(new_n15126_));
  NAND2_X1   g14934(.A1(new_n15124_), .A2(new_n15077_), .ZN(new_n15127_));
  OAI21_X1   g14935(.A1(new_n15055_), .A2(new_n15066_), .B(new_n14552_), .ZN(new_n15128_));
  NAND2_X1   g14936(.A1(new_n15120_), .A2(new_n15044_), .ZN(new_n15129_));
  OAI21_X1   g14937(.A1(new_n15062_), .A2(new_n14550_), .B(new_n14398_), .ZN(new_n15130_));
  NAND4_X1   g14938(.A1(new_n15119_), .A2(new_n15129_), .A3(new_n15060_), .A4(new_n15130_), .ZN(new_n15131_));
  AOI21_X1   g14939(.A1(new_n15131_), .A2(new_n15128_), .B(new_n14565_), .ZN(new_n15132_));
  INV_X1     g14940(.I(new_n15129_), .ZN(new_n15133_));
  NAND2_X1   g14941(.A1(new_n15060_), .A2(new_n15130_), .ZN(new_n15134_));
  NOR3_X1    g14942(.A1(new_n15133_), .A2(new_n15055_), .A3(new_n15134_), .ZN(new_n15135_));
  NOR3_X1    g14943(.A1(new_n15135_), .A2(new_n15122_), .A3(\a[32] ), .ZN(new_n15136_));
  NOR2_X1    g14944(.A1(new_n15132_), .A2(new_n15136_), .ZN(new_n15137_));
  AOI21_X1   g14945(.A1(new_n15073_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n15138_));
  AOI21_X1   g14946(.A1(new_n15127_), .A2(new_n15138_), .B(new_n15137_), .ZN(new_n15139_));
  OAI21_X1   g14947(.A1(new_n15139_), .A2(new_n15126_), .B(\asqrt[18] ), .ZN(new_n15140_));
  OAI21_X1   g14948(.A1(\asqrt[63] ), .A2(new_n15054_), .B(new_n15121_), .ZN(\asqrt[15] ));
  NOR3_X1    g14949(.A1(new_n14645_), .A2(new_n14564_), .A3(new_n14570_), .ZN(new_n15142_));
  NAND3_X1   g14950(.A1(\asqrt[15] ), .A2(new_n14583_), .A3(new_n14630_), .ZN(new_n15143_));
  AOI22_X1   g14951(.A1(new_n15143_), .A2(new_n14645_), .B1(\asqrt[15] ), .B2(new_n15142_), .ZN(new_n15144_));
  INV_X1     g14952(.I(new_n15144_), .ZN(new_n15145_));
  OAI21_X1   g14953(.A1(new_n15125_), .A2(new_n14017_), .B(new_n13353_), .ZN(new_n15146_));
  OAI21_X1   g14954(.A1(new_n15146_), .A2(new_n15139_), .B(new_n15145_), .ZN(new_n15147_));
  AOI21_X1   g14955(.A1(new_n15147_), .A2(new_n15140_), .B(new_n12913_), .ZN(new_n15148_));
  NOR2_X1    g14956(.A1(new_n14582_), .A2(new_n14580_), .ZN(new_n15149_));
  NOR2_X1    g14957(.A1(new_n14574_), .A2(new_n14584_), .ZN(new_n15150_));
  INV_X1     g14958(.I(new_n15150_), .ZN(new_n15151_));
  NAND4_X1   g14959(.A1(\asqrt[15] ), .A2(new_n14575_), .A3(new_n15149_), .A4(new_n15151_), .ZN(new_n15152_));
  NOR3_X1    g14960(.A1(new_n15067_), .A2(new_n14634_), .A3(new_n15150_), .ZN(new_n15153_));
  OAI21_X1   g14961(.A1(new_n15153_), .A2(new_n15149_), .B(new_n15152_), .ZN(new_n15154_));
  INV_X1     g14962(.I(new_n15154_), .ZN(new_n15155_));
  AOI21_X1   g14963(.A1(new_n15119_), .A2(new_n15121_), .B(new_n15068_), .ZN(new_n15156_));
  OAI21_X1   g14964(.A1(new_n15156_), .A2(new_n15071_), .B(\asqrt[16] ), .ZN(new_n15157_));
  INV_X1     g14965(.I(new_n15157_), .ZN(new_n15158_));
  NOR2_X1    g14966(.A1(new_n15156_), .A2(new_n15075_), .ZN(new_n15159_));
  INV_X1     g14967(.I(\a[31] ), .ZN(new_n15160_));
  AOI21_X1   g14968(.A1(\asqrt[15] ), .A2(new_n15068_), .B(new_n15160_), .ZN(new_n15161_));
  NOR3_X1    g14969(.A1(new_n15159_), .A2(new_n15161_), .A3(new_n15122_), .ZN(new_n15162_));
  OAI21_X1   g14970(.A1(new_n15162_), .A2(new_n15158_), .B(\asqrt[17] ), .ZN(new_n15163_));
  AOI21_X1   g14971(.A1(\asqrt[15] ), .A2(\a[30] ), .B(new_n15071_), .ZN(new_n15164_));
  OAI21_X1   g14972(.A1(new_n15164_), .A2(new_n14601_), .B(new_n14017_), .ZN(new_n15165_));
  OAI22_X1   g14973(.A1(new_n15162_), .A2(new_n15165_), .B1(new_n15132_), .B2(new_n15136_), .ZN(new_n15166_));
  AOI21_X1   g14974(.A1(new_n15166_), .A2(new_n15163_), .B(new_n13353_), .ZN(new_n15167_));
  AOI21_X1   g14975(.A1(new_n15119_), .A2(new_n15121_), .B(\a[30] ), .ZN(new_n15168_));
  OAI21_X1   g14976(.A1(new_n15160_), .A2(new_n15168_), .B(new_n15128_), .ZN(new_n15169_));
  OAI21_X1   g14977(.A1(new_n15169_), .A2(new_n15159_), .B(new_n15157_), .ZN(new_n15170_));
  AOI21_X1   g14978(.A1(new_n15170_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n15171_));
  AOI21_X1   g14979(.A1(new_n15171_), .A2(new_n15166_), .B(new_n15144_), .ZN(new_n15172_));
  NOR3_X1    g14980(.A1(new_n15172_), .A2(new_n15167_), .A3(\asqrt[19] ), .ZN(new_n15173_));
  NOR2_X1    g14981(.A1(new_n15173_), .A2(new_n15155_), .ZN(new_n15174_));
  OAI21_X1   g14982(.A1(new_n15174_), .A2(new_n15148_), .B(\asqrt[20] ), .ZN(new_n15175_));
  NOR2_X1    g14983(.A1(new_n14647_), .A2(new_n14639_), .ZN(new_n15176_));
  NOR3_X1    g14984(.A1(new_n15067_), .A2(new_n14586_), .A3(new_n15176_), .ZN(new_n15177_));
  INV_X1     g14985(.I(new_n15177_), .ZN(new_n15178_));
  NOR3_X1    g14986(.A1(new_n15176_), .A2(new_n14586_), .A3(new_n14644_), .ZN(new_n15179_));
  AOI22_X1   g14987(.A1(new_n15178_), .A2(new_n14644_), .B1(\asqrt[15] ), .B2(new_n15179_), .ZN(new_n15180_));
  INV_X1     g14988(.I(new_n15180_), .ZN(new_n15181_));
  OAI21_X1   g14989(.A1(new_n15172_), .A2(new_n15167_), .B(\asqrt[19] ), .ZN(new_n15182_));
  NAND2_X1   g14990(.A1(new_n15182_), .A2(new_n12364_), .ZN(new_n15183_));
  OAI21_X1   g14991(.A1(new_n15174_), .A2(new_n15183_), .B(new_n15181_), .ZN(new_n15184_));
  AOI21_X1   g14992(.A1(new_n15184_), .A2(new_n15175_), .B(new_n11736_), .ZN(new_n15185_));
  NOR3_X1    g14993(.A1(new_n14596_), .A2(new_n14605_), .A3(new_n14603_), .ZN(new_n15186_));
  NOR3_X1    g14994(.A1(new_n15067_), .A2(new_n14596_), .A3(new_n14605_), .ZN(new_n15187_));
  INV_X1     g14995(.I(new_n15187_), .ZN(new_n15188_));
  AOI22_X1   g14996(.A1(new_n15188_), .A2(new_n14603_), .B1(\asqrt[15] ), .B2(new_n15186_), .ZN(new_n15189_));
  OAI21_X1   g14997(.A1(new_n15155_), .A2(new_n15173_), .B(new_n15182_), .ZN(new_n15190_));
  AOI21_X1   g14998(.A1(new_n15190_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n15191_));
  AOI21_X1   g14999(.A1(new_n15191_), .A2(new_n15184_), .B(new_n15189_), .ZN(new_n15192_));
  OAI21_X1   g15000(.A1(new_n15192_), .A2(new_n15185_), .B(\asqrt[22] ), .ZN(new_n15193_));
  INV_X1     g15001(.I(new_n15193_), .ZN(new_n15194_));
  NAND2_X1   g15002(.A1(new_n14650_), .A2(new_n14642_), .ZN(new_n15195_));
  NAND3_X1   g15003(.A1(\asqrt[15] ), .A2(new_n14607_), .A3(new_n15195_), .ZN(new_n15196_));
  AND3_X2    g15004(.A1(new_n14607_), .A2(new_n14612_), .A3(new_n15195_), .Z(new_n15197_));
  AOI22_X1   g15005(.A1(new_n15196_), .A2(new_n14613_), .B1(\asqrt[15] ), .B2(new_n15197_), .ZN(new_n15198_));
  NOR3_X1    g15006(.A1(new_n15192_), .A2(new_n15185_), .A3(\asqrt[22] ), .ZN(new_n15199_));
  NOR2_X1    g15007(.A1(new_n15199_), .A2(new_n15198_), .ZN(new_n15200_));
  OAI21_X1   g15008(.A1(new_n15200_), .A2(new_n15194_), .B(\asqrt[23] ), .ZN(new_n15201_));
  INV_X1     g15009(.I(new_n14620_), .ZN(new_n15202_));
  NOR3_X1    g15010(.A1(new_n14616_), .A2(new_n14661_), .A3(new_n15202_), .ZN(new_n15203_));
  NOR3_X1    g15011(.A1(new_n15067_), .A2(new_n14616_), .A3(new_n14661_), .ZN(new_n15204_));
  INV_X1     g15012(.I(new_n15204_), .ZN(new_n15205_));
  AOI22_X1   g15013(.A1(new_n15205_), .A2(new_n15202_), .B1(\asqrt[15] ), .B2(new_n15203_), .ZN(new_n15206_));
  INV_X1     g15014(.I(new_n15206_), .ZN(new_n15207_));
  NAND2_X1   g15015(.A1(new_n15193_), .A2(new_n10812_), .ZN(new_n15208_));
  OAI21_X1   g15016(.A1(new_n15200_), .A2(new_n15208_), .B(new_n15207_), .ZN(new_n15209_));
  AOI21_X1   g15017(.A1(new_n15209_), .A2(new_n15201_), .B(new_n10221_), .ZN(new_n15210_));
  INV_X1     g15018(.I(new_n14686_), .ZN(new_n15211_));
  NAND3_X1   g15019(.A1(\asqrt[15] ), .A2(new_n14624_), .A3(new_n15211_), .ZN(new_n15212_));
  AND3_X2    g15020(.A1(new_n15211_), .A2(new_n14624_), .A3(new_n14628_), .Z(new_n15213_));
  AOI22_X1   g15021(.A1(new_n15212_), .A2(new_n14629_), .B1(\asqrt[15] ), .B2(new_n15213_), .ZN(new_n15214_));
  OAI21_X1   g15022(.A1(new_n15198_), .A2(new_n15199_), .B(new_n15193_), .ZN(new_n15215_));
  AOI21_X1   g15023(.A1(new_n15215_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n15216_));
  AOI21_X1   g15024(.A1(new_n15216_), .A2(new_n15209_), .B(new_n15214_), .ZN(new_n15217_));
  OAI21_X1   g15025(.A1(new_n15217_), .A2(new_n15210_), .B(\asqrt[25] ), .ZN(new_n15218_));
  INV_X1     g15026(.I(new_n15218_), .ZN(new_n15219_));
  INV_X1     g15027(.I(new_n14689_), .ZN(new_n15220_));
  NOR3_X1    g15028(.A1(new_n15220_), .A2(new_n14655_), .A3(new_n14688_), .ZN(new_n15221_));
  NOR3_X1    g15029(.A1(new_n15067_), .A2(new_n14655_), .A3(new_n15220_), .ZN(new_n15222_));
  INV_X1     g15030(.I(new_n15222_), .ZN(new_n15223_));
  AOI22_X1   g15031(.A1(new_n15223_), .A2(new_n14688_), .B1(\asqrt[15] ), .B2(new_n15221_), .ZN(new_n15224_));
  NOR3_X1    g15032(.A1(new_n15217_), .A2(new_n15210_), .A3(\asqrt[25] ), .ZN(new_n15225_));
  NOR2_X1    g15033(.A1(new_n15225_), .A2(new_n15224_), .ZN(new_n15226_));
  OAI21_X1   g15034(.A1(new_n15226_), .A2(new_n15219_), .B(\asqrt[26] ), .ZN(new_n15227_));
  INV_X1     g15035(.I(new_n14670_), .ZN(new_n15228_));
  NOR3_X1    g15036(.A1(new_n15067_), .A2(new_n14666_), .A3(new_n14671_), .ZN(new_n15229_));
  INV_X1     g15037(.I(new_n15229_), .ZN(new_n15230_));
  NOR3_X1    g15038(.A1(new_n14666_), .A2(new_n15228_), .A3(new_n14671_), .ZN(new_n15231_));
  AOI22_X1   g15039(.A1(new_n15230_), .A2(new_n15228_), .B1(\asqrt[15] ), .B2(new_n15231_), .ZN(new_n15232_));
  INV_X1     g15040(.I(new_n15232_), .ZN(new_n15233_));
  NAND2_X1   g15041(.A1(new_n15218_), .A2(new_n9317_), .ZN(new_n15234_));
  OAI21_X1   g15042(.A1(new_n15226_), .A2(new_n15234_), .B(new_n15233_), .ZN(new_n15235_));
  AOI21_X1   g15043(.A1(new_n15235_), .A2(new_n15227_), .B(new_n8826_), .ZN(new_n15236_));
  OAI21_X1   g15044(.A1(new_n14672_), .A2(new_n14678_), .B(new_n14676_), .ZN(new_n15237_));
  AOI21_X1   g15045(.A1(\asqrt[26] ), .A2(new_n14691_), .B(new_n15237_), .ZN(new_n15238_));
  OAI21_X1   g15046(.A1(new_n14672_), .A2(new_n14678_), .B(new_n14673_), .ZN(new_n15239_));
  NOR2_X1    g15047(.A1(new_n15067_), .A2(new_n15239_), .ZN(new_n15240_));
  INV_X1     g15048(.I(new_n15240_), .ZN(new_n15241_));
  AOI22_X1   g15049(.A1(new_n15241_), .A2(new_n14677_), .B1(\asqrt[15] ), .B2(new_n15238_), .ZN(new_n15242_));
  OAI21_X1   g15050(.A1(new_n15224_), .A2(new_n15225_), .B(new_n15218_), .ZN(new_n15243_));
  AOI21_X1   g15051(.A1(new_n15243_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n15244_));
  AOI21_X1   g15052(.A1(new_n15244_), .A2(new_n15235_), .B(new_n15242_), .ZN(new_n15245_));
  OAI21_X1   g15053(.A1(new_n15245_), .A2(new_n15236_), .B(\asqrt[28] ), .ZN(new_n15246_));
  INV_X1     g15054(.I(new_n15246_), .ZN(new_n15247_));
  INV_X1     g15055(.I(new_n14685_), .ZN(new_n15248_));
  INV_X1     g15056(.I(new_n14679_), .ZN(new_n15249_));
  INV_X1     g15057(.I(new_n14692_), .ZN(new_n15250_));
  NOR2_X1    g15058(.A1(new_n15250_), .A2(new_n15249_), .ZN(new_n15251_));
  NOR3_X1    g15059(.A1(new_n15067_), .A2(new_n14680_), .A3(new_n15251_), .ZN(new_n15252_));
  INV_X1     g15060(.I(new_n15252_), .ZN(new_n15253_));
  NOR3_X1    g15061(.A1(new_n15251_), .A2(new_n14680_), .A3(new_n15248_), .ZN(new_n15254_));
  AOI22_X1   g15062(.A1(new_n15253_), .A2(new_n15248_), .B1(\asqrt[15] ), .B2(new_n15254_), .ZN(new_n15255_));
  NOR3_X1    g15063(.A1(new_n15245_), .A2(new_n15236_), .A3(\asqrt[28] ), .ZN(new_n15256_));
  NOR2_X1    g15064(.A1(new_n15256_), .A2(new_n15255_), .ZN(new_n15257_));
  OAI21_X1   g15065(.A1(new_n15257_), .A2(new_n15247_), .B(\asqrt[29] ), .ZN(new_n15258_));
  INV_X1     g15066(.I(new_n14700_), .ZN(new_n15259_));
  NOR3_X1    g15067(.A1(new_n14695_), .A2(new_n15259_), .A3(new_n14737_), .ZN(new_n15260_));
  NOR3_X1    g15068(.A1(new_n15067_), .A2(new_n14695_), .A3(new_n14737_), .ZN(new_n15261_));
  INV_X1     g15069(.I(new_n15261_), .ZN(new_n15262_));
  AOI22_X1   g15070(.A1(new_n15262_), .A2(new_n15259_), .B1(\asqrt[15] ), .B2(new_n15260_), .ZN(new_n15263_));
  INV_X1     g15071(.I(new_n15263_), .ZN(new_n15264_));
  NAND2_X1   g15072(.A1(new_n15246_), .A2(new_n8036_), .ZN(new_n15265_));
  OAI21_X1   g15073(.A1(new_n15257_), .A2(new_n15265_), .B(new_n15264_), .ZN(new_n15266_));
  AOI21_X1   g15074(.A1(new_n15266_), .A2(new_n15258_), .B(new_n7539_), .ZN(new_n15267_));
  NOR2_X1    g15075(.A1(new_n14710_), .A2(new_n14702_), .ZN(new_n15268_));
  INV_X1     g15076(.I(new_n15268_), .ZN(new_n15269_));
  NAND3_X1   g15077(.A1(\asqrt[15] ), .A2(new_n14703_), .A3(new_n15269_), .ZN(new_n15270_));
  AND3_X2    g15078(.A1(new_n15269_), .A2(new_n14703_), .A3(new_n14708_), .Z(new_n15271_));
  AOI22_X1   g15079(.A1(new_n15270_), .A2(new_n14709_), .B1(\asqrt[15] ), .B2(new_n15271_), .ZN(new_n15272_));
  OAI21_X1   g15080(.A1(new_n15255_), .A2(new_n15256_), .B(new_n15246_), .ZN(new_n15273_));
  AOI21_X1   g15081(.A1(new_n15273_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n15274_));
  AOI21_X1   g15082(.A1(new_n15274_), .A2(new_n15266_), .B(new_n15272_), .ZN(new_n15275_));
  OAI21_X1   g15083(.A1(new_n15275_), .A2(new_n15267_), .B(\asqrt[31] ), .ZN(new_n15276_));
  INV_X1     g15084(.I(new_n15276_), .ZN(new_n15277_));
  NOR2_X1    g15085(.A1(new_n14721_), .A2(new_n14714_), .ZN(new_n15278_));
  NOR3_X1    g15086(.A1(new_n15278_), .A2(new_n14712_), .A3(new_n14720_), .ZN(new_n15279_));
  NOR3_X1    g15087(.A1(new_n15067_), .A2(new_n14712_), .A3(new_n15278_), .ZN(new_n15280_));
  INV_X1     g15088(.I(new_n15280_), .ZN(new_n15281_));
  AOI22_X1   g15089(.A1(new_n15281_), .A2(new_n14720_), .B1(\asqrt[15] ), .B2(new_n15279_), .ZN(new_n15282_));
  NOR3_X1    g15090(.A1(new_n15275_), .A2(new_n15267_), .A3(\asqrt[31] ), .ZN(new_n15283_));
  NOR2_X1    g15091(.A1(new_n15283_), .A2(new_n15282_), .ZN(new_n15284_));
  OAI21_X1   g15092(.A1(new_n15284_), .A2(new_n15277_), .B(\asqrt[32] ), .ZN(new_n15285_));
  INV_X1     g15093(.I(new_n14727_), .ZN(new_n15286_));
  NOR3_X1    g15094(.A1(new_n15067_), .A2(new_n14723_), .A3(new_n14769_), .ZN(new_n15287_));
  INV_X1     g15095(.I(new_n15287_), .ZN(new_n15288_));
  NOR3_X1    g15096(.A1(new_n14723_), .A2(new_n15286_), .A3(new_n14769_), .ZN(new_n15289_));
  AOI22_X1   g15097(.A1(new_n15288_), .A2(new_n15286_), .B1(\asqrt[15] ), .B2(new_n15289_), .ZN(new_n15290_));
  INV_X1     g15098(.I(new_n15290_), .ZN(new_n15291_));
  NAND2_X1   g15099(.A1(new_n15276_), .A2(new_n6824_), .ZN(new_n15292_));
  OAI21_X1   g15100(.A1(new_n15284_), .A2(new_n15292_), .B(new_n15291_), .ZN(new_n15293_));
  AOI21_X1   g15101(.A1(new_n15293_), .A2(new_n15285_), .B(new_n6356_), .ZN(new_n15294_));
  NOR2_X1    g15102(.A1(new_n14742_), .A2(new_n14729_), .ZN(new_n15295_));
  INV_X1     g15103(.I(new_n15295_), .ZN(new_n15296_));
  AND3_X2    g15104(.A1(new_n15296_), .A2(new_n14730_), .A3(new_n14735_), .Z(new_n15297_));
  NAND3_X1   g15105(.A1(\asqrt[15] ), .A2(new_n14730_), .A3(new_n15296_), .ZN(new_n15298_));
  AOI22_X1   g15106(.A1(new_n15298_), .A2(new_n14736_), .B1(\asqrt[15] ), .B2(new_n15297_), .ZN(new_n15299_));
  OAI21_X1   g15107(.A1(new_n15282_), .A2(new_n15283_), .B(new_n15276_), .ZN(new_n15300_));
  AOI21_X1   g15108(.A1(new_n15300_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n15301_));
  AOI21_X1   g15109(.A1(new_n15301_), .A2(new_n15293_), .B(new_n15299_), .ZN(new_n15302_));
  OAI21_X1   g15110(.A1(new_n15302_), .A2(new_n15294_), .B(\asqrt[34] ), .ZN(new_n15303_));
  INV_X1     g15111(.I(new_n15303_), .ZN(new_n15304_));
  NOR2_X1    g15112(.A1(new_n14753_), .A2(new_n14746_), .ZN(new_n15305_));
  NOR3_X1    g15113(.A1(new_n15067_), .A2(new_n14744_), .A3(new_n15305_), .ZN(new_n15306_));
  INV_X1     g15114(.I(new_n15306_), .ZN(new_n15307_));
  NOR3_X1    g15115(.A1(new_n15305_), .A2(new_n14744_), .A3(new_n14752_), .ZN(new_n15308_));
  AOI22_X1   g15116(.A1(new_n15307_), .A2(new_n14752_), .B1(\asqrt[15] ), .B2(new_n15308_), .ZN(new_n15309_));
  NOR3_X1    g15117(.A1(new_n15302_), .A2(new_n15294_), .A3(\asqrt[34] ), .ZN(new_n15310_));
  NOR2_X1    g15118(.A1(new_n15310_), .A2(new_n15309_), .ZN(new_n15311_));
  OAI21_X1   g15119(.A1(new_n15311_), .A2(new_n15304_), .B(\asqrt[35] ), .ZN(new_n15312_));
  INV_X1     g15120(.I(new_n14759_), .ZN(new_n15313_));
  NOR3_X1    g15121(.A1(new_n14755_), .A2(new_n15313_), .A3(new_n14819_), .ZN(new_n15314_));
  NOR3_X1    g15122(.A1(new_n15067_), .A2(new_n14755_), .A3(new_n14819_), .ZN(new_n15315_));
  INV_X1     g15123(.I(new_n15315_), .ZN(new_n15316_));
  AOI22_X1   g15124(.A1(new_n15316_), .A2(new_n15313_), .B1(\asqrt[15] ), .B2(new_n15314_), .ZN(new_n15317_));
  INV_X1     g15125(.I(new_n15317_), .ZN(new_n15318_));
  NAND2_X1   g15126(.A1(new_n15303_), .A2(new_n5708_), .ZN(new_n15319_));
  OAI21_X1   g15127(.A1(new_n15311_), .A2(new_n15319_), .B(new_n15318_), .ZN(new_n15320_));
  AOI21_X1   g15128(.A1(new_n15320_), .A2(new_n15312_), .B(new_n5277_), .ZN(new_n15321_));
  NOR2_X1    g15129(.A1(new_n14774_), .A2(new_n14761_), .ZN(new_n15322_));
  INV_X1     g15130(.I(new_n15322_), .ZN(new_n15323_));
  NAND3_X1   g15131(.A1(\asqrt[15] ), .A2(new_n14762_), .A3(new_n15323_), .ZN(new_n15324_));
  AND3_X2    g15132(.A1(new_n15323_), .A2(new_n14762_), .A3(new_n14767_), .Z(new_n15325_));
  AOI22_X1   g15133(.A1(new_n15324_), .A2(new_n14768_), .B1(\asqrt[15] ), .B2(new_n15325_), .ZN(new_n15326_));
  OAI21_X1   g15134(.A1(new_n15309_), .A2(new_n15310_), .B(new_n15303_), .ZN(new_n15327_));
  AOI21_X1   g15135(.A1(new_n15327_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n15328_));
  AOI21_X1   g15136(.A1(new_n15328_), .A2(new_n15320_), .B(new_n15326_), .ZN(new_n15329_));
  OAI21_X1   g15137(.A1(new_n15329_), .A2(new_n15321_), .B(\asqrt[37] ), .ZN(new_n15330_));
  INV_X1     g15138(.I(new_n15330_), .ZN(new_n15331_));
  NOR2_X1    g15139(.A1(new_n14778_), .A2(new_n14785_), .ZN(new_n15332_));
  NOR3_X1    g15140(.A1(new_n15332_), .A2(new_n14792_), .A3(new_n14784_), .ZN(new_n15333_));
  NOR3_X1    g15141(.A1(new_n15067_), .A2(new_n14792_), .A3(new_n15332_), .ZN(new_n15334_));
  INV_X1     g15142(.I(new_n15334_), .ZN(new_n15335_));
  AOI22_X1   g15143(.A1(new_n15335_), .A2(new_n14784_), .B1(\asqrt[15] ), .B2(new_n15333_), .ZN(new_n15336_));
  NOR3_X1    g15144(.A1(new_n15329_), .A2(new_n15321_), .A3(\asqrt[37] ), .ZN(new_n15337_));
  NOR2_X1    g15145(.A1(new_n15337_), .A2(new_n15336_), .ZN(new_n15338_));
  OAI21_X1   g15146(.A1(new_n15338_), .A2(new_n15331_), .B(\asqrt[38] ), .ZN(new_n15339_));
  INV_X1     g15147(.I(new_n14791_), .ZN(new_n15340_));
  NOR3_X1    g15148(.A1(new_n15067_), .A2(new_n14787_), .A3(new_n14836_), .ZN(new_n15341_));
  INV_X1     g15149(.I(new_n15341_), .ZN(new_n15342_));
  NOR3_X1    g15150(.A1(new_n14787_), .A2(new_n15340_), .A3(new_n14836_), .ZN(new_n15343_));
  AOI22_X1   g15151(.A1(new_n15342_), .A2(new_n15340_), .B1(\asqrt[15] ), .B2(new_n15343_), .ZN(new_n15344_));
  INV_X1     g15152(.I(new_n15344_), .ZN(new_n15345_));
  NAND2_X1   g15153(.A1(new_n15330_), .A2(new_n4696_), .ZN(new_n15346_));
  OAI21_X1   g15154(.A1(new_n15338_), .A2(new_n15346_), .B(new_n15345_), .ZN(new_n15347_));
  AOI21_X1   g15155(.A1(new_n15347_), .A2(new_n15339_), .B(new_n4298_), .ZN(new_n15348_));
  NOR3_X1    g15156(.A1(new_n14796_), .A2(new_n14818_), .A3(new_n14802_), .ZN(new_n15349_));
  NOR3_X1    g15157(.A1(new_n15067_), .A2(new_n14796_), .A3(new_n14802_), .ZN(new_n15350_));
  INV_X1     g15158(.I(new_n15350_), .ZN(new_n15351_));
  AOI22_X1   g15159(.A1(new_n15351_), .A2(new_n14818_), .B1(\asqrt[15] ), .B2(new_n15349_), .ZN(new_n15352_));
  OAI21_X1   g15160(.A1(new_n15336_), .A2(new_n15337_), .B(new_n15330_), .ZN(new_n15353_));
  AOI21_X1   g15161(.A1(new_n15353_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n15354_));
  AOI21_X1   g15162(.A1(new_n15354_), .A2(new_n15347_), .B(new_n15352_), .ZN(new_n15355_));
  OAI21_X1   g15163(.A1(new_n15355_), .A2(new_n15348_), .B(\asqrt[40] ), .ZN(new_n15356_));
  INV_X1     g15164(.I(new_n15356_), .ZN(new_n15357_));
  NOR2_X1    g15165(.A1(new_n14803_), .A2(new_n14811_), .ZN(new_n15358_));
  NOR3_X1    g15166(.A1(new_n15067_), .A2(new_n14826_), .A3(new_n15358_), .ZN(new_n15359_));
  INV_X1     g15167(.I(new_n15359_), .ZN(new_n15360_));
  NOR3_X1    g15168(.A1(new_n15358_), .A2(new_n14826_), .A3(new_n14810_), .ZN(new_n15361_));
  AOI22_X1   g15169(.A1(new_n15360_), .A2(new_n14810_), .B1(\asqrt[15] ), .B2(new_n15361_), .ZN(new_n15362_));
  NOR3_X1    g15170(.A1(new_n15355_), .A2(new_n15348_), .A3(\asqrt[40] ), .ZN(new_n15363_));
  NOR2_X1    g15171(.A1(new_n15363_), .A2(new_n15362_), .ZN(new_n15364_));
  OAI21_X1   g15172(.A1(new_n15364_), .A2(new_n15357_), .B(\asqrt[41] ), .ZN(new_n15365_));
  INV_X1     g15173(.I(new_n14817_), .ZN(new_n15366_));
  NOR3_X1    g15174(.A1(new_n14813_), .A2(new_n15366_), .A3(new_n14849_), .ZN(new_n15367_));
  NOR3_X1    g15175(.A1(new_n15067_), .A2(new_n14813_), .A3(new_n14849_), .ZN(new_n15368_));
  INV_X1     g15176(.I(new_n15368_), .ZN(new_n15369_));
  AOI22_X1   g15177(.A1(new_n15369_), .A2(new_n15366_), .B1(\asqrt[15] ), .B2(new_n15367_), .ZN(new_n15370_));
  INV_X1     g15178(.I(new_n15370_), .ZN(new_n15371_));
  NAND2_X1   g15179(.A1(new_n15356_), .A2(new_n3782_), .ZN(new_n15372_));
  OAI21_X1   g15180(.A1(new_n15364_), .A2(new_n15372_), .B(new_n15371_), .ZN(new_n15373_));
  AOI21_X1   g15181(.A1(new_n15373_), .A2(new_n15365_), .B(new_n3419_), .ZN(new_n15374_));
  NOR3_X1    g15182(.A1(new_n15067_), .A2(new_n15087_), .A3(new_n15088_), .ZN(new_n15375_));
  INV_X1     g15183(.I(new_n15375_), .ZN(new_n15376_));
  NOR3_X1    g15184(.A1(new_n15087_), .A2(new_n14835_), .A3(new_n15088_), .ZN(new_n15377_));
  AOI22_X1   g15185(.A1(new_n15376_), .A2(new_n14835_), .B1(\asqrt[15] ), .B2(new_n15377_), .ZN(new_n15378_));
  OAI21_X1   g15186(.A1(new_n15362_), .A2(new_n15363_), .B(new_n15356_), .ZN(new_n15379_));
  AOI21_X1   g15187(.A1(new_n15379_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n15380_));
  AOI21_X1   g15188(.A1(new_n15380_), .A2(new_n15373_), .B(new_n15378_), .ZN(new_n15381_));
  OAI21_X1   g15189(.A1(new_n15381_), .A2(new_n15374_), .B(\asqrt[43] ), .ZN(new_n15382_));
  INV_X1     g15190(.I(new_n15382_), .ZN(new_n15383_));
  INV_X1     g15191(.I(new_n14848_), .ZN(new_n15384_));
  NAND2_X1   g15192(.A1(new_n14829_), .A2(new_n3419_), .ZN(new_n15385_));
  NOR2_X1    g15193(.A1(new_n15089_), .A2(new_n15385_), .ZN(new_n15386_));
  NOR3_X1    g15194(.A1(new_n15386_), .A2(new_n14843_), .A3(new_n15384_), .ZN(new_n15387_));
  NOR3_X1    g15195(.A1(new_n15067_), .A2(new_n14843_), .A3(new_n15386_), .ZN(new_n15388_));
  INV_X1     g15196(.I(new_n15388_), .ZN(new_n15389_));
  AOI22_X1   g15197(.A1(new_n15389_), .A2(new_n15384_), .B1(\asqrt[15] ), .B2(new_n15387_), .ZN(new_n15390_));
  NOR3_X1    g15198(.A1(new_n15381_), .A2(new_n15374_), .A3(\asqrt[43] ), .ZN(new_n15391_));
  NOR2_X1    g15199(.A1(new_n15391_), .A2(new_n15390_), .ZN(new_n15392_));
  OAI21_X1   g15200(.A1(new_n15392_), .A2(new_n15383_), .B(\asqrt[44] ), .ZN(new_n15393_));
  NOR3_X1    g15201(.A1(new_n15067_), .A2(new_n14854_), .A3(new_n14859_), .ZN(new_n15394_));
  INV_X1     g15202(.I(new_n15394_), .ZN(new_n15395_));
  NOR3_X1    g15203(.A1(new_n14854_), .A2(new_n14859_), .A3(new_n15086_), .ZN(new_n15396_));
  AOI22_X1   g15204(.A1(new_n15395_), .A2(new_n15086_), .B1(\asqrt[15] ), .B2(new_n15396_), .ZN(new_n15397_));
  INV_X1     g15205(.I(new_n15397_), .ZN(new_n15398_));
  NAND2_X1   g15206(.A1(new_n15382_), .A2(new_n2954_), .ZN(new_n15399_));
  OAI21_X1   g15207(.A1(new_n15392_), .A2(new_n15399_), .B(new_n15398_), .ZN(new_n15400_));
  AOI21_X1   g15208(.A1(new_n15400_), .A2(new_n15393_), .B(new_n2641_), .ZN(new_n15401_));
  INV_X1     g15209(.I(new_n14861_), .ZN(new_n15402_));
  NOR2_X1    g15210(.A1(new_n14860_), .A2(new_n14868_), .ZN(new_n15403_));
  NOR3_X1    g15211(.A1(new_n15402_), .A2(new_n15403_), .A3(new_n14867_), .ZN(new_n15404_));
  NOR3_X1    g15212(.A1(new_n15067_), .A2(new_n15402_), .A3(new_n15403_), .ZN(new_n15405_));
  INV_X1     g15213(.I(new_n15405_), .ZN(new_n15406_));
  AOI22_X1   g15214(.A1(new_n15406_), .A2(new_n14867_), .B1(\asqrt[15] ), .B2(new_n15404_), .ZN(new_n15407_));
  OAI21_X1   g15215(.A1(new_n15390_), .A2(new_n15391_), .B(new_n15382_), .ZN(new_n15408_));
  AOI21_X1   g15216(.A1(new_n15408_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n15409_));
  AOI21_X1   g15217(.A1(new_n15409_), .A2(new_n15400_), .B(new_n15407_), .ZN(new_n15410_));
  OAI21_X1   g15218(.A1(new_n15410_), .A2(new_n15401_), .B(\asqrt[46] ), .ZN(new_n15411_));
  INV_X1     g15219(.I(new_n15411_), .ZN(new_n15412_));
  INV_X1     g15220(.I(new_n14875_), .ZN(new_n15413_));
  INV_X1     g15221(.I(new_n14869_), .ZN(new_n15414_));
  INV_X1     g15222(.I(new_n14877_), .ZN(new_n15415_));
  NOR2_X1    g15223(.A1(new_n15415_), .A2(new_n15414_), .ZN(new_n15416_));
  NOR3_X1    g15224(.A1(new_n15067_), .A2(new_n14870_), .A3(new_n15416_), .ZN(new_n15417_));
  INV_X1     g15225(.I(new_n15417_), .ZN(new_n15418_));
  NOR3_X1    g15226(.A1(new_n15416_), .A2(new_n14870_), .A3(new_n15413_), .ZN(new_n15419_));
  AOI22_X1   g15227(.A1(new_n15418_), .A2(new_n15413_), .B1(\asqrt[15] ), .B2(new_n15419_), .ZN(new_n15420_));
  NOR3_X1    g15228(.A1(new_n15410_), .A2(new_n15401_), .A3(\asqrt[46] ), .ZN(new_n15421_));
  NOR2_X1    g15229(.A1(new_n15421_), .A2(new_n15420_), .ZN(new_n15422_));
  OAI21_X1   g15230(.A1(new_n15422_), .A2(new_n15412_), .B(\asqrt[47] ), .ZN(new_n15423_));
  NOR3_X1    g15231(.A1(new_n14880_), .A2(new_n15085_), .A3(new_n14885_), .ZN(new_n15424_));
  NOR3_X1    g15232(.A1(new_n15067_), .A2(new_n14880_), .A3(new_n14885_), .ZN(new_n15425_));
  INV_X1     g15233(.I(new_n15425_), .ZN(new_n15426_));
  AOI22_X1   g15234(.A1(new_n15426_), .A2(new_n15085_), .B1(\asqrt[15] ), .B2(new_n15424_), .ZN(new_n15427_));
  INV_X1     g15235(.I(new_n15427_), .ZN(new_n15428_));
  NAND2_X1   g15236(.A1(new_n15411_), .A2(new_n2229_), .ZN(new_n15429_));
  OAI21_X1   g15237(.A1(new_n15422_), .A2(new_n15429_), .B(new_n15428_), .ZN(new_n15430_));
  AOI21_X1   g15238(.A1(new_n15430_), .A2(new_n15423_), .B(new_n1956_), .ZN(new_n15431_));
  INV_X1     g15239(.I(new_n14887_), .ZN(new_n15432_));
  NOR2_X1    g15240(.A1(new_n14886_), .A2(new_n14894_), .ZN(new_n15433_));
  NOR3_X1    g15241(.A1(new_n15067_), .A2(new_n15432_), .A3(new_n15433_), .ZN(new_n15434_));
  INV_X1     g15242(.I(new_n15434_), .ZN(new_n15435_));
  NOR3_X1    g15243(.A1(new_n15432_), .A2(new_n15433_), .A3(new_n14893_), .ZN(new_n15436_));
  AOI22_X1   g15244(.A1(new_n15435_), .A2(new_n14893_), .B1(\asqrt[15] ), .B2(new_n15436_), .ZN(new_n15437_));
  OAI21_X1   g15245(.A1(new_n15420_), .A2(new_n15421_), .B(new_n15411_), .ZN(new_n15438_));
  AOI21_X1   g15246(.A1(new_n15438_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n15439_));
  AOI21_X1   g15247(.A1(new_n15439_), .A2(new_n15430_), .B(new_n15437_), .ZN(new_n15440_));
  OAI21_X1   g15248(.A1(new_n15440_), .A2(new_n15431_), .B(\asqrt[49] ), .ZN(new_n15441_));
  INV_X1     g15249(.I(new_n15441_), .ZN(new_n15442_));
  INV_X1     g15250(.I(new_n14901_), .ZN(new_n15443_));
  INV_X1     g15251(.I(new_n14895_), .ZN(new_n15444_));
  INV_X1     g15252(.I(new_n14903_), .ZN(new_n15445_));
  NOR2_X1    g15253(.A1(new_n15445_), .A2(new_n15444_), .ZN(new_n15446_));
  NOR3_X1    g15254(.A1(new_n15446_), .A2(new_n14896_), .A3(new_n15443_), .ZN(new_n15447_));
  NOR3_X1    g15255(.A1(new_n15067_), .A2(new_n14896_), .A3(new_n15446_), .ZN(new_n15448_));
  INV_X1     g15256(.I(new_n15448_), .ZN(new_n15449_));
  AOI22_X1   g15257(.A1(new_n15449_), .A2(new_n15443_), .B1(\asqrt[15] ), .B2(new_n15447_), .ZN(new_n15450_));
  NOR3_X1    g15258(.A1(new_n15440_), .A2(new_n15431_), .A3(\asqrt[49] ), .ZN(new_n15451_));
  NOR2_X1    g15259(.A1(new_n15451_), .A2(new_n15450_), .ZN(new_n15452_));
  OAI21_X1   g15260(.A1(new_n15452_), .A2(new_n15442_), .B(\asqrt[50] ), .ZN(new_n15453_));
  NOR3_X1    g15261(.A1(new_n15067_), .A2(new_n14906_), .A3(new_n14911_), .ZN(new_n15454_));
  INV_X1     g15262(.I(new_n15454_), .ZN(new_n15455_));
  NOR3_X1    g15263(.A1(new_n14906_), .A2(new_n15084_), .A3(new_n14911_), .ZN(new_n15456_));
  AOI22_X1   g15264(.A1(new_n15455_), .A2(new_n15084_), .B1(\asqrt[15] ), .B2(new_n15456_), .ZN(new_n15457_));
  INV_X1     g15265(.I(new_n15457_), .ZN(new_n15458_));
  NAND2_X1   g15266(.A1(new_n15441_), .A2(new_n1612_), .ZN(new_n15459_));
  OAI21_X1   g15267(.A1(new_n15452_), .A2(new_n15459_), .B(new_n15458_), .ZN(new_n15460_));
  AOI21_X1   g15268(.A1(new_n15460_), .A2(new_n15453_), .B(new_n1376_), .ZN(new_n15461_));
  INV_X1     g15269(.I(new_n14913_), .ZN(new_n15462_));
  NOR2_X1    g15270(.A1(new_n14912_), .A2(new_n14920_), .ZN(new_n15463_));
  NOR3_X1    g15271(.A1(new_n15462_), .A2(new_n14919_), .A3(new_n15463_), .ZN(new_n15464_));
  NOR3_X1    g15272(.A1(new_n15067_), .A2(new_n15462_), .A3(new_n15463_), .ZN(new_n15465_));
  INV_X1     g15273(.I(new_n15465_), .ZN(new_n15466_));
  AOI22_X1   g15274(.A1(new_n15466_), .A2(new_n14919_), .B1(\asqrt[15] ), .B2(new_n15464_), .ZN(new_n15467_));
  OAI21_X1   g15275(.A1(new_n15450_), .A2(new_n15451_), .B(new_n15441_), .ZN(new_n15468_));
  AOI21_X1   g15276(.A1(new_n15468_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n15469_));
  AOI21_X1   g15277(.A1(new_n15469_), .A2(new_n15460_), .B(new_n15467_), .ZN(new_n15470_));
  OAI21_X1   g15278(.A1(new_n15470_), .A2(new_n15461_), .B(\asqrt[52] ), .ZN(new_n15471_));
  INV_X1     g15279(.I(new_n15471_), .ZN(new_n15472_));
  INV_X1     g15280(.I(new_n14927_), .ZN(new_n15473_));
  INV_X1     g15281(.I(new_n14921_), .ZN(new_n15474_));
  INV_X1     g15282(.I(new_n14929_), .ZN(new_n15475_));
  NOR2_X1    g15283(.A1(new_n15475_), .A2(new_n15474_), .ZN(new_n15476_));
  NOR3_X1    g15284(.A1(new_n15067_), .A2(new_n14922_), .A3(new_n15476_), .ZN(new_n15477_));
  INV_X1     g15285(.I(new_n15477_), .ZN(new_n15478_));
  NOR3_X1    g15286(.A1(new_n15476_), .A2(new_n14922_), .A3(new_n15473_), .ZN(new_n15479_));
  AOI22_X1   g15287(.A1(new_n15478_), .A2(new_n15473_), .B1(\asqrt[15] ), .B2(new_n15479_), .ZN(new_n15480_));
  NOR3_X1    g15288(.A1(new_n15470_), .A2(new_n15461_), .A3(\asqrt[52] ), .ZN(new_n15481_));
  NOR2_X1    g15289(.A1(new_n15481_), .A2(new_n15480_), .ZN(new_n15482_));
  OAI21_X1   g15290(.A1(new_n15482_), .A2(new_n15472_), .B(\asqrt[53] ), .ZN(new_n15483_));
  NOR3_X1    g15291(.A1(new_n14932_), .A2(new_n15083_), .A3(new_n14974_), .ZN(new_n15484_));
  NOR3_X1    g15292(.A1(new_n15067_), .A2(new_n14932_), .A3(new_n14974_), .ZN(new_n15485_));
  INV_X1     g15293(.I(new_n15485_), .ZN(new_n15486_));
  AOI22_X1   g15294(.A1(new_n15486_), .A2(new_n15083_), .B1(\asqrt[15] ), .B2(new_n15484_), .ZN(new_n15487_));
  INV_X1     g15295(.I(new_n15487_), .ZN(new_n15488_));
  NAND2_X1   g15296(.A1(new_n15471_), .A2(new_n1103_), .ZN(new_n15489_));
  OAI21_X1   g15297(.A1(new_n15482_), .A2(new_n15489_), .B(new_n15488_), .ZN(new_n15490_));
  AOI21_X1   g15298(.A1(new_n15490_), .A2(new_n15483_), .B(new_n904_), .ZN(new_n15491_));
  INV_X1     g15299(.I(new_n14940_), .ZN(new_n15492_));
  NOR2_X1    g15300(.A1(new_n14947_), .A2(new_n14939_), .ZN(new_n15493_));
  NOR3_X1    g15301(.A1(new_n15067_), .A2(new_n15492_), .A3(new_n15493_), .ZN(new_n15494_));
  INV_X1     g15302(.I(new_n15494_), .ZN(new_n15495_));
  NOR3_X1    g15303(.A1(new_n15492_), .A2(new_n14946_), .A3(new_n15493_), .ZN(new_n15496_));
  AOI22_X1   g15304(.A1(new_n15495_), .A2(new_n14946_), .B1(\asqrt[15] ), .B2(new_n15496_), .ZN(new_n15497_));
  OAI21_X1   g15305(.A1(new_n15480_), .A2(new_n15481_), .B(new_n15471_), .ZN(new_n15498_));
  AOI21_X1   g15306(.A1(new_n15498_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n15499_));
  AOI21_X1   g15307(.A1(new_n15499_), .A2(new_n15490_), .B(new_n15497_), .ZN(new_n15500_));
  OAI21_X1   g15308(.A1(new_n15500_), .A2(new_n15491_), .B(\asqrt[55] ), .ZN(new_n15501_));
  INV_X1     g15309(.I(new_n15501_), .ZN(new_n15502_));
  NOR2_X1    g15310(.A1(new_n14958_), .A2(new_n14951_), .ZN(new_n15503_));
  NOR3_X1    g15311(.A1(new_n15503_), .A2(new_n14949_), .A3(new_n14957_), .ZN(new_n15504_));
  NOR3_X1    g15312(.A1(new_n15067_), .A2(new_n14949_), .A3(new_n15503_), .ZN(new_n15505_));
  INV_X1     g15313(.I(new_n15505_), .ZN(new_n15506_));
  AOI22_X1   g15314(.A1(new_n15506_), .A2(new_n14957_), .B1(\asqrt[15] ), .B2(new_n15504_), .ZN(new_n15507_));
  NOR3_X1    g15315(.A1(new_n15500_), .A2(new_n15491_), .A3(\asqrt[55] ), .ZN(new_n15508_));
  NOR2_X1    g15316(.A1(new_n15508_), .A2(new_n15507_), .ZN(new_n15509_));
  OAI21_X1   g15317(.A1(new_n15509_), .A2(new_n15502_), .B(\asqrt[56] ), .ZN(new_n15510_));
  NOR3_X1    g15318(.A1(new_n15067_), .A2(new_n14960_), .A3(new_n15006_), .ZN(new_n15511_));
  INV_X1     g15319(.I(new_n15511_), .ZN(new_n15512_));
  NOR3_X1    g15320(.A1(new_n14960_), .A2(new_n15082_), .A3(new_n15006_), .ZN(new_n15513_));
  AOI22_X1   g15321(.A1(new_n15512_), .A2(new_n15082_), .B1(\asqrt[15] ), .B2(new_n15513_), .ZN(new_n15514_));
  INV_X1     g15322(.I(new_n15514_), .ZN(new_n15515_));
  NAND2_X1   g15323(.A1(new_n15501_), .A2(new_n703_), .ZN(new_n15516_));
  OAI21_X1   g15324(.A1(new_n15509_), .A2(new_n15516_), .B(new_n15515_), .ZN(new_n15517_));
  AOI21_X1   g15325(.A1(new_n15517_), .A2(new_n15510_), .B(new_n531_), .ZN(new_n15518_));
  INV_X1     g15326(.I(new_n14967_), .ZN(new_n15519_));
  NOR2_X1    g15327(.A1(new_n14979_), .A2(new_n14966_), .ZN(new_n15520_));
  NOR3_X1    g15328(.A1(new_n15519_), .A2(new_n14973_), .A3(new_n15520_), .ZN(new_n15521_));
  NOR3_X1    g15329(.A1(new_n15067_), .A2(new_n15519_), .A3(new_n15520_), .ZN(new_n15522_));
  INV_X1     g15330(.I(new_n15522_), .ZN(new_n15523_));
  AOI22_X1   g15331(.A1(new_n15523_), .A2(new_n14973_), .B1(\asqrt[15] ), .B2(new_n15521_), .ZN(new_n15524_));
  OAI21_X1   g15332(.A1(new_n15507_), .A2(new_n15508_), .B(new_n15501_), .ZN(new_n15525_));
  AOI21_X1   g15333(.A1(new_n15525_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n15526_));
  AOI21_X1   g15334(.A1(new_n15526_), .A2(new_n15517_), .B(new_n15524_), .ZN(new_n15527_));
  OAI21_X1   g15335(.A1(new_n15527_), .A2(new_n15518_), .B(\asqrt[58] ), .ZN(new_n15528_));
  NOR2_X1    g15336(.A1(new_n14990_), .A2(new_n14983_), .ZN(new_n15529_));
  NOR3_X1    g15337(.A1(new_n15067_), .A2(new_n14981_), .A3(new_n15529_), .ZN(new_n15530_));
  INV_X1     g15338(.I(new_n15530_), .ZN(new_n15531_));
  NOR3_X1    g15339(.A1(new_n15529_), .A2(new_n14981_), .A3(new_n14989_), .ZN(new_n15532_));
  AOI22_X1   g15340(.A1(new_n15531_), .A2(new_n14989_), .B1(\asqrt[15] ), .B2(new_n15532_), .ZN(new_n15533_));
  INV_X1     g15341(.I(new_n15533_), .ZN(new_n15534_));
  INV_X1     g15342(.I(new_n15507_), .ZN(new_n15535_));
  INV_X1     g15343(.I(new_n15480_), .ZN(new_n15536_));
  INV_X1     g15344(.I(new_n15450_), .ZN(new_n15537_));
  INV_X1     g15345(.I(new_n15420_), .ZN(new_n15538_));
  INV_X1     g15346(.I(new_n15390_), .ZN(new_n15539_));
  INV_X1     g15347(.I(new_n15362_), .ZN(new_n15540_));
  INV_X1     g15348(.I(new_n15336_), .ZN(new_n15541_));
  INV_X1     g15349(.I(new_n15309_), .ZN(new_n15542_));
  INV_X1     g15350(.I(new_n15282_), .ZN(new_n15543_));
  INV_X1     g15351(.I(new_n15255_), .ZN(new_n15544_));
  INV_X1     g15352(.I(new_n15224_), .ZN(new_n15545_));
  INV_X1     g15353(.I(new_n15198_), .ZN(new_n15546_));
  NAND2_X1   g15354(.A1(new_n15140_), .A2(new_n12913_), .ZN(new_n15547_));
  OAI21_X1   g15355(.A1(new_n15547_), .A2(new_n15172_), .B(new_n15154_), .ZN(new_n15548_));
  AOI21_X1   g15356(.A1(new_n15548_), .A2(new_n15182_), .B(new_n12364_), .ZN(new_n15549_));
  NOR2_X1    g15357(.A1(new_n15148_), .A2(\asqrt[20] ), .ZN(new_n15550_));
  AOI21_X1   g15358(.A1(new_n15550_), .A2(new_n15548_), .B(new_n15180_), .ZN(new_n15551_));
  OAI21_X1   g15359(.A1(new_n15551_), .A2(new_n15549_), .B(\asqrt[21] ), .ZN(new_n15552_));
  NAND2_X1   g15360(.A1(new_n15552_), .A2(new_n11326_), .ZN(new_n15553_));
  OAI21_X1   g15361(.A1(new_n15553_), .A2(new_n15192_), .B(new_n15546_), .ZN(new_n15554_));
  NAND3_X1   g15362(.A1(new_n15554_), .A2(new_n10812_), .A3(new_n15193_), .ZN(new_n15555_));
  AOI22_X1   g15363(.A1(new_n15555_), .A2(new_n15207_), .B1(\asqrt[23] ), .B2(new_n15215_), .ZN(new_n15556_));
  OAI21_X1   g15364(.A1(new_n15556_), .A2(new_n10221_), .B(new_n9846_), .ZN(new_n15557_));
  OAI21_X1   g15365(.A1(new_n15557_), .A2(new_n15217_), .B(new_n15545_), .ZN(new_n15558_));
  AOI21_X1   g15366(.A1(new_n15558_), .A2(new_n15218_), .B(new_n9317_), .ZN(new_n15559_));
  AOI21_X1   g15367(.A1(new_n15554_), .A2(new_n15193_), .B(new_n10812_), .ZN(new_n15560_));
  NOR3_X1    g15368(.A1(new_n15551_), .A2(new_n15549_), .A3(\asqrt[21] ), .ZN(new_n15561_));
  OAI21_X1   g15369(.A1(new_n15189_), .A2(new_n15561_), .B(new_n15552_), .ZN(new_n15562_));
  AOI21_X1   g15370(.A1(new_n15562_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n15563_));
  AOI21_X1   g15371(.A1(new_n15563_), .A2(new_n15554_), .B(new_n15206_), .ZN(new_n15564_));
  NOR3_X1    g15372(.A1(new_n15564_), .A2(\asqrt[24] ), .A3(new_n15560_), .ZN(new_n15565_));
  OAI22_X1   g15373(.A1(new_n15565_), .A2(new_n15214_), .B1(new_n15556_), .B2(new_n10221_), .ZN(new_n15566_));
  AOI21_X1   g15374(.A1(new_n15566_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n15567_));
  AOI21_X1   g15375(.A1(new_n15567_), .A2(new_n15558_), .B(new_n15232_), .ZN(new_n15568_));
  OAI21_X1   g15376(.A1(new_n15568_), .A2(new_n15559_), .B(\asqrt[27] ), .ZN(new_n15569_));
  NAND2_X1   g15377(.A1(new_n15569_), .A2(new_n8483_), .ZN(new_n15570_));
  OAI21_X1   g15378(.A1(new_n15570_), .A2(new_n15245_), .B(new_n15544_), .ZN(new_n15571_));
  AOI21_X1   g15379(.A1(new_n15571_), .A2(new_n15246_), .B(new_n8036_), .ZN(new_n15572_));
  NOR3_X1    g15380(.A1(new_n15568_), .A2(\asqrt[27] ), .A3(new_n15559_), .ZN(new_n15573_));
  OAI21_X1   g15381(.A1(new_n15242_), .A2(new_n15573_), .B(new_n15569_), .ZN(new_n15574_));
  AOI21_X1   g15382(.A1(new_n15574_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n15575_));
  AOI21_X1   g15383(.A1(new_n15575_), .A2(new_n15571_), .B(new_n15263_), .ZN(new_n15576_));
  OAI21_X1   g15384(.A1(new_n15576_), .A2(new_n15572_), .B(\asqrt[30] ), .ZN(new_n15577_));
  NAND2_X1   g15385(.A1(new_n15577_), .A2(new_n7229_), .ZN(new_n15578_));
  OAI21_X1   g15386(.A1(new_n15578_), .A2(new_n15275_), .B(new_n15543_), .ZN(new_n15579_));
  AOI21_X1   g15387(.A1(new_n15579_), .A2(new_n15276_), .B(new_n6824_), .ZN(new_n15580_));
  NOR3_X1    g15388(.A1(new_n15576_), .A2(\asqrt[30] ), .A3(new_n15572_), .ZN(new_n15581_));
  OAI21_X1   g15389(.A1(new_n15272_), .A2(new_n15581_), .B(new_n15577_), .ZN(new_n15582_));
  AOI21_X1   g15390(.A1(new_n15582_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n15583_));
  AOI21_X1   g15391(.A1(new_n15583_), .A2(new_n15579_), .B(new_n15290_), .ZN(new_n15584_));
  OAI21_X1   g15392(.A1(new_n15584_), .A2(new_n15580_), .B(\asqrt[33] ), .ZN(new_n15585_));
  NAND2_X1   g15393(.A1(new_n15585_), .A2(new_n6077_), .ZN(new_n15586_));
  OAI21_X1   g15394(.A1(new_n15586_), .A2(new_n15302_), .B(new_n15542_), .ZN(new_n15587_));
  AOI21_X1   g15395(.A1(new_n15587_), .A2(new_n15303_), .B(new_n5708_), .ZN(new_n15588_));
  NOR3_X1    g15396(.A1(new_n15584_), .A2(\asqrt[33] ), .A3(new_n15580_), .ZN(new_n15589_));
  OAI21_X1   g15397(.A1(new_n15299_), .A2(new_n15589_), .B(new_n15585_), .ZN(new_n15590_));
  AOI21_X1   g15398(.A1(new_n15590_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n15591_));
  AOI21_X1   g15399(.A1(new_n15591_), .A2(new_n15587_), .B(new_n15317_), .ZN(new_n15592_));
  OAI21_X1   g15400(.A1(new_n15592_), .A2(new_n15588_), .B(\asqrt[36] ), .ZN(new_n15593_));
  NAND2_X1   g15401(.A1(new_n15593_), .A2(new_n5024_), .ZN(new_n15594_));
  OAI21_X1   g15402(.A1(new_n15594_), .A2(new_n15329_), .B(new_n15541_), .ZN(new_n15595_));
  AOI21_X1   g15403(.A1(new_n15595_), .A2(new_n15330_), .B(new_n4696_), .ZN(new_n15596_));
  NOR3_X1    g15404(.A1(new_n15592_), .A2(\asqrt[36] ), .A3(new_n15588_), .ZN(new_n15597_));
  OAI21_X1   g15405(.A1(new_n15326_), .A2(new_n15597_), .B(new_n15593_), .ZN(new_n15598_));
  AOI21_X1   g15406(.A1(new_n15598_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n15599_));
  AOI21_X1   g15407(.A1(new_n15599_), .A2(new_n15595_), .B(new_n15344_), .ZN(new_n15600_));
  OAI21_X1   g15408(.A1(new_n15600_), .A2(new_n15596_), .B(\asqrt[39] ), .ZN(new_n15601_));
  NAND2_X1   g15409(.A1(new_n15601_), .A2(new_n4071_), .ZN(new_n15602_));
  OAI21_X1   g15410(.A1(new_n15602_), .A2(new_n15355_), .B(new_n15540_), .ZN(new_n15603_));
  AOI21_X1   g15411(.A1(new_n15603_), .A2(new_n15356_), .B(new_n3782_), .ZN(new_n15604_));
  NOR3_X1    g15412(.A1(new_n15600_), .A2(\asqrt[39] ), .A3(new_n15596_), .ZN(new_n15605_));
  OAI21_X1   g15413(.A1(new_n15352_), .A2(new_n15605_), .B(new_n15601_), .ZN(new_n15606_));
  AOI21_X1   g15414(.A1(new_n15606_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n15607_));
  AOI21_X1   g15415(.A1(new_n15607_), .A2(new_n15603_), .B(new_n15370_), .ZN(new_n15608_));
  OAI21_X1   g15416(.A1(new_n15608_), .A2(new_n15604_), .B(\asqrt[42] ), .ZN(new_n15609_));
  NAND2_X1   g15417(.A1(new_n15609_), .A2(new_n3218_), .ZN(new_n15610_));
  OAI21_X1   g15418(.A1(new_n15610_), .A2(new_n15381_), .B(new_n15539_), .ZN(new_n15611_));
  AOI21_X1   g15419(.A1(new_n15611_), .A2(new_n15382_), .B(new_n2954_), .ZN(new_n15612_));
  NOR3_X1    g15420(.A1(new_n15608_), .A2(\asqrt[42] ), .A3(new_n15604_), .ZN(new_n15613_));
  OAI21_X1   g15421(.A1(new_n15378_), .A2(new_n15613_), .B(new_n15609_), .ZN(new_n15614_));
  AOI21_X1   g15422(.A1(new_n15614_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n15615_));
  AOI21_X1   g15423(.A1(new_n15615_), .A2(new_n15611_), .B(new_n15397_), .ZN(new_n15616_));
  OAI21_X1   g15424(.A1(new_n15616_), .A2(new_n15612_), .B(\asqrt[45] ), .ZN(new_n15617_));
  NAND2_X1   g15425(.A1(new_n15617_), .A2(new_n2465_), .ZN(new_n15618_));
  OAI21_X1   g15426(.A1(new_n15618_), .A2(new_n15410_), .B(new_n15538_), .ZN(new_n15619_));
  AOI21_X1   g15427(.A1(new_n15619_), .A2(new_n15411_), .B(new_n2229_), .ZN(new_n15620_));
  NOR3_X1    g15428(.A1(new_n15616_), .A2(\asqrt[45] ), .A3(new_n15612_), .ZN(new_n15621_));
  OAI21_X1   g15429(.A1(new_n15407_), .A2(new_n15621_), .B(new_n15617_), .ZN(new_n15622_));
  AOI21_X1   g15430(.A1(new_n15622_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n15623_));
  AOI21_X1   g15431(.A1(new_n15623_), .A2(new_n15619_), .B(new_n15427_), .ZN(new_n15624_));
  OAI21_X1   g15432(.A1(new_n15624_), .A2(new_n15620_), .B(\asqrt[48] ), .ZN(new_n15625_));
  NAND2_X1   g15433(.A1(new_n15625_), .A2(new_n1806_), .ZN(new_n15626_));
  OAI21_X1   g15434(.A1(new_n15626_), .A2(new_n15440_), .B(new_n15537_), .ZN(new_n15627_));
  AOI21_X1   g15435(.A1(new_n15627_), .A2(new_n15441_), .B(new_n1612_), .ZN(new_n15628_));
  NOR3_X1    g15436(.A1(new_n15624_), .A2(\asqrt[48] ), .A3(new_n15620_), .ZN(new_n15629_));
  OAI21_X1   g15437(.A1(new_n15437_), .A2(new_n15629_), .B(new_n15625_), .ZN(new_n15630_));
  AOI21_X1   g15438(.A1(new_n15630_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n15631_));
  AOI21_X1   g15439(.A1(new_n15631_), .A2(new_n15627_), .B(new_n15457_), .ZN(new_n15632_));
  OAI21_X1   g15440(.A1(new_n15632_), .A2(new_n15628_), .B(\asqrt[51] ), .ZN(new_n15633_));
  NAND2_X1   g15441(.A1(new_n15633_), .A2(new_n1256_), .ZN(new_n15634_));
  OAI21_X1   g15442(.A1(new_n15634_), .A2(new_n15470_), .B(new_n15536_), .ZN(new_n15635_));
  NAND3_X1   g15443(.A1(new_n15635_), .A2(new_n1103_), .A3(new_n15471_), .ZN(new_n15636_));
  AOI22_X1   g15444(.A1(new_n15636_), .A2(new_n15488_), .B1(\asqrt[53] ), .B2(new_n15498_), .ZN(new_n15637_));
  OAI21_X1   g15445(.A1(new_n15637_), .A2(new_n904_), .B(new_n823_), .ZN(new_n15638_));
  OAI21_X1   g15446(.A1(new_n15638_), .A2(new_n15500_), .B(new_n15535_), .ZN(new_n15639_));
  NAND3_X1   g15447(.A1(new_n15639_), .A2(new_n703_), .A3(new_n15501_), .ZN(new_n15640_));
  AOI22_X1   g15448(.A1(new_n15640_), .A2(new_n15515_), .B1(\asqrt[56] ), .B2(new_n15525_), .ZN(new_n15641_));
  OAI21_X1   g15449(.A1(new_n15641_), .A2(new_n531_), .B(new_n436_), .ZN(new_n15642_));
  OAI21_X1   g15450(.A1(new_n15642_), .A2(new_n15527_), .B(new_n15534_), .ZN(new_n15643_));
  AOI21_X1   g15451(.A1(new_n15643_), .A2(new_n15528_), .B(new_n327_), .ZN(new_n15644_));
  NOR3_X1    g15452(.A1(new_n14992_), .A2(new_n15081_), .A3(new_n15038_), .ZN(new_n15645_));
  NOR3_X1    g15453(.A1(new_n15067_), .A2(new_n14992_), .A3(new_n15038_), .ZN(new_n15646_));
  INV_X1     g15454(.I(new_n15646_), .ZN(new_n15647_));
  AOI22_X1   g15455(.A1(new_n15647_), .A2(new_n15081_), .B1(\asqrt[15] ), .B2(new_n15645_), .ZN(new_n15648_));
  NAND2_X1   g15456(.A1(new_n15528_), .A2(new_n327_), .ZN(new_n15649_));
  INV_X1     g15457(.I(new_n15649_), .ZN(new_n15650_));
  AOI21_X1   g15458(.A1(new_n15650_), .A2(new_n15643_), .B(new_n15648_), .ZN(new_n15651_));
  OAI21_X1   g15459(.A1(new_n15651_), .A2(new_n15644_), .B(\asqrt[60] ), .ZN(new_n15652_));
  INV_X1     g15460(.I(new_n14999_), .ZN(new_n15653_));
  NOR2_X1    g15461(.A1(new_n15011_), .A2(new_n14998_), .ZN(new_n15654_));
  NOR3_X1    g15462(.A1(new_n15067_), .A2(new_n15653_), .A3(new_n15654_), .ZN(new_n15655_));
  INV_X1     g15463(.I(new_n15655_), .ZN(new_n15656_));
  NOR3_X1    g15464(.A1(new_n15653_), .A2(new_n15005_), .A3(new_n15654_), .ZN(new_n15657_));
  AOI22_X1   g15465(.A1(new_n15656_), .A2(new_n15005_), .B1(\asqrt[15] ), .B2(new_n15657_), .ZN(new_n15658_));
  INV_X1     g15466(.I(new_n15658_), .ZN(new_n15659_));
  INV_X1     g15467(.I(new_n15528_), .ZN(new_n15660_));
  NOR3_X1    g15468(.A1(new_n15527_), .A2(new_n15518_), .A3(\asqrt[58] ), .ZN(new_n15661_));
  NOR2_X1    g15469(.A1(new_n15661_), .A2(new_n15533_), .ZN(new_n15662_));
  OAI21_X1   g15470(.A1(new_n15662_), .A2(new_n15660_), .B(\asqrt[59] ), .ZN(new_n15663_));
  NAND2_X1   g15471(.A1(new_n15663_), .A2(new_n306_), .ZN(new_n15664_));
  OAI21_X1   g15472(.A1(new_n15664_), .A2(new_n15651_), .B(new_n15659_), .ZN(new_n15665_));
  AOI21_X1   g15473(.A1(new_n15665_), .A2(new_n15652_), .B(new_n218_), .ZN(new_n15666_));
  NOR2_X1    g15474(.A1(new_n15015_), .A2(new_n15022_), .ZN(new_n15667_));
  NOR3_X1    g15475(.A1(new_n15667_), .A2(new_n15013_), .A3(new_n15021_), .ZN(new_n15668_));
  NOR3_X1    g15476(.A1(new_n15067_), .A2(new_n15013_), .A3(new_n15667_), .ZN(new_n15669_));
  INV_X1     g15477(.I(new_n15669_), .ZN(new_n15670_));
  AOI22_X1   g15478(.A1(new_n15670_), .A2(new_n15021_), .B1(\asqrt[15] ), .B2(new_n15668_), .ZN(new_n15671_));
  INV_X1     g15479(.I(new_n15648_), .ZN(new_n15672_));
  OAI21_X1   g15480(.A1(new_n15662_), .A2(new_n15649_), .B(new_n15672_), .ZN(new_n15673_));
  AOI21_X1   g15481(.A1(new_n15673_), .A2(new_n15663_), .B(new_n306_), .ZN(new_n15674_));
  NOR2_X1    g15482(.A1(new_n15674_), .A2(\asqrt[61] ), .ZN(new_n15675_));
  AOI21_X1   g15483(.A1(new_n15675_), .A2(new_n15665_), .B(new_n15671_), .ZN(new_n15676_));
  OAI21_X1   g15484(.A1(new_n15676_), .A2(new_n15666_), .B(\asqrt[62] ), .ZN(new_n15677_));
  NOR3_X1    g15485(.A1(new_n15067_), .A2(new_n15024_), .A3(new_n15078_), .ZN(new_n15678_));
  INV_X1     g15486(.I(new_n15678_), .ZN(new_n15679_));
  NOR3_X1    g15487(.A1(new_n15024_), .A2(new_n15080_), .A3(new_n15078_), .ZN(new_n15680_));
  AOI22_X1   g15488(.A1(new_n15679_), .A2(new_n15080_), .B1(\asqrt[15] ), .B2(new_n15680_), .ZN(new_n15681_));
  INV_X1     g15489(.I(new_n15681_), .ZN(new_n15682_));
  OAI21_X1   g15490(.A1(new_n15533_), .A2(new_n15661_), .B(new_n15528_), .ZN(new_n15683_));
  AOI21_X1   g15491(.A1(new_n15683_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n15684_));
  AOI21_X1   g15492(.A1(new_n15684_), .A2(new_n15673_), .B(new_n15658_), .ZN(new_n15685_));
  OAI21_X1   g15493(.A1(new_n15685_), .A2(new_n15674_), .B(\asqrt[61] ), .ZN(new_n15686_));
  NAND2_X1   g15494(.A1(new_n15686_), .A2(new_n207_), .ZN(new_n15687_));
  OAI21_X1   g15495(.A1(new_n15687_), .A2(new_n15676_), .B(new_n15682_), .ZN(new_n15688_));
  NAND4_X1   g15496(.A1(\asqrt[15] ), .A2(new_n15031_), .A3(new_n15036_), .A4(new_n15117_), .ZN(new_n15689_));
  NAND2_X1   g15497(.A1(new_n15031_), .A2(new_n15117_), .ZN(new_n15690_));
  OAI21_X1   g15498(.A1(new_n15067_), .A2(new_n15690_), .B(new_n15037_), .ZN(new_n15691_));
  NAND2_X1   g15499(.A1(new_n15689_), .A2(new_n15691_), .ZN(new_n15692_));
  NOR2_X1    g15500(.A1(new_n15118_), .A2(new_n15057_), .ZN(new_n15693_));
  NAND2_X1   g15501(.A1(\asqrt[15] ), .A2(new_n15693_), .ZN(new_n15694_));
  NAND3_X1   g15502(.A1(new_n15692_), .A2(new_n15129_), .A3(new_n15694_), .ZN(new_n15695_));
  AOI21_X1   g15503(.A1(new_n15688_), .A2(new_n15677_), .B(new_n15695_), .ZN(new_n15696_));
  NOR3_X1    g15504(.A1(new_n15685_), .A2(new_n15674_), .A3(\asqrt[61] ), .ZN(new_n15697_));
  OAI21_X1   g15505(.A1(new_n15671_), .A2(new_n15697_), .B(new_n15686_), .ZN(new_n15698_));
  AOI21_X1   g15506(.A1(new_n15698_), .A2(\asqrt[62] ), .B(new_n15692_), .ZN(new_n15699_));
  OAI21_X1   g15507(.A1(new_n15067_), .A2(new_n15057_), .B(new_n15118_), .ZN(new_n15700_));
  NOR2_X1    g15508(.A1(new_n15693_), .A2(new_n193_), .ZN(new_n15701_));
  NAND2_X1   g15509(.A1(new_n15700_), .A2(new_n15701_), .ZN(new_n15702_));
  INV_X1     g15510(.I(new_n15702_), .ZN(new_n15703_));
  AND3_X2    g15511(.A1(new_n15048_), .A2(new_n15046_), .A3(new_n15063_), .Z(new_n15704_));
  NAND4_X1   g15512(.A1(new_n15119_), .A2(new_n15129_), .A3(new_n15060_), .A4(new_n15704_), .ZN(new_n15705_));
  INV_X1     g15513(.I(new_n15705_), .ZN(new_n15706_));
  NOR2_X1    g15514(.A1(new_n15703_), .A2(new_n15706_), .ZN(new_n15707_));
  INV_X1     g15515(.I(new_n15707_), .ZN(new_n15708_));
  AOI21_X1   g15516(.A1(new_n15699_), .A2(new_n15688_), .B(new_n15708_), .ZN(new_n15709_));
  OAI21_X1   g15517(.A1(\asqrt[63] ), .A2(new_n15696_), .B(new_n15709_), .ZN(\asqrt[14] ));
  NOR2_X1    g15518(.A1(\a[26] ), .A2(\a[27] ), .ZN(new_n15711_));
  INV_X1     g15519(.I(new_n15711_), .ZN(new_n15712_));
  NOR2_X1    g15520(.A1(new_n15712_), .A2(\a[28] ), .ZN(new_n15713_));
  INV_X1     g15521(.I(new_n15713_), .ZN(new_n15714_));
  NAND2_X1   g15522(.A1(new_n15688_), .A2(new_n15677_), .ZN(new_n15715_));
  INV_X1     g15523(.I(new_n15695_), .ZN(new_n15716_));
  AOI21_X1   g15524(.A1(new_n15715_), .A2(new_n15716_), .B(\asqrt[63] ), .ZN(new_n15717_));
  INV_X1     g15525(.I(new_n15671_), .ZN(new_n15718_));
  NAND3_X1   g15526(.A1(new_n15643_), .A2(new_n327_), .A3(new_n15528_), .ZN(new_n15719_));
  AOI22_X1   g15527(.A1(new_n15719_), .A2(new_n15672_), .B1(new_n15683_), .B2(\asqrt[59] ), .ZN(new_n15720_));
  OAI21_X1   g15528(.A1(new_n15720_), .A2(new_n306_), .B(new_n218_), .ZN(new_n15721_));
  OAI21_X1   g15529(.A1(new_n15721_), .A2(new_n15685_), .B(new_n15718_), .ZN(new_n15722_));
  NOR2_X1    g15530(.A1(new_n15666_), .A2(\asqrt[62] ), .ZN(new_n15723_));
  AOI21_X1   g15531(.A1(new_n15723_), .A2(new_n15722_), .B(new_n15681_), .ZN(new_n15724_));
  INV_X1     g15532(.I(new_n15692_), .ZN(new_n15725_));
  NAND2_X1   g15533(.A1(new_n15677_), .A2(new_n15725_), .ZN(new_n15726_));
  OAI21_X1   g15534(.A1(new_n15726_), .A2(new_n15724_), .B(new_n15707_), .ZN(new_n15727_));
  OAI21_X1   g15535(.A1(new_n15717_), .A2(new_n15727_), .B(\a[28] ), .ZN(new_n15728_));
  AOI21_X1   g15536(.A1(new_n15728_), .A2(new_n15714_), .B(new_n15067_), .ZN(new_n15729_));
  INV_X1     g15537(.I(\a[28] ), .ZN(new_n15730_));
  NAND3_X1   g15538(.A1(new_n15722_), .A2(new_n207_), .A3(new_n15686_), .ZN(new_n15731_));
  AOI22_X1   g15539(.A1(new_n15731_), .A2(new_n15682_), .B1(new_n15698_), .B2(\asqrt[62] ), .ZN(new_n15732_));
  OAI21_X1   g15540(.A1(new_n15732_), .A2(new_n15695_), .B(new_n193_), .ZN(new_n15733_));
  AOI21_X1   g15541(.A1(new_n15733_), .A2(new_n15709_), .B(new_n15730_), .ZN(new_n15734_));
  NAND4_X1   g15542(.A1(new_n15129_), .A2(new_n15060_), .A3(new_n15063_), .A4(new_n15714_), .ZN(new_n15735_));
  NOR2_X1    g15543(.A1(new_n15735_), .A2(new_n15055_), .ZN(new_n15736_));
  INV_X1     g15544(.I(new_n15736_), .ZN(new_n15737_));
  NOR2_X1    g15545(.A1(new_n15734_), .A2(new_n15737_), .ZN(new_n15738_));
  AOI21_X1   g15546(.A1(new_n15733_), .A2(new_n15709_), .B(new_n15070_), .ZN(new_n15739_));
  INV_X1     g15547(.I(\a[29] ), .ZN(new_n15740_));
  AOI21_X1   g15548(.A1(\asqrt[14] ), .A2(new_n15730_), .B(new_n15740_), .ZN(new_n15741_));
  NOR3_X1    g15549(.A1(new_n15738_), .A2(new_n15741_), .A3(new_n15739_), .ZN(new_n15742_));
  OAI21_X1   g15550(.A1(new_n15742_), .A2(new_n15729_), .B(\asqrt[16] ), .ZN(new_n15743_));
  OAI21_X1   g15551(.A1(new_n15717_), .A2(new_n15727_), .B(new_n15069_), .ZN(new_n15744_));
  NAND2_X1   g15552(.A1(new_n15699_), .A2(new_n15688_), .ZN(new_n15745_));
  NOR3_X1    g15553(.A1(new_n15703_), .A2(new_n15067_), .A3(new_n15706_), .ZN(new_n15746_));
  NAND3_X1   g15554(.A1(new_n15733_), .A2(new_n15745_), .A3(new_n15746_), .ZN(new_n15747_));
  AOI21_X1   g15555(.A1(new_n15747_), .A2(new_n15744_), .B(new_n15068_), .ZN(new_n15748_));
  NAND2_X1   g15556(.A1(new_n15745_), .A2(new_n15746_), .ZN(new_n15749_));
  NOR2_X1    g15557(.A1(new_n15749_), .A2(new_n15717_), .ZN(new_n15750_));
  NOR3_X1    g15558(.A1(new_n15750_), .A2(new_n15739_), .A3(\a[30] ), .ZN(new_n15751_));
  AOI21_X1   g15559(.A1(\asqrt[14] ), .A2(\a[28] ), .B(new_n15713_), .ZN(new_n15752_));
  OAI21_X1   g15560(.A1(new_n15752_), .A2(new_n15067_), .B(new_n14601_), .ZN(new_n15753_));
  OAI22_X1   g15561(.A1(new_n15742_), .A2(new_n15753_), .B1(new_n15748_), .B2(new_n15751_), .ZN(new_n15754_));
  AOI21_X1   g15562(.A1(new_n15754_), .A2(new_n15743_), .B(new_n14017_), .ZN(new_n15755_));
  NOR3_X1    g15563(.A1(new_n15158_), .A2(new_n15159_), .A3(new_n15124_), .ZN(new_n15756_));
  NAND3_X1   g15564(.A1(\asqrt[14] ), .A2(new_n15157_), .A3(new_n15077_), .ZN(new_n15757_));
  AOI22_X1   g15565(.A1(new_n15757_), .A2(new_n15124_), .B1(\asqrt[14] ), .B2(new_n15756_), .ZN(new_n15758_));
  OAI21_X1   g15566(.A1(new_n15734_), .A2(new_n15713_), .B(\asqrt[15] ), .ZN(new_n15759_));
  AOI21_X1   g15567(.A1(new_n15733_), .A2(new_n15709_), .B(\a[28] ), .ZN(new_n15760_));
  OAI21_X1   g15568(.A1(new_n15740_), .A2(new_n15760_), .B(new_n15744_), .ZN(new_n15761_));
  OAI21_X1   g15569(.A1(new_n15761_), .A2(new_n15738_), .B(new_n15759_), .ZN(new_n15762_));
  AOI21_X1   g15570(.A1(new_n15762_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n15763_));
  AOI21_X1   g15571(.A1(new_n15763_), .A2(new_n15754_), .B(new_n15758_), .ZN(new_n15764_));
  OAI21_X1   g15572(.A1(new_n15764_), .A2(new_n15755_), .B(\asqrt[18] ), .ZN(new_n15765_));
  INV_X1     g15573(.I(new_n15765_), .ZN(new_n15766_));
  NOR2_X1    g15574(.A1(new_n15162_), .A2(new_n15165_), .ZN(new_n15767_));
  INV_X1     g15575(.I(new_n15767_), .ZN(new_n15768_));
  NAND4_X1   g15576(.A1(\asqrt[14] ), .A2(new_n15163_), .A3(new_n15137_), .A4(new_n15768_), .ZN(new_n15769_));
  INV_X1     g15577(.I(\asqrt[14] ), .ZN(new_n15770_));
  NOR3_X1    g15578(.A1(new_n15770_), .A2(new_n15126_), .A3(new_n15767_), .ZN(new_n15771_));
  OAI21_X1   g15579(.A1(new_n15771_), .A2(new_n15137_), .B(new_n15769_), .ZN(new_n15772_));
  INV_X1     g15580(.I(new_n15772_), .ZN(new_n15773_));
  NOR3_X1    g15581(.A1(new_n15764_), .A2(new_n15755_), .A3(\asqrt[18] ), .ZN(new_n15774_));
  NOR2_X1    g15582(.A1(new_n15774_), .A2(new_n15773_), .ZN(new_n15775_));
  OAI21_X1   g15583(.A1(new_n15775_), .A2(new_n15766_), .B(\asqrt[19] ), .ZN(new_n15776_));
  NAND2_X1   g15584(.A1(new_n15171_), .A2(new_n15166_), .ZN(new_n15777_));
  NAND3_X1   g15585(.A1(\asqrt[14] ), .A2(new_n15140_), .A3(new_n15777_), .ZN(new_n15778_));
  AND3_X2    g15586(.A1(new_n15140_), .A2(new_n15144_), .A3(new_n15777_), .Z(new_n15779_));
  AOI22_X1   g15587(.A1(new_n15778_), .A2(new_n15145_), .B1(\asqrt[14] ), .B2(new_n15779_), .ZN(new_n15780_));
  INV_X1     g15588(.I(new_n15780_), .ZN(new_n15781_));
  NAND2_X1   g15589(.A1(new_n15765_), .A2(new_n12913_), .ZN(new_n15782_));
  OAI21_X1   g15590(.A1(new_n15775_), .A2(new_n15782_), .B(new_n15781_), .ZN(new_n15783_));
  AOI21_X1   g15591(.A1(new_n15783_), .A2(new_n15776_), .B(new_n12364_), .ZN(new_n15784_));
  NOR3_X1    g15592(.A1(new_n15148_), .A2(new_n15154_), .A3(new_n15173_), .ZN(new_n15785_));
  NOR3_X1    g15593(.A1(new_n15770_), .A2(new_n15148_), .A3(new_n15173_), .ZN(new_n15786_));
  INV_X1     g15594(.I(new_n15786_), .ZN(new_n15787_));
  AOI22_X1   g15595(.A1(new_n15787_), .A2(new_n15154_), .B1(\asqrt[14] ), .B2(new_n15785_), .ZN(new_n15788_));
  OAI21_X1   g15596(.A1(new_n15773_), .A2(new_n15774_), .B(new_n15765_), .ZN(new_n15789_));
  AOI21_X1   g15597(.A1(new_n15789_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n15790_));
  AOI21_X1   g15598(.A1(new_n15790_), .A2(new_n15783_), .B(new_n15788_), .ZN(new_n15791_));
  OAI21_X1   g15599(.A1(new_n15791_), .A2(new_n15784_), .B(\asqrt[21] ), .ZN(new_n15792_));
  INV_X1     g15600(.I(new_n15792_), .ZN(new_n15793_));
  NAND2_X1   g15601(.A1(new_n15550_), .A2(new_n15548_), .ZN(new_n15794_));
  NAND3_X1   g15602(.A1(\asqrt[14] ), .A2(new_n15175_), .A3(new_n15794_), .ZN(new_n15795_));
  AND3_X2    g15603(.A1(new_n15794_), .A2(new_n15175_), .A3(new_n15180_), .Z(new_n15796_));
  AOI22_X1   g15604(.A1(new_n15795_), .A2(new_n15181_), .B1(\asqrt[14] ), .B2(new_n15796_), .ZN(new_n15797_));
  NOR3_X1    g15605(.A1(new_n15791_), .A2(new_n15784_), .A3(\asqrt[21] ), .ZN(new_n15798_));
  NOR2_X1    g15606(.A1(new_n15798_), .A2(new_n15797_), .ZN(new_n15799_));
  OAI21_X1   g15607(.A1(new_n15799_), .A2(new_n15793_), .B(\asqrt[22] ), .ZN(new_n15800_));
  INV_X1     g15608(.I(new_n15189_), .ZN(new_n15801_));
  NOR3_X1    g15609(.A1(new_n15561_), .A2(new_n15185_), .A3(new_n15801_), .ZN(new_n15802_));
  NOR3_X1    g15610(.A1(new_n15770_), .A2(new_n15185_), .A3(new_n15561_), .ZN(new_n15803_));
  INV_X1     g15611(.I(new_n15803_), .ZN(new_n15804_));
  AOI22_X1   g15612(.A1(new_n15804_), .A2(new_n15801_), .B1(\asqrt[14] ), .B2(new_n15802_), .ZN(new_n15805_));
  INV_X1     g15613(.I(new_n15805_), .ZN(new_n15806_));
  NAND2_X1   g15614(.A1(new_n15792_), .A2(new_n11326_), .ZN(new_n15807_));
  OAI21_X1   g15615(.A1(new_n15799_), .A2(new_n15807_), .B(new_n15806_), .ZN(new_n15808_));
  AOI21_X1   g15616(.A1(new_n15808_), .A2(new_n15800_), .B(new_n10812_), .ZN(new_n15809_));
  NOR3_X1    g15617(.A1(new_n15770_), .A2(new_n15194_), .A3(new_n15199_), .ZN(new_n15810_));
  INV_X1     g15618(.I(new_n15810_), .ZN(new_n15811_));
  NOR3_X1    g15619(.A1(new_n15194_), .A2(new_n15546_), .A3(new_n15199_), .ZN(new_n15812_));
  AOI22_X1   g15620(.A1(new_n15811_), .A2(new_n15546_), .B1(\asqrt[14] ), .B2(new_n15812_), .ZN(new_n15813_));
  OAI21_X1   g15621(.A1(new_n15797_), .A2(new_n15798_), .B(new_n15792_), .ZN(new_n15814_));
  AOI21_X1   g15622(.A1(new_n15814_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n15815_));
  AOI21_X1   g15623(.A1(new_n15815_), .A2(new_n15808_), .B(new_n15813_), .ZN(new_n15816_));
  OAI21_X1   g15624(.A1(new_n15816_), .A2(new_n15809_), .B(\asqrt[24] ), .ZN(new_n15817_));
  INV_X1     g15625(.I(new_n15817_), .ZN(new_n15818_));
  INV_X1     g15626(.I(new_n15555_), .ZN(new_n15819_));
  NOR3_X1    g15627(.A1(new_n15819_), .A2(new_n15560_), .A3(new_n15207_), .ZN(new_n15820_));
  NOR3_X1    g15628(.A1(new_n15770_), .A2(new_n15560_), .A3(new_n15819_), .ZN(new_n15821_));
  INV_X1     g15629(.I(new_n15821_), .ZN(new_n15822_));
  AOI22_X1   g15630(.A1(new_n15822_), .A2(new_n15207_), .B1(\asqrt[14] ), .B2(new_n15820_), .ZN(new_n15823_));
  NOR3_X1    g15631(.A1(new_n15816_), .A2(new_n15809_), .A3(\asqrt[24] ), .ZN(new_n15824_));
  NOR2_X1    g15632(.A1(new_n15824_), .A2(new_n15823_), .ZN(new_n15825_));
  OAI21_X1   g15633(.A1(new_n15825_), .A2(new_n15818_), .B(\asqrt[25] ), .ZN(new_n15826_));
  INV_X1     g15634(.I(new_n15214_), .ZN(new_n15827_));
  NOR3_X1    g15635(.A1(new_n15770_), .A2(new_n15210_), .A3(new_n15565_), .ZN(new_n15828_));
  INV_X1     g15636(.I(new_n15828_), .ZN(new_n15829_));
  NOR3_X1    g15637(.A1(new_n15565_), .A2(new_n15210_), .A3(new_n15827_), .ZN(new_n15830_));
  AOI22_X1   g15638(.A1(new_n15829_), .A2(new_n15827_), .B1(\asqrt[14] ), .B2(new_n15830_), .ZN(new_n15831_));
  INV_X1     g15639(.I(new_n15831_), .ZN(new_n15832_));
  NAND2_X1   g15640(.A1(new_n15817_), .A2(new_n9846_), .ZN(new_n15833_));
  OAI21_X1   g15641(.A1(new_n15825_), .A2(new_n15833_), .B(new_n15832_), .ZN(new_n15834_));
  AOI21_X1   g15642(.A1(new_n15834_), .A2(new_n15826_), .B(new_n9317_), .ZN(new_n15835_));
  NOR3_X1    g15643(.A1(new_n15219_), .A2(new_n15545_), .A3(new_n15225_), .ZN(new_n15836_));
  NOR3_X1    g15644(.A1(new_n15770_), .A2(new_n15219_), .A3(new_n15225_), .ZN(new_n15837_));
  INV_X1     g15645(.I(new_n15837_), .ZN(new_n15838_));
  AOI22_X1   g15646(.A1(new_n15838_), .A2(new_n15545_), .B1(\asqrt[14] ), .B2(new_n15836_), .ZN(new_n15839_));
  OAI21_X1   g15647(.A1(new_n15823_), .A2(new_n15824_), .B(new_n15817_), .ZN(new_n15840_));
  AOI21_X1   g15648(.A1(new_n15840_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n15841_));
  AOI21_X1   g15649(.A1(new_n15841_), .A2(new_n15834_), .B(new_n15839_), .ZN(new_n15842_));
  OAI21_X1   g15650(.A1(new_n15842_), .A2(new_n15835_), .B(\asqrt[27] ), .ZN(new_n15843_));
  INV_X1     g15651(.I(new_n15843_), .ZN(new_n15844_));
  NOR2_X1    g15652(.A1(new_n15226_), .A2(new_n15234_), .ZN(new_n15845_));
  NOR3_X1    g15653(.A1(new_n15770_), .A2(new_n15559_), .A3(new_n15845_), .ZN(new_n15846_));
  INV_X1     g15654(.I(new_n15846_), .ZN(new_n15847_));
  NOR3_X1    g15655(.A1(new_n15845_), .A2(new_n15559_), .A3(new_n15233_), .ZN(new_n15848_));
  AOI22_X1   g15656(.A1(new_n15847_), .A2(new_n15233_), .B1(\asqrt[14] ), .B2(new_n15848_), .ZN(new_n15849_));
  NOR3_X1    g15657(.A1(new_n15842_), .A2(new_n15835_), .A3(\asqrt[27] ), .ZN(new_n15850_));
  NOR2_X1    g15658(.A1(new_n15850_), .A2(new_n15849_), .ZN(new_n15851_));
  OAI21_X1   g15659(.A1(new_n15851_), .A2(new_n15844_), .B(\asqrt[28] ), .ZN(new_n15852_));
  INV_X1     g15660(.I(new_n15242_), .ZN(new_n15853_));
  NOR3_X1    g15661(.A1(new_n15573_), .A2(new_n15236_), .A3(new_n15853_), .ZN(new_n15854_));
  NOR3_X1    g15662(.A1(new_n15770_), .A2(new_n15236_), .A3(new_n15573_), .ZN(new_n15855_));
  INV_X1     g15663(.I(new_n15855_), .ZN(new_n15856_));
  AOI22_X1   g15664(.A1(new_n15856_), .A2(new_n15853_), .B1(\asqrt[14] ), .B2(new_n15854_), .ZN(new_n15857_));
  INV_X1     g15665(.I(new_n15857_), .ZN(new_n15858_));
  NAND2_X1   g15666(.A1(new_n15843_), .A2(new_n8483_), .ZN(new_n15859_));
  OAI21_X1   g15667(.A1(new_n15851_), .A2(new_n15859_), .B(new_n15858_), .ZN(new_n15860_));
  AOI21_X1   g15668(.A1(new_n15860_), .A2(new_n15852_), .B(new_n8036_), .ZN(new_n15861_));
  NOR3_X1    g15669(.A1(new_n15770_), .A2(new_n15247_), .A3(new_n15256_), .ZN(new_n15862_));
  INV_X1     g15670(.I(new_n15862_), .ZN(new_n15863_));
  NOR3_X1    g15671(.A1(new_n15247_), .A2(new_n15544_), .A3(new_n15256_), .ZN(new_n15864_));
  AOI22_X1   g15672(.A1(new_n15863_), .A2(new_n15544_), .B1(\asqrt[14] ), .B2(new_n15864_), .ZN(new_n15865_));
  OAI21_X1   g15673(.A1(new_n15849_), .A2(new_n15850_), .B(new_n15843_), .ZN(new_n15866_));
  AOI21_X1   g15674(.A1(new_n15866_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n15867_));
  AOI21_X1   g15675(.A1(new_n15867_), .A2(new_n15860_), .B(new_n15865_), .ZN(new_n15868_));
  OAI21_X1   g15676(.A1(new_n15868_), .A2(new_n15861_), .B(\asqrt[30] ), .ZN(new_n15869_));
  INV_X1     g15677(.I(new_n15869_), .ZN(new_n15870_));
  NOR2_X1    g15678(.A1(new_n15257_), .A2(new_n15265_), .ZN(new_n15871_));
  NOR3_X1    g15679(.A1(new_n15871_), .A2(new_n15572_), .A3(new_n15264_), .ZN(new_n15872_));
  NOR3_X1    g15680(.A1(new_n15770_), .A2(new_n15572_), .A3(new_n15871_), .ZN(new_n15873_));
  INV_X1     g15681(.I(new_n15873_), .ZN(new_n15874_));
  AOI22_X1   g15682(.A1(new_n15874_), .A2(new_n15264_), .B1(\asqrt[14] ), .B2(new_n15872_), .ZN(new_n15875_));
  NOR3_X1    g15683(.A1(new_n15868_), .A2(new_n15861_), .A3(\asqrt[30] ), .ZN(new_n15876_));
  NOR2_X1    g15684(.A1(new_n15876_), .A2(new_n15875_), .ZN(new_n15877_));
  OAI21_X1   g15685(.A1(new_n15877_), .A2(new_n15870_), .B(\asqrt[31] ), .ZN(new_n15878_));
  INV_X1     g15686(.I(new_n15272_), .ZN(new_n15879_));
  NOR3_X1    g15687(.A1(new_n15770_), .A2(new_n15267_), .A3(new_n15581_), .ZN(new_n15880_));
  INV_X1     g15688(.I(new_n15880_), .ZN(new_n15881_));
  NOR3_X1    g15689(.A1(new_n15581_), .A2(new_n15267_), .A3(new_n15879_), .ZN(new_n15882_));
  AOI22_X1   g15690(.A1(new_n15881_), .A2(new_n15879_), .B1(\asqrt[14] ), .B2(new_n15882_), .ZN(new_n15883_));
  INV_X1     g15691(.I(new_n15883_), .ZN(new_n15884_));
  NAND2_X1   g15692(.A1(new_n15869_), .A2(new_n7229_), .ZN(new_n15885_));
  OAI21_X1   g15693(.A1(new_n15877_), .A2(new_n15885_), .B(new_n15884_), .ZN(new_n15886_));
  AOI21_X1   g15694(.A1(new_n15886_), .A2(new_n15878_), .B(new_n6824_), .ZN(new_n15887_));
  NOR3_X1    g15695(.A1(new_n15277_), .A2(new_n15543_), .A3(new_n15283_), .ZN(new_n15888_));
  NOR3_X1    g15696(.A1(new_n15770_), .A2(new_n15277_), .A3(new_n15283_), .ZN(new_n15889_));
  INV_X1     g15697(.I(new_n15889_), .ZN(new_n15890_));
  AOI22_X1   g15698(.A1(new_n15890_), .A2(new_n15543_), .B1(\asqrt[14] ), .B2(new_n15888_), .ZN(new_n15891_));
  OAI21_X1   g15699(.A1(new_n15875_), .A2(new_n15876_), .B(new_n15869_), .ZN(new_n15892_));
  AOI21_X1   g15700(.A1(new_n15892_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n15893_));
  AOI21_X1   g15701(.A1(new_n15893_), .A2(new_n15886_), .B(new_n15891_), .ZN(new_n15894_));
  OAI21_X1   g15702(.A1(new_n15894_), .A2(new_n15887_), .B(\asqrt[33] ), .ZN(new_n15895_));
  INV_X1     g15703(.I(new_n15895_), .ZN(new_n15896_));
  NOR2_X1    g15704(.A1(new_n15284_), .A2(new_n15292_), .ZN(new_n15897_));
  NOR3_X1    g15705(.A1(new_n15770_), .A2(new_n15580_), .A3(new_n15897_), .ZN(new_n15898_));
  INV_X1     g15706(.I(new_n15898_), .ZN(new_n15899_));
  NOR3_X1    g15707(.A1(new_n15897_), .A2(new_n15580_), .A3(new_n15291_), .ZN(new_n15900_));
  AOI22_X1   g15708(.A1(new_n15899_), .A2(new_n15291_), .B1(\asqrt[14] ), .B2(new_n15900_), .ZN(new_n15901_));
  NOR3_X1    g15709(.A1(new_n15894_), .A2(new_n15887_), .A3(\asqrt[33] ), .ZN(new_n15902_));
  NOR2_X1    g15710(.A1(new_n15902_), .A2(new_n15901_), .ZN(new_n15903_));
  OAI21_X1   g15711(.A1(new_n15903_), .A2(new_n15896_), .B(\asqrt[34] ), .ZN(new_n15904_));
  INV_X1     g15712(.I(new_n15299_), .ZN(new_n15905_));
  NOR3_X1    g15713(.A1(new_n15589_), .A2(new_n15294_), .A3(new_n15905_), .ZN(new_n15906_));
  NOR3_X1    g15714(.A1(new_n15770_), .A2(new_n15294_), .A3(new_n15589_), .ZN(new_n15907_));
  INV_X1     g15715(.I(new_n15907_), .ZN(new_n15908_));
  AOI22_X1   g15716(.A1(new_n15908_), .A2(new_n15905_), .B1(\asqrt[14] ), .B2(new_n15906_), .ZN(new_n15909_));
  INV_X1     g15717(.I(new_n15909_), .ZN(new_n15910_));
  NAND2_X1   g15718(.A1(new_n15895_), .A2(new_n6077_), .ZN(new_n15911_));
  OAI21_X1   g15719(.A1(new_n15903_), .A2(new_n15911_), .B(new_n15910_), .ZN(new_n15912_));
  AOI21_X1   g15720(.A1(new_n15912_), .A2(new_n15904_), .B(new_n5708_), .ZN(new_n15913_));
  NOR3_X1    g15721(.A1(new_n15770_), .A2(new_n15304_), .A3(new_n15310_), .ZN(new_n15914_));
  INV_X1     g15722(.I(new_n15914_), .ZN(new_n15915_));
  NOR3_X1    g15723(.A1(new_n15304_), .A2(new_n15542_), .A3(new_n15310_), .ZN(new_n15916_));
  AOI22_X1   g15724(.A1(new_n15915_), .A2(new_n15542_), .B1(\asqrt[14] ), .B2(new_n15916_), .ZN(new_n15917_));
  OAI21_X1   g15725(.A1(new_n15901_), .A2(new_n15902_), .B(new_n15895_), .ZN(new_n15918_));
  AOI21_X1   g15726(.A1(new_n15918_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n15919_));
  AOI21_X1   g15727(.A1(new_n15919_), .A2(new_n15912_), .B(new_n15917_), .ZN(new_n15920_));
  OAI21_X1   g15728(.A1(new_n15920_), .A2(new_n15913_), .B(\asqrt[36] ), .ZN(new_n15921_));
  INV_X1     g15729(.I(new_n15921_), .ZN(new_n15922_));
  NOR2_X1    g15730(.A1(new_n15311_), .A2(new_n15319_), .ZN(new_n15923_));
  NOR3_X1    g15731(.A1(new_n15923_), .A2(new_n15588_), .A3(new_n15318_), .ZN(new_n15924_));
  NOR3_X1    g15732(.A1(new_n15770_), .A2(new_n15588_), .A3(new_n15923_), .ZN(new_n15925_));
  INV_X1     g15733(.I(new_n15925_), .ZN(new_n15926_));
  AOI22_X1   g15734(.A1(new_n15926_), .A2(new_n15318_), .B1(\asqrt[14] ), .B2(new_n15924_), .ZN(new_n15927_));
  NOR3_X1    g15735(.A1(new_n15920_), .A2(new_n15913_), .A3(\asqrt[36] ), .ZN(new_n15928_));
  NOR2_X1    g15736(.A1(new_n15928_), .A2(new_n15927_), .ZN(new_n15929_));
  OAI21_X1   g15737(.A1(new_n15929_), .A2(new_n15922_), .B(\asqrt[37] ), .ZN(new_n15930_));
  INV_X1     g15738(.I(new_n15326_), .ZN(new_n15931_));
  NOR3_X1    g15739(.A1(new_n15770_), .A2(new_n15321_), .A3(new_n15597_), .ZN(new_n15932_));
  INV_X1     g15740(.I(new_n15932_), .ZN(new_n15933_));
  NOR3_X1    g15741(.A1(new_n15597_), .A2(new_n15321_), .A3(new_n15931_), .ZN(new_n15934_));
  AOI22_X1   g15742(.A1(new_n15933_), .A2(new_n15931_), .B1(\asqrt[14] ), .B2(new_n15934_), .ZN(new_n15935_));
  INV_X1     g15743(.I(new_n15935_), .ZN(new_n15936_));
  NAND2_X1   g15744(.A1(new_n15921_), .A2(new_n5024_), .ZN(new_n15937_));
  OAI21_X1   g15745(.A1(new_n15929_), .A2(new_n15937_), .B(new_n15936_), .ZN(new_n15938_));
  AOI21_X1   g15746(.A1(new_n15938_), .A2(new_n15930_), .B(new_n4696_), .ZN(new_n15939_));
  NOR3_X1    g15747(.A1(new_n15331_), .A2(new_n15541_), .A3(new_n15337_), .ZN(new_n15940_));
  NOR3_X1    g15748(.A1(new_n15770_), .A2(new_n15331_), .A3(new_n15337_), .ZN(new_n15941_));
  INV_X1     g15749(.I(new_n15941_), .ZN(new_n15942_));
  AOI22_X1   g15750(.A1(new_n15942_), .A2(new_n15541_), .B1(\asqrt[14] ), .B2(new_n15940_), .ZN(new_n15943_));
  OAI21_X1   g15751(.A1(new_n15927_), .A2(new_n15928_), .B(new_n15921_), .ZN(new_n15944_));
  AOI21_X1   g15752(.A1(new_n15944_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n15945_));
  AOI21_X1   g15753(.A1(new_n15945_), .A2(new_n15938_), .B(new_n15943_), .ZN(new_n15946_));
  OAI21_X1   g15754(.A1(new_n15946_), .A2(new_n15939_), .B(\asqrt[39] ), .ZN(new_n15947_));
  INV_X1     g15755(.I(new_n15947_), .ZN(new_n15948_));
  NOR2_X1    g15756(.A1(new_n15338_), .A2(new_n15346_), .ZN(new_n15949_));
  NOR3_X1    g15757(.A1(new_n15770_), .A2(new_n15596_), .A3(new_n15949_), .ZN(new_n15950_));
  INV_X1     g15758(.I(new_n15950_), .ZN(new_n15951_));
  NOR3_X1    g15759(.A1(new_n15949_), .A2(new_n15596_), .A3(new_n15345_), .ZN(new_n15952_));
  AOI22_X1   g15760(.A1(new_n15951_), .A2(new_n15345_), .B1(\asqrt[14] ), .B2(new_n15952_), .ZN(new_n15953_));
  NOR3_X1    g15761(.A1(new_n15946_), .A2(new_n15939_), .A3(\asqrt[39] ), .ZN(new_n15954_));
  NOR2_X1    g15762(.A1(new_n15954_), .A2(new_n15953_), .ZN(new_n15955_));
  OAI21_X1   g15763(.A1(new_n15955_), .A2(new_n15948_), .B(\asqrt[40] ), .ZN(new_n15956_));
  INV_X1     g15764(.I(new_n15352_), .ZN(new_n15957_));
  NOR3_X1    g15765(.A1(new_n15605_), .A2(new_n15348_), .A3(new_n15957_), .ZN(new_n15958_));
  NOR3_X1    g15766(.A1(new_n15770_), .A2(new_n15348_), .A3(new_n15605_), .ZN(new_n15959_));
  INV_X1     g15767(.I(new_n15959_), .ZN(new_n15960_));
  AOI22_X1   g15768(.A1(new_n15960_), .A2(new_n15957_), .B1(\asqrt[14] ), .B2(new_n15958_), .ZN(new_n15961_));
  INV_X1     g15769(.I(new_n15961_), .ZN(new_n15962_));
  NAND2_X1   g15770(.A1(new_n15947_), .A2(new_n4071_), .ZN(new_n15963_));
  OAI21_X1   g15771(.A1(new_n15955_), .A2(new_n15963_), .B(new_n15962_), .ZN(new_n15964_));
  AOI21_X1   g15772(.A1(new_n15964_), .A2(new_n15956_), .B(new_n3782_), .ZN(new_n15965_));
  NOR3_X1    g15773(.A1(new_n15770_), .A2(new_n15357_), .A3(new_n15363_), .ZN(new_n15966_));
  INV_X1     g15774(.I(new_n15966_), .ZN(new_n15967_));
  NOR3_X1    g15775(.A1(new_n15357_), .A2(new_n15540_), .A3(new_n15363_), .ZN(new_n15968_));
  AOI22_X1   g15776(.A1(new_n15967_), .A2(new_n15540_), .B1(\asqrt[14] ), .B2(new_n15968_), .ZN(new_n15969_));
  OAI21_X1   g15777(.A1(new_n15953_), .A2(new_n15954_), .B(new_n15947_), .ZN(new_n15970_));
  AOI21_X1   g15778(.A1(new_n15970_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n15971_));
  AOI21_X1   g15779(.A1(new_n15971_), .A2(new_n15964_), .B(new_n15969_), .ZN(new_n15972_));
  OAI21_X1   g15780(.A1(new_n15972_), .A2(new_n15965_), .B(\asqrt[42] ), .ZN(new_n15973_));
  INV_X1     g15781(.I(new_n15973_), .ZN(new_n15974_));
  NOR2_X1    g15782(.A1(new_n15364_), .A2(new_n15372_), .ZN(new_n15975_));
  NOR3_X1    g15783(.A1(new_n15975_), .A2(new_n15604_), .A3(new_n15371_), .ZN(new_n15976_));
  NOR3_X1    g15784(.A1(new_n15770_), .A2(new_n15604_), .A3(new_n15975_), .ZN(new_n15977_));
  INV_X1     g15785(.I(new_n15977_), .ZN(new_n15978_));
  AOI22_X1   g15786(.A1(new_n15978_), .A2(new_n15371_), .B1(\asqrt[14] ), .B2(new_n15976_), .ZN(new_n15979_));
  NOR3_X1    g15787(.A1(new_n15972_), .A2(new_n15965_), .A3(\asqrt[42] ), .ZN(new_n15980_));
  NOR2_X1    g15788(.A1(new_n15980_), .A2(new_n15979_), .ZN(new_n15981_));
  OAI21_X1   g15789(.A1(new_n15981_), .A2(new_n15974_), .B(\asqrt[43] ), .ZN(new_n15982_));
  INV_X1     g15790(.I(new_n15378_), .ZN(new_n15983_));
  NOR3_X1    g15791(.A1(new_n15770_), .A2(new_n15374_), .A3(new_n15613_), .ZN(new_n15984_));
  INV_X1     g15792(.I(new_n15984_), .ZN(new_n15985_));
  NOR3_X1    g15793(.A1(new_n15613_), .A2(new_n15374_), .A3(new_n15983_), .ZN(new_n15986_));
  AOI22_X1   g15794(.A1(new_n15985_), .A2(new_n15983_), .B1(\asqrt[14] ), .B2(new_n15986_), .ZN(new_n15987_));
  INV_X1     g15795(.I(new_n15987_), .ZN(new_n15988_));
  NAND2_X1   g15796(.A1(new_n15973_), .A2(new_n3218_), .ZN(new_n15989_));
  OAI21_X1   g15797(.A1(new_n15981_), .A2(new_n15989_), .B(new_n15988_), .ZN(new_n15990_));
  AOI21_X1   g15798(.A1(new_n15990_), .A2(new_n15982_), .B(new_n2954_), .ZN(new_n15991_));
  NOR3_X1    g15799(.A1(new_n15383_), .A2(new_n15539_), .A3(new_n15391_), .ZN(new_n15992_));
  NOR3_X1    g15800(.A1(new_n15770_), .A2(new_n15383_), .A3(new_n15391_), .ZN(new_n15993_));
  INV_X1     g15801(.I(new_n15993_), .ZN(new_n15994_));
  AOI22_X1   g15802(.A1(new_n15994_), .A2(new_n15539_), .B1(\asqrt[14] ), .B2(new_n15992_), .ZN(new_n15995_));
  OAI21_X1   g15803(.A1(new_n15979_), .A2(new_n15980_), .B(new_n15973_), .ZN(new_n15996_));
  AOI21_X1   g15804(.A1(new_n15996_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n15997_));
  AOI21_X1   g15805(.A1(new_n15997_), .A2(new_n15990_), .B(new_n15995_), .ZN(new_n15998_));
  OAI21_X1   g15806(.A1(new_n15998_), .A2(new_n15991_), .B(\asqrt[45] ), .ZN(new_n15999_));
  INV_X1     g15807(.I(new_n15999_), .ZN(new_n16000_));
  NOR2_X1    g15808(.A1(new_n15392_), .A2(new_n15399_), .ZN(new_n16001_));
  NOR3_X1    g15809(.A1(new_n15770_), .A2(new_n15612_), .A3(new_n16001_), .ZN(new_n16002_));
  INV_X1     g15810(.I(new_n16002_), .ZN(new_n16003_));
  NOR3_X1    g15811(.A1(new_n16001_), .A2(new_n15612_), .A3(new_n15398_), .ZN(new_n16004_));
  AOI22_X1   g15812(.A1(new_n16003_), .A2(new_n15398_), .B1(\asqrt[14] ), .B2(new_n16004_), .ZN(new_n16005_));
  NOR3_X1    g15813(.A1(new_n15998_), .A2(new_n15991_), .A3(\asqrt[45] ), .ZN(new_n16006_));
  NOR2_X1    g15814(.A1(new_n16006_), .A2(new_n16005_), .ZN(new_n16007_));
  OAI21_X1   g15815(.A1(new_n16007_), .A2(new_n16000_), .B(\asqrt[46] ), .ZN(new_n16008_));
  INV_X1     g15816(.I(new_n15407_), .ZN(new_n16009_));
  NOR3_X1    g15817(.A1(new_n15621_), .A2(new_n15401_), .A3(new_n16009_), .ZN(new_n16010_));
  NOR3_X1    g15818(.A1(new_n15770_), .A2(new_n15401_), .A3(new_n15621_), .ZN(new_n16011_));
  INV_X1     g15819(.I(new_n16011_), .ZN(new_n16012_));
  AOI22_X1   g15820(.A1(new_n16012_), .A2(new_n16009_), .B1(\asqrt[14] ), .B2(new_n16010_), .ZN(new_n16013_));
  INV_X1     g15821(.I(new_n16013_), .ZN(new_n16014_));
  NAND2_X1   g15822(.A1(new_n15999_), .A2(new_n2465_), .ZN(new_n16015_));
  OAI21_X1   g15823(.A1(new_n16007_), .A2(new_n16015_), .B(new_n16014_), .ZN(new_n16016_));
  AOI21_X1   g15824(.A1(new_n16016_), .A2(new_n16008_), .B(new_n2229_), .ZN(new_n16017_));
  NOR3_X1    g15825(.A1(new_n15770_), .A2(new_n15412_), .A3(new_n15421_), .ZN(new_n16018_));
  INV_X1     g15826(.I(new_n16018_), .ZN(new_n16019_));
  NOR3_X1    g15827(.A1(new_n15412_), .A2(new_n15538_), .A3(new_n15421_), .ZN(new_n16020_));
  AOI22_X1   g15828(.A1(new_n16019_), .A2(new_n15538_), .B1(\asqrt[14] ), .B2(new_n16020_), .ZN(new_n16021_));
  OAI21_X1   g15829(.A1(new_n16005_), .A2(new_n16006_), .B(new_n15999_), .ZN(new_n16022_));
  AOI21_X1   g15830(.A1(new_n16022_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n16023_));
  AOI21_X1   g15831(.A1(new_n16023_), .A2(new_n16016_), .B(new_n16021_), .ZN(new_n16024_));
  OAI21_X1   g15832(.A1(new_n16024_), .A2(new_n16017_), .B(\asqrt[48] ), .ZN(new_n16025_));
  INV_X1     g15833(.I(new_n16025_), .ZN(new_n16026_));
  NOR2_X1    g15834(.A1(new_n15422_), .A2(new_n15429_), .ZN(new_n16027_));
  NOR3_X1    g15835(.A1(new_n16027_), .A2(new_n15620_), .A3(new_n15428_), .ZN(new_n16028_));
  NOR3_X1    g15836(.A1(new_n15770_), .A2(new_n15620_), .A3(new_n16027_), .ZN(new_n16029_));
  INV_X1     g15837(.I(new_n16029_), .ZN(new_n16030_));
  AOI22_X1   g15838(.A1(new_n16030_), .A2(new_n15428_), .B1(\asqrt[14] ), .B2(new_n16028_), .ZN(new_n16031_));
  NOR3_X1    g15839(.A1(new_n16024_), .A2(new_n16017_), .A3(\asqrt[48] ), .ZN(new_n16032_));
  NOR2_X1    g15840(.A1(new_n16032_), .A2(new_n16031_), .ZN(new_n16033_));
  OAI21_X1   g15841(.A1(new_n16033_), .A2(new_n16026_), .B(\asqrt[49] ), .ZN(new_n16034_));
  INV_X1     g15842(.I(new_n15437_), .ZN(new_n16035_));
  NOR3_X1    g15843(.A1(new_n15770_), .A2(new_n15431_), .A3(new_n15629_), .ZN(new_n16036_));
  INV_X1     g15844(.I(new_n16036_), .ZN(new_n16037_));
  NOR3_X1    g15845(.A1(new_n15629_), .A2(new_n15431_), .A3(new_n16035_), .ZN(new_n16038_));
  AOI22_X1   g15846(.A1(new_n16037_), .A2(new_n16035_), .B1(\asqrt[14] ), .B2(new_n16038_), .ZN(new_n16039_));
  INV_X1     g15847(.I(new_n16039_), .ZN(new_n16040_));
  NAND2_X1   g15848(.A1(new_n16025_), .A2(new_n1806_), .ZN(new_n16041_));
  OAI21_X1   g15849(.A1(new_n16033_), .A2(new_n16041_), .B(new_n16040_), .ZN(new_n16042_));
  AOI21_X1   g15850(.A1(new_n16042_), .A2(new_n16034_), .B(new_n1612_), .ZN(new_n16043_));
  NOR3_X1    g15851(.A1(new_n15442_), .A2(new_n15537_), .A3(new_n15451_), .ZN(new_n16044_));
  NOR3_X1    g15852(.A1(new_n15770_), .A2(new_n15442_), .A3(new_n15451_), .ZN(new_n16045_));
  INV_X1     g15853(.I(new_n16045_), .ZN(new_n16046_));
  AOI22_X1   g15854(.A1(new_n16046_), .A2(new_n15537_), .B1(\asqrt[14] ), .B2(new_n16044_), .ZN(new_n16047_));
  OAI21_X1   g15855(.A1(new_n16031_), .A2(new_n16032_), .B(new_n16025_), .ZN(new_n16048_));
  AOI21_X1   g15856(.A1(new_n16048_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n16049_));
  AOI21_X1   g15857(.A1(new_n16049_), .A2(new_n16042_), .B(new_n16047_), .ZN(new_n16050_));
  OAI21_X1   g15858(.A1(new_n16050_), .A2(new_n16043_), .B(\asqrt[51] ), .ZN(new_n16051_));
  INV_X1     g15859(.I(new_n16051_), .ZN(new_n16052_));
  NOR2_X1    g15860(.A1(new_n15452_), .A2(new_n15459_), .ZN(new_n16053_));
  NOR3_X1    g15861(.A1(new_n15770_), .A2(new_n15628_), .A3(new_n16053_), .ZN(new_n16054_));
  INV_X1     g15862(.I(new_n16054_), .ZN(new_n16055_));
  NOR3_X1    g15863(.A1(new_n16053_), .A2(new_n15628_), .A3(new_n15458_), .ZN(new_n16056_));
  AOI22_X1   g15864(.A1(new_n16055_), .A2(new_n15458_), .B1(\asqrt[14] ), .B2(new_n16056_), .ZN(new_n16057_));
  NOR3_X1    g15865(.A1(new_n16050_), .A2(new_n16043_), .A3(\asqrt[51] ), .ZN(new_n16058_));
  NOR2_X1    g15866(.A1(new_n16058_), .A2(new_n16057_), .ZN(new_n16059_));
  OAI21_X1   g15867(.A1(new_n16059_), .A2(new_n16052_), .B(\asqrt[52] ), .ZN(new_n16060_));
  INV_X1     g15868(.I(new_n15467_), .ZN(new_n16061_));
  NAND2_X1   g15869(.A1(new_n15469_), .A2(new_n15460_), .ZN(new_n16062_));
  INV_X1     g15870(.I(new_n16062_), .ZN(new_n16063_));
  NOR3_X1    g15871(.A1(new_n16063_), .A2(new_n15461_), .A3(new_n16061_), .ZN(new_n16064_));
  NOR3_X1    g15872(.A1(new_n15770_), .A2(new_n15461_), .A3(new_n16063_), .ZN(new_n16065_));
  INV_X1     g15873(.I(new_n16065_), .ZN(new_n16066_));
  AOI22_X1   g15874(.A1(new_n16066_), .A2(new_n16061_), .B1(\asqrt[14] ), .B2(new_n16064_), .ZN(new_n16067_));
  INV_X1     g15875(.I(new_n16067_), .ZN(new_n16068_));
  NAND2_X1   g15876(.A1(new_n16051_), .A2(new_n1256_), .ZN(new_n16069_));
  OAI21_X1   g15877(.A1(new_n16059_), .A2(new_n16069_), .B(new_n16068_), .ZN(new_n16070_));
  AOI21_X1   g15878(.A1(new_n16070_), .A2(new_n16060_), .B(new_n1103_), .ZN(new_n16071_));
  NOR3_X1    g15879(.A1(new_n15770_), .A2(new_n15472_), .A3(new_n15481_), .ZN(new_n16072_));
  INV_X1     g15880(.I(new_n16072_), .ZN(new_n16073_));
  NOR3_X1    g15881(.A1(new_n15472_), .A2(new_n15536_), .A3(new_n15481_), .ZN(new_n16074_));
  AOI22_X1   g15882(.A1(new_n16073_), .A2(new_n15536_), .B1(\asqrt[14] ), .B2(new_n16074_), .ZN(new_n16075_));
  OAI21_X1   g15883(.A1(new_n16057_), .A2(new_n16058_), .B(new_n16051_), .ZN(new_n16076_));
  AOI21_X1   g15884(.A1(new_n16076_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n16077_));
  AOI21_X1   g15885(.A1(new_n16077_), .A2(new_n16070_), .B(new_n16075_), .ZN(new_n16078_));
  OAI21_X1   g15886(.A1(new_n16078_), .A2(new_n16071_), .B(\asqrt[54] ), .ZN(new_n16079_));
  INV_X1     g15887(.I(new_n16079_), .ZN(new_n16080_));
  INV_X1     g15888(.I(new_n15483_), .ZN(new_n16081_));
  INV_X1     g15889(.I(new_n15636_), .ZN(new_n16082_));
  NOR3_X1    g15890(.A1(new_n16081_), .A2(new_n16082_), .A3(new_n15488_), .ZN(new_n16083_));
  NOR3_X1    g15891(.A1(new_n15770_), .A2(new_n16081_), .A3(new_n16082_), .ZN(new_n16084_));
  INV_X1     g15892(.I(new_n16084_), .ZN(new_n16085_));
  AOI22_X1   g15893(.A1(new_n16085_), .A2(new_n15488_), .B1(\asqrt[14] ), .B2(new_n16083_), .ZN(new_n16086_));
  NOR3_X1    g15894(.A1(new_n16078_), .A2(new_n16071_), .A3(\asqrt[54] ), .ZN(new_n16087_));
  NOR2_X1    g15895(.A1(new_n16087_), .A2(new_n16086_), .ZN(new_n16088_));
  OAI21_X1   g15896(.A1(new_n16088_), .A2(new_n16080_), .B(\asqrt[55] ), .ZN(new_n16089_));
  INV_X1     g15897(.I(new_n15497_), .ZN(new_n16090_));
  INV_X1     g15898(.I(new_n15490_), .ZN(new_n16091_));
  INV_X1     g15899(.I(new_n15499_), .ZN(new_n16092_));
  NOR2_X1    g15900(.A1(new_n16092_), .A2(new_n16091_), .ZN(new_n16093_));
  NOR3_X1    g15901(.A1(new_n15770_), .A2(new_n15491_), .A3(new_n16093_), .ZN(new_n16094_));
  INV_X1     g15902(.I(new_n16094_), .ZN(new_n16095_));
  NOR3_X1    g15903(.A1(new_n16093_), .A2(new_n15491_), .A3(new_n16090_), .ZN(new_n16096_));
  AOI22_X1   g15904(.A1(new_n16095_), .A2(new_n16090_), .B1(\asqrt[14] ), .B2(new_n16096_), .ZN(new_n16097_));
  INV_X1     g15905(.I(new_n16097_), .ZN(new_n16098_));
  NAND2_X1   g15906(.A1(new_n16079_), .A2(new_n823_), .ZN(new_n16099_));
  OAI21_X1   g15907(.A1(new_n16088_), .A2(new_n16099_), .B(new_n16098_), .ZN(new_n16100_));
  AOI21_X1   g15908(.A1(new_n16100_), .A2(new_n16089_), .B(new_n703_), .ZN(new_n16101_));
  NOR3_X1    g15909(.A1(new_n15502_), .A2(new_n15535_), .A3(new_n15508_), .ZN(new_n16102_));
  NOR3_X1    g15910(.A1(new_n15770_), .A2(new_n15502_), .A3(new_n15508_), .ZN(new_n16103_));
  INV_X1     g15911(.I(new_n16103_), .ZN(new_n16104_));
  AOI22_X1   g15912(.A1(new_n16104_), .A2(new_n15535_), .B1(\asqrt[14] ), .B2(new_n16102_), .ZN(new_n16105_));
  OAI21_X1   g15913(.A1(new_n16086_), .A2(new_n16087_), .B(new_n16079_), .ZN(new_n16106_));
  AOI21_X1   g15914(.A1(new_n16106_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n16107_));
  AOI21_X1   g15915(.A1(new_n16107_), .A2(new_n16100_), .B(new_n16105_), .ZN(new_n16108_));
  OAI21_X1   g15916(.A1(new_n16108_), .A2(new_n16101_), .B(\asqrt[57] ), .ZN(new_n16109_));
  INV_X1     g15917(.I(new_n16109_), .ZN(new_n16110_));
  INV_X1     g15918(.I(new_n15510_), .ZN(new_n16111_));
  INV_X1     g15919(.I(new_n15640_), .ZN(new_n16112_));
  NOR3_X1    g15920(.A1(new_n15770_), .A2(new_n16111_), .A3(new_n16112_), .ZN(new_n16113_));
  INV_X1     g15921(.I(new_n16113_), .ZN(new_n16114_));
  NOR3_X1    g15922(.A1(new_n16111_), .A2(new_n16112_), .A3(new_n15515_), .ZN(new_n16115_));
  AOI22_X1   g15923(.A1(new_n16114_), .A2(new_n15515_), .B1(\asqrt[14] ), .B2(new_n16115_), .ZN(new_n16116_));
  NOR3_X1    g15924(.A1(new_n16108_), .A2(new_n16101_), .A3(\asqrt[57] ), .ZN(new_n16117_));
  NOR2_X1    g15925(.A1(new_n16117_), .A2(new_n16116_), .ZN(new_n16118_));
  OAI21_X1   g15926(.A1(new_n16118_), .A2(new_n16110_), .B(\asqrt[58] ), .ZN(new_n16119_));
  INV_X1     g15927(.I(new_n15524_), .ZN(new_n16120_));
  INV_X1     g15928(.I(new_n15517_), .ZN(new_n16121_));
  INV_X1     g15929(.I(new_n15526_), .ZN(new_n16122_));
  OAI21_X1   g15930(.A1(new_n16122_), .A2(new_n16121_), .B(new_n15524_), .ZN(new_n16123_));
  NOR2_X1    g15931(.A1(new_n16123_), .A2(new_n15518_), .ZN(new_n16124_));
  NOR2_X1    g15932(.A1(new_n16122_), .A2(new_n16121_), .ZN(new_n16125_));
  NOR3_X1    g15933(.A1(new_n15770_), .A2(new_n15518_), .A3(new_n16125_), .ZN(new_n16126_));
  INV_X1     g15934(.I(new_n16126_), .ZN(new_n16127_));
  AOI22_X1   g15935(.A1(new_n16127_), .A2(new_n16120_), .B1(\asqrt[14] ), .B2(new_n16124_), .ZN(new_n16128_));
  INV_X1     g15936(.I(new_n16128_), .ZN(new_n16129_));
  NAND2_X1   g15937(.A1(new_n16109_), .A2(new_n436_), .ZN(new_n16130_));
  OAI21_X1   g15938(.A1(new_n16118_), .A2(new_n16130_), .B(new_n16129_), .ZN(new_n16131_));
  AOI21_X1   g15939(.A1(new_n16131_), .A2(new_n16119_), .B(new_n327_), .ZN(new_n16132_));
  NOR3_X1    g15940(.A1(new_n15770_), .A2(new_n15660_), .A3(new_n15661_), .ZN(new_n16133_));
  INV_X1     g15941(.I(new_n16133_), .ZN(new_n16134_));
  NOR3_X1    g15942(.A1(new_n15660_), .A2(new_n15534_), .A3(new_n15661_), .ZN(new_n16135_));
  AOI22_X1   g15943(.A1(new_n16134_), .A2(new_n15534_), .B1(\asqrt[14] ), .B2(new_n16135_), .ZN(new_n16136_));
  OAI21_X1   g15944(.A1(new_n16116_), .A2(new_n16117_), .B(new_n16109_), .ZN(new_n16137_));
  AOI21_X1   g15945(.A1(new_n16137_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n16138_));
  AOI21_X1   g15946(.A1(new_n16138_), .A2(new_n16131_), .B(new_n16136_), .ZN(new_n16139_));
  OAI21_X1   g15947(.A1(new_n16139_), .A2(new_n16132_), .B(\asqrt[60] ), .ZN(new_n16140_));
  INV_X1     g15948(.I(new_n16140_), .ZN(new_n16141_));
  INV_X1     g15949(.I(new_n15719_), .ZN(new_n16142_));
  NOR3_X1    g15950(.A1(new_n16142_), .A2(new_n15644_), .A3(new_n15672_), .ZN(new_n16143_));
  NOR3_X1    g15951(.A1(new_n15770_), .A2(new_n15644_), .A3(new_n16142_), .ZN(new_n16144_));
  INV_X1     g15952(.I(new_n16144_), .ZN(new_n16145_));
  AOI22_X1   g15953(.A1(new_n16145_), .A2(new_n15672_), .B1(\asqrt[14] ), .B2(new_n16143_), .ZN(new_n16146_));
  NOR3_X1    g15954(.A1(new_n16139_), .A2(new_n16132_), .A3(\asqrt[60] ), .ZN(new_n16147_));
  NOR2_X1    g15955(.A1(new_n16147_), .A2(new_n16146_), .ZN(new_n16148_));
  OAI21_X1   g15956(.A1(new_n16148_), .A2(new_n16141_), .B(\asqrt[61] ), .ZN(new_n16149_));
  NAND2_X1   g15957(.A1(new_n15684_), .A2(new_n15673_), .ZN(new_n16150_));
  NAND3_X1   g15958(.A1(\asqrt[14] ), .A2(new_n15652_), .A3(new_n16150_), .ZN(new_n16151_));
  AND3_X2    g15959(.A1(new_n15652_), .A2(new_n15658_), .A3(new_n16150_), .Z(new_n16152_));
  AOI22_X1   g15960(.A1(new_n16151_), .A2(new_n15659_), .B1(\asqrt[14] ), .B2(new_n16152_), .ZN(new_n16153_));
  INV_X1     g15961(.I(new_n16153_), .ZN(new_n16154_));
  NAND2_X1   g15962(.A1(new_n16140_), .A2(new_n218_), .ZN(new_n16155_));
  OAI21_X1   g15963(.A1(new_n16148_), .A2(new_n16155_), .B(new_n16154_), .ZN(new_n16156_));
  AOI21_X1   g15964(.A1(new_n16156_), .A2(new_n16149_), .B(new_n207_), .ZN(new_n16157_));
  NOR3_X1    g15965(.A1(new_n15666_), .A2(new_n15718_), .A3(new_n15697_), .ZN(new_n16158_));
  NOR3_X1    g15966(.A1(new_n15770_), .A2(new_n15666_), .A3(new_n15697_), .ZN(new_n16159_));
  INV_X1     g15967(.I(new_n16159_), .ZN(new_n16160_));
  AOI22_X1   g15968(.A1(new_n16160_), .A2(new_n15718_), .B1(\asqrt[14] ), .B2(new_n16158_), .ZN(new_n16161_));
  OAI21_X1   g15969(.A1(new_n16146_), .A2(new_n16147_), .B(new_n16140_), .ZN(new_n16162_));
  AOI21_X1   g15970(.A1(new_n16162_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n16163_));
  AOI21_X1   g15971(.A1(new_n16163_), .A2(new_n16156_), .B(new_n16161_), .ZN(new_n16164_));
  INV_X1     g15972(.I(new_n15677_), .ZN(new_n16165_));
  INV_X1     g15973(.I(new_n15731_), .ZN(new_n16166_));
  NOR3_X1    g15974(.A1(new_n16165_), .A2(new_n16166_), .A3(new_n15682_), .ZN(new_n16167_));
  NAND2_X1   g15975(.A1(\asqrt[14] ), .A2(new_n16167_), .ZN(new_n16168_));
  INV_X1     g15976(.I(new_n16168_), .ZN(new_n16169_));
  NOR2_X1    g15977(.A1(new_n16165_), .A2(new_n16166_), .ZN(new_n16170_));
  AOI21_X1   g15978(.A1(\asqrt[14] ), .A2(new_n16170_), .B(new_n15681_), .ZN(new_n16171_));
  NOR2_X1    g15979(.A1(new_n16169_), .A2(new_n16171_), .ZN(new_n16172_));
  INV_X1     g15980(.I(new_n16172_), .ZN(new_n16173_));
  NAND3_X1   g15981(.A1(\asqrt[14] ), .A2(new_n15715_), .A3(new_n15692_), .ZN(new_n16174_));
  AND3_X2    g15982(.A1(new_n16173_), .A2(new_n15745_), .A3(new_n16174_), .Z(new_n16175_));
  OAI21_X1   g15983(.A1(new_n16164_), .A2(new_n16157_), .B(new_n16175_), .ZN(new_n16176_));
  NAND2_X1   g15984(.A1(new_n16176_), .A2(new_n193_), .ZN(new_n16177_));
  INV_X1     g15985(.I(new_n16146_), .ZN(new_n16178_));
  INV_X1     g15986(.I(new_n16116_), .ZN(new_n16179_));
  INV_X1     g15987(.I(new_n16086_), .ZN(new_n16180_));
  INV_X1     g15988(.I(new_n16057_), .ZN(new_n16181_));
  INV_X1     g15989(.I(new_n16031_), .ZN(new_n16182_));
  INV_X1     g15990(.I(new_n16005_), .ZN(new_n16183_));
  INV_X1     g15991(.I(new_n15979_), .ZN(new_n16184_));
  INV_X1     g15992(.I(new_n15953_), .ZN(new_n16185_));
  INV_X1     g15993(.I(new_n15927_), .ZN(new_n16186_));
  INV_X1     g15994(.I(new_n15901_), .ZN(new_n16187_));
  INV_X1     g15995(.I(new_n15875_), .ZN(new_n16188_));
  INV_X1     g15996(.I(new_n15849_), .ZN(new_n16189_));
  INV_X1     g15997(.I(new_n15823_), .ZN(new_n16190_));
  INV_X1     g15998(.I(new_n15797_), .ZN(new_n16191_));
  NAND2_X1   g15999(.A1(new_n15728_), .A2(new_n15736_), .ZN(new_n16192_));
  OAI21_X1   g16000(.A1(new_n15717_), .A2(new_n15727_), .B(new_n15730_), .ZN(new_n16193_));
  NAND2_X1   g16001(.A1(new_n16193_), .A2(\a[29] ), .ZN(new_n16194_));
  NAND3_X1   g16002(.A1(new_n16192_), .A2(new_n16194_), .A3(new_n15744_), .ZN(new_n16195_));
  AOI21_X1   g16003(.A1(new_n16195_), .A2(new_n15759_), .B(new_n14601_), .ZN(new_n16196_));
  OAI21_X1   g16004(.A1(new_n15750_), .A2(new_n15739_), .B(\a[30] ), .ZN(new_n16197_));
  NAND3_X1   g16005(.A1(new_n15747_), .A2(new_n15744_), .A3(new_n15068_), .ZN(new_n16198_));
  NAND2_X1   g16006(.A1(new_n15728_), .A2(new_n15714_), .ZN(new_n16199_));
  AOI21_X1   g16007(.A1(new_n16199_), .A2(\asqrt[15] ), .B(\asqrt[16] ), .ZN(new_n16200_));
  AOI22_X1   g16008(.A1(new_n16195_), .A2(new_n16200_), .B1(new_n16197_), .B2(new_n16198_), .ZN(new_n16201_));
  OAI21_X1   g16009(.A1(new_n16201_), .A2(new_n16196_), .B(\asqrt[17] ), .ZN(new_n16202_));
  NAND2_X1   g16010(.A1(new_n16202_), .A2(new_n13353_), .ZN(new_n16203_));
  OAI21_X1   g16011(.A1(new_n16203_), .A2(new_n15764_), .B(new_n15772_), .ZN(new_n16204_));
  AOI21_X1   g16012(.A1(new_n16204_), .A2(new_n15765_), .B(new_n12913_), .ZN(new_n16205_));
  INV_X1     g16013(.I(new_n15758_), .ZN(new_n16206_));
  AOI21_X1   g16014(.A1(\a[29] ), .A2(new_n16193_), .B(new_n15739_), .ZN(new_n16207_));
  AOI21_X1   g16015(.A1(new_n16207_), .A2(new_n16192_), .B(new_n15729_), .ZN(new_n16208_));
  OAI21_X1   g16016(.A1(new_n16208_), .A2(new_n14601_), .B(new_n14017_), .ZN(new_n16209_));
  OAI21_X1   g16017(.A1(new_n16209_), .A2(new_n16201_), .B(new_n16206_), .ZN(new_n16210_));
  NAND2_X1   g16018(.A1(new_n16210_), .A2(new_n16202_), .ZN(new_n16211_));
  AOI21_X1   g16019(.A1(new_n16211_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n16212_));
  AOI21_X1   g16020(.A1(new_n16212_), .A2(new_n16204_), .B(new_n15780_), .ZN(new_n16213_));
  OAI21_X1   g16021(.A1(new_n16213_), .A2(new_n16205_), .B(\asqrt[20] ), .ZN(new_n16214_));
  NAND2_X1   g16022(.A1(new_n16214_), .A2(new_n11736_), .ZN(new_n16215_));
  OAI21_X1   g16023(.A1(new_n16215_), .A2(new_n15791_), .B(new_n16191_), .ZN(new_n16216_));
  NAND3_X1   g16024(.A1(new_n16216_), .A2(new_n11326_), .A3(new_n15792_), .ZN(new_n16217_));
  AOI22_X1   g16025(.A1(new_n16217_), .A2(new_n15806_), .B1(new_n15814_), .B2(\asqrt[22] ), .ZN(new_n16218_));
  OAI21_X1   g16026(.A1(new_n16218_), .A2(new_n10812_), .B(new_n10221_), .ZN(new_n16219_));
  OAI21_X1   g16027(.A1(new_n16219_), .A2(new_n15816_), .B(new_n16190_), .ZN(new_n16220_));
  AOI21_X1   g16028(.A1(new_n16220_), .A2(new_n15817_), .B(new_n9846_), .ZN(new_n16221_));
  AOI21_X1   g16029(.A1(new_n16216_), .A2(new_n15792_), .B(new_n11326_), .ZN(new_n16222_));
  NOR3_X1    g16030(.A1(new_n16213_), .A2(new_n16205_), .A3(\asqrt[20] ), .ZN(new_n16223_));
  OAI21_X1   g16031(.A1(new_n15788_), .A2(new_n16223_), .B(new_n16214_), .ZN(new_n16224_));
  AOI21_X1   g16032(.A1(new_n16224_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n16225_));
  AOI21_X1   g16033(.A1(new_n16225_), .A2(new_n16216_), .B(new_n15805_), .ZN(new_n16226_));
  NOR3_X1    g16034(.A1(new_n16226_), .A2(\asqrt[23] ), .A3(new_n16222_), .ZN(new_n16227_));
  OAI22_X1   g16035(.A1(new_n16227_), .A2(new_n15813_), .B1(new_n16218_), .B2(new_n10812_), .ZN(new_n16228_));
  AOI21_X1   g16036(.A1(new_n16228_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n16229_));
  AOI21_X1   g16037(.A1(new_n16229_), .A2(new_n16220_), .B(new_n15831_), .ZN(new_n16230_));
  OAI21_X1   g16038(.A1(new_n16230_), .A2(new_n16221_), .B(\asqrt[26] ), .ZN(new_n16231_));
  NAND2_X1   g16039(.A1(new_n16231_), .A2(new_n8826_), .ZN(new_n16232_));
  OAI21_X1   g16040(.A1(new_n16232_), .A2(new_n15842_), .B(new_n16189_), .ZN(new_n16233_));
  AOI21_X1   g16041(.A1(new_n16233_), .A2(new_n15843_), .B(new_n8483_), .ZN(new_n16234_));
  NOR3_X1    g16042(.A1(new_n16230_), .A2(\asqrt[26] ), .A3(new_n16221_), .ZN(new_n16235_));
  OAI21_X1   g16043(.A1(new_n15839_), .A2(new_n16235_), .B(new_n16231_), .ZN(new_n16236_));
  AOI21_X1   g16044(.A1(new_n16236_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n16237_));
  AOI21_X1   g16045(.A1(new_n16237_), .A2(new_n16233_), .B(new_n15857_), .ZN(new_n16238_));
  OAI21_X1   g16046(.A1(new_n16238_), .A2(new_n16234_), .B(\asqrt[29] ), .ZN(new_n16239_));
  NAND2_X1   g16047(.A1(new_n16239_), .A2(new_n7539_), .ZN(new_n16240_));
  OAI21_X1   g16048(.A1(new_n16240_), .A2(new_n15868_), .B(new_n16188_), .ZN(new_n16241_));
  AOI21_X1   g16049(.A1(new_n16241_), .A2(new_n15869_), .B(new_n7229_), .ZN(new_n16242_));
  NOR3_X1    g16050(.A1(new_n16238_), .A2(\asqrt[29] ), .A3(new_n16234_), .ZN(new_n16243_));
  OAI21_X1   g16051(.A1(new_n15865_), .A2(new_n16243_), .B(new_n16239_), .ZN(new_n16244_));
  AOI21_X1   g16052(.A1(new_n16244_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n16245_));
  AOI21_X1   g16053(.A1(new_n16245_), .A2(new_n16241_), .B(new_n15883_), .ZN(new_n16246_));
  OAI21_X1   g16054(.A1(new_n16246_), .A2(new_n16242_), .B(\asqrt[32] ), .ZN(new_n16247_));
  NAND2_X1   g16055(.A1(new_n16247_), .A2(new_n6356_), .ZN(new_n16248_));
  OAI21_X1   g16056(.A1(new_n16248_), .A2(new_n15894_), .B(new_n16187_), .ZN(new_n16249_));
  AOI21_X1   g16057(.A1(new_n16249_), .A2(new_n15895_), .B(new_n6077_), .ZN(new_n16250_));
  NOR3_X1    g16058(.A1(new_n16246_), .A2(\asqrt[32] ), .A3(new_n16242_), .ZN(new_n16251_));
  OAI21_X1   g16059(.A1(new_n15891_), .A2(new_n16251_), .B(new_n16247_), .ZN(new_n16252_));
  AOI21_X1   g16060(.A1(new_n16252_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n16253_));
  AOI21_X1   g16061(.A1(new_n16253_), .A2(new_n16249_), .B(new_n15909_), .ZN(new_n16254_));
  OAI21_X1   g16062(.A1(new_n16254_), .A2(new_n16250_), .B(\asqrt[35] ), .ZN(new_n16255_));
  NAND2_X1   g16063(.A1(new_n16255_), .A2(new_n5277_), .ZN(new_n16256_));
  OAI21_X1   g16064(.A1(new_n16256_), .A2(new_n15920_), .B(new_n16186_), .ZN(new_n16257_));
  AOI21_X1   g16065(.A1(new_n16257_), .A2(new_n15921_), .B(new_n5024_), .ZN(new_n16258_));
  NOR3_X1    g16066(.A1(new_n16254_), .A2(\asqrt[35] ), .A3(new_n16250_), .ZN(new_n16259_));
  OAI21_X1   g16067(.A1(new_n15917_), .A2(new_n16259_), .B(new_n16255_), .ZN(new_n16260_));
  AOI21_X1   g16068(.A1(new_n16260_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n16261_));
  AOI21_X1   g16069(.A1(new_n16261_), .A2(new_n16257_), .B(new_n15935_), .ZN(new_n16262_));
  OAI21_X1   g16070(.A1(new_n16262_), .A2(new_n16258_), .B(\asqrt[38] ), .ZN(new_n16263_));
  NAND2_X1   g16071(.A1(new_n16263_), .A2(new_n4298_), .ZN(new_n16264_));
  OAI21_X1   g16072(.A1(new_n16264_), .A2(new_n15946_), .B(new_n16185_), .ZN(new_n16265_));
  AOI21_X1   g16073(.A1(new_n16265_), .A2(new_n15947_), .B(new_n4071_), .ZN(new_n16266_));
  NOR3_X1    g16074(.A1(new_n16262_), .A2(\asqrt[38] ), .A3(new_n16258_), .ZN(new_n16267_));
  OAI21_X1   g16075(.A1(new_n15943_), .A2(new_n16267_), .B(new_n16263_), .ZN(new_n16268_));
  AOI21_X1   g16076(.A1(new_n16268_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n16269_));
  AOI21_X1   g16077(.A1(new_n16269_), .A2(new_n16265_), .B(new_n15961_), .ZN(new_n16270_));
  OAI21_X1   g16078(.A1(new_n16270_), .A2(new_n16266_), .B(\asqrt[41] ), .ZN(new_n16271_));
  NAND2_X1   g16079(.A1(new_n16271_), .A2(new_n3419_), .ZN(new_n16272_));
  OAI21_X1   g16080(.A1(new_n16272_), .A2(new_n15972_), .B(new_n16184_), .ZN(new_n16273_));
  AOI21_X1   g16081(.A1(new_n16273_), .A2(new_n15973_), .B(new_n3218_), .ZN(new_n16274_));
  NOR3_X1    g16082(.A1(new_n16270_), .A2(\asqrt[41] ), .A3(new_n16266_), .ZN(new_n16275_));
  OAI21_X1   g16083(.A1(new_n15969_), .A2(new_n16275_), .B(new_n16271_), .ZN(new_n16276_));
  AOI21_X1   g16084(.A1(new_n16276_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n16277_));
  AOI21_X1   g16085(.A1(new_n16277_), .A2(new_n16273_), .B(new_n15987_), .ZN(new_n16278_));
  OAI21_X1   g16086(.A1(new_n16278_), .A2(new_n16274_), .B(\asqrt[44] ), .ZN(new_n16279_));
  NAND2_X1   g16087(.A1(new_n16279_), .A2(new_n2641_), .ZN(new_n16280_));
  OAI21_X1   g16088(.A1(new_n16280_), .A2(new_n15998_), .B(new_n16183_), .ZN(new_n16281_));
  AOI21_X1   g16089(.A1(new_n16281_), .A2(new_n15999_), .B(new_n2465_), .ZN(new_n16282_));
  NOR3_X1    g16090(.A1(new_n16278_), .A2(\asqrt[44] ), .A3(new_n16274_), .ZN(new_n16283_));
  OAI21_X1   g16091(.A1(new_n15995_), .A2(new_n16283_), .B(new_n16279_), .ZN(new_n16284_));
  AOI21_X1   g16092(.A1(new_n16284_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n16285_));
  AOI21_X1   g16093(.A1(new_n16285_), .A2(new_n16281_), .B(new_n16013_), .ZN(new_n16286_));
  OAI21_X1   g16094(.A1(new_n16286_), .A2(new_n16282_), .B(\asqrt[47] ), .ZN(new_n16287_));
  NAND2_X1   g16095(.A1(new_n16287_), .A2(new_n1956_), .ZN(new_n16288_));
  OAI21_X1   g16096(.A1(new_n16288_), .A2(new_n16024_), .B(new_n16182_), .ZN(new_n16289_));
  AOI21_X1   g16097(.A1(new_n16289_), .A2(new_n16025_), .B(new_n1806_), .ZN(new_n16290_));
  NOR3_X1    g16098(.A1(new_n16286_), .A2(\asqrt[47] ), .A3(new_n16282_), .ZN(new_n16291_));
  OAI21_X1   g16099(.A1(new_n16021_), .A2(new_n16291_), .B(new_n16287_), .ZN(new_n16292_));
  AOI21_X1   g16100(.A1(new_n16292_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n16293_));
  AOI21_X1   g16101(.A1(new_n16293_), .A2(new_n16289_), .B(new_n16039_), .ZN(new_n16294_));
  OAI21_X1   g16102(.A1(new_n16294_), .A2(new_n16290_), .B(\asqrt[50] ), .ZN(new_n16295_));
  NAND2_X1   g16103(.A1(new_n16295_), .A2(new_n1376_), .ZN(new_n16296_));
  OAI21_X1   g16104(.A1(new_n16296_), .A2(new_n16050_), .B(new_n16181_), .ZN(new_n16297_));
  AOI21_X1   g16105(.A1(new_n16297_), .A2(new_n16051_), .B(new_n1256_), .ZN(new_n16298_));
  NOR3_X1    g16106(.A1(new_n16294_), .A2(\asqrt[50] ), .A3(new_n16290_), .ZN(new_n16299_));
  OAI21_X1   g16107(.A1(new_n16047_), .A2(new_n16299_), .B(new_n16295_), .ZN(new_n16300_));
  AOI21_X1   g16108(.A1(new_n16300_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n16301_));
  AOI21_X1   g16109(.A1(new_n16301_), .A2(new_n16297_), .B(new_n16067_), .ZN(new_n16302_));
  OAI21_X1   g16110(.A1(new_n16302_), .A2(new_n16298_), .B(\asqrt[53] ), .ZN(new_n16303_));
  NAND2_X1   g16111(.A1(new_n16303_), .A2(new_n904_), .ZN(new_n16304_));
  OAI21_X1   g16112(.A1(new_n16304_), .A2(new_n16078_), .B(new_n16180_), .ZN(new_n16305_));
  AOI21_X1   g16113(.A1(new_n16305_), .A2(new_n16079_), .B(new_n823_), .ZN(new_n16306_));
  NOR3_X1    g16114(.A1(new_n16302_), .A2(\asqrt[53] ), .A3(new_n16298_), .ZN(new_n16307_));
  OAI21_X1   g16115(.A1(new_n16075_), .A2(new_n16307_), .B(new_n16303_), .ZN(new_n16308_));
  AOI21_X1   g16116(.A1(new_n16308_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n16309_));
  AOI21_X1   g16117(.A1(new_n16309_), .A2(new_n16305_), .B(new_n16097_), .ZN(new_n16310_));
  OAI21_X1   g16118(.A1(new_n16310_), .A2(new_n16306_), .B(\asqrt[56] ), .ZN(new_n16311_));
  NAND2_X1   g16119(.A1(new_n16311_), .A2(new_n531_), .ZN(new_n16312_));
  OAI21_X1   g16120(.A1(new_n16312_), .A2(new_n16108_), .B(new_n16179_), .ZN(new_n16313_));
  AOI21_X1   g16121(.A1(new_n16313_), .A2(new_n16109_), .B(new_n436_), .ZN(new_n16314_));
  NOR3_X1    g16122(.A1(new_n16310_), .A2(\asqrt[56] ), .A3(new_n16306_), .ZN(new_n16315_));
  OAI21_X1   g16123(.A1(new_n16105_), .A2(new_n16315_), .B(new_n16311_), .ZN(new_n16316_));
  AOI21_X1   g16124(.A1(new_n16316_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n16317_));
  AOI21_X1   g16125(.A1(new_n16317_), .A2(new_n16313_), .B(new_n16128_), .ZN(new_n16318_));
  OAI21_X1   g16126(.A1(new_n16318_), .A2(new_n16314_), .B(\asqrt[59] ), .ZN(new_n16319_));
  NAND2_X1   g16127(.A1(new_n16319_), .A2(new_n306_), .ZN(new_n16320_));
  OAI21_X1   g16128(.A1(new_n16320_), .A2(new_n16139_), .B(new_n16178_), .ZN(new_n16321_));
  NOR3_X1    g16129(.A1(new_n16318_), .A2(\asqrt[59] ), .A3(new_n16314_), .ZN(new_n16322_));
  OAI21_X1   g16130(.A1(new_n16136_), .A2(new_n16322_), .B(new_n16319_), .ZN(new_n16323_));
  AOI21_X1   g16131(.A1(new_n16323_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n16324_));
  AOI21_X1   g16132(.A1(new_n16324_), .A2(new_n16321_), .B(new_n16153_), .ZN(new_n16325_));
  INV_X1     g16133(.I(new_n16161_), .ZN(new_n16326_));
  NAND2_X1   g16134(.A1(new_n16149_), .A2(new_n207_), .ZN(new_n16327_));
  OAI21_X1   g16135(.A1(new_n16327_), .A2(new_n16325_), .B(new_n16326_), .ZN(new_n16328_));
  NOR2_X1    g16136(.A1(new_n16157_), .A2(new_n16173_), .ZN(new_n16329_));
  NAND2_X1   g16137(.A1(\asqrt[14] ), .A2(new_n15692_), .ZN(new_n16330_));
  OAI21_X1   g16138(.A1(new_n15732_), .A2(new_n15725_), .B(\asqrt[63] ), .ZN(new_n16331_));
  AOI21_X1   g16139(.A1(new_n16330_), .A2(new_n15732_), .B(new_n16331_), .ZN(new_n16332_));
  AND2_X2    g16140(.A1(new_n15689_), .A2(new_n15705_), .Z(new_n16333_));
  NAND4_X1   g16141(.A1(new_n15745_), .A2(new_n15691_), .A3(new_n15702_), .A4(new_n16333_), .ZN(new_n16334_));
  NOR2_X1    g16142(.A1(new_n16334_), .A2(new_n15717_), .ZN(new_n16335_));
  NOR2_X1    g16143(.A1(new_n16332_), .A2(new_n16335_), .ZN(new_n16336_));
  INV_X1     g16144(.I(new_n16336_), .ZN(new_n16337_));
  AOI21_X1   g16145(.A1(new_n16329_), .A2(new_n16328_), .B(new_n16337_), .ZN(new_n16338_));
  NAND2_X1   g16146(.A1(new_n16177_), .A2(new_n16338_), .ZN(\asqrt[13] ));
  NOR2_X1    g16147(.A1(\a[24] ), .A2(\a[25] ), .ZN(new_n16340_));
  INV_X1     g16148(.I(new_n16340_), .ZN(new_n16341_));
  NOR2_X1    g16149(.A1(new_n16341_), .A2(\a[26] ), .ZN(new_n16342_));
  INV_X1     g16150(.I(new_n16342_), .ZN(new_n16343_));
  AOI21_X1   g16151(.A1(new_n16321_), .A2(new_n16140_), .B(new_n218_), .ZN(new_n16344_));
  OAI21_X1   g16152(.A1(new_n16325_), .A2(new_n16344_), .B(\asqrt[62] ), .ZN(new_n16345_));
  NOR3_X1    g16153(.A1(new_n16325_), .A2(\asqrt[62] ), .A3(new_n16344_), .ZN(new_n16346_));
  OAI21_X1   g16154(.A1(new_n16161_), .A2(new_n16346_), .B(new_n16345_), .ZN(new_n16347_));
  AOI21_X1   g16155(.A1(new_n16347_), .A2(new_n16175_), .B(\asqrt[63] ), .ZN(new_n16348_));
  NAND2_X1   g16156(.A1(new_n16345_), .A2(new_n16172_), .ZN(new_n16349_));
  OAI21_X1   g16157(.A1(new_n16349_), .A2(new_n16164_), .B(new_n16336_), .ZN(new_n16350_));
  OAI21_X1   g16158(.A1(new_n16348_), .A2(new_n16350_), .B(\a[26] ), .ZN(new_n16351_));
  AOI21_X1   g16159(.A1(new_n16351_), .A2(new_n16343_), .B(new_n15770_), .ZN(new_n16352_));
  INV_X1     g16160(.I(\a[26] ), .ZN(new_n16353_));
  AOI21_X1   g16161(.A1(new_n16177_), .A2(new_n16338_), .B(new_n16353_), .ZN(new_n16354_));
  NAND4_X1   g16162(.A1(new_n15745_), .A2(new_n15702_), .A3(new_n15705_), .A4(new_n16343_), .ZN(new_n16355_));
  NOR2_X1    g16163(.A1(new_n16355_), .A2(new_n15717_), .ZN(new_n16356_));
  INV_X1     g16164(.I(new_n16356_), .ZN(new_n16357_));
  NOR2_X1    g16165(.A1(new_n16354_), .A2(new_n16357_), .ZN(new_n16358_));
  AOI21_X1   g16166(.A1(new_n16177_), .A2(new_n16338_), .B(new_n15712_), .ZN(new_n16359_));
  INV_X1     g16167(.I(\a[27] ), .ZN(new_n16360_));
  AOI21_X1   g16168(.A1(\asqrt[13] ), .A2(new_n16353_), .B(new_n16360_), .ZN(new_n16361_));
  NOR3_X1    g16169(.A1(new_n16358_), .A2(new_n16361_), .A3(new_n16359_), .ZN(new_n16362_));
  OAI21_X1   g16170(.A1(new_n16362_), .A2(new_n16352_), .B(\asqrt[15] ), .ZN(new_n16363_));
  OAI21_X1   g16171(.A1(new_n16348_), .A2(new_n16350_), .B(new_n15711_), .ZN(new_n16364_));
  NAND2_X1   g16172(.A1(new_n16329_), .A2(new_n16328_), .ZN(new_n16365_));
  NOR3_X1    g16173(.A1(new_n16332_), .A2(new_n15770_), .A3(new_n16335_), .ZN(new_n16366_));
  NAND3_X1   g16174(.A1(new_n16177_), .A2(new_n16365_), .A3(new_n16366_), .ZN(new_n16367_));
  AOI21_X1   g16175(.A1(new_n16364_), .A2(new_n16367_), .B(new_n15730_), .ZN(new_n16368_));
  AND3_X2    g16176(.A1(new_n16177_), .A2(new_n16365_), .A3(new_n16366_), .Z(new_n16369_));
  NOR3_X1    g16177(.A1(new_n16369_), .A2(\a[28] ), .A3(new_n16359_), .ZN(new_n16370_));
  OAI21_X1   g16178(.A1(new_n16354_), .A2(new_n16342_), .B(\asqrt[14] ), .ZN(new_n16371_));
  NAND2_X1   g16179(.A1(new_n16371_), .A2(new_n15067_), .ZN(new_n16372_));
  OAI22_X1   g16180(.A1(new_n16362_), .A2(new_n16372_), .B1(new_n16368_), .B2(new_n16370_), .ZN(new_n16373_));
  AOI21_X1   g16181(.A1(new_n16373_), .A2(new_n16363_), .B(new_n14601_), .ZN(new_n16374_));
  NOR3_X1    g16182(.A1(new_n16207_), .A2(new_n15729_), .A3(new_n15738_), .ZN(new_n16375_));
  NAND3_X1   g16183(.A1(\asqrt[13] ), .A2(new_n15759_), .A3(new_n16192_), .ZN(new_n16376_));
  AOI22_X1   g16184(.A1(new_n16376_), .A2(new_n16207_), .B1(\asqrt[13] ), .B2(new_n16375_), .ZN(new_n16377_));
  AOI21_X1   g16185(.A1(new_n16177_), .A2(new_n16338_), .B(\a[26] ), .ZN(new_n16378_));
  OAI21_X1   g16186(.A1(new_n16360_), .A2(new_n16378_), .B(new_n16364_), .ZN(new_n16379_));
  OAI21_X1   g16187(.A1(new_n16379_), .A2(new_n16358_), .B(new_n16371_), .ZN(new_n16380_));
  AOI21_X1   g16188(.A1(new_n16380_), .A2(\asqrt[15] ), .B(\asqrt[16] ), .ZN(new_n16381_));
  AOI21_X1   g16189(.A1(new_n16381_), .A2(new_n16373_), .B(new_n16377_), .ZN(new_n16382_));
  OAI21_X1   g16190(.A1(new_n16382_), .A2(new_n16374_), .B(\asqrt[17] ), .ZN(new_n16383_));
  INV_X1     g16191(.I(new_n16383_), .ZN(new_n16384_));
  NOR2_X1    g16192(.A1(new_n15751_), .A2(new_n15748_), .ZN(new_n16385_));
  NOR2_X1    g16193(.A1(new_n15742_), .A2(new_n15753_), .ZN(new_n16386_));
  INV_X1     g16194(.I(new_n16386_), .ZN(new_n16387_));
  NAND4_X1   g16195(.A1(\asqrt[13] ), .A2(new_n15743_), .A3(new_n16385_), .A4(new_n16387_), .ZN(new_n16388_));
  INV_X1     g16196(.I(\asqrt[13] ), .ZN(new_n16389_));
  NOR3_X1    g16197(.A1(new_n16389_), .A2(new_n16196_), .A3(new_n16386_), .ZN(new_n16390_));
  OAI21_X1   g16198(.A1(new_n16390_), .A2(new_n16385_), .B(new_n16388_), .ZN(new_n16391_));
  INV_X1     g16199(.I(new_n16391_), .ZN(new_n16392_));
  NOR3_X1    g16200(.A1(new_n16382_), .A2(new_n16374_), .A3(\asqrt[17] ), .ZN(new_n16393_));
  NOR2_X1    g16201(.A1(new_n16393_), .A2(new_n16392_), .ZN(new_n16394_));
  OAI21_X1   g16202(.A1(new_n16394_), .A2(new_n16384_), .B(\asqrt[18] ), .ZN(new_n16395_));
  NOR2_X1    g16203(.A1(new_n16209_), .A2(new_n16201_), .ZN(new_n16396_));
  NOR3_X1    g16204(.A1(new_n16389_), .A2(new_n15755_), .A3(new_n16396_), .ZN(new_n16397_));
  INV_X1     g16205(.I(new_n16397_), .ZN(new_n16398_));
  NOR3_X1    g16206(.A1(new_n16396_), .A2(new_n15755_), .A3(new_n16206_), .ZN(new_n16399_));
  AOI22_X1   g16207(.A1(new_n16398_), .A2(new_n16206_), .B1(\asqrt[13] ), .B2(new_n16399_), .ZN(new_n16400_));
  INV_X1     g16208(.I(new_n16400_), .ZN(new_n16401_));
  NAND2_X1   g16209(.A1(new_n16383_), .A2(new_n13353_), .ZN(new_n16402_));
  OAI21_X1   g16210(.A1(new_n16394_), .A2(new_n16402_), .B(new_n16401_), .ZN(new_n16403_));
  AOI21_X1   g16211(.A1(new_n16403_), .A2(new_n16395_), .B(new_n12913_), .ZN(new_n16404_));
  NOR3_X1    g16212(.A1(new_n15766_), .A2(new_n15774_), .A3(new_n15772_), .ZN(new_n16405_));
  NOR3_X1    g16213(.A1(new_n16389_), .A2(new_n15766_), .A3(new_n15774_), .ZN(new_n16406_));
  INV_X1     g16214(.I(new_n16406_), .ZN(new_n16407_));
  AOI22_X1   g16215(.A1(new_n16407_), .A2(new_n15772_), .B1(\asqrt[13] ), .B2(new_n16405_), .ZN(new_n16408_));
  OAI21_X1   g16216(.A1(new_n16392_), .A2(new_n16393_), .B(new_n16383_), .ZN(new_n16409_));
  AOI21_X1   g16217(.A1(new_n16409_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n16410_));
  AOI21_X1   g16218(.A1(new_n16410_), .A2(new_n16403_), .B(new_n16408_), .ZN(new_n16411_));
  OAI21_X1   g16219(.A1(new_n16411_), .A2(new_n16404_), .B(\asqrt[20] ), .ZN(new_n16412_));
  NAND2_X1   g16220(.A1(new_n16212_), .A2(new_n16204_), .ZN(new_n16413_));
  NAND3_X1   g16221(.A1(\asqrt[13] ), .A2(new_n15776_), .A3(new_n16413_), .ZN(new_n16414_));
  AND3_X2    g16222(.A1(new_n15776_), .A2(new_n15780_), .A3(new_n16413_), .Z(new_n16415_));
  AOI22_X1   g16223(.A1(new_n16414_), .A2(new_n15781_), .B1(\asqrt[13] ), .B2(new_n16415_), .ZN(new_n16416_));
  INV_X1     g16224(.I(new_n16416_), .ZN(new_n16417_));
  NAND2_X1   g16225(.A1(new_n16351_), .A2(new_n16356_), .ZN(new_n16418_));
  OAI21_X1   g16226(.A1(new_n16348_), .A2(new_n16350_), .B(new_n16353_), .ZN(new_n16419_));
  NAND2_X1   g16227(.A1(new_n16419_), .A2(\a[27] ), .ZN(new_n16420_));
  NAND3_X1   g16228(.A1(new_n16418_), .A2(new_n16420_), .A3(new_n16364_), .ZN(new_n16421_));
  AOI21_X1   g16229(.A1(new_n16421_), .A2(new_n16371_), .B(new_n15067_), .ZN(new_n16422_));
  OAI21_X1   g16230(.A1(new_n16369_), .A2(new_n16359_), .B(\a[28] ), .ZN(new_n16423_));
  NAND3_X1   g16231(.A1(new_n16364_), .A2(new_n16367_), .A3(new_n15730_), .ZN(new_n16424_));
  NAND2_X1   g16232(.A1(new_n16351_), .A2(new_n16343_), .ZN(new_n16425_));
  AOI21_X1   g16233(.A1(new_n16425_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n16426_));
  AOI22_X1   g16234(.A1(new_n16421_), .A2(new_n16426_), .B1(new_n16423_), .B2(new_n16424_), .ZN(new_n16427_));
  OAI21_X1   g16235(.A1(new_n16427_), .A2(new_n16422_), .B(\asqrt[16] ), .ZN(new_n16428_));
  NAND2_X1   g16236(.A1(new_n16428_), .A2(new_n14017_), .ZN(new_n16429_));
  OAI21_X1   g16237(.A1(new_n16429_), .A2(new_n16382_), .B(new_n16391_), .ZN(new_n16430_));
  AOI21_X1   g16238(.A1(new_n16430_), .A2(new_n16383_), .B(new_n13353_), .ZN(new_n16431_));
  INV_X1     g16239(.I(new_n16377_), .ZN(new_n16432_));
  AOI21_X1   g16240(.A1(\a[27] ), .A2(new_n16419_), .B(new_n16359_), .ZN(new_n16433_));
  AOI21_X1   g16241(.A1(new_n16433_), .A2(new_n16418_), .B(new_n16352_), .ZN(new_n16434_));
  OAI21_X1   g16242(.A1(new_n16434_), .A2(new_n15067_), .B(new_n14601_), .ZN(new_n16435_));
  OAI21_X1   g16243(.A1(new_n16435_), .A2(new_n16427_), .B(new_n16432_), .ZN(new_n16436_));
  NAND2_X1   g16244(.A1(new_n16436_), .A2(new_n16428_), .ZN(new_n16437_));
  AOI21_X1   g16245(.A1(new_n16437_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n16438_));
  AOI21_X1   g16246(.A1(new_n16438_), .A2(new_n16430_), .B(new_n16400_), .ZN(new_n16439_));
  OAI21_X1   g16247(.A1(new_n16439_), .A2(new_n16431_), .B(\asqrt[19] ), .ZN(new_n16440_));
  NAND2_X1   g16248(.A1(new_n16440_), .A2(new_n12364_), .ZN(new_n16441_));
  OAI21_X1   g16249(.A1(new_n16441_), .A2(new_n16411_), .B(new_n16417_), .ZN(new_n16442_));
  AOI21_X1   g16250(.A1(new_n16442_), .A2(new_n16412_), .B(new_n11736_), .ZN(new_n16443_));
  INV_X1     g16251(.I(new_n15788_), .ZN(new_n16444_));
  NOR3_X1    g16252(.A1(new_n15784_), .A2(new_n16223_), .A3(new_n16444_), .ZN(new_n16445_));
  NOR3_X1    g16253(.A1(new_n16389_), .A2(new_n15784_), .A3(new_n16223_), .ZN(new_n16446_));
  INV_X1     g16254(.I(new_n16446_), .ZN(new_n16447_));
  AOI22_X1   g16255(.A1(new_n16447_), .A2(new_n16444_), .B1(\asqrt[13] ), .B2(new_n16445_), .ZN(new_n16448_));
  NOR3_X1    g16256(.A1(new_n16439_), .A2(new_n16431_), .A3(\asqrt[19] ), .ZN(new_n16449_));
  OAI21_X1   g16257(.A1(new_n16408_), .A2(new_n16449_), .B(new_n16440_), .ZN(new_n16450_));
  AOI21_X1   g16258(.A1(new_n16450_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n16451_));
  AOI21_X1   g16259(.A1(new_n16451_), .A2(new_n16442_), .B(new_n16448_), .ZN(new_n16452_));
  OAI21_X1   g16260(.A1(new_n16452_), .A2(new_n16443_), .B(\asqrt[22] ), .ZN(new_n16453_));
  INV_X1     g16261(.I(new_n16453_), .ZN(new_n16454_));
  NOR3_X1    g16262(.A1(new_n16389_), .A2(new_n15793_), .A3(new_n15798_), .ZN(new_n16455_));
  INV_X1     g16263(.I(new_n16455_), .ZN(new_n16456_));
  NOR3_X1    g16264(.A1(new_n15793_), .A2(new_n16191_), .A3(new_n15798_), .ZN(new_n16457_));
  AOI22_X1   g16265(.A1(new_n16456_), .A2(new_n16191_), .B1(\asqrt[13] ), .B2(new_n16457_), .ZN(new_n16458_));
  NOR3_X1    g16266(.A1(new_n16452_), .A2(\asqrt[22] ), .A3(new_n16443_), .ZN(new_n16459_));
  NOR2_X1    g16267(.A1(new_n16459_), .A2(new_n16458_), .ZN(new_n16460_));
  OAI21_X1   g16268(.A1(new_n16460_), .A2(new_n16454_), .B(\asqrt[23] ), .ZN(new_n16461_));
  AND3_X2    g16269(.A1(new_n15800_), .A2(new_n15805_), .A3(new_n16217_), .Z(new_n16462_));
  NAND3_X1   g16270(.A1(\asqrt[13] ), .A2(new_n15800_), .A3(new_n16217_), .ZN(new_n16463_));
  AOI22_X1   g16271(.A1(new_n16463_), .A2(new_n15806_), .B1(\asqrt[13] ), .B2(new_n16462_), .ZN(new_n16464_));
  INV_X1     g16272(.I(new_n16464_), .ZN(new_n16465_));
  NAND2_X1   g16273(.A1(new_n16453_), .A2(new_n10812_), .ZN(new_n16466_));
  OAI21_X1   g16274(.A1(new_n16460_), .A2(new_n16466_), .B(new_n16465_), .ZN(new_n16467_));
  AOI21_X1   g16275(.A1(new_n16467_), .A2(new_n16461_), .B(new_n10221_), .ZN(new_n16468_));
  INV_X1     g16276(.I(new_n15813_), .ZN(new_n16469_));
  NOR3_X1    g16277(.A1(new_n16389_), .A2(new_n15809_), .A3(new_n16227_), .ZN(new_n16470_));
  INV_X1     g16278(.I(new_n16470_), .ZN(new_n16471_));
  NOR3_X1    g16279(.A1(new_n15809_), .A2(new_n16227_), .A3(new_n16469_), .ZN(new_n16472_));
  AOI22_X1   g16280(.A1(new_n16471_), .A2(new_n16469_), .B1(\asqrt[13] ), .B2(new_n16472_), .ZN(new_n16473_));
  NOR3_X1    g16281(.A1(new_n16411_), .A2(new_n16404_), .A3(\asqrt[20] ), .ZN(new_n16474_));
  OAI21_X1   g16282(.A1(new_n16416_), .A2(new_n16474_), .B(new_n16412_), .ZN(new_n16475_));
  INV_X1     g16283(.I(new_n16448_), .ZN(new_n16476_));
  NAND3_X1   g16284(.A1(new_n16442_), .A2(new_n11736_), .A3(new_n16412_), .ZN(new_n16477_));
  AOI22_X1   g16285(.A1(new_n16477_), .A2(new_n16476_), .B1(new_n16475_), .B2(\asqrt[21] ), .ZN(new_n16478_));
  OAI22_X1   g16286(.A1(new_n16459_), .A2(new_n16458_), .B1(new_n16478_), .B2(new_n11326_), .ZN(new_n16479_));
  AOI21_X1   g16287(.A1(new_n16479_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n16480_));
  AOI21_X1   g16288(.A1(new_n16480_), .A2(new_n16467_), .B(new_n16473_), .ZN(new_n16481_));
  OAI21_X1   g16289(.A1(new_n16481_), .A2(new_n16468_), .B(\asqrt[25] ), .ZN(new_n16482_));
  INV_X1     g16290(.I(new_n16482_), .ZN(new_n16483_));
  NOR3_X1    g16291(.A1(new_n15818_), .A2(new_n16190_), .A3(new_n15824_), .ZN(new_n16484_));
  NOR3_X1    g16292(.A1(new_n16389_), .A2(new_n15818_), .A3(new_n15824_), .ZN(new_n16485_));
  INV_X1     g16293(.I(new_n16485_), .ZN(new_n16486_));
  AOI22_X1   g16294(.A1(new_n16486_), .A2(new_n16190_), .B1(\asqrt[13] ), .B2(new_n16484_), .ZN(new_n16487_));
  NOR3_X1    g16295(.A1(new_n16481_), .A2(new_n16468_), .A3(\asqrt[25] ), .ZN(new_n16488_));
  NOR2_X1    g16296(.A1(new_n16488_), .A2(new_n16487_), .ZN(new_n16489_));
  OAI21_X1   g16297(.A1(new_n16489_), .A2(new_n16483_), .B(\asqrt[26] ), .ZN(new_n16490_));
  NOR2_X1    g16298(.A1(new_n15825_), .A2(new_n15833_), .ZN(new_n16491_));
  NOR3_X1    g16299(.A1(new_n16389_), .A2(new_n16221_), .A3(new_n16491_), .ZN(new_n16492_));
  INV_X1     g16300(.I(new_n16492_), .ZN(new_n16493_));
  NOR3_X1    g16301(.A1(new_n16491_), .A2(new_n16221_), .A3(new_n15832_), .ZN(new_n16494_));
  AOI22_X1   g16302(.A1(new_n16493_), .A2(new_n15832_), .B1(\asqrt[13] ), .B2(new_n16494_), .ZN(new_n16495_));
  INV_X1     g16303(.I(new_n16495_), .ZN(new_n16496_));
  NAND2_X1   g16304(.A1(new_n16482_), .A2(new_n9317_), .ZN(new_n16497_));
  OAI21_X1   g16305(.A1(new_n16489_), .A2(new_n16497_), .B(new_n16496_), .ZN(new_n16498_));
  AOI21_X1   g16306(.A1(new_n16498_), .A2(new_n16490_), .B(new_n8826_), .ZN(new_n16499_));
  INV_X1     g16307(.I(new_n15839_), .ZN(new_n16500_));
  NOR3_X1    g16308(.A1(new_n15835_), .A2(new_n16235_), .A3(new_n16500_), .ZN(new_n16501_));
  NOR3_X1    g16309(.A1(new_n16389_), .A2(new_n15835_), .A3(new_n16235_), .ZN(new_n16502_));
  INV_X1     g16310(.I(new_n16502_), .ZN(new_n16503_));
  AOI22_X1   g16311(.A1(new_n16503_), .A2(new_n16500_), .B1(\asqrt[13] ), .B2(new_n16501_), .ZN(new_n16504_));
  OAI21_X1   g16312(.A1(new_n16487_), .A2(new_n16488_), .B(new_n16482_), .ZN(new_n16505_));
  AOI21_X1   g16313(.A1(new_n16505_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n16506_));
  AOI21_X1   g16314(.A1(new_n16506_), .A2(new_n16498_), .B(new_n16504_), .ZN(new_n16507_));
  OAI21_X1   g16315(.A1(new_n16507_), .A2(new_n16499_), .B(\asqrt[28] ), .ZN(new_n16508_));
  INV_X1     g16316(.I(new_n16508_), .ZN(new_n16509_));
  INV_X1     g16317(.I(new_n16507_), .ZN(new_n16510_));
  NOR3_X1    g16318(.A1(new_n16389_), .A2(new_n15844_), .A3(new_n15850_), .ZN(new_n16511_));
  INV_X1     g16319(.I(new_n16511_), .ZN(new_n16512_));
  NOR3_X1    g16320(.A1(new_n15844_), .A2(new_n16189_), .A3(new_n15850_), .ZN(new_n16513_));
  AOI22_X1   g16321(.A1(new_n16512_), .A2(new_n16189_), .B1(\asqrt[13] ), .B2(new_n16513_), .ZN(new_n16514_));
  NOR2_X1    g16322(.A1(new_n16499_), .A2(\asqrt[28] ), .ZN(new_n16515_));
  AOI21_X1   g16323(.A1(new_n16510_), .A2(new_n16515_), .B(new_n16514_), .ZN(new_n16516_));
  OAI21_X1   g16324(.A1(new_n16516_), .A2(new_n16509_), .B(\asqrt[29] ), .ZN(new_n16517_));
  NOR2_X1    g16325(.A1(new_n15851_), .A2(new_n15859_), .ZN(new_n16518_));
  NOR3_X1    g16326(.A1(new_n16518_), .A2(new_n16234_), .A3(new_n15858_), .ZN(new_n16519_));
  NOR3_X1    g16327(.A1(new_n16389_), .A2(new_n16234_), .A3(new_n16518_), .ZN(new_n16520_));
  INV_X1     g16328(.I(new_n16520_), .ZN(new_n16521_));
  AOI22_X1   g16329(.A1(new_n16521_), .A2(new_n15858_), .B1(\asqrt[13] ), .B2(new_n16519_), .ZN(new_n16522_));
  INV_X1     g16330(.I(new_n16522_), .ZN(new_n16523_));
  NAND2_X1   g16331(.A1(new_n16508_), .A2(new_n8036_), .ZN(new_n16524_));
  OAI21_X1   g16332(.A1(new_n16524_), .A2(new_n16516_), .B(new_n16523_), .ZN(new_n16525_));
  AOI21_X1   g16333(.A1(new_n16525_), .A2(new_n16517_), .B(new_n7539_), .ZN(new_n16526_));
  INV_X1     g16334(.I(new_n16526_), .ZN(new_n16527_));
  INV_X1     g16335(.I(new_n16525_), .ZN(new_n16528_));
  INV_X1     g16336(.I(new_n15865_), .ZN(new_n16529_));
  NOR3_X1    g16337(.A1(new_n16389_), .A2(new_n15861_), .A3(new_n16243_), .ZN(new_n16530_));
  INV_X1     g16338(.I(new_n16530_), .ZN(new_n16531_));
  NOR3_X1    g16339(.A1(new_n15861_), .A2(new_n16243_), .A3(new_n16529_), .ZN(new_n16532_));
  AOI22_X1   g16340(.A1(new_n16531_), .A2(new_n16529_), .B1(\asqrt[13] ), .B2(new_n16532_), .ZN(new_n16533_));
  INV_X1     g16341(.I(new_n16533_), .ZN(new_n16534_));
  NAND2_X1   g16342(.A1(new_n16517_), .A2(new_n7539_), .ZN(new_n16535_));
  OAI21_X1   g16343(.A1(new_n16535_), .A2(new_n16528_), .B(new_n16534_), .ZN(new_n16536_));
  AOI21_X1   g16344(.A1(new_n16536_), .A2(new_n16527_), .B(new_n7229_), .ZN(new_n16537_));
  NOR3_X1    g16345(.A1(new_n15870_), .A2(new_n16188_), .A3(new_n15876_), .ZN(new_n16538_));
  NOR3_X1    g16346(.A1(new_n16389_), .A2(new_n15870_), .A3(new_n15876_), .ZN(new_n16539_));
  INV_X1     g16347(.I(new_n16539_), .ZN(new_n16540_));
  AOI22_X1   g16348(.A1(new_n16540_), .A2(new_n16188_), .B1(\asqrt[13] ), .B2(new_n16538_), .ZN(new_n16541_));
  NOR2_X1    g16349(.A1(new_n16526_), .A2(\asqrt[31] ), .ZN(new_n16542_));
  AOI21_X1   g16350(.A1(new_n16542_), .A2(new_n16536_), .B(new_n16541_), .ZN(new_n16543_));
  OAI21_X1   g16351(.A1(new_n16543_), .A2(new_n16537_), .B(\asqrt[32] ), .ZN(new_n16544_));
  NOR2_X1    g16352(.A1(new_n15877_), .A2(new_n15885_), .ZN(new_n16545_));
  NOR3_X1    g16353(.A1(new_n16389_), .A2(new_n16242_), .A3(new_n16545_), .ZN(new_n16546_));
  INV_X1     g16354(.I(new_n16546_), .ZN(new_n16547_));
  NOR3_X1    g16355(.A1(new_n16545_), .A2(new_n16242_), .A3(new_n15884_), .ZN(new_n16548_));
  AOI22_X1   g16356(.A1(new_n16547_), .A2(new_n15884_), .B1(\asqrt[13] ), .B2(new_n16548_), .ZN(new_n16549_));
  INV_X1     g16357(.I(new_n16549_), .ZN(new_n16550_));
  NOR3_X1    g16358(.A1(new_n16507_), .A2(new_n16499_), .A3(\asqrt[28] ), .ZN(new_n16551_));
  OAI21_X1   g16359(.A1(new_n16514_), .A2(new_n16551_), .B(new_n16508_), .ZN(new_n16552_));
  AOI21_X1   g16360(.A1(new_n16552_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n16553_));
  AOI21_X1   g16361(.A1(new_n16553_), .A2(new_n16525_), .B(new_n16533_), .ZN(new_n16554_));
  OAI21_X1   g16362(.A1(new_n16554_), .A2(new_n16526_), .B(\asqrt[31] ), .ZN(new_n16555_));
  NAND2_X1   g16363(.A1(new_n16555_), .A2(new_n6824_), .ZN(new_n16556_));
  OAI21_X1   g16364(.A1(new_n16556_), .A2(new_n16543_), .B(new_n16550_), .ZN(new_n16557_));
  AOI21_X1   g16365(.A1(new_n16557_), .A2(new_n16544_), .B(new_n6356_), .ZN(new_n16558_));
  INV_X1     g16366(.I(new_n16558_), .ZN(new_n16559_));
  INV_X1     g16367(.I(new_n16557_), .ZN(new_n16560_));
  INV_X1     g16368(.I(new_n15891_), .ZN(new_n16561_));
  NOR3_X1    g16369(.A1(new_n15887_), .A2(new_n16251_), .A3(new_n16561_), .ZN(new_n16562_));
  NOR3_X1    g16370(.A1(new_n16389_), .A2(new_n15887_), .A3(new_n16251_), .ZN(new_n16563_));
  INV_X1     g16371(.I(new_n16563_), .ZN(new_n16564_));
  AOI22_X1   g16372(.A1(new_n16564_), .A2(new_n16561_), .B1(\asqrt[13] ), .B2(new_n16562_), .ZN(new_n16565_));
  INV_X1     g16373(.I(new_n16565_), .ZN(new_n16566_));
  NAND2_X1   g16374(.A1(new_n16544_), .A2(new_n6356_), .ZN(new_n16567_));
  OAI21_X1   g16375(.A1(new_n16567_), .A2(new_n16560_), .B(new_n16566_), .ZN(new_n16568_));
  AOI21_X1   g16376(.A1(new_n16568_), .A2(new_n16559_), .B(new_n6077_), .ZN(new_n16569_));
  NOR3_X1    g16377(.A1(new_n16389_), .A2(new_n15896_), .A3(new_n15902_), .ZN(new_n16570_));
  INV_X1     g16378(.I(new_n16570_), .ZN(new_n16571_));
  NOR3_X1    g16379(.A1(new_n15896_), .A2(new_n16187_), .A3(new_n15902_), .ZN(new_n16572_));
  AOI22_X1   g16380(.A1(new_n16571_), .A2(new_n16187_), .B1(\asqrt[13] ), .B2(new_n16572_), .ZN(new_n16573_));
  NOR2_X1    g16381(.A1(new_n16558_), .A2(\asqrt[34] ), .ZN(new_n16574_));
  AOI21_X1   g16382(.A1(new_n16574_), .A2(new_n16568_), .B(new_n16573_), .ZN(new_n16575_));
  OAI21_X1   g16383(.A1(new_n16575_), .A2(new_n16569_), .B(\asqrt[35] ), .ZN(new_n16576_));
  NOR2_X1    g16384(.A1(new_n15903_), .A2(new_n15911_), .ZN(new_n16577_));
  NOR3_X1    g16385(.A1(new_n16577_), .A2(new_n16250_), .A3(new_n15910_), .ZN(new_n16578_));
  NOR3_X1    g16386(.A1(new_n16389_), .A2(new_n16250_), .A3(new_n16577_), .ZN(new_n16579_));
  INV_X1     g16387(.I(new_n16579_), .ZN(new_n16580_));
  AOI22_X1   g16388(.A1(new_n16580_), .A2(new_n15910_), .B1(\asqrt[13] ), .B2(new_n16578_), .ZN(new_n16581_));
  INV_X1     g16389(.I(new_n16581_), .ZN(new_n16582_));
  NOR3_X1    g16390(.A1(new_n16554_), .A2(\asqrt[31] ), .A3(new_n16526_), .ZN(new_n16583_));
  OAI21_X1   g16391(.A1(new_n16541_), .A2(new_n16583_), .B(new_n16555_), .ZN(new_n16584_));
  AOI21_X1   g16392(.A1(new_n16584_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n16585_));
  AOI21_X1   g16393(.A1(new_n16585_), .A2(new_n16557_), .B(new_n16565_), .ZN(new_n16586_));
  OAI21_X1   g16394(.A1(new_n16586_), .A2(new_n16558_), .B(\asqrt[34] ), .ZN(new_n16587_));
  NAND2_X1   g16395(.A1(new_n16587_), .A2(new_n5708_), .ZN(new_n16588_));
  OAI21_X1   g16396(.A1(new_n16588_), .A2(new_n16575_), .B(new_n16582_), .ZN(new_n16589_));
  NAND2_X1   g16397(.A1(new_n16589_), .A2(new_n16576_), .ZN(new_n16590_));
  NAND2_X1   g16398(.A1(new_n16590_), .A2(\asqrt[36] ), .ZN(new_n16591_));
  INV_X1     g16399(.I(new_n16589_), .ZN(new_n16592_));
  INV_X1     g16400(.I(new_n15917_), .ZN(new_n16593_));
  NOR3_X1    g16401(.A1(new_n16389_), .A2(new_n15913_), .A3(new_n16259_), .ZN(new_n16594_));
  INV_X1     g16402(.I(new_n16594_), .ZN(new_n16595_));
  NOR3_X1    g16403(.A1(new_n15913_), .A2(new_n16259_), .A3(new_n16593_), .ZN(new_n16596_));
  AOI22_X1   g16404(.A1(new_n16595_), .A2(new_n16593_), .B1(\asqrt[13] ), .B2(new_n16596_), .ZN(new_n16597_));
  INV_X1     g16405(.I(new_n16597_), .ZN(new_n16598_));
  NAND2_X1   g16406(.A1(new_n16576_), .A2(new_n5277_), .ZN(new_n16599_));
  OAI21_X1   g16407(.A1(new_n16592_), .A2(new_n16599_), .B(new_n16598_), .ZN(new_n16600_));
  AOI21_X1   g16408(.A1(new_n16600_), .A2(new_n16591_), .B(new_n5024_), .ZN(new_n16601_));
  NOR3_X1    g16409(.A1(new_n15922_), .A2(new_n16186_), .A3(new_n15928_), .ZN(new_n16602_));
  NOR3_X1    g16410(.A1(new_n16389_), .A2(new_n15922_), .A3(new_n15928_), .ZN(new_n16603_));
  INV_X1     g16411(.I(new_n16603_), .ZN(new_n16604_));
  AOI22_X1   g16412(.A1(new_n16604_), .A2(new_n16186_), .B1(\asqrt[13] ), .B2(new_n16602_), .ZN(new_n16605_));
  AOI21_X1   g16413(.A1(new_n16589_), .A2(new_n16576_), .B(new_n5277_), .ZN(new_n16606_));
  NOR2_X1    g16414(.A1(new_n16606_), .A2(\asqrt[37] ), .ZN(new_n16607_));
  AOI21_X1   g16415(.A1(new_n16607_), .A2(new_n16600_), .B(new_n16605_), .ZN(new_n16608_));
  OAI21_X1   g16416(.A1(new_n16608_), .A2(new_n16601_), .B(\asqrt[38] ), .ZN(new_n16609_));
  INV_X1     g16417(.I(new_n16609_), .ZN(new_n16610_));
  NOR2_X1    g16418(.A1(new_n15929_), .A2(new_n15937_), .ZN(new_n16611_));
  NOR3_X1    g16419(.A1(new_n16389_), .A2(new_n16258_), .A3(new_n16611_), .ZN(new_n16612_));
  INV_X1     g16420(.I(new_n16612_), .ZN(new_n16613_));
  NOR3_X1    g16421(.A1(new_n16611_), .A2(new_n16258_), .A3(new_n15936_), .ZN(new_n16614_));
  AOI22_X1   g16422(.A1(new_n16613_), .A2(new_n15936_), .B1(\asqrt[13] ), .B2(new_n16614_), .ZN(new_n16615_));
  NOR3_X1    g16423(.A1(new_n16608_), .A2(new_n16601_), .A3(\asqrt[38] ), .ZN(new_n16616_));
  NOR2_X1    g16424(.A1(new_n16616_), .A2(new_n16615_), .ZN(new_n16617_));
  OAI21_X1   g16425(.A1(new_n16617_), .A2(new_n16610_), .B(\asqrt[39] ), .ZN(new_n16618_));
  INV_X1     g16426(.I(new_n15943_), .ZN(new_n16619_));
  NOR3_X1    g16427(.A1(new_n15939_), .A2(new_n16267_), .A3(new_n16619_), .ZN(new_n16620_));
  NOR3_X1    g16428(.A1(new_n16389_), .A2(new_n15939_), .A3(new_n16267_), .ZN(new_n16621_));
  INV_X1     g16429(.I(new_n16621_), .ZN(new_n16622_));
  AOI22_X1   g16430(.A1(new_n16622_), .A2(new_n16619_), .B1(\asqrt[13] ), .B2(new_n16620_), .ZN(new_n16623_));
  INV_X1     g16431(.I(new_n16623_), .ZN(new_n16624_));
  NAND2_X1   g16432(.A1(new_n16609_), .A2(new_n4298_), .ZN(new_n16625_));
  OAI21_X1   g16433(.A1(new_n16617_), .A2(new_n16625_), .B(new_n16624_), .ZN(new_n16626_));
  AOI21_X1   g16434(.A1(new_n16626_), .A2(new_n16618_), .B(new_n4071_), .ZN(new_n16627_));
  NOR3_X1    g16435(.A1(new_n16389_), .A2(new_n15948_), .A3(new_n15954_), .ZN(new_n16628_));
  INV_X1     g16436(.I(new_n16628_), .ZN(new_n16629_));
  NOR3_X1    g16437(.A1(new_n15948_), .A2(new_n16185_), .A3(new_n15954_), .ZN(new_n16630_));
  AOI22_X1   g16438(.A1(new_n16629_), .A2(new_n16185_), .B1(\asqrt[13] ), .B2(new_n16630_), .ZN(new_n16631_));
  INV_X1     g16439(.I(new_n16615_), .ZN(new_n16632_));
  NOR3_X1    g16440(.A1(new_n16586_), .A2(\asqrt[34] ), .A3(new_n16558_), .ZN(new_n16633_));
  OAI21_X1   g16441(.A1(new_n16573_), .A2(new_n16633_), .B(new_n16587_), .ZN(new_n16634_));
  AOI21_X1   g16442(.A1(new_n16634_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n16635_));
  AOI21_X1   g16443(.A1(new_n16635_), .A2(new_n16589_), .B(new_n16597_), .ZN(new_n16636_));
  OAI21_X1   g16444(.A1(new_n16636_), .A2(new_n16606_), .B(\asqrt[37] ), .ZN(new_n16637_));
  NAND2_X1   g16445(.A1(new_n16637_), .A2(new_n4696_), .ZN(new_n16638_));
  OAI21_X1   g16446(.A1(new_n16638_), .A2(new_n16608_), .B(new_n16632_), .ZN(new_n16639_));
  AOI21_X1   g16447(.A1(new_n16639_), .A2(new_n16609_), .B(new_n4298_), .ZN(new_n16640_));
  NOR2_X1    g16448(.A1(new_n16640_), .A2(\asqrt[40] ), .ZN(new_n16641_));
  AOI21_X1   g16449(.A1(new_n16641_), .A2(new_n16626_), .B(new_n16631_), .ZN(new_n16642_));
  OAI21_X1   g16450(.A1(new_n16642_), .A2(new_n16627_), .B(\asqrt[41] ), .ZN(new_n16643_));
  NOR2_X1    g16451(.A1(new_n15955_), .A2(new_n15963_), .ZN(new_n16644_));
  NOR3_X1    g16452(.A1(new_n16644_), .A2(new_n16266_), .A3(new_n15962_), .ZN(new_n16645_));
  NOR3_X1    g16453(.A1(new_n16389_), .A2(new_n16266_), .A3(new_n16644_), .ZN(new_n16646_));
  INV_X1     g16454(.I(new_n16646_), .ZN(new_n16647_));
  AOI22_X1   g16455(.A1(new_n16647_), .A2(new_n15962_), .B1(\asqrt[13] ), .B2(new_n16645_), .ZN(new_n16648_));
  INV_X1     g16456(.I(new_n16648_), .ZN(new_n16649_));
  NOR3_X1    g16457(.A1(new_n16636_), .A2(\asqrt[37] ), .A3(new_n16606_), .ZN(new_n16650_));
  OAI21_X1   g16458(.A1(new_n16605_), .A2(new_n16650_), .B(new_n16637_), .ZN(new_n16651_));
  AOI21_X1   g16459(.A1(new_n16651_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n16652_));
  AOI21_X1   g16460(.A1(new_n16652_), .A2(new_n16639_), .B(new_n16623_), .ZN(new_n16653_));
  OAI21_X1   g16461(.A1(new_n16653_), .A2(new_n16640_), .B(\asqrt[40] ), .ZN(new_n16654_));
  NAND2_X1   g16462(.A1(new_n16654_), .A2(new_n3782_), .ZN(new_n16655_));
  OAI21_X1   g16463(.A1(new_n16655_), .A2(new_n16642_), .B(new_n16649_), .ZN(new_n16656_));
  AOI21_X1   g16464(.A1(new_n16656_), .A2(new_n16643_), .B(new_n3419_), .ZN(new_n16657_));
  INV_X1     g16465(.I(new_n15969_), .ZN(new_n16658_));
  NOR3_X1    g16466(.A1(new_n16389_), .A2(new_n15965_), .A3(new_n16275_), .ZN(new_n16659_));
  INV_X1     g16467(.I(new_n16659_), .ZN(new_n16660_));
  NOR3_X1    g16468(.A1(new_n15965_), .A2(new_n16275_), .A3(new_n16658_), .ZN(new_n16661_));
  AOI22_X1   g16469(.A1(new_n16660_), .A2(new_n16658_), .B1(\asqrt[13] ), .B2(new_n16661_), .ZN(new_n16662_));
  NOR3_X1    g16470(.A1(new_n16653_), .A2(\asqrt[40] ), .A3(new_n16640_), .ZN(new_n16663_));
  OAI21_X1   g16471(.A1(new_n16631_), .A2(new_n16663_), .B(new_n16654_), .ZN(new_n16664_));
  AOI21_X1   g16472(.A1(new_n16664_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n16665_));
  AOI21_X1   g16473(.A1(new_n16665_), .A2(new_n16656_), .B(new_n16662_), .ZN(new_n16666_));
  OAI21_X1   g16474(.A1(new_n16666_), .A2(new_n16657_), .B(\asqrt[43] ), .ZN(new_n16667_));
  INV_X1     g16475(.I(new_n16667_), .ZN(new_n16668_));
  NOR3_X1    g16476(.A1(new_n15974_), .A2(new_n16184_), .A3(new_n15980_), .ZN(new_n16669_));
  NOR3_X1    g16477(.A1(new_n16389_), .A2(new_n15974_), .A3(new_n15980_), .ZN(new_n16670_));
  INV_X1     g16478(.I(new_n16670_), .ZN(new_n16671_));
  AOI22_X1   g16479(.A1(new_n16671_), .A2(new_n16184_), .B1(\asqrt[13] ), .B2(new_n16669_), .ZN(new_n16672_));
  NOR3_X1    g16480(.A1(new_n16666_), .A2(\asqrt[43] ), .A3(new_n16657_), .ZN(new_n16673_));
  NOR2_X1    g16481(.A1(new_n16673_), .A2(new_n16672_), .ZN(new_n16674_));
  OAI21_X1   g16482(.A1(new_n16674_), .A2(new_n16668_), .B(\asqrt[44] ), .ZN(new_n16675_));
  NOR2_X1    g16483(.A1(new_n15981_), .A2(new_n15989_), .ZN(new_n16676_));
  NOR3_X1    g16484(.A1(new_n16389_), .A2(new_n16274_), .A3(new_n16676_), .ZN(new_n16677_));
  INV_X1     g16485(.I(new_n16677_), .ZN(new_n16678_));
  NOR3_X1    g16486(.A1(new_n16676_), .A2(new_n16274_), .A3(new_n15988_), .ZN(new_n16679_));
  AOI22_X1   g16487(.A1(new_n16678_), .A2(new_n15988_), .B1(\asqrt[13] ), .B2(new_n16679_), .ZN(new_n16680_));
  INV_X1     g16488(.I(new_n16680_), .ZN(new_n16681_));
  NAND2_X1   g16489(.A1(new_n16667_), .A2(new_n2954_), .ZN(new_n16682_));
  OAI21_X1   g16490(.A1(new_n16674_), .A2(new_n16682_), .B(new_n16681_), .ZN(new_n16683_));
  AOI21_X1   g16491(.A1(new_n16683_), .A2(new_n16675_), .B(new_n2641_), .ZN(new_n16684_));
  INV_X1     g16492(.I(new_n15995_), .ZN(new_n16685_));
  NOR3_X1    g16493(.A1(new_n15991_), .A2(new_n16283_), .A3(new_n16685_), .ZN(new_n16686_));
  NOR3_X1    g16494(.A1(new_n16389_), .A2(new_n15991_), .A3(new_n16283_), .ZN(new_n16687_));
  INV_X1     g16495(.I(new_n16687_), .ZN(new_n16688_));
  AOI22_X1   g16496(.A1(new_n16688_), .A2(new_n16685_), .B1(\asqrt[13] ), .B2(new_n16686_), .ZN(new_n16689_));
  OAI21_X1   g16497(.A1(new_n16672_), .A2(new_n16673_), .B(new_n16667_), .ZN(new_n16690_));
  AOI21_X1   g16498(.A1(new_n16690_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n16691_));
  AOI21_X1   g16499(.A1(new_n16691_), .A2(new_n16683_), .B(new_n16689_), .ZN(new_n16692_));
  OAI21_X1   g16500(.A1(new_n16692_), .A2(new_n16684_), .B(\asqrt[46] ), .ZN(new_n16693_));
  INV_X1     g16501(.I(new_n16693_), .ZN(new_n16694_));
  NOR3_X1    g16502(.A1(new_n16389_), .A2(new_n16000_), .A3(new_n16006_), .ZN(new_n16695_));
  INV_X1     g16503(.I(new_n16695_), .ZN(new_n16696_));
  NOR3_X1    g16504(.A1(new_n16000_), .A2(new_n16183_), .A3(new_n16006_), .ZN(new_n16697_));
  AOI22_X1   g16505(.A1(new_n16696_), .A2(new_n16183_), .B1(\asqrt[13] ), .B2(new_n16697_), .ZN(new_n16698_));
  NOR3_X1    g16506(.A1(new_n16692_), .A2(new_n16684_), .A3(\asqrt[46] ), .ZN(new_n16699_));
  NOR2_X1    g16507(.A1(new_n16699_), .A2(new_n16698_), .ZN(new_n16700_));
  OAI21_X1   g16508(.A1(new_n16700_), .A2(new_n16694_), .B(\asqrt[47] ), .ZN(new_n16701_));
  NOR2_X1    g16509(.A1(new_n16007_), .A2(new_n16015_), .ZN(new_n16702_));
  NOR3_X1    g16510(.A1(new_n16702_), .A2(new_n16282_), .A3(new_n16014_), .ZN(new_n16703_));
  NOR3_X1    g16511(.A1(new_n16389_), .A2(new_n16282_), .A3(new_n16702_), .ZN(new_n16704_));
  INV_X1     g16512(.I(new_n16704_), .ZN(new_n16705_));
  AOI22_X1   g16513(.A1(new_n16705_), .A2(new_n16014_), .B1(\asqrt[13] ), .B2(new_n16703_), .ZN(new_n16706_));
  INV_X1     g16514(.I(new_n16706_), .ZN(new_n16707_));
  NAND2_X1   g16515(.A1(new_n16693_), .A2(new_n2229_), .ZN(new_n16708_));
  OAI21_X1   g16516(.A1(new_n16700_), .A2(new_n16708_), .B(new_n16707_), .ZN(new_n16709_));
  AOI21_X1   g16517(.A1(new_n16709_), .A2(new_n16701_), .B(new_n1956_), .ZN(new_n16710_));
  INV_X1     g16518(.I(new_n16021_), .ZN(new_n16711_));
  NOR3_X1    g16519(.A1(new_n16389_), .A2(new_n16017_), .A3(new_n16291_), .ZN(new_n16712_));
  INV_X1     g16520(.I(new_n16712_), .ZN(new_n16713_));
  NOR3_X1    g16521(.A1(new_n16017_), .A2(new_n16291_), .A3(new_n16711_), .ZN(new_n16714_));
  AOI22_X1   g16522(.A1(new_n16713_), .A2(new_n16711_), .B1(\asqrt[13] ), .B2(new_n16714_), .ZN(new_n16715_));
  OAI21_X1   g16523(.A1(new_n16698_), .A2(new_n16699_), .B(new_n16693_), .ZN(new_n16716_));
  AOI21_X1   g16524(.A1(new_n16716_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n16717_));
  AOI21_X1   g16525(.A1(new_n16717_), .A2(new_n16709_), .B(new_n16715_), .ZN(new_n16718_));
  OAI21_X1   g16526(.A1(new_n16718_), .A2(new_n16710_), .B(\asqrt[49] ), .ZN(new_n16719_));
  INV_X1     g16527(.I(new_n16719_), .ZN(new_n16720_));
  NOR3_X1    g16528(.A1(new_n16026_), .A2(new_n16182_), .A3(new_n16032_), .ZN(new_n16721_));
  NOR3_X1    g16529(.A1(new_n16389_), .A2(new_n16026_), .A3(new_n16032_), .ZN(new_n16722_));
  INV_X1     g16530(.I(new_n16722_), .ZN(new_n16723_));
  AOI22_X1   g16531(.A1(new_n16723_), .A2(new_n16182_), .B1(\asqrt[13] ), .B2(new_n16721_), .ZN(new_n16724_));
  NOR3_X1    g16532(.A1(new_n16718_), .A2(new_n16710_), .A3(\asqrt[49] ), .ZN(new_n16725_));
  NOR2_X1    g16533(.A1(new_n16725_), .A2(new_n16724_), .ZN(new_n16726_));
  OAI21_X1   g16534(.A1(new_n16726_), .A2(new_n16720_), .B(\asqrt[50] ), .ZN(new_n16727_));
  NOR2_X1    g16535(.A1(new_n16033_), .A2(new_n16041_), .ZN(new_n16728_));
  NOR3_X1    g16536(.A1(new_n16389_), .A2(new_n16290_), .A3(new_n16728_), .ZN(new_n16729_));
  INV_X1     g16537(.I(new_n16729_), .ZN(new_n16730_));
  NOR3_X1    g16538(.A1(new_n16728_), .A2(new_n16290_), .A3(new_n16040_), .ZN(new_n16731_));
  AOI22_X1   g16539(.A1(new_n16730_), .A2(new_n16040_), .B1(\asqrt[13] ), .B2(new_n16731_), .ZN(new_n16732_));
  INV_X1     g16540(.I(new_n16732_), .ZN(new_n16733_));
  NAND2_X1   g16541(.A1(new_n16719_), .A2(new_n1612_), .ZN(new_n16734_));
  OAI21_X1   g16542(.A1(new_n16726_), .A2(new_n16734_), .B(new_n16733_), .ZN(new_n16735_));
  AOI21_X1   g16543(.A1(new_n16735_), .A2(new_n16727_), .B(new_n1376_), .ZN(new_n16736_));
  INV_X1     g16544(.I(new_n16047_), .ZN(new_n16737_));
  NOR3_X1    g16545(.A1(new_n16043_), .A2(new_n16299_), .A3(new_n16737_), .ZN(new_n16738_));
  NOR3_X1    g16546(.A1(new_n16389_), .A2(new_n16043_), .A3(new_n16299_), .ZN(new_n16739_));
  INV_X1     g16547(.I(new_n16739_), .ZN(new_n16740_));
  AOI22_X1   g16548(.A1(new_n16740_), .A2(new_n16737_), .B1(\asqrt[13] ), .B2(new_n16738_), .ZN(new_n16741_));
  OAI21_X1   g16549(.A1(new_n16724_), .A2(new_n16725_), .B(new_n16719_), .ZN(new_n16742_));
  AOI21_X1   g16550(.A1(new_n16742_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n16743_));
  AOI21_X1   g16551(.A1(new_n16743_), .A2(new_n16735_), .B(new_n16741_), .ZN(new_n16744_));
  OAI21_X1   g16552(.A1(new_n16744_), .A2(new_n16736_), .B(\asqrt[52] ), .ZN(new_n16745_));
  INV_X1     g16553(.I(new_n16745_), .ZN(new_n16746_));
  INV_X1     g16554(.I(new_n16744_), .ZN(new_n16747_));
  NOR3_X1    g16555(.A1(new_n16389_), .A2(new_n16052_), .A3(new_n16058_), .ZN(new_n16748_));
  INV_X1     g16556(.I(new_n16748_), .ZN(new_n16749_));
  NOR3_X1    g16557(.A1(new_n16052_), .A2(new_n16181_), .A3(new_n16058_), .ZN(new_n16750_));
  AOI22_X1   g16558(.A1(new_n16749_), .A2(new_n16181_), .B1(\asqrt[13] ), .B2(new_n16750_), .ZN(new_n16751_));
  NOR2_X1    g16559(.A1(new_n16736_), .A2(\asqrt[52] ), .ZN(new_n16752_));
  AOI21_X1   g16560(.A1(new_n16747_), .A2(new_n16752_), .B(new_n16751_), .ZN(new_n16753_));
  OAI21_X1   g16561(.A1(new_n16753_), .A2(new_n16746_), .B(\asqrt[53] ), .ZN(new_n16754_));
  NOR2_X1    g16562(.A1(new_n16059_), .A2(new_n16069_), .ZN(new_n16755_));
  NOR3_X1    g16563(.A1(new_n16755_), .A2(new_n16298_), .A3(new_n16068_), .ZN(new_n16756_));
  NOR3_X1    g16564(.A1(new_n16389_), .A2(new_n16298_), .A3(new_n16755_), .ZN(new_n16757_));
  INV_X1     g16565(.I(new_n16757_), .ZN(new_n16758_));
  AOI22_X1   g16566(.A1(new_n16758_), .A2(new_n16068_), .B1(\asqrt[13] ), .B2(new_n16756_), .ZN(new_n16759_));
  INV_X1     g16567(.I(new_n16759_), .ZN(new_n16760_));
  NAND2_X1   g16568(.A1(new_n16745_), .A2(new_n1103_), .ZN(new_n16761_));
  OAI21_X1   g16569(.A1(new_n16761_), .A2(new_n16753_), .B(new_n16760_), .ZN(new_n16762_));
  AOI21_X1   g16570(.A1(new_n16762_), .A2(new_n16754_), .B(new_n904_), .ZN(new_n16763_));
  INV_X1     g16571(.I(new_n16763_), .ZN(new_n16764_));
  INV_X1     g16572(.I(new_n16762_), .ZN(new_n16765_));
  INV_X1     g16573(.I(new_n16075_), .ZN(new_n16766_));
  NOR3_X1    g16574(.A1(new_n16389_), .A2(new_n16071_), .A3(new_n16307_), .ZN(new_n16767_));
  INV_X1     g16575(.I(new_n16767_), .ZN(new_n16768_));
  NOR3_X1    g16576(.A1(new_n16071_), .A2(new_n16307_), .A3(new_n16766_), .ZN(new_n16769_));
  AOI22_X1   g16577(.A1(new_n16768_), .A2(new_n16766_), .B1(\asqrt[13] ), .B2(new_n16769_), .ZN(new_n16770_));
  INV_X1     g16578(.I(new_n16770_), .ZN(new_n16771_));
  NAND2_X1   g16579(.A1(new_n16754_), .A2(new_n904_), .ZN(new_n16772_));
  OAI21_X1   g16580(.A1(new_n16772_), .A2(new_n16765_), .B(new_n16771_), .ZN(new_n16773_));
  AOI21_X1   g16581(.A1(new_n16773_), .A2(new_n16764_), .B(new_n823_), .ZN(new_n16774_));
  NOR3_X1    g16582(.A1(new_n16080_), .A2(new_n16180_), .A3(new_n16087_), .ZN(new_n16775_));
  NOR3_X1    g16583(.A1(new_n16389_), .A2(new_n16080_), .A3(new_n16087_), .ZN(new_n16776_));
  INV_X1     g16584(.I(new_n16776_), .ZN(new_n16777_));
  AOI22_X1   g16585(.A1(new_n16777_), .A2(new_n16180_), .B1(\asqrt[13] ), .B2(new_n16775_), .ZN(new_n16778_));
  NOR2_X1    g16586(.A1(new_n16763_), .A2(\asqrt[55] ), .ZN(new_n16779_));
  AOI21_X1   g16587(.A1(new_n16779_), .A2(new_n16773_), .B(new_n16778_), .ZN(new_n16780_));
  OAI21_X1   g16588(.A1(new_n16780_), .A2(new_n16774_), .B(\asqrt[56] ), .ZN(new_n16781_));
  NOR2_X1    g16589(.A1(new_n16088_), .A2(new_n16099_), .ZN(new_n16782_));
  NOR3_X1    g16590(.A1(new_n16389_), .A2(new_n16306_), .A3(new_n16782_), .ZN(new_n16783_));
  INV_X1     g16591(.I(new_n16783_), .ZN(new_n16784_));
  NOR3_X1    g16592(.A1(new_n16782_), .A2(new_n16306_), .A3(new_n16098_), .ZN(new_n16785_));
  AOI22_X1   g16593(.A1(new_n16784_), .A2(new_n16098_), .B1(\asqrt[13] ), .B2(new_n16785_), .ZN(new_n16786_));
  INV_X1     g16594(.I(new_n16786_), .ZN(new_n16787_));
  NOR3_X1    g16595(.A1(new_n16744_), .A2(new_n16736_), .A3(\asqrt[52] ), .ZN(new_n16788_));
  OAI21_X1   g16596(.A1(new_n16751_), .A2(new_n16788_), .B(new_n16745_), .ZN(new_n16789_));
  AOI21_X1   g16597(.A1(new_n16789_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n16790_));
  AOI21_X1   g16598(.A1(new_n16790_), .A2(new_n16762_), .B(new_n16770_), .ZN(new_n16791_));
  OAI21_X1   g16599(.A1(new_n16791_), .A2(new_n16763_), .B(\asqrt[55] ), .ZN(new_n16792_));
  NAND2_X1   g16600(.A1(new_n16792_), .A2(new_n703_), .ZN(new_n16793_));
  OAI21_X1   g16601(.A1(new_n16793_), .A2(new_n16780_), .B(new_n16787_), .ZN(new_n16794_));
  AOI21_X1   g16602(.A1(new_n16794_), .A2(new_n16781_), .B(new_n531_), .ZN(new_n16795_));
  INV_X1     g16603(.I(new_n16795_), .ZN(new_n16796_));
  INV_X1     g16604(.I(new_n16794_), .ZN(new_n16797_));
  INV_X1     g16605(.I(new_n16105_), .ZN(new_n16798_));
  NOR3_X1    g16606(.A1(new_n16101_), .A2(new_n16315_), .A3(new_n16798_), .ZN(new_n16799_));
  NOR3_X1    g16607(.A1(new_n16389_), .A2(new_n16101_), .A3(new_n16315_), .ZN(new_n16800_));
  INV_X1     g16608(.I(new_n16800_), .ZN(new_n16801_));
  AOI22_X1   g16609(.A1(new_n16801_), .A2(new_n16798_), .B1(\asqrt[13] ), .B2(new_n16799_), .ZN(new_n16802_));
  INV_X1     g16610(.I(new_n16802_), .ZN(new_n16803_));
  NAND2_X1   g16611(.A1(new_n16781_), .A2(new_n531_), .ZN(new_n16804_));
  OAI21_X1   g16612(.A1(new_n16804_), .A2(new_n16797_), .B(new_n16803_), .ZN(new_n16805_));
  AOI21_X1   g16613(.A1(new_n16805_), .A2(new_n16796_), .B(new_n436_), .ZN(new_n16806_));
  NOR3_X1    g16614(.A1(new_n16389_), .A2(new_n16110_), .A3(new_n16117_), .ZN(new_n16807_));
  INV_X1     g16615(.I(new_n16807_), .ZN(new_n16808_));
  NOR3_X1    g16616(.A1(new_n16110_), .A2(new_n16179_), .A3(new_n16117_), .ZN(new_n16809_));
  AOI22_X1   g16617(.A1(new_n16808_), .A2(new_n16179_), .B1(\asqrt[13] ), .B2(new_n16809_), .ZN(new_n16810_));
  NOR2_X1    g16618(.A1(new_n16795_), .A2(\asqrt[58] ), .ZN(new_n16811_));
  AOI21_X1   g16619(.A1(new_n16811_), .A2(new_n16805_), .B(new_n16810_), .ZN(new_n16812_));
  OAI21_X1   g16620(.A1(new_n16812_), .A2(new_n16806_), .B(\asqrt[59] ), .ZN(new_n16813_));
  NOR2_X1    g16621(.A1(new_n16118_), .A2(new_n16130_), .ZN(new_n16814_));
  NOR3_X1    g16622(.A1(new_n16814_), .A2(new_n16314_), .A3(new_n16129_), .ZN(new_n16815_));
  NOR3_X1    g16623(.A1(new_n16389_), .A2(new_n16314_), .A3(new_n16814_), .ZN(new_n16816_));
  INV_X1     g16624(.I(new_n16816_), .ZN(new_n16817_));
  AOI22_X1   g16625(.A1(new_n16817_), .A2(new_n16129_), .B1(\asqrt[13] ), .B2(new_n16815_), .ZN(new_n16818_));
  INV_X1     g16626(.I(new_n16818_), .ZN(new_n16819_));
  NOR3_X1    g16627(.A1(new_n16791_), .A2(\asqrt[55] ), .A3(new_n16763_), .ZN(new_n16820_));
  OAI21_X1   g16628(.A1(new_n16778_), .A2(new_n16820_), .B(new_n16792_), .ZN(new_n16821_));
  AOI21_X1   g16629(.A1(new_n16821_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n16822_));
  AOI21_X1   g16630(.A1(new_n16822_), .A2(new_n16794_), .B(new_n16802_), .ZN(new_n16823_));
  OAI21_X1   g16631(.A1(new_n16823_), .A2(new_n16795_), .B(\asqrt[58] ), .ZN(new_n16824_));
  NAND2_X1   g16632(.A1(new_n16824_), .A2(new_n327_), .ZN(new_n16825_));
  OAI21_X1   g16633(.A1(new_n16825_), .A2(new_n16812_), .B(new_n16819_), .ZN(new_n16826_));
  AOI21_X1   g16634(.A1(new_n16826_), .A2(new_n16813_), .B(new_n306_), .ZN(new_n16827_));
  INV_X1     g16635(.I(new_n16827_), .ZN(new_n16828_));
  INV_X1     g16636(.I(new_n16826_), .ZN(new_n16829_));
  INV_X1     g16637(.I(new_n16136_), .ZN(new_n16830_));
  NOR3_X1    g16638(.A1(new_n16389_), .A2(new_n16132_), .A3(new_n16322_), .ZN(new_n16831_));
  INV_X1     g16639(.I(new_n16831_), .ZN(new_n16832_));
  NOR3_X1    g16640(.A1(new_n16132_), .A2(new_n16322_), .A3(new_n16830_), .ZN(new_n16833_));
  AOI22_X1   g16641(.A1(new_n16832_), .A2(new_n16830_), .B1(\asqrt[13] ), .B2(new_n16833_), .ZN(new_n16834_));
  INV_X1     g16642(.I(new_n16834_), .ZN(new_n16835_));
  NAND2_X1   g16643(.A1(new_n16813_), .A2(new_n306_), .ZN(new_n16836_));
  OAI21_X1   g16644(.A1(new_n16829_), .A2(new_n16836_), .B(new_n16835_), .ZN(new_n16837_));
  AOI21_X1   g16645(.A1(new_n16837_), .A2(new_n16828_), .B(new_n218_), .ZN(new_n16838_));
  NOR3_X1    g16646(.A1(new_n16141_), .A2(new_n16178_), .A3(new_n16147_), .ZN(new_n16839_));
  NOR3_X1    g16647(.A1(new_n16389_), .A2(new_n16141_), .A3(new_n16147_), .ZN(new_n16840_));
  INV_X1     g16648(.I(new_n16840_), .ZN(new_n16841_));
  AOI22_X1   g16649(.A1(new_n16841_), .A2(new_n16178_), .B1(\asqrt[13] ), .B2(new_n16839_), .ZN(new_n16842_));
  NOR2_X1    g16650(.A1(new_n16827_), .A2(\asqrt[61] ), .ZN(new_n16843_));
  AOI21_X1   g16651(.A1(new_n16843_), .A2(new_n16837_), .B(new_n16842_), .ZN(new_n16844_));
  OAI21_X1   g16652(.A1(new_n16844_), .A2(new_n16838_), .B(\asqrt[62] ), .ZN(new_n16845_));
  NOR2_X1    g16653(.A1(new_n16148_), .A2(new_n16155_), .ZN(new_n16846_));
  NOR3_X1    g16654(.A1(new_n16389_), .A2(new_n16344_), .A3(new_n16846_), .ZN(new_n16847_));
  INV_X1     g16655(.I(new_n16847_), .ZN(new_n16848_));
  NOR3_X1    g16656(.A1(new_n16846_), .A2(new_n16344_), .A3(new_n16154_), .ZN(new_n16849_));
  AOI22_X1   g16657(.A1(new_n16848_), .A2(new_n16154_), .B1(\asqrt[13] ), .B2(new_n16849_), .ZN(new_n16850_));
  INV_X1     g16658(.I(new_n16850_), .ZN(new_n16851_));
  NOR3_X1    g16659(.A1(new_n16823_), .A2(\asqrt[58] ), .A3(new_n16795_), .ZN(new_n16852_));
  OAI21_X1   g16660(.A1(new_n16810_), .A2(new_n16852_), .B(new_n16824_), .ZN(new_n16853_));
  AOI21_X1   g16661(.A1(new_n16853_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n16854_));
  AOI21_X1   g16662(.A1(new_n16854_), .A2(new_n16826_), .B(new_n16834_), .ZN(new_n16855_));
  OAI21_X1   g16663(.A1(new_n16855_), .A2(new_n16827_), .B(\asqrt[61] ), .ZN(new_n16856_));
  NAND2_X1   g16664(.A1(new_n16856_), .A2(new_n207_), .ZN(new_n16857_));
  OAI21_X1   g16665(.A1(new_n16857_), .A2(new_n16844_), .B(new_n16851_), .ZN(new_n16858_));
  INV_X1     g16666(.I(new_n16346_), .ZN(new_n16859_));
  NAND4_X1   g16667(.A1(\asqrt[13] ), .A2(new_n16345_), .A3(new_n16161_), .A4(new_n16859_), .ZN(new_n16860_));
  NAND2_X1   g16668(.A1(new_n16859_), .A2(new_n16345_), .ZN(new_n16861_));
  OAI21_X1   g16669(.A1(new_n16389_), .A2(new_n16861_), .B(new_n16326_), .ZN(new_n16862_));
  NAND2_X1   g16670(.A1(new_n16862_), .A2(new_n16860_), .ZN(new_n16863_));
  INV_X1     g16671(.I(new_n16365_), .ZN(new_n16864_));
  AOI21_X1   g16672(.A1(new_n16328_), .A2(new_n16345_), .B(new_n16172_), .ZN(new_n16865_));
  AOI21_X1   g16673(.A1(\asqrt[13] ), .A2(new_n16865_), .B(new_n16864_), .ZN(new_n16866_));
  NAND2_X1   g16674(.A1(new_n16863_), .A2(new_n16866_), .ZN(new_n16867_));
  AOI21_X1   g16675(.A1(new_n16858_), .A2(new_n16845_), .B(new_n16867_), .ZN(new_n16868_));
  NOR2_X1    g16676(.A1(new_n16868_), .A2(\asqrt[63] ), .ZN(new_n16869_));
  INV_X1     g16677(.I(new_n16858_), .ZN(new_n16870_));
  INV_X1     g16678(.I(new_n16863_), .ZN(new_n16871_));
  NAND2_X1   g16679(.A1(new_n16845_), .A2(new_n16871_), .ZN(new_n16872_));
  AOI21_X1   g16680(.A1(\asqrt[13] ), .A2(new_n16173_), .B(new_n16347_), .ZN(new_n16873_));
  OR3_X2     g16681(.A1(new_n16873_), .A2(new_n193_), .A3(new_n16865_), .Z(new_n16874_));
  OAI21_X1   g16682(.A1(new_n15717_), .A2(new_n16334_), .B(new_n16168_), .ZN(new_n16875_));
  NOR4_X1    g16683(.A1(new_n16864_), .A2(new_n16171_), .A3(new_n16332_), .A4(new_n16875_), .ZN(new_n16876_));
  NAND2_X1   g16684(.A1(new_n16876_), .A2(new_n16177_), .ZN(new_n16877_));
  NAND2_X1   g16685(.A1(new_n16874_), .A2(new_n16877_), .ZN(new_n16878_));
  INV_X1     g16686(.I(new_n16878_), .ZN(new_n16879_));
  OAI21_X1   g16687(.A1(new_n16870_), .A2(new_n16872_), .B(new_n16879_), .ZN(new_n16880_));
  NOR2_X1    g16688(.A1(new_n16869_), .A2(new_n16880_), .ZN(new_n16881_));
  INV_X1     g16689(.I(\a[24] ), .ZN(new_n16882_));
  NOR2_X1    g16690(.A1(\a[22] ), .A2(\a[23] ), .ZN(new_n16883_));
  INV_X1     g16691(.I(new_n16883_), .ZN(new_n16884_));
  NOR2_X1    g16692(.A1(new_n16884_), .A2(\a[24] ), .ZN(new_n16885_));
  INV_X1     g16693(.I(new_n16885_), .ZN(new_n16886_));
  OAI21_X1   g16694(.A1(new_n16881_), .A2(new_n16882_), .B(new_n16886_), .ZN(new_n16887_));
  NOR3_X1    g16695(.A1(new_n16332_), .A2(new_n16335_), .A3(new_n16885_), .ZN(new_n16888_));
  NAND3_X1   g16696(.A1(new_n16177_), .A2(new_n16365_), .A3(new_n16888_), .ZN(new_n16889_));
  INV_X1     g16697(.I(new_n16889_), .ZN(new_n16890_));
  OAI21_X1   g16698(.A1(new_n16881_), .A2(new_n16882_), .B(new_n16890_), .ZN(new_n16891_));
  NOR3_X1    g16699(.A1(new_n16855_), .A2(\asqrt[61] ), .A3(new_n16827_), .ZN(new_n16892_));
  OAI21_X1   g16700(.A1(new_n16842_), .A2(new_n16892_), .B(new_n16856_), .ZN(new_n16893_));
  INV_X1     g16701(.I(new_n16842_), .ZN(new_n16894_));
  INV_X1     g16702(.I(new_n16810_), .ZN(new_n16895_));
  INV_X1     g16703(.I(new_n16778_), .ZN(new_n16896_));
  INV_X1     g16704(.I(new_n16751_), .ZN(new_n16897_));
  INV_X1     g16705(.I(new_n16724_), .ZN(new_n16898_));
  INV_X1     g16706(.I(new_n16698_), .ZN(new_n16899_));
  INV_X1     g16707(.I(new_n16672_), .ZN(new_n16900_));
  INV_X1     g16708(.I(new_n16643_), .ZN(new_n16901_));
  NOR3_X1    g16709(.A1(new_n16642_), .A2(new_n16627_), .A3(\asqrt[41] ), .ZN(new_n16902_));
  NOR2_X1    g16710(.A1(new_n16902_), .A2(new_n16648_), .ZN(new_n16903_));
  OAI21_X1   g16711(.A1(new_n16903_), .A2(new_n16901_), .B(\asqrt[42] ), .ZN(new_n16904_));
  NAND2_X1   g16712(.A1(new_n16904_), .A2(new_n3218_), .ZN(new_n16905_));
  OAI21_X1   g16713(.A1(new_n16905_), .A2(new_n16666_), .B(new_n16900_), .ZN(new_n16906_));
  NAND3_X1   g16714(.A1(new_n16906_), .A2(new_n2954_), .A3(new_n16667_), .ZN(new_n16907_));
  AOI22_X1   g16715(.A1(new_n16907_), .A2(new_n16681_), .B1(\asqrt[44] ), .B2(new_n16690_), .ZN(new_n16908_));
  OAI21_X1   g16716(.A1(new_n16908_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n16909_));
  OAI21_X1   g16717(.A1(new_n16909_), .A2(new_n16692_), .B(new_n16899_), .ZN(new_n16910_));
  NAND3_X1   g16718(.A1(new_n16910_), .A2(new_n2229_), .A3(new_n16693_), .ZN(new_n16911_));
  AOI22_X1   g16719(.A1(new_n16911_), .A2(new_n16707_), .B1(\asqrt[47] ), .B2(new_n16716_), .ZN(new_n16912_));
  OAI21_X1   g16720(.A1(new_n16912_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n16913_));
  OAI21_X1   g16721(.A1(new_n16913_), .A2(new_n16718_), .B(new_n16898_), .ZN(new_n16914_));
  NAND3_X1   g16722(.A1(new_n16914_), .A2(new_n1612_), .A3(new_n16719_), .ZN(new_n16915_));
  AOI22_X1   g16723(.A1(new_n16915_), .A2(new_n16733_), .B1(\asqrt[50] ), .B2(new_n16742_), .ZN(new_n16916_));
  OAI21_X1   g16724(.A1(new_n16916_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n16917_));
  OAI21_X1   g16725(.A1(new_n16917_), .A2(new_n16744_), .B(new_n16897_), .ZN(new_n16918_));
  NAND3_X1   g16726(.A1(new_n16918_), .A2(new_n1103_), .A3(new_n16745_), .ZN(new_n16919_));
  AOI22_X1   g16727(.A1(new_n16919_), .A2(new_n16760_), .B1(\asqrt[53] ), .B2(new_n16789_), .ZN(new_n16920_));
  OAI21_X1   g16728(.A1(new_n16920_), .A2(new_n904_), .B(new_n823_), .ZN(new_n16921_));
  OAI21_X1   g16729(.A1(new_n16921_), .A2(new_n16791_), .B(new_n16896_), .ZN(new_n16922_));
  NAND3_X1   g16730(.A1(new_n16922_), .A2(new_n703_), .A3(new_n16792_), .ZN(new_n16923_));
  AOI22_X1   g16731(.A1(new_n16923_), .A2(new_n16787_), .B1(\asqrt[56] ), .B2(new_n16821_), .ZN(new_n16924_));
  OAI21_X1   g16732(.A1(new_n16924_), .A2(new_n531_), .B(new_n436_), .ZN(new_n16925_));
  OAI21_X1   g16733(.A1(new_n16925_), .A2(new_n16823_), .B(new_n16895_), .ZN(new_n16926_));
  NAND3_X1   g16734(.A1(new_n16926_), .A2(new_n327_), .A3(new_n16824_), .ZN(new_n16927_));
  AOI22_X1   g16735(.A1(new_n16927_), .A2(new_n16819_), .B1(new_n16853_), .B2(\asqrt[59] ), .ZN(new_n16928_));
  OAI21_X1   g16736(.A1(new_n16928_), .A2(new_n306_), .B(new_n218_), .ZN(new_n16929_));
  OAI21_X1   g16737(.A1(new_n16929_), .A2(new_n16855_), .B(new_n16894_), .ZN(new_n16930_));
  NAND3_X1   g16738(.A1(new_n16930_), .A2(new_n207_), .A3(new_n16856_), .ZN(new_n16931_));
  AOI22_X1   g16739(.A1(new_n16931_), .A2(new_n16851_), .B1(new_n16893_), .B2(\asqrt[62] ), .ZN(new_n16932_));
  OAI21_X1   g16740(.A1(new_n16932_), .A2(new_n16867_), .B(new_n193_), .ZN(new_n16933_));
  AOI21_X1   g16741(.A1(new_n16893_), .A2(\asqrt[62] ), .B(new_n16863_), .ZN(new_n16934_));
  AOI21_X1   g16742(.A1(new_n16934_), .A2(new_n16858_), .B(new_n16878_), .ZN(new_n16935_));
  AOI21_X1   g16743(.A1(new_n16933_), .A2(new_n16935_), .B(new_n16341_), .ZN(new_n16936_));
  OAI21_X1   g16744(.A1(new_n16869_), .A2(new_n16880_), .B(new_n16882_), .ZN(new_n16937_));
  AOI21_X1   g16745(.A1(\a[25] ), .A2(new_n16937_), .B(new_n16936_), .ZN(new_n16938_));
  AOI22_X1   g16746(.A1(new_n16938_), .A2(new_n16891_), .B1(\asqrt[13] ), .B2(new_n16887_), .ZN(new_n16939_));
  NOR2_X1    g16747(.A1(new_n16939_), .A2(new_n15770_), .ZN(new_n16940_));
  NAND2_X1   g16748(.A1(new_n16938_), .A2(new_n16891_), .ZN(new_n16941_));
  OAI21_X1   g16749(.A1(new_n16869_), .A2(new_n16880_), .B(new_n16340_), .ZN(new_n16942_));
  NAND2_X1   g16750(.A1(new_n16934_), .A2(new_n16858_), .ZN(new_n16943_));
  OAI21_X1   g16751(.A1(new_n16876_), .A2(new_n16338_), .B(new_n16177_), .ZN(new_n16944_));
  NAND4_X1   g16752(.A1(new_n16933_), .A2(new_n16943_), .A3(new_n16874_), .A4(new_n16944_), .ZN(new_n16945_));
  AOI21_X1   g16753(.A1(new_n16945_), .A2(new_n16942_), .B(new_n16353_), .ZN(new_n16946_));
  INV_X1     g16754(.I(new_n16943_), .ZN(new_n16947_));
  NAND2_X1   g16755(.A1(new_n16874_), .A2(new_n16944_), .ZN(new_n16948_));
  NOR3_X1    g16756(.A1(new_n16947_), .A2(new_n16869_), .A3(new_n16948_), .ZN(new_n16949_));
  NOR3_X1    g16757(.A1(new_n16949_), .A2(new_n16936_), .A3(\a[26] ), .ZN(new_n16950_));
  NOR2_X1    g16758(.A1(new_n16946_), .A2(new_n16950_), .ZN(new_n16951_));
  AOI21_X1   g16759(.A1(new_n16887_), .A2(\asqrt[13] ), .B(\asqrt[14] ), .ZN(new_n16952_));
  AOI21_X1   g16760(.A1(new_n16941_), .A2(new_n16952_), .B(new_n16951_), .ZN(new_n16953_));
  OAI21_X1   g16761(.A1(new_n16953_), .A2(new_n16940_), .B(\asqrt[15] ), .ZN(new_n16954_));
  OAI21_X1   g16762(.A1(\asqrt[63] ), .A2(new_n16868_), .B(new_n16935_), .ZN(\asqrt[12] ));
  NOR3_X1    g16763(.A1(new_n16433_), .A2(new_n16352_), .A3(new_n16358_), .ZN(new_n16956_));
  NAND3_X1   g16764(.A1(\asqrt[12] ), .A2(new_n16371_), .A3(new_n16418_), .ZN(new_n16957_));
  AOI22_X1   g16765(.A1(new_n16957_), .A2(new_n16433_), .B1(\asqrt[12] ), .B2(new_n16956_), .ZN(new_n16958_));
  INV_X1     g16766(.I(new_n16958_), .ZN(new_n16959_));
  OAI21_X1   g16767(.A1(new_n16939_), .A2(new_n15770_), .B(new_n15067_), .ZN(new_n16960_));
  OAI21_X1   g16768(.A1(new_n16960_), .A2(new_n16953_), .B(new_n16959_), .ZN(new_n16961_));
  AOI21_X1   g16769(.A1(new_n16961_), .A2(new_n16954_), .B(new_n14601_), .ZN(new_n16962_));
  NOR2_X1    g16770(.A1(new_n16370_), .A2(new_n16368_), .ZN(new_n16963_));
  NOR2_X1    g16771(.A1(new_n16362_), .A2(new_n16372_), .ZN(new_n16964_));
  INV_X1     g16772(.I(new_n16964_), .ZN(new_n16965_));
  NAND4_X1   g16773(.A1(\asqrt[12] ), .A2(new_n16363_), .A3(new_n16963_), .A4(new_n16965_), .ZN(new_n16966_));
  NOR3_X1    g16774(.A1(new_n16881_), .A2(new_n16422_), .A3(new_n16964_), .ZN(new_n16967_));
  OAI21_X1   g16775(.A1(new_n16967_), .A2(new_n16963_), .B(new_n16966_), .ZN(new_n16968_));
  INV_X1     g16776(.I(new_n16968_), .ZN(new_n16969_));
  AOI21_X1   g16777(.A1(new_n16933_), .A2(new_n16935_), .B(new_n16882_), .ZN(new_n16970_));
  OAI21_X1   g16778(.A1(new_n16970_), .A2(new_n16885_), .B(\asqrt[13] ), .ZN(new_n16971_));
  INV_X1     g16779(.I(new_n16971_), .ZN(new_n16972_));
  NOR2_X1    g16780(.A1(new_n16970_), .A2(new_n16889_), .ZN(new_n16973_));
  INV_X1     g16781(.I(\a[25] ), .ZN(new_n16974_));
  AOI21_X1   g16782(.A1(\asqrt[12] ), .A2(new_n16882_), .B(new_n16974_), .ZN(new_n16975_));
  NOR3_X1    g16783(.A1(new_n16973_), .A2(new_n16975_), .A3(new_n16936_), .ZN(new_n16976_));
  OAI21_X1   g16784(.A1(new_n16976_), .A2(new_n16972_), .B(\asqrt[14] ), .ZN(new_n16977_));
  AOI21_X1   g16785(.A1(\asqrt[12] ), .A2(\a[24] ), .B(new_n16885_), .ZN(new_n16978_));
  OAI21_X1   g16786(.A1(new_n16978_), .A2(new_n16389_), .B(new_n15770_), .ZN(new_n16979_));
  OAI22_X1   g16787(.A1(new_n16976_), .A2(new_n16979_), .B1(new_n16946_), .B2(new_n16950_), .ZN(new_n16980_));
  AOI21_X1   g16788(.A1(new_n16980_), .A2(new_n16977_), .B(new_n15067_), .ZN(new_n16981_));
  AOI21_X1   g16789(.A1(new_n16933_), .A2(new_n16935_), .B(\a[24] ), .ZN(new_n16982_));
  OAI21_X1   g16790(.A1(new_n16974_), .A2(new_n16982_), .B(new_n16942_), .ZN(new_n16983_));
  OAI21_X1   g16791(.A1(new_n16983_), .A2(new_n16973_), .B(new_n16971_), .ZN(new_n16984_));
  AOI21_X1   g16792(.A1(new_n16984_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n16985_));
  AOI21_X1   g16793(.A1(new_n16985_), .A2(new_n16980_), .B(new_n16958_), .ZN(new_n16986_));
  NOR3_X1    g16794(.A1(new_n16986_), .A2(new_n16981_), .A3(\asqrt[16] ), .ZN(new_n16987_));
  NOR2_X1    g16795(.A1(new_n16987_), .A2(new_n16969_), .ZN(new_n16988_));
  OAI21_X1   g16796(.A1(new_n16988_), .A2(new_n16962_), .B(\asqrt[17] ), .ZN(new_n16989_));
  NOR2_X1    g16797(.A1(new_n16435_), .A2(new_n16427_), .ZN(new_n16990_));
  NOR3_X1    g16798(.A1(new_n16881_), .A2(new_n16374_), .A3(new_n16990_), .ZN(new_n16991_));
  INV_X1     g16799(.I(new_n16991_), .ZN(new_n16992_));
  NOR3_X1    g16800(.A1(new_n16990_), .A2(new_n16374_), .A3(new_n16432_), .ZN(new_n16993_));
  AOI22_X1   g16801(.A1(new_n16992_), .A2(new_n16432_), .B1(\asqrt[12] ), .B2(new_n16993_), .ZN(new_n16994_));
  INV_X1     g16802(.I(new_n16994_), .ZN(new_n16995_));
  OAI21_X1   g16803(.A1(new_n16986_), .A2(new_n16981_), .B(\asqrt[16] ), .ZN(new_n16996_));
  NAND2_X1   g16804(.A1(new_n16996_), .A2(new_n14017_), .ZN(new_n16997_));
  OAI21_X1   g16805(.A1(new_n16988_), .A2(new_n16997_), .B(new_n16995_), .ZN(new_n16998_));
  AOI21_X1   g16806(.A1(new_n16998_), .A2(new_n16989_), .B(new_n13353_), .ZN(new_n16999_));
  NOR3_X1    g16807(.A1(new_n16384_), .A2(new_n16393_), .A3(new_n16391_), .ZN(new_n17000_));
  NOR3_X1    g16808(.A1(new_n16881_), .A2(new_n16384_), .A3(new_n16393_), .ZN(new_n17001_));
  INV_X1     g16809(.I(new_n17001_), .ZN(new_n17002_));
  AOI22_X1   g16810(.A1(new_n17002_), .A2(new_n16391_), .B1(\asqrt[12] ), .B2(new_n17000_), .ZN(new_n17003_));
  OAI21_X1   g16811(.A1(new_n16969_), .A2(new_n16987_), .B(new_n16996_), .ZN(new_n17004_));
  AOI21_X1   g16812(.A1(new_n17004_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n17005_));
  AOI21_X1   g16813(.A1(new_n17005_), .A2(new_n16998_), .B(new_n17003_), .ZN(new_n17006_));
  OAI21_X1   g16814(.A1(new_n17006_), .A2(new_n16999_), .B(\asqrt[19] ), .ZN(new_n17007_));
  INV_X1     g16815(.I(new_n17007_), .ZN(new_n17008_));
  NAND2_X1   g16816(.A1(new_n16438_), .A2(new_n16430_), .ZN(new_n17009_));
  NAND3_X1   g16817(.A1(\asqrt[12] ), .A2(new_n16395_), .A3(new_n17009_), .ZN(new_n17010_));
  AND3_X2    g16818(.A1(new_n16395_), .A2(new_n16400_), .A3(new_n17009_), .Z(new_n17011_));
  AOI22_X1   g16819(.A1(new_n17010_), .A2(new_n16401_), .B1(\asqrt[12] ), .B2(new_n17011_), .ZN(new_n17012_));
  NOR3_X1    g16820(.A1(new_n17006_), .A2(new_n16999_), .A3(\asqrt[19] ), .ZN(new_n17013_));
  NOR2_X1    g16821(.A1(new_n17013_), .A2(new_n17012_), .ZN(new_n17014_));
  OAI21_X1   g16822(.A1(new_n17014_), .A2(new_n17008_), .B(\asqrt[20] ), .ZN(new_n17015_));
  INV_X1     g16823(.I(new_n16408_), .ZN(new_n17016_));
  NOR3_X1    g16824(.A1(new_n16404_), .A2(new_n16449_), .A3(new_n17016_), .ZN(new_n17017_));
  NOR3_X1    g16825(.A1(new_n16881_), .A2(new_n16404_), .A3(new_n16449_), .ZN(new_n17018_));
  INV_X1     g16826(.I(new_n17018_), .ZN(new_n17019_));
  AOI22_X1   g16827(.A1(new_n17019_), .A2(new_n17016_), .B1(\asqrt[12] ), .B2(new_n17017_), .ZN(new_n17020_));
  INV_X1     g16828(.I(new_n17020_), .ZN(new_n17021_));
  NAND2_X1   g16829(.A1(new_n17007_), .A2(new_n12364_), .ZN(new_n17022_));
  OAI21_X1   g16830(.A1(new_n17014_), .A2(new_n17022_), .B(new_n17021_), .ZN(new_n17023_));
  AOI21_X1   g16831(.A1(new_n17023_), .A2(new_n17015_), .B(new_n11736_), .ZN(new_n17024_));
  INV_X1     g16832(.I(new_n16474_), .ZN(new_n17025_));
  NAND3_X1   g16833(.A1(\asqrt[12] ), .A2(new_n16412_), .A3(new_n17025_), .ZN(new_n17026_));
  AND3_X2    g16834(.A1(new_n17025_), .A2(new_n16412_), .A3(new_n16416_), .Z(new_n17027_));
  AOI22_X1   g16835(.A1(new_n17026_), .A2(new_n16417_), .B1(\asqrt[12] ), .B2(new_n17027_), .ZN(new_n17028_));
  OAI21_X1   g16836(.A1(new_n17012_), .A2(new_n17013_), .B(new_n17007_), .ZN(new_n17029_));
  AOI21_X1   g16837(.A1(new_n17029_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n17030_));
  AOI21_X1   g16838(.A1(new_n17030_), .A2(new_n17023_), .B(new_n17028_), .ZN(new_n17031_));
  OAI21_X1   g16839(.A1(new_n17031_), .A2(new_n17024_), .B(\asqrt[22] ), .ZN(new_n17032_));
  INV_X1     g16840(.I(new_n17032_), .ZN(new_n17033_));
  INV_X1     g16841(.I(new_n16477_), .ZN(new_n17034_));
  NOR3_X1    g16842(.A1(new_n17034_), .A2(new_n16443_), .A3(new_n16476_), .ZN(new_n17035_));
  NOR3_X1    g16843(.A1(new_n16881_), .A2(new_n16443_), .A3(new_n17034_), .ZN(new_n17036_));
  INV_X1     g16844(.I(new_n17036_), .ZN(new_n17037_));
  AOI22_X1   g16845(.A1(new_n17037_), .A2(new_n16476_), .B1(\asqrt[12] ), .B2(new_n17035_), .ZN(new_n17038_));
  NOR3_X1    g16846(.A1(new_n17031_), .A2(new_n17024_), .A3(\asqrt[22] ), .ZN(new_n17039_));
  NOR2_X1    g16847(.A1(new_n17039_), .A2(new_n17038_), .ZN(new_n17040_));
  OAI21_X1   g16848(.A1(new_n17040_), .A2(new_n17033_), .B(\asqrt[23] ), .ZN(new_n17041_));
  INV_X1     g16849(.I(new_n16458_), .ZN(new_n17042_));
  NOR3_X1    g16850(.A1(new_n16881_), .A2(new_n16454_), .A3(new_n16459_), .ZN(new_n17043_));
  INV_X1     g16851(.I(new_n17043_), .ZN(new_n17044_));
  NOR3_X1    g16852(.A1(new_n16454_), .A2(new_n17042_), .A3(new_n16459_), .ZN(new_n17045_));
  AOI22_X1   g16853(.A1(new_n17044_), .A2(new_n17042_), .B1(\asqrt[12] ), .B2(new_n17045_), .ZN(new_n17046_));
  INV_X1     g16854(.I(new_n17046_), .ZN(new_n17047_));
  NAND2_X1   g16855(.A1(new_n17032_), .A2(new_n10812_), .ZN(new_n17048_));
  OAI21_X1   g16856(.A1(new_n17040_), .A2(new_n17048_), .B(new_n17047_), .ZN(new_n17049_));
  AOI21_X1   g16857(.A1(new_n17049_), .A2(new_n17041_), .B(new_n10221_), .ZN(new_n17050_));
  OAI21_X1   g16858(.A1(new_n16460_), .A2(new_n16466_), .B(new_n16464_), .ZN(new_n17051_));
  AOI21_X1   g16859(.A1(\asqrt[23] ), .A2(new_n16479_), .B(new_n17051_), .ZN(new_n17052_));
  OAI21_X1   g16860(.A1(new_n16460_), .A2(new_n16466_), .B(new_n16461_), .ZN(new_n17053_));
  NOR2_X1    g16861(.A1(new_n16881_), .A2(new_n17053_), .ZN(new_n17054_));
  INV_X1     g16862(.I(new_n17054_), .ZN(new_n17055_));
  AOI22_X1   g16863(.A1(new_n17055_), .A2(new_n16465_), .B1(\asqrt[12] ), .B2(new_n17052_), .ZN(new_n17056_));
  OAI21_X1   g16864(.A1(new_n17038_), .A2(new_n17039_), .B(new_n17032_), .ZN(new_n17057_));
  AOI21_X1   g16865(.A1(new_n17057_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n17058_));
  AOI21_X1   g16866(.A1(new_n17058_), .A2(new_n17049_), .B(new_n17056_), .ZN(new_n17059_));
  OAI21_X1   g16867(.A1(new_n17059_), .A2(new_n17050_), .B(\asqrt[25] ), .ZN(new_n17060_));
  INV_X1     g16868(.I(new_n17060_), .ZN(new_n17061_));
  INV_X1     g16869(.I(new_n16473_), .ZN(new_n17062_));
  INV_X1     g16870(.I(new_n16467_), .ZN(new_n17063_));
  INV_X1     g16871(.I(new_n16480_), .ZN(new_n17064_));
  NOR2_X1    g16872(.A1(new_n17064_), .A2(new_n17063_), .ZN(new_n17065_));
  NOR3_X1    g16873(.A1(new_n16881_), .A2(new_n16468_), .A3(new_n17065_), .ZN(new_n17066_));
  INV_X1     g16874(.I(new_n17066_), .ZN(new_n17067_));
  NOR3_X1    g16875(.A1(new_n17065_), .A2(new_n16468_), .A3(new_n17062_), .ZN(new_n17068_));
  AOI22_X1   g16876(.A1(new_n17067_), .A2(new_n17062_), .B1(\asqrt[12] ), .B2(new_n17068_), .ZN(new_n17069_));
  NOR3_X1    g16877(.A1(new_n17059_), .A2(new_n17050_), .A3(\asqrt[25] ), .ZN(new_n17070_));
  NOR2_X1    g16878(.A1(new_n17070_), .A2(new_n17069_), .ZN(new_n17071_));
  OAI21_X1   g16879(.A1(new_n17071_), .A2(new_n17061_), .B(\asqrt[26] ), .ZN(new_n17072_));
  INV_X1     g16880(.I(new_n16487_), .ZN(new_n17073_));
  NOR3_X1    g16881(.A1(new_n16483_), .A2(new_n17073_), .A3(new_n16488_), .ZN(new_n17074_));
  NOR3_X1    g16882(.A1(new_n16881_), .A2(new_n16483_), .A3(new_n16488_), .ZN(new_n17075_));
  INV_X1     g16883(.I(new_n17075_), .ZN(new_n17076_));
  AOI22_X1   g16884(.A1(new_n17076_), .A2(new_n17073_), .B1(\asqrt[12] ), .B2(new_n17074_), .ZN(new_n17077_));
  INV_X1     g16885(.I(new_n17077_), .ZN(new_n17078_));
  NAND2_X1   g16886(.A1(new_n17060_), .A2(new_n9317_), .ZN(new_n17079_));
  OAI21_X1   g16887(.A1(new_n17071_), .A2(new_n17079_), .B(new_n17078_), .ZN(new_n17080_));
  AOI21_X1   g16888(.A1(new_n17080_), .A2(new_n17072_), .B(new_n8826_), .ZN(new_n17081_));
  NOR2_X1    g16889(.A1(new_n16489_), .A2(new_n16497_), .ZN(new_n17082_));
  INV_X1     g16890(.I(new_n17082_), .ZN(new_n17083_));
  NAND3_X1   g16891(.A1(\asqrt[12] ), .A2(new_n16490_), .A3(new_n17083_), .ZN(new_n17084_));
  AND3_X2    g16892(.A1(new_n17083_), .A2(new_n16490_), .A3(new_n16495_), .Z(new_n17085_));
  AOI22_X1   g16893(.A1(new_n17084_), .A2(new_n16496_), .B1(\asqrt[12] ), .B2(new_n17085_), .ZN(new_n17086_));
  OAI21_X1   g16894(.A1(new_n17069_), .A2(new_n17070_), .B(new_n17060_), .ZN(new_n17087_));
  AOI21_X1   g16895(.A1(new_n17087_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n17088_));
  AOI21_X1   g16896(.A1(new_n17088_), .A2(new_n17080_), .B(new_n17086_), .ZN(new_n17089_));
  OAI21_X1   g16897(.A1(new_n17089_), .A2(new_n17081_), .B(\asqrt[28] ), .ZN(new_n17090_));
  INV_X1     g16898(.I(new_n17090_), .ZN(new_n17091_));
  INV_X1     g16899(.I(new_n16504_), .ZN(new_n17092_));
  INV_X1     g16900(.I(new_n16498_), .ZN(new_n17093_));
  INV_X1     g16901(.I(new_n16506_), .ZN(new_n17094_));
  NOR2_X1    g16902(.A1(new_n17094_), .A2(new_n17093_), .ZN(new_n17095_));
  NOR3_X1    g16903(.A1(new_n17095_), .A2(new_n16499_), .A3(new_n17092_), .ZN(new_n17096_));
  NOR3_X1    g16904(.A1(new_n16881_), .A2(new_n16499_), .A3(new_n17095_), .ZN(new_n17097_));
  INV_X1     g16905(.I(new_n17097_), .ZN(new_n17098_));
  AOI22_X1   g16906(.A1(new_n17098_), .A2(new_n17092_), .B1(\asqrt[12] ), .B2(new_n17096_), .ZN(new_n17099_));
  NOR3_X1    g16907(.A1(new_n17089_), .A2(new_n17081_), .A3(\asqrt[28] ), .ZN(new_n17100_));
  NOR2_X1    g16908(.A1(new_n17100_), .A2(new_n17099_), .ZN(new_n17101_));
  OAI21_X1   g16909(.A1(new_n17101_), .A2(new_n17091_), .B(\asqrt[29] ), .ZN(new_n17102_));
  INV_X1     g16910(.I(new_n16514_), .ZN(new_n17103_));
  NOR3_X1    g16911(.A1(new_n16881_), .A2(new_n16509_), .A3(new_n16551_), .ZN(new_n17104_));
  INV_X1     g16912(.I(new_n17104_), .ZN(new_n17105_));
  NOR3_X1    g16913(.A1(new_n16509_), .A2(new_n17103_), .A3(new_n16551_), .ZN(new_n17106_));
  AOI22_X1   g16914(.A1(new_n17105_), .A2(new_n17103_), .B1(\asqrt[12] ), .B2(new_n17106_), .ZN(new_n17107_));
  INV_X1     g16915(.I(new_n17107_), .ZN(new_n17108_));
  NAND2_X1   g16916(.A1(new_n17090_), .A2(new_n8036_), .ZN(new_n17109_));
  OAI21_X1   g16917(.A1(new_n17101_), .A2(new_n17109_), .B(new_n17108_), .ZN(new_n17110_));
  AOI21_X1   g16918(.A1(new_n17110_), .A2(new_n17102_), .B(new_n7539_), .ZN(new_n17111_));
  NOR2_X1    g16919(.A1(new_n16524_), .A2(new_n16516_), .ZN(new_n17112_));
  INV_X1     g16920(.I(new_n17112_), .ZN(new_n17113_));
  AND3_X2    g16921(.A1(new_n17113_), .A2(new_n16517_), .A3(new_n16522_), .Z(new_n17114_));
  NAND3_X1   g16922(.A1(\asqrt[12] ), .A2(new_n16517_), .A3(new_n17113_), .ZN(new_n17115_));
  AOI22_X1   g16923(.A1(new_n17115_), .A2(new_n16523_), .B1(\asqrt[12] ), .B2(new_n17114_), .ZN(new_n17116_));
  OAI21_X1   g16924(.A1(new_n17099_), .A2(new_n17100_), .B(new_n17090_), .ZN(new_n17117_));
  AOI21_X1   g16925(.A1(new_n17117_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n17118_));
  AOI21_X1   g16926(.A1(new_n17118_), .A2(new_n17110_), .B(new_n17116_), .ZN(new_n17119_));
  OAI21_X1   g16927(.A1(new_n17119_), .A2(new_n17111_), .B(\asqrt[31] ), .ZN(new_n17120_));
  INV_X1     g16928(.I(new_n17120_), .ZN(new_n17121_));
  NOR2_X1    g16929(.A1(new_n16535_), .A2(new_n16528_), .ZN(new_n17122_));
  NOR3_X1    g16930(.A1(new_n16881_), .A2(new_n16526_), .A3(new_n17122_), .ZN(new_n17123_));
  INV_X1     g16931(.I(new_n17123_), .ZN(new_n17124_));
  NOR3_X1    g16932(.A1(new_n17122_), .A2(new_n16526_), .A3(new_n16534_), .ZN(new_n17125_));
  AOI22_X1   g16933(.A1(new_n17124_), .A2(new_n16534_), .B1(\asqrt[12] ), .B2(new_n17125_), .ZN(new_n17126_));
  NOR3_X1    g16934(.A1(new_n17119_), .A2(new_n17111_), .A3(\asqrt[31] ), .ZN(new_n17127_));
  NOR2_X1    g16935(.A1(new_n17127_), .A2(new_n17126_), .ZN(new_n17128_));
  OAI21_X1   g16936(.A1(new_n17128_), .A2(new_n17121_), .B(\asqrt[32] ), .ZN(new_n17129_));
  INV_X1     g16937(.I(new_n16541_), .ZN(new_n17130_));
  NOR3_X1    g16938(.A1(new_n16537_), .A2(new_n17130_), .A3(new_n16583_), .ZN(new_n17131_));
  NOR3_X1    g16939(.A1(new_n16881_), .A2(new_n16537_), .A3(new_n16583_), .ZN(new_n17132_));
  INV_X1     g16940(.I(new_n17132_), .ZN(new_n17133_));
  AOI22_X1   g16941(.A1(new_n17133_), .A2(new_n17130_), .B1(\asqrt[12] ), .B2(new_n17131_), .ZN(new_n17134_));
  INV_X1     g16942(.I(new_n17134_), .ZN(new_n17135_));
  NAND2_X1   g16943(.A1(new_n17120_), .A2(new_n6824_), .ZN(new_n17136_));
  OAI21_X1   g16944(.A1(new_n17128_), .A2(new_n17136_), .B(new_n17135_), .ZN(new_n17137_));
  AOI21_X1   g16945(.A1(new_n17137_), .A2(new_n17129_), .B(new_n6356_), .ZN(new_n17138_));
  NOR2_X1    g16946(.A1(new_n16556_), .A2(new_n16543_), .ZN(new_n17139_));
  INV_X1     g16947(.I(new_n17139_), .ZN(new_n17140_));
  NAND3_X1   g16948(.A1(\asqrt[12] ), .A2(new_n16544_), .A3(new_n17140_), .ZN(new_n17141_));
  AND3_X2    g16949(.A1(new_n17140_), .A2(new_n16544_), .A3(new_n16549_), .Z(new_n17142_));
  AOI22_X1   g16950(.A1(new_n17141_), .A2(new_n16550_), .B1(\asqrt[12] ), .B2(new_n17142_), .ZN(new_n17143_));
  OAI21_X1   g16951(.A1(new_n17126_), .A2(new_n17127_), .B(new_n17120_), .ZN(new_n17144_));
  AOI21_X1   g16952(.A1(new_n17144_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n17145_));
  AOI21_X1   g16953(.A1(new_n17145_), .A2(new_n17137_), .B(new_n17143_), .ZN(new_n17146_));
  OAI21_X1   g16954(.A1(new_n17146_), .A2(new_n17138_), .B(\asqrt[34] ), .ZN(new_n17147_));
  INV_X1     g16955(.I(new_n17147_), .ZN(new_n17148_));
  NOR2_X1    g16956(.A1(new_n16567_), .A2(new_n16560_), .ZN(new_n17149_));
  NOR3_X1    g16957(.A1(new_n17149_), .A2(new_n16558_), .A3(new_n16566_), .ZN(new_n17150_));
  NOR3_X1    g16958(.A1(new_n16881_), .A2(new_n16558_), .A3(new_n17149_), .ZN(new_n17151_));
  INV_X1     g16959(.I(new_n17151_), .ZN(new_n17152_));
  AOI22_X1   g16960(.A1(new_n17152_), .A2(new_n16566_), .B1(\asqrt[12] ), .B2(new_n17150_), .ZN(new_n17153_));
  NOR3_X1    g16961(.A1(new_n17146_), .A2(new_n17138_), .A3(\asqrt[34] ), .ZN(new_n17154_));
  NOR2_X1    g16962(.A1(new_n17154_), .A2(new_n17153_), .ZN(new_n17155_));
  OAI21_X1   g16963(.A1(new_n17155_), .A2(new_n17148_), .B(\asqrt[35] ), .ZN(new_n17156_));
  INV_X1     g16964(.I(new_n16573_), .ZN(new_n17157_));
  NOR3_X1    g16965(.A1(new_n16881_), .A2(new_n16569_), .A3(new_n16633_), .ZN(new_n17158_));
  INV_X1     g16966(.I(new_n17158_), .ZN(new_n17159_));
  NOR3_X1    g16967(.A1(new_n16569_), .A2(new_n17157_), .A3(new_n16633_), .ZN(new_n17160_));
  AOI22_X1   g16968(.A1(new_n17159_), .A2(new_n17157_), .B1(\asqrt[12] ), .B2(new_n17160_), .ZN(new_n17161_));
  INV_X1     g16969(.I(new_n17161_), .ZN(new_n17162_));
  NAND2_X1   g16970(.A1(new_n17147_), .A2(new_n5708_), .ZN(new_n17163_));
  OAI21_X1   g16971(.A1(new_n17155_), .A2(new_n17163_), .B(new_n17162_), .ZN(new_n17164_));
  AOI21_X1   g16972(.A1(new_n17164_), .A2(new_n17156_), .B(new_n5277_), .ZN(new_n17165_));
  NOR2_X1    g16973(.A1(new_n16588_), .A2(new_n16575_), .ZN(new_n17166_));
  INV_X1     g16974(.I(new_n17166_), .ZN(new_n17167_));
  AND3_X2    g16975(.A1(new_n17167_), .A2(new_n16576_), .A3(new_n16581_), .Z(new_n17168_));
  NAND3_X1   g16976(.A1(\asqrt[12] ), .A2(new_n16576_), .A3(new_n17167_), .ZN(new_n17169_));
  AOI22_X1   g16977(.A1(new_n17169_), .A2(new_n16582_), .B1(\asqrt[12] ), .B2(new_n17168_), .ZN(new_n17170_));
  OAI21_X1   g16978(.A1(new_n17153_), .A2(new_n17154_), .B(new_n17147_), .ZN(new_n17171_));
  AOI21_X1   g16979(.A1(new_n17171_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n17172_));
  AOI21_X1   g16980(.A1(new_n17172_), .A2(new_n17164_), .B(new_n17170_), .ZN(new_n17173_));
  OAI21_X1   g16981(.A1(new_n17173_), .A2(new_n17165_), .B(\asqrt[37] ), .ZN(new_n17174_));
  INV_X1     g16982(.I(new_n17174_), .ZN(new_n17175_));
  NOR2_X1    g16983(.A1(new_n16592_), .A2(new_n16599_), .ZN(new_n17176_));
  NOR3_X1    g16984(.A1(new_n16881_), .A2(new_n16606_), .A3(new_n17176_), .ZN(new_n17177_));
  INV_X1     g16985(.I(new_n17177_), .ZN(new_n17178_));
  NOR3_X1    g16986(.A1(new_n17176_), .A2(new_n16606_), .A3(new_n16598_), .ZN(new_n17179_));
  AOI22_X1   g16987(.A1(new_n17178_), .A2(new_n16598_), .B1(\asqrt[12] ), .B2(new_n17179_), .ZN(new_n17180_));
  NOR3_X1    g16988(.A1(new_n17173_), .A2(new_n17165_), .A3(\asqrt[37] ), .ZN(new_n17181_));
  NOR2_X1    g16989(.A1(new_n17181_), .A2(new_n17180_), .ZN(new_n17182_));
  OAI21_X1   g16990(.A1(new_n17182_), .A2(new_n17175_), .B(\asqrt[38] ), .ZN(new_n17183_));
  INV_X1     g16991(.I(new_n16605_), .ZN(new_n17184_));
  NOR3_X1    g16992(.A1(new_n16601_), .A2(new_n17184_), .A3(new_n16650_), .ZN(new_n17185_));
  NOR3_X1    g16993(.A1(new_n16881_), .A2(new_n16601_), .A3(new_n16650_), .ZN(new_n17186_));
  INV_X1     g16994(.I(new_n17186_), .ZN(new_n17187_));
  AOI22_X1   g16995(.A1(new_n17187_), .A2(new_n17184_), .B1(\asqrt[12] ), .B2(new_n17185_), .ZN(new_n17188_));
  INV_X1     g16996(.I(new_n17188_), .ZN(new_n17189_));
  NAND2_X1   g16997(.A1(new_n17174_), .A2(new_n4696_), .ZN(new_n17190_));
  OAI21_X1   g16998(.A1(new_n17182_), .A2(new_n17190_), .B(new_n17189_), .ZN(new_n17191_));
  AOI21_X1   g16999(.A1(new_n17191_), .A2(new_n17183_), .B(new_n4298_), .ZN(new_n17192_));
  NOR3_X1    g17000(.A1(new_n16881_), .A2(new_n16610_), .A3(new_n16616_), .ZN(new_n17193_));
  INV_X1     g17001(.I(new_n17193_), .ZN(new_n17194_));
  NOR3_X1    g17002(.A1(new_n16610_), .A2(new_n16632_), .A3(new_n16616_), .ZN(new_n17195_));
  AOI22_X1   g17003(.A1(new_n17194_), .A2(new_n16632_), .B1(\asqrt[12] ), .B2(new_n17195_), .ZN(new_n17196_));
  OAI21_X1   g17004(.A1(new_n17180_), .A2(new_n17181_), .B(new_n17174_), .ZN(new_n17197_));
  AOI21_X1   g17005(.A1(new_n17197_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n17198_));
  AOI21_X1   g17006(.A1(new_n17198_), .A2(new_n17191_), .B(new_n17196_), .ZN(new_n17199_));
  OAI21_X1   g17007(.A1(new_n17199_), .A2(new_n17192_), .B(\asqrt[40] ), .ZN(new_n17200_));
  INV_X1     g17008(.I(new_n17200_), .ZN(new_n17201_));
  NOR2_X1    g17009(.A1(new_n16617_), .A2(new_n16625_), .ZN(new_n17202_));
  NOR3_X1    g17010(.A1(new_n17202_), .A2(new_n16640_), .A3(new_n16624_), .ZN(new_n17203_));
  NOR3_X1    g17011(.A1(new_n16881_), .A2(new_n16640_), .A3(new_n17202_), .ZN(new_n17204_));
  INV_X1     g17012(.I(new_n17204_), .ZN(new_n17205_));
  AOI22_X1   g17013(.A1(new_n17205_), .A2(new_n16624_), .B1(\asqrt[12] ), .B2(new_n17203_), .ZN(new_n17206_));
  NOR3_X1    g17014(.A1(new_n17199_), .A2(new_n17192_), .A3(\asqrt[40] ), .ZN(new_n17207_));
  NOR2_X1    g17015(.A1(new_n17207_), .A2(new_n17206_), .ZN(new_n17208_));
  OAI21_X1   g17016(.A1(new_n17208_), .A2(new_n17201_), .B(\asqrt[41] ), .ZN(new_n17209_));
  INV_X1     g17017(.I(new_n16631_), .ZN(new_n17210_));
  NOR3_X1    g17018(.A1(new_n16881_), .A2(new_n16627_), .A3(new_n16663_), .ZN(new_n17211_));
  INV_X1     g17019(.I(new_n17211_), .ZN(new_n17212_));
  NOR3_X1    g17020(.A1(new_n16627_), .A2(new_n17210_), .A3(new_n16663_), .ZN(new_n17213_));
  AOI22_X1   g17021(.A1(new_n17212_), .A2(new_n17210_), .B1(\asqrt[12] ), .B2(new_n17213_), .ZN(new_n17214_));
  INV_X1     g17022(.I(new_n17214_), .ZN(new_n17215_));
  NAND2_X1   g17023(.A1(new_n17200_), .A2(new_n3782_), .ZN(new_n17216_));
  OAI21_X1   g17024(.A1(new_n17208_), .A2(new_n17216_), .B(new_n17215_), .ZN(new_n17217_));
  AOI21_X1   g17025(.A1(new_n17217_), .A2(new_n17209_), .B(new_n3419_), .ZN(new_n17218_));
  NOR3_X1    g17026(.A1(new_n16901_), .A2(new_n16649_), .A3(new_n16902_), .ZN(new_n17219_));
  NOR3_X1    g17027(.A1(new_n16881_), .A2(new_n16901_), .A3(new_n16902_), .ZN(new_n17220_));
  INV_X1     g17028(.I(new_n17220_), .ZN(new_n17221_));
  AOI22_X1   g17029(.A1(new_n17221_), .A2(new_n16649_), .B1(\asqrt[12] ), .B2(new_n17219_), .ZN(new_n17222_));
  OAI21_X1   g17030(.A1(new_n17206_), .A2(new_n17207_), .B(new_n17200_), .ZN(new_n17223_));
  AOI21_X1   g17031(.A1(new_n17223_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n17224_));
  AOI21_X1   g17032(.A1(new_n17224_), .A2(new_n17217_), .B(new_n17222_), .ZN(new_n17225_));
  OAI21_X1   g17033(.A1(new_n17225_), .A2(new_n17218_), .B(\asqrt[43] ), .ZN(new_n17226_));
  INV_X1     g17034(.I(new_n17226_), .ZN(new_n17227_));
  INV_X1     g17035(.I(new_n16662_), .ZN(new_n17228_));
  NAND2_X1   g17036(.A1(new_n16643_), .A2(new_n3419_), .ZN(new_n17229_));
  NOR2_X1    g17037(.A1(new_n16903_), .A2(new_n17229_), .ZN(new_n17230_));
  NOR3_X1    g17038(.A1(new_n16881_), .A2(new_n16657_), .A3(new_n17230_), .ZN(new_n17231_));
  INV_X1     g17039(.I(new_n17231_), .ZN(new_n17232_));
  NOR3_X1    g17040(.A1(new_n17230_), .A2(new_n16657_), .A3(new_n17228_), .ZN(new_n17233_));
  AOI22_X1   g17041(.A1(new_n17232_), .A2(new_n17228_), .B1(\asqrt[12] ), .B2(new_n17233_), .ZN(new_n17234_));
  NOR3_X1    g17042(.A1(new_n17225_), .A2(new_n17218_), .A3(\asqrt[43] ), .ZN(new_n17235_));
  NOR2_X1    g17043(.A1(new_n17235_), .A2(new_n17234_), .ZN(new_n17236_));
  OAI21_X1   g17044(.A1(new_n17236_), .A2(new_n17227_), .B(\asqrt[44] ), .ZN(new_n17237_));
  NOR3_X1    g17045(.A1(new_n16668_), .A2(new_n16673_), .A3(new_n16900_), .ZN(new_n17238_));
  NOR3_X1    g17046(.A1(new_n16881_), .A2(new_n16668_), .A3(new_n16673_), .ZN(new_n17239_));
  INV_X1     g17047(.I(new_n17239_), .ZN(new_n17240_));
  AOI22_X1   g17048(.A1(new_n17240_), .A2(new_n16900_), .B1(\asqrt[12] ), .B2(new_n17238_), .ZN(new_n17241_));
  INV_X1     g17049(.I(new_n17241_), .ZN(new_n17242_));
  NAND2_X1   g17050(.A1(new_n17226_), .A2(new_n2954_), .ZN(new_n17243_));
  OAI21_X1   g17051(.A1(new_n17236_), .A2(new_n17243_), .B(new_n17242_), .ZN(new_n17244_));
  AOI21_X1   g17052(.A1(new_n17244_), .A2(new_n17237_), .B(new_n2641_), .ZN(new_n17245_));
  INV_X1     g17053(.I(new_n16675_), .ZN(new_n17246_));
  NOR2_X1    g17054(.A1(new_n16674_), .A2(new_n16682_), .ZN(new_n17247_));
  NOR3_X1    g17055(.A1(new_n16881_), .A2(new_n17246_), .A3(new_n17247_), .ZN(new_n17248_));
  INV_X1     g17056(.I(new_n17248_), .ZN(new_n17249_));
  NOR3_X1    g17057(.A1(new_n17246_), .A2(new_n17247_), .A3(new_n16681_), .ZN(new_n17250_));
  AOI22_X1   g17058(.A1(new_n17249_), .A2(new_n16681_), .B1(\asqrt[12] ), .B2(new_n17250_), .ZN(new_n17251_));
  OAI21_X1   g17059(.A1(new_n17234_), .A2(new_n17235_), .B(new_n17226_), .ZN(new_n17252_));
  AOI21_X1   g17060(.A1(new_n17252_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n17253_));
  AOI21_X1   g17061(.A1(new_n17253_), .A2(new_n17244_), .B(new_n17251_), .ZN(new_n17254_));
  OAI21_X1   g17062(.A1(new_n17254_), .A2(new_n17245_), .B(\asqrt[46] ), .ZN(new_n17255_));
  INV_X1     g17063(.I(new_n17255_), .ZN(new_n17256_));
  INV_X1     g17064(.I(new_n16689_), .ZN(new_n17257_));
  INV_X1     g17065(.I(new_n16683_), .ZN(new_n17258_));
  INV_X1     g17066(.I(new_n16691_), .ZN(new_n17259_));
  NOR2_X1    g17067(.A1(new_n17259_), .A2(new_n17258_), .ZN(new_n17260_));
  NOR3_X1    g17068(.A1(new_n17260_), .A2(new_n16684_), .A3(new_n17257_), .ZN(new_n17261_));
  NOR3_X1    g17069(.A1(new_n16881_), .A2(new_n16684_), .A3(new_n17260_), .ZN(new_n17262_));
  INV_X1     g17070(.I(new_n17262_), .ZN(new_n17263_));
  AOI22_X1   g17071(.A1(new_n17263_), .A2(new_n17257_), .B1(\asqrt[12] ), .B2(new_n17261_), .ZN(new_n17264_));
  NOR3_X1    g17072(.A1(new_n17254_), .A2(new_n17245_), .A3(\asqrt[46] ), .ZN(new_n17265_));
  NOR2_X1    g17073(.A1(new_n17265_), .A2(new_n17264_), .ZN(new_n17266_));
  OAI21_X1   g17074(.A1(new_n17266_), .A2(new_n17256_), .B(\asqrt[47] ), .ZN(new_n17267_));
  NOR3_X1    g17075(.A1(new_n16881_), .A2(new_n16694_), .A3(new_n16699_), .ZN(new_n17268_));
  INV_X1     g17076(.I(new_n17268_), .ZN(new_n17269_));
  NOR3_X1    g17077(.A1(new_n16694_), .A2(new_n16899_), .A3(new_n16699_), .ZN(new_n17270_));
  AOI22_X1   g17078(.A1(new_n17269_), .A2(new_n16899_), .B1(\asqrt[12] ), .B2(new_n17270_), .ZN(new_n17271_));
  INV_X1     g17079(.I(new_n17271_), .ZN(new_n17272_));
  NAND2_X1   g17080(.A1(new_n17255_), .A2(new_n2229_), .ZN(new_n17273_));
  OAI21_X1   g17081(.A1(new_n17266_), .A2(new_n17273_), .B(new_n17272_), .ZN(new_n17274_));
  AOI21_X1   g17082(.A1(new_n17274_), .A2(new_n17267_), .B(new_n1956_), .ZN(new_n17275_));
  INV_X1     g17083(.I(new_n16701_), .ZN(new_n17276_));
  NOR2_X1    g17084(.A1(new_n16700_), .A2(new_n16708_), .ZN(new_n17277_));
  NOR3_X1    g17085(.A1(new_n17276_), .A2(new_n17277_), .A3(new_n16707_), .ZN(new_n17278_));
  NOR3_X1    g17086(.A1(new_n16881_), .A2(new_n17276_), .A3(new_n17277_), .ZN(new_n17279_));
  INV_X1     g17087(.I(new_n17279_), .ZN(new_n17280_));
  AOI22_X1   g17088(.A1(new_n17280_), .A2(new_n16707_), .B1(\asqrt[12] ), .B2(new_n17278_), .ZN(new_n17281_));
  OAI21_X1   g17089(.A1(new_n17264_), .A2(new_n17265_), .B(new_n17255_), .ZN(new_n17282_));
  AOI21_X1   g17090(.A1(new_n17282_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n17283_));
  AOI21_X1   g17091(.A1(new_n17283_), .A2(new_n17274_), .B(new_n17281_), .ZN(new_n17284_));
  OAI21_X1   g17092(.A1(new_n17284_), .A2(new_n17275_), .B(\asqrt[49] ), .ZN(new_n17285_));
  INV_X1     g17093(.I(new_n17285_), .ZN(new_n17286_));
  INV_X1     g17094(.I(new_n16715_), .ZN(new_n17287_));
  INV_X1     g17095(.I(new_n16709_), .ZN(new_n17288_));
  INV_X1     g17096(.I(new_n16717_), .ZN(new_n17289_));
  NOR2_X1    g17097(.A1(new_n17289_), .A2(new_n17288_), .ZN(new_n17290_));
  NOR3_X1    g17098(.A1(new_n16881_), .A2(new_n16710_), .A3(new_n17290_), .ZN(new_n17291_));
  INV_X1     g17099(.I(new_n17291_), .ZN(new_n17292_));
  NOR3_X1    g17100(.A1(new_n17290_), .A2(new_n16710_), .A3(new_n17287_), .ZN(new_n17293_));
  AOI22_X1   g17101(.A1(new_n17292_), .A2(new_n17287_), .B1(\asqrt[12] ), .B2(new_n17293_), .ZN(new_n17294_));
  NOR3_X1    g17102(.A1(new_n17284_), .A2(new_n17275_), .A3(\asqrt[49] ), .ZN(new_n17295_));
  NOR2_X1    g17103(.A1(new_n17295_), .A2(new_n17294_), .ZN(new_n17296_));
  OAI21_X1   g17104(.A1(new_n17296_), .A2(new_n17286_), .B(\asqrt[50] ), .ZN(new_n17297_));
  NOR3_X1    g17105(.A1(new_n16720_), .A2(new_n16898_), .A3(new_n16725_), .ZN(new_n17298_));
  NOR3_X1    g17106(.A1(new_n16881_), .A2(new_n16720_), .A3(new_n16725_), .ZN(new_n17299_));
  INV_X1     g17107(.I(new_n17299_), .ZN(new_n17300_));
  AOI22_X1   g17108(.A1(new_n17300_), .A2(new_n16898_), .B1(\asqrt[12] ), .B2(new_n17298_), .ZN(new_n17301_));
  INV_X1     g17109(.I(new_n17301_), .ZN(new_n17302_));
  NAND2_X1   g17110(.A1(new_n17285_), .A2(new_n1612_), .ZN(new_n17303_));
  OAI21_X1   g17111(.A1(new_n17296_), .A2(new_n17303_), .B(new_n17302_), .ZN(new_n17304_));
  AOI21_X1   g17112(.A1(new_n17304_), .A2(new_n17297_), .B(new_n1376_), .ZN(new_n17305_));
  INV_X1     g17113(.I(new_n16727_), .ZN(new_n17306_));
  NOR2_X1    g17114(.A1(new_n16726_), .A2(new_n16734_), .ZN(new_n17307_));
  NOR3_X1    g17115(.A1(new_n16881_), .A2(new_n17306_), .A3(new_n17307_), .ZN(new_n17308_));
  INV_X1     g17116(.I(new_n17308_), .ZN(new_n17309_));
  NOR3_X1    g17117(.A1(new_n17306_), .A2(new_n16733_), .A3(new_n17307_), .ZN(new_n17310_));
  AOI22_X1   g17118(.A1(new_n17309_), .A2(new_n16733_), .B1(\asqrt[12] ), .B2(new_n17310_), .ZN(new_n17311_));
  OAI21_X1   g17119(.A1(new_n17294_), .A2(new_n17295_), .B(new_n17285_), .ZN(new_n17312_));
  AOI21_X1   g17120(.A1(new_n17312_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n17313_));
  AOI21_X1   g17121(.A1(new_n17313_), .A2(new_n17304_), .B(new_n17311_), .ZN(new_n17314_));
  OAI21_X1   g17122(.A1(new_n17314_), .A2(new_n17305_), .B(\asqrt[52] ), .ZN(new_n17315_));
  INV_X1     g17123(.I(new_n17315_), .ZN(new_n17316_));
  INV_X1     g17124(.I(new_n16741_), .ZN(new_n17317_));
  INV_X1     g17125(.I(new_n16735_), .ZN(new_n17318_));
  INV_X1     g17126(.I(new_n16743_), .ZN(new_n17319_));
  NOR2_X1    g17127(.A1(new_n17319_), .A2(new_n17318_), .ZN(new_n17320_));
  NOR3_X1    g17128(.A1(new_n17320_), .A2(new_n16736_), .A3(new_n17317_), .ZN(new_n17321_));
  NOR3_X1    g17129(.A1(new_n16881_), .A2(new_n16736_), .A3(new_n17320_), .ZN(new_n17322_));
  INV_X1     g17130(.I(new_n17322_), .ZN(new_n17323_));
  AOI22_X1   g17131(.A1(new_n17323_), .A2(new_n17317_), .B1(\asqrt[12] ), .B2(new_n17321_), .ZN(new_n17324_));
  NOR3_X1    g17132(.A1(new_n17314_), .A2(new_n17305_), .A3(\asqrt[52] ), .ZN(new_n17325_));
  NOR2_X1    g17133(.A1(new_n17325_), .A2(new_n17324_), .ZN(new_n17326_));
  OAI21_X1   g17134(.A1(new_n17326_), .A2(new_n17316_), .B(\asqrt[53] ), .ZN(new_n17327_));
  NOR3_X1    g17135(.A1(new_n16881_), .A2(new_n16746_), .A3(new_n16788_), .ZN(new_n17328_));
  INV_X1     g17136(.I(new_n17328_), .ZN(new_n17329_));
  NOR3_X1    g17137(.A1(new_n16746_), .A2(new_n16897_), .A3(new_n16788_), .ZN(new_n17330_));
  AOI22_X1   g17138(.A1(new_n17329_), .A2(new_n16897_), .B1(\asqrt[12] ), .B2(new_n17330_), .ZN(new_n17331_));
  INV_X1     g17139(.I(new_n17331_), .ZN(new_n17332_));
  NAND2_X1   g17140(.A1(new_n17315_), .A2(new_n1103_), .ZN(new_n17333_));
  OAI21_X1   g17141(.A1(new_n17326_), .A2(new_n17333_), .B(new_n17332_), .ZN(new_n17334_));
  AOI21_X1   g17142(.A1(new_n17334_), .A2(new_n17327_), .B(new_n904_), .ZN(new_n17335_));
  INV_X1     g17143(.I(new_n16754_), .ZN(new_n17336_));
  NOR2_X1    g17144(.A1(new_n16761_), .A2(new_n16753_), .ZN(new_n17337_));
  NOR3_X1    g17145(.A1(new_n17336_), .A2(new_n16760_), .A3(new_n17337_), .ZN(new_n17338_));
  NOR3_X1    g17146(.A1(new_n16881_), .A2(new_n17336_), .A3(new_n17337_), .ZN(new_n17339_));
  INV_X1     g17147(.I(new_n17339_), .ZN(new_n17340_));
  AOI22_X1   g17148(.A1(new_n17340_), .A2(new_n16760_), .B1(\asqrt[12] ), .B2(new_n17338_), .ZN(new_n17341_));
  OAI21_X1   g17149(.A1(new_n17324_), .A2(new_n17325_), .B(new_n17315_), .ZN(new_n17342_));
  AOI21_X1   g17150(.A1(new_n17342_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n17343_));
  AOI21_X1   g17151(.A1(new_n17343_), .A2(new_n17334_), .B(new_n17341_), .ZN(new_n17344_));
  OAI21_X1   g17152(.A1(new_n17344_), .A2(new_n17335_), .B(\asqrt[55] ), .ZN(new_n17345_));
  INV_X1     g17153(.I(new_n17345_), .ZN(new_n17346_));
  NOR2_X1    g17154(.A1(new_n16772_), .A2(new_n16765_), .ZN(new_n17347_));
  NOR3_X1    g17155(.A1(new_n16881_), .A2(new_n16763_), .A3(new_n17347_), .ZN(new_n17348_));
  INV_X1     g17156(.I(new_n17348_), .ZN(new_n17349_));
  NOR3_X1    g17157(.A1(new_n17347_), .A2(new_n16763_), .A3(new_n16771_), .ZN(new_n17350_));
  AOI22_X1   g17158(.A1(new_n17349_), .A2(new_n16771_), .B1(\asqrt[12] ), .B2(new_n17350_), .ZN(new_n17351_));
  NOR3_X1    g17159(.A1(new_n17344_), .A2(new_n17335_), .A3(\asqrt[55] ), .ZN(new_n17352_));
  NOR2_X1    g17160(.A1(new_n17352_), .A2(new_n17351_), .ZN(new_n17353_));
  OAI21_X1   g17161(.A1(new_n17353_), .A2(new_n17346_), .B(\asqrt[56] ), .ZN(new_n17354_));
  NOR3_X1    g17162(.A1(new_n16774_), .A2(new_n16896_), .A3(new_n16820_), .ZN(new_n17355_));
  NOR3_X1    g17163(.A1(new_n16881_), .A2(new_n16774_), .A3(new_n16820_), .ZN(new_n17356_));
  INV_X1     g17164(.I(new_n17356_), .ZN(new_n17357_));
  AOI22_X1   g17165(.A1(new_n17357_), .A2(new_n16896_), .B1(\asqrt[12] ), .B2(new_n17355_), .ZN(new_n17358_));
  INV_X1     g17166(.I(new_n17358_), .ZN(new_n17359_));
  NAND2_X1   g17167(.A1(new_n17345_), .A2(new_n703_), .ZN(new_n17360_));
  OAI21_X1   g17168(.A1(new_n17353_), .A2(new_n17360_), .B(new_n17359_), .ZN(new_n17361_));
  AOI21_X1   g17169(.A1(new_n17361_), .A2(new_n17354_), .B(new_n531_), .ZN(new_n17362_));
  INV_X1     g17170(.I(new_n16781_), .ZN(new_n17363_));
  NOR2_X1    g17171(.A1(new_n16793_), .A2(new_n16780_), .ZN(new_n17364_));
  NOR3_X1    g17172(.A1(new_n16881_), .A2(new_n17363_), .A3(new_n17364_), .ZN(new_n17365_));
  INV_X1     g17173(.I(new_n17365_), .ZN(new_n17366_));
  NOR3_X1    g17174(.A1(new_n17363_), .A2(new_n16787_), .A3(new_n17364_), .ZN(new_n17367_));
  AOI22_X1   g17175(.A1(new_n17366_), .A2(new_n16787_), .B1(\asqrt[12] ), .B2(new_n17367_), .ZN(new_n17368_));
  OAI21_X1   g17176(.A1(new_n17351_), .A2(new_n17352_), .B(new_n17345_), .ZN(new_n17369_));
  AOI21_X1   g17177(.A1(new_n17369_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n17370_));
  AOI21_X1   g17178(.A1(new_n17370_), .A2(new_n17361_), .B(new_n17368_), .ZN(new_n17371_));
  OAI21_X1   g17179(.A1(new_n17371_), .A2(new_n17362_), .B(\asqrt[58] ), .ZN(new_n17372_));
  NOR2_X1    g17180(.A1(new_n16804_), .A2(new_n16797_), .ZN(new_n17373_));
  NOR3_X1    g17181(.A1(new_n17373_), .A2(new_n16795_), .A3(new_n16803_), .ZN(new_n17374_));
  NOR3_X1    g17182(.A1(new_n16881_), .A2(new_n16795_), .A3(new_n17373_), .ZN(new_n17375_));
  INV_X1     g17183(.I(new_n17375_), .ZN(new_n17376_));
  AOI22_X1   g17184(.A1(new_n17376_), .A2(new_n16803_), .B1(\asqrt[12] ), .B2(new_n17374_), .ZN(new_n17377_));
  INV_X1     g17185(.I(new_n17377_), .ZN(new_n17378_));
  INV_X1     g17186(.I(new_n17351_), .ZN(new_n17379_));
  INV_X1     g17187(.I(new_n17324_), .ZN(new_n17380_));
  INV_X1     g17188(.I(new_n17294_), .ZN(new_n17381_));
  INV_X1     g17189(.I(new_n17264_), .ZN(new_n17382_));
  INV_X1     g17190(.I(new_n17234_), .ZN(new_n17383_));
  INV_X1     g17191(.I(new_n17206_), .ZN(new_n17384_));
  INV_X1     g17192(.I(new_n17180_), .ZN(new_n17385_));
  INV_X1     g17193(.I(new_n17153_), .ZN(new_n17386_));
  INV_X1     g17194(.I(new_n17126_), .ZN(new_n17387_));
  INV_X1     g17195(.I(new_n17099_), .ZN(new_n17388_));
  INV_X1     g17196(.I(new_n17069_), .ZN(new_n17389_));
  INV_X1     g17197(.I(new_n17038_), .ZN(new_n17390_));
  INV_X1     g17198(.I(new_n17012_), .ZN(new_n17391_));
  NAND2_X1   g17199(.A1(new_n16954_), .A2(new_n14601_), .ZN(new_n17392_));
  OAI21_X1   g17200(.A1(new_n17392_), .A2(new_n16986_), .B(new_n16968_), .ZN(new_n17393_));
  AOI21_X1   g17201(.A1(new_n17393_), .A2(new_n16996_), .B(new_n14017_), .ZN(new_n17394_));
  NOR2_X1    g17202(.A1(new_n16962_), .A2(\asqrt[17] ), .ZN(new_n17395_));
  AOI21_X1   g17203(.A1(new_n17395_), .A2(new_n17393_), .B(new_n16994_), .ZN(new_n17396_));
  OAI21_X1   g17204(.A1(new_n17396_), .A2(new_n17394_), .B(\asqrt[18] ), .ZN(new_n17397_));
  NAND2_X1   g17205(.A1(new_n17397_), .A2(new_n12913_), .ZN(new_n17398_));
  OAI21_X1   g17206(.A1(new_n17398_), .A2(new_n17006_), .B(new_n17391_), .ZN(new_n17399_));
  NAND3_X1   g17207(.A1(new_n17399_), .A2(new_n12364_), .A3(new_n17007_), .ZN(new_n17400_));
  AOI22_X1   g17208(.A1(new_n17400_), .A2(new_n17021_), .B1(\asqrt[20] ), .B2(new_n17029_), .ZN(new_n17401_));
  OAI21_X1   g17209(.A1(new_n17401_), .A2(new_n11736_), .B(new_n11326_), .ZN(new_n17402_));
  OAI21_X1   g17210(.A1(new_n17402_), .A2(new_n17031_), .B(new_n17390_), .ZN(new_n17403_));
  AOI21_X1   g17211(.A1(new_n17403_), .A2(new_n17032_), .B(new_n10812_), .ZN(new_n17404_));
  AOI21_X1   g17212(.A1(new_n17399_), .A2(new_n17007_), .B(new_n12364_), .ZN(new_n17405_));
  NOR3_X1    g17213(.A1(new_n17396_), .A2(new_n17394_), .A3(\asqrt[18] ), .ZN(new_n17406_));
  OAI21_X1   g17214(.A1(new_n17003_), .A2(new_n17406_), .B(new_n17397_), .ZN(new_n17407_));
  AOI21_X1   g17215(.A1(new_n17407_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n17408_));
  AOI21_X1   g17216(.A1(new_n17408_), .A2(new_n17399_), .B(new_n17020_), .ZN(new_n17409_));
  NOR3_X1    g17217(.A1(new_n17409_), .A2(\asqrt[21] ), .A3(new_n17405_), .ZN(new_n17410_));
  OAI22_X1   g17218(.A1(new_n17410_), .A2(new_n17028_), .B1(new_n17401_), .B2(new_n11736_), .ZN(new_n17411_));
  AOI21_X1   g17219(.A1(new_n17411_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n17412_));
  AOI21_X1   g17220(.A1(new_n17412_), .A2(new_n17403_), .B(new_n17046_), .ZN(new_n17413_));
  OAI21_X1   g17221(.A1(new_n17413_), .A2(new_n17404_), .B(\asqrt[24] ), .ZN(new_n17414_));
  NAND2_X1   g17222(.A1(new_n17414_), .A2(new_n9846_), .ZN(new_n17415_));
  OAI21_X1   g17223(.A1(new_n17415_), .A2(new_n17059_), .B(new_n17389_), .ZN(new_n17416_));
  AOI21_X1   g17224(.A1(new_n17416_), .A2(new_n17060_), .B(new_n9317_), .ZN(new_n17417_));
  NOR3_X1    g17225(.A1(new_n17413_), .A2(\asqrt[24] ), .A3(new_n17404_), .ZN(new_n17418_));
  OAI21_X1   g17226(.A1(new_n17056_), .A2(new_n17418_), .B(new_n17414_), .ZN(new_n17419_));
  AOI21_X1   g17227(.A1(new_n17419_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n17420_));
  AOI21_X1   g17228(.A1(new_n17420_), .A2(new_n17416_), .B(new_n17077_), .ZN(new_n17421_));
  OAI21_X1   g17229(.A1(new_n17421_), .A2(new_n17417_), .B(\asqrt[27] ), .ZN(new_n17422_));
  NAND2_X1   g17230(.A1(new_n17422_), .A2(new_n8483_), .ZN(new_n17423_));
  OAI21_X1   g17231(.A1(new_n17423_), .A2(new_n17089_), .B(new_n17388_), .ZN(new_n17424_));
  AOI21_X1   g17232(.A1(new_n17424_), .A2(new_n17090_), .B(new_n8036_), .ZN(new_n17425_));
  NOR3_X1    g17233(.A1(new_n17421_), .A2(\asqrt[27] ), .A3(new_n17417_), .ZN(new_n17426_));
  OAI21_X1   g17234(.A1(new_n17086_), .A2(new_n17426_), .B(new_n17422_), .ZN(new_n17427_));
  AOI21_X1   g17235(.A1(new_n17427_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n17428_));
  AOI21_X1   g17236(.A1(new_n17428_), .A2(new_n17424_), .B(new_n17107_), .ZN(new_n17429_));
  OAI21_X1   g17237(.A1(new_n17429_), .A2(new_n17425_), .B(\asqrt[30] ), .ZN(new_n17430_));
  NAND2_X1   g17238(.A1(new_n17430_), .A2(new_n7229_), .ZN(new_n17431_));
  OAI21_X1   g17239(.A1(new_n17431_), .A2(new_n17119_), .B(new_n17387_), .ZN(new_n17432_));
  AOI21_X1   g17240(.A1(new_n17432_), .A2(new_n17120_), .B(new_n6824_), .ZN(new_n17433_));
  NOR3_X1    g17241(.A1(new_n17429_), .A2(\asqrt[30] ), .A3(new_n17425_), .ZN(new_n17434_));
  OAI21_X1   g17242(.A1(new_n17116_), .A2(new_n17434_), .B(new_n17430_), .ZN(new_n17435_));
  AOI21_X1   g17243(.A1(new_n17435_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n17436_));
  AOI21_X1   g17244(.A1(new_n17436_), .A2(new_n17432_), .B(new_n17134_), .ZN(new_n17437_));
  OAI21_X1   g17245(.A1(new_n17437_), .A2(new_n17433_), .B(\asqrt[33] ), .ZN(new_n17438_));
  NAND2_X1   g17246(.A1(new_n17438_), .A2(new_n6077_), .ZN(new_n17439_));
  OAI21_X1   g17247(.A1(new_n17439_), .A2(new_n17146_), .B(new_n17386_), .ZN(new_n17440_));
  AOI21_X1   g17248(.A1(new_n17440_), .A2(new_n17147_), .B(new_n5708_), .ZN(new_n17441_));
  NOR3_X1    g17249(.A1(new_n17437_), .A2(\asqrt[33] ), .A3(new_n17433_), .ZN(new_n17442_));
  OAI21_X1   g17250(.A1(new_n17143_), .A2(new_n17442_), .B(new_n17438_), .ZN(new_n17443_));
  AOI21_X1   g17251(.A1(new_n17443_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n17444_));
  AOI21_X1   g17252(.A1(new_n17444_), .A2(new_n17440_), .B(new_n17161_), .ZN(new_n17445_));
  OAI21_X1   g17253(.A1(new_n17445_), .A2(new_n17441_), .B(\asqrt[36] ), .ZN(new_n17446_));
  NAND2_X1   g17254(.A1(new_n17446_), .A2(new_n5024_), .ZN(new_n17447_));
  OAI21_X1   g17255(.A1(new_n17447_), .A2(new_n17173_), .B(new_n17385_), .ZN(new_n17448_));
  AOI21_X1   g17256(.A1(new_n17448_), .A2(new_n17174_), .B(new_n4696_), .ZN(new_n17449_));
  NOR3_X1    g17257(.A1(new_n17445_), .A2(\asqrt[36] ), .A3(new_n17441_), .ZN(new_n17450_));
  OAI21_X1   g17258(.A1(new_n17170_), .A2(new_n17450_), .B(new_n17446_), .ZN(new_n17451_));
  AOI21_X1   g17259(.A1(new_n17451_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n17452_));
  AOI21_X1   g17260(.A1(new_n17452_), .A2(new_n17448_), .B(new_n17188_), .ZN(new_n17453_));
  OAI21_X1   g17261(.A1(new_n17453_), .A2(new_n17449_), .B(\asqrt[39] ), .ZN(new_n17454_));
  NAND2_X1   g17262(.A1(new_n17454_), .A2(new_n4071_), .ZN(new_n17455_));
  OAI21_X1   g17263(.A1(new_n17455_), .A2(new_n17199_), .B(new_n17384_), .ZN(new_n17456_));
  AOI21_X1   g17264(.A1(new_n17456_), .A2(new_n17200_), .B(new_n3782_), .ZN(new_n17457_));
  NOR3_X1    g17265(.A1(new_n17453_), .A2(\asqrt[39] ), .A3(new_n17449_), .ZN(new_n17458_));
  OAI21_X1   g17266(.A1(new_n17196_), .A2(new_n17458_), .B(new_n17454_), .ZN(new_n17459_));
  AOI21_X1   g17267(.A1(new_n17459_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n17460_));
  AOI21_X1   g17268(.A1(new_n17460_), .A2(new_n17456_), .B(new_n17214_), .ZN(new_n17461_));
  OAI21_X1   g17269(.A1(new_n17461_), .A2(new_n17457_), .B(\asqrt[42] ), .ZN(new_n17462_));
  NAND2_X1   g17270(.A1(new_n17462_), .A2(new_n3218_), .ZN(new_n17463_));
  OAI21_X1   g17271(.A1(new_n17463_), .A2(new_n17225_), .B(new_n17383_), .ZN(new_n17464_));
  AOI21_X1   g17272(.A1(new_n17464_), .A2(new_n17226_), .B(new_n2954_), .ZN(new_n17465_));
  NOR3_X1    g17273(.A1(new_n17461_), .A2(\asqrt[42] ), .A3(new_n17457_), .ZN(new_n17466_));
  OAI21_X1   g17274(.A1(new_n17222_), .A2(new_n17466_), .B(new_n17462_), .ZN(new_n17467_));
  AOI21_X1   g17275(.A1(new_n17467_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n17468_));
  AOI21_X1   g17276(.A1(new_n17468_), .A2(new_n17464_), .B(new_n17241_), .ZN(new_n17469_));
  OAI21_X1   g17277(.A1(new_n17469_), .A2(new_n17465_), .B(\asqrt[45] ), .ZN(new_n17470_));
  NAND2_X1   g17278(.A1(new_n17470_), .A2(new_n2465_), .ZN(new_n17471_));
  OAI21_X1   g17279(.A1(new_n17471_), .A2(new_n17254_), .B(new_n17382_), .ZN(new_n17472_));
  AOI21_X1   g17280(.A1(new_n17472_), .A2(new_n17255_), .B(new_n2229_), .ZN(new_n17473_));
  NOR3_X1    g17281(.A1(new_n17469_), .A2(\asqrt[45] ), .A3(new_n17465_), .ZN(new_n17474_));
  OAI21_X1   g17282(.A1(new_n17251_), .A2(new_n17474_), .B(new_n17470_), .ZN(new_n17475_));
  AOI21_X1   g17283(.A1(new_n17475_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n17476_));
  AOI21_X1   g17284(.A1(new_n17476_), .A2(new_n17472_), .B(new_n17271_), .ZN(new_n17477_));
  OAI21_X1   g17285(.A1(new_n17477_), .A2(new_n17473_), .B(\asqrt[48] ), .ZN(new_n17478_));
  NAND2_X1   g17286(.A1(new_n17478_), .A2(new_n1806_), .ZN(new_n17479_));
  OAI21_X1   g17287(.A1(new_n17479_), .A2(new_n17284_), .B(new_n17381_), .ZN(new_n17480_));
  AOI21_X1   g17288(.A1(new_n17480_), .A2(new_n17285_), .B(new_n1612_), .ZN(new_n17481_));
  NOR3_X1    g17289(.A1(new_n17477_), .A2(\asqrt[48] ), .A3(new_n17473_), .ZN(new_n17482_));
  OAI21_X1   g17290(.A1(new_n17281_), .A2(new_n17482_), .B(new_n17478_), .ZN(new_n17483_));
  AOI21_X1   g17291(.A1(new_n17483_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n17484_));
  AOI21_X1   g17292(.A1(new_n17484_), .A2(new_n17480_), .B(new_n17301_), .ZN(new_n17485_));
  OAI21_X1   g17293(.A1(new_n17485_), .A2(new_n17481_), .B(\asqrt[51] ), .ZN(new_n17486_));
  NAND2_X1   g17294(.A1(new_n17486_), .A2(new_n1256_), .ZN(new_n17487_));
  OAI21_X1   g17295(.A1(new_n17487_), .A2(new_n17314_), .B(new_n17380_), .ZN(new_n17488_));
  NAND3_X1   g17296(.A1(new_n17488_), .A2(new_n1103_), .A3(new_n17315_), .ZN(new_n17489_));
  AOI22_X1   g17297(.A1(new_n17489_), .A2(new_n17332_), .B1(\asqrt[53] ), .B2(new_n17342_), .ZN(new_n17490_));
  OAI21_X1   g17298(.A1(new_n17490_), .A2(new_n904_), .B(new_n823_), .ZN(new_n17491_));
  OAI21_X1   g17299(.A1(new_n17491_), .A2(new_n17344_), .B(new_n17379_), .ZN(new_n17492_));
  NAND3_X1   g17300(.A1(new_n17492_), .A2(new_n703_), .A3(new_n17345_), .ZN(new_n17493_));
  AOI22_X1   g17301(.A1(new_n17493_), .A2(new_n17359_), .B1(\asqrt[56] ), .B2(new_n17369_), .ZN(new_n17494_));
  OAI21_X1   g17302(.A1(new_n17494_), .A2(new_n531_), .B(new_n436_), .ZN(new_n17495_));
  OAI21_X1   g17303(.A1(new_n17495_), .A2(new_n17371_), .B(new_n17378_), .ZN(new_n17496_));
  AOI21_X1   g17304(.A1(new_n17496_), .A2(new_n17372_), .B(new_n327_), .ZN(new_n17497_));
  NOR3_X1    g17305(.A1(new_n16881_), .A2(new_n16806_), .A3(new_n16852_), .ZN(new_n17498_));
  INV_X1     g17306(.I(new_n17498_), .ZN(new_n17499_));
  NOR3_X1    g17307(.A1(new_n16806_), .A2(new_n16895_), .A3(new_n16852_), .ZN(new_n17500_));
  AOI22_X1   g17308(.A1(new_n17499_), .A2(new_n16895_), .B1(\asqrt[12] ), .B2(new_n17500_), .ZN(new_n17501_));
  NAND2_X1   g17309(.A1(new_n17372_), .A2(new_n327_), .ZN(new_n17502_));
  INV_X1     g17310(.I(new_n17502_), .ZN(new_n17503_));
  AOI21_X1   g17311(.A1(new_n17503_), .A2(new_n17496_), .B(new_n17501_), .ZN(new_n17504_));
  OAI21_X1   g17312(.A1(new_n17504_), .A2(new_n17497_), .B(\asqrt[60] ), .ZN(new_n17505_));
  INV_X1     g17313(.I(new_n16813_), .ZN(new_n17506_));
  NOR2_X1    g17314(.A1(new_n16825_), .A2(new_n16812_), .ZN(new_n17507_));
  NOR3_X1    g17315(.A1(new_n17506_), .A2(new_n16819_), .A3(new_n17507_), .ZN(new_n17508_));
  NOR3_X1    g17316(.A1(new_n16881_), .A2(new_n17506_), .A3(new_n17507_), .ZN(new_n17509_));
  INV_X1     g17317(.I(new_n17509_), .ZN(new_n17510_));
  AOI22_X1   g17318(.A1(new_n17510_), .A2(new_n16819_), .B1(\asqrt[12] ), .B2(new_n17508_), .ZN(new_n17511_));
  INV_X1     g17319(.I(new_n17511_), .ZN(new_n17512_));
  INV_X1     g17320(.I(new_n17372_), .ZN(new_n17513_));
  NOR3_X1    g17321(.A1(new_n17371_), .A2(new_n17362_), .A3(\asqrt[58] ), .ZN(new_n17514_));
  NOR2_X1    g17322(.A1(new_n17514_), .A2(new_n17377_), .ZN(new_n17515_));
  OAI21_X1   g17323(.A1(new_n17515_), .A2(new_n17513_), .B(\asqrt[59] ), .ZN(new_n17516_));
  NAND2_X1   g17324(.A1(new_n17516_), .A2(new_n306_), .ZN(new_n17517_));
  OAI21_X1   g17325(.A1(new_n17517_), .A2(new_n17504_), .B(new_n17512_), .ZN(new_n17518_));
  AOI21_X1   g17326(.A1(new_n17518_), .A2(new_n17505_), .B(new_n218_), .ZN(new_n17519_));
  NOR2_X1    g17327(.A1(new_n16829_), .A2(new_n16836_), .ZN(new_n17520_));
  NOR3_X1    g17328(.A1(new_n16881_), .A2(new_n16827_), .A3(new_n17520_), .ZN(new_n17521_));
  INV_X1     g17329(.I(new_n17521_), .ZN(new_n17522_));
  NOR3_X1    g17330(.A1(new_n17520_), .A2(new_n16827_), .A3(new_n16835_), .ZN(new_n17523_));
  AOI22_X1   g17331(.A1(new_n17522_), .A2(new_n16835_), .B1(\asqrt[12] ), .B2(new_n17523_), .ZN(new_n17524_));
  INV_X1     g17332(.I(new_n17501_), .ZN(new_n17525_));
  OAI21_X1   g17333(.A1(new_n17515_), .A2(new_n17502_), .B(new_n17525_), .ZN(new_n17526_));
  AOI21_X1   g17334(.A1(new_n17526_), .A2(new_n17516_), .B(new_n306_), .ZN(new_n17527_));
  NOR2_X1    g17335(.A1(new_n17527_), .A2(\asqrt[61] ), .ZN(new_n17528_));
  AOI21_X1   g17336(.A1(new_n17528_), .A2(new_n17518_), .B(new_n17524_), .ZN(new_n17529_));
  OAI21_X1   g17337(.A1(new_n17529_), .A2(new_n17519_), .B(\asqrt[62] ), .ZN(new_n17530_));
  NOR3_X1    g17338(.A1(new_n16838_), .A2(new_n16894_), .A3(new_n16892_), .ZN(new_n17531_));
  NOR3_X1    g17339(.A1(new_n16881_), .A2(new_n16838_), .A3(new_n16892_), .ZN(new_n17532_));
  INV_X1     g17340(.I(new_n17532_), .ZN(new_n17533_));
  AOI22_X1   g17341(.A1(new_n17533_), .A2(new_n16894_), .B1(\asqrt[12] ), .B2(new_n17531_), .ZN(new_n17534_));
  INV_X1     g17342(.I(new_n17534_), .ZN(new_n17535_));
  OAI21_X1   g17343(.A1(new_n17377_), .A2(new_n17514_), .B(new_n17372_), .ZN(new_n17536_));
  AOI21_X1   g17344(.A1(new_n17536_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n17537_));
  AOI21_X1   g17345(.A1(new_n17537_), .A2(new_n17526_), .B(new_n17511_), .ZN(new_n17538_));
  OAI21_X1   g17346(.A1(new_n17538_), .A2(new_n17527_), .B(\asqrt[61] ), .ZN(new_n17539_));
  NAND2_X1   g17347(.A1(new_n17539_), .A2(new_n207_), .ZN(new_n17540_));
  OAI21_X1   g17348(.A1(new_n17540_), .A2(new_n17529_), .B(new_n17535_), .ZN(new_n17541_));
  NAND4_X1   g17349(.A1(\asqrt[12] ), .A2(new_n16845_), .A3(new_n16850_), .A4(new_n16931_), .ZN(new_n17542_));
  NAND2_X1   g17350(.A1(new_n16845_), .A2(new_n16931_), .ZN(new_n17543_));
  OAI21_X1   g17351(.A1(new_n16881_), .A2(new_n17543_), .B(new_n16851_), .ZN(new_n17544_));
  NAND2_X1   g17352(.A1(new_n17542_), .A2(new_n17544_), .ZN(new_n17545_));
  NOR2_X1    g17353(.A1(new_n16932_), .A2(new_n16871_), .ZN(new_n17546_));
  NAND2_X1   g17354(.A1(\asqrt[12] ), .A2(new_n17546_), .ZN(new_n17547_));
  NAND3_X1   g17355(.A1(new_n17545_), .A2(new_n16943_), .A3(new_n17547_), .ZN(new_n17548_));
  AOI21_X1   g17356(.A1(new_n17541_), .A2(new_n17530_), .B(new_n17548_), .ZN(new_n17549_));
  NOR3_X1    g17357(.A1(new_n17538_), .A2(new_n17527_), .A3(\asqrt[61] ), .ZN(new_n17550_));
  OAI21_X1   g17358(.A1(new_n17524_), .A2(new_n17550_), .B(new_n17539_), .ZN(new_n17551_));
  AOI21_X1   g17359(.A1(new_n17551_), .A2(\asqrt[62] ), .B(new_n17545_), .ZN(new_n17552_));
  OAI21_X1   g17360(.A1(new_n16881_), .A2(new_n16871_), .B(new_n16932_), .ZN(new_n17553_));
  NOR2_X1    g17361(.A1(new_n17546_), .A2(new_n193_), .ZN(new_n17554_));
  NAND2_X1   g17362(.A1(new_n17553_), .A2(new_n17554_), .ZN(new_n17555_));
  INV_X1     g17363(.I(new_n17555_), .ZN(new_n17556_));
  AND3_X2    g17364(.A1(new_n16862_), .A2(new_n16860_), .A3(new_n16877_), .Z(new_n17557_));
  NAND4_X1   g17365(.A1(new_n16933_), .A2(new_n16943_), .A3(new_n16874_), .A4(new_n17557_), .ZN(new_n17558_));
  INV_X1     g17366(.I(new_n17558_), .ZN(new_n17559_));
  NOR2_X1    g17367(.A1(new_n17556_), .A2(new_n17559_), .ZN(new_n17560_));
  INV_X1     g17368(.I(new_n17560_), .ZN(new_n17561_));
  AOI21_X1   g17369(.A1(new_n17552_), .A2(new_n17541_), .B(new_n17561_), .ZN(new_n17562_));
  OAI21_X1   g17370(.A1(\asqrt[63] ), .A2(new_n17549_), .B(new_n17562_), .ZN(\asqrt[11] ));
  NOR2_X1    g17371(.A1(\a[20] ), .A2(\a[21] ), .ZN(new_n17564_));
  INV_X1     g17372(.I(new_n17564_), .ZN(new_n17565_));
  NOR2_X1    g17373(.A1(new_n17565_), .A2(\a[22] ), .ZN(new_n17566_));
  INV_X1     g17374(.I(new_n17566_), .ZN(new_n17567_));
  NAND2_X1   g17375(.A1(new_n17541_), .A2(new_n17530_), .ZN(new_n17568_));
  INV_X1     g17376(.I(new_n17548_), .ZN(new_n17569_));
  AOI21_X1   g17377(.A1(new_n17568_), .A2(new_n17569_), .B(\asqrt[63] ), .ZN(new_n17570_));
  INV_X1     g17378(.I(new_n17524_), .ZN(new_n17571_));
  NAND3_X1   g17379(.A1(new_n17496_), .A2(new_n327_), .A3(new_n17372_), .ZN(new_n17572_));
  AOI22_X1   g17380(.A1(new_n17572_), .A2(new_n17525_), .B1(new_n17536_), .B2(\asqrt[59] ), .ZN(new_n17573_));
  OAI21_X1   g17381(.A1(new_n17573_), .A2(new_n306_), .B(new_n218_), .ZN(new_n17574_));
  OAI21_X1   g17382(.A1(new_n17574_), .A2(new_n17538_), .B(new_n17571_), .ZN(new_n17575_));
  NOR2_X1    g17383(.A1(new_n17519_), .A2(\asqrt[62] ), .ZN(new_n17576_));
  AOI21_X1   g17384(.A1(new_n17576_), .A2(new_n17575_), .B(new_n17534_), .ZN(new_n17577_));
  INV_X1     g17385(.I(new_n17545_), .ZN(new_n17578_));
  NAND2_X1   g17386(.A1(new_n17530_), .A2(new_n17578_), .ZN(new_n17579_));
  OAI21_X1   g17387(.A1(new_n17579_), .A2(new_n17577_), .B(new_n17560_), .ZN(new_n17580_));
  OAI21_X1   g17388(.A1(new_n17570_), .A2(new_n17580_), .B(\a[22] ), .ZN(new_n17581_));
  AOI21_X1   g17389(.A1(new_n17581_), .A2(new_n17567_), .B(new_n16881_), .ZN(new_n17582_));
  INV_X1     g17390(.I(\a[22] ), .ZN(new_n17583_));
  NAND3_X1   g17391(.A1(new_n17575_), .A2(new_n207_), .A3(new_n17539_), .ZN(new_n17584_));
  AOI22_X1   g17392(.A1(new_n17584_), .A2(new_n17535_), .B1(new_n17551_), .B2(\asqrt[62] ), .ZN(new_n17585_));
  OAI21_X1   g17393(.A1(new_n17585_), .A2(new_n17548_), .B(new_n193_), .ZN(new_n17586_));
  AOI21_X1   g17394(.A1(new_n17586_), .A2(new_n17562_), .B(new_n17583_), .ZN(new_n17587_));
  NAND4_X1   g17395(.A1(new_n16943_), .A2(new_n16874_), .A3(new_n16877_), .A4(new_n17567_), .ZN(new_n17588_));
  NOR2_X1    g17396(.A1(new_n17588_), .A2(new_n16869_), .ZN(new_n17589_));
  INV_X1     g17397(.I(new_n17589_), .ZN(new_n17590_));
  NOR2_X1    g17398(.A1(new_n17587_), .A2(new_n17590_), .ZN(new_n17591_));
  AOI21_X1   g17399(.A1(new_n17586_), .A2(new_n17562_), .B(new_n16884_), .ZN(new_n17592_));
  INV_X1     g17400(.I(\a[23] ), .ZN(new_n17593_));
  AOI21_X1   g17401(.A1(\asqrt[11] ), .A2(new_n17583_), .B(new_n17593_), .ZN(new_n17594_));
  NOR3_X1    g17402(.A1(new_n17591_), .A2(new_n17594_), .A3(new_n17592_), .ZN(new_n17595_));
  OAI21_X1   g17403(.A1(new_n17595_), .A2(new_n17582_), .B(\asqrt[13] ), .ZN(new_n17596_));
  OAI21_X1   g17404(.A1(new_n17570_), .A2(new_n17580_), .B(new_n16883_), .ZN(new_n17597_));
  NAND2_X1   g17405(.A1(new_n17552_), .A2(new_n17541_), .ZN(new_n17598_));
  NOR3_X1    g17406(.A1(new_n17556_), .A2(new_n16881_), .A3(new_n17559_), .ZN(new_n17599_));
  NAND3_X1   g17407(.A1(new_n17586_), .A2(new_n17598_), .A3(new_n17599_), .ZN(new_n17600_));
  AOI21_X1   g17408(.A1(new_n17600_), .A2(new_n17597_), .B(new_n16882_), .ZN(new_n17601_));
  NAND2_X1   g17409(.A1(new_n17598_), .A2(new_n17599_), .ZN(new_n17602_));
  NOR2_X1    g17410(.A1(new_n17602_), .A2(new_n17570_), .ZN(new_n17603_));
  NOR3_X1    g17411(.A1(new_n17603_), .A2(new_n17592_), .A3(\a[24] ), .ZN(new_n17604_));
  AOI21_X1   g17412(.A1(\asqrt[11] ), .A2(\a[22] ), .B(new_n17566_), .ZN(new_n17605_));
  OAI21_X1   g17413(.A1(new_n17605_), .A2(new_n16881_), .B(new_n16389_), .ZN(new_n17606_));
  OAI22_X1   g17414(.A1(new_n17595_), .A2(new_n17606_), .B1(new_n17601_), .B2(new_n17604_), .ZN(new_n17607_));
  AOI21_X1   g17415(.A1(new_n17607_), .A2(new_n17596_), .B(new_n15770_), .ZN(new_n17608_));
  NOR3_X1    g17416(.A1(new_n16972_), .A2(new_n16973_), .A3(new_n16938_), .ZN(new_n17609_));
  NAND3_X1   g17417(.A1(\asqrt[11] ), .A2(new_n16971_), .A3(new_n16891_), .ZN(new_n17610_));
  AOI22_X1   g17418(.A1(new_n17610_), .A2(new_n16938_), .B1(\asqrt[11] ), .B2(new_n17609_), .ZN(new_n17611_));
  OAI21_X1   g17419(.A1(new_n17587_), .A2(new_n17566_), .B(\asqrt[12] ), .ZN(new_n17612_));
  AOI21_X1   g17420(.A1(new_n17586_), .A2(new_n17562_), .B(\a[22] ), .ZN(new_n17613_));
  OAI21_X1   g17421(.A1(new_n17593_), .A2(new_n17613_), .B(new_n17597_), .ZN(new_n17614_));
  OAI21_X1   g17422(.A1(new_n17614_), .A2(new_n17591_), .B(new_n17612_), .ZN(new_n17615_));
  AOI21_X1   g17423(.A1(new_n17615_), .A2(\asqrt[13] ), .B(\asqrt[14] ), .ZN(new_n17616_));
  AOI21_X1   g17424(.A1(new_n17616_), .A2(new_n17607_), .B(new_n17611_), .ZN(new_n17617_));
  OAI21_X1   g17425(.A1(new_n17617_), .A2(new_n17608_), .B(\asqrt[15] ), .ZN(new_n17618_));
  INV_X1     g17426(.I(new_n17618_), .ZN(new_n17619_));
  NOR2_X1    g17427(.A1(new_n16976_), .A2(new_n16979_), .ZN(new_n17620_));
  INV_X1     g17428(.I(new_n17620_), .ZN(new_n17621_));
  NAND4_X1   g17429(.A1(\asqrt[11] ), .A2(new_n16977_), .A3(new_n16951_), .A4(new_n17621_), .ZN(new_n17622_));
  INV_X1     g17430(.I(\asqrt[11] ), .ZN(new_n17623_));
  NOR3_X1    g17431(.A1(new_n17623_), .A2(new_n16940_), .A3(new_n17620_), .ZN(new_n17624_));
  OAI21_X1   g17432(.A1(new_n17624_), .A2(new_n16951_), .B(new_n17622_), .ZN(new_n17625_));
  INV_X1     g17433(.I(new_n17625_), .ZN(new_n17626_));
  NOR3_X1    g17434(.A1(new_n17617_), .A2(new_n17608_), .A3(\asqrt[15] ), .ZN(new_n17627_));
  NOR2_X1    g17435(.A1(new_n17627_), .A2(new_n17626_), .ZN(new_n17628_));
  OAI21_X1   g17436(.A1(new_n17628_), .A2(new_n17619_), .B(\asqrt[16] ), .ZN(new_n17629_));
  NAND2_X1   g17437(.A1(new_n16985_), .A2(new_n16980_), .ZN(new_n17630_));
  NAND3_X1   g17438(.A1(\asqrt[11] ), .A2(new_n16954_), .A3(new_n17630_), .ZN(new_n17631_));
  AND3_X2    g17439(.A1(new_n16954_), .A2(new_n16958_), .A3(new_n17630_), .Z(new_n17632_));
  AOI22_X1   g17440(.A1(new_n17631_), .A2(new_n16959_), .B1(\asqrt[11] ), .B2(new_n17632_), .ZN(new_n17633_));
  INV_X1     g17441(.I(new_n17633_), .ZN(new_n17634_));
  NAND2_X1   g17442(.A1(new_n17618_), .A2(new_n14601_), .ZN(new_n17635_));
  OAI21_X1   g17443(.A1(new_n17628_), .A2(new_n17635_), .B(new_n17634_), .ZN(new_n17636_));
  AOI21_X1   g17444(.A1(new_n17636_), .A2(new_n17629_), .B(new_n14017_), .ZN(new_n17637_));
  NOR3_X1    g17445(.A1(new_n16962_), .A2(new_n16968_), .A3(new_n16987_), .ZN(new_n17638_));
  NOR3_X1    g17446(.A1(new_n17623_), .A2(new_n16962_), .A3(new_n16987_), .ZN(new_n17639_));
  INV_X1     g17447(.I(new_n17639_), .ZN(new_n17640_));
  AOI22_X1   g17448(.A1(new_n17640_), .A2(new_n16968_), .B1(\asqrt[11] ), .B2(new_n17638_), .ZN(new_n17641_));
  OAI21_X1   g17449(.A1(new_n17626_), .A2(new_n17627_), .B(new_n17618_), .ZN(new_n17642_));
  AOI21_X1   g17450(.A1(new_n17642_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n17643_));
  AOI21_X1   g17451(.A1(new_n17643_), .A2(new_n17636_), .B(new_n17641_), .ZN(new_n17644_));
  OAI21_X1   g17452(.A1(new_n17644_), .A2(new_n17637_), .B(\asqrt[18] ), .ZN(new_n17645_));
  INV_X1     g17453(.I(new_n17645_), .ZN(new_n17646_));
  NAND2_X1   g17454(.A1(new_n17395_), .A2(new_n17393_), .ZN(new_n17647_));
  NAND3_X1   g17455(.A1(\asqrt[11] ), .A2(new_n16989_), .A3(new_n17647_), .ZN(new_n17648_));
  AND3_X2    g17456(.A1(new_n17647_), .A2(new_n16989_), .A3(new_n16994_), .Z(new_n17649_));
  AOI22_X1   g17457(.A1(new_n17648_), .A2(new_n16995_), .B1(\asqrt[11] ), .B2(new_n17649_), .ZN(new_n17650_));
  NOR3_X1    g17458(.A1(new_n17644_), .A2(new_n17637_), .A3(\asqrt[18] ), .ZN(new_n17651_));
  NOR2_X1    g17459(.A1(new_n17651_), .A2(new_n17650_), .ZN(new_n17652_));
  OAI21_X1   g17460(.A1(new_n17652_), .A2(new_n17646_), .B(\asqrt[19] ), .ZN(new_n17653_));
  INV_X1     g17461(.I(new_n17003_), .ZN(new_n17654_));
  NOR3_X1    g17462(.A1(new_n17406_), .A2(new_n16999_), .A3(new_n17654_), .ZN(new_n17655_));
  NOR3_X1    g17463(.A1(new_n17623_), .A2(new_n16999_), .A3(new_n17406_), .ZN(new_n17656_));
  INV_X1     g17464(.I(new_n17656_), .ZN(new_n17657_));
  AOI22_X1   g17465(.A1(new_n17657_), .A2(new_n17654_), .B1(\asqrt[11] ), .B2(new_n17655_), .ZN(new_n17658_));
  INV_X1     g17466(.I(new_n17658_), .ZN(new_n17659_));
  NAND2_X1   g17467(.A1(new_n17645_), .A2(new_n12913_), .ZN(new_n17660_));
  OAI21_X1   g17468(.A1(new_n17652_), .A2(new_n17660_), .B(new_n17659_), .ZN(new_n17661_));
  AOI21_X1   g17469(.A1(new_n17661_), .A2(new_n17653_), .B(new_n12364_), .ZN(new_n17662_));
  NOR3_X1    g17470(.A1(new_n17623_), .A2(new_n17008_), .A3(new_n17013_), .ZN(new_n17663_));
  INV_X1     g17471(.I(new_n17663_), .ZN(new_n17664_));
  NOR3_X1    g17472(.A1(new_n17008_), .A2(new_n17391_), .A3(new_n17013_), .ZN(new_n17665_));
  AOI22_X1   g17473(.A1(new_n17664_), .A2(new_n17391_), .B1(\asqrt[11] ), .B2(new_n17665_), .ZN(new_n17666_));
  OAI21_X1   g17474(.A1(new_n17650_), .A2(new_n17651_), .B(new_n17645_), .ZN(new_n17667_));
  AOI21_X1   g17475(.A1(new_n17667_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n17668_));
  AOI21_X1   g17476(.A1(new_n17668_), .A2(new_n17661_), .B(new_n17666_), .ZN(new_n17669_));
  OAI21_X1   g17477(.A1(new_n17669_), .A2(new_n17662_), .B(\asqrt[21] ), .ZN(new_n17670_));
  INV_X1     g17478(.I(new_n17670_), .ZN(new_n17671_));
  AND3_X2    g17479(.A1(new_n17015_), .A2(new_n17020_), .A3(new_n17400_), .Z(new_n17672_));
  NAND3_X1   g17480(.A1(\asqrt[11] ), .A2(new_n17015_), .A3(new_n17400_), .ZN(new_n17673_));
  AOI22_X1   g17481(.A1(new_n17673_), .A2(new_n17021_), .B1(\asqrt[11] ), .B2(new_n17672_), .ZN(new_n17674_));
  NOR3_X1    g17482(.A1(new_n17669_), .A2(new_n17662_), .A3(\asqrt[21] ), .ZN(new_n17675_));
  NOR2_X1    g17483(.A1(new_n17675_), .A2(new_n17674_), .ZN(new_n17676_));
  OAI21_X1   g17484(.A1(new_n17676_), .A2(new_n17671_), .B(\asqrt[22] ), .ZN(new_n17677_));
  INV_X1     g17485(.I(new_n17028_), .ZN(new_n17678_));
  NOR3_X1    g17486(.A1(new_n17623_), .A2(new_n17024_), .A3(new_n17410_), .ZN(new_n17679_));
  INV_X1     g17487(.I(new_n17679_), .ZN(new_n17680_));
  NOR3_X1    g17488(.A1(new_n17410_), .A2(new_n17024_), .A3(new_n17678_), .ZN(new_n17681_));
  AOI22_X1   g17489(.A1(new_n17680_), .A2(new_n17678_), .B1(\asqrt[11] ), .B2(new_n17681_), .ZN(new_n17682_));
  INV_X1     g17490(.I(new_n17682_), .ZN(new_n17683_));
  NAND2_X1   g17491(.A1(new_n17670_), .A2(new_n11326_), .ZN(new_n17684_));
  OAI21_X1   g17492(.A1(new_n17676_), .A2(new_n17684_), .B(new_n17683_), .ZN(new_n17685_));
  AOI21_X1   g17493(.A1(new_n17685_), .A2(new_n17677_), .B(new_n10812_), .ZN(new_n17686_));
  NOR3_X1    g17494(.A1(new_n17033_), .A2(new_n17390_), .A3(new_n17039_), .ZN(new_n17687_));
  NOR3_X1    g17495(.A1(new_n17623_), .A2(new_n17033_), .A3(new_n17039_), .ZN(new_n17688_));
  INV_X1     g17496(.I(new_n17688_), .ZN(new_n17689_));
  AOI22_X1   g17497(.A1(new_n17689_), .A2(new_n17390_), .B1(\asqrt[11] ), .B2(new_n17687_), .ZN(new_n17690_));
  OAI21_X1   g17498(.A1(new_n17674_), .A2(new_n17675_), .B(new_n17670_), .ZN(new_n17691_));
  AOI21_X1   g17499(.A1(new_n17691_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n17692_));
  AOI21_X1   g17500(.A1(new_n17692_), .A2(new_n17685_), .B(new_n17690_), .ZN(new_n17693_));
  OAI21_X1   g17501(.A1(new_n17693_), .A2(new_n17686_), .B(\asqrt[24] ), .ZN(new_n17694_));
  INV_X1     g17502(.I(new_n17694_), .ZN(new_n17695_));
  NOR2_X1    g17503(.A1(new_n17040_), .A2(new_n17048_), .ZN(new_n17696_));
  NOR3_X1    g17504(.A1(new_n17623_), .A2(new_n17404_), .A3(new_n17696_), .ZN(new_n17697_));
  INV_X1     g17505(.I(new_n17697_), .ZN(new_n17698_));
  NOR3_X1    g17506(.A1(new_n17696_), .A2(new_n17404_), .A3(new_n17047_), .ZN(new_n17699_));
  AOI22_X1   g17507(.A1(new_n17698_), .A2(new_n17047_), .B1(\asqrt[11] ), .B2(new_n17699_), .ZN(new_n17700_));
  NOR3_X1    g17508(.A1(new_n17693_), .A2(new_n17686_), .A3(\asqrt[24] ), .ZN(new_n17701_));
  NOR2_X1    g17509(.A1(new_n17701_), .A2(new_n17700_), .ZN(new_n17702_));
  OAI21_X1   g17510(.A1(new_n17702_), .A2(new_n17695_), .B(\asqrt[25] ), .ZN(new_n17703_));
  INV_X1     g17511(.I(new_n17056_), .ZN(new_n17704_));
  NOR3_X1    g17512(.A1(new_n17418_), .A2(new_n17050_), .A3(new_n17704_), .ZN(new_n17705_));
  NOR3_X1    g17513(.A1(new_n17623_), .A2(new_n17050_), .A3(new_n17418_), .ZN(new_n17706_));
  INV_X1     g17514(.I(new_n17706_), .ZN(new_n17707_));
  AOI22_X1   g17515(.A1(new_n17707_), .A2(new_n17704_), .B1(\asqrt[11] ), .B2(new_n17705_), .ZN(new_n17708_));
  INV_X1     g17516(.I(new_n17708_), .ZN(new_n17709_));
  NAND2_X1   g17517(.A1(new_n17694_), .A2(new_n9846_), .ZN(new_n17710_));
  OAI21_X1   g17518(.A1(new_n17702_), .A2(new_n17710_), .B(new_n17709_), .ZN(new_n17711_));
  AOI21_X1   g17519(.A1(new_n17711_), .A2(new_n17703_), .B(new_n9317_), .ZN(new_n17712_));
  NOR3_X1    g17520(.A1(new_n17623_), .A2(new_n17061_), .A3(new_n17070_), .ZN(new_n17713_));
  INV_X1     g17521(.I(new_n17713_), .ZN(new_n17714_));
  NOR3_X1    g17522(.A1(new_n17061_), .A2(new_n17389_), .A3(new_n17070_), .ZN(new_n17715_));
  AOI22_X1   g17523(.A1(new_n17714_), .A2(new_n17389_), .B1(\asqrt[11] ), .B2(new_n17715_), .ZN(new_n17716_));
  OAI21_X1   g17524(.A1(new_n17700_), .A2(new_n17701_), .B(new_n17694_), .ZN(new_n17717_));
  AOI21_X1   g17525(.A1(new_n17717_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n17718_));
  AOI21_X1   g17526(.A1(new_n17718_), .A2(new_n17711_), .B(new_n17716_), .ZN(new_n17719_));
  OAI21_X1   g17527(.A1(new_n17719_), .A2(new_n17712_), .B(\asqrt[27] ), .ZN(new_n17720_));
  INV_X1     g17528(.I(new_n17720_), .ZN(new_n17721_));
  NOR2_X1    g17529(.A1(new_n17071_), .A2(new_n17079_), .ZN(new_n17722_));
  NOR3_X1    g17530(.A1(new_n17722_), .A2(new_n17417_), .A3(new_n17078_), .ZN(new_n17723_));
  NOR3_X1    g17531(.A1(new_n17623_), .A2(new_n17417_), .A3(new_n17722_), .ZN(new_n17724_));
  INV_X1     g17532(.I(new_n17724_), .ZN(new_n17725_));
  AOI22_X1   g17533(.A1(new_n17725_), .A2(new_n17078_), .B1(\asqrt[11] ), .B2(new_n17723_), .ZN(new_n17726_));
  NOR3_X1    g17534(.A1(new_n17719_), .A2(new_n17712_), .A3(\asqrt[27] ), .ZN(new_n17727_));
  NOR2_X1    g17535(.A1(new_n17727_), .A2(new_n17726_), .ZN(new_n17728_));
  OAI21_X1   g17536(.A1(new_n17728_), .A2(new_n17721_), .B(\asqrt[28] ), .ZN(new_n17729_));
  INV_X1     g17537(.I(new_n17086_), .ZN(new_n17730_));
  NOR3_X1    g17538(.A1(new_n17623_), .A2(new_n17081_), .A3(new_n17426_), .ZN(new_n17731_));
  INV_X1     g17539(.I(new_n17731_), .ZN(new_n17732_));
  NOR3_X1    g17540(.A1(new_n17426_), .A2(new_n17081_), .A3(new_n17730_), .ZN(new_n17733_));
  AOI22_X1   g17541(.A1(new_n17732_), .A2(new_n17730_), .B1(\asqrt[11] ), .B2(new_n17733_), .ZN(new_n17734_));
  INV_X1     g17542(.I(new_n17734_), .ZN(new_n17735_));
  NAND2_X1   g17543(.A1(new_n17720_), .A2(new_n8483_), .ZN(new_n17736_));
  OAI21_X1   g17544(.A1(new_n17728_), .A2(new_n17736_), .B(new_n17735_), .ZN(new_n17737_));
  AOI21_X1   g17545(.A1(new_n17737_), .A2(new_n17729_), .B(new_n8036_), .ZN(new_n17738_));
  NOR3_X1    g17546(.A1(new_n17091_), .A2(new_n17388_), .A3(new_n17100_), .ZN(new_n17739_));
  NOR3_X1    g17547(.A1(new_n17623_), .A2(new_n17091_), .A3(new_n17100_), .ZN(new_n17740_));
  INV_X1     g17548(.I(new_n17740_), .ZN(new_n17741_));
  AOI22_X1   g17549(.A1(new_n17741_), .A2(new_n17388_), .B1(\asqrt[11] ), .B2(new_n17739_), .ZN(new_n17742_));
  OAI21_X1   g17550(.A1(new_n17726_), .A2(new_n17727_), .B(new_n17720_), .ZN(new_n17743_));
  AOI21_X1   g17551(.A1(new_n17743_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n17744_));
  AOI21_X1   g17552(.A1(new_n17744_), .A2(new_n17737_), .B(new_n17742_), .ZN(new_n17745_));
  OAI21_X1   g17553(.A1(new_n17745_), .A2(new_n17738_), .B(\asqrt[30] ), .ZN(new_n17746_));
  INV_X1     g17554(.I(new_n17746_), .ZN(new_n17747_));
  NOR2_X1    g17555(.A1(new_n17101_), .A2(new_n17109_), .ZN(new_n17748_));
  NOR3_X1    g17556(.A1(new_n17623_), .A2(new_n17425_), .A3(new_n17748_), .ZN(new_n17749_));
  INV_X1     g17557(.I(new_n17749_), .ZN(new_n17750_));
  NOR3_X1    g17558(.A1(new_n17748_), .A2(new_n17425_), .A3(new_n17108_), .ZN(new_n17751_));
  AOI22_X1   g17559(.A1(new_n17750_), .A2(new_n17108_), .B1(\asqrt[11] ), .B2(new_n17751_), .ZN(new_n17752_));
  NOR3_X1    g17560(.A1(new_n17745_), .A2(new_n17738_), .A3(\asqrt[30] ), .ZN(new_n17753_));
  NOR2_X1    g17561(.A1(new_n17753_), .A2(new_n17752_), .ZN(new_n17754_));
  OAI21_X1   g17562(.A1(new_n17754_), .A2(new_n17747_), .B(\asqrt[31] ), .ZN(new_n17755_));
  INV_X1     g17563(.I(new_n17116_), .ZN(new_n17756_));
  NOR3_X1    g17564(.A1(new_n17434_), .A2(new_n17111_), .A3(new_n17756_), .ZN(new_n17757_));
  NOR3_X1    g17565(.A1(new_n17623_), .A2(new_n17111_), .A3(new_n17434_), .ZN(new_n17758_));
  INV_X1     g17566(.I(new_n17758_), .ZN(new_n17759_));
  AOI22_X1   g17567(.A1(new_n17759_), .A2(new_n17756_), .B1(\asqrt[11] ), .B2(new_n17757_), .ZN(new_n17760_));
  INV_X1     g17568(.I(new_n17760_), .ZN(new_n17761_));
  NAND2_X1   g17569(.A1(new_n17746_), .A2(new_n7229_), .ZN(new_n17762_));
  OAI21_X1   g17570(.A1(new_n17754_), .A2(new_n17762_), .B(new_n17761_), .ZN(new_n17763_));
  AOI21_X1   g17571(.A1(new_n17763_), .A2(new_n17755_), .B(new_n6824_), .ZN(new_n17764_));
  NOR3_X1    g17572(.A1(new_n17623_), .A2(new_n17121_), .A3(new_n17127_), .ZN(new_n17765_));
  INV_X1     g17573(.I(new_n17765_), .ZN(new_n17766_));
  NOR3_X1    g17574(.A1(new_n17121_), .A2(new_n17387_), .A3(new_n17127_), .ZN(new_n17767_));
  AOI22_X1   g17575(.A1(new_n17766_), .A2(new_n17387_), .B1(\asqrt[11] ), .B2(new_n17767_), .ZN(new_n17768_));
  OAI21_X1   g17576(.A1(new_n17752_), .A2(new_n17753_), .B(new_n17746_), .ZN(new_n17769_));
  AOI21_X1   g17577(.A1(new_n17769_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n17770_));
  AOI21_X1   g17578(.A1(new_n17770_), .A2(new_n17763_), .B(new_n17768_), .ZN(new_n17771_));
  OAI21_X1   g17579(.A1(new_n17771_), .A2(new_n17764_), .B(\asqrt[33] ), .ZN(new_n17772_));
  INV_X1     g17580(.I(new_n17772_), .ZN(new_n17773_));
  NOR2_X1    g17581(.A1(new_n17128_), .A2(new_n17136_), .ZN(new_n17774_));
  NOR3_X1    g17582(.A1(new_n17774_), .A2(new_n17433_), .A3(new_n17135_), .ZN(new_n17775_));
  NOR3_X1    g17583(.A1(new_n17623_), .A2(new_n17433_), .A3(new_n17774_), .ZN(new_n17776_));
  INV_X1     g17584(.I(new_n17776_), .ZN(new_n17777_));
  AOI22_X1   g17585(.A1(new_n17777_), .A2(new_n17135_), .B1(\asqrt[11] ), .B2(new_n17775_), .ZN(new_n17778_));
  NOR3_X1    g17586(.A1(new_n17771_), .A2(new_n17764_), .A3(\asqrt[33] ), .ZN(new_n17779_));
  NOR2_X1    g17587(.A1(new_n17779_), .A2(new_n17778_), .ZN(new_n17780_));
  OAI21_X1   g17588(.A1(new_n17780_), .A2(new_n17773_), .B(\asqrt[34] ), .ZN(new_n17781_));
  INV_X1     g17589(.I(new_n17143_), .ZN(new_n17782_));
  NOR3_X1    g17590(.A1(new_n17623_), .A2(new_n17138_), .A3(new_n17442_), .ZN(new_n17783_));
  INV_X1     g17591(.I(new_n17783_), .ZN(new_n17784_));
  NOR3_X1    g17592(.A1(new_n17442_), .A2(new_n17138_), .A3(new_n17782_), .ZN(new_n17785_));
  AOI22_X1   g17593(.A1(new_n17784_), .A2(new_n17782_), .B1(\asqrt[11] ), .B2(new_n17785_), .ZN(new_n17786_));
  INV_X1     g17594(.I(new_n17786_), .ZN(new_n17787_));
  NAND2_X1   g17595(.A1(new_n17772_), .A2(new_n6077_), .ZN(new_n17788_));
  OAI21_X1   g17596(.A1(new_n17780_), .A2(new_n17788_), .B(new_n17787_), .ZN(new_n17789_));
  AOI21_X1   g17597(.A1(new_n17789_), .A2(new_n17781_), .B(new_n5708_), .ZN(new_n17790_));
  NOR3_X1    g17598(.A1(new_n17148_), .A2(new_n17386_), .A3(new_n17154_), .ZN(new_n17791_));
  NOR3_X1    g17599(.A1(new_n17623_), .A2(new_n17148_), .A3(new_n17154_), .ZN(new_n17792_));
  INV_X1     g17600(.I(new_n17792_), .ZN(new_n17793_));
  AOI22_X1   g17601(.A1(new_n17793_), .A2(new_n17386_), .B1(\asqrt[11] ), .B2(new_n17791_), .ZN(new_n17794_));
  OAI21_X1   g17602(.A1(new_n17778_), .A2(new_n17779_), .B(new_n17772_), .ZN(new_n17795_));
  AOI21_X1   g17603(.A1(new_n17795_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n17796_));
  AOI21_X1   g17604(.A1(new_n17796_), .A2(new_n17789_), .B(new_n17794_), .ZN(new_n17797_));
  OAI21_X1   g17605(.A1(new_n17797_), .A2(new_n17790_), .B(\asqrt[36] ), .ZN(new_n17798_));
  INV_X1     g17606(.I(new_n17798_), .ZN(new_n17799_));
  NOR2_X1    g17607(.A1(new_n17155_), .A2(new_n17163_), .ZN(new_n17800_));
  NOR3_X1    g17608(.A1(new_n17623_), .A2(new_n17441_), .A3(new_n17800_), .ZN(new_n17801_));
  INV_X1     g17609(.I(new_n17801_), .ZN(new_n17802_));
  NOR3_X1    g17610(.A1(new_n17800_), .A2(new_n17441_), .A3(new_n17162_), .ZN(new_n17803_));
  AOI22_X1   g17611(.A1(new_n17802_), .A2(new_n17162_), .B1(\asqrt[11] ), .B2(new_n17803_), .ZN(new_n17804_));
  NOR3_X1    g17612(.A1(new_n17797_), .A2(new_n17790_), .A3(\asqrt[36] ), .ZN(new_n17805_));
  NOR2_X1    g17613(.A1(new_n17805_), .A2(new_n17804_), .ZN(new_n17806_));
  OAI21_X1   g17614(.A1(new_n17806_), .A2(new_n17799_), .B(\asqrt[37] ), .ZN(new_n17807_));
  INV_X1     g17615(.I(new_n17170_), .ZN(new_n17808_));
  NOR3_X1    g17616(.A1(new_n17450_), .A2(new_n17165_), .A3(new_n17808_), .ZN(new_n17809_));
  NOR3_X1    g17617(.A1(new_n17623_), .A2(new_n17165_), .A3(new_n17450_), .ZN(new_n17810_));
  INV_X1     g17618(.I(new_n17810_), .ZN(new_n17811_));
  AOI22_X1   g17619(.A1(new_n17811_), .A2(new_n17808_), .B1(\asqrt[11] ), .B2(new_n17809_), .ZN(new_n17812_));
  INV_X1     g17620(.I(new_n17812_), .ZN(new_n17813_));
  NAND2_X1   g17621(.A1(new_n17798_), .A2(new_n5024_), .ZN(new_n17814_));
  OAI21_X1   g17622(.A1(new_n17806_), .A2(new_n17814_), .B(new_n17813_), .ZN(new_n17815_));
  AOI21_X1   g17623(.A1(new_n17815_), .A2(new_n17807_), .B(new_n4696_), .ZN(new_n17816_));
  NOR3_X1    g17624(.A1(new_n17623_), .A2(new_n17175_), .A3(new_n17181_), .ZN(new_n17817_));
  INV_X1     g17625(.I(new_n17817_), .ZN(new_n17818_));
  NOR3_X1    g17626(.A1(new_n17175_), .A2(new_n17385_), .A3(new_n17181_), .ZN(new_n17819_));
  AOI22_X1   g17627(.A1(new_n17818_), .A2(new_n17385_), .B1(\asqrt[11] ), .B2(new_n17819_), .ZN(new_n17820_));
  OAI21_X1   g17628(.A1(new_n17804_), .A2(new_n17805_), .B(new_n17798_), .ZN(new_n17821_));
  AOI21_X1   g17629(.A1(new_n17821_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n17822_));
  AOI21_X1   g17630(.A1(new_n17822_), .A2(new_n17815_), .B(new_n17820_), .ZN(new_n17823_));
  OAI21_X1   g17631(.A1(new_n17823_), .A2(new_n17816_), .B(\asqrt[39] ), .ZN(new_n17824_));
  INV_X1     g17632(.I(new_n17824_), .ZN(new_n17825_));
  NOR2_X1    g17633(.A1(new_n17182_), .A2(new_n17190_), .ZN(new_n17826_));
  NOR3_X1    g17634(.A1(new_n17826_), .A2(new_n17449_), .A3(new_n17189_), .ZN(new_n17827_));
  NOR3_X1    g17635(.A1(new_n17623_), .A2(new_n17449_), .A3(new_n17826_), .ZN(new_n17828_));
  INV_X1     g17636(.I(new_n17828_), .ZN(new_n17829_));
  AOI22_X1   g17637(.A1(new_n17829_), .A2(new_n17189_), .B1(\asqrt[11] ), .B2(new_n17827_), .ZN(new_n17830_));
  NOR3_X1    g17638(.A1(new_n17823_), .A2(new_n17816_), .A3(\asqrt[39] ), .ZN(new_n17831_));
  NOR2_X1    g17639(.A1(new_n17831_), .A2(new_n17830_), .ZN(new_n17832_));
  OAI21_X1   g17640(.A1(new_n17832_), .A2(new_n17825_), .B(\asqrt[40] ), .ZN(new_n17833_));
  INV_X1     g17641(.I(new_n17196_), .ZN(new_n17834_));
  NOR3_X1    g17642(.A1(new_n17623_), .A2(new_n17192_), .A3(new_n17458_), .ZN(new_n17835_));
  INV_X1     g17643(.I(new_n17835_), .ZN(new_n17836_));
  NOR3_X1    g17644(.A1(new_n17458_), .A2(new_n17192_), .A3(new_n17834_), .ZN(new_n17837_));
  AOI22_X1   g17645(.A1(new_n17836_), .A2(new_n17834_), .B1(\asqrt[11] ), .B2(new_n17837_), .ZN(new_n17838_));
  INV_X1     g17646(.I(new_n17838_), .ZN(new_n17839_));
  NAND2_X1   g17647(.A1(new_n17824_), .A2(new_n4071_), .ZN(new_n17840_));
  OAI21_X1   g17648(.A1(new_n17832_), .A2(new_n17840_), .B(new_n17839_), .ZN(new_n17841_));
  AOI21_X1   g17649(.A1(new_n17841_), .A2(new_n17833_), .B(new_n3782_), .ZN(new_n17842_));
  NOR3_X1    g17650(.A1(new_n17201_), .A2(new_n17384_), .A3(new_n17207_), .ZN(new_n17843_));
  NOR3_X1    g17651(.A1(new_n17623_), .A2(new_n17201_), .A3(new_n17207_), .ZN(new_n17844_));
  INV_X1     g17652(.I(new_n17844_), .ZN(new_n17845_));
  AOI22_X1   g17653(.A1(new_n17845_), .A2(new_n17384_), .B1(\asqrt[11] ), .B2(new_n17843_), .ZN(new_n17846_));
  OAI21_X1   g17654(.A1(new_n17830_), .A2(new_n17831_), .B(new_n17824_), .ZN(new_n17847_));
  AOI21_X1   g17655(.A1(new_n17847_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n17848_));
  AOI21_X1   g17656(.A1(new_n17848_), .A2(new_n17841_), .B(new_n17846_), .ZN(new_n17849_));
  OAI21_X1   g17657(.A1(new_n17849_), .A2(new_n17842_), .B(\asqrt[42] ), .ZN(new_n17850_));
  INV_X1     g17658(.I(new_n17850_), .ZN(new_n17851_));
  NOR2_X1    g17659(.A1(new_n17208_), .A2(new_n17216_), .ZN(new_n17852_));
  NOR3_X1    g17660(.A1(new_n17623_), .A2(new_n17457_), .A3(new_n17852_), .ZN(new_n17853_));
  INV_X1     g17661(.I(new_n17853_), .ZN(new_n17854_));
  NOR3_X1    g17662(.A1(new_n17852_), .A2(new_n17457_), .A3(new_n17215_), .ZN(new_n17855_));
  AOI22_X1   g17663(.A1(new_n17854_), .A2(new_n17215_), .B1(\asqrt[11] ), .B2(new_n17855_), .ZN(new_n17856_));
  NOR3_X1    g17664(.A1(new_n17849_), .A2(new_n17842_), .A3(\asqrt[42] ), .ZN(new_n17857_));
  NOR2_X1    g17665(.A1(new_n17857_), .A2(new_n17856_), .ZN(new_n17858_));
  OAI21_X1   g17666(.A1(new_n17858_), .A2(new_n17851_), .B(\asqrt[43] ), .ZN(new_n17859_));
  INV_X1     g17667(.I(new_n17222_), .ZN(new_n17860_));
  NOR3_X1    g17668(.A1(new_n17466_), .A2(new_n17218_), .A3(new_n17860_), .ZN(new_n17861_));
  NOR3_X1    g17669(.A1(new_n17623_), .A2(new_n17218_), .A3(new_n17466_), .ZN(new_n17862_));
  INV_X1     g17670(.I(new_n17862_), .ZN(new_n17863_));
  AOI22_X1   g17671(.A1(new_n17863_), .A2(new_n17860_), .B1(\asqrt[11] ), .B2(new_n17861_), .ZN(new_n17864_));
  INV_X1     g17672(.I(new_n17864_), .ZN(new_n17865_));
  NAND2_X1   g17673(.A1(new_n17850_), .A2(new_n3218_), .ZN(new_n17866_));
  OAI21_X1   g17674(.A1(new_n17858_), .A2(new_n17866_), .B(new_n17865_), .ZN(new_n17867_));
  AOI21_X1   g17675(.A1(new_n17867_), .A2(new_n17859_), .B(new_n2954_), .ZN(new_n17868_));
  NOR3_X1    g17676(.A1(new_n17623_), .A2(new_n17227_), .A3(new_n17235_), .ZN(new_n17869_));
  INV_X1     g17677(.I(new_n17869_), .ZN(new_n17870_));
  NOR3_X1    g17678(.A1(new_n17227_), .A2(new_n17383_), .A3(new_n17235_), .ZN(new_n17871_));
  AOI22_X1   g17679(.A1(new_n17870_), .A2(new_n17383_), .B1(\asqrt[11] ), .B2(new_n17871_), .ZN(new_n17872_));
  OAI21_X1   g17680(.A1(new_n17856_), .A2(new_n17857_), .B(new_n17850_), .ZN(new_n17873_));
  AOI21_X1   g17681(.A1(new_n17873_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n17874_));
  AOI21_X1   g17682(.A1(new_n17874_), .A2(new_n17867_), .B(new_n17872_), .ZN(new_n17875_));
  OAI21_X1   g17683(.A1(new_n17875_), .A2(new_n17868_), .B(\asqrt[45] ), .ZN(new_n17876_));
  INV_X1     g17684(.I(new_n17876_), .ZN(new_n17877_));
  NOR2_X1    g17685(.A1(new_n17236_), .A2(new_n17243_), .ZN(new_n17878_));
  NOR3_X1    g17686(.A1(new_n17878_), .A2(new_n17465_), .A3(new_n17242_), .ZN(new_n17879_));
  NOR3_X1    g17687(.A1(new_n17623_), .A2(new_n17465_), .A3(new_n17878_), .ZN(new_n17880_));
  INV_X1     g17688(.I(new_n17880_), .ZN(new_n17881_));
  AOI22_X1   g17689(.A1(new_n17881_), .A2(new_n17242_), .B1(\asqrt[11] ), .B2(new_n17879_), .ZN(new_n17882_));
  NOR3_X1    g17690(.A1(new_n17875_), .A2(new_n17868_), .A3(\asqrt[45] ), .ZN(new_n17883_));
  NOR2_X1    g17691(.A1(new_n17883_), .A2(new_n17882_), .ZN(new_n17884_));
  OAI21_X1   g17692(.A1(new_n17884_), .A2(new_n17877_), .B(\asqrt[46] ), .ZN(new_n17885_));
  INV_X1     g17693(.I(new_n17251_), .ZN(new_n17886_));
  NOR3_X1    g17694(.A1(new_n17623_), .A2(new_n17245_), .A3(new_n17474_), .ZN(new_n17887_));
  INV_X1     g17695(.I(new_n17887_), .ZN(new_n17888_));
  NOR3_X1    g17696(.A1(new_n17474_), .A2(new_n17245_), .A3(new_n17886_), .ZN(new_n17889_));
  AOI22_X1   g17697(.A1(new_n17888_), .A2(new_n17886_), .B1(\asqrt[11] ), .B2(new_n17889_), .ZN(new_n17890_));
  INV_X1     g17698(.I(new_n17890_), .ZN(new_n17891_));
  NAND2_X1   g17699(.A1(new_n17876_), .A2(new_n2465_), .ZN(new_n17892_));
  OAI21_X1   g17700(.A1(new_n17884_), .A2(new_n17892_), .B(new_n17891_), .ZN(new_n17893_));
  AOI21_X1   g17701(.A1(new_n17893_), .A2(new_n17885_), .B(new_n2229_), .ZN(new_n17894_));
  NOR3_X1    g17702(.A1(new_n17256_), .A2(new_n17382_), .A3(new_n17265_), .ZN(new_n17895_));
  NOR3_X1    g17703(.A1(new_n17623_), .A2(new_n17256_), .A3(new_n17265_), .ZN(new_n17896_));
  INV_X1     g17704(.I(new_n17896_), .ZN(new_n17897_));
  AOI22_X1   g17705(.A1(new_n17897_), .A2(new_n17382_), .B1(\asqrt[11] ), .B2(new_n17895_), .ZN(new_n17898_));
  OAI21_X1   g17706(.A1(new_n17882_), .A2(new_n17883_), .B(new_n17876_), .ZN(new_n17899_));
  AOI21_X1   g17707(.A1(new_n17899_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n17900_));
  AOI21_X1   g17708(.A1(new_n17900_), .A2(new_n17893_), .B(new_n17898_), .ZN(new_n17901_));
  OAI21_X1   g17709(.A1(new_n17901_), .A2(new_n17894_), .B(\asqrt[48] ), .ZN(new_n17902_));
  INV_X1     g17710(.I(new_n17902_), .ZN(new_n17903_));
  NOR2_X1    g17711(.A1(new_n17266_), .A2(new_n17273_), .ZN(new_n17904_));
  NOR3_X1    g17712(.A1(new_n17623_), .A2(new_n17473_), .A3(new_n17904_), .ZN(new_n17905_));
  INV_X1     g17713(.I(new_n17905_), .ZN(new_n17906_));
  NOR3_X1    g17714(.A1(new_n17904_), .A2(new_n17473_), .A3(new_n17272_), .ZN(new_n17907_));
  AOI22_X1   g17715(.A1(new_n17906_), .A2(new_n17272_), .B1(\asqrt[11] ), .B2(new_n17907_), .ZN(new_n17908_));
  NOR3_X1    g17716(.A1(new_n17901_), .A2(new_n17894_), .A3(\asqrt[48] ), .ZN(new_n17909_));
  NOR2_X1    g17717(.A1(new_n17909_), .A2(new_n17908_), .ZN(new_n17910_));
  OAI21_X1   g17718(.A1(new_n17910_), .A2(new_n17903_), .B(\asqrt[49] ), .ZN(new_n17911_));
  INV_X1     g17719(.I(new_n17281_), .ZN(new_n17912_));
  NOR3_X1    g17720(.A1(new_n17482_), .A2(new_n17275_), .A3(new_n17912_), .ZN(new_n17913_));
  NOR3_X1    g17721(.A1(new_n17623_), .A2(new_n17275_), .A3(new_n17482_), .ZN(new_n17914_));
  INV_X1     g17722(.I(new_n17914_), .ZN(new_n17915_));
  AOI22_X1   g17723(.A1(new_n17915_), .A2(new_n17912_), .B1(\asqrt[11] ), .B2(new_n17913_), .ZN(new_n17916_));
  INV_X1     g17724(.I(new_n17916_), .ZN(new_n17917_));
  NAND2_X1   g17725(.A1(new_n17902_), .A2(new_n1806_), .ZN(new_n17918_));
  OAI21_X1   g17726(.A1(new_n17910_), .A2(new_n17918_), .B(new_n17917_), .ZN(new_n17919_));
  AOI21_X1   g17727(.A1(new_n17919_), .A2(new_n17911_), .B(new_n1612_), .ZN(new_n17920_));
  NOR3_X1    g17728(.A1(new_n17623_), .A2(new_n17286_), .A3(new_n17295_), .ZN(new_n17921_));
  INV_X1     g17729(.I(new_n17921_), .ZN(new_n17922_));
  NOR3_X1    g17730(.A1(new_n17286_), .A2(new_n17381_), .A3(new_n17295_), .ZN(new_n17923_));
  AOI22_X1   g17731(.A1(new_n17922_), .A2(new_n17381_), .B1(\asqrt[11] ), .B2(new_n17923_), .ZN(new_n17924_));
  OAI21_X1   g17732(.A1(new_n17908_), .A2(new_n17909_), .B(new_n17902_), .ZN(new_n17925_));
  AOI21_X1   g17733(.A1(new_n17925_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n17926_));
  AOI21_X1   g17734(.A1(new_n17926_), .A2(new_n17919_), .B(new_n17924_), .ZN(new_n17927_));
  OAI21_X1   g17735(.A1(new_n17927_), .A2(new_n17920_), .B(\asqrt[51] ), .ZN(new_n17928_));
  INV_X1     g17736(.I(new_n17928_), .ZN(new_n17929_));
  NOR2_X1    g17737(.A1(new_n17296_), .A2(new_n17303_), .ZN(new_n17930_));
  NOR3_X1    g17738(.A1(new_n17930_), .A2(new_n17481_), .A3(new_n17302_), .ZN(new_n17931_));
  NOR3_X1    g17739(.A1(new_n17623_), .A2(new_n17481_), .A3(new_n17930_), .ZN(new_n17932_));
  INV_X1     g17740(.I(new_n17932_), .ZN(new_n17933_));
  AOI22_X1   g17741(.A1(new_n17933_), .A2(new_n17302_), .B1(\asqrt[11] ), .B2(new_n17931_), .ZN(new_n17934_));
  NOR3_X1    g17742(.A1(new_n17927_), .A2(new_n17920_), .A3(\asqrt[51] ), .ZN(new_n17935_));
  NOR2_X1    g17743(.A1(new_n17935_), .A2(new_n17934_), .ZN(new_n17936_));
  OAI21_X1   g17744(.A1(new_n17936_), .A2(new_n17929_), .B(\asqrt[52] ), .ZN(new_n17937_));
  INV_X1     g17745(.I(new_n17311_), .ZN(new_n17938_));
  NAND2_X1   g17746(.A1(new_n17313_), .A2(new_n17304_), .ZN(new_n17939_));
  INV_X1     g17747(.I(new_n17939_), .ZN(new_n17940_));
  NOR3_X1    g17748(.A1(new_n17623_), .A2(new_n17305_), .A3(new_n17940_), .ZN(new_n17941_));
  INV_X1     g17749(.I(new_n17941_), .ZN(new_n17942_));
  NOR3_X1    g17750(.A1(new_n17940_), .A2(new_n17305_), .A3(new_n17938_), .ZN(new_n17943_));
  AOI22_X1   g17751(.A1(new_n17942_), .A2(new_n17938_), .B1(\asqrt[11] ), .B2(new_n17943_), .ZN(new_n17944_));
  INV_X1     g17752(.I(new_n17944_), .ZN(new_n17945_));
  NAND2_X1   g17753(.A1(new_n17928_), .A2(new_n1256_), .ZN(new_n17946_));
  OAI21_X1   g17754(.A1(new_n17936_), .A2(new_n17946_), .B(new_n17945_), .ZN(new_n17947_));
  AOI21_X1   g17755(.A1(new_n17947_), .A2(new_n17937_), .B(new_n1103_), .ZN(new_n17948_));
  NOR3_X1    g17756(.A1(new_n17316_), .A2(new_n17380_), .A3(new_n17325_), .ZN(new_n17949_));
  NOR3_X1    g17757(.A1(new_n17623_), .A2(new_n17316_), .A3(new_n17325_), .ZN(new_n17950_));
  INV_X1     g17758(.I(new_n17950_), .ZN(new_n17951_));
  AOI22_X1   g17759(.A1(new_n17951_), .A2(new_n17380_), .B1(\asqrt[11] ), .B2(new_n17949_), .ZN(new_n17952_));
  OAI21_X1   g17760(.A1(new_n17934_), .A2(new_n17935_), .B(new_n17928_), .ZN(new_n17953_));
  AOI21_X1   g17761(.A1(new_n17953_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n17954_));
  AOI21_X1   g17762(.A1(new_n17954_), .A2(new_n17947_), .B(new_n17952_), .ZN(new_n17955_));
  OAI21_X1   g17763(.A1(new_n17955_), .A2(new_n17948_), .B(\asqrt[54] ), .ZN(new_n17956_));
  INV_X1     g17764(.I(new_n17956_), .ZN(new_n17957_));
  INV_X1     g17765(.I(new_n17327_), .ZN(new_n17958_));
  INV_X1     g17766(.I(new_n17489_), .ZN(new_n17959_));
  NOR3_X1    g17767(.A1(new_n17623_), .A2(new_n17958_), .A3(new_n17959_), .ZN(new_n17960_));
  INV_X1     g17768(.I(new_n17960_), .ZN(new_n17961_));
  NOR3_X1    g17769(.A1(new_n17958_), .A2(new_n17959_), .A3(new_n17332_), .ZN(new_n17962_));
  AOI22_X1   g17770(.A1(new_n17961_), .A2(new_n17332_), .B1(\asqrt[11] ), .B2(new_n17962_), .ZN(new_n17963_));
  NOR3_X1    g17771(.A1(new_n17955_), .A2(new_n17948_), .A3(\asqrt[54] ), .ZN(new_n17964_));
  NOR2_X1    g17772(.A1(new_n17964_), .A2(new_n17963_), .ZN(new_n17965_));
  OAI21_X1   g17773(.A1(new_n17965_), .A2(new_n17957_), .B(\asqrt[55] ), .ZN(new_n17966_));
  INV_X1     g17774(.I(new_n17341_), .ZN(new_n17967_));
  INV_X1     g17775(.I(new_n17334_), .ZN(new_n17968_));
  INV_X1     g17776(.I(new_n17343_), .ZN(new_n17969_));
  OAI21_X1   g17777(.A1(new_n17969_), .A2(new_n17968_), .B(new_n17341_), .ZN(new_n17970_));
  NOR2_X1    g17778(.A1(new_n17970_), .A2(new_n17335_), .ZN(new_n17971_));
  NOR2_X1    g17779(.A1(new_n17969_), .A2(new_n17968_), .ZN(new_n17972_));
  NOR3_X1    g17780(.A1(new_n17623_), .A2(new_n17335_), .A3(new_n17972_), .ZN(new_n17973_));
  INV_X1     g17781(.I(new_n17973_), .ZN(new_n17974_));
  AOI22_X1   g17782(.A1(new_n17974_), .A2(new_n17967_), .B1(\asqrt[11] ), .B2(new_n17971_), .ZN(new_n17975_));
  INV_X1     g17783(.I(new_n17975_), .ZN(new_n17976_));
  NAND2_X1   g17784(.A1(new_n17956_), .A2(new_n823_), .ZN(new_n17977_));
  OAI21_X1   g17785(.A1(new_n17965_), .A2(new_n17977_), .B(new_n17976_), .ZN(new_n17978_));
  AOI21_X1   g17786(.A1(new_n17978_), .A2(new_n17966_), .B(new_n703_), .ZN(new_n17979_));
  NOR3_X1    g17787(.A1(new_n17623_), .A2(new_n17346_), .A3(new_n17352_), .ZN(new_n17980_));
  INV_X1     g17788(.I(new_n17980_), .ZN(new_n17981_));
  NOR3_X1    g17789(.A1(new_n17346_), .A2(new_n17379_), .A3(new_n17352_), .ZN(new_n17982_));
  AOI22_X1   g17790(.A1(new_n17981_), .A2(new_n17379_), .B1(\asqrt[11] ), .B2(new_n17982_), .ZN(new_n17983_));
  OAI21_X1   g17791(.A1(new_n17963_), .A2(new_n17964_), .B(new_n17956_), .ZN(new_n17984_));
  AOI21_X1   g17792(.A1(new_n17984_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n17985_));
  AOI21_X1   g17793(.A1(new_n17985_), .A2(new_n17978_), .B(new_n17983_), .ZN(new_n17986_));
  OAI21_X1   g17794(.A1(new_n17986_), .A2(new_n17979_), .B(\asqrt[57] ), .ZN(new_n17987_));
  INV_X1     g17795(.I(new_n17987_), .ZN(new_n17988_));
  INV_X1     g17796(.I(new_n17354_), .ZN(new_n17989_));
  INV_X1     g17797(.I(new_n17493_), .ZN(new_n17990_));
  NOR3_X1    g17798(.A1(new_n17989_), .A2(new_n17990_), .A3(new_n17359_), .ZN(new_n17991_));
  NOR3_X1    g17799(.A1(new_n17623_), .A2(new_n17989_), .A3(new_n17990_), .ZN(new_n17992_));
  INV_X1     g17800(.I(new_n17992_), .ZN(new_n17993_));
  AOI22_X1   g17801(.A1(new_n17993_), .A2(new_n17359_), .B1(\asqrt[11] ), .B2(new_n17991_), .ZN(new_n17994_));
  NOR3_X1    g17802(.A1(new_n17986_), .A2(new_n17979_), .A3(\asqrt[57] ), .ZN(new_n17995_));
  NOR2_X1    g17803(.A1(new_n17995_), .A2(new_n17994_), .ZN(new_n17996_));
  OAI21_X1   g17804(.A1(new_n17996_), .A2(new_n17988_), .B(\asqrt[58] ), .ZN(new_n17997_));
  INV_X1     g17805(.I(new_n17368_), .ZN(new_n17998_));
  INV_X1     g17806(.I(new_n17361_), .ZN(new_n17999_));
  INV_X1     g17807(.I(new_n17370_), .ZN(new_n18000_));
  NOR2_X1    g17808(.A1(new_n18000_), .A2(new_n17999_), .ZN(new_n18001_));
  NOR3_X1    g17809(.A1(new_n17623_), .A2(new_n17362_), .A3(new_n18001_), .ZN(new_n18002_));
  INV_X1     g17810(.I(new_n18002_), .ZN(new_n18003_));
  NOR3_X1    g17811(.A1(new_n18001_), .A2(new_n17362_), .A3(new_n17998_), .ZN(new_n18004_));
  AOI22_X1   g17812(.A1(new_n18003_), .A2(new_n17998_), .B1(\asqrt[11] ), .B2(new_n18004_), .ZN(new_n18005_));
  INV_X1     g17813(.I(new_n18005_), .ZN(new_n18006_));
  NAND2_X1   g17814(.A1(new_n17987_), .A2(new_n436_), .ZN(new_n18007_));
  OAI21_X1   g17815(.A1(new_n17996_), .A2(new_n18007_), .B(new_n18006_), .ZN(new_n18008_));
  AOI21_X1   g17816(.A1(new_n18008_), .A2(new_n17997_), .B(new_n327_), .ZN(new_n18009_));
  NOR3_X1    g17817(.A1(new_n17513_), .A2(new_n17378_), .A3(new_n17514_), .ZN(new_n18010_));
  NOR3_X1    g17818(.A1(new_n17623_), .A2(new_n17513_), .A3(new_n17514_), .ZN(new_n18011_));
  INV_X1     g17819(.I(new_n18011_), .ZN(new_n18012_));
  AOI22_X1   g17820(.A1(new_n18012_), .A2(new_n17378_), .B1(\asqrt[11] ), .B2(new_n18010_), .ZN(new_n18013_));
  OAI21_X1   g17821(.A1(new_n17994_), .A2(new_n17995_), .B(new_n17987_), .ZN(new_n18014_));
  AOI21_X1   g17822(.A1(new_n18014_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n18015_));
  AOI21_X1   g17823(.A1(new_n18015_), .A2(new_n18008_), .B(new_n18013_), .ZN(new_n18016_));
  OAI21_X1   g17824(.A1(new_n18016_), .A2(new_n18009_), .B(\asqrt[60] ), .ZN(new_n18017_));
  INV_X1     g17825(.I(new_n18017_), .ZN(new_n18018_));
  INV_X1     g17826(.I(new_n17572_), .ZN(new_n18019_));
  NOR3_X1    g17827(.A1(new_n17623_), .A2(new_n17497_), .A3(new_n18019_), .ZN(new_n18020_));
  INV_X1     g17828(.I(new_n18020_), .ZN(new_n18021_));
  NOR3_X1    g17829(.A1(new_n18019_), .A2(new_n17497_), .A3(new_n17525_), .ZN(new_n18022_));
  AOI22_X1   g17830(.A1(new_n18021_), .A2(new_n17525_), .B1(\asqrt[11] ), .B2(new_n18022_), .ZN(new_n18023_));
  NOR3_X1    g17831(.A1(new_n18016_), .A2(new_n18009_), .A3(\asqrt[60] ), .ZN(new_n18024_));
  NOR2_X1    g17832(.A1(new_n18024_), .A2(new_n18023_), .ZN(new_n18025_));
  OAI21_X1   g17833(.A1(new_n18025_), .A2(new_n18018_), .B(\asqrt[61] ), .ZN(new_n18026_));
  NAND2_X1   g17834(.A1(new_n17537_), .A2(new_n17526_), .ZN(new_n18027_));
  AND3_X2    g17835(.A1(new_n17505_), .A2(new_n17511_), .A3(new_n18027_), .Z(new_n18028_));
  NAND3_X1   g17836(.A1(\asqrt[11] ), .A2(new_n17505_), .A3(new_n18027_), .ZN(new_n18029_));
  AOI22_X1   g17837(.A1(new_n18029_), .A2(new_n17512_), .B1(\asqrt[11] ), .B2(new_n18028_), .ZN(new_n18030_));
  INV_X1     g17838(.I(new_n18030_), .ZN(new_n18031_));
  NAND2_X1   g17839(.A1(new_n18017_), .A2(new_n218_), .ZN(new_n18032_));
  OAI21_X1   g17840(.A1(new_n18025_), .A2(new_n18032_), .B(new_n18031_), .ZN(new_n18033_));
  AOI21_X1   g17841(.A1(new_n18033_), .A2(new_n18026_), .B(new_n207_), .ZN(new_n18034_));
  NOR3_X1    g17842(.A1(new_n17623_), .A2(new_n17519_), .A3(new_n17550_), .ZN(new_n18035_));
  INV_X1     g17843(.I(new_n18035_), .ZN(new_n18036_));
  NOR3_X1    g17844(.A1(new_n17519_), .A2(new_n17571_), .A3(new_n17550_), .ZN(new_n18037_));
  AOI22_X1   g17845(.A1(new_n18036_), .A2(new_n17571_), .B1(\asqrt[11] ), .B2(new_n18037_), .ZN(new_n18038_));
  OAI21_X1   g17846(.A1(new_n18023_), .A2(new_n18024_), .B(new_n18017_), .ZN(new_n18039_));
  AOI21_X1   g17847(.A1(new_n18039_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n18040_));
  AOI21_X1   g17848(.A1(new_n18040_), .A2(new_n18033_), .B(new_n18038_), .ZN(new_n18041_));
  INV_X1     g17849(.I(new_n17530_), .ZN(new_n18042_));
  INV_X1     g17850(.I(new_n17584_), .ZN(new_n18043_));
  NOR3_X1    g17851(.A1(new_n18042_), .A2(new_n18043_), .A3(new_n17535_), .ZN(new_n18044_));
  NAND2_X1   g17852(.A1(\asqrt[11] ), .A2(new_n18044_), .ZN(new_n18045_));
  INV_X1     g17853(.I(new_n18045_), .ZN(new_n18046_));
  NOR2_X1    g17854(.A1(new_n18042_), .A2(new_n18043_), .ZN(new_n18047_));
  AOI21_X1   g17855(.A1(\asqrt[11] ), .A2(new_n18047_), .B(new_n17534_), .ZN(new_n18048_));
  NOR2_X1    g17856(.A1(new_n18046_), .A2(new_n18048_), .ZN(new_n18049_));
  INV_X1     g17857(.I(new_n18049_), .ZN(new_n18050_));
  NAND3_X1   g17858(.A1(\asqrt[11] ), .A2(new_n17568_), .A3(new_n17545_), .ZN(new_n18051_));
  AND3_X2    g17859(.A1(new_n18050_), .A2(new_n17598_), .A3(new_n18051_), .Z(new_n18052_));
  OAI21_X1   g17860(.A1(new_n18041_), .A2(new_n18034_), .B(new_n18052_), .ZN(new_n18053_));
  NAND2_X1   g17861(.A1(new_n18053_), .A2(new_n193_), .ZN(new_n18054_));
  INV_X1     g17862(.I(new_n18023_), .ZN(new_n18055_));
  INV_X1     g17863(.I(new_n17994_), .ZN(new_n18056_));
  INV_X1     g17864(.I(new_n17963_), .ZN(new_n18057_));
  INV_X1     g17865(.I(new_n17934_), .ZN(new_n18058_));
  INV_X1     g17866(.I(new_n17908_), .ZN(new_n18059_));
  INV_X1     g17867(.I(new_n17882_), .ZN(new_n18060_));
  INV_X1     g17868(.I(new_n17856_), .ZN(new_n18061_));
  INV_X1     g17869(.I(new_n17830_), .ZN(new_n18062_));
  INV_X1     g17870(.I(new_n17804_), .ZN(new_n18063_));
  INV_X1     g17871(.I(new_n17778_), .ZN(new_n18064_));
  INV_X1     g17872(.I(new_n17752_), .ZN(new_n18065_));
  INV_X1     g17873(.I(new_n17726_), .ZN(new_n18066_));
  INV_X1     g17874(.I(new_n17700_), .ZN(new_n18067_));
  INV_X1     g17875(.I(new_n17674_), .ZN(new_n18068_));
  INV_X1     g17876(.I(new_n17650_), .ZN(new_n18069_));
  NAND2_X1   g17877(.A1(new_n17581_), .A2(new_n17589_), .ZN(new_n18070_));
  OAI21_X1   g17878(.A1(new_n17570_), .A2(new_n17580_), .B(new_n17583_), .ZN(new_n18071_));
  NAND2_X1   g17879(.A1(new_n18071_), .A2(\a[23] ), .ZN(new_n18072_));
  NAND3_X1   g17880(.A1(new_n18070_), .A2(new_n18072_), .A3(new_n17597_), .ZN(new_n18073_));
  AOI21_X1   g17881(.A1(new_n18073_), .A2(new_n17612_), .B(new_n16389_), .ZN(new_n18074_));
  OAI21_X1   g17882(.A1(new_n17603_), .A2(new_n17592_), .B(\a[24] ), .ZN(new_n18075_));
  NAND3_X1   g17883(.A1(new_n17600_), .A2(new_n17597_), .A3(new_n16882_), .ZN(new_n18076_));
  NAND2_X1   g17884(.A1(new_n17581_), .A2(new_n17567_), .ZN(new_n18077_));
  AOI21_X1   g17885(.A1(new_n18077_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n18078_));
  AOI22_X1   g17886(.A1(new_n18073_), .A2(new_n18078_), .B1(new_n18075_), .B2(new_n18076_), .ZN(new_n18079_));
  OAI21_X1   g17887(.A1(new_n18079_), .A2(new_n18074_), .B(\asqrt[14] ), .ZN(new_n18080_));
  NAND2_X1   g17888(.A1(new_n18080_), .A2(new_n15067_), .ZN(new_n18081_));
  OAI21_X1   g17889(.A1(new_n18081_), .A2(new_n17617_), .B(new_n17625_), .ZN(new_n18082_));
  AOI21_X1   g17890(.A1(new_n18082_), .A2(new_n17618_), .B(new_n14601_), .ZN(new_n18083_));
  INV_X1     g17891(.I(new_n17611_), .ZN(new_n18084_));
  AOI21_X1   g17892(.A1(\a[23] ), .A2(new_n18071_), .B(new_n17592_), .ZN(new_n18085_));
  AOI21_X1   g17893(.A1(new_n18085_), .A2(new_n18070_), .B(new_n17582_), .ZN(new_n18086_));
  OAI21_X1   g17894(.A1(new_n18086_), .A2(new_n16389_), .B(new_n15770_), .ZN(new_n18087_));
  OAI21_X1   g17895(.A1(new_n18087_), .A2(new_n18079_), .B(new_n18084_), .ZN(new_n18088_));
  NAND2_X1   g17896(.A1(new_n18088_), .A2(new_n18080_), .ZN(new_n18089_));
  AOI21_X1   g17897(.A1(new_n18089_), .A2(\asqrt[15] ), .B(\asqrt[16] ), .ZN(new_n18090_));
  AOI21_X1   g17898(.A1(new_n18090_), .A2(new_n18082_), .B(new_n17633_), .ZN(new_n18091_));
  OAI21_X1   g17899(.A1(new_n18091_), .A2(new_n18083_), .B(\asqrt[17] ), .ZN(new_n18092_));
  NAND2_X1   g17900(.A1(new_n18092_), .A2(new_n13353_), .ZN(new_n18093_));
  OAI21_X1   g17901(.A1(new_n18093_), .A2(new_n17644_), .B(new_n18069_), .ZN(new_n18094_));
  NAND3_X1   g17902(.A1(new_n18094_), .A2(new_n12913_), .A3(new_n17645_), .ZN(new_n18095_));
  AOI22_X1   g17903(.A1(new_n18095_), .A2(new_n17659_), .B1(new_n17667_), .B2(\asqrt[19] ), .ZN(new_n18096_));
  OAI21_X1   g17904(.A1(new_n18096_), .A2(new_n12364_), .B(new_n11736_), .ZN(new_n18097_));
  OAI21_X1   g17905(.A1(new_n18097_), .A2(new_n17669_), .B(new_n18068_), .ZN(new_n18098_));
  AOI21_X1   g17906(.A1(new_n18098_), .A2(new_n17670_), .B(new_n11326_), .ZN(new_n18099_));
  AOI21_X1   g17907(.A1(new_n18094_), .A2(new_n17645_), .B(new_n12913_), .ZN(new_n18100_));
  NOR3_X1    g17908(.A1(new_n18091_), .A2(new_n18083_), .A3(\asqrt[17] ), .ZN(new_n18101_));
  OAI21_X1   g17909(.A1(new_n17641_), .A2(new_n18101_), .B(new_n18092_), .ZN(new_n18102_));
  AOI21_X1   g17910(.A1(new_n18102_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n18103_));
  AOI21_X1   g17911(.A1(new_n18103_), .A2(new_n18094_), .B(new_n17658_), .ZN(new_n18104_));
  NOR3_X1    g17912(.A1(new_n18104_), .A2(\asqrt[20] ), .A3(new_n18100_), .ZN(new_n18105_));
  OAI22_X1   g17913(.A1(new_n18105_), .A2(new_n17666_), .B1(new_n18096_), .B2(new_n12364_), .ZN(new_n18106_));
  AOI21_X1   g17914(.A1(new_n18106_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n18107_));
  AOI21_X1   g17915(.A1(new_n18107_), .A2(new_n18098_), .B(new_n17682_), .ZN(new_n18108_));
  OAI21_X1   g17916(.A1(new_n18108_), .A2(new_n18099_), .B(\asqrt[23] ), .ZN(new_n18109_));
  NAND2_X1   g17917(.A1(new_n18109_), .A2(new_n10221_), .ZN(new_n18110_));
  OAI21_X1   g17918(.A1(new_n18110_), .A2(new_n17693_), .B(new_n18067_), .ZN(new_n18111_));
  AOI21_X1   g17919(.A1(new_n18111_), .A2(new_n17694_), .B(new_n9846_), .ZN(new_n18112_));
  NOR3_X1    g17920(.A1(new_n18108_), .A2(\asqrt[23] ), .A3(new_n18099_), .ZN(new_n18113_));
  OAI21_X1   g17921(.A1(new_n17690_), .A2(new_n18113_), .B(new_n18109_), .ZN(new_n18114_));
  AOI21_X1   g17922(.A1(new_n18114_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n18115_));
  AOI21_X1   g17923(.A1(new_n18115_), .A2(new_n18111_), .B(new_n17708_), .ZN(new_n18116_));
  OAI21_X1   g17924(.A1(new_n18116_), .A2(new_n18112_), .B(\asqrt[26] ), .ZN(new_n18117_));
  NAND2_X1   g17925(.A1(new_n18117_), .A2(new_n8826_), .ZN(new_n18118_));
  OAI21_X1   g17926(.A1(new_n18118_), .A2(new_n17719_), .B(new_n18066_), .ZN(new_n18119_));
  AOI21_X1   g17927(.A1(new_n18119_), .A2(new_n17720_), .B(new_n8483_), .ZN(new_n18120_));
  NOR3_X1    g17928(.A1(new_n18116_), .A2(\asqrt[26] ), .A3(new_n18112_), .ZN(new_n18121_));
  OAI21_X1   g17929(.A1(new_n17716_), .A2(new_n18121_), .B(new_n18117_), .ZN(new_n18122_));
  AOI21_X1   g17930(.A1(new_n18122_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n18123_));
  AOI21_X1   g17931(.A1(new_n18123_), .A2(new_n18119_), .B(new_n17734_), .ZN(new_n18124_));
  OAI21_X1   g17932(.A1(new_n18124_), .A2(new_n18120_), .B(\asqrt[29] ), .ZN(new_n18125_));
  NAND2_X1   g17933(.A1(new_n18125_), .A2(new_n7539_), .ZN(new_n18126_));
  OAI21_X1   g17934(.A1(new_n18126_), .A2(new_n17745_), .B(new_n18065_), .ZN(new_n18127_));
  AOI21_X1   g17935(.A1(new_n18127_), .A2(new_n17746_), .B(new_n7229_), .ZN(new_n18128_));
  NOR3_X1    g17936(.A1(new_n18124_), .A2(\asqrt[29] ), .A3(new_n18120_), .ZN(new_n18129_));
  OAI21_X1   g17937(.A1(new_n17742_), .A2(new_n18129_), .B(new_n18125_), .ZN(new_n18130_));
  AOI21_X1   g17938(.A1(new_n18130_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n18131_));
  AOI21_X1   g17939(.A1(new_n18131_), .A2(new_n18127_), .B(new_n17760_), .ZN(new_n18132_));
  OAI21_X1   g17940(.A1(new_n18132_), .A2(new_n18128_), .B(\asqrt[32] ), .ZN(new_n18133_));
  NAND2_X1   g17941(.A1(new_n18133_), .A2(new_n6356_), .ZN(new_n18134_));
  OAI21_X1   g17942(.A1(new_n18134_), .A2(new_n17771_), .B(new_n18064_), .ZN(new_n18135_));
  AOI21_X1   g17943(.A1(new_n18135_), .A2(new_n17772_), .B(new_n6077_), .ZN(new_n18136_));
  NOR3_X1    g17944(.A1(new_n18132_), .A2(\asqrt[32] ), .A3(new_n18128_), .ZN(new_n18137_));
  OAI21_X1   g17945(.A1(new_n17768_), .A2(new_n18137_), .B(new_n18133_), .ZN(new_n18138_));
  AOI21_X1   g17946(.A1(new_n18138_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n18139_));
  AOI21_X1   g17947(.A1(new_n18139_), .A2(new_n18135_), .B(new_n17786_), .ZN(new_n18140_));
  OAI21_X1   g17948(.A1(new_n18140_), .A2(new_n18136_), .B(\asqrt[35] ), .ZN(new_n18141_));
  NAND2_X1   g17949(.A1(new_n18141_), .A2(new_n5277_), .ZN(new_n18142_));
  OAI21_X1   g17950(.A1(new_n18142_), .A2(new_n17797_), .B(new_n18063_), .ZN(new_n18143_));
  AOI21_X1   g17951(.A1(new_n18143_), .A2(new_n17798_), .B(new_n5024_), .ZN(new_n18144_));
  NOR3_X1    g17952(.A1(new_n18140_), .A2(\asqrt[35] ), .A3(new_n18136_), .ZN(new_n18145_));
  OAI21_X1   g17953(.A1(new_n17794_), .A2(new_n18145_), .B(new_n18141_), .ZN(new_n18146_));
  AOI21_X1   g17954(.A1(new_n18146_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n18147_));
  AOI21_X1   g17955(.A1(new_n18147_), .A2(new_n18143_), .B(new_n17812_), .ZN(new_n18148_));
  OAI21_X1   g17956(.A1(new_n18148_), .A2(new_n18144_), .B(\asqrt[38] ), .ZN(new_n18149_));
  NAND2_X1   g17957(.A1(new_n18149_), .A2(new_n4298_), .ZN(new_n18150_));
  OAI21_X1   g17958(.A1(new_n18150_), .A2(new_n17823_), .B(new_n18062_), .ZN(new_n18151_));
  AOI21_X1   g17959(.A1(new_n18151_), .A2(new_n17824_), .B(new_n4071_), .ZN(new_n18152_));
  NOR3_X1    g17960(.A1(new_n18148_), .A2(\asqrt[38] ), .A3(new_n18144_), .ZN(new_n18153_));
  OAI21_X1   g17961(.A1(new_n17820_), .A2(new_n18153_), .B(new_n18149_), .ZN(new_n18154_));
  AOI21_X1   g17962(.A1(new_n18154_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n18155_));
  AOI21_X1   g17963(.A1(new_n18155_), .A2(new_n18151_), .B(new_n17838_), .ZN(new_n18156_));
  OAI21_X1   g17964(.A1(new_n18156_), .A2(new_n18152_), .B(\asqrt[41] ), .ZN(new_n18157_));
  NAND2_X1   g17965(.A1(new_n18157_), .A2(new_n3419_), .ZN(new_n18158_));
  OAI21_X1   g17966(.A1(new_n18158_), .A2(new_n17849_), .B(new_n18061_), .ZN(new_n18159_));
  AOI21_X1   g17967(.A1(new_n18159_), .A2(new_n17850_), .B(new_n3218_), .ZN(new_n18160_));
  NOR3_X1    g17968(.A1(new_n18156_), .A2(\asqrt[41] ), .A3(new_n18152_), .ZN(new_n18161_));
  OAI21_X1   g17969(.A1(new_n17846_), .A2(new_n18161_), .B(new_n18157_), .ZN(new_n18162_));
  AOI21_X1   g17970(.A1(new_n18162_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n18163_));
  AOI21_X1   g17971(.A1(new_n18163_), .A2(new_n18159_), .B(new_n17864_), .ZN(new_n18164_));
  OAI21_X1   g17972(.A1(new_n18164_), .A2(new_n18160_), .B(\asqrt[44] ), .ZN(new_n18165_));
  NAND2_X1   g17973(.A1(new_n18165_), .A2(new_n2641_), .ZN(new_n18166_));
  OAI21_X1   g17974(.A1(new_n18166_), .A2(new_n17875_), .B(new_n18060_), .ZN(new_n18167_));
  AOI21_X1   g17975(.A1(new_n18167_), .A2(new_n17876_), .B(new_n2465_), .ZN(new_n18168_));
  NOR3_X1    g17976(.A1(new_n18164_), .A2(\asqrt[44] ), .A3(new_n18160_), .ZN(new_n18169_));
  OAI21_X1   g17977(.A1(new_n17872_), .A2(new_n18169_), .B(new_n18165_), .ZN(new_n18170_));
  AOI21_X1   g17978(.A1(new_n18170_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n18171_));
  AOI21_X1   g17979(.A1(new_n18171_), .A2(new_n18167_), .B(new_n17890_), .ZN(new_n18172_));
  OAI21_X1   g17980(.A1(new_n18172_), .A2(new_n18168_), .B(\asqrt[47] ), .ZN(new_n18173_));
  NAND2_X1   g17981(.A1(new_n18173_), .A2(new_n1956_), .ZN(new_n18174_));
  OAI21_X1   g17982(.A1(new_n18174_), .A2(new_n17901_), .B(new_n18059_), .ZN(new_n18175_));
  AOI21_X1   g17983(.A1(new_n18175_), .A2(new_n17902_), .B(new_n1806_), .ZN(new_n18176_));
  NOR3_X1    g17984(.A1(new_n18172_), .A2(\asqrt[47] ), .A3(new_n18168_), .ZN(new_n18177_));
  OAI21_X1   g17985(.A1(new_n17898_), .A2(new_n18177_), .B(new_n18173_), .ZN(new_n18178_));
  AOI21_X1   g17986(.A1(new_n18178_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n18179_));
  AOI21_X1   g17987(.A1(new_n18179_), .A2(new_n18175_), .B(new_n17916_), .ZN(new_n18180_));
  OAI21_X1   g17988(.A1(new_n18180_), .A2(new_n18176_), .B(\asqrt[50] ), .ZN(new_n18181_));
  NAND2_X1   g17989(.A1(new_n18181_), .A2(new_n1376_), .ZN(new_n18182_));
  OAI21_X1   g17990(.A1(new_n18182_), .A2(new_n17927_), .B(new_n18058_), .ZN(new_n18183_));
  AOI21_X1   g17991(.A1(new_n18183_), .A2(new_n17928_), .B(new_n1256_), .ZN(new_n18184_));
  NOR3_X1    g17992(.A1(new_n18180_), .A2(\asqrt[50] ), .A3(new_n18176_), .ZN(new_n18185_));
  OAI21_X1   g17993(.A1(new_n17924_), .A2(new_n18185_), .B(new_n18181_), .ZN(new_n18186_));
  AOI21_X1   g17994(.A1(new_n18186_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n18187_));
  AOI21_X1   g17995(.A1(new_n18187_), .A2(new_n18183_), .B(new_n17944_), .ZN(new_n18188_));
  OAI21_X1   g17996(.A1(new_n18188_), .A2(new_n18184_), .B(\asqrt[53] ), .ZN(new_n18189_));
  NAND2_X1   g17997(.A1(new_n18189_), .A2(new_n904_), .ZN(new_n18190_));
  OAI21_X1   g17998(.A1(new_n18190_), .A2(new_n17955_), .B(new_n18057_), .ZN(new_n18191_));
  AOI21_X1   g17999(.A1(new_n18191_), .A2(new_n17956_), .B(new_n823_), .ZN(new_n18192_));
  NOR3_X1    g18000(.A1(new_n18188_), .A2(\asqrt[53] ), .A3(new_n18184_), .ZN(new_n18193_));
  OAI21_X1   g18001(.A1(new_n17952_), .A2(new_n18193_), .B(new_n18189_), .ZN(new_n18194_));
  AOI21_X1   g18002(.A1(new_n18194_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n18195_));
  AOI21_X1   g18003(.A1(new_n18195_), .A2(new_n18191_), .B(new_n17975_), .ZN(new_n18196_));
  OAI21_X1   g18004(.A1(new_n18196_), .A2(new_n18192_), .B(\asqrt[56] ), .ZN(new_n18197_));
  NAND2_X1   g18005(.A1(new_n18197_), .A2(new_n531_), .ZN(new_n18198_));
  OAI21_X1   g18006(.A1(new_n18198_), .A2(new_n17986_), .B(new_n18056_), .ZN(new_n18199_));
  AOI21_X1   g18007(.A1(new_n18199_), .A2(new_n17987_), .B(new_n436_), .ZN(new_n18200_));
  NOR3_X1    g18008(.A1(new_n18196_), .A2(\asqrt[56] ), .A3(new_n18192_), .ZN(new_n18201_));
  OAI21_X1   g18009(.A1(new_n17983_), .A2(new_n18201_), .B(new_n18197_), .ZN(new_n18202_));
  AOI21_X1   g18010(.A1(new_n18202_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n18203_));
  AOI21_X1   g18011(.A1(new_n18203_), .A2(new_n18199_), .B(new_n18005_), .ZN(new_n18204_));
  OAI21_X1   g18012(.A1(new_n18204_), .A2(new_n18200_), .B(\asqrt[59] ), .ZN(new_n18205_));
  NAND2_X1   g18013(.A1(new_n18205_), .A2(new_n306_), .ZN(new_n18206_));
  OAI21_X1   g18014(.A1(new_n18206_), .A2(new_n18016_), .B(new_n18055_), .ZN(new_n18207_));
  NOR3_X1    g18015(.A1(new_n18204_), .A2(\asqrt[59] ), .A3(new_n18200_), .ZN(new_n18208_));
  OAI21_X1   g18016(.A1(new_n18013_), .A2(new_n18208_), .B(new_n18205_), .ZN(new_n18209_));
  AOI21_X1   g18017(.A1(new_n18209_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n18210_));
  AOI21_X1   g18018(.A1(new_n18210_), .A2(new_n18207_), .B(new_n18030_), .ZN(new_n18211_));
  INV_X1     g18019(.I(new_n18038_), .ZN(new_n18212_));
  NAND2_X1   g18020(.A1(new_n18026_), .A2(new_n207_), .ZN(new_n18213_));
  OAI21_X1   g18021(.A1(new_n18213_), .A2(new_n18211_), .B(new_n18212_), .ZN(new_n18214_));
  NOR2_X1    g18022(.A1(new_n18034_), .A2(new_n18050_), .ZN(new_n18215_));
  NAND2_X1   g18023(.A1(\asqrt[11] ), .A2(new_n17545_), .ZN(new_n18216_));
  OAI21_X1   g18024(.A1(new_n17585_), .A2(new_n17578_), .B(\asqrt[63] ), .ZN(new_n18217_));
  AOI21_X1   g18025(.A1(new_n18216_), .A2(new_n17585_), .B(new_n18217_), .ZN(new_n18218_));
  AND2_X2    g18026(.A1(new_n17542_), .A2(new_n17558_), .Z(new_n18219_));
  NAND4_X1   g18027(.A1(new_n17598_), .A2(new_n17544_), .A3(new_n17555_), .A4(new_n18219_), .ZN(new_n18220_));
  NOR2_X1    g18028(.A1(new_n18220_), .A2(new_n17570_), .ZN(new_n18221_));
  NOR2_X1    g18029(.A1(new_n18218_), .A2(new_n18221_), .ZN(new_n18222_));
  INV_X1     g18030(.I(new_n18222_), .ZN(new_n18223_));
  AOI21_X1   g18031(.A1(new_n18215_), .A2(new_n18214_), .B(new_n18223_), .ZN(new_n18224_));
  NAND2_X1   g18032(.A1(new_n18054_), .A2(new_n18224_), .ZN(\asqrt[10] ));
  NOR2_X1    g18033(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n18226_));
  INV_X1     g18034(.I(new_n18226_), .ZN(new_n18227_));
  NOR2_X1    g18035(.A1(new_n18227_), .A2(\a[20] ), .ZN(new_n18228_));
  INV_X1     g18036(.I(new_n18228_), .ZN(new_n18229_));
  AOI21_X1   g18037(.A1(new_n18207_), .A2(new_n18017_), .B(new_n218_), .ZN(new_n18230_));
  OAI21_X1   g18038(.A1(new_n18211_), .A2(new_n18230_), .B(\asqrt[62] ), .ZN(new_n18231_));
  NOR3_X1    g18039(.A1(new_n18211_), .A2(\asqrt[62] ), .A3(new_n18230_), .ZN(new_n18232_));
  OAI21_X1   g18040(.A1(new_n18038_), .A2(new_n18232_), .B(new_n18231_), .ZN(new_n18233_));
  AOI21_X1   g18041(.A1(new_n18233_), .A2(new_n18052_), .B(\asqrt[63] ), .ZN(new_n18234_));
  NAND2_X1   g18042(.A1(new_n18231_), .A2(new_n18049_), .ZN(new_n18235_));
  OAI21_X1   g18043(.A1(new_n18235_), .A2(new_n18041_), .B(new_n18222_), .ZN(new_n18236_));
  OAI21_X1   g18044(.A1(new_n18234_), .A2(new_n18236_), .B(\a[20] ), .ZN(new_n18237_));
  AOI21_X1   g18045(.A1(new_n18237_), .A2(new_n18229_), .B(new_n17623_), .ZN(new_n18238_));
  INV_X1     g18046(.I(\a[20] ), .ZN(new_n18239_));
  AOI21_X1   g18047(.A1(new_n18054_), .A2(new_n18224_), .B(new_n18239_), .ZN(new_n18240_));
  NAND4_X1   g18048(.A1(new_n17598_), .A2(new_n17555_), .A3(new_n17558_), .A4(new_n18229_), .ZN(new_n18241_));
  NOR2_X1    g18049(.A1(new_n18241_), .A2(new_n17570_), .ZN(new_n18242_));
  INV_X1     g18050(.I(new_n18242_), .ZN(new_n18243_));
  NOR2_X1    g18051(.A1(new_n18240_), .A2(new_n18243_), .ZN(new_n18244_));
  AOI21_X1   g18052(.A1(new_n18054_), .A2(new_n18224_), .B(new_n17565_), .ZN(new_n18245_));
  INV_X1     g18053(.I(\a[21] ), .ZN(new_n18246_));
  AOI21_X1   g18054(.A1(\asqrt[10] ), .A2(new_n18239_), .B(new_n18246_), .ZN(new_n18247_));
  NOR3_X1    g18055(.A1(new_n18244_), .A2(new_n18247_), .A3(new_n18245_), .ZN(new_n18248_));
  OAI21_X1   g18056(.A1(new_n18248_), .A2(new_n18238_), .B(\asqrt[12] ), .ZN(new_n18249_));
  OAI21_X1   g18057(.A1(new_n18234_), .A2(new_n18236_), .B(new_n17564_), .ZN(new_n18250_));
  NAND2_X1   g18058(.A1(new_n18215_), .A2(new_n18214_), .ZN(new_n18251_));
  NOR3_X1    g18059(.A1(new_n18218_), .A2(new_n17623_), .A3(new_n18221_), .ZN(new_n18252_));
  NAND3_X1   g18060(.A1(new_n18054_), .A2(new_n18251_), .A3(new_n18252_), .ZN(new_n18253_));
  AOI21_X1   g18061(.A1(new_n18250_), .A2(new_n18253_), .B(new_n17583_), .ZN(new_n18254_));
  AND3_X2    g18062(.A1(new_n18054_), .A2(new_n18251_), .A3(new_n18252_), .Z(new_n18255_));
  NOR3_X1    g18063(.A1(new_n18255_), .A2(\a[22] ), .A3(new_n18245_), .ZN(new_n18256_));
  OAI21_X1   g18064(.A1(new_n18240_), .A2(new_n18228_), .B(\asqrt[11] ), .ZN(new_n18257_));
  NAND2_X1   g18065(.A1(new_n18257_), .A2(new_n16881_), .ZN(new_n18258_));
  OAI22_X1   g18066(.A1(new_n18248_), .A2(new_n18258_), .B1(new_n18254_), .B2(new_n18256_), .ZN(new_n18259_));
  AOI21_X1   g18067(.A1(new_n18259_), .A2(new_n18249_), .B(new_n16389_), .ZN(new_n18260_));
  NOR3_X1    g18068(.A1(new_n18085_), .A2(new_n17582_), .A3(new_n17591_), .ZN(new_n18261_));
  NAND3_X1   g18069(.A1(\asqrt[10] ), .A2(new_n17612_), .A3(new_n18070_), .ZN(new_n18262_));
  AOI22_X1   g18070(.A1(new_n18262_), .A2(new_n18085_), .B1(\asqrt[10] ), .B2(new_n18261_), .ZN(new_n18263_));
  AOI21_X1   g18071(.A1(new_n18054_), .A2(new_n18224_), .B(\a[20] ), .ZN(new_n18264_));
  OAI21_X1   g18072(.A1(new_n18246_), .A2(new_n18264_), .B(new_n18250_), .ZN(new_n18265_));
  OAI21_X1   g18073(.A1(new_n18265_), .A2(new_n18244_), .B(new_n18257_), .ZN(new_n18266_));
  AOI21_X1   g18074(.A1(new_n18266_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n18267_));
  AOI21_X1   g18075(.A1(new_n18267_), .A2(new_n18259_), .B(new_n18263_), .ZN(new_n18268_));
  OAI21_X1   g18076(.A1(new_n18268_), .A2(new_n18260_), .B(\asqrt[14] ), .ZN(new_n18269_));
  INV_X1     g18077(.I(new_n18269_), .ZN(new_n18270_));
  NOR2_X1    g18078(.A1(new_n17604_), .A2(new_n17601_), .ZN(new_n18271_));
  NOR2_X1    g18079(.A1(new_n17595_), .A2(new_n17606_), .ZN(new_n18272_));
  INV_X1     g18080(.I(new_n18272_), .ZN(new_n18273_));
  NAND4_X1   g18081(.A1(\asqrt[10] ), .A2(new_n17596_), .A3(new_n18271_), .A4(new_n18273_), .ZN(new_n18274_));
  INV_X1     g18082(.I(\asqrt[10] ), .ZN(new_n18275_));
  NOR3_X1    g18083(.A1(new_n18275_), .A2(new_n18074_), .A3(new_n18272_), .ZN(new_n18276_));
  OAI21_X1   g18084(.A1(new_n18276_), .A2(new_n18271_), .B(new_n18274_), .ZN(new_n18277_));
  INV_X1     g18085(.I(new_n18277_), .ZN(new_n18278_));
  NOR3_X1    g18086(.A1(new_n18268_), .A2(new_n18260_), .A3(\asqrt[14] ), .ZN(new_n18279_));
  NOR2_X1    g18087(.A1(new_n18279_), .A2(new_n18278_), .ZN(new_n18280_));
  OAI21_X1   g18088(.A1(new_n18280_), .A2(new_n18270_), .B(\asqrt[15] ), .ZN(new_n18281_));
  NOR2_X1    g18089(.A1(new_n18087_), .A2(new_n18079_), .ZN(new_n18282_));
  NOR3_X1    g18090(.A1(new_n18275_), .A2(new_n17608_), .A3(new_n18282_), .ZN(new_n18283_));
  INV_X1     g18091(.I(new_n18283_), .ZN(new_n18284_));
  NOR3_X1    g18092(.A1(new_n18282_), .A2(new_n17608_), .A3(new_n18084_), .ZN(new_n18285_));
  AOI22_X1   g18093(.A1(new_n18284_), .A2(new_n18084_), .B1(\asqrt[10] ), .B2(new_n18285_), .ZN(new_n18286_));
  INV_X1     g18094(.I(new_n18286_), .ZN(new_n18287_));
  NAND2_X1   g18095(.A1(new_n18269_), .A2(new_n15067_), .ZN(new_n18288_));
  OAI21_X1   g18096(.A1(new_n18280_), .A2(new_n18288_), .B(new_n18287_), .ZN(new_n18289_));
  AOI21_X1   g18097(.A1(new_n18289_), .A2(new_n18281_), .B(new_n14601_), .ZN(new_n18290_));
  NOR3_X1    g18098(.A1(new_n17619_), .A2(new_n17627_), .A3(new_n17625_), .ZN(new_n18291_));
  NOR3_X1    g18099(.A1(new_n18275_), .A2(new_n17619_), .A3(new_n17627_), .ZN(new_n18292_));
  INV_X1     g18100(.I(new_n18292_), .ZN(new_n18293_));
  AOI22_X1   g18101(.A1(new_n18293_), .A2(new_n17625_), .B1(\asqrt[10] ), .B2(new_n18291_), .ZN(new_n18294_));
  OAI21_X1   g18102(.A1(new_n18278_), .A2(new_n18279_), .B(new_n18269_), .ZN(new_n18295_));
  AOI21_X1   g18103(.A1(new_n18295_), .A2(\asqrt[15] ), .B(\asqrt[16] ), .ZN(new_n18296_));
  AOI21_X1   g18104(.A1(new_n18296_), .A2(new_n18289_), .B(new_n18294_), .ZN(new_n18297_));
  OAI21_X1   g18105(.A1(new_n18297_), .A2(new_n18290_), .B(\asqrt[17] ), .ZN(new_n18298_));
  NAND2_X1   g18106(.A1(new_n18090_), .A2(new_n18082_), .ZN(new_n18299_));
  NAND3_X1   g18107(.A1(\asqrt[10] ), .A2(new_n17629_), .A3(new_n18299_), .ZN(new_n18300_));
  AND3_X2    g18108(.A1(new_n17629_), .A2(new_n17633_), .A3(new_n18299_), .Z(new_n18301_));
  AOI22_X1   g18109(.A1(new_n18300_), .A2(new_n17634_), .B1(\asqrt[10] ), .B2(new_n18301_), .ZN(new_n18302_));
  INV_X1     g18110(.I(new_n18302_), .ZN(new_n18303_));
  NAND2_X1   g18111(.A1(new_n18237_), .A2(new_n18242_), .ZN(new_n18304_));
  OAI21_X1   g18112(.A1(new_n18234_), .A2(new_n18236_), .B(new_n18239_), .ZN(new_n18305_));
  NAND2_X1   g18113(.A1(new_n18305_), .A2(\a[21] ), .ZN(new_n18306_));
  NAND3_X1   g18114(.A1(new_n18304_), .A2(new_n18306_), .A3(new_n18250_), .ZN(new_n18307_));
  AOI21_X1   g18115(.A1(new_n18307_), .A2(new_n18257_), .B(new_n16881_), .ZN(new_n18308_));
  OAI21_X1   g18116(.A1(new_n18255_), .A2(new_n18245_), .B(\a[22] ), .ZN(new_n18309_));
  NAND3_X1   g18117(.A1(new_n18250_), .A2(new_n18253_), .A3(new_n17583_), .ZN(new_n18310_));
  NAND2_X1   g18118(.A1(new_n18237_), .A2(new_n18229_), .ZN(new_n18311_));
  AOI21_X1   g18119(.A1(new_n18311_), .A2(\asqrt[11] ), .B(\asqrt[12] ), .ZN(new_n18312_));
  AOI22_X1   g18120(.A1(new_n18307_), .A2(new_n18312_), .B1(new_n18309_), .B2(new_n18310_), .ZN(new_n18313_));
  OAI21_X1   g18121(.A1(new_n18313_), .A2(new_n18308_), .B(\asqrt[13] ), .ZN(new_n18314_));
  NAND2_X1   g18122(.A1(new_n18314_), .A2(new_n15770_), .ZN(new_n18315_));
  OAI21_X1   g18123(.A1(new_n18315_), .A2(new_n18268_), .B(new_n18277_), .ZN(new_n18316_));
  AOI21_X1   g18124(.A1(new_n18316_), .A2(new_n18269_), .B(new_n15067_), .ZN(new_n18317_));
  INV_X1     g18125(.I(new_n18263_), .ZN(new_n18318_));
  AOI21_X1   g18126(.A1(\a[21] ), .A2(new_n18305_), .B(new_n18245_), .ZN(new_n18319_));
  AOI21_X1   g18127(.A1(new_n18319_), .A2(new_n18304_), .B(new_n18238_), .ZN(new_n18320_));
  OAI21_X1   g18128(.A1(new_n18320_), .A2(new_n16881_), .B(new_n16389_), .ZN(new_n18321_));
  OAI21_X1   g18129(.A1(new_n18321_), .A2(new_n18313_), .B(new_n18318_), .ZN(new_n18322_));
  NAND2_X1   g18130(.A1(new_n18322_), .A2(new_n18314_), .ZN(new_n18323_));
  AOI21_X1   g18131(.A1(new_n18323_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n18324_));
  AOI21_X1   g18132(.A1(new_n18324_), .A2(new_n18316_), .B(new_n18286_), .ZN(new_n18325_));
  OAI21_X1   g18133(.A1(new_n18325_), .A2(new_n18317_), .B(\asqrt[16] ), .ZN(new_n18326_));
  NAND2_X1   g18134(.A1(new_n18326_), .A2(new_n14017_), .ZN(new_n18327_));
  OAI21_X1   g18135(.A1(new_n18327_), .A2(new_n18297_), .B(new_n18303_), .ZN(new_n18328_));
  AOI21_X1   g18136(.A1(new_n18328_), .A2(new_n18298_), .B(new_n13353_), .ZN(new_n18329_));
  INV_X1     g18137(.I(new_n17641_), .ZN(new_n18330_));
  NOR3_X1    g18138(.A1(new_n17637_), .A2(new_n18101_), .A3(new_n18330_), .ZN(new_n18331_));
  NOR3_X1    g18139(.A1(new_n18275_), .A2(new_n17637_), .A3(new_n18101_), .ZN(new_n18332_));
  INV_X1     g18140(.I(new_n18332_), .ZN(new_n18333_));
  AOI22_X1   g18141(.A1(new_n18333_), .A2(new_n18330_), .B1(\asqrt[10] ), .B2(new_n18331_), .ZN(new_n18334_));
  NOR3_X1    g18142(.A1(new_n18325_), .A2(new_n18317_), .A3(\asqrt[16] ), .ZN(new_n18335_));
  OAI21_X1   g18143(.A1(new_n18294_), .A2(new_n18335_), .B(new_n18326_), .ZN(new_n18336_));
  AOI21_X1   g18144(.A1(new_n18336_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n18337_));
  AOI21_X1   g18145(.A1(new_n18337_), .A2(new_n18328_), .B(new_n18334_), .ZN(new_n18338_));
  OAI21_X1   g18146(.A1(new_n18338_), .A2(new_n18329_), .B(\asqrt[19] ), .ZN(new_n18339_));
  INV_X1     g18147(.I(new_n18339_), .ZN(new_n18340_));
  NOR3_X1    g18148(.A1(new_n18275_), .A2(new_n17646_), .A3(new_n17651_), .ZN(new_n18341_));
  INV_X1     g18149(.I(new_n18341_), .ZN(new_n18342_));
  NOR3_X1    g18150(.A1(new_n17646_), .A2(new_n18069_), .A3(new_n17651_), .ZN(new_n18343_));
  AOI22_X1   g18151(.A1(new_n18342_), .A2(new_n18069_), .B1(\asqrt[10] ), .B2(new_n18343_), .ZN(new_n18344_));
  NOR3_X1    g18152(.A1(new_n18338_), .A2(\asqrt[19] ), .A3(new_n18329_), .ZN(new_n18345_));
  NOR2_X1    g18153(.A1(new_n18345_), .A2(new_n18344_), .ZN(new_n18346_));
  OAI21_X1   g18154(.A1(new_n18346_), .A2(new_n18340_), .B(\asqrt[20] ), .ZN(new_n18347_));
  AND3_X2    g18155(.A1(new_n17653_), .A2(new_n17658_), .A3(new_n18095_), .Z(new_n18348_));
  NAND3_X1   g18156(.A1(\asqrt[10] ), .A2(new_n17653_), .A3(new_n18095_), .ZN(new_n18349_));
  AOI22_X1   g18157(.A1(new_n18349_), .A2(new_n17659_), .B1(\asqrt[10] ), .B2(new_n18348_), .ZN(new_n18350_));
  INV_X1     g18158(.I(new_n18350_), .ZN(new_n18351_));
  NAND2_X1   g18159(.A1(new_n18339_), .A2(new_n12364_), .ZN(new_n18352_));
  OAI21_X1   g18160(.A1(new_n18346_), .A2(new_n18352_), .B(new_n18351_), .ZN(new_n18353_));
  AOI21_X1   g18161(.A1(new_n18353_), .A2(new_n18347_), .B(new_n11736_), .ZN(new_n18354_));
  INV_X1     g18162(.I(new_n17666_), .ZN(new_n18355_));
  NOR3_X1    g18163(.A1(new_n18275_), .A2(new_n17662_), .A3(new_n18105_), .ZN(new_n18356_));
  INV_X1     g18164(.I(new_n18356_), .ZN(new_n18357_));
  NOR3_X1    g18165(.A1(new_n17662_), .A2(new_n18105_), .A3(new_n18355_), .ZN(new_n18358_));
  AOI22_X1   g18166(.A1(new_n18357_), .A2(new_n18355_), .B1(\asqrt[10] ), .B2(new_n18358_), .ZN(new_n18359_));
  NOR3_X1    g18167(.A1(new_n18297_), .A2(new_n18290_), .A3(\asqrt[17] ), .ZN(new_n18360_));
  OAI21_X1   g18168(.A1(new_n18302_), .A2(new_n18360_), .B(new_n18298_), .ZN(new_n18361_));
  INV_X1     g18169(.I(new_n18334_), .ZN(new_n18362_));
  NAND3_X1   g18170(.A1(new_n18328_), .A2(new_n13353_), .A3(new_n18298_), .ZN(new_n18363_));
  AOI22_X1   g18171(.A1(new_n18363_), .A2(new_n18362_), .B1(new_n18361_), .B2(\asqrt[18] ), .ZN(new_n18364_));
  OAI22_X1   g18172(.A1(new_n18345_), .A2(new_n18344_), .B1(new_n18364_), .B2(new_n12913_), .ZN(new_n18365_));
  AOI21_X1   g18173(.A1(new_n18365_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n18366_));
  AOI21_X1   g18174(.A1(new_n18366_), .A2(new_n18353_), .B(new_n18359_), .ZN(new_n18367_));
  OAI21_X1   g18175(.A1(new_n18367_), .A2(new_n18354_), .B(\asqrt[22] ), .ZN(new_n18368_));
  INV_X1     g18176(.I(new_n18368_), .ZN(new_n18369_));
  NOR3_X1    g18177(.A1(new_n17671_), .A2(new_n18068_), .A3(new_n17675_), .ZN(new_n18370_));
  NOR3_X1    g18178(.A1(new_n18275_), .A2(new_n17671_), .A3(new_n17675_), .ZN(new_n18371_));
  INV_X1     g18179(.I(new_n18371_), .ZN(new_n18372_));
  AOI22_X1   g18180(.A1(new_n18372_), .A2(new_n18068_), .B1(\asqrt[10] ), .B2(new_n18370_), .ZN(new_n18373_));
  NOR3_X1    g18181(.A1(new_n18367_), .A2(new_n18354_), .A3(\asqrt[22] ), .ZN(new_n18374_));
  NOR2_X1    g18182(.A1(new_n18374_), .A2(new_n18373_), .ZN(new_n18375_));
  OAI21_X1   g18183(.A1(new_n18375_), .A2(new_n18369_), .B(\asqrt[23] ), .ZN(new_n18376_));
  NOR2_X1    g18184(.A1(new_n17676_), .A2(new_n17684_), .ZN(new_n18377_));
  NOR3_X1    g18185(.A1(new_n18275_), .A2(new_n18099_), .A3(new_n18377_), .ZN(new_n18378_));
  INV_X1     g18186(.I(new_n18378_), .ZN(new_n18379_));
  NOR3_X1    g18187(.A1(new_n18377_), .A2(new_n18099_), .A3(new_n17683_), .ZN(new_n18380_));
  AOI22_X1   g18188(.A1(new_n18379_), .A2(new_n17683_), .B1(\asqrt[10] ), .B2(new_n18380_), .ZN(new_n18381_));
  INV_X1     g18189(.I(new_n18381_), .ZN(new_n18382_));
  NAND2_X1   g18190(.A1(new_n18368_), .A2(new_n10812_), .ZN(new_n18383_));
  OAI21_X1   g18191(.A1(new_n18375_), .A2(new_n18383_), .B(new_n18382_), .ZN(new_n18384_));
  AOI21_X1   g18192(.A1(new_n18384_), .A2(new_n18376_), .B(new_n10221_), .ZN(new_n18385_));
  INV_X1     g18193(.I(new_n17690_), .ZN(new_n18386_));
  NOR3_X1    g18194(.A1(new_n17686_), .A2(new_n18113_), .A3(new_n18386_), .ZN(new_n18387_));
  NOR3_X1    g18195(.A1(new_n18275_), .A2(new_n17686_), .A3(new_n18113_), .ZN(new_n18388_));
  INV_X1     g18196(.I(new_n18388_), .ZN(new_n18389_));
  AOI22_X1   g18197(.A1(new_n18389_), .A2(new_n18386_), .B1(\asqrt[10] ), .B2(new_n18387_), .ZN(new_n18390_));
  OAI21_X1   g18198(.A1(new_n18373_), .A2(new_n18374_), .B(new_n18368_), .ZN(new_n18391_));
  AOI21_X1   g18199(.A1(new_n18391_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n18392_));
  AOI21_X1   g18200(.A1(new_n18392_), .A2(new_n18384_), .B(new_n18390_), .ZN(new_n18393_));
  OAI21_X1   g18201(.A1(new_n18393_), .A2(new_n18385_), .B(\asqrt[25] ), .ZN(new_n18394_));
  INV_X1     g18202(.I(new_n18394_), .ZN(new_n18395_));
  NOR3_X1    g18203(.A1(new_n18275_), .A2(new_n17695_), .A3(new_n17701_), .ZN(new_n18396_));
  INV_X1     g18204(.I(new_n18396_), .ZN(new_n18397_));
  NOR3_X1    g18205(.A1(new_n17695_), .A2(new_n18067_), .A3(new_n17701_), .ZN(new_n18398_));
  AOI22_X1   g18206(.A1(new_n18397_), .A2(new_n18067_), .B1(\asqrt[10] ), .B2(new_n18398_), .ZN(new_n18399_));
  NOR3_X1    g18207(.A1(new_n18393_), .A2(new_n18385_), .A3(\asqrt[25] ), .ZN(new_n18400_));
  NOR2_X1    g18208(.A1(new_n18400_), .A2(new_n18399_), .ZN(new_n18401_));
  OAI21_X1   g18209(.A1(new_n18401_), .A2(new_n18395_), .B(\asqrt[26] ), .ZN(new_n18402_));
  NOR2_X1    g18210(.A1(new_n17702_), .A2(new_n17710_), .ZN(new_n18403_));
  NOR3_X1    g18211(.A1(new_n18403_), .A2(new_n18112_), .A3(new_n17709_), .ZN(new_n18404_));
  NOR3_X1    g18212(.A1(new_n18275_), .A2(new_n18112_), .A3(new_n18403_), .ZN(new_n18405_));
  INV_X1     g18213(.I(new_n18405_), .ZN(new_n18406_));
  AOI22_X1   g18214(.A1(new_n18406_), .A2(new_n17709_), .B1(\asqrt[10] ), .B2(new_n18404_), .ZN(new_n18407_));
  INV_X1     g18215(.I(new_n18407_), .ZN(new_n18408_));
  NAND2_X1   g18216(.A1(new_n18394_), .A2(new_n9317_), .ZN(new_n18409_));
  OAI21_X1   g18217(.A1(new_n18401_), .A2(new_n18409_), .B(new_n18408_), .ZN(new_n18410_));
  AOI21_X1   g18218(.A1(new_n18410_), .A2(new_n18402_), .B(new_n8826_), .ZN(new_n18411_));
  INV_X1     g18219(.I(new_n17716_), .ZN(new_n18412_));
  NOR3_X1    g18220(.A1(new_n18275_), .A2(new_n17712_), .A3(new_n18121_), .ZN(new_n18413_));
  INV_X1     g18221(.I(new_n18413_), .ZN(new_n18414_));
  NOR3_X1    g18222(.A1(new_n17712_), .A2(new_n18121_), .A3(new_n18412_), .ZN(new_n18415_));
  AOI22_X1   g18223(.A1(new_n18414_), .A2(new_n18412_), .B1(\asqrt[10] ), .B2(new_n18415_), .ZN(new_n18416_));
  OAI21_X1   g18224(.A1(new_n18399_), .A2(new_n18400_), .B(new_n18394_), .ZN(new_n18417_));
  AOI21_X1   g18225(.A1(new_n18417_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n18418_));
  AOI21_X1   g18226(.A1(new_n18418_), .A2(new_n18410_), .B(new_n18416_), .ZN(new_n18419_));
  OAI21_X1   g18227(.A1(new_n18419_), .A2(new_n18411_), .B(\asqrt[28] ), .ZN(new_n18420_));
  INV_X1     g18228(.I(new_n18420_), .ZN(new_n18421_));
  INV_X1     g18229(.I(new_n18419_), .ZN(new_n18422_));
  NOR3_X1    g18230(.A1(new_n17721_), .A2(new_n18066_), .A3(new_n17727_), .ZN(new_n18423_));
  NOR3_X1    g18231(.A1(new_n18275_), .A2(new_n17721_), .A3(new_n17727_), .ZN(new_n18424_));
  INV_X1     g18232(.I(new_n18424_), .ZN(new_n18425_));
  AOI22_X1   g18233(.A1(new_n18425_), .A2(new_n18066_), .B1(\asqrt[10] ), .B2(new_n18423_), .ZN(new_n18426_));
  NOR2_X1    g18234(.A1(new_n18411_), .A2(\asqrt[28] ), .ZN(new_n18427_));
  AOI21_X1   g18235(.A1(new_n18422_), .A2(new_n18427_), .B(new_n18426_), .ZN(new_n18428_));
  OAI21_X1   g18236(.A1(new_n18428_), .A2(new_n18421_), .B(\asqrt[29] ), .ZN(new_n18429_));
  NOR2_X1    g18237(.A1(new_n17728_), .A2(new_n17736_), .ZN(new_n18430_));
  NOR3_X1    g18238(.A1(new_n18275_), .A2(new_n18120_), .A3(new_n18430_), .ZN(new_n18431_));
  INV_X1     g18239(.I(new_n18431_), .ZN(new_n18432_));
  NOR3_X1    g18240(.A1(new_n18430_), .A2(new_n18120_), .A3(new_n17735_), .ZN(new_n18433_));
  AOI22_X1   g18241(.A1(new_n18432_), .A2(new_n17735_), .B1(\asqrt[10] ), .B2(new_n18433_), .ZN(new_n18434_));
  INV_X1     g18242(.I(new_n18434_), .ZN(new_n18435_));
  NAND2_X1   g18243(.A1(new_n18420_), .A2(new_n8036_), .ZN(new_n18436_));
  OAI21_X1   g18244(.A1(new_n18436_), .A2(new_n18428_), .B(new_n18435_), .ZN(new_n18437_));
  AOI21_X1   g18245(.A1(new_n18437_), .A2(new_n18429_), .B(new_n7539_), .ZN(new_n18438_));
  INV_X1     g18246(.I(new_n18438_), .ZN(new_n18439_));
  INV_X1     g18247(.I(new_n18437_), .ZN(new_n18440_));
  INV_X1     g18248(.I(new_n17742_), .ZN(new_n18441_));
  NOR3_X1    g18249(.A1(new_n17738_), .A2(new_n18129_), .A3(new_n18441_), .ZN(new_n18442_));
  NOR3_X1    g18250(.A1(new_n18275_), .A2(new_n17738_), .A3(new_n18129_), .ZN(new_n18443_));
  INV_X1     g18251(.I(new_n18443_), .ZN(new_n18444_));
  AOI22_X1   g18252(.A1(new_n18444_), .A2(new_n18441_), .B1(\asqrt[10] ), .B2(new_n18442_), .ZN(new_n18445_));
  INV_X1     g18253(.I(new_n18445_), .ZN(new_n18446_));
  NAND2_X1   g18254(.A1(new_n18429_), .A2(new_n7539_), .ZN(new_n18447_));
  OAI21_X1   g18255(.A1(new_n18447_), .A2(new_n18440_), .B(new_n18446_), .ZN(new_n18448_));
  AOI21_X1   g18256(.A1(new_n18448_), .A2(new_n18439_), .B(new_n7229_), .ZN(new_n18449_));
  NOR3_X1    g18257(.A1(new_n18275_), .A2(new_n17747_), .A3(new_n17753_), .ZN(new_n18450_));
  INV_X1     g18258(.I(new_n18450_), .ZN(new_n18451_));
  NOR3_X1    g18259(.A1(new_n17747_), .A2(new_n18065_), .A3(new_n17753_), .ZN(new_n18452_));
  AOI22_X1   g18260(.A1(new_n18451_), .A2(new_n18065_), .B1(\asqrt[10] ), .B2(new_n18452_), .ZN(new_n18453_));
  NOR2_X1    g18261(.A1(new_n18438_), .A2(\asqrt[31] ), .ZN(new_n18454_));
  AOI21_X1   g18262(.A1(new_n18454_), .A2(new_n18448_), .B(new_n18453_), .ZN(new_n18455_));
  OAI21_X1   g18263(.A1(new_n18455_), .A2(new_n18449_), .B(\asqrt[32] ), .ZN(new_n18456_));
  NOR2_X1    g18264(.A1(new_n17754_), .A2(new_n17762_), .ZN(new_n18457_));
  NOR3_X1    g18265(.A1(new_n18457_), .A2(new_n18128_), .A3(new_n17761_), .ZN(new_n18458_));
  NOR3_X1    g18266(.A1(new_n18275_), .A2(new_n18128_), .A3(new_n18457_), .ZN(new_n18459_));
  INV_X1     g18267(.I(new_n18459_), .ZN(new_n18460_));
  AOI22_X1   g18268(.A1(new_n18460_), .A2(new_n17761_), .B1(\asqrt[10] ), .B2(new_n18458_), .ZN(new_n18461_));
  INV_X1     g18269(.I(new_n18461_), .ZN(new_n18462_));
  NOR3_X1    g18270(.A1(new_n18419_), .A2(new_n18411_), .A3(\asqrt[28] ), .ZN(new_n18463_));
  OAI21_X1   g18271(.A1(new_n18426_), .A2(new_n18463_), .B(new_n18420_), .ZN(new_n18464_));
  AOI21_X1   g18272(.A1(new_n18464_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n18465_));
  AOI21_X1   g18273(.A1(new_n18465_), .A2(new_n18437_), .B(new_n18445_), .ZN(new_n18466_));
  OAI21_X1   g18274(.A1(new_n18466_), .A2(new_n18438_), .B(\asqrt[31] ), .ZN(new_n18467_));
  NAND2_X1   g18275(.A1(new_n18467_), .A2(new_n6824_), .ZN(new_n18468_));
  OAI21_X1   g18276(.A1(new_n18468_), .A2(new_n18455_), .B(new_n18462_), .ZN(new_n18469_));
  AOI21_X1   g18277(.A1(new_n18469_), .A2(new_n18456_), .B(new_n6356_), .ZN(new_n18470_));
  INV_X1     g18278(.I(new_n18470_), .ZN(new_n18471_));
  INV_X1     g18279(.I(new_n18469_), .ZN(new_n18472_));
  INV_X1     g18280(.I(new_n17768_), .ZN(new_n18473_));
  NOR3_X1    g18281(.A1(new_n18275_), .A2(new_n17764_), .A3(new_n18137_), .ZN(new_n18474_));
  INV_X1     g18282(.I(new_n18474_), .ZN(new_n18475_));
  NOR3_X1    g18283(.A1(new_n17764_), .A2(new_n18137_), .A3(new_n18473_), .ZN(new_n18476_));
  AOI22_X1   g18284(.A1(new_n18475_), .A2(new_n18473_), .B1(\asqrt[10] ), .B2(new_n18476_), .ZN(new_n18477_));
  INV_X1     g18285(.I(new_n18477_), .ZN(new_n18478_));
  NAND2_X1   g18286(.A1(new_n18456_), .A2(new_n6356_), .ZN(new_n18479_));
  OAI21_X1   g18287(.A1(new_n18479_), .A2(new_n18472_), .B(new_n18478_), .ZN(new_n18480_));
  AOI21_X1   g18288(.A1(new_n18480_), .A2(new_n18471_), .B(new_n6077_), .ZN(new_n18481_));
  NOR3_X1    g18289(.A1(new_n17773_), .A2(new_n18064_), .A3(new_n17779_), .ZN(new_n18482_));
  NOR3_X1    g18290(.A1(new_n18275_), .A2(new_n17773_), .A3(new_n17779_), .ZN(new_n18483_));
  INV_X1     g18291(.I(new_n18483_), .ZN(new_n18484_));
  AOI22_X1   g18292(.A1(new_n18484_), .A2(new_n18064_), .B1(\asqrt[10] ), .B2(new_n18482_), .ZN(new_n18485_));
  NOR2_X1    g18293(.A1(new_n18470_), .A2(\asqrt[34] ), .ZN(new_n18486_));
  AOI21_X1   g18294(.A1(new_n18486_), .A2(new_n18480_), .B(new_n18485_), .ZN(new_n18487_));
  OAI21_X1   g18295(.A1(new_n18487_), .A2(new_n18481_), .B(\asqrt[35] ), .ZN(new_n18488_));
  NOR2_X1    g18296(.A1(new_n17780_), .A2(new_n17788_), .ZN(new_n18489_));
  NOR3_X1    g18297(.A1(new_n18275_), .A2(new_n18136_), .A3(new_n18489_), .ZN(new_n18490_));
  INV_X1     g18298(.I(new_n18490_), .ZN(new_n18491_));
  NOR3_X1    g18299(.A1(new_n18489_), .A2(new_n18136_), .A3(new_n17787_), .ZN(new_n18492_));
  AOI22_X1   g18300(.A1(new_n18491_), .A2(new_n17787_), .B1(\asqrt[10] ), .B2(new_n18492_), .ZN(new_n18493_));
  INV_X1     g18301(.I(new_n18493_), .ZN(new_n18494_));
  NOR3_X1    g18302(.A1(new_n18466_), .A2(\asqrt[31] ), .A3(new_n18438_), .ZN(new_n18495_));
  OAI21_X1   g18303(.A1(new_n18453_), .A2(new_n18495_), .B(new_n18467_), .ZN(new_n18496_));
  AOI21_X1   g18304(.A1(new_n18496_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n18497_));
  AOI21_X1   g18305(.A1(new_n18497_), .A2(new_n18469_), .B(new_n18477_), .ZN(new_n18498_));
  OAI21_X1   g18306(.A1(new_n18498_), .A2(new_n18470_), .B(\asqrt[34] ), .ZN(new_n18499_));
  NAND2_X1   g18307(.A1(new_n18499_), .A2(new_n5708_), .ZN(new_n18500_));
  OAI21_X1   g18308(.A1(new_n18500_), .A2(new_n18487_), .B(new_n18494_), .ZN(new_n18501_));
  NAND2_X1   g18309(.A1(new_n18501_), .A2(new_n18488_), .ZN(new_n18502_));
  NAND2_X1   g18310(.A1(new_n18502_), .A2(\asqrt[36] ), .ZN(new_n18503_));
  INV_X1     g18311(.I(new_n18501_), .ZN(new_n18504_));
  INV_X1     g18312(.I(new_n17794_), .ZN(new_n18505_));
  NOR3_X1    g18313(.A1(new_n17790_), .A2(new_n18145_), .A3(new_n18505_), .ZN(new_n18506_));
  NOR3_X1    g18314(.A1(new_n18275_), .A2(new_n17790_), .A3(new_n18145_), .ZN(new_n18507_));
  INV_X1     g18315(.I(new_n18507_), .ZN(new_n18508_));
  AOI22_X1   g18316(.A1(new_n18508_), .A2(new_n18505_), .B1(\asqrt[10] ), .B2(new_n18506_), .ZN(new_n18509_));
  INV_X1     g18317(.I(new_n18509_), .ZN(new_n18510_));
  NAND2_X1   g18318(.A1(new_n18488_), .A2(new_n5277_), .ZN(new_n18511_));
  OAI21_X1   g18319(.A1(new_n18504_), .A2(new_n18511_), .B(new_n18510_), .ZN(new_n18512_));
  AOI21_X1   g18320(.A1(new_n18512_), .A2(new_n18503_), .B(new_n5024_), .ZN(new_n18513_));
  NOR3_X1    g18321(.A1(new_n18275_), .A2(new_n17799_), .A3(new_n17805_), .ZN(new_n18514_));
  INV_X1     g18322(.I(new_n18514_), .ZN(new_n18515_));
  NOR3_X1    g18323(.A1(new_n17799_), .A2(new_n18063_), .A3(new_n17805_), .ZN(new_n18516_));
  AOI22_X1   g18324(.A1(new_n18515_), .A2(new_n18063_), .B1(\asqrt[10] ), .B2(new_n18516_), .ZN(new_n18517_));
  AOI21_X1   g18325(.A1(new_n18501_), .A2(new_n18488_), .B(new_n5277_), .ZN(new_n18518_));
  NOR2_X1    g18326(.A1(new_n18518_), .A2(\asqrt[37] ), .ZN(new_n18519_));
  AOI21_X1   g18327(.A1(new_n18519_), .A2(new_n18512_), .B(new_n18517_), .ZN(new_n18520_));
  OAI21_X1   g18328(.A1(new_n18520_), .A2(new_n18513_), .B(\asqrt[38] ), .ZN(new_n18521_));
  INV_X1     g18329(.I(new_n18521_), .ZN(new_n18522_));
  NOR2_X1    g18330(.A1(new_n17806_), .A2(new_n17814_), .ZN(new_n18523_));
  NOR3_X1    g18331(.A1(new_n18523_), .A2(new_n18144_), .A3(new_n17813_), .ZN(new_n18524_));
  NOR3_X1    g18332(.A1(new_n18275_), .A2(new_n18144_), .A3(new_n18523_), .ZN(new_n18525_));
  INV_X1     g18333(.I(new_n18525_), .ZN(new_n18526_));
  AOI22_X1   g18334(.A1(new_n18526_), .A2(new_n17813_), .B1(\asqrt[10] ), .B2(new_n18524_), .ZN(new_n18527_));
  NOR3_X1    g18335(.A1(new_n18520_), .A2(new_n18513_), .A3(\asqrt[38] ), .ZN(new_n18528_));
  NOR2_X1    g18336(.A1(new_n18528_), .A2(new_n18527_), .ZN(new_n18529_));
  OAI21_X1   g18337(.A1(new_n18529_), .A2(new_n18522_), .B(\asqrt[39] ), .ZN(new_n18530_));
  INV_X1     g18338(.I(new_n17820_), .ZN(new_n18531_));
  NOR3_X1    g18339(.A1(new_n18275_), .A2(new_n17816_), .A3(new_n18153_), .ZN(new_n18532_));
  INV_X1     g18340(.I(new_n18532_), .ZN(new_n18533_));
  NOR3_X1    g18341(.A1(new_n17816_), .A2(new_n18153_), .A3(new_n18531_), .ZN(new_n18534_));
  AOI22_X1   g18342(.A1(new_n18533_), .A2(new_n18531_), .B1(\asqrt[10] ), .B2(new_n18534_), .ZN(new_n18535_));
  INV_X1     g18343(.I(new_n18535_), .ZN(new_n18536_));
  NAND2_X1   g18344(.A1(new_n18521_), .A2(new_n4298_), .ZN(new_n18537_));
  OAI21_X1   g18345(.A1(new_n18529_), .A2(new_n18537_), .B(new_n18536_), .ZN(new_n18538_));
  AOI21_X1   g18346(.A1(new_n18538_), .A2(new_n18530_), .B(new_n4071_), .ZN(new_n18539_));
  NOR3_X1    g18347(.A1(new_n17825_), .A2(new_n18062_), .A3(new_n17831_), .ZN(new_n18540_));
  NOR3_X1    g18348(.A1(new_n18275_), .A2(new_n17825_), .A3(new_n17831_), .ZN(new_n18541_));
  INV_X1     g18349(.I(new_n18541_), .ZN(new_n18542_));
  AOI22_X1   g18350(.A1(new_n18542_), .A2(new_n18062_), .B1(\asqrt[10] ), .B2(new_n18540_), .ZN(new_n18543_));
  INV_X1     g18351(.I(new_n18527_), .ZN(new_n18544_));
  NOR3_X1    g18352(.A1(new_n18498_), .A2(\asqrt[34] ), .A3(new_n18470_), .ZN(new_n18545_));
  OAI21_X1   g18353(.A1(new_n18485_), .A2(new_n18545_), .B(new_n18499_), .ZN(new_n18546_));
  AOI21_X1   g18354(.A1(new_n18546_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n18547_));
  AOI21_X1   g18355(.A1(new_n18547_), .A2(new_n18501_), .B(new_n18509_), .ZN(new_n18548_));
  OAI21_X1   g18356(.A1(new_n18548_), .A2(new_n18518_), .B(\asqrt[37] ), .ZN(new_n18549_));
  NAND2_X1   g18357(.A1(new_n18549_), .A2(new_n4696_), .ZN(new_n18550_));
  OAI21_X1   g18358(.A1(new_n18550_), .A2(new_n18520_), .B(new_n18544_), .ZN(new_n18551_));
  AOI21_X1   g18359(.A1(new_n18551_), .A2(new_n18521_), .B(new_n4298_), .ZN(new_n18552_));
  NOR2_X1    g18360(.A1(new_n18552_), .A2(\asqrt[40] ), .ZN(new_n18553_));
  AOI21_X1   g18361(.A1(new_n18553_), .A2(new_n18538_), .B(new_n18543_), .ZN(new_n18554_));
  OAI21_X1   g18362(.A1(new_n18554_), .A2(new_n18539_), .B(\asqrt[41] ), .ZN(new_n18555_));
  NOR2_X1    g18363(.A1(new_n17832_), .A2(new_n17840_), .ZN(new_n18556_));
  NOR3_X1    g18364(.A1(new_n18275_), .A2(new_n18152_), .A3(new_n18556_), .ZN(new_n18557_));
  INV_X1     g18365(.I(new_n18557_), .ZN(new_n18558_));
  NOR3_X1    g18366(.A1(new_n18556_), .A2(new_n18152_), .A3(new_n17839_), .ZN(new_n18559_));
  AOI22_X1   g18367(.A1(new_n18558_), .A2(new_n17839_), .B1(\asqrt[10] ), .B2(new_n18559_), .ZN(new_n18560_));
  INV_X1     g18368(.I(new_n18560_), .ZN(new_n18561_));
  NOR3_X1    g18369(.A1(new_n18548_), .A2(\asqrt[37] ), .A3(new_n18518_), .ZN(new_n18562_));
  OAI21_X1   g18370(.A1(new_n18517_), .A2(new_n18562_), .B(new_n18549_), .ZN(new_n18563_));
  AOI21_X1   g18371(.A1(new_n18563_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n18564_));
  AOI21_X1   g18372(.A1(new_n18564_), .A2(new_n18551_), .B(new_n18535_), .ZN(new_n18565_));
  OAI21_X1   g18373(.A1(new_n18565_), .A2(new_n18552_), .B(\asqrt[40] ), .ZN(new_n18566_));
  NAND2_X1   g18374(.A1(new_n18566_), .A2(new_n3782_), .ZN(new_n18567_));
  OAI21_X1   g18375(.A1(new_n18567_), .A2(new_n18554_), .B(new_n18561_), .ZN(new_n18568_));
  AOI21_X1   g18376(.A1(new_n18568_), .A2(new_n18555_), .B(new_n3419_), .ZN(new_n18569_));
  INV_X1     g18377(.I(new_n17846_), .ZN(new_n18570_));
  NOR3_X1    g18378(.A1(new_n17842_), .A2(new_n18161_), .A3(new_n18570_), .ZN(new_n18571_));
  NOR3_X1    g18379(.A1(new_n18275_), .A2(new_n17842_), .A3(new_n18161_), .ZN(new_n18572_));
  INV_X1     g18380(.I(new_n18572_), .ZN(new_n18573_));
  AOI22_X1   g18381(.A1(new_n18573_), .A2(new_n18570_), .B1(\asqrt[10] ), .B2(new_n18571_), .ZN(new_n18574_));
  NOR3_X1    g18382(.A1(new_n18565_), .A2(\asqrt[40] ), .A3(new_n18552_), .ZN(new_n18575_));
  OAI21_X1   g18383(.A1(new_n18543_), .A2(new_n18575_), .B(new_n18566_), .ZN(new_n18576_));
  AOI21_X1   g18384(.A1(new_n18576_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n18577_));
  AOI21_X1   g18385(.A1(new_n18577_), .A2(new_n18568_), .B(new_n18574_), .ZN(new_n18578_));
  OAI21_X1   g18386(.A1(new_n18578_), .A2(new_n18569_), .B(\asqrt[43] ), .ZN(new_n18579_));
  INV_X1     g18387(.I(new_n18579_), .ZN(new_n18580_));
  NOR3_X1    g18388(.A1(new_n18275_), .A2(new_n17851_), .A3(new_n17857_), .ZN(new_n18581_));
  INV_X1     g18389(.I(new_n18581_), .ZN(new_n18582_));
  NOR3_X1    g18390(.A1(new_n17851_), .A2(new_n18061_), .A3(new_n17857_), .ZN(new_n18583_));
  AOI22_X1   g18391(.A1(new_n18582_), .A2(new_n18061_), .B1(\asqrt[10] ), .B2(new_n18583_), .ZN(new_n18584_));
  NOR3_X1    g18392(.A1(new_n18578_), .A2(\asqrt[43] ), .A3(new_n18569_), .ZN(new_n18585_));
  NOR2_X1    g18393(.A1(new_n18585_), .A2(new_n18584_), .ZN(new_n18586_));
  OAI21_X1   g18394(.A1(new_n18586_), .A2(new_n18580_), .B(\asqrt[44] ), .ZN(new_n18587_));
  NOR2_X1    g18395(.A1(new_n17858_), .A2(new_n17866_), .ZN(new_n18588_));
  NOR3_X1    g18396(.A1(new_n18588_), .A2(new_n18160_), .A3(new_n17865_), .ZN(new_n18589_));
  NOR3_X1    g18397(.A1(new_n18275_), .A2(new_n18160_), .A3(new_n18588_), .ZN(new_n18590_));
  INV_X1     g18398(.I(new_n18590_), .ZN(new_n18591_));
  AOI22_X1   g18399(.A1(new_n18591_), .A2(new_n17865_), .B1(\asqrt[10] ), .B2(new_n18589_), .ZN(new_n18592_));
  INV_X1     g18400(.I(new_n18592_), .ZN(new_n18593_));
  NAND2_X1   g18401(.A1(new_n18579_), .A2(new_n2954_), .ZN(new_n18594_));
  OAI21_X1   g18402(.A1(new_n18586_), .A2(new_n18594_), .B(new_n18593_), .ZN(new_n18595_));
  AOI21_X1   g18403(.A1(new_n18595_), .A2(new_n18587_), .B(new_n2641_), .ZN(new_n18596_));
  INV_X1     g18404(.I(new_n17872_), .ZN(new_n18597_));
  NOR3_X1    g18405(.A1(new_n18275_), .A2(new_n17868_), .A3(new_n18169_), .ZN(new_n18598_));
  INV_X1     g18406(.I(new_n18598_), .ZN(new_n18599_));
  NOR3_X1    g18407(.A1(new_n17868_), .A2(new_n18169_), .A3(new_n18597_), .ZN(new_n18600_));
  AOI22_X1   g18408(.A1(new_n18599_), .A2(new_n18597_), .B1(\asqrt[10] ), .B2(new_n18600_), .ZN(new_n18601_));
  OAI21_X1   g18409(.A1(new_n18584_), .A2(new_n18585_), .B(new_n18579_), .ZN(new_n18602_));
  AOI21_X1   g18410(.A1(new_n18602_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n18603_));
  AOI21_X1   g18411(.A1(new_n18603_), .A2(new_n18595_), .B(new_n18601_), .ZN(new_n18604_));
  OAI21_X1   g18412(.A1(new_n18604_), .A2(new_n18596_), .B(\asqrt[46] ), .ZN(new_n18605_));
  INV_X1     g18413(.I(new_n18605_), .ZN(new_n18606_));
  NOR3_X1    g18414(.A1(new_n17877_), .A2(new_n18060_), .A3(new_n17883_), .ZN(new_n18607_));
  NOR3_X1    g18415(.A1(new_n18275_), .A2(new_n17877_), .A3(new_n17883_), .ZN(new_n18608_));
  INV_X1     g18416(.I(new_n18608_), .ZN(new_n18609_));
  AOI22_X1   g18417(.A1(new_n18609_), .A2(new_n18060_), .B1(\asqrt[10] ), .B2(new_n18607_), .ZN(new_n18610_));
  NOR3_X1    g18418(.A1(new_n18604_), .A2(new_n18596_), .A3(\asqrt[46] ), .ZN(new_n18611_));
  NOR2_X1    g18419(.A1(new_n18611_), .A2(new_n18610_), .ZN(new_n18612_));
  OAI21_X1   g18420(.A1(new_n18612_), .A2(new_n18606_), .B(\asqrt[47] ), .ZN(new_n18613_));
  NOR2_X1    g18421(.A1(new_n17884_), .A2(new_n17892_), .ZN(new_n18614_));
  NOR3_X1    g18422(.A1(new_n18275_), .A2(new_n18168_), .A3(new_n18614_), .ZN(new_n18615_));
  INV_X1     g18423(.I(new_n18615_), .ZN(new_n18616_));
  NOR3_X1    g18424(.A1(new_n18614_), .A2(new_n18168_), .A3(new_n17891_), .ZN(new_n18617_));
  AOI22_X1   g18425(.A1(new_n18616_), .A2(new_n17891_), .B1(\asqrt[10] ), .B2(new_n18617_), .ZN(new_n18618_));
  INV_X1     g18426(.I(new_n18618_), .ZN(new_n18619_));
  NAND2_X1   g18427(.A1(new_n18605_), .A2(new_n2229_), .ZN(new_n18620_));
  OAI21_X1   g18428(.A1(new_n18612_), .A2(new_n18620_), .B(new_n18619_), .ZN(new_n18621_));
  AOI21_X1   g18429(.A1(new_n18621_), .A2(new_n18613_), .B(new_n1956_), .ZN(new_n18622_));
  INV_X1     g18430(.I(new_n17898_), .ZN(new_n18623_));
  NOR3_X1    g18431(.A1(new_n17894_), .A2(new_n18177_), .A3(new_n18623_), .ZN(new_n18624_));
  NOR3_X1    g18432(.A1(new_n18275_), .A2(new_n17894_), .A3(new_n18177_), .ZN(new_n18625_));
  INV_X1     g18433(.I(new_n18625_), .ZN(new_n18626_));
  AOI22_X1   g18434(.A1(new_n18626_), .A2(new_n18623_), .B1(\asqrt[10] ), .B2(new_n18624_), .ZN(new_n18627_));
  OAI21_X1   g18435(.A1(new_n18610_), .A2(new_n18611_), .B(new_n18605_), .ZN(new_n18628_));
  AOI21_X1   g18436(.A1(new_n18628_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n18629_));
  AOI21_X1   g18437(.A1(new_n18629_), .A2(new_n18621_), .B(new_n18627_), .ZN(new_n18630_));
  OAI21_X1   g18438(.A1(new_n18630_), .A2(new_n18622_), .B(\asqrt[49] ), .ZN(new_n18631_));
  INV_X1     g18439(.I(new_n18631_), .ZN(new_n18632_));
  NOR3_X1    g18440(.A1(new_n18275_), .A2(new_n17903_), .A3(new_n17909_), .ZN(new_n18633_));
  INV_X1     g18441(.I(new_n18633_), .ZN(new_n18634_));
  NOR3_X1    g18442(.A1(new_n17903_), .A2(new_n18059_), .A3(new_n17909_), .ZN(new_n18635_));
  AOI22_X1   g18443(.A1(new_n18634_), .A2(new_n18059_), .B1(\asqrt[10] ), .B2(new_n18635_), .ZN(new_n18636_));
  NOR3_X1    g18444(.A1(new_n18630_), .A2(new_n18622_), .A3(\asqrt[49] ), .ZN(new_n18637_));
  NOR2_X1    g18445(.A1(new_n18637_), .A2(new_n18636_), .ZN(new_n18638_));
  OAI21_X1   g18446(.A1(new_n18638_), .A2(new_n18632_), .B(\asqrt[50] ), .ZN(new_n18639_));
  NOR2_X1    g18447(.A1(new_n17910_), .A2(new_n17918_), .ZN(new_n18640_));
  NOR3_X1    g18448(.A1(new_n18640_), .A2(new_n18176_), .A3(new_n17917_), .ZN(new_n18641_));
  NOR3_X1    g18449(.A1(new_n18275_), .A2(new_n18176_), .A3(new_n18640_), .ZN(new_n18642_));
  INV_X1     g18450(.I(new_n18642_), .ZN(new_n18643_));
  AOI22_X1   g18451(.A1(new_n18643_), .A2(new_n17917_), .B1(\asqrt[10] ), .B2(new_n18641_), .ZN(new_n18644_));
  INV_X1     g18452(.I(new_n18644_), .ZN(new_n18645_));
  NAND2_X1   g18453(.A1(new_n18631_), .A2(new_n1612_), .ZN(new_n18646_));
  OAI21_X1   g18454(.A1(new_n18638_), .A2(new_n18646_), .B(new_n18645_), .ZN(new_n18647_));
  AOI21_X1   g18455(.A1(new_n18647_), .A2(new_n18639_), .B(new_n1376_), .ZN(new_n18648_));
  INV_X1     g18456(.I(new_n17924_), .ZN(new_n18649_));
  NOR3_X1    g18457(.A1(new_n18275_), .A2(new_n17920_), .A3(new_n18185_), .ZN(new_n18650_));
  INV_X1     g18458(.I(new_n18650_), .ZN(new_n18651_));
  NOR3_X1    g18459(.A1(new_n17920_), .A2(new_n18185_), .A3(new_n18649_), .ZN(new_n18652_));
  AOI22_X1   g18460(.A1(new_n18651_), .A2(new_n18649_), .B1(\asqrt[10] ), .B2(new_n18652_), .ZN(new_n18653_));
  OAI21_X1   g18461(.A1(new_n18636_), .A2(new_n18637_), .B(new_n18631_), .ZN(new_n18654_));
  AOI21_X1   g18462(.A1(new_n18654_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n18655_));
  AOI21_X1   g18463(.A1(new_n18655_), .A2(new_n18647_), .B(new_n18653_), .ZN(new_n18656_));
  OAI21_X1   g18464(.A1(new_n18656_), .A2(new_n18648_), .B(\asqrt[52] ), .ZN(new_n18657_));
  INV_X1     g18465(.I(new_n18657_), .ZN(new_n18658_));
  INV_X1     g18466(.I(new_n18656_), .ZN(new_n18659_));
  NOR3_X1    g18467(.A1(new_n17929_), .A2(new_n18058_), .A3(new_n17935_), .ZN(new_n18660_));
  NOR3_X1    g18468(.A1(new_n18275_), .A2(new_n17929_), .A3(new_n17935_), .ZN(new_n18661_));
  INV_X1     g18469(.I(new_n18661_), .ZN(new_n18662_));
  AOI22_X1   g18470(.A1(new_n18662_), .A2(new_n18058_), .B1(\asqrt[10] ), .B2(new_n18660_), .ZN(new_n18663_));
  NOR2_X1    g18471(.A1(new_n18648_), .A2(\asqrt[52] ), .ZN(new_n18664_));
  AOI21_X1   g18472(.A1(new_n18659_), .A2(new_n18664_), .B(new_n18663_), .ZN(new_n18665_));
  OAI21_X1   g18473(.A1(new_n18665_), .A2(new_n18658_), .B(\asqrt[53] ), .ZN(new_n18666_));
  NOR2_X1    g18474(.A1(new_n17936_), .A2(new_n17946_), .ZN(new_n18667_));
  NOR3_X1    g18475(.A1(new_n18275_), .A2(new_n18184_), .A3(new_n18667_), .ZN(new_n18668_));
  INV_X1     g18476(.I(new_n18668_), .ZN(new_n18669_));
  NOR3_X1    g18477(.A1(new_n18667_), .A2(new_n18184_), .A3(new_n17945_), .ZN(new_n18670_));
  AOI22_X1   g18478(.A1(new_n18669_), .A2(new_n17945_), .B1(\asqrt[10] ), .B2(new_n18670_), .ZN(new_n18671_));
  INV_X1     g18479(.I(new_n18671_), .ZN(new_n18672_));
  NAND2_X1   g18480(.A1(new_n18657_), .A2(new_n1103_), .ZN(new_n18673_));
  OAI21_X1   g18481(.A1(new_n18673_), .A2(new_n18665_), .B(new_n18672_), .ZN(new_n18674_));
  AOI21_X1   g18482(.A1(new_n18674_), .A2(new_n18666_), .B(new_n904_), .ZN(new_n18675_));
  INV_X1     g18483(.I(new_n18675_), .ZN(new_n18676_));
  INV_X1     g18484(.I(new_n18674_), .ZN(new_n18677_));
  INV_X1     g18485(.I(new_n17952_), .ZN(new_n18678_));
  NOR3_X1    g18486(.A1(new_n17948_), .A2(new_n18193_), .A3(new_n18678_), .ZN(new_n18679_));
  NOR3_X1    g18487(.A1(new_n18275_), .A2(new_n17948_), .A3(new_n18193_), .ZN(new_n18680_));
  INV_X1     g18488(.I(new_n18680_), .ZN(new_n18681_));
  AOI22_X1   g18489(.A1(new_n18681_), .A2(new_n18678_), .B1(\asqrt[10] ), .B2(new_n18679_), .ZN(new_n18682_));
  INV_X1     g18490(.I(new_n18682_), .ZN(new_n18683_));
  NAND2_X1   g18491(.A1(new_n18666_), .A2(new_n904_), .ZN(new_n18684_));
  OAI21_X1   g18492(.A1(new_n18684_), .A2(new_n18677_), .B(new_n18683_), .ZN(new_n18685_));
  AOI21_X1   g18493(.A1(new_n18685_), .A2(new_n18676_), .B(new_n823_), .ZN(new_n18686_));
  NOR3_X1    g18494(.A1(new_n18275_), .A2(new_n17957_), .A3(new_n17964_), .ZN(new_n18687_));
  INV_X1     g18495(.I(new_n18687_), .ZN(new_n18688_));
  NOR3_X1    g18496(.A1(new_n17957_), .A2(new_n18057_), .A3(new_n17964_), .ZN(new_n18689_));
  AOI22_X1   g18497(.A1(new_n18688_), .A2(new_n18057_), .B1(\asqrt[10] ), .B2(new_n18689_), .ZN(new_n18690_));
  NOR2_X1    g18498(.A1(new_n18675_), .A2(\asqrt[55] ), .ZN(new_n18691_));
  AOI21_X1   g18499(.A1(new_n18691_), .A2(new_n18685_), .B(new_n18690_), .ZN(new_n18692_));
  OAI21_X1   g18500(.A1(new_n18692_), .A2(new_n18686_), .B(\asqrt[56] ), .ZN(new_n18693_));
  NOR2_X1    g18501(.A1(new_n17965_), .A2(new_n17977_), .ZN(new_n18694_));
  NOR3_X1    g18502(.A1(new_n18694_), .A2(new_n18192_), .A3(new_n17976_), .ZN(new_n18695_));
  NOR3_X1    g18503(.A1(new_n18275_), .A2(new_n18192_), .A3(new_n18694_), .ZN(new_n18696_));
  INV_X1     g18504(.I(new_n18696_), .ZN(new_n18697_));
  AOI22_X1   g18505(.A1(new_n18697_), .A2(new_n17976_), .B1(\asqrt[10] ), .B2(new_n18695_), .ZN(new_n18698_));
  INV_X1     g18506(.I(new_n18698_), .ZN(new_n18699_));
  NOR3_X1    g18507(.A1(new_n18656_), .A2(new_n18648_), .A3(\asqrt[52] ), .ZN(new_n18700_));
  OAI21_X1   g18508(.A1(new_n18663_), .A2(new_n18700_), .B(new_n18657_), .ZN(new_n18701_));
  AOI21_X1   g18509(.A1(new_n18701_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n18702_));
  AOI21_X1   g18510(.A1(new_n18702_), .A2(new_n18674_), .B(new_n18682_), .ZN(new_n18703_));
  OAI21_X1   g18511(.A1(new_n18703_), .A2(new_n18675_), .B(\asqrt[55] ), .ZN(new_n18704_));
  NAND2_X1   g18512(.A1(new_n18704_), .A2(new_n703_), .ZN(new_n18705_));
  OAI21_X1   g18513(.A1(new_n18705_), .A2(new_n18692_), .B(new_n18699_), .ZN(new_n18706_));
  AOI21_X1   g18514(.A1(new_n18706_), .A2(new_n18693_), .B(new_n531_), .ZN(new_n18707_));
  INV_X1     g18515(.I(new_n18707_), .ZN(new_n18708_));
  INV_X1     g18516(.I(new_n18706_), .ZN(new_n18709_));
  INV_X1     g18517(.I(new_n17983_), .ZN(new_n18710_));
  NOR3_X1    g18518(.A1(new_n18275_), .A2(new_n17979_), .A3(new_n18201_), .ZN(new_n18711_));
  INV_X1     g18519(.I(new_n18711_), .ZN(new_n18712_));
  NOR3_X1    g18520(.A1(new_n17979_), .A2(new_n18201_), .A3(new_n18710_), .ZN(new_n18713_));
  AOI22_X1   g18521(.A1(new_n18712_), .A2(new_n18710_), .B1(\asqrt[10] ), .B2(new_n18713_), .ZN(new_n18714_));
  INV_X1     g18522(.I(new_n18714_), .ZN(new_n18715_));
  NAND2_X1   g18523(.A1(new_n18693_), .A2(new_n531_), .ZN(new_n18716_));
  OAI21_X1   g18524(.A1(new_n18716_), .A2(new_n18709_), .B(new_n18715_), .ZN(new_n18717_));
  AOI21_X1   g18525(.A1(new_n18717_), .A2(new_n18708_), .B(new_n436_), .ZN(new_n18718_));
  NOR3_X1    g18526(.A1(new_n17988_), .A2(new_n18056_), .A3(new_n17995_), .ZN(new_n18719_));
  NOR3_X1    g18527(.A1(new_n18275_), .A2(new_n17988_), .A3(new_n17995_), .ZN(new_n18720_));
  INV_X1     g18528(.I(new_n18720_), .ZN(new_n18721_));
  AOI22_X1   g18529(.A1(new_n18721_), .A2(new_n18056_), .B1(\asqrt[10] ), .B2(new_n18719_), .ZN(new_n18722_));
  NOR2_X1    g18530(.A1(new_n18707_), .A2(\asqrt[58] ), .ZN(new_n18723_));
  AOI21_X1   g18531(.A1(new_n18723_), .A2(new_n18717_), .B(new_n18722_), .ZN(new_n18724_));
  OAI21_X1   g18532(.A1(new_n18724_), .A2(new_n18718_), .B(\asqrt[59] ), .ZN(new_n18725_));
  NOR2_X1    g18533(.A1(new_n17996_), .A2(new_n18007_), .ZN(new_n18726_));
  NOR3_X1    g18534(.A1(new_n18275_), .A2(new_n18200_), .A3(new_n18726_), .ZN(new_n18727_));
  INV_X1     g18535(.I(new_n18727_), .ZN(new_n18728_));
  NOR3_X1    g18536(.A1(new_n18726_), .A2(new_n18200_), .A3(new_n18006_), .ZN(new_n18729_));
  AOI22_X1   g18537(.A1(new_n18728_), .A2(new_n18006_), .B1(\asqrt[10] ), .B2(new_n18729_), .ZN(new_n18730_));
  INV_X1     g18538(.I(new_n18730_), .ZN(new_n18731_));
  NOR3_X1    g18539(.A1(new_n18703_), .A2(\asqrt[55] ), .A3(new_n18675_), .ZN(new_n18732_));
  OAI21_X1   g18540(.A1(new_n18690_), .A2(new_n18732_), .B(new_n18704_), .ZN(new_n18733_));
  AOI21_X1   g18541(.A1(new_n18733_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n18734_));
  AOI21_X1   g18542(.A1(new_n18734_), .A2(new_n18706_), .B(new_n18714_), .ZN(new_n18735_));
  OAI21_X1   g18543(.A1(new_n18735_), .A2(new_n18707_), .B(\asqrt[58] ), .ZN(new_n18736_));
  NAND2_X1   g18544(.A1(new_n18736_), .A2(new_n327_), .ZN(new_n18737_));
  OAI21_X1   g18545(.A1(new_n18737_), .A2(new_n18724_), .B(new_n18731_), .ZN(new_n18738_));
  AOI21_X1   g18546(.A1(new_n18738_), .A2(new_n18725_), .B(new_n306_), .ZN(new_n18739_));
  INV_X1     g18547(.I(new_n18739_), .ZN(new_n18740_));
  INV_X1     g18548(.I(new_n18738_), .ZN(new_n18741_));
  INV_X1     g18549(.I(new_n18013_), .ZN(new_n18742_));
  NOR3_X1    g18550(.A1(new_n18009_), .A2(new_n18208_), .A3(new_n18742_), .ZN(new_n18743_));
  NOR3_X1    g18551(.A1(new_n18275_), .A2(new_n18009_), .A3(new_n18208_), .ZN(new_n18744_));
  INV_X1     g18552(.I(new_n18744_), .ZN(new_n18745_));
  AOI22_X1   g18553(.A1(new_n18745_), .A2(new_n18742_), .B1(\asqrt[10] ), .B2(new_n18743_), .ZN(new_n18746_));
  INV_X1     g18554(.I(new_n18746_), .ZN(new_n18747_));
  NAND2_X1   g18555(.A1(new_n18725_), .A2(new_n306_), .ZN(new_n18748_));
  OAI21_X1   g18556(.A1(new_n18741_), .A2(new_n18748_), .B(new_n18747_), .ZN(new_n18749_));
  AOI21_X1   g18557(.A1(new_n18749_), .A2(new_n18740_), .B(new_n218_), .ZN(new_n18750_));
  NOR3_X1    g18558(.A1(new_n18275_), .A2(new_n18018_), .A3(new_n18024_), .ZN(new_n18751_));
  INV_X1     g18559(.I(new_n18751_), .ZN(new_n18752_));
  NOR3_X1    g18560(.A1(new_n18018_), .A2(new_n18055_), .A3(new_n18024_), .ZN(new_n18753_));
  AOI22_X1   g18561(.A1(new_n18752_), .A2(new_n18055_), .B1(\asqrt[10] ), .B2(new_n18753_), .ZN(new_n18754_));
  NOR2_X1    g18562(.A1(new_n18739_), .A2(\asqrt[61] ), .ZN(new_n18755_));
  AOI21_X1   g18563(.A1(new_n18755_), .A2(new_n18749_), .B(new_n18754_), .ZN(new_n18756_));
  OAI21_X1   g18564(.A1(new_n18756_), .A2(new_n18750_), .B(\asqrt[62] ), .ZN(new_n18757_));
  NOR2_X1    g18565(.A1(new_n18025_), .A2(new_n18032_), .ZN(new_n18758_));
  NOR3_X1    g18566(.A1(new_n18758_), .A2(new_n18230_), .A3(new_n18031_), .ZN(new_n18759_));
  NOR3_X1    g18567(.A1(new_n18275_), .A2(new_n18230_), .A3(new_n18758_), .ZN(new_n18760_));
  INV_X1     g18568(.I(new_n18760_), .ZN(new_n18761_));
  AOI22_X1   g18569(.A1(new_n18761_), .A2(new_n18031_), .B1(\asqrt[10] ), .B2(new_n18759_), .ZN(new_n18762_));
  INV_X1     g18570(.I(new_n18762_), .ZN(new_n18763_));
  NOR3_X1    g18571(.A1(new_n18735_), .A2(\asqrt[58] ), .A3(new_n18707_), .ZN(new_n18764_));
  OAI21_X1   g18572(.A1(new_n18722_), .A2(new_n18764_), .B(new_n18736_), .ZN(new_n18765_));
  AOI21_X1   g18573(.A1(new_n18765_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n18766_));
  AOI21_X1   g18574(.A1(new_n18766_), .A2(new_n18738_), .B(new_n18746_), .ZN(new_n18767_));
  OAI21_X1   g18575(.A1(new_n18767_), .A2(new_n18739_), .B(\asqrt[61] ), .ZN(new_n18768_));
  NAND2_X1   g18576(.A1(new_n18768_), .A2(new_n207_), .ZN(new_n18769_));
  OAI21_X1   g18577(.A1(new_n18769_), .A2(new_n18756_), .B(new_n18763_), .ZN(new_n18770_));
  INV_X1     g18578(.I(new_n18232_), .ZN(new_n18771_));
  NAND4_X1   g18579(.A1(\asqrt[10] ), .A2(new_n18231_), .A3(new_n18038_), .A4(new_n18771_), .ZN(new_n18772_));
  NAND2_X1   g18580(.A1(new_n18771_), .A2(new_n18231_), .ZN(new_n18773_));
  OAI21_X1   g18581(.A1(new_n18275_), .A2(new_n18773_), .B(new_n18212_), .ZN(new_n18774_));
  NAND2_X1   g18582(.A1(new_n18774_), .A2(new_n18772_), .ZN(new_n18775_));
  AOI21_X1   g18583(.A1(new_n18214_), .A2(new_n18231_), .B(new_n18049_), .ZN(new_n18776_));
  NAND2_X1   g18584(.A1(\asqrt[10] ), .A2(new_n18776_), .ZN(new_n18777_));
  NAND3_X1   g18585(.A1(new_n18775_), .A2(new_n18251_), .A3(new_n18777_), .ZN(new_n18778_));
  AOI21_X1   g18586(.A1(new_n18770_), .A2(new_n18757_), .B(new_n18778_), .ZN(new_n18779_));
  NOR2_X1    g18587(.A1(new_n18779_), .A2(\asqrt[63] ), .ZN(new_n18780_));
  INV_X1     g18588(.I(new_n18770_), .ZN(new_n18781_));
  INV_X1     g18589(.I(new_n18775_), .ZN(new_n18782_));
  NAND2_X1   g18590(.A1(new_n18757_), .A2(new_n18782_), .ZN(new_n18783_));
  AOI21_X1   g18591(.A1(\asqrt[10] ), .A2(new_n18050_), .B(new_n18233_), .ZN(new_n18784_));
  OR3_X2     g18592(.A1(new_n18784_), .A2(new_n193_), .A3(new_n18776_), .Z(new_n18785_));
  NOR4_X1    g18593(.A1(new_n18218_), .A2(new_n18046_), .A3(new_n18048_), .A4(new_n18221_), .ZN(new_n18786_));
  AND2_X2    g18594(.A1(new_n18251_), .A2(new_n18786_), .Z(new_n18787_));
  NAND2_X1   g18595(.A1(new_n18787_), .A2(new_n18054_), .ZN(new_n18788_));
  NAND2_X1   g18596(.A1(new_n18785_), .A2(new_n18788_), .ZN(new_n18789_));
  INV_X1     g18597(.I(new_n18789_), .ZN(new_n18790_));
  OAI21_X1   g18598(.A1(new_n18781_), .A2(new_n18783_), .B(new_n18790_), .ZN(new_n18791_));
  NOR2_X1    g18599(.A1(new_n18780_), .A2(new_n18791_), .ZN(new_n18792_));
  INV_X1     g18600(.I(\a[18] ), .ZN(new_n18793_));
  NOR2_X1    g18601(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n18794_));
  INV_X1     g18602(.I(new_n18794_), .ZN(new_n18795_));
  NOR2_X1    g18603(.A1(new_n18795_), .A2(\a[18] ), .ZN(new_n18796_));
  INV_X1     g18604(.I(new_n18796_), .ZN(new_n18797_));
  OAI21_X1   g18605(.A1(new_n18792_), .A2(new_n18793_), .B(new_n18797_), .ZN(new_n18798_));
  NOR3_X1    g18606(.A1(new_n18218_), .A2(new_n18221_), .A3(new_n18796_), .ZN(new_n18799_));
  NAND3_X1   g18607(.A1(new_n18054_), .A2(new_n18251_), .A3(new_n18799_), .ZN(new_n18800_));
  INV_X1     g18608(.I(new_n18800_), .ZN(new_n18801_));
  OAI21_X1   g18609(.A1(new_n18792_), .A2(new_n18793_), .B(new_n18801_), .ZN(new_n18802_));
  NOR3_X1    g18610(.A1(new_n18767_), .A2(\asqrt[61] ), .A3(new_n18739_), .ZN(new_n18803_));
  OAI21_X1   g18611(.A1(new_n18754_), .A2(new_n18803_), .B(new_n18768_), .ZN(new_n18804_));
  INV_X1     g18612(.I(new_n18754_), .ZN(new_n18805_));
  INV_X1     g18613(.I(new_n18722_), .ZN(new_n18806_));
  INV_X1     g18614(.I(new_n18690_), .ZN(new_n18807_));
  INV_X1     g18615(.I(new_n18663_), .ZN(new_n18808_));
  INV_X1     g18616(.I(new_n18636_), .ZN(new_n18809_));
  INV_X1     g18617(.I(new_n18610_), .ZN(new_n18810_));
  INV_X1     g18618(.I(new_n18584_), .ZN(new_n18811_));
  INV_X1     g18619(.I(new_n18555_), .ZN(new_n18812_));
  NOR3_X1    g18620(.A1(new_n18554_), .A2(new_n18539_), .A3(\asqrt[41] ), .ZN(new_n18813_));
  NOR2_X1    g18621(.A1(new_n18813_), .A2(new_n18560_), .ZN(new_n18814_));
  OAI21_X1   g18622(.A1(new_n18814_), .A2(new_n18812_), .B(\asqrt[42] ), .ZN(new_n18815_));
  NAND2_X1   g18623(.A1(new_n18815_), .A2(new_n3218_), .ZN(new_n18816_));
  OAI21_X1   g18624(.A1(new_n18816_), .A2(new_n18578_), .B(new_n18811_), .ZN(new_n18817_));
  NAND3_X1   g18625(.A1(new_n18817_), .A2(new_n2954_), .A3(new_n18579_), .ZN(new_n18818_));
  AOI22_X1   g18626(.A1(new_n18818_), .A2(new_n18593_), .B1(\asqrt[44] ), .B2(new_n18602_), .ZN(new_n18819_));
  OAI21_X1   g18627(.A1(new_n18819_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n18820_));
  OAI21_X1   g18628(.A1(new_n18820_), .A2(new_n18604_), .B(new_n18810_), .ZN(new_n18821_));
  NAND3_X1   g18629(.A1(new_n18821_), .A2(new_n2229_), .A3(new_n18605_), .ZN(new_n18822_));
  AOI22_X1   g18630(.A1(new_n18822_), .A2(new_n18619_), .B1(\asqrt[47] ), .B2(new_n18628_), .ZN(new_n18823_));
  OAI21_X1   g18631(.A1(new_n18823_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n18824_));
  OAI21_X1   g18632(.A1(new_n18824_), .A2(new_n18630_), .B(new_n18809_), .ZN(new_n18825_));
  NAND3_X1   g18633(.A1(new_n18825_), .A2(new_n1612_), .A3(new_n18631_), .ZN(new_n18826_));
  AOI22_X1   g18634(.A1(new_n18826_), .A2(new_n18645_), .B1(\asqrt[50] ), .B2(new_n18654_), .ZN(new_n18827_));
  OAI21_X1   g18635(.A1(new_n18827_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n18828_));
  OAI21_X1   g18636(.A1(new_n18828_), .A2(new_n18656_), .B(new_n18808_), .ZN(new_n18829_));
  NAND3_X1   g18637(.A1(new_n18829_), .A2(new_n1103_), .A3(new_n18657_), .ZN(new_n18830_));
  AOI22_X1   g18638(.A1(new_n18830_), .A2(new_n18672_), .B1(\asqrt[53] ), .B2(new_n18701_), .ZN(new_n18831_));
  OAI21_X1   g18639(.A1(new_n18831_), .A2(new_n904_), .B(new_n823_), .ZN(new_n18832_));
  OAI21_X1   g18640(.A1(new_n18832_), .A2(new_n18703_), .B(new_n18807_), .ZN(new_n18833_));
  NAND3_X1   g18641(.A1(new_n18833_), .A2(new_n703_), .A3(new_n18704_), .ZN(new_n18834_));
  AOI22_X1   g18642(.A1(new_n18834_), .A2(new_n18699_), .B1(\asqrt[56] ), .B2(new_n18733_), .ZN(new_n18835_));
  OAI21_X1   g18643(.A1(new_n18835_), .A2(new_n531_), .B(new_n436_), .ZN(new_n18836_));
  OAI21_X1   g18644(.A1(new_n18836_), .A2(new_n18735_), .B(new_n18806_), .ZN(new_n18837_));
  NAND3_X1   g18645(.A1(new_n18837_), .A2(new_n327_), .A3(new_n18736_), .ZN(new_n18838_));
  AOI22_X1   g18646(.A1(new_n18838_), .A2(new_n18731_), .B1(new_n18765_), .B2(\asqrt[59] ), .ZN(new_n18839_));
  OAI21_X1   g18647(.A1(new_n18839_), .A2(new_n306_), .B(new_n218_), .ZN(new_n18840_));
  OAI21_X1   g18648(.A1(new_n18840_), .A2(new_n18767_), .B(new_n18805_), .ZN(new_n18841_));
  NAND3_X1   g18649(.A1(new_n18841_), .A2(new_n207_), .A3(new_n18768_), .ZN(new_n18842_));
  AOI22_X1   g18650(.A1(new_n18842_), .A2(new_n18763_), .B1(new_n18804_), .B2(\asqrt[62] ), .ZN(new_n18843_));
  OAI21_X1   g18651(.A1(new_n18843_), .A2(new_n18778_), .B(new_n193_), .ZN(new_n18844_));
  AOI21_X1   g18652(.A1(new_n18804_), .A2(\asqrt[62] ), .B(new_n18775_), .ZN(new_n18845_));
  AOI21_X1   g18653(.A1(new_n18845_), .A2(new_n18770_), .B(new_n18789_), .ZN(new_n18846_));
  AOI21_X1   g18654(.A1(new_n18844_), .A2(new_n18846_), .B(new_n18227_), .ZN(new_n18847_));
  OAI21_X1   g18655(.A1(new_n18780_), .A2(new_n18791_), .B(new_n18793_), .ZN(new_n18848_));
  AOI21_X1   g18656(.A1(\a[19] ), .A2(new_n18848_), .B(new_n18847_), .ZN(new_n18849_));
  AOI22_X1   g18657(.A1(new_n18849_), .A2(new_n18802_), .B1(\asqrt[10] ), .B2(new_n18798_), .ZN(new_n18850_));
  NOR2_X1    g18658(.A1(new_n18850_), .A2(new_n17623_), .ZN(new_n18851_));
  NAND2_X1   g18659(.A1(new_n18849_), .A2(new_n18802_), .ZN(new_n18852_));
  OAI21_X1   g18660(.A1(new_n18780_), .A2(new_n18791_), .B(new_n18226_), .ZN(new_n18853_));
  NAND2_X1   g18661(.A1(new_n18845_), .A2(new_n18770_), .ZN(new_n18854_));
  OAI21_X1   g18662(.A1(new_n18787_), .A2(new_n18224_), .B(new_n18054_), .ZN(new_n18855_));
  NAND4_X1   g18663(.A1(new_n18844_), .A2(new_n18854_), .A3(new_n18785_), .A4(new_n18855_), .ZN(new_n18856_));
  AOI21_X1   g18664(.A1(new_n18856_), .A2(new_n18853_), .B(new_n18239_), .ZN(new_n18857_));
  INV_X1     g18665(.I(new_n18854_), .ZN(new_n18858_));
  NAND2_X1   g18666(.A1(new_n18785_), .A2(new_n18855_), .ZN(new_n18859_));
  NOR3_X1    g18667(.A1(new_n18858_), .A2(new_n18780_), .A3(new_n18859_), .ZN(new_n18860_));
  NOR3_X1    g18668(.A1(new_n18860_), .A2(new_n18847_), .A3(\a[20] ), .ZN(new_n18861_));
  NOR2_X1    g18669(.A1(new_n18857_), .A2(new_n18861_), .ZN(new_n18862_));
  AOI21_X1   g18670(.A1(new_n18798_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n18863_));
  AOI21_X1   g18671(.A1(new_n18852_), .A2(new_n18863_), .B(new_n18862_), .ZN(new_n18864_));
  OAI21_X1   g18672(.A1(new_n18864_), .A2(new_n18851_), .B(\asqrt[12] ), .ZN(new_n18865_));
  OAI21_X1   g18673(.A1(\asqrt[63] ), .A2(new_n18779_), .B(new_n18846_), .ZN(\asqrt[9] ));
  NOR3_X1    g18674(.A1(new_n18319_), .A2(new_n18238_), .A3(new_n18244_), .ZN(new_n18867_));
  NAND3_X1   g18675(.A1(\asqrt[9] ), .A2(new_n18257_), .A3(new_n18304_), .ZN(new_n18868_));
  AOI22_X1   g18676(.A1(new_n18868_), .A2(new_n18319_), .B1(\asqrt[9] ), .B2(new_n18867_), .ZN(new_n18869_));
  INV_X1     g18677(.I(new_n18869_), .ZN(new_n18870_));
  OAI21_X1   g18678(.A1(new_n18850_), .A2(new_n17623_), .B(new_n16881_), .ZN(new_n18871_));
  OAI21_X1   g18679(.A1(new_n18871_), .A2(new_n18864_), .B(new_n18870_), .ZN(new_n18872_));
  AOI21_X1   g18680(.A1(new_n18872_), .A2(new_n18865_), .B(new_n16389_), .ZN(new_n18873_));
  NOR2_X1    g18681(.A1(new_n18256_), .A2(new_n18254_), .ZN(new_n18874_));
  NOR2_X1    g18682(.A1(new_n18248_), .A2(new_n18258_), .ZN(new_n18875_));
  INV_X1     g18683(.I(new_n18875_), .ZN(new_n18876_));
  NAND4_X1   g18684(.A1(\asqrt[9] ), .A2(new_n18249_), .A3(new_n18874_), .A4(new_n18876_), .ZN(new_n18877_));
  NOR3_X1    g18685(.A1(new_n18792_), .A2(new_n18308_), .A3(new_n18875_), .ZN(new_n18878_));
  OAI21_X1   g18686(.A1(new_n18878_), .A2(new_n18874_), .B(new_n18877_), .ZN(new_n18879_));
  INV_X1     g18687(.I(new_n18879_), .ZN(new_n18880_));
  AOI21_X1   g18688(.A1(new_n18844_), .A2(new_n18846_), .B(new_n18793_), .ZN(new_n18881_));
  OAI21_X1   g18689(.A1(new_n18881_), .A2(new_n18796_), .B(\asqrt[10] ), .ZN(new_n18882_));
  INV_X1     g18690(.I(new_n18882_), .ZN(new_n18883_));
  NOR2_X1    g18691(.A1(new_n18881_), .A2(new_n18800_), .ZN(new_n18884_));
  INV_X1     g18692(.I(\a[19] ), .ZN(new_n18885_));
  AOI21_X1   g18693(.A1(\asqrt[9] ), .A2(new_n18793_), .B(new_n18885_), .ZN(new_n18886_));
  NOR3_X1    g18694(.A1(new_n18884_), .A2(new_n18886_), .A3(new_n18847_), .ZN(new_n18887_));
  OAI21_X1   g18695(.A1(new_n18887_), .A2(new_n18883_), .B(\asqrt[11] ), .ZN(new_n18888_));
  AOI21_X1   g18696(.A1(\asqrt[9] ), .A2(\a[18] ), .B(new_n18796_), .ZN(new_n18889_));
  OAI21_X1   g18697(.A1(new_n18889_), .A2(new_n18275_), .B(new_n17623_), .ZN(new_n18890_));
  OAI22_X1   g18698(.A1(new_n18887_), .A2(new_n18890_), .B1(new_n18857_), .B2(new_n18861_), .ZN(new_n18891_));
  AOI21_X1   g18699(.A1(new_n18891_), .A2(new_n18888_), .B(new_n16881_), .ZN(new_n18892_));
  AOI21_X1   g18700(.A1(new_n18844_), .A2(new_n18846_), .B(\a[18] ), .ZN(new_n18893_));
  OAI21_X1   g18701(.A1(new_n18885_), .A2(new_n18893_), .B(new_n18853_), .ZN(new_n18894_));
  OAI21_X1   g18702(.A1(new_n18894_), .A2(new_n18884_), .B(new_n18882_), .ZN(new_n18895_));
  AOI21_X1   g18703(.A1(new_n18895_), .A2(\asqrt[11] ), .B(\asqrt[12] ), .ZN(new_n18896_));
  AOI21_X1   g18704(.A1(new_n18896_), .A2(new_n18891_), .B(new_n18869_), .ZN(new_n18897_));
  NOR3_X1    g18705(.A1(new_n18897_), .A2(new_n18892_), .A3(\asqrt[13] ), .ZN(new_n18898_));
  NOR2_X1    g18706(.A1(new_n18898_), .A2(new_n18880_), .ZN(new_n18899_));
  OAI21_X1   g18707(.A1(new_n18899_), .A2(new_n18873_), .B(\asqrt[14] ), .ZN(new_n18900_));
  NOR2_X1    g18708(.A1(new_n18321_), .A2(new_n18313_), .ZN(new_n18901_));
  NOR3_X1    g18709(.A1(new_n18792_), .A2(new_n18260_), .A3(new_n18901_), .ZN(new_n18902_));
  INV_X1     g18710(.I(new_n18902_), .ZN(new_n18903_));
  NOR3_X1    g18711(.A1(new_n18901_), .A2(new_n18260_), .A3(new_n18318_), .ZN(new_n18904_));
  AOI22_X1   g18712(.A1(new_n18903_), .A2(new_n18318_), .B1(\asqrt[9] ), .B2(new_n18904_), .ZN(new_n18905_));
  INV_X1     g18713(.I(new_n18905_), .ZN(new_n18906_));
  OAI21_X1   g18714(.A1(new_n18897_), .A2(new_n18892_), .B(\asqrt[13] ), .ZN(new_n18907_));
  NAND2_X1   g18715(.A1(new_n18907_), .A2(new_n15770_), .ZN(new_n18908_));
  OAI21_X1   g18716(.A1(new_n18899_), .A2(new_n18908_), .B(new_n18906_), .ZN(new_n18909_));
  AOI21_X1   g18717(.A1(new_n18909_), .A2(new_n18900_), .B(new_n15067_), .ZN(new_n18910_));
  NOR3_X1    g18718(.A1(new_n18270_), .A2(new_n18279_), .A3(new_n18277_), .ZN(new_n18911_));
  NOR3_X1    g18719(.A1(new_n18792_), .A2(new_n18270_), .A3(new_n18279_), .ZN(new_n18912_));
  INV_X1     g18720(.I(new_n18912_), .ZN(new_n18913_));
  AOI22_X1   g18721(.A1(new_n18913_), .A2(new_n18277_), .B1(\asqrt[9] ), .B2(new_n18911_), .ZN(new_n18914_));
  OAI21_X1   g18722(.A1(new_n18880_), .A2(new_n18898_), .B(new_n18907_), .ZN(new_n18915_));
  AOI21_X1   g18723(.A1(new_n18915_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n18916_));
  AOI21_X1   g18724(.A1(new_n18916_), .A2(new_n18909_), .B(new_n18914_), .ZN(new_n18917_));
  OAI21_X1   g18725(.A1(new_n18917_), .A2(new_n18910_), .B(\asqrt[16] ), .ZN(new_n18918_));
  INV_X1     g18726(.I(new_n18918_), .ZN(new_n18919_));
  NAND2_X1   g18727(.A1(new_n18324_), .A2(new_n18316_), .ZN(new_n18920_));
  NAND3_X1   g18728(.A1(\asqrt[9] ), .A2(new_n18281_), .A3(new_n18920_), .ZN(new_n18921_));
  AND3_X2    g18729(.A1(new_n18281_), .A2(new_n18286_), .A3(new_n18920_), .Z(new_n18922_));
  AOI22_X1   g18730(.A1(new_n18921_), .A2(new_n18287_), .B1(\asqrt[9] ), .B2(new_n18922_), .ZN(new_n18923_));
  NOR3_X1    g18731(.A1(new_n18917_), .A2(new_n18910_), .A3(\asqrt[16] ), .ZN(new_n18924_));
  NOR2_X1    g18732(.A1(new_n18924_), .A2(new_n18923_), .ZN(new_n18925_));
  OAI21_X1   g18733(.A1(new_n18925_), .A2(new_n18919_), .B(\asqrt[17] ), .ZN(new_n18926_));
  INV_X1     g18734(.I(new_n18294_), .ZN(new_n18927_));
  NOR3_X1    g18735(.A1(new_n18290_), .A2(new_n18335_), .A3(new_n18927_), .ZN(new_n18928_));
  NOR3_X1    g18736(.A1(new_n18792_), .A2(new_n18290_), .A3(new_n18335_), .ZN(new_n18929_));
  INV_X1     g18737(.I(new_n18929_), .ZN(new_n18930_));
  AOI22_X1   g18738(.A1(new_n18930_), .A2(new_n18927_), .B1(\asqrt[9] ), .B2(new_n18928_), .ZN(new_n18931_));
  INV_X1     g18739(.I(new_n18931_), .ZN(new_n18932_));
  NAND2_X1   g18740(.A1(new_n18918_), .A2(new_n14017_), .ZN(new_n18933_));
  OAI21_X1   g18741(.A1(new_n18925_), .A2(new_n18933_), .B(new_n18932_), .ZN(new_n18934_));
  AOI21_X1   g18742(.A1(new_n18934_), .A2(new_n18926_), .B(new_n13353_), .ZN(new_n18935_));
  INV_X1     g18743(.I(new_n18360_), .ZN(new_n18936_));
  NAND3_X1   g18744(.A1(\asqrt[9] ), .A2(new_n18298_), .A3(new_n18936_), .ZN(new_n18937_));
  AND3_X2    g18745(.A1(new_n18936_), .A2(new_n18298_), .A3(new_n18302_), .Z(new_n18938_));
  AOI22_X1   g18746(.A1(new_n18937_), .A2(new_n18303_), .B1(\asqrt[9] ), .B2(new_n18938_), .ZN(new_n18939_));
  OAI21_X1   g18747(.A1(new_n18923_), .A2(new_n18924_), .B(new_n18918_), .ZN(new_n18940_));
  AOI21_X1   g18748(.A1(new_n18940_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n18941_));
  AOI21_X1   g18749(.A1(new_n18941_), .A2(new_n18934_), .B(new_n18939_), .ZN(new_n18942_));
  OAI21_X1   g18750(.A1(new_n18942_), .A2(new_n18935_), .B(\asqrt[19] ), .ZN(new_n18943_));
  INV_X1     g18751(.I(new_n18943_), .ZN(new_n18944_));
  INV_X1     g18752(.I(new_n18363_), .ZN(new_n18945_));
  NOR3_X1    g18753(.A1(new_n18945_), .A2(new_n18329_), .A3(new_n18362_), .ZN(new_n18946_));
  NOR3_X1    g18754(.A1(new_n18792_), .A2(new_n18329_), .A3(new_n18945_), .ZN(new_n18947_));
  INV_X1     g18755(.I(new_n18947_), .ZN(new_n18948_));
  AOI22_X1   g18756(.A1(new_n18948_), .A2(new_n18362_), .B1(\asqrt[9] ), .B2(new_n18946_), .ZN(new_n18949_));
  NOR3_X1    g18757(.A1(new_n18942_), .A2(new_n18935_), .A3(\asqrt[19] ), .ZN(new_n18950_));
  NOR2_X1    g18758(.A1(new_n18950_), .A2(new_n18949_), .ZN(new_n18951_));
  OAI21_X1   g18759(.A1(new_n18951_), .A2(new_n18944_), .B(\asqrt[20] ), .ZN(new_n18952_));
  INV_X1     g18760(.I(new_n18344_), .ZN(new_n18953_));
  NOR3_X1    g18761(.A1(new_n18792_), .A2(new_n18340_), .A3(new_n18345_), .ZN(new_n18954_));
  INV_X1     g18762(.I(new_n18954_), .ZN(new_n18955_));
  NOR3_X1    g18763(.A1(new_n18340_), .A2(new_n18953_), .A3(new_n18345_), .ZN(new_n18956_));
  AOI22_X1   g18764(.A1(new_n18955_), .A2(new_n18953_), .B1(\asqrt[9] ), .B2(new_n18956_), .ZN(new_n18957_));
  INV_X1     g18765(.I(new_n18957_), .ZN(new_n18958_));
  NAND2_X1   g18766(.A1(new_n18943_), .A2(new_n12364_), .ZN(new_n18959_));
  OAI21_X1   g18767(.A1(new_n18951_), .A2(new_n18959_), .B(new_n18958_), .ZN(new_n18960_));
  AOI21_X1   g18768(.A1(new_n18960_), .A2(new_n18952_), .B(new_n11736_), .ZN(new_n18961_));
  OAI21_X1   g18769(.A1(new_n18346_), .A2(new_n18352_), .B(new_n18350_), .ZN(new_n18962_));
  AOI21_X1   g18770(.A1(\asqrt[20] ), .A2(new_n18365_), .B(new_n18962_), .ZN(new_n18963_));
  OAI21_X1   g18771(.A1(new_n18346_), .A2(new_n18352_), .B(new_n18347_), .ZN(new_n18964_));
  NOR2_X1    g18772(.A1(new_n18792_), .A2(new_n18964_), .ZN(new_n18965_));
  INV_X1     g18773(.I(new_n18965_), .ZN(new_n18966_));
  AOI22_X1   g18774(.A1(new_n18966_), .A2(new_n18351_), .B1(\asqrt[9] ), .B2(new_n18963_), .ZN(new_n18967_));
  OAI21_X1   g18775(.A1(new_n18949_), .A2(new_n18950_), .B(new_n18943_), .ZN(new_n18968_));
  AOI21_X1   g18776(.A1(new_n18968_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n18969_));
  AOI21_X1   g18777(.A1(new_n18969_), .A2(new_n18960_), .B(new_n18967_), .ZN(new_n18970_));
  OAI21_X1   g18778(.A1(new_n18970_), .A2(new_n18961_), .B(\asqrt[22] ), .ZN(new_n18971_));
  INV_X1     g18779(.I(new_n18971_), .ZN(new_n18972_));
  INV_X1     g18780(.I(new_n18359_), .ZN(new_n18973_));
  INV_X1     g18781(.I(new_n18353_), .ZN(new_n18974_));
  INV_X1     g18782(.I(new_n18366_), .ZN(new_n18975_));
  NOR2_X1    g18783(.A1(new_n18975_), .A2(new_n18974_), .ZN(new_n18976_));
  NOR3_X1    g18784(.A1(new_n18792_), .A2(new_n18354_), .A3(new_n18976_), .ZN(new_n18977_));
  INV_X1     g18785(.I(new_n18977_), .ZN(new_n18978_));
  NOR3_X1    g18786(.A1(new_n18976_), .A2(new_n18354_), .A3(new_n18973_), .ZN(new_n18979_));
  AOI22_X1   g18787(.A1(new_n18978_), .A2(new_n18973_), .B1(\asqrt[9] ), .B2(new_n18979_), .ZN(new_n18980_));
  NOR3_X1    g18788(.A1(new_n18970_), .A2(new_n18961_), .A3(\asqrt[22] ), .ZN(new_n18981_));
  NOR2_X1    g18789(.A1(new_n18981_), .A2(new_n18980_), .ZN(new_n18982_));
  OAI21_X1   g18790(.A1(new_n18982_), .A2(new_n18972_), .B(\asqrt[23] ), .ZN(new_n18983_));
  INV_X1     g18791(.I(new_n18373_), .ZN(new_n18984_));
  NOR3_X1    g18792(.A1(new_n18369_), .A2(new_n18984_), .A3(new_n18374_), .ZN(new_n18985_));
  NOR3_X1    g18793(.A1(new_n18792_), .A2(new_n18369_), .A3(new_n18374_), .ZN(new_n18986_));
  INV_X1     g18794(.I(new_n18986_), .ZN(new_n18987_));
  AOI22_X1   g18795(.A1(new_n18987_), .A2(new_n18984_), .B1(\asqrt[9] ), .B2(new_n18985_), .ZN(new_n18988_));
  INV_X1     g18796(.I(new_n18988_), .ZN(new_n18989_));
  NAND2_X1   g18797(.A1(new_n18971_), .A2(new_n10812_), .ZN(new_n18990_));
  OAI21_X1   g18798(.A1(new_n18982_), .A2(new_n18990_), .B(new_n18989_), .ZN(new_n18991_));
  AOI21_X1   g18799(.A1(new_n18991_), .A2(new_n18983_), .B(new_n10221_), .ZN(new_n18992_));
  NOR2_X1    g18800(.A1(new_n18375_), .A2(new_n18383_), .ZN(new_n18993_));
  INV_X1     g18801(.I(new_n18993_), .ZN(new_n18994_));
  NAND3_X1   g18802(.A1(\asqrt[9] ), .A2(new_n18376_), .A3(new_n18994_), .ZN(new_n18995_));
  AND3_X2    g18803(.A1(new_n18994_), .A2(new_n18376_), .A3(new_n18381_), .Z(new_n18996_));
  AOI22_X1   g18804(.A1(new_n18995_), .A2(new_n18382_), .B1(\asqrt[9] ), .B2(new_n18996_), .ZN(new_n18997_));
  OAI21_X1   g18805(.A1(new_n18980_), .A2(new_n18981_), .B(new_n18971_), .ZN(new_n18998_));
  AOI21_X1   g18806(.A1(new_n18998_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n18999_));
  AOI21_X1   g18807(.A1(new_n18999_), .A2(new_n18991_), .B(new_n18997_), .ZN(new_n19000_));
  OAI21_X1   g18808(.A1(new_n19000_), .A2(new_n18992_), .B(\asqrt[25] ), .ZN(new_n19001_));
  INV_X1     g18809(.I(new_n19001_), .ZN(new_n19002_));
  INV_X1     g18810(.I(new_n18390_), .ZN(new_n19003_));
  INV_X1     g18811(.I(new_n18384_), .ZN(new_n19004_));
  INV_X1     g18812(.I(new_n18392_), .ZN(new_n19005_));
  NOR2_X1    g18813(.A1(new_n19005_), .A2(new_n19004_), .ZN(new_n19006_));
  NOR3_X1    g18814(.A1(new_n19006_), .A2(new_n18385_), .A3(new_n19003_), .ZN(new_n19007_));
  NOR3_X1    g18815(.A1(new_n18792_), .A2(new_n18385_), .A3(new_n19006_), .ZN(new_n19008_));
  INV_X1     g18816(.I(new_n19008_), .ZN(new_n19009_));
  AOI22_X1   g18817(.A1(new_n19009_), .A2(new_n19003_), .B1(\asqrt[9] ), .B2(new_n19007_), .ZN(new_n19010_));
  NOR3_X1    g18818(.A1(new_n19000_), .A2(new_n18992_), .A3(\asqrt[25] ), .ZN(new_n19011_));
  NOR2_X1    g18819(.A1(new_n19011_), .A2(new_n19010_), .ZN(new_n19012_));
  OAI21_X1   g18820(.A1(new_n19012_), .A2(new_n19002_), .B(\asqrt[26] ), .ZN(new_n19013_));
  INV_X1     g18821(.I(new_n18399_), .ZN(new_n19014_));
  NOR3_X1    g18822(.A1(new_n18792_), .A2(new_n18395_), .A3(new_n18400_), .ZN(new_n19015_));
  INV_X1     g18823(.I(new_n19015_), .ZN(new_n19016_));
  NOR3_X1    g18824(.A1(new_n18395_), .A2(new_n19014_), .A3(new_n18400_), .ZN(new_n19017_));
  AOI22_X1   g18825(.A1(new_n19016_), .A2(new_n19014_), .B1(\asqrt[9] ), .B2(new_n19017_), .ZN(new_n19018_));
  INV_X1     g18826(.I(new_n19018_), .ZN(new_n19019_));
  NAND2_X1   g18827(.A1(new_n19001_), .A2(new_n9317_), .ZN(new_n19020_));
  OAI21_X1   g18828(.A1(new_n19012_), .A2(new_n19020_), .B(new_n19019_), .ZN(new_n19021_));
  AOI21_X1   g18829(.A1(new_n19021_), .A2(new_n19013_), .B(new_n8826_), .ZN(new_n19022_));
  NOR2_X1    g18830(.A1(new_n18401_), .A2(new_n18409_), .ZN(new_n19023_));
  INV_X1     g18831(.I(new_n19023_), .ZN(new_n19024_));
  AND3_X2    g18832(.A1(new_n19024_), .A2(new_n18402_), .A3(new_n18407_), .Z(new_n19025_));
  NAND3_X1   g18833(.A1(\asqrt[9] ), .A2(new_n18402_), .A3(new_n19024_), .ZN(new_n19026_));
  AOI22_X1   g18834(.A1(new_n19026_), .A2(new_n18408_), .B1(\asqrt[9] ), .B2(new_n19025_), .ZN(new_n19027_));
  OAI21_X1   g18835(.A1(new_n19010_), .A2(new_n19011_), .B(new_n19001_), .ZN(new_n19028_));
  AOI21_X1   g18836(.A1(new_n19028_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n19029_));
  AOI21_X1   g18837(.A1(new_n19029_), .A2(new_n19021_), .B(new_n19027_), .ZN(new_n19030_));
  OAI21_X1   g18838(.A1(new_n19030_), .A2(new_n19022_), .B(\asqrt[28] ), .ZN(new_n19031_));
  INV_X1     g18839(.I(new_n19031_), .ZN(new_n19032_));
  INV_X1     g18840(.I(new_n18416_), .ZN(new_n19033_));
  INV_X1     g18841(.I(new_n18410_), .ZN(new_n19034_));
  INV_X1     g18842(.I(new_n18418_), .ZN(new_n19035_));
  NOR2_X1    g18843(.A1(new_n19035_), .A2(new_n19034_), .ZN(new_n19036_));
  NOR3_X1    g18844(.A1(new_n18792_), .A2(new_n18411_), .A3(new_n19036_), .ZN(new_n19037_));
  INV_X1     g18845(.I(new_n19037_), .ZN(new_n19038_));
  NOR3_X1    g18846(.A1(new_n19036_), .A2(new_n18411_), .A3(new_n19033_), .ZN(new_n19039_));
  AOI22_X1   g18847(.A1(new_n19038_), .A2(new_n19033_), .B1(\asqrt[9] ), .B2(new_n19039_), .ZN(new_n19040_));
  NOR3_X1    g18848(.A1(new_n19030_), .A2(new_n19022_), .A3(\asqrt[28] ), .ZN(new_n19041_));
  NOR2_X1    g18849(.A1(new_n19041_), .A2(new_n19040_), .ZN(new_n19042_));
  OAI21_X1   g18850(.A1(new_n19042_), .A2(new_n19032_), .B(\asqrt[29] ), .ZN(new_n19043_));
  INV_X1     g18851(.I(new_n18426_), .ZN(new_n19044_));
  NOR3_X1    g18852(.A1(new_n18421_), .A2(new_n19044_), .A3(new_n18463_), .ZN(new_n19045_));
  NOR3_X1    g18853(.A1(new_n18792_), .A2(new_n18421_), .A3(new_n18463_), .ZN(new_n19046_));
  INV_X1     g18854(.I(new_n19046_), .ZN(new_n19047_));
  AOI22_X1   g18855(.A1(new_n19047_), .A2(new_n19044_), .B1(\asqrt[9] ), .B2(new_n19045_), .ZN(new_n19048_));
  INV_X1     g18856(.I(new_n19048_), .ZN(new_n19049_));
  NAND2_X1   g18857(.A1(new_n19031_), .A2(new_n8036_), .ZN(new_n19050_));
  OAI21_X1   g18858(.A1(new_n19042_), .A2(new_n19050_), .B(new_n19049_), .ZN(new_n19051_));
  AOI21_X1   g18859(.A1(new_n19051_), .A2(new_n19043_), .B(new_n7539_), .ZN(new_n19052_));
  NOR2_X1    g18860(.A1(new_n18436_), .A2(new_n18428_), .ZN(new_n19053_));
  INV_X1     g18861(.I(new_n19053_), .ZN(new_n19054_));
  NAND3_X1   g18862(.A1(\asqrt[9] ), .A2(new_n18429_), .A3(new_n19054_), .ZN(new_n19055_));
  AND3_X2    g18863(.A1(new_n19054_), .A2(new_n18429_), .A3(new_n18434_), .Z(new_n19056_));
  AOI22_X1   g18864(.A1(new_n19055_), .A2(new_n18435_), .B1(\asqrt[9] ), .B2(new_n19056_), .ZN(new_n19057_));
  OAI21_X1   g18865(.A1(new_n19040_), .A2(new_n19041_), .B(new_n19031_), .ZN(new_n19058_));
  AOI21_X1   g18866(.A1(new_n19058_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n19059_));
  AOI21_X1   g18867(.A1(new_n19059_), .A2(new_n19051_), .B(new_n19057_), .ZN(new_n19060_));
  OAI21_X1   g18868(.A1(new_n19060_), .A2(new_n19052_), .B(\asqrt[31] ), .ZN(new_n19061_));
  INV_X1     g18869(.I(new_n19061_), .ZN(new_n19062_));
  NOR2_X1    g18870(.A1(new_n18447_), .A2(new_n18440_), .ZN(new_n19063_));
  NOR3_X1    g18871(.A1(new_n19063_), .A2(new_n18438_), .A3(new_n18446_), .ZN(new_n19064_));
  NOR3_X1    g18872(.A1(new_n18792_), .A2(new_n18438_), .A3(new_n19063_), .ZN(new_n19065_));
  INV_X1     g18873(.I(new_n19065_), .ZN(new_n19066_));
  AOI22_X1   g18874(.A1(new_n19066_), .A2(new_n18446_), .B1(\asqrt[9] ), .B2(new_n19064_), .ZN(new_n19067_));
  NOR3_X1    g18875(.A1(new_n19060_), .A2(new_n19052_), .A3(\asqrt[31] ), .ZN(new_n19068_));
  NOR2_X1    g18876(.A1(new_n19068_), .A2(new_n19067_), .ZN(new_n19069_));
  OAI21_X1   g18877(.A1(new_n19069_), .A2(new_n19062_), .B(\asqrt[32] ), .ZN(new_n19070_));
  INV_X1     g18878(.I(new_n18453_), .ZN(new_n19071_));
  NOR3_X1    g18879(.A1(new_n18792_), .A2(new_n18449_), .A3(new_n18495_), .ZN(new_n19072_));
  INV_X1     g18880(.I(new_n19072_), .ZN(new_n19073_));
  NOR3_X1    g18881(.A1(new_n18449_), .A2(new_n19071_), .A3(new_n18495_), .ZN(new_n19074_));
  AOI22_X1   g18882(.A1(new_n19073_), .A2(new_n19071_), .B1(\asqrt[9] ), .B2(new_n19074_), .ZN(new_n19075_));
  INV_X1     g18883(.I(new_n19075_), .ZN(new_n19076_));
  NAND2_X1   g18884(.A1(new_n19061_), .A2(new_n6824_), .ZN(new_n19077_));
  OAI21_X1   g18885(.A1(new_n19069_), .A2(new_n19077_), .B(new_n19076_), .ZN(new_n19078_));
  AOI21_X1   g18886(.A1(new_n19078_), .A2(new_n19070_), .B(new_n6356_), .ZN(new_n19079_));
  NOR2_X1    g18887(.A1(new_n18468_), .A2(new_n18455_), .ZN(new_n19080_));
  INV_X1     g18888(.I(new_n19080_), .ZN(new_n19081_));
  AND3_X2    g18889(.A1(new_n19081_), .A2(new_n18456_), .A3(new_n18461_), .Z(new_n19082_));
  NAND3_X1   g18890(.A1(\asqrt[9] ), .A2(new_n18456_), .A3(new_n19081_), .ZN(new_n19083_));
  AOI22_X1   g18891(.A1(new_n19083_), .A2(new_n18462_), .B1(\asqrt[9] ), .B2(new_n19082_), .ZN(new_n19084_));
  OAI21_X1   g18892(.A1(new_n19067_), .A2(new_n19068_), .B(new_n19061_), .ZN(new_n19085_));
  AOI21_X1   g18893(.A1(new_n19085_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n19086_));
  AOI21_X1   g18894(.A1(new_n19086_), .A2(new_n19078_), .B(new_n19084_), .ZN(new_n19087_));
  OAI21_X1   g18895(.A1(new_n19087_), .A2(new_n19079_), .B(\asqrt[34] ), .ZN(new_n19088_));
  INV_X1     g18896(.I(new_n19088_), .ZN(new_n19089_));
  NOR2_X1    g18897(.A1(new_n18479_), .A2(new_n18472_), .ZN(new_n19090_));
  NOR3_X1    g18898(.A1(new_n18792_), .A2(new_n18470_), .A3(new_n19090_), .ZN(new_n19091_));
  INV_X1     g18899(.I(new_n19091_), .ZN(new_n19092_));
  NOR3_X1    g18900(.A1(new_n19090_), .A2(new_n18470_), .A3(new_n18478_), .ZN(new_n19093_));
  AOI22_X1   g18901(.A1(new_n19092_), .A2(new_n18478_), .B1(\asqrt[9] ), .B2(new_n19093_), .ZN(new_n19094_));
  NOR3_X1    g18902(.A1(new_n19087_), .A2(new_n19079_), .A3(\asqrt[34] ), .ZN(new_n19095_));
  NOR2_X1    g18903(.A1(new_n19095_), .A2(new_n19094_), .ZN(new_n19096_));
  OAI21_X1   g18904(.A1(new_n19096_), .A2(new_n19089_), .B(\asqrt[35] ), .ZN(new_n19097_));
  INV_X1     g18905(.I(new_n18485_), .ZN(new_n19098_));
  NOR3_X1    g18906(.A1(new_n18481_), .A2(new_n19098_), .A3(new_n18545_), .ZN(new_n19099_));
  NOR3_X1    g18907(.A1(new_n18792_), .A2(new_n18481_), .A3(new_n18545_), .ZN(new_n19100_));
  INV_X1     g18908(.I(new_n19100_), .ZN(new_n19101_));
  AOI22_X1   g18909(.A1(new_n19101_), .A2(new_n19098_), .B1(\asqrt[9] ), .B2(new_n19099_), .ZN(new_n19102_));
  INV_X1     g18910(.I(new_n19102_), .ZN(new_n19103_));
  NAND2_X1   g18911(.A1(new_n19088_), .A2(new_n5708_), .ZN(new_n19104_));
  OAI21_X1   g18912(.A1(new_n19096_), .A2(new_n19104_), .B(new_n19103_), .ZN(new_n19105_));
  AOI21_X1   g18913(.A1(new_n19105_), .A2(new_n19097_), .B(new_n5277_), .ZN(new_n19106_));
  NOR2_X1    g18914(.A1(new_n18500_), .A2(new_n18487_), .ZN(new_n19107_));
  INV_X1     g18915(.I(new_n19107_), .ZN(new_n19108_));
  NAND3_X1   g18916(.A1(\asqrt[9] ), .A2(new_n18488_), .A3(new_n19108_), .ZN(new_n19109_));
  AND3_X2    g18917(.A1(new_n19108_), .A2(new_n18488_), .A3(new_n18493_), .Z(new_n19110_));
  AOI22_X1   g18918(.A1(new_n19109_), .A2(new_n18494_), .B1(\asqrt[9] ), .B2(new_n19110_), .ZN(new_n19111_));
  OAI21_X1   g18919(.A1(new_n19094_), .A2(new_n19095_), .B(new_n19088_), .ZN(new_n19112_));
  AOI21_X1   g18920(.A1(new_n19112_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n19113_));
  AOI21_X1   g18921(.A1(new_n19113_), .A2(new_n19105_), .B(new_n19111_), .ZN(new_n19114_));
  OAI21_X1   g18922(.A1(new_n19114_), .A2(new_n19106_), .B(\asqrt[37] ), .ZN(new_n19115_));
  INV_X1     g18923(.I(new_n19115_), .ZN(new_n19116_));
  NOR2_X1    g18924(.A1(new_n18504_), .A2(new_n18511_), .ZN(new_n19117_));
  NOR3_X1    g18925(.A1(new_n19117_), .A2(new_n18518_), .A3(new_n18510_), .ZN(new_n19118_));
  NOR3_X1    g18926(.A1(new_n18792_), .A2(new_n18518_), .A3(new_n19117_), .ZN(new_n19119_));
  INV_X1     g18927(.I(new_n19119_), .ZN(new_n19120_));
  AOI22_X1   g18928(.A1(new_n19120_), .A2(new_n18510_), .B1(\asqrt[9] ), .B2(new_n19118_), .ZN(new_n19121_));
  NOR3_X1    g18929(.A1(new_n19114_), .A2(new_n19106_), .A3(\asqrt[37] ), .ZN(new_n19122_));
  NOR2_X1    g18930(.A1(new_n19122_), .A2(new_n19121_), .ZN(new_n19123_));
  OAI21_X1   g18931(.A1(new_n19123_), .A2(new_n19116_), .B(\asqrt[38] ), .ZN(new_n19124_));
  INV_X1     g18932(.I(new_n18517_), .ZN(new_n19125_));
  NOR3_X1    g18933(.A1(new_n18792_), .A2(new_n18513_), .A3(new_n18562_), .ZN(new_n19126_));
  INV_X1     g18934(.I(new_n19126_), .ZN(new_n19127_));
  NOR3_X1    g18935(.A1(new_n18513_), .A2(new_n19125_), .A3(new_n18562_), .ZN(new_n19128_));
  AOI22_X1   g18936(.A1(new_n19127_), .A2(new_n19125_), .B1(\asqrt[9] ), .B2(new_n19128_), .ZN(new_n19129_));
  INV_X1     g18937(.I(new_n19129_), .ZN(new_n19130_));
  NAND2_X1   g18938(.A1(new_n19115_), .A2(new_n4696_), .ZN(new_n19131_));
  OAI21_X1   g18939(.A1(new_n19123_), .A2(new_n19131_), .B(new_n19130_), .ZN(new_n19132_));
  AOI21_X1   g18940(.A1(new_n19132_), .A2(new_n19124_), .B(new_n4298_), .ZN(new_n19133_));
  NOR3_X1    g18941(.A1(new_n18522_), .A2(new_n18544_), .A3(new_n18528_), .ZN(new_n19134_));
  NOR3_X1    g18942(.A1(new_n18792_), .A2(new_n18522_), .A3(new_n18528_), .ZN(new_n19135_));
  INV_X1     g18943(.I(new_n19135_), .ZN(new_n19136_));
  AOI22_X1   g18944(.A1(new_n19136_), .A2(new_n18544_), .B1(\asqrt[9] ), .B2(new_n19134_), .ZN(new_n19137_));
  OAI21_X1   g18945(.A1(new_n19121_), .A2(new_n19122_), .B(new_n19115_), .ZN(new_n19138_));
  AOI21_X1   g18946(.A1(new_n19138_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n19139_));
  AOI21_X1   g18947(.A1(new_n19139_), .A2(new_n19132_), .B(new_n19137_), .ZN(new_n19140_));
  OAI21_X1   g18948(.A1(new_n19140_), .A2(new_n19133_), .B(\asqrt[40] ), .ZN(new_n19141_));
  INV_X1     g18949(.I(new_n19141_), .ZN(new_n19142_));
  NOR2_X1    g18950(.A1(new_n18529_), .A2(new_n18537_), .ZN(new_n19143_));
  NOR3_X1    g18951(.A1(new_n18792_), .A2(new_n18552_), .A3(new_n19143_), .ZN(new_n19144_));
  INV_X1     g18952(.I(new_n19144_), .ZN(new_n19145_));
  NOR3_X1    g18953(.A1(new_n19143_), .A2(new_n18552_), .A3(new_n18536_), .ZN(new_n19146_));
  AOI22_X1   g18954(.A1(new_n19145_), .A2(new_n18536_), .B1(\asqrt[9] ), .B2(new_n19146_), .ZN(new_n19147_));
  NOR3_X1    g18955(.A1(new_n19140_), .A2(new_n19133_), .A3(\asqrt[40] ), .ZN(new_n19148_));
  NOR2_X1    g18956(.A1(new_n19148_), .A2(new_n19147_), .ZN(new_n19149_));
  OAI21_X1   g18957(.A1(new_n19149_), .A2(new_n19142_), .B(\asqrt[41] ), .ZN(new_n19150_));
  INV_X1     g18958(.I(new_n18543_), .ZN(new_n19151_));
  NOR3_X1    g18959(.A1(new_n18539_), .A2(new_n19151_), .A3(new_n18575_), .ZN(new_n19152_));
  NOR3_X1    g18960(.A1(new_n18792_), .A2(new_n18539_), .A3(new_n18575_), .ZN(new_n19153_));
  INV_X1     g18961(.I(new_n19153_), .ZN(new_n19154_));
  AOI22_X1   g18962(.A1(new_n19154_), .A2(new_n19151_), .B1(\asqrt[9] ), .B2(new_n19152_), .ZN(new_n19155_));
  INV_X1     g18963(.I(new_n19155_), .ZN(new_n19156_));
  NAND2_X1   g18964(.A1(new_n19141_), .A2(new_n3782_), .ZN(new_n19157_));
  OAI21_X1   g18965(.A1(new_n19149_), .A2(new_n19157_), .B(new_n19156_), .ZN(new_n19158_));
  AOI21_X1   g18966(.A1(new_n19158_), .A2(new_n19150_), .B(new_n3419_), .ZN(new_n19159_));
  NOR3_X1    g18967(.A1(new_n18792_), .A2(new_n18812_), .A3(new_n18813_), .ZN(new_n19160_));
  INV_X1     g18968(.I(new_n19160_), .ZN(new_n19161_));
  NOR3_X1    g18969(.A1(new_n18812_), .A2(new_n18561_), .A3(new_n18813_), .ZN(new_n19162_));
  AOI22_X1   g18970(.A1(new_n19161_), .A2(new_n18561_), .B1(\asqrt[9] ), .B2(new_n19162_), .ZN(new_n19163_));
  OAI21_X1   g18971(.A1(new_n19147_), .A2(new_n19148_), .B(new_n19141_), .ZN(new_n19164_));
  AOI21_X1   g18972(.A1(new_n19164_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n19165_));
  AOI21_X1   g18973(.A1(new_n19165_), .A2(new_n19158_), .B(new_n19163_), .ZN(new_n19166_));
  OAI21_X1   g18974(.A1(new_n19166_), .A2(new_n19159_), .B(\asqrt[43] ), .ZN(new_n19167_));
  INV_X1     g18975(.I(new_n19167_), .ZN(new_n19168_));
  INV_X1     g18976(.I(new_n18574_), .ZN(new_n19169_));
  NAND2_X1   g18977(.A1(new_n18555_), .A2(new_n3419_), .ZN(new_n19170_));
  NOR2_X1    g18978(.A1(new_n18814_), .A2(new_n19170_), .ZN(new_n19171_));
  NOR3_X1    g18979(.A1(new_n19171_), .A2(new_n18569_), .A3(new_n19169_), .ZN(new_n19172_));
  NOR3_X1    g18980(.A1(new_n18792_), .A2(new_n18569_), .A3(new_n19171_), .ZN(new_n19173_));
  INV_X1     g18981(.I(new_n19173_), .ZN(new_n19174_));
  AOI22_X1   g18982(.A1(new_n19174_), .A2(new_n19169_), .B1(\asqrt[9] ), .B2(new_n19172_), .ZN(new_n19175_));
  NOR3_X1    g18983(.A1(new_n19166_), .A2(new_n19159_), .A3(\asqrt[43] ), .ZN(new_n19176_));
  NOR2_X1    g18984(.A1(new_n19176_), .A2(new_n19175_), .ZN(new_n19177_));
  OAI21_X1   g18985(.A1(new_n19177_), .A2(new_n19168_), .B(\asqrt[44] ), .ZN(new_n19178_));
  NOR3_X1    g18986(.A1(new_n18792_), .A2(new_n18580_), .A3(new_n18585_), .ZN(new_n19179_));
  INV_X1     g18987(.I(new_n19179_), .ZN(new_n19180_));
  NOR3_X1    g18988(.A1(new_n18580_), .A2(new_n18585_), .A3(new_n18811_), .ZN(new_n19181_));
  AOI22_X1   g18989(.A1(new_n19180_), .A2(new_n18811_), .B1(\asqrt[9] ), .B2(new_n19181_), .ZN(new_n19182_));
  INV_X1     g18990(.I(new_n19182_), .ZN(new_n19183_));
  NAND2_X1   g18991(.A1(new_n19167_), .A2(new_n2954_), .ZN(new_n19184_));
  OAI21_X1   g18992(.A1(new_n19177_), .A2(new_n19184_), .B(new_n19183_), .ZN(new_n19185_));
  AOI21_X1   g18993(.A1(new_n19185_), .A2(new_n19178_), .B(new_n2641_), .ZN(new_n19186_));
  INV_X1     g18994(.I(new_n18587_), .ZN(new_n19187_));
  NOR2_X1    g18995(.A1(new_n18586_), .A2(new_n18594_), .ZN(new_n19188_));
  NOR3_X1    g18996(.A1(new_n19187_), .A2(new_n19188_), .A3(new_n18593_), .ZN(new_n19189_));
  NOR3_X1    g18997(.A1(new_n18792_), .A2(new_n19187_), .A3(new_n19188_), .ZN(new_n19190_));
  INV_X1     g18998(.I(new_n19190_), .ZN(new_n19191_));
  AOI22_X1   g18999(.A1(new_n19191_), .A2(new_n18593_), .B1(\asqrt[9] ), .B2(new_n19189_), .ZN(new_n19192_));
  OAI21_X1   g19000(.A1(new_n19175_), .A2(new_n19176_), .B(new_n19167_), .ZN(new_n19193_));
  AOI21_X1   g19001(.A1(new_n19193_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n19194_));
  AOI21_X1   g19002(.A1(new_n19194_), .A2(new_n19185_), .B(new_n19192_), .ZN(new_n19195_));
  OAI21_X1   g19003(.A1(new_n19195_), .A2(new_n19186_), .B(\asqrt[46] ), .ZN(new_n19196_));
  INV_X1     g19004(.I(new_n19196_), .ZN(new_n19197_));
  INV_X1     g19005(.I(new_n18601_), .ZN(new_n19198_));
  INV_X1     g19006(.I(new_n18595_), .ZN(new_n19199_));
  INV_X1     g19007(.I(new_n18603_), .ZN(new_n19200_));
  NOR2_X1    g19008(.A1(new_n19200_), .A2(new_n19199_), .ZN(new_n19201_));
  NOR3_X1    g19009(.A1(new_n18792_), .A2(new_n18596_), .A3(new_n19201_), .ZN(new_n19202_));
  INV_X1     g19010(.I(new_n19202_), .ZN(new_n19203_));
  NOR3_X1    g19011(.A1(new_n19201_), .A2(new_n18596_), .A3(new_n19198_), .ZN(new_n19204_));
  AOI22_X1   g19012(.A1(new_n19203_), .A2(new_n19198_), .B1(\asqrt[9] ), .B2(new_n19204_), .ZN(new_n19205_));
  NOR3_X1    g19013(.A1(new_n19195_), .A2(new_n19186_), .A3(\asqrt[46] ), .ZN(new_n19206_));
  NOR2_X1    g19014(.A1(new_n19206_), .A2(new_n19205_), .ZN(new_n19207_));
  OAI21_X1   g19015(.A1(new_n19207_), .A2(new_n19197_), .B(\asqrt[47] ), .ZN(new_n19208_));
  NOR3_X1    g19016(.A1(new_n18606_), .A2(new_n18810_), .A3(new_n18611_), .ZN(new_n19209_));
  NOR3_X1    g19017(.A1(new_n18792_), .A2(new_n18606_), .A3(new_n18611_), .ZN(new_n19210_));
  INV_X1     g19018(.I(new_n19210_), .ZN(new_n19211_));
  AOI22_X1   g19019(.A1(new_n19211_), .A2(new_n18810_), .B1(\asqrt[9] ), .B2(new_n19209_), .ZN(new_n19212_));
  INV_X1     g19020(.I(new_n19212_), .ZN(new_n19213_));
  NAND2_X1   g19021(.A1(new_n19196_), .A2(new_n2229_), .ZN(new_n19214_));
  OAI21_X1   g19022(.A1(new_n19207_), .A2(new_n19214_), .B(new_n19213_), .ZN(new_n19215_));
  AOI21_X1   g19023(.A1(new_n19215_), .A2(new_n19208_), .B(new_n1956_), .ZN(new_n19216_));
  INV_X1     g19024(.I(new_n18613_), .ZN(new_n19217_));
  NOR2_X1    g19025(.A1(new_n18612_), .A2(new_n18620_), .ZN(new_n19218_));
  NOR3_X1    g19026(.A1(new_n18792_), .A2(new_n19217_), .A3(new_n19218_), .ZN(new_n19219_));
  INV_X1     g19027(.I(new_n19219_), .ZN(new_n19220_));
  NOR3_X1    g19028(.A1(new_n19217_), .A2(new_n19218_), .A3(new_n18619_), .ZN(new_n19221_));
  AOI22_X1   g19029(.A1(new_n19220_), .A2(new_n18619_), .B1(\asqrt[9] ), .B2(new_n19221_), .ZN(new_n19222_));
  OAI21_X1   g19030(.A1(new_n19205_), .A2(new_n19206_), .B(new_n19196_), .ZN(new_n19223_));
  AOI21_X1   g19031(.A1(new_n19223_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n19224_));
  AOI21_X1   g19032(.A1(new_n19224_), .A2(new_n19215_), .B(new_n19222_), .ZN(new_n19225_));
  OAI21_X1   g19033(.A1(new_n19225_), .A2(new_n19216_), .B(\asqrt[49] ), .ZN(new_n19226_));
  INV_X1     g19034(.I(new_n19226_), .ZN(new_n19227_));
  INV_X1     g19035(.I(new_n18627_), .ZN(new_n19228_));
  INV_X1     g19036(.I(new_n18621_), .ZN(new_n19229_));
  INV_X1     g19037(.I(new_n18629_), .ZN(new_n19230_));
  NOR2_X1    g19038(.A1(new_n19230_), .A2(new_n19229_), .ZN(new_n19231_));
  NOR3_X1    g19039(.A1(new_n19231_), .A2(new_n18622_), .A3(new_n19228_), .ZN(new_n19232_));
  NOR3_X1    g19040(.A1(new_n18792_), .A2(new_n18622_), .A3(new_n19231_), .ZN(new_n19233_));
  INV_X1     g19041(.I(new_n19233_), .ZN(new_n19234_));
  AOI22_X1   g19042(.A1(new_n19234_), .A2(new_n19228_), .B1(\asqrt[9] ), .B2(new_n19232_), .ZN(new_n19235_));
  NOR3_X1    g19043(.A1(new_n19225_), .A2(new_n19216_), .A3(\asqrt[49] ), .ZN(new_n19236_));
  NOR2_X1    g19044(.A1(new_n19236_), .A2(new_n19235_), .ZN(new_n19237_));
  OAI21_X1   g19045(.A1(new_n19237_), .A2(new_n19227_), .B(\asqrt[50] ), .ZN(new_n19238_));
  NOR3_X1    g19046(.A1(new_n18792_), .A2(new_n18632_), .A3(new_n18637_), .ZN(new_n19239_));
  INV_X1     g19047(.I(new_n19239_), .ZN(new_n19240_));
  NOR3_X1    g19048(.A1(new_n18632_), .A2(new_n18809_), .A3(new_n18637_), .ZN(new_n19241_));
  AOI22_X1   g19049(.A1(new_n19240_), .A2(new_n18809_), .B1(\asqrt[9] ), .B2(new_n19241_), .ZN(new_n19242_));
  INV_X1     g19050(.I(new_n19242_), .ZN(new_n19243_));
  NAND2_X1   g19051(.A1(new_n19226_), .A2(new_n1612_), .ZN(new_n19244_));
  OAI21_X1   g19052(.A1(new_n19237_), .A2(new_n19244_), .B(new_n19243_), .ZN(new_n19245_));
  AOI21_X1   g19053(.A1(new_n19245_), .A2(new_n19238_), .B(new_n1376_), .ZN(new_n19246_));
  INV_X1     g19054(.I(new_n18639_), .ZN(new_n19247_));
  NOR2_X1    g19055(.A1(new_n18638_), .A2(new_n18646_), .ZN(new_n19248_));
  NOR3_X1    g19056(.A1(new_n19247_), .A2(new_n18645_), .A3(new_n19248_), .ZN(new_n19249_));
  NOR3_X1    g19057(.A1(new_n18792_), .A2(new_n19247_), .A3(new_n19248_), .ZN(new_n19250_));
  INV_X1     g19058(.I(new_n19250_), .ZN(new_n19251_));
  AOI22_X1   g19059(.A1(new_n19251_), .A2(new_n18645_), .B1(\asqrt[9] ), .B2(new_n19249_), .ZN(new_n19252_));
  OAI21_X1   g19060(.A1(new_n19235_), .A2(new_n19236_), .B(new_n19226_), .ZN(new_n19253_));
  AOI21_X1   g19061(.A1(new_n19253_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n19254_));
  AOI21_X1   g19062(.A1(new_n19254_), .A2(new_n19245_), .B(new_n19252_), .ZN(new_n19255_));
  OAI21_X1   g19063(.A1(new_n19255_), .A2(new_n19246_), .B(\asqrt[52] ), .ZN(new_n19256_));
  INV_X1     g19064(.I(new_n19256_), .ZN(new_n19257_));
  INV_X1     g19065(.I(new_n18653_), .ZN(new_n19258_));
  INV_X1     g19066(.I(new_n18647_), .ZN(new_n19259_));
  INV_X1     g19067(.I(new_n18655_), .ZN(new_n19260_));
  NOR2_X1    g19068(.A1(new_n19260_), .A2(new_n19259_), .ZN(new_n19261_));
  NOR3_X1    g19069(.A1(new_n18792_), .A2(new_n18648_), .A3(new_n19261_), .ZN(new_n19262_));
  INV_X1     g19070(.I(new_n19262_), .ZN(new_n19263_));
  NOR3_X1    g19071(.A1(new_n19261_), .A2(new_n18648_), .A3(new_n19258_), .ZN(new_n19264_));
  AOI22_X1   g19072(.A1(new_n19263_), .A2(new_n19258_), .B1(\asqrt[9] ), .B2(new_n19264_), .ZN(new_n19265_));
  NOR3_X1    g19073(.A1(new_n19255_), .A2(new_n19246_), .A3(\asqrt[52] ), .ZN(new_n19266_));
  NOR2_X1    g19074(.A1(new_n19266_), .A2(new_n19265_), .ZN(new_n19267_));
  OAI21_X1   g19075(.A1(new_n19267_), .A2(new_n19257_), .B(\asqrt[53] ), .ZN(new_n19268_));
  NOR3_X1    g19076(.A1(new_n18658_), .A2(new_n18808_), .A3(new_n18700_), .ZN(new_n19269_));
  NOR3_X1    g19077(.A1(new_n18792_), .A2(new_n18658_), .A3(new_n18700_), .ZN(new_n19270_));
  INV_X1     g19078(.I(new_n19270_), .ZN(new_n19271_));
  AOI22_X1   g19079(.A1(new_n19271_), .A2(new_n18808_), .B1(\asqrt[9] ), .B2(new_n19269_), .ZN(new_n19272_));
  INV_X1     g19080(.I(new_n19272_), .ZN(new_n19273_));
  NAND2_X1   g19081(.A1(new_n19256_), .A2(new_n1103_), .ZN(new_n19274_));
  OAI21_X1   g19082(.A1(new_n19267_), .A2(new_n19274_), .B(new_n19273_), .ZN(new_n19275_));
  AOI21_X1   g19083(.A1(new_n19275_), .A2(new_n19268_), .B(new_n904_), .ZN(new_n19276_));
  INV_X1     g19084(.I(new_n18666_), .ZN(new_n19277_));
  NOR2_X1    g19085(.A1(new_n18673_), .A2(new_n18665_), .ZN(new_n19278_));
  NOR3_X1    g19086(.A1(new_n18792_), .A2(new_n19277_), .A3(new_n19278_), .ZN(new_n19279_));
  INV_X1     g19087(.I(new_n19279_), .ZN(new_n19280_));
  NOR3_X1    g19088(.A1(new_n19277_), .A2(new_n18672_), .A3(new_n19278_), .ZN(new_n19281_));
  AOI22_X1   g19089(.A1(new_n19280_), .A2(new_n18672_), .B1(\asqrt[9] ), .B2(new_n19281_), .ZN(new_n19282_));
  OAI21_X1   g19090(.A1(new_n19265_), .A2(new_n19266_), .B(new_n19256_), .ZN(new_n19283_));
  AOI21_X1   g19091(.A1(new_n19283_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n19284_));
  AOI21_X1   g19092(.A1(new_n19284_), .A2(new_n19275_), .B(new_n19282_), .ZN(new_n19285_));
  OAI21_X1   g19093(.A1(new_n19285_), .A2(new_n19276_), .B(\asqrt[55] ), .ZN(new_n19286_));
  INV_X1     g19094(.I(new_n19286_), .ZN(new_n19287_));
  NOR2_X1    g19095(.A1(new_n18684_), .A2(new_n18677_), .ZN(new_n19288_));
  NOR3_X1    g19096(.A1(new_n19288_), .A2(new_n18675_), .A3(new_n18683_), .ZN(new_n19289_));
  NOR3_X1    g19097(.A1(new_n18792_), .A2(new_n18675_), .A3(new_n19288_), .ZN(new_n19290_));
  INV_X1     g19098(.I(new_n19290_), .ZN(new_n19291_));
  AOI22_X1   g19099(.A1(new_n19291_), .A2(new_n18683_), .B1(\asqrt[9] ), .B2(new_n19289_), .ZN(new_n19292_));
  NOR3_X1    g19100(.A1(new_n19285_), .A2(new_n19276_), .A3(\asqrt[55] ), .ZN(new_n19293_));
  NOR2_X1    g19101(.A1(new_n19293_), .A2(new_n19292_), .ZN(new_n19294_));
  OAI21_X1   g19102(.A1(new_n19294_), .A2(new_n19287_), .B(\asqrt[56] ), .ZN(new_n19295_));
  NOR3_X1    g19103(.A1(new_n18792_), .A2(new_n18686_), .A3(new_n18732_), .ZN(new_n19296_));
  INV_X1     g19104(.I(new_n19296_), .ZN(new_n19297_));
  NOR3_X1    g19105(.A1(new_n18686_), .A2(new_n18807_), .A3(new_n18732_), .ZN(new_n19298_));
  AOI22_X1   g19106(.A1(new_n19297_), .A2(new_n18807_), .B1(\asqrt[9] ), .B2(new_n19298_), .ZN(new_n19299_));
  INV_X1     g19107(.I(new_n19299_), .ZN(new_n19300_));
  NAND2_X1   g19108(.A1(new_n19286_), .A2(new_n703_), .ZN(new_n19301_));
  OAI21_X1   g19109(.A1(new_n19294_), .A2(new_n19301_), .B(new_n19300_), .ZN(new_n19302_));
  AOI21_X1   g19110(.A1(new_n19302_), .A2(new_n19295_), .B(new_n531_), .ZN(new_n19303_));
  INV_X1     g19111(.I(new_n18693_), .ZN(new_n19304_));
  NOR2_X1    g19112(.A1(new_n18705_), .A2(new_n18692_), .ZN(new_n19305_));
  NOR3_X1    g19113(.A1(new_n19304_), .A2(new_n18699_), .A3(new_n19305_), .ZN(new_n19306_));
  NOR3_X1    g19114(.A1(new_n18792_), .A2(new_n19304_), .A3(new_n19305_), .ZN(new_n19307_));
  INV_X1     g19115(.I(new_n19307_), .ZN(new_n19308_));
  AOI22_X1   g19116(.A1(new_n19308_), .A2(new_n18699_), .B1(\asqrt[9] ), .B2(new_n19306_), .ZN(new_n19309_));
  OAI21_X1   g19117(.A1(new_n19292_), .A2(new_n19293_), .B(new_n19286_), .ZN(new_n19310_));
  AOI21_X1   g19118(.A1(new_n19310_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n19311_));
  AOI21_X1   g19119(.A1(new_n19311_), .A2(new_n19302_), .B(new_n19309_), .ZN(new_n19312_));
  OAI21_X1   g19120(.A1(new_n19312_), .A2(new_n19303_), .B(\asqrt[58] ), .ZN(new_n19313_));
  NOR2_X1    g19121(.A1(new_n18716_), .A2(new_n18709_), .ZN(new_n19314_));
  NOR3_X1    g19122(.A1(new_n18792_), .A2(new_n18707_), .A3(new_n19314_), .ZN(new_n19315_));
  INV_X1     g19123(.I(new_n19315_), .ZN(new_n19316_));
  NOR3_X1    g19124(.A1(new_n19314_), .A2(new_n18707_), .A3(new_n18715_), .ZN(new_n19317_));
  AOI22_X1   g19125(.A1(new_n19316_), .A2(new_n18715_), .B1(\asqrt[9] ), .B2(new_n19317_), .ZN(new_n19318_));
  INV_X1     g19126(.I(new_n19318_), .ZN(new_n19319_));
  INV_X1     g19127(.I(new_n19292_), .ZN(new_n19320_));
  INV_X1     g19128(.I(new_n19265_), .ZN(new_n19321_));
  INV_X1     g19129(.I(new_n19235_), .ZN(new_n19322_));
  INV_X1     g19130(.I(new_n19205_), .ZN(new_n19323_));
  INV_X1     g19131(.I(new_n19175_), .ZN(new_n19324_));
  INV_X1     g19132(.I(new_n19147_), .ZN(new_n19325_));
  INV_X1     g19133(.I(new_n19121_), .ZN(new_n19326_));
  INV_X1     g19134(.I(new_n19094_), .ZN(new_n19327_));
  INV_X1     g19135(.I(new_n19067_), .ZN(new_n19328_));
  INV_X1     g19136(.I(new_n19040_), .ZN(new_n19329_));
  INV_X1     g19137(.I(new_n19010_), .ZN(new_n19330_));
  INV_X1     g19138(.I(new_n18980_), .ZN(new_n19331_));
  INV_X1     g19139(.I(new_n18949_), .ZN(new_n19332_));
  INV_X1     g19140(.I(new_n18923_), .ZN(new_n19333_));
  NAND2_X1   g19141(.A1(new_n18865_), .A2(new_n16389_), .ZN(new_n19334_));
  OAI21_X1   g19142(.A1(new_n19334_), .A2(new_n18897_), .B(new_n18879_), .ZN(new_n19335_));
  AOI21_X1   g19143(.A1(new_n19335_), .A2(new_n18907_), .B(new_n15770_), .ZN(new_n19336_));
  NOR2_X1    g19144(.A1(new_n18873_), .A2(\asqrt[14] ), .ZN(new_n19337_));
  AOI21_X1   g19145(.A1(new_n19337_), .A2(new_n19335_), .B(new_n18905_), .ZN(new_n19338_));
  OAI21_X1   g19146(.A1(new_n19338_), .A2(new_n19336_), .B(\asqrt[15] ), .ZN(new_n19339_));
  NAND2_X1   g19147(.A1(new_n19339_), .A2(new_n14601_), .ZN(new_n19340_));
  OAI21_X1   g19148(.A1(new_n19340_), .A2(new_n18917_), .B(new_n19333_), .ZN(new_n19341_));
  NAND3_X1   g19149(.A1(new_n19341_), .A2(new_n14017_), .A3(new_n18918_), .ZN(new_n19342_));
  AOI22_X1   g19150(.A1(new_n19342_), .A2(new_n18932_), .B1(\asqrt[17] ), .B2(new_n18940_), .ZN(new_n19343_));
  OAI21_X1   g19151(.A1(new_n19343_), .A2(new_n13353_), .B(new_n12913_), .ZN(new_n19344_));
  OAI21_X1   g19152(.A1(new_n19344_), .A2(new_n18942_), .B(new_n19332_), .ZN(new_n19345_));
  AOI21_X1   g19153(.A1(new_n19345_), .A2(new_n18943_), .B(new_n12364_), .ZN(new_n19346_));
  AOI21_X1   g19154(.A1(new_n19341_), .A2(new_n18918_), .B(new_n14017_), .ZN(new_n19347_));
  NOR3_X1    g19155(.A1(new_n19338_), .A2(new_n19336_), .A3(\asqrt[15] ), .ZN(new_n19348_));
  OAI21_X1   g19156(.A1(new_n18914_), .A2(new_n19348_), .B(new_n19339_), .ZN(new_n19349_));
  AOI21_X1   g19157(.A1(new_n19349_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n19350_));
  AOI21_X1   g19158(.A1(new_n19350_), .A2(new_n19341_), .B(new_n18931_), .ZN(new_n19351_));
  NOR3_X1    g19159(.A1(new_n19351_), .A2(\asqrt[18] ), .A3(new_n19347_), .ZN(new_n19352_));
  OAI22_X1   g19160(.A1(new_n19352_), .A2(new_n18939_), .B1(new_n19343_), .B2(new_n13353_), .ZN(new_n19353_));
  AOI21_X1   g19161(.A1(new_n19353_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n19354_));
  AOI21_X1   g19162(.A1(new_n19354_), .A2(new_n19345_), .B(new_n18957_), .ZN(new_n19355_));
  OAI21_X1   g19163(.A1(new_n19355_), .A2(new_n19346_), .B(\asqrt[21] ), .ZN(new_n19356_));
  NAND2_X1   g19164(.A1(new_n19356_), .A2(new_n11326_), .ZN(new_n19357_));
  OAI21_X1   g19165(.A1(new_n19357_), .A2(new_n18970_), .B(new_n19331_), .ZN(new_n19358_));
  AOI21_X1   g19166(.A1(new_n19358_), .A2(new_n18971_), .B(new_n10812_), .ZN(new_n19359_));
  NOR3_X1    g19167(.A1(new_n19355_), .A2(\asqrt[21] ), .A3(new_n19346_), .ZN(new_n19360_));
  OAI21_X1   g19168(.A1(new_n18967_), .A2(new_n19360_), .B(new_n19356_), .ZN(new_n19361_));
  AOI21_X1   g19169(.A1(new_n19361_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n19362_));
  AOI21_X1   g19170(.A1(new_n19362_), .A2(new_n19358_), .B(new_n18988_), .ZN(new_n19363_));
  OAI21_X1   g19171(.A1(new_n19363_), .A2(new_n19359_), .B(\asqrt[24] ), .ZN(new_n19364_));
  NAND2_X1   g19172(.A1(new_n19364_), .A2(new_n9846_), .ZN(new_n19365_));
  OAI21_X1   g19173(.A1(new_n19365_), .A2(new_n19000_), .B(new_n19330_), .ZN(new_n19366_));
  AOI21_X1   g19174(.A1(new_n19366_), .A2(new_n19001_), .B(new_n9317_), .ZN(new_n19367_));
  NOR3_X1    g19175(.A1(new_n19363_), .A2(\asqrt[24] ), .A3(new_n19359_), .ZN(new_n19368_));
  OAI21_X1   g19176(.A1(new_n18997_), .A2(new_n19368_), .B(new_n19364_), .ZN(new_n19369_));
  AOI21_X1   g19177(.A1(new_n19369_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n19370_));
  AOI21_X1   g19178(.A1(new_n19370_), .A2(new_n19366_), .B(new_n19018_), .ZN(new_n19371_));
  OAI21_X1   g19179(.A1(new_n19371_), .A2(new_n19367_), .B(\asqrt[27] ), .ZN(new_n19372_));
  NAND2_X1   g19180(.A1(new_n19372_), .A2(new_n8483_), .ZN(new_n19373_));
  OAI21_X1   g19181(.A1(new_n19373_), .A2(new_n19030_), .B(new_n19329_), .ZN(new_n19374_));
  AOI21_X1   g19182(.A1(new_n19374_), .A2(new_n19031_), .B(new_n8036_), .ZN(new_n19375_));
  NOR3_X1    g19183(.A1(new_n19371_), .A2(\asqrt[27] ), .A3(new_n19367_), .ZN(new_n19376_));
  OAI21_X1   g19184(.A1(new_n19027_), .A2(new_n19376_), .B(new_n19372_), .ZN(new_n19377_));
  AOI21_X1   g19185(.A1(new_n19377_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n19378_));
  AOI21_X1   g19186(.A1(new_n19378_), .A2(new_n19374_), .B(new_n19048_), .ZN(new_n19379_));
  OAI21_X1   g19187(.A1(new_n19379_), .A2(new_n19375_), .B(\asqrt[30] ), .ZN(new_n19380_));
  NAND2_X1   g19188(.A1(new_n19380_), .A2(new_n7229_), .ZN(new_n19381_));
  OAI21_X1   g19189(.A1(new_n19381_), .A2(new_n19060_), .B(new_n19328_), .ZN(new_n19382_));
  AOI21_X1   g19190(.A1(new_n19382_), .A2(new_n19061_), .B(new_n6824_), .ZN(new_n19383_));
  NOR3_X1    g19191(.A1(new_n19379_), .A2(\asqrt[30] ), .A3(new_n19375_), .ZN(new_n19384_));
  OAI21_X1   g19192(.A1(new_n19057_), .A2(new_n19384_), .B(new_n19380_), .ZN(new_n19385_));
  AOI21_X1   g19193(.A1(new_n19385_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n19386_));
  AOI21_X1   g19194(.A1(new_n19386_), .A2(new_n19382_), .B(new_n19075_), .ZN(new_n19387_));
  OAI21_X1   g19195(.A1(new_n19387_), .A2(new_n19383_), .B(\asqrt[33] ), .ZN(new_n19388_));
  NAND2_X1   g19196(.A1(new_n19388_), .A2(new_n6077_), .ZN(new_n19389_));
  OAI21_X1   g19197(.A1(new_n19389_), .A2(new_n19087_), .B(new_n19327_), .ZN(new_n19390_));
  AOI21_X1   g19198(.A1(new_n19390_), .A2(new_n19088_), .B(new_n5708_), .ZN(new_n19391_));
  NOR3_X1    g19199(.A1(new_n19387_), .A2(\asqrt[33] ), .A3(new_n19383_), .ZN(new_n19392_));
  OAI21_X1   g19200(.A1(new_n19084_), .A2(new_n19392_), .B(new_n19388_), .ZN(new_n19393_));
  AOI21_X1   g19201(.A1(new_n19393_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n19394_));
  AOI21_X1   g19202(.A1(new_n19394_), .A2(new_n19390_), .B(new_n19102_), .ZN(new_n19395_));
  OAI21_X1   g19203(.A1(new_n19395_), .A2(new_n19391_), .B(\asqrt[36] ), .ZN(new_n19396_));
  NAND2_X1   g19204(.A1(new_n19396_), .A2(new_n5024_), .ZN(new_n19397_));
  OAI21_X1   g19205(.A1(new_n19397_), .A2(new_n19114_), .B(new_n19326_), .ZN(new_n19398_));
  AOI21_X1   g19206(.A1(new_n19398_), .A2(new_n19115_), .B(new_n4696_), .ZN(new_n19399_));
  NOR3_X1    g19207(.A1(new_n19395_), .A2(\asqrt[36] ), .A3(new_n19391_), .ZN(new_n19400_));
  OAI21_X1   g19208(.A1(new_n19111_), .A2(new_n19400_), .B(new_n19396_), .ZN(new_n19401_));
  AOI21_X1   g19209(.A1(new_n19401_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n19402_));
  AOI21_X1   g19210(.A1(new_n19402_), .A2(new_n19398_), .B(new_n19129_), .ZN(new_n19403_));
  OAI21_X1   g19211(.A1(new_n19403_), .A2(new_n19399_), .B(\asqrt[39] ), .ZN(new_n19404_));
  NAND2_X1   g19212(.A1(new_n19404_), .A2(new_n4071_), .ZN(new_n19405_));
  OAI21_X1   g19213(.A1(new_n19405_), .A2(new_n19140_), .B(new_n19325_), .ZN(new_n19406_));
  AOI21_X1   g19214(.A1(new_n19406_), .A2(new_n19141_), .B(new_n3782_), .ZN(new_n19407_));
  NOR3_X1    g19215(.A1(new_n19403_), .A2(\asqrt[39] ), .A3(new_n19399_), .ZN(new_n19408_));
  OAI21_X1   g19216(.A1(new_n19137_), .A2(new_n19408_), .B(new_n19404_), .ZN(new_n19409_));
  AOI21_X1   g19217(.A1(new_n19409_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n19410_));
  AOI21_X1   g19218(.A1(new_n19410_), .A2(new_n19406_), .B(new_n19155_), .ZN(new_n19411_));
  OAI21_X1   g19219(.A1(new_n19411_), .A2(new_n19407_), .B(\asqrt[42] ), .ZN(new_n19412_));
  NAND2_X1   g19220(.A1(new_n19412_), .A2(new_n3218_), .ZN(new_n19413_));
  OAI21_X1   g19221(.A1(new_n19413_), .A2(new_n19166_), .B(new_n19324_), .ZN(new_n19414_));
  AOI21_X1   g19222(.A1(new_n19414_), .A2(new_n19167_), .B(new_n2954_), .ZN(new_n19415_));
  NOR3_X1    g19223(.A1(new_n19411_), .A2(\asqrt[42] ), .A3(new_n19407_), .ZN(new_n19416_));
  OAI21_X1   g19224(.A1(new_n19163_), .A2(new_n19416_), .B(new_n19412_), .ZN(new_n19417_));
  AOI21_X1   g19225(.A1(new_n19417_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n19418_));
  AOI21_X1   g19226(.A1(new_n19418_), .A2(new_n19414_), .B(new_n19182_), .ZN(new_n19419_));
  OAI21_X1   g19227(.A1(new_n19419_), .A2(new_n19415_), .B(\asqrt[45] ), .ZN(new_n19420_));
  NAND2_X1   g19228(.A1(new_n19420_), .A2(new_n2465_), .ZN(new_n19421_));
  OAI21_X1   g19229(.A1(new_n19421_), .A2(new_n19195_), .B(new_n19323_), .ZN(new_n19422_));
  AOI21_X1   g19230(.A1(new_n19422_), .A2(new_n19196_), .B(new_n2229_), .ZN(new_n19423_));
  NOR3_X1    g19231(.A1(new_n19419_), .A2(\asqrt[45] ), .A3(new_n19415_), .ZN(new_n19424_));
  OAI21_X1   g19232(.A1(new_n19192_), .A2(new_n19424_), .B(new_n19420_), .ZN(new_n19425_));
  AOI21_X1   g19233(.A1(new_n19425_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n19426_));
  AOI21_X1   g19234(.A1(new_n19426_), .A2(new_n19422_), .B(new_n19212_), .ZN(new_n19427_));
  OAI21_X1   g19235(.A1(new_n19427_), .A2(new_n19423_), .B(\asqrt[48] ), .ZN(new_n19428_));
  NAND2_X1   g19236(.A1(new_n19428_), .A2(new_n1806_), .ZN(new_n19429_));
  OAI21_X1   g19237(.A1(new_n19429_), .A2(new_n19225_), .B(new_n19322_), .ZN(new_n19430_));
  AOI21_X1   g19238(.A1(new_n19430_), .A2(new_n19226_), .B(new_n1612_), .ZN(new_n19431_));
  NOR3_X1    g19239(.A1(new_n19427_), .A2(\asqrt[48] ), .A3(new_n19423_), .ZN(new_n19432_));
  OAI21_X1   g19240(.A1(new_n19222_), .A2(new_n19432_), .B(new_n19428_), .ZN(new_n19433_));
  AOI21_X1   g19241(.A1(new_n19433_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n19434_));
  AOI21_X1   g19242(.A1(new_n19434_), .A2(new_n19430_), .B(new_n19242_), .ZN(new_n19435_));
  OAI21_X1   g19243(.A1(new_n19435_), .A2(new_n19431_), .B(\asqrt[51] ), .ZN(new_n19436_));
  NAND2_X1   g19244(.A1(new_n19436_), .A2(new_n1256_), .ZN(new_n19437_));
  OAI21_X1   g19245(.A1(new_n19437_), .A2(new_n19255_), .B(new_n19321_), .ZN(new_n19438_));
  NAND3_X1   g19246(.A1(new_n19438_), .A2(new_n1103_), .A3(new_n19256_), .ZN(new_n19439_));
  AOI22_X1   g19247(.A1(new_n19439_), .A2(new_n19273_), .B1(\asqrt[53] ), .B2(new_n19283_), .ZN(new_n19440_));
  OAI21_X1   g19248(.A1(new_n19440_), .A2(new_n904_), .B(new_n823_), .ZN(new_n19441_));
  OAI21_X1   g19249(.A1(new_n19441_), .A2(new_n19285_), .B(new_n19320_), .ZN(new_n19442_));
  NAND3_X1   g19250(.A1(new_n19442_), .A2(new_n703_), .A3(new_n19286_), .ZN(new_n19443_));
  AOI22_X1   g19251(.A1(new_n19443_), .A2(new_n19300_), .B1(\asqrt[56] ), .B2(new_n19310_), .ZN(new_n19444_));
  OAI21_X1   g19252(.A1(new_n19444_), .A2(new_n531_), .B(new_n436_), .ZN(new_n19445_));
  OAI21_X1   g19253(.A1(new_n19445_), .A2(new_n19312_), .B(new_n19319_), .ZN(new_n19446_));
  AOI21_X1   g19254(.A1(new_n19446_), .A2(new_n19313_), .B(new_n327_), .ZN(new_n19447_));
  NOR3_X1    g19255(.A1(new_n18718_), .A2(new_n18806_), .A3(new_n18764_), .ZN(new_n19448_));
  NOR3_X1    g19256(.A1(new_n18792_), .A2(new_n18718_), .A3(new_n18764_), .ZN(new_n19449_));
  INV_X1     g19257(.I(new_n19449_), .ZN(new_n19450_));
  AOI22_X1   g19258(.A1(new_n19450_), .A2(new_n18806_), .B1(\asqrt[9] ), .B2(new_n19448_), .ZN(new_n19451_));
  NAND2_X1   g19259(.A1(new_n19313_), .A2(new_n327_), .ZN(new_n19452_));
  INV_X1     g19260(.I(new_n19452_), .ZN(new_n19453_));
  AOI21_X1   g19261(.A1(new_n19453_), .A2(new_n19446_), .B(new_n19451_), .ZN(new_n19454_));
  OAI21_X1   g19262(.A1(new_n19454_), .A2(new_n19447_), .B(\asqrt[60] ), .ZN(new_n19455_));
  INV_X1     g19263(.I(new_n18725_), .ZN(new_n19456_));
  NOR2_X1    g19264(.A1(new_n18737_), .A2(new_n18724_), .ZN(new_n19457_));
  NOR3_X1    g19265(.A1(new_n18792_), .A2(new_n19456_), .A3(new_n19457_), .ZN(new_n19458_));
  INV_X1     g19266(.I(new_n19458_), .ZN(new_n19459_));
  NOR3_X1    g19267(.A1(new_n19456_), .A2(new_n18731_), .A3(new_n19457_), .ZN(new_n19460_));
  AOI22_X1   g19268(.A1(new_n19459_), .A2(new_n18731_), .B1(\asqrt[9] ), .B2(new_n19460_), .ZN(new_n19461_));
  INV_X1     g19269(.I(new_n19461_), .ZN(new_n19462_));
  INV_X1     g19270(.I(new_n19313_), .ZN(new_n19463_));
  NOR3_X1    g19271(.A1(new_n19312_), .A2(new_n19303_), .A3(\asqrt[58] ), .ZN(new_n19464_));
  NOR2_X1    g19272(.A1(new_n19464_), .A2(new_n19318_), .ZN(new_n19465_));
  OAI21_X1   g19273(.A1(new_n19465_), .A2(new_n19463_), .B(\asqrt[59] ), .ZN(new_n19466_));
  NAND2_X1   g19274(.A1(new_n19466_), .A2(new_n306_), .ZN(new_n19467_));
  OAI21_X1   g19275(.A1(new_n19467_), .A2(new_n19454_), .B(new_n19462_), .ZN(new_n19468_));
  AOI21_X1   g19276(.A1(new_n19468_), .A2(new_n19455_), .B(new_n218_), .ZN(new_n19469_));
  NOR2_X1    g19277(.A1(new_n18741_), .A2(new_n18748_), .ZN(new_n19470_));
  NOR3_X1    g19278(.A1(new_n19470_), .A2(new_n18739_), .A3(new_n18747_), .ZN(new_n19471_));
  NOR3_X1    g19279(.A1(new_n18792_), .A2(new_n18739_), .A3(new_n19470_), .ZN(new_n19472_));
  INV_X1     g19280(.I(new_n19472_), .ZN(new_n19473_));
  AOI22_X1   g19281(.A1(new_n19473_), .A2(new_n18747_), .B1(\asqrt[9] ), .B2(new_n19471_), .ZN(new_n19474_));
  INV_X1     g19282(.I(new_n19451_), .ZN(new_n19475_));
  OAI21_X1   g19283(.A1(new_n19465_), .A2(new_n19452_), .B(new_n19475_), .ZN(new_n19476_));
  AOI21_X1   g19284(.A1(new_n19476_), .A2(new_n19466_), .B(new_n306_), .ZN(new_n19477_));
  NOR2_X1    g19285(.A1(new_n19477_), .A2(\asqrt[61] ), .ZN(new_n19478_));
  AOI21_X1   g19286(.A1(new_n19478_), .A2(new_n19468_), .B(new_n19474_), .ZN(new_n19479_));
  OAI21_X1   g19287(.A1(new_n19479_), .A2(new_n19469_), .B(\asqrt[62] ), .ZN(new_n19480_));
  NOR3_X1    g19288(.A1(new_n18792_), .A2(new_n18750_), .A3(new_n18803_), .ZN(new_n19481_));
  INV_X1     g19289(.I(new_n19481_), .ZN(new_n19482_));
  NOR3_X1    g19290(.A1(new_n18750_), .A2(new_n18805_), .A3(new_n18803_), .ZN(new_n19483_));
  AOI22_X1   g19291(.A1(new_n19482_), .A2(new_n18805_), .B1(\asqrt[9] ), .B2(new_n19483_), .ZN(new_n19484_));
  INV_X1     g19292(.I(new_n19484_), .ZN(new_n19485_));
  OAI21_X1   g19293(.A1(new_n19318_), .A2(new_n19464_), .B(new_n19313_), .ZN(new_n19486_));
  AOI21_X1   g19294(.A1(new_n19486_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n19487_));
  AOI21_X1   g19295(.A1(new_n19487_), .A2(new_n19476_), .B(new_n19461_), .ZN(new_n19488_));
  OAI21_X1   g19296(.A1(new_n19488_), .A2(new_n19477_), .B(\asqrt[61] ), .ZN(new_n19489_));
  NAND2_X1   g19297(.A1(new_n19489_), .A2(new_n207_), .ZN(new_n19490_));
  OAI21_X1   g19298(.A1(new_n19490_), .A2(new_n19479_), .B(new_n19485_), .ZN(new_n19491_));
  NAND4_X1   g19299(.A1(\asqrt[9] ), .A2(new_n18757_), .A3(new_n18762_), .A4(new_n18842_), .ZN(new_n19492_));
  NAND2_X1   g19300(.A1(new_n18757_), .A2(new_n18842_), .ZN(new_n19493_));
  OAI21_X1   g19301(.A1(new_n18792_), .A2(new_n19493_), .B(new_n18763_), .ZN(new_n19494_));
  NAND2_X1   g19302(.A1(new_n19492_), .A2(new_n19494_), .ZN(new_n19495_));
  NOR2_X1    g19303(.A1(new_n18843_), .A2(new_n18782_), .ZN(new_n19496_));
  NAND2_X1   g19304(.A1(\asqrt[9] ), .A2(new_n19496_), .ZN(new_n19497_));
  NAND3_X1   g19305(.A1(new_n19495_), .A2(new_n18854_), .A3(new_n19497_), .ZN(new_n19498_));
  AOI21_X1   g19306(.A1(new_n19491_), .A2(new_n19480_), .B(new_n19498_), .ZN(new_n19499_));
  NOR3_X1    g19307(.A1(new_n19488_), .A2(new_n19477_), .A3(\asqrt[61] ), .ZN(new_n19500_));
  OAI21_X1   g19308(.A1(new_n19474_), .A2(new_n19500_), .B(new_n19489_), .ZN(new_n19501_));
  AOI21_X1   g19309(.A1(new_n19501_), .A2(\asqrt[62] ), .B(new_n19495_), .ZN(new_n19502_));
  OAI21_X1   g19310(.A1(new_n18792_), .A2(new_n18782_), .B(new_n18843_), .ZN(new_n19503_));
  NOR2_X1    g19311(.A1(new_n19496_), .A2(new_n193_), .ZN(new_n19504_));
  NAND2_X1   g19312(.A1(new_n19503_), .A2(new_n19504_), .ZN(new_n19505_));
  INV_X1     g19313(.I(new_n19505_), .ZN(new_n19506_));
  AND3_X2    g19314(.A1(new_n18774_), .A2(new_n18772_), .A3(new_n18788_), .Z(new_n19507_));
  NAND4_X1   g19315(.A1(new_n18844_), .A2(new_n18854_), .A3(new_n18785_), .A4(new_n19507_), .ZN(new_n19508_));
  INV_X1     g19316(.I(new_n19508_), .ZN(new_n19509_));
  NOR2_X1    g19317(.A1(new_n19506_), .A2(new_n19509_), .ZN(new_n19510_));
  INV_X1     g19318(.I(new_n19510_), .ZN(new_n19511_));
  AOI21_X1   g19319(.A1(new_n19502_), .A2(new_n19491_), .B(new_n19511_), .ZN(new_n19512_));
  OAI21_X1   g19320(.A1(\asqrt[63] ), .A2(new_n19499_), .B(new_n19512_), .ZN(\asqrt[8] ));
  NOR2_X1    g19321(.A1(\a[14] ), .A2(\a[15] ), .ZN(new_n19514_));
  INV_X1     g19322(.I(new_n19514_), .ZN(new_n19515_));
  NOR2_X1    g19323(.A1(new_n19515_), .A2(\a[16] ), .ZN(new_n19516_));
  INV_X1     g19324(.I(new_n19516_), .ZN(new_n19517_));
  NAND2_X1   g19325(.A1(new_n19491_), .A2(new_n19480_), .ZN(new_n19518_));
  INV_X1     g19326(.I(new_n19498_), .ZN(new_n19519_));
  AOI21_X1   g19327(.A1(new_n19518_), .A2(new_n19519_), .B(\asqrt[63] ), .ZN(new_n19520_));
  INV_X1     g19328(.I(new_n19474_), .ZN(new_n19521_));
  NAND3_X1   g19329(.A1(new_n19446_), .A2(new_n327_), .A3(new_n19313_), .ZN(new_n19522_));
  AOI22_X1   g19330(.A1(new_n19522_), .A2(new_n19475_), .B1(new_n19486_), .B2(\asqrt[59] ), .ZN(new_n19523_));
  OAI21_X1   g19331(.A1(new_n19523_), .A2(new_n306_), .B(new_n218_), .ZN(new_n19524_));
  OAI21_X1   g19332(.A1(new_n19524_), .A2(new_n19488_), .B(new_n19521_), .ZN(new_n19525_));
  NOR2_X1    g19333(.A1(new_n19469_), .A2(\asqrt[62] ), .ZN(new_n19526_));
  AOI21_X1   g19334(.A1(new_n19526_), .A2(new_n19525_), .B(new_n19484_), .ZN(new_n19527_));
  INV_X1     g19335(.I(new_n19495_), .ZN(new_n19528_));
  NAND2_X1   g19336(.A1(new_n19480_), .A2(new_n19528_), .ZN(new_n19529_));
  OAI21_X1   g19337(.A1(new_n19529_), .A2(new_n19527_), .B(new_n19510_), .ZN(new_n19530_));
  OAI21_X1   g19338(.A1(new_n19520_), .A2(new_n19530_), .B(\a[16] ), .ZN(new_n19531_));
  AOI21_X1   g19339(.A1(new_n19531_), .A2(new_n19517_), .B(new_n18792_), .ZN(new_n19532_));
  INV_X1     g19340(.I(\a[16] ), .ZN(new_n19533_));
  NAND3_X1   g19341(.A1(new_n19525_), .A2(new_n207_), .A3(new_n19489_), .ZN(new_n19534_));
  AOI22_X1   g19342(.A1(new_n19534_), .A2(new_n19485_), .B1(new_n19501_), .B2(\asqrt[62] ), .ZN(new_n19535_));
  OAI21_X1   g19343(.A1(new_n19535_), .A2(new_n19498_), .B(new_n193_), .ZN(new_n19536_));
  AOI21_X1   g19344(.A1(new_n19536_), .A2(new_n19512_), .B(new_n19533_), .ZN(new_n19537_));
  NAND4_X1   g19345(.A1(new_n18854_), .A2(new_n18785_), .A3(new_n18788_), .A4(new_n19517_), .ZN(new_n19538_));
  NOR2_X1    g19346(.A1(new_n19538_), .A2(new_n18780_), .ZN(new_n19539_));
  INV_X1     g19347(.I(new_n19539_), .ZN(new_n19540_));
  NOR2_X1    g19348(.A1(new_n19537_), .A2(new_n19540_), .ZN(new_n19541_));
  AOI21_X1   g19349(.A1(new_n19536_), .A2(new_n19512_), .B(new_n18795_), .ZN(new_n19542_));
  INV_X1     g19350(.I(\a[17] ), .ZN(new_n19543_));
  AOI21_X1   g19351(.A1(\asqrt[8] ), .A2(new_n19533_), .B(new_n19543_), .ZN(new_n19544_));
  NOR3_X1    g19352(.A1(new_n19541_), .A2(new_n19544_), .A3(new_n19542_), .ZN(new_n19545_));
  OAI21_X1   g19353(.A1(new_n19545_), .A2(new_n19532_), .B(\asqrt[10] ), .ZN(new_n19546_));
  OAI21_X1   g19354(.A1(new_n19520_), .A2(new_n19530_), .B(new_n18794_), .ZN(new_n19547_));
  NAND2_X1   g19355(.A1(new_n19502_), .A2(new_n19491_), .ZN(new_n19548_));
  NOR3_X1    g19356(.A1(new_n19506_), .A2(new_n18792_), .A3(new_n19509_), .ZN(new_n19549_));
  NAND3_X1   g19357(.A1(new_n19536_), .A2(new_n19548_), .A3(new_n19549_), .ZN(new_n19550_));
  AOI21_X1   g19358(.A1(new_n19550_), .A2(new_n19547_), .B(new_n18793_), .ZN(new_n19551_));
  NAND2_X1   g19359(.A1(new_n19548_), .A2(new_n19549_), .ZN(new_n19552_));
  NOR2_X1    g19360(.A1(new_n19552_), .A2(new_n19520_), .ZN(new_n19553_));
  NOR3_X1    g19361(.A1(new_n19553_), .A2(new_n19542_), .A3(\a[18] ), .ZN(new_n19554_));
  AOI21_X1   g19362(.A1(\asqrt[8] ), .A2(\a[16] ), .B(new_n19516_), .ZN(new_n19555_));
  OAI21_X1   g19363(.A1(new_n19555_), .A2(new_n18792_), .B(new_n18275_), .ZN(new_n19556_));
  OAI22_X1   g19364(.A1(new_n19545_), .A2(new_n19556_), .B1(new_n19551_), .B2(new_n19554_), .ZN(new_n19557_));
  AOI21_X1   g19365(.A1(new_n19557_), .A2(new_n19546_), .B(new_n17623_), .ZN(new_n19558_));
  NOR3_X1    g19366(.A1(new_n18883_), .A2(new_n18884_), .A3(new_n18849_), .ZN(new_n19559_));
  NAND3_X1   g19367(.A1(\asqrt[8] ), .A2(new_n18882_), .A3(new_n18802_), .ZN(new_n19560_));
  AOI22_X1   g19368(.A1(new_n19560_), .A2(new_n18849_), .B1(\asqrt[8] ), .B2(new_n19559_), .ZN(new_n19561_));
  OAI21_X1   g19369(.A1(new_n19537_), .A2(new_n19516_), .B(\asqrt[9] ), .ZN(new_n19562_));
  AOI21_X1   g19370(.A1(new_n19536_), .A2(new_n19512_), .B(\a[16] ), .ZN(new_n19563_));
  OAI21_X1   g19371(.A1(new_n19543_), .A2(new_n19563_), .B(new_n19547_), .ZN(new_n19564_));
  OAI21_X1   g19372(.A1(new_n19564_), .A2(new_n19541_), .B(new_n19562_), .ZN(new_n19565_));
  AOI21_X1   g19373(.A1(new_n19565_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n19566_));
  AOI21_X1   g19374(.A1(new_n19566_), .A2(new_n19557_), .B(new_n19561_), .ZN(new_n19567_));
  OAI21_X1   g19375(.A1(new_n19567_), .A2(new_n19558_), .B(\asqrt[12] ), .ZN(new_n19568_));
  INV_X1     g19376(.I(new_n19568_), .ZN(new_n19569_));
  NOR2_X1    g19377(.A1(new_n18887_), .A2(new_n18890_), .ZN(new_n19570_));
  INV_X1     g19378(.I(new_n19570_), .ZN(new_n19571_));
  NAND4_X1   g19379(.A1(\asqrt[8] ), .A2(new_n18888_), .A3(new_n18862_), .A4(new_n19571_), .ZN(new_n19572_));
  INV_X1     g19380(.I(\asqrt[8] ), .ZN(new_n19573_));
  NOR3_X1    g19381(.A1(new_n19573_), .A2(new_n18851_), .A3(new_n19570_), .ZN(new_n19574_));
  OAI21_X1   g19382(.A1(new_n19574_), .A2(new_n18862_), .B(new_n19572_), .ZN(new_n19575_));
  INV_X1     g19383(.I(new_n19575_), .ZN(new_n19576_));
  NOR3_X1    g19384(.A1(new_n19567_), .A2(new_n19558_), .A3(\asqrt[12] ), .ZN(new_n19577_));
  NOR2_X1    g19385(.A1(new_n19577_), .A2(new_n19576_), .ZN(new_n19578_));
  OAI21_X1   g19386(.A1(new_n19578_), .A2(new_n19569_), .B(\asqrt[13] ), .ZN(new_n19579_));
  NAND2_X1   g19387(.A1(new_n18896_), .A2(new_n18891_), .ZN(new_n19580_));
  NAND3_X1   g19388(.A1(\asqrt[8] ), .A2(new_n18865_), .A3(new_n19580_), .ZN(new_n19581_));
  AND3_X2    g19389(.A1(new_n18865_), .A2(new_n18869_), .A3(new_n19580_), .Z(new_n19582_));
  AOI22_X1   g19390(.A1(new_n19581_), .A2(new_n18870_), .B1(\asqrt[8] ), .B2(new_n19582_), .ZN(new_n19583_));
  INV_X1     g19391(.I(new_n19583_), .ZN(new_n19584_));
  NAND2_X1   g19392(.A1(new_n19568_), .A2(new_n16389_), .ZN(new_n19585_));
  OAI21_X1   g19393(.A1(new_n19578_), .A2(new_n19585_), .B(new_n19584_), .ZN(new_n19586_));
  AOI21_X1   g19394(.A1(new_n19586_), .A2(new_n19579_), .B(new_n15770_), .ZN(new_n19587_));
  NOR3_X1    g19395(.A1(new_n18873_), .A2(new_n18879_), .A3(new_n18898_), .ZN(new_n19588_));
  NOR3_X1    g19396(.A1(new_n19573_), .A2(new_n18873_), .A3(new_n18898_), .ZN(new_n19589_));
  INV_X1     g19397(.I(new_n19589_), .ZN(new_n19590_));
  AOI22_X1   g19398(.A1(new_n19590_), .A2(new_n18879_), .B1(\asqrt[8] ), .B2(new_n19588_), .ZN(new_n19591_));
  OAI21_X1   g19399(.A1(new_n19576_), .A2(new_n19577_), .B(new_n19568_), .ZN(new_n19592_));
  AOI21_X1   g19400(.A1(new_n19592_), .A2(\asqrt[13] ), .B(\asqrt[14] ), .ZN(new_n19593_));
  AOI21_X1   g19401(.A1(new_n19593_), .A2(new_n19586_), .B(new_n19591_), .ZN(new_n19594_));
  OAI21_X1   g19402(.A1(new_n19594_), .A2(new_n19587_), .B(\asqrt[15] ), .ZN(new_n19595_));
  INV_X1     g19403(.I(new_n19595_), .ZN(new_n19596_));
  NAND2_X1   g19404(.A1(new_n19337_), .A2(new_n19335_), .ZN(new_n19597_));
  NAND3_X1   g19405(.A1(\asqrt[8] ), .A2(new_n18900_), .A3(new_n19597_), .ZN(new_n19598_));
  AND3_X2    g19406(.A1(new_n19597_), .A2(new_n18900_), .A3(new_n18905_), .Z(new_n19599_));
  AOI22_X1   g19407(.A1(new_n19598_), .A2(new_n18906_), .B1(\asqrt[8] ), .B2(new_n19599_), .ZN(new_n19600_));
  NOR3_X1    g19408(.A1(new_n19594_), .A2(new_n19587_), .A3(\asqrt[15] ), .ZN(new_n19601_));
  NOR2_X1    g19409(.A1(new_n19601_), .A2(new_n19600_), .ZN(new_n19602_));
  OAI21_X1   g19410(.A1(new_n19602_), .A2(new_n19596_), .B(\asqrt[16] ), .ZN(new_n19603_));
  INV_X1     g19411(.I(new_n18914_), .ZN(new_n19604_));
  NOR3_X1    g19412(.A1(new_n19348_), .A2(new_n18910_), .A3(new_n19604_), .ZN(new_n19605_));
  NOR3_X1    g19413(.A1(new_n19573_), .A2(new_n18910_), .A3(new_n19348_), .ZN(new_n19606_));
  INV_X1     g19414(.I(new_n19606_), .ZN(new_n19607_));
  AOI22_X1   g19415(.A1(new_n19607_), .A2(new_n19604_), .B1(\asqrt[8] ), .B2(new_n19605_), .ZN(new_n19608_));
  INV_X1     g19416(.I(new_n19608_), .ZN(new_n19609_));
  NAND2_X1   g19417(.A1(new_n19595_), .A2(new_n14601_), .ZN(new_n19610_));
  OAI21_X1   g19418(.A1(new_n19602_), .A2(new_n19610_), .B(new_n19609_), .ZN(new_n19611_));
  AOI21_X1   g19419(.A1(new_n19611_), .A2(new_n19603_), .B(new_n14017_), .ZN(new_n19612_));
  NOR3_X1    g19420(.A1(new_n19573_), .A2(new_n18919_), .A3(new_n18924_), .ZN(new_n19613_));
  INV_X1     g19421(.I(new_n19613_), .ZN(new_n19614_));
  NOR3_X1    g19422(.A1(new_n18919_), .A2(new_n19333_), .A3(new_n18924_), .ZN(new_n19615_));
  AOI22_X1   g19423(.A1(new_n19614_), .A2(new_n19333_), .B1(\asqrt[8] ), .B2(new_n19615_), .ZN(new_n19616_));
  OAI21_X1   g19424(.A1(new_n19600_), .A2(new_n19601_), .B(new_n19595_), .ZN(new_n19617_));
  AOI21_X1   g19425(.A1(new_n19617_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n19618_));
  AOI21_X1   g19426(.A1(new_n19618_), .A2(new_n19611_), .B(new_n19616_), .ZN(new_n19619_));
  OAI21_X1   g19427(.A1(new_n19619_), .A2(new_n19612_), .B(\asqrt[18] ), .ZN(new_n19620_));
  INV_X1     g19428(.I(new_n19620_), .ZN(new_n19621_));
  AND3_X2    g19429(.A1(new_n18926_), .A2(new_n18931_), .A3(new_n19342_), .Z(new_n19622_));
  NAND3_X1   g19430(.A1(\asqrt[8] ), .A2(new_n18926_), .A3(new_n19342_), .ZN(new_n19623_));
  AOI22_X1   g19431(.A1(new_n19623_), .A2(new_n18932_), .B1(\asqrt[8] ), .B2(new_n19622_), .ZN(new_n19624_));
  NOR3_X1    g19432(.A1(new_n19619_), .A2(new_n19612_), .A3(\asqrt[18] ), .ZN(new_n19625_));
  NOR2_X1    g19433(.A1(new_n19625_), .A2(new_n19624_), .ZN(new_n19626_));
  OAI21_X1   g19434(.A1(new_n19626_), .A2(new_n19621_), .B(\asqrt[19] ), .ZN(new_n19627_));
  INV_X1     g19435(.I(new_n18939_), .ZN(new_n19628_));
  NOR3_X1    g19436(.A1(new_n19573_), .A2(new_n18935_), .A3(new_n19352_), .ZN(new_n19629_));
  INV_X1     g19437(.I(new_n19629_), .ZN(new_n19630_));
  NOR3_X1    g19438(.A1(new_n19352_), .A2(new_n18935_), .A3(new_n19628_), .ZN(new_n19631_));
  AOI22_X1   g19439(.A1(new_n19630_), .A2(new_n19628_), .B1(\asqrt[8] ), .B2(new_n19631_), .ZN(new_n19632_));
  INV_X1     g19440(.I(new_n19632_), .ZN(new_n19633_));
  NAND2_X1   g19441(.A1(new_n19620_), .A2(new_n12913_), .ZN(new_n19634_));
  OAI21_X1   g19442(.A1(new_n19626_), .A2(new_n19634_), .B(new_n19633_), .ZN(new_n19635_));
  AOI21_X1   g19443(.A1(new_n19635_), .A2(new_n19627_), .B(new_n12364_), .ZN(new_n19636_));
  NOR3_X1    g19444(.A1(new_n18944_), .A2(new_n19332_), .A3(new_n18950_), .ZN(new_n19637_));
  NOR3_X1    g19445(.A1(new_n19573_), .A2(new_n18944_), .A3(new_n18950_), .ZN(new_n19638_));
  INV_X1     g19446(.I(new_n19638_), .ZN(new_n19639_));
  AOI22_X1   g19447(.A1(new_n19639_), .A2(new_n19332_), .B1(\asqrt[8] ), .B2(new_n19637_), .ZN(new_n19640_));
  OAI21_X1   g19448(.A1(new_n19624_), .A2(new_n19625_), .B(new_n19620_), .ZN(new_n19641_));
  AOI21_X1   g19449(.A1(new_n19641_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n19642_));
  AOI21_X1   g19450(.A1(new_n19642_), .A2(new_n19635_), .B(new_n19640_), .ZN(new_n19643_));
  OAI21_X1   g19451(.A1(new_n19643_), .A2(new_n19636_), .B(\asqrt[21] ), .ZN(new_n19644_));
  INV_X1     g19452(.I(new_n19644_), .ZN(new_n19645_));
  NOR2_X1    g19453(.A1(new_n18951_), .A2(new_n18959_), .ZN(new_n19646_));
  NOR3_X1    g19454(.A1(new_n19573_), .A2(new_n19346_), .A3(new_n19646_), .ZN(new_n19647_));
  INV_X1     g19455(.I(new_n19647_), .ZN(new_n19648_));
  NOR3_X1    g19456(.A1(new_n19646_), .A2(new_n19346_), .A3(new_n18958_), .ZN(new_n19649_));
  AOI22_X1   g19457(.A1(new_n19648_), .A2(new_n18958_), .B1(\asqrt[8] ), .B2(new_n19649_), .ZN(new_n19650_));
  NOR3_X1    g19458(.A1(new_n19643_), .A2(new_n19636_), .A3(\asqrt[21] ), .ZN(new_n19651_));
  NOR2_X1    g19459(.A1(new_n19651_), .A2(new_n19650_), .ZN(new_n19652_));
  OAI21_X1   g19460(.A1(new_n19652_), .A2(new_n19645_), .B(\asqrt[22] ), .ZN(new_n19653_));
  INV_X1     g19461(.I(new_n18967_), .ZN(new_n19654_));
  NOR3_X1    g19462(.A1(new_n19360_), .A2(new_n18961_), .A3(new_n19654_), .ZN(new_n19655_));
  NOR3_X1    g19463(.A1(new_n19573_), .A2(new_n18961_), .A3(new_n19360_), .ZN(new_n19656_));
  INV_X1     g19464(.I(new_n19656_), .ZN(new_n19657_));
  AOI22_X1   g19465(.A1(new_n19657_), .A2(new_n19654_), .B1(\asqrt[8] ), .B2(new_n19655_), .ZN(new_n19658_));
  INV_X1     g19466(.I(new_n19658_), .ZN(new_n19659_));
  NAND2_X1   g19467(.A1(new_n19644_), .A2(new_n11326_), .ZN(new_n19660_));
  OAI21_X1   g19468(.A1(new_n19652_), .A2(new_n19660_), .B(new_n19659_), .ZN(new_n19661_));
  AOI21_X1   g19469(.A1(new_n19661_), .A2(new_n19653_), .B(new_n10812_), .ZN(new_n19662_));
  NOR3_X1    g19470(.A1(new_n19573_), .A2(new_n18972_), .A3(new_n18981_), .ZN(new_n19663_));
  INV_X1     g19471(.I(new_n19663_), .ZN(new_n19664_));
  NOR3_X1    g19472(.A1(new_n18972_), .A2(new_n19331_), .A3(new_n18981_), .ZN(new_n19665_));
  AOI22_X1   g19473(.A1(new_n19664_), .A2(new_n19331_), .B1(\asqrt[8] ), .B2(new_n19665_), .ZN(new_n19666_));
  OAI21_X1   g19474(.A1(new_n19650_), .A2(new_n19651_), .B(new_n19644_), .ZN(new_n19667_));
  AOI21_X1   g19475(.A1(new_n19667_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n19668_));
  AOI21_X1   g19476(.A1(new_n19668_), .A2(new_n19661_), .B(new_n19666_), .ZN(new_n19669_));
  OAI21_X1   g19477(.A1(new_n19669_), .A2(new_n19662_), .B(\asqrt[24] ), .ZN(new_n19670_));
  INV_X1     g19478(.I(new_n19670_), .ZN(new_n19671_));
  NOR2_X1    g19479(.A1(new_n18982_), .A2(new_n18990_), .ZN(new_n19672_));
  NOR3_X1    g19480(.A1(new_n19672_), .A2(new_n19359_), .A3(new_n18989_), .ZN(new_n19673_));
  NOR3_X1    g19481(.A1(new_n19573_), .A2(new_n19359_), .A3(new_n19672_), .ZN(new_n19674_));
  INV_X1     g19482(.I(new_n19674_), .ZN(new_n19675_));
  AOI22_X1   g19483(.A1(new_n19675_), .A2(new_n18989_), .B1(\asqrt[8] ), .B2(new_n19673_), .ZN(new_n19676_));
  NOR3_X1    g19484(.A1(new_n19669_), .A2(new_n19662_), .A3(\asqrt[24] ), .ZN(new_n19677_));
  NOR2_X1    g19485(.A1(new_n19677_), .A2(new_n19676_), .ZN(new_n19678_));
  OAI21_X1   g19486(.A1(new_n19678_), .A2(new_n19671_), .B(\asqrt[25] ), .ZN(new_n19679_));
  INV_X1     g19487(.I(new_n18997_), .ZN(new_n19680_));
  NOR3_X1    g19488(.A1(new_n19573_), .A2(new_n18992_), .A3(new_n19368_), .ZN(new_n19681_));
  INV_X1     g19489(.I(new_n19681_), .ZN(new_n19682_));
  NOR3_X1    g19490(.A1(new_n19368_), .A2(new_n18992_), .A3(new_n19680_), .ZN(new_n19683_));
  AOI22_X1   g19491(.A1(new_n19682_), .A2(new_n19680_), .B1(\asqrt[8] ), .B2(new_n19683_), .ZN(new_n19684_));
  INV_X1     g19492(.I(new_n19684_), .ZN(new_n19685_));
  NAND2_X1   g19493(.A1(new_n19670_), .A2(new_n9846_), .ZN(new_n19686_));
  OAI21_X1   g19494(.A1(new_n19678_), .A2(new_n19686_), .B(new_n19685_), .ZN(new_n19687_));
  AOI21_X1   g19495(.A1(new_n19687_), .A2(new_n19679_), .B(new_n9317_), .ZN(new_n19688_));
  NOR3_X1    g19496(.A1(new_n19002_), .A2(new_n19330_), .A3(new_n19011_), .ZN(new_n19689_));
  NOR3_X1    g19497(.A1(new_n19573_), .A2(new_n19002_), .A3(new_n19011_), .ZN(new_n19690_));
  INV_X1     g19498(.I(new_n19690_), .ZN(new_n19691_));
  AOI22_X1   g19499(.A1(new_n19691_), .A2(new_n19330_), .B1(\asqrt[8] ), .B2(new_n19689_), .ZN(new_n19692_));
  OAI21_X1   g19500(.A1(new_n19676_), .A2(new_n19677_), .B(new_n19670_), .ZN(new_n19693_));
  AOI21_X1   g19501(.A1(new_n19693_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n19694_));
  AOI21_X1   g19502(.A1(new_n19694_), .A2(new_n19687_), .B(new_n19692_), .ZN(new_n19695_));
  OAI21_X1   g19503(.A1(new_n19695_), .A2(new_n19688_), .B(\asqrt[27] ), .ZN(new_n19696_));
  INV_X1     g19504(.I(new_n19696_), .ZN(new_n19697_));
  NOR2_X1    g19505(.A1(new_n19012_), .A2(new_n19020_), .ZN(new_n19698_));
  NOR3_X1    g19506(.A1(new_n19573_), .A2(new_n19367_), .A3(new_n19698_), .ZN(new_n19699_));
  INV_X1     g19507(.I(new_n19699_), .ZN(new_n19700_));
  NOR3_X1    g19508(.A1(new_n19698_), .A2(new_n19367_), .A3(new_n19019_), .ZN(new_n19701_));
  AOI22_X1   g19509(.A1(new_n19700_), .A2(new_n19019_), .B1(\asqrt[8] ), .B2(new_n19701_), .ZN(new_n19702_));
  NOR3_X1    g19510(.A1(new_n19695_), .A2(new_n19688_), .A3(\asqrt[27] ), .ZN(new_n19703_));
  NOR2_X1    g19511(.A1(new_n19703_), .A2(new_n19702_), .ZN(new_n19704_));
  OAI21_X1   g19512(.A1(new_n19704_), .A2(new_n19697_), .B(\asqrt[28] ), .ZN(new_n19705_));
  INV_X1     g19513(.I(new_n19027_), .ZN(new_n19706_));
  NOR3_X1    g19514(.A1(new_n19376_), .A2(new_n19022_), .A3(new_n19706_), .ZN(new_n19707_));
  NOR3_X1    g19515(.A1(new_n19573_), .A2(new_n19022_), .A3(new_n19376_), .ZN(new_n19708_));
  INV_X1     g19516(.I(new_n19708_), .ZN(new_n19709_));
  AOI22_X1   g19517(.A1(new_n19709_), .A2(new_n19706_), .B1(\asqrt[8] ), .B2(new_n19707_), .ZN(new_n19710_));
  INV_X1     g19518(.I(new_n19710_), .ZN(new_n19711_));
  NAND2_X1   g19519(.A1(new_n19696_), .A2(new_n8483_), .ZN(new_n19712_));
  OAI21_X1   g19520(.A1(new_n19704_), .A2(new_n19712_), .B(new_n19711_), .ZN(new_n19713_));
  AOI21_X1   g19521(.A1(new_n19713_), .A2(new_n19705_), .B(new_n8036_), .ZN(new_n19714_));
  NOR3_X1    g19522(.A1(new_n19573_), .A2(new_n19032_), .A3(new_n19041_), .ZN(new_n19715_));
  INV_X1     g19523(.I(new_n19715_), .ZN(new_n19716_));
  NOR3_X1    g19524(.A1(new_n19032_), .A2(new_n19329_), .A3(new_n19041_), .ZN(new_n19717_));
  AOI22_X1   g19525(.A1(new_n19716_), .A2(new_n19329_), .B1(\asqrt[8] ), .B2(new_n19717_), .ZN(new_n19718_));
  OAI21_X1   g19526(.A1(new_n19702_), .A2(new_n19703_), .B(new_n19696_), .ZN(new_n19719_));
  AOI21_X1   g19527(.A1(new_n19719_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n19720_));
  AOI21_X1   g19528(.A1(new_n19720_), .A2(new_n19713_), .B(new_n19718_), .ZN(new_n19721_));
  OAI21_X1   g19529(.A1(new_n19721_), .A2(new_n19714_), .B(\asqrt[30] ), .ZN(new_n19722_));
  INV_X1     g19530(.I(new_n19722_), .ZN(new_n19723_));
  NOR2_X1    g19531(.A1(new_n19042_), .A2(new_n19050_), .ZN(new_n19724_));
  NOR3_X1    g19532(.A1(new_n19724_), .A2(new_n19375_), .A3(new_n19049_), .ZN(new_n19725_));
  NOR3_X1    g19533(.A1(new_n19573_), .A2(new_n19375_), .A3(new_n19724_), .ZN(new_n19726_));
  INV_X1     g19534(.I(new_n19726_), .ZN(new_n19727_));
  AOI22_X1   g19535(.A1(new_n19727_), .A2(new_n19049_), .B1(\asqrt[8] ), .B2(new_n19725_), .ZN(new_n19728_));
  NOR3_X1    g19536(.A1(new_n19721_), .A2(new_n19714_), .A3(\asqrt[30] ), .ZN(new_n19729_));
  NOR2_X1    g19537(.A1(new_n19729_), .A2(new_n19728_), .ZN(new_n19730_));
  OAI21_X1   g19538(.A1(new_n19730_), .A2(new_n19723_), .B(\asqrt[31] ), .ZN(new_n19731_));
  INV_X1     g19539(.I(new_n19057_), .ZN(new_n19732_));
  NOR3_X1    g19540(.A1(new_n19573_), .A2(new_n19052_), .A3(new_n19384_), .ZN(new_n19733_));
  INV_X1     g19541(.I(new_n19733_), .ZN(new_n19734_));
  NOR3_X1    g19542(.A1(new_n19384_), .A2(new_n19052_), .A3(new_n19732_), .ZN(new_n19735_));
  AOI22_X1   g19543(.A1(new_n19734_), .A2(new_n19732_), .B1(\asqrt[8] ), .B2(new_n19735_), .ZN(new_n19736_));
  INV_X1     g19544(.I(new_n19736_), .ZN(new_n19737_));
  NAND2_X1   g19545(.A1(new_n19722_), .A2(new_n7229_), .ZN(new_n19738_));
  OAI21_X1   g19546(.A1(new_n19730_), .A2(new_n19738_), .B(new_n19737_), .ZN(new_n19739_));
  AOI21_X1   g19547(.A1(new_n19739_), .A2(new_n19731_), .B(new_n6824_), .ZN(new_n19740_));
  NOR3_X1    g19548(.A1(new_n19062_), .A2(new_n19328_), .A3(new_n19068_), .ZN(new_n19741_));
  NOR3_X1    g19549(.A1(new_n19573_), .A2(new_n19062_), .A3(new_n19068_), .ZN(new_n19742_));
  INV_X1     g19550(.I(new_n19742_), .ZN(new_n19743_));
  AOI22_X1   g19551(.A1(new_n19743_), .A2(new_n19328_), .B1(\asqrt[8] ), .B2(new_n19741_), .ZN(new_n19744_));
  OAI21_X1   g19552(.A1(new_n19728_), .A2(new_n19729_), .B(new_n19722_), .ZN(new_n19745_));
  AOI21_X1   g19553(.A1(new_n19745_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n19746_));
  AOI21_X1   g19554(.A1(new_n19746_), .A2(new_n19739_), .B(new_n19744_), .ZN(new_n19747_));
  OAI21_X1   g19555(.A1(new_n19747_), .A2(new_n19740_), .B(\asqrt[33] ), .ZN(new_n19748_));
  INV_X1     g19556(.I(new_n19748_), .ZN(new_n19749_));
  NOR2_X1    g19557(.A1(new_n19069_), .A2(new_n19077_), .ZN(new_n19750_));
  NOR3_X1    g19558(.A1(new_n19573_), .A2(new_n19383_), .A3(new_n19750_), .ZN(new_n19751_));
  INV_X1     g19559(.I(new_n19751_), .ZN(new_n19752_));
  NOR3_X1    g19560(.A1(new_n19750_), .A2(new_n19383_), .A3(new_n19076_), .ZN(new_n19753_));
  AOI22_X1   g19561(.A1(new_n19752_), .A2(new_n19076_), .B1(\asqrt[8] ), .B2(new_n19753_), .ZN(new_n19754_));
  NOR3_X1    g19562(.A1(new_n19747_), .A2(new_n19740_), .A3(\asqrt[33] ), .ZN(new_n19755_));
  NOR2_X1    g19563(.A1(new_n19755_), .A2(new_n19754_), .ZN(new_n19756_));
  OAI21_X1   g19564(.A1(new_n19756_), .A2(new_n19749_), .B(\asqrt[34] ), .ZN(new_n19757_));
  INV_X1     g19565(.I(new_n19084_), .ZN(new_n19758_));
  NOR3_X1    g19566(.A1(new_n19392_), .A2(new_n19079_), .A3(new_n19758_), .ZN(new_n19759_));
  NOR3_X1    g19567(.A1(new_n19573_), .A2(new_n19079_), .A3(new_n19392_), .ZN(new_n19760_));
  INV_X1     g19568(.I(new_n19760_), .ZN(new_n19761_));
  AOI22_X1   g19569(.A1(new_n19761_), .A2(new_n19758_), .B1(\asqrt[8] ), .B2(new_n19759_), .ZN(new_n19762_));
  INV_X1     g19570(.I(new_n19762_), .ZN(new_n19763_));
  NAND2_X1   g19571(.A1(new_n19748_), .A2(new_n6077_), .ZN(new_n19764_));
  OAI21_X1   g19572(.A1(new_n19756_), .A2(new_n19764_), .B(new_n19763_), .ZN(new_n19765_));
  AOI21_X1   g19573(.A1(new_n19765_), .A2(new_n19757_), .B(new_n5708_), .ZN(new_n19766_));
  NOR3_X1    g19574(.A1(new_n19573_), .A2(new_n19089_), .A3(new_n19095_), .ZN(new_n19767_));
  INV_X1     g19575(.I(new_n19767_), .ZN(new_n19768_));
  NOR3_X1    g19576(.A1(new_n19089_), .A2(new_n19327_), .A3(new_n19095_), .ZN(new_n19769_));
  AOI22_X1   g19577(.A1(new_n19768_), .A2(new_n19327_), .B1(\asqrt[8] ), .B2(new_n19769_), .ZN(new_n19770_));
  OAI21_X1   g19578(.A1(new_n19754_), .A2(new_n19755_), .B(new_n19748_), .ZN(new_n19771_));
  AOI21_X1   g19579(.A1(new_n19771_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n19772_));
  AOI21_X1   g19580(.A1(new_n19772_), .A2(new_n19765_), .B(new_n19770_), .ZN(new_n19773_));
  OAI21_X1   g19581(.A1(new_n19773_), .A2(new_n19766_), .B(\asqrt[36] ), .ZN(new_n19774_));
  INV_X1     g19582(.I(new_n19774_), .ZN(new_n19775_));
  NOR2_X1    g19583(.A1(new_n19096_), .A2(new_n19104_), .ZN(new_n19776_));
  NOR3_X1    g19584(.A1(new_n19776_), .A2(new_n19391_), .A3(new_n19103_), .ZN(new_n19777_));
  NOR3_X1    g19585(.A1(new_n19573_), .A2(new_n19391_), .A3(new_n19776_), .ZN(new_n19778_));
  INV_X1     g19586(.I(new_n19778_), .ZN(new_n19779_));
  AOI22_X1   g19587(.A1(new_n19779_), .A2(new_n19103_), .B1(\asqrt[8] ), .B2(new_n19777_), .ZN(new_n19780_));
  NOR3_X1    g19588(.A1(new_n19773_), .A2(new_n19766_), .A3(\asqrt[36] ), .ZN(new_n19781_));
  NOR2_X1    g19589(.A1(new_n19781_), .A2(new_n19780_), .ZN(new_n19782_));
  OAI21_X1   g19590(.A1(new_n19782_), .A2(new_n19775_), .B(\asqrt[37] ), .ZN(new_n19783_));
  INV_X1     g19591(.I(new_n19111_), .ZN(new_n19784_));
  NOR3_X1    g19592(.A1(new_n19573_), .A2(new_n19106_), .A3(new_n19400_), .ZN(new_n19785_));
  INV_X1     g19593(.I(new_n19785_), .ZN(new_n19786_));
  NOR3_X1    g19594(.A1(new_n19400_), .A2(new_n19106_), .A3(new_n19784_), .ZN(new_n19787_));
  AOI22_X1   g19595(.A1(new_n19786_), .A2(new_n19784_), .B1(\asqrt[8] ), .B2(new_n19787_), .ZN(new_n19788_));
  INV_X1     g19596(.I(new_n19788_), .ZN(new_n19789_));
  NAND2_X1   g19597(.A1(new_n19774_), .A2(new_n5024_), .ZN(new_n19790_));
  OAI21_X1   g19598(.A1(new_n19782_), .A2(new_n19790_), .B(new_n19789_), .ZN(new_n19791_));
  AOI21_X1   g19599(.A1(new_n19791_), .A2(new_n19783_), .B(new_n4696_), .ZN(new_n19792_));
  NOR3_X1    g19600(.A1(new_n19116_), .A2(new_n19326_), .A3(new_n19122_), .ZN(new_n19793_));
  NOR3_X1    g19601(.A1(new_n19573_), .A2(new_n19116_), .A3(new_n19122_), .ZN(new_n19794_));
  INV_X1     g19602(.I(new_n19794_), .ZN(new_n19795_));
  AOI22_X1   g19603(.A1(new_n19795_), .A2(new_n19326_), .B1(\asqrt[8] ), .B2(new_n19793_), .ZN(new_n19796_));
  OAI21_X1   g19604(.A1(new_n19780_), .A2(new_n19781_), .B(new_n19774_), .ZN(new_n19797_));
  AOI21_X1   g19605(.A1(new_n19797_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n19798_));
  AOI21_X1   g19606(.A1(new_n19798_), .A2(new_n19791_), .B(new_n19796_), .ZN(new_n19799_));
  OAI21_X1   g19607(.A1(new_n19799_), .A2(new_n19792_), .B(\asqrt[39] ), .ZN(new_n19800_));
  INV_X1     g19608(.I(new_n19800_), .ZN(new_n19801_));
  NOR2_X1    g19609(.A1(new_n19123_), .A2(new_n19131_), .ZN(new_n19802_));
  NOR3_X1    g19610(.A1(new_n19573_), .A2(new_n19399_), .A3(new_n19802_), .ZN(new_n19803_));
  INV_X1     g19611(.I(new_n19803_), .ZN(new_n19804_));
  NOR3_X1    g19612(.A1(new_n19802_), .A2(new_n19399_), .A3(new_n19130_), .ZN(new_n19805_));
  AOI22_X1   g19613(.A1(new_n19804_), .A2(new_n19130_), .B1(\asqrt[8] ), .B2(new_n19805_), .ZN(new_n19806_));
  NOR3_X1    g19614(.A1(new_n19799_), .A2(new_n19792_), .A3(\asqrt[39] ), .ZN(new_n19807_));
  NOR2_X1    g19615(.A1(new_n19807_), .A2(new_n19806_), .ZN(new_n19808_));
  OAI21_X1   g19616(.A1(new_n19808_), .A2(new_n19801_), .B(\asqrt[40] ), .ZN(new_n19809_));
  INV_X1     g19617(.I(new_n19137_), .ZN(new_n19810_));
  NOR3_X1    g19618(.A1(new_n19408_), .A2(new_n19133_), .A3(new_n19810_), .ZN(new_n19811_));
  NOR3_X1    g19619(.A1(new_n19573_), .A2(new_n19133_), .A3(new_n19408_), .ZN(new_n19812_));
  INV_X1     g19620(.I(new_n19812_), .ZN(new_n19813_));
  AOI22_X1   g19621(.A1(new_n19813_), .A2(new_n19810_), .B1(\asqrt[8] ), .B2(new_n19811_), .ZN(new_n19814_));
  INV_X1     g19622(.I(new_n19814_), .ZN(new_n19815_));
  NAND2_X1   g19623(.A1(new_n19800_), .A2(new_n4071_), .ZN(new_n19816_));
  OAI21_X1   g19624(.A1(new_n19808_), .A2(new_n19816_), .B(new_n19815_), .ZN(new_n19817_));
  AOI21_X1   g19625(.A1(new_n19817_), .A2(new_n19809_), .B(new_n3782_), .ZN(new_n19818_));
  NOR3_X1    g19626(.A1(new_n19573_), .A2(new_n19142_), .A3(new_n19148_), .ZN(new_n19819_));
  INV_X1     g19627(.I(new_n19819_), .ZN(new_n19820_));
  NOR3_X1    g19628(.A1(new_n19142_), .A2(new_n19325_), .A3(new_n19148_), .ZN(new_n19821_));
  AOI22_X1   g19629(.A1(new_n19820_), .A2(new_n19325_), .B1(\asqrt[8] ), .B2(new_n19821_), .ZN(new_n19822_));
  OAI21_X1   g19630(.A1(new_n19806_), .A2(new_n19807_), .B(new_n19800_), .ZN(new_n19823_));
  AOI21_X1   g19631(.A1(new_n19823_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n19824_));
  AOI21_X1   g19632(.A1(new_n19824_), .A2(new_n19817_), .B(new_n19822_), .ZN(new_n19825_));
  OAI21_X1   g19633(.A1(new_n19825_), .A2(new_n19818_), .B(\asqrt[42] ), .ZN(new_n19826_));
  INV_X1     g19634(.I(new_n19826_), .ZN(new_n19827_));
  NOR2_X1    g19635(.A1(new_n19149_), .A2(new_n19157_), .ZN(new_n19828_));
  NOR3_X1    g19636(.A1(new_n19828_), .A2(new_n19407_), .A3(new_n19156_), .ZN(new_n19829_));
  NOR3_X1    g19637(.A1(new_n19573_), .A2(new_n19407_), .A3(new_n19828_), .ZN(new_n19830_));
  INV_X1     g19638(.I(new_n19830_), .ZN(new_n19831_));
  AOI22_X1   g19639(.A1(new_n19831_), .A2(new_n19156_), .B1(\asqrt[8] ), .B2(new_n19829_), .ZN(new_n19832_));
  NOR3_X1    g19640(.A1(new_n19825_), .A2(new_n19818_), .A3(\asqrt[42] ), .ZN(new_n19833_));
  NOR2_X1    g19641(.A1(new_n19833_), .A2(new_n19832_), .ZN(new_n19834_));
  OAI21_X1   g19642(.A1(new_n19834_), .A2(new_n19827_), .B(\asqrt[43] ), .ZN(new_n19835_));
  INV_X1     g19643(.I(new_n19163_), .ZN(new_n19836_));
  NOR3_X1    g19644(.A1(new_n19573_), .A2(new_n19159_), .A3(new_n19416_), .ZN(new_n19837_));
  INV_X1     g19645(.I(new_n19837_), .ZN(new_n19838_));
  NOR3_X1    g19646(.A1(new_n19416_), .A2(new_n19159_), .A3(new_n19836_), .ZN(new_n19839_));
  AOI22_X1   g19647(.A1(new_n19838_), .A2(new_n19836_), .B1(\asqrt[8] ), .B2(new_n19839_), .ZN(new_n19840_));
  INV_X1     g19648(.I(new_n19840_), .ZN(new_n19841_));
  NAND2_X1   g19649(.A1(new_n19826_), .A2(new_n3218_), .ZN(new_n19842_));
  OAI21_X1   g19650(.A1(new_n19834_), .A2(new_n19842_), .B(new_n19841_), .ZN(new_n19843_));
  AOI21_X1   g19651(.A1(new_n19843_), .A2(new_n19835_), .B(new_n2954_), .ZN(new_n19844_));
  NOR3_X1    g19652(.A1(new_n19168_), .A2(new_n19324_), .A3(new_n19176_), .ZN(new_n19845_));
  NOR3_X1    g19653(.A1(new_n19573_), .A2(new_n19168_), .A3(new_n19176_), .ZN(new_n19846_));
  INV_X1     g19654(.I(new_n19846_), .ZN(new_n19847_));
  AOI22_X1   g19655(.A1(new_n19847_), .A2(new_n19324_), .B1(\asqrt[8] ), .B2(new_n19845_), .ZN(new_n19848_));
  OAI21_X1   g19656(.A1(new_n19832_), .A2(new_n19833_), .B(new_n19826_), .ZN(new_n19849_));
  AOI21_X1   g19657(.A1(new_n19849_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n19850_));
  AOI21_X1   g19658(.A1(new_n19850_), .A2(new_n19843_), .B(new_n19848_), .ZN(new_n19851_));
  OAI21_X1   g19659(.A1(new_n19851_), .A2(new_n19844_), .B(\asqrt[45] ), .ZN(new_n19852_));
  INV_X1     g19660(.I(new_n19852_), .ZN(new_n19853_));
  NOR2_X1    g19661(.A1(new_n19177_), .A2(new_n19184_), .ZN(new_n19854_));
  NOR3_X1    g19662(.A1(new_n19573_), .A2(new_n19415_), .A3(new_n19854_), .ZN(new_n19855_));
  INV_X1     g19663(.I(new_n19855_), .ZN(new_n19856_));
  NOR3_X1    g19664(.A1(new_n19854_), .A2(new_n19415_), .A3(new_n19183_), .ZN(new_n19857_));
  AOI22_X1   g19665(.A1(new_n19856_), .A2(new_n19183_), .B1(\asqrt[8] ), .B2(new_n19857_), .ZN(new_n19858_));
  NOR3_X1    g19666(.A1(new_n19851_), .A2(new_n19844_), .A3(\asqrt[45] ), .ZN(new_n19859_));
  NOR2_X1    g19667(.A1(new_n19859_), .A2(new_n19858_), .ZN(new_n19860_));
  OAI21_X1   g19668(.A1(new_n19860_), .A2(new_n19853_), .B(\asqrt[46] ), .ZN(new_n19861_));
  INV_X1     g19669(.I(new_n19192_), .ZN(new_n19862_));
  NOR3_X1    g19670(.A1(new_n19424_), .A2(new_n19186_), .A3(new_n19862_), .ZN(new_n19863_));
  NOR3_X1    g19671(.A1(new_n19573_), .A2(new_n19186_), .A3(new_n19424_), .ZN(new_n19864_));
  INV_X1     g19672(.I(new_n19864_), .ZN(new_n19865_));
  AOI22_X1   g19673(.A1(new_n19865_), .A2(new_n19862_), .B1(\asqrt[8] ), .B2(new_n19863_), .ZN(new_n19866_));
  INV_X1     g19674(.I(new_n19866_), .ZN(new_n19867_));
  NAND2_X1   g19675(.A1(new_n19852_), .A2(new_n2465_), .ZN(new_n19868_));
  OAI21_X1   g19676(.A1(new_n19860_), .A2(new_n19868_), .B(new_n19867_), .ZN(new_n19869_));
  AOI21_X1   g19677(.A1(new_n19869_), .A2(new_n19861_), .B(new_n2229_), .ZN(new_n19870_));
  NOR3_X1    g19678(.A1(new_n19573_), .A2(new_n19197_), .A3(new_n19206_), .ZN(new_n19871_));
  INV_X1     g19679(.I(new_n19871_), .ZN(new_n19872_));
  NOR3_X1    g19680(.A1(new_n19197_), .A2(new_n19323_), .A3(new_n19206_), .ZN(new_n19873_));
  AOI22_X1   g19681(.A1(new_n19872_), .A2(new_n19323_), .B1(\asqrt[8] ), .B2(new_n19873_), .ZN(new_n19874_));
  OAI21_X1   g19682(.A1(new_n19858_), .A2(new_n19859_), .B(new_n19852_), .ZN(new_n19875_));
  AOI21_X1   g19683(.A1(new_n19875_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n19876_));
  AOI21_X1   g19684(.A1(new_n19876_), .A2(new_n19869_), .B(new_n19874_), .ZN(new_n19877_));
  OAI21_X1   g19685(.A1(new_n19877_), .A2(new_n19870_), .B(\asqrt[48] ), .ZN(new_n19878_));
  INV_X1     g19686(.I(new_n19878_), .ZN(new_n19879_));
  NOR2_X1    g19687(.A1(new_n19207_), .A2(new_n19214_), .ZN(new_n19880_));
  NOR3_X1    g19688(.A1(new_n19880_), .A2(new_n19423_), .A3(new_n19213_), .ZN(new_n19881_));
  NOR3_X1    g19689(.A1(new_n19573_), .A2(new_n19423_), .A3(new_n19880_), .ZN(new_n19882_));
  INV_X1     g19690(.I(new_n19882_), .ZN(new_n19883_));
  AOI22_X1   g19691(.A1(new_n19883_), .A2(new_n19213_), .B1(\asqrt[8] ), .B2(new_n19881_), .ZN(new_n19884_));
  NOR3_X1    g19692(.A1(new_n19877_), .A2(new_n19870_), .A3(\asqrt[48] ), .ZN(new_n19885_));
  NOR2_X1    g19693(.A1(new_n19885_), .A2(new_n19884_), .ZN(new_n19886_));
  OAI21_X1   g19694(.A1(new_n19886_), .A2(new_n19879_), .B(\asqrt[49] ), .ZN(new_n19887_));
  INV_X1     g19695(.I(new_n19222_), .ZN(new_n19888_));
  NOR3_X1    g19696(.A1(new_n19573_), .A2(new_n19216_), .A3(new_n19432_), .ZN(new_n19889_));
  INV_X1     g19697(.I(new_n19889_), .ZN(new_n19890_));
  NOR3_X1    g19698(.A1(new_n19432_), .A2(new_n19216_), .A3(new_n19888_), .ZN(new_n19891_));
  AOI22_X1   g19699(.A1(new_n19890_), .A2(new_n19888_), .B1(\asqrt[8] ), .B2(new_n19891_), .ZN(new_n19892_));
  INV_X1     g19700(.I(new_n19892_), .ZN(new_n19893_));
  NAND2_X1   g19701(.A1(new_n19878_), .A2(new_n1806_), .ZN(new_n19894_));
  OAI21_X1   g19702(.A1(new_n19886_), .A2(new_n19894_), .B(new_n19893_), .ZN(new_n19895_));
  AOI21_X1   g19703(.A1(new_n19895_), .A2(new_n19887_), .B(new_n1612_), .ZN(new_n19896_));
  NOR3_X1    g19704(.A1(new_n19227_), .A2(new_n19322_), .A3(new_n19236_), .ZN(new_n19897_));
  NOR3_X1    g19705(.A1(new_n19573_), .A2(new_n19227_), .A3(new_n19236_), .ZN(new_n19898_));
  INV_X1     g19706(.I(new_n19898_), .ZN(new_n19899_));
  AOI22_X1   g19707(.A1(new_n19899_), .A2(new_n19322_), .B1(\asqrt[8] ), .B2(new_n19897_), .ZN(new_n19900_));
  OAI21_X1   g19708(.A1(new_n19884_), .A2(new_n19885_), .B(new_n19878_), .ZN(new_n19901_));
  AOI21_X1   g19709(.A1(new_n19901_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n19902_));
  AOI21_X1   g19710(.A1(new_n19902_), .A2(new_n19895_), .B(new_n19900_), .ZN(new_n19903_));
  OAI21_X1   g19711(.A1(new_n19903_), .A2(new_n19896_), .B(\asqrt[51] ), .ZN(new_n19904_));
  INV_X1     g19712(.I(new_n19904_), .ZN(new_n19905_));
  NOR2_X1    g19713(.A1(new_n19237_), .A2(new_n19244_), .ZN(new_n19906_));
  NOR3_X1    g19714(.A1(new_n19573_), .A2(new_n19431_), .A3(new_n19906_), .ZN(new_n19907_));
  INV_X1     g19715(.I(new_n19907_), .ZN(new_n19908_));
  NOR3_X1    g19716(.A1(new_n19906_), .A2(new_n19431_), .A3(new_n19243_), .ZN(new_n19909_));
  AOI22_X1   g19717(.A1(new_n19908_), .A2(new_n19243_), .B1(\asqrt[8] ), .B2(new_n19909_), .ZN(new_n19910_));
  NOR3_X1    g19718(.A1(new_n19903_), .A2(new_n19896_), .A3(\asqrt[51] ), .ZN(new_n19911_));
  NOR2_X1    g19719(.A1(new_n19911_), .A2(new_n19910_), .ZN(new_n19912_));
  OAI21_X1   g19720(.A1(new_n19912_), .A2(new_n19905_), .B(\asqrt[52] ), .ZN(new_n19913_));
  INV_X1     g19721(.I(new_n19252_), .ZN(new_n19914_));
  NAND2_X1   g19722(.A1(new_n19254_), .A2(new_n19245_), .ZN(new_n19915_));
  INV_X1     g19723(.I(new_n19915_), .ZN(new_n19916_));
  NOR3_X1    g19724(.A1(new_n19916_), .A2(new_n19246_), .A3(new_n19914_), .ZN(new_n19917_));
  NOR3_X1    g19725(.A1(new_n19573_), .A2(new_n19246_), .A3(new_n19916_), .ZN(new_n19918_));
  INV_X1     g19726(.I(new_n19918_), .ZN(new_n19919_));
  AOI22_X1   g19727(.A1(new_n19919_), .A2(new_n19914_), .B1(\asqrt[8] ), .B2(new_n19917_), .ZN(new_n19920_));
  INV_X1     g19728(.I(new_n19920_), .ZN(new_n19921_));
  NAND2_X1   g19729(.A1(new_n19904_), .A2(new_n1256_), .ZN(new_n19922_));
  OAI21_X1   g19730(.A1(new_n19912_), .A2(new_n19922_), .B(new_n19921_), .ZN(new_n19923_));
  AOI21_X1   g19731(.A1(new_n19923_), .A2(new_n19913_), .B(new_n1103_), .ZN(new_n19924_));
  NOR3_X1    g19732(.A1(new_n19573_), .A2(new_n19257_), .A3(new_n19266_), .ZN(new_n19925_));
  INV_X1     g19733(.I(new_n19925_), .ZN(new_n19926_));
  NOR3_X1    g19734(.A1(new_n19257_), .A2(new_n19321_), .A3(new_n19266_), .ZN(new_n19927_));
  AOI22_X1   g19735(.A1(new_n19926_), .A2(new_n19321_), .B1(\asqrt[8] ), .B2(new_n19927_), .ZN(new_n19928_));
  OAI21_X1   g19736(.A1(new_n19910_), .A2(new_n19911_), .B(new_n19904_), .ZN(new_n19929_));
  AOI21_X1   g19737(.A1(new_n19929_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n19930_));
  AOI21_X1   g19738(.A1(new_n19930_), .A2(new_n19923_), .B(new_n19928_), .ZN(new_n19931_));
  OAI21_X1   g19739(.A1(new_n19931_), .A2(new_n19924_), .B(\asqrt[54] ), .ZN(new_n19932_));
  INV_X1     g19740(.I(new_n19932_), .ZN(new_n19933_));
  INV_X1     g19741(.I(new_n19268_), .ZN(new_n19934_));
  INV_X1     g19742(.I(new_n19439_), .ZN(new_n19935_));
  NOR3_X1    g19743(.A1(new_n19934_), .A2(new_n19935_), .A3(new_n19273_), .ZN(new_n19936_));
  NOR3_X1    g19744(.A1(new_n19573_), .A2(new_n19934_), .A3(new_n19935_), .ZN(new_n19937_));
  INV_X1     g19745(.I(new_n19937_), .ZN(new_n19938_));
  AOI22_X1   g19746(.A1(new_n19938_), .A2(new_n19273_), .B1(\asqrt[8] ), .B2(new_n19936_), .ZN(new_n19939_));
  NOR3_X1    g19747(.A1(new_n19931_), .A2(new_n19924_), .A3(\asqrt[54] ), .ZN(new_n19940_));
  NOR2_X1    g19748(.A1(new_n19940_), .A2(new_n19939_), .ZN(new_n19941_));
  OAI21_X1   g19749(.A1(new_n19941_), .A2(new_n19933_), .B(\asqrt[55] ), .ZN(new_n19942_));
  INV_X1     g19750(.I(new_n19282_), .ZN(new_n19943_));
  INV_X1     g19751(.I(new_n19275_), .ZN(new_n19944_));
  INV_X1     g19752(.I(new_n19284_), .ZN(new_n19945_));
  NOR2_X1    g19753(.A1(new_n19945_), .A2(new_n19944_), .ZN(new_n19946_));
  NOR3_X1    g19754(.A1(new_n19573_), .A2(new_n19276_), .A3(new_n19946_), .ZN(new_n19947_));
  INV_X1     g19755(.I(new_n19947_), .ZN(new_n19948_));
  NOR3_X1    g19756(.A1(new_n19946_), .A2(new_n19276_), .A3(new_n19943_), .ZN(new_n19949_));
  AOI22_X1   g19757(.A1(new_n19948_), .A2(new_n19943_), .B1(\asqrt[8] ), .B2(new_n19949_), .ZN(new_n19950_));
  INV_X1     g19758(.I(new_n19950_), .ZN(new_n19951_));
  NAND2_X1   g19759(.A1(new_n19932_), .A2(new_n823_), .ZN(new_n19952_));
  OAI21_X1   g19760(.A1(new_n19941_), .A2(new_n19952_), .B(new_n19951_), .ZN(new_n19953_));
  AOI21_X1   g19761(.A1(new_n19953_), .A2(new_n19942_), .B(new_n703_), .ZN(new_n19954_));
  NOR3_X1    g19762(.A1(new_n19287_), .A2(new_n19320_), .A3(new_n19293_), .ZN(new_n19955_));
  NOR3_X1    g19763(.A1(new_n19573_), .A2(new_n19287_), .A3(new_n19293_), .ZN(new_n19956_));
  INV_X1     g19764(.I(new_n19956_), .ZN(new_n19957_));
  AOI22_X1   g19765(.A1(new_n19957_), .A2(new_n19320_), .B1(\asqrt[8] ), .B2(new_n19955_), .ZN(new_n19958_));
  OAI21_X1   g19766(.A1(new_n19939_), .A2(new_n19940_), .B(new_n19932_), .ZN(new_n19959_));
  AOI21_X1   g19767(.A1(new_n19959_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n19960_));
  AOI21_X1   g19768(.A1(new_n19960_), .A2(new_n19953_), .B(new_n19958_), .ZN(new_n19961_));
  OAI21_X1   g19769(.A1(new_n19961_), .A2(new_n19954_), .B(\asqrt[57] ), .ZN(new_n19962_));
  INV_X1     g19770(.I(new_n19962_), .ZN(new_n19963_));
  INV_X1     g19771(.I(new_n19295_), .ZN(new_n19964_));
  INV_X1     g19772(.I(new_n19443_), .ZN(new_n19965_));
  NOR3_X1    g19773(.A1(new_n19573_), .A2(new_n19964_), .A3(new_n19965_), .ZN(new_n19966_));
  INV_X1     g19774(.I(new_n19966_), .ZN(new_n19967_));
  NOR3_X1    g19775(.A1(new_n19964_), .A2(new_n19965_), .A3(new_n19300_), .ZN(new_n19968_));
  AOI22_X1   g19776(.A1(new_n19967_), .A2(new_n19300_), .B1(\asqrt[8] ), .B2(new_n19968_), .ZN(new_n19969_));
  NOR3_X1    g19777(.A1(new_n19961_), .A2(new_n19954_), .A3(\asqrt[57] ), .ZN(new_n19970_));
  NOR2_X1    g19778(.A1(new_n19970_), .A2(new_n19969_), .ZN(new_n19971_));
  OAI21_X1   g19779(.A1(new_n19971_), .A2(new_n19963_), .B(\asqrt[58] ), .ZN(new_n19972_));
  INV_X1     g19780(.I(new_n19309_), .ZN(new_n19973_));
  INV_X1     g19781(.I(new_n19302_), .ZN(new_n19974_));
  INV_X1     g19782(.I(new_n19311_), .ZN(new_n19975_));
  OAI21_X1   g19783(.A1(new_n19975_), .A2(new_n19974_), .B(new_n19309_), .ZN(new_n19976_));
  NOR2_X1    g19784(.A1(new_n19976_), .A2(new_n19303_), .ZN(new_n19977_));
  NOR2_X1    g19785(.A1(new_n19975_), .A2(new_n19974_), .ZN(new_n19978_));
  NOR3_X1    g19786(.A1(new_n19573_), .A2(new_n19303_), .A3(new_n19978_), .ZN(new_n19979_));
  INV_X1     g19787(.I(new_n19979_), .ZN(new_n19980_));
  AOI22_X1   g19788(.A1(new_n19980_), .A2(new_n19973_), .B1(\asqrt[8] ), .B2(new_n19977_), .ZN(new_n19981_));
  INV_X1     g19789(.I(new_n19981_), .ZN(new_n19982_));
  NAND2_X1   g19790(.A1(new_n19962_), .A2(new_n436_), .ZN(new_n19983_));
  OAI21_X1   g19791(.A1(new_n19971_), .A2(new_n19983_), .B(new_n19982_), .ZN(new_n19984_));
  AOI21_X1   g19792(.A1(new_n19984_), .A2(new_n19972_), .B(new_n327_), .ZN(new_n19985_));
  NOR3_X1    g19793(.A1(new_n19573_), .A2(new_n19463_), .A3(new_n19464_), .ZN(new_n19986_));
  INV_X1     g19794(.I(new_n19986_), .ZN(new_n19987_));
  NOR3_X1    g19795(.A1(new_n19463_), .A2(new_n19319_), .A3(new_n19464_), .ZN(new_n19988_));
  AOI22_X1   g19796(.A1(new_n19987_), .A2(new_n19319_), .B1(\asqrt[8] ), .B2(new_n19988_), .ZN(new_n19989_));
  OAI21_X1   g19797(.A1(new_n19969_), .A2(new_n19970_), .B(new_n19962_), .ZN(new_n19990_));
  AOI21_X1   g19798(.A1(new_n19990_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n19991_));
  AOI21_X1   g19799(.A1(new_n19991_), .A2(new_n19984_), .B(new_n19989_), .ZN(new_n19992_));
  OAI21_X1   g19800(.A1(new_n19992_), .A2(new_n19985_), .B(\asqrt[60] ), .ZN(new_n19993_));
  INV_X1     g19801(.I(new_n19993_), .ZN(new_n19994_));
  INV_X1     g19802(.I(new_n19522_), .ZN(new_n19995_));
  NOR3_X1    g19803(.A1(new_n19995_), .A2(new_n19447_), .A3(new_n19475_), .ZN(new_n19996_));
  NOR3_X1    g19804(.A1(new_n19573_), .A2(new_n19447_), .A3(new_n19995_), .ZN(new_n19997_));
  INV_X1     g19805(.I(new_n19997_), .ZN(new_n19998_));
  AOI22_X1   g19806(.A1(new_n19998_), .A2(new_n19475_), .B1(\asqrt[8] ), .B2(new_n19996_), .ZN(new_n19999_));
  NOR3_X1    g19807(.A1(new_n19992_), .A2(new_n19985_), .A3(\asqrt[60] ), .ZN(new_n20000_));
  NOR2_X1    g19808(.A1(new_n20000_), .A2(new_n19999_), .ZN(new_n20001_));
  OAI21_X1   g19809(.A1(new_n20001_), .A2(new_n19994_), .B(\asqrt[61] ), .ZN(new_n20002_));
  NAND2_X1   g19810(.A1(new_n19487_), .A2(new_n19476_), .ZN(new_n20003_));
  NAND3_X1   g19811(.A1(\asqrt[8] ), .A2(new_n19455_), .A3(new_n20003_), .ZN(new_n20004_));
  AND3_X2    g19812(.A1(new_n19455_), .A2(new_n19461_), .A3(new_n20003_), .Z(new_n20005_));
  AOI22_X1   g19813(.A1(new_n20004_), .A2(new_n19462_), .B1(\asqrt[8] ), .B2(new_n20005_), .ZN(new_n20006_));
  INV_X1     g19814(.I(new_n20006_), .ZN(new_n20007_));
  NAND2_X1   g19815(.A1(new_n19993_), .A2(new_n218_), .ZN(new_n20008_));
  OAI21_X1   g19816(.A1(new_n20001_), .A2(new_n20008_), .B(new_n20007_), .ZN(new_n20009_));
  AOI21_X1   g19817(.A1(new_n20009_), .A2(new_n20002_), .B(new_n207_), .ZN(new_n20010_));
  NOR3_X1    g19818(.A1(new_n19469_), .A2(new_n19521_), .A3(new_n19500_), .ZN(new_n20011_));
  NOR3_X1    g19819(.A1(new_n19573_), .A2(new_n19469_), .A3(new_n19500_), .ZN(new_n20012_));
  INV_X1     g19820(.I(new_n20012_), .ZN(new_n20013_));
  AOI22_X1   g19821(.A1(new_n20013_), .A2(new_n19521_), .B1(\asqrt[8] ), .B2(new_n20011_), .ZN(new_n20014_));
  OAI21_X1   g19822(.A1(new_n19999_), .A2(new_n20000_), .B(new_n19993_), .ZN(new_n20015_));
  AOI21_X1   g19823(.A1(new_n20015_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n20016_));
  AOI21_X1   g19824(.A1(new_n20016_), .A2(new_n20009_), .B(new_n20014_), .ZN(new_n20017_));
  INV_X1     g19825(.I(new_n19480_), .ZN(new_n20018_));
  INV_X1     g19826(.I(new_n19534_), .ZN(new_n20019_));
  NOR3_X1    g19827(.A1(new_n20018_), .A2(new_n20019_), .A3(new_n19485_), .ZN(new_n20020_));
  NAND2_X1   g19828(.A1(\asqrt[8] ), .A2(new_n20020_), .ZN(new_n20021_));
  INV_X1     g19829(.I(new_n20021_), .ZN(new_n20022_));
  NOR2_X1    g19830(.A1(new_n20018_), .A2(new_n20019_), .ZN(new_n20023_));
  AOI21_X1   g19831(.A1(\asqrt[8] ), .A2(new_n20023_), .B(new_n19484_), .ZN(new_n20024_));
  NOR2_X1    g19832(.A1(new_n20022_), .A2(new_n20024_), .ZN(new_n20025_));
  INV_X1     g19833(.I(new_n20025_), .ZN(new_n20026_));
  NAND3_X1   g19834(.A1(\asqrt[8] ), .A2(new_n19518_), .A3(new_n19495_), .ZN(new_n20027_));
  AND3_X2    g19835(.A1(new_n20026_), .A2(new_n19548_), .A3(new_n20027_), .Z(new_n20028_));
  OAI21_X1   g19836(.A1(new_n20017_), .A2(new_n20010_), .B(new_n20028_), .ZN(new_n20029_));
  NAND2_X1   g19837(.A1(new_n20029_), .A2(new_n193_), .ZN(new_n20030_));
  INV_X1     g19838(.I(new_n19999_), .ZN(new_n20031_));
  INV_X1     g19839(.I(new_n19969_), .ZN(new_n20032_));
  INV_X1     g19840(.I(new_n19939_), .ZN(new_n20033_));
  INV_X1     g19841(.I(new_n19910_), .ZN(new_n20034_));
  INV_X1     g19842(.I(new_n19884_), .ZN(new_n20035_));
  INV_X1     g19843(.I(new_n19858_), .ZN(new_n20036_));
  INV_X1     g19844(.I(new_n19832_), .ZN(new_n20037_));
  INV_X1     g19845(.I(new_n19806_), .ZN(new_n20038_));
  INV_X1     g19846(.I(new_n19780_), .ZN(new_n20039_));
  INV_X1     g19847(.I(new_n19754_), .ZN(new_n20040_));
  INV_X1     g19848(.I(new_n19728_), .ZN(new_n20041_));
  INV_X1     g19849(.I(new_n19702_), .ZN(new_n20042_));
  INV_X1     g19850(.I(new_n19676_), .ZN(new_n20043_));
  INV_X1     g19851(.I(new_n19650_), .ZN(new_n20044_));
  INV_X1     g19852(.I(new_n19624_), .ZN(new_n20045_));
  INV_X1     g19853(.I(new_n19600_), .ZN(new_n20046_));
  NAND2_X1   g19854(.A1(new_n19531_), .A2(new_n19539_), .ZN(new_n20047_));
  OAI21_X1   g19855(.A1(new_n19520_), .A2(new_n19530_), .B(new_n19533_), .ZN(new_n20048_));
  NAND2_X1   g19856(.A1(new_n20048_), .A2(\a[17] ), .ZN(new_n20049_));
  NAND3_X1   g19857(.A1(new_n20047_), .A2(new_n20049_), .A3(new_n19547_), .ZN(new_n20050_));
  AOI21_X1   g19858(.A1(new_n20050_), .A2(new_n19562_), .B(new_n18275_), .ZN(new_n20051_));
  OAI21_X1   g19859(.A1(new_n19553_), .A2(new_n19542_), .B(\a[18] ), .ZN(new_n20052_));
  NAND3_X1   g19860(.A1(new_n19550_), .A2(new_n19547_), .A3(new_n18793_), .ZN(new_n20053_));
  NAND2_X1   g19861(.A1(new_n19531_), .A2(new_n19517_), .ZN(new_n20054_));
  AOI21_X1   g19862(.A1(new_n20054_), .A2(\asqrt[9] ), .B(\asqrt[10] ), .ZN(new_n20055_));
  AOI22_X1   g19863(.A1(new_n20050_), .A2(new_n20055_), .B1(new_n20052_), .B2(new_n20053_), .ZN(new_n20056_));
  OAI21_X1   g19864(.A1(new_n20056_), .A2(new_n20051_), .B(\asqrt[11] ), .ZN(new_n20057_));
  NAND2_X1   g19865(.A1(new_n20057_), .A2(new_n16881_), .ZN(new_n20058_));
  OAI21_X1   g19866(.A1(new_n20058_), .A2(new_n19567_), .B(new_n19575_), .ZN(new_n20059_));
  AOI21_X1   g19867(.A1(new_n20059_), .A2(new_n19568_), .B(new_n16389_), .ZN(new_n20060_));
  INV_X1     g19868(.I(new_n19561_), .ZN(new_n20061_));
  AOI21_X1   g19869(.A1(\a[17] ), .A2(new_n20048_), .B(new_n19542_), .ZN(new_n20062_));
  AOI21_X1   g19870(.A1(new_n20062_), .A2(new_n20047_), .B(new_n19532_), .ZN(new_n20063_));
  OAI21_X1   g19871(.A1(new_n20063_), .A2(new_n18275_), .B(new_n17623_), .ZN(new_n20064_));
  OAI21_X1   g19872(.A1(new_n20064_), .A2(new_n20056_), .B(new_n20061_), .ZN(new_n20065_));
  NAND2_X1   g19873(.A1(new_n20065_), .A2(new_n20057_), .ZN(new_n20066_));
  AOI21_X1   g19874(.A1(new_n20066_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n20067_));
  AOI21_X1   g19875(.A1(new_n20067_), .A2(new_n20059_), .B(new_n19583_), .ZN(new_n20068_));
  OAI21_X1   g19876(.A1(new_n20068_), .A2(new_n20060_), .B(\asqrt[14] ), .ZN(new_n20069_));
  NAND2_X1   g19877(.A1(new_n20069_), .A2(new_n15067_), .ZN(new_n20070_));
  OAI21_X1   g19878(.A1(new_n20070_), .A2(new_n19594_), .B(new_n20046_), .ZN(new_n20071_));
  NAND3_X1   g19879(.A1(new_n20071_), .A2(new_n14601_), .A3(new_n19595_), .ZN(new_n20072_));
  AOI22_X1   g19880(.A1(new_n20072_), .A2(new_n19609_), .B1(new_n19617_), .B2(\asqrt[16] ), .ZN(new_n20073_));
  OAI21_X1   g19881(.A1(new_n20073_), .A2(new_n14017_), .B(new_n13353_), .ZN(new_n20074_));
  OAI21_X1   g19882(.A1(new_n20074_), .A2(new_n19619_), .B(new_n20045_), .ZN(new_n20075_));
  AOI21_X1   g19883(.A1(new_n20075_), .A2(new_n19620_), .B(new_n12913_), .ZN(new_n20076_));
  AOI21_X1   g19884(.A1(new_n20071_), .A2(new_n19595_), .B(new_n14601_), .ZN(new_n20077_));
  NOR3_X1    g19885(.A1(new_n20068_), .A2(new_n20060_), .A3(\asqrt[14] ), .ZN(new_n20078_));
  OAI21_X1   g19886(.A1(new_n19591_), .A2(new_n20078_), .B(new_n20069_), .ZN(new_n20079_));
  AOI21_X1   g19887(.A1(new_n20079_), .A2(\asqrt[15] ), .B(\asqrt[16] ), .ZN(new_n20080_));
  AOI21_X1   g19888(.A1(new_n20080_), .A2(new_n20071_), .B(new_n19608_), .ZN(new_n20081_));
  NOR3_X1    g19889(.A1(new_n20081_), .A2(\asqrt[17] ), .A3(new_n20077_), .ZN(new_n20082_));
  OAI22_X1   g19890(.A1(new_n20082_), .A2(new_n19616_), .B1(new_n20073_), .B2(new_n14017_), .ZN(new_n20083_));
  AOI21_X1   g19891(.A1(new_n20083_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n20084_));
  AOI21_X1   g19892(.A1(new_n20084_), .A2(new_n20075_), .B(new_n19632_), .ZN(new_n20085_));
  OAI21_X1   g19893(.A1(new_n20085_), .A2(new_n20076_), .B(\asqrt[20] ), .ZN(new_n20086_));
  NAND2_X1   g19894(.A1(new_n20086_), .A2(new_n11736_), .ZN(new_n20087_));
  OAI21_X1   g19895(.A1(new_n20087_), .A2(new_n19643_), .B(new_n20044_), .ZN(new_n20088_));
  AOI21_X1   g19896(.A1(new_n20088_), .A2(new_n19644_), .B(new_n11326_), .ZN(new_n20089_));
  NOR3_X1    g19897(.A1(new_n20085_), .A2(\asqrt[20] ), .A3(new_n20076_), .ZN(new_n20090_));
  OAI21_X1   g19898(.A1(new_n19640_), .A2(new_n20090_), .B(new_n20086_), .ZN(new_n20091_));
  AOI21_X1   g19899(.A1(new_n20091_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n20092_));
  AOI21_X1   g19900(.A1(new_n20092_), .A2(new_n20088_), .B(new_n19658_), .ZN(new_n20093_));
  OAI21_X1   g19901(.A1(new_n20093_), .A2(new_n20089_), .B(\asqrt[23] ), .ZN(new_n20094_));
  NAND2_X1   g19902(.A1(new_n20094_), .A2(new_n10221_), .ZN(new_n20095_));
  OAI21_X1   g19903(.A1(new_n20095_), .A2(new_n19669_), .B(new_n20043_), .ZN(new_n20096_));
  AOI21_X1   g19904(.A1(new_n20096_), .A2(new_n19670_), .B(new_n9846_), .ZN(new_n20097_));
  NOR3_X1    g19905(.A1(new_n20093_), .A2(\asqrt[23] ), .A3(new_n20089_), .ZN(new_n20098_));
  OAI21_X1   g19906(.A1(new_n19666_), .A2(new_n20098_), .B(new_n20094_), .ZN(new_n20099_));
  AOI21_X1   g19907(.A1(new_n20099_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n20100_));
  AOI21_X1   g19908(.A1(new_n20100_), .A2(new_n20096_), .B(new_n19684_), .ZN(new_n20101_));
  OAI21_X1   g19909(.A1(new_n20101_), .A2(new_n20097_), .B(\asqrt[26] ), .ZN(new_n20102_));
  NAND2_X1   g19910(.A1(new_n20102_), .A2(new_n8826_), .ZN(new_n20103_));
  OAI21_X1   g19911(.A1(new_n20103_), .A2(new_n19695_), .B(new_n20042_), .ZN(new_n20104_));
  AOI21_X1   g19912(.A1(new_n20104_), .A2(new_n19696_), .B(new_n8483_), .ZN(new_n20105_));
  NOR3_X1    g19913(.A1(new_n20101_), .A2(\asqrt[26] ), .A3(new_n20097_), .ZN(new_n20106_));
  OAI21_X1   g19914(.A1(new_n19692_), .A2(new_n20106_), .B(new_n20102_), .ZN(new_n20107_));
  AOI21_X1   g19915(.A1(new_n20107_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n20108_));
  AOI21_X1   g19916(.A1(new_n20108_), .A2(new_n20104_), .B(new_n19710_), .ZN(new_n20109_));
  OAI21_X1   g19917(.A1(new_n20109_), .A2(new_n20105_), .B(\asqrt[29] ), .ZN(new_n20110_));
  NAND2_X1   g19918(.A1(new_n20110_), .A2(new_n7539_), .ZN(new_n20111_));
  OAI21_X1   g19919(.A1(new_n20111_), .A2(new_n19721_), .B(new_n20041_), .ZN(new_n20112_));
  AOI21_X1   g19920(.A1(new_n20112_), .A2(new_n19722_), .B(new_n7229_), .ZN(new_n20113_));
  NOR3_X1    g19921(.A1(new_n20109_), .A2(\asqrt[29] ), .A3(new_n20105_), .ZN(new_n20114_));
  OAI21_X1   g19922(.A1(new_n19718_), .A2(new_n20114_), .B(new_n20110_), .ZN(new_n20115_));
  AOI21_X1   g19923(.A1(new_n20115_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n20116_));
  AOI21_X1   g19924(.A1(new_n20116_), .A2(new_n20112_), .B(new_n19736_), .ZN(new_n20117_));
  OAI21_X1   g19925(.A1(new_n20117_), .A2(new_n20113_), .B(\asqrt[32] ), .ZN(new_n20118_));
  NAND2_X1   g19926(.A1(new_n20118_), .A2(new_n6356_), .ZN(new_n20119_));
  OAI21_X1   g19927(.A1(new_n20119_), .A2(new_n19747_), .B(new_n20040_), .ZN(new_n20120_));
  AOI21_X1   g19928(.A1(new_n20120_), .A2(new_n19748_), .B(new_n6077_), .ZN(new_n20121_));
  NOR3_X1    g19929(.A1(new_n20117_), .A2(\asqrt[32] ), .A3(new_n20113_), .ZN(new_n20122_));
  OAI21_X1   g19930(.A1(new_n19744_), .A2(new_n20122_), .B(new_n20118_), .ZN(new_n20123_));
  AOI21_X1   g19931(.A1(new_n20123_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n20124_));
  AOI21_X1   g19932(.A1(new_n20124_), .A2(new_n20120_), .B(new_n19762_), .ZN(new_n20125_));
  OAI21_X1   g19933(.A1(new_n20125_), .A2(new_n20121_), .B(\asqrt[35] ), .ZN(new_n20126_));
  NAND2_X1   g19934(.A1(new_n20126_), .A2(new_n5277_), .ZN(new_n20127_));
  OAI21_X1   g19935(.A1(new_n20127_), .A2(new_n19773_), .B(new_n20039_), .ZN(new_n20128_));
  AOI21_X1   g19936(.A1(new_n20128_), .A2(new_n19774_), .B(new_n5024_), .ZN(new_n20129_));
  NOR3_X1    g19937(.A1(new_n20125_), .A2(\asqrt[35] ), .A3(new_n20121_), .ZN(new_n20130_));
  OAI21_X1   g19938(.A1(new_n19770_), .A2(new_n20130_), .B(new_n20126_), .ZN(new_n20131_));
  AOI21_X1   g19939(.A1(new_n20131_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n20132_));
  AOI21_X1   g19940(.A1(new_n20132_), .A2(new_n20128_), .B(new_n19788_), .ZN(new_n20133_));
  OAI21_X1   g19941(.A1(new_n20133_), .A2(new_n20129_), .B(\asqrt[38] ), .ZN(new_n20134_));
  NAND2_X1   g19942(.A1(new_n20134_), .A2(new_n4298_), .ZN(new_n20135_));
  OAI21_X1   g19943(.A1(new_n20135_), .A2(new_n19799_), .B(new_n20038_), .ZN(new_n20136_));
  AOI21_X1   g19944(.A1(new_n20136_), .A2(new_n19800_), .B(new_n4071_), .ZN(new_n20137_));
  NOR3_X1    g19945(.A1(new_n20133_), .A2(\asqrt[38] ), .A3(new_n20129_), .ZN(new_n20138_));
  OAI21_X1   g19946(.A1(new_n19796_), .A2(new_n20138_), .B(new_n20134_), .ZN(new_n20139_));
  AOI21_X1   g19947(.A1(new_n20139_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n20140_));
  AOI21_X1   g19948(.A1(new_n20140_), .A2(new_n20136_), .B(new_n19814_), .ZN(new_n20141_));
  OAI21_X1   g19949(.A1(new_n20141_), .A2(new_n20137_), .B(\asqrt[41] ), .ZN(new_n20142_));
  NAND2_X1   g19950(.A1(new_n20142_), .A2(new_n3419_), .ZN(new_n20143_));
  OAI21_X1   g19951(.A1(new_n20143_), .A2(new_n19825_), .B(new_n20037_), .ZN(new_n20144_));
  AOI21_X1   g19952(.A1(new_n20144_), .A2(new_n19826_), .B(new_n3218_), .ZN(new_n20145_));
  NOR3_X1    g19953(.A1(new_n20141_), .A2(\asqrt[41] ), .A3(new_n20137_), .ZN(new_n20146_));
  OAI21_X1   g19954(.A1(new_n19822_), .A2(new_n20146_), .B(new_n20142_), .ZN(new_n20147_));
  AOI21_X1   g19955(.A1(new_n20147_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n20148_));
  AOI21_X1   g19956(.A1(new_n20148_), .A2(new_n20144_), .B(new_n19840_), .ZN(new_n20149_));
  OAI21_X1   g19957(.A1(new_n20149_), .A2(new_n20145_), .B(\asqrt[44] ), .ZN(new_n20150_));
  NAND2_X1   g19958(.A1(new_n20150_), .A2(new_n2641_), .ZN(new_n20151_));
  OAI21_X1   g19959(.A1(new_n20151_), .A2(new_n19851_), .B(new_n20036_), .ZN(new_n20152_));
  AOI21_X1   g19960(.A1(new_n20152_), .A2(new_n19852_), .B(new_n2465_), .ZN(new_n20153_));
  NOR3_X1    g19961(.A1(new_n20149_), .A2(\asqrt[44] ), .A3(new_n20145_), .ZN(new_n20154_));
  OAI21_X1   g19962(.A1(new_n19848_), .A2(new_n20154_), .B(new_n20150_), .ZN(new_n20155_));
  AOI21_X1   g19963(.A1(new_n20155_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n20156_));
  AOI21_X1   g19964(.A1(new_n20156_), .A2(new_n20152_), .B(new_n19866_), .ZN(new_n20157_));
  OAI21_X1   g19965(.A1(new_n20157_), .A2(new_n20153_), .B(\asqrt[47] ), .ZN(new_n20158_));
  NAND2_X1   g19966(.A1(new_n20158_), .A2(new_n1956_), .ZN(new_n20159_));
  OAI21_X1   g19967(.A1(new_n20159_), .A2(new_n19877_), .B(new_n20035_), .ZN(new_n20160_));
  AOI21_X1   g19968(.A1(new_n20160_), .A2(new_n19878_), .B(new_n1806_), .ZN(new_n20161_));
  NOR3_X1    g19969(.A1(new_n20157_), .A2(\asqrt[47] ), .A3(new_n20153_), .ZN(new_n20162_));
  OAI21_X1   g19970(.A1(new_n19874_), .A2(new_n20162_), .B(new_n20158_), .ZN(new_n20163_));
  AOI21_X1   g19971(.A1(new_n20163_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n20164_));
  AOI21_X1   g19972(.A1(new_n20164_), .A2(new_n20160_), .B(new_n19892_), .ZN(new_n20165_));
  OAI21_X1   g19973(.A1(new_n20165_), .A2(new_n20161_), .B(\asqrt[50] ), .ZN(new_n20166_));
  NAND2_X1   g19974(.A1(new_n20166_), .A2(new_n1376_), .ZN(new_n20167_));
  OAI21_X1   g19975(.A1(new_n20167_), .A2(new_n19903_), .B(new_n20034_), .ZN(new_n20168_));
  AOI21_X1   g19976(.A1(new_n20168_), .A2(new_n19904_), .B(new_n1256_), .ZN(new_n20169_));
  NOR3_X1    g19977(.A1(new_n20165_), .A2(\asqrt[50] ), .A3(new_n20161_), .ZN(new_n20170_));
  OAI21_X1   g19978(.A1(new_n19900_), .A2(new_n20170_), .B(new_n20166_), .ZN(new_n20171_));
  AOI21_X1   g19979(.A1(new_n20171_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n20172_));
  AOI21_X1   g19980(.A1(new_n20172_), .A2(new_n20168_), .B(new_n19920_), .ZN(new_n20173_));
  OAI21_X1   g19981(.A1(new_n20173_), .A2(new_n20169_), .B(\asqrt[53] ), .ZN(new_n20174_));
  NAND2_X1   g19982(.A1(new_n20174_), .A2(new_n904_), .ZN(new_n20175_));
  OAI21_X1   g19983(.A1(new_n20175_), .A2(new_n19931_), .B(new_n20033_), .ZN(new_n20176_));
  AOI21_X1   g19984(.A1(new_n20176_), .A2(new_n19932_), .B(new_n823_), .ZN(new_n20177_));
  NOR3_X1    g19985(.A1(new_n20173_), .A2(\asqrt[53] ), .A3(new_n20169_), .ZN(new_n20178_));
  OAI21_X1   g19986(.A1(new_n19928_), .A2(new_n20178_), .B(new_n20174_), .ZN(new_n20179_));
  AOI21_X1   g19987(.A1(new_n20179_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n20180_));
  AOI21_X1   g19988(.A1(new_n20180_), .A2(new_n20176_), .B(new_n19950_), .ZN(new_n20181_));
  OAI21_X1   g19989(.A1(new_n20181_), .A2(new_n20177_), .B(\asqrt[56] ), .ZN(new_n20182_));
  NAND2_X1   g19990(.A1(new_n20182_), .A2(new_n531_), .ZN(new_n20183_));
  OAI21_X1   g19991(.A1(new_n20183_), .A2(new_n19961_), .B(new_n20032_), .ZN(new_n20184_));
  AOI21_X1   g19992(.A1(new_n20184_), .A2(new_n19962_), .B(new_n436_), .ZN(new_n20185_));
  NOR3_X1    g19993(.A1(new_n20181_), .A2(\asqrt[56] ), .A3(new_n20177_), .ZN(new_n20186_));
  OAI21_X1   g19994(.A1(new_n19958_), .A2(new_n20186_), .B(new_n20182_), .ZN(new_n20187_));
  AOI21_X1   g19995(.A1(new_n20187_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n20188_));
  AOI21_X1   g19996(.A1(new_n20188_), .A2(new_n20184_), .B(new_n19981_), .ZN(new_n20189_));
  OAI21_X1   g19997(.A1(new_n20189_), .A2(new_n20185_), .B(\asqrt[59] ), .ZN(new_n20190_));
  NAND2_X1   g19998(.A1(new_n20190_), .A2(new_n306_), .ZN(new_n20191_));
  OAI21_X1   g19999(.A1(new_n20191_), .A2(new_n19992_), .B(new_n20031_), .ZN(new_n20192_));
  NOR3_X1    g20000(.A1(new_n20189_), .A2(\asqrt[59] ), .A3(new_n20185_), .ZN(new_n20193_));
  OAI21_X1   g20001(.A1(new_n19989_), .A2(new_n20193_), .B(new_n20190_), .ZN(new_n20194_));
  AOI21_X1   g20002(.A1(new_n20194_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n20195_));
  AOI21_X1   g20003(.A1(new_n20195_), .A2(new_n20192_), .B(new_n20006_), .ZN(new_n20196_));
  INV_X1     g20004(.I(new_n20014_), .ZN(new_n20197_));
  NAND2_X1   g20005(.A1(new_n20002_), .A2(new_n207_), .ZN(new_n20198_));
  OAI21_X1   g20006(.A1(new_n20198_), .A2(new_n20196_), .B(new_n20197_), .ZN(new_n20199_));
  NOR2_X1    g20007(.A1(new_n20010_), .A2(new_n20026_), .ZN(new_n20200_));
  AOI21_X1   g20008(.A1(\asqrt[8] ), .A2(new_n19495_), .B(new_n19518_), .ZN(new_n20201_));
  OAI21_X1   g20009(.A1(new_n19535_), .A2(new_n19528_), .B(\asqrt[63] ), .ZN(new_n20202_));
  NOR2_X1    g20010(.A1(new_n20201_), .A2(new_n20202_), .ZN(new_n20203_));
  AND2_X2    g20011(.A1(new_n19492_), .A2(new_n19508_), .Z(new_n20204_));
  NAND4_X1   g20012(.A1(new_n19548_), .A2(new_n19494_), .A3(new_n19505_), .A4(new_n20204_), .ZN(new_n20205_));
  NOR2_X1    g20013(.A1(new_n20205_), .A2(new_n19520_), .ZN(new_n20206_));
  NOR2_X1    g20014(.A1(new_n20203_), .A2(new_n20206_), .ZN(new_n20207_));
  INV_X1     g20015(.I(new_n20207_), .ZN(new_n20208_));
  AOI21_X1   g20016(.A1(new_n20200_), .A2(new_n20199_), .B(new_n20208_), .ZN(new_n20209_));
  NAND2_X1   g20017(.A1(new_n20030_), .A2(new_n20209_), .ZN(\asqrt[7] ));
  NOR2_X1    g20018(.A1(\a[12] ), .A2(\a[13] ), .ZN(new_n20211_));
  INV_X1     g20019(.I(new_n20211_), .ZN(new_n20212_));
  NOR2_X1    g20020(.A1(new_n20212_), .A2(\a[14] ), .ZN(new_n20213_));
  INV_X1     g20021(.I(new_n20213_), .ZN(new_n20214_));
  AOI21_X1   g20022(.A1(new_n20192_), .A2(new_n19993_), .B(new_n218_), .ZN(new_n20215_));
  OAI21_X1   g20023(.A1(new_n20196_), .A2(new_n20215_), .B(\asqrt[62] ), .ZN(new_n20216_));
  NOR3_X1    g20024(.A1(new_n20196_), .A2(\asqrt[62] ), .A3(new_n20215_), .ZN(new_n20217_));
  OAI21_X1   g20025(.A1(new_n20014_), .A2(new_n20217_), .B(new_n20216_), .ZN(new_n20218_));
  AOI21_X1   g20026(.A1(new_n20218_), .A2(new_n20028_), .B(\asqrt[63] ), .ZN(new_n20219_));
  NAND2_X1   g20027(.A1(new_n20216_), .A2(new_n20025_), .ZN(new_n20220_));
  OAI21_X1   g20028(.A1(new_n20220_), .A2(new_n20017_), .B(new_n20207_), .ZN(new_n20221_));
  OAI21_X1   g20029(.A1(new_n20219_), .A2(new_n20221_), .B(\a[14] ), .ZN(new_n20222_));
  AOI21_X1   g20030(.A1(new_n20222_), .A2(new_n20214_), .B(new_n19573_), .ZN(new_n20223_));
  INV_X1     g20031(.I(\a[14] ), .ZN(new_n20224_));
  AOI21_X1   g20032(.A1(new_n20030_), .A2(new_n20209_), .B(new_n20224_), .ZN(new_n20225_));
  NAND4_X1   g20033(.A1(new_n19548_), .A2(new_n19505_), .A3(new_n19508_), .A4(new_n20214_), .ZN(new_n20226_));
  NOR2_X1    g20034(.A1(new_n20226_), .A2(new_n19520_), .ZN(new_n20227_));
  INV_X1     g20035(.I(new_n20227_), .ZN(new_n20228_));
  NOR2_X1    g20036(.A1(new_n20225_), .A2(new_n20228_), .ZN(new_n20229_));
  AOI21_X1   g20037(.A1(new_n20030_), .A2(new_n20209_), .B(new_n19515_), .ZN(new_n20230_));
  INV_X1     g20038(.I(\a[15] ), .ZN(new_n20231_));
  AOI21_X1   g20039(.A1(\asqrt[7] ), .A2(new_n20224_), .B(new_n20231_), .ZN(new_n20232_));
  NOR3_X1    g20040(.A1(new_n20229_), .A2(new_n20232_), .A3(new_n20230_), .ZN(new_n20233_));
  OAI21_X1   g20041(.A1(new_n20233_), .A2(new_n20223_), .B(\asqrt[9] ), .ZN(new_n20234_));
  OAI21_X1   g20042(.A1(new_n20219_), .A2(new_n20221_), .B(new_n19514_), .ZN(new_n20235_));
  NOR2_X1    g20043(.A1(new_n20220_), .A2(new_n20017_), .ZN(new_n20236_));
  INV_X1     g20044(.I(new_n20203_), .ZN(new_n20237_));
  NOR2_X1    g20045(.A1(new_n19573_), .A2(new_n20206_), .ZN(new_n20238_));
  NAND2_X1   g20046(.A1(new_n20237_), .A2(new_n20238_), .ZN(new_n20239_));
  NOR3_X1    g20047(.A1(new_n20219_), .A2(new_n20236_), .A3(new_n20239_), .ZN(new_n20240_));
  INV_X1     g20048(.I(new_n20240_), .ZN(new_n20241_));
  AOI21_X1   g20049(.A1(new_n20241_), .A2(new_n20235_), .B(new_n19533_), .ZN(new_n20242_));
  NOR3_X1    g20050(.A1(new_n20240_), .A2(new_n20230_), .A3(\a[16] ), .ZN(new_n20243_));
  OAI21_X1   g20051(.A1(new_n20225_), .A2(new_n20213_), .B(\asqrt[8] ), .ZN(new_n20244_));
  NAND2_X1   g20052(.A1(new_n20244_), .A2(new_n18792_), .ZN(new_n20245_));
  OAI22_X1   g20053(.A1(new_n20233_), .A2(new_n20245_), .B1(new_n20242_), .B2(new_n20243_), .ZN(new_n20246_));
  AOI21_X1   g20054(.A1(new_n20246_), .A2(new_n20234_), .B(new_n18275_), .ZN(new_n20247_));
  NOR3_X1    g20055(.A1(new_n20062_), .A2(new_n19532_), .A3(new_n19541_), .ZN(new_n20248_));
  NAND3_X1   g20056(.A1(\asqrt[7] ), .A2(new_n19562_), .A3(new_n20047_), .ZN(new_n20249_));
  AOI22_X1   g20057(.A1(new_n20249_), .A2(new_n20062_), .B1(\asqrt[7] ), .B2(new_n20248_), .ZN(new_n20250_));
  AOI21_X1   g20058(.A1(new_n20030_), .A2(new_n20209_), .B(\a[14] ), .ZN(new_n20251_));
  OAI21_X1   g20059(.A1(new_n20231_), .A2(new_n20251_), .B(new_n20235_), .ZN(new_n20252_));
  OAI21_X1   g20060(.A1(new_n20252_), .A2(new_n20229_), .B(new_n20244_), .ZN(new_n20253_));
  AOI21_X1   g20061(.A1(new_n20253_), .A2(\asqrt[9] ), .B(\asqrt[10] ), .ZN(new_n20254_));
  AOI21_X1   g20062(.A1(new_n20254_), .A2(new_n20246_), .B(new_n20250_), .ZN(new_n20255_));
  OAI21_X1   g20063(.A1(new_n20255_), .A2(new_n20247_), .B(\asqrt[11] ), .ZN(new_n20256_));
  INV_X1     g20064(.I(new_n20256_), .ZN(new_n20257_));
  NOR2_X1    g20065(.A1(new_n19554_), .A2(new_n19551_), .ZN(new_n20258_));
  NOR2_X1    g20066(.A1(new_n19545_), .A2(new_n19556_), .ZN(new_n20259_));
  INV_X1     g20067(.I(new_n20259_), .ZN(new_n20260_));
  NAND4_X1   g20068(.A1(\asqrt[7] ), .A2(new_n19546_), .A3(new_n20258_), .A4(new_n20260_), .ZN(new_n20261_));
  INV_X1     g20069(.I(\asqrt[7] ), .ZN(new_n20262_));
  NOR3_X1    g20070(.A1(new_n20262_), .A2(new_n20051_), .A3(new_n20259_), .ZN(new_n20263_));
  OAI21_X1   g20071(.A1(new_n20263_), .A2(new_n20258_), .B(new_n20261_), .ZN(new_n20264_));
  INV_X1     g20072(.I(new_n20264_), .ZN(new_n20265_));
  NOR3_X1    g20073(.A1(new_n20255_), .A2(new_n20247_), .A3(\asqrt[11] ), .ZN(new_n20266_));
  NOR2_X1    g20074(.A1(new_n20266_), .A2(new_n20265_), .ZN(new_n20267_));
  OAI21_X1   g20075(.A1(new_n20267_), .A2(new_n20257_), .B(\asqrt[12] ), .ZN(new_n20268_));
  NOR2_X1    g20076(.A1(new_n20064_), .A2(new_n20056_), .ZN(new_n20269_));
  NOR3_X1    g20077(.A1(new_n20262_), .A2(new_n19558_), .A3(new_n20269_), .ZN(new_n20270_));
  INV_X1     g20078(.I(new_n20270_), .ZN(new_n20271_));
  NOR3_X1    g20079(.A1(new_n20269_), .A2(new_n19558_), .A3(new_n20061_), .ZN(new_n20272_));
  AOI22_X1   g20080(.A1(new_n20271_), .A2(new_n20061_), .B1(\asqrt[7] ), .B2(new_n20272_), .ZN(new_n20273_));
  INV_X1     g20081(.I(new_n20273_), .ZN(new_n20274_));
  NAND2_X1   g20082(.A1(new_n20256_), .A2(new_n16881_), .ZN(new_n20275_));
  OAI21_X1   g20083(.A1(new_n20267_), .A2(new_n20275_), .B(new_n20274_), .ZN(new_n20276_));
  AOI21_X1   g20084(.A1(new_n20276_), .A2(new_n20268_), .B(new_n16389_), .ZN(new_n20277_));
  NOR3_X1    g20085(.A1(new_n19569_), .A2(new_n19577_), .A3(new_n19575_), .ZN(new_n20278_));
  NOR3_X1    g20086(.A1(new_n20262_), .A2(new_n19569_), .A3(new_n19577_), .ZN(new_n20279_));
  INV_X1     g20087(.I(new_n20279_), .ZN(new_n20280_));
  AOI22_X1   g20088(.A1(new_n20280_), .A2(new_n19575_), .B1(\asqrt[7] ), .B2(new_n20278_), .ZN(new_n20281_));
  OAI21_X1   g20089(.A1(new_n20265_), .A2(new_n20266_), .B(new_n20256_), .ZN(new_n20282_));
  AOI21_X1   g20090(.A1(new_n20282_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n20283_));
  AOI21_X1   g20091(.A1(new_n20283_), .A2(new_n20276_), .B(new_n20281_), .ZN(new_n20284_));
  OAI21_X1   g20092(.A1(new_n20284_), .A2(new_n20277_), .B(\asqrt[14] ), .ZN(new_n20285_));
  NAND2_X1   g20093(.A1(new_n20067_), .A2(new_n20059_), .ZN(new_n20286_));
  NAND3_X1   g20094(.A1(\asqrt[7] ), .A2(new_n19579_), .A3(new_n20286_), .ZN(new_n20287_));
  AND3_X2    g20095(.A1(new_n19579_), .A2(new_n19583_), .A3(new_n20286_), .Z(new_n20288_));
  AOI22_X1   g20096(.A1(new_n20287_), .A2(new_n19584_), .B1(\asqrt[7] ), .B2(new_n20288_), .ZN(new_n20289_));
  INV_X1     g20097(.I(new_n20289_), .ZN(new_n20290_));
  NAND2_X1   g20098(.A1(new_n20222_), .A2(new_n20227_), .ZN(new_n20291_));
  OAI21_X1   g20099(.A1(new_n20219_), .A2(new_n20221_), .B(new_n20224_), .ZN(new_n20292_));
  NAND2_X1   g20100(.A1(new_n20292_), .A2(\a[15] ), .ZN(new_n20293_));
  NAND3_X1   g20101(.A1(new_n20291_), .A2(new_n20293_), .A3(new_n20235_), .ZN(new_n20294_));
  AOI21_X1   g20102(.A1(new_n20294_), .A2(new_n20244_), .B(new_n18792_), .ZN(new_n20295_));
  OAI21_X1   g20103(.A1(new_n20240_), .A2(new_n20230_), .B(\a[16] ), .ZN(new_n20296_));
  NAND3_X1   g20104(.A1(new_n20241_), .A2(new_n20235_), .A3(new_n19533_), .ZN(new_n20297_));
  NAND2_X1   g20105(.A1(new_n20222_), .A2(new_n20214_), .ZN(new_n20298_));
  AOI21_X1   g20106(.A1(new_n20298_), .A2(\asqrt[8] ), .B(\asqrt[9] ), .ZN(new_n20299_));
  AOI22_X1   g20107(.A1(new_n20294_), .A2(new_n20299_), .B1(new_n20296_), .B2(new_n20297_), .ZN(new_n20300_));
  OAI21_X1   g20108(.A1(new_n20300_), .A2(new_n20295_), .B(\asqrt[10] ), .ZN(new_n20301_));
  NAND2_X1   g20109(.A1(new_n20301_), .A2(new_n17623_), .ZN(new_n20302_));
  OAI21_X1   g20110(.A1(new_n20302_), .A2(new_n20255_), .B(new_n20264_), .ZN(new_n20303_));
  AOI21_X1   g20111(.A1(new_n20303_), .A2(new_n20256_), .B(new_n16881_), .ZN(new_n20304_));
  INV_X1     g20112(.I(new_n20250_), .ZN(new_n20305_));
  AOI21_X1   g20113(.A1(\a[15] ), .A2(new_n20292_), .B(new_n20230_), .ZN(new_n20306_));
  AOI21_X1   g20114(.A1(new_n20306_), .A2(new_n20291_), .B(new_n20223_), .ZN(new_n20307_));
  OAI21_X1   g20115(.A1(new_n20307_), .A2(new_n18792_), .B(new_n18275_), .ZN(new_n20308_));
  OAI21_X1   g20116(.A1(new_n20308_), .A2(new_n20300_), .B(new_n20305_), .ZN(new_n20309_));
  NAND2_X1   g20117(.A1(new_n20309_), .A2(new_n20301_), .ZN(new_n20310_));
  AOI21_X1   g20118(.A1(new_n20310_), .A2(\asqrt[11] ), .B(\asqrt[12] ), .ZN(new_n20311_));
  AOI21_X1   g20119(.A1(new_n20311_), .A2(new_n20303_), .B(new_n20273_), .ZN(new_n20312_));
  OAI21_X1   g20120(.A1(new_n20312_), .A2(new_n20304_), .B(\asqrt[13] ), .ZN(new_n20313_));
  NAND2_X1   g20121(.A1(new_n20313_), .A2(new_n15770_), .ZN(new_n20314_));
  OAI21_X1   g20122(.A1(new_n20314_), .A2(new_n20284_), .B(new_n20290_), .ZN(new_n20315_));
  AOI21_X1   g20123(.A1(new_n20315_), .A2(new_n20285_), .B(new_n15067_), .ZN(new_n20316_));
  INV_X1     g20124(.I(new_n19591_), .ZN(new_n20317_));
  NOR3_X1    g20125(.A1(new_n19587_), .A2(new_n20078_), .A3(new_n20317_), .ZN(new_n20318_));
  NOR3_X1    g20126(.A1(new_n20262_), .A2(new_n19587_), .A3(new_n20078_), .ZN(new_n20319_));
  INV_X1     g20127(.I(new_n20319_), .ZN(new_n20320_));
  AOI22_X1   g20128(.A1(new_n20320_), .A2(new_n20317_), .B1(\asqrt[7] ), .B2(new_n20318_), .ZN(new_n20321_));
  NOR3_X1    g20129(.A1(new_n20312_), .A2(new_n20304_), .A3(\asqrt[13] ), .ZN(new_n20322_));
  OAI21_X1   g20130(.A1(new_n20281_), .A2(new_n20322_), .B(new_n20313_), .ZN(new_n20323_));
  AOI21_X1   g20131(.A1(new_n20323_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n20324_));
  AOI21_X1   g20132(.A1(new_n20324_), .A2(new_n20315_), .B(new_n20321_), .ZN(new_n20325_));
  OAI21_X1   g20133(.A1(new_n20325_), .A2(new_n20316_), .B(\asqrt[16] ), .ZN(new_n20326_));
  INV_X1     g20134(.I(new_n20326_), .ZN(new_n20327_));
  NOR3_X1    g20135(.A1(new_n20262_), .A2(new_n19596_), .A3(new_n19601_), .ZN(new_n20328_));
  INV_X1     g20136(.I(new_n20328_), .ZN(new_n20329_));
  NOR3_X1    g20137(.A1(new_n19596_), .A2(new_n20046_), .A3(new_n19601_), .ZN(new_n20330_));
  AOI22_X1   g20138(.A1(new_n20329_), .A2(new_n20046_), .B1(\asqrt[7] ), .B2(new_n20330_), .ZN(new_n20331_));
  NOR3_X1    g20139(.A1(new_n20325_), .A2(\asqrt[16] ), .A3(new_n20316_), .ZN(new_n20332_));
  NOR2_X1    g20140(.A1(new_n20332_), .A2(new_n20331_), .ZN(new_n20333_));
  OAI21_X1   g20141(.A1(new_n20333_), .A2(new_n20327_), .B(\asqrt[17] ), .ZN(new_n20334_));
  AND3_X2    g20142(.A1(new_n19603_), .A2(new_n19608_), .A3(new_n20072_), .Z(new_n20335_));
  NAND3_X1   g20143(.A1(\asqrt[7] ), .A2(new_n19603_), .A3(new_n20072_), .ZN(new_n20336_));
  AOI22_X1   g20144(.A1(new_n20336_), .A2(new_n19609_), .B1(\asqrt[7] ), .B2(new_n20335_), .ZN(new_n20337_));
  INV_X1     g20145(.I(new_n20337_), .ZN(new_n20338_));
  NAND2_X1   g20146(.A1(new_n20326_), .A2(new_n14017_), .ZN(new_n20339_));
  OAI21_X1   g20147(.A1(new_n20333_), .A2(new_n20339_), .B(new_n20338_), .ZN(new_n20340_));
  AOI21_X1   g20148(.A1(new_n20340_), .A2(new_n20334_), .B(new_n13353_), .ZN(new_n20341_));
  INV_X1     g20149(.I(new_n19616_), .ZN(new_n20342_));
  NOR3_X1    g20150(.A1(new_n20262_), .A2(new_n19612_), .A3(new_n20082_), .ZN(new_n20343_));
  INV_X1     g20151(.I(new_n20343_), .ZN(new_n20344_));
  NOR3_X1    g20152(.A1(new_n19612_), .A2(new_n20082_), .A3(new_n20342_), .ZN(new_n20345_));
  AOI22_X1   g20153(.A1(new_n20344_), .A2(new_n20342_), .B1(\asqrt[7] ), .B2(new_n20345_), .ZN(new_n20346_));
  NOR3_X1    g20154(.A1(new_n20284_), .A2(new_n20277_), .A3(\asqrt[14] ), .ZN(new_n20347_));
  OAI21_X1   g20155(.A1(new_n20289_), .A2(new_n20347_), .B(new_n20285_), .ZN(new_n20348_));
  INV_X1     g20156(.I(new_n20321_), .ZN(new_n20349_));
  NAND3_X1   g20157(.A1(new_n20315_), .A2(new_n15067_), .A3(new_n20285_), .ZN(new_n20350_));
  AOI22_X1   g20158(.A1(new_n20350_), .A2(new_n20349_), .B1(new_n20348_), .B2(\asqrt[15] ), .ZN(new_n20351_));
  OAI22_X1   g20159(.A1(new_n20332_), .A2(new_n20331_), .B1(new_n20351_), .B2(new_n14601_), .ZN(new_n20352_));
  AOI21_X1   g20160(.A1(new_n20352_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n20353_));
  AOI21_X1   g20161(.A1(new_n20353_), .A2(new_n20340_), .B(new_n20346_), .ZN(new_n20354_));
  OAI21_X1   g20162(.A1(new_n20354_), .A2(new_n20341_), .B(\asqrt[19] ), .ZN(new_n20355_));
  INV_X1     g20163(.I(new_n20355_), .ZN(new_n20356_));
  NOR3_X1    g20164(.A1(new_n19621_), .A2(new_n20045_), .A3(new_n19625_), .ZN(new_n20357_));
  NOR3_X1    g20165(.A1(new_n20262_), .A2(new_n19621_), .A3(new_n19625_), .ZN(new_n20358_));
  INV_X1     g20166(.I(new_n20358_), .ZN(new_n20359_));
  AOI22_X1   g20167(.A1(new_n20359_), .A2(new_n20045_), .B1(\asqrt[7] ), .B2(new_n20357_), .ZN(new_n20360_));
  NOR3_X1    g20168(.A1(new_n20354_), .A2(new_n20341_), .A3(\asqrt[19] ), .ZN(new_n20361_));
  NOR2_X1    g20169(.A1(new_n20361_), .A2(new_n20360_), .ZN(new_n20362_));
  OAI21_X1   g20170(.A1(new_n20362_), .A2(new_n20356_), .B(\asqrt[20] ), .ZN(new_n20363_));
  NOR2_X1    g20171(.A1(new_n19626_), .A2(new_n19634_), .ZN(new_n20364_));
  NOR3_X1    g20172(.A1(new_n20262_), .A2(new_n20076_), .A3(new_n20364_), .ZN(new_n20365_));
  INV_X1     g20173(.I(new_n20365_), .ZN(new_n20366_));
  NOR3_X1    g20174(.A1(new_n20364_), .A2(new_n20076_), .A3(new_n19633_), .ZN(new_n20367_));
  AOI22_X1   g20175(.A1(new_n20366_), .A2(new_n19633_), .B1(\asqrt[7] ), .B2(new_n20367_), .ZN(new_n20368_));
  INV_X1     g20176(.I(new_n20368_), .ZN(new_n20369_));
  NAND2_X1   g20177(.A1(new_n20355_), .A2(new_n12364_), .ZN(new_n20370_));
  OAI21_X1   g20178(.A1(new_n20362_), .A2(new_n20370_), .B(new_n20369_), .ZN(new_n20371_));
  AOI21_X1   g20179(.A1(new_n20371_), .A2(new_n20363_), .B(new_n11736_), .ZN(new_n20372_));
  INV_X1     g20180(.I(new_n19640_), .ZN(new_n20373_));
  NOR3_X1    g20181(.A1(new_n19636_), .A2(new_n20090_), .A3(new_n20373_), .ZN(new_n20374_));
  NOR3_X1    g20182(.A1(new_n20262_), .A2(new_n19636_), .A3(new_n20090_), .ZN(new_n20375_));
  INV_X1     g20183(.I(new_n20375_), .ZN(new_n20376_));
  AOI22_X1   g20184(.A1(new_n20376_), .A2(new_n20373_), .B1(\asqrt[7] ), .B2(new_n20374_), .ZN(new_n20377_));
  OAI21_X1   g20185(.A1(new_n20360_), .A2(new_n20361_), .B(new_n20355_), .ZN(new_n20378_));
  AOI21_X1   g20186(.A1(new_n20378_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n20379_));
  AOI21_X1   g20187(.A1(new_n20379_), .A2(new_n20371_), .B(new_n20377_), .ZN(new_n20380_));
  OAI21_X1   g20188(.A1(new_n20380_), .A2(new_n20372_), .B(\asqrt[22] ), .ZN(new_n20381_));
  INV_X1     g20189(.I(new_n20381_), .ZN(new_n20382_));
  NOR3_X1    g20190(.A1(new_n20262_), .A2(new_n19645_), .A3(new_n19651_), .ZN(new_n20383_));
  INV_X1     g20191(.I(new_n20383_), .ZN(new_n20384_));
  NOR3_X1    g20192(.A1(new_n19645_), .A2(new_n20044_), .A3(new_n19651_), .ZN(new_n20385_));
  AOI22_X1   g20193(.A1(new_n20384_), .A2(new_n20044_), .B1(\asqrt[7] ), .B2(new_n20385_), .ZN(new_n20386_));
  NOR3_X1    g20194(.A1(new_n20380_), .A2(new_n20372_), .A3(\asqrt[22] ), .ZN(new_n20387_));
  NOR2_X1    g20195(.A1(new_n20387_), .A2(new_n20386_), .ZN(new_n20388_));
  OAI21_X1   g20196(.A1(new_n20388_), .A2(new_n20382_), .B(\asqrt[23] ), .ZN(new_n20389_));
  NOR2_X1    g20197(.A1(new_n19652_), .A2(new_n19660_), .ZN(new_n20390_));
  NOR3_X1    g20198(.A1(new_n20390_), .A2(new_n20089_), .A3(new_n19659_), .ZN(new_n20391_));
  NOR3_X1    g20199(.A1(new_n20262_), .A2(new_n20089_), .A3(new_n20390_), .ZN(new_n20392_));
  INV_X1     g20200(.I(new_n20392_), .ZN(new_n20393_));
  AOI22_X1   g20201(.A1(new_n20393_), .A2(new_n19659_), .B1(\asqrt[7] ), .B2(new_n20391_), .ZN(new_n20394_));
  INV_X1     g20202(.I(new_n20394_), .ZN(new_n20395_));
  NAND2_X1   g20203(.A1(new_n20381_), .A2(new_n10812_), .ZN(new_n20396_));
  OAI21_X1   g20204(.A1(new_n20388_), .A2(new_n20396_), .B(new_n20395_), .ZN(new_n20397_));
  AOI21_X1   g20205(.A1(new_n20397_), .A2(new_n20389_), .B(new_n10221_), .ZN(new_n20398_));
  INV_X1     g20206(.I(new_n19666_), .ZN(new_n20399_));
  NOR3_X1    g20207(.A1(new_n20262_), .A2(new_n19662_), .A3(new_n20098_), .ZN(new_n20400_));
  INV_X1     g20208(.I(new_n20400_), .ZN(new_n20401_));
  NOR3_X1    g20209(.A1(new_n19662_), .A2(new_n20098_), .A3(new_n20399_), .ZN(new_n20402_));
  AOI22_X1   g20210(.A1(new_n20401_), .A2(new_n20399_), .B1(\asqrt[7] ), .B2(new_n20402_), .ZN(new_n20403_));
  OAI21_X1   g20211(.A1(new_n20386_), .A2(new_n20387_), .B(new_n20381_), .ZN(new_n20404_));
  AOI21_X1   g20212(.A1(new_n20404_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n20405_));
  AOI21_X1   g20213(.A1(new_n20405_), .A2(new_n20397_), .B(new_n20403_), .ZN(new_n20406_));
  OAI21_X1   g20214(.A1(new_n20406_), .A2(new_n20398_), .B(\asqrt[25] ), .ZN(new_n20407_));
  INV_X1     g20215(.I(new_n20407_), .ZN(new_n20408_));
  NOR3_X1    g20216(.A1(new_n19671_), .A2(new_n20043_), .A3(new_n19677_), .ZN(new_n20409_));
  NOR3_X1    g20217(.A1(new_n20262_), .A2(new_n19671_), .A3(new_n19677_), .ZN(new_n20410_));
  INV_X1     g20218(.I(new_n20410_), .ZN(new_n20411_));
  AOI22_X1   g20219(.A1(new_n20411_), .A2(new_n20043_), .B1(\asqrt[7] ), .B2(new_n20409_), .ZN(new_n20412_));
  NOR3_X1    g20220(.A1(new_n20406_), .A2(new_n20398_), .A3(\asqrt[25] ), .ZN(new_n20413_));
  NOR2_X1    g20221(.A1(new_n20413_), .A2(new_n20412_), .ZN(new_n20414_));
  OAI21_X1   g20222(.A1(new_n20414_), .A2(new_n20408_), .B(\asqrt[26] ), .ZN(new_n20415_));
  NOR2_X1    g20223(.A1(new_n19678_), .A2(new_n19686_), .ZN(new_n20416_));
  NOR3_X1    g20224(.A1(new_n20262_), .A2(new_n20097_), .A3(new_n20416_), .ZN(new_n20417_));
  INV_X1     g20225(.I(new_n20417_), .ZN(new_n20418_));
  NOR3_X1    g20226(.A1(new_n20416_), .A2(new_n20097_), .A3(new_n19685_), .ZN(new_n20419_));
  AOI22_X1   g20227(.A1(new_n20418_), .A2(new_n19685_), .B1(\asqrt[7] ), .B2(new_n20419_), .ZN(new_n20420_));
  INV_X1     g20228(.I(new_n20420_), .ZN(new_n20421_));
  NAND2_X1   g20229(.A1(new_n20407_), .A2(new_n9317_), .ZN(new_n20422_));
  OAI21_X1   g20230(.A1(new_n20414_), .A2(new_n20422_), .B(new_n20421_), .ZN(new_n20423_));
  AOI21_X1   g20231(.A1(new_n20423_), .A2(new_n20415_), .B(new_n8826_), .ZN(new_n20424_));
  INV_X1     g20232(.I(new_n19692_), .ZN(new_n20425_));
  NOR3_X1    g20233(.A1(new_n19688_), .A2(new_n20106_), .A3(new_n20425_), .ZN(new_n20426_));
  NOR3_X1    g20234(.A1(new_n20262_), .A2(new_n19688_), .A3(new_n20106_), .ZN(new_n20427_));
  INV_X1     g20235(.I(new_n20427_), .ZN(new_n20428_));
  AOI22_X1   g20236(.A1(new_n20428_), .A2(new_n20425_), .B1(\asqrt[7] ), .B2(new_n20426_), .ZN(new_n20429_));
  OAI21_X1   g20237(.A1(new_n20412_), .A2(new_n20413_), .B(new_n20407_), .ZN(new_n20430_));
  AOI21_X1   g20238(.A1(new_n20430_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n20431_));
  AOI21_X1   g20239(.A1(new_n20431_), .A2(new_n20423_), .B(new_n20429_), .ZN(new_n20432_));
  OAI21_X1   g20240(.A1(new_n20432_), .A2(new_n20424_), .B(\asqrt[28] ), .ZN(new_n20433_));
  INV_X1     g20241(.I(new_n20433_), .ZN(new_n20434_));
  INV_X1     g20242(.I(new_n20432_), .ZN(new_n20435_));
  NOR3_X1    g20243(.A1(new_n20262_), .A2(new_n19697_), .A3(new_n19703_), .ZN(new_n20436_));
  INV_X1     g20244(.I(new_n20436_), .ZN(new_n20437_));
  NOR3_X1    g20245(.A1(new_n19697_), .A2(new_n20042_), .A3(new_n19703_), .ZN(new_n20438_));
  AOI22_X1   g20246(.A1(new_n20437_), .A2(new_n20042_), .B1(\asqrt[7] ), .B2(new_n20438_), .ZN(new_n20439_));
  NOR2_X1    g20247(.A1(new_n20424_), .A2(\asqrt[28] ), .ZN(new_n20440_));
  AOI21_X1   g20248(.A1(new_n20435_), .A2(new_n20440_), .B(new_n20439_), .ZN(new_n20441_));
  OAI21_X1   g20249(.A1(new_n20441_), .A2(new_n20434_), .B(\asqrt[29] ), .ZN(new_n20442_));
  NOR2_X1    g20250(.A1(new_n19704_), .A2(new_n19712_), .ZN(new_n20443_));
  NOR3_X1    g20251(.A1(new_n20443_), .A2(new_n20105_), .A3(new_n19711_), .ZN(new_n20444_));
  NOR3_X1    g20252(.A1(new_n20262_), .A2(new_n20105_), .A3(new_n20443_), .ZN(new_n20445_));
  INV_X1     g20253(.I(new_n20445_), .ZN(new_n20446_));
  AOI22_X1   g20254(.A1(new_n20446_), .A2(new_n19711_), .B1(\asqrt[7] ), .B2(new_n20444_), .ZN(new_n20447_));
  INV_X1     g20255(.I(new_n20447_), .ZN(new_n20448_));
  NAND2_X1   g20256(.A1(new_n20433_), .A2(new_n8036_), .ZN(new_n20449_));
  OAI21_X1   g20257(.A1(new_n20449_), .A2(new_n20441_), .B(new_n20448_), .ZN(new_n20450_));
  AOI21_X1   g20258(.A1(new_n20450_), .A2(new_n20442_), .B(new_n7539_), .ZN(new_n20451_));
  INV_X1     g20259(.I(new_n20451_), .ZN(new_n20452_));
  INV_X1     g20260(.I(new_n20450_), .ZN(new_n20453_));
  INV_X1     g20261(.I(new_n19718_), .ZN(new_n20454_));
  NOR3_X1    g20262(.A1(new_n20262_), .A2(new_n19714_), .A3(new_n20114_), .ZN(new_n20455_));
  INV_X1     g20263(.I(new_n20455_), .ZN(new_n20456_));
  NOR3_X1    g20264(.A1(new_n19714_), .A2(new_n20114_), .A3(new_n20454_), .ZN(new_n20457_));
  AOI22_X1   g20265(.A1(new_n20456_), .A2(new_n20454_), .B1(\asqrt[7] ), .B2(new_n20457_), .ZN(new_n20458_));
  INV_X1     g20266(.I(new_n20458_), .ZN(new_n20459_));
  NAND2_X1   g20267(.A1(new_n20442_), .A2(new_n7539_), .ZN(new_n20460_));
  OAI21_X1   g20268(.A1(new_n20460_), .A2(new_n20453_), .B(new_n20459_), .ZN(new_n20461_));
  AOI21_X1   g20269(.A1(new_n20461_), .A2(new_n20452_), .B(new_n7229_), .ZN(new_n20462_));
  NOR3_X1    g20270(.A1(new_n19723_), .A2(new_n20041_), .A3(new_n19729_), .ZN(new_n20463_));
  NOR3_X1    g20271(.A1(new_n20262_), .A2(new_n19723_), .A3(new_n19729_), .ZN(new_n20464_));
  INV_X1     g20272(.I(new_n20464_), .ZN(new_n20465_));
  AOI22_X1   g20273(.A1(new_n20465_), .A2(new_n20041_), .B1(\asqrt[7] ), .B2(new_n20463_), .ZN(new_n20466_));
  NOR2_X1    g20274(.A1(new_n20451_), .A2(\asqrt[31] ), .ZN(new_n20467_));
  AOI21_X1   g20275(.A1(new_n20467_), .A2(new_n20461_), .B(new_n20466_), .ZN(new_n20468_));
  OAI21_X1   g20276(.A1(new_n20468_), .A2(new_n20462_), .B(\asqrt[32] ), .ZN(new_n20469_));
  NOR2_X1    g20277(.A1(new_n19730_), .A2(new_n19738_), .ZN(new_n20470_));
  NOR3_X1    g20278(.A1(new_n20262_), .A2(new_n20113_), .A3(new_n20470_), .ZN(new_n20471_));
  INV_X1     g20279(.I(new_n20471_), .ZN(new_n20472_));
  NOR3_X1    g20280(.A1(new_n20470_), .A2(new_n20113_), .A3(new_n19737_), .ZN(new_n20473_));
  AOI22_X1   g20281(.A1(new_n20472_), .A2(new_n19737_), .B1(\asqrt[7] ), .B2(new_n20473_), .ZN(new_n20474_));
  INV_X1     g20282(.I(new_n20474_), .ZN(new_n20475_));
  NOR3_X1    g20283(.A1(new_n20432_), .A2(new_n20424_), .A3(\asqrt[28] ), .ZN(new_n20476_));
  OAI21_X1   g20284(.A1(new_n20439_), .A2(new_n20476_), .B(new_n20433_), .ZN(new_n20477_));
  AOI21_X1   g20285(.A1(new_n20477_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n20478_));
  AOI21_X1   g20286(.A1(new_n20478_), .A2(new_n20450_), .B(new_n20458_), .ZN(new_n20479_));
  OAI21_X1   g20287(.A1(new_n20479_), .A2(new_n20451_), .B(\asqrt[31] ), .ZN(new_n20480_));
  NAND2_X1   g20288(.A1(new_n20480_), .A2(new_n6824_), .ZN(new_n20481_));
  OAI21_X1   g20289(.A1(new_n20481_), .A2(new_n20468_), .B(new_n20475_), .ZN(new_n20482_));
  AOI21_X1   g20290(.A1(new_n20482_), .A2(new_n20469_), .B(new_n6356_), .ZN(new_n20483_));
  INV_X1     g20291(.I(new_n20483_), .ZN(new_n20484_));
  INV_X1     g20292(.I(new_n20482_), .ZN(new_n20485_));
  INV_X1     g20293(.I(new_n19744_), .ZN(new_n20486_));
  NOR3_X1    g20294(.A1(new_n19740_), .A2(new_n20122_), .A3(new_n20486_), .ZN(new_n20487_));
  NOR3_X1    g20295(.A1(new_n20262_), .A2(new_n19740_), .A3(new_n20122_), .ZN(new_n20488_));
  INV_X1     g20296(.I(new_n20488_), .ZN(new_n20489_));
  AOI22_X1   g20297(.A1(new_n20489_), .A2(new_n20486_), .B1(\asqrt[7] ), .B2(new_n20487_), .ZN(new_n20490_));
  INV_X1     g20298(.I(new_n20490_), .ZN(new_n20491_));
  NAND2_X1   g20299(.A1(new_n20469_), .A2(new_n6356_), .ZN(new_n20492_));
  OAI21_X1   g20300(.A1(new_n20492_), .A2(new_n20485_), .B(new_n20491_), .ZN(new_n20493_));
  AOI21_X1   g20301(.A1(new_n20493_), .A2(new_n20484_), .B(new_n6077_), .ZN(new_n20494_));
  NOR3_X1    g20302(.A1(new_n20262_), .A2(new_n19749_), .A3(new_n19755_), .ZN(new_n20495_));
  INV_X1     g20303(.I(new_n20495_), .ZN(new_n20496_));
  NOR3_X1    g20304(.A1(new_n19749_), .A2(new_n20040_), .A3(new_n19755_), .ZN(new_n20497_));
  AOI22_X1   g20305(.A1(new_n20496_), .A2(new_n20040_), .B1(\asqrt[7] ), .B2(new_n20497_), .ZN(new_n20498_));
  NOR2_X1    g20306(.A1(new_n20483_), .A2(\asqrt[34] ), .ZN(new_n20499_));
  AOI21_X1   g20307(.A1(new_n20499_), .A2(new_n20493_), .B(new_n20498_), .ZN(new_n20500_));
  OAI21_X1   g20308(.A1(new_n20500_), .A2(new_n20494_), .B(\asqrt[35] ), .ZN(new_n20501_));
  NOR2_X1    g20309(.A1(new_n19756_), .A2(new_n19764_), .ZN(new_n20502_));
  NOR3_X1    g20310(.A1(new_n20502_), .A2(new_n20121_), .A3(new_n19763_), .ZN(new_n20503_));
  NOR3_X1    g20311(.A1(new_n20262_), .A2(new_n20121_), .A3(new_n20502_), .ZN(new_n20504_));
  INV_X1     g20312(.I(new_n20504_), .ZN(new_n20505_));
  AOI22_X1   g20313(.A1(new_n20505_), .A2(new_n19763_), .B1(\asqrt[7] ), .B2(new_n20503_), .ZN(new_n20506_));
  INV_X1     g20314(.I(new_n20506_), .ZN(new_n20507_));
  NOR3_X1    g20315(.A1(new_n20479_), .A2(\asqrt[31] ), .A3(new_n20451_), .ZN(new_n20508_));
  OAI21_X1   g20316(.A1(new_n20466_), .A2(new_n20508_), .B(new_n20480_), .ZN(new_n20509_));
  AOI21_X1   g20317(.A1(new_n20509_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n20510_));
  AOI21_X1   g20318(.A1(new_n20510_), .A2(new_n20482_), .B(new_n20490_), .ZN(new_n20511_));
  OAI21_X1   g20319(.A1(new_n20511_), .A2(new_n20483_), .B(\asqrt[34] ), .ZN(new_n20512_));
  NAND2_X1   g20320(.A1(new_n20512_), .A2(new_n5708_), .ZN(new_n20513_));
  OAI21_X1   g20321(.A1(new_n20513_), .A2(new_n20500_), .B(new_n20507_), .ZN(new_n20514_));
  NAND2_X1   g20322(.A1(new_n20514_), .A2(new_n20501_), .ZN(new_n20515_));
  NAND2_X1   g20323(.A1(new_n20515_), .A2(\asqrt[36] ), .ZN(new_n20516_));
  INV_X1     g20324(.I(new_n20514_), .ZN(new_n20517_));
  INV_X1     g20325(.I(new_n19770_), .ZN(new_n20518_));
  NOR3_X1    g20326(.A1(new_n20262_), .A2(new_n19766_), .A3(new_n20130_), .ZN(new_n20519_));
  INV_X1     g20327(.I(new_n20519_), .ZN(new_n20520_));
  NOR3_X1    g20328(.A1(new_n19766_), .A2(new_n20130_), .A3(new_n20518_), .ZN(new_n20521_));
  AOI22_X1   g20329(.A1(new_n20520_), .A2(new_n20518_), .B1(\asqrt[7] ), .B2(new_n20521_), .ZN(new_n20522_));
  INV_X1     g20330(.I(new_n20522_), .ZN(new_n20523_));
  NAND2_X1   g20331(.A1(new_n20501_), .A2(new_n5277_), .ZN(new_n20524_));
  OAI21_X1   g20332(.A1(new_n20517_), .A2(new_n20524_), .B(new_n20523_), .ZN(new_n20525_));
  AOI21_X1   g20333(.A1(new_n20525_), .A2(new_n20516_), .B(new_n5024_), .ZN(new_n20526_));
  NOR3_X1    g20334(.A1(new_n19775_), .A2(new_n20039_), .A3(new_n19781_), .ZN(new_n20527_));
  NOR3_X1    g20335(.A1(new_n20262_), .A2(new_n19775_), .A3(new_n19781_), .ZN(new_n20528_));
  INV_X1     g20336(.I(new_n20528_), .ZN(new_n20529_));
  AOI22_X1   g20337(.A1(new_n20529_), .A2(new_n20039_), .B1(\asqrt[7] ), .B2(new_n20527_), .ZN(new_n20530_));
  AOI21_X1   g20338(.A1(new_n20514_), .A2(new_n20501_), .B(new_n5277_), .ZN(new_n20531_));
  NOR2_X1    g20339(.A1(new_n20531_), .A2(\asqrt[37] ), .ZN(new_n20532_));
  AOI21_X1   g20340(.A1(new_n20532_), .A2(new_n20525_), .B(new_n20530_), .ZN(new_n20533_));
  OAI21_X1   g20341(.A1(new_n20533_), .A2(new_n20526_), .B(\asqrt[38] ), .ZN(new_n20534_));
  INV_X1     g20342(.I(new_n20534_), .ZN(new_n20535_));
  NOR2_X1    g20343(.A1(new_n19782_), .A2(new_n19790_), .ZN(new_n20536_));
  NOR3_X1    g20344(.A1(new_n20262_), .A2(new_n20129_), .A3(new_n20536_), .ZN(new_n20537_));
  INV_X1     g20345(.I(new_n20537_), .ZN(new_n20538_));
  NOR3_X1    g20346(.A1(new_n20536_), .A2(new_n20129_), .A3(new_n19789_), .ZN(new_n20539_));
  AOI22_X1   g20347(.A1(new_n20538_), .A2(new_n19789_), .B1(\asqrt[7] ), .B2(new_n20539_), .ZN(new_n20540_));
  NOR3_X1    g20348(.A1(new_n20533_), .A2(new_n20526_), .A3(\asqrt[38] ), .ZN(new_n20541_));
  NOR2_X1    g20349(.A1(new_n20541_), .A2(new_n20540_), .ZN(new_n20542_));
  OAI21_X1   g20350(.A1(new_n20542_), .A2(new_n20535_), .B(\asqrt[39] ), .ZN(new_n20543_));
  INV_X1     g20351(.I(new_n19796_), .ZN(new_n20544_));
  NOR3_X1    g20352(.A1(new_n19792_), .A2(new_n20138_), .A3(new_n20544_), .ZN(new_n20545_));
  NOR3_X1    g20353(.A1(new_n20262_), .A2(new_n19792_), .A3(new_n20138_), .ZN(new_n20546_));
  INV_X1     g20354(.I(new_n20546_), .ZN(new_n20547_));
  AOI22_X1   g20355(.A1(new_n20547_), .A2(new_n20544_), .B1(\asqrt[7] ), .B2(new_n20545_), .ZN(new_n20548_));
  INV_X1     g20356(.I(new_n20548_), .ZN(new_n20549_));
  NAND2_X1   g20357(.A1(new_n20534_), .A2(new_n4298_), .ZN(new_n20550_));
  OAI21_X1   g20358(.A1(new_n20542_), .A2(new_n20550_), .B(new_n20549_), .ZN(new_n20551_));
  AOI21_X1   g20359(.A1(new_n20551_), .A2(new_n20543_), .B(new_n4071_), .ZN(new_n20552_));
  NOR3_X1    g20360(.A1(new_n20262_), .A2(new_n19801_), .A3(new_n19807_), .ZN(new_n20553_));
  INV_X1     g20361(.I(new_n20553_), .ZN(new_n20554_));
  NOR3_X1    g20362(.A1(new_n19801_), .A2(new_n20038_), .A3(new_n19807_), .ZN(new_n20555_));
  AOI22_X1   g20363(.A1(new_n20554_), .A2(new_n20038_), .B1(\asqrt[7] ), .B2(new_n20555_), .ZN(new_n20556_));
  INV_X1     g20364(.I(new_n20540_), .ZN(new_n20557_));
  NOR3_X1    g20365(.A1(new_n20511_), .A2(\asqrt[34] ), .A3(new_n20483_), .ZN(new_n20558_));
  OAI21_X1   g20366(.A1(new_n20498_), .A2(new_n20558_), .B(new_n20512_), .ZN(new_n20559_));
  AOI21_X1   g20367(.A1(new_n20559_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n20560_));
  AOI21_X1   g20368(.A1(new_n20560_), .A2(new_n20514_), .B(new_n20522_), .ZN(new_n20561_));
  OAI21_X1   g20369(.A1(new_n20561_), .A2(new_n20531_), .B(\asqrt[37] ), .ZN(new_n20562_));
  NAND2_X1   g20370(.A1(new_n20562_), .A2(new_n4696_), .ZN(new_n20563_));
  OAI21_X1   g20371(.A1(new_n20563_), .A2(new_n20533_), .B(new_n20557_), .ZN(new_n20564_));
  AOI21_X1   g20372(.A1(new_n20564_), .A2(new_n20534_), .B(new_n4298_), .ZN(new_n20565_));
  NOR2_X1    g20373(.A1(new_n20565_), .A2(\asqrt[40] ), .ZN(new_n20566_));
  AOI21_X1   g20374(.A1(new_n20566_), .A2(new_n20551_), .B(new_n20556_), .ZN(new_n20567_));
  OAI21_X1   g20375(.A1(new_n20567_), .A2(new_n20552_), .B(\asqrt[41] ), .ZN(new_n20568_));
  NOR2_X1    g20376(.A1(new_n19808_), .A2(new_n19816_), .ZN(new_n20569_));
  NOR3_X1    g20377(.A1(new_n20569_), .A2(new_n20137_), .A3(new_n19815_), .ZN(new_n20570_));
  NOR3_X1    g20378(.A1(new_n20262_), .A2(new_n20137_), .A3(new_n20569_), .ZN(new_n20571_));
  INV_X1     g20379(.I(new_n20571_), .ZN(new_n20572_));
  AOI22_X1   g20380(.A1(new_n20572_), .A2(new_n19815_), .B1(\asqrt[7] ), .B2(new_n20570_), .ZN(new_n20573_));
  INV_X1     g20381(.I(new_n20573_), .ZN(new_n20574_));
  NOR3_X1    g20382(.A1(new_n20561_), .A2(\asqrt[37] ), .A3(new_n20531_), .ZN(new_n20575_));
  OAI21_X1   g20383(.A1(new_n20530_), .A2(new_n20575_), .B(new_n20562_), .ZN(new_n20576_));
  AOI21_X1   g20384(.A1(new_n20576_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n20577_));
  AOI21_X1   g20385(.A1(new_n20577_), .A2(new_n20564_), .B(new_n20548_), .ZN(new_n20578_));
  OAI21_X1   g20386(.A1(new_n20578_), .A2(new_n20565_), .B(\asqrt[40] ), .ZN(new_n20579_));
  NAND2_X1   g20387(.A1(new_n20579_), .A2(new_n3782_), .ZN(new_n20580_));
  OAI21_X1   g20388(.A1(new_n20580_), .A2(new_n20567_), .B(new_n20574_), .ZN(new_n20581_));
  AOI21_X1   g20389(.A1(new_n20581_), .A2(new_n20568_), .B(new_n3419_), .ZN(new_n20582_));
  INV_X1     g20390(.I(new_n19822_), .ZN(new_n20583_));
  NOR3_X1    g20391(.A1(new_n20262_), .A2(new_n19818_), .A3(new_n20146_), .ZN(new_n20584_));
  INV_X1     g20392(.I(new_n20584_), .ZN(new_n20585_));
  NOR3_X1    g20393(.A1(new_n19818_), .A2(new_n20146_), .A3(new_n20583_), .ZN(new_n20586_));
  AOI22_X1   g20394(.A1(new_n20585_), .A2(new_n20583_), .B1(\asqrt[7] ), .B2(new_n20586_), .ZN(new_n20587_));
  NOR3_X1    g20395(.A1(new_n20578_), .A2(\asqrt[40] ), .A3(new_n20565_), .ZN(new_n20588_));
  OAI21_X1   g20396(.A1(new_n20556_), .A2(new_n20588_), .B(new_n20579_), .ZN(new_n20589_));
  AOI21_X1   g20397(.A1(new_n20589_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n20590_));
  AOI21_X1   g20398(.A1(new_n20590_), .A2(new_n20581_), .B(new_n20587_), .ZN(new_n20591_));
  OAI21_X1   g20399(.A1(new_n20591_), .A2(new_n20582_), .B(\asqrt[43] ), .ZN(new_n20592_));
  INV_X1     g20400(.I(new_n20592_), .ZN(new_n20593_));
  NOR3_X1    g20401(.A1(new_n19827_), .A2(new_n20037_), .A3(new_n19833_), .ZN(new_n20594_));
  NOR3_X1    g20402(.A1(new_n20262_), .A2(new_n19827_), .A3(new_n19833_), .ZN(new_n20595_));
  INV_X1     g20403(.I(new_n20595_), .ZN(new_n20596_));
  AOI22_X1   g20404(.A1(new_n20596_), .A2(new_n20037_), .B1(\asqrt[7] ), .B2(new_n20594_), .ZN(new_n20597_));
  NOR3_X1    g20405(.A1(new_n20591_), .A2(\asqrt[43] ), .A3(new_n20582_), .ZN(new_n20598_));
  NOR2_X1    g20406(.A1(new_n20598_), .A2(new_n20597_), .ZN(new_n20599_));
  OAI21_X1   g20407(.A1(new_n20599_), .A2(new_n20593_), .B(\asqrt[44] ), .ZN(new_n20600_));
  NOR2_X1    g20408(.A1(new_n19834_), .A2(new_n19842_), .ZN(new_n20601_));
  NOR3_X1    g20409(.A1(new_n20262_), .A2(new_n20145_), .A3(new_n20601_), .ZN(new_n20602_));
  INV_X1     g20410(.I(new_n20602_), .ZN(new_n20603_));
  NOR3_X1    g20411(.A1(new_n20601_), .A2(new_n20145_), .A3(new_n19841_), .ZN(new_n20604_));
  AOI22_X1   g20412(.A1(new_n20603_), .A2(new_n19841_), .B1(\asqrt[7] ), .B2(new_n20604_), .ZN(new_n20605_));
  INV_X1     g20413(.I(new_n20605_), .ZN(new_n20606_));
  NAND2_X1   g20414(.A1(new_n20592_), .A2(new_n2954_), .ZN(new_n20607_));
  OAI21_X1   g20415(.A1(new_n20599_), .A2(new_n20607_), .B(new_n20606_), .ZN(new_n20608_));
  AOI21_X1   g20416(.A1(new_n20608_), .A2(new_n20600_), .B(new_n2641_), .ZN(new_n20609_));
  INV_X1     g20417(.I(new_n19848_), .ZN(new_n20610_));
  NOR3_X1    g20418(.A1(new_n19844_), .A2(new_n20154_), .A3(new_n20610_), .ZN(new_n20611_));
  NOR3_X1    g20419(.A1(new_n20262_), .A2(new_n19844_), .A3(new_n20154_), .ZN(new_n20612_));
  INV_X1     g20420(.I(new_n20612_), .ZN(new_n20613_));
  AOI22_X1   g20421(.A1(new_n20613_), .A2(new_n20610_), .B1(\asqrt[7] ), .B2(new_n20611_), .ZN(new_n20614_));
  OAI21_X1   g20422(.A1(new_n20597_), .A2(new_n20598_), .B(new_n20592_), .ZN(new_n20615_));
  AOI21_X1   g20423(.A1(new_n20615_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n20616_));
  AOI21_X1   g20424(.A1(new_n20616_), .A2(new_n20608_), .B(new_n20614_), .ZN(new_n20617_));
  OAI21_X1   g20425(.A1(new_n20617_), .A2(new_n20609_), .B(\asqrt[46] ), .ZN(new_n20618_));
  INV_X1     g20426(.I(new_n20618_), .ZN(new_n20619_));
  NOR3_X1    g20427(.A1(new_n20262_), .A2(new_n19853_), .A3(new_n19859_), .ZN(new_n20620_));
  INV_X1     g20428(.I(new_n20620_), .ZN(new_n20621_));
  NOR3_X1    g20429(.A1(new_n19853_), .A2(new_n20036_), .A3(new_n19859_), .ZN(new_n20622_));
  AOI22_X1   g20430(.A1(new_n20621_), .A2(new_n20036_), .B1(\asqrt[7] ), .B2(new_n20622_), .ZN(new_n20623_));
  NOR3_X1    g20431(.A1(new_n20617_), .A2(new_n20609_), .A3(\asqrt[46] ), .ZN(new_n20624_));
  NOR2_X1    g20432(.A1(new_n20624_), .A2(new_n20623_), .ZN(new_n20625_));
  OAI21_X1   g20433(.A1(new_n20625_), .A2(new_n20619_), .B(\asqrt[47] ), .ZN(new_n20626_));
  NOR2_X1    g20434(.A1(new_n19860_), .A2(new_n19868_), .ZN(new_n20627_));
  NOR3_X1    g20435(.A1(new_n20627_), .A2(new_n20153_), .A3(new_n19867_), .ZN(new_n20628_));
  NOR3_X1    g20436(.A1(new_n20262_), .A2(new_n20153_), .A3(new_n20627_), .ZN(new_n20629_));
  INV_X1     g20437(.I(new_n20629_), .ZN(new_n20630_));
  AOI22_X1   g20438(.A1(new_n20630_), .A2(new_n19867_), .B1(\asqrt[7] ), .B2(new_n20628_), .ZN(new_n20631_));
  INV_X1     g20439(.I(new_n20631_), .ZN(new_n20632_));
  NAND2_X1   g20440(.A1(new_n20618_), .A2(new_n2229_), .ZN(new_n20633_));
  OAI21_X1   g20441(.A1(new_n20625_), .A2(new_n20633_), .B(new_n20632_), .ZN(new_n20634_));
  AOI21_X1   g20442(.A1(new_n20634_), .A2(new_n20626_), .B(new_n1956_), .ZN(new_n20635_));
  INV_X1     g20443(.I(new_n19874_), .ZN(new_n20636_));
  NOR3_X1    g20444(.A1(new_n20262_), .A2(new_n19870_), .A3(new_n20162_), .ZN(new_n20637_));
  INV_X1     g20445(.I(new_n20637_), .ZN(new_n20638_));
  NOR3_X1    g20446(.A1(new_n19870_), .A2(new_n20162_), .A3(new_n20636_), .ZN(new_n20639_));
  AOI22_X1   g20447(.A1(new_n20638_), .A2(new_n20636_), .B1(\asqrt[7] ), .B2(new_n20639_), .ZN(new_n20640_));
  OAI21_X1   g20448(.A1(new_n20623_), .A2(new_n20624_), .B(new_n20618_), .ZN(new_n20641_));
  AOI21_X1   g20449(.A1(new_n20641_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n20642_));
  AOI21_X1   g20450(.A1(new_n20642_), .A2(new_n20634_), .B(new_n20640_), .ZN(new_n20643_));
  OAI21_X1   g20451(.A1(new_n20643_), .A2(new_n20635_), .B(\asqrt[49] ), .ZN(new_n20644_));
  INV_X1     g20452(.I(new_n20644_), .ZN(new_n20645_));
  NOR3_X1    g20453(.A1(new_n19879_), .A2(new_n20035_), .A3(new_n19885_), .ZN(new_n20646_));
  NOR3_X1    g20454(.A1(new_n20262_), .A2(new_n19879_), .A3(new_n19885_), .ZN(new_n20647_));
  INV_X1     g20455(.I(new_n20647_), .ZN(new_n20648_));
  AOI22_X1   g20456(.A1(new_n20648_), .A2(new_n20035_), .B1(\asqrt[7] ), .B2(new_n20646_), .ZN(new_n20649_));
  NOR3_X1    g20457(.A1(new_n20643_), .A2(new_n20635_), .A3(\asqrt[49] ), .ZN(new_n20650_));
  NOR2_X1    g20458(.A1(new_n20650_), .A2(new_n20649_), .ZN(new_n20651_));
  OAI21_X1   g20459(.A1(new_n20651_), .A2(new_n20645_), .B(\asqrt[50] ), .ZN(new_n20652_));
  NOR2_X1    g20460(.A1(new_n19886_), .A2(new_n19894_), .ZN(new_n20653_));
  NOR3_X1    g20461(.A1(new_n20262_), .A2(new_n20161_), .A3(new_n20653_), .ZN(new_n20654_));
  INV_X1     g20462(.I(new_n20654_), .ZN(new_n20655_));
  NOR3_X1    g20463(.A1(new_n20653_), .A2(new_n20161_), .A3(new_n19893_), .ZN(new_n20656_));
  AOI22_X1   g20464(.A1(new_n20655_), .A2(new_n19893_), .B1(\asqrt[7] ), .B2(new_n20656_), .ZN(new_n20657_));
  INV_X1     g20465(.I(new_n20657_), .ZN(new_n20658_));
  NAND2_X1   g20466(.A1(new_n20644_), .A2(new_n1612_), .ZN(new_n20659_));
  OAI21_X1   g20467(.A1(new_n20651_), .A2(new_n20659_), .B(new_n20658_), .ZN(new_n20660_));
  AOI21_X1   g20468(.A1(new_n20660_), .A2(new_n20652_), .B(new_n1376_), .ZN(new_n20661_));
  INV_X1     g20469(.I(new_n19900_), .ZN(new_n20662_));
  NOR3_X1    g20470(.A1(new_n19896_), .A2(new_n20170_), .A3(new_n20662_), .ZN(new_n20663_));
  NOR3_X1    g20471(.A1(new_n20262_), .A2(new_n19896_), .A3(new_n20170_), .ZN(new_n20664_));
  INV_X1     g20472(.I(new_n20664_), .ZN(new_n20665_));
  AOI22_X1   g20473(.A1(new_n20665_), .A2(new_n20662_), .B1(\asqrt[7] ), .B2(new_n20663_), .ZN(new_n20666_));
  OAI21_X1   g20474(.A1(new_n20649_), .A2(new_n20650_), .B(new_n20644_), .ZN(new_n20667_));
  AOI21_X1   g20475(.A1(new_n20667_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n20668_));
  AOI21_X1   g20476(.A1(new_n20668_), .A2(new_n20660_), .B(new_n20666_), .ZN(new_n20669_));
  OAI21_X1   g20477(.A1(new_n20669_), .A2(new_n20661_), .B(\asqrt[52] ), .ZN(new_n20670_));
  INV_X1     g20478(.I(new_n20670_), .ZN(new_n20671_));
  INV_X1     g20479(.I(new_n20669_), .ZN(new_n20672_));
  NOR3_X1    g20480(.A1(new_n20262_), .A2(new_n19905_), .A3(new_n19911_), .ZN(new_n20673_));
  INV_X1     g20481(.I(new_n20673_), .ZN(new_n20674_));
  NOR3_X1    g20482(.A1(new_n19905_), .A2(new_n20034_), .A3(new_n19911_), .ZN(new_n20675_));
  AOI22_X1   g20483(.A1(new_n20674_), .A2(new_n20034_), .B1(\asqrt[7] ), .B2(new_n20675_), .ZN(new_n20676_));
  NOR2_X1    g20484(.A1(new_n20661_), .A2(\asqrt[52] ), .ZN(new_n20677_));
  AOI21_X1   g20485(.A1(new_n20672_), .A2(new_n20677_), .B(new_n20676_), .ZN(new_n20678_));
  OAI21_X1   g20486(.A1(new_n20678_), .A2(new_n20671_), .B(\asqrt[53] ), .ZN(new_n20679_));
  NOR2_X1    g20487(.A1(new_n19912_), .A2(new_n19922_), .ZN(new_n20680_));
  NOR3_X1    g20488(.A1(new_n20680_), .A2(new_n20169_), .A3(new_n19921_), .ZN(new_n20681_));
  NOR3_X1    g20489(.A1(new_n20262_), .A2(new_n20169_), .A3(new_n20680_), .ZN(new_n20682_));
  INV_X1     g20490(.I(new_n20682_), .ZN(new_n20683_));
  AOI22_X1   g20491(.A1(new_n20683_), .A2(new_n19921_), .B1(\asqrt[7] ), .B2(new_n20681_), .ZN(new_n20684_));
  INV_X1     g20492(.I(new_n20684_), .ZN(new_n20685_));
  NAND2_X1   g20493(.A1(new_n20670_), .A2(new_n1103_), .ZN(new_n20686_));
  OAI21_X1   g20494(.A1(new_n20686_), .A2(new_n20678_), .B(new_n20685_), .ZN(new_n20687_));
  AOI21_X1   g20495(.A1(new_n20687_), .A2(new_n20679_), .B(new_n904_), .ZN(new_n20688_));
  INV_X1     g20496(.I(new_n20688_), .ZN(new_n20689_));
  INV_X1     g20497(.I(new_n20687_), .ZN(new_n20690_));
  INV_X1     g20498(.I(new_n19928_), .ZN(new_n20691_));
  NOR3_X1    g20499(.A1(new_n20262_), .A2(new_n19924_), .A3(new_n20178_), .ZN(new_n20692_));
  INV_X1     g20500(.I(new_n20692_), .ZN(new_n20693_));
  NOR3_X1    g20501(.A1(new_n19924_), .A2(new_n20178_), .A3(new_n20691_), .ZN(new_n20694_));
  AOI22_X1   g20502(.A1(new_n20693_), .A2(new_n20691_), .B1(\asqrt[7] ), .B2(new_n20694_), .ZN(new_n20695_));
  INV_X1     g20503(.I(new_n20695_), .ZN(new_n20696_));
  NAND2_X1   g20504(.A1(new_n20679_), .A2(new_n904_), .ZN(new_n20697_));
  OAI21_X1   g20505(.A1(new_n20697_), .A2(new_n20690_), .B(new_n20696_), .ZN(new_n20698_));
  AOI21_X1   g20506(.A1(new_n20698_), .A2(new_n20689_), .B(new_n823_), .ZN(new_n20699_));
  NOR3_X1    g20507(.A1(new_n19933_), .A2(new_n20033_), .A3(new_n19940_), .ZN(new_n20700_));
  NOR3_X1    g20508(.A1(new_n20262_), .A2(new_n19933_), .A3(new_n19940_), .ZN(new_n20701_));
  INV_X1     g20509(.I(new_n20701_), .ZN(new_n20702_));
  AOI22_X1   g20510(.A1(new_n20702_), .A2(new_n20033_), .B1(\asqrt[7] ), .B2(new_n20700_), .ZN(new_n20703_));
  NOR2_X1    g20511(.A1(new_n20688_), .A2(\asqrt[55] ), .ZN(new_n20704_));
  AOI21_X1   g20512(.A1(new_n20704_), .A2(new_n20698_), .B(new_n20703_), .ZN(new_n20705_));
  OAI21_X1   g20513(.A1(new_n20705_), .A2(new_n20699_), .B(\asqrt[56] ), .ZN(new_n20706_));
  NOR2_X1    g20514(.A1(new_n19941_), .A2(new_n19952_), .ZN(new_n20707_));
  NOR3_X1    g20515(.A1(new_n20262_), .A2(new_n20177_), .A3(new_n20707_), .ZN(new_n20708_));
  INV_X1     g20516(.I(new_n20708_), .ZN(new_n20709_));
  NOR3_X1    g20517(.A1(new_n20707_), .A2(new_n20177_), .A3(new_n19951_), .ZN(new_n20710_));
  AOI22_X1   g20518(.A1(new_n20709_), .A2(new_n19951_), .B1(\asqrt[7] ), .B2(new_n20710_), .ZN(new_n20711_));
  INV_X1     g20519(.I(new_n20711_), .ZN(new_n20712_));
  NOR3_X1    g20520(.A1(new_n20669_), .A2(new_n20661_), .A3(\asqrt[52] ), .ZN(new_n20713_));
  OAI21_X1   g20521(.A1(new_n20676_), .A2(new_n20713_), .B(new_n20670_), .ZN(new_n20714_));
  AOI21_X1   g20522(.A1(new_n20714_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n20715_));
  AOI21_X1   g20523(.A1(new_n20715_), .A2(new_n20687_), .B(new_n20695_), .ZN(new_n20716_));
  OAI21_X1   g20524(.A1(new_n20716_), .A2(new_n20688_), .B(\asqrt[55] ), .ZN(new_n20717_));
  NAND2_X1   g20525(.A1(new_n20717_), .A2(new_n703_), .ZN(new_n20718_));
  OAI21_X1   g20526(.A1(new_n20718_), .A2(new_n20705_), .B(new_n20712_), .ZN(new_n20719_));
  AOI21_X1   g20527(.A1(new_n20719_), .A2(new_n20706_), .B(new_n531_), .ZN(new_n20720_));
  INV_X1     g20528(.I(new_n20720_), .ZN(new_n20721_));
  INV_X1     g20529(.I(new_n20719_), .ZN(new_n20722_));
  INV_X1     g20530(.I(new_n19958_), .ZN(new_n20723_));
  NOR3_X1    g20531(.A1(new_n19954_), .A2(new_n20186_), .A3(new_n20723_), .ZN(new_n20724_));
  NOR3_X1    g20532(.A1(new_n20262_), .A2(new_n19954_), .A3(new_n20186_), .ZN(new_n20725_));
  INV_X1     g20533(.I(new_n20725_), .ZN(new_n20726_));
  AOI22_X1   g20534(.A1(new_n20726_), .A2(new_n20723_), .B1(\asqrt[7] ), .B2(new_n20724_), .ZN(new_n20727_));
  INV_X1     g20535(.I(new_n20727_), .ZN(new_n20728_));
  NAND2_X1   g20536(.A1(new_n20706_), .A2(new_n531_), .ZN(new_n20729_));
  OAI21_X1   g20537(.A1(new_n20729_), .A2(new_n20722_), .B(new_n20728_), .ZN(new_n20730_));
  AOI21_X1   g20538(.A1(new_n20730_), .A2(new_n20721_), .B(new_n436_), .ZN(new_n20731_));
  NOR3_X1    g20539(.A1(new_n20262_), .A2(new_n19963_), .A3(new_n19970_), .ZN(new_n20732_));
  INV_X1     g20540(.I(new_n20732_), .ZN(new_n20733_));
  NOR3_X1    g20541(.A1(new_n19963_), .A2(new_n20032_), .A3(new_n19970_), .ZN(new_n20734_));
  AOI22_X1   g20542(.A1(new_n20733_), .A2(new_n20032_), .B1(\asqrt[7] ), .B2(new_n20734_), .ZN(new_n20735_));
  NOR2_X1    g20543(.A1(new_n20720_), .A2(\asqrt[58] ), .ZN(new_n20736_));
  AOI21_X1   g20544(.A1(new_n20736_), .A2(new_n20730_), .B(new_n20735_), .ZN(new_n20737_));
  OAI21_X1   g20545(.A1(new_n20737_), .A2(new_n20731_), .B(\asqrt[59] ), .ZN(new_n20738_));
  NOR2_X1    g20546(.A1(new_n19971_), .A2(new_n19983_), .ZN(new_n20739_));
  NOR3_X1    g20547(.A1(new_n20739_), .A2(new_n20185_), .A3(new_n19982_), .ZN(new_n20740_));
  NOR3_X1    g20548(.A1(new_n20262_), .A2(new_n20185_), .A3(new_n20739_), .ZN(new_n20741_));
  INV_X1     g20549(.I(new_n20741_), .ZN(new_n20742_));
  AOI22_X1   g20550(.A1(new_n20742_), .A2(new_n19982_), .B1(\asqrt[7] ), .B2(new_n20740_), .ZN(new_n20743_));
  INV_X1     g20551(.I(new_n20743_), .ZN(new_n20744_));
  NOR3_X1    g20552(.A1(new_n20716_), .A2(\asqrt[55] ), .A3(new_n20688_), .ZN(new_n20745_));
  OAI21_X1   g20553(.A1(new_n20703_), .A2(new_n20745_), .B(new_n20717_), .ZN(new_n20746_));
  AOI21_X1   g20554(.A1(new_n20746_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n20747_));
  AOI21_X1   g20555(.A1(new_n20747_), .A2(new_n20719_), .B(new_n20727_), .ZN(new_n20748_));
  OAI21_X1   g20556(.A1(new_n20748_), .A2(new_n20720_), .B(\asqrt[58] ), .ZN(new_n20749_));
  NAND2_X1   g20557(.A1(new_n20749_), .A2(new_n327_), .ZN(new_n20750_));
  OAI21_X1   g20558(.A1(new_n20750_), .A2(new_n20737_), .B(new_n20744_), .ZN(new_n20751_));
  AOI21_X1   g20559(.A1(new_n20751_), .A2(new_n20738_), .B(new_n306_), .ZN(new_n20752_));
  INV_X1     g20560(.I(new_n20752_), .ZN(new_n20753_));
  INV_X1     g20561(.I(new_n20751_), .ZN(new_n20754_));
  INV_X1     g20562(.I(new_n19989_), .ZN(new_n20755_));
  NOR3_X1    g20563(.A1(new_n20262_), .A2(new_n19985_), .A3(new_n20193_), .ZN(new_n20756_));
  INV_X1     g20564(.I(new_n20756_), .ZN(new_n20757_));
  NOR3_X1    g20565(.A1(new_n19985_), .A2(new_n20193_), .A3(new_n20755_), .ZN(new_n20758_));
  AOI22_X1   g20566(.A1(new_n20757_), .A2(new_n20755_), .B1(\asqrt[7] ), .B2(new_n20758_), .ZN(new_n20759_));
  INV_X1     g20567(.I(new_n20759_), .ZN(new_n20760_));
  NAND2_X1   g20568(.A1(new_n20738_), .A2(new_n306_), .ZN(new_n20761_));
  OAI21_X1   g20569(.A1(new_n20754_), .A2(new_n20761_), .B(new_n20760_), .ZN(new_n20762_));
  AOI21_X1   g20570(.A1(new_n20762_), .A2(new_n20753_), .B(new_n218_), .ZN(new_n20763_));
  NOR3_X1    g20571(.A1(new_n19994_), .A2(new_n20031_), .A3(new_n20000_), .ZN(new_n20764_));
  NOR3_X1    g20572(.A1(new_n20262_), .A2(new_n19994_), .A3(new_n20000_), .ZN(new_n20765_));
  INV_X1     g20573(.I(new_n20765_), .ZN(new_n20766_));
  AOI22_X1   g20574(.A1(new_n20766_), .A2(new_n20031_), .B1(\asqrt[7] ), .B2(new_n20764_), .ZN(new_n20767_));
  NOR2_X1    g20575(.A1(new_n20752_), .A2(\asqrt[61] ), .ZN(new_n20768_));
  AOI21_X1   g20576(.A1(new_n20768_), .A2(new_n20762_), .B(new_n20767_), .ZN(new_n20769_));
  OAI21_X1   g20577(.A1(new_n20769_), .A2(new_n20763_), .B(\asqrt[62] ), .ZN(new_n20770_));
  NOR2_X1    g20578(.A1(new_n20001_), .A2(new_n20008_), .ZN(new_n20771_));
  NOR3_X1    g20579(.A1(new_n20262_), .A2(new_n20215_), .A3(new_n20771_), .ZN(new_n20772_));
  INV_X1     g20580(.I(new_n20772_), .ZN(new_n20773_));
  NOR3_X1    g20581(.A1(new_n20771_), .A2(new_n20215_), .A3(new_n20007_), .ZN(new_n20774_));
  AOI22_X1   g20582(.A1(new_n20773_), .A2(new_n20007_), .B1(\asqrt[7] ), .B2(new_n20774_), .ZN(new_n20775_));
  INV_X1     g20583(.I(new_n20775_), .ZN(new_n20776_));
  NOR3_X1    g20584(.A1(new_n20748_), .A2(\asqrt[58] ), .A3(new_n20720_), .ZN(new_n20777_));
  OAI21_X1   g20585(.A1(new_n20735_), .A2(new_n20777_), .B(new_n20749_), .ZN(new_n20778_));
  AOI21_X1   g20586(.A1(new_n20778_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n20779_));
  AOI21_X1   g20587(.A1(new_n20779_), .A2(new_n20751_), .B(new_n20759_), .ZN(new_n20780_));
  OAI21_X1   g20588(.A1(new_n20780_), .A2(new_n20752_), .B(\asqrt[61] ), .ZN(new_n20781_));
  NAND2_X1   g20589(.A1(new_n20781_), .A2(new_n207_), .ZN(new_n20782_));
  OAI21_X1   g20590(.A1(new_n20782_), .A2(new_n20769_), .B(new_n20776_), .ZN(new_n20783_));
  INV_X1     g20591(.I(new_n20217_), .ZN(new_n20784_));
  NAND4_X1   g20592(.A1(\asqrt[7] ), .A2(new_n20216_), .A3(new_n20014_), .A4(new_n20784_), .ZN(new_n20785_));
  NAND2_X1   g20593(.A1(new_n20784_), .A2(new_n20216_), .ZN(new_n20786_));
  OAI21_X1   g20594(.A1(new_n20262_), .A2(new_n20786_), .B(new_n20197_), .ZN(new_n20787_));
  NAND2_X1   g20595(.A1(new_n20787_), .A2(new_n20785_), .ZN(new_n20788_));
  AOI21_X1   g20596(.A1(new_n20199_), .A2(new_n20216_), .B(new_n20025_), .ZN(new_n20789_));
  AOI21_X1   g20597(.A1(\asqrt[7] ), .A2(new_n20789_), .B(new_n20236_), .ZN(new_n20790_));
  NAND2_X1   g20598(.A1(new_n20788_), .A2(new_n20790_), .ZN(new_n20791_));
  AOI21_X1   g20599(.A1(new_n20783_), .A2(new_n20770_), .B(new_n20791_), .ZN(new_n20792_));
  NOR2_X1    g20600(.A1(new_n20792_), .A2(\asqrt[63] ), .ZN(new_n20793_));
  INV_X1     g20601(.I(new_n20783_), .ZN(new_n20794_));
  INV_X1     g20602(.I(new_n20788_), .ZN(new_n20795_));
  NAND2_X1   g20603(.A1(new_n20770_), .A2(new_n20795_), .ZN(new_n20796_));
  AOI21_X1   g20604(.A1(\asqrt[7] ), .A2(new_n20026_), .B(new_n20218_), .ZN(new_n20797_));
  OR3_X2     g20605(.A1(new_n20797_), .A2(new_n193_), .A3(new_n20789_), .Z(new_n20798_));
  INV_X1     g20606(.I(new_n20206_), .ZN(new_n20799_));
  NAND2_X1   g20607(.A1(new_n20799_), .A2(new_n20021_), .ZN(new_n20800_));
  NOR4_X1    g20608(.A1(new_n20236_), .A2(new_n20024_), .A3(new_n20203_), .A4(new_n20800_), .ZN(new_n20801_));
  NAND2_X1   g20609(.A1(new_n20801_), .A2(new_n20030_), .ZN(new_n20802_));
  NAND2_X1   g20610(.A1(new_n20798_), .A2(new_n20802_), .ZN(new_n20803_));
  INV_X1     g20611(.I(new_n20803_), .ZN(new_n20804_));
  OAI21_X1   g20612(.A1(new_n20794_), .A2(new_n20796_), .B(new_n20804_), .ZN(new_n20805_));
  NOR2_X1    g20613(.A1(new_n20793_), .A2(new_n20805_), .ZN(new_n20806_));
  INV_X1     g20614(.I(\a[12] ), .ZN(new_n20807_));
  NOR2_X1    g20615(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n20808_));
  INV_X1     g20616(.I(new_n20808_), .ZN(new_n20809_));
  NOR2_X1    g20617(.A1(new_n20809_), .A2(\a[12] ), .ZN(new_n20810_));
  INV_X1     g20618(.I(new_n20810_), .ZN(new_n20811_));
  OAI21_X1   g20619(.A1(new_n20806_), .A2(new_n20807_), .B(new_n20811_), .ZN(new_n20812_));
  NAND2_X1   g20620(.A1(new_n20799_), .A2(new_n20811_), .ZN(new_n20813_));
  NOR4_X1    g20621(.A1(new_n20219_), .A2(new_n20236_), .A3(new_n20203_), .A4(new_n20813_), .ZN(new_n20814_));
  OAI21_X1   g20622(.A1(new_n20806_), .A2(new_n20807_), .B(new_n20814_), .ZN(new_n20815_));
  NOR3_X1    g20623(.A1(new_n20780_), .A2(\asqrt[61] ), .A3(new_n20752_), .ZN(new_n20816_));
  OAI21_X1   g20624(.A1(new_n20767_), .A2(new_n20816_), .B(new_n20781_), .ZN(new_n20817_));
  INV_X1     g20625(.I(new_n20767_), .ZN(new_n20818_));
  INV_X1     g20626(.I(new_n20735_), .ZN(new_n20819_));
  INV_X1     g20627(.I(new_n20703_), .ZN(new_n20820_));
  INV_X1     g20628(.I(new_n20676_), .ZN(new_n20821_));
  INV_X1     g20629(.I(new_n20649_), .ZN(new_n20822_));
  INV_X1     g20630(.I(new_n20623_), .ZN(new_n20823_));
  INV_X1     g20631(.I(new_n20597_), .ZN(new_n20824_));
  INV_X1     g20632(.I(new_n20568_), .ZN(new_n20825_));
  NOR3_X1    g20633(.A1(new_n20567_), .A2(new_n20552_), .A3(\asqrt[41] ), .ZN(new_n20826_));
  NOR2_X1    g20634(.A1(new_n20826_), .A2(new_n20573_), .ZN(new_n20827_));
  OAI21_X1   g20635(.A1(new_n20827_), .A2(new_n20825_), .B(\asqrt[42] ), .ZN(new_n20828_));
  NAND2_X1   g20636(.A1(new_n20828_), .A2(new_n3218_), .ZN(new_n20829_));
  OAI21_X1   g20637(.A1(new_n20829_), .A2(new_n20591_), .B(new_n20824_), .ZN(new_n20830_));
  NAND3_X1   g20638(.A1(new_n20830_), .A2(new_n2954_), .A3(new_n20592_), .ZN(new_n20831_));
  AOI22_X1   g20639(.A1(new_n20831_), .A2(new_n20606_), .B1(\asqrt[44] ), .B2(new_n20615_), .ZN(new_n20832_));
  OAI21_X1   g20640(.A1(new_n20832_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n20833_));
  OAI21_X1   g20641(.A1(new_n20833_), .A2(new_n20617_), .B(new_n20823_), .ZN(new_n20834_));
  NAND3_X1   g20642(.A1(new_n20834_), .A2(new_n2229_), .A3(new_n20618_), .ZN(new_n20835_));
  AOI22_X1   g20643(.A1(new_n20835_), .A2(new_n20632_), .B1(\asqrt[47] ), .B2(new_n20641_), .ZN(new_n20836_));
  OAI21_X1   g20644(.A1(new_n20836_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n20837_));
  OAI21_X1   g20645(.A1(new_n20837_), .A2(new_n20643_), .B(new_n20822_), .ZN(new_n20838_));
  NAND3_X1   g20646(.A1(new_n20838_), .A2(new_n1612_), .A3(new_n20644_), .ZN(new_n20839_));
  AOI22_X1   g20647(.A1(new_n20839_), .A2(new_n20658_), .B1(\asqrt[50] ), .B2(new_n20667_), .ZN(new_n20840_));
  OAI21_X1   g20648(.A1(new_n20840_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n20841_));
  OAI21_X1   g20649(.A1(new_n20841_), .A2(new_n20669_), .B(new_n20821_), .ZN(new_n20842_));
  NAND3_X1   g20650(.A1(new_n20842_), .A2(new_n1103_), .A3(new_n20670_), .ZN(new_n20843_));
  AOI22_X1   g20651(.A1(new_n20843_), .A2(new_n20685_), .B1(\asqrt[53] ), .B2(new_n20714_), .ZN(new_n20844_));
  OAI21_X1   g20652(.A1(new_n20844_), .A2(new_n904_), .B(new_n823_), .ZN(new_n20845_));
  OAI21_X1   g20653(.A1(new_n20845_), .A2(new_n20716_), .B(new_n20820_), .ZN(new_n20846_));
  NAND3_X1   g20654(.A1(new_n20846_), .A2(new_n703_), .A3(new_n20717_), .ZN(new_n20847_));
  AOI22_X1   g20655(.A1(new_n20847_), .A2(new_n20712_), .B1(\asqrt[56] ), .B2(new_n20746_), .ZN(new_n20848_));
  OAI21_X1   g20656(.A1(new_n20848_), .A2(new_n531_), .B(new_n436_), .ZN(new_n20849_));
  OAI21_X1   g20657(.A1(new_n20849_), .A2(new_n20748_), .B(new_n20819_), .ZN(new_n20850_));
  NAND3_X1   g20658(.A1(new_n20850_), .A2(new_n327_), .A3(new_n20749_), .ZN(new_n20851_));
  AOI22_X1   g20659(.A1(new_n20851_), .A2(new_n20744_), .B1(new_n20778_), .B2(\asqrt[59] ), .ZN(new_n20852_));
  OAI21_X1   g20660(.A1(new_n20852_), .A2(new_n306_), .B(new_n218_), .ZN(new_n20853_));
  OAI21_X1   g20661(.A1(new_n20853_), .A2(new_n20780_), .B(new_n20818_), .ZN(new_n20854_));
  NAND3_X1   g20662(.A1(new_n20854_), .A2(new_n207_), .A3(new_n20781_), .ZN(new_n20855_));
  AOI22_X1   g20663(.A1(new_n20855_), .A2(new_n20776_), .B1(new_n20817_), .B2(\asqrt[62] ), .ZN(new_n20856_));
  OAI21_X1   g20664(.A1(new_n20856_), .A2(new_n20791_), .B(new_n193_), .ZN(new_n20857_));
  AOI21_X1   g20665(.A1(new_n20817_), .A2(\asqrt[62] ), .B(new_n20788_), .ZN(new_n20858_));
  AOI21_X1   g20666(.A1(new_n20858_), .A2(new_n20783_), .B(new_n20803_), .ZN(new_n20859_));
  AOI21_X1   g20667(.A1(new_n20857_), .A2(new_n20859_), .B(new_n20212_), .ZN(new_n20860_));
  OAI21_X1   g20668(.A1(new_n20793_), .A2(new_n20805_), .B(new_n20807_), .ZN(new_n20861_));
  AOI21_X1   g20669(.A1(\a[13] ), .A2(new_n20861_), .B(new_n20860_), .ZN(new_n20862_));
  AOI22_X1   g20670(.A1(new_n20862_), .A2(new_n20815_), .B1(\asqrt[7] ), .B2(new_n20812_), .ZN(new_n20863_));
  NOR2_X1    g20671(.A1(new_n20863_), .A2(new_n19573_), .ZN(new_n20864_));
  NAND2_X1   g20672(.A1(new_n20862_), .A2(new_n20815_), .ZN(new_n20865_));
  OAI21_X1   g20673(.A1(new_n20793_), .A2(new_n20805_), .B(new_n20211_), .ZN(new_n20866_));
  NAND2_X1   g20674(.A1(new_n20858_), .A2(new_n20783_), .ZN(new_n20867_));
  OAI21_X1   g20675(.A1(new_n20801_), .A2(new_n20209_), .B(new_n20030_), .ZN(new_n20868_));
  NAND4_X1   g20676(.A1(new_n20857_), .A2(new_n20867_), .A3(new_n20798_), .A4(new_n20868_), .ZN(new_n20869_));
  AOI21_X1   g20677(.A1(new_n20869_), .A2(new_n20866_), .B(new_n20224_), .ZN(new_n20870_));
  INV_X1     g20678(.I(new_n20867_), .ZN(new_n20871_));
  NAND2_X1   g20679(.A1(new_n20798_), .A2(new_n20868_), .ZN(new_n20872_));
  NOR3_X1    g20680(.A1(new_n20871_), .A2(new_n20793_), .A3(new_n20872_), .ZN(new_n20873_));
  NOR3_X1    g20681(.A1(new_n20873_), .A2(new_n20860_), .A3(\a[14] ), .ZN(new_n20874_));
  NOR2_X1    g20682(.A1(new_n20870_), .A2(new_n20874_), .ZN(new_n20875_));
  AOI21_X1   g20683(.A1(new_n20812_), .A2(\asqrt[7] ), .B(\asqrt[8] ), .ZN(new_n20876_));
  AOI21_X1   g20684(.A1(new_n20865_), .A2(new_n20876_), .B(new_n20875_), .ZN(new_n20877_));
  OAI21_X1   g20685(.A1(new_n20877_), .A2(new_n20864_), .B(\asqrt[9] ), .ZN(new_n20878_));
  OAI21_X1   g20686(.A1(\asqrt[63] ), .A2(new_n20792_), .B(new_n20859_), .ZN(\asqrt[6] ));
  NOR3_X1    g20687(.A1(new_n20306_), .A2(new_n20223_), .A3(new_n20229_), .ZN(new_n20880_));
  NAND3_X1   g20688(.A1(\asqrt[6] ), .A2(new_n20244_), .A3(new_n20291_), .ZN(new_n20881_));
  AOI22_X1   g20689(.A1(new_n20881_), .A2(new_n20306_), .B1(\asqrt[6] ), .B2(new_n20880_), .ZN(new_n20882_));
  INV_X1     g20690(.I(new_n20882_), .ZN(new_n20883_));
  OAI21_X1   g20691(.A1(new_n20863_), .A2(new_n19573_), .B(new_n18792_), .ZN(new_n20884_));
  OAI21_X1   g20692(.A1(new_n20884_), .A2(new_n20877_), .B(new_n20883_), .ZN(new_n20885_));
  AOI21_X1   g20693(.A1(new_n20885_), .A2(new_n20878_), .B(new_n18275_), .ZN(new_n20886_));
  NOR2_X1    g20694(.A1(new_n20242_), .A2(new_n20243_), .ZN(new_n20887_));
  NOR2_X1    g20695(.A1(new_n20233_), .A2(new_n20245_), .ZN(new_n20888_));
  INV_X1     g20696(.I(new_n20888_), .ZN(new_n20889_));
  NAND4_X1   g20697(.A1(\asqrt[6] ), .A2(new_n20234_), .A3(new_n20887_), .A4(new_n20889_), .ZN(new_n20890_));
  NOR3_X1    g20698(.A1(new_n20806_), .A2(new_n20295_), .A3(new_n20888_), .ZN(new_n20891_));
  OAI21_X1   g20699(.A1(new_n20891_), .A2(new_n20887_), .B(new_n20890_), .ZN(new_n20892_));
  INV_X1     g20700(.I(new_n20892_), .ZN(new_n20893_));
  AOI21_X1   g20701(.A1(new_n20857_), .A2(new_n20859_), .B(new_n20807_), .ZN(new_n20894_));
  OAI21_X1   g20702(.A1(new_n20894_), .A2(new_n20810_), .B(\asqrt[7] ), .ZN(new_n20895_));
  INV_X1     g20703(.I(new_n20895_), .ZN(new_n20896_));
  INV_X1     g20704(.I(new_n20814_), .ZN(new_n20897_));
  NOR2_X1    g20705(.A1(new_n20894_), .A2(new_n20897_), .ZN(new_n20898_));
  INV_X1     g20706(.I(\a[13] ), .ZN(new_n20899_));
  AOI21_X1   g20707(.A1(\asqrt[6] ), .A2(new_n20807_), .B(new_n20899_), .ZN(new_n20900_));
  NOR3_X1    g20708(.A1(new_n20898_), .A2(new_n20900_), .A3(new_n20860_), .ZN(new_n20901_));
  OAI21_X1   g20709(.A1(new_n20901_), .A2(new_n20896_), .B(\asqrt[8] ), .ZN(new_n20902_));
  AOI21_X1   g20710(.A1(\asqrt[6] ), .A2(\a[12] ), .B(new_n20810_), .ZN(new_n20903_));
  OAI21_X1   g20711(.A1(new_n20903_), .A2(new_n20262_), .B(new_n19573_), .ZN(new_n20904_));
  OAI22_X1   g20712(.A1(new_n20901_), .A2(new_n20904_), .B1(new_n20870_), .B2(new_n20874_), .ZN(new_n20905_));
  AOI21_X1   g20713(.A1(new_n20905_), .A2(new_n20902_), .B(new_n18792_), .ZN(new_n20906_));
  AOI21_X1   g20714(.A1(new_n20857_), .A2(new_n20859_), .B(\a[12] ), .ZN(new_n20907_));
  OAI21_X1   g20715(.A1(new_n20899_), .A2(new_n20907_), .B(new_n20866_), .ZN(new_n20908_));
  OAI21_X1   g20716(.A1(new_n20908_), .A2(new_n20898_), .B(new_n20895_), .ZN(new_n20909_));
  AOI21_X1   g20717(.A1(new_n20909_), .A2(\asqrt[8] ), .B(\asqrt[9] ), .ZN(new_n20910_));
  AOI21_X1   g20718(.A1(new_n20910_), .A2(new_n20905_), .B(new_n20882_), .ZN(new_n20911_));
  NOR3_X1    g20719(.A1(new_n20911_), .A2(new_n20906_), .A3(\asqrt[10] ), .ZN(new_n20912_));
  NOR2_X1    g20720(.A1(new_n20912_), .A2(new_n20893_), .ZN(new_n20913_));
  OAI21_X1   g20721(.A1(new_n20913_), .A2(new_n20886_), .B(\asqrt[11] ), .ZN(new_n20914_));
  NOR2_X1    g20722(.A1(new_n20308_), .A2(new_n20300_), .ZN(new_n20915_));
  NOR3_X1    g20723(.A1(new_n20806_), .A2(new_n20247_), .A3(new_n20915_), .ZN(new_n20916_));
  INV_X1     g20724(.I(new_n20916_), .ZN(new_n20917_));
  NOR3_X1    g20725(.A1(new_n20915_), .A2(new_n20247_), .A3(new_n20305_), .ZN(new_n20918_));
  AOI22_X1   g20726(.A1(new_n20917_), .A2(new_n20305_), .B1(\asqrt[6] ), .B2(new_n20918_), .ZN(new_n20919_));
  INV_X1     g20727(.I(new_n20919_), .ZN(new_n20920_));
  OAI21_X1   g20728(.A1(new_n20911_), .A2(new_n20906_), .B(\asqrt[10] ), .ZN(new_n20921_));
  NAND2_X1   g20729(.A1(new_n20921_), .A2(new_n17623_), .ZN(new_n20922_));
  OAI21_X1   g20730(.A1(new_n20913_), .A2(new_n20922_), .B(new_n20920_), .ZN(new_n20923_));
  AOI21_X1   g20731(.A1(new_n20923_), .A2(new_n20914_), .B(new_n16881_), .ZN(new_n20924_));
  NOR3_X1    g20732(.A1(new_n20257_), .A2(new_n20266_), .A3(new_n20264_), .ZN(new_n20925_));
  NOR3_X1    g20733(.A1(new_n20806_), .A2(new_n20257_), .A3(new_n20266_), .ZN(new_n20926_));
  INV_X1     g20734(.I(new_n20926_), .ZN(new_n20927_));
  AOI22_X1   g20735(.A1(new_n20927_), .A2(new_n20264_), .B1(\asqrt[6] ), .B2(new_n20925_), .ZN(new_n20928_));
  OAI21_X1   g20736(.A1(new_n20893_), .A2(new_n20912_), .B(new_n20921_), .ZN(new_n20929_));
  AOI21_X1   g20737(.A1(new_n20929_), .A2(\asqrt[11] ), .B(\asqrt[12] ), .ZN(new_n20930_));
  AOI21_X1   g20738(.A1(new_n20930_), .A2(new_n20923_), .B(new_n20928_), .ZN(new_n20931_));
  OAI21_X1   g20739(.A1(new_n20931_), .A2(new_n20924_), .B(\asqrt[13] ), .ZN(new_n20932_));
  INV_X1     g20740(.I(new_n20932_), .ZN(new_n20933_));
  NAND2_X1   g20741(.A1(new_n20311_), .A2(new_n20303_), .ZN(new_n20934_));
  NAND3_X1   g20742(.A1(\asqrt[6] ), .A2(new_n20268_), .A3(new_n20934_), .ZN(new_n20935_));
  AND3_X2    g20743(.A1(new_n20268_), .A2(new_n20273_), .A3(new_n20934_), .Z(new_n20936_));
  AOI22_X1   g20744(.A1(new_n20935_), .A2(new_n20274_), .B1(\asqrt[6] ), .B2(new_n20936_), .ZN(new_n20937_));
  NOR3_X1    g20745(.A1(new_n20931_), .A2(new_n20924_), .A3(\asqrt[13] ), .ZN(new_n20938_));
  NOR2_X1    g20746(.A1(new_n20938_), .A2(new_n20937_), .ZN(new_n20939_));
  OAI21_X1   g20747(.A1(new_n20939_), .A2(new_n20933_), .B(\asqrt[14] ), .ZN(new_n20940_));
  INV_X1     g20748(.I(new_n20281_), .ZN(new_n20941_));
  NOR3_X1    g20749(.A1(new_n20277_), .A2(new_n20322_), .A3(new_n20941_), .ZN(new_n20942_));
  NOR3_X1    g20750(.A1(new_n20806_), .A2(new_n20277_), .A3(new_n20322_), .ZN(new_n20943_));
  INV_X1     g20751(.I(new_n20943_), .ZN(new_n20944_));
  AOI22_X1   g20752(.A1(new_n20944_), .A2(new_n20941_), .B1(\asqrt[6] ), .B2(new_n20942_), .ZN(new_n20945_));
  INV_X1     g20753(.I(new_n20945_), .ZN(new_n20946_));
  NAND2_X1   g20754(.A1(new_n20932_), .A2(new_n15770_), .ZN(new_n20947_));
  OAI21_X1   g20755(.A1(new_n20939_), .A2(new_n20947_), .B(new_n20946_), .ZN(new_n20948_));
  AOI21_X1   g20756(.A1(new_n20948_), .A2(new_n20940_), .B(new_n15067_), .ZN(new_n20949_));
  INV_X1     g20757(.I(new_n20347_), .ZN(new_n20950_));
  NAND3_X1   g20758(.A1(\asqrt[6] ), .A2(new_n20285_), .A3(new_n20950_), .ZN(new_n20951_));
  AND3_X2    g20759(.A1(new_n20950_), .A2(new_n20285_), .A3(new_n20289_), .Z(new_n20952_));
  AOI22_X1   g20760(.A1(new_n20951_), .A2(new_n20290_), .B1(\asqrt[6] ), .B2(new_n20952_), .ZN(new_n20953_));
  OAI21_X1   g20761(.A1(new_n20937_), .A2(new_n20938_), .B(new_n20932_), .ZN(new_n20954_));
  AOI21_X1   g20762(.A1(new_n20954_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n20955_));
  AOI21_X1   g20763(.A1(new_n20955_), .A2(new_n20948_), .B(new_n20953_), .ZN(new_n20956_));
  OAI21_X1   g20764(.A1(new_n20956_), .A2(new_n20949_), .B(\asqrt[16] ), .ZN(new_n20957_));
  INV_X1     g20765(.I(new_n20957_), .ZN(new_n20958_));
  INV_X1     g20766(.I(new_n20350_), .ZN(new_n20959_));
  NOR3_X1    g20767(.A1(new_n20959_), .A2(new_n20316_), .A3(new_n20349_), .ZN(new_n20960_));
  NOR3_X1    g20768(.A1(new_n20806_), .A2(new_n20316_), .A3(new_n20959_), .ZN(new_n20961_));
  INV_X1     g20769(.I(new_n20961_), .ZN(new_n20962_));
  AOI22_X1   g20770(.A1(new_n20962_), .A2(new_n20349_), .B1(\asqrt[6] ), .B2(new_n20960_), .ZN(new_n20963_));
  NOR3_X1    g20771(.A1(new_n20956_), .A2(new_n20949_), .A3(\asqrt[16] ), .ZN(new_n20964_));
  NOR2_X1    g20772(.A1(new_n20964_), .A2(new_n20963_), .ZN(new_n20965_));
  OAI21_X1   g20773(.A1(new_n20965_), .A2(new_n20958_), .B(\asqrt[17] ), .ZN(new_n20966_));
  INV_X1     g20774(.I(new_n20331_), .ZN(new_n20967_));
  NOR3_X1    g20775(.A1(new_n20806_), .A2(new_n20327_), .A3(new_n20332_), .ZN(new_n20968_));
  INV_X1     g20776(.I(new_n20968_), .ZN(new_n20969_));
  NOR3_X1    g20777(.A1(new_n20327_), .A2(new_n20967_), .A3(new_n20332_), .ZN(new_n20970_));
  AOI22_X1   g20778(.A1(new_n20969_), .A2(new_n20967_), .B1(\asqrt[6] ), .B2(new_n20970_), .ZN(new_n20971_));
  INV_X1     g20779(.I(new_n20971_), .ZN(new_n20972_));
  NAND2_X1   g20780(.A1(new_n20957_), .A2(new_n14017_), .ZN(new_n20973_));
  OAI21_X1   g20781(.A1(new_n20965_), .A2(new_n20973_), .B(new_n20972_), .ZN(new_n20974_));
  AOI21_X1   g20782(.A1(new_n20974_), .A2(new_n20966_), .B(new_n13353_), .ZN(new_n20975_));
  OAI21_X1   g20783(.A1(new_n20333_), .A2(new_n20339_), .B(new_n20337_), .ZN(new_n20976_));
  AOI21_X1   g20784(.A1(\asqrt[17] ), .A2(new_n20352_), .B(new_n20976_), .ZN(new_n20977_));
  OAI21_X1   g20785(.A1(new_n20333_), .A2(new_n20339_), .B(new_n20334_), .ZN(new_n20978_));
  NOR2_X1    g20786(.A1(new_n20806_), .A2(new_n20978_), .ZN(new_n20979_));
  INV_X1     g20787(.I(new_n20979_), .ZN(new_n20980_));
  AOI22_X1   g20788(.A1(new_n20980_), .A2(new_n20338_), .B1(\asqrt[6] ), .B2(new_n20977_), .ZN(new_n20981_));
  OAI21_X1   g20789(.A1(new_n20963_), .A2(new_n20964_), .B(new_n20957_), .ZN(new_n20982_));
  AOI21_X1   g20790(.A1(new_n20982_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n20983_));
  AOI21_X1   g20791(.A1(new_n20983_), .A2(new_n20974_), .B(new_n20981_), .ZN(new_n20984_));
  OAI21_X1   g20792(.A1(new_n20984_), .A2(new_n20975_), .B(\asqrt[19] ), .ZN(new_n20985_));
  INV_X1     g20793(.I(new_n20985_), .ZN(new_n20986_));
  INV_X1     g20794(.I(new_n20346_), .ZN(new_n20987_));
  INV_X1     g20795(.I(new_n20340_), .ZN(new_n20988_));
  INV_X1     g20796(.I(new_n20353_), .ZN(new_n20989_));
  NOR2_X1    g20797(.A1(new_n20989_), .A2(new_n20988_), .ZN(new_n20990_));
  NOR3_X1    g20798(.A1(new_n20806_), .A2(new_n20341_), .A3(new_n20990_), .ZN(new_n20991_));
  INV_X1     g20799(.I(new_n20991_), .ZN(new_n20992_));
  NOR3_X1    g20800(.A1(new_n20990_), .A2(new_n20341_), .A3(new_n20987_), .ZN(new_n20993_));
  AOI22_X1   g20801(.A1(new_n20992_), .A2(new_n20987_), .B1(\asqrt[6] ), .B2(new_n20993_), .ZN(new_n20994_));
  NOR3_X1    g20802(.A1(new_n20984_), .A2(new_n20975_), .A3(\asqrt[19] ), .ZN(new_n20995_));
  NOR2_X1    g20803(.A1(new_n20995_), .A2(new_n20994_), .ZN(new_n20996_));
  OAI21_X1   g20804(.A1(new_n20996_), .A2(new_n20986_), .B(\asqrt[20] ), .ZN(new_n20997_));
  INV_X1     g20805(.I(new_n20360_), .ZN(new_n20998_));
  NOR3_X1    g20806(.A1(new_n20356_), .A2(new_n20998_), .A3(new_n20361_), .ZN(new_n20999_));
  NOR3_X1    g20807(.A1(new_n20806_), .A2(new_n20356_), .A3(new_n20361_), .ZN(new_n21000_));
  INV_X1     g20808(.I(new_n21000_), .ZN(new_n21001_));
  AOI22_X1   g20809(.A1(new_n21001_), .A2(new_n20998_), .B1(\asqrt[6] ), .B2(new_n20999_), .ZN(new_n21002_));
  INV_X1     g20810(.I(new_n21002_), .ZN(new_n21003_));
  NAND2_X1   g20811(.A1(new_n20985_), .A2(new_n12364_), .ZN(new_n21004_));
  OAI21_X1   g20812(.A1(new_n20996_), .A2(new_n21004_), .B(new_n21003_), .ZN(new_n21005_));
  AOI21_X1   g20813(.A1(new_n21005_), .A2(new_n20997_), .B(new_n11736_), .ZN(new_n21006_));
  NOR2_X1    g20814(.A1(new_n20362_), .A2(new_n20370_), .ZN(new_n21007_));
  INV_X1     g20815(.I(new_n21007_), .ZN(new_n21008_));
  NAND3_X1   g20816(.A1(\asqrt[6] ), .A2(new_n20363_), .A3(new_n21008_), .ZN(new_n21009_));
  AND3_X2    g20817(.A1(new_n21008_), .A2(new_n20363_), .A3(new_n20368_), .Z(new_n21010_));
  AOI22_X1   g20818(.A1(new_n21009_), .A2(new_n20369_), .B1(\asqrt[6] ), .B2(new_n21010_), .ZN(new_n21011_));
  OAI21_X1   g20819(.A1(new_n20994_), .A2(new_n20995_), .B(new_n20985_), .ZN(new_n21012_));
  AOI21_X1   g20820(.A1(new_n21012_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n21013_));
  AOI21_X1   g20821(.A1(new_n21013_), .A2(new_n21005_), .B(new_n21011_), .ZN(new_n21014_));
  OAI21_X1   g20822(.A1(new_n21014_), .A2(new_n21006_), .B(\asqrt[22] ), .ZN(new_n21015_));
  INV_X1     g20823(.I(new_n21015_), .ZN(new_n21016_));
  INV_X1     g20824(.I(new_n20377_), .ZN(new_n21017_));
  INV_X1     g20825(.I(new_n20371_), .ZN(new_n21018_));
  INV_X1     g20826(.I(new_n20379_), .ZN(new_n21019_));
  NOR2_X1    g20827(.A1(new_n21019_), .A2(new_n21018_), .ZN(new_n21020_));
  NOR3_X1    g20828(.A1(new_n21020_), .A2(new_n20372_), .A3(new_n21017_), .ZN(new_n21021_));
  NOR3_X1    g20829(.A1(new_n20806_), .A2(new_n20372_), .A3(new_n21020_), .ZN(new_n21022_));
  INV_X1     g20830(.I(new_n21022_), .ZN(new_n21023_));
  AOI22_X1   g20831(.A1(new_n21023_), .A2(new_n21017_), .B1(\asqrt[6] ), .B2(new_n21021_), .ZN(new_n21024_));
  NOR3_X1    g20832(.A1(new_n21014_), .A2(new_n21006_), .A3(\asqrt[22] ), .ZN(new_n21025_));
  NOR2_X1    g20833(.A1(new_n21025_), .A2(new_n21024_), .ZN(new_n21026_));
  OAI21_X1   g20834(.A1(new_n21026_), .A2(new_n21016_), .B(\asqrt[23] ), .ZN(new_n21027_));
  INV_X1     g20835(.I(new_n20386_), .ZN(new_n21028_));
  NOR3_X1    g20836(.A1(new_n20806_), .A2(new_n20382_), .A3(new_n20387_), .ZN(new_n21029_));
  INV_X1     g20837(.I(new_n21029_), .ZN(new_n21030_));
  NOR3_X1    g20838(.A1(new_n20382_), .A2(new_n21028_), .A3(new_n20387_), .ZN(new_n21031_));
  AOI22_X1   g20839(.A1(new_n21030_), .A2(new_n21028_), .B1(\asqrt[6] ), .B2(new_n21031_), .ZN(new_n21032_));
  INV_X1     g20840(.I(new_n21032_), .ZN(new_n21033_));
  NAND2_X1   g20841(.A1(new_n21015_), .A2(new_n10812_), .ZN(new_n21034_));
  OAI21_X1   g20842(.A1(new_n21026_), .A2(new_n21034_), .B(new_n21033_), .ZN(new_n21035_));
  AOI21_X1   g20843(.A1(new_n21035_), .A2(new_n21027_), .B(new_n10221_), .ZN(new_n21036_));
  NOR2_X1    g20844(.A1(new_n20388_), .A2(new_n20396_), .ZN(new_n21037_));
  INV_X1     g20845(.I(new_n21037_), .ZN(new_n21038_));
  AND3_X2    g20846(.A1(new_n21038_), .A2(new_n20389_), .A3(new_n20394_), .Z(new_n21039_));
  NAND3_X1   g20847(.A1(\asqrt[6] ), .A2(new_n20389_), .A3(new_n21038_), .ZN(new_n21040_));
  AOI22_X1   g20848(.A1(new_n21040_), .A2(new_n20395_), .B1(\asqrt[6] ), .B2(new_n21039_), .ZN(new_n21041_));
  OAI21_X1   g20849(.A1(new_n21024_), .A2(new_n21025_), .B(new_n21015_), .ZN(new_n21042_));
  AOI21_X1   g20850(.A1(new_n21042_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n21043_));
  AOI21_X1   g20851(.A1(new_n21043_), .A2(new_n21035_), .B(new_n21041_), .ZN(new_n21044_));
  OAI21_X1   g20852(.A1(new_n21044_), .A2(new_n21036_), .B(\asqrt[25] ), .ZN(new_n21045_));
  INV_X1     g20853(.I(new_n21045_), .ZN(new_n21046_));
  INV_X1     g20854(.I(new_n20403_), .ZN(new_n21047_));
  INV_X1     g20855(.I(new_n20397_), .ZN(new_n21048_));
  INV_X1     g20856(.I(new_n20405_), .ZN(new_n21049_));
  NOR2_X1    g20857(.A1(new_n21049_), .A2(new_n21048_), .ZN(new_n21050_));
  NOR3_X1    g20858(.A1(new_n20806_), .A2(new_n20398_), .A3(new_n21050_), .ZN(new_n21051_));
  INV_X1     g20859(.I(new_n21051_), .ZN(new_n21052_));
  NOR3_X1    g20860(.A1(new_n21050_), .A2(new_n20398_), .A3(new_n21047_), .ZN(new_n21053_));
  AOI22_X1   g20861(.A1(new_n21052_), .A2(new_n21047_), .B1(\asqrt[6] ), .B2(new_n21053_), .ZN(new_n21054_));
  NOR3_X1    g20862(.A1(new_n21044_), .A2(new_n21036_), .A3(\asqrt[25] ), .ZN(new_n21055_));
  NOR2_X1    g20863(.A1(new_n21055_), .A2(new_n21054_), .ZN(new_n21056_));
  OAI21_X1   g20864(.A1(new_n21056_), .A2(new_n21046_), .B(\asqrt[26] ), .ZN(new_n21057_));
  INV_X1     g20865(.I(new_n20412_), .ZN(new_n21058_));
  NOR3_X1    g20866(.A1(new_n20408_), .A2(new_n21058_), .A3(new_n20413_), .ZN(new_n21059_));
  NOR3_X1    g20867(.A1(new_n20806_), .A2(new_n20408_), .A3(new_n20413_), .ZN(new_n21060_));
  INV_X1     g20868(.I(new_n21060_), .ZN(new_n21061_));
  AOI22_X1   g20869(.A1(new_n21061_), .A2(new_n21058_), .B1(\asqrt[6] ), .B2(new_n21059_), .ZN(new_n21062_));
  INV_X1     g20870(.I(new_n21062_), .ZN(new_n21063_));
  NAND2_X1   g20871(.A1(new_n21045_), .A2(new_n9317_), .ZN(new_n21064_));
  OAI21_X1   g20872(.A1(new_n21056_), .A2(new_n21064_), .B(new_n21063_), .ZN(new_n21065_));
  AOI21_X1   g20873(.A1(new_n21065_), .A2(new_n21057_), .B(new_n8826_), .ZN(new_n21066_));
  NOR2_X1    g20874(.A1(new_n20414_), .A2(new_n20422_), .ZN(new_n21067_));
  INV_X1     g20875(.I(new_n21067_), .ZN(new_n21068_));
  NAND3_X1   g20876(.A1(\asqrt[6] ), .A2(new_n20415_), .A3(new_n21068_), .ZN(new_n21069_));
  AND3_X2    g20877(.A1(new_n21068_), .A2(new_n20415_), .A3(new_n20420_), .Z(new_n21070_));
  AOI22_X1   g20878(.A1(new_n21069_), .A2(new_n20421_), .B1(\asqrt[6] ), .B2(new_n21070_), .ZN(new_n21071_));
  OAI21_X1   g20879(.A1(new_n21054_), .A2(new_n21055_), .B(new_n21045_), .ZN(new_n21072_));
  AOI21_X1   g20880(.A1(new_n21072_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n21073_));
  AOI21_X1   g20881(.A1(new_n21073_), .A2(new_n21065_), .B(new_n21071_), .ZN(new_n21074_));
  OAI21_X1   g20882(.A1(new_n21074_), .A2(new_n21066_), .B(\asqrt[28] ), .ZN(new_n21075_));
  INV_X1     g20883(.I(new_n21075_), .ZN(new_n21076_));
  INV_X1     g20884(.I(new_n20429_), .ZN(new_n21077_));
  INV_X1     g20885(.I(new_n20423_), .ZN(new_n21078_));
  INV_X1     g20886(.I(new_n20431_), .ZN(new_n21079_));
  NOR2_X1    g20887(.A1(new_n21079_), .A2(new_n21078_), .ZN(new_n21080_));
  NOR3_X1    g20888(.A1(new_n21080_), .A2(new_n20424_), .A3(new_n21077_), .ZN(new_n21081_));
  NOR3_X1    g20889(.A1(new_n20806_), .A2(new_n20424_), .A3(new_n21080_), .ZN(new_n21082_));
  INV_X1     g20890(.I(new_n21082_), .ZN(new_n21083_));
  AOI22_X1   g20891(.A1(new_n21083_), .A2(new_n21077_), .B1(\asqrt[6] ), .B2(new_n21081_), .ZN(new_n21084_));
  NOR3_X1    g20892(.A1(new_n21074_), .A2(new_n21066_), .A3(\asqrt[28] ), .ZN(new_n21085_));
  NOR2_X1    g20893(.A1(new_n21085_), .A2(new_n21084_), .ZN(new_n21086_));
  OAI21_X1   g20894(.A1(new_n21086_), .A2(new_n21076_), .B(\asqrt[29] ), .ZN(new_n21087_));
  INV_X1     g20895(.I(new_n20439_), .ZN(new_n21088_));
  NOR3_X1    g20896(.A1(new_n20806_), .A2(new_n20434_), .A3(new_n20476_), .ZN(new_n21089_));
  INV_X1     g20897(.I(new_n21089_), .ZN(new_n21090_));
  NOR3_X1    g20898(.A1(new_n20434_), .A2(new_n21088_), .A3(new_n20476_), .ZN(new_n21091_));
  AOI22_X1   g20899(.A1(new_n21090_), .A2(new_n21088_), .B1(\asqrt[6] ), .B2(new_n21091_), .ZN(new_n21092_));
  INV_X1     g20900(.I(new_n21092_), .ZN(new_n21093_));
  NAND2_X1   g20901(.A1(new_n21075_), .A2(new_n8036_), .ZN(new_n21094_));
  OAI21_X1   g20902(.A1(new_n21086_), .A2(new_n21094_), .B(new_n21093_), .ZN(new_n21095_));
  AOI21_X1   g20903(.A1(new_n21095_), .A2(new_n21087_), .B(new_n7539_), .ZN(new_n21096_));
  NOR2_X1    g20904(.A1(new_n20449_), .A2(new_n20441_), .ZN(new_n21097_));
  INV_X1     g20905(.I(new_n21097_), .ZN(new_n21098_));
  AND3_X2    g20906(.A1(new_n21098_), .A2(new_n20442_), .A3(new_n20447_), .Z(new_n21099_));
  NAND3_X1   g20907(.A1(\asqrt[6] ), .A2(new_n20442_), .A3(new_n21098_), .ZN(new_n21100_));
  AOI22_X1   g20908(.A1(new_n21100_), .A2(new_n20448_), .B1(\asqrt[6] ), .B2(new_n21099_), .ZN(new_n21101_));
  OAI21_X1   g20909(.A1(new_n21084_), .A2(new_n21085_), .B(new_n21075_), .ZN(new_n21102_));
  AOI21_X1   g20910(.A1(new_n21102_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n21103_));
  AOI21_X1   g20911(.A1(new_n21103_), .A2(new_n21095_), .B(new_n21101_), .ZN(new_n21104_));
  OAI21_X1   g20912(.A1(new_n21104_), .A2(new_n21096_), .B(\asqrt[31] ), .ZN(new_n21105_));
  INV_X1     g20913(.I(new_n21105_), .ZN(new_n21106_));
  NOR2_X1    g20914(.A1(new_n20460_), .A2(new_n20453_), .ZN(new_n21107_));
  NOR3_X1    g20915(.A1(new_n20806_), .A2(new_n20451_), .A3(new_n21107_), .ZN(new_n21108_));
  INV_X1     g20916(.I(new_n21108_), .ZN(new_n21109_));
  NOR3_X1    g20917(.A1(new_n21107_), .A2(new_n20451_), .A3(new_n20459_), .ZN(new_n21110_));
  AOI22_X1   g20918(.A1(new_n21109_), .A2(new_n20459_), .B1(\asqrt[6] ), .B2(new_n21110_), .ZN(new_n21111_));
  NOR3_X1    g20919(.A1(new_n21104_), .A2(new_n21096_), .A3(\asqrt[31] ), .ZN(new_n21112_));
  NOR2_X1    g20920(.A1(new_n21112_), .A2(new_n21111_), .ZN(new_n21113_));
  OAI21_X1   g20921(.A1(new_n21113_), .A2(new_n21106_), .B(\asqrt[32] ), .ZN(new_n21114_));
  INV_X1     g20922(.I(new_n20466_), .ZN(new_n21115_));
  NOR3_X1    g20923(.A1(new_n20462_), .A2(new_n21115_), .A3(new_n20508_), .ZN(new_n21116_));
  NOR3_X1    g20924(.A1(new_n20806_), .A2(new_n20462_), .A3(new_n20508_), .ZN(new_n21117_));
  INV_X1     g20925(.I(new_n21117_), .ZN(new_n21118_));
  AOI22_X1   g20926(.A1(new_n21118_), .A2(new_n21115_), .B1(\asqrt[6] ), .B2(new_n21116_), .ZN(new_n21119_));
  INV_X1     g20927(.I(new_n21119_), .ZN(new_n21120_));
  NAND2_X1   g20928(.A1(new_n21105_), .A2(new_n6824_), .ZN(new_n21121_));
  OAI21_X1   g20929(.A1(new_n21113_), .A2(new_n21121_), .B(new_n21120_), .ZN(new_n21122_));
  AOI21_X1   g20930(.A1(new_n21122_), .A2(new_n21114_), .B(new_n6356_), .ZN(new_n21123_));
  NOR2_X1    g20931(.A1(new_n20481_), .A2(new_n20468_), .ZN(new_n21124_));
  INV_X1     g20932(.I(new_n21124_), .ZN(new_n21125_));
  NAND3_X1   g20933(.A1(\asqrt[6] ), .A2(new_n20469_), .A3(new_n21125_), .ZN(new_n21126_));
  AND3_X2    g20934(.A1(new_n21125_), .A2(new_n20469_), .A3(new_n20474_), .Z(new_n21127_));
  AOI22_X1   g20935(.A1(new_n21126_), .A2(new_n20475_), .B1(\asqrt[6] ), .B2(new_n21127_), .ZN(new_n21128_));
  OAI21_X1   g20936(.A1(new_n21111_), .A2(new_n21112_), .B(new_n21105_), .ZN(new_n21129_));
  AOI21_X1   g20937(.A1(new_n21129_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n21130_));
  AOI21_X1   g20938(.A1(new_n21130_), .A2(new_n21122_), .B(new_n21128_), .ZN(new_n21131_));
  OAI21_X1   g20939(.A1(new_n21131_), .A2(new_n21123_), .B(\asqrt[34] ), .ZN(new_n21132_));
  INV_X1     g20940(.I(new_n21132_), .ZN(new_n21133_));
  NOR2_X1    g20941(.A1(new_n20492_), .A2(new_n20485_), .ZN(new_n21134_));
  NOR3_X1    g20942(.A1(new_n21134_), .A2(new_n20483_), .A3(new_n20491_), .ZN(new_n21135_));
  NOR3_X1    g20943(.A1(new_n20806_), .A2(new_n20483_), .A3(new_n21134_), .ZN(new_n21136_));
  INV_X1     g20944(.I(new_n21136_), .ZN(new_n21137_));
  AOI22_X1   g20945(.A1(new_n21137_), .A2(new_n20491_), .B1(\asqrt[6] ), .B2(new_n21135_), .ZN(new_n21138_));
  NOR3_X1    g20946(.A1(new_n21131_), .A2(new_n21123_), .A3(\asqrt[34] ), .ZN(new_n21139_));
  NOR2_X1    g20947(.A1(new_n21139_), .A2(new_n21138_), .ZN(new_n21140_));
  OAI21_X1   g20948(.A1(new_n21140_), .A2(new_n21133_), .B(\asqrt[35] ), .ZN(new_n21141_));
  INV_X1     g20949(.I(new_n20498_), .ZN(new_n21142_));
  NOR3_X1    g20950(.A1(new_n20806_), .A2(new_n20494_), .A3(new_n20558_), .ZN(new_n21143_));
  INV_X1     g20951(.I(new_n21143_), .ZN(new_n21144_));
  NOR3_X1    g20952(.A1(new_n20494_), .A2(new_n21142_), .A3(new_n20558_), .ZN(new_n21145_));
  AOI22_X1   g20953(.A1(new_n21144_), .A2(new_n21142_), .B1(\asqrt[6] ), .B2(new_n21145_), .ZN(new_n21146_));
  INV_X1     g20954(.I(new_n21146_), .ZN(new_n21147_));
  NAND2_X1   g20955(.A1(new_n21132_), .A2(new_n5708_), .ZN(new_n21148_));
  OAI21_X1   g20956(.A1(new_n21140_), .A2(new_n21148_), .B(new_n21147_), .ZN(new_n21149_));
  AOI21_X1   g20957(.A1(new_n21149_), .A2(new_n21141_), .B(new_n5277_), .ZN(new_n21150_));
  NOR2_X1    g20958(.A1(new_n20513_), .A2(new_n20500_), .ZN(new_n21151_));
  INV_X1     g20959(.I(new_n21151_), .ZN(new_n21152_));
  AND3_X2    g20960(.A1(new_n21152_), .A2(new_n20501_), .A3(new_n20506_), .Z(new_n21153_));
  NAND3_X1   g20961(.A1(\asqrt[6] ), .A2(new_n20501_), .A3(new_n21152_), .ZN(new_n21154_));
  AOI22_X1   g20962(.A1(new_n21154_), .A2(new_n20507_), .B1(\asqrt[6] ), .B2(new_n21153_), .ZN(new_n21155_));
  OAI21_X1   g20963(.A1(new_n21138_), .A2(new_n21139_), .B(new_n21132_), .ZN(new_n21156_));
  AOI21_X1   g20964(.A1(new_n21156_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n21157_));
  AOI21_X1   g20965(.A1(new_n21157_), .A2(new_n21149_), .B(new_n21155_), .ZN(new_n21158_));
  OAI21_X1   g20966(.A1(new_n21158_), .A2(new_n21150_), .B(\asqrt[37] ), .ZN(new_n21159_));
  INV_X1     g20967(.I(new_n21159_), .ZN(new_n21160_));
  NOR2_X1    g20968(.A1(new_n20517_), .A2(new_n20524_), .ZN(new_n21161_));
  NOR3_X1    g20969(.A1(new_n20806_), .A2(new_n20531_), .A3(new_n21161_), .ZN(new_n21162_));
  INV_X1     g20970(.I(new_n21162_), .ZN(new_n21163_));
  NOR3_X1    g20971(.A1(new_n21161_), .A2(new_n20531_), .A3(new_n20523_), .ZN(new_n21164_));
  AOI22_X1   g20972(.A1(new_n21163_), .A2(new_n20523_), .B1(\asqrt[6] ), .B2(new_n21164_), .ZN(new_n21165_));
  NOR3_X1    g20973(.A1(new_n21158_), .A2(new_n21150_), .A3(\asqrt[37] ), .ZN(new_n21166_));
  NOR2_X1    g20974(.A1(new_n21166_), .A2(new_n21165_), .ZN(new_n21167_));
  OAI21_X1   g20975(.A1(new_n21167_), .A2(new_n21160_), .B(\asqrt[38] ), .ZN(new_n21168_));
  INV_X1     g20976(.I(new_n20530_), .ZN(new_n21169_));
  NOR3_X1    g20977(.A1(new_n20526_), .A2(new_n21169_), .A3(new_n20575_), .ZN(new_n21170_));
  NOR3_X1    g20978(.A1(new_n20806_), .A2(new_n20526_), .A3(new_n20575_), .ZN(new_n21171_));
  INV_X1     g20979(.I(new_n21171_), .ZN(new_n21172_));
  AOI22_X1   g20980(.A1(new_n21172_), .A2(new_n21169_), .B1(\asqrt[6] ), .B2(new_n21170_), .ZN(new_n21173_));
  INV_X1     g20981(.I(new_n21173_), .ZN(new_n21174_));
  NAND2_X1   g20982(.A1(new_n21159_), .A2(new_n4696_), .ZN(new_n21175_));
  OAI21_X1   g20983(.A1(new_n21167_), .A2(new_n21175_), .B(new_n21174_), .ZN(new_n21176_));
  AOI21_X1   g20984(.A1(new_n21176_), .A2(new_n21168_), .B(new_n4298_), .ZN(new_n21177_));
  NOR3_X1    g20985(.A1(new_n20806_), .A2(new_n20535_), .A3(new_n20541_), .ZN(new_n21178_));
  INV_X1     g20986(.I(new_n21178_), .ZN(new_n21179_));
  NOR3_X1    g20987(.A1(new_n20535_), .A2(new_n20557_), .A3(new_n20541_), .ZN(new_n21180_));
  AOI22_X1   g20988(.A1(new_n21179_), .A2(new_n20557_), .B1(\asqrt[6] ), .B2(new_n21180_), .ZN(new_n21181_));
  OAI21_X1   g20989(.A1(new_n21165_), .A2(new_n21166_), .B(new_n21159_), .ZN(new_n21182_));
  AOI21_X1   g20990(.A1(new_n21182_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n21183_));
  AOI21_X1   g20991(.A1(new_n21183_), .A2(new_n21176_), .B(new_n21181_), .ZN(new_n21184_));
  OAI21_X1   g20992(.A1(new_n21184_), .A2(new_n21177_), .B(\asqrt[40] ), .ZN(new_n21185_));
  INV_X1     g20993(.I(new_n21185_), .ZN(new_n21186_));
  NOR2_X1    g20994(.A1(new_n20542_), .A2(new_n20550_), .ZN(new_n21187_));
  NOR3_X1    g20995(.A1(new_n21187_), .A2(new_n20565_), .A3(new_n20549_), .ZN(new_n21188_));
  NOR3_X1    g20996(.A1(new_n20806_), .A2(new_n20565_), .A3(new_n21187_), .ZN(new_n21189_));
  INV_X1     g20997(.I(new_n21189_), .ZN(new_n21190_));
  AOI22_X1   g20998(.A1(new_n21190_), .A2(new_n20549_), .B1(\asqrt[6] ), .B2(new_n21188_), .ZN(new_n21191_));
  NOR3_X1    g20999(.A1(new_n21184_), .A2(new_n21177_), .A3(\asqrt[40] ), .ZN(new_n21192_));
  NOR2_X1    g21000(.A1(new_n21192_), .A2(new_n21191_), .ZN(new_n21193_));
  OAI21_X1   g21001(.A1(new_n21193_), .A2(new_n21186_), .B(\asqrt[41] ), .ZN(new_n21194_));
  INV_X1     g21002(.I(new_n20556_), .ZN(new_n21195_));
  NOR3_X1    g21003(.A1(new_n20806_), .A2(new_n20552_), .A3(new_n20588_), .ZN(new_n21196_));
  INV_X1     g21004(.I(new_n21196_), .ZN(new_n21197_));
  NOR3_X1    g21005(.A1(new_n20552_), .A2(new_n21195_), .A3(new_n20588_), .ZN(new_n21198_));
  AOI22_X1   g21006(.A1(new_n21197_), .A2(new_n21195_), .B1(\asqrt[6] ), .B2(new_n21198_), .ZN(new_n21199_));
  INV_X1     g21007(.I(new_n21199_), .ZN(new_n21200_));
  NAND2_X1   g21008(.A1(new_n21185_), .A2(new_n3782_), .ZN(new_n21201_));
  OAI21_X1   g21009(.A1(new_n21193_), .A2(new_n21201_), .B(new_n21200_), .ZN(new_n21202_));
  AOI21_X1   g21010(.A1(new_n21202_), .A2(new_n21194_), .B(new_n3419_), .ZN(new_n21203_));
  NOR3_X1    g21011(.A1(new_n20825_), .A2(new_n20574_), .A3(new_n20826_), .ZN(new_n21204_));
  NOR3_X1    g21012(.A1(new_n20806_), .A2(new_n20825_), .A3(new_n20826_), .ZN(new_n21205_));
  INV_X1     g21013(.I(new_n21205_), .ZN(new_n21206_));
  AOI22_X1   g21014(.A1(new_n21206_), .A2(new_n20574_), .B1(\asqrt[6] ), .B2(new_n21204_), .ZN(new_n21207_));
  OAI21_X1   g21015(.A1(new_n21191_), .A2(new_n21192_), .B(new_n21185_), .ZN(new_n21208_));
  AOI21_X1   g21016(.A1(new_n21208_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n21209_));
  AOI21_X1   g21017(.A1(new_n21209_), .A2(new_n21202_), .B(new_n21207_), .ZN(new_n21210_));
  OAI21_X1   g21018(.A1(new_n21210_), .A2(new_n21203_), .B(\asqrt[43] ), .ZN(new_n21211_));
  INV_X1     g21019(.I(new_n21211_), .ZN(new_n21212_));
  INV_X1     g21020(.I(new_n20587_), .ZN(new_n21213_));
  NAND2_X1   g21021(.A1(new_n20568_), .A2(new_n3419_), .ZN(new_n21214_));
  NOR2_X1    g21022(.A1(new_n20827_), .A2(new_n21214_), .ZN(new_n21215_));
  NOR3_X1    g21023(.A1(new_n20806_), .A2(new_n20582_), .A3(new_n21215_), .ZN(new_n21216_));
  INV_X1     g21024(.I(new_n21216_), .ZN(new_n21217_));
  NOR3_X1    g21025(.A1(new_n21215_), .A2(new_n20582_), .A3(new_n21213_), .ZN(new_n21218_));
  AOI22_X1   g21026(.A1(new_n21217_), .A2(new_n21213_), .B1(\asqrt[6] ), .B2(new_n21218_), .ZN(new_n21219_));
  NOR3_X1    g21027(.A1(new_n21210_), .A2(new_n21203_), .A3(\asqrt[43] ), .ZN(new_n21220_));
  NOR2_X1    g21028(.A1(new_n21220_), .A2(new_n21219_), .ZN(new_n21221_));
  OAI21_X1   g21029(.A1(new_n21221_), .A2(new_n21212_), .B(\asqrt[44] ), .ZN(new_n21222_));
  NOR3_X1    g21030(.A1(new_n20593_), .A2(new_n20598_), .A3(new_n20824_), .ZN(new_n21223_));
  NOR3_X1    g21031(.A1(new_n20806_), .A2(new_n20593_), .A3(new_n20598_), .ZN(new_n21224_));
  INV_X1     g21032(.I(new_n21224_), .ZN(new_n21225_));
  AOI22_X1   g21033(.A1(new_n21225_), .A2(new_n20824_), .B1(\asqrt[6] ), .B2(new_n21223_), .ZN(new_n21226_));
  INV_X1     g21034(.I(new_n21226_), .ZN(new_n21227_));
  NAND2_X1   g21035(.A1(new_n21211_), .A2(new_n2954_), .ZN(new_n21228_));
  OAI21_X1   g21036(.A1(new_n21221_), .A2(new_n21228_), .B(new_n21227_), .ZN(new_n21229_));
  AOI21_X1   g21037(.A1(new_n21229_), .A2(new_n21222_), .B(new_n2641_), .ZN(new_n21230_));
  INV_X1     g21038(.I(new_n20600_), .ZN(new_n21231_));
  NOR2_X1    g21039(.A1(new_n20599_), .A2(new_n20607_), .ZN(new_n21232_));
  NOR3_X1    g21040(.A1(new_n20806_), .A2(new_n21231_), .A3(new_n21232_), .ZN(new_n21233_));
  INV_X1     g21041(.I(new_n21233_), .ZN(new_n21234_));
  NOR3_X1    g21042(.A1(new_n21231_), .A2(new_n21232_), .A3(new_n20606_), .ZN(new_n21235_));
  AOI22_X1   g21043(.A1(new_n21234_), .A2(new_n20606_), .B1(\asqrt[6] ), .B2(new_n21235_), .ZN(new_n21236_));
  OAI21_X1   g21044(.A1(new_n21219_), .A2(new_n21220_), .B(new_n21211_), .ZN(new_n21237_));
  AOI21_X1   g21045(.A1(new_n21237_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n21238_));
  AOI21_X1   g21046(.A1(new_n21238_), .A2(new_n21229_), .B(new_n21236_), .ZN(new_n21239_));
  OAI21_X1   g21047(.A1(new_n21239_), .A2(new_n21230_), .B(\asqrt[46] ), .ZN(new_n21240_));
  INV_X1     g21048(.I(new_n21240_), .ZN(new_n21241_));
  INV_X1     g21049(.I(new_n20614_), .ZN(new_n21242_));
  INV_X1     g21050(.I(new_n20608_), .ZN(new_n21243_));
  INV_X1     g21051(.I(new_n20616_), .ZN(new_n21244_));
  NOR2_X1    g21052(.A1(new_n21244_), .A2(new_n21243_), .ZN(new_n21245_));
  NOR3_X1    g21053(.A1(new_n21245_), .A2(new_n20609_), .A3(new_n21242_), .ZN(new_n21246_));
  NOR3_X1    g21054(.A1(new_n20806_), .A2(new_n20609_), .A3(new_n21245_), .ZN(new_n21247_));
  INV_X1     g21055(.I(new_n21247_), .ZN(new_n21248_));
  AOI22_X1   g21056(.A1(new_n21248_), .A2(new_n21242_), .B1(\asqrt[6] ), .B2(new_n21246_), .ZN(new_n21249_));
  NOR3_X1    g21057(.A1(new_n21239_), .A2(new_n21230_), .A3(\asqrt[46] ), .ZN(new_n21250_));
  NOR2_X1    g21058(.A1(new_n21250_), .A2(new_n21249_), .ZN(new_n21251_));
  OAI21_X1   g21059(.A1(new_n21251_), .A2(new_n21241_), .B(\asqrt[47] ), .ZN(new_n21252_));
  NOR3_X1    g21060(.A1(new_n20806_), .A2(new_n20619_), .A3(new_n20624_), .ZN(new_n21253_));
  INV_X1     g21061(.I(new_n21253_), .ZN(new_n21254_));
  NOR3_X1    g21062(.A1(new_n20619_), .A2(new_n20823_), .A3(new_n20624_), .ZN(new_n21255_));
  AOI22_X1   g21063(.A1(new_n21254_), .A2(new_n20823_), .B1(\asqrt[6] ), .B2(new_n21255_), .ZN(new_n21256_));
  INV_X1     g21064(.I(new_n21256_), .ZN(new_n21257_));
  NAND2_X1   g21065(.A1(new_n21240_), .A2(new_n2229_), .ZN(new_n21258_));
  OAI21_X1   g21066(.A1(new_n21251_), .A2(new_n21258_), .B(new_n21257_), .ZN(new_n21259_));
  AOI21_X1   g21067(.A1(new_n21259_), .A2(new_n21252_), .B(new_n1956_), .ZN(new_n21260_));
  INV_X1     g21068(.I(new_n20626_), .ZN(new_n21261_));
  NOR2_X1    g21069(.A1(new_n20625_), .A2(new_n20633_), .ZN(new_n21262_));
  NOR3_X1    g21070(.A1(new_n21261_), .A2(new_n21262_), .A3(new_n20632_), .ZN(new_n21263_));
  NOR3_X1    g21071(.A1(new_n20806_), .A2(new_n21261_), .A3(new_n21262_), .ZN(new_n21264_));
  INV_X1     g21072(.I(new_n21264_), .ZN(new_n21265_));
  AOI22_X1   g21073(.A1(new_n21265_), .A2(new_n20632_), .B1(\asqrt[6] ), .B2(new_n21263_), .ZN(new_n21266_));
  OAI21_X1   g21074(.A1(new_n21249_), .A2(new_n21250_), .B(new_n21240_), .ZN(new_n21267_));
  AOI21_X1   g21075(.A1(new_n21267_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n21268_));
  AOI21_X1   g21076(.A1(new_n21268_), .A2(new_n21259_), .B(new_n21266_), .ZN(new_n21269_));
  OAI21_X1   g21077(.A1(new_n21269_), .A2(new_n21260_), .B(\asqrt[49] ), .ZN(new_n21270_));
  INV_X1     g21078(.I(new_n21270_), .ZN(new_n21271_));
  INV_X1     g21079(.I(new_n20640_), .ZN(new_n21272_));
  INV_X1     g21080(.I(new_n20634_), .ZN(new_n21273_));
  INV_X1     g21081(.I(new_n20642_), .ZN(new_n21274_));
  NOR2_X1    g21082(.A1(new_n21274_), .A2(new_n21273_), .ZN(new_n21275_));
  NOR3_X1    g21083(.A1(new_n20806_), .A2(new_n20635_), .A3(new_n21275_), .ZN(new_n21276_));
  INV_X1     g21084(.I(new_n21276_), .ZN(new_n21277_));
  NOR3_X1    g21085(.A1(new_n21275_), .A2(new_n20635_), .A3(new_n21272_), .ZN(new_n21278_));
  AOI22_X1   g21086(.A1(new_n21277_), .A2(new_n21272_), .B1(\asqrt[6] ), .B2(new_n21278_), .ZN(new_n21279_));
  NOR3_X1    g21087(.A1(new_n21269_), .A2(new_n21260_), .A3(\asqrt[49] ), .ZN(new_n21280_));
  NOR2_X1    g21088(.A1(new_n21280_), .A2(new_n21279_), .ZN(new_n21281_));
  OAI21_X1   g21089(.A1(new_n21281_), .A2(new_n21271_), .B(\asqrt[50] ), .ZN(new_n21282_));
  NOR3_X1    g21090(.A1(new_n20645_), .A2(new_n20822_), .A3(new_n20650_), .ZN(new_n21283_));
  NOR3_X1    g21091(.A1(new_n20806_), .A2(new_n20645_), .A3(new_n20650_), .ZN(new_n21284_));
  INV_X1     g21092(.I(new_n21284_), .ZN(new_n21285_));
  AOI22_X1   g21093(.A1(new_n21285_), .A2(new_n20822_), .B1(\asqrt[6] ), .B2(new_n21283_), .ZN(new_n21286_));
  INV_X1     g21094(.I(new_n21286_), .ZN(new_n21287_));
  NAND2_X1   g21095(.A1(new_n21270_), .A2(new_n1612_), .ZN(new_n21288_));
  OAI21_X1   g21096(.A1(new_n21281_), .A2(new_n21288_), .B(new_n21287_), .ZN(new_n21289_));
  AOI21_X1   g21097(.A1(new_n21289_), .A2(new_n21282_), .B(new_n1376_), .ZN(new_n21290_));
  INV_X1     g21098(.I(new_n20652_), .ZN(new_n21291_));
  NOR2_X1    g21099(.A1(new_n20651_), .A2(new_n20659_), .ZN(new_n21292_));
  NOR3_X1    g21100(.A1(new_n20806_), .A2(new_n21291_), .A3(new_n21292_), .ZN(new_n21293_));
  INV_X1     g21101(.I(new_n21293_), .ZN(new_n21294_));
  NOR3_X1    g21102(.A1(new_n21291_), .A2(new_n20658_), .A3(new_n21292_), .ZN(new_n21295_));
  AOI22_X1   g21103(.A1(new_n21294_), .A2(new_n20658_), .B1(\asqrt[6] ), .B2(new_n21295_), .ZN(new_n21296_));
  OAI21_X1   g21104(.A1(new_n21279_), .A2(new_n21280_), .B(new_n21270_), .ZN(new_n21297_));
  AOI21_X1   g21105(.A1(new_n21297_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n21298_));
  AOI21_X1   g21106(.A1(new_n21298_), .A2(new_n21289_), .B(new_n21296_), .ZN(new_n21299_));
  OAI21_X1   g21107(.A1(new_n21299_), .A2(new_n21290_), .B(\asqrt[52] ), .ZN(new_n21300_));
  INV_X1     g21108(.I(new_n21300_), .ZN(new_n21301_));
  INV_X1     g21109(.I(new_n20666_), .ZN(new_n21302_));
  INV_X1     g21110(.I(new_n20660_), .ZN(new_n21303_));
  INV_X1     g21111(.I(new_n20668_), .ZN(new_n21304_));
  NOR2_X1    g21112(.A1(new_n21304_), .A2(new_n21303_), .ZN(new_n21305_));
  NOR3_X1    g21113(.A1(new_n21305_), .A2(new_n20661_), .A3(new_n21302_), .ZN(new_n21306_));
  NOR3_X1    g21114(.A1(new_n20806_), .A2(new_n20661_), .A3(new_n21305_), .ZN(new_n21307_));
  INV_X1     g21115(.I(new_n21307_), .ZN(new_n21308_));
  AOI22_X1   g21116(.A1(new_n21308_), .A2(new_n21302_), .B1(\asqrt[6] ), .B2(new_n21306_), .ZN(new_n21309_));
  NOR3_X1    g21117(.A1(new_n21299_), .A2(new_n21290_), .A3(\asqrt[52] ), .ZN(new_n21310_));
  NOR2_X1    g21118(.A1(new_n21310_), .A2(new_n21309_), .ZN(new_n21311_));
  OAI21_X1   g21119(.A1(new_n21311_), .A2(new_n21301_), .B(\asqrt[53] ), .ZN(new_n21312_));
  NOR3_X1    g21120(.A1(new_n20806_), .A2(new_n20671_), .A3(new_n20713_), .ZN(new_n21313_));
  INV_X1     g21121(.I(new_n21313_), .ZN(new_n21314_));
  NOR3_X1    g21122(.A1(new_n20671_), .A2(new_n20821_), .A3(new_n20713_), .ZN(new_n21315_));
  AOI22_X1   g21123(.A1(new_n21314_), .A2(new_n20821_), .B1(\asqrt[6] ), .B2(new_n21315_), .ZN(new_n21316_));
  INV_X1     g21124(.I(new_n21316_), .ZN(new_n21317_));
  NAND2_X1   g21125(.A1(new_n21300_), .A2(new_n1103_), .ZN(new_n21318_));
  OAI21_X1   g21126(.A1(new_n21311_), .A2(new_n21318_), .B(new_n21317_), .ZN(new_n21319_));
  AOI21_X1   g21127(.A1(new_n21319_), .A2(new_n21312_), .B(new_n904_), .ZN(new_n21320_));
  INV_X1     g21128(.I(new_n20679_), .ZN(new_n21321_));
  NOR2_X1    g21129(.A1(new_n20686_), .A2(new_n20678_), .ZN(new_n21322_));
  NOR3_X1    g21130(.A1(new_n21321_), .A2(new_n20685_), .A3(new_n21322_), .ZN(new_n21323_));
  NOR3_X1    g21131(.A1(new_n20806_), .A2(new_n21321_), .A3(new_n21322_), .ZN(new_n21324_));
  INV_X1     g21132(.I(new_n21324_), .ZN(new_n21325_));
  AOI22_X1   g21133(.A1(new_n21325_), .A2(new_n20685_), .B1(\asqrt[6] ), .B2(new_n21323_), .ZN(new_n21326_));
  OAI21_X1   g21134(.A1(new_n21309_), .A2(new_n21310_), .B(new_n21300_), .ZN(new_n21327_));
  AOI21_X1   g21135(.A1(new_n21327_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n21328_));
  AOI21_X1   g21136(.A1(new_n21328_), .A2(new_n21319_), .B(new_n21326_), .ZN(new_n21329_));
  OAI21_X1   g21137(.A1(new_n21329_), .A2(new_n21320_), .B(\asqrt[55] ), .ZN(new_n21330_));
  INV_X1     g21138(.I(new_n21330_), .ZN(new_n21331_));
  NOR2_X1    g21139(.A1(new_n20697_), .A2(new_n20690_), .ZN(new_n21332_));
  NOR3_X1    g21140(.A1(new_n20806_), .A2(new_n20688_), .A3(new_n21332_), .ZN(new_n21333_));
  INV_X1     g21141(.I(new_n21333_), .ZN(new_n21334_));
  NOR3_X1    g21142(.A1(new_n21332_), .A2(new_n20688_), .A3(new_n20696_), .ZN(new_n21335_));
  AOI22_X1   g21143(.A1(new_n21334_), .A2(new_n20696_), .B1(\asqrt[6] ), .B2(new_n21335_), .ZN(new_n21336_));
  NOR3_X1    g21144(.A1(new_n21329_), .A2(new_n21320_), .A3(\asqrt[55] ), .ZN(new_n21337_));
  NOR2_X1    g21145(.A1(new_n21337_), .A2(new_n21336_), .ZN(new_n21338_));
  OAI21_X1   g21146(.A1(new_n21338_), .A2(new_n21331_), .B(\asqrt[56] ), .ZN(new_n21339_));
  NOR3_X1    g21147(.A1(new_n20699_), .A2(new_n20820_), .A3(new_n20745_), .ZN(new_n21340_));
  NOR3_X1    g21148(.A1(new_n20806_), .A2(new_n20699_), .A3(new_n20745_), .ZN(new_n21341_));
  INV_X1     g21149(.I(new_n21341_), .ZN(new_n21342_));
  AOI22_X1   g21150(.A1(new_n21342_), .A2(new_n20820_), .B1(\asqrt[6] ), .B2(new_n21340_), .ZN(new_n21343_));
  INV_X1     g21151(.I(new_n21343_), .ZN(new_n21344_));
  NAND2_X1   g21152(.A1(new_n21330_), .A2(new_n703_), .ZN(new_n21345_));
  OAI21_X1   g21153(.A1(new_n21338_), .A2(new_n21345_), .B(new_n21344_), .ZN(new_n21346_));
  AOI21_X1   g21154(.A1(new_n21346_), .A2(new_n21339_), .B(new_n531_), .ZN(new_n21347_));
  INV_X1     g21155(.I(new_n20706_), .ZN(new_n21348_));
  NOR2_X1    g21156(.A1(new_n20718_), .A2(new_n20705_), .ZN(new_n21349_));
  NOR3_X1    g21157(.A1(new_n20806_), .A2(new_n21348_), .A3(new_n21349_), .ZN(new_n21350_));
  INV_X1     g21158(.I(new_n21350_), .ZN(new_n21351_));
  NOR3_X1    g21159(.A1(new_n21348_), .A2(new_n20712_), .A3(new_n21349_), .ZN(new_n21352_));
  AOI22_X1   g21160(.A1(new_n21351_), .A2(new_n20712_), .B1(\asqrt[6] ), .B2(new_n21352_), .ZN(new_n21353_));
  OAI21_X1   g21161(.A1(new_n21336_), .A2(new_n21337_), .B(new_n21330_), .ZN(new_n21354_));
  AOI21_X1   g21162(.A1(new_n21354_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n21355_));
  AOI21_X1   g21163(.A1(new_n21355_), .A2(new_n21346_), .B(new_n21353_), .ZN(new_n21356_));
  OAI21_X1   g21164(.A1(new_n21356_), .A2(new_n21347_), .B(\asqrt[58] ), .ZN(new_n21357_));
  NOR2_X1    g21165(.A1(new_n20729_), .A2(new_n20722_), .ZN(new_n21358_));
  NOR3_X1    g21166(.A1(new_n21358_), .A2(new_n20720_), .A3(new_n20728_), .ZN(new_n21359_));
  NOR3_X1    g21167(.A1(new_n20806_), .A2(new_n20720_), .A3(new_n21358_), .ZN(new_n21360_));
  INV_X1     g21168(.I(new_n21360_), .ZN(new_n21361_));
  AOI22_X1   g21169(.A1(new_n21361_), .A2(new_n20728_), .B1(\asqrt[6] ), .B2(new_n21359_), .ZN(new_n21362_));
  INV_X1     g21170(.I(new_n21362_), .ZN(new_n21363_));
  INV_X1     g21171(.I(new_n21336_), .ZN(new_n21364_));
  INV_X1     g21172(.I(new_n21309_), .ZN(new_n21365_));
  INV_X1     g21173(.I(new_n21279_), .ZN(new_n21366_));
  INV_X1     g21174(.I(new_n21249_), .ZN(new_n21367_));
  INV_X1     g21175(.I(new_n21219_), .ZN(new_n21368_));
  INV_X1     g21176(.I(new_n21191_), .ZN(new_n21369_));
  INV_X1     g21177(.I(new_n21165_), .ZN(new_n21370_));
  INV_X1     g21178(.I(new_n21138_), .ZN(new_n21371_));
  INV_X1     g21179(.I(new_n21111_), .ZN(new_n21372_));
  INV_X1     g21180(.I(new_n21084_), .ZN(new_n21373_));
  INV_X1     g21181(.I(new_n21054_), .ZN(new_n21374_));
  INV_X1     g21182(.I(new_n21024_), .ZN(new_n21375_));
  INV_X1     g21183(.I(new_n20994_), .ZN(new_n21376_));
  INV_X1     g21184(.I(new_n20963_), .ZN(new_n21377_));
  INV_X1     g21185(.I(new_n20937_), .ZN(new_n21378_));
  NAND2_X1   g21186(.A1(new_n20878_), .A2(new_n18275_), .ZN(new_n21379_));
  OAI21_X1   g21187(.A1(new_n21379_), .A2(new_n20911_), .B(new_n20892_), .ZN(new_n21380_));
  AOI21_X1   g21188(.A1(new_n21380_), .A2(new_n20921_), .B(new_n17623_), .ZN(new_n21381_));
  NOR2_X1    g21189(.A1(new_n20886_), .A2(\asqrt[11] ), .ZN(new_n21382_));
  AOI21_X1   g21190(.A1(new_n21382_), .A2(new_n21380_), .B(new_n20919_), .ZN(new_n21383_));
  OAI21_X1   g21191(.A1(new_n21383_), .A2(new_n21381_), .B(\asqrt[12] ), .ZN(new_n21384_));
  NAND2_X1   g21192(.A1(new_n21384_), .A2(new_n16389_), .ZN(new_n21385_));
  OAI21_X1   g21193(.A1(new_n21385_), .A2(new_n20931_), .B(new_n21378_), .ZN(new_n21386_));
  NAND3_X1   g21194(.A1(new_n21386_), .A2(new_n15770_), .A3(new_n20932_), .ZN(new_n21387_));
  AOI22_X1   g21195(.A1(new_n21387_), .A2(new_n20946_), .B1(\asqrt[14] ), .B2(new_n20954_), .ZN(new_n21388_));
  OAI21_X1   g21196(.A1(new_n21388_), .A2(new_n15067_), .B(new_n14601_), .ZN(new_n21389_));
  OAI21_X1   g21197(.A1(new_n21389_), .A2(new_n20956_), .B(new_n21377_), .ZN(new_n21390_));
  AOI21_X1   g21198(.A1(new_n21390_), .A2(new_n20957_), .B(new_n14017_), .ZN(new_n21391_));
  AOI21_X1   g21199(.A1(new_n21386_), .A2(new_n20932_), .B(new_n15770_), .ZN(new_n21392_));
  NOR3_X1    g21200(.A1(new_n21383_), .A2(new_n21381_), .A3(\asqrt[12] ), .ZN(new_n21393_));
  OAI21_X1   g21201(.A1(new_n20928_), .A2(new_n21393_), .B(new_n21384_), .ZN(new_n21394_));
  AOI21_X1   g21202(.A1(new_n21394_), .A2(\asqrt[13] ), .B(\asqrt[14] ), .ZN(new_n21395_));
  AOI21_X1   g21203(.A1(new_n21395_), .A2(new_n21386_), .B(new_n20945_), .ZN(new_n21396_));
  NOR3_X1    g21204(.A1(new_n21396_), .A2(\asqrt[15] ), .A3(new_n21392_), .ZN(new_n21397_));
  OAI22_X1   g21205(.A1(new_n21397_), .A2(new_n20953_), .B1(new_n21388_), .B2(new_n15067_), .ZN(new_n21398_));
  AOI21_X1   g21206(.A1(new_n21398_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n21399_));
  AOI21_X1   g21207(.A1(new_n21399_), .A2(new_n21390_), .B(new_n20971_), .ZN(new_n21400_));
  OAI21_X1   g21208(.A1(new_n21400_), .A2(new_n21391_), .B(\asqrt[18] ), .ZN(new_n21401_));
  NAND2_X1   g21209(.A1(new_n21401_), .A2(new_n12913_), .ZN(new_n21402_));
  OAI21_X1   g21210(.A1(new_n21402_), .A2(new_n20984_), .B(new_n21376_), .ZN(new_n21403_));
  AOI21_X1   g21211(.A1(new_n21403_), .A2(new_n20985_), .B(new_n12364_), .ZN(new_n21404_));
  NOR3_X1    g21212(.A1(new_n21400_), .A2(\asqrt[18] ), .A3(new_n21391_), .ZN(new_n21405_));
  OAI21_X1   g21213(.A1(new_n20981_), .A2(new_n21405_), .B(new_n21401_), .ZN(new_n21406_));
  AOI21_X1   g21214(.A1(new_n21406_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n21407_));
  AOI21_X1   g21215(.A1(new_n21407_), .A2(new_n21403_), .B(new_n21002_), .ZN(new_n21408_));
  OAI21_X1   g21216(.A1(new_n21408_), .A2(new_n21404_), .B(\asqrt[21] ), .ZN(new_n21409_));
  NAND2_X1   g21217(.A1(new_n21409_), .A2(new_n11326_), .ZN(new_n21410_));
  OAI21_X1   g21218(.A1(new_n21410_), .A2(new_n21014_), .B(new_n21375_), .ZN(new_n21411_));
  AOI21_X1   g21219(.A1(new_n21411_), .A2(new_n21015_), .B(new_n10812_), .ZN(new_n21412_));
  NOR3_X1    g21220(.A1(new_n21408_), .A2(\asqrt[21] ), .A3(new_n21404_), .ZN(new_n21413_));
  OAI21_X1   g21221(.A1(new_n21011_), .A2(new_n21413_), .B(new_n21409_), .ZN(new_n21414_));
  AOI21_X1   g21222(.A1(new_n21414_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n21415_));
  AOI21_X1   g21223(.A1(new_n21415_), .A2(new_n21411_), .B(new_n21032_), .ZN(new_n21416_));
  OAI21_X1   g21224(.A1(new_n21416_), .A2(new_n21412_), .B(\asqrt[24] ), .ZN(new_n21417_));
  NAND2_X1   g21225(.A1(new_n21417_), .A2(new_n9846_), .ZN(new_n21418_));
  OAI21_X1   g21226(.A1(new_n21418_), .A2(new_n21044_), .B(new_n21374_), .ZN(new_n21419_));
  AOI21_X1   g21227(.A1(new_n21419_), .A2(new_n21045_), .B(new_n9317_), .ZN(new_n21420_));
  NOR3_X1    g21228(.A1(new_n21416_), .A2(\asqrt[24] ), .A3(new_n21412_), .ZN(new_n21421_));
  OAI21_X1   g21229(.A1(new_n21041_), .A2(new_n21421_), .B(new_n21417_), .ZN(new_n21422_));
  AOI21_X1   g21230(.A1(new_n21422_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n21423_));
  AOI21_X1   g21231(.A1(new_n21423_), .A2(new_n21419_), .B(new_n21062_), .ZN(new_n21424_));
  OAI21_X1   g21232(.A1(new_n21424_), .A2(new_n21420_), .B(\asqrt[27] ), .ZN(new_n21425_));
  NAND2_X1   g21233(.A1(new_n21425_), .A2(new_n8483_), .ZN(new_n21426_));
  OAI21_X1   g21234(.A1(new_n21426_), .A2(new_n21074_), .B(new_n21373_), .ZN(new_n21427_));
  AOI21_X1   g21235(.A1(new_n21427_), .A2(new_n21075_), .B(new_n8036_), .ZN(new_n21428_));
  NOR3_X1    g21236(.A1(new_n21424_), .A2(\asqrt[27] ), .A3(new_n21420_), .ZN(new_n21429_));
  OAI21_X1   g21237(.A1(new_n21071_), .A2(new_n21429_), .B(new_n21425_), .ZN(new_n21430_));
  AOI21_X1   g21238(.A1(new_n21430_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n21431_));
  AOI21_X1   g21239(.A1(new_n21431_), .A2(new_n21427_), .B(new_n21092_), .ZN(new_n21432_));
  OAI21_X1   g21240(.A1(new_n21432_), .A2(new_n21428_), .B(\asqrt[30] ), .ZN(new_n21433_));
  NAND2_X1   g21241(.A1(new_n21433_), .A2(new_n7229_), .ZN(new_n21434_));
  OAI21_X1   g21242(.A1(new_n21434_), .A2(new_n21104_), .B(new_n21372_), .ZN(new_n21435_));
  AOI21_X1   g21243(.A1(new_n21435_), .A2(new_n21105_), .B(new_n6824_), .ZN(new_n21436_));
  NOR3_X1    g21244(.A1(new_n21432_), .A2(\asqrt[30] ), .A3(new_n21428_), .ZN(new_n21437_));
  OAI21_X1   g21245(.A1(new_n21101_), .A2(new_n21437_), .B(new_n21433_), .ZN(new_n21438_));
  AOI21_X1   g21246(.A1(new_n21438_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n21439_));
  AOI21_X1   g21247(.A1(new_n21439_), .A2(new_n21435_), .B(new_n21119_), .ZN(new_n21440_));
  OAI21_X1   g21248(.A1(new_n21440_), .A2(new_n21436_), .B(\asqrt[33] ), .ZN(new_n21441_));
  NAND2_X1   g21249(.A1(new_n21441_), .A2(new_n6077_), .ZN(new_n21442_));
  OAI21_X1   g21250(.A1(new_n21442_), .A2(new_n21131_), .B(new_n21371_), .ZN(new_n21443_));
  AOI21_X1   g21251(.A1(new_n21443_), .A2(new_n21132_), .B(new_n5708_), .ZN(new_n21444_));
  NOR3_X1    g21252(.A1(new_n21440_), .A2(\asqrt[33] ), .A3(new_n21436_), .ZN(new_n21445_));
  OAI21_X1   g21253(.A1(new_n21128_), .A2(new_n21445_), .B(new_n21441_), .ZN(new_n21446_));
  AOI21_X1   g21254(.A1(new_n21446_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n21447_));
  AOI21_X1   g21255(.A1(new_n21447_), .A2(new_n21443_), .B(new_n21146_), .ZN(new_n21448_));
  OAI21_X1   g21256(.A1(new_n21448_), .A2(new_n21444_), .B(\asqrt[36] ), .ZN(new_n21449_));
  NAND2_X1   g21257(.A1(new_n21449_), .A2(new_n5024_), .ZN(new_n21450_));
  OAI21_X1   g21258(.A1(new_n21450_), .A2(new_n21158_), .B(new_n21370_), .ZN(new_n21451_));
  AOI21_X1   g21259(.A1(new_n21451_), .A2(new_n21159_), .B(new_n4696_), .ZN(new_n21452_));
  NOR3_X1    g21260(.A1(new_n21448_), .A2(\asqrt[36] ), .A3(new_n21444_), .ZN(new_n21453_));
  OAI21_X1   g21261(.A1(new_n21155_), .A2(new_n21453_), .B(new_n21449_), .ZN(new_n21454_));
  AOI21_X1   g21262(.A1(new_n21454_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n21455_));
  AOI21_X1   g21263(.A1(new_n21455_), .A2(new_n21451_), .B(new_n21173_), .ZN(new_n21456_));
  OAI21_X1   g21264(.A1(new_n21456_), .A2(new_n21452_), .B(\asqrt[39] ), .ZN(new_n21457_));
  NAND2_X1   g21265(.A1(new_n21457_), .A2(new_n4071_), .ZN(new_n21458_));
  OAI21_X1   g21266(.A1(new_n21458_), .A2(new_n21184_), .B(new_n21369_), .ZN(new_n21459_));
  AOI21_X1   g21267(.A1(new_n21459_), .A2(new_n21185_), .B(new_n3782_), .ZN(new_n21460_));
  NOR3_X1    g21268(.A1(new_n21456_), .A2(\asqrt[39] ), .A3(new_n21452_), .ZN(new_n21461_));
  OAI21_X1   g21269(.A1(new_n21181_), .A2(new_n21461_), .B(new_n21457_), .ZN(new_n21462_));
  AOI21_X1   g21270(.A1(new_n21462_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n21463_));
  AOI21_X1   g21271(.A1(new_n21463_), .A2(new_n21459_), .B(new_n21199_), .ZN(new_n21464_));
  OAI21_X1   g21272(.A1(new_n21464_), .A2(new_n21460_), .B(\asqrt[42] ), .ZN(new_n21465_));
  NAND2_X1   g21273(.A1(new_n21465_), .A2(new_n3218_), .ZN(new_n21466_));
  OAI21_X1   g21274(.A1(new_n21466_), .A2(new_n21210_), .B(new_n21368_), .ZN(new_n21467_));
  AOI21_X1   g21275(.A1(new_n21467_), .A2(new_n21211_), .B(new_n2954_), .ZN(new_n21468_));
  NOR3_X1    g21276(.A1(new_n21464_), .A2(\asqrt[42] ), .A3(new_n21460_), .ZN(new_n21469_));
  OAI21_X1   g21277(.A1(new_n21207_), .A2(new_n21469_), .B(new_n21465_), .ZN(new_n21470_));
  AOI21_X1   g21278(.A1(new_n21470_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n21471_));
  AOI21_X1   g21279(.A1(new_n21471_), .A2(new_n21467_), .B(new_n21226_), .ZN(new_n21472_));
  OAI21_X1   g21280(.A1(new_n21472_), .A2(new_n21468_), .B(\asqrt[45] ), .ZN(new_n21473_));
  NAND2_X1   g21281(.A1(new_n21473_), .A2(new_n2465_), .ZN(new_n21474_));
  OAI21_X1   g21282(.A1(new_n21474_), .A2(new_n21239_), .B(new_n21367_), .ZN(new_n21475_));
  AOI21_X1   g21283(.A1(new_n21475_), .A2(new_n21240_), .B(new_n2229_), .ZN(new_n21476_));
  NOR3_X1    g21284(.A1(new_n21472_), .A2(\asqrt[45] ), .A3(new_n21468_), .ZN(new_n21477_));
  OAI21_X1   g21285(.A1(new_n21236_), .A2(new_n21477_), .B(new_n21473_), .ZN(new_n21478_));
  AOI21_X1   g21286(.A1(new_n21478_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n21479_));
  AOI21_X1   g21287(.A1(new_n21479_), .A2(new_n21475_), .B(new_n21256_), .ZN(new_n21480_));
  OAI21_X1   g21288(.A1(new_n21480_), .A2(new_n21476_), .B(\asqrt[48] ), .ZN(new_n21481_));
  NAND2_X1   g21289(.A1(new_n21481_), .A2(new_n1806_), .ZN(new_n21482_));
  OAI21_X1   g21290(.A1(new_n21482_), .A2(new_n21269_), .B(new_n21366_), .ZN(new_n21483_));
  AOI21_X1   g21291(.A1(new_n21483_), .A2(new_n21270_), .B(new_n1612_), .ZN(new_n21484_));
  NOR3_X1    g21292(.A1(new_n21480_), .A2(\asqrt[48] ), .A3(new_n21476_), .ZN(new_n21485_));
  OAI21_X1   g21293(.A1(new_n21266_), .A2(new_n21485_), .B(new_n21481_), .ZN(new_n21486_));
  AOI21_X1   g21294(.A1(new_n21486_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n21487_));
  AOI21_X1   g21295(.A1(new_n21487_), .A2(new_n21483_), .B(new_n21286_), .ZN(new_n21488_));
  OAI21_X1   g21296(.A1(new_n21488_), .A2(new_n21484_), .B(\asqrt[51] ), .ZN(new_n21489_));
  NAND2_X1   g21297(.A1(new_n21489_), .A2(new_n1256_), .ZN(new_n21490_));
  OAI21_X1   g21298(.A1(new_n21490_), .A2(new_n21299_), .B(new_n21365_), .ZN(new_n21491_));
  NAND3_X1   g21299(.A1(new_n21491_), .A2(new_n1103_), .A3(new_n21300_), .ZN(new_n21492_));
  AOI22_X1   g21300(.A1(new_n21492_), .A2(new_n21317_), .B1(\asqrt[53] ), .B2(new_n21327_), .ZN(new_n21493_));
  OAI21_X1   g21301(.A1(new_n21493_), .A2(new_n904_), .B(new_n823_), .ZN(new_n21494_));
  OAI21_X1   g21302(.A1(new_n21494_), .A2(new_n21329_), .B(new_n21364_), .ZN(new_n21495_));
  NAND3_X1   g21303(.A1(new_n21495_), .A2(new_n703_), .A3(new_n21330_), .ZN(new_n21496_));
  AOI22_X1   g21304(.A1(new_n21496_), .A2(new_n21344_), .B1(\asqrt[56] ), .B2(new_n21354_), .ZN(new_n21497_));
  OAI21_X1   g21305(.A1(new_n21497_), .A2(new_n531_), .B(new_n436_), .ZN(new_n21498_));
  OAI21_X1   g21306(.A1(new_n21498_), .A2(new_n21356_), .B(new_n21363_), .ZN(new_n21499_));
  AOI21_X1   g21307(.A1(new_n21499_), .A2(new_n21357_), .B(new_n327_), .ZN(new_n21500_));
  NOR3_X1    g21308(.A1(new_n20806_), .A2(new_n20731_), .A3(new_n20777_), .ZN(new_n21501_));
  INV_X1     g21309(.I(new_n21501_), .ZN(new_n21502_));
  NOR3_X1    g21310(.A1(new_n20731_), .A2(new_n20819_), .A3(new_n20777_), .ZN(new_n21503_));
  AOI22_X1   g21311(.A1(new_n21502_), .A2(new_n20819_), .B1(\asqrt[6] ), .B2(new_n21503_), .ZN(new_n21504_));
  NAND2_X1   g21312(.A1(new_n21357_), .A2(new_n327_), .ZN(new_n21505_));
  INV_X1     g21313(.I(new_n21505_), .ZN(new_n21506_));
  AOI21_X1   g21314(.A1(new_n21506_), .A2(new_n21499_), .B(new_n21504_), .ZN(new_n21507_));
  OAI21_X1   g21315(.A1(new_n21507_), .A2(new_n21500_), .B(\asqrt[60] ), .ZN(new_n21508_));
  INV_X1     g21316(.I(new_n20738_), .ZN(new_n21509_));
  NOR2_X1    g21317(.A1(new_n20750_), .A2(new_n20737_), .ZN(new_n21510_));
  NOR3_X1    g21318(.A1(new_n21509_), .A2(new_n20744_), .A3(new_n21510_), .ZN(new_n21511_));
  NOR3_X1    g21319(.A1(new_n20806_), .A2(new_n21509_), .A3(new_n21510_), .ZN(new_n21512_));
  INV_X1     g21320(.I(new_n21512_), .ZN(new_n21513_));
  AOI22_X1   g21321(.A1(new_n21513_), .A2(new_n20744_), .B1(\asqrt[6] ), .B2(new_n21511_), .ZN(new_n21514_));
  INV_X1     g21322(.I(new_n21514_), .ZN(new_n21515_));
  INV_X1     g21323(.I(new_n21357_), .ZN(new_n21516_));
  NOR3_X1    g21324(.A1(new_n21356_), .A2(new_n21347_), .A3(\asqrt[58] ), .ZN(new_n21517_));
  NOR2_X1    g21325(.A1(new_n21517_), .A2(new_n21362_), .ZN(new_n21518_));
  OAI21_X1   g21326(.A1(new_n21518_), .A2(new_n21516_), .B(\asqrt[59] ), .ZN(new_n21519_));
  NAND2_X1   g21327(.A1(new_n21519_), .A2(new_n306_), .ZN(new_n21520_));
  OAI21_X1   g21328(.A1(new_n21520_), .A2(new_n21507_), .B(new_n21515_), .ZN(new_n21521_));
  AOI21_X1   g21329(.A1(new_n21521_), .A2(new_n21508_), .B(new_n218_), .ZN(new_n21522_));
  NOR2_X1    g21330(.A1(new_n20754_), .A2(new_n20761_), .ZN(new_n21523_));
  NOR3_X1    g21331(.A1(new_n20806_), .A2(new_n20752_), .A3(new_n21523_), .ZN(new_n21524_));
  INV_X1     g21332(.I(new_n21524_), .ZN(new_n21525_));
  NOR3_X1    g21333(.A1(new_n21523_), .A2(new_n20752_), .A3(new_n20760_), .ZN(new_n21526_));
  AOI22_X1   g21334(.A1(new_n21525_), .A2(new_n20760_), .B1(\asqrt[6] ), .B2(new_n21526_), .ZN(new_n21527_));
  INV_X1     g21335(.I(new_n21504_), .ZN(new_n21528_));
  OAI21_X1   g21336(.A1(new_n21518_), .A2(new_n21505_), .B(new_n21528_), .ZN(new_n21529_));
  AOI21_X1   g21337(.A1(new_n21529_), .A2(new_n21519_), .B(new_n306_), .ZN(new_n21530_));
  NOR2_X1    g21338(.A1(new_n21530_), .A2(\asqrt[61] ), .ZN(new_n21531_));
  AOI21_X1   g21339(.A1(new_n21531_), .A2(new_n21521_), .B(new_n21527_), .ZN(new_n21532_));
  OAI21_X1   g21340(.A1(new_n21532_), .A2(new_n21522_), .B(\asqrt[62] ), .ZN(new_n21533_));
  NOR3_X1    g21341(.A1(new_n20763_), .A2(new_n20818_), .A3(new_n20816_), .ZN(new_n21534_));
  NOR3_X1    g21342(.A1(new_n20806_), .A2(new_n20763_), .A3(new_n20816_), .ZN(new_n21535_));
  INV_X1     g21343(.I(new_n21535_), .ZN(new_n21536_));
  AOI22_X1   g21344(.A1(new_n21536_), .A2(new_n20818_), .B1(\asqrt[6] ), .B2(new_n21534_), .ZN(new_n21537_));
  INV_X1     g21345(.I(new_n21537_), .ZN(new_n21538_));
  OAI21_X1   g21346(.A1(new_n21362_), .A2(new_n21517_), .B(new_n21357_), .ZN(new_n21539_));
  AOI21_X1   g21347(.A1(new_n21539_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n21540_));
  AOI21_X1   g21348(.A1(new_n21540_), .A2(new_n21529_), .B(new_n21514_), .ZN(new_n21541_));
  OAI21_X1   g21349(.A1(new_n21541_), .A2(new_n21530_), .B(\asqrt[61] ), .ZN(new_n21542_));
  NAND2_X1   g21350(.A1(new_n21542_), .A2(new_n207_), .ZN(new_n21543_));
  OAI21_X1   g21351(.A1(new_n21543_), .A2(new_n21532_), .B(new_n21538_), .ZN(new_n21544_));
  NAND2_X1   g21352(.A1(new_n20770_), .A2(new_n20855_), .ZN(new_n21545_));
  OAI21_X1   g21353(.A1(new_n20806_), .A2(new_n21545_), .B(new_n20776_), .ZN(new_n21546_));
  NAND4_X1   g21354(.A1(\asqrt[6] ), .A2(new_n20770_), .A3(new_n20775_), .A4(new_n20855_), .ZN(new_n21547_));
  NAND2_X1   g21355(.A1(new_n21547_), .A2(new_n21546_), .ZN(new_n21548_));
  NOR2_X1    g21356(.A1(new_n20856_), .A2(new_n20795_), .ZN(new_n21549_));
  NAND2_X1   g21357(.A1(\asqrt[6] ), .A2(new_n21549_), .ZN(new_n21550_));
  NAND3_X1   g21358(.A1(new_n21548_), .A2(new_n20867_), .A3(new_n21550_), .ZN(new_n21551_));
  AOI21_X1   g21359(.A1(new_n21544_), .A2(new_n21533_), .B(new_n21551_), .ZN(new_n21552_));
  NOR3_X1    g21360(.A1(new_n21541_), .A2(new_n21530_), .A3(\asqrt[61] ), .ZN(new_n21553_));
  OAI21_X1   g21361(.A1(new_n21527_), .A2(new_n21553_), .B(new_n21542_), .ZN(new_n21554_));
  AOI21_X1   g21362(.A1(new_n21554_), .A2(\asqrt[62] ), .B(new_n21548_), .ZN(new_n21555_));
  OAI21_X1   g21363(.A1(new_n20806_), .A2(new_n20795_), .B(new_n20856_), .ZN(new_n21556_));
  NOR2_X1    g21364(.A1(new_n21549_), .A2(new_n193_), .ZN(new_n21557_));
  NAND2_X1   g21365(.A1(new_n21556_), .A2(new_n21557_), .ZN(new_n21558_));
  INV_X1     g21366(.I(new_n21558_), .ZN(new_n21559_));
  AOI21_X1   g21367(.A1(new_n21555_), .A2(new_n21544_), .B(new_n21559_), .ZN(new_n21560_));
  OAI21_X1   g21368(.A1(\asqrt[63] ), .A2(new_n21552_), .B(new_n21560_), .ZN(\asqrt[5] ));
  NOR2_X1    g21369(.A1(\a[8] ), .A2(\a[9] ), .ZN(new_n21562_));
  INV_X1     g21370(.I(new_n21562_), .ZN(new_n21563_));
  NOR2_X1    g21371(.A1(new_n21563_), .A2(\a[10] ), .ZN(new_n21564_));
  INV_X1     g21372(.I(new_n21564_), .ZN(new_n21565_));
  NAND2_X1   g21373(.A1(new_n21544_), .A2(new_n21533_), .ZN(new_n21566_));
  INV_X1     g21374(.I(new_n21551_), .ZN(new_n21567_));
  AOI21_X1   g21375(.A1(new_n21566_), .A2(new_n21567_), .B(\asqrt[63] ), .ZN(new_n21568_));
  INV_X1     g21376(.I(new_n21527_), .ZN(new_n21569_));
  NAND3_X1   g21377(.A1(new_n21499_), .A2(new_n327_), .A3(new_n21357_), .ZN(new_n21570_));
  AOI22_X1   g21378(.A1(new_n21570_), .A2(new_n21528_), .B1(new_n21539_), .B2(\asqrt[59] ), .ZN(new_n21571_));
  OAI21_X1   g21379(.A1(new_n21571_), .A2(new_n306_), .B(new_n218_), .ZN(new_n21572_));
  OAI21_X1   g21380(.A1(new_n21572_), .A2(new_n21541_), .B(new_n21569_), .ZN(new_n21573_));
  NOR2_X1    g21381(.A1(new_n21522_), .A2(\asqrt[62] ), .ZN(new_n21574_));
  AOI21_X1   g21382(.A1(new_n21574_), .A2(new_n21573_), .B(new_n21537_), .ZN(new_n21575_));
  INV_X1     g21383(.I(new_n21548_), .ZN(new_n21576_));
  NAND2_X1   g21384(.A1(new_n21533_), .A2(new_n21576_), .ZN(new_n21577_));
  OAI21_X1   g21385(.A1(new_n21577_), .A2(new_n21575_), .B(new_n21558_), .ZN(new_n21578_));
  OAI21_X1   g21386(.A1(new_n21568_), .A2(new_n21578_), .B(\a[10] ), .ZN(new_n21579_));
  AOI21_X1   g21387(.A1(new_n21579_), .A2(new_n21565_), .B(new_n20806_), .ZN(new_n21580_));
  INV_X1     g21388(.I(\a[10] ), .ZN(new_n21581_));
  NAND3_X1   g21389(.A1(new_n21573_), .A2(new_n207_), .A3(new_n21542_), .ZN(new_n21582_));
  AOI22_X1   g21390(.A1(new_n21582_), .A2(new_n21538_), .B1(new_n21554_), .B2(\asqrt[62] ), .ZN(new_n21583_));
  OAI21_X1   g21391(.A1(new_n21583_), .A2(new_n21551_), .B(new_n193_), .ZN(new_n21584_));
  AOI21_X1   g21392(.A1(new_n21584_), .A2(new_n21560_), .B(new_n21581_), .ZN(new_n21585_));
  NAND4_X1   g21393(.A1(new_n20867_), .A2(new_n20798_), .A3(new_n20802_), .A4(new_n21565_), .ZN(new_n21586_));
  NOR2_X1    g21394(.A1(new_n21586_), .A2(new_n20793_), .ZN(new_n21587_));
  INV_X1     g21395(.I(new_n21587_), .ZN(new_n21588_));
  NOR2_X1    g21396(.A1(new_n21585_), .A2(new_n21588_), .ZN(new_n21589_));
  AOI21_X1   g21397(.A1(new_n21584_), .A2(new_n21560_), .B(new_n20809_), .ZN(new_n21590_));
  INV_X1     g21398(.I(\a[11] ), .ZN(new_n21591_));
  AOI21_X1   g21399(.A1(\asqrt[5] ), .A2(new_n21581_), .B(new_n21591_), .ZN(new_n21592_));
  NOR3_X1    g21400(.A1(new_n21589_), .A2(new_n21592_), .A3(new_n21590_), .ZN(new_n21593_));
  OAI21_X1   g21401(.A1(new_n21593_), .A2(new_n21580_), .B(\asqrt[7] ), .ZN(new_n21594_));
  OAI21_X1   g21402(.A1(new_n21568_), .A2(new_n21578_), .B(new_n20808_), .ZN(new_n21595_));
  NAND2_X1   g21403(.A1(new_n21555_), .A2(new_n21544_), .ZN(new_n21596_));
  NAND4_X1   g21404(.A1(new_n21584_), .A2(\asqrt[6] ), .A3(new_n21596_), .A4(new_n21558_), .ZN(new_n21597_));
  AOI21_X1   g21405(.A1(new_n21597_), .A2(new_n21595_), .B(new_n20807_), .ZN(new_n21598_));
  NAND3_X1   g21406(.A1(new_n21596_), .A2(\asqrt[6] ), .A3(new_n21558_), .ZN(new_n21599_));
  NOR2_X1    g21407(.A1(new_n21599_), .A2(new_n21568_), .ZN(new_n21600_));
  NOR3_X1    g21408(.A1(new_n21600_), .A2(new_n21590_), .A3(\a[12] ), .ZN(new_n21601_));
  AOI21_X1   g21409(.A1(\asqrt[5] ), .A2(\a[10] ), .B(new_n21564_), .ZN(new_n21602_));
  OAI21_X1   g21410(.A1(new_n21602_), .A2(new_n20806_), .B(new_n20262_), .ZN(new_n21603_));
  OAI22_X1   g21411(.A1(new_n21593_), .A2(new_n21603_), .B1(new_n21598_), .B2(new_n21601_), .ZN(new_n21604_));
  AOI21_X1   g21412(.A1(new_n21604_), .A2(new_n21594_), .B(new_n19573_), .ZN(new_n21605_));
  NOR3_X1    g21413(.A1(new_n20896_), .A2(new_n20898_), .A3(new_n20862_), .ZN(new_n21606_));
  NAND3_X1   g21414(.A1(\asqrt[5] ), .A2(new_n20895_), .A3(new_n20815_), .ZN(new_n21607_));
  AOI22_X1   g21415(.A1(new_n21607_), .A2(new_n20862_), .B1(\asqrt[5] ), .B2(new_n21606_), .ZN(new_n21608_));
  OAI21_X1   g21416(.A1(new_n21585_), .A2(new_n21564_), .B(\asqrt[6] ), .ZN(new_n21609_));
  AOI21_X1   g21417(.A1(new_n21584_), .A2(new_n21560_), .B(\a[10] ), .ZN(new_n21610_));
  OAI21_X1   g21418(.A1(new_n21591_), .A2(new_n21610_), .B(new_n21595_), .ZN(new_n21611_));
  OAI21_X1   g21419(.A1(new_n21611_), .A2(new_n21589_), .B(new_n21609_), .ZN(new_n21612_));
  AOI21_X1   g21420(.A1(new_n21612_), .A2(\asqrt[7] ), .B(\asqrt[8] ), .ZN(new_n21613_));
  AOI21_X1   g21421(.A1(new_n21613_), .A2(new_n21604_), .B(new_n21608_), .ZN(new_n21614_));
  OAI21_X1   g21422(.A1(new_n21614_), .A2(new_n21605_), .B(\asqrt[9] ), .ZN(new_n21615_));
  INV_X1     g21423(.I(new_n21615_), .ZN(new_n21616_));
  NOR2_X1    g21424(.A1(new_n20901_), .A2(new_n20904_), .ZN(new_n21617_));
  INV_X1     g21425(.I(new_n21617_), .ZN(new_n21618_));
  NAND4_X1   g21426(.A1(\asqrt[5] ), .A2(new_n20902_), .A3(new_n20875_), .A4(new_n21618_), .ZN(new_n21619_));
  INV_X1     g21427(.I(\asqrt[5] ), .ZN(new_n21620_));
  NOR3_X1    g21428(.A1(new_n21620_), .A2(new_n20864_), .A3(new_n21617_), .ZN(new_n21621_));
  OAI21_X1   g21429(.A1(new_n21621_), .A2(new_n20875_), .B(new_n21619_), .ZN(new_n21622_));
  INV_X1     g21430(.I(new_n21622_), .ZN(new_n21623_));
  NOR3_X1    g21431(.A1(new_n21614_), .A2(new_n21605_), .A3(\asqrt[9] ), .ZN(new_n21624_));
  NOR2_X1    g21432(.A1(new_n21624_), .A2(new_n21623_), .ZN(new_n21625_));
  OAI21_X1   g21433(.A1(new_n21625_), .A2(new_n21616_), .B(\asqrt[10] ), .ZN(new_n21626_));
  NAND2_X1   g21434(.A1(new_n20910_), .A2(new_n20905_), .ZN(new_n21627_));
  NAND3_X1   g21435(.A1(\asqrt[5] ), .A2(new_n20878_), .A3(new_n21627_), .ZN(new_n21628_));
  AND3_X2    g21436(.A1(new_n20878_), .A2(new_n20882_), .A3(new_n21627_), .Z(new_n21629_));
  AOI22_X1   g21437(.A1(new_n21628_), .A2(new_n20883_), .B1(\asqrt[5] ), .B2(new_n21629_), .ZN(new_n21630_));
  INV_X1     g21438(.I(new_n21630_), .ZN(new_n21631_));
  NAND2_X1   g21439(.A1(new_n21615_), .A2(new_n18275_), .ZN(new_n21632_));
  OAI21_X1   g21440(.A1(new_n21625_), .A2(new_n21632_), .B(new_n21631_), .ZN(new_n21633_));
  AOI21_X1   g21441(.A1(new_n21633_), .A2(new_n21626_), .B(new_n17623_), .ZN(new_n21634_));
  NOR3_X1    g21442(.A1(new_n20886_), .A2(new_n20892_), .A3(new_n20912_), .ZN(new_n21635_));
  NOR3_X1    g21443(.A1(new_n21620_), .A2(new_n20886_), .A3(new_n20912_), .ZN(new_n21636_));
  INV_X1     g21444(.I(new_n21636_), .ZN(new_n21637_));
  AOI22_X1   g21445(.A1(new_n21637_), .A2(new_n20892_), .B1(\asqrt[5] ), .B2(new_n21635_), .ZN(new_n21638_));
  OAI21_X1   g21446(.A1(new_n21623_), .A2(new_n21624_), .B(new_n21615_), .ZN(new_n21639_));
  AOI21_X1   g21447(.A1(new_n21639_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n21640_));
  AOI21_X1   g21448(.A1(new_n21640_), .A2(new_n21633_), .B(new_n21638_), .ZN(new_n21641_));
  OAI21_X1   g21449(.A1(new_n21641_), .A2(new_n21634_), .B(\asqrt[12] ), .ZN(new_n21642_));
  INV_X1     g21450(.I(new_n21642_), .ZN(new_n21643_));
  NAND2_X1   g21451(.A1(new_n21382_), .A2(new_n21380_), .ZN(new_n21644_));
  NAND3_X1   g21452(.A1(\asqrt[5] ), .A2(new_n20914_), .A3(new_n21644_), .ZN(new_n21645_));
  AND3_X2    g21453(.A1(new_n21644_), .A2(new_n20914_), .A3(new_n20919_), .Z(new_n21646_));
  AOI22_X1   g21454(.A1(new_n21645_), .A2(new_n20920_), .B1(\asqrt[5] ), .B2(new_n21646_), .ZN(new_n21647_));
  NOR3_X1    g21455(.A1(new_n21641_), .A2(new_n21634_), .A3(\asqrt[12] ), .ZN(new_n21648_));
  NOR2_X1    g21456(.A1(new_n21648_), .A2(new_n21647_), .ZN(new_n21649_));
  OAI21_X1   g21457(.A1(new_n21649_), .A2(new_n21643_), .B(\asqrt[13] ), .ZN(new_n21650_));
  INV_X1     g21458(.I(new_n20928_), .ZN(new_n21651_));
  NOR3_X1    g21459(.A1(new_n21393_), .A2(new_n20924_), .A3(new_n21651_), .ZN(new_n21652_));
  NOR3_X1    g21460(.A1(new_n21620_), .A2(new_n20924_), .A3(new_n21393_), .ZN(new_n21653_));
  INV_X1     g21461(.I(new_n21653_), .ZN(new_n21654_));
  AOI22_X1   g21462(.A1(new_n21654_), .A2(new_n21651_), .B1(\asqrt[5] ), .B2(new_n21652_), .ZN(new_n21655_));
  INV_X1     g21463(.I(new_n21655_), .ZN(new_n21656_));
  NAND2_X1   g21464(.A1(new_n21642_), .A2(new_n16389_), .ZN(new_n21657_));
  OAI21_X1   g21465(.A1(new_n21649_), .A2(new_n21657_), .B(new_n21656_), .ZN(new_n21658_));
  AOI21_X1   g21466(.A1(new_n21658_), .A2(new_n21650_), .B(new_n15770_), .ZN(new_n21659_));
  NOR3_X1    g21467(.A1(new_n21620_), .A2(new_n20933_), .A3(new_n20938_), .ZN(new_n21660_));
  INV_X1     g21468(.I(new_n21660_), .ZN(new_n21661_));
  NOR3_X1    g21469(.A1(new_n20933_), .A2(new_n21378_), .A3(new_n20938_), .ZN(new_n21662_));
  AOI22_X1   g21470(.A1(new_n21661_), .A2(new_n21378_), .B1(\asqrt[5] ), .B2(new_n21662_), .ZN(new_n21663_));
  OAI21_X1   g21471(.A1(new_n21647_), .A2(new_n21648_), .B(new_n21642_), .ZN(new_n21664_));
  AOI21_X1   g21472(.A1(new_n21664_), .A2(\asqrt[13] ), .B(\asqrt[14] ), .ZN(new_n21665_));
  AOI21_X1   g21473(.A1(new_n21665_), .A2(new_n21658_), .B(new_n21663_), .ZN(new_n21666_));
  OAI21_X1   g21474(.A1(new_n21666_), .A2(new_n21659_), .B(\asqrt[15] ), .ZN(new_n21667_));
  INV_X1     g21475(.I(new_n21667_), .ZN(new_n21668_));
  INV_X1     g21476(.I(new_n21387_), .ZN(new_n21669_));
  NOR3_X1    g21477(.A1(new_n21669_), .A2(new_n21392_), .A3(new_n20946_), .ZN(new_n21670_));
  NOR3_X1    g21478(.A1(new_n21620_), .A2(new_n21392_), .A3(new_n21669_), .ZN(new_n21671_));
  INV_X1     g21479(.I(new_n21671_), .ZN(new_n21672_));
  AOI22_X1   g21480(.A1(new_n21672_), .A2(new_n20946_), .B1(\asqrt[5] ), .B2(new_n21670_), .ZN(new_n21673_));
  NOR3_X1    g21481(.A1(new_n21666_), .A2(new_n21659_), .A3(\asqrt[15] ), .ZN(new_n21674_));
  NOR2_X1    g21482(.A1(new_n21674_), .A2(new_n21673_), .ZN(new_n21675_));
  OAI21_X1   g21483(.A1(new_n21675_), .A2(new_n21668_), .B(\asqrt[16] ), .ZN(new_n21676_));
  INV_X1     g21484(.I(new_n20953_), .ZN(new_n21677_));
  NOR3_X1    g21485(.A1(new_n21620_), .A2(new_n20949_), .A3(new_n21397_), .ZN(new_n21678_));
  INV_X1     g21486(.I(new_n21678_), .ZN(new_n21679_));
  NOR3_X1    g21487(.A1(new_n21397_), .A2(new_n20949_), .A3(new_n21677_), .ZN(new_n21680_));
  AOI22_X1   g21488(.A1(new_n21679_), .A2(new_n21677_), .B1(\asqrt[5] ), .B2(new_n21680_), .ZN(new_n21681_));
  INV_X1     g21489(.I(new_n21681_), .ZN(new_n21682_));
  NAND2_X1   g21490(.A1(new_n21667_), .A2(new_n14601_), .ZN(new_n21683_));
  OAI21_X1   g21491(.A1(new_n21675_), .A2(new_n21683_), .B(new_n21682_), .ZN(new_n21684_));
  AOI21_X1   g21492(.A1(new_n21684_), .A2(new_n21676_), .B(new_n14017_), .ZN(new_n21685_));
  NOR3_X1    g21493(.A1(new_n20958_), .A2(new_n21377_), .A3(new_n20964_), .ZN(new_n21686_));
  NOR3_X1    g21494(.A1(new_n21620_), .A2(new_n20958_), .A3(new_n20964_), .ZN(new_n21687_));
  INV_X1     g21495(.I(new_n21687_), .ZN(new_n21688_));
  AOI22_X1   g21496(.A1(new_n21688_), .A2(new_n21377_), .B1(\asqrt[5] ), .B2(new_n21686_), .ZN(new_n21689_));
  OAI21_X1   g21497(.A1(new_n21673_), .A2(new_n21674_), .B(new_n21667_), .ZN(new_n21690_));
  AOI21_X1   g21498(.A1(new_n21690_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n21691_));
  AOI21_X1   g21499(.A1(new_n21691_), .A2(new_n21684_), .B(new_n21689_), .ZN(new_n21692_));
  OAI21_X1   g21500(.A1(new_n21692_), .A2(new_n21685_), .B(\asqrt[18] ), .ZN(new_n21693_));
  INV_X1     g21501(.I(new_n21693_), .ZN(new_n21694_));
  NOR2_X1    g21502(.A1(new_n20965_), .A2(new_n20973_), .ZN(new_n21695_));
  NOR3_X1    g21503(.A1(new_n21620_), .A2(new_n21391_), .A3(new_n21695_), .ZN(new_n21696_));
  INV_X1     g21504(.I(new_n21696_), .ZN(new_n21697_));
  NOR3_X1    g21505(.A1(new_n21695_), .A2(new_n21391_), .A3(new_n20972_), .ZN(new_n21698_));
  AOI22_X1   g21506(.A1(new_n21697_), .A2(new_n20972_), .B1(\asqrt[5] ), .B2(new_n21698_), .ZN(new_n21699_));
  NOR3_X1    g21507(.A1(new_n21692_), .A2(new_n21685_), .A3(\asqrt[18] ), .ZN(new_n21700_));
  NOR2_X1    g21508(.A1(new_n21700_), .A2(new_n21699_), .ZN(new_n21701_));
  OAI21_X1   g21509(.A1(new_n21701_), .A2(new_n21694_), .B(\asqrt[19] ), .ZN(new_n21702_));
  INV_X1     g21510(.I(new_n20981_), .ZN(new_n21703_));
  NOR3_X1    g21511(.A1(new_n21405_), .A2(new_n20975_), .A3(new_n21703_), .ZN(new_n21704_));
  NOR3_X1    g21512(.A1(new_n21620_), .A2(new_n20975_), .A3(new_n21405_), .ZN(new_n21705_));
  INV_X1     g21513(.I(new_n21705_), .ZN(new_n21706_));
  AOI22_X1   g21514(.A1(new_n21706_), .A2(new_n21703_), .B1(\asqrt[5] ), .B2(new_n21704_), .ZN(new_n21707_));
  INV_X1     g21515(.I(new_n21707_), .ZN(new_n21708_));
  NAND2_X1   g21516(.A1(new_n21693_), .A2(new_n12913_), .ZN(new_n21709_));
  OAI21_X1   g21517(.A1(new_n21701_), .A2(new_n21709_), .B(new_n21708_), .ZN(new_n21710_));
  AOI21_X1   g21518(.A1(new_n21710_), .A2(new_n21702_), .B(new_n12364_), .ZN(new_n21711_));
  NOR3_X1    g21519(.A1(new_n21620_), .A2(new_n20986_), .A3(new_n20995_), .ZN(new_n21712_));
  INV_X1     g21520(.I(new_n21712_), .ZN(new_n21713_));
  NOR3_X1    g21521(.A1(new_n20986_), .A2(new_n21376_), .A3(new_n20995_), .ZN(new_n21714_));
  AOI22_X1   g21522(.A1(new_n21713_), .A2(new_n21376_), .B1(\asqrt[5] ), .B2(new_n21714_), .ZN(new_n21715_));
  OAI21_X1   g21523(.A1(new_n21699_), .A2(new_n21700_), .B(new_n21693_), .ZN(new_n21716_));
  AOI21_X1   g21524(.A1(new_n21716_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n21717_));
  AOI21_X1   g21525(.A1(new_n21717_), .A2(new_n21710_), .B(new_n21715_), .ZN(new_n21718_));
  OAI21_X1   g21526(.A1(new_n21718_), .A2(new_n21711_), .B(\asqrt[21] ), .ZN(new_n21719_));
  INV_X1     g21527(.I(new_n21719_), .ZN(new_n21720_));
  NOR2_X1    g21528(.A1(new_n20996_), .A2(new_n21004_), .ZN(new_n21721_));
  NOR3_X1    g21529(.A1(new_n21721_), .A2(new_n21404_), .A3(new_n21003_), .ZN(new_n21722_));
  NOR3_X1    g21530(.A1(new_n21620_), .A2(new_n21404_), .A3(new_n21721_), .ZN(new_n21723_));
  INV_X1     g21531(.I(new_n21723_), .ZN(new_n21724_));
  AOI22_X1   g21532(.A1(new_n21724_), .A2(new_n21003_), .B1(\asqrt[5] ), .B2(new_n21722_), .ZN(new_n21725_));
  NOR3_X1    g21533(.A1(new_n21718_), .A2(new_n21711_), .A3(\asqrt[21] ), .ZN(new_n21726_));
  NOR2_X1    g21534(.A1(new_n21726_), .A2(new_n21725_), .ZN(new_n21727_));
  OAI21_X1   g21535(.A1(new_n21727_), .A2(new_n21720_), .B(\asqrt[22] ), .ZN(new_n21728_));
  INV_X1     g21536(.I(new_n21011_), .ZN(new_n21729_));
  NOR3_X1    g21537(.A1(new_n21620_), .A2(new_n21006_), .A3(new_n21413_), .ZN(new_n21730_));
  INV_X1     g21538(.I(new_n21730_), .ZN(new_n21731_));
  NOR3_X1    g21539(.A1(new_n21413_), .A2(new_n21006_), .A3(new_n21729_), .ZN(new_n21732_));
  AOI22_X1   g21540(.A1(new_n21731_), .A2(new_n21729_), .B1(\asqrt[5] ), .B2(new_n21732_), .ZN(new_n21733_));
  INV_X1     g21541(.I(new_n21733_), .ZN(new_n21734_));
  NAND2_X1   g21542(.A1(new_n21719_), .A2(new_n11326_), .ZN(new_n21735_));
  OAI21_X1   g21543(.A1(new_n21727_), .A2(new_n21735_), .B(new_n21734_), .ZN(new_n21736_));
  AOI21_X1   g21544(.A1(new_n21736_), .A2(new_n21728_), .B(new_n10812_), .ZN(new_n21737_));
  NOR3_X1    g21545(.A1(new_n21016_), .A2(new_n21375_), .A3(new_n21025_), .ZN(new_n21738_));
  NOR3_X1    g21546(.A1(new_n21620_), .A2(new_n21016_), .A3(new_n21025_), .ZN(new_n21739_));
  INV_X1     g21547(.I(new_n21739_), .ZN(new_n21740_));
  AOI22_X1   g21548(.A1(new_n21740_), .A2(new_n21375_), .B1(\asqrt[5] ), .B2(new_n21738_), .ZN(new_n21741_));
  OAI21_X1   g21549(.A1(new_n21725_), .A2(new_n21726_), .B(new_n21719_), .ZN(new_n21742_));
  AOI21_X1   g21550(.A1(new_n21742_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n21743_));
  AOI21_X1   g21551(.A1(new_n21743_), .A2(new_n21736_), .B(new_n21741_), .ZN(new_n21744_));
  OAI21_X1   g21552(.A1(new_n21744_), .A2(new_n21737_), .B(\asqrt[24] ), .ZN(new_n21745_));
  INV_X1     g21553(.I(new_n21745_), .ZN(new_n21746_));
  NOR2_X1    g21554(.A1(new_n21026_), .A2(new_n21034_), .ZN(new_n21747_));
  NOR3_X1    g21555(.A1(new_n21620_), .A2(new_n21412_), .A3(new_n21747_), .ZN(new_n21748_));
  INV_X1     g21556(.I(new_n21748_), .ZN(new_n21749_));
  NOR3_X1    g21557(.A1(new_n21747_), .A2(new_n21412_), .A3(new_n21033_), .ZN(new_n21750_));
  AOI22_X1   g21558(.A1(new_n21749_), .A2(new_n21033_), .B1(\asqrt[5] ), .B2(new_n21750_), .ZN(new_n21751_));
  NOR3_X1    g21559(.A1(new_n21744_), .A2(new_n21737_), .A3(\asqrt[24] ), .ZN(new_n21752_));
  NOR2_X1    g21560(.A1(new_n21752_), .A2(new_n21751_), .ZN(new_n21753_));
  OAI21_X1   g21561(.A1(new_n21753_), .A2(new_n21746_), .B(\asqrt[25] ), .ZN(new_n21754_));
  INV_X1     g21562(.I(new_n21041_), .ZN(new_n21755_));
  NOR3_X1    g21563(.A1(new_n21421_), .A2(new_n21036_), .A3(new_n21755_), .ZN(new_n21756_));
  NOR3_X1    g21564(.A1(new_n21620_), .A2(new_n21036_), .A3(new_n21421_), .ZN(new_n21757_));
  INV_X1     g21565(.I(new_n21757_), .ZN(new_n21758_));
  AOI22_X1   g21566(.A1(new_n21758_), .A2(new_n21755_), .B1(\asqrt[5] ), .B2(new_n21756_), .ZN(new_n21759_));
  INV_X1     g21567(.I(new_n21759_), .ZN(new_n21760_));
  NAND2_X1   g21568(.A1(new_n21745_), .A2(new_n9846_), .ZN(new_n21761_));
  OAI21_X1   g21569(.A1(new_n21753_), .A2(new_n21761_), .B(new_n21760_), .ZN(new_n21762_));
  AOI21_X1   g21570(.A1(new_n21762_), .A2(new_n21754_), .B(new_n9317_), .ZN(new_n21763_));
  NOR3_X1    g21571(.A1(new_n21620_), .A2(new_n21046_), .A3(new_n21055_), .ZN(new_n21764_));
  INV_X1     g21572(.I(new_n21764_), .ZN(new_n21765_));
  NOR3_X1    g21573(.A1(new_n21046_), .A2(new_n21374_), .A3(new_n21055_), .ZN(new_n21766_));
  AOI22_X1   g21574(.A1(new_n21765_), .A2(new_n21374_), .B1(\asqrt[5] ), .B2(new_n21766_), .ZN(new_n21767_));
  OAI21_X1   g21575(.A1(new_n21751_), .A2(new_n21752_), .B(new_n21745_), .ZN(new_n21768_));
  AOI21_X1   g21576(.A1(new_n21768_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n21769_));
  AOI21_X1   g21577(.A1(new_n21769_), .A2(new_n21762_), .B(new_n21767_), .ZN(new_n21770_));
  OAI21_X1   g21578(.A1(new_n21770_), .A2(new_n21763_), .B(\asqrt[27] ), .ZN(new_n21771_));
  INV_X1     g21579(.I(new_n21771_), .ZN(new_n21772_));
  NOR2_X1    g21580(.A1(new_n21056_), .A2(new_n21064_), .ZN(new_n21773_));
  NOR3_X1    g21581(.A1(new_n21773_), .A2(new_n21420_), .A3(new_n21063_), .ZN(new_n21774_));
  NOR3_X1    g21582(.A1(new_n21620_), .A2(new_n21420_), .A3(new_n21773_), .ZN(new_n21775_));
  INV_X1     g21583(.I(new_n21775_), .ZN(new_n21776_));
  AOI22_X1   g21584(.A1(new_n21776_), .A2(new_n21063_), .B1(\asqrt[5] ), .B2(new_n21774_), .ZN(new_n21777_));
  NOR3_X1    g21585(.A1(new_n21770_), .A2(new_n21763_), .A3(\asqrt[27] ), .ZN(new_n21778_));
  NOR2_X1    g21586(.A1(new_n21778_), .A2(new_n21777_), .ZN(new_n21779_));
  OAI21_X1   g21587(.A1(new_n21779_), .A2(new_n21772_), .B(\asqrt[28] ), .ZN(new_n21780_));
  INV_X1     g21588(.I(new_n21071_), .ZN(new_n21781_));
  NOR3_X1    g21589(.A1(new_n21620_), .A2(new_n21066_), .A3(new_n21429_), .ZN(new_n21782_));
  INV_X1     g21590(.I(new_n21782_), .ZN(new_n21783_));
  NOR3_X1    g21591(.A1(new_n21429_), .A2(new_n21066_), .A3(new_n21781_), .ZN(new_n21784_));
  AOI22_X1   g21592(.A1(new_n21783_), .A2(new_n21781_), .B1(\asqrt[5] ), .B2(new_n21784_), .ZN(new_n21785_));
  INV_X1     g21593(.I(new_n21785_), .ZN(new_n21786_));
  NAND2_X1   g21594(.A1(new_n21771_), .A2(new_n8483_), .ZN(new_n21787_));
  OAI21_X1   g21595(.A1(new_n21779_), .A2(new_n21787_), .B(new_n21786_), .ZN(new_n21788_));
  AOI21_X1   g21596(.A1(new_n21788_), .A2(new_n21780_), .B(new_n8036_), .ZN(new_n21789_));
  NOR3_X1    g21597(.A1(new_n21076_), .A2(new_n21373_), .A3(new_n21085_), .ZN(new_n21790_));
  NOR3_X1    g21598(.A1(new_n21620_), .A2(new_n21076_), .A3(new_n21085_), .ZN(new_n21791_));
  INV_X1     g21599(.I(new_n21791_), .ZN(new_n21792_));
  AOI22_X1   g21600(.A1(new_n21792_), .A2(new_n21373_), .B1(\asqrt[5] ), .B2(new_n21790_), .ZN(new_n21793_));
  OAI21_X1   g21601(.A1(new_n21777_), .A2(new_n21778_), .B(new_n21771_), .ZN(new_n21794_));
  AOI21_X1   g21602(.A1(new_n21794_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n21795_));
  AOI21_X1   g21603(.A1(new_n21795_), .A2(new_n21788_), .B(new_n21793_), .ZN(new_n21796_));
  OAI21_X1   g21604(.A1(new_n21796_), .A2(new_n21789_), .B(\asqrt[30] ), .ZN(new_n21797_));
  INV_X1     g21605(.I(new_n21797_), .ZN(new_n21798_));
  NOR2_X1    g21606(.A1(new_n21086_), .A2(new_n21094_), .ZN(new_n21799_));
  NOR3_X1    g21607(.A1(new_n21620_), .A2(new_n21428_), .A3(new_n21799_), .ZN(new_n21800_));
  INV_X1     g21608(.I(new_n21800_), .ZN(new_n21801_));
  NOR3_X1    g21609(.A1(new_n21799_), .A2(new_n21428_), .A3(new_n21093_), .ZN(new_n21802_));
  AOI22_X1   g21610(.A1(new_n21801_), .A2(new_n21093_), .B1(\asqrt[5] ), .B2(new_n21802_), .ZN(new_n21803_));
  NOR3_X1    g21611(.A1(new_n21796_), .A2(new_n21789_), .A3(\asqrt[30] ), .ZN(new_n21804_));
  NOR2_X1    g21612(.A1(new_n21804_), .A2(new_n21803_), .ZN(new_n21805_));
  OAI21_X1   g21613(.A1(new_n21805_), .A2(new_n21798_), .B(\asqrt[31] ), .ZN(new_n21806_));
  INV_X1     g21614(.I(new_n21101_), .ZN(new_n21807_));
  NOR3_X1    g21615(.A1(new_n21437_), .A2(new_n21096_), .A3(new_n21807_), .ZN(new_n21808_));
  NOR3_X1    g21616(.A1(new_n21620_), .A2(new_n21096_), .A3(new_n21437_), .ZN(new_n21809_));
  INV_X1     g21617(.I(new_n21809_), .ZN(new_n21810_));
  AOI22_X1   g21618(.A1(new_n21810_), .A2(new_n21807_), .B1(\asqrt[5] ), .B2(new_n21808_), .ZN(new_n21811_));
  INV_X1     g21619(.I(new_n21811_), .ZN(new_n21812_));
  NAND2_X1   g21620(.A1(new_n21797_), .A2(new_n7229_), .ZN(new_n21813_));
  OAI21_X1   g21621(.A1(new_n21805_), .A2(new_n21813_), .B(new_n21812_), .ZN(new_n21814_));
  AOI21_X1   g21622(.A1(new_n21814_), .A2(new_n21806_), .B(new_n6824_), .ZN(new_n21815_));
  NOR3_X1    g21623(.A1(new_n21620_), .A2(new_n21106_), .A3(new_n21112_), .ZN(new_n21816_));
  INV_X1     g21624(.I(new_n21816_), .ZN(new_n21817_));
  NOR3_X1    g21625(.A1(new_n21106_), .A2(new_n21372_), .A3(new_n21112_), .ZN(new_n21818_));
  AOI22_X1   g21626(.A1(new_n21817_), .A2(new_n21372_), .B1(\asqrt[5] ), .B2(new_n21818_), .ZN(new_n21819_));
  OAI21_X1   g21627(.A1(new_n21803_), .A2(new_n21804_), .B(new_n21797_), .ZN(new_n21820_));
  AOI21_X1   g21628(.A1(new_n21820_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n21821_));
  AOI21_X1   g21629(.A1(new_n21821_), .A2(new_n21814_), .B(new_n21819_), .ZN(new_n21822_));
  OAI21_X1   g21630(.A1(new_n21822_), .A2(new_n21815_), .B(\asqrt[33] ), .ZN(new_n21823_));
  INV_X1     g21631(.I(new_n21823_), .ZN(new_n21824_));
  NOR2_X1    g21632(.A1(new_n21113_), .A2(new_n21121_), .ZN(new_n21825_));
  NOR3_X1    g21633(.A1(new_n21825_), .A2(new_n21436_), .A3(new_n21120_), .ZN(new_n21826_));
  NOR3_X1    g21634(.A1(new_n21620_), .A2(new_n21436_), .A3(new_n21825_), .ZN(new_n21827_));
  INV_X1     g21635(.I(new_n21827_), .ZN(new_n21828_));
  AOI22_X1   g21636(.A1(new_n21828_), .A2(new_n21120_), .B1(\asqrt[5] ), .B2(new_n21826_), .ZN(new_n21829_));
  NOR3_X1    g21637(.A1(new_n21822_), .A2(new_n21815_), .A3(\asqrt[33] ), .ZN(new_n21830_));
  NOR2_X1    g21638(.A1(new_n21830_), .A2(new_n21829_), .ZN(new_n21831_));
  OAI21_X1   g21639(.A1(new_n21831_), .A2(new_n21824_), .B(\asqrt[34] ), .ZN(new_n21832_));
  INV_X1     g21640(.I(new_n21128_), .ZN(new_n21833_));
  NOR3_X1    g21641(.A1(new_n21620_), .A2(new_n21123_), .A3(new_n21445_), .ZN(new_n21834_));
  INV_X1     g21642(.I(new_n21834_), .ZN(new_n21835_));
  NOR3_X1    g21643(.A1(new_n21445_), .A2(new_n21123_), .A3(new_n21833_), .ZN(new_n21836_));
  AOI22_X1   g21644(.A1(new_n21835_), .A2(new_n21833_), .B1(\asqrt[5] ), .B2(new_n21836_), .ZN(new_n21837_));
  INV_X1     g21645(.I(new_n21837_), .ZN(new_n21838_));
  NAND2_X1   g21646(.A1(new_n21823_), .A2(new_n6077_), .ZN(new_n21839_));
  OAI21_X1   g21647(.A1(new_n21831_), .A2(new_n21839_), .B(new_n21838_), .ZN(new_n21840_));
  AOI21_X1   g21648(.A1(new_n21840_), .A2(new_n21832_), .B(new_n5708_), .ZN(new_n21841_));
  NOR3_X1    g21649(.A1(new_n21133_), .A2(new_n21371_), .A3(new_n21139_), .ZN(new_n21842_));
  NOR3_X1    g21650(.A1(new_n21620_), .A2(new_n21133_), .A3(new_n21139_), .ZN(new_n21843_));
  INV_X1     g21651(.I(new_n21843_), .ZN(new_n21844_));
  AOI22_X1   g21652(.A1(new_n21844_), .A2(new_n21371_), .B1(\asqrt[5] ), .B2(new_n21842_), .ZN(new_n21845_));
  OAI21_X1   g21653(.A1(new_n21829_), .A2(new_n21830_), .B(new_n21823_), .ZN(new_n21846_));
  AOI21_X1   g21654(.A1(new_n21846_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n21847_));
  AOI21_X1   g21655(.A1(new_n21847_), .A2(new_n21840_), .B(new_n21845_), .ZN(new_n21848_));
  OAI21_X1   g21656(.A1(new_n21848_), .A2(new_n21841_), .B(\asqrt[36] ), .ZN(new_n21849_));
  INV_X1     g21657(.I(new_n21849_), .ZN(new_n21850_));
  NOR2_X1    g21658(.A1(new_n21140_), .A2(new_n21148_), .ZN(new_n21851_));
  NOR3_X1    g21659(.A1(new_n21620_), .A2(new_n21444_), .A3(new_n21851_), .ZN(new_n21852_));
  INV_X1     g21660(.I(new_n21852_), .ZN(new_n21853_));
  NOR3_X1    g21661(.A1(new_n21851_), .A2(new_n21444_), .A3(new_n21147_), .ZN(new_n21854_));
  AOI22_X1   g21662(.A1(new_n21853_), .A2(new_n21147_), .B1(\asqrt[5] ), .B2(new_n21854_), .ZN(new_n21855_));
  NOR3_X1    g21663(.A1(new_n21848_), .A2(new_n21841_), .A3(\asqrt[36] ), .ZN(new_n21856_));
  NOR2_X1    g21664(.A1(new_n21856_), .A2(new_n21855_), .ZN(new_n21857_));
  OAI21_X1   g21665(.A1(new_n21857_), .A2(new_n21850_), .B(\asqrt[37] ), .ZN(new_n21858_));
  INV_X1     g21666(.I(new_n21155_), .ZN(new_n21859_));
  NOR3_X1    g21667(.A1(new_n21453_), .A2(new_n21150_), .A3(new_n21859_), .ZN(new_n21860_));
  NOR3_X1    g21668(.A1(new_n21620_), .A2(new_n21150_), .A3(new_n21453_), .ZN(new_n21861_));
  INV_X1     g21669(.I(new_n21861_), .ZN(new_n21862_));
  AOI22_X1   g21670(.A1(new_n21862_), .A2(new_n21859_), .B1(\asqrt[5] ), .B2(new_n21860_), .ZN(new_n21863_));
  INV_X1     g21671(.I(new_n21863_), .ZN(new_n21864_));
  NAND2_X1   g21672(.A1(new_n21849_), .A2(new_n5024_), .ZN(new_n21865_));
  OAI21_X1   g21673(.A1(new_n21857_), .A2(new_n21865_), .B(new_n21864_), .ZN(new_n21866_));
  AOI21_X1   g21674(.A1(new_n21866_), .A2(new_n21858_), .B(new_n4696_), .ZN(new_n21867_));
  NOR3_X1    g21675(.A1(new_n21620_), .A2(new_n21160_), .A3(new_n21166_), .ZN(new_n21868_));
  INV_X1     g21676(.I(new_n21868_), .ZN(new_n21869_));
  NOR3_X1    g21677(.A1(new_n21160_), .A2(new_n21370_), .A3(new_n21166_), .ZN(new_n21870_));
  AOI22_X1   g21678(.A1(new_n21869_), .A2(new_n21370_), .B1(\asqrt[5] ), .B2(new_n21870_), .ZN(new_n21871_));
  OAI21_X1   g21679(.A1(new_n21855_), .A2(new_n21856_), .B(new_n21849_), .ZN(new_n21872_));
  AOI21_X1   g21680(.A1(new_n21872_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n21873_));
  AOI21_X1   g21681(.A1(new_n21873_), .A2(new_n21866_), .B(new_n21871_), .ZN(new_n21874_));
  OAI21_X1   g21682(.A1(new_n21874_), .A2(new_n21867_), .B(\asqrt[39] ), .ZN(new_n21875_));
  INV_X1     g21683(.I(new_n21875_), .ZN(new_n21876_));
  NOR2_X1    g21684(.A1(new_n21167_), .A2(new_n21175_), .ZN(new_n21877_));
  NOR3_X1    g21685(.A1(new_n21877_), .A2(new_n21452_), .A3(new_n21174_), .ZN(new_n21878_));
  NOR3_X1    g21686(.A1(new_n21620_), .A2(new_n21452_), .A3(new_n21877_), .ZN(new_n21879_));
  INV_X1     g21687(.I(new_n21879_), .ZN(new_n21880_));
  AOI22_X1   g21688(.A1(new_n21880_), .A2(new_n21174_), .B1(\asqrt[5] ), .B2(new_n21878_), .ZN(new_n21881_));
  NOR3_X1    g21689(.A1(new_n21874_), .A2(new_n21867_), .A3(\asqrt[39] ), .ZN(new_n21882_));
  NOR2_X1    g21690(.A1(new_n21882_), .A2(new_n21881_), .ZN(new_n21883_));
  OAI21_X1   g21691(.A1(new_n21883_), .A2(new_n21876_), .B(\asqrt[40] ), .ZN(new_n21884_));
  INV_X1     g21692(.I(new_n21181_), .ZN(new_n21885_));
  NOR3_X1    g21693(.A1(new_n21620_), .A2(new_n21177_), .A3(new_n21461_), .ZN(new_n21886_));
  INV_X1     g21694(.I(new_n21886_), .ZN(new_n21887_));
  NOR3_X1    g21695(.A1(new_n21461_), .A2(new_n21177_), .A3(new_n21885_), .ZN(new_n21888_));
  AOI22_X1   g21696(.A1(new_n21887_), .A2(new_n21885_), .B1(\asqrt[5] ), .B2(new_n21888_), .ZN(new_n21889_));
  INV_X1     g21697(.I(new_n21889_), .ZN(new_n21890_));
  NAND2_X1   g21698(.A1(new_n21875_), .A2(new_n4071_), .ZN(new_n21891_));
  OAI21_X1   g21699(.A1(new_n21883_), .A2(new_n21891_), .B(new_n21890_), .ZN(new_n21892_));
  AOI21_X1   g21700(.A1(new_n21892_), .A2(new_n21884_), .B(new_n3782_), .ZN(new_n21893_));
  NOR3_X1    g21701(.A1(new_n21186_), .A2(new_n21369_), .A3(new_n21192_), .ZN(new_n21894_));
  NOR3_X1    g21702(.A1(new_n21620_), .A2(new_n21186_), .A3(new_n21192_), .ZN(new_n21895_));
  INV_X1     g21703(.I(new_n21895_), .ZN(new_n21896_));
  AOI22_X1   g21704(.A1(new_n21896_), .A2(new_n21369_), .B1(\asqrt[5] ), .B2(new_n21894_), .ZN(new_n21897_));
  OAI21_X1   g21705(.A1(new_n21881_), .A2(new_n21882_), .B(new_n21875_), .ZN(new_n21898_));
  AOI21_X1   g21706(.A1(new_n21898_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n21899_));
  AOI21_X1   g21707(.A1(new_n21899_), .A2(new_n21892_), .B(new_n21897_), .ZN(new_n21900_));
  OAI21_X1   g21708(.A1(new_n21900_), .A2(new_n21893_), .B(\asqrt[42] ), .ZN(new_n21901_));
  INV_X1     g21709(.I(new_n21901_), .ZN(new_n21902_));
  NOR2_X1    g21710(.A1(new_n21193_), .A2(new_n21201_), .ZN(new_n21903_));
  NOR3_X1    g21711(.A1(new_n21620_), .A2(new_n21460_), .A3(new_n21903_), .ZN(new_n21904_));
  INV_X1     g21712(.I(new_n21904_), .ZN(new_n21905_));
  NOR3_X1    g21713(.A1(new_n21903_), .A2(new_n21460_), .A3(new_n21200_), .ZN(new_n21906_));
  AOI22_X1   g21714(.A1(new_n21905_), .A2(new_n21200_), .B1(\asqrt[5] ), .B2(new_n21906_), .ZN(new_n21907_));
  NOR3_X1    g21715(.A1(new_n21900_), .A2(new_n21893_), .A3(\asqrt[42] ), .ZN(new_n21908_));
  NOR2_X1    g21716(.A1(new_n21908_), .A2(new_n21907_), .ZN(new_n21909_));
  OAI21_X1   g21717(.A1(new_n21909_), .A2(new_n21902_), .B(\asqrt[43] ), .ZN(new_n21910_));
  INV_X1     g21718(.I(new_n21207_), .ZN(new_n21911_));
  NOR3_X1    g21719(.A1(new_n21469_), .A2(new_n21203_), .A3(new_n21911_), .ZN(new_n21912_));
  NOR3_X1    g21720(.A1(new_n21620_), .A2(new_n21203_), .A3(new_n21469_), .ZN(new_n21913_));
  INV_X1     g21721(.I(new_n21913_), .ZN(new_n21914_));
  AOI22_X1   g21722(.A1(new_n21914_), .A2(new_n21911_), .B1(\asqrt[5] ), .B2(new_n21912_), .ZN(new_n21915_));
  INV_X1     g21723(.I(new_n21915_), .ZN(new_n21916_));
  NAND2_X1   g21724(.A1(new_n21901_), .A2(new_n3218_), .ZN(new_n21917_));
  OAI21_X1   g21725(.A1(new_n21909_), .A2(new_n21917_), .B(new_n21916_), .ZN(new_n21918_));
  AOI21_X1   g21726(.A1(new_n21918_), .A2(new_n21910_), .B(new_n2954_), .ZN(new_n21919_));
  NOR3_X1    g21727(.A1(new_n21620_), .A2(new_n21212_), .A3(new_n21220_), .ZN(new_n21920_));
  INV_X1     g21728(.I(new_n21920_), .ZN(new_n21921_));
  NOR3_X1    g21729(.A1(new_n21212_), .A2(new_n21368_), .A3(new_n21220_), .ZN(new_n21922_));
  AOI22_X1   g21730(.A1(new_n21921_), .A2(new_n21368_), .B1(\asqrt[5] ), .B2(new_n21922_), .ZN(new_n21923_));
  OAI21_X1   g21731(.A1(new_n21907_), .A2(new_n21908_), .B(new_n21901_), .ZN(new_n21924_));
  AOI21_X1   g21732(.A1(new_n21924_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n21925_));
  AOI21_X1   g21733(.A1(new_n21925_), .A2(new_n21918_), .B(new_n21923_), .ZN(new_n21926_));
  OAI21_X1   g21734(.A1(new_n21926_), .A2(new_n21919_), .B(\asqrt[45] ), .ZN(new_n21927_));
  INV_X1     g21735(.I(new_n21927_), .ZN(new_n21928_));
  NOR2_X1    g21736(.A1(new_n21221_), .A2(new_n21228_), .ZN(new_n21929_));
  NOR3_X1    g21737(.A1(new_n21929_), .A2(new_n21468_), .A3(new_n21227_), .ZN(new_n21930_));
  NOR3_X1    g21738(.A1(new_n21620_), .A2(new_n21468_), .A3(new_n21929_), .ZN(new_n21931_));
  INV_X1     g21739(.I(new_n21931_), .ZN(new_n21932_));
  AOI22_X1   g21740(.A1(new_n21932_), .A2(new_n21227_), .B1(\asqrt[5] ), .B2(new_n21930_), .ZN(new_n21933_));
  NOR3_X1    g21741(.A1(new_n21926_), .A2(new_n21919_), .A3(\asqrt[45] ), .ZN(new_n21934_));
  NOR2_X1    g21742(.A1(new_n21934_), .A2(new_n21933_), .ZN(new_n21935_));
  OAI21_X1   g21743(.A1(new_n21935_), .A2(new_n21928_), .B(\asqrt[46] ), .ZN(new_n21936_));
  INV_X1     g21744(.I(new_n21236_), .ZN(new_n21937_));
  NOR3_X1    g21745(.A1(new_n21620_), .A2(new_n21230_), .A3(new_n21477_), .ZN(new_n21938_));
  INV_X1     g21746(.I(new_n21938_), .ZN(new_n21939_));
  NOR3_X1    g21747(.A1(new_n21477_), .A2(new_n21230_), .A3(new_n21937_), .ZN(new_n21940_));
  AOI22_X1   g21748(.A1(new_n21939_), .A2(new_n21937_), .B1(\asqrt[5] ), .B2(new_n21940_), .ZN(new_n21941_));
  INV_X1     g21749(.I(new_n21941_), .ZN(new_n21942_));
  NAND2_X1   g21750(.A1(new_n21927_), .A2(new_n2465_), .ZN(new_n21943_));
  OAI21_X1   g21751(.A1(new_n21935_), .A2(new_n21943_), .B(new_n21942_), .ZN(new_n21944_));
  AOI21_X1   g21752(.A1(new_n21944_), .A2(new_n21936_), .B(new_n2229_), .ZN(new_n21945_));
  NOR3_X1    g21753(.A1(new_n21241_), .A2(new_n21367_), .A3(new_n21250_), .ZN(new_n21946_));
  NOR3_X1    g21754(.A1(new_n21620_), .A2(new_n21241_), .A3(new_n21250_), .ZN(new_n21947_));
  INV_X1     g21755(.I(new_n21947_), .ZN(new_n21948_));
  AOI22_X1   g21756(.A1(new_n21948_), .A2(new_n21367_), .B1(\asqrt[5] ), .B2(new_n21946_), .ZN(new_n21949_));
  OAI21_X1   g21757(.A1(new_n21933_), .A2(new_n21934_), .B(new_n21927_), .ZN(new_n21950_));
  AOI21_X1   g21758(.A1(new_n21950_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n21951_));
  AOI21_X1   g21759(.A1(new_n21951_), .A2(new_n21944_), .B(new_n21949_), .ZN(new_n21952_));
  OAI21_X1   g21760(.A1(new_n21952_), .A2(new_n21945_), .B(\asqrt[48] ), .ZN(new_n21953_));
  INV_X1     g21761(.I(new_n21953_), .ZN(new_n21954_));
  NOR2_X1    g21762(.A1(new_n21251_), .A2(new_n21258_), .ZN(new_n21955_));
  NOR3_X1    g21763(.A1(new_n21620_), .A2(new_n21476_), .A3(new_n21955_), .ZN(new_n21956_));
  INV_X1     g21764(.I(new_n21956_), .ZN(new_n21957_));
  NOR3_X1    g21765(.A1(new_n21955_), .A2(new_n21476_), .A3(new_n21257_), .ZN(new_n21958_));
  AOI22_X1   g21766(.A1(new_n21957_), .A2(new_n21257_), .B1(\asqrt[5] ), .B2(new_n21958_), .ZN(new_n21959_));
  NOR3_X1    g21767(.A1(new_n21952_), .A2(new_n21945_), .A3(\asqrt[48] ), .ZN(new_n21960_));
  NOR2_X1    g21768(.A1(new_n21960_), .A2(new_n21959_), .ZN(new_n21961_));
  OAI21_X1   g21769(.A1(new_n21961_), .A2(new_n21954_), .B(\asqrt[49] ), .ZN(new_n21962_));
  INV_X1     g21770(.I(new_n21266_), .ZN(new_n21963_));
  NOR3_X1    g21771(.A1(new_n21485_), .A2(new_n21260_), .A3(new_n21963_), .ZN(new_n21964_));
  NOR3_X1    g21772(.A1(new_n21620_), .A2(new_n21260_), .A3(new_n21485_), .ZN(new_n21965_));
  INV_X1     g21773(.I(new_n21965_), .ZN(new_n21966_));
  AOI22_X1   g21774(.A1(new_n21966_), .A2(new_n21963_), .B1(\asqrt[5] ), .B2(new_n21964_), .ZN(new_n21967_));
  INV_X1     g21775(.I(new_n21967_), .ZN(new_n21968_));
  NAND2_X1   g21776(.A1(new_n21953_), .A2(new_n1806_), .ZN(new_n21969_));
  OAI21_X1   g21777(.A1(new_n21961_), .A2(new_n21969_), .B(new_n21968_), .ZN(new_n21970_));
  AOI21_X1   g21778(.A1(new_n21970_), .A2(new_n21962_), .B(new_n1612_), .ZN(new_n21971_));
  NOR3_X1    g21779(.A1(new_n21620_), .A2(new_n21271_), .A3(new_n21280_), .ZN(new_n21972_));
  INV_X1     g21780(.I(new_n21972_), .ZN(new_n21973_));
  NOR3_X1    g21781(.A1(new_n21271_), .A2(new_n21366_), .A3(new_n21280_), .ZN(new_n21974_));
  AOI22_X1   g21782(.A1(new_n21973_), .A2(new_n21366_), .B1(\asqrt[5] ), .B2(new_n21974_), .ZN(new_n21975_));
  OAI21_X1   g21783(.A1(new_n21959_), .A2(new_n21960_), .B(new_n21953_), .ZN(new_n21976_));
  AOI21_X1   g21784(.A1(new_n21976_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n21977_));
  AOI21_X1   g21785(.A1(new_n21977_), .A2(new_n21970_), .B(new_n21975_), .ZN(new_n21978_));
  OAI21_X1   g21786(.A1(new_n21978_), .A2(new_n21971_), .B(\asqrt[51] ), .ZN(new_n21979_));
  INV_X1     g21787(.I(new_n21979_), .ZN(new_n21980_));
  NOR2_X1    g21788(.A1(new_n21281_), .A2(new_n21288_), .ZN(new_n21981_));
  NOR3_X1    g21789(.A1(new_n21981_), .A2(new_n21484_), .A3(new_n21287_), .ZN(new_n21982_));
  NOR3_X1    g21790(.A1(new_n21620_), .A2(new_n21484_), .A3(new_n21981_), .ZN(new_n21983_));
  INV_X1     g21791(.I(new_n21983_), .ZN(new_n21984_));
  AOI22_X1   g21792(.A1(new_n21984_), .A2(new_n21287_), .B1(\asqrt[5] ), .B2(new_n21982_), .ZN(new_n21985_));
  NOR3_X1    g21793(.A1(new_n21978_), .A2(new_n21971_), .A3(\asqrt[51] ), .ZN(new_n21986_));
  NOR2_X1    g21794(.A1(new_n21986_), .A2(new_n21985_), .ZN(new_n21987_));
  OAI21_X1   g21795(.A1(new_n21987_), .A2(new_n21980_), .B(\asqrt[52] ), .ZN(new_n21988_));
  INV_X1     g21796(.I(new_n21296_), .ZN(new_n21989_));
  NAND2_X1   g21797(.A1(new_n21298_), .A2(new_n21289_), .ZN(new_n21990_));
  INV_X1     g21798(.I(new_n21990_), .ZN(new_n21991_));
  NOR3_X1    g21799(.A1(new_n21620_), .A2(new_n21290_), .A3(new_n21991_), .ZN(new_n21992_));
  INV_X1     g21800(.I(new_n21992_), .ZN(new_n21993_));
  NOR3_X1    g21801(.A1(new_n21991_), .A2(new_n21290_), .A3(new_n21989_), .ZN(new_n21994_));
  AOI22_X1   g21802(.A1(new_n21993_), .A2(new_n21989_), .B1(\asqrt[5] ), .B2(new_n21994_), .ZN(new_n21995_));
  INV_X1     g21803(.I(new_n21995_), .ZN(new_n21996_));
  NAND2_X1   g21804(.A1(new_n21979_), .A2(new_n1256_), .ZN(new_n21997_));
  OAI21_X1   g21805(.A1(new_n21987_), .A2(new_n21997_), .B(new_n21996_), .ZN(new_n21998_));
  AOI21_X1   g21806(.A1(new_n21998_), .A2(new_n21988_), .B(new_n1103_), .ZN(new_n21999_));
  NOR3_X1    g21807(.A1(new_n21301_), .A2(new_n21365_), .A3(new_n21310_), .ZN(new_n22000_));
  NOR3_X1    g21808(.A1(new_n21620_), .A2(new_n21301_), .A3(new_n21310_), .ZN(new_n22001_));
  INV_X1     g21809(.I(new_n22001_), .ZN(new_n22002_));
  AOI22_X1   g21810(.A1(new_n22002_), .A2(new_n21365_), .B1(\asqrt[5] ), .B2(new_n22000_), .ZN(new_n22003_));
  OAI21_X1   g21811(.A1(new_n21985_), .A2(new_n21986_), .B(new_n21979_), .ZN(new_n22004_));
  AOI21_X1   g21812(.A1(new_n22004_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n22005_));
  AOI21_X1   g21813(.A1(new_n22005_), .A2(new_n21998_), .B(new_n22003_), .ZN(new_n22006_));
  OAI21_X1   g21814(.A1(new_n22006_), .A2(new_n21999_), .B(\asqrt[54] ), .ZN(new_n22007_));
  INV_X1     g21815(.I(new_n22007_), .ZN(new_n22008_));
  INV_X1     g21816(.I(new_n21312_), .ZN(new_n22009_));
  INV_X1     g21817(.I(new_n21492_), .ZN(new_n22010_));
  NOR3_X1    g21818(.A1(new_n21620_), .A2(new_n22009_), .A3(new_n22010_), .ZN(new_n22011_));
  INV_X1     g21819(.I(new_n22011_), .ZN(new_n22012_));
  NOR3_X1    g21820(.A1(new_n22009_), .A2(new_n22010_), .A3(new_n21317_), .ZN(new_n22013_));
  AOI22_X1   g21821(.A1(new_n22012_), .A2(new_n21317_), .B1(\asqrt[5] ), .B2(new_n22013_), .ZN(new_n22014_));
  NOR3_X1    g21822(.A1(new_n22006_), .A2(new_n21999_), .A3(\asqrt[54] ), .ZN(new_n22015_));
  NOR2_X1    g21823(.A1(new_n22015_), .A2(new_n22014_), .ZN(new_n22016_));
  OAI21_X1   g21824(.A1(new_n22016_), .A2(new_n22008_), .B(\asqrt[55] ), .ZN(new_n22017_));
  INV_X1     g21825(.I(new_n21326_), .ZN(new_n22018_));
  INV_X1     g21826(.I(new_n21319_), .ZN(new_n22019_));
  INV_X1     g21827(.I(new_n21328_), .ZN(new_n22020_));
  OAI21_X1   g21828(.A1(new_n22020_), .A2(new_n22019_), .B(new_n21326_), .ZN(new_n22021_));
  NOR2_X1    g21829(.A1(new_n22021_), .A2(new_n21320_), .ZN(new_n22022_));
  NOR2_X1    g21830(.A1(new_n22020_), .A2(new_n22019_), .ZN(new_n22023_));
  NOR3_X1    g21831(.A1(new_n21620_), .A2(new_n21320_), .A3(new_n22023_), .ZN(new_n22024_));
  INV_X1     g21832(.I(new_n22024_), .ZN(new_n22025_));
  AOI22_X1   g21833(.A1(new_n22025_), .A2(new_n22018_), .B1(\asqrt[5] ), .B2(new_n22022_), .ZN(new_n22026_));
  INV_X1     g21834(.I(new_n22026_), .ZN(new_n22027_));
  NAND2_X1   g21835(.A1(new_n22007_), .A2(new_n823_), .ZN(new_n22028_));
  OAI21_X1   g21836(.A1(new_n22016_), .A2(new_n22028_), .B(new_n22027_), .ZN(new_n22029_));
  AOI21_X1   g21837(.A1(new_n22029_), .A2(new_n22017_), .B(new_n703_), .ZN(new_n22030_));
  NOR3_X1    g21838(.A1(new_n21620_), .A2(new_n21331_), .A3(new_n21337_), .ZN(new_n22031_));
  INV_X1     g21839(.I(new_n22031_), .ZN(new_n22032_));
  NOR3_X1    g21840(.A1(new_n21331_), .A2(new_n21364_), .A3(new_n21337_), .ZN(new_n22033_));
  AOI22_X1   g21841(.A1(new_n22032_), .A2(new_n21364_), .B1(\asqrt[5] ), .B2(new_n22033_), .ZN(new_n22034_));
  OAI21_X1   g21842(.A1(new_n22014_), .A2(new_n22015_), .B(new_n22007_), .ZN(new_n22035_));
  AOI21_X1   g21843(.A1(new_n22035_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n22036_));
  AOI21_X1   g21844(.A1(new_n22036_), .A2(new_n22029_), .B(new_n22034_), .ZN(new_n22037_));
  OAI21_X1   g21845(.A1(new_n22037_), .A2(new_n22030_), .B(\asqrt[57] ), .ZN(new_n22038_));
  INV_X1     g21846(.I(new_n22038_), .ZN(new_n22039_));
  INV_X1     g21847(.I(new_n21339_), .ZN(new_n22040_));
  INV_X1     g21848(.I(new_n21496_), .ZN(new_n22041_));
  NOR3_X1    g21849(.A1(new_n22040_), .A2(new_n22041_), .A3(new_n21344_), .ZN(new_n22042_));
  NOR3_X1    g21850(.A1(new_n21620_), .A2(new_n22040_), .A3(new_n22041_), .ZN(new_n22043_));
  INV_X1     g21851(.I(new_n22043_), .ZN(new_n22044_));
  AOI22_X1   g21852(.A1(new_n22044_), .A2(new_n21344_), .B1(\asqrt[5] ), .B2(new_n22042_), .ZN(new_n22045_));
  NOR3_X1    g21853(.A1(new_n22037_), .A2(new_n22030_), .A3(\asqrt[57] ), .ZN(new_n22046_));
  NOR2_X1    g21854(.A1(new_n22046_), .A2(new_n22045_), .ZN(new_n22047_));
  OAI21_X1   g21855(.A1(new_n22047_), .A2(new_n22039_), .B(\asqrt[58] ), .ZN(new_n22048_));
  INV_X1     g21856(.I(new_n21353_), .ZN(new_n22049_));
  INV_X1     g21857(.I(new_n21346_), .ZN(new_n22050_));
  INV_X1     g21858(.I(new_n21355_), .ZN(new_n22051_));
  NOR2_X1    g21859(.A1(new_n22051_), .A2(new_n22050_), .ZN(new_n22052_));
  NOR3_X1    g21860(.A1(new_n21620_), .A2(new_n21347_), .A3(new_n22052_), .ZN(new_n22053_));
  INV_X1     g21861(.I(new_n22053_), .ZN(new_n22054_));
  NOR3_X1    g21862(.A1(new_n22052_), .A2(new_n21347_), .A3(new_n22049_), .ZN(new_n22055_));
  AOI22_X1   g21863(.A1(new_n22054_), .A2(new_n22049_), .B1(\asqrt[5] ), .B2(new_n22055_), .ZN(new_n22056_));
  INV_X1     g21864(.I(new_n22056_), .ZN(new_n22057_));
  NAND2_X1   g21865(.A1(new_n22038_), .A2(new_n436_), .ZN(new_n22058_));
  OAI21_X1   g21866(.A1(new_n22047_), .A2(new_n22058_), .B(new_n22057_), .ZN(new_n22059_));
  AOI21_X1   g21867(.A1(new_n22059_), .A2(new_n22048_), .B(new_n327_), .ZN(new_n22060_));
  NOR3_X1    g21868(.A1(new_n21516_), .A2(new_n21363_), .A3(new_n21517_), .ZN(new_n22061_));
  NOR3_X1    g21869(.A1(new_n21620_), .A2(new_n21516_), .A3(new_n21517_), .ZN(new_n22062_));
  INV_X1     g21870(.I(new_n22062_), .ZN(new_n22063_));
  AOI22_X1   g21871(.A1(new_n22063_), .A2(new_n21363_), .B1(\asqrt[5] ), .B2(new_n22061_), .ZN(new_n22064_));
  OAI21_X1   g21872(.A1(new_n22045_), .A2(new_n22046_), .B(new_n22038_), .ZN(new_n22065_));
  AOI21_X1   g21873(.A1(new_n22065_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n22066_));
  AOI21_X1   g21874(.A1(new_n22066_), .A2(new_n22059_), .B(new_n22064_), .ZN(new_n22067_));
  OAI21_X1   g21875(.A1(new_n22067_), .A2(new_n22060_), .B(\asqrt[60] ), .ZN(new_n22068_));
  INV_X1     g21876(.I(new_n22068_), .ZN(new_n22069_));
  INV_X1     g21877(.I(new_n21570_), .ZN(new_n22070_));
  NOR3_X1    g21878(.A1(new_n21620_), .A2(new_n21500_), .A3(new_n22070_), .ZN(new_n22071_));
  INV_X1     g21879(.I(new_n22071_), .ZN(new_n22072_));
  NOR3_X1    g21880(.A1(new_n22070_), .A2(new_n21500_), .A3(new_n21528_), .ZN(new_n22073_));
  AOI22_X1   g21881(.A1(new_n22072_), .A2(new_n21528_), .B1(\asqrt[5] ), .B2(new_n22073_), .ZN(new_n22074_));
  NOR3_X1    g21882(.A1(new_n22067_), .A2(new_n22060_), .A3(\asqrt[60] ), .ZN(new_n22075_));
  NOR2_X1    g21883(.A1(new_n22075_), .A2(new_n22074_), .ZN(new_n22076_));
  OAI21_X1   g21884(.A1(new_n22076_), .A2(new_n22069_), .B(\asqrt[61] ), .ZN(new_n22077_));
  NAND2_X1   g21885(.A1(new_n21540_), .A2(new_n21529_), .ZN(new_n22078_));
  AND3_X2    g21886(.A1(new_n21508_), .A2(new_n21514_), .A3(new_n22078_), .Z(new_n22079_));
  NAND3_X1   g21887(.A1(\asqrt[5] ), .A2(new_n21508_), .A3(new_n22078_), .ZN(new_n22080_));
  AOI22_X1   g21888(.A1(new_n22080_), .A2(new_n21515_), .B1(\asqrt[5] ), .B2(new_n22079_), .ZN(new_n22081_));
  INV_X1     g21889(.I(new_n22081_), .ZN(new_n22082_));
  NAND2_X1   g21890(.A1(new_n22068_), .A2(new_n218_), .ZN(new_n22083_));
  OAI21_X1   g21891(.A1(new_n22076_), .A2(new_n22083_), .B(new_n22082_), .ZN(new_n22084_));
  AOI21_X1   g21892(.A1(new_n22084_), .A2(new_n22077_), .B(new_n207_), .ZN(new_n22085_));
  NOR3_X1    g21893(.A1(new_n21620_), .A2(new_n21522_), .A3(new_n21553_), .ZN(new_n22086_));
  INV_X1     g21894(.I(new_n22086_), .ZN(new_n22087_));
  NOR3_X1    g21895(.A1(new_n21522_), .A2(new_n21569_), .A3(new_n21553_), .ZN(new_n22088_));
  AOI22_X1   g21896(.A1(new_n22087_), .A2(new_n21569_), .B1(\asqrt[5] ), .B2(new_n22088_), .ZN(new_n22089_));
  OAI21_X1   g21897(.A1(new_n22074_), .A2(new_n22075_), .B(new_n22068_), .ZN(new_n22090_));
  AOI21_X1   g21898(.A1(new_n22090_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n22091_));
  AOI21_X1   g21899(.A1(new_n22091_), .A2(new_n22084_), .B(new_n22089_), .ZN(new_n22092_));
  INV_X1     g21900(.I(new_n21533_), .ZN(new_n22093_));
  INV_X1     g21901(.I(new_n21582_), .ZN(new_n22094_));
  NOR3_X1    g21902(.A1(new_n22093_), .A2(new_n22094_), .A3(new_n21538_), .ZN(new_n22095_));
  NOR3_X1    g21903(.A1(new_n21620_), .A2(new_n22093_), .A3(new_n22094_), .ZN(new_n22096_));
  INV_X1     g21904(.I(new_n22096_), .ZN(new_n22097_));
  AOI22_X1   g21905(.A1(new_n22097_), .A2(new_n21538_), .B1(\asqrt[5] ), .B2(new_n22095_), .ZN(new_n22098_));
  INV_X1     g21906(.I(new_n22098_), .ZN(new_n22099_));
  NOR2_X1    g21907(.A1(new_n21583_), .A2(new_n21576_), .ZN(new_n22100_));
  NAND2_X1   g21908(.A1(\asqrt[5] ), .A2(new_n22100_), .ZN(new_n22101_));
  AND3_X2    g21909(.A1(new_n22099_), .A2(new_n21596_), .A3(new_n22101_), .Z(new_n22102_));
  OAI21_X1   g21910(.A1(new_n22092_), .A2(new_n22085_), .B(new_n22102_), .ZN(new_n22103_));
  NAND2_X1   g21911(.A1(new_n22103_), .A2(new_n193_), .ZN(new_n22104_));
  INV_X1     g21912(.I(new_n22074_), .ZN(new_n22105_));
  INV_X1     g21913(.I(new_n22045_), .ZN(new_n22106_));
  INV_X1     g21914(.I(new_n22014_), .ZN(new_n22107_));
  INV_X1     g21915(.I(new_n21985_), .ZN(new_n22108_));
  INV_X1     g21916(.I(new_n21959_), .ZN(new_n22109_));
  INV_X1     g21917(.I(new_n21933_), .ZN(new_n22110_));
  INV_X1     g21918(.I(new_n21907_), .ZN(new_n22111_));
  INV_X1     g21919(.I(new_n21881_), .ZN(new_n22112_));
  INV_X1     g21920(.I(new_n21855_), .ZN(new_n22113_));
  INV_X1     g21921(.I(new_n21829_), .ZN(new_n22114_));
  INV_X1     g21922(.I(new_n21803_), .ZN(new_n22115_));
  INV_X1     g21923(.I(new_n21777_), .ZN(new_n22116_));
  INV_X1     g21924(.I(new_n21751_), .ZN(new_n22117_));
  INV_X1     g21925(.I(new_n21725_), .ZN(new_n22118_));
  INV_X1     g21926(.I(new_n21699_), .ZN(new_n22119_));
  INV_X1     g21927(.I(new_n21673_), .ZN(new_n22120_));
  INV_X1     g21928(.I(new_n21647_), .ZN(new_n22121_));
  NAND2_X1   g21929(.A1(new_n21579_), .A2(new_n21587_), .ZN(new_n22122_));
  OAI21_X1   g21930(.A1(new_n21568_), .A2(new_n21578_), .B(new_n21581_), .ZN(new_n22123_));
  NAND2_X1   g21931(.A1(new_n22123_), .A2(\a[11] ), .ZN(new_n22124_));
  NAND3_X1   g21932(.A1(new_n22122_), .A2(new_n22124_), .A3(new_n21595_), .ZN(new_n22125_));
  AOI21_X1   g21933(.A1(new_n22125_), .A2(new_n21609_), .B(new_n20262_), .ZN(new_n22126_));
  OAI21_X1   g21934(.A1(new_n21600_), .A2(new_n21590_), .B(\a[12] ), .ZN(new_n22127_));
  NAND3_X1   g21935(.A1(new_n21597_), .A2(new_n21595_), .A3(new_n20807_), .ZN(new_n22128_));
  NAND2_X1   g21936(.A1(new_n21579_), .A2(new_n21565_), .ZN(new_n22129_));
  AOI21_X1   g21937(.A1(new_n22129_), .A2(\asqrt[6] ), .B(\asqrt[7] ), .ZN(new_n22130_));
  AOI22_X1   g21938(.A1(new_n22125_), .A2(new_n22130_), .B1(new_n22127_), .B2(new_n22128_), .ZN(new_n22131_));
  OAI21_X1   g21939(.A1(new_n22131_), .A2(new_n22126_), .B(\asqrt[8] ), .ZN(new_n22132_));
  NAND2_X1   g21940(.A1(new_n22132_), .A2(new_n18792_), .ZN(new_n22133_));
  OAI21_X1   g21941(.A1(new_n22133_), .A2(new_n21614_), .B(new_n21622_), .ZN(new_n22134_));
  AOI21_X1   g21942(.A1(new_n22134_), .A2(new_n21615_), .B(new_n18275_), .ZN(new_n22135_));
  INV_X1     g21943(.I(new_n21608_), .ZN(new_n22136_));
  AOI21_X1   g21944(.A1(\a[11] ), .A2(new_n22123_), .B(new_n21590_), .ZN(new_n22137_));
  AOI21_X1   g21945(.A1(new_n22137_), .A2(new_n22122_), .B(new_n21580_), .ZN(new_n22138_));
  OAI21_X1   g21946(.A1(new_n22138_), .A2(new_n20262_), .B(new_n19573_), .ZN(new_n22139_));
  OAI21_X1   g21947(.A1(new_n22139_), .A2(new_n22131_), .B(new_n22136_), .ZN(new_n22140_));
  NAND2_X1   g21948(.A1(new_n22140_), .A2(new_n22132_), .ZN(new_n22141_));
  AOI21_X1   g21949(.A1(new_n22141_), .A2(\asqrt[9] ), .B(\asqrt[10] ), .ZN(new_n22142_));
  AOI21_X1   g21950(.A1(new_n22142_), .A2(new_n22134_), .B(new_n21630_), .ZN(new_n22143_));
  OAI21_X1   g21951(.A1(new_n22143_), .A2(new_n22135_), .B(\asqrt[11] ), .ZN(new_n22144_));
  NAND2_X1   g21952(.A1(new_n22144_), .A2(new_n16881_), .ZN(new_n22145_));
  OAI21_X1   g21953(.A1(new_n22145_), .A2(new_n21641_), .B(new_n22121_), .ZN(new_n22146_));
  NAND3_X1   g21954(.A1(new_n22146_), .A2(new_n16389_), .A3(new_n21642_), .ZN(new_n22147_));
  AOI22_X1   g21955(.A1(new_n22147_), .A2(new_n21656_), .B1(new_n21664_), .B2(\asqrt[13] ), .ZN(new_n22148_));
  OAI21_X1   g21956(.A1(new_n22148_), .A2(new_n15770_), .B(new_n15067_), .ZN(new_n22149_));
  OAI21_X1   g21957(.A1(new_n22149_), .A2(new_n21666_), .B(new_n22120_), .ZN(new_n22150_));
  AOI21_X1   g21958(.A1(new_n22150_), .A2(new_n21667_), .B(new_n14601_), .ZN(new_n22151_));
  AOI21_X1   g21959(.A1(new_n22146_), .A2(new_n21642_), .B(new_n16389_), .ZN(new_n22152_));
  NOR3_X1    g21960(.A1(new_n22143_), .A2(new_n22135_), .A3(\asqrt[11] ), .ZN(new_n22153_));
  OAI21_X1   g21961(.A1(new_n21638_), .A2(new_n22153_), .B(new_n22144_), .ZN(new_n22154_));
  AOI21_X1   g21962(.A1(new_n22154_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n22155_));
  AOI21_X1   g21963(.A1(new_n22155_), .A2(new_n22146_), .B(new_n21655_), .ZN(new_n22156_));
  NOR3_X1    g21964(.A1(new_n22156_), .A2(\asqrt[14] ), .A3(new_n22152_), .ZN(new_n22157_));
  OAI22_X1   g21965(.A1(new_n22157_), .A2(new_n21663_), .B1(new_n22148_), .B2(new_n15770_), .ZN(new_n22158_));
  AOI21_X1   g21966(.A1(new_n22158_), .A2(\asqrt[15] ), .B(\asqrt[16] ), .ZN(new_n22159_));
  AOI21_X1   g21967(.A1(new_n22159_), .A2(new_n22150_), .B(new_n21681_), .ZN(new_n22160_));
  OAI21_X1   g21968(.A1(new_n22160_), .A2(new_n22151_), .B(\asqrt[17] ), .ZN(new_n22161_));
  NAND2_X1   g21969(.A1(new_n22161_), .A2(new_n13353_), .ZN(new_n22162_));
  OAI21_X1   g21970(.A1(new_n22162_), .A2(new_n21692_), .B(new_n22119_), .ZN(new_n22163_));
  AOI21_X1   g21971(.A1(new_n22163_), .A2(new_n21693_), .B(new_n12913_), .ZN(new_n22164_));
  NOR3_X1    g21972(.A1(new_n22160_), .A2(\asqrt[17] ), .A3(new_n22151_), .ZN(new_n22165_));
  OAI21_X1   g21973(.A1(new_n21689_), .A2(new_n22165_), .B(new_n22161_), .ZN(new_n22166_));
  AOI21_X1   g21974(.A1(new_n22166_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n22167_));
  AOI21_X1   g21975(.A1(new_n22167_), .A2(new_n22163_), .B(new_n21707_), .ZN(new_n22168_));
  OAI21_X1   g21976(.A1(new_n22168_), .A2(new_n22164_), .B(\asqrt[20] ), .ZN(new_n22169_));
  NAND2_X1   g21977(.A1(new_n22169_), .A2(new_n11736_), .ZN(new_n22170_));
  OAI21_X1   g21978(.A1(new_n22170_), .A2(new_n21718_), .B(new_n22118_), .ZN(new_n22171_));
  AOI21_X1   g21979(.A1(new_n22171_), .A2(new_n21719_), .B(new_n11326_), .ZN(new_n22172_));
  NOR3_X1    g21980(.A1(new_n22168_), .A2(\asqrt[20] ), .A3(new_n22164_), .ZN(new_n22173_));
  OAI21_X1   g21981(.A1(new_n21715_), .A2(new_n22173_), .B(new_n22169_), .ZN(new_n22174_));
  AOI21_X1   g21982(.A1(new_n22174_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n22175_));
  AOI21_X1   g21983(.A1(new_n22175_), .A2(new_n22171_), .B(new_n21733_), .ZN(new_n22176_));
  OAI21_X1   g21984(.A1(new_n22176_), .A2(new_n22172_), .B(\asqrt[23] ), .ZN(new_n22177_));
  NAND2_X1   g21985(.A1(new_n22177_), .A2(new_n10221_), .ZN(new_n22178_));
  OAI21_X1   g21986(.A1(new_n22178_), .A2(new_n21744_), .B(new_n22117_), .ZN(new_n22179_));
  AOI21_X1   g21987(.A1(new_n22179_), .A2(new_n21745_), .B(new_n9846_), .ZN(new_n22180_));
  NOR3_X1    g21988(.A1(new_n22176_), .A2(\asqrt[23] ), .A3(new_n22172_), .ZN(new_n22181_));
  OAI21_X1   g21989(.A1(new_n21741_), .A2(new_n22181_), .B(new_n22177_), .ZN(new_n22182_));
  AOI21_X1   g21990(.A1(new_n22182_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n22183_));
  AOI21_X1   g21991(.A1(new_n22183_), .A2(new_n22179_), .B(new_n21759_), .ZN(new_n22184_));
  OAI21_X1   g21992(.A1(new_n22184_), .A2(new_n22180_), .B(\asqrt[26] ), .ZN(new_n22185_));
  NAND2_X1   g21993(.A1(new_n22185_), .A2(new_n8826_), .ZN(new_n22186_));
  OAI21_X1   g21994(.A1(new_n22186_), .A2(new_n21770_), .B(new_n22116_), .ZN(new_n22187_));
  AOI21_X1   g21995(.A1(new_n22187_), .A2(new_n21771_), .B(new_n8483_), .ZN(new_n22188_));
  NOR3_X1    g21996(.A1(new_n22184_), .A2(\asqrt[26] ), .A3(new_n22180_), .ZN(new_n22189_));
  OAI21_X1   g21997(.A1(new_n21767_), .A2(new_n22189_), .B(new_n22185_), .ZN(new_n22190_));
  AOI21_X1   g21998(.A1(new_n22190_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n22191_));
  AOI21_X1   g21999(.A1(new_n22191_), .A2(new_n22187_), .B(new_n21785_), .ZN(new_n22192_));
  OAI21_X1   g22000(.A1(new_n22192_), .A2(new_n22188_), .B(\asqrt[29] ), .ZN(new_n22193_));
  NAND2_X1   g22001(.A1(new_n22193_), .A2(new_n7539_), .ZN(new_n22194_));
  OAI21_X1   g22002(.A1(new_n22194_), .A2(new_n21796_), .B(new_n22115_), .ZN(new_n22195_));
  AOI21_X1   g22003(.A1(new_n22195_), .A2(new_n21797_), .B(new_n7229_), .ZN(new_n22196_));
  NOR3_X1    g22004(.A1(new_n22192_), .A2(\asqrt[29] ), .A3(new_n22188_), .ZN(new_n22197_));
  OAI21_X1   g22005(.A1(new_n21793_), .A2(new_n22197_), .B(new_n22193_), .ZN(new_n22198_));
  AOI21_X1   g22006(.A1(new_n22198_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n22199_));
  AOI21_X1   g22007(.A1(new_n22199_), .A2(new_n22195_), .B(new_n21811_), .ZN(new_n22200_));
  OAI21_X1   g22008(.A1(new_n22200_), .A2(new_n22196_), .B(\asqrt[32] ), .ZN(new_n22201_));
  NAND2_X1   g22009(.A1(new_n22201_), .A2(new_n6356_), .ZN(new_n22202_));
  OAI21_X1   g22010(.A1(new_n22202_), .A2(new_n21822_), .B(new_n22114_), .ZN(new_n22203_));
  AOI21_X1   g22011(.A1(new_n22203_), .A2(new_n21823_), .B(new_n6077_), .ZN(new_n22204_));
  NOR3_X1    g22012(.A1(new_n22200_), .A2(\asqrt[32] ), .A3(new_n22196_), .ZN(new_n22205_));
  OAI21_X1   g22013(.A1(new_n21819_), .A2(new_n22205_), .B(new_n22201_), .ZN(new_n22206_));
  AOI21_X1   g22014(.A1(new_n22206_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n22207_));
  AOI21_X1   g22015(.A1(new_n22207_), .A2(new_n22203_), .B(new_n21837_), .ZN(new_n22208_));
  OAI21_X1   g22016(.A1(new_n22208_), .A2(new_n22204_), .B(\asqrt[35] ), .ZN(new_n22209_));
  NAND2_X1   g22017(.A1(new_n22209_), .A2(new_n5277_), .ZN(new_n22210_));
  OAI21_X1   g22018(.A1(new_n22210_), .A2(new_n21848_), .B(new_n22113_), .ZN(new_n22211_));
  AOI21_X1   g22019(.A1(new_n22211_), .A2(new_n21849_), .B(new_n5024_), .ZN(new_n22212_));
  NOR3_X1    g22020(.A1(new_n22208_), .A2(\asqrt[35] ), .A3(new_n22204_), .ZN(new_n22213_));
  OAI21_X1   g22021(.A1(new_n21845_), .A2(new_n22213_), .B(new_n22209_), .ZN(new_n22214_));
  AOI21_X1   g22022(.A1(new_n22214_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n22215_));
  AOI21_X1   g22023(.A1(new_n22215_), .A2(new_n22211_), .B(new_n21863_), .ZN(new_n22216_));
  OAI21_X1   g22024(.A1(new_n22216_), .A2(new_n22212_), .B(\asqrt[38] ), .ZN(new_n22217_));
  NAND2_X1   g22025(.A1(new_n22217_), .A2(new_n4298_), .ZN(new_n22218_));
  OAI21_X1   g22026(.A1(new_n22218_), .A2(new_n21874_), .B(new_n22112_), .ZN(new_n22219_));
  AOI21_X1   g22027(.A1(new_n22219_), .A2(new_n21875_), .B(new_n4071_), .ZN(new_n22220_));
  NOR3_X1    g22028(.A1(new_n22216_), .A2(\asqrt[38] ), .A3(new_n22212_), .ZN(new_n22221_));
  OAI21_X1   g22029(.A1(new_n21871_), .A2(new_n22221_), .B(new_n22217_), .ZN(new_n22222_));
  AOI21_X1   g22030(.A1(new_n22222_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n22223_));
  AOI21_X1   g22031(.A1(new_n22223_), .A2(new_n22219_), .B(new_n21889_), .ZN(new_n22224_));
  OAI21_X1   g22032(.A1(new_n22224_), .A2(new_n22220_), .B(\asqrt[41] ), .ZN(new_n22225_));
  NAND2_X1   g22033(.A1(new_n22225_), .A2(new_n3419_), .ZN(new_n22226_));
  OAI21_X1   g22034(.A1(new_n22226_), .A2(new_n21900_), .B(new_n22111_), .ZN(new_n22227_));
  AOI21_X1   g22035(.A1(new_n22227_), .A2(new_n21901_), .B(new_n3218_), .ZN(new_n22228_));
  NOR3_X1    g22036(.A1(new_n22224_), .A2(\asqrt[41] ), .A3(new_n22220_), .ZN(new_n22229_));
  OAI21_X1   g22037(.A1(new_n21897_), .A2(new_n22229_), .B(new_n22225_), .ZN(new_n22230_));
  AOI21_X1   g22038(.A1(new_n22230_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n22231_));
  AOI21_X1   g22039(.A1(new_n22231_), .A2(new_n22227_), .B(new_n21915_), .ZN(new_n22232_));
  OAI21_X1   g22040(.A1(new_n22232_), .A2(new_n22228_), .B(\asqrt[44] ), .ZN(new_n22233_));
  NAND2_X1   g22041(.A1(new_n22233_), .A2(new_n2641_), .ZN(new_n22234_));
  OAI21_X1   g22042(.A1(new_n22234_), .A2(new_n21926_), .B(new_n22110_), .ZN(new_n22235_));
  AOI21_X1   g22043(.A1(new_n22235_), .A2(new_n21927_), .B(new_n2465_), .ZN(new_n22236_));
  NOR3_X1    g22044(.A1(new_n22232_), .A2(\asqrt[44] ), .A3(new_n22228_), .ZN(new_n22237_));
  OAI21_X1   g22045(.A1(new_n21923_), .A2(new_n22237_), .B(new_n22233_), .ZN(new_n22238_));
  AOI21_X1   g22046(.A1(new_n22238_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n22239_));
  AOI21_X1   g22047(.A1(new_n22239_), .A2(new_n22235_), .B(new_n21941_), .ZN(new_n22240_));
  OAI21_X1   g22048(.A1(new_n22240_), .A2(new_n22236_), .B(\asqrt[47] ), .ZN(new_n22241_));
  NAND2_X1   g22049(.A1(new_n22241_), .A2(new_n1956_), .ZN(new_n22242_));
  OAI21_X1   g22050(.A1(new_n22242_), .A2(new_n21952_), .B(new_n22109_), .ZN(new_n22243_));
  AOI21_X1   g22051(.A1(new_n22243_), .A2(new_n21953_), .B(new_n1806_), .ZN(new_n22244_));
  NOR3_X1    g22052(.A1(new_n22240_), .A2(\asqrt[47] ), .A3(new_n22236_), .ZN(new_n22245_));
  OAI21_X1   g22053(.A1(new_n21949_), .A2(new_n22245_), .B(new_n22241_), .ZN(new_n22246_));
  AOI21_X1   g22054(.A1(new_n22246_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n22247_));
  AOI21_X1   g22055(.A1(new_n22247_), .A2(new_n22243_), .B(new_n21967_), .ZN(new_n22248_));
  OAI21_X1   g22056(.A1(new_n22248_), .A2(new_n22244_), .B(\asqrt[50] ), .ZN(new_n22249_));
  NAND2_X1   g22057(.A1(new_n22249_), .A2(new_n1376_), .ZN(new_n22250_));
  OAI21_X1   g22058(.A1(new_n22250_), .A2(new_n21978_), .B(new_n22108_), .ZN(new_n22251_));
  AOI21_X1   g22059(.A1(new_n22251_), .A2(new_n21979_), .B(new_n1256_), .ZN(new_n22252_));
  NOR3_X1    g22060(.A1(new_n22248_), .A2(\asqrt[50] ), .A3(new_n22244_), .ZN(new_n22253_));
  OAI21_X1   g22061(.A1(new_n21975_), .A2(new_n22253_), .B(new_n22249_), .ZN(new_n22254_));
  AOI21_X1   g22062(.A1(new_n22254_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n22255_));
  AOI21_X1   g22063(.A1(new_n22255_), .A2(new_n22251_), .B(new_n21995_), .ZN(new_n22256_));
  OAI21_X1   g22064(.A1(new_n22256_), .A2(new_n22252_), .B(\asqrt[53] ), .ZN(new_n22257_));
  NAND2_X1   g22065(.A1(new_n22257_), .A2(new_n904_), .ZN(new_n22258_));
  OAI21_X1   g22066(.A1(new_n22258_), .A2(new_n22006_), .B(new_n22107_), .ZN(new_n22259_));
  AOI21_X1   g22067(.A1(new_n22259_), .A2(new_n22007_), .B(new_n823_), .ZN(new_n22260_));
  NOR3_X1    g22068(.A1(new_n22256_), .A2(\asqrt[53] ), .A3(new_n22252_), .ZN(new_n22261_));
  OAI21_X1   g22069(.A1(new_n22003_), .A2(new_n22261_), .B(new_n22257_), .ZN(new_n22262_));
  AOI21_X1   g22070(.A1(new_n22262_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n22263_));
  AOI21_X1   g22071(.A1(new_n22263_), .A2(new_n22259_), .B(new_n22026_), .ZN(new_n22264_));
  OAI21_X1   g22072(.A1(new_n22264_), .A2(new_n22260_), .B(\asqrt[56] ), .ZN(new_n22265_));
  NAND2_X1   g22073(.A1(new_n22265_), .A2(new_n531_), .ZN(new_n22266_));
  OAI21_X1   g22074(.A1(new_n22266_), .A2(new_n22037_), .B(new_n22106_), .ZN(new_n22267_));
  AOI21_X1   g22075(.A1(new_n22267_), .A2(new_n22038_), .B(new_n436_), .ZN(new_n22268_));
  NOR3_X1    g22076(.A1(new_n22264_), .A2(\asqrt[56] ), .A3(new_n22260_), .ZN(new_n22269_));
  OAI21_X1   g22077(.A1(new_n22034_), .A2(new_n22269_), .B(new_n22265_), .ZN(new_n22270_));
  AOI21_X1   g22078(.A1(new_n22270_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n22271_));
  AOI21_X1   g22079(.A1(new_n22271_), .A2(new_n22267_), .B(new_n22056_), .ZN(new_n22272_));
  OAI21_X1   g22080(.A1(new_n22272_), .A2(new_n22268_), .B(\asqrt[59] ), .ZN(new_n22273_));
  NAND2_X1   g22081(.A1(new_n22273_), .A2(new_n306_), .ZN(new_n22274_));
  OAI21_X1   g22082(.A1(new_n22274_), .A2(new_n22067_), .B(new_n22105_), .ZN(new_n22275_));
  NOR3_X1    g22083(.A1(new_n22272_), .A2(\asqrt[59] ), .A3(new_n22268_), .ZN(new_n22276_));
  OAI21_X1   g22084(.A1(new_n22064_), .A2(new_n22276_), .B(new_n22273_), .ZN(new_n22277_));
  AOI21_X1   g22085(.A1(new_n22277_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n22278_));
  AOI21_X1   g22086(.A1(new_n22278_), .A2(new_n22275_), .B(new_n22081_), .ZN(new_n22279_));
  INV_X1     g22087(.I(new_n22089_), .ZN(new_n22280_));
  NAND2_X1   g22088(.A1(new_n22077_), .A2(new_n207_), .ZN(new_n22281_));
  OAI21_X1   g22089(.A1(new_n22281_), .A2(new_n22279_), .B(new_n22280_), .ZN(new_n22282_));
  NOR2_X1    g22090(.A1(new_n22085_), .A2(new_n22099_), .ZN(new_n22283_));
  AOI21_X1   g22091(.A1(\asqrt[5] ), .A2(new_n21548_), .B(new_n21566_), .ZN(new_n22284_));
  NOR2_X1    g22092(.A1(new_n22100_), .A2(new_n193_), .ZN(new_n22285_));
  INV_X1     g22093(.I(new_n22285_), .ZN(new_n22286_));
  NOR2_X1    g22094(.A1(new_n22284_), .A2(new_n22286_), .ZN(new_n22287_));
  AOI21_X1   g22095(.A1(new_n22283_), .A2(new_n22282_), .B(new_n22287_), .ZN(new_n22288_));
  NAND2_X1   g22096(.A1(new_n22104_), .A2(new_n22288_), .ZN(\asqrt[4] ));
  NOR2_X1    g22097(.A1(\a[6] ), .A2(\a[7] ), .ZN(new_n22290_));
  INV_X1     g22098(.I(new_n22290_), .ZN(new_n22291_));
  NOR2_X1    g22099(.A1(new_n22291_), .A2(\a[8] ), .ZN(new_n22292_));
  INV_X1     g22100(.I(new_n22292_), .ZN(new_n22293_));
  AOI21_X1   g22101(.A1(new_n22275_), .A2(new_n22068_), .B(new_n218_), .ZN(new_n22294_));
  OAI21_X1   g22102(.A1(new_n22279_), .A2(new_n22294_), .B(\asqrt[62] ), .ZN(new_n22295_));
  NOR3_X1    g22103(.A1(new_n22279_), .A2(\asqrt[62] ), .A3(new_n22294_), .ZN(new_n22296_));
  OAI21_X1   g22104(.A1(new_n22089_), .A2(new_n22296_), .B(new_n22295_), .ZN(new_n22297_));
  AOI21_X1   g22105(.A1(new_n22297_), .A2(new_n22102_), .B(\asqrt[63] ), .ZN(new_n22298_));
  NAND2_X1   g22106(.A1(new_n22295_), .A2(new_n22098_), .ZN(new_n22299_));
  OAI22_X1   g22107(.A1(new_n22299_), .A2(new_n22092_), .B1(new_n22284_), .B2(new_n22286_), .ZN(new_n22300_));
  OAI21_X1   g22108(.A1(new_n22298_), .A2(new_n22300_), .B(\a[8] ), .ZN(new_n22301_));
  AOI21_X1   g22109(.A1(new_n22301_), .A2(new_n22293_), .B(new_n21620_), .ZN(new_n22302_));
  INV_X1     g22110(.I(\a[8] ), .ZN(new_n22303_));
  AOI21_X1   g22111(.A1(new_n22104_), .A2(new_n22288_), .B(new_n22303_), .ZN(new_n22304_));
  NAND4_X1   g22112(.A1(new_n21584_), .A2(new_n21596_), .A3(new_n21558_), .A4(new_n22293_), .ZN(new_n22305_));
  NOR2_X1    g22113(.A1(new_n22304_), .A2(new_n22305_), .ZN(new_n22306_));
  AOI21_X1   g22114(.A1(new_n22104_), .A2(new_n22288_), .B(new_n21563_), .ZN(new_n22307_));
  INV_X1     g22115(.I(\a[9] ), .ZN(new_n22308_));
  AOI21_X1   g22116(.A1(\asqrt[4] ), .A2(new_n22303_), .B(new_n22308_), .ZN(new_n22309_));
  NOR3_X1    g22117(.A1(new_n22306_), .A2(new_n22309_), .A3(new_n22307_), .ZN(new_n22310_));
  OAI21_X1   g22118(.A1(new_n22310_), .A2(new_n22302_), .B(\asqrt[6] ), .ZN(new_n22311_));
  OAI21_X1   g22119(.A1(new_n22298_), .A2(new_n22300_), .B(new_n21562_), .ZN(new_n22312_));
  NOR2_X1    g22120(.A1(new_n22299_), .A2(new_n22092_), .ZN(new_n22313_));
  NOR3_X1    g22121(.A1(new_n22313_), .A2(new_n21620_), .A3(new_n22287_), .ZN(new_n22314_));
  NAND2_X1   g22122(.A1(new_n22314_), .A2(new_n22104_), .ZN(new_n22315_));
  AOI21_X1   g22123(.A1(new_n22315_), .A2(new_n22312_), .B(new_n21581_), .ZN(new_n22316_));
  NOR4_X1    g22124(.A1(new_n22298_), .A2(new_n21620_), .A3(new_n22313_), .A4(new_n22287_), .ZN(new_n22317_));
  NOR3_X1    g22125(.A1(new_n22317_), .A2(new_n22307_), .A3(\a[10] ), .ZN(new_n22318_));
  OAI21_X1   g22126(.A1(new_n22304_), .A2(new_n22292_), .B(\asqrt[5] ), .ZN(new_n22319_));
  NAND2_X1   g22127(.A1(new_n22319_), .A2(new_n20806_), .ZN(new_n22320_));
  OAI22_X1   g22128(.A1(new_n22310_), .A2(new_n22320_), .B1(new_n22316_), .B2(new_n22318_), .ZN(new_n22321_));
  AOI21_X1   g22129(.A1(new_n22321_), .A2(new_n22311_), .B(new_n20262_), .ZN(new_n22322_));
  NOR3_X1    g22130(.A1(new_n22137_), .A2(new_n21580_), .A3(new_n21589_), .ZN(new_n22323_));
  NAND3_X1   g22131(.A1(\asqrt[4] ), .A2(new_n21609_), .A3(new_n22122_), .ZN(new_n22324_));
  AOI22_X1   g22132(.A1(new_n22324_), .A2(new_n22137_), .B1(\asqrt[4] ), .B2(new_n22323_), .ZN(new_n22325_));
  AOI21_X1   g22133(.A1(new_n22104_), .A2(new_n22288_), .B(\a[8] ), .ZN(new_n22326_));
  OAI21_X1   g22134(.A1(new_n22308_), .A2(new_n22326_), .B(new_n22312_), .ZN(new_n22327_));
  OAI21_X1   g22135(.A1(new_n22327_), .A2(new_n22306_), .B(new_n22319_), .ZN(new_n22328_));
  AOI21_X1   g22136(.A1(new_n22328_), .A2(\asqrt[6] ), .B(\asqrt[7] ), .ZN(new_n22329_));
  AOI21_X1   g22137(.A1(new_n22329_), .A2(new_n22321_), .B(new_n22325_), .ZN(new_n22330_));
  OAI21_X1   g22138(.A1(new_n22330_), .A2(new_n22322_), .B(\asqrt[8] ), .ZN(new_n22331_));
  INV_X1     g22139(.I(new_n22331_), .ZN(new_n22332_));
  NOR2_X1    g22140(.A1(new_n21601_), .A2(new_n21598_), .ZN(new_n22333_));
  NOR2_X1    g22141(.A1(new_n21593_), .A2(new_n21603_), .ZN(new_n22334_));
  INV_X1     g22142(.I(new_n22334_), .ZN(new_n22335_));
  NAND4_X1   g22143(.A1(\asqrt[4] ), .A2(new_n21594_), .A3(new_n22333_), .A4(new_n22335_), .ZN(new_n22336_));
  INV_X1     g22144(.I(\asqrt[4] ), .ZN(new_n22337_));
  NOR3_X1    g22145(.A1(new_n22337_), .A2(new_n22126_), .A3(new_n22334_), .ZN(new_n22338_));
  OAI21_X1   g22146(.A1(new_n22338_), .A2(new_n22333_), .B(new_n22336_), .ZN(new_n22339_));
  INV_X1     g22147(.I(new_n22339_), .ZN(new_n22340_));
  NOR3_X1    g22148(.A1(new_n22330_), .A2(new_n22322_), .A3(\asqrt[8] ), .ZN(new_n22341_));
  NOR2_X1    g22149(.A1(new_n22341_), .A2(new_n22340_), .ZN(new_n22342_));
  OAI21_X1   g22150(.A1(new_n22342_), .A2(new_n22332_), .B(\asqrt[9] ), .ZN(new_n22343_));
  NOR2_X1    g22151(.A1(new_n22139_), .A2(new_n22131_), .ZN(new_n22344_));
  NOR3_X1    g22152(.A1(new_n22337_), .A2(new_n21605_), .A3(new_n22344_), .ZN(new_n22345_));
  INV_X1     g22153(.I(new_n22345_), .ZN(new_n22346_));
  NOR3_X1    g22154(.A1(new_n22344_), .A2(new_n21605_), .A3(new_n22136_), .ZN(new_n22347_));
  AOI22_X1   g22155(.A1(new_n22346_), .A2(new_n22136_), .B1(\asqrt[4] ), .B2(new_n22347_), .ZN(new_n22348_));
  INV_X1     g22156(.I(new_n22348_), .ZN(new_n22349_));
  NAND2_X1   g22157(.A1(new_n22331_), .A2(new_n18792_), .ZN(new_n22350_));
  OAI21_X1   g22158(.A1(new_n22342_), .A2(new_n22350_), .B(new_n22349_), .ZN(new_n22351_));
  AOI21_X1   g22159(.A1(new_n22351_), .A2(new_n22343_), .B(new_n18275_), .ZN(new_n22352_));
  NOR3_X1    g22160(.A1(new_n21616_), .A2(new_n21624_), .A3(new_n21622_), .ZN(new_n22353_));
  NOR3_X1    g22161(.A1(new_n22337_), .A2(new_n21616_), .A3(new_n21624_), .ZN(new_n22354_));
  INV_X1     g22162(.I(new_n22354_), .ZN(new_n22355_));
  AOI22_X1   g22163(.A1(new_n22355_), .A2(new_n21622_), .B1(\asqrt[4] ), .B2(new_n22353_), .ZN(new_n22356_));
  OAI21_X1   g22164(.A1(new_n22340_), .A2(new_n22341_), .B(new_n22331_), .ZN(new_n22357_));
  AOI21_X1   g22165(.A1(new_n22357_), .A2(\asqrt[9] ), .B(\asqrt[10] ), .ZN(new_n22358_));
  AOI21_X1   g22166(.A1(new_n22358_), .A2(new_n22351_), .B(new_n22356_), .ZN(new_n22359_));
  OAI21_X1   g22167(.A1(new_n22359_), .A2(new_n22352_), .B(\asqrt[11] ), .ZN(new_n22360_));
  NAND2_X1   g22168(.A1(new_n22142_), .A2(new_n22134_), .ZN(new_n22361_));
  NAND3_X1   g22169(.A1(\asqrt[4] ), .A2(new_n21626_), .A3(new_n22361_), .ZN(new_n22362_));
  AND3_X2    g22170(.A1(new_n21626_), .A2(new_n21630_), .A3(new_n22361_), .Z(new_n22363_));
  AOI22_X1   g22171(.A1(new_n22362_), .A2(new_n21631_), .B1(\asqrt[4] ), .B2(new_n22363_), .ZN(new_n22364_));
  INV_X1     g22172(.I(new_n22364_), .ZN(new_n22365_));
  INV_X1     g22173(.I(new_n22305_), .ZN(new_n22366_));
  NAND2_X1   g22174(.A1(new_n22301_), .A2(new_n22366_), .ZN(new_n22367_));
  OAI21_X1   g22175(.A1(new_n22298_), .A2(new_n22300_), .B(new_n22303_), .ZN(new_n22368_));
  NAND2_X1   g22176(.A1(new_n22368_), .A2(\a[9] ), .ZN(new_n22369_));
  NAND3_X1   g22177(.A1(new_n22367_), .A2(new_n22369_), .A3(new_n22312_), .ZN(new_n22370_));
  AOI21_X1   g22178(.A1(new_n22370_), .A2(new_n22319_), .B(new_n20806_), .ZN(new_n22371_));
  OAI21_X1   g22179(.A1(new_n22317_), .A2(new_n22307_), .B(\a[10] ), .ZN(new_n22372_));
  NAND3_X1   g22180(.A1(new_n22315_), .A2(new_n21581_), .A3(new_n22312_), .ZN(new_n22373_));
  NAND2_X1   g22181(.A1(new_n22301_), .A2(new_n22293_), .ZN(new_n22374_));
  AOI21_X1   g22182(.A1(new_n22374_), .A2(\asqrt[5] ), .B(\asqrt[6] ), .ZN(new_n22375_));
  AOI22_X1   g22183(.A1(new_n22370_), .A2(new_n22375_), .B1(new_n22372_), .B2(new_n22373_), .ZN(new_n22376_));
  OAI21_X1   g22184(.A1(new_n22376_), .A2(new_n22371_), .B(\asqrt[7] ), .ZN(new_n22377_));
  NAND2_X1   g22185(.A1(new_n22377_), .A2(new_n19573_), .ZN(new_n22378_));
  OAI21_X1   g22186(.A1(new_n22378_), .A2(new_n22330_), .B(new_n22339_), .ZN(new_n22379_));
  AOI21_X1   g22187(.A1(new_n22379_), .A2(new_n22331_), .B(new_n18792_), .ZN(new_n22380_));
  INV_X1     g22188(.I(new_n22325_), .ZN(new_n22381_));
  AOI21_X1   g22189(.A1(\a[9] ), .A2(new_n22368_), .B(new_n22307_), .ZN(new_n22382_));
  AOI21_X1   g22190(.A1(new_n22382_), .A2(new_n22367_), .B(new_n22302_), .ZN(new_n22383_));
  OAI21_X1   g22191(.A1(new_n22383_), .A2(new_n20806_), .B(new_n20262_), .ZN(new_n22384_));
  OAI21_X1   g22192(.A1(new_n22384_), .A2(new_n22376_), .B(new_n22381_), .ZN(new_n22385_));
  NAND2_X1   g22193(.A1(new_n22385_), .A2(new_n22377_), .ZN(new_n22386_));
  AOI21_X1   g22194(.A1(new_n22386_), .A2(\asqrt[8] ), .B(\asqrt[9] ), .ZN(new_n22387_));
  AOI21_X1   g22195(.A1(new_n22387_), .A2(new_n22379_), .B(new_n22348_), .ZN(new_n22388_));
  OAI21_X1   g22196(.A1(new_n22388_), .A2(new_n22380_), .B(\asqrt[10] ), .ZN(new_n22389_));
  NAND2_X1   g22197(.A1(new_n22389_), .A2(new_n17623_), .ZN(new_n22390_));
  OAI21_X1   g22198(.A1(new_n22390_), .A2(new_n22359_), .B(new_n22365_), .ZN(new_n22391_));
  AOI21_X1   g22199(.A1(new_n22391_), .A2(new_n22360_), .B(new_n16881_), .ZN(new_n22392_));
  INV_X1     g22200(.I(new_n21638_), .ZN(new_n22393_));
  NOR3_X1    g22201(.A1(new_n21634_), .A2(new_n22153_), .A3(new_n22393_), .ZN(new_n22394_));
  NOR3_X1    g22202(.A1(new_n22337_), .A2(new_n21634_), .A3(new_n22153_), .ZN(new_n22395_));
  INV_X1     g22203(.I(new_n22395_), .ZN(new_n22396_));
  AOI22_X1   g22204(.A1(new_n22396_), .A2(new_n22393_), .B1(\asqrt[4] ), .B2(new_n22394_), .ZN(new_n22397_));
  NOR3_X1    g22205(.A1(new_n22388_), .A2(new_n22380_), .A3(\asqrt[10] ), .ZN(new_n22398_));
  OAI21_X1   g22206(.A1(new_n22356_), .A2(new_n22398_), .B(new_n22389_), .ZN(new_n22399_));
  AOI21_X1   g22207(.A1(new_n22399_), .A2(\asqrt[11] ), .B(\asqrt[12] ), .ZN(new_n22400_));
  AOI21_X1   g22208(.A1(new_n22400_), .A2(new_n22391_), .B(new_n22397_), .ZN(new_n22401_));
  OAI21_X1   g22209(.A1(new_n22401_), .A2(new_n22392_), .B(\asqrt[13] ), .ZN(new_n22402_));
  INV_X1     g22210(.I(new_n22402_), .ZN(new_n22403_));
  NOR3_X1    g22211(.A1(new_n22337_), .A2(new_n21643_), .A3(new_n21648_), .ZN(new_n22404_));
  INV_X1     g22212(.I(new_n22404_), .ZN(new_n22405_));
  NOR3_X1    g22213(.A1(new_n21643_), .A2(new_n22121_), .A3(new_n21648_), .ZN(new_n22406_));
  AOI22_X1   g22214(.A1(new_n22405_), .A2(new_n22121_), .B1(\asqrt[4] ), .B2(new_n22406_), .ZN(new_n22407_));
  NOR3_X1    g22215(.A1(new_n22401_), .A2(\asqrt[13] ), .A3(new_n22392_), .ZN(new_n22408_));
  NOR2_X1    g22216(.A1(new_n22408_), .A2(new_n22407_), .ZN(new_n22409_));
  OAI21_X1   g22217(.A1(new_n22409_), .A2(new_n22403_), .B(\asqrt[14] ), .ZN(new_n22410_));
  INV_X1     g22218(.I(new_n22147_), .ZN(new_n22411_));
  NOR3_X1    g22219(.A1(new_n22411_), .A2(new_n22152_), .A3(new_n21656_), .ZN(new_n22412_));
  NOR3_X1    g22220(.A1(new_n22337_), .A2(new_n22152_), .A3(new_n22411_), .ZN(new_n22413_));
  INV_X1     g22221(.I(new_n22413_), .ZN(new_n22414_));
  AOI22_X1   g22222(.A1(new_n22414_), .A2(new_n21656_), .B1(\asqrt[4] ), .B2(new_n22412_), .ZN(new_n22415_));
  INV_X1     g22223(.I(new_n22415_), .ZN(new_n22416_));
  NAND2_X1   g22224(.A1(new_n22402_), .A2(new_n15770_), .ZN(new_n22417_));
  OAI21_X1   g22225(.A1(new_n22409_), .A2(new_n22417_), .B(new_n22416_), .ZN(new_n22418_));
  AOI21_X1   g22226(.A1(new_n22418_), .A2(new_n22410_), .B(new_n15067_), .ZN(new_n22419_));
  INV_X1     g22227(.I(new_n21663_), .ZN(new_n22420_));
  NOR3_X1    g22228(.A1(new_n22337_), .A2(new_n21659_), .A3(new_n22157_), .ZN(new_n22421_));
  INV_X1     g22229(.I(new_n22421_), .ZN(new_n22422_));
  NOR3_X1    g22230(.A1(new_n21659_), .A2(new_n22157_), .A3(new_n22420_), .ZN(new_n22423_));
  AOI22_X1   g22231(.A1(new_n22422_), .A2(new_n22420_), .B1(\asqrt[4] ), .B2(new_n22423_), .ZN(new_n22424_));
  NOR3_X1    g22232(.A1(new_n22359_), .A2(new_n22352_), .A3(\asqrt[11] ), .ZN(new_n22425_));
  OAI21_X1   g22233(.A1(new_n22364_), .A2(new_n22425_), .B(new_n22360_), .ZN(new_n22426_));
  INV_X1     g22234(.I(new_n22397_), .ZN(new_n22427_));
  NAND3_X1   g22235(.A1(new_n22391_), .A2(new_n16881_), .A3(new_n22360_), .ZN(new_n22428_));
  AOI22_X1   g22236(.A1(new_n22428_), .A2(new_n22427_), .B1(new_n22426_), .B2(\asqrt[12] ), .ZN(new_n22429_));
  OAI22_X1   g22237(.A1(new_n22408_), .A2(new_n22407_), .B1(new_n22429_), .B2(new_n16389_), .ZN(new_n22430_));
  AOI21_X1   g22238(.A1(new_n22430_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n22431_));
  AOI21_X1   g22239(.A1(new_n22431_), .A2(new_n22418_), .B(new_n22424_), .ZN(new_n22432_));
  OAI21_X1   g22240(.A1(new_n22432_), .A2(new_n22419_), .B(\asqrt[16] ), .ZN(new_n22433_));
  INV_X1     g22241(.I(new_n22433_), .ZN(new_n22434_));
  NOR3_X1    g22242(.A1(new_n21668_), .A2(new_n22120_), .A3(new_n21674_), .ZN(new_n22435_));
  NOR3_X1    g22243(.A1(new_n22337_), .A2(new_n21668_), .A3(new_n21674_), .ZN(new_n22436_));
  INV_X1     g22244(.I(new_n22436_), .ZN(new_n22437_));
  AOI22_X1   g22245(.A1(new_n22437_), .A2(new_n22120_), .B1(\asqrt[4] ), .B2(new_n22435_), .ZN(new_n22438_));
  NOR3_X1    g22246(.A1(new_n22432_), .A2(new_n22419_), .A3(\asqrt[16] ), .ZN(new_n22439_));
  NOR2_X1    g22247(.A1(new_n22439_), .A2(new_n22438_), .ZN(new_n22440_));
  OAI21_X1   g22248(.A1(new_n22440_), .A2(new_n22434_), .B(\asqrt[17] ), .ZN(new_n22441_));
  NOR2_X1    g22249(.A1(new_n21675_), .A2(new_n21683_), .ZN(new_n22442_));
  NOR3_X1    g22250(.A1(new_n22337_), .A2(new_n22151_), .A3(new_n22442_), .ZN(new_n22443_));
  INV_X1     g22251(.I(new_n22443_), .ZN(new_n22444_));
  NOR3_X1    g22252(.A1(new_n22442_), .A2(new_n22151_), .A3(new_n21682_), .ZN(new_n22445_));
  AOI22_X1   g22253(.A1(new_n22444_), .A2(new_n21682_), .B1(\asqrt[4] ), .B2(new_n22445_), .ZN(new_n22446_));
  INV_X1     g22254(.I(new_n22446_), .ZN(new_n22447_));
  NAND2_X1   g22255(.A1(new_n22433_), .A2(new_n14017_), .ZN(new_n22448_));
  OAI21_X1   g22256(.A1(new_n22440_), .A2(new_n22448_), .B(new_n22447_), .ZN(new_n22449_));
  AOI21_X1   g22257(.A1(new_n22449_), .A2(new_n22441_), .B(new_n13353_), .ZN(new_n22450_));
  INV_X1     g22258(.I(new_n21689_), .ZN(new_n22451_));
  NOR3_X1    g22259(.A1(new_n21685_), .A2(new_n22165_), .A3(new_n22451_), .ZN(new_n22452_));
  NOR3_X1    g22260(.A1(new_n22337_), .A2(new_n21685_), .A3(new_n22165_), .ZN(new_n22453_));
  INV_X1     g22261(.I(new_n22453_), .ZN(new_n22454_));
  AOI22_X1   g22262(.A1(new_n22454_), .A2(new_n22451_), .B1(\asqrt[4] ), .B2(new_n22452_), .ZN(new_n22455_));
  OAI21_X1   g22263(.A1(new_n22438_), .A2(new_n22439_), .B(new_n22433_), .ZN(new_n22456_));
  AOI21_X1   g22264(.A1(new_n22456_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n22457_));
  AOI21_X1   g22265(.A1(new_n22457_), .A2(new_n22449_), .B(new_n22455_), .ZN(new_n22458_));
  OAI21_X1   g22266(.A1(new_n22458_), .A2(new_n22450_), .B(\asqrt[19] ), .ZN(new_n22459_));
  INV_X1     g22267(.I(new_n22459_), .ZN(new_n22460_));
  NOR3_X1    g22268(.A1(new_n22337_), .A2(new_n21694_), .A3(new_n21700_), .ZN(new_n22461_));
  INV_X1     g22269(.I(new_n22461_), .ZN(new_n22462_));
  NOR3_X1    g22270(.A1(new_n21694_), .A2(new_n22119_), .A3(new_n21700_), .ZN(new_n22463_));
  AOI22_X1   g22271(.A1(new_n22462_), .A2(new_n22119_), .B1(\asqrt[4] ), .B2(new_n22463_), .ZN(new_n22464_));
  NOR3_X1    g22272(.A1(new_n22458_), .A2(new_n22450_), .A3(\asqrt[19] ), .ZN(new_n22465_));
  NOR2_X1    g22273(.A1(new_n22465_), .A2(new_n22464_), .ZN(new_n22466_));
  OAI21_X1   g22274(.A1(new_n22466_), .A2(new_n22460_), .B(\asqrt[20] ), .ZN(new_n22467_));
  NOR2_X1    g22275(.A1(new_n21701_), .A2(new_n21709_), .ZN(new_n22468_));
  NOR3_X1    g22276(.A1(new_n22468_), .A2(new_n22164_), .A3(new_n21708_), .ZN(new_n22469_));
  NOR3_X1    g22277(.A1(new_n22337_), .A2(new_n22164_), .A3(new_n22468_), .ZN(new_n22470_));
  INV_X1     g22278(.I(new_n22470_), .ZN(new_n22471_));
  AOI22_X1   g22279(.A1(new_n22471_), .A2(new_n21708_), .B1(\asqrt[4] ), .B2(new_n22469_), .ZN(new_n22472_));
  INV_X1     g22280(.I(new_n22472_), .ZN(new_n22473_));
  NAND2_X1   g22281(.A1(new_n22459_), .A2(new_n12364_), .ZN(new_n22474_));
  OAI21_X1   g22282(.A1(new_n22466_), .A2(new_n22474_), .B(new_n22473_), .ZN(new_n22475_));
  AOI21_X1   g22283(.A1(new_n22475_), .A2(new_n22467_), .B(new_n11736_), .ZN(new_n22476_));
  INV_X1     g22284(.I(new_n21715_), .ZN(new_n22477_));
  NOR3_X1    g22285(.A1(new_n22337_), .A2(new_n21711_), .A3(new_n22173_), .ZN(new_n22478_));
  INV_X1     g22286(.I(new_n22478_), .ZN(new_n22479_));
  NOR3_X1    g22287(.A1(new_n21711_), .A2(new_n22173_), .A3(new_n22477_), .ZN(new_n22480_));
  AOI22_X1   g22288(.A1(new_n22479_), .A2(new_n22477_), .B1(\asqrt[4] ), .B2(new_n22480_), .ZN(new_n22481_));
  OAI21_X1   g22289(.A1(new_n22464_), .A2(new_n22465_), .B(new_n22459_), .ZN(new_n22482_));
  AOI21_X1   g22290(.A1(new_n22482_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n22483_));
  AOI21_X1   g22291(.A1(new_n22483_), .A2(new_n22475_), .B(new_n22481_), .ZN(new_n22484_));
  OAI21_X1   g22292(.A1(new_n22484_), .A2(new_n22476_), .B(\asqrt[22] ), .ZN(new_n22485_));
  INV_X1     g22293(.I(new_n22485_), .ZN(new_n22486_));
  NOR3_X1    g22294(.A1(new_n21720_), .A2(new_n22118_), .A3(new_n21726_), .ZN(new_n22487_));
  NOR3_X1    g22295(.A1(new_n22337_), .A2(new_n21720_), .A3(new_n21726_), .ZN(new_n22488_));
  INV_X1     g22296(.I(new_n22488_), .ZN(new_n22489_));
  AOI22_X1   g22297(.A1(new_n22489_), .A2(new_n22118_), .B1(\asqrt[4] ), .B2(new_n22487_), .ZN(new_n22490_));
  NOR3_X1    g22298(.A1(new_n22484_), .A2(new_n22476_), .A3(\asqrt[22] ), .ZN(new_n22491_));
  NOR2_X1    g22299(.A1(new_n22491_), .A2(new_n22490_), .ZN(new_n22492_));
  OAI21_X1   g22300(.A1(new_n22492_), .A2(new_n22486_), .B(\asqrt[23] ), .ZN(new_n22493_));
  NOR2_X1    g22301(.A1(new_n21727_), .A2(new_n21735_), .ZN(new_n22494_));
  NOR3_X1    g22302(.A1(new_n22337_), .A2(new_n22172_), .A3(new_n22494_), .ZN(new_n22495_));
  INV_X1     g22303(.I(new_n22495_), .ZN(new_n22496_));
  NOR3_X1    g22304(.A1(new_n22494_), .A2(new_n22172_), .A3(new_n21734_), .ZN(new_n22497_));
  AOI22_X1   g22305(.A1(new_n22496_), .A2(new_n21734_), .B1(\asqrt[4] ), .B2(new_n22497_), .ZN(new_n22498_));
  INV_X1     g22306(.I(new_n22498_), .ZN(new_n22499_));
  NAND2_X1   g22307(.A1(new_n22485_), .A2(new_n10812_), .ZN(new_n22500_));
  OAI21_X1   g22308(.A1(new_n22492_), .A2(new_n22500_), .B(new_n22499_), .ZN(new_n22501_));
  AOI21_X1   g22309(.A1(new_n22501_), .A2(new_n22493_), .B(new_n10221_), .ZN(new_n22502_));
  INV_X1     g22310(.I(new_n21741_), .ZN(new_n22503_));
  NOR3_X1    g22311(.A1(new_n21737_), .A2(new_n22181_), .A3(new_n22503_), .ZN(new_n22504_));
  NOR3_X1    g22312(.A1(new_n22337_), .A2(new_n21737_), .A3(new_n22181_), .ZN(new_n22505_));
  INV_X1     g22313(.I(new_n22505_), .ZN(new_n22506_));
  AOI22_X1   g22314(.A1(new_n22506_), .A2(new_n22503_), .B1(\asqrt[4] ), .B2(new_n22504_), .ZN(new_n22507_));
  OAI21_X1   g22315(.A1(new_n22490_), .A2(new_n22491_), .B(new_n22485_), .ZN(new_n22508_));
  AOI21_X1   g22316(.A1(new_n22508_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n22509_));
  AOI21_X1   g22317(.A1(new_n22509_), .A2(new_n22501_), .B(new_n22507_), .ZN(new_n22510_));
  OAI21_X1   g22318(.A1(new_n22510_), .A2(new_n22502_), .B(\asqrt[25] ), .ZN(new_n22511_));
  INV_X1     g22319(.I(new_n22511_), .ZN(new_n22512_));
  NOR3_X1    g22320(.A1(new_n22337_), .A2(new_n21746_), .A3(new_n21752_), .ZN(new_n22513_));
  INV_X1     g22321(.I(new_n22513_), .ZN(new_n22514_));
  NOR3_X1    g22322(.A1(new_n21746_), .A2(new_n22117_), .A3(new_n21752_), .ZN(new_n22515_));
  AOI22_X1   g22323(.A1(new_n22514_), .A2(new_n22117_), .B1(\asqrt[4] ), .B2(new_n22515_), .ZN(new_n22516_));
  NOR3_X1    g22324(.A1(new_n22510_), .A2(new_n22502_), .A3(\asqrt[25] ), .ZN(new_n22517_));
  NOR2_X1    g22325(.A1(new_n22517_), .A2(new_n22516_), .ZN(new_n22518_));
  OAI21_X1   g22326(.A1(new_n22518_), .A2(new_n22512_), .B(\asqrt[26] ), .ZN(new_n22519_));
  NOR2_X1    g22327(.A1(new_n21753_), .A2(new_n21761_), .ZN(new_n22520_));
  NOR3_X1    g22328(.A1(new_n22520_), .A2(new_n22180_), .A3(new_n21760_), .ZN(new_n22521_));
  NOR3_X1    g22329(.A1(new_n22337_), .A2(new_n22180_), .A3(new_n22520_), .ZN(new_n22522_));
  INV_X1     g22330(.I(new_n22522_), .ZN(new_n22523_));
  AOI22_X1   g22331(.A1(new_n22523_), .A2(new_n21760_), .B1(\asqrt[4] ), .B2(new_n22521_), .ZN(new_n22524_));
  INV_X1     g22332(.I(new_n22524_), .ZN(new_n22525_));
  NAND2_X1   g22333(.A1(new_n22511_), .A2(new_n9317_), .ZN(new_n22526_));
  OAI21_X1   g22334(.A1(new_n22518_), .A2(new_n22526_), .B(new_n22525_), .ZN(new_n22527_));
  AOI21_X1   g22335(.A1(new_n22527_), .A2(new_n22519_), .B(new_n8826_), .ZN(new_n22528_));
  INV_X1     g22336(.I(new_n21767_), .ZN(new_n22529_));
  NOR3_X1    g22337(.A1(new_n22337_), .A2(new_n21763_), .A3(new_n22189_), .ZN(new_n22530_));
  INV_X1     g22338(.I(new_n22530_), .ZN(new_n22531_));
  NOR3_X1    g22339(.A1(new_n21763_), .A2(new_n22189_), .A3(new_n22529_), .ZN(new_n22532_));
  AOI22_X1   g22340(.A1(new_n22531_), .A2(new_n22529_), .B1(\asqrt[4] ), .B2(new_n22532_), .ZN(new_n22533_));
  OAI21_X1   g22341(.A1(new_n22516_), .A2(new_n22517_), .B(new_n22511_), .ZN(new_n22534_));
  AOI21_X1   g22342(.A1(new_n22534_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n22535_));
  AOI21_X1   g22343(.A1(new_n22535_), .A2(new_n22527_), .B(new_n22533_), .ZN(new_n22536_));
  OAI21_X1   g22344(.A1(new_n22536_), .A2(new_n22528_), .B(\asqrt[28] ), .ZN(new_n22537_));
  INV_X1     g22345(.I(new_n22537_), .ZN(new_n22538_));
  INV_X1     g22346(.I(new_n22536_), .ZN(new_n22539_));
  NOR3_X1    g22347(.A1(new_n21772_), .A2(new_n22116_), .A3(new_n21778_), .ZN(new_n22540_));
  NOR3_X1    g22348(.A1(new_n22337_), .A2(new_n21772_), .A3(new_n21778_), .ZN(new_n22541_));
  INV_X1     g22349(.I(new_n22541_), .ZN(new_n22542_));
  AOI22_X1   g22350(.A1(new_n22542_), .A2(new_n22116_), .B1(\asqrt[4] ), .B2(new_n22540_), .ZN(new_n22543_));
  NOR2_X1    g22351(.A1(new_n22528_), .A2(\asqrt[28] ), .ZN(new_n22544_));
  AOI21_X1   g22352(.A1(new_n22539_), .A2(new_n22544_), .B(new_n22543_), .ZN(new_n22545_));
  OAI21_X1   g22353(.A1(new_n22545_), .A2(new_n22538_), .B(\asqrt[29] ), .ZN(new_n22546_));
  NOR2_X1    g22354(.A1(new_n21779_), .A2(new_n21787_), .ZN(new_n22547_));
  NOR3_X1    g22355(.A1(new_n22337_), .A2(new_n22188_), .A3(new_n22547_), .ZN(new_n22548_));
  INV_X1     g22356(.I(new_n22548_), .ZN(new_n22549_));
  NOR3_X1    g22357(.A1(new_n22547_), .A2(new_n22188_), .A3(new_n21786_), .ZN(new_n22550_));
  AOI22_X1   g22358(.A1(new_n22549_), .A2(new_n21786_), .B1(\asqrt[4] ), .B2(new_n22550_), .ZN(new_n22551_));
  INV_X1     g22359(.I(new_n22551_), .ZN(new_n22552_));
  NAND2_X1   g22360(.A1(new_n22537_), .A2(new_n8036_), .ZN(new_n22553_));
  OAI21_X1   g22361(.A1(new_n22553_), .A2(new_n22545_), .B(new_n22552_), .ZN(new_n22554_));
  AOI21_X1   g22362(.A1(new_n22554_), .A2(new_n22546_), .B(new_n7539_), .ZN(new_n22555_));
  INV_X1     g22363(.I(new_n22555_), .ZN(new_n22556_));
  INV_X1     g22364(.I(new_n22554_), .ZN(new_n22557_));
  INV_X1     g22365(.I(new_n21793_), .ZN(new_n22558_));
  NOR3_X1    g22366(.A1(new_n21789_), .A2(new_n22197_), .A3(new_n22558_), .ZN(new_n22559_));
  NOR3_X1    g22367(.A1(new_n22337_), .A2(new_n21789_), .A3(new_n22197_), .ZN(new_n22560_));
  INV_X1     g22368(.I(new_n22560_), .ZN(new_n22561_));
  AOI22_X1   g22369(.A1(new_n22561_), .A2(new_n22558_), .B1(\asqrt[4] ), .B2(new_n22559_), .ZN(new_n22562_));
  INV_X1     g22370(.I(new_n22562_), .ZN(new_n22563_));
  NAND2_X1   g22371(.A1(new_n22546_), .A2(new_n7539_), .ZN(new_n22564_));
  OAI21_X1   g22372(.A1(new_n22564_), .A2(new_n22557_), .B(new_n22563_), .ZN(new_n22565_));
  AOI21_X1   g22373(.A1(new_n22565_), .A2(new_n22556_), .B(new_n7229_), .ZN(new_n22566_));
  NOR3_X1    g22374(.A1(new_n22337_), .A2(new_n21798_), .A3(new_n21804_), .ZN(new_n22567_));
  INV_X1     g22375(.I(new_n22567_), .ZN(new_n22568_));
  NOR3_X1    g22376(.A1(new_n21798_), .A2(new_n22115_), .A3(new_n21804_), .ZN(new_n22569_));
  AOI22_X1   g22377(.A1(new_n22568_), .A2(new_n22115_), .B1(\asqrt[4] ), .B2(new_n22569_), .ZN(new_n22570_));
  NOR2_X1    g22378(.A1(new_n22555_), .A2(\asqrt[31] ), .ZN(new_n22571_));
  AOI21_X1   g22379(.A1(new_n22571_), .A2(new_n22565_), .B(new_n22570_), .ZN(new_n22572_));
  OAI21_X1   g22380(.A1(new_n22572_), .A2(new_n22566_), .B(\asqrt[32] ), .ZN(new_n22573_));
  NOR2_X1    g22381(.A1(new_n21805_), .A2(new_n21813_), .ZN(new_n22574_));
  NOR3_X1    g22382(.A1(new_n22574_), .A2(new_n22196_), .A3(new_n21812_), .ZN(new_n22575_));
  NOR3_X1    g22383(.A1(new_n22337_), .A2(new_n22196_), .A3(new_n22574_), .ZN(new_n22576_));
  INV_X1     g22384(.I(new_n22576_), .ZN(new_n22577_));
  AOI22_X1   g22385(.A1(new_n22577_), .A2(new_n21812_), .B1(\asqrt[4] ), .B2(new_n22575_), .ZN(new_n22578_));
  INV_X1     g22386(.I(new_n22578_), .ZN(new_n22579_));
  NOR3_X1    g22387(.A1(new_n22536_), .A2(new_n22528_), .A3(\asqrt[28] ), .ZN(new_n22580_));
  OAI21_X1   g22388(.A1(new_n22543_), .A2(new_n22580_), .B(new_n22537_), .ZN(new_n22581_));
  AOI21_X1   g22389(.A1(new_n22581_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n22582_));
  AOI21_X1   g22390(.A1(new_n22582_), .A2(new_n22554_), .B(new_n22562_), .ZN(new_n22583_));
  OAI21_X1   g22391(.A1(new_n22583_), .A2(new_n22555_), .B(\asqrt[31] ), .ZN(new_n22584_));
  NAND2_X1   g22392(.A1(new_n22584_), .A2(new_n6824_), .ZN(new_n22585_));
  OAI21_X1   g22393(.A1(new_n22585_), .A2(new_n22572_), .B(new_n22579_), .ZN(new_n22586_));
  AOI21_X1   g22394(.A1(new_n22586_), .A2(new_n22573_), .B(new_n6356_), .ZN(new_n22587_));
  INV_X1     g22395(.I(new_n22587_), .ZN(new_n22588_));
  INV_X1     g22396(.I(new_n22586_), .ZN(new_n22589_));
  INV_X1     g22397(.I(new_n21819_), .ZN(new_n22590_));
  NOR3_X1    g22398(.A1(new_n22337_), .A2(new_n21815_), .A3(new_n22205_), .ZN(new_n22591_));
  INV_X1     g22399(.I(new_n22591_), .ZN(new_n22592_));
  NOR3_X1    g22400(.A1(new_n21815_), .A2(new_n22205_), .A3(new_n22590_), .ZN(new_n22593_));
  AOI22_X1   g22401(.A1(new_n22592_), .A2(new_n22590_), .B1(\asqrt[4] ), .B2(new_n22593_), .ZN(new_n22594_));
  INV_X1     g22402(.I(new_n22594_), .ZN(new_n22595_));
  NAND2_X1   g22403(.A1(new_n22573_), .A2(new_n6356_), .ZN(new_n22596_));
  OAI21_X1   g22404(.A1(new_n22596_), .A2(new_n22589_), .B(new_n22595_), .ZN(new_n22597_));
  AOI21_X1   g22405(.A1(new_n22597_), .A2(new_n22588_), .B(new_n6077_), .ZN(new_n22598_));
  NOR3_X1    g22406(.A1(new_n21824_), .A2(new_n22114_), .A3(new_n21830_), .ZN(new_n22599_));
  NOR3_X1    g22407(.A1(new_n22337_), .A2(new_n21824_), .A3(new_n21830_), .ZN(new_n22600_));
  INV_X1     g22408(.I(new_n22600_), .ZN(new_n22601_));
  AOI22_X1   g22409(.A1(new_n22601_), .A2(new_n22114_), .B1(\asqrt[4] ), .B2(new_n22599_), .ZN(new_n22602_));
  NOR2_X1    g22410(.A1(new_n22587_), .A2(\asqrt[34] ), .ZN(new_n22603_));
  AOI21_X1   g22411(.A1(new_n22603_), .A2(new_n22597_), .B(new_n22602_), .ZN(new_n22604_));
  OAI21_X1   g22412(.A1(new_n22604_), .A2(new_n22598_), .B(\asqrt[35] ), .ZN(new_n22605_));
  NOR2_X1    g22413(.A1(new_n21831_), .A2(new_n21839_), .ZN(new_n22606_));
  NOR3_X1    g22414(.A1(new_n22337_), .A2(new_n22204_), .A3(new_n22606_), .ZN(new_n22607_));
  INV_X1     g22415(.I(new_n22607_), .ZN(new_n22608_));
  NOR3_X1    g22416(.A1(new_n22606_), .A2(new_n22204_), .A3(new_n21838_), .ZN(new_n22609_));
  AOI22_X1   g22417(.A1(new_n22608_), .A2(new_n21838_), .B1(\asqrt[4] ), .B2(new_n22609_), .ZN(new_n22610_));
  INV_X1     g22418(.I(new_n22610_), .ZN(new_n22611_));
  NOR3_X1    g22419(.A1(new_n22583_), .A2(\asqrt[31] ), .A3(new_n22555_), .ZN(new_n22612_));
  OAI21_X1   g22420(.A1(new_n22570_), .A2(new_n22612_), .B(new_n22584_), .ZN(new_n22613_));
  AOI21_X1   g22421(.A1(new_n22613_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n22614_));
  AOI21_X1   g22422(.A1(new_n22614_), .A2(new_n22586_), .B(new_n22594_), .ZN(new_n22615_));
  OAI21_X1   g22423(.A1(new_n22615_), .A2(new_n22587_), .B(\asqrt[34] ), .ZN(new_n22616_));
  NAND2_X1   g22424(.A1(new_n22616_), .A2(new_n5708_), .ZN(new_n22617_));
  OAI21_X1   g22425(.A1(new_n22617_), .A2(new_n22604_), .B(new_n22611_), .ZN(new_n22618_));
  NAND2_X1   g22426(.A1(new_n22618_), .A2(new_n22605_), .ZN(new_n22619_));
  NAND2_X1   g22427(.A1(new_n22619_), .A2(\asqrt[36] ), .ZN(new_n22620_));
  INV_X1     g22428(.I(new_n22618_), .ZN(new_n22621_));
  INV_X1     g22429(.I(new_n21845_), .ZN(new_n22622_));
  NOR3_X1    g22430(.A1(new_n21841_), .A2(new_n22213_), .A3(new_n22622_), .ZN(new_n22623_));
  NOR3_X1    g22431(.A1(new_n22337_), .A2(new_n21841_), .A3(new_n22213_), .ZN(new_n22624_));
  INV_X1     g22432(.I(new_n22624_), .ZN(new_n22625_));
  AOI22_X1   g22433(.A1(new_n22625_), .A2(new_n22622_), .B1(\asqrt[4] ), .B2(new_n22623_), .ZN(new_n22626_));
  INV_X1     g22434(.I(new_n22626_), .ZN(new_n22627_));
  NAND2_X1   g22435(.A1(new_n22605_), .A2(new_n5277_), .ZN(new_n22628_));
  OAI21_X1   g22436(.A1(new_n22621_), .A2(new_n22628_), .B(new_n22627_), .ZN(new_n22629_));
  AOI21_X1   g22437(.A1(new_n22629_), .A2(new_n22620_), .B(new_n5024_), .ZN(new_n22630_));
  NOR3_X1    g22438(.A1(new_n22337_), .A2(new_n21850_), .A3(new_n21856_), .ZN(new_n22631_));
  INV_X1     g22439(.I(new_n22631_), .ZN(new_n22632_));
  NOR3_X1    g22440(.A1(new_n21850_), .A2(new_n22113_), .A3(new_n21856_), .ZN(new_n22633_));
  AOI22_X1   g22441(.A1(new_n22632_), .A2(new_n22113_), .B1(\asqrt[4] ), .B2(new_n22633_), .ZN(new_n22634_));
  AOI21_X1   g22442(.A1(new_n22618_), .A2(new_n22605_), .B(new_n5277_), .ZN(new_n22635_));
  NOR2_X1    g22443(.A1(new_n22635_), .A2(\asqrt[37] ), .ZN(new_n22636_));
  AOI21_X1   g22444(.A1(new_n22636_), .A2(new_n22629_), .B(new_n22634_), .ZN(new_n22637_));
  OAI21_X1   g22445(.A1(new_n22637_), .A2(new_n22630_), .B(\asqrt[38] ), .ZN(new_n22638_));
  INV_X1     g22446(.I(new_n22638_), .ZN(new_n22639_));
  NOR2_X1    g22447(.A1(new_n21857_), .A2(new_n21865_), .ZN(new_n22640_));
  NOR3_X1    g22448(.A1(new_n22640_), .A2(new_n22212_), .A3(new_n21864_), .ZN(new_n22641_));
  NOR3_X1    g22449(.A1(new_n22337_), .A2(new_n22212_), .A3(new_n22640_), .ZN(new_n22642_));
  INV_X1     g22450(.I(new_n22642_), .ZN(new_n22643_));
  AOI22_X1   g22451(.A1(new_n22643_), .A2(new_n21864_), .B1(\asqrt[4] ), .B2(new_n22641_), .ZN(new_n22644_));
  NOR3_X1    g22452(.A1(new_n22637_), .A2(new_n22630_), .A3(\asqrt[38] ), .ZN(new_n22645_));
  NOR2_X1    g22453(.A1(new_n22645_), .A2(new_n22644_), .ZN(new_n22646_));
  OAI21_X1   g22454(.A1(new_n22646_), .A2(new_n22639_), .B(\asqrt[39] ), .ZN(new_n22647_));
  INV_X1     g22455(.I(new_n21871_), .ZN(new_n22648_));
  NOR3_X1    g22456(.A1(new_n22337_), .A2(new_n21867_), .A3(new_n22221_), .ZN(new_n22649_));
  INV_X1     g22457(.I(new_n22649_), .ZN(new_n22650_));
  NOR3_X1    g22458(.A1(new_n21867_), .A2(new_n22221_), .A3(new_n22648_), .ZN(new_n22651_));
  AOI22_X1   g22459(.A1(new_n22650_), .A2(new_n22648_), .B1(\asqrt[4] ), .B2(new_n22651_), .ZN(new_n22652_));
  INV_X1     g22460(.I(new_n22652_), .ZN(new_n22653_));
  NAND2_X1   g22461(.A1(new_n22638_), .A2(new_n4298_), .ZN(new_n22654_));
  OAI21_X1   g22462(.A1(new_n22646_), .A2(new_n22654_), .B(new_n22653_), .ZN(new_n22655_));
  AOI21_X1   g22463(.A1(new_n22655_), .A2(new_n22647_), .B(new_n4071_), .ZN(new_n22656_));
  NOR3_X1    g22464(.A1(new_n21876_), .A2(new_n22112_), .A3(new_n21882_), .ZN(new_n22657_));
  NOR3_X1    g22465(.A1(new_n22337_), .A2(new_n21876_), .A3(new_n21882_), .ZN(new_n22658_));
  INV_X1     g22466(.I(new_n22658_), .ZN(new_n22659_));
  AOI22_X1   g22467(.A1(new_n22659_), .A2(new_n22112_), .B1(\asqrt[4] ), .B2(new_n22657_), .ZN(new_n22660_));
  INV_X1     g22468(.I(new_n22644_), .ZN(new_n22661_));
  NOR3_X1    g22469(.A1(new_n22615_), .A2(\asqrt[34] ), .A3(new_n22587_), .ZN(new_n22662_));
  OAI21_X1   g22470(.A1(new_n22602_), .A2(new_n22662_), .B(new_n22616_), .ZN(new_n22663_));
  AOI21_X1   g22471(.A1(new_n22663_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n22664_));
  AOI21_X1   g22472(.A1(new_n22664_), .A2(new_n22618_), .B(new_n22626_), .ZN(new_n22665_));
  OAI21_X1   g22473(.A1(new_n22665_), .A2(new_n22635_), .B(\asqrt[37] ), .ZN(new_n22666_));
  NAND2_X1   g22474(.A1(new_n22666_), .A2(new_n4696_), .ZN(new_n22667_));
  OAI21_X1   g22475(.A1(new_n22667_), .A2(new_n22637_), .B(new_n22661_), .ZN(new_n22668_));
  AOI21_X1   g22476(.A1(new_n22668_), .A2(new_n22638_), .B(new_n4298_), .ZN(new_n22669_));
  NOR2_X1    g22477(.A1(new_n22669_), .A2(\asqrt[40] ), .ZN(new_n22670_));
  AOI21_X1   g22478(.A1(new_n22670_), .A2(new_n22655_), .B(new_n22660_), .ZN(new_n22671_));
  OAI21_X1   g22479(.A1(new_n22671_), .A2(new_n22656_), .B(\asqrt[41] ), .ZN(new_n22672_));
  NOR2_X1    g22480(.A1(new_n21883_), .A2(new_n21891_), .ZN(new_n22673_));
  NOR3_X1    g22481(.A1(new_n22337_), .A2(new_n22220_), .A3(new_n22673_), .ZN(new_n22674_));
  INV_X1     g22482(.I(new_n22674_), .ZN(new_n22675_));
  NOR3_X1    g22483(.A1(new_n22673_), .A2(new_n22220_), .A3(new_n21890_), .ZN(new_n22676_));
  AOI22_X1   g22484(.A1(new_n22675_), .A2(new_n21890_), .B1(\asqrt[4] ), .B2(new_n22676_), .ZN(new_n22677_));
  INV_X1     g22485(.I(new_n22677_), .ZN(new_n22678_));
  NOR3_X1    g22486(.A1(new_n22665_), .A2(\asqrt[37] ), .A3(new_n22635_), .ZN(new_n22679_));
  OAI21_X1   g22487(.A1(new_n22634_), .A2(new_n22679_), .B(new_n22666_), .ZN(new_n22680_));
  AOI21_X1   g22488(.A1(new_n22680_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n22681_));
  AOI21_X1   g22489(.A1(new_n22681_), .A2(new_n22668_), .B(new_n22652_), .ZN(new_n22682_));
  OAI21_X1   g22490(.A1(new_n22682_), .A2(new_n22669_), .B(\asqrt[40] ), .ZN(new_n22683_));
  NAND2_X1   g22491(.A1(new_n22683_), .A2(new_n3782_), .ZN(new_n22684_));
  OAI21_X1   g22492(.A1(new_n22684_), .A2(new_n22671_), .B(new_n22678_), .ZN(new_n22685_));
  AOI21_X1   g22493(.A1(new_n22685_), .A2(new_n22672_), .B(new_n3419_), .ZN(new_n22686_));
  INV_X1     g22494(.I(new_n21897_), .ZN(new_n22687_));
  NOR3_X1    g22495(.A1(new_n21893_), .A2(new_n22229_), .A3(new_n22687_), .ZN(new_n22688_));
  NOR3_X1    g22496(.A1(new_n22337_), .A2(new_n21893_), .A3(new_n22229_), .ZN(new_n22689_));
  INV_X1     g22497(.I(new_n22689_), .ZN(new_n22690_));
  AOI22_X1   g22498(.A1(new_n22690_), .A2(new_n22687_), .B1(\asqrt[4] ), .B2(new_n22688_), .ZN(new_n22691_));
  NOR3_X1    g22499(.A1(new_n22682_), .A2(\asqrt[40] ), .A3(new_n22669_), .ZN(new_n22692_));
  OAI21_X1   g22500(.A1(new_n22660_), .A2(new_n22692_), .B(new_n22683_), .ZN(new_n22693_));
  AOI21_X1   g22501(.A1(new_n22693_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n22694_));
  AOI21_X1   g22502(.A1(new_n22694_), .A2(new_n22685_), .B(new_n22691_), .ZN(new_n22695_));
  OAI21_X1   g22503(.A1(new_n22695_), .A2(new_n22686_), .B(\asqrt[43] ), .ZN(new_n22696_));
  INV_X1     g22504(.I(new_n22696_), .ZN(new_n22697_));
  NOR3_X1    g22505(.A1(new_n22337_), .A2(new_n21902_), .A3(new_n21908_), .ZN(new_n22698_));
  INV_X1     g22506(.I(new_n22698_), .ZN(new_n22699_));
  NOR3_X1    g22507(.A1(new_n21902_), .A2(new_n22111_), .A3(new_n21908_), .ZN(new_n22700_));
  AOI22_X1   g22508(.A1(new_n22699_), .A2(new_n22111_), .B1(\asqrt[4] ), .B2(new_n22700_), .ZN(new_n22701_));
  NOR3_X1    g22509(.A1(new_n22695_), .A2(\asqrt[43] ), .A3(new_n22686_), .ZN(new_n22702_));
  NOR2_X1    g22510(.A1(new_n22702_), .A2(new_n22701_), .ZN(new_n22703_));
  OAI21_X1   g22511(.A1(new_n22703_), .A2(new_n22697_), .B(\asqrt[44] ), .ZN(new_n22704_));
  NOR2_X1    g22512(.A1(new_n21909_), .A2(new_n21917_), .ZN(new_n22705_));
  NOR3_X1    g22513(.A1(new_n22705_), .A2(new_n22228_), .A3(new_n21916_), .ZN(new_n22706_));
  NOR3_X1    g22514(.A1(new_n22337_), .A2(new_n22228_), .A3(new_n22705_), .ZN(new_n22707_));
  INV_X1     g22515(.I(new_n22707_), .ZN(new_n22708_));
  AOI22_X1   g22516(.A1(new_n22708_), .A2(new_n21916_), .B1(\asqrt[4] ), .B2(new_n22706_), .ZN(new_n22709_));
  INV_X1     g22517(.I(new_n22709_), .ZN(new_n22710_));
  NAND2_X1   g22518(.A1(new_n22696_), .A2(new_n2954_), .ZN(new_n22711_));
  OAI21_X1   g22519(.A1(new_n22703_), .A2(new_n22711_), .B(new_n22710_), .ZN(new_n22712_));
  AOI21_X1   g22520(.A1(new_n22712_), .A2(new_n22704_), .B(new_n2641_), .ZN(new_n22713_));
  INV_X1     g22521(.I(new_n21923_), .ZN(new_n22714_));
  NOR3_X1    g22522(.A1(new_n22337_), .A2(new_n21919_), .A3(new_n22237_), .ZN(new_n22715_));
  INV_X1     g22523(.I(new_n22715_), .ZN(new_n22716_));
  NOR3_X1    g22524(.A1(new_n21919_), .A2(new_n22237_), .A3(new_n22714_), .ZN(new_n22717_));
  AOI22_X1   g22525(.A1(new_n22716_), .A2(new_n22714_), .B1(\asqrt[4] ), .B2(new_n22717_), .ZN(new_n22718_));
  OAI21_X1   g22526(.A1(new_n22701_), .A2(new_n22702_), .B(new_n22696_), .ZN(new_n22719_));
  AOI21_X1   g22527(.A1(new_n22719_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n22720_));
  AOI21_X1   g22528(.A1(new_n22720_), .A2(new_n22712_), .B(new_n22718_), .ZN(new_n22721_));
  OAI21_X1   g22529(.A1(new_n22721_), .A2(new_n22713_), .B(\asqrt[46] ), .ZN(new_n22722_));
  INV_X1     g22530(.I(new_n22722_), .ZN(new_n22723_));
  NOR3_X1    g22531(.A1(new_n21928_), .A2(new_n22110_), .A3(new_n21934_), .ZN(new_n22724_));
  NOR3_X1    g22532(.A1(new_n22337_), .A2(new_n21928_), .A3(new_n21934_), .ZN(new_n22725_));
  INV_X1     g22533(.I(new_n22725_), .ZN(new_n22726_));
  AOI22_X1   g22534(.A1(new_n22726_), .A2(new_n22110_), .B1(\asqrt[4] ), .B2(new_n22724_), .ZN(new_n22727_));
  NOR3_X1    g22535(.A1(new_n22721_), .A2(new_n22713_), .A3(\asqrt[46] ), .ZN(new_n22728_));
  NOR2_X1    g22536(.A1(new_n22728_), .A2(new_n22727_), .ZN(new_n22729_));
  OAI21_X1   g22537(.A1(new_n22729_), .A2(new_n22723_), .B(\asqrt[47] ), .ZN(new_n22730_));
  NOR2_X1    g22538(.A1(new_n21935_), .A2(new_n21943_), .ZN(new_n22731_));
  NOR3_X1    g22539(.A1(new_n22337_), .A2(new_n22236_), .A3(new_n22731_), .ZN(new_n22732_));
  INV_X1     g22540(.I(new_n22732_), .ZN(new_n22733_));
  NOR3_X1    g22541(.A1(new_n22731_), .A2(new_n22236_), .A3(new_n21942_), .ZN(new_n22734_));
  AOI22_X1   g22542(.A1(new_n22733_), .A2(new_n21942_), .B1(\asqrt[4] ), .B2(new_n22734_), .ZN(new_n22735_));
  INV_X1     g22543(.I(new_n22735_), .ZN(new_n22736_));
  NAND2_X1   g22544(.A1(new_n22722_), .A2(new_n2229_), .ZN(new_n22737_));
  OAI21_X1   g22545(.A1(new_n22729_), .A2(new_n22737_), .B(new_n22736_), .ZN(new_n22738_));
  AOI21_X1   g22546(.A1(new_n22738_), .A2(new_n22730_), .B(new_n1956_), .ZN(new_n22739_));
  INV_X1     g22547(.I(new_n21949_), .ZN(new_n22740_));
  NOR3_X1    g22548(.A1(new_n21945_), .A2(new_n22245_), .A3(new_n22740_), .ZN(new_n22741_));
  NOR3_X1    g22549(.A1(new_n22337_), .A2(new_n21945_), .A3(new_n22245_), .ZN(new_n22742_));
  INV_X1     g22550(.I(new_n22742_), .ZN(new_n22743_));
  AOI22_X1   g22551(.A1(new_n22743_), .A2(new_n22740_), .B1(\asqrt[4] ), .B2(new_n22741_), .ZN(new_n22744_));
  OAI21_X1   g22552(.A1(new_n22727_), .A2(new_n22728_), .B(new_n22722_), .ZN(new_n22745_));
  AOI21_X1   g22553(.A1(new_n22745_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n22746_));
  AOI21_X1   g22554(.A1(new_n22746_), .A2(new_n22738_), .B(new_n22744_), .ZN(new_n22747_));
  OAI21_X1   g22555(.A1(new_n22747_), .A2(new_n22739_), .B(\asqrt[49] ), .ZN(new_n22748_));
  INV_X1     g22556(.I(new_n22748_), .ZN(new_n22749_));
  NOR3_X1    g22557(.A1(new_n22337_), .A2(new_n21954_), .A3(new_n21960_), .ZN(new_n22750_));
  INV_X1     g22558(.I(new_n22750_), .ZN(new_n22751_));
  NOR3_X1    g22559(.A1(new_n21954_), .A2(new_n22109_), .A3(new_n21960_), .ZN(new_n22752_));
  AOI22_X1   g22560(.A1(new_n22751_), .A2(new_n22109_), .B1(\asqrt[4] ), .B2(new_n22752_), .ZN(new_n22753_));
  NOR3_X1    g22561(.A1(new_n22747_), .A2(new_n22739_), .A3(\asqrt[49] ), .ZN(new_n22754_));
  NOR2_X1    g22562(.A1(new_n22754_), .A2(new_n22753_), .ZN(new_n22755_));
  OAI21_X1   g22563(.A1(new_n22755_), .A2(new_n22749_), .B(\asqrt[50] ), .ZN(new_n22756_));
  NOR2_X1    g22564(.A1(new_n21961_), .A2(new_n21969_), .ZN(new_n22757_));
  NOR3_X1    g22565(.A1(new_n22757_), .A2(new_n22244_), .A3(new_n21968_), .ZN(new_n22758_));
  NOR3_X1    g22566(.A1(new_n22337_), .A2(new_n22244_), .A3(new_n22757_), .ZN(new_n22759_));
  INV_X1     g22567(.I(new_n22759_), .ZN(new_n22760_));
  AOI22_X1   g22568(.A1(new_n22760_), .A2(new_n21968_), .B1(\asqrt[4] ), .B2(new_n22758_), .ZN(new_n22761_));
  INV_X1     g22569(.I(new_n22761_), .ZN(new_n22762_));
  NAND2_X1   g22570(.A1(new_n22748_), .A2(new_n1612_), .ZN(new_n22763_));
  OAI21_X1   g22571(.A1(new_n22755_), .A2(new_n22763_), .B(new_n22762_), .ZN(new_n22764_));
  AOI21_X1   g22572(.A1(new_n22764_), .A2(new_n22756_), .B(new_n1376_), .ZN(new_n22765_));
  INV_X1     g22573(.I(new_n21975_), .ZN(new_n22766_));
  NOR3_X1    g22574(.A1(new_n22337_), .A2(new_n21971_), .A3(new_n22253_), .ZN(new_n22767_));
  INV_X1     g22575(.I(new_n22767_), .ZN(new_n22768_));
  NOR3_X1    g22576(.A1(new_n21971_), .A2(new_n22253_), .A3(new_n22766_), .ZN(new_n22769_));
  AOI22_X1   g22577(.A1(new_n22768_), .A2(new_n22766_), .B1(\asqrt[4] ), .B2(new_n22769_), .ZN(new_n22770_));
  OAI21_X1   g22578(.A1(new_n22753_), .A2(new_n22754_), .B(new_n22748_), .ZN(new_n22771_));
  AOI21_X1   g22579(.A1(new_n22771_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n22772_));
  AOI21_X1   g22580(.A1(new_n22772_), .A2(new_n22764_), .B(new_n22770_), .ZN(new_n22773_));
  OAI21_X1   g22581(.A1(new_n22773_), .A2(new_n22765_), .B(\asqrt[52] ), .ZN(new_n22774_));
  INV_X1     g22582(.I(new_n22774_), .ZN(new_n22775_));
  INV_X1     g22583(.I(new_n22773_), .ZN(new_n22776_));
  NOR3_X1    g22584(.A1(new_n21980_), .A2(new_n22108_), .A3(new_n21986_), .ZN(new_n22777_));
  NOR3_X1    g22585(.A1(new_n22337_), .A2(new_n21980_), .A3(new_n21986_), .ZN(new_n22778_));
  INV_X1     g22586(.I(new_n22778_), .ZN(new_n22779_));
  AOI22_X1   g22587(.A1(new_n22779_), .A2(new_n22108_), .B1(\asqrt[4] ), .B2(new_n22777_), .ZN(new_n22780_));
  NOR2_X1    g22588(.A1(new_n22765_), .A2(\asqrt[52] ), .ZN(new_n22781_));
  AOI21_X1   g22589(.A1(new_n22776_), .A2(new_n22781_), .B(new_n22780_), .ZN(new_n22782_));
  OAI21_X1   g22590(.A1(new_n22782_), .A2(new_n22775_), .B(\asqrt[53] ), .ZN(new_n22783_));
  NOR2_X1    g22591(.A1(new_n21987_), .A2(new_n21997_), .ZN(new_n22784_));
  NOR3_X1    g22592(.A1(new_n22337_), .A2(new_n22252_), .A3(new_n22784_), .ZN(new_n22785_));
  INV_X1     g22593(.I(new_n22785_), .ZN(new_n22786_));
  NOR3_X1    g22594(.A1(new_n22784_), .A2(new_n22252_), .A3(new_n21996_), .ZN(new_n22787_));
  AOI22_X1   g22595(.A1(new_n22786_), .A2(new_n21996_), .B1(\asqrt[4] ), .B2(new_n22787_), .ZN(new_n22788_));
  INV_X1     g22596(.I(new_n22788_), .ZN(new_n22789_));
  NAND2_X1   g22597(.A1(new_n22774_), .A2(new_n1103_), .ZN(new_n22790_));
  OAI21_X1   g22598(.A1(new_n22790_), .A2(new_n22782_), .B(new_n22789_), .ZN(new_n22791_));
  AOI21_X1   g22599(.A1(new_n22791_), .A2(new_n22783_), .B(new_n904_), .ZN(new_n22792_));
  INV_X1     g22600(.I(new_n22792_), .ZN(new_n22793_));
  INV_X1     g22601(.I(new_n22791_), .ZN(new_n22794_));
  INV_X1     g22602(.I(new_n22003_), .ZN(new_n22795_));
  NOR3_X1    g22603(.A1(new_n21999_), .A2(new_n22261_), .A3(new_n22795_), .ZN(new_n22796_));
  NOR3_X1    g22604(.A1(new_n22337_), .A2(new_n21999_), .A3(new_n22261_), .ZN(new_n22797_));
  INV_X1     g22605(.I(new_n22797_), .ZN(new_n22798_));
  AOI22_X1   g22606(.A1(new_n22798_), .A2(new_n22795_), .B1(\asqrt[4] ), .B2(new_n22796_), .ZN(new_n22799_));
  INV_X1     g22607(.I(new_n22799_), .ZN(new_n22800_));
  NAND2_X1   g22608(.A1(new_n22783_), .A2(new_n904_), .ZN(new_n22801_));
  OAI21_X1   g22609(.A1(new_n22801_), .A2(new_n22794_), .B(new_n22800_), .ZN(new_n22802_));
  AOI21_X1   g22610(.A1(new_n22802_), .A2(new_n22793_), .B(new_n823_), .ZN(new_n22803_));
  NOR3_X1    g22611(.A1(new_n22337_), .A2(new_n22008_), .A3(new_n22015_), .ZN(new_n22804_));
  INV_X1     g22612(.I(new_n22804_), .ZN(new_n22805_));
  NOR3_X1    g22613(.A1(new_n22008_), .A2(new_n22107_), .A3(new_n22015_), .ZN(new_n22806_));
  AOI22_X1   g22614(.A1(new_n22805_), .A2(new_n22107_), .B1(\asqrt[4] ), .B2(new_n22806_), .ZN(new_n22807_));
  NOR2_X1    g22615(.A1(new_n22792_), .A2(\asqrt[55] ), .ZN(new_n22808_));
  AOI21_X1   g22616(.A1(new_n22808_), .A2(new_n22802_), .B(new_n22807_), .ZN(new_n22809_));
  OAI21_X1   g22617(.A1(new_n22809_), .A2(new_n22803_), .B(\asqrt[56] ), .ZN(new_n22810_));
  NOR2_X1    g22618(.A1(new_n22016_), .A2(new_n22028_), .ZN(new_n22811_));
  NOR3_X1    g22619(.A1(new_n22811_), .A2(new_n22260_), .A3(new_n22027_), .ZN(new_n22812_));
  NOR3_X1    g22620(.A1(new_n22337_), .A2(new_n22260_), .A3(new_n22811_), .ZN(new_n22813_));
  INV_X1     g22621(.I(new_n22813_), .ZN(new_n22814_));
  AOI22_X1   g22622(.A1(new_n22814_), .A2(new_n22027_), .B1(\asqrt[4] ), .B2(new_n22812_), .ZN(new_n22815_));
  INV_X1     g22623(.I(new_n22815_), .ZN(new_n22816_));
  NOR3_X1    g22624(.A1(new_n22773_), .A2(new_n22765_), .A3(\asqrt[52] ), .ZN(new_n22817_));
  OAI21_X1   g22625(.A1(new_n22780_), .A2(new_n22817_), .B(new_n22774_), .ZN(new_n22818_));
  AOI21_X1   g22626(.A1(new_n22818_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n22819_));
  AOI21_X1   g22627(.A1(new_n22819_), .A2(new_n22791_), .B(new_n22799_), .ZN(new_n22820_));
  OAI21_X1   g22628(.A1(new_n22820_), .A2(new_n22792_), .B(\asqrt[55] ), .ZN(new_n22821_));
  NAND2_X1   g22629(.A1(new_n22821_), .A2(new_n703_), .ZN(new_n22822_));
  OAI21_X1   g22630(.A1(new_n22822_), .A2(new_n22809_), .B(new_n22816_), .ZN(new_n22823_));
  AOI21_X1   g22631(.A1(new_n22823_), .A2(new_n22810_), .B(new_n531_), .ZN(new_n22824_));
  INV_X1     g22632(.I(new_n22824_), .ZN(new_n22825_));
  INV_X1     g22633(.I(new_n22823_), .ZN(new_n22826_));
  INV_X1     g22634(.I(new_n22034_), .ZN(new_n22827_));
  NOR3_X1    g22635(.A1(new_n22337_), .A2(new_n22030_), .A3(new_n22269_), .ZN(new_n22828_));
  INV_X1     g22636(.I(new_n22828_), .ZN(new_n22829_));
  NOR3_X1    g22637(.A1(new_n22030_), .A2(new_n22269_), .A3(new_n22827_), .ZN(new_n22830_));
  AOI22_X1   g22638(.A1(new_n22829_), .A2(new_n22827_), .B1(\asqrt[4] ), .B2(new_n22830_), .ZN(new_n22831_));
  INV_X1     g22639(.I(new_n22831_), .ZN(new_n22832_));
  NAND2_X1   g22640(.A1(new_n22810_), .A2(new_n531_), .ZN(new_n22833_));
  OAI21_X1   g22641(.A1(new_n22833_), .A2(new_n22826_), .B(new_n22832_), .ZN(new_n22834_));
  AOI21_X1   g22642(.A1(new_n22834_), .A2(new_n22825_), .B(new_n436_), .ZN(new_n22835_));
  NOR3_X1    g22643(.A1(new_n22039_), .A2(new_n22106_), .A3(new_n22046_), .ZN(new_n22836_));
  NOR3_X1    g22644(.A1(new_n22337_), .A2(new_n22039_), .A3(new_n22046_), .ZN(new_n22837_));
  INV_X1     g22645(.I(new_n22837_), .ZN(new_n22838_));
  AOI22_X1   g22646(.A1(new_n22838_), .A2(new_n22106_), .B1(\asqrt[4] ), .B2(new_n22836_), .ZN(new_n22839_));
  NOR2_X1    g22647(.A1(new_n22824_), .A2(\asqrt[58] ), .ZN(new_n22840_));
  AOI21_X1   g22648(.A1(new_n22840_), .A2(new_n22834_), .B(new_n22839_), .ZN(new_n22841_));
  OAI21_X1   g22649(.A1(new_n22841_), .A2(new_n22835_), .B(\asqrt[59] ), .ZN(new_n22842_));
  NOR2_X1    g22650(.A1(new_n22047_), .A2(new_n22058_), .ZN(new_n22843_));
  NOR3_X1    g22651(.A1(new_n22337_), .A2(new_n22268_), .A3(new_n22843_), .ZN(new_n22844_));
  INV_X1     g22652(.I(new_n22844_), .ZN(new_n22845_));
  NOR3_X1    g22653(.A1(new_n22843_), .A2(new_n22268_), .A3(new_n22057_), .ZN(new_n22846_));
  AOI22_X1   g22654(.A1(new_n22845_), .A2(new_n22057_), .B1(\asqrt[4] ), .B2(new_n22846_), .ZN(new_n22847_));
  INV_X1     g22655(.I(new_n22847_), .ZN(new_n22848_));
  NOR3_X1    g22656(.A1(new_n22820_), .A2(\asqrt[55] ), .A3(new_n22792_), .ZN(new_n22849_));
  OAI21_X1   g22657(.A1(new_n22807_), .A2(new_n22849_), .B(new_n22821_), .ZN(new_n22850_));
  AOI21_X1   g22658(.A1(new_n22850_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n22851_));
  AOI21_X1   g22659(.A1(new_n22851_), .A2(new_n22823_), .B(new_n22831_), .ZN(new_n22852_));
  OAI21_X1   g22660(.A1(new_n22852_), .A2(new_n22824_), .B(\asqrt[58] ), .ZN(new_n22853_));
  NAND2_X1   g22661(.A1(new_n22853_), .A2(new_n327_), .ZN(new_n22854_));
  OAI21_X1   g22662(.A1(new_n22854_), .A2(new_n22841_), .B(new_n22848_), .ZN(new_n22855_));
  AOI21_X1   g22663(.A1(new_n22855_), .A2(new_n22842_), .B(new_n306_), .ZN(new_n22856_));
  INV_X1     g22664(.I(new_n22856_), .ZN(new_n22857_));
  INV_X1     g22665(.I(new_n22855_), .ZN(new_n22858_));
  INV_X1     g22666(.I(new_n22064_), .ZN(new_n22859_));
  NOR3_X1    g22667(.A1(new_n22060_), .A2(new_n22276_), .A3(new_n22859_), .ZN(new_n22860_));
  NOR3_X1    g22668(.A1(new_n22337_), .A2(new_n22060_), .A3(new_n22276_), .ZN(new_n22861_));
  INV_X1     g22669(.I(new_n22861_), .ZN(new_n22862_));
  AOI22_X1   g22670(.A1(new_n22862_), .A2(new_n22859_), .B1(\asqrt[4] ), .B2(new_n22860_), .ZN(new_n22863_));
  INV_X1     g22671(.I(new_n22863_), .ZN(new_n22864_));
  NAND2_X1   g22672(.A1(new_n22842_), .A2(new_n306_), .ZN(new_n22865_));
  OAI21_X1   g22673(.A1(new_n22858_), .A2(new_n22865_), .B(new_n22864_), .ZN(new_n22866_));
  AOI21_X1   g22674(.A1(new_n22866_), .A2(new_n22857_), .B(new_n218_), .ZN(new_n22867_));
  NOR3_X1    g22675(.A1(new_n22337_), .A2(new_n22069_), .A3(new_n22075_), .ZN(new_n22868_));
  INV_X1     g22676(.I(new_n22868_), .ZN(new_n22869_));
  NOR3_X1    g22677(.A1(new_n22069_), .A2(new_n22105_), .A3(new_n22075_), .ZN(new_n22870_));
  AOI22_X1   g22678(.A1(new_n22869_), .A2(new_n22105_), .B1(\asqrt[4] ), .B2(new_n22870_), .ZN(new_n22871_));
  NOR2_X1    g22679(.A1(new_n22856_), .A2(\asqrt[61] ), .ZN(new_n22872_));
  AOI21_X1   g22680(.A1(new_n22872_), .A2(new_n22866_), .B(new_n22871_), .ZN(new_n22873_));
  OAI21_X1   g22681(.A1(new_n22873_), .A2(new_n22867_), .B(\asqrt[62] ), .ZN(new_n22874_));
  NOR2_X1    g22682(.A1(new_n22076_), .A2(new_n22083_), .ZN(new_n22875_));
  NOR3_X1    g22683(.A1(new_n22875_), .A2(new_n22294_), .A3(new_n22082_), .ZN(new_n22876_));
  NOR3_X1    g22684(.A1(new_n22337_), .A2(new_n22294_), .A3(new_n22875_), .ZN(new_n22877_));
  INV_X1     g22685(.I(new_n22877_), .ZN(new_n22878_));
  AOI22_X1   g22686(.A1(new_n22878_), .A2(new_n22082_), .B1(\asqrt[4] ), .B2(new_n22876_), .ZN(new_n22879_));
  INV_X1     g22687(.I(new_n22879_), .ZN(new_n22880_));
  NOR3_X1    g22688(.A1(new_n22852_), .A2(\asqrt[58] ), .A3(new_n22824_), .ZN(new_n22881_));
  OAI21_X1   g22689(.A1(new_n22839_), .A2(new_n22881_), .B(new_n22853_), .ZN(new_n22882_));
  AOI21_X1   g22690(.A1(new_n22882_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n22883_));
  AOI21_X1   g22691(.A1(new_n22883_), .A2(new_n22855_), .B(new_n22863_), .ZN(new_n22884_));
  OAI21_X1   g22692(.A1(new_n22884_), .A2(new_n22856_), .B(\asqrt[61] ), .ZN(new_n22885_));
  NAND2_X1   g22693(.A1(new_n22885_), .A2(new_n207_), .ZN(new_n22886_));
  OAI21_X1   g22694(.A1(new_n22886_), .A2(new_n22873_), .B(new_n22880_), .ZN(new_n22887_));
  INV_X1     g22695(.I(new_n22296_), .ZN(new_n22888_));
  NAND2_X1   g22696(.A1(new_n22888_), .A2(new_n22295_), .ZN(new_n22889_));
  OAI21_X1   g22697(.A1(new_n22337_), .A2(new_n22889_), .B(new_n22280_), .ZN(new_n22890_));
  NAND4_X1   g22698(.A1(\asqrt[4] ), .A2(new_n22295_), .A3(new_n22089_), .A4(new_n22888_), .ZN(new_n22891_));
  NAND2_X1   g22699(.A1(new_n22890_), .A2(new_n22891_), .ZN(new_n22892_));
  INV_X1     g22700(.I(new_n22297_), .ZN(new_n22893_));
  NOR2_X1    g22701(.A1(new_n22893_), .A2(new_n22098_), .ZN(new_n22894_));
  AOI21_X1   g22702(.A1(\asqrt[4] ), .A2(new_n22894_), .B(new_n22313_), .ZN(new_n22895_));
  NAND2_X1   g22703(.A1(new_n22892_), .A2(new_n22895_), .ZN(new_n22896_));
  AOI21_X1   g22704(.A1(new_n22887_), .A2(new_n22874_), .B(new_n22896_), .ZN(new_n22897_));
  NOR2_X1    g22705(.A1(new_n22897_), .A2(\asqrt[63] ), .ZN(new_n22898_));
  INV_X1     g22706(.I(new_n22887_), .ZN(new_n22899_));
  INV_X1     g22707(.I(new_n22892_), .ZN(new_n22900_));
  NAND2_X1   g22708(.A1(new_n22874_), .A2(new_n22900_), .ZN(new_n22901_));
  OAI21_X1   g22709(.A1(new_n22337_), .A2(new_n22098_), .B(new_n22893_), .ZN(new_n22902_));
  NOR2_X1    g22710(.A1(new_n22894_), .A2(new_n193_), .ZN(new_n22903_));
  NAND2_X1   g22711(.A1(new_n22902_), .A2(new_n22903_), .ZN(new_n22904_));
  OAI21_X1   g22712(.A1(new_n22899_), .A2(new_n22901_), .B(new_n22904_), .ZN(new_n22905_));
  NOR2_X1    g22713(.A1(new_n22898_), .A2(new_n22905_), .ZN(new_n22906_));
  INV_X1     g22714(.I(\a[4] ), .ZN(new_n22907_));
  NOR2_X1    g22715(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n22908_));
  INV_X1     g22716(.I(new_n22908_), .ZN(new_n22909_));
  NOR2_X1    g22717(.A1(new_n22909_), .A2(\a[4] ), .ZN(new_n22910_));
  INV_X1     g22718(.I(new_n22910_), .ZN(new_n22911_));
  INV_X1     g22719(.I(\a[6] ), .ZN(new_n22912_));
  NOR2_X1    g22720(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n22913_));
  INV_X1     g22721(.I(new_n22913_), .ZN(new_n22914_));
  NOR2_X1    g22722(.A1(new_n22914_), .A2(\a[6] ), .ZN(new_n22915_));
  INV_X1     g22723(.I(new_n22915_), .ZN(new_n22916_));
  OAI21_X1   g22724(.A1(new_n22906_), .A2(new_n22912_), .B(new_n22916_), .ZN(new_n22917_));
  NOR4_X1    g22725(.A1(new_n22298_), .A2(new_n22313_), .A3(new_n22287_), .A4(new_n22915_), .ZN(new_n22918_));
  OAI21_X1   g22726(.A1(new_n22906_), .A2(new_n22912_), .B(new_n22918_), .ZN(new_n22919_));
  NOR3_X1    g22727(.A1(new_n22884_), .A2(\asqrt[61] ), .A3(new_n22856_), .ZN(new_n22920_));
  OAI21_X1   g22728(.A1(new_n22871_), .A2(new_n22920_), .B(new_n22885_), .ZN(new_n22921_));
  INV_X1     g22729(.I(new_n22871_), .ZN(new_n22922_));
  INV_X1     g22730(.I(new_n22839_), .ZN(new_n22923_));
  INV_X1     g22731(.I(new_n22807_), .ZN(new_n22924_));
  INV_X1     g22732(.I(new_n22780_), .ZN(new_n22925_));
  INV_X1     g22733(.I(new_n22753_), .ZN(new_n22926_));
  INV_X1     g22734(.I(new_n22727_), .ZN(new_n22927_));
  INV_X1     g22735(.I(new_n22701_), .ZN(new_n22928_));
  INV_X1     g22736(.I(new_n22672_), .ZN(new_n22929_));
  NOR3_X1    g22737(.A1(new_n22671_), .A2(new_n22656_), .A3(\asqrt[41] ), .ZN(new_n22930_));
  NOR2_X1    g22738(.A1(new_n22930_), .A2(new_n22677_), .ZN(new_n22931_));
  OAI21_X1   g22739(.A1(new_n22931_), .A2(new_n22929_), .B(\asqrt[42] ), .ZN(new_n22932_));
  NAND2_X1   g22740(.A1(new_n22932_), .A2(new_n3218_), .ZN(new_n22933_));
  OAI21_X1   g22741(.A1(new_n22933_), .A2(new_n22695_), .B(new_n22928_), .ZN(new_n22934_));
  NAND3_X1   g22742(.A1(new_n22934_), .A2(new_n2954_), .A3(new_n22696_), .ZN(new_n22935_));
  AOI22_X1   g22743(.A1(new_n22935_), .A2(new_n22710_), .B1(\asqrt[44] ), .B2(new_n22719_), .ZN(new_n22936_));
  OAI21_X1   g22744(.A1(new_n22936_), .A2(new_n2641_), .B(new_n2465_), .ZN(new_n22937_));
  OAI21_X1   g22745(.A1(new_n22937_), .A2(new_n22721_), .B(new_n22927_), .ZN(new_n22938_));
  NAND3_X1   g22746(.A1(new_n22938_), .A2(new_n2229_), .A3(new_n22722_), .ZN(new_n22939_));
  AOI22_X1   g22747(.A1(new_n22939_), .A2(new_n22736_), .B1(\asqrt[47] ), .B2(new_n22745_), .ZN(new_n22940_));
  OAI21_X1   g22748(.A1(new_n22940_), .A2(new_n1956_), .B(new_n1806_), .ZN(new_n22941_));
  OAI21_X1   g22749(.A1(new_n22941_), .A2(new_n22747_), .B(new_n22926_), .ZN(new_n22942_));
  NAND3_X1   g22750(.A1(new_n22942_), .A2(new_n1612_), .A3(new_n22748_), .ZN(new_n22943_));
  AOI22_X1   g22751(.A1(new_n22943_), .A2(new_n22762_), .B1(\asqrt[50] ), .B2(new_n22771_), .ZN(new_n22944_));
  OAI21_X1   g22752(.A1(new_n22944_), .A2(new_n1376_), .B(new_n1256_), .ZN(new_n22945_));
  OAI21_X1   g22753(.A1(new_n22945_), .A2(new_n22773_), .B(new_n22925_), .ZN(new_n22946_));
  NAND3_X1   g22754(.A1(new_n22946_), .A2(new_n1103_), .A3(new_n22774_), .ZN(new_n22947_));
  AOI22_X1   g22755(.A1(new_n22947_), .A2(new_n22789_), .B1(\asqrt[53] ), .B2(new_n22818_), .ZN(new_n22948_));
  OAI21_X1   g22756(.A1(new_n22948_), .A2(new_n904_), .B(new_n823_), .ZN(new_n22949_));
  OAI21_X1   g22757(.A1(new_n22949_), .A2(new_n22820_), .B(new_n22924_), .ZN(new_n22950_));
  NAND3_X1   g22758(.A1(new_n22950_), .A2(new_n703_), .A3(new_n22821_), .ZN(new_n22951_));
  AOI22_X1   g22759(.A1(new_n22951_), .A2(new_n22816_), .B1(\asqrt[56] ), .B2(new_n22850_), .ZN(new_n22952_));
  OAI21_X1   g22760(.A1(new_n22952_), .A2(new_n531_), .B(new_n436_), .ZN(new_n22953_));
  OAI21_X1   g22761(.A1(new_n22953_), .A2(new_n22852_), .B(new_n22923_), .ZN(new_n22954_));
  NAND3_X1   g22762(.A1(new_n22954_), .A2(new_n327_), .A3(new_n22853_), .ZN(new_n22955_));
  AOI22_X1   g22763(.A1(new_n22955_), .A2(new_n22848_), .B1(new_n22882_), .B2(\asqrt[59] ), .ZN(new_n22956_));
  OAI21_X1   g22764(.A1(new_n22956_), .A2(new_n306_), .B(new_n218_), .ZN(new_n22957_));
  OAI21_X1   g22765(.A1(new_n22957_), .A2(new_n22884_), .B(new_n22922_), .ZN(new_n22958_));
  NAND3_X1   g22766(.A1(new_n22958_), .A2(new_n207_), .A3(new_n22885_), .ZN(new_n22959_));
  AOI22_X1   g22767(.A1(new_n22959_), .A2(new_n22880_), .B1(new_n22921_), .B2(\asqrt[62] ), .ZN(new_n22960_));
  OAI21_X1   g22768(.A1(new_n22960_), .A2(new_n22896_), .B(new_n193_), .ZN(new_n22961_));
  AOI21_X1   g22769(.A1(new_n22921_), .A2(\asqrt[62] ), .B(new_n22892_), .ZN(new_n22962_));
  INV_X1     g22770(.I(new_n22904_), .ZN(new_n22963_));
  AOI21_X1   g22771(.A1(new_n22962_), .A2(new_n22887_), .B(new_n22963_), .ZN(new_n22964_));
  AOI21_X1   g22772(.A1(new_n22961_), .A2(new_n22964_), .B(new_n22291_), .ZN(new_n22965_));
  OAI21_X1   g22773(.A1(new_n22898_), .A2(new_n22905_), .B(new_n22912_), .ZN(new_n22966_));
  AOI21_X1   g22774(.A1(\a[7] ), .A2(new_n22966_), .B(new_n22965_), .ZN(new_n22967_));
  AOI22_X1   g22775(.A1(new_n22967_), .A2(new_n22919_), .B1(\asqrt[4] ), .B2(new_n22917_), .ZN(new_n22968_));
  NOR2_X1    g22776(.A1(new_n22968_), .A2(new_n21620_), .ZN(new_n22969_));
  NAND2_X1   g22777(.A1(new_n22967_), .A2(new_n22919_), .ZN(new_n22970_));
  OAI21_X1   g22778(.A1(new_n22898_), .A2(new_n22905_), .B(new_n22290_), .ZN(new_n22971_));
  NAND2_X1   g22779(.A1(new_n22962_), .A2(new_n22887_), .ZN(new_n22972_));
  NAND4_X1   g22780(.A1(new_n22961_), .A2(\asqrt[4] ), .A3(new_n22972_), .A4(new_n22904_), .ZN(new_n22973_));
  AOI21_X1   g22781(.A1(new_n22973_), .A2(new_n22971_), .B(new_n22303_), .ZN(new_n22974_));
  INV_X1     g22782(.I(new_n22972_), .ZN(new_n22975_));
  NAND2_X1   g22783(.A1(new_n22904_), .A2(\asqrt[4] ), .ZN(new_n22976_));
  NOR3_X1    g22784(.A1(new_n22975_), .A2(new_n22898_), .A3(new_n22976_), .ZN(new_n22977_));
  NOR3_X1    g22785(.A1(new_n22977_), .A2(new_n22965_), .A3(\a[8] ), .ZN(new_n22978_));
  NOR2_X1    g22786(.A1(new_n22974_), .A2(new_n22978_), .ZN(new_n22979_));
  AOI21_X1   g22787(.A1(new_n22917_), .A2(\asqrt[4] ), .B(\asqrt[5] ), .ZN(new_n22980_));
  AOI21_X1   g22788(.A1(new_n22970_), .A2(new_n22980_), .B(new_n22979_), .ZN(new_n22981_));
  OAI21_X1   g22789(.A1(new_n22981_), .A2(new_n22969_), .B(\asqrt[6] ), .ZN(new_n22982_));
  OAI21_X1   g22790(.A1(\asqrt[63] ), .A2(new_n22897_), .B(new_n22964_), .ZN(\asqrt[3] ));
  NOR3_X1    g22791(.A1(new_n22382_), .A2(new_n22302_), .A3(new_n22306_), .ZN(new_n22984_));
  NAND3_X1   g22792(.A1(\asqrt[3] ), .A2(new_n22319_), .A3(new_n22367_), .ZN(new_n22985_));
  AOI22_X1   g22793(.A1(new_n22985_), .A2(new_n22382_), .B1(\asqrt[3] ), .B2(new_n22984_), .ZN(new_n22986_));
  INV_X1     g22794(.I(new_n22986_), .ZN(new_n22987_));
  OAI21_X1   g22795(.A1(new_n22968_), .A2(new_n21620_), .B(new_n20806_), .ZN(new_n22988_));
  OAI21_X1   g22796(.A1(new_n22988_), .A2(new_n22981_), .B(new_n22987_), .ZN(new_n22989_));
  AOI21_X1   g22797(.A1(new_n22989_), .A2(new_n22982_), .B(new_n20262_), .ZN(new_n22990_));
  NOR2_X1    g22798(.A1(new_n22316_), .A2(new_n22318_), .ZN(new_n22991_));
  NOR2_X1    g22799(.A1(new_n22310_), .A2(new_n22320_), .ZN(new_n22992_));
  INV_X1     g22800(.I(new_n22992_), .ZN(new_n22993_));
  NAND4_X1   g22801(.A1(\asqrt[3] ), .A2(new_n22311_), .A3(new_n22991_), .A4(new_n22993_), .ZN(new_n22994_));
  NOR3_X1    g22802(.A1(new_n22906_), .A2(new_n22371_), .A3(new_n22992_), .ZN(new_n22995_));
  OAI21_X1   g22803(.A1(new_n22995_), .A2(new_n22991_), .B(new_n22994_), .ZN(new_n22996_));
  INV_X1     g22804(.I(new_n22996_), .ZN(new_n22997_));
  AOI21_X1   g22805(.A1(new_n22961_), .A2(new_n22964_), .B(new_n22912_), .ZN(new_n22998_));
  OAI21_X1   g22806(.A1(new_n22998_), .A2(new_n22915_), .B(\asqrt[4] ), .ZN(new_n22999_));
  INV_X1     g22807(.I(new_n22999_), .ZN(new_n23000_));
  INV_X1     g22808(.I(new_n22918_), .ZN(new_n23001_));
  NOR2_X1    g22809(.A1(new_n22998_), .A2(new_n23001_), .ZN(new_n23002_));
  INV_X1     g22810(.I(\a[7] ), .ZN(new_n23003_));
  AOI21_X1   g22811(.A1(\asqrt[3] ), .A2(new_n22912_), .B(new_n23003_), .ZN(new_n23004_));
  NOR3_X1    g22812(.A1(new_n23002_), .A2(new_n23004_), .A3(new_n22965_), .ZN(new_n23005_));
  OAI21_X1   g22813(.A1(new_n23005_), .A2(new_n23000_), .B(\asqrt[5] ), .ZN(new_n23006_));
  AOI21_X1   g22814(.A1(\asqrt[3] ), .A2(\a[6] ), .B(new_n22915_), .ZN(new_n23007_));
  OAI21_X1   g22815(.A1(new_n23007_), .A2(new_n22337_), .B(new_n21620_), .ZN(new_n23008_));
  OAI22_X1   g22816(.A1(new_n23005_), .A2(new_n23008_), .B1(new_n22974_), .B2(new_n22978_), .ZN(new_n23009_));
  AOI21_X1   g22817(.A1(new_n23009_), .A2(new_n23006_), .B(new_n20806_), .ZN(new_n23010_));
  AOI21_X1   g22818(.A1(new_n22961_), .A2(new_n22964_), .B(\a[6] ), .ZN(new_n23011_));
  OAI21_X1   g22819(.A1(new_n23003_), .A2(new_n23011_), .B(new_n22971_), .ZN(new_n23012_));
  OAI21_X1   g22820(.A1(new_n23012_), .A2(new_n23002_), .B(new_n22999_), .ZN(new_n23013_));
  AOI21_X1   g22821(.A1(new_n23013_), .A2(\asqrt[5] ), .B(\asqrt[6] ), .ZN(new_n23014_));
  AOI21_X1   g22822(.A1(new_n23014_), .A2(new_n23009_), .B(new_n22986_), .ZN(new_n23015_));
  NOR3_X1    g22823(.A1(new_n23015_), .A2(new_n23010_), .A3(\asqrt[7] ), .ZN(new_n23016_));
  NOR2_X1    g22824(.A1(new_n23016_), .A2(new_n22997_), .ZN(new_n23017_));
  OAI21_X1   g22825(.A1(new_n23017_), .A2(new_n22990_), .B(\asqrt[8] ), .ZN(new_n23018_));
  NOR2_X1    g22826(.A1(new_n22384_), .A2(new_n22376_), .ZN(new_n23019_));
  NOR3_X1    g22827(.A1(new_n22906_), .A2(new_n22322_), .A3(new_n23019_), .ZN(new_n23020_));
  INV_X1     g22828(.I(new_n23020_), .ZN(new_n23021_));
  NOR3_X1    g22829(.A1(new_n23019_), .A2(new_n22322_), .A3(new_n22381_), .ZN(new_n23022_));
  AOI22_X1   g22830(.A1(new_n23021_), .A2(new_n22381_), .B1(\asqrt[3] ), .B2(new_n23022_), .ZN(new_n23023_));
  INV_X1     g22831(.I(new_n23023_), .ZN(new_n23024_));
  OAI21_X1   g22832(.A1(new_n23015_), .A2(new_n23010_), .B(\asqrt[7] ), .ZN(new_n23025_));
  NAND2_X1   g22833(.A1(new_n23025_), .A2(new_n19573_), .ZN(new_n23026_));
  OAI21_X1   g22834(.A1(new_n23017_), .A2(new_n23026_), .B(new_n23024_), .ZN(new_n23027_));
  AOI21_X1   g22835(.A1(new_n23027_), .A2(new_n23018_), .B(new_n18792_), .ZN(new_n23028_));
  NOR3_X1    g22836(.A1(new_n22332_), .A2(new_n22341_), .A3(new_n22339_), .ZN(new_n23029_));
  NOR3_X1    g22837(.A1(new_n22906_), .A2(new_n22332_), .A3(new_n22341_), .ZN(new_n23030_));
  INV_X1     g22838(.I(new_n23030_), .ZN(new_n23031_));
  AOI22_X1   g22839(.A1(new_n23031_), .A2(new_n22339_), .B1(\asqrt[3] ), .B2(new_n23029_), .ZN(new_n23032_));
  OAI21_X1   g22840(.A1(new_n22997_), .A2(new_n23016_), .B(new_n23025_), .ZN(new_n23033_));
  AOI21_X1   g22841(.A1(new_n23033_), .A2(\asqrt[8] ), .B(\asqrt[9] ), .ZN(new_n23034_));
  AOI21_X1   g22842(.A1(new_n23034_), .A2(new_n23027_), .B(new_n23032_), .ZN(new_n23035_));
  OAI21_X1   g22843(.A1(new_n23035_), .A2(new_n23028_), .B(\asqrt[10] ), .ZN(new_n23036_));
  INV_X1     g22844(.I(new_n23036_), .ZN(new_n23037_));
  NAND2_X1   g22845(.A1(new_n22387_), .A2(new_n22379_), .ZN(new_n23038_));
  NAND3_X1   g22846(.A1(\asqrt[3] ), .A2(new_n22343_), .A3(new_n23038_), .ZN(new_n23039_));
  AND3_X2    g22847(.A1(new_n22343_), .A2(new_n22348_), .A3(new_n23038_), .Z(new_n23040_));
  AOI22_X1   g22848(.A1(new_n23039_), .A2(new_n22349_), .B1(\asqrt[3] ), .B2(new_n23040_), .ZN(new_n23041_));
  NOR3_X1    g22849(.A1(new_n23035_), .A2(new_n23028_), .A3(\asqrt[10] ), .ZN(new_n23042_));
  NOR2_X1    g22850(.A1(new_n23042_), .A2(new_n23041_), .ZN(new_n23043_));
  OAI21_X1   g22851(.A1(new_n23043_), .A2(new_n23037_), .B(\asqrt[11] ), .ZN(new_n23044_));
  INV_X1     g22852(.I(new_n22356_), .ZN(new_n23045_));
  NOR3_X1    g22853(.A1(new_n22352_), .A2(new_n22398_), .A3(new_n23045_), .ZN(new_n23046_));
  NOR3_X1    g22854(.A1(new_n22906_), .A2(new_n22352_), .A3(new_n22398_), .ZN(new_n23047_));
  INV_X1     g22855(.I(new_n23047_), .ZN(new_n23048_));
  AOI22_X1   g22856(.A1(new_n23048_), .A2(new_n23045_), .B1(\asqrt[3] ), .B2(new_n23046_), .ZN(new_n23049_));
  INV_X1     g22857(.I(new_n23049_), .ZN(new_n23050_));
  NAND2_X1   g22858(.A1(new_n23036_), .A2(new_n17623_), .ZN(new_n23051_));
  OAI21_X1   g22859(.A1(new_n23043_), .A2(new_n23051_), .B(new_n23050_), .ZN(new_n23052_));
  AOI21_X1   g22860(.A1(new_n23052_), .A2(new_n23044_), .B(new_n16881_), .ZN(new_n23053_));
  INV_X1     g22861(.I(new_n22425_), .ZN(new_n23054_));
  NAND3_X1   g22862(.A1(\asqrt[3] ), .A2(new_n22360_), .A3(new_n23054_), .ZN(new_n23055_));
  AND3_X2    g22863(.A1(new_n23054_), .A2(new_n22360_), .A3(new_n22364_), .Z(new_n23056_));
  AOI22_X1   g22864(.A1(new_n23055_), .A2(new_n22365_), .B1(\asqrt[3] ), .B2(new_n23056_), .ZN(new_n23057_));
  OAI21_X1   g22865(.A1(new_n23041_), .A2(new_n23042_), .B(new_n23036_), .ZN(new_n23058_));
  AOI21_X1   g22866(.A1(new_n23058_), .A2(\asqrt[11] ), .B(\asqrt[12] ), .ZN(new_n23059_));
  AOI21_X1   g22867(.A1(new_n23059_), .A2(new_n23052_), .B(new_n23057_), .ZN(new_n23060_));
  OAI21_X1   g22868(.A1(new_n23060_), .A2(new_n23053_), .B(\asqrt[13] ), .ZN(new_n23061_));
  INV_X1     g22869(.I(new_n23061_), .ZN(new_n23062_));
  INV_X1     g22870(.I(new_n22392_), .ZN(new_n23063_));
  AND3_X2    g22871(.A1(new_n23063_), .A2(new_n22397_), .A3(new_n22428_), .Z(new_n23064_));
  NAND3_X1   g22872(.A1(\asqrt[3] ), .A2(new_n23063_), .A3(new_n22428_), .ZN(new_n23065_));
  AOI22_X1   g22873(.A1(new_n23065_), .A2(new_n22427_), .B1(\asqrt[3] ), .B2(new_n23064_), .ZN(new_n23066_));
  NOR3_X1    g22874(.A1(new_n23060_), .A2(new_n23053_), .A3(\asqrt[13] ), .ZN(new_n23067_));
  NOR2_X1    g22875(.A1(new_n23067_), .A2(new_n23066_), .ZN(new_n23068_));
  OAI21_X1   g22876(.A1(new_n23068_), .A2(new_n23062_), .B(\asqrt[14] ), .ZN(new_n23069_));
  INV_X1     g22877(.I(new_n22407_), .ZN(new_n23070_));
  NOR3_X1    g22878(.A1(new_n22906_), .A2(new_n22403_), .A3(new_n22408_), .ZN(new_n23071_));
  INV_X1     g22879(.I(new_n23071_), .ZN(new_n23072_));
  NOR3_X1    g22880(.A1(new_n22403_), .A2(new_n23070_), .A3(new_n22408_), .ZN(new_n23073_));
  AOI22_X1   g22881(.A1(new_n23072_), .A2(new_n23070_), .B1(\asqrt[3] ), .B2(new_n23073_), .ZN(new_n23074_));
  INV_X1     g22882(.I(new_n23074_), .ZN(new_n23075_));
  NAND2_X1   g22883(.A1(new_n23061_), .A2(new_n15770_), .ZN(new_n23076_));
  OAI21_X1   g22884(.A1(new_n23068_), .A2(new_n23076_), .B(new_n23075_), .ZN(new_n23077_));
  AOI21_X1   g22885(.A1(new_n23077_), .A2(new_n23069_), .B(new_n15067_), .ZN(new_n23078_));
  OAI21_X1   g22886(.A1(new_n22409_), .A2(new_n22417_), .B(new_n22415_), .ZN(new_n23079_));
  AOI21_X1   g22887(.A1(\asqrt[14] ), .A2(new_n22430_), .B(new_n23079_), .ZN(new_n23080_));
  OAI21_X1   g22888(.A1(new_n22409_), .A2(new_n22417_), .B(new_n22410_), .ZN(new_n23081_));
  NOR2_X1    g22889(.A1(new_n22906_), .A2(new_n23081_), .ZN(new_n23082_));
  INV_X1     g22890(.I(new_n23082_), .ZN(new_n23083_));
  AOI22_X1   g22891(.A1(new_n23083_), .A2(new_n22416_), .B1(\asqrt[3] ), .B2(new_n23080_), .ZN(new_n23084_));
  OAI21_X1   g22892(.A1(new_n23066_), .A2(new_n23067_), .B(new_n23061_), .ZN(new_n23085_));
  AOI21_X1   g22893(.A1(new_n23085_), .A2(\asqrt[14] ), .B(\asqrt[15] ), .ZN(new_n23086_));
  AOI21_X1   g22894(.A1(new_n23086_), .A2(new_n23077_), .B(new_n23084_), .ZN(new_n23087_));
  OAI21_X1   g22895(.A1(new_n23087_), .A2(new_n23078_), .B(\asqrt[16] ), .ZN(new_n23088_));
  INV_X1     g22896(.I(new_n23088_), .ZN(new_n23089_));
  INV_X1     g22897(.I(new_n22424_), .ZN(new_n23090_));
  INV_X1     g22898(.I(new_n22418_), .ZN(new_n23091_));
  INV_X1     g22899(.I(new_n22431_), .ZN(new_n23092_));
  NOR2_X1    g22900(.A1(new_n23092_), .A2(new_n23091_), .ZN(new_n23093_));
  NOR3_X1    g22901(.A1(new_n22906_), .A2(new_n22419_), .A3(new_n23093_), .ZN(new_n23094_));
  INV_X1     g22902(.I(new_n23094_), .ZN(new_n23095_));
  NOR3_X1    g22903(.A1(new_n23093_), .A2(new_n22419_), .A3(new_n23090_), .ZN(new_n23096_));
  AOI22_X1   g22904(.A1(new_n23095_), .A2(new_n23090_), .B1(\asqrt[3] ), .B2(new_n23096_), .ZN(new_n23097_));
  NOR3_X1    g22905(.A1(new_n23087_), .A2(new_n23078_), .A3(\asqrt[16] ), .ZN(new_n23098_));
  NOR2_X1    g22906(.A1(new_n23098_), .A2(new_n23097_), .ZN(new_n23099_));
  OAI21_X1   g22907(.A1(new_n23099_), .A2(new_n23089_), .B(\asqrt[17] ), .ZN(new_n23100_));
  INV_X1     g22908(.I(new_n22438_), .ZN(new_n23101_));
  NOR3_X1    g22909(.A1(new_n22434_), .A2(new_n23101_), .A3(new_n22439_), .ZN(new_n23102_));
  NOR3_X1    g22910(.A1(new_n22906_), .A2(new_n22434_), .A3(new_n22439_), .ZN(new_n23103_));
  INV_X1     g22911(.I(new_n23103_), .ZN(new_n23104_));
  AOI22_X1   g22912(.A1(new_n23104_), .A2(new_n23101_), .B1(\asqrt[3] ), .B2(new_n23102_), .ZN(new_n23105_));
  INV_X1     g22913(.I(new_n23105_), .ZN(new_n23106_));
  NAND2_X1   g22914(.A1(new_n23088_), .A2(new_n14017_), .ZN(new_n23107_));
  OAI21_X1   g22915(.A1(new_n23099_), .A2(new_n23107_), .B(new_n23106_), .ZN(new_n23108_));
  AOI21_X1   g22916(.A1(new_n23108_), .A2(new_n23100_), .B(new_n13353_), .ZN(new_n23109_));
  NOR2_X1    g22917(.A1(new_n22440_), .A2(new_n22448_), .ZN(new_n23110_));
  INV_X1     g22918(.I(new_n23110_), .ZN(new_n23111_));
  NAND3_X1   g22919(.A1(\asqrt[3] ), .A2(new_n22441_), .A3(new_n23111_), .ZN(new_n23112_));
  AND3_X2    g22920(.A1(new_n23111_), .A2(new_n22441_), .A3(new_n22446_), .Z(new_n23113_));
  AOI22_X1   g22921(.A1(new_n23112_), .A2(new_n22447_), .B1(\asqrt[3] ), .B2(new_n23113_), .ZN(new_n23114_));
  OAI21_X1   g22922(.A1(new_n23097_), .A2(new_n23098_), .B(new_n23088_), .ZN(new_n23115_));
  AOI21_X1   g22923(.A1(new_n23115_), .A2(\asqrt[17] ), .B(\asqrt[18] ), .ZN(new_n23116_));
  AOI21_X1   g22924(.A1(new_n23116_), .A2(new_n23108_), .B(new_n23114_), .ZN(new_n23117_));
  OAI21_X1   g22925(.A1(new_n23117_), .A2(new_n23109_), .B(\asqrt[19] ), .ZN(new_n23118_));
  INV_X1     g22926(.I(new_n23118_), .ZN(new_n23119_));
  INV_X1     g22927(.I(new_n22455_), .ZN(new_n23120_));
  INV_X1     g22928(.I(new_n22449_), .ZN(new_n23121_));
  INV_X1     g22929(.I(new_n22457_), .ZN(new_n23122_));
  NOR2_X1    g22930(.A1(new_n23122_), .A2(new_n23121_), .ZN(new_n23123_));
  NOR3_X1    g22931(.A1(new_n23123_), .A2(new_n22450_), .A3(new_n23120_), .ZN(new_n23124_));
  NOR3_X1    g22932(.A1(new_n22906_), .A2(new_n22450_), .A3(new_n23123_), .ZN(new_n23125_));
  INV_X1     g22933(.I(new_n23125_), .ZN(new_n23126_));
  AOI22_X1   g22934(.A1(new_n23126_), .A2(new_n23120_), .B1(\asqrt[3] ), .B2(new_n23124_), .ZN(new_n23127_));
  NOR3_X1    g22935(.A1(new_n23117_), .A2(new_n23109_), .A3(\asqrt[19] ), .ZN(new_n23128_));
  NOR2_X1    g22936(.A1(new_n23128_), .A2(new_n23127_), .ZN(new_n23129_));
  OAI21_X1   g22937(.A1(new_n23129_), .A2(new_n23119_), .B(\asqrt[20] ), .ZN(new_n23130_));
  INV_X1     g22938(.I(new_n22464_), .ZN(new_n23131_));
  NOR3_X1    g22939(.A1(new_n22906_), .A2(new_n22460_), .A3(new_n22465_), .ZN(new_n23132_));
  INV_X1     g22940(.I(new_n23132_), .ZN(new_n23133_));
  NOR3_X1    g22941(.A1(new_n22460_), .A2(new_n23131_), .A3(new_n22465_), .ZN(new_n23134_));
  AOI22_X1   g22942(.A1(new_n23133_), .A2(new_n23131_), .B1(\asqrt[3] ), .B2(new_n23134_), .ZN(new_n23135_));
  INV_X1     g22943(.I(new_n23135_), .ZN(new_n23136_));
  NAND2_X1   g22944(.A1(new_n23118_), .A2(new_n12364_), .ZN(new_n23137_));
  OAI21_X1   g22945(.A1(new_n23129_), .A2(new_n23137_), .B(new_n23136_), .ZN(new_n23138_));
  AOI21_X1   g22946(.A1(new_n23138_), .A2(new_n23130_), .B(new_n11736_), .ZN(new_n23139_));
  NOR2_X1    g22947(.A1(new_n22466_), .A2(new_n22474_), .ZN(new_n23140_));
  INV_X1     g22948(.I(new_n23140_), .ZN(new_n23141_));
  AND3_X2    g22949(.A1(new_n23141_), .A2(new_n22467_), .A3(new_n22472_), .Z(new_n23142_));
  NAND3_X1   g22950(.A1(\asqrt[3] ), .A2(new_n22467_), .A3(new_n23141_), .ZN(new_n23143_));
  AOI22_X1   g22951(.A1(new_n23143_), .A2(new_n22473_), .B1(\asqrt[3] ), .B2(new_n23142_), .ZN(new_n23144_));
  OAI21_X1   g22952(.A1(new_n23127_), .A2(new_n23128_), .B(new_n23118_), .ZN(new_n23145_));
  AOI21_X1   g22953(.A1(new_n23145_), .A2(\asqrt[20] ), .B(\asqrt[21] ), .ZN(new_n23146_));
  AOI21_X1   g22954(.A1(new_n23146_), .A2(new_n23138_), .B(new_n23144_), .ZN(new_n23147_));
  OAI21_X1   g22955(.A1(new_n23147_), .A2(new_n23139_), .B(\asqrt[22] ), .ZN(new_n23148_));
  INV_X1     g22956(.I(new_n23148_), .ZN(new_n23149_));
  INV_X1     g22957(.I(new_n22481_), .ZN(new_n23150_));
  INV_X1     g22958(.I(new_n22475_), .ZN(new_n23151_));
  INV_X1     g22959(.I(new_n22483_), .ZN(new_n23152_));
  NOR2_X1    g22960(.A1(new_n23152_), .A2(new_n23151_), .ZN(new_n23153_));
  NOR3_X1    g22961(.A1(new_n22906_), .A2(new_n22476_), .A3(new_n23153_), .ZN(new_n23154_));
  INV_X1     g22962(.I(new_n23154_), .ZN(new_n23155_));
  NOR3_X1    g22963(.A1(new_n23153_), .A2(new_n22476_), .A3(new_n23150_), .ZN(new_n23156_));
  AOI22_X1   g22964(.A1(new_n23155_), .A2(new_n23150_), .B1(\asqrt[3] ), .B2(new_n23156_), .ZN(new_n23157_));
  NOR3_X1    g22965(.A1(new_n23147_), .A2(new_n23139_), .A3(\asqrt[22] ), .ZN(new_n23158_));
  NOR2_X1    g22966(.A1(new_n23158_), .A2(new_n23157_), .ZN(new_n23159_));
  OAI21_X1   g22967(.A1(new_n23159_), .A2(new_n23149_), .B(\asqrt[23] ), .ZN(new_n23160_));
  INV_X1     g22968(.I(new_n22490_), .ZN(new_n23161_));
  NOR3_X1    g22969(.A1(new_n22486_), .A2(new_n23161_), .A3(new_n22491_), .ZN(new_n23162_));
  NOR3_X1    g22970(.A1(new_n22906_), .A2(new_n22486_), .A3(new_n22491_), .ZN(new_n23163_));
  INV_X1     g22971(.I(new_n23163_), .ZN(new_n23164_));
  AOI22_X1   g22972(.A1(new_n23164_), .A2(new_n23161_), .B1(\asqrt[3] ), .B2(new_n23162_), .ZN(new_n23165_));
  INV_X1     g22973(.I(new_n23165_), .ZN(new_n23166_));
  NAND2_X1   g22974(.A1(new_n23148_), .A2(new_n10812_), .ZN(new_n23167_));
  OAI21_X1   g22975(.A1(new_n23159_), .A2(new_n23167_), .B(new_n23166_), .ZN(new_n23168_));
  AOI21_X1   g22976(.A1(new_n23168_), .A2(new_n23160_), .B(new_n10221_), .ZN(new_n23169_));
  NOR2_X1    g22977(.A1(new_n22492_), .A2(new_n22500_), .ZN(new_n23170_));
  INV_X1     g22978(.I(new_n23170_), .ZN(new_n23171_));
  NAND3_X1   g22979(.A1(\asqrt[3] ), .A2(new_n22493_), .A3(new_n23171_), .ZN(new_n23172_));
  AND3_X2    g22980(.A1(new_n23171_), .A2(new_n22493_), .A3(new_n22498_), .Z(new_n23173_));
  AOI22_X1   g22981(.A1(new_n23172_), .A2(new_n22499_), .B1(\asqrt[3] ), .B2(new_n23173_), .ZN(new_n23174_));
  OAI21_X1   g22982(.A1(new_n23157_), .A2(new_n23158_), .B(new_n23148_), .ZN(new_n23175_));
  AOI21_X1   g22983(.A1(new_n23175_), .A2(\asqrt[23] ), .B(\asqrt[24] ), .ZN(new_n23176_));
  AOI21_X1   g22984(.A1(new_n23176_), .A2(new_n23168_), .B(new_n23174_), .ZN(new_n23177_));
  OAI21_X1   g22985(.A1(new_n23177_), .A2(new_n23169_), .B(\asqrt[25] ), .ZN(new_n23178_));
  INV_X1     g22986(.I(new_n23178_), .ZN(new_n23179_));
  INV_X1     g22987(.I(new_n22507_), .ZN(new_n23180_));
  INV_X1     g22988(.I(new_n22501_), .ZN(new_n23181_));
  INV_X1     g22989(.I(new_n22509_), .ZN(new_n23182_));
  NOR2_X1    g22990(.A1(new_n23182_), .A2(new_n23181_), .ZN(new_n23183_));
  NOR3_X1    g22991(.A1(new_n23183_), .A2(new_n22502_), .A3(new_n23180_), .ZN(new_n23184_));
  NOR3_X1    g22992(.A1(new_n22906_), .A2(new_n22502_), .A3(new_n23183_), .ZN(new_n23185_));
  INV_X1     g22993(.I(new_n23185_), .ZN(new_n23186_));
  AOI22_X1   g22994(.A1(new_n23186_), .A2(new_n23180_), .B1(\asqrt[3] ), .B2(new_n23184_), .ZN(new_n23187_));
  NOR3_X1    g22995(.A1(new_n23177_), .A2(new_n23169_), .A3(\asqrt[25] ), .ZN(new_n23188_));
  NOR2_X1    g22996(.A1(new_n23188_), .A2(new_n23187_), .ZN(new_n23189_));
  OAI21_X1   g22997(.A1(new_n23189_), .A2(new_n23179_), .B(\asqrt[26] ), .ZN(new_n23190_));
  INV_X1     g22998(.I(new_n22516_), .ZN(new_n23191_));
  NOR3_X1    g22999(.A1(new_n22906_), .A2(new_n22512_), .A3(new_n22517_), .ZN(new_n23192_));
  INV_X1     g23000(.I(new_n23192_), .ZN(new_n23193_));
  NOR3_X1    g23001(.A1(new_n22512_), .A2(new_n23191_), .A3(new_n22517_), .ZN(new_n23194_));
  AOI22_X1   g23002(.A1(new_n23193_), .A2(new_n23191_), .B1(\asqrt[3] ), .B2(new_n23194_), .ZN(new_n23195_));
  INV_X1     g23003(.I(new_n23195_), .ZN(new_n23196_));
  NAND2_X1   g23004(.A1(new_n23178_), .A2(new_n9317_), .ZN(new_n23197_));
  OAI21_X1   g23005(.A1(new_n23189_), .A2(new_n23197_), .B(new_n23196_), .ZN(new_n23198_));
  AOI21_X1   g23006(.A1(new_n23198_), .A2(new_n23190_), .B(new_n8826_), .ZN(new_n23199_));
  NOR2_X1    g23007(.A1(new_n22518_), .A2(new_n22526_), .ZN(new_n23200_));
  INV_X1     g23008(.I(new_n23200_), .ZN(new_n23201_));
  AND3_X2    g23009(.A1(new_n23201_), .A2(new_n22519_), .A3(new_n22524_), .Z(new_n23202_));
  NAND3_X1   g23010(.A1(\asqrt[3] ), .A2(new_n22519_), .A3(new_n23201_), .ZN(new_n23203_));
  AOI22_X1   g23011(.A1(new_n23203_), .A2(new_n22525_), .B1(\asqrt[3] ), .B2(new_n23202_), .ZN(new_n23204_));
  OAI21_X1   g23012(.A1(new_n23187_), .A2(new_n23188_), .B(new_n23178_), .ZN(new_n23205_));
  AOI21_X1   g23013(.A1(new_n23205_), .A2(\asqrt[26] ), .B(\asqrt[27] ), .ZN(new_n23206_));
  AOI21_X1   g23014(.A1(new_n23206_), .A2(new_n23198_), .B(new_n23204_), .ZN(new_n23207_));
  OAI21_X1   g23015(.A1(new_n23207_), .A2(new_n23199_), .B(\asqrt[28] ), .ZN(new_n23208_));
  INV_X1     g23016(.I(new_n23208_), .ZN(new_n23209_));
  INV_X1     g23017(.I(new_n22533_), .ZN(new_n23210_));
  INV_X1     g23018(.I(new_n22527_), .ZN(new_n23211_));
  INV_X1     g23019(.I(new_n22535_), .ZN(new_n23212_));
  NOR2_X1    g23020(.A1(new_n23212_), .A2(new_n23211_), .ZN(new_n23213_));
  NOR3_X1    g23021(.A1(new_n22906_), .A2(new_n22528_), .A3(new_n23213_), .ZN(new_n23214_));
  INV_X1     g23022(.I(new_n23214_), .ZN(new_n23215_));
  NOR3_X1    g23023(.A1(new_n23213_), .A2(new_n22528_), .A3(new_n23210_), .ZN(new_n23216_));
  AOI22_X1   g23024(.A1(new_n23215_), .A2(new_n23210_), .B1(\asqrt[3] ), .B2(new_n23216_), .ZN(new_n23217_));
  NOR3_X1    g23025(.A1(new_n23207_), .A2(new_n23199_), .A3(\asqrt[28] ), .ZN(new_n23218_));
  NOR2_X1    g23026(.A1(new_n23218_), .A2(new_n23217_), .ZN(new_n23219_));
  OAI21_X1   g23027(.A1(new_n23219_), .A2(new_n23209_), .B(\asqrt[29] ), .ZN(new_n23220_));
  INV_X1     g23028(.I(new_n22543_), .ZN(new_n23221_));
  NOR3_X1    g23029(.A1(new_n22538_), .A2(new_n23221_), .A3(new_n22580_), .ZN(new_n23222_));
  NOR3_X1    g23030(.A1(new_n22906_), .A2(new_n22538_), .A3(new_n22580_), .ZN(new_n23223_));
  INV_X1     g23031(.I(new_n23223_), .ZN(new_n23224_));
  AOI22_X1   g23032(.A1(new_n23224_), .A2(new_n23221_), .B1(\asqrt[3] ), .B2(new_n23222_), .ZN(new_n23225_));
  INV_X1     g23033(.I(new_n23225_), .ZN(new_n23226_));
  NAND2_X1   g23034(.A1(new_n23208_), .A2(new_n8036_), .ZN(new_n23227_));
  OAI21_X1   g23035(.A1(new_n23219_), .A2(new_n23227_), .B(new_n23226_), .ZN(new_n23228_));
  AOI21_X1   g23036(.A1(new_n23228_), .A2(new_n23220_), .B(new_n7539_), .ZN(new_n23229_));
  NOR2_X1    g23037(.A1(new_n22553_), .A2(new_n22545_), .ZN(new_n23230_));
  INV_X1     g23038(.I(new_n23230_), .ZN(new_n23231_));
  NAND3_X1   g23039(.A1(\asqrt[3] ), .A2(new_n22546_), .A3(new_n23231_), .ZN(new_n23232_));
  AND3_X2    g23040(.A1(new_n23231_), .A2(new_n22546_), .A3(new_n22551_), .Z(new_n23233_));
  AOI22_X1   g23041(.A1(new_n23232_), .A2(new_n22552_), .B1(\asqrt[3] ), .B2(new_n23233_), .ZN(new_n23234_));
  OAI21_X1   g23042(.A1(new_n23217_), .A2(new_n23218_), .B(new_n23208_), .ZN(new_n23235_));
  AOI21_X1   g23043(.A1(new_n23235_), .A2(\asqrt[29] ), .B(\asqrt[30] ), .ZN(new_n23236_));
  AOI21_X1   g23044(.A1(new_n23236_), .A2(new_n23228_), .B(new_n23234_), .ZN(new_n23237_));
  OAI21_X1   g23045(.A1(new_n23237_), .A2(new_n23229_), .B(\asqrt[31] ), .ZN(new_n23238_));
  INV_X1     g23046(.I(new_n23238_), .ZN(new_n23239_));
  NOR2_X1    g23047(.A1(new_n22564_), .A2(new_n22557_), .ZN(new_n23240_));
  NOR3_X1    g23048(.A1(new_n23240_), .A2(new_n22555_), .A3(new_n22563_), .ZN(new_n23241_));
  NOR3_X1    g23049(.A1(new_n22906_), .A2(new_n22555_), .A3(new_n23240_), .ZN(new_n23242_));
  INV_X1     g23050(.I(new_n23242_), .ZN(new_n23243_));
  AOI22_X1   g23051(.A1(new_n23243_), .A2(new_n22563_), .B1(\asqrt[3] ), .B2(new_n23241_), .ZN(new_n23244_));
  NOR3_X1    g23052(.A1(new_n23237_), .A2(new_n23229_), .A3(\asqrt[31] ), .ZN(new_n23245_));
  NOR2_X1    g23053(.A1(new_n23245_), .A2(new_n23244_), .ZN(new_n23246_));
  OAI21_X1   g23054(.A1(new_n23246_), .A2(new_n23239_), .B(\asqrt[32] ), .ZN(new_n23247_));
  INV_X1     g23055(.I(new_n22570_), .ZN(new_n23248_));
  NOR3_X1    g23056(.A1(new_n22906_), .A2(new_n22566_), .A3(new_n22612_), .ZN(new_n23249_));
  INV_X1     g23057(.I(new_n23249_), .ZN(new_n23250_));
  NOR3_X1    g23058(.A1(new_n22566_), .A2(new_n23248_), .A3(new_n22612_), .ZN(new_n23251_));
  AOI22_X1   g23059(.A1(new_n23250_), .A2(new_n23248_), .B1(\asqrt[3] ), .B2(new_n23251_), .ZN(new_n23252_));
  INV_X1     g23060(.I(new_n23252_), .ZN(new_n23253_));
  NAND2_X1   g23061(.A1(new_n23238_), .A2(new_n6824_), .ZN(new_n23254_));
  OAI21_X1   g23062(.A1(new_n23246_), .A2(new_n23254_), .B(new_n23253_), .ZN(new_n23255_));
  AOI21_X1   g23063(.A1(new_n23255_), .A2(new_n23247_), .B(new_n6356_), .ZN(new_n23256_));
  NOR2_X1    g23064(.A1(new_n22585_), .A2(new_n22572_), .ZN(new_n23257_));
  INV_X1     g23065(.I(new_n23257_), .ZN(new_n23258_));
  AND3_X2    g23066(.A1(new_n23258_), .A2(new_n22573_), .A3(new_n22578_), .Z(new_n23259_));
  NAND3_X1   g23067(.A1(\asqrt[3] ), .A2(new_n22573_), .A3(new_n23258_), .ZN(new_n23260_));
  AOI22_X1   g23068(.A1(new_n23260_), .A2(new_n22579_), .B1(\asqrt[3] ), .B2(new_n23259_), .ZN(new_n23261_));
  OAI21_X1   g23069(.A1(new_n23244_), .A2(new_n23245_), .B(new_n23238_), .ZN(new_n23262_));
  AOI21_X1   g23070(.A1(new_n23262_), .A2(\asqrt[32] ), .B(\asqrt[33] ), .ZN(new_n23263_));
  AOI21_X1   g23071(.A1(new_n23263_), .A2(new_n23255_), .B(new_n23261_), .ZN(new_n23264_));
  OAI21_X1   g23072(.A1(new_n23264_), .A2(new_n23256_), .B(\asqrt[34] ), .ZN(new_n23265_));
  INV_X1     g23073(.I(new_n23265_), .ZN(new_n23266_));
  NOR2_X1    g23074(.A1(new_n22596_), .A2(new_n22589_), .ZN(new_n23267_));
  NOR3_X1    g23075(.A1(new_n22906_), .A2(new_n22587_), .A3(new_n23267_), .ZN(new_n23268_));
  INV_X1     g23076(.I(new_n23268_), .ZN(new_n23269_));
  NOR3_X1    g23077(.A1(new_n23267_), .A2(new_n22587_), .A3(new_n22595_), .ZN(new_n23270_));
  AOI22_X1   g23078(.A1(new_n23269_), .A2(new_n22595_), .B1(\asqrt[3] ), .B2(new_n23270_), .ZN(new_n23271_));
  NOR3_X1    g23079(.A1(new_n23264_), .A2(new_n23256_), .A3(\asqrt[34] ), .ZN(new_n23272_));
  NOR2_X1    g23080(.A1(new_n23272_), .A2(new_n23271_), .ZN(new_n23273_));
  OAI21_X1   g23081(.A1(new_n23273_), .A2(new_n23266_), .B(\asqrt[35] ), .ZN(new_n23274_));
  INV_X1     g23082(.I(new_n22602_), .ZN(new_n23275_));
  NOR3_X1    g23083(.A1(new_n22598_), .A2(new_n23275_), .A3(new_n22662_), .ZN(new_n23276_));
  NOR3_X1    g23084(.A1(new_n22906_), .A2(new_n22598_), .A3(new_n22662_), .ZN(new_n23277_));
  INV_X1     g23085(.I(new_n23277_), .ZN(new_n23278_));
  AOI22_X1   g23086(.A1(new_n23278_), .A2(new_n23275_), .B1(\asqrt[3] ), .B2(new_n23276_), .ZN(new_n23279_));
  INV_X1     g23087(.I(new_n23279_), .ZN(new_n23280_));
  NAND2_X1   g23088(.A1(new_n23265_), .A2(new_n5708_), .ZN(new_n23281_));
  OAI21_X1   g23089(.A1(new_n23273_), .A2(new_n23281_), .B(new_n23280_), .ZN(new_n23282_));
  AOI21_X1   g23090(.A1(new_n23282_), .A2(new_n23274_), .B(new_n5277_), .ZN(new_n23283_));
  NOR2_X1    g23091(.A1(new_n22617_), .A2(new_n22604_), .ZN(new_n23284_));
  INV_X1     g23092(.I(new_n23284_), .ZN(new_n23285_));
  NAND3_X1   g23093(.A1(\asqrt[3] ), .A2(new_n22605_), .A3(new_n23285_), .ZN(new_n23286_));
  AND3_X2    g23094(.A1(new_n23285_), .A2(new_n22605_), .A3(new_n22610_), .Z(new_n23287_));
  AOI22_X1   g23095(.A1(new_n23286_), .A2(new_n22611_), .B1(\asqrt[3] ), .B2(new_n23287_), .ZN(new_n23288_));
  OAI21_X1   g23096(.A1(new_n23271_), .A2(new_n23272_), .B(new_n23265_), .ZN(new_n23289_));
  AOI21_X1   g23097(.A1(new_n23289_), .A2(\asqrt[35] ), .B(\asqrt[36] ), .ZN(new_n23290_));
  AOI21_X1   g23098(.A1(new_n23290_), .A2(new_n23282_), .B(new_n23288_), .ZN(new_n23291_));
  OAI21_X1   g23099(.A1(new_n23291_), .A2(new_n23283_), .B(\asqrt[37] ), .ZN(new_n23292_));
  INV_X1     g23100(.I(new_n23292_), .ZN(new_n23293_));
  NOR2_X1    g23101(.A1(new_n22621_), .A2(new_n22628_), .ZN(new_n23294_));
  NOR3_X1    g23102(.A1(new_n23294_), .A2(new_n22635_), .A3(new_n22627_), .ZN(new_n23295_));
  NOR3_X1    g23103(.A1(new_n22906_), .A2(new_n22635_), .A3(new_n23294_), .ZN(new_n23296_));
  INV_X1     g23104(.I(new_n23296_), .ZN(new_n23297_));
  AOI22_X1   g23105(.A1(new_n23297_), .A2(new_n22627_), .B1(\asqrt[3] ), .B2(new_n23295_), .ZN(new_n23298_));
  NOR3_X1    g23106(.A1(new_n23291_), .A2(new_n23283_), .A3(\asqrt[37] ), .ZN(new_n23299_));
  NOR2_X1    g23107(.A1(new_n23299_), .A2(new_n23298_), .ZN(new_n23300_));
  OAI21_X1   g23108(.A1(new_n23300_), .A2(new_n23293_), .B(\asqrt[38] ), .ZN(new_n23301_));
  INV_X1     g23109(.I(new_n22634_), .ZN(new_n23302_));
  NOR3_X1    g23110(.A1(new_n22906_), .A2(new_n22630_), .A3(new_n22679_), .ZN(new_n23303_));
  INV_X1     g23111(.I(new_n23303_), .ZN(new_n23304_));
  NOR3_X1    g23112(.A1(new_n22630_), .A2(new_n23302_), .A3(new_n22679_), .ZN(new_n23305_));
  AOI22_X1   g23113(.A1(new_n23304_), .A2(new_n23302_), .B1(\asqrt[3] ), .B2(new_n23305_), .ZN(new_n23306_));
  INV_X1     g23114(.I(new_n23306_), .ZN(new_n23307_));
  NAND2_X1   g23115(.A1(new_n23292_), .A2(new_n4696_), .ZN(new_n23308_));
  OAI21_X1   g23116(.A1(new_n23300_), .A2(new_n23308_), .B(new_n23307_), .ZN(new_n23309_));
  AOI21_X1   g23117(.A1(new_n23309_), .A2(new_n23301_), .B(new_n4298_), .ZN(new_n23310_));
  NOR3_X1    g23118(.A1(new_n22639_), .A2(new_n22661_), .A3(new_n22645_), .ZN(new_n23311_));
  NOR3_X1    g23119(.A1(new_n22906_), .A2(new_n22639_), .A3(new_n22645_), .ZN(new_n23312_));
  INV_X1     g23120(.I(new_n23312_), .ZN(new_n23313_));
  AOI22_X1   g23121(.A1(new_n23313_), .A2(new_n22661_), .B1(\asqrt[3] ), .B2(new_n23311_), .ZN(new_n23314_));
  OAI21_X1   g23122(.A1(new_n23298_), .A2(new_n23299_), .B(new_n23292_), .ZN(new_n23315_));
  AOI21_X1   g23123(.A1(new_n23315_), .A2(\asqrt[38] ), .B(\asqrt[39] ), .ZN(new_n23316_));
  AOI21_X1   g23124(.A1(new_n23316_), .A2(new_n23309_), .B(new_n23314_), .ZN(new_n23317_));
  OAI21_X1   g23125(.A1(new_n23317_), .A2(new_n23310_), .B(\asqrt[40] ), .ZN(new_n23318_));
  INV_X1     g23126(.I(new_n23318_), .ZN(new_n23319_));
  NOR2_X1    g23127(.A1(new_n22646_), .A2(new_n22654_), .ZN(new_n23320_));
  NOR3_X1    g23128(.A1(new_n22906_), .A2(new_n22669_), .A3(new_n23320_), .ZN(new_n23321_));
  INV_X1     g23129(.I(new_n23321_), .ZN(new_n23322_));
  NOR3_X1    g23130(.A1(new_n23320_), .A2(new_n22669_), .A3(new_n22653_), .ZN(new_n23323_));
  AOI22_X1   g23131(.A1(new_n23322_), .A2(new_n22653_), .B1(\asqrt[3] ), .B2(new_n23323_), .ZN(new_n23324_));
  NOR3_X1    g23132(.A1(new_n23317_), .A2(new_n23310_), .A3(\asqrt[40] ), .ZN(new_n23325_));
  NOR2_X1    g23133(.A1(new_n23325_), .A2(new_n23324_), .ZN(new_n23326_));
  OAI21_X1   g23134(.A1(new_n23326_), .A2(new_n23319_), .B(\asqrt[41] ), .ZN(new_n23327_));
  INV_X1     g23135(.I(new_n22660_), .ZN(new_n23328_));
  NOR3_X1    g23136(.A1(new_n22656_), .A2(new_n23328_), .A3(new_n22692_), .ZN(new_n23329_));
  NOR3_X1    g23137(.A1(new_n22906_), .A2(new_n22656_), .A3(new_n22692_), .ZN(new_n23330_));
  INV_X1     g23138(.I(new_n23330_), .ZN(new_n23331_));
  AOI22_X1   g23139(.A1(new_n23331_), .A2(new_n23328_), .B1(\asqrt[3] ), .B2(new_n23329_), .ZN(new_n23332_));
  INV_X1     g23140(.I(new_n23332_), .ZN(new_n23333_));
  NAND2_X1   g23141(.A1(new_n23318_), .A2(new_n3782_), .ZN(new_n23334_));
  OAI21_X1   g23142(.A1(new_n23326_), .A2(new_n23334_), .B(new_n23333_), .ZN(new_n23335_));
  AOI21_X1   g23143(.A1(new_n23335_), .A2(new_n23327_), .B(new_n3419_), .ZN(new_n23336_));
  NOR3_X1    g23144(.A1(new_n22906_), .A2(new_n22929_), .A3(new_n22930_), .ZN(new_n23337_));
  INV_X1     g23145(.I(new_n23337_), .ZN(new_n23338_));
  NOR3_X1    g23146(.A1(new_n22929_), .A2(new_n22678_), .A3(new_n22930_), .ZN(new_n23339_));
  AOI22_X1   g23147(.A1(new_n23338_), .A2(new_n22678_), .B1(\asqrt[3] ), .B2(new_n23339_), .ZN(new_n23340_));
  OAI21_X1   g23148(.A1(new_n23324_), .A2(new_n23325_), .B(new_n23318_), .ZN(new_n23341_));
  AOI21_X1   g23149(.A1(new_n23341_), .A2(\asqrt[41] ), .B(\asqrt[42] ), .ZN(new_n23342_));
  AOI21_X1   g23150(.A1(new_n23342_), .A2(new_n23335_), .B(new_n23340_), .ZN(new_n23343_));
  OAI21_X1   g23151(.A1(new_n23343_), .A2(new_n23336_), .B(\asqrt[43] ), .ZN(new_n23344_));
  INV_X1     g23152(.I(new_n23344_), .ZN(new_n23345_));
  INV_X1     g23153(.I(new_n22691_), .ZN(new_n23346_));
  NAND2_X1   g23154(.A1(new_n22672_), .A2(new_n3419_), .ZN(new_n23347_));
  NOR2_X1    g23155(.A1(new_n22931_), .A2(new_n23347_), .ZN(new_n23348_));
  NOR3_X1    g23156(.A1(new_n23348_), .A2(new_n22686_), .A3(new_n23346_), .ZN(new_n23349_));
  NOR3_X1    g23157(.A1(new_n22906_), .A2(new_n22686_), .A3(new_n23348_), .ZN(new_n23350_));
  INV_X1     g23158(.I(new_n23350_), .ZN(new_n23351_));
  AOI22_X1   g23159(.A1(new_n23351_), .A2(new_n23346_), .B1(\asqrt[3] ), .B2(new_n23349_), .ZN(new_n23352_));
  NOR3_X1    g23160(.A1(new_n23343_), .A2(new_n23336_), .A3(\asqrt[43] ), .ZN(new_n23353_));
  NOR2_X1    g23161(.A1(new_n23353_), .A2(new_n23352_), .ZN(new_n23354_));
  OAI21_X1   g23162(.A1(new_n23354_), .A2(new_n23345_), .B(\asqrt[44] ), .ZN(new_n23355_));
  NOR3_X1    g23163(.A1(new_n22906_), .A2(new_n22697_), .A3(new_n22702_), .ZN(new_n23356_));
  INV_X1     g23164(.I(new_n23356_), .ZN(new_n23357_));
  NOR3_X1    g23165(.A1(new_n22697_), .A2(new_n22702_), .A3(new_n22928_), .ZN(new_n23358_));
  AOI22_X1   g23166(.A1(new_n23357_), .A2(new_n22928_), .B1(\asqrt[3] ), .B2(new_n23358_), .ZN(new_n23359_));
  INV_X1     g23167(.I(new_n23359_), .ZN(new_n23360_));
  NAND2_X1   g23168(.A1(new_n23344_), .A2(new_n2954_), .ZN(new_n23361_));
  OAI21_X1   g23169(.A1(new_n23354_), .A2(new_n23361_), .B(new_n23360_), .ZN(new_n23362_));
  AOI21_X1   g23170(.A1(new_n23362_), .A2(new_n23355_), .B(new_n2641_), .ZN(new_n23363_));
  INV_X1     g23171(.I(new_n22704_), .ZN(new_n23364_));
  NOR2_X1    g23172(.A1(new_n22703_), .A2(new_n22711_), .ZN(new_n23365_));
  NOR3_X1    g23173(.A1(new_n23364_), .A2(new_n23365_), .A3(new_n22710_), .ZN(new_n23366_));
  NOR3_X1    g23174(.A1(new_n22906_), .A2(new_n23364_), .A3(new_n23365_), .ZN(new_n23367_));
  INV_X1     g23175(.I(new_n23367_), .ZN(new_n23368_));
  AOI22_X1   g23176(.A1(new_n23368_), .A2(new_n22710_), .B1(\asqrt[3] ), .B2(new_n23366_), .ZN(new_n23369_));
  OAI21_X1   g23177(.A1(new_n23352_), .A2(new_n23353_), .B(new_n23344_), .ZN(new_n23370_));
  AOI21_X1   g23178(.A1(new_n23370_), .A2(\asqrt[44] ), .B(\asqrt[45] ), .ZN(new_n23371_));
  AOI21_X1   g23179(.A1(new_n23371_), .A2(new_n23362_), .B(new_n23369_), .ZN(new_n23372_));
  OAI21_X1   g23180(.A1(new_n23372_), .A2(new_n23363_), .B(\asqrt[46] ), .ZN(new_n23373_));
  INV_X1     g23181(.I(new_n23373_), .ZN(new_n23374_));
  INV_X1     g23182(.I(new_n22718_), .ZN(new_n23375_));
  INV_X1     g23183(.I(new_n22712_), .ZN(new_n23376_));
  INV_X1     g23184(.I(new_n22720_), .ZN(new_n23377_));
  NOR2_X1    g23185(.A1(new_n23377_), .A2(new_n23376_), .ZN(new_n23378_));
  NOR3_X1    g23186(.A1(new_n22906_), .A2(new_n22713_), .A3(new_n23378_), .ZN(new_n23379_));
  INV_X1     g23187(.I(new_n23379_), .ZN(new_n23380_));
  NOR3_X1    g23188(.A1(new_n23378_), .A2(new_n22713_), .A3(new_n23375_), .ZN(new_n23381_));
  AOI22_X1   g23189(.A1(new_n23380_), .A2(new_n23375_), .B1(\asqrt[3] ), .B2(new_n23381_), .ZN(new_n23382_));
  NOR3_X1    g23190(.A1(new_n23372_), .A2(new_n23363_), .A3(\asqrt[46] ), .ZN(new_n23383_));
  NOR2_X1    g23191(.A1(new_n23383_), .A2(new_n23382_), .ZN(new_n23384_));
  OAI21_X1   g23192(.A1(new_n23384_), .A2(new_n23374_), .B(\asqrt[47] ), .ZN(new_n23385_));
  NOR3_X1    g23193(.A1(new_n22723_), .A2(new_n22927_), .A3(new_n22728_), .ZN(new_n23386_));
  NOR3_X1    g23194(.A1(new_n22906_), .A2(new_n22723_), .A3(new_n22728_), .ZN(new_n23387_));
  INV_X1     g23195(.I(new_n23387_), .ZN(new_n23388_));
  AOI22_X1   g23196(.A1(new_n23388_), .A2(new_n22927_), .B1(\asqrt[3] ), .B2(new_n23386_), .ZN(new_n23389_));
  INV_X1     g23197(.I(new_n23389_), .ZN(new_n23390_));
  NAND2_X1   g23198(.A1(new_n23373_), .A2(new_n2229_), .ZN(new_n23391_));
  OAI21_X1   g23199(.A1(new_n23384_), .A2(new_n23391_), .B(new_n23390_), .ZN(new_n23392_));
  AOI21_X1   g23200(.A1(new_n23392_), .A2(new_n23385_), .B(new_n1956_), .ZN(new_n23393_));
  INV_X1     g23201(.I(new_n22730_), .ZN(new_n23394_));
  NOR2_X1    g23202(.A1(new_n22729_), .A2(new_n22737_), .ZN(new_n23395_));
  NOR3_X1    g23203(.A1(new_n22906_), .A2(new_n23394_), .A3(new_n23395_), .ZN(new_n23396_));
  INV_X1     g23204(.I(new_n23396_), .ZN(new_n23397_));
  NOR3_X1    g23205(.A1(new_n23394_), .A2(new_n23395_), .A3(new_n22736_), .ZN(new_n23398_));
  AOI22_X1   g23206(.A1(new_n23397_), .A2(new_n22736_), .B1(\asqrt[3] ), .B2(new_n23398_), .ZN(new_n23399_));
  OAI21_X1   g23207(.A1(new_n23382_), .A2(new_n23383_), .B(new_n23373_), .ZN(new_n23400_));
  AOI21_X1   g23208(.A1(new_n23400_), .A2(\asqrt[47] ), .B(\asqrt[48] ), .ZN(new_n23401_));
  AOI21_X1   g23209(.A1(new_n23401_), .A2(new_n23392_), .B(new_n23399_), .ZN(new_n23402_));
  OAI21_X1   g23210(.A1(new_n23402_), .A2(new_n23393_), .B(\asqrt[49] ), .ZN(new_n23403_));
  INV_X1     g23211(.I(new_n23403_), .ZN(new_n23404_));
  INV_X1     g23212(.I(new_n22744_), .ZN(new_n23405_));
  INV_X1     g23213(.I(new_n22738_), .ZN(new_n23406_));
  INV_X1     g23214(.I(new_n22746_), .ZN(new_n23407_));
  NOR2_X1    g23215(.A1(new_n23407_), .A2(new_n23406_), .ZN(new_n23408_));
  NOR3_X1    g23216(.A1(new_n23408_), .A2(new_n22739_), .A3(new_n23405_), .ZN(new_n23409_));
  NOR3_X1    g23217(.A1(new_n22906_), .A2(new_n22739_), .A3(new_n23408_), .ZN(new_n23410_));
  INV_X1     g23218(.I(new_n23410_), .ZN(new_n23411_));
  AOI22_X1   g23219(.A1(new_n23411_), .A2(new_n23405_), .B1(\asqrt[3] ), .B2(new_n23409_), .ZN(new_n23412_));
  NOR3_X1    g23220(.A1(new_n23402_), .A2(new_n23393_), .A3(\asqrt[49] ), .ZN(new_n23413_));
  NOR2_X1    g23221(.A1(new_n23413_), .A2(new_n23412_), .ZN(new_n23414_));
  OAI21_X1   g23222(.A1(new_n23414_), .A2(new_n23404_), .B(\asqrt[50] ), .ZN(new_n23415_));
  NOR3_X1    g23223(.A1(new_n22906_), .A2(new_n22749_), .A3(new_n22754_), .ZN(new_n23416_));
  INV_X1     g23224(.I(new_n23416_), .ZN(new_n23417_));
  NOR3_X1    g23225(.A1(new_n22749_), .A2(new_n22926_), .A3(new_n22754_), .ZN(new_n23418_));
  AOI22_X1   g23226(.A1(new_n23417_), .A2(new_n22926_), .B1(\asqrt[3] ), .B2(new_n23418_), .ZN(new_n23419_));
  INV_X1     g23227(.I(new_n23419_), .ZN(new_n23420_));
  NAND2_X1   g23228(.A1(new_n23403_), .A2(new_n1612_), .ZN(new_n23421_));
  OAI21_X1   g23229(.A1(new_n23414_), .A2(new_n23421_), .B(new_n23420_), .ZN(new_n23422_));
  AOI21_X1   g23230(.A1(new_n23422_), .A2(new_n23415_), .B(new_n1376_), .ZN(new_n23423_));
  INV_X1     g23231(.I(new_n22756_), .ZN(new_n23424_));
  NOR2_X1    g23232(.A1(new_n22755_), .A2(new_n22763_), .ZN(new_n23425_));
  NOR3_X1    g23233(.A1(new_n23424_), .A2(new_n22762_), .A3(new_n23425_), .ZN(new_n23426_));
  NOR3_X1    g23234(.A1(new_n22906_), .A2(new_n23424_), .A3(new_n23425_), .ZN(new_n23427_));
  INV_X1     g23235(.I(new_n23427_), .ZN(new_n23428_));
  AOI22_X1   g23236(.A1(new_n23428_), .A2(new_n22762_), .B1(\asqrt[3] ), .B2(new_n23426_), .ZN(new_n23429_));
  OAI21_X1   g23237(.A1(new_n23412_), .A2(new_n23413_), .B(new_n23403_), .ZN(new_n23430_));
  AOI21_X1   g23238(.A1(new_n23430_), .A2(\asqrt[50] ), .B(\asqrt[51] ), .ZN(new_n23431_));
  AOI21_X1   g23239(.A1(new_n23431_), .A2(new_n23422_), .B(new_n23429_), .ZN(new_n23432_));
  OAI21_X1   g23240(.A1(new_n23432_), .A2(new_n23423_), .B(\asqrt[52] ), .ZN(new_n23433_));
  INV_X1     g23241(.I(new_n23433_), .ZN(new_n23434_));
  INV_X1     g23242(.I(new_n22770_), .ZN(new_n23435_));
  INV_X1     g23243(.I(new_n22764_), .ZN(new_n23436_));
  INV_X1     g23244(.I(new_n22772_), .ZN(new_n23437_));
  NOR2_X1    g23245(.A1(new_n23437_), .A2(new_n23436_), .ZN(new_n23438_));
  NOR3_X1    g23246(.A1(new_n22906_), .A2(new_n22765_), .A3(new_n23438_), .ZN(new_n23439_));
  INV_X1     g23247(.I(new_n23439_), .ZN(new_n23440_));
  NOR3_X1    g23248(.A1(new_n23438_), .A2(new_n22765_), .A3(new_n23435_), .ZN(new_n23441_));
  AOI22_X1   g23249(.A1(new_n23440_), .A2(new_n23435_), .B1(\asqrt[3] ), .B2(new_n23441_), .ZN(new_n23442_));
  NOR3_X1    g23250(.A1(new_n23432_), .A2(new_n23423_), .A3(\asqrt[52] ), .ZN(new_n23443_));
  NOR2_X1    g23251(.A1(new_n23443_), .A2(new_n23442_), .ZN(new_n23444_));
  OAI21_X1   g23252(.A1(new_n23444_), .A2(new_n23434_), .B(\asqrt[53] ), .ZN(new_n23445_));
  NOR3_X1    g23253(.A1(new_n22775_), .A2(new_n22925_), .A3(new_n22817_), .ZN(new_n23446_));
  NOR3_X1    g23254(.A1(new_n22906_), .A2(new_n22775_), .A3(new_n22817_), .ZN(new_n23447_));
  INV_X1     g23255(.I(new_n23447_), .ZN(new_n23448_));
  AOI22_X1   g23256(.A1(new_n23448_), .A2(new_n22925_), .B1(\asqrt[3] ), .B2(new_n23446_), .ZN(new_n23449_));
  INV_X1     g23257(.I(new_n23449_), .ZN(new_n23450_));
  NAND2_X1   g23258(.A1(new_n23433_), .A2(new_n1103_), .ZN(new_n23451_));
  OAI21_X1   g23259(.A1(new_n23444_), .A2(new_n23451_), .B(new_n23450_), .ZN(new_n23452_));
  AOI21_X1   g23260(.A1(new_n23452_), .A2(new_n23445_), .B(new_n904_), .ZN(new_n23453_));
  INV_X1     g23261(.I(new_n22783_), .ZN(new_n23454_));
  NOR2_X1    g23262(.A1(new_n22790_), .A2(new_n22782_), .ZN(new_n23455_));
  NOR3_X1    g23263(.A1(new_n22906_), .A2(new_n23454_), .A3(new_n23455_), .ZN(new_n23456_));
  INV_X1     g23264(.I(new_n23456_), .ZN(new_n23457_));
  NOR3_X1    g23265(.A1(new_n23454_), .A2(new_n22789_), .A3(new_n23455_), .ZN(new_n23458_));
  AOI22_X1   g23266(.A1(new_n23457_), .A2(new_n22789_), .B1(\asqrt[3] ), .B2(new_n23458_), .ZN(new_n23459_));
  OAI21_X1   g23267(.A1(new_n23442_), .A2(new_n23443_), .B(new_n23433_), .ZN(new_n23460_));
  AOI21_X1   g23268(.A1(new_n23460_), .A2(\asqrt[53] ), .B(\asqrt[54] ), .ZN(new_n23461_));
  AOI21_X1   g23269(.A1(new_n23461_), .A2(new_n23452_), .B(new_n23459_), .ZN(new_n23462_));
  OAI21_X1   g23270(.A1(new_n23462_), .A2(new_n23453_), .B(\asqrt[55] ), .ZN(new_n23463_));
  INV_X1     g23271(.I(new_n23463_), .ZN(new_n23464_));
  NOR2_X1    g23272(.A1(new_n22801_), .A2(new_n22794_), .ZN(new_n23465_));
  NOR3_X1    g23273(.A1(new_n23465_), .A2(new_n22792_), .A3(new_n22800_), .ZN(new_n23466_));
  NOR3_X1    g23274(.A1(new_n22906_), .A2(new_n22792_), .A3(new_n23465_), .ZN(new_n23467_));
  INV_X1     g23275(.I(new_n23467_), .ZN(new_n23468_));
  AOI22_X1   g23276(.A1(new_n23468_), .A2(new_n22800_), .B1(\asqrt[3] ), .B2(new_n23466_), .ZN(new_n23469_));
  NOR3_X1    g23277(.A1(new_n23462_), .A2(new_n23453_), .A3(\asqrt[55] ), .ZN(new_n23470_));
  NOR2_X1    g23278(.A1(new_n23470_), .A2(new_n23469_), .ZN(new_n23471_));
  OAI21_X1   g23279(.A1(new_n23471_), .A2(new_n23464_), .B(\asqrt[56] ), .ZN(new_n23472_));
  NOR3_X1    g23280(.A1(new_n22906_), .A2(new_n22803_), .A3(new_n22849_), .ZN(new_n23473_));
  INV_X1     g23281(.I(new_n23473_), .ZN(new_n23474_));
  NOR3_X1    g23282(.A1(new_n22803_), .A2(new_n22924_), .A3(new_n22849_), .ZN(new_n23475_));
  AOI22_X1   g23283(.A1(new_n23474_), .A2(new_n22924_), .B1(\asqrt[3] ), .B2(new_n23475_), .ZN(new_n23476_));
  INV_X1     g23284(.I(new_n23476_), .ZN(new_n23477_));
  NAND2_X1   g23285(.A1(new_n23463_), .A2(new_n703_), .ZN(new_n23478_));
  OAI21_X1   g23286(.A1(new_n23471_), .A2(new_n23478_), .B(new_n23477_), .ZN(new_n23479_));
  AOI21_X1   g23287(.A1(new_n23479_), .A2(new_n23472_), .B(new_n531_), .ZN(new_n23480_));
  INV_X1     g23288(.I(new_n22810_), .ZN(new_n23481_));
  NOR2_X1    g23289(.A1(new_n22822_), .A2(new_n22809_), .ZN(new_n23482_));
  NOR3_X1    g23290(.A1(new_n23481_), .A2(new_n22816_), .A3(new_n23482_), .ZN(new_n23483_));
  NOR3_X1    g23291(.A1(new_n22906_), .A2(new_n23481_), .A3(new_n23482_), .ZN(new_n23484_));
  INV_X1     g23292(.I(new_n23484_), .ZN(new_n23485_));
  AOI22_X1   g23293(.A1(new_n23485_), .A2(new_n22816_), .B1(\asqrt[3] ), .B2(new_n23483_), .ZN(new_n23486_));
  OAI21_X1   g23294(.A1(new_n23469_), .A2(new_n23470_), .B(new_n23463_), .ZN(new_n23487_));
  AOI21_X1   g23295(.A1(new_n23487_), .A2(\asqrt[56] ), .B(\asqrt[57] ), .ZN(new_n23488_));
  AOI21_X1   g23296(.A1(new_n23488_), .A2(new_n23479_), .B(new_n23486_), .ZN(new_n23489_));
  OAI21_X1   g23297(.A1(new_n23489_), .A2(new_n23480_), .B(\asqrt[58] ), .ZN(new_n23490_));
  NOR2_X1    g23298(.A1(new_n22833_), .A2(new_n22826_), .ZN(new_n23491_));
  NOR3_X1    g23299(.A1(new_n22906_), .A2(new_n22824_), .A3(new_n23491_), .ZN(new_n23492_));
  INV_X1     g23300(.I(new_n23492_), .ZN(new_n23493_));
  NOR3_X1    g23301(.A1(new_n23491_), .A2(new_n22824_), .A3(new_n22832_), .ZN(new_n23494_));
  AOI22_X1   g23302(.A1(new_n23493_), .A2(new_n22832_), .B1(\asqrt[3] ), .B2(new_n23494_), .ZN(new_n23495_));
  INV_X1     g23303(.I(new_n23495_), .ZN(new_n23496_));
  INV_X1     g23304(.I(new_n23469_), .ZN(new_n23497_));
  INV_X1     g23305(.I(new_n23442_), .ZN(new_n23498_));
  INV_X1     g23306(.I(new_n23412_), .ZN(new_n23499_));
  INV_X1     g23307(.I(new_n23382_), .ZN(new_n23500_));
  INV_X1     g23308(.I(new_n23352_), .ZN(new_n23501_));
  INV_X1     g23309(.I(new_n23324_), .ZN(new_n23502_));
  INV_X1     g23310(.I(new_n23298_), .ZN(new_n23503_));
  INV_X1     g23311(.I(new_n23271_), .ZN(new_n23504_));
  INV_X1     g23312(.I(new_n23244_), .ZN(new_n23505_));
  INV_X1     g23313(.I(new_n23217_), .ZN(new_n23506_));
  INV_X1     g23314(.I(new_n23187_), .ZN(new_n23507_));
  INV_X1     g23315(.I(new_n23157_), .ZN(new_n23508_));
  INV_X1     g23316(.I(new_n23127_), .ZN(new_n23509_));
  INV_X1     g23317(.I(new_n23097_), .ZN(new_n23510_));
  INV_X1     g23318(.I(new_n23066_), .ZN(new_n23511_));
  INV_X1     g23319(.I(new_n23041_), .ZN(new_n23512_));
  NAND2_X1   g23320(.A1(new_n22982_), .A2(new_n20262_), .ZN(new_n23513_));
  OAI21_X1   g23321(.A1(new_n23513_), .A2(new_n23015_), .B(new_n22996_), .ZN(new_n23514_));
  AOI21_X1   g23322(.A1(new_n23514_), .A2(new_n23025_), .B(new_n19573_), .ZN(new_n23515_));
  NOR2_X1    g23323(.A1(new_n22990_), .A2(\asqrt[8] ), .ZN(new_n23516_));
  AOI21_X1   g23324(.A1(new_n23516_), .A2(new_n23514_), .B(new_n23023_), .ZN(new_n23517_));
  OAI21_X1   g23325(.A1(new_n23517_), .A2(new_n23515_), .B(\asqrt[9] ), .ZN(new_n23518_));
  NAND2_X1   g23326(.A1(new_n23518_), .A2(new_n18275_), .ZN(new_n23519_));
  OAI21_X1   g23327(.A1(new_n23519_), .A2(new_n23035_), .B(new_n23512_), .ZN(new_n23520_));
  NAND3_X1   g23328(.A1(new_n23520_), .A2(new_n17623_), .A3(new_n23036_), .ZN(new_n23521_));
  AOI22_X1   g23329(.A1(new_n23521_), .A2(new_n23050_), .B1(\asqrt[11] ), .B2(new_n23058_), .ZN(new_n23522_));
  OAI21_X1   g23330(.A1(new_n23522_), .A2(new_n16881_), .B(new_n16389_), .ZN(new_n23523_));
  OAI21_X1   g23331(.A1(new_n23523_), .A2(new_n23060_), .B(new_n23511_), .ZN(new_n23524_));
  AOI21_X1   g23332(.A1(new_n23524_), .A2(new_n23061_), .B(new_n15770_), .ZN(new_n23525_));
  AOI21_X1   g23333(.A1(new_n23520_), .A2(new_n23036_), .B(new_n17623_), .ZN(new_n23526_));
  NOR3_X1    g23334(.A1(new_n23517_), .A2(new_n23515_), .A3(\asqrt[9] ), .ZN(new_n23527_));
  OAI21_X1   g23335(.A1(new_n23032_), .A2(new_n23527_), .B(new_n23518_), .ZN(new_n23528_));
  AOI21_X1   g23336(.A1(new_n23528_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n23529_));
  AOI21_X1   g23337(.A1(new_n23529_), .A2(new_n23520_), .B(new_n23049_), .ZN(new_n23530_));
  NOR3_X1    g23338(.A1(new_n23530_), .A2(\asqrt[12] ), .A3(new_n23526_), .ZN(new_n23531_));
  OAI22_X1   g23339(.A1(new_n23531_), .A2(new_n23057_), .B1(new_n23522_), .B2(new_n16881_), .ZN(new_n23532_));
  AOI21_X1   g23340(.A1(new_n23532_), .A2(\asqrt[13] ), .B(\asqrt[14] ), .ZN(new_n23533_));
  AOI21_X1   g23341(.A1(new_n23533_), .A2(new_n23524_), .B(new_n23074_), .ZN(new_n23534_));
  OAI21_X1   g23342(.A1(new_n23534_), .A2(new_n23525_), .B(\asqrt[15] ), .ZN(new_n23535_));
  NAND2_X1   g23343(.A1(new_n23535_), .A2(new_n14601_), .ZN(new_n23536_));
  OAI21_X1   g23344(.A1(new_n23536_), .A2(new_n23087_), .B(new_n23510_), .ZN(new_n23537_));
  AOI21_X1   g23345(.A1(new_n23537_), .A2(new_n23088_), .B(new_n14017_), .ZN(new_n23538_));
  NOR3_X1    g23346(.A1(new_n23534_), .A2(\asqrt[15] ), .A3(new_n23525_), .ZN(new_n23539_));
  OAI21_X1   g23347(.A1(new_n23084_), .A2(new_n23539_), .B(new_n23535_), .ZN(new_n23540_));
  AOI21_X1   g23348(.A1(new_n23540_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n23541_));
  AOI21_X1   g23349(.A1(new_n23541_), .A2(new_n23537_), .B(new_n23105_), .ZN(new_n23542_));
  OAI21_X1   g23350(.A1(new_n23542_), .A2(new_n23538_), .B(\asqrt[18] ), .ZN(new_n23543_));
  NAND2_X1   g23351(.A1(new_n23543_), .A2(new_n12913_), .ZN(new_n23544_));
  OAI21_X1   g23352(.A1(new_n23544_), .A2(new_n23117_), .B(new_n23509_), .ZN(new_n23545_));
  AOI21_X1   g23353(.A1(new_n23545_), .A2(new_n23118_), .B(new_n12364_), .ZN(new_n23546_));
  NOR3_X1    g23354(.A1(new_n23542_), .A2(\asqrt[18] ), .A3(new_n23538_), .ZN(new_n23547_));
  OAI21_X1   g23355(.A1(new_n23114_), .A2(new_n23547_), .B(new_n23543_), .ZN(new_n23548_));
  AOI21_X1   g23356(.A1(new_n23548_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n23549_));
  AOI21_X1   g23357(.A1(new_n23549_), .A2(new_n23545_), .B(new_n23135_), .ZN(new_n23550_));
  OAI21_X1   g23358(.A1(new_n23550_), .A2(new_n23546_), .B(\asqrt[21] ), .ZN(new_n23551_));
  NAND2_X1   g23359(.A1(new_n23551_), .A2(new_n11326_), .ZN(new_n23552_));
  OAI21_X1   g23360(.A1(new_n23552_), .A2(new_n23147_), .B(new_n23508_), .ZN(new_n23553_));
  AOI21_X1   g23361(.A1(new_n23553_), .A2(new_n23148_), .B(new_n10812_), .ZN(new_n23554_));
  NOR3_X1    g23362(.A1(new_n23550_), .A2(\asqrt[21] ), .A3(new_n23546_), .ZN(new_n23555_));
  OAI21_X1   g23363(.A1(new_n23144_), .A2(new_n23555_), .B(new_n23551_), .ZN(new_n23556_));
  AOI21_X1   g23364(.A1(new_n23556_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n23557_));
  AOI21_X1   g23365(.A1(new_n23557_), .A2(new_n23553_), .B(new_n23165_), .ZN(new_n23558_));
  OAI21_X1   g23366(.A1(new_n23558_), .A2(new_n23554_), .B(\asqrt[24] ), .ZN(new_n23559_));
  NAND2_X1   g23367(.A1(new_n23559_), .A2(new_n9846_), .ZN(new_n23560_));
  OAI21_X1   g23368(.A1(new_n23560_), .A2(new_n23177_), .B(new_n23507_), .ZN(new_n23561_));
  AOI21_X1   g23369(.A1(new_n23561_), .A2(new_n23178_), .B(new_n9317_), .ZN(new_n23562_));
  NOR3_X1    g23370(.A1(new_n23558_), .A2(\asqrt[24] ), .A3(new_n23554_), .ZN(new_n23563_));
  OAI21_X1   g23371(.A1(new_n23174_), .A2(new_n23563_), .B(new_n23559_), .ZN(new_n23564_));
  AOI21_X1   g23372(.A1(new_n23564_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n23565_));
  AOI21_X1   g23373(.A1(new_n23565_), .A2(new_n23561_), .B(new_n23195_), .ZN(new_n23566_));
  OAI21_X1   g23374(.A1(new_n23566_), .A2(new_n23562_), .B(\asqrt[27] ), .ZN(new_n23567_));
  NAND2_X1   g23375(.A1(new_n23567_), .A2(new_n8483_), .ZN(new_n23568_));
  OAI21_X1   g23376(.A1(new_n23568_), .A2(new_n23207_), .B(new_n23506_), .ZN(new_n23569_));
  AOI21_X1   g23377(.A1(new_n23569_), .A2(new_n23208_), .B(new_n8036_), .ZN(new_n23570_));
  NOR3_X1    g23378(.A1(new_n23566_), .A2(\asqrt[27] ), .A3(new_n23562_), .ZN(new_n23571_));
  OAI21_X1   g23379(.A1(new_n23204_), .A2(new_n23571_), .B(new_n23567_), .ZN(new_n23572_));
  AOI21_X1   g23380(.A1(new_n23572_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n23573_));
  AOI21_X1   g23381(.A1(new_n23573_), .A2(new_n23569_), .B(new_n23225_), .ZN(new_n23574_));
  OAI21_X1   g23382(.A1(new_n23574_), .A2(new_n23570_), .B(\asqrt[30] ), .ZN(new_n23575_));
  NAND2_X1   g23383(.A1(new_n23575_), .A2(new_n7229_), .ZN(new_n23576_));
  OAI21_X1   g23384(.A1(new_n23576_), .A2(new_n23237_), .B(new_n23505_), .ZN(new_n23577_));
  AOI21_X1   g23385(.A1(new_n23577_), .A2(new_n23238_), .B(new_n6824_), .ZN(new_n23578_));
  NOR3_X1    g23386(.A1(new_n23574_), .A2(\asqrt[30] ), .A3(new_n23570_), .ZN(new_n23579_));
  OAI21_X1   g23387(.A1(new_n23234_), .A2(new_n23579_), .B(new_n23575_), .ZN(new_n23580_));
  AOI21_X1   g23388(.A1(new_n23580_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n23581_));
  AOI21_X1   g23389(.A1(new_n23581_), .A2(new_n23577_), .B(new_n23252_), .ZN(new_n23582_));
  OAI21_X1   g23390(.A1(new_n23582_), .A2(new_n23578_), .B(\asqrt[33] ), .ZN(new_n23583_));
  NAND2_X1   g23391(.A1(new_n23583_), .A2(new_n6077_), .ZN(new_n23584_));
  OAI21_X1   g23392(.A1(new_n23584_), .A2(new_n23264_), .B(new_n23504_), .ZN(new_n23585_));
  AOI21_X1   g23393(.A1(new_n23585_), .A2(new_n23265_), .B(new_n5708_), .ZN(new_n23586_));
  NOR3_X1    g23394(.A1(new_n23582_), .A2(\asqrt[33] ), .A3(new_n23578_), .ZN(new_n23587_));
  OAI21_X1   g23395(.A1(new_n23261_), .A2(new_n23587_), .B(new_n23583_), .ZN(new_n23588_));
  AOI21_X1   g23396(.A1(new_n23588_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n23589_));
  AOI21_X1   g23397(.A1(new_n23589_), .A2(new_n23585_), .B(new_n23279_), .ZN(new_n23590_));
  OAI21_X1   g23398(.A1(new_n23590_), .A2(new_n23586_), .B(\asqrt[36] ), .ZN(new_n23591_));
  NAND2_X1   g23399(.A1(new_n23591_), .A2(new_n5024_), .ZN(new_n23592_));
  OAI21_X1   g23400(.A1(new_n23592_), .A2(new_n23291_), .B(new_n23503_), .ZN(new_n23593_));
  AOI21_X1   g23401(.A1(new_n23593_), .A2(new_n23292_), .B(new_n4696_), .ZN(new_n23594_));
  NOR3_X1    g23402(.A1(new_n23590_), .A2(\asqrt[36] ), .A3(new_n23586_), .ZN(new_n23595_));
  OAI21_X1   g23403(.A1(new_n23288_), .A2(new_n23595_), .B(new_n23591_), .ZN(new_n23596_));
  AOI21_X1   g23404(.A1(new_n23596_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n23597_));
  AOI21_X1   g23405(.A1(new_n23597_), .A2(new_n23593_), .B(new_n23306_), .ZN(new_n23598_));
  OAI21_X1   g23406(.A1(new_n23598_), .A2(new_n23594_), .B(\asqrt[39] ), .ZN(new_n23599_));
  NAND2_X1   g23407(.A1(new_n23599_), .A2(new_n4071_), .ZN(new_n23600_));
  OAI21_X1   g23408(.A1(new_n23600_), .A2(new_n23317_), .B(new_n23502_), .ZN(new_n23601_));
  AOI21_X1   g23409(.A1(new_n23601_), .A2(new_n23318_), .B(new_n3782_), .ZN(new_n23602_));
  NOR3_X1    g23410(.A1(new_n23598_), .A2(\asqrt[39] ), .A3(new_n23594_), .ZN(new_n23603_));
  OAI21_X1   g23411(.A1(new_n23314_), .A2(new_n23603_), .B(new_n23599_), .ZN(new_n23604_));
  AOI21_X1   g23412(.A1(new_n23604_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n23605_));
  AOI21_X1   g23413(.A1(new_n23605_), .A2(new_n23601_), .B(new_n23332_), .ZN(new_n23606_));
  OAI21_X1   g23414(.A1(new_n23606_), .A2(new_n23602_), .B(\asqrt[42] ), .ZN(new_n23607_));
  NAND2_X1   g23415(.A1(new_n23607_), .A2(new_n3218_), .ZN(new_n23608_));
  OAI21_X1   g23416(.A1(new_n23608_), .A2(new_n23343_), .B(new_n23501_), .ZN(new_n23609_));
  AOI21_X1   g23417(.A1(new_n23609_), .A2(new_n23344_), .B(new_n2954_), .ZN(new_n23610_));
  NOR3_X1    g23418(.A1(new_n23606_), .A2(\asqrt[42] ), .A3(new_n23602_), .ZN(new_n23611_));
  OAI21_X1   g23419(.A1(new_n23340_), .A2(new_n23611_), .B(new_n23607_), .ZN(new_n23612_));
  AOI21_X1   g23420(.A1(new_n23612_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n23613_));
  AOI21_X1   g23421(.A1(new_n23613_), .A2(new_n23609_), .B(new_n23359_), .ZN(new_n23614_));
  OAI21_X1   g23422(.A1(new_n23614_), .A2(new_n23610_), .B(\asqrt[45] ), .ZN(new_n23615_));
  NAND2_X1   g23423(.A1(new_n23615_), .A2(new_n2465_), .ZN(new_n23616_));
  OAI21_X1   g23424(.A1(new_n23616_), .A2(new_n23372_), .B(new_n23500_), .ZN(new_n23617_));
  AOI21_X1   g23425(.A1(new_n23617_), .A2(new_n23373_), .B(new_n2229_), .ZN(new_n23618_));
  NOR3_X1    g23426(.A1(new_n23614_), .A2(\asqrt[45] ), .A3(new_n23610_), .ZN(new_n23619_));
  OAI21_X1   g23427(.A1(new_n23369_), .A2(new_n23619_), .B(new_n23615_), .ZN(new_n23620_));
  AOI21_X1   g23428(.A1(new_n23620_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n23621_));
  AOI21_X1   g23429(.A1(new_n23621_), .A2(new_n23617_), .B(new_n23389_), .ZN(new_n23622_));
  OAI21_X1   g23430(.A1(new_n23622_), .A2(new_n23618_), .B(\asqrt[48] ), .ZN(new_n23623_));
  NAND2_X1   g23431(.A1(new_n23623_), .A2(new_n1806_), .ZN(new_n23624_));
  OAI21_X1   g23432(.A1(new_n23624_), .A2(new_n23402_), .B(new_n23499_), .ZN(new_n23625_));
  AOI21_X1   g23433(.A1(new_n23625_), .A2(new_n23403_), .B(new_n1612_), .ZN(new_n23626_));
  NOR3_X1    g23434(.A1(new_n23622_), .A2(\asqrt[48] ), .A3(new_n23618_), .ZN(new_n23627_));
  OAI21_X1   g23435(.A1(new_n23399_), .A2(new_n23627_), .B(new_n23623_), .ZN(new_n23628_));
  AOI21_X1   g23436(.A1(new_n23628_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n23629_));
  AOI21_X1   g23437(.A1(new_n23629_), .A2(new_n23625_), .B(new_n23419_), .ZN(new_n23630_));
  OAI21_X1   g23438(.A1(new_n23630_), .A2(new_n23626_), .B(\asqrt[51] ), .ZN(new_n23631_));
  NAND2_X1   g23439(.A1(new_n23631_), .A2(new_n1256_), .ZN(new_n23632_));
  OAI21_X1   g23440(.A1(new_n23632_), .A2(new_n23432_), .B(new_n23498_), .ZN(new_n23633_));
  NAND3_X1   g23441(.A1(new_n23633_), .A2(new_n1103_), .A3(new_n23433_), .ZN(new_n23634_));
  AOI22_X1   g23442(.A1(new_n23634_), .A2(new_n23450_), .B1(\asqrt[53] ), .B2(new_n23460_), .ZN(new_n23635_));
  OAI21_X1   g23443(.A1(new_n23635_), .A2(new_n904_), .B(new_n823_), .ZN(new_n23636_));
  OAI21_X1   g23444(.A1(new_n23636_), .A2(new_n23462_), .B(new_n23497_), .ZN(new_n23637_));
  NAND3_X1   g23445(.A1(new_n23637_), .A2(new_n703_), .A3(new_n23463_), .ZN(new_n23638_));
  AOI22_X1   g23446(.A1(new_n23638_), .A2(new_n23477_), .B1(\asqrt[56] ), .B2(new_n23487_), .ZN(new_n23639_));
  OAI21_X1   g23447(.A1(new_n23639_), .A2(new_n531_), .B(new_n436_), .ZN(new_n23640_));
  OAI21_X1   g23448(.A1(new_n23640_), .A2(new_n23489_), .B(new_n23496_), .ZN(new_n23641_));
  AOI21_X1   g23449(.A1(new_n23641_), .A2(new_n23490_), .B(new_n327_), .ZN(new_n23642_));
  NOR3_X1    g23450(.A1(new_n22835_), .A2(new_n22923_), .A3(new_n22881_), .ZN(new_n23643_));
  NOR3_X1    g23451(.A1(new_n22906_), .A2(new_n22835_), .A3(new_n22881_), .ZN(new_n23644_));
  INV_X1     g23452(.I(new_n23644_), .ZN(new_n23645_));
  AOI22_X1   g23453(.A1(new_n23645_), .A2(new_n22923_), .B1(\asqrt[3] ), .B2(new_n23643_), .ZN(new_n23646_));
  NAND2_X1   g23454(.A1(new_n23490_), .A2(new_n327_), .ZN(new_n23647_));
  INV_X1     g23455(.I(new_n23647_), .ZN(new_n23648_));
  AOI21_X1   g23456(.A1(new_n23648_), .A2(new_n23641_), .B(new_n23646_), .ZN(new_n23649_));
  OAI21_X1   g23457(.A1(new_n23649_), .A2(new_n23642_), .B(\asqrt[60] ), .ZN(new_n23650_));
  INV_X1     g23458(.I(new_n22842_), .ZN(new_n23651_));
  NOR2_X1    g23459(.A1(new_n22854_), .A2(new_n22841_), .ZN(new_n23652_));
  NOR3_X1    g23460(.A1(new_n22906_), .A2(new_n23651_), .A3(new_n23652_), .ZN(new_n23653_));
  INV_X1     g23461(.I(new_n23653_), .ZN(new_n23654_));
  NOR3_X1    g23462(.A1(new_n23651_), .A2(new_n22848_), .A3(new_n23652_), .ZN(new_n23655_));
  AOI22_X1   g23463(.A1(new_n23654_), .A2(new_n22848_), .B1(\asqrt[3] ), .B2(new_n23655_), .ZN(new_n23656_));
  INV_X1     g23464(.I(new_n23656_), .ZN(new_n23657_));
  INV_X1     g23465(.I(new_n23490_), .ZN(new_n23658_));
  NOR3_X1    g23466(.A1(new_n23489_), .A2(new_n23480_), .A3(\asqrt[58] ), .ZN(new_n23659_));
  NOR2_X1    g23467(.A1(new_n23659_), .A2(new_n23495_), .ZN(new_n23660_));
  OAI21_X1   g23468(.A1(new_n23660_), .A2(new_n23658_), .B(\asqrt[59] ), .ZN(new_n23661_));
  NAND2_X1   g23469(.A1(new_n23661_), .A2(new_n306_), .ZN(new_n23662_));
  OAI21_X1   g23470(.A1(new_n23662_), .A2(new_n23649_), .B(new_n23657_), .ZN(new_n23663_));
  AOI21_X1   g23471(.A1(new_n23663_), .A2(new_n23650_), .B(new_n218_), .ZN(new_n23664_));
  NOR2_X1    g23472(.A1(new_n22858_), .A2(new_n22865_), .ZN(new_n23665_));
  NOR3_X1    g23473(.A1(new_n23665_), .A2(new_n22856_), .A3(new_n22864_), .ZN(new_n23666_));
  NOR3_X1    g23474(.A1(new_n22906_), .A2(new_n22856_), .A3(new_n23665_), .ZN(new_n23667_));
  INV_X1     g23475(.I(new_n23667_), .ZN(new_n23668_));
  AOI22_X1   g23476(.A1(new_n23668_), .A2(new_n22864_), .B1(\asqrt[3] ), .B2(new_n23666_), .ZN(new_n23669_));
  INV_X1     g23477(.I(new_n23646_), .ZN(new_n23670_));
  OAI21_X1   g23478(.A1(new_n23660_), .A2(new_n23647_), .B(new_n23670_), .ZN(new_n23671_));
  AOI21_X1   g23479(.A1(new_n23671_), .A2(new_n23661_), .B(new_n306_), .ZN(new_n23672_));
  NOR2_X1    g23480(.A1(new_n23672_), .A2(\asqrt[61] ), .ZN(new_n23673_));
  AOI21_X1   g23481(.A1(new_n23673_), .A2(new_n23663_), .B(new_n23669_), .ZN(new_n23674_));
  OAI21_X1   g23482(.A1(new_n23674_), .A2(new_n23664_), .B(\asqrt[62] ), .ZN(new_n23675_));
  NOR3_X1    g23483(.A1(new_n22906_), .A2(new_n22867_), .A3(new_n22920_), .ZN(new_n23676_));
  INV_X1     g23484(.I(new_n23676_), .ZN(new_n23677_));
  NOR3_X1    g23485(.A1(new_n22867_), .A2(new_n22922_), .A3(new_n22920_), .ZN(new_n23678_));
  AOI22_X1   g23486(.A1(new_n23677_), .A2(new_n22922_), .B1(\asqrt[3] ), .B2(new_n23678_), .ZN(new_n23679_));
  INV_X1     g23487(.I(new_n23679_), .ZN(new_n23680_));
  OAI21_X1   g23488(.A1(new_n23495_), .A2(new_n23659_), .B(new_n23490_), .ZN(new_n23681_));
  AOI21_X1   g23489(.A1(new_n23681_), .A2(\asqrt[59] ), .B(\asqrt[60] ), .ZN(new_n23682_));
  AOI21_X1   g23490(.A1(new_n23682_), .A2(new_n23671_), .B(new_n23656_), .ZN(new_n23683_));
  OAI21_X1   g23491(.A1(new_n23683_), .A2(new_n23672_), .B(\asqrt[61] ), .ZN(new_n23684_));
  NAND2_X1   g23492(.A1(new_n23684_), .A2(new_n207_), .ZN(new_n23685_));
  OAI21_X1   g23493(.A1(new_n23685_), .A2(new_n23674_), .B(new_n23680_), .ZN(new_n23686_));
  NAND2_X1   g23494(.A1(new_n23686_), .A2(new_n23675_), .ZN(new_n23687_));
  NAND4_X1   g23495(.A1(\asqrt[3] ), .A2(new_n22874_), .A3(new_n22879_), .A4(new_n22959_), .ZN(new_n23688_));
  NAND2_X1   g23496(.A1(new_n22874_), .A2(new_n22959_), .ZN(new_n23689_));
  OAI21_X1   g23497(.A1(new_n22906_), .A2(new_n23689_), .B(new_n22880_), .ZN(new_n23690_));
  NAND2_X1   g23498(.A1(new_n23688_), .A2(new_n23690_), .ZN(new_n23691_));
  NOR2_X1    g23499(.A1(new_n22960_), .A2(new_n22900_), .ZN(new_n23692_));
  NAND2_X1   g23500(.A1(\asqrt[3] ), .A2(new_n23692_), .ZN(new_n23693_));
  NAND3_X1   g23501(.A1(new_n23691_), .A2(new_n22972_), .A3(new_n23693_), .ZN(new_n23694_));
  INV_X1     g23502(.I(new_n23694_), .ZN(new_n23695_));
  AOI21_X1   g23503(.A1(new_n23687_), .A2(new_n23695_), .B(\asqrt[63] ), .ZN(new_n23696_));
  INV_X1     g23504(.I(new_n23669_), .ZN(new_n23697_));
  NAND3_X1   g23505(.A1(new_n23641_), .A2(new_n327_), .A3(new_n23490_), .ZN(new_n23698_));
  AOI22_X1   g23506(.A1(new_n23698_), .A2(new_n23670_), .B1(new_n23681_), .B2(\asqrt[59] ), .ZN(new_n23699_));
  OAI21_X1   g23507(.A1(new_n23699_), .A2(new_n306_), .B(new_n218_), .ZN(new_n23700_));
  OAI21_X1   g23508(.A1(new_n23700_), .A2(new_n23683_), .B(new_n23697_), .ZN(new_n23701_));
  NOR2_X1    g23509(.A1(new_n23664_), .A2(\asqrt[62] ), .ZN(new_n23702_));
  AOI21_X1   g23510(.A1(new_n23702_), .A2(new_n23701_), .B(new_n23679_), .ZN(new_n23703_));
  INV_X1     g23511(.I(new_n23691_), .ZN(new_n23704_));
  NAND2_X1   g23512(.A1(new_n23675_), .A2(new_n23704_), .ZN(new_n23705_));
  INV_X1     g23513(.I(new_n22960_), .ZN(new_n23706_));
  NOR2_X1    g23514(.A1(new_n22906_), .A2(new_n22900_), .ZN(new_n23707_));
  NOR2_X1    g23515(.A1(new_n23692_), .A2(new_n193_), .ZN(new_n23708_));
  OAI21_X1   g23516(.A1(new_n23707_), .A2(new_n23706_), .B(new_n23708_), .ZN(new_n23709_));
  OAI21_X1   g23517(.A1(new_n23705_), .A2(new_n23703_), .B(new_n23709_), .ZN(new_n23710_));
  OAI21_X1   g23518(.A1(new_n23696_), .A2(new_n23710_), .B(\a[4] ), .ZN(new_n23711_));
  AOI21_X1   g23519(.A1(new_n23711_), .A2(new_n22911_), .B(new_n22906_), .ZN(new_n23712_));
  NOR3_X1    g23520(.A1(new_n23683_), .A2(new_n23672_), .A3(\asqrt[61] ), .ZN(new_n23713_));
  OAI21_X1   g23521(.A1(new_n23669_), .A2(new_n23713_), .B(new_n23684_), .ZN(new_n23714_));
  NAND3_X1   g23522(.A1(new_n23701_), .A2(new_n207_), .A3(new_n23684_), .ZN(new_n23715_));
  AOI22_X1   g23523(.A1(new_n23715_), .A2(new_n23680_), .B1(new_n23714_), .B2(\asqrt[62] ), .ZN(new_n23716_));
  OAI21_X1   g23524(.A1(new_n23716_), .A2(new_n23694_), .B(new_n193_), .ZN(new_n23717_));
  AOI21_X1   g23525(.A1(new_n23714_), .A2(\asqrt[62] ), .B(new_n23691_), .ZN(new_n23718_));
  INV_X1     g23526(.I(new_n23709_), .ZN(new_n23719_));
  AOI21_X1   g23527(.A1(new_n23718_), .A2(new_n23686_), .B(new_n23719_), .ZN(new_n23720_));
  AOI21_X1   g23528(.A1(new_n23717_), .A2(new_n23720_), .B(new_n22907_), .ZN(new_n23721_));
  NOR4_X1    g23529(.A1(new_n22975_), .A2(new_n22898_), .A3(new_n22963_), .A4(new_n22910_), .ZN(new_n23722_));
  INV_X1     g23530(.I(new_n23722_), .ZN(new_n23723_));
  NOR2_X1    g23531(.A1(new_n23721_), .A2(new_n23723_), .ZN(new_n23724_));
  AOI21_X1   g23532(.A1(new_n23717_), .A2(new_n23720_), .B(new_n22914_), .ZN(new_n23725_));
  INV_X1     g23533(.I(\a[5] ), .ZN(new_n23726_));
  AOI21_X1   g23534(.A1(new_n23686_), .A2(new_n23675_), .B(new_n23694_), .ZN(new_n23727_));
  OAI21_X1   g23535(.A1(\asqrt[63] ), .A2(new_n23727_), .B(new_n23720_), .ZN(\asqrt[2] ));
  AOI21_X1   g23536(.A1(\asqrt[2] ), .A2(new_n22907_), .B(new_n23726_), .ZN(new_n23729_));
  NOR3_X1    g23537(.A1(new_n23724_), .A2(new_n23729_), .A3(new_n23725_), .ZN(new_n23730_));
  OAI21_X1   g23538(.A1(new_n23730_), .A2(new_n23712_), .B(\asqrt[4] ), .ZN(new_n23731_));
  OAI21_X1   g23539(.A1(new_n23696_), .A2(new_n23710_), .B(new_n22913_), .ZN(new_n23732_));
  NAND2_X1   g23540(.A1(new_n23718_), .A2(new_n23686_), .ZN(new_n23733_));
  NAND4_X1   g23541(.A1(new_n23717_), .A2(\asqrt[3] ), .A3(new_n23733_), .A4(new_n23709_), .ZN(new_n23734_));
  AOI21_X1   g23542(.A1(new_n23734_), .A2(new_n23732_), .B(new_n22912_), .ZN(new_n23735_));
  NAND3_X1   g23543(.A1(new_n23733_), .A2(\asqrt[3] ), .A3(new_n23709_), .ZN(new_n23736_));
  NOR2_X1    g23544(.A1(new_n23736_), .A2(new_n23696_), .ZN(new_n23737_));
  NOR3_X1    g23545(.A1(new_n23737_), .A2(new_n23725_), .A3(\a[6] ), .ZN(new_n23738_));
  AOI21_X1   g23546(.A1(\asqrt[2] ), .A2(\a[4] ), .B(new_n22910_), .ZN(new_n23739_));
  OAI21_X1   g23547(.A1(new_n23739_), .A2(new_n22906_), .B(new_n22337_), .ZN(new_n23740_));
  OAI22_X1   g23548(.A1(new_n23730_), .A2(new_n23740_), .B1(new_n23735_), .B2(new_n23738_), .ZN(new_n23741_));
  AOI21_X1   g23549(.A1(new_n23741_), .A2(new_n23731_), .B(new_n21620_), .ZN(new_n23742_));
  NOR3_X1    g23550(.A1(new_n23000_), .A2(new_n23002_), .A3(new_n22967_), .ZN(new_n23743_));
  NAND3_X1   g23551(.A1(\asqrt[2] ), .A2(new_n22999_), .A3(new_n22919_), .ZN(new_n23744_));
  AOI22_X1   g23552(.A1(new_n23744_), .A2(new_n22967_), .B1(\asqrt[2] ), .B2(new_n23743_), .ZN(new_n23745_));
  OAI21_X1   g23553(.A1(new_n23721_), .A2(new_n22910_), .B(\asqrt[3] ), .ZN(new_n23746_));
  AOI21_X1   g23554(.A1(new_n23717_), .A2(new_n23720_), .B(\a[4] ), .ZN(new_n23747_));
  OAI21_X1   g23555(.A1(new_n23726_), .A2(new_n23747_), .B(new_n23732_), .ZN(new_n23748_));
  OAI21_X1   g23556(.A1(new_n23748_), .A2(new_n23724_), .B(new_n23746_), .ZN(new_n23749_));
  AOI21_X1   g23557(.A1(new_n23749_), .A2(\asqrt[4] ), .B(\asqrt[5] ), .ZN(new_n23750_));
  AOI21_X1   g23558(.A1(new_n23750_), .A2(new_n23741_), .B(new_n23745_), .ZN(new_n23751_));
  OAI21_X1   g23559(.A1(new_n23751_), .A2(new_n23742_), .B(\asqrt[6] ), .ZN(new_n23752_));
  INV_X1     g23560(.I(new_n23752_), .ZN(new_n23753_));
  NOR2_X1    g23561(.A1(new_n23005_), .A2(new_n23008_), .ZN(new_n23754_));
  INV_X1     g23562(.I(new_n23754_), .ZN(new_n23755_));
  NAND4_X1   g23563(.A1(\asqrt[2] ), .A2(new_n23006_), .A3(new_n22979_), .A4(new_n23755_), .ZN(new_n23756_));
  INV_X1     g23564(.I(\asqrt[2] ), .ZN(new_n23757_));
  NOR3_X1    g23565(.A1(new_n23757_), .A2(new_n22969_), .A3(new_n23754_), .ZN(new_n23758_));
  OAI21_X1   g23566(.A1(new_n23758_), .A2(new_n22979_), .B(new_n23756_), .ZN(new_n23759_));
  INV_X1     g23567(.I(new_n23759_), .ZN(new_n23760_));
  NOR3_X1    g23568(.A1(new_n23751_), .A2(new_n23742_), .A3(\asqrt[6] ), .ZN(new_n23761_));
  NOR2_X1    g23569(.A1(new_n23761_), .A2(new_n23760_), .ZN(new_n23762_));
  OAI21_X1   g23570(.A1(new_n23762_), .A2(new_n23753_), .B(\asqrt[7] ), .ZN(new_n23763_));
  NAND2_X1   g23571(.A1(new_n23014_), .A2(new_n23009_), .ZN(new_n23764_));
  NAND3_X1   g23572(.A1(\asqrt[2] ), .A2(new_n22982_), .A3(new_n23764_), .ZN(new_n23765_));
  AND3_X2    g23573(.A1(new_n22982_), .A2(new_n22986_), .A3(new_n23764_), .Z(new_n23766_));
  AOI22_X1   g23574(.A1(new_n23765_), .A2(new_n22987_), .B1(\asqrt[2] ), .B2(new_n23766_), .ZN(new_n23767_));
  INV_X1     g23575(.I(new_n23767_), .ZN(new_n23768_));
  NAND2_X1   g23576(.A1(new_n23752_), .A2(new_n20262_), .ZN(new_n23769_));
  OAI21_X1   g23577(.A1(new_n23762_), .A2(new_n23769_), .B(new_n23768_), .ZN(new_n23770_));
  AOI21_X1   g23578(.A1(new_n23770_), .A2(new_n23763_), .B(new_n19573_), .ZN(new_n23771_));
  NOR3_X1    g23579(.A1(new_n22990_), .A2(new_n22996_), .A3(new_n23016_), .ZN(new_n23772_));
  NOR3_X1    g23580(.A1(new_n23757_), .A2(new_n22990_), .A3(new_n23016_), .ZN(new_n23773_));
  INV_X1     g23581(.I(new_n23773_), .ZN(new_n23774_));
  AOI22_X1   g23582(.A1(new_n23774_), .A2(new_n22996_), .B1(\asqrt[2] ), .B2(new_n23772_), .ZN(new_n23775_));
  OAI21_X1   g23583(.A1(new_n23760_), .A2(new_n23761_), .B(new_n23752_), .ZN(new_n23776_));
  AOI21_X1   g23584(.A1(new_n23776_), .A2(\asqrt[7] ), .B(\asqrt[8] ), .ZN(new_n23777_));
  AOI21_X1   g23585(.A1(new_n23777_), .A2(new_n23770_), .B(new_n23775_), .ZN(new_n23778_));
  OAI21_X1   g23586(.A1(new_n23778_), .A2(new_n23771_), .B(\asqrt[9] ), .ZN(new_n23779_));
  INV_X1     g23587(.I(new_n23779_), .ZN(new_n23780_));
  NAND2_X1   g23588(.A1(new_n23516_), .A2(new_n23514_), .ZN(new_n23781_));
  NAND3_X1   g23589(.A1(\asqrt[2] ), .A2(new_n23018_), .A3(new_n23781_), .ZN(new_n23782_));
  AND3_X2    g23590(.A1(new_n23781_), .A2(new_n23018_), .A3(new_n23023_), .Z(new_n23783_));
  AOI22_X1   g23591(.A1(new_n23782_), .A2(new_n23024_), .B1(\asqrt[2] ), .B2(new_n23783_), .ZN(new_n23784_));
  NOR3_X1    g23592(.A1(new_n23778_), .A2(new_n23771_), .A3(\asqrt[9] ), .ZN(new_n23785_));
  NOR2_X1    g23593(.A1(new_n23785_), .A2(new_n23784_), .ZN(new_n23786_));
  OAI21_X1   g23594(.A1(new_n23786_), .A2(new_n23780_), .B(\asqrt[10] ), .ZN(new_n23787_));
  INV_X1     g23595(.I(new_n23032_), .ZN(new_n23788_));
  NOR3_X1    g23596(.A1(new_n23527_), .A2(new_n23028_), .A3(new_n23788_), .ZN(new_n23789_));
  NOR3_X1    g23597(.A1(new_n23757_), .A2(new_n23028_), .A3(new_n23527_), .ZN(new_n23790_));
  INV_X1     g23598(.I(new_n23790_), .ZN(new_n23791_));
  AOI22_X1   g23599(.A1(new_n23791_), .A2(new_n23788_), .B1(\asqrt[2] ), .B2(new_n23789_), .ZN(new_n23792_));
  INV_X1     g23600(.I(new_n23792_), .ZN(new_n23793_));
  NAND2_X1   g23601(.A1(new_n23779_), .A2(new_n18275_), .ZN(new_n23794_));
  OAI21_X1   g23602(.A1(new_n23786_), .A2(new_n23794_), .B(new_n23793_), .ZN(new_n23795_));
  AOI21_X1   g23603(.A1(new_n23795_), .A2(new_n23787_), .B(new_n17623_), .ZN(new_n23796_));
  NOR3_X1    g23604(.A1(new_n23757_), .A2(new_n23037_), .A3(new_n23042_), .ZN(new_n23797_));
  INV_X1     g23605(.I(new_n23797_), .ZN(new_n23798_));
  NOR3_X1    g23606(.A1(new_n23037_), .A2(new_n23512_), .A3(new_n23042_), .ZN(new_n23799_));
  AOI22_X1   g23607(.A1(new_n23798_), .A2(new_n23512_), .B1(\asqrt[2] ), .B2(new_n23799_), .ZN(new_n23800_));
  OAI21_X1   g23608(.A1(new_n23784_), .A2(new_n23785_), .B(new_n23779_), .ZN(new_n23801_));
  AOI21_X1   g23609(.A1(new_n23801_), .A2(\asqrt[10] ), .B(\asqrt[11] ), .ZN(new_n23802_));
  AOI21_X1   g23610(.A1(new_n23802_), .A2(new_n23795_), .B(new_n23800_), .ZN(new_n23803_));
  OAI21_X1   g23611(.A1(new_n23803_), .A2(new_n23796_), .B(\asqrt[12] ), .ZN(new_n23804_));
  INV_X1     g23612(.I(new_n23804_), .ZN(new_n23805_));
  AND3_X2    g23613(.A1(new_n23044_), .A2(new_n23049_), .A3(new_n23521_), .Z(new_n23806_));
  NAND3_X1   g23614(.A1(\asqrt[2] ), .A2(new_n23044_), .A3(new_n23521_), .ZN(new_n23807_));
  AOI22_X1   g23615(.A1(new_n23807_), .A2(new_n23050_), .B1(\asqrt[2] ), .B2(new_n23806_), .ZN(new_n23808_));
  NOR3_X1    g23616(.A1(new_n23803_), .A2(new_n23796_), .A3(\asqrt[12] ), .ZN(new_n23809_));
  NOR2_X1    g23617(.A1(new_n23809_), .A2(new_n23808_), .ZN(new_n23810_));
  OAI21_X1   g23618(.A1(new_n23810_), .A2(new_n23805_), .B(\asqrt[13] ), .ZN(new_n23811_));
  INV_X1     g23619(.I(new_n23057_), .ZN(new_n23812_));
  NOR3_X1    g23620(.A1(new_n23757_), .A2(new_n23053_), .A3(new_n23531_), .ZN(new_n23813_));
  INV_X1     g23621(.I(new_n23813_), .ZN(new_n23814_));
  NOR3_X1    g23622(.A1(new_n23531_), .A2(new_n23053_), .A3(new_n23812_), .ZN(new_n23815_));
  AOI22_X1   g23623(.A1(new_n23814_), .A2(new_n23812_), .B1(\asqrt[2] ), .B2(new_n23815_), .ZN(new_n23816_));
  INV_X1     g23624(.I(new_n23816_), .ZN(new_n23817_));
  NAND2_X1   g23625(.A1(new_n23804_), .A2(new_n16389_), .ZN(new_n23818_));
  OAI21_X1   g23626(.A1(new_n23810_), .A2(new_n23818_), .B(new_n23817_), .ZN(new_n23819_));
  AOI21_X1   g23627(.A1(new_n23819_), .A2(new_n23811_), .B(new_n15770_), .ZN(new_n23820_));
  NOR3_X1    g23628(.A1(new_n23062_), .A2(new_n23511_), .A3(new_n23067_), .ZN(new_n23821_));
  NOR3_X1    g23629(.A1(new_n23757_), .A2(new_n23062_), .A3(new_n23067_), .ZN(new_n23822_));
  INV_X1     g23630(.I(new_n23822_), .ZN(new_n23823_));
  AOI22_X1   g23631(.A1(new_n23823_), .A2(new_n23511_), .B1(\asqrt[2] ), .B2(new_n23821_), .ZN(new_n23824_));
  OAI21_X1   g23632(.A1(new_n23808_), .A2(new_n23809_), .B(new_n23804_), .ZN(new_n23825_));
  AOI21_X1   g23633(.A1(new_n23825_), .A2(\asqrt[13] ), .B(\asqrt[14] ), .ZN(new_n23826_));
  AOI21_X1   g23634(.A1(new_n23826_), .A2(new_n23819_), .B(new_n23824_), .ZN(new_n23827_));
  OAI21_X1   g23635(.A1(new_n23827_), .A2(new_n23820_), .B(\asqrt[15] ), .ZN(new_n23828_));
  INV_X1     g23636(.I(new_n23828_), .ZN(new_n23829_));
  NOR2_X1    g23637(.A1(new_n23068_), .A2(new_n23076_), .ZN(new_n23830_));
  NOR3_X1    g23638(.A1(new_n23757_), .A2(new_n23525_), .A3(new_n23830_), .ZN(new_n23831_));
  INV_X1     g23639(.I(new_n23831_), .ZN(new_n23832_));
  NOR3_X1    g23640(.A1(new_n23830_), .A2(new_n23525_), .A3(new_n23075_), .ZN(new_n23833_));
  AOI22_X1   g23641(.A1(new_n23832_), .A2(new_n23075_), .B1(\asqrt[2] ), .B2(new_n23833_), .ZN(new_n23834_));
  NOR3_X1    g23642(.A1(new_n23827_), .A2(new_n23820_), .A3(\asqrt[15] ), .ZN(new_n23835_));
  NOR2_X1    g23643(.A1(new_n23835_), .A2(new_n23834_), .ZN(new_n23836_));
  OAI21_X1   g23644(.A1(new_n23836_), .A2(new_n23829_), .B(\asqrt[16] ), .ZN(new_n23837_));
  INV_X1     g23645(.I(new_n23084_), .ZN(new_n23838_));
  NOR3_X1    g23646(.A1(new_n23539_), .A2(new_n23078_), .A3(new_n23838_), .ZN(new_n23839_));
  NOR3_X1    g23647(.A1(new_n23757_), .A2(new_n23078_), .A3(new_n23539_), .ZN(new_n23840_));
  INV_X1     g23648(.I(new_n23840_), .ZN(new_n23841_));
  AOI22_X1   g23649(.A1(new_n23841_), .A2(new_n23838_), .B1(\asqrt[2] ), .B2(new_n23839_), .ZN(new_n23842_));
  INV_X1     g23650(.I(new_n23842_), .ZN(new_n23843_));
  NAND2_X1   g23651(.A1(new_n23828_), .A2(new_n14601_), .ZN(new_n23844_));
  OAI21_X1   g23652(.A1(new_n23836_), .A2(new_n23844_), .B(new_n23843_), .ZN(new_n23845_));
  AOI21_X1   g23653(.A1(new_n23845_), .A2(new_n23837_), .B(new_n14017_), .ZN(new_n23846_));
  NOR3_X1    g23654(.A1(new_n23757_), .A2(new_n23089_), .A3(new_n23098_), .ZN(new_n23847_));
  INV_X1     g23655(.I(new_n23847_), .ZN(new_n23848_));
  NOR3_X1    g23656(.A1(new_n23089_), .A2(new_n23510_), .A3(new_n23098_), .ZN(new_n23849_));
  AOI22_X1   g23657(.A1(new_n23848_), .A2(new_n23510_), .B1(\asqrt[2] ), .B2(new_n23849_), .ZN(new_n23850_));
  OAI21_X1   g23658(.A1(new_n23834_), .A2(new_n23835_), .B(new_n23828_), .ZN(new_n23851_));
  AOI21_X1   g23659(.A1(new_n23851_), .A2(\asqrt[16] ), .B(\asqrt[17] ), .ZN(new_n23852_));
  AOI21_X1   g23660(.A1(new_n23852_), .A2(new_n23845_), .B(new_n23850_), .ZN(new_n23853_));
  OAI21_X1   g23661(.A1(new_n23853_), .A2(new_n23846_), .B(\asqrt[18] ), .ZN(new_n23854_));
  INV_X1     g23662(.I(new_n23854_), .ZN(new_n23855_));
  NOR2_X1    g23663(.A1(new_n23099_), .A2(new_n23107_), .ZN(new_n23856_));
  NOR3_X1    g23664(.A1(new_n23856_), .A2(new_n23538_), .A3(new_n23106_), .ZN(new_n23857_));
  NOR3_X1    g23665(.A1(new_n23757_), .A2(new_n23538_), .A3(new_n23856_), .ZN(new_n23858_));
  INV_X1     g23666(.I(new_n23858_), .ZN(new_n23859_));
  AOI22_X1   g23667(.A1(new_n23859_), .A2(new_n23106_), .B1(\asqrt[2] ), .B2(new_n23857_), .ZN(new_n23860_));
  NOR3_X1    g23668(.A1(new_n23853_), .A2(new_n23846_), .A3(\asqrt[18] ), .ZN(new_n23861_));
  NOR2_X1    g23669(.A1(new_n23861_), .A2(new_n23860_), .ZN(new_n23862_));
  OAI21_X1   g23670(.A1(new_n23862_), .A2(new_n23855_), .B(\asqrt[19] ), .ZN(new_n23863_));
  INV_X1     g23671(.I(new_n23114_), .ZN(new_n23864_));
  NOR3_X1    g23672(.A1(new_n23757_), .A2(new_n23109_), .A3(new_n23547_), .ZN(new_n23865_));
  INV_X1     g23673(.I(new_n23865_), .ZN(new_n23866_));
  NOR3_X1    g23674(.A1(new_n23547_), .A2(new_n23109_), .A3(new_n23864_), .ZN(new_n23867_));
  AOI22_X1   g23675(.A1(new_n23866_), .A2(new_n23864_), .B1(\asqrt[2] ), .B2(new_n23867_), .ZN(new_n23868_));
  INV_X1     g23676(.I(new_n23868_), .ZN(new_n23869_));
  NAND2_X1   g23677(.A1(new_n23854_), .A2(new_n12913_), .ZN(new_n23870_));
  OAI21_X1   g23678(.A1(new_n23862_), .A2(new_n23870_), .B(new_n23869_), .ZN(new_n23871_));
  AOI21_X1   g23679(.A1(new_n23871_), .A2(new_n23863_), .B(new_n12364_), .ZN(new_n23872_));
  NOR3_X1    g23680(.A1(new_n23119_), .A2(new_n23509_), .A3(new_n23128_), .ZN(new_n23873_));
  NOR3_X1    g23681(.A1(new_n23757_), .A2(new_n23119_), .A3(new_n23128_), .ZN(new_n23874_));
  INV_X1     g23682(.I(new_n23874_), .ZN(new_n23875_));
  AOI22_X1   g23683(.A1(new_n23875_), .A2(new_n23509_), .B1(\asqrt[2] ), .B2(new_n23873_), .ZN(new_n23876_));
  OAI21_X1   g23684(.A1(new_n23860_), .A2(new_n23861_), .B(new_n23854_), .ZN(new_n23877_));
  AOI21_X1   g23685(.A1(new_n23877_), .A2(\asqrt[19] ), .B(\asqrt[20] ), .ZN(new_n23878_));
  AOI21_X1   g23686(.A1(new_n23878_), .A2(new_n23871_), .B(new_n23876_), .ZN(new_n23879_));
  OAI21_X1   g23687(.A1(new_n23879_), .A2(new_n23872_), .B(\asqrt[21] ), .ZN(new_n23880_));
  INV_X1     g23688(.I(new_n23880_), .ZN(new_n23881_));
  NOR2_X1    g23689(.A1(new_n23129_), .A2(new_n23137_), .ZN(new_n23882_));
  NOR3_X1    g23690(.A1(new_n23757_), .A2(new_n23546_), .A3(new_n23882_), .ZN(new_n23883_));
  INV_X1     g23691(.I(new_n23883_), .ZN(new_n23884_));
  NOR3_X1    g23692(.A1(new_n23882_), .A2(new_n23546_), .A3(new_n23136_), .ZN(new_n23885_));
  AOI22_X1   g23693(.A1(new_n23884_), .A2(new_n23136_), .B1(\asqrt[2] ), .B2(new_n23885_), .ZN(new_n23886_));
  NOR3_X1    g23694(.A1(new_n23879_), .A2(new_n23872_), .A3(\asqrt[21] ), .ZN(new_n23887_));
  NOR2_X1    g23695(.A1(new_n23887_), .A2(new_n23886_), .ZN(new_n23888_));
  OAI21_X1   g23696(.A1(new_n23888_), .A2(new_n23881_), .B(\asqrt[22] ), .ZN(new_n23889_));
  INV_X1     g23697(.I(new_n23144_), .ZN(new_n23890_));
  NOR3_X1    g23698(.A1(new_n23555_), .A2(new_n23139_), .A3(new_n23890_), .ZN(new_n23891_));
  NOR3_X1    g23699(.A1(new_n23757_), .A2(new_n23139_), .A3(new_n23555_), .ZN(new_n23892_));
  INV_X1     g23700(.I(new_n23892_), .ZN(new_n23893_));
  AOI22_X1   g23701(.A1(new_n23893_), .A2(new_n23890_), .B1(\asqrt[2] ), .B2(new_n23891_), .ZN(new_n23894_));
  INV_X1     g23702(.I(new_n23894_), .ZN(new_n23895_));
  NAND2_X1   g23703(.A1(new_n23880_), .A2(new_n11326_), .ZN(new_n23896_));
  OAI21_X1   g23704(.A1(new_n23888_), .A2(new_n23896_), .B(new_n23895_), .ZN(new_n23897_));
  AOI21_X1   g23705(.A1(new_n23897_), .A2(new_n23889_), .B(new_n10812_), .ZN(new_n23898_));
  NOR3_X1    g23706(.A1(new_n23757_), .A2(new_n23149_), .A3(new_n23158_), .ZN(new_n23899_));
  INV_X1     g23707(.I(new_n23899_), .ZN(new_n23900_));
  NOR3_X1    g23708(.A1(new_n23149_), .A2(new_n23508_), .A3(new_n23158_), .ZN(new_n23901_));
  AOI22_X1   g23709(.A1(new_n23900_), .A2(new_n23508_), .B1(\asqrt[2] ), .B2(new_n23901_), .ZN(new_n23902_));
  OAI21_X1   g23710(.A1(new_n23886_), .A2(new_n23887_), .B(new_n23880_), .ZN(new_n23903_));
  AOI21_X1   g23711(.A1(new_n23903_), .A2(\asqrt[22] ), .B(\asqrt[23] ), .ZN(new_n23904_));
  AOI21_X1   g23712(.A1(new_n23904_), .A2(new_n23897_), .B(new_n23902_), .ZN(new_n23905_));
  OAI21_X1   g23713(.A1(new_n23905_), .A2(new_n23898_), .B(\asqrt[24] ), .ZN(new_n23906_));
  INV_X1     g23714(.I(new_n23906_), .ZN(new_n23907_));
  NOR2_X1    g23715(.A1(new_n23159_), .A2(new_n23167_), .ZN(new_n23908_));
  NOR3_X1    g23716(.A1(new_n23908_), .A2(new_n23554_), .A3(new_n23166_), .ZN(new_n23909_));
  NOR3_X1    g23717(.A1(new_n23757_), .A2(new_n23554_), .A3(new_n23908_), .ZN(new_n23910_));
  INV_X1     g23718(.I(new_n23910_), .ZN(new_n23911_));
  AOI22_X1   g23719(.A1(new_n23911_), .A2(new_n23166_), .B1(\asqrt[2] ), .B2(new_n23909_), .ZN(new_n23912_));
  NOR3_X1    g23720(.A1(new_n23905_), .A2(new_n23898_), .A3(\asqrt[24] ), .ZN(new_n23913_));
  NOR2_X1    g23721(.A1(new_n23913_), .A2(new_n23912_), .ZN(new_n23914_));
  OAI21_X1   g23722(.A1(new_n23914_), .A2(new_n23907_), .B(\asqrt[25] ), .ZN(new_n23915_));
  INV_X1     g23723(.I(new_n23174_), .ZN(new_n23916_));
  NOR3_X1    g23724(.A1(new_n23757_), .A2(new_n23169_), .A3(new_n23563_), .ZN(new_n23917_));
  INV_X1     g23725(.I(new_n23917_), .ZN(new_n23918_));
  NOR3_X1    g23726(.A1(new_n23563_), .A2(new_n23169_), .A3(new_n23916_), .ZN(new_n23919_));
  AOI22_X1   g23727(.A1(new_n23918_), .A2(new_n23916_), .B1(\asqrt[2] ), .B2(new_n23919_), .ZN(new_n23920_));
  INV_X1     g23728(.I(new_n23920_), .ZN(new_n23921_));
  NAND2_X1   g23729(.A1(new_n23906_), .A2(new_n9846_), .ZN(new_n23922_));
  OAI21_X1   g23730(.A1(new_n23914_), .A2(new_n23922_), .B(new_n23921_), .ZN(new_n23923_));
  AOI21_X1   g23731(.A1(new_n23923_), .A2(new_n23915_), .B(new_n9317_), .ZN(new_n23924_));
  NOR3_X1    g23732(.A1(new_n23179_), .A2(new_n23507_), .A3(new_n23188_), .ZN(new_n23925_));
  NOR3_X1    g23733(.A1(new_n23757_), .A2(new_n23179_), .A3(new_n23188_), .ZN(new_n23926_));
  INV_X1     g23734(.I(new_n23926_), .ZN(new_n23927_));
  AOI22_X1   g23735(.A1(new_n23927_), .A2(new_n23507_), .B1(\asqrt[2] ), .B2(new_n23925_), .ZN(new_n23928_));
  OAI21_X1   g23736(.A1(new_n23912_), .A2(new_n23913_), .B(new_n23906_), .ZN(new_n23929_));
  AOI21_X1   g23737(.A1(new_n23929_), .A2(\asqrt[25] ), .B(\asqrt[26] ), .ZN(new_n23930_));
  AOI21_X1   g23738(.A1(new_n23930_), .A2(new_n23923_), .B(new_n23928_), .ZN(new_n23931_));
  OAI21_X1   g23739(.A1(new_n23931_), .A2(new_n23924_), .B(\asqrt[27] ), .ZN(new_n23932_));
  INV_X1     g23740(.I(new_n23932_), .ZN(new_n23933_));
  NOR2_X1    g23741(.A1(new_n23189_), .A2(new_n23197_), .ZN(new_n23934_));
  NOR3_X1    g23742(.A1(new_n23757_), .A2(new_n23562_), .A3(new_n23934_), .ZN(new_n23935_));
  INV_X1     g23743(.I(new_n23935_), .ZN(new_n23936_));
  NOR3_X1    g23744(.A1(new_n23934_), .A2(new_n23562_), .A3(new_n23196_), .ZN(new_n23937_));
  AOI22_X1   g23745(.A1(new_n23936_), .A2(new_n23196_), .B1(\asqrt[2] ), .B2(new_n23937_), .ZN(new_n23938_));
  NOR3_X1    g23746(.A1(new_n23931_), .A2(new_n23924_), .A3(\asqrt[27] ), .ZN(new_n23939_));
  NOR2_X1    g23747(.A1(new_n23939_), .A2(new_n23938_), .ZN(new_n23940_));
  OAI21_X1   g23748(.A1(new_n23940_), .A2(new_n23933_), .B(\asqrt[28] ), .ZN(new_n23941_));
  INV_X1     g23749(.I(new_n23204_), .ZN(new_n23942_));
  NOR3_X1    g23750(.A1(new_n23571_), .A2(new_n23199_), .A3(new_n23942_), .ZN(new_n23943_));
  NOR3_X1    g23751(.A1(new_n23757_), .A2(new_n23199_), .A3(new_n23571_), .ZN(new_n23944_));
  INV_X1     g23752(.I(new_n23944_), .ZN(new_n23945_));
  AOI22_X1   g23753(.A1(new_n23945_), .A2(new_n23942_), .B1(\asqrt[2] ), .B2(new_n23943_), .ZN(new_n23946_));
  INV_X1     g23754(.I(new_n23946_), .ZN(new_n23947_));
  NAND2_X1   g23755(.A1(new_n23932_), .A2(new_n8483_), .ZN(new_n23948_));
  OAI21_X1   g23756(.A1(new_n23940_), .A2(new_n23948_), .B(new_n23947_), .ZN(new_n23949_));
  AOI21_X1   g23757(.A1(new_n23949_), .A2(new_n23941_), .B(new_n8036_), .ZN(new_n23950_));
  NOR3_X1    g23758(.A1(new_n23757_), .A2(new_n23209_), .A3(new_n23218_), .ZN(new_n23951_));
  INV_X1     g23759(.I(new_n23951_), .ZN(new_n23952_));
  NOR3_X1    g23760(.A1(new_n23209_), .A2(new_n23506_), .A3(new_n23218_), .ZN(new_n23953_));
  AOI22_X1   g23761(.A1(new_n23952_), .A2(new_n23506_), .B1(\asqrt[2] ), .B2(new_n23953_), .ZN(new_n23954_));
  OAI21_X1   g23762(.A1(new_n23938_), .A2(new_n23939_), .B(new_n23932_), .ZN(new_n23955_));
  AOI21_X1   g23763(.A1(new_n23955_), .A2(\asqrt[28] ), .B(\asqrt[29] ), .ZN(new_n23956_));
  AOI21_X1   g23764(.A1(new_n23956_), .A2(new_n23949_), .B(new_n23954_), .ZN(new_n23957_));
  OAI21_X1   g23765(.A1(new_n23957_), .A2(new_n23950_), .B(\asqrt[30] ), .ZN(new_n23958_));
  INV_X1     g23766(.I(new_n23958_), .ZN(new_n23959_));
  NOR2_X1    g23767(.A1(new_n23219_), .A2(new_n23227_), .ZN(new_n23960_));
  NOR3_X1    g23768(.A1(new_n23960_), .A2(new_n23570_), .A3(new_n23226_), .ZN(new_n23961_));
  NOR3_X1    g23769(.A1(new_n23757_), .A2(new_n23570_), .A3(new_n23960_), .ZN(new_n23962_));
  INV_X1     g23770(.I(new_n23962_), .ZN(new_n23963_));
  AOI22_X1   g23771(.A1(new_n23963_), .A2(new_n23226_), .B1(\asqrt[2] ), .B2(new_n23961_), .ZN(new_n23964_));
  NOR3_X1    g23772(.A1(new_n23957_), .A2(new_n23950_), .A3(\asqrt[30] ), .ZN(new_n23965_));
  NOR2_X1    g23773(.A1(new_n23965_), .A2(new_n23964_), .ZN(new_n23966_));
  OAI21_X1   g23774(.A1(new_n23966_), .A2(new_n23959_), .B(\asqrt[31] ), .ZN(new_n23967_));
  INV_X1     g23775(.I(new_n23234_), .ZN(new_n23968_));
  NOR3_X1    g23776(.A1(new_n23757_), .A2(new_n23229_), .A3(new_n23579_), .ZN(new_n23969_));
  INV_X1     g23777(.I(new_n23969_), .ZN(new_n23970_));
  NOR3_X1    g23778(.A1(new_n23579_), .A2(new_n23229_), .A3(new_n23968_), .ZN(new_n23971_));
  AOI22_X1   g23779(.A1(new_n23970_), .A2(new_n23968_), .B1(\asqrt[2] ), .B2(new_n23971_), .ZN(new_n23972_));
  INV_X1     g23780(.I(new_n23972_), .ZN(new_n23973_));
  NAND2_X1   g23781(.A1(new_n23958_), .A2(new_n7229_), .ZN(new_n23974_));
  OAI21_X1   g23782(.A1(new_n23966_), .A2(new_n23974_), .B(new_n23973_), .ZN(new_n23975_));
  AOI21_X1   g23783(.A1(new_n23975_), .A2(new_n23967_), .B(new_n6824_), .ZN(new_n23976_));
  NOR3_X1    g23784(.A1(new_n23239_), .A2(new_n23505_), .A3(new_n23245_), .ZN(new_n23977_));
  NOR3_X1    g23785(.A1(new_n23757_), .A2(new_n23239_), .A3(new_n23245_), .ZN(new_n23978_));
  INV_X1     g23786(.I(new_n23978_), .ZN(new_n23979_));
  AOI22_X1   g23787(.A1(new_n23979_), .A2(new_n23505_), .B1(\asqrt[2] ), .B2(new_n23977_), .ZN(new_n23980_));
  OAI21_X1   g23788(.A1(new_n23964_), .A2(new_n23965_), .B(new_n23958_), .ZN(new_n23981_));
  AOI21_X1   g23789(.A1(new_n23981_), .A2(\asqrt[31] ), .B(\asqrt[32] ), .ZN(new_n23982_));
  AOI21_X1   g23790(.A1(new_n23982_), .A2(new_n23975_), .B(new_n23980_), .ZN(new_n23983_));
  OAI21_X1   g23791(.A1(new_n23983_), .A2(new_n23976_), .B(\asqrt[33] ), .ZN(new_n23984_));
  INV_X1     g23792(.I(new_n23984_), .ZN(new_n23985_));
  NOR2_X1    g23793(.A1(new_n23246_), .A2(new_n23254_), .ZN(new_n23986_));
  NOR3_X1    g23794(.A1(new_n23757_), .A2(new_n23578_), .A3(new_n23986_), .ZN(new_n23987_));
  INV_X1     g23795(.I(new_n23987_), .ZN(new_n23988_));
  NOR3_X1    g23796(.A1(new_n23986_), .A2(new_n23578_), .A3(new_n23253_), .ZN(new_n23989_));
  AOI22_X1   g23797(.A1(new_n23988_), .A2(new_n23253_), .B1(\asqrt[2] ), .B2(new_n23989_), .ZN(new_n23990_));
  NOR3_X1    g23798(.A1(new_n23983_), .A2(new_n23976_), .A3(\asqrt[33] ), .ZN(new_n23991_));
  NOR2_X1    g23799(.A1(new_n23991_), .A2(new_n23990_), .ZN(new_n23992_));
  OAI21_X1   g23800(.A1(new_n23992_), .A2(new_n23985_), .B(\asqrt[34] ), .ZN(new_n23993_));
  INV_X1     g23801(.I(new_n23261_), .ZN(new_n23994_));
  NOR3_X1    g23802(.A1(new_n23587_), .A2(new_n23256_), .A3(new_n23994_), .ZN(new_n23995_));
  NOR3_X1    g23803(.A1(new_n23757_), .A2(new_n23256_), .A3(new_n23587_), .ZN(new_n23996_));
  INV_X1     g23804(.I(new_n23996_), .ZN(new_n23997_));
  AOI22_X1   g23805(.A1(new_n23997_), .A2(new_n23994_), .B1(\asqrt[2] ), .B2(new_n23995_), .ZN(new_n23998_));
  INV_X1     g23806(.I(new_n23998_), .ZN(new_n23999_));
  NAND2_X1   g23807(.A1(new_n23984_), .A2(new_n6077_), .ZN(new_n24000_));
  OAI21_X1   g23808(.A1(new_n23992_), .A2(new_n24000_), .B(new_n23999_), .ZN(new_n24001_));
  AOI21_X1   g23809(.A1(new_n24001_), .A2(new_n23993_), .B(new_n5708_), .ZN(new_n24002_));
  NOR3_X1    g23810(.A1(new_n23757_), .A2(new_n23266_), .A3(new_n23272_), .ZN(new_n24003_));
  INV_X1     g23811(.I(new_n24003_), .ZN(new_n24004_));
  NOR3_X1    g23812(.A1(new_n23266_), .A2(new_n23504_), .A3(new_n23272_), .ZN(new_n24005_));
  AOI22_X1   g23813(.A1(new_n24004_), .A2(new_n23504_), .B1(\asqrt[2] ), .B2(new_n24005_), .ZN(new_n24006_));
  OAI21_X1   g23814(.A1(new_n23990_), .A2(new_n23991_), .B(new_n23984_), .ZN(new_n24007_));
  AOI21_X1   g23815(.A1(new_n24007_), .A2(\asqrt[34] ), .B(\asqrt[35] ), .ZN(new_n24008_));
  AOI21_X1   g23816(.A1(new_n24008_), .A2(new_n24001_), .B(new_n24006_), .ZN(new_n24009_));
  OAI21_X1   g23817(.A1(new_n24009_), .A2(new_n24002_), .B(\asqrt[36] ), .ZN(new_n24010_));
  INV_X1     g23818(.I(new_n24010_), .ZN(new_n24011_));
  NOR2_X1    g23819(.A1(new_n23273_), .A2(new_n23281_), .ZN(new_n24012_));
  NOR3_X1    g23820(.A1(new_n24012_), .A2(new_n23586_), .A3(new_n23280_), .ZN(new_n24013_));
  NOR3_X1    g23821(.A1(new_n23757_), .A2(new_n23586_), .A3(new_n24012_), .ZN(new_n24014_));
  INV_X1     g23822(.I(new_n24014_), .ZN(new_n24015_));
  AOI22_X1   g23823(.A1(new_n24015_), .A2(new_n23280_), .B1(\asqrt[2] ), .B2(new_n24013_), .ZN(new_n24016_));
  NOR3_X1    g23824(.A1(new_n24009_), .A2(new_n24002_), .A3(\asqrt[36] ), .ZN(new_n24017_));
  NOR2_X1    g23825(.A1(new_n24017_), .A2(new_n24016_), .ZN(new_n24018_));
  OAI21_X1   g23826(.A1(new_n24018_), .A2(new_n24011_), .B(\asqrt[37] ), .ZN(new_n24019_));
  INV_X1     g23827(.I(new_n23288_), .ZN(new_n24020_));
  NOR3_X1    g23828(.A1(new_n23757_), .A2(new_n23283_), .A3(new_n23595_), .ZN(new_n24021_));
  INV_X1     g23829(.I(new_n24021_), .ZN(new_n24022_));
  NOR3_X1    g23830(.A1(new_n23595_), .A2(new_n23283_), .A3(new_n24020_), .ZN(new_n24023_));
  AOI22_X1   g23831(.A1(new_n24022_), .A2(new_n24020_), .B1(\asqrt[2] ), .B2(new_n24023_), .ZN(new_n24024_));
  INV_X1     g23832(.I(new_n24024_), .ZN(new_n24025_));
  NAND2_X1   g23833(.A1(new_n24010_), .A2(new_n5024_), .ZN(new_n24026_));
  OAI21_X1   g23834(.A1(new_n24018_), .A2(new_n24026_), .B(new_n24025_), .ZN(new_n24027_));
  AOI21_X1   g23835(.A1(new_n24027_), .A2(new_n24019_), .B(new_n4696_), .ZN(new_n24028_));
  NOR3_X1    g23836(.A1(new_n23293_), .A2(new_n23503_), .A3(new_n23299_), .ZN(new_n24029_));
  NOR3_X1    g23837(.A1(new_n23757_), .A2(new_n23293_), .A3(new_n23299_), .ZN(new_n24030_));
  INV_X1     g23838(.I(new_n24030_), .ZN(new_n24031_));
  AOI22_X1   g23839(.A1(new_n24031_), .A2(new_n23503_), .B1(\asqrt[2] ), .B2(new_n24029_), .ZN(new_n24032_));
  OAI21_X1   g23840(.A1(new_n24016_), .A2(new_n24017_), .B(new_n24010_), .ZN(new_n24033_));
  AOI21_X1   g23841(.A1(new_n24033_), .A2(\asqrt[37] ), .B(\asqrt[38] ), .ZN(new_n24034_));
  AOI21_X1   g23842(.A1(new_n24034_), .A2(new_n24027_), .B(new_n24032_), .ZN(new_n24035_));
  OAI21_X1   g23843(.A1(new_n24035_), .A2(new_n24028_), .B(\asqrt[39] ), .ZN(new_n24036_));
  INV_X1     g23844(.I(new_n24036_), .ZN(new_n24037_));
  NOR2_X1    g23845(.A1(new_n23300_), .A2(new_n23308_), .ZN(new_n24038_));
  NOR3_X1    g23846(.A1(new_n23757_), .A2(new_n23594_), .A3(new_n24038_), .ZN(new_n24039_));
  INV_X1     g23847(.I(new_n24039_), .ZN(new_n24040_));
  NOR3_X1    g23848(.A1(new_n24038_), .A2(new_n23594_), .A3(new_n23307_), .ZN(new_n24041_));
  AOI22_X1   g23849(.A1(new_n24040_), .A2(new_n23307_), .B1(\asqrt[2] ), .B2(new_n24041_), .ZN(new_n24042_));
  NOR3_X1    g23850(.A1(new_n24035_), .A2(new_n24028_), .A3(\asqrt[39] ), .ZN(new_n24043_));
  NOR2_X1    g23851(.A1(new_n24043_), .A2(new_n24042_), .ZN(new_n24044_));
  OAI21_X1   g23852(.A1(new_n24044_), .A2(new_n24037_), .B(\asqrt[40] ), .ZN(new_n24045_));
  INV_X1     g23853(.I(new_n23314_), .ZN(new_n24046_));
  NOR3_X1    g23854(.A1(new_n23603_), .A2(new_n23310_), .A3(new_n24046_), .ZN(new_n24047_));
  NOR3_X1    g23855(.A1(new_n23757_), .A2(new_n23310_), .A3(new_n23603_), .ZN(new_n24048_));
  INV_X1     g23856(.I(new_n24048_), .ZN(new_n24049_));
  AOI22_X1   g23857(.A1(new_n24049_), .A2(new_n24046_), .B1(\asqrt[2] ), .B2(new_n24047_), .ZN(new_n24050_));
  INV_X1     g23858(.I(new_n24050_), .ZN(new_n24051_));
  NAND2_X1   g23859(.A1(new_n24036_), .A2(new_n4071_), .ZN(new_n24052_));
  OAI21_X1   g23860(.A1(new_n24044_), .A2(new_n24052_), .B(new_n24051_), .ZN(new_n24053_));
  AOI21_X1   g23861(.A1(new_n24053_), .A2(new_n24045_), .B(new_n3782_), .ZN(new_n24054_));
  NOR3_X1    g23862(.A1(new_n23757_), .A2(new_n23319_), .A3(new_n23325_), .ZN(new_n24055_));
  INV_X1     g23863(.I(new_n24055_), .ZN(new_n24056_));
  NOR3_X1    g23864(.A1(new_n23319_), .A2(new_n23502_), .A3(new_n23325_), .ZN(new_n24057_));
  AOI22_X1   g23865(.A1(new_n24056_), .A2(new_n23502_), .B1(\asqrt[2] ), .B2(new_n24057_), .ZN(new_n24058_));
  OAI21_X1   g23866(.A1(new_n24042_), .A2(new_n24043_), .B(new_n24036_), .ZN(new_n24059_));
  AOI21_X1   g23867(.A1(new_n24059_), .A2(\asqrt[40] ), .B(\asqrt[41] ), .ZN(new_n24060_));
  AOI21_X1   g23868(.A1(new_n24060_), .A2(new_n24053_), .B(new_n24058_), .ZN(new_n24061_));
  OAI21_X1   g23869(.A1(new_n24061_), .A2(new_n24054_), .B(\asqrt[42] ), .ZN(new_n24062_));
  INV_X1     g23870(.I(new_n24062_), .ZN(new_n24063_));
  NOR2_X1    g23871(.A1(new_n23326_), .A2(new_n23334_), .ZN(new_n24064_));
  NOR3_X1    g23872(.A1(new_n24064_), .A2(new_n23602_), .A3(new_n23333_), .ZN(new_n24065_));
  NOR3_X1    g23873(.A1(new_n23757_), .A2(new_n23602_), .A3(new_n24064_), .ZN(new_n24066_));
  INV_X1     g23874(.I(new_n24066_), .ZN(new_n24067_));
  AOI22_X1   g23875(.A1(new_n24067_), .A2(new_n23333_), .B1(\asqrt[2] ), .B2(new_n24065_), .ZN(new_n24068_));
  NOR3_X1    g23876(.A1(new_n24061_), .A2(new_n24054_), .A3(\asqrt[42] ), .ZN(new_n24069_));
  NOR2_X1    g23877(.A1(new_n24069_), .A2(new_n24068_), .ZN(new_n24070_));
  OAI21_X1   g23878(.A1(new_n24070_), .A2(new_n24063_), .B(\asqrt[43] ), .ZN(new_n24071_));
  INV_X1     g23879(.I(new_n23340_), .ZN(new_n24072_));
  NOR3_X1    g23880(.A1(new_n23757_), .A2(new_n23336_), .A3(new_n23611_), .ZN(new_n24073_));
  INV_X1     g23881(.I(new_n24073_), .ZN(new_n24074_));
  NOR3_X1    g23882(.A1(new_n23611_), .A2(new_n23336_), .A3(new_n24072_), .ZN(new_n24075_));
  AOI22_X1   g23883(.A1(new_n24074_), .A2(new_n24072_), .B1(\asqrt[2] ), .B2(new_n24075_), .ZN(new_n24076_));
  INV_X1     g23884(.I(new_n24076_), .ZN(new_n24077_));
  NAND2_X1   g23885(.A1(new_n24062_), .A2(new_n3218_), .ZN(new_n24078_));
  OAI21_X1   g23886(.A1(new_n24070_), .A2(new_n24078_), .B(new_n24077_), .ZN(new_n24079_));
  AOI21_X1   g23887(.A1(new_n24079_), .A2(new_n24071_), .B(new_n2954_), .ZN(new_n24080_));
  NOR3_X1    g23888(.A1(new_n23345_), .A2(new_n23501_), .A3(new_n23353_), .ZN(new_n24081_));
  NOR3_X1    g23889(.A1(new_n23757_), .A2(new_n23345_), .A3(new_n23353_), .ZN(new_n24082_));
  INV_X1     g23890(.I(new_n24082_), .ZN(new_n24083_));
  AOI22_X1   g23891(.A1(new_n24083_), .A2(new_n23501_), .B1(\asqrt[2] ), .B2(new_n24081_), .ZN(new_n24084_));
  OAI21_X1   g23892(.A1(new_n24068_), .A2(new_n24069_), .B(new_n24062_), .ZN(new_n24085_));
  AOI21_X1   g23893(.A1(new_n24085_), .A2(\asqrt[43] ), .B(\asqrt[44] ), .ZN(new_n24086_));
  AOI21_X1   g23894(.A1(new_n24086_), .A2(new_n24079_), .B(new_n24084_), .ZN(new_n24087_));
  OAI21_X1   g23895(.A1(new_n24087_), .A2(new_n24080_), .B(\asqrt[45] ), .ZN(new_n24088_));
  INV_X1     g23896(.I(new_n24088_), .ZN(new_n24089_));
  NOR2_X1    g23897(.A1(new_n23354_), .A2(new_n23361_), .ZN(new_n24090_));
  NOR3_X1    g23898(.A1(new_n23757_), .A2(new_n23610_), .A3(new_n24090_), .ZN(new_n24091_));
  INV_X1     g23899(.I(new_n24091_), .ZN(new_n24092_));
  NOR3_X1    g23900(.A1(new_n24090_), .A2(new_n23610_), .A3(new_n23360_), .ZN(new_n24093_));
  AOI22_X1   g23901(.A1(new_n24092_), .A2(new_n23360_), .B1(\asqrt[2] ), .B2(new_n24093_), .ZN(new_n24094_));
  NOR3_X1    g23902(.A1(new_n24087_), .A2(new_n24080_), .A3(\asqrt[45] ), .ZN(new_n24095_));
  NOR2_X1    g23903(.A1(new_n24095_), .A2(new_n24094_), .ZN(new_n24096_));
  OAI21_X1   g23904(.A1(new_n24096_), .A2(new_n24089_), .B(\asqrt[46] ), .ZN(new_n24097_));
  INV_X1     g23905(.I(new_n23369_), .ZN(new_n24098_));
  NOR3_X1    g23906(.A1(new_n23619_), .A2(new_n23363_), .A3(new_n24098_), .ZN(new_n24099_));
  NOR3_X1    g23907(.A1(new_n23757_), .A2(new_n23363_), .A3(new_n23619_), .ZN(new_n24100_));
  INV_X1     g23908(.I(new_n24100_), .ZN(new_n24101_));
  AOI22_X1   g23909(.A1(new_n24101_), .A2(new_n24098_), .B1(\asqrt[2] ), .B2(new_n24099_), .ZN(new_n24102_));
  INV_X1     g23910(.I(new_n24102_), .ZN(new_n24103_));
  NAND2_X1   g23911(.A1(new_n24088_), .A2(new_n2465_), .ZN(new_n24104_));
  OAI21_X1   g23912(.A1(new_n24096_), .A2(new_n24104_), .B(new_n24103_), .ZN(new_n24105_));
  AOI21_X1   g23913(.A1(new_n24105_), .A2(new_n24097_), .B(new_n2229_), .ZN(new_n24106_));
  NOR3_X1    g23914(.A1(new_n23757_), .A2(new_n23374_), .A3(new_n23383_), .ZN(new_n24107_));
  INV_X1     g23915(.I(new_n24107_), .ZN(new_n24108_));
  NOR3_X1    g23916(.A1(new_n23374_), .A2(new_n23500_), .A3(new_n23383_), .ZN(new_n24109_));
  AOI22_X1   g23917(.A1(new_n24108_), .A2(new_n23500_), .B1(\asqrt[2] ), .B2(new_n24109_), .ZN(new_n24110_));
  OAI21_X1   g23918(.A1(new_n24094_), .A2(new_n24095_), .B(new_n24088_), .ZN(new_n24111_));
  AOI21_X1   g23919(.A1(new_n24111_), .A2(\asqrt[46] ), .B(\asqrt[47] ), .ZN(new_n24112_));
  AOI21_X1   g23920(.A1(new_n24112_), .A2(new_n24105_), .B(new_n24110_), .ZN(new_n24113_));
  OAI21_X1   g23921(.A1(new_n24113_), .A2(new_n24106_), .B(\asqrt[48] ), .ZN(new_n24114_));
  INV_X1     g23922(.I(new_n24114_), .ZN(new_n24115_));
  NOR2_X1    g23923(.A1(new_n23384_), .A2(new_n23391_), .ZN(new_n24116_));
  NOR3_X1    g23924(.A1(new_n24116_), .A2(new_n23618_), .A3(new_n23390_), .ZN(new_n24117_));
  NOR3_X1    g23925(.A1(new_n23757_), .A2(new_n23618_), .A3(new_n24116_), .ZN(new_n24118_));
  INV_X1     g23926(.I(new_n24118_), .ZN(new_n24119_));
  AOI22_X1   g23927(.A1(new_n24119_), .A2(new_n23390_), .B1(\asqrt[2] ), .B2(new_n24117_), .ZN(new_n24120_));
  NOR3_X1    g23928(.A1(new_n24113_), .A2(new_n24106_), .A3(\asqrt[48] ), .ZN(new_n24121_));
  NOR2_X1    g23929(.A1(new_n24121_), .A2(new_n24120_), .ZN(new_n24122_));
  OAI21_X1   g23930(.A1(new_n24122_), .A2(new_n24115_), .B(\asqrt[49] ), .ZN(new_n24123_));
  INV_X1     g23931(.I(new_n23399_), .ZN(new_n24124_));
  NOR3_X1    g23932(.A1(new_n23757_), .A2(new_n23393_), .A3(new_n23627_), .ZN(new_n24125_));
  INV_X1     g23933(.I(new_n24125_), .ZN(new_n24126_));
  NOR3_X1    g23934(.A1(new_n23627_), .A2(new_n23393_), .A3(new_n24124_), .ZN(new_n24127_));
  AOI22_X1   g23935(.A1(new_n24126_), .A2(new_n24124_), .B1(\asqrt[2] ), .B2(new_n24127_), .ZN(new_n24128_));
  INV_X1     g23936(.I(new_n24128_), .ZN(new_n24129_));
  NAND2_X1   g23937(.A1(new_n24114_), .A2(new_n1806_), .ZN(new_n24130_));
  OAI21_X1   g23938(.A1(new_n24122_), .A2(new_n24130_), .B(new_n24129_), .ZN(new_n24131_));
  AOI21_X1   g23939(.A1(new_n24131_), .A2(new_n24123_), .B(new_n1612_), .ZN(new_n24132_));
  NOR3_X1    g23940(.A1(new_n23404_), .A2(new_n23499_), .A3(new_n23413_), .ZN(new_n24133_));
  NOR3_X1    g23941(.A1(new_n23757_), .A2(new_n23404_), .A3(new_n23413_), .ZN(new_n24134_));
  INV_X1     g23942(.I(new_n24134_), .ZN(new_n24135_));
  AOI22_X1   g23943(.A1(new_n24135_), .A2(new_n23499_), .B1(\asqrt[2] ), .B2(new_n24133_), .ZN(new_n24136_));
  OAI21_X1   g23944(.A1(new_n24120_), .A2(new_n24121_), .B(new_n24114_), .ZN(new_n24137_));
  AOI21_X1   g23945(.A1(new_n24137_), .A2(\asqrt[49] ), .B(\asqrt[50] ), .ZN(new_n24138_));
  AOI21_X1   g23946(.A1(new_n24138_), .A2(new_n24131_), .B(new_n24136_), .ZN(new_n24139_));
  OAI21_X1   g23947(.A1(new_n24139_), .A2(new_n24132_), .B(\asqrt[51] ), .ZN(new_n24140_));
  INV_X1     g23948(.I(new_n24140_), .ZN(new_n24141_));
  NOR2_X1    g23949(.A1(new_n23414_), .A2(new_n23421_), .ZN(new_n24142_));
  NOR3_X1    g23950(.A1(new_n23757_), .A2(new_n23626_), .A3(new_n24142_), .ZN(new_n24143_));
  INV_X1     g23951(.I(new_n24143_), .ZN(new_n24144_));
  NOR3_X1    g23952(.A1(new_n24142_), .A2(new_n23626_), .A3(new_n23420_), .ZN(new_n24145_));
  AOI22_X1   g23953(.A1(new_n24144_), .A2(new_n23420_), .B1(\asqrt[2] ), .B2(new_n24145_), .ZN(new_n24146_));
  NOR3_X1    g23954(.A1(new_n24139_), .A2(new_n24132_), .A3(\asqrt[51] ), .ZN(new_n24147_));
  NOR2_X1    g23955(.A1(new_n24147_), .A2(new_n24146_), .ZN(new_n24148_));
  OAI21_X1   g23956(.A1(new_n24148_), .A2(new_n24141_), .B(\asqrt[52] ), .ZN(new_n24149_));
  INV_X1     g23957(.I(new_n23429_), .ZN(new_n24150_));
  NAND2_X1   g23958(.A1(new_n23431_), .A2(new_n23422_), .ZN(new_n24151_));
  INV_X1     g23959(.I(new_n24151_), .ZN(new_n24152_));
  NOR3_X1    g23960(.A1(new_n24152_), .A2(new_n23423_), .A3(new_n24150_), .ZN(new_n24153_));
  NOR3_X1    g23961(.A1(new_n23757_), .A2(new_n23423_), .A3(new_n24152_), .ZN(new_n24154_));
  INV_X1     g23962(.I(new_n24154_), .ZN(new_n24155_));
  AOI22_X1   g23963(.A1(new_n24155_), .A2(new_n24150_), .B1(\asqrt[2] ), .B2(new_n24153_), .ZN(new_n24156_));
  INV_X1     g23964(.I(new_n24156_), .ZN(new_n24157_));
  NAND2_X1   g23965(.A1(new_n24140_), .A2(new_n1256_), .ZN(new_n24158_));
  OAI21_X1   g23966(.A1(new_n24148_), .A2(new_n24158_), .B(new_n24157_), .ZN(new_n24159_));
  AOI21_X1   g23967(.A1(new_n24159_), .A2(new_n24149_), .B(new_n1103_), .ZN(new_n24160_));
  NOR3_X1    g23968(.A1(new_n23757_), .A2(new_n23434_), .A3(new_n23443_), .ZN(new_n24161_));
  INV_X1     g23969(.I(new_n24161_), .ZN(new_n24162_));
  NOR3_X1    g23970(.A1(new_n23434_), .A2(new_n23498_), .A3(new_n23443_), .ZN(new_n24163_));
  AOI22_X1   g23971(.A1(new_n24162_), .A2(new_n23498_), .B1(\asqrt[2] ), .B2(new_n24163_), .ZN(new_n24164_));
  OAI21_X1   g23972(.A1(new_n24146_), .A2(new_n24147_), .B(new_n24140_), .ZN(new_n24165_));
  AOI21_X1   g23973(.A1(new_n24165_), .A2(\asqrt[52] ), .B(\asqrt[53] ), .ZN(new_n24166_));
  AOI21_X1   g23974(.A1(new_n24166_), .A2(new_n24159_), .B(new_n24164_), .ZN(new_n24167_));
  OAI21_X1   g23975(.A1(new_n24167_), .A2(new_n24160_), .B(\asqrt[54] ), .ZN(new_n24168_));
  INV_X1     g23976(.I(new_n24168_), .ZN(new_n24169_));
  INV_X1     g23977(.I(new_n23445_), .ZN(new_n24170_));
  INV_X1     g23978(.I(new_n23634_), .ZN(new_n24171_));
  NOR3_X1    g23979(.A1(new_n24170_), .A2(new_n24171_), .A3(new_n23450_), .ZN(new_n24172_));
  NOR3_X1    g23980(.A1(new_n23757_), .A2(new_n24170_), .A3(new_n24171_), .ZN(new_n24173_));
  INV_X1     g23981(.I(new_n24173_), .ZN(new_n24174_));
  AOI22_X1   g23982(.A1(new_n24174_), .A2(new_n23450_), .B1(\asqrt[2] ), .B2(new_n24172_), .ZN(new_n24175_));
  NOR3_X1    g23983(.A1(new_n24167_), .A2(new_n24160_), .A3(\asqrt[54] ), .ZN(new_n24176_));
  NOR2_X1    g23984(.A1(new_n24176_), .A2(new_n24175_), .ZN(new_n24177_));
  OAI21_X1   g23985(.A1(new_n24177_), .A2(new_n24169_), .B(\asqrt[55] ), .ZN(new_n24178_));
  INV_X1     g23986(.I(new_n23459_), .ZN(new_n24179_));
  INV_X1     g23987(.I(new_n23452_), .ZN(new_n24180_));
  INV_X1     g23988(.I(new_n23461_), .ZN(new_n24181_));
  NOR2_X1    g23989(.A1(new_n24181_), .A2(new_n24180_), .ZN(new_n24182_));
  NOR3_X1    g23990(.A1(new_n23757_), .A2(new_n23453_), .A3(new_n24182_), .ZN(new_n24183_));
  INV_X1     g23991(.I(new_n24183_), .ZN(new_n24184_));
  NOR3_X1    g23992(.A1(new_n24182_), .A2(new_n23453_), .A3(new_n24179_), .ZN(new_n24185_));
  AOI22_X1   g23993(.A1(new_n24184_), .A2(new_n24179_), .B1(\asqrt[2] ), .B2(new_n24185_), .ZN(new_n24186_));
  INV_X1     g23994(.I(new_n24186_), .ZN(new_n24187_));
  NAND2_X1   g23995(.A1(new_n24168_), .A2(new_n823_), .ZN(new_n24188_));
  OAI21_X1   g23996(.A1(new_n24177_), .A2(new_n24188_), .B(new_n24187_), .ZN(new_n24189_));
  AOI21_X1   g23997(.A1(new_n24189_), .A2(new_n24178_), .B(new_n703_), .ZN(new_n24190_));
  NOR3_X1    g23998(.A1(new_n23464_), .A2(new_n23497_), .A3(new_n23470_), .ZN(new_n24191_));
  NOR3_X1    g23999(.A1(new_n23757_), .A2(new_n23464_), .A3(new_n23470_), .ZN(new_n24192_));
  INV_X1     g24000(.I(new_n24192_), .ZN(new_n24193_));
  AOI22_X1   g24001(.A1(new_n24193_), .A2(new_n23497_), .B1(\asqrt[2] ), .B2(new_n24191_), .ZN(new_n24194_));
  OAI21_X1   g24002(.A1(new_n24175_), .A2(new_n24176_), .B(new_n24168_), .ZN(new_n24195_));
  AOI21_X1   g24003(.A1(new_n24195_), .A2(\asqrt[55] ), .B(\asqrt[56] ), .ZN(new_n24196_));
  AOI21_X1   g24004(.A1(new_n24196_), .A2(new_n24189_), .B(new_n24194_), .ZN(new_n24197_));
  OAI21_X1   g24005(.A1(new_n24197_), .A2(new_n24190_), .B(\asqrt[57] ), .ZN(new_n24198_));
  INV_X1     g24006(.I(new_n24198_), .ZN(new_n24199_));
  INV_X1     g24007(.I(new_n23472_), .ZN(new_n24200_));
  INV_X1     g24008(.I(new_n23638_), .ZN(new_n24201_));
  NOR3_X1    g24009(.A1(new_n23757_), .A2(new_n24200_), .A3(new_n24201_), .ZN(new_n24202_));
  INV_X1     g24010(.I(new_n24202_), .ZN(new_n24203_));
  NOR3_X1    g24011(.A1(new_n24200_), .A2(new_n24201_), .A3(new_n23477_), .ZN(new_n24204_));
  AOI22_X1   g24012(.A1(new_n24203_), .A2(new_n23477_), .B1(\asqrt[2] ), .B2(new_n24204_), .ZN(new_n24205_));
  NOR3_X1    g24013(.A1(new_n24197_), .A2(new_n24190_), .A3(\asqrt[57] ), .ZN(new_n24206_));
  NOR2_X1    g24014(.A1(new_n24206_), .A2(new_n24205_), .ZN(new_n24207_));
  OAI21_X1   g24015(.A1(new_n24207_), .A2(new_n24199_), .B(\asqrt[58] ), .ZN(new_n24208_));
  INV_X1     g24016(.I(new_n23486_), .ZN(new_n24209_));
  INV_X1     g24017(.I(new_n23479_), .ZN(new_n24210_));
  INV_X1     g24018(.I(new_n23488_), .ZN(new_n24211_));
  OAI21_X1   g24019(.A1(new_n24211_), .A2(new_n24210_), .B(new_n23486_), .ZN(new_n24212_));
  NOR2_X1    g24020(.A1(new_n24212_), .A2(new_n23480_), .ZN(new_n24213_));
  NOR2_X1    g24021(.A1(new_n24211_), .A2(new_n24210_), .ZN(new_n24214_));
  NOR3_X1    g24022(.A1(new_n23757_), .A2(new_n23480_), .A3(new_n24214_), .ZN(new_n24215_));
  INV_X1     g24023(.I(new_n24215_), .ZN(new_n24216_));
  AOI22_X1   g24024(.A1(new_n24216_), .A2(new_n24209_), .B1(\asqrt[2] ), .B2(new_n24213_), .ZN(new_n24217_));
  INV_X1     g24025(.I(new_n24217_), .ZN(new_n24218_));
  NAND2_X1   g24026(.A1(new_n24198_), .A2(new_n436_), .ZN(new_n24219_));
  OAI21_X1   g24027(.A1(new_n24207_), .A2(new_n24219_), .B(new_n24218_), .ZN(new_n24220_));
  AOI21_X1   g24028(.A1(new_n24220_), .A2(new_n24208_), .B(new_n327_), .ZN(new_n24221_));
  NOR3_X1    g24029(.A1(new_n23757_), .A2(new_n23658_), .A3(new_n23659_), .ZN(new_n24222_));
  INV_X1     g24030(.I(new_n24222_), .ZN(new_n24223_));
  NOR3_X1    g24031(.A1(new_n23658_), .A2(new_n23496_), .A3(new_n23659_), .ZN(new_n24224_));
  AOI22_X1   g24032(.A1(new_n24223_), .A2(new_n23496_), .B1(\asqrt[2] ), .B2(new_n24224_), .ZN(new_n24225_));
  OAI21_X1   g24033(.A1(new_n24205_), .A2(new_n24206_), .B(new_n24198_), .ZN(new_n24226_));
  AOI21_X1   g24034(.A1(new_n24226_), .A2(\asqrt[58] ), .B(\asqrt[59] ), .ZN(new_n24227_));
  AOI21_X1   g24035(.A1(new_n24227_), .A2(new_n24220_), .B(new_n24225_), .ZN(new_n24228_));
  OAI21_X1   g24036(.A1(new_n24228_), .A2(new_n24221_), .B(\asqrt[60] ), .ZN(new_n24229_));
  INV_X1     g24037(.I(new_n23698_), .ZN(new_n24230_));
  NOR3_X1    g24038(.A1(new_n24230_), .A2(new_n23642_), .A3(new_n23670_), .ZN(new_n24231_));
  NOR3_X1    g24039(.A1(new_n23757_), .A2(new_n23642_), .A3(new_n24230_), .ZN(new_n24232_));
  INV_X1     g24040(.I(new_n24232_), .ZN(new_n24233_));
  AOI22_X1   g24041(.A1(new_n24233_), .A2(new_n23670_), .B1(\asqrt[2] ), .B2(new_n24231_), .ZN(new_n24234_));
  INV_X1     g24042(.I(new_n24234_), .ZN(new_n24235_));
  INV_X1     g24043(.I(new_n24205_), .ZN(new_n24236_));
  INV_X1     g24044(.I(new_n24175_), .ZN(new_n24237_));
  INV_X1     g24045(.I(new_n24146_), .ZN(new_n24238_));
  INV_X1     g24046(.I(new_n24120_), .ZN(new_n24239_));
  INV_X1     g24047(.I(new_n24094_), .ZN(new_n24240_));
  INV_X1     g24048(.I(new_n24068_), .ZN(new_n24241_));
  INV_X1     g24049(.I(new_n24042_), .ZN(new_n24242_));
  INV_X1     g24050(.I(new_n24016_), .ZN(new_n24243_));
  INV_X1     g24051(.I(new_n23990_), .ZN(new_n24244_));
  INV_X1     g24052(.I(new_n23964_), .ZN(new_n24245_));
  INV_X1     g24053(.I(new_n23938_), .ZN(new_n24246_));
  INV_X1     g24054(.I(new_n23912_), .ZN(new_n24247_));
  INV_X1     g24055(.I(new_n23886_), .ZN(new_n24248_));
  INV_X1     g24056(.I(new_n23860_), .ZN(new_n24249_));
  INV_X1     g24057(.I(new_n23834_), .ZN(new_n24250_));
  INV_X1     g24058(.I(new_n23808_), .ZN(new_n24251_));
  INV_X1     g24059(.I(new_n23784_), .ZN(new_n24252_));
  NAND2_X1   g24060(.A1(new_n23711_), .A2(new_n23722_), .ZN(new_n24253_));
  OAI21_X1   g24061(.A1(new_n23696_), .A2(new_n23710_), .B(new_n22907_), .ZN(new_n24254_));
  NAND2_X1   g24062(.A1(new_n24254_), .A2(\a[5] ), .ZN(new_n24255_));
  NAND3_X1   g24063(.A1(new_n24253_), .A2(new_n24255_), .A3(new_n23732_), .ZN(new_n24256_));
  AOI21_X1   g24064(.A1(new_n24256_), .A2(new_n23746_), .B(new_n22337_), .ZN(new_n24257_));
  OAI21_X1   g24065(.A1(new_n23737_), .A2(new_n23725_), .B(\a[6] ), .ZN(new_n24258_));
  NAND3_X1   g24066(.A1(new_n23734_), .A2(new_n23732_), .A3(new_n22912_), .ZN(new_n24259_));
  NAND2_X1   g24067(.A1(new_n23711_), .A2(new_n22911_), .ZN(new_n24260_));
  AOI21_X1   g24068(.A1(new_n24260_), .A2(\asqrt[3] ), .B(\asqrt[4] ), .ZN(new_n24261_));
  AOI22_X1   g24069(.A1(new_n24256_), .A2(new_n24261_), .B1(new_n24258_), .B2(new_n24259_), .ZN(new_n24262_));
  OAI21_X1   g24070(.A1(new_n24262_), .A2(new_n24257_), .B(\asqrt[5] ), .ZN(new_n24263_));
  NAND2_X1   g24071(.A1(new_n24263_), .A2(new_n20806_), .ZN(new_n24264_));
  OAI21_X1   g24072(.A1(new_n24264_), .A2(new_n23751_), .B(new_n23759_), .ZN(new_n24265_));
  AOI21_X1   g24073(.A1(new_n24265_), .A2(new_n23752_), .B(new_n20262_), .ZN(new_n24266_));
  INV_X1     g24074(.I(new_n23745_), .ZN(new_n24267_));
  AOI21_X1   g24075(.A1(\a[5] ), .A2(new_n24254_), .B(new_n23725_), .ZN(new_n24268_));
  AOI21_X1   g24076(.A1(new_n24268_), .A2(new_n24253_), .B(new_n23712_), .ZN(new_n24269_));
  OAI21_X1   g24077(.A1(new_n24269_), .A2(new_n22337_), .B(new_n21620_), .ZN(new_n24270_));
  OAI21_X1   g24078(.A1(new_n24270_), .A2(new_n24262_), .B(new_n24267_), .ZN(new_n24271_));
  NAND2_X1   g24079(.A1(new_n24271_), .A2(new_n24263_), .ZN(new_n24272_));
  AOI21_X1   g24080(.A1(new_n24272_), .A2(\asqrt[6] ), .B(\asqrt[7] ), .ZN(new_n24273_));
  AOI21_X1   g24081(.A1(new_n24273_), .A2(new_n24265_), .B(new_n23767_), .ZN(new_n24274_));
  OAI21_X1   g24082(.A1(new_n24274_), .A2(new_n24266_), .B(\asqrt[8] ), .ZN(new_n24275_));
  NAND2_X1   g24083(.A1(new_n24275_), .A2(new_n18792_), .ZN(new_n24276_));
  OAI21_X1   g24084(.A1(new_n24276_), .A2(new_n23778_), .B(new_n24252_), .ZN(new_n24277_));
  NAND3_X1   g24085(.A1(new_n24277_), .A2(new_n18275_), .A3(new_n23779_), .ZN(new_n24278_));
  AOI22_X1   g24086(.A1(new_n24278_), .A2(new_n23793_), .B1(new_n23801_), .B2(\asqrt[10] ), .ZN(new_n24279_));
  OAI21_X1   g24087(.A1(new_n24279_), .A2(new_n17623_), .B(new_n16881_), .ZN(new_n24280_));
  OAI21_X1   g24088(.A1(new_n24280_), .A2(new_n23803_), .B(new_n24251_), .ZN(new_n24281_));
  AOI21_X1   g24089(.A1(new_n24281_), .A2(new_n23804_), .B(new_n16389_), .ZN(new_n24282_));
  AOI21_X1   g24090(.A1(new_n24277_), .A2(new_n23779_), .B(new_n18275_), .ZN(new_n24283_));
  NOR3_X1    g24091(.A1(new_n24274_), .A2(new_n24266_), .A3(\asqrt[8] ), .ZN(new_n24284_));
  OAI21_X1   g24092(.A1(new_n23775_), .A2(new_n24284_), .B(new_n24275_), .ZN(new_n24285_));
  AOI21_X1   g24093(.A1(new_n24285_), .A2(\asqrt[9] ), .B(\asqrt[10] ), .ZN(new_n24286_));
  AOI21_X1   g24094(.A1(new_n24286_), .A2(new_n24277_), .B(new_n23792_), .ZN(new_n24287_));
  NOR3_X1    g24095(.A1(new_n24287_), .A2(\asqrt[11] ), .A3(new_n24283_), .ZN(new_n24288_));
  OAI22_X1   g24096(.A1(new_n24288_), .A2(new_n23800_), .B1(new_n24279_), .B2(new_n17623_), .ZN(new_n24289_));
  AOI21_X1   g24097(.A1(new_n24289_), .A2(\asqrt[12] ), .B(\asqrt[13] ), .ZN(new_n24290_));
  AOI21_X1   g24098(.A1(new_n24290_), .A2(new_n24281_), .B(new_n23816_), .ZN(new_n24291_));
  OAI21_X1   g24099(.A1(new_n24291_), .A2(new_n24282_), .B(\asqrt[14] ), .ZN(new_n24292_));
  NAND2_X1   g24100(.A1(new_n24292_), .A2(new_n15067_), .ZN(new_n24293_));
  OAI21_X1   g24101(.A1(new_n24293_), .A2(new_n23827_), .B(new_n24250_), .ZN(new_n24294_));
  AOI21_X1   g24102(.A1(new_n24294_), .A2(new_n23828_), .B(new_n14601_), .ZN(new_n24295_));
  NOR3_X1    g24103(.A1(new_n24291_), .A2(\asqrt[14] ), .A3(new_n24282_), .ZN(new_n24296_));
  OAI21_X1   g24104(.A1(new_n23824_), .A2(new_n24296_), .B(new_n24292_), .ZN(new_n24297_));
  AOI21_X1   g24105(.A1(new_n24297_), .A2(\asqrt[15] ), .B(\asqrt[16] ), .ZN(new_n24298_));
  AOI21_X1   g24106(.A1(new_n24298_), .A2(new_n24294_), .B(new_n23842_), .ZN(new_n24299_));
  OAI21_X1   g24107(.A1(new_n24299_), .A2(new_n24295_), .B(\asqrt[17] ), .ZN(new_n24300_));
  NAND2_X1   g24108(.A1(new_n24300_), .A2(new_n13353_), .ZN(new_n24301_));
  OAI21_X1   g24109(.A1(new_n24301_), .A2(new_n23853_), .B(new_n24249_), .ZN(new_n24302_));
  AOI21_X1   g24110(.A1(new_n24302_), .A2(new_n23854_), .B(new_n12913_), .ZN(new_n24303_));
  NOR3_X1    g24111(.A1(new_n24299_), .A2(\asqrt[17] ), .A3(new_n24295_), .ZN(new_n24304_));
  OAI21_X1   g24112(.A1(new_n23850_), .A2(new_n24304_), .B(new_n24300_), .ZN(new_n24305_));
  AOI21_X1   g24113(.A1(new_n24305_), .A2(\asqrt[18] ), .B(\asqrt[19] ), .ZN(new_n24306_));
  AOI21_X1   g24114(.A1(new_n24306_), .A2(new_n24302_), .B(new_n23868_), .ZN(new_n24307_));
  OAI21_X1   g24115(.A1(new_n24307_), .A2(new_n24303_), .B(\asqrt[20] ), .ZN(new_n24308_));
  NAND2_X1   g24116(.A1(new_n24308_), .A2(new_n11736_), .ZN(new_n24309_));
  OAI21_X1   g24117(.A1(new_n24309_), .A2(new_n23879_), .B(new_n24248_), .ZN(new_n24310_));
  AOI21_X1   g24118(.A1(new_n24310_), .A2(new_n23880_), .B(new_n11326_), .ZN(new_n24311_));
  NOR3_X1    g24119(.A1(new_n24307_), .A2(\asqrt[20] ), .A3(new_n24303_), .ZN(new_n24312_));
  OAI21_X1   g24120(.A1(new_n23876_), .A2(new_n24312_), .B(new_n24308_), .ZN(new_n24313_));
  AOI21_X1   g24121(.A1(new_n24313_), .A2(\asqrt[21] ), .B(\asqrt[22] ), .ZN(new_n24314_));
  AOI21_X1   g24122(.A1(new_n24314_), .A2(new_n24310_), .B(new_n23894_), .ZN(new_n24315_));
  OAI21_X1   g24123(.A1(new_n24315_), .A2(new_n24311_), .B(\asqrt[23] ), .ZN(new_n24316_));
  NAND2_X1   g24124(.A1(new_n24316_), .A2(new_n10221_), .ZN(new_n24317_));
  OAI21_X1   g24125(.A1(new_n24317_), .A2(new_n23905_), .B(new_n24247_), .ZN(new_n24318_));
  AOI21_X1   g24126(.A1(new_n24318_), .A2(new_n23906_), .B(new_n9846_), .ZN(new_n24319_));
  NOR3_X1    g24127(.A1(new_n24315_), .A2(\asqrt[23] ), .A3(new_n24311_), .ZN(new_n24320_));
  OAI21_X1   g24128(.A1(new_n23902_), .A2(new_n24320_), .B(new_n24316_), .ZN(new_n24321_));
  AOI21_X1   g24129(.A1(new_n24321_), .A2(\asqrt[24] ), .B(\asqrt[25] ), .ZN(new_n24322_));
  AOI21_X1   g24130(.A1(new_n24322_), .A2(new_n24318_), .B(new_n23920_), .ZN(new_n24323_));
  OAI21_X1   g24131(.A1(new_n24323_), .A2(new_n24319_), .B(\asqrt[26] ), .ZN(new_n24324_));
  NAND2_X1   g24132(.A1(new_n24324_), .A2(new_n8826_), .ZN(new_n24325_));
  OAI21_X1   g24133(.A1(new_n24325_), .A2(new_n23931_), .B(new_n24246_), .ZN(new_n24326_));
  AOI21_X1   g24134(.A1(new_n24326_), .A2(new_n23932_), .B(new_n8483_), .ZN(new_n24327_));
  NOR3_X1    g24135(.A1(new_n24323_), .A2(\asqrt[26] ), .A3(new_n24319_), .ZN(new_n24328_));
  OAI21_X1   g24136(.A1(new_n23928_), .A2(new_n24328_), .B(new_n24324_), .ZN(new_n24329_));
  AOI21_X1   g24137(.A1(new_n24329_), .A2(\asqrt[27] ), .B(\asqrt[28] ), .ZN(new_n24330_));
  AOI21_X1   g24138(.A1(new_n24330_), .A2(new_n24326_), .B(new_n23946_), .ZN(new_n24331_));
  OAI21_X1   g24139(.A1(new_n24331_), .A2(new_n24327_), .B(\asqrt[29] ), .ZN(new_n24332_));
  NAND2_X1   g24140(.A1(new_n24332_), .A2(new_n7539_), .ZN(new_n24333_));
  OAI21_X1   g24141(.A1(new_n24333_), .A2(new_n23957_), .B(new_n24245_), .ZN(new_n24334_));
  AOI21_X1   g24142(.A1(new_n24334_), .A2(new_n23958_), .B(new_n7229_), .ZN(new_n24335_));
  NOR3_X1    g24143(.A1(new_n24331_), .A2(\asqrt[29] ), .A3(new_n24327_), .ZN(new_n24336_));
  OAI21_X1   g24144(.A1(new_n23954_), .A2(new_n24336_), .B(new_n24332_), .ZN(new_n24337_));
  AOI21_X1   g24145(.A1(new_n24337_), .A2(\asqrt[30] ), .B(\asqrt[31] ), .ZN(new_n24338_));
  AOI21_X1   g24146(.A1(new_n24338_), .A2(new_n24334_), .B(new_n23972_), .ZN(new_n24339_));
  OAI21_X1   g24147(.A1(new_n24339_), .A2(new_n24335_), .B(\asqrt[32] ), .ZN(new_n24340_));
  NAND2_X1   g24148(.A1(new_n24340_), .A2(new_n6356_), .ZN(new_n24341_));
  OAI21_X1   g24149(.A1(new_n24341_), .A2(new_n23983_), .B(new_n24244_), .ZN(new_n24342_));
  AOI21_X1   g24150(.A1(new_n24342_), .A2(new_n23984_), .B(new_n6077_), .ZN(new_n24343_));
  NOR3_X1    g24151(.A1(new_n24339_), .A2(\asqrt[32] ), .A3(new_n24335_), .ZN(new_n24344_));
  OAI21_X1   g24152(.A1(new_n23980_), .A2(new_n24344_), .B(new_n24340_), .ZN(new_n24345_));
  AOI21_X1   g24153(.A1(new_n24345_), .A2(\asqrt[33] ), .B(\asqrt[34] ), .ZN(new_n24346_));
  AOI21_X1   g24154(.A1(new_n24346_), .A2(new_n24342_), .B(new_n23998_), .ZN(new_n24347_));
  OAI21_X1   g24155(.A1(new_n24347_), .A2(new_n24343_), .B(\asqrt[35] ), .ZN(new_n24348_));
  NAND2_X1   g24156(.A1(new_n24348_), .A2(new_n5277_), .ZN(new_n24349_));
  OAI21_X1   g24157(.A1(new_n24349_), .A2(new_n24009_), .B(new_n24243_), .ZN(new_n24350_));
  AOI21_X1   g24158(.A1(new_n24350_), .A2(new_n24010_), .B(new_n5024_), .ZN(new_n24351_));
  NOR3_X1    g24159(.A1(new_n24347_), .A2(\asqrt[35] ), .A3(new_n24343_), .ZN(new_n24352_));
  OAI21_X1   g24160(.A1(new_n24006_), .A2(new_n24352_), .B(new_n24348_), .ZN(new_n24353_));
  AOI21_X1   g24161(.A1(new_n24353_), .A2(\asqrt[36] ), .B(\asqrt[37] ), .ZN(new_n24354_));
  AOI21_X1   g24162(.A1(new_n24354_), .A2(new_n24350_), .B(new_n24024_), .ZN(new_n24355_));
  OAI21_X1   g24163(.A1(new_n24355_), .A2(new_n24351_), .B(\asqrt[38] ), .ZN(new_n24356_));
  NAND2_X1   g24164(.A1(new_n24356_), .A2(new_n4298_), .ZN(new_n24357_));
  OAI21_X1   g24165(.A1(new_n24357_), .A2(new_n24035_), .B(new_n24242_), .ZN(new_n24358_));
  AOI21_X1   g24166(.A1(new_n24358_), .A2(new_n24036_), .B(new_n4071_), .ZN(new_n24359_));
  NOR3_X1    g24167(.A1(new_n24355_), .A2(\asqrt[38] ), .A3(new_n24351_), .ZN(new_n24360_));
  OAI21_X1   g24168(.A1(new_n24032_), .A2(new_n24360_), .B(new_n24356_), .ZN(new_n24361_));
  AOI21_X1   g24169(.A1(new_n24361_), .A2(\asqrt[39] ), .B(\asqrt[40] ), .ZN(new_n24362_));
  AOI21_X1   g24170(.A1(new_n24362_), .A2(new_n24358_), .B(new_n24050_), .ZN(new_n24363_));
  OAI21_X1   g24171(.A1(new_n24363_), .A2(new_n24359_), .B(\asqrt[41] ), .ZN(new_n24364_));
  NAND2_X1   g24172(.A1(new_n24364_), .A2(new_n3419_), .ZN(new_n24365_));
  OAI21_X1   g24173(.A1(new_n24365_), .A2(new_n24061_), .B(new_n24241_), .ZN(new_n24366_));
  AOI21_X1   g24174(.A1(new_n24366_), .A2(new_n24062_), .B(new_n3218_), .ZN(new_n24367_));
  NOR3_X1    g24175(.A1(new_n24363_), .A2(\asqrt[41] ), .A3(new_n24359_), .ZN(new_n24368_));
  OAI21_X1   g24176(.A1(new_n24058_), .A2(new_n24368_), .B(new_n24364_), .ZN(new_n24369_));
  AOI21_X1   g24177(.A1(new_n24369_), .A2(\asqrt[42] ), .B(\asqrt[43] ), .ZN(new_n24370_));
  AOI21_X1   g24178(.A1(new_n24370_), .A2(new_n24366_), .B(new_n24076_), .ZN(new_n24371_));
  OAI21_X1   g24179(.A1(new_n24371_), .A2(new_n24367_), .B(\asqrt[44] ), .ZN(new_n24372_));
  NAND2_X1   g24180(.A1(new_n24372_), .A2(new_n2641_), .ZN(new_n24373_));
  OAI21_X1   g24181(.A1(new_n24373_), .A2(new_n24087_), .B(new_n24240_), .ZN(new_n24374_));
  AOI21_X1   g24182(.A1(new_n24374_), .A2(new_n24088_), .B(new_n2465_), .ZN(new_n24375_));
  NOR3_X1    g24183(.A1(new_n24371_), .A2(\asqrt[44] ), .A3(new_n24367_), .ZN(new_n24376_));
  OAI21_X1   g24184(.A1(new_n24084_), .A2(new_n24376_), .B(new_n24372_), .ZN(new_n24377_));
  AOI21_X1   g24185(.A1(new_n24377_), .A2(\asqrt[45] ), .B(\asqrt[46] ), .ZN(new_n24378_));
  AOI21_X1   g24186(.A1(new_n24378_), .A2(new_n24374_), .B(new_n24102_), .ZN(new_n24379_));
  OAI21_X1   g24187(.A1(new_n24379_), .A2(new_n24375_), .B(\asqrt[47] ), .ZN(new_n24380_));
  NAND2_X1   g24188(.A1(new_n24380_), .A2(new_n1956_), .ZN(new_n24381_));
  OAI21_X1   g24189(.A1(new_n24381_), .A2(new_n24113_), .B(new_n24239_), .ZN(new_n24382_));
  AOI21_X1   g24190(.A1(new_n24382_), .A2(new_n24114_), .B(new_n1806_), .ZN(new_n24383_));
  NOR3_X1    g24191(.A1(new_n24379_), .A2(\asqrt[47] ), .A3(new_n24375_), .ZN(new_n24384_));
  OAI21_X1   g24192(.A1(new_n24110_), .A2(new_n24384_), .B(new_n24380_), .ZN(new_n24385_));
  AOI21_X1   g24193(.A1(new_n24385_), .A2(\asqrt[48] ), .B(\asqrt[49] ), .ZN(new_n24386_));
  AOI21_X1   g24194(.A1(new_n24386_), .A2(new_n24382_), .B(new_n24128_), .ZN(new_n24387_));
  OAI21_X1   g24195(.A1(new_n24387_), .A2(new_n24383_), .B(\asqrt[50] ), .ZN(new_n24388_));
  NAND2_X1   g24196(.A1(new_n24388_), .A2(new_n1376_), .ZN(new_n24389_));
  OAI21_X1   g24197(.A1(new_n24389_), .A2(new_n24139_), .B(new_n24238_), .ZN(new_n24390_));
  AOI21_X1   g24198(.A1(new_n24390_), .A2(new_n24140_), .B(new_n1256_), .ZN(new_n24391_));
  NOR3_X1    g24199(.A1(new_n24387_), .A2(\asqrt[50] ), .A3(new_n24383_), .ZN(new_n24392_));
  OAI21_X1   g24200(.A1(new_n24136_), .A2(new_n24392_), .B(new_n24388_), .ZN(new_n24393_));
  AOI21_X1   g24201(.A1(new_n24393_), .A2(\asqrt[51] ), .B(\asqrt[52] ), .ZN(new_n24394_));
  AOI21_X1   g24202(.A1(new_n24394_), .A2(new_n24390_), .B(new_n24156_), .ZN(new_n24395_));
  OAI21_X1   g24203(.A1(new_n24395_), .A2(new_n24391_), .B(\asqrt[53] ), .ZN(new_n24396_));
  NAND2_X1   g24204(.A1(new_n24396_), .A2(new_n904_), .ZN(new_n24397_));
  OAI21_X1   g24205(.A1(new_n24397_), .A2(new_n24167_), .B(new_n24237_), .ZN(new_n24398_));
  AOI21_X1   g24206(.A1(new_n24398_), .A2(new_n24168_), .B(new_n823_), .ZN(new_n24399_));
  NOR3_X1    g24207(.A1(new_n24395_), .A2(\asqrt[53] ), .A3(new_n24391_), .ZN(new_n24400_));
  OAI21_X1   g24208(.A1(new_n24164_), .A2(new_n24400_), .B(new_n24396_), .ZN(new_n24401_));
  AOI21_X1   g24209(.A1(new_n24401_), .A2(\asqrt[54] ), .B(\asqrt[55] ), .ZN(new_n24402_));
  AOI21_X1   g24210(.A1(new_n24402_), .A2(new_n24398_), .B(new_n24186_), .ZN(new_n24403_));
  OAI21_X1   g24211(.A1(new_n24403_), .A2(new_n24399_), .B(\asqrt[56] ), .ZN(new_n24404_));
  NAND2_X1   g24212(.A1(new_n24404_), .A2(new_n531_), .ZN(new_n24405_));
  OAI21_X1   g24213(.A1(new_n24405_), .A2(new_n24197_), .B(new_n24236_), .ZN(new_n24406_));
  AOI21_X1   g24214(.A1(new_n24406_), .A2(new_n24198_), .B(new_n436_), .ZN(new_n24407_));
  NOR3_X1    g24215(.A1(new_n24403_), .A2(\asqrt[56] ), .A3(new_n24399_), .ZN(new_n24408_));
  OAI21_X1   g24216(.A1(new_n24194_), .A2(new_n24408_), .B(new_n24404_), .ZN(new_n24409_));
  AOI21_X1   g24217(.A1(new_n24409_), .A2(\asqrt[57] ), .B(\asqrt[58] ), .ZN(new_n24410_));
  AOI21_X1   g24218(.A1(new_n24410_), .A2(new_n24406_), .B(new_n24217_), .ZN(new_n24411_));
  OAI21_X1   g24219(.A1(new_n24411_), .A2(new_n24407_), .B(\asqrt[59] ), .ZN(new_n24412_));
  NAND2_X1   g24220(.A1(new_n24412_), .A2(new_n306_), .ZN(new_n24413_));
  OAI21_X1   g24221(.A1(new_n24413_), .A2(new_n24228_), .B(new_n24235_), .ZN(new_n24414_));
  AOI21_X1   g24222(.A1(new_n24414_), .A2(new_n24229_), .B(new_n218_), .ZN(new_n24415_));
  NAND2_X1   g24223(.A1(new_n23682_), .A2(new_n23671_), .ZN(new_n24416_));
  NAND3_X1   g24224(.A1(\asqrt[2] ), .A2(new_n23650_), .A3(new_n24416_), .ZN(new_n24417_));
  AND3_X2    g24225(.A1(new_n23650_), .A2(new_n23656_), .A3(new_n24416_), .Z(new_n24418_));
  AOI22_X1   g24226(.A1(new_n24417_), .A2(new_n23657_), .B1(\asqrt[2] ), .B2(new_n24418_), .ZN(new_n24419_));
  NOR3_X1    g24227(.A1(new_n24411_), .A2(\asqrt[59] ), .A3(new_n24407_), .ZN(new_n24420_));
  OAI21_X1   g24228(.A1(new_n24225_), .A2(new_n24420_), .B(new_n24412_), .ZN(new_n24421_));
  AOI21_X1   g24229(.A1(new_n24421_), .A2(\asqrt[60] ), .B(\asqrt[61] ), .ZN(new_n24422_));
  AOI21_X1   g24230(.A1(new_n24422_), .A2(new_n24414_), .B(new_n24419_), .ZN(new_n24423_));
  OAI21_X1   g24231(.A1(new_n24423_), .A2(new_n24415_), .B(\asqrt[62] ), .ZN(new_n24424_));
  NOR3_X1    g24232(.A1(new_n23664_), .A2(new_n23697_), .A3(new_n23713_), .ZN(new_n24425_));
  NOR3_X1    g24233(.A1(new_n23757_), .A2(new_n23664_), .A3(new_n23713_), .ZN(new_n24426_));
  INV_X1     g24234(.I(new_n24426_), .ZN(new_n24427_));
  AOI22_X1   g24235(.A1(new_n24427_), .A2(new_n23697_), .B1(\asqrt[2] ), .B2(new_n24425_), .ZN(new_n24428_));
  NOR3_X1    g24236(.A1(new_n24423_), .A2(\asqrt[62] ), .A3(new_n24415_), .ZN(new_n24429_));
  OAI21_X1   g24237(.A1(new_n24428_), .A2(new_n24429_), .B(new_n24424_), .ZN(new_n24430_));
  INV_X1     g24238(.I(new_n23675_), .ZN(new_n24431_));
  INV_X1     g24239(.I(new_n23715_), .ZN(new_n24432_));
  NOR3_X1    g24240(.A1(new_n23757_), .A2(new_n24431_), .A3(new_n24432_), .ZN(new_n24433_));
  INV_X1     g24241(.I(new_n24433_), .ZN(new_n24434_));
  NOR3_X1    g24242(.A1(new_n24431_), .A2(new_n24432_), .A3(new_n23680_), .ZN(new_n24435_));
  AOI22_X1   g24243(.A1(new_n24434_), .A2(new_n23680_), .B1(\asqrt[2] ), .B2(new_n24435_), .ZN(new_n24436_));
  INV_X1     g24244(.I(new_n24436_), .ZN(new_n24437_));
  NOR2_X1    g24245(.A1(new_n23716_), .A2(new_n23704_), .ZN(new_n24438_));
  NAND2_X1   g24246(.A1(\asqrt[2] ), .A2(new_n24438_), .ZN(new_n24439_));
  AND3_X2    g24247(.A1(new_n24437_), .A2(new_n23733_), .A3(new_n24439_), .Z(new_n24440_));
  AOI21_X1   g24248(.A1(new_n24430_), .A2(new_n24440_), .B(\asqrt[63] ), .ZN(new_n24441_));
  NOR3_X1    g24249(.A1(new_n24228_), .A2(new_n24221_), .A3(\asqrt[60] ), .ZN(new_n24442_));
  NOR2_X1    g24250(.A1(new_n24442_), .A2(new_n24234_), .ZN(new_n24443_));
  INV_X1     g24251(.I(new_n24419_), .ZN(new_n24444_));
  NAND2_X1   g24252(.A1(new_n24229_), .A2(new_n218_), .ZN(new_n24445_));
  OAI21_X1   g24253(.A1(new_n24443_), .A2(new_n24445_), .B(new_n24444_), .ZN(new_n24446_));
  OAI21_X1   g24254(.A1(new_n24234_), .A2(new_n24442_), .B(new_n24229_), .ZN(new_n24447_));
  AOI21_X1   g24255(.A1(new_n24447_), .A2(\asqrt[61] ), .B(\asqrt[62] ), .ZN(new_n24448_));
  AOI21_X1   g24256(.A1(new_n24448_), .A2(new_n24446_), .B(new_n24428_), .ZN(new_n24449_));
  AOI21_X1   g24257(.A1(\asqrt[2] ), .A2(new_n23691_), .B(new_n23687_), .ZN(new_n24450_));
  NOR2_X1    g24258(.A1(new_n24438_), .A2(new_n193_), .ZN(new_n24451_));
  INV_X1     g24259(.I(new_n24451_), .ZN(new_n24452_));
  NAND2_X1   g24260(.A1(new_n24424_), .A2(new_n24436_), .ZN(new_n24453_));
  OAI22_X1   g24261(.A1(new_n24453_), .A2(new_n24449_), .B1(new_n24450_), .B2(new_n24452_), .ZN(new_n24454_));
  OAI21_X1   g24262(.A1(new_n24441_), .A2(new_n24454_), .B(new_n22908_), .ZN(new_n24455_));
  INV_X1     g24263(.I(new_n24229_), .ZN(new_n24456_));
  OAI21_X1   g24264(.A1(new_n24443_), .A2(new_n24456_), .B(\asqrt[61] ), .ZN(new_n24457_));
  AOI21_X1   g24265(.A1(new_n24446_), .A2(new_n24457_), .B(new_n207_), .ZN(new_n24458_));
  OAI21_X1   g24266(.A1(new_n24449_), .A2(new_n24458_), .B(new_n24440_), .ZN(new_n24459_));
  NAND2_X1   g24267(.A1(new_n24459_), .A2(new_n193_), .ZN(new_n24460_));
  INV_X1     g24268(.I(new_n24428_), .ZN(new_n24461_));
  NAND2_X1   g24269(.A1(new_n24457_), .A2(new_n207_), .ZN(new_n24462_));
  OAI21_X1   g24270(.A1(new_n24462_), .A2(new_n24423_), .B(new_n24461_), .ZN(new_n24463_));
  NOR2_X1    g24271(.A1(new_n24458_), .A2(new_n24437_), .ZN(new_n24464_));
  NAND2_X1   g24272(.A1(new_n24464_), .A2(new_n24463_), .ZN(new_n24465_));
  NOR2_X1    g24273(.A1(new_n24450_), .A2(new_n24452_), .ZN(new_n24466_));
  NOR2_X1    g24274(.A1(new_n24466_), .A2(new_n23757_), .ZN(new_n24467_));
  NAND3_X1   g24275(.A1(new_n24460_), .A2(new_n24465_), .A3(new_n24467_), .ZN(new_n24468_));
  AND3_X2    g24276(.A1(new_n24455_), .A2(new_n24468_), .A3(new_n22907_), .Z(new_n24469_));
  AOI21_X1   g24277(.A1(new_n24455_), .A2(new_n24468_), .B(new_n22907_), .ZN(new_n24470_));
  NOR2_X1    g24278(.A1(new_n24469_), .A2(new_n24470_), .ZN(new_n24471_));
  AOI21_X1   g24279(.A1(new_n24464_), .A2(new_n24463_), .B(new_n24466_), .ZN(new_n24472_));
  AOI21_X1   g24280(.A1(new_n24460_), .A2(new_n24472_), .B(new_n22909_), .ZN(new_n24473_));
  INV_X1     g24281(.I(\a[2] ), .ZN(new_n24474_));
  OAI21_X1   g24282(.A1(\a[0] ), .A2(\a[1] ), .B(new_n24474_), .ZN(new_n24475_));
  NOR2_X1    g24283(.A1(new_n24466_), .A2(new_n24474_), .ZN(new_n24476_));
  INV_X1     g24284(.I(new_n24476_), .ZN(new_n24477_));
  AOI21_X1   g24285(.A1(new_n24464_), .A2(new_n24463_), .B(new_n24477_), .ZN(new_n24478_));
  INV_X1     g24286(.I(new_n24478_), .ZN(new_n24479_));
  OAI21_X1   g24287(.A1(new_n24479_), .A2(new_n24441_), .B(new_n24475_), .ZN(new_n24480_));
  INV_X1     g24288(.I(\a[3] ), .ZN(new_n24481_));
  NAND2_X1   g24289(.A1(new_n24460_), .A2(new_n24472_), .ZN(\asqrt[1] ));
  AOI21_X1   g24290(.A1(\asqrt[1] ), .A2(new_n24474_), .B(new_n24481_), .ZN(new_n24483_));
  OAI21_X1   g24291(.A1(new_n24483_), .A2(new_n24473_), .B(new_n24480_), .ZN(new_n24484_));
  NAND2_X1   g24292(.A1(new_n24460_), .A2(new_n24478_), .ZN(new_n24485_));
  NAND3_X1   g24293(.A1(new_n24455_), .A2(new_n24485_), .A3(new_n24475_), .ZN(new_n24486_));
  OAI21_X1   g24294(.A1(new_n24486_), .A2(new_n24483_), .B(new_n23757_), .ZN(new_n24487_));
  NAND2_X1   g24295(.A1(new_n24487_), .A2(new_n24484_), .ZN(new_n24488_));
  OAI21_X1   g24296(.A1(new_n24488_), .A2(new_n24471_), .B(new_n22906_), .ZN(new_n24489_));
  NOR3_X1    g24297(.A1(new_n24268_), .A2(new_n23712_), .A3(new_n23724_), .ZN(new_n24490_));
  NAND3_X1   g24298(.A1(\asqrt[1] ), .A2(new_n23746_), .A3(new_n24253_), .ZN(new_n24491_));
  AOI22_X1   g24299(.A1(new_n24491_), .A2(new_n24268_), .B1(\asqrt[1] ), .B2(new_n24490_), .ZN(new_n24492_));
  AOI21_X1   g24300(.A1(new_n24488_), .A2(new_n24471_), .B(new_n24492_), .ZN(new_n24493_));
  AOI21_X1   g24301(.A1(new_n24493_), .A2(new_n24489_), .B(\asqrt[4] ), .ZN(new_n24494_));
  NOR2_X1    g24302(.A1(new_n23738_), .A2(new_n23735_), .ZN(new_n24495_));
  NOR2_X1    g24303(.A1(new_n23730_), .A2(new_n23740_), .ZN(new_n24496_));
  INV_X1     g24304(.I(new_n24496_), .ZN(new_n24497_));
  NAND4_X1   g24305(.A1(\asqrt[1] ), .A2(new_n23731_), .A3(new_n24495_), .A4(new_n24497_), .ZN(new_n24498_));
  INV_X1     g24306(.I(\asqrt[1] ), .ZN(new_n24499_));
  NOR3_X1    g24307(.A1(new_n24499_), .A2(new_n24257_), .A3(new_n24496_), .ZN(new_n24500_));
  OAI21_X1   g24308(.A1(new_n24500_), .A2(new_n24495_), .B(new_n24498_), .ZN(new_n24501_));
  INV_X1     g24309(.I(new_n24501_), .ZN(new_n24502_));
  INV_X1     g24310(.I(new_n24492_), .ZN(new_n24503_));
  NAND2_X1   g24311(.A1(new_n24488_), .A2(new_n24471_), .ZN(new_n24504_));
  AOI21_X1   g24312(.A1(new_n24489_), .A2(new_n24504_), .B(new_n24503_), .ZN(new_n24505_));
  NOR3_X1    g24313(.A1(new_n24494_), .A2(new_n24505_), .A3(new_n24502_), .ZN(new_n24506_));
  NOR2_X1    g24314(.A1(new_n24506_), .A2(\asqrt[5] ), .ZN(new_n24507_));
  NOR2_X1    g24315(.A1(new_n24270_), .A2(new_n24262_), .ZN(new_n24508_));
  NOR3_X1    g24316(.A1(new_n24499_), .A2(new_n23742_), .A3(new_n24508_), .ZN(new_n24509_));
  INV_X1     g24317(.I(new_n24509_), .ZN(new_n24510_));
  NOR3_X1    g24318(.A1(new_n24508_), .A2(new_n23742_), .A3(new_n24267_), .ZN(new_n24511_));
  AOI22_X1   g24319(.A1(new_n24510_), .A2(new_n24267_), .B1(\asqrt[1] ), .B2(new_n24511_), .ZN(new_n24512_));
  INV_X1     g24320(.I(new_n24512_), .ZN(new_n24513_));
  OAI21_X1   g24321(.A1(new_n24494_), .A2(new_n24505_), .B(new_n24502_), .ZN(new_n24514_));
  NAND2_X1   g24322(.A1(new_n24514_), .A2(new_n24513_), .ZN(new_n24515_));
  OAI21_X1   g24323(.A1(new_n24507_), .A2(new_n24515_), .B(new_n20806_), .ZN(new_n24516_));
  NOR3_X1    g24324(.A1(new_n23753_), .A2(new_n23761_), .A3(new_n23759_), .ZN(new_n24517_));
  NOR3_X1    g24325(.A1(new_n24499_), .A2(new_n23753_), .A3(new_n23761_), .ZN(new_n24518_));
  INV_X1     g24326(.I(new_n24518_), .ZN(new_n24519_));
  AOI22_X1   g24327(.A1(new_n24519_), .A2(new_n23759_), .B1(\asqrt[1] ), .B2(new_n24517_), .ZN(new_n24520_));
  OAI21_X1   g24328(.A1(\asqrt[5] ), .A2(new_n24506_), .B(new_n24514_), .ZN(new_n24521_));
  AOI21_X1   g24329(.A1(new_n24521_), .A2(new_n24512_), .B(new_n24520_), .ZN(new_n24522_));
  AOI21_X1   g24330(.A1(new_n24522_), .A2(new_n24516_), .B(\asqrt[7] ), .ZN(new_n24523_));
  NAND2_X1   g24331(.A1(new_n24273_), .A2(new_n24265_), .ZN(new_n24524_));
  NAND3_X1   g24332(.A1(\asqrt[1] ), .A2(new_n23763_), .A3(new_n24524_), .ZN(new_n24525_));
  AND3_X2    g24333(.A1(new_n23763_), .A2(new_n23767_), .A3(new_n24524_), .Z(new_n24526_));
  AOI22_X1   g24334(.A1(new_n24525_), .A2(new_n23768_), .B1(\asqrt[1] ), .B2(new_n24526_), .ZN(new_n24527_));
  INV_X1     g24335(.I(new_n24520_), .ZN(new_n24528_));
  INV_X1     g24336(.I(new_n24514_), .ZN(new_n24529_));
  OAI21_X1   g24337(.A1(new_n24507_), .A2(new_n24529_), .B(new_n24512_), .ZN(new_n24530_));
  AOI21_X1   g24338(.A1(new_n24516_), .A2(new_n24530_), .B(new_n24528_), .ZN(new_n24531_));
  NOR3_X1    g24339(.A1(new_n24523_), .A2(new_n24531_), .A3(new_n24527_), .ZN(new_n24532_));
  NOR2_X1    g24340(.A1(new_n24532_), .A2(\asqrt[8] ), .ZN(new_n24533_));
  INV_X1     g24341(.I(new_n23775_), .ZN(new_n24534_));
  NOR3_X1    g24342(.A1(new_n23771_), .A2(new_n24284_), .A3(new_n24534_), .ZN(new_n24535_));
  NOR3_X1    g24343(.A1(new_n24499_), .A2(new_n23771_), .A3(new_n24284_), .ZN(new_n24536_));
  INV_X1     g24344(.I(new_n24536_), .ZN(new_n24537_));
  AOI22_X1   g24345(.A1(new_n24537_), .A2(new_n24534_), .B1(\asqrt[1] ), .B2(new_n24535_), .ZN(new_n24538_));
  INV_X1     g24346(.I(new_n24538_), .ZN(new_n24539_));
  OAI21_X1   g24347(.A1(new_n24523_), .A2(new_n24531_), .B(new_n24527_), .ZN(new_n24540_));
  NAND2_X1   g24348(.A1(new_n24540_), .A2(new_n24539_), .ZN(new_n24541_));
  OAI21_X1   g24349(.A1(new_n24533_), .A2(new_n24541_), .B(new_n18792_), .ZN(new_n24542_));
  NOR3_X1    g24350(.A1(new_n24499_), .A2(new_n23780_), .A3(new_n23785_), .ZN(new_n24543_));
  INV_X1     g24351(.I(new_n24543_), .ZN(new_n24544_));
  NOR3_X1    g24352(.A1(new_n23780_), .A2(new_n24252_), .A3(new_n23785_), .ZN(new_n24545_));
  AOI22_X1   g24353(.A1(new_n24544_), .A2(new_n24252_), .B1(\asqrt[1] ), .B2(new_n24545_), .ZN(new_n24546_));
  OAI21_X1   g24354(.A1(\asqrt[8] ), .A2(new_n24532_), .B(new_n24540_), .ZN(new_n24547_));
  AOI21_X1   g24355(.A1(new_n24547_), .A2(new_n24538_), .B(new_n24546_), .ZN(new_n24548_));
  AOI21_X1   g24356(.A1(new_n24548_), .A2(new_n24542_), .B(\asqrt[10] ), .ZN(new_n24549_));
  AND3_X2    g24357(.A1(new_n23787_), .A2(new_n23792_), .A3(new_n24278_), .Z(new_n24550_));
  NAND3_X1   g24358(.A1(\asqrt[1] ), .A2(new_n23787_), .A3(new_n24278_), .ZN(new_n24551_));
  AOI22_X1   g24359(.A1(new_n24551_), .A2(new_n23793_), .B1(\asqrt[1] ), .B2(new_n24550_), .ZN(new_n24552_));
  INV_X1     g24360(.I(new_n24546_), .ZN(new_n24553_));
  INV_X1     g24361(.I(new_n24540_), .ZN(new_n24554_));
  OAI21_X1   g24362(.A1(new_n24533_), .A2(new_n24554_), .B(new_n24538_), .ZN(new_n24555_));
  AOI21_X1   g24363(.A1(new_n24542_), .A2(new_n24555_), .B(new_n24553_), .ZN(new_n24556_));
  NOR3_X1    g24364(.A1(new_n24549_), .A2(new_n24556_), .A3(new_n24552_), .ZN(new_n24557_));
  NOR2_X1    g24365(.A1(new_n24557_), .A2(\asqrt[11] ), .ZN(new_n24558_));
  INV_X1     g24366(.I(new_n23800_), .ZN(new_n24559_));
  NOR3_X1    g24367(.A1(new_n24499_), .A2(new_n23796_), .A3(new_n24288_), .ZN(new_n24560_));
  INV_X1     g24368(.I(new_n24560_), .ZN(new_n24561_));
  NOR3_X1    g24369(.A1(new_n23796_), .A2(new_n24288_), .A3(new_n24559_), .ZN(new_n24562_));
  AOI22_X1   g24370(.A1(new_n24561_), .A2(new_n24559_), .B1(\asqrt[1] ), .B2(new_n24562_), .ZN(new_n24563_));
  INV_X1     g24371(.I(new_n24563_), .ZN(new_n24564_));
  OAI21_X1   g24372(.A1(new_n24549_), .A2(new_n24556_), .B(new_n24552_), .ZN(new_n24565_));
  NAND2_X1   g24373(.A1(new_n24565_), .A2(new_n24564_), .ZN(new_n24566_));
  OAI21_X1   g24374(.A1(new_n24558_), .A2(new_n24566_), .B(new_n16881_), .ZN(new_n24567_));
  NOR3_X1    g24375(.A1(new_n23805_), .A2(new_n24251_), .A3(new_n23809_), .ZN(new_n24568_));
  NOR3_X1    g24376(.A1(new_n24499_), .A2(new_n23805_), .A3(new_n23809_), .ZN(new_n24569_));
  INV_X1     g24377(.I(new_n24569_), .ZN(new_n24570_));
  AOI22_X1   g24378(.A1(new_n24570_), .A2(new_n24251_), .B1(\asqrt[1] ), .B2(new_n24568_), .ZN(new_n24571_));
  OAI21_X1   g24379(.A1(\asqrt[11] ), .A2(new_n24557_), .B(new_n24565_), .ZN(new_n24572_));
  AOI21_X1   g24380(.A1(new_n24572_), .A2(new_n24563_), .B(new_n24571_), .ZN(new_n24573_));
  AOI21_X1   g24381(.A1(new_n24573_), .A2(new_n24567_), .B(\asqrt[13] ), .ZN(new_n24574_));
  NOR2_X1    g24382(.A1(new_n23810_), .A2(new_n23818_), .ZN(new_n24575_));
  NOR3_X1    g24383(.A1(new_n24499_), .A2(new_n24282_), .A3(new_n24575_), .ZN(new_n24576_));
  INV_X1     g24384(.I(new_n24576_), .ZN(new_n24577_));
  NOR3_X1    g24385(.A1(new_n24575_), .A2(new_n24282_), .A3(new_n23817_), .ZN(new_n24578_));
  AOI22_X1   g24386(.A1(new_n24577_), .A2(new_n23817_), .B1(\asqrt[1] ), .B2(new_n24578_), .ZN(new_n24579_));
  INV_X1     g24387(.I(new_n24571_), .ZN(new_n24580_));
  INV_X1     g24388(.I(new_n24565_), .ZN(new_n24581_));
  OAI21_X1   g24389(.A1(new_n24558_), .A2(new_n24581_), .B(new_n24563_), .ZN(new_n24582_));
  AOI21_X1   g24390(.A1(new_n24567_), .A2(new_n24582_), .B(new_n24580_), .ZN(new_n24583_));
  NOR3_X1    g24391(.A1(new_n24574_), .A2(new_n24583_), .A3(new_n24579_), .ZN(new_n24584_));
  NOR2_X1    g24392(.A1(new_n24584_), .A2(\asqrt[14] ), .ZN(new_n24585_));
  INV_X1     g24393(.I(new_n23824_), .ZN(new_n24586_));
  NOR3_X1    g24394(.A1(new_n23820_), .A2(new_n24296_), .A3(new_n24586_), .ZN(new_n24587_));
  NOR3_X1    g24395(.A1(new_n24499_), .A2(new_n23820_), .A3(new_n24296_), .ZN(new_n24588_));
  INV_X1     g24396(.I(new_n24588_), .ZN(new_n24589_));
  AOI22_X1   g24397(.A1(new_n24589_), .A2(new_n24586_), .B1(\asqrt[1] ), .B2(new_n24587_), .ZN(new_n24590_));
  INV_X1     g24398(.I(new_n24590_), .ZN(new_n24591_));
  OAI21_X1   g24399(.A1(new_n24574_), .A2(new_n24583_), .B(new_n24579_), .ZN(new_n24592_));
  NAND2_X1   g24400(.A1(new_n24592_), .A2(new_n24591_), .ZN(new_n24593_));
  OAI21_X1   g24401(.A1(new_n24585_), .A2(new_n24593_), .B(new_n15067_), .ZN(new_n24594_));
  NOR3_X1    g24402(.A1(new_n24499_), .A2(new_n23829_), .A3(new_n23835_), .ZN(new_n24595_));
  INV_X1     g24403(.I(new_n24595_), .ZN(new_n24596_));
  NOR3_X1    g24404(.A1(new_n23829_), .A2(new_n24250_), .A3(new_n23835_), .ZN(new_n24597_));
  AOI22_X1   g24405(.A1(new_n24596_), .A2(new_n24250_), .B1(\asqrt[1] ), .B2(new_n24597_), .ZN(new_n24598_));
  OAI21_X1   g24406(.A1(\asqrt[14] ), .A2(new_n24584_), .B(new_n24592_), .ZN(new_n24599_));
  AOI21_X1   g24407(.A1(new_n24599_), .A2(new_n24590_), .B(new_n24598_), .ZN(new_n24600_));
  AOI21_X1   g24408(.A1(new_n24600_), .A2(new_n24594_), .B(\asqrt[16] ), .ZN(new_n24601_));
  NOR2_X1    g24409(.A1(new_n23836_), .A2(new_n23844_), .ZN(new_n24602_));
  NOR3_X1    g24410(.A1(new_n24602_), .A2(new_n24295_), .A3(new_n23843_), .ZN(new_n24603_));
  NOR3_X1    g24411(.A1(new_n24499_), .A2(new_n24295_), .A3(new_n24602_), .ZN(new_n24604_));
  INV_X1     g24412(.I(new_n24604_), .ZN(new_n24605_));
  AOI22_X1   g24413(.A1(new_n24605_), .A2(new_n23843_), .B1(\asqrt[1] ), .B2(new_n24603_), .ZN(new_n24606_));
  INV_X1     g24414(.I(new_n24598_), .ZN(new_n24607_));
  INV_X1     g24415(.I(new_n24592_), .ZN(new_n24608_));
  OAI21_X1   g24416(.A1(new_n24585_), .A2(new_n24608_), .B(new_n24590_), .ZN(new_n24609_));
  AOI21_X1   g24417(.A1(new_n24594_), .A2(new_n24609_), .B(new_n24607_), .ZN(new_n24610_));
  NOR3_X1    g24418(.A1(new_n24601_), .A2(new_n24610_), .A3(new_n24606_), .ZN(new_n24611_));
  NOR2_X1    g24419(.A1(new_n24611_), .A2(\asqrt[17] ), .ZN(new_n24612_));
  INV_X1     g24420(.I(new_n23850_), .ZN(new_n24613_));
  NOR3_X1    g24421(.A1(new_n24499_), .A2(new_n23846_), .A3(new_n24304_), .ZN(new_n24614_));
  INV_X1     g24422(.I(new_n24614_), .ZN(new_n24615_));
  NOR3_X1    g24423(.A1(new_n23846_), .A2(new_n24304_), .A3(new_n24613_), .ZN(new_n24616_));
  AOI22_X1   g24424(.A1(new_n24615_), .A2(new_n24613_), .B1(\asqrt[1] ), .B2(new_n24616_), .ZN(new_n24617_));
  INV_X1     g24425(.I(new_n24617_), .ZN(new_n24618_));
  OAI21_X1   g24426(.A1(new_n24601_), .A2(new_n24610_), .B(new_n24606_), .ZN(new_n24619_));
  NAND2_X1   g24427(.A1(new_n24619_), .A2(new_n24618_), .ZN(new_n24620_));
  OAI21_X1   g24428(.A1(new_n24612_), .A2(new_n24620_), .B(new_n13353_), .ZN(new_n24621_));
  NOR3_X1    g24429(.A1(new_n23855_), .A2(new_n24249_), .A3(new_n23861_), .ZN(new_n24622_));
  NOR3_X1    g24430(.A1(new_n24499_), .A2(new_n23855_), .A3(new_n23861_), .ZN(new_n24623_));
  INV_X1     g24431(.I(new_n24623_), .ZN(new_n24624_));
  AOI22_X1   g24432(.A1(new_n24624_), .A2(new_n24249_), .B1(\asqrt[1] ), .B2(new_n24622_), .ZN(new_n24625_));
  OAI21_X1   g24433(.A1(\asqrt[17] ), .A2(new_n24611_), .B(new_n24619_), .ZN(new_n24626_));
  AOI21_X1   g24434(.A1(new_n24626_), .A2(new_n24617_), .B(new_n24625_), .ZN(new_n24627_));
  AOI21_X1   g24435(.A1(new_n24627_), .A2(new_n24621_), .B(\asqrt[19] ), .ZN(new_n24628_));
  NOR2_X1    g24436(.A1(new_n23862_), .A2(new_n23870_), .ZN(new_n24629_));
  NOR3_X1    g24437(.A1(new_n24499_), .A2(new_n24303_), .A3(new_n24629_), .ZN(new_n24630_));
  INV_X1     g24438(.I(new_n24630_), .ZN(new_n24631_));
  NOR3_X1    g24439(.A1(new_n24629_), .A2(new_n24303_), .A3(new_n23869_), .ZN(new_n24632_));
  AOI22_X1   g24440(.A1(new_n24631_), .A2(new_n23869_), .B1(\asqrt[1] ), .B2(new_n24632_), .ZN(new_n24633_));
  INV_X1     g24441(.I(new_n24625_), .ZN(new_n24634_));
  INV_X1     g24442(.I(new_n24619_), .ZN(new_n24635_));
  OAI21_X1   g24443(.A1(new_n24612_), .A2(new_n24635_), .B(new_n24617_), .ZN(new_n24636_));
  AOI21_X1   g24444(.A1(new_n24621_), .A2(new_n24636_), .B(new_n24634_), .ZN(new_n24637_));
  NOR3_X1    g24445(.A1(new_n24628_), .A2(new_n24637_), .A3(new_n24633_), .ZN(new_n24638_));
  NOR2_X1    g24446(.A1(new_n24638_), .A2(\asqrt[20] ), .ZN(new_n24639_));
  INV_X1     g24447(.I(new_n23876_), .ZN(new_n24640_));
  NOR3_X1    g24448(.A1(new_n23872_), .A2(new_n24312_), .A3(new_n24640_), .ZN(new_n24641_));
  NOR3_X1    g24449(.A1(new_n24499_), .A2(new_n23872_), .A3(new_n24312_), .ZN(new_n24642_));
  INV_X1     g24450(.I(new_n24642_), .ZN(new_n24643_));
  AOI22_X1   g24451(.A1(new_n24643_), .A2(new_n24640_), .B1(\asqrt[1] ), .B2(new_n24641_), .ZN(new_n24644_));
  INV_X1     g24452(.I(new_n24644_), .ZN(new_n24645_));
  OAI21_X1   g24453(.A1(new_n24628_), .A2(new_n24637_), .B(new_n24633_), .ZN(new_n24646_));
  NAND2_X1   g24454(.A1(new_n24646_), .A2(new_n24645_), .ZN(new_n24647_));
  OAI21_X1   g24455(.A1(new_n24639_), .A2(new_n24647_), .B(new_n11736_), .ZN(new_n24648_));
  NOR3_X1    g24456(.A1(new_n24499_), .A2(new_n23881_), .A3(new_n23887_), .ZN(new_n24649_));
  INV_X1     g24457(.I(new_n24649_), .ZN(new_n24650_));
  NOR3_X1    g24458(.A1(new_n23881_), .A2(new_n24248_), .A3(new_n23887_), .ZN(new_n24651_));
  AOI22_X1   g24459(.A1(new_n24650_), .A2(new_n24248_), .B1(\asqrt[1] ), .B2(new_n24651_), .ZN(new_n24652_));
  OAI21_X1   g24460(.A1(\asqrt[20] ), .A2(new_n24638_), .B(new_n24646_), .ZN(new_n24653_));
  AOI21_X1   g24461(.A1(new_n24653_), .A2(new_n24644_), .B(new_n24652_), .ZN(new_n24654_));
  AOI21_X1   g24462(.A1(new_n24654_), .A2(new_n24648_), .B(\asqrt[22] ), .ZN(new_n24655_));
  NOR2_X1    g24463(.A1(new_n23888_), .A2(new_n23896_), .ZN(new_n24656_));
  NOR3_X1    g24464(.A1(new_n24656_), .A2(new_n24311_), .A3(new_n23895_), .ZN(new_n24657_));
  NOR3_X1    g24465(.A1(new_n24499_), .A2(new_n24311_), .A3(new_n24656_), .ZN(new_n24658_));
  INV_X1     g24466(.I(new_n24658_), .ZN(new_n24659_));
  AOI22_X1   g24467(.A1(new_n24659_), .A2(new_n23895_), .B1(\asqrt[1] ), .B2(new_n24657_), .ZN(new_n24660_));
  INV_X1     g24468(.I(new_n24652_), .ZN(new_n24661_));
  INV_X1     g24469(.I(new_n24646_), .ZN(new_n24662_));
  OAI21_X1   g24470(.A1(new_n24639_), .A2(new_n24662_), .B(new_n24644_), .ZN(new_n24663_));
  AOI21_X1   g24471(.A1(new_n24648_), .A2(new_n24663_), .B(new_n24661_), .ZN(new_n24664_));
  NOR3_X1    g24472(.A1(new_n24655_), .A2(new_n24664_), .A3(new_n24660_), .ZN(new_n24665_));
  NOR2_X1    g24473(.A1(new_n24665_), .A2(\asqrt[23] ), .ZN(new_n24666_));
  INV_X1     g24474(.I(new_n23902_), .ZN(new_n24667_));
  NOR3_X1    g24475(.A1(new_n24499_), .A2(new_n23898_), .A3(new_n24320_), .ZN(new_n24668_));
  INV_X1     g24476(.I(new_n24668_), .ZN(new_n24669_));
  NOR3_X1    g24477(.A1(new_n23898_), .A2(new_n24320_), .A3(new_n24667_), .ZN(new_n24670_));
  AOI22_X1   g24478(.A1(new_n24669_), .A2(new_n24667_), .B1(\asqrt[1] ), .B2(new_n24670_), .ZN(new_n24671_));
  INV_X1     g24479(.I(new_n24671_), .ZN(new_n24672_));
  OAI21_X1   g24480(.A1(new_n24655_), .A2(new_n24664_), .B(new_n24660_), .ZN(new_n24673_));
  NAND2_X1   g24481(.A1(new_n24673_), .A2(new_n24672_), .ZN(new_n24674_));
  OAI21_X1   g24482(.A1(new_n24666_), .A2(new_n24674_), .B(new_n10221_), .ZN(new_n24675_));
  NOR3_X1    g24483(.A1(new_n23907_), .A2(new_n24247_), .A3(new_n23913_), .ZN(new_n24676_));
  NOR3_X1    g24484(.A1(new_n24499_), .A2(new_n23907_), .A3(new_n23913_), .ZN(new_n24677_));
  INV_X1     g24485(.I(new_n24677_), .ZN(new_n24678_));
  AOI22_X1   g24486(.A1(new_n24678_), .A2(new_n24247_), .B1(\asqrt[1] ), .B2(new_n24676_), .ZN(new_n24679_));
  OAI21_X1   g24487(.A1(\asqrt[23] ), .A2(new_n24665_), .B(new_n24673_), .ZN(new_n24680_));
  AOI21_X1   g24488(.A1(new_n24680_), .A2(new_n24671_), .B(new_n24679_), .ZN(new_n24681_));
  AOI21_X1   g24489(.A1(new_n24681_), .A2(new_n24675_), .B(\asqrt[25] ), .ZN(new_n24682_));
  NOR2_X1    g24490(.A1(new_n23914_), .A2(new_n23922_), .ZN(new_n24683_));
  NOR3_X1    g24491(.A1(new_n24499_), .A2(new_n24319_), .A3(new_n24683_), .ZN(new_n24684_));
  INV_X1     g24492(.I(new_n24684_), .ZN(new_n24685_));
  NOR3_X1    g24493(.A1(new_n24683_), .A2(new_n24319_), .A3(new_n23921_), .ZN(new_n24686_));
  AOI22_X1   g24494(.A1(new_n24685_), .A2(new_n23921_), .B1(\asqrt[1] ), .B2(new_n24686_), .ZN(new_n24687_));
  INV_X1     g24495(.I(new_n24679_), .ZN(new_n24688_));
  INV_X1     g24496(.I(new_n24673_), .ZN(new_n24689_));
  OAI21_X1   g24497(.A1(new_n24666_), .A2(new_n24689_), .B(new_n24671_), .ZN(new_n24690_));
  AOI21_X1   g24498(.A1(new_n24675_), .A2(new_n24690_), .B(new_n24688_), .ZN(new_n24691_));
  NOR3_X1    g24499(.A1(new_n24682_), .A2(new_n24691_), .A3(new_n24687_), .ZN(new_n24692_));
  NOR2_X1    g24500(.A1(new_n24692_), .A2(\asqrt[26] ), .ZN(new_n24693_));
  INV_X1     g24501(.I(new_n23928_), .ZN(new_n24694_));
  NOR3_X1    g24502(.A1(new_n23924_), .A2(new_n24328_), .A3(new_n24694_), .ZN(new_n24695_));
  NOR3_X1    g24503(.A1(new_n24499_), .A2(new_n23924_), .A3(new_n24328_), .ZN(new_n24696_));
  INV_X1     g24504(.I(new_n24696_), .ZN(new_n24697_));
  AOI22_X1   g24505(.A1(new_n24697_), .A2(new_n24694_), .B1(\asqrt[1] ), .B2(new_n24695_), .ZN(new_n24698_));
  INV_X1     g24506(.I(new_n24698_), .ZN(new_n24699_));
  OAI21_X1   g24507(.A1(new_n24682_), .A2(new_n24691_), .B(new_n24687_), .ZN(new_n24700_));
  NAND2_X1   g24508(.A1(new_n24700_), .A2(new_n24699_), .ZN(new_n24701_));
  OAI21_X1   g24509(.A1(new_n24693_), .A2(new_n24701_), .B(new_n8826_), .ZN(new_n24702_));
  NOR3_X1    g24510(.A1(new_n24499_), .A2(new_n23933_), .A3(new_n23939_), .ZN(new_n24703_));
  INV_X1     g24511(.I(new_n24703_), .ZN(new_n24704_));
  NOR3_X1    g24512(.A1(new_n23933_), .A2(new_n24246_), .A3(new_n23939_), .ZN(new_n24705_));
  AOI22_X1   g24513(.A1(new_n24704_), .A2(new_n24246_), .B1(\asqrt[1] ), .B2(new_n24705_), .ZN(new_n24706_));
  OAI21_X1   g24514(.A1(\asqrt[26] ), .A2(new_n24692_), .B(new_n24700_), .ZN(new_n24707_));
  AOI21_X1   g24515(.A1(new_n24707_), .A2(new_n24698_), .B(new_n24706_), .ZN(new_n24708_));
  AOI21_X1   g24516(.A1(new_n24708_), .A2(new_n24702_), .B(\asqrt[28] ), .ZN(new_n24709_));
  NOR2_X1    g24517(.A1(new_n23940_), .A2(new_n23948_), .ZN(new_n24710_));
  NOR3_X1    g24518(.A1(new_n24710_), .A2(new_n24327_), .A3(new_n23947_), .ZN(new_n24711_));
  NOR3_X1    g24519(.A1(new_n24499_), .A2(new_n24327_), .A3(new_n24710_), .ZN(new_n24712_));
  INV_X1     g24520(.I(new_n24712_), .ZN(new_n24713_));
  AOI22_X1   g24521(.A1(new_n24713_), .A2(new_n23947_), .B1(\asqrt[1] ), .B2(new_n24711_), .ZN(new_n24714_));
  INV_X1     g24522(.I(new_n24706_), .ZN(new_n24715_));
  INV_X1     g24523(.I(new_n24700_), .ZN(new_n24716_));
  OAI21_X1   g24524(.A1(new_n24693_), .A2(new_n24716_), .B(new_n24698_), .ZN(new_n24717_));
  AOI21_X1   g24525(.A1(new_n24702_), .A2(new_n24717_), .B(new_n24715_), .ZN(new_n24718_));
  NOR3_X1    g24526(.A1(new_n24709_), .A2(new_n24718_), .A3(new_n24714_), .ZN(new_n24719_));
  NOR2_X1    g24527(.A1(new_n24719_), .A2(\asqrt[29] ), .ZN(new_n24720_));
  INV_X1     g24528(.I(new_n23954_), .ZN(new_n24721_));
  NOR3_X1    g24529(.A1(new_n24499_), .A2(new_n23950_), .A3(new_n24336_), .ZN(new_n24722_));
  INV_X1     g24530(.I(new_n24722_), .ZN(new_n24723_));
  NOR3_X1    g24531(.A1(new_n23950_), .A2(new_n24336_), .A3(new_n24721_), .ZN(new_n24724_));
  AOI22_X1   g24532(.A1(new_n24723_), .A2(new_n24721_), .B1(\asqrt[1] ), .B2(new_n24724_), .ZN(new_n24725_));
  INV_X1     g24533(.I(new_n24725_), .ZN(new_n24726_));
  OAI21_X1   g24534(.A1(new_n24709_), .A2(new_n24718_), .B(new_n24714_), .ZN(new_n24727_));
  NAND2_X1   g24535(.A1(new_n24727_), .A2(new_n24726_), .ZN(new_n24728_));
  OAI21_X1   g24536(.A1(new_n24720_), .A2(new_n24728_), .B(new_n7539_), .ZN(new_n24729_));
  NOR3_X1    g24537(.A1(new_n23959_), .A2(new_n24245_), .A3(new_n23965_), .ZN(new_n24730_));
  NOR3_X1    g24538(.A1(new_n24499_), .A2(new_n23959_), .A3(new_n23965_), .ZN(new_n24731_));
  INV_X1     g24539(.I(new_n24731_), .ZN(new_n24732_));
  AOI22_X1   g24540(.A1(new_n24732_), .A2(new_n24245_), .B1(\asqrt[1] ), .B2(new_n24730_), .ZN(new_n24733_));
  OAI21_X1   g24541(.A1(\asqrt[29] ), .A2(new_n24719_), .B(new_n24727_), .ZN(new_n24734_));
  AOI21_X1   g24542(.A1(new_n24734_), .A2(new_n24725_), .B(new_n24733_), .ZN(new_n24735_));
  AOI21_X1   g24543(.A1(new_n24735_), .A2(new_n24729_), .B(\asqrt[31] ), .ZN(new_n24736_));
  NOR2_X1    g24544(.A1(new_n23966_), .A2(new_n23974_), .ZN(new_n24737_));
  NOR3_X1    g24545(.A1(new_n24499_), .A2(new_n24335_), .A3(new_n24737_), .ZN(new_n24738_));
  INV_X1     g24546(.I(new_n24738_), .ZN(new_n24739_));
  NOR3_X1    g24547(.A1(new_n24737_), .A2(new_n24335_), .A3(new_n23973_), .ZN(new_n24740_));
  AOI22_X1   g24548(.A1(new_n24739_), .A2(new_n23973_), .B1(\asqrt[1] ), .B2(new_n24740_), .ZN(new_n24741_));
  INV_X1     g24549(.I(new_n24733_), .ZN(new_n24742_));
  INV_X1     g24550(.I(new_n24727_), .ZN(new_n24743_));
  OAI21_X1   g24551(.A1(new_n24720_), .A2(new_n24743_), .B(new_n24725_), .ZN(new_n24744_));
  AOI21_X1   g24552(.A1(new_n24729_), .A2(new_n24744_), .B(new_n24742_), .ZN(new_n24745_));
  NOR3_X1    g24553(.A1(new_n24736_), .A2(new_n24745_), .A3(new_n24741_), .ZN(new_n24746_));
  NOR2_X1    g24554(.A1(new_n24746_), .A2(\asqrt[32] ), .ZN(new_n24747_));
  INV_X1     g24555(.I(new_n23980_), .ZN(new_n24748_));
  NOR3_X1    g24556(.A1(new_n23976_), .A2(new_n24344_), .A3(new_n24748_), .ZN(new_n24749_));
  NOR3_X1    g24557(.A1(new_n24499_), .A2(new_n23976_), .A3(new_n24344_), .ZN(new_n24750_));
  INV_X1     g24558(.I(new_n24750_), .ZN(new_n24751_));
  AOI22_X1   g24559(.A1(new_n24751_), .A2(new_n24748_), .B1(\asqrt[1] ), .B2(new_n24749_), .ZN(new_n24752_));
  INV_X1     g24560(.I(new_n24752_), .ZN(new_n24753_));
  OAI21_X1   g24561(.A1(new_n24736_), .A2(new_n24745_), .B(new_n24741_), .ZN(new_n24754_));
  NAND2_X1   g24562(.A1(new_n24754_), .A2(new_n24753_), .ZN(new_n24755_));
  OAI21_X1   g24563(.A1(new_n24747_), .A2(new_n24755_), .B(new_n6356_), .ZN(new_n24756_));
  NOR3_X1    g24564(.A1(new_n24499_), .A2(new_n23985_), .A3(new_n23991_), .ZN(new_n24757_));
  INV_X1     g24565(.I(new_n24757_), .ZN(new_n24758_));
  NOR3_X1    g24566(.A1(new_n23985_), .A2(new_n24244_), .A3(new_n23991_), .ZN(new_n24759_));
  AOI22_X1   g24567(.A1(new_n24758_), .A2(new_n24244_), .B1(\asqrt[1] ), .B2(new_n24759_), .ZN(new_n24760_));
  OAI21_X1   g24568(.A1(\asqrt[32] ), .A2(new_n24746_), .B(new_n24754_), .ZN(new_n24761_));
  AOI21_X1   g24569(.A1(new_n24761_), .A2(new_n24752_), .B(new_n24760_), .ZN(new_n24762_));
  AOI21_X1   g24570(.A1(new_n24762_), .A2(new_n24756_), .B(\asqrt[34] ), .ZN(new_n24763_));
  NOR2_X1    g24571(.A1(new_n23992_), .A2(new_n24000_), .ZN(new_n24764_));
  NOR3_X1    g24572(.A1(new_n24764_), .A2(new_n24343_), .A3(new_n23999_), .ZN(new_n24765_));
  NOR3_X1    g24573(.A1(new_n24499_), .A2(new_n24343_), .A3(new_n24764_), .ZN(new_n24766_));
  INV_X1     g24574(.I(new_n24766_), .ZN(new_n24767_));
  AOI22_X1   g24575(.A1(new_n24767_), .A2(new_n23999_), .B1(\asqrt[1] ), .B2(new_n24765_), .ZN(new_n24768_));
  INV_X1     g24576(.I(new_n24760_), .ZN(new_n24769_));
  INV_X1     g24577(.I(new_n24754_), .ZN(new_n24770_));
  OAI21_X1   g24578(.A1(new_n24747_), .A2(new_n24770_), .B(new_n24752_), .ZN(new_n24771_));
  AOI21_X1   g24579(.A1(new_n24756_), .A2(new_n24771_), .B(new_n24769_), .ZN(new_n24772_));
  NOR3_X1    g24580(.A1(new_n24763_), .A2(new_n24772_), .A3(new_n24768_), .ZN(new_n24773_));
  NOR2_X1    g24581(.A1(new_n24773_), .A2(\asqrt[35] ), .ZN(new_n24774_));
  INV_X1     g24582(.I(new_n24006_), .ZN(new_n24775_));
  NOR3_X1    g24583(.A1(new_n24499_), .A2(new_n24002_), .A3(new_n24352_), .ZN(new_n24776_));
  INV_X1     g24584(.I(new_n24776_), .ZN(new_n24777_));
  NOR3_X1    g24585(.A1(new_n24002_), .A2(new_n24352_), .A3(new_n24775_), .ZN(new_n24778_));
  AOI22_X1   g24586(.A1(new_n24777_), .A2(new_n24775_), .B1(\asqrt[1] ), .B2(new_n24778_), .ZN(new_n24779_));
  INV_X1     g24587(.I(new_n24779_), .ZN(new_n24780_));
  OAI21_X1   g24588(.A1(new_n24763_), .A2(new_n24772_), .B(new_n24768_), .ZN(new_n24781_));
  NAND2_X1   g24589(.A1(new_n24781_), .A2(new_n24780_), .ZN(new_n24782_));
  OAI21_X1   g24590(.A1(new_n24774_), .A2(new_n24782_), .B(new_n5277_), .ZN(new_n24783_));
  NOR3_X1    g24591(.A1(new_n24011_), .A2(new_n24243_), .A3(new_n24017_), .ZN(new_n24784_));
  NOR3_X1    g24592(.A1(new_n24499_), .A2(new_n24011_), .A3(new_n24017_), .ZN(new_n24785_));
  INV_X1     g24593(.I(new_n24785_), .ZN(new_n24786_));
  AOI22_X1   g24594(.A1(new_n24786_), .A2(new_n24243_), .B1(\asqrt[1] ), .B2(new_n24784_), .ZN(new_n24787_));
  OAI21_X1   g24595(.A1(\asqrt[35] ), .A2(new_n24773_), .B(new_n24781_), .ZN(new_n24788_));
  AOI21_X1   g24596(.A1(new_n24788_), .A2(new_n24779_), .B(new_n24787_), .ZN(new_n24789_));
  AOI21_X1   g24597(.A1(new_n24789_), .A2(new_n24783_), .B(\asqrt[37] ), .ZN(new_n24790_));
  NOR2_X1    g24598(.A1(new_n24018_), .A2(new_n24026_), .ZN(new_n24791_));
  NOR3_X1    g24599(.A1(new_n24499_), .A2(new_n24351_), .A3(new_n24791_), .ZN(new_n24792_));
  INV_X1     g24600(.I(new_n24792_), .ZN(new_n24793_));
  NOR3_X1    g24601(.A1(new_n24791_), .A2(new_n24351_), .A3(new_n24025_), .ZN(new_n24794_));
  AOI22_X1   g24602(.A1(new_n24793_), .A2(new_n24025_), .B1(\asqrt[1] ), .B2(new_n24794_), .ZN(new_n24795_));
  INV_X1     g24603(.I(new_n24787_), .ZN(new_n24796_));
  INV_X1     g24604(.I(new_n24781_), .ZN(new_n24797_));
  OAI21_X1   g24605(.A1(new_n24774_), .A2(new_n24797_), .B(new_n24779_), .ZN(new_n24798_));
  AOI21_X1   g24606(.A1(new_n24783_), .A2(new_n24798_), .B(new_n24796_), .ZN(new_n24799_));
  NOR3_X1    g24607(.A1(new_n24790_), .A2(new_n24799_), .A3(new_n24795_), .ZN(new_n24800_));
  NOR2_X1    g24608(.A1(new_n24800_), .A2(\asqrt[38] ), .ZN(new_n24801_));
  INV_X1     g24609(.I(new_n24032_), .ZN(new_n24802_));
  NOR3_X1    g24610(.A1(new_n24028_), .A2(new_n24360_), .A3(new_n24802_), .ZN(new_n24803_));
  NOR3_X1    g24611(.A1(new_n24499_), .A2(new_n24028_), .A3(new_n24360_), .ZN(new_n24804_));
  INV_X1     g24612(.I(new_n24804_), .ZN(new_n24805_));
  AOI22_X1   g24613(.A1(new_n24805_), .A2(new_n24802_), .B1(\asqrt[1] ), .B2(new_n24803_), .ZN(new_n24806_));
  INV_X1     g24614(.I(new_n24806_), .ZN(new_n24807_));
  OAI21_X1   g24615(.A1(new_n24790_), .A2(new_n24799_), .B(new_n24795_), .ZN(new_n24808_));
  NAND2_X1   g24616(.A1(new_n24808_), .A2(new_n24807_), .ZN(new_n24809_));
  OAI21_X1   g24617(.A1(new_n24801_), .A2(new_n24809_), .B(new_n4298_), .ZN(new_n24810_));
  NOR3_X1    g24618(.A1(new_n24499_), .A2(new_n24037_), .A3(new_n24043_), .ZN(new_n24811_));
  INV_X1     g24619(.I(new_n24811_), .ZN(new_n24812_));
  NOR3_X1    g24620(.A1(new_n24037_), .A2(new_n24242_), .A3(new_n24043_), .ZN(new_n24813_));
  AOI22_X1   g24621(.A1(new_n24812_), .A2(new_n24242_), .B1(\asqrt[1] ), .B2(new_n24813_), .ZN(new_n24814_));
  OAI21_X1   g24622(.A1(\asqrt[38] ), .A2(new_n24800_), .B(new_n24808_), .ZN(new_n24815_));
  AOI21_X1   g24623(.A1(new_n24815_), .A2(new_n24806_), .B(new_n24814_), .ZN(new_n24816_));
  AOI21_X1   g24624(.A1(new_n24816_), .A2(new_n24810_), .B(\asqrt[40] ), .ZN(new_n24817_));
  NOR2_X1    g24625(.A1(new_n24044_), .A2(new_n24052_), .ZN(new_n24818_));
  NOR3_X1    g24626(.A1(new_n24818_), .A2(new_n24359_), .A3(new_n24051_), .ZN(new_n24819_));
  NOR3_X1    g24627(.A1(new_n24499_), .A2(new_n24359_), .A3(new_n24818_), .ZN(new_n24820_));
  INV_X1     g24628(.I(new_n24820_), .ZN(new_n24821_));
  AOI22_X1   g24629(.A1(new_n24821_), .A2(new_n24051_), .B1(\asqrt[1] ), .B2(new_n24819_), .ZN(new_n24822_));
  INV_X1     g24630(.I(new_n24814_), .ZN(new_n24823_));
  INV_X1     g24631(.I(new_n24808_), .ZN(new_n24824_));
  OAI21_X1   g24632(.A1(new_n24801_), .A2(new_n24824_), .B(new_n24806_), .ZN(new_n24825_));
  AOI21_X1   g24633(.A1(new_n24810_), .A2(new_n24825_), .B(new_n24823_), .ZN(new_n24826_));
  NOR3_X1    g24634(.A1(new_n24817_), .A2(new_n24826_), .A3(new_n24822_), .ZN(new_n24827_));
  NOR2_X1    g24635(.A1(new_n24827_), .A2(\asqrt[41] ), .ZN(new_n24828_));
  INV_X1     g24636(.I(new_n24058_), .ZN(new_n24829_));
  NOR3_X1    g24637(.A1(new_n24499_), .A2(new_n24054_), .A3(new_n24368_), .ZN(new_n24830_));
  INV_X1     g24638(.I(new_n24830_), .ZN(new_n24831_));
  NOR3_X1    g24639(.A1(new_n24054_), .A2(new_n24368_), .A3(new_n24829_), .ZN(new_n24832_));
  AOI22_X1   g24640(.A1(new_n24831_), .A2(new_n24829_), .B1(\asqrt[1] ), .B2(new_n24832_), .ZN(new_n24833_));
  INV_X1     g24641(.I(new_n24833_), .ZN(new_n24834_));
  OAI21_X1   g24642(.A1(new_n24817_), .A2(new_n24826_), .B(new_n24822_), .ZN(new_n24835_));
  NAND2_X1   g24643(.A1(new_n24835_), .A2(new_n24834_), .ZN(new_n24836_));
  OAI21_X1   g24644(.A1(new_n24828_), .A2(new_n24836_), .B(new_n3419_), .ZN(new_n24837_));
  NOR3_X1    g24645(.A1(new_n24063_), .A2(new_n24241_), .A3(new_n24069_), .ZN(new_n24838_));
  NOR3_X1    g24646(.A1(new_n24499_), .A2(new_n24063_), .A3(new_n24069_), .ZN(new_n24839_));
  INV_X1     g24647(.I(new_n24839_), .ZN(new_n24840_));
  AOI22_X1   g24648(.A1(new_n24840_), .A2(new_n24241_), .B1(\asqrt[1] ), .B2(new_n24838_), .ZN(new_n24841_));
  OAI21_X1   g24649(.A1(\asqrt[41] ), .A2(new_n24827_), .B(new_n24835_), .ZN(new_n24842_));
  AOI21_X1   g24650(.A1(new_n24842_), .A2(new_n24833_), .B(new_n24841_), .ZN(new_n24843_));
  AOI21_X1   g24651(.A1(new_n24843_), .A2(new_n24837_), .B(\asqrt[43] ), .ZN(new_n24844_));
  NOR2_X1    g24652(.A1(new_n24070_), .A2(new_n24078_), .ZN(new_n24845_));
  NOR3_X1    g24653(.A1(new_n24499_), .A2(new_n24367_), .A3(new_n24845_), .ZN(new_n24846_));
  INV_X1     g24654(.I(new_n24846_), .ZN(new_n24847_));
  NOR3_X1    g24655(.A1(new_n24845_), .A2(new_n24367_), .A3(new_n24077_), .ZN(new_n24848_));
  AOI22_X1   g24656(.A1(new_n24847_), .A2(new_n24077_), .B1(\asqrt[1] ), .B2(new_n24848_), .ZN(new_n24849_));
  INV_X1     g24657(.I(new_n24841_), .ZN(new_n24850_));
  INV_X1     g24658(.I(new_n24835_), .ZN(new_n24851_));
  OAI21_X1   g24659(.A1(new_n24828_), .A2(new_n24851_), .B(new_n24833_), .ZN(new_n24852_));
  AOI21_X1   g24660(.A1(new_n24837_), .A2(new_n24852_), .B(new_n24850_), .ZN(new_n24853_));
  NOR3_X1    g24661(.A1(new_n24844_), .A2(new_n24853_), .A3(new_n24849_), .ZN(new_n24854_));
  NOR2_X1    g24662(.A1(new_n24854_), .A2(\asqrt[44] ), .ZN(new_n24855_));
  INV_X1     g24663(.I(new_n24084_), .ZN(new_n24856_));
  NOR3_X1    g24664(.A1(new_n24080_), .A2(new_n24376_), .A3(new_n24856_), .ZN(new_n24857_));
  NOR3_X1    g24665(.A1(new_n24499_), .A2(new_n24080_), .A3(new_n24376_), .ZN(new_n24858_));
  INV_X1     g24666(.I(new_n24858_), .ZN(new_n24859_));
  AOI22_X1   g24667(.A1(new_n24859_), .A2(new_n24856_), .B1(\asqrt[1] ), .B2(new_n24857_), .ZN(new_n24860_));
  INV_X1     g24668(.I(new_n24860_), .ZN(new_n24861_));
  OAI21_X1   g24669(.A1(new_n24844_), .A2(new_n24853_), .B(new_n24849_), .ZN(new_n24862_));
  NAND2_X1   g24670(.A1(new_n24862_), .A2(new_n24861_), .ZN(new_n24863_));
  OAI21_X1   g24671(.A1(new_n24855_), .A2(new_n24863_), .B(new_n2641_), .ZN(new_n24864_));
  NOR3_X1    g24672(.A1(new_n24499_), .A2(new_n24089_), .A3(new_n24095_), .ZN(new_n24865_));
  INV_X1     g24673(.I(new_n24865_), .ZN(new_n24866_));
  NOR3_X1    g24674(.A1(new_n24089_), .A2(new_n24240_), .A3(new_n24095_), .ZN(new_n24867_));
  AOI22_X1   g24675(.A1(new_n24866_), .A2(new_n24240_), .B1(\asqrt[1] ), .B2(new_n24867_), .ZN(new_n24868_));
  OAI21_X1   g24676(.A1(\asqrt[44] ), .A2(new_n24854_), .B(new_n24862_), .ZN(new_n24869_));
  AOI21_X1   g24677(.A1(new_n24869_), .A2(new_n24860_), .B(new_n24868_), .ZN(new_n24870_));
  AOI21_X1   g24678(.A1(new_n24870_), .A2(new_n24864_), .B(\asqrt[46] ), .ZN(new_n24871_));
  NOR2_X1    g24679(.A1(new_n24096_), .A2(new_n24104_), .ZN(new_n24872_));
  NOR3_X1    g24680(.A1(new_n24872_), .A2(new_n24375_), .A3(new_n24103_), .ZN(new_n24873_));
  NOR3_X1    g24681(.A1(new_n24499_), .A2(new_n24375_), .A3(new_n24872_), .ZN(new_n24874_));
  INV_X1     g24682(.I(new_n24874_), .ZN(new_n24875_));
  AOI22_X1   g24683(.A1(new_n24875_), .A2(new_n24103_), .B1(\asqrt[1] ), .B2(new_n24873_), .ZN(new_n24876_));
  INV_X1     g24684(.I(new_n24868_), .ZN(new_n24877_));
  INV_X1     g24685(.I(new_n24862_), .ZN(new_n24878_));
  OAI21_X1   g24686(.A1(new_n24855_), .A2(new_n24878_), .B(new_n24860_), .ZN(new_n24879_));
  AOI21_X1   g24687(.A1(new_n24864_), .A2(new_n24879_), .B(new_n24877_), .ZN(new_n24880_));
  NOR3_X1    g24688(.A1(new_n24871_), .A2(new_n24880_), .A3(new_n24876_), .ZN(new_n24881_));
  NOR2_X1    g24689(.A1(new_n24881_), .A2(\asqrt[47] ), .ZN(new_n24882_));
  INV_X1     g24690(.I(new_n24110_), .ZN(new_n24883_));
  NOR3_X1    g24691(.A1(new_n24499_), .A2(new_n24106_), .A3(new_n24384_), .ZN(new_n24884_));
  INV_X1     g24692(.I(new_n24884_), .ZN(new_n24885_));
  NOR3_X1    g24693(.A1(new_n24106_), .A2(new_n24384_), .A3(new_n24883_), .ZN(new_n24886_));
  AOI22_X1   g24694(.A1(new_n24885_), .A2(new_n24883_), .B1(\asqrt[1] ), .B2(new_n24886_), .ZN(new_n24887_));
  INV_X1     g24695(.I(new_n24887_), .ZN(new_n24888_));
  OAI21_X1   g24696(.A1(new_n24871_), .A2(new_n24880_), .B(new_n24876_), .ZN(new_n24889_));
  NAND2_X1   g24697(.A1(new_n24889_), .A2(new_n24888_), .ZN(new_n24890_));
  OAI21_X1   g24698(.A1(new_n24882_), .A2(new_n24890_), .B(new_n1956_), .ZN(new_n24891_));
  NOR3_X1    g24699(.A1(new_n24115_), .A2(new_n24239_), .A3(new_n24121_), .ZN(new_n24892_));
  NOR3_X1    g24700(.A1(new_n24499_), .A2(new_n24115_), .A3(new_n24121_), .ZN(new_n24893_));
  INV_X1     g24701(.I(new_n24893_), .ZN(new_n24894_));
  AOI22_X1   g24702(.A1(new_n24894_), .A2(new_n24239_), .B1(\asqrt[1] ), .B2(new_n24892_), .ZN(new_n24895_));
  OAI21_X1   g24703(.A1(\asqrt[47] ), .A2(new_n24881_), .B(new_n24889_), .ZN(new_n24896_));
  AOI21_X1   g24704(.A1(new_n24896_), .A2(new_n24887_), .B(new_n24895_), .ZN(new_n24897_));
  AOI21_X1   g24705(.A1(new_n24897_), .A2(new_n24891_), .B(\asqrt[49] ), .ZN(new_n24898_));
  NOR2_X1    g24706(.A1(new_n24122_), .A2(new_n24130_), .ZN(new_n24899_));
  NOR3_X1    g24707(.A1(new_n24499_), .A2(new_n24383_), .A3(new_n24899_), .ZN(new_n24900_));
  INV_X1     g24708(.I(new_n24900_), .ZN(new_n24901_));
  NOR3_X1    g24709(.A1(new_n24899_), .A2(new_n24383_), .A3(new_n24129_), .ZN(new_n24902_));
  AOI22_X1   g24710(.A1(new_n24901_), .A2(new_n24129_), .B1(\asqrt[1] ), .B2(new_n24902_), .ZN(new_n24903_));
  INV_X1     g24711(.I(new_n24895_), .ZN(new_n24904_));
  INV_X1     g24712(.I(new_n24889_), .ZN(new_n24905_));
  OAI21_X1   g24713(.A1(new_n24882_), .A2(new_n24905_), .B(new_n24887_), .ZN(new_n24906_));
  AOI21_X1   g24714(.A1(new_n24891_), .A2(new_n24906_), .B(new_n24904_), .ZN(new_n24907_));
  NOR3_X1    g24715(.A1(new_n24898_), .A2(new_n24907_), .A3(new_n24903_), .ZN(new_n24908_));
  NOR2_X1    g24716(.A1(new_n24908_), .A2(\asqrt[50] ), .ZN(new_n24909_));
  INV_X1     g24717(.I(new_n24136_), .ZN(new_n24910_));
  NOR3_X1    g24718(.A1(new_n24132_), .A2(new_n24392_), .A3(new_n24910_), .ZN(new_n24911_));
  NOR3_X1    g24719(.A1(new_n24499_), .A2(new_n24132_), .A3(new_n24392_), .ZN(new_n24912_));
  INV_X1     g24720(.I(new_n24912_), .ZN(new_n24913_));
  AOI22_X1   g24721(.A1(new_n24913_), .A2(new_n24910_), .B1(\asqrt[1] ), .B2(new_n24911_), .ZN(new_n24914_));
  INV_X1     g24722(.I(new_n24914_), .ZN(new_n24915_));
  OAI21_X1   g24723(.A1(new_n24898_), .A2(new_n24907_), .B(new_n24903_), .ZN(new_n24916_));
  NAND2_X1   g24724(.A1(new_n24916_), .A2(new_n24915_), .ZN(new_n24917_));
  OAI21_X1   g24725(.A1(new_n24909_), .A2(new_n24917_), .B(new_n1376_), .ZN(new_n24918_));
  NOR3_X1    g24726(.A1(new_n24499_), .A2(new_n24141_), .A3(new_n24147_), .ZN(new_n24919_));
  INV_X1     g24727(.I(new_n24919_), .ZN(new_n24920_));
  NOR3_X1    g24728(.A1(new_n24141_), .A2(new_n24238_), .A3(new_n24147_), .ZN(new_n24921_));
  AOI22_X1   g24729(.A1(new_n24920_), .A2(new_n24238_), .B1(\asqrt[1] ), .B2(new_n24921_), .ZN(new_n24922_));
  OAI21_X1   g24730(.A1(\asqrt[50] ), .A2(new_n24908_), .B(new_n24916_), .ZN(new_n24923_));
  AOI21_X1   g24731(.A1(new_n24923_), .A2(new_n24914_), .B(new_n24922_), .ZN(new_n24924_));
  AOI21_X1   g24732(.A1(new_n24924_), .A2(new_n24918_), .B(\asqrt[52] ), .ZN(new_n24925_));
  NOR2_X1    g24733(.A1(new_n24148_), .A2(new_n24158_), .ZN(new_n24926_));
  NOR3_X1    g24734(.A1(new_n24926_), .A2(new_n24391_), .A3(new_n24157_), .ZN(new_n24927_));
  NOR3_X1    g24735(.A1(new_n24499_), .A2(new_n24391_), .A3(new_n24926_), .ZN(new_n24928_));
  INV_X1     g24736(.I(new_n24928_), .ZN(new_n24929_));
  AOI22_X1   g24737(.A1(new_n24929_), .A2(new_n24157_), .B1(\asqrt[1] ), .B2(new_n24927_), .ZN(new_n24930_));
  INV_X1     g24738(.I(new_n24922_), .ZN(new_n24931_));
  INV_X1     g24739(.I(new_n24916_), .ZN(new_n24932_));
  OAI21_X1   g24740(.A1(new_n24909_), .A2(new_n24932_), .B(new_n24914_), .ZN(new_n24933_));
  AOI21_X1   g24741(.A1(new_n24918_), .A2(new_n24933_), .B(new_n24931_), .ZN(new_n24934_));
  NOR3_X1    g24742(.A1(new_n24925_), .A2(new_n24934_), .A3(new_n24930_), .ZN(new_n24935_));
  NOR2_X1    g24743(.A1(new_n24935_), .A2(\asqrt[53] ), .ZN(new_n24936_));
  INV_X1     g24744(.I(new_n24164_), .ZN(new_n24937_));
  NOR3_X1    g24745(.A1(new_n24499_), .A2(new_n24160_), .A3(new_n24400_), .ZN(new_n24938_));
  INV_X1     g24746(.I(new_n24938_), .ZN(new_n24939_));
  NOR3_X1    g24747(.A1(new_n24160_), .A2(new_n24400_), .A3(new_n24937_), .ZN(new_n24940_));
  AOI22_X1   g24748(.A1(new_n24939_), .A2(new_n24937_), .B1(\asqrt[1] ), .B2(new_n24940_), .ZN(new_n24941_));
  INV_X1     g24749(.I(new_n24941_), .ZN(new_n24942_));
  OAI21_X1   g24750(.A1(new_n24925_), .A2(new_n24934_), .B(new_n24930_), .ZN(new_n24943_));
  NAND2_X1   g24751(.A1(new_n24943_), .A2(new_n24942_), .ZN(new_n24944_));
  OAI21_X1   g24752(.A1(new_n24936_), .A2(new_n24944_), .B(new_n904_), .ZN(new_n24945_));
  NOR3_X1    g24753(.A1(new_n24169_), .A2(new_n24237_), .A3(new_n24176_), .ZN(new_n24946_));
  NOR3_X1    g24754(.A1(new_n24499_), .A2(new_n24169_), .A3(new_n24176_), .ZN(new_n24947_));
  INV_X1     g24755(.I(new_n24947_), .ZN(new_n24948_));
  AOI22_X1   g24756(.A1(new_n24948_), .A2(new_n24237_), .B1(\asqrt[1] ), .B2(new_n24946_), .ZN(new_n24949_));
  OAI21_X1   g24757(.A1(\asqrt[53] ), .A2(new_n24935_), .B(new_n24943_), .ZN(new_n24950_));
  AOI21_X1   g24758(.A1(new_n24950_), .A2(new_n24941_), .B(new_n24949_), .ZN(new_n24951_));
  AOI21_X1   g24759(.A1(new_n24951_), .A2(new_n24945_), .B(\asqrt[55] ), .ZN(new_n24952_));
  NOR2_X1    g24760(.A1(new_n24177_), .A2(new_n24188_), .ZN(new_n24953_));
  NOR3_X1    g24761(.A1(new_n24499_), .A2(new_n24399_), .A3(new_n24953_), .ZN(new_n24954_));
  INV_X1     g24762(.I(new_n24954_), .ZN(new_n24955_));
  NOR3_X1    g24763(.A1(new_n24953_), .A2(new_n24399_), .A3(new_n24187_), .ZN(new_n24956_));
  AOI22_X1   g24764(.A1(new_n24955_), .A2(new_n24187_), .B1(\asqrt[1] ), .B2(new_n24956_), .ZN(new_n24957_));
  INV_X1     g24765(.I(new_n24949_), .ZN(new_n24958_));
  INV_X1     g24766(.I(new_n24943_), .ZN(new_n24959_));
  OAI21_X1   g24767(.A1(new_n24936_), .A2(new_n24959_), .B(new_n24941_), .ZN(new_n24960_));
  AOI21_X1   g24768(.A1(new_n24945_), .A2(new_n24960_), .B(new_n24958_), .ZN(new_n24961_));
  NOR3_X1    g24769(.A1(new_n24952_), .A2(new_n24961_), .A3(new_n24957_), .ZN(new_n24962_));
  NOR2_X1    g24770(.A1(new_n24962_), .A2(\asqrt[56] ), .ZN(new_n24963_));
  INV_X1     g24771(.I(new_n24194_), .ZN(new_n24964_));
  NOR3_X1    g24772(.A1(new_n24190_), .A2(new_n24408_), .A3(new_n24964_), .ZN(new_n24965_));
  NOR3_X1    g24773(.A1(new_n24499_), .A2(new_n24190_), .A3(new_n24408_), .ZN(new_n24966_));
  INV_X1     g24774(.I(new_n24966_), .ZN(new_n24967_));
  AOI22_X1   g24775(.A1(new_n24967_), .A2(new_n24964_), .B1(\asqrt[1] ), .B2(new_n24965_), .ZN(new_n24968_));
  INV_X1     g24776(.I(new_n24968_), .ZN(new_n24969_));
  OAI21_X1   g24777(.A1(new_n24952_), .A2(new_n24961_), .B(new_n24957_), .ZN(new_n24970_));
  NAND2_X1   g24778(.A1(new_n24970_), .A2(new_n24969_), .ZN(new_n24971_));
  OAI21_X1   g24779(.A1(new_n24963_), .A2(new_n24971_), .B(new_n531_), .ZN(new_n24972_));
  NOR3_X1    g24780(.A1(new_n24499_), .A2(new_n24199_), .A3(new_n24206_), .ZN(new_n24973_));
  INV_X1     g24781(.I(new_n24973_), .ZN(new_n24974_));
  NOR3_X1    g24782(.A1(new_n24199_), .A2(new_n24236_), .A3(new_n24206_), .ZN(new_n24975_));
  AOI22_X1   g24783(.A1(new_n24974_), .A2(new_n24236_), .B1(\asqrt[1] ), .B2(new_n24975_), .ZN(new_n24976_));
  OAI21_X1   g24784(.A1(\asqrt[56] ), .A2(new_n24962_), .B(new_n24970_), .ZN(new_n24977_));
  AOI21_X1   g24785(.A1(new_n24977_), .A2(new_n24968_), .B(new_n24976_), .ZN(new_n24978_));
  NAND2_X1   g24786(.A1(new_n24978_), .A2(new_n24972_), .ZN(new_n24979_));
  NAND2_X1   g24787(.A1(new_n24979_), .A2(new_n436_), .ZN(new_n24980_));
  NOR2_X1    g24788(.A1(new_n24207_), .A2(new_n24219_), .ZN(new_n24981_));
  NOR3_X1    g24789(.A1(new_n24981_), .A2(new_n24407_), .A3(new_n24218_), .ZN(new_n24982_));
  NOR3_X1    g24790(.A1(new_n24499_), .A2(new_n24407_), .A3(new_n24981_), .ZN(new_n24983_));
  INV_X1     g24791(.I(new_n24983_), .ZN(new_n24984_));
  AOI22_X1   g24792(.A1(new_n24984_), .A2(new_n24218_), .B1(\asqrt[1] ), .B2(new_n24982_), .ZN(new_n24985_));
  INV_X1     g24793(.I(new_n24976_), .ZN(new_n24986_));
  INV_X1     g24794(.I(new_n24970_), .ZN(new_n24987_));
  OAI21_X1   g24795(.A1(new_n24963_), .A2(new_n24987_), .B(new_n24968_), .ZN(new_n24988_));
  AOI21_X1   g24796(.A1(new_n24972_), .A2(new_n24988_), .B(new_n24986_), .ZN(new_n24989_));
  NOR2_X1    g24797(.A1(new_n24989_), .A2(new_n24985_), .ZN(new_n24990_));
  NAND2_X1   g24798(.A1(new_n24980_), .A2(new_n24990_), .ZN(new_n24991_));
  NAND2_X1   g24799(.A1(new_n24991_), .A2(new_n327_), .ZN(new_n24992_));
  INV_X1     g24800(.I(new_n24225_), .ZN(new_n24993_));
  NOR3_X1    g24801(.A1(new_n24499_), .A2(new_n24221_), .A3(new_n24420_), .ZN(new_n24994_));
  INV_X1     g24802(.I(new_n24994_), .ZN(new_n24995_));
  NOR3_X1    g24803(.A1(new_n24221_), .A2(new_n24420_), .A3(new_n24993_), .ZN(new_n24996_));
  AOI22_X1   g24804(.A1(new_n24995_), .A2(new_n24993_), .B1(\asqrt[1] ), .B2(new_n24996_), .ZN(new_n24997_));
  INV_X1     g24805(.I(new_n24997_), .ZN(new_n24998_));
  AOI21_X1   g24806(.A1(new_n24978_), .A2(new_n24972_), .B(\asqrt[58] ), .ZN(new_n24999_));
  OAI21_X1   g24807(.A1(new_n24999_), .A2(new_n24989_), .B(new_n24985_), .ZN(new_n25000_));
  NAND2_X1   g24808(.A1(new_n25000_), .A2(new_n24998_), .ZN(new_n25001_));
  INV_X1     g24809(.I(new_n25001_), .ZN(new_n25002_));
  AOI21_X1   g24810(.A1(new_n25002_), .A2(new_n24992_), .B(\asqrt[60] ), .ZN(new_n25003_));
  NOR3_X1    g24811(.A1(new_n24456_), .A2(new_n24235_), .A3(new_n24442_), .ZN(new_n25004_));
  NOR3_X1    g24812(.A1(new_n24499_), .A2(new_n24456_), .A3(new_n24442_), .ZN(new_n25005_));
  INV_X1     g24813(.I(new_n25005_), .ZN(new_n25006_));
  AOI22_X1   g24814(.A1(new_n25006_), .A2(new_n24235_), .B1(\asqrt[1] ), .B2(new_n25004_), .ZN(new_n25007_));
  INV_X1     g24815(.I(new_n25007_), .ZN(new_n25008_));
  AOI21_X1   g24816(.A1(new_n24980_), .A2(new_n24990_), .B(\asqrt[59] ), .ZN(new_n25009_));
  INV_X1     g24817(.I(new_n25000_), .ZN(new_n25010_));
  OAI21_X1   g24818(.A1(new_n25009_), .A2(new_n25010_), .B(new_n24997_), .ZN(new_n25011_));
  NAND2_X1   g24819(.A1(new_n25011_), .A2(new_n25008_), .ZN(new_n25012_));
  OAI21_X1   g24820(.A1(new_n25012_), .A2(new_n25003_), .B(new_n218_), .ZN(new_n25013_));
  NOR2_X1    g24821(.A1(new_n24443_), .A2(new_n24445_), .ZN(new_n25014_));
  NOR3_X1    g24822(.A1(new_n24499_), .A2(new_n24415_), .A3(new_n25014_), .ZN(new_n25015_));
  INV_X1     g24823(.I(new_n25015_), .ZN(new_n25016_));
  NOR3_X1    g24824(.A1(new_n25014_), .A2(new_n24415_), .A3(new_n24444_), .ZN(new_n25017_));
  AOI22_X1   g24825(.A1(new_n25016_), .A2(new_n24444_), .B1(\asqrt[1] ), .B2(new_n25017_), .ZN(new_n25018_));
  OAI21_X1   g24826(.A1(new_n25001_), .A2(new_n25009_), .B(new_n306_), .ZN(new_n25019_));
  AOI21_X1   g24827(.A1(new_n25019_), .A2(new_n25011_), .B(new_n25008_), .ZN(new_n25020_));
  NOR2_X1    g24828(.A1(new_n25020_), .A2(new_n25018_), .ZN(new_n25021_));
  AOI21_X1   g24829(.A1(new_n25021_), .A2(new_n25013_), .B(\asqrt[62] ), .ZN(new_n25022_));
  NOR3_X1    g24830(.A1(new_n24999_), .A2(new_n24989_), .A3(new_n24985_), .ZN(new_n25023_));
  OAI21_X1   g24831(.A1(\asqrt[59] ), .A2(new_n25023_), .B(new_n25000_), .ZN(new_n25024_));
  AOI21_X1   g24832(.A1(new_n25024_), .A2(new_n24997_), .B(new_n25007_), .ZN(new_n25025_));
  AOI21_X1   g24833(.A1(new_n25025_), .A2(new_n25019_), .B(\asqrt[61] ), .ZN(new_n25026_));
  OAI21_X1   g24834(.A1(new_n25026_), .A2(new_n25020_), .B(new_n25018_), .ZN(new_n25027_));
  NOR4_X1    g24835(.A1(new_n24499_), .A2(new_n24458_), .A3(new_n24461_), .A4(new_n24429_), .ZN(new_n25028_));
  OR3_X2     g24836(.A1(new_n24499_), .A2(new_n24458_), .A3(new_n24429_), .Z(new_n25029_));
  AOI21_X1   g24837(.A1(new_n25029_), .A2(new_n24461_), .B(new_n25028_), .ZN(new_n25030_));
  AOI21_X1   g24838(.A1(new_n24463_), .A2(new_n24424_), .B(new_n24436_), .ZN(new_n25031_));
  NAND2_X1   g24839(.A1(\asqrt[1] ), .A2(new_n25031_), .ZN(new_n25032_));
  NAND2_X1   g24840(.A1(new_n25032_), .A2(new_n24465_), .ZN(new_n25033_));
  NOR2_X1    g24841(.A1(new_n25030_), .A2(new_n25033_), .ZN(new_n25034_));
  NAND2_X1   g24842(.A1(new_n25027_), .A2(new_n25034_), .ZN(new_n25035_));
  OAI21_X1   g24843(.A1(new_n25035_), .A2(new_n25022_), .B(new_n193_), .ZN(new_n25036_));
  INV_X1     g24844(.I(new_n25018_), .ZN(new_n25037_));
  NAND2_X1   g24845(.A1(new_n25019_), .A2(new_n25011_), .ZN(new_n25038_));
  NAND2_X1   g24846(.A1(new_n25038_), .A2(new_n25007_), .ZN(new_n25039_));
  AOI21_X1   g24847(.A1(new_n25013_), .A2(new_n25039_), .B(new_n25037_), .ZN(new_n25040_));
  OAI21_X1   g24848(.A1(new_n25022_), .A2(new_n25040_), .B(new_n25030_), .ZN(new_n25041_));
  NOR2_X1    g24849(.A1(new_n24499_), .A2(new_n24436_), .ZN(new_n25042_));
  NOR2_X1    g24850(.A1(new_n25031_), .A2(new_n193_), .ZN(new_n25043_));
  OAI21_X1   g24851(.A1(new_n25042_), .A2(new_n24430_), .B(new_n25043_), .ZN(new_n25044_));
  NAND3_X1   g24852(.A1(new_n25036_), .A2(new_n25041_), .A3(new_n25044_), .ZN(\asqrt[0] ));
endmodule


