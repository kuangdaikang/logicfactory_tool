// Benchmark "voter" written by ABC on Fri Sep 15 11:27:45 2023

module voter ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] ,
    \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] ,
    \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] ,
    \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
    \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] ,
    \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] ,
    \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] ,
    \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] ,
    \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] ,
    \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
    \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] ,
    \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] ,
    \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] ,
    \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] ,
    \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] ,
    \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
    \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] ,
    \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] ,
    \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] ,
    \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] ,
    \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] ,
    \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
    \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] ,
    \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] ,
    \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] ,
    \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] ,
    \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] ,
    \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
    \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] ,
    \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] ,
    \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] ,
    \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] ,
    \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] ,
    \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
    \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] ,
    \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] ,
    \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] ,
    \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] ,
    \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] ,
    \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
    \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] ,
    \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] ,
    \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] ,
    \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] ,
    \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] ,
    \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
    \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] ,
    \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] ,
    \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] ,
    \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] ,
    \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] ,
    \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
    \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] ,
    \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] ,
    \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] ,
    \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] ,
    \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] ,
    \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
    \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] ,
    \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] ,
    \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] ,
    \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] ,
    \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] ,
    \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
    \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] ,
    \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] ,
    \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] ,
    \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] ,
    \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] ,
    \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
    \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] ,
    \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] ,
    \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] ,
    \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] ,
    \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] ,
    \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
    \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] ,
    \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] ,
    \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] ,
    \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] ,
    \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] ,
    \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
    \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] ,
    \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] ,
    \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] ,
    \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] ,
    \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] ,
    \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
    \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] ,
    \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] ,
    \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] ,
    \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] ,
    \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] ,
    \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
    \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] ,
    \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] ,
    \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] ,
    \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] ,
    \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] ,
    \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
    \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] ,
    \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] ,
    \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] ,
    \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] ,
    \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] ,
    \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
    \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] ,
    \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] ,
    \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] ,
    \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] ,
    \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] ,
    \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
    \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] ,
    \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] ,
    \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] ,
    \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] ,
    \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] ,
    \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
    \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] ,
    \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] ,
    \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] ,
    \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] ,
    \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] ,
    \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
    \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] ,
    \A[1000] ,
    maj  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] ,
    \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] ,
    \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] ,
    \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] ,
    \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
    \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] ,
    \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] ,
    \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] ,
    \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] ,
    \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] ,
    \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
    \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] ,
    \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] ,
    \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] ,
    \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] ,
    \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] ,
    \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
    \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] ,
    \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] ,
    \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] ,
    \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] ,
    \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] ,
    \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
    \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] ,
    \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] ,
    \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] ,
    \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] ,
    \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] ,
    \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
    \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] ,
    \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] ,
    \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] ,
    \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] ,
    \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] ,
    \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
    \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] ,
    \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] ,
    \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] ,
    \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] ,
    \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] ,
    \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
    \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] ,
    \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] ,
    \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] ,
    \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] ,
    \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] ,
    \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
    \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] ,
    \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] ,
    \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] ,
    \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] ,
    \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] ,
    \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
    \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] ,
    \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] ,
    \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] ,
    \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] ,
    \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] ,
    \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
    \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] ,
    \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] ,
    \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] ,
    \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] ,
    \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] ,
    \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
    \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] ,
    \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] ,
    \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] ,
    \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] ,
    \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] ,
    \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
    \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] ,
    \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] ,
    \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] ,
    \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] ,
    \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] ,
    \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
    \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] ,
    \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] ,
    \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] ,
    \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] ,
    \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] ,
    \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
    \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] ,
    \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] ,
    \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] ,
    \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] ,
    \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] ,
    \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
    \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] ,
    \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] ,
    \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] ,
    \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] ,
    \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] ,
    \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
    \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] ,
    \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] ,
    \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] ,
    \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] ,
    \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] ,
    \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
    \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] ,
    \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] ,
    \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] ,
    \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] ,
    \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] ,
    \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
    \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] ,
    \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] ,
    \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] ,
    \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] ,
    \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] ,
    \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
    \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] ,
    \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] ,
    \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] ,
    \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] ,
    \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] ,
    \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
    \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] ,
    \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] ,
    \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] ,
    \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] ,
    \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] ,
    \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
    \A[999] , \A[1000] ;
  output maj;
  wire new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_,
    new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_,
    new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_,
    new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_,
    new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_,
    new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_,
    new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_,
    new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_,
    new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_,
    new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_,
    new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_,
    new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_,
    new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_,
    new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_,
    new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_,
    new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_,
    new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_,
    new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_,
    new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_,
    new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_,
    new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_,
    new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_,
    new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_,
    new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_,
    new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_,
    new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_,
    new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_,
    new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_,
    new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_,
    new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_,
    new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_,
    new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_,
    new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_,
    new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_,
    new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_,
    new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_,
    new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_,
    new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_,
    new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_,
    new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_,
    new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_,
    new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_,
    new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_,
    new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_,
    new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_,
    new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_,
    new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_,
    new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_,
    new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_,
    new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_,
    new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_,
    new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_,
    new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_,
    new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_,
    new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_,
    new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_,
    new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_,
    new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_,
    new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_,
    new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_,
    new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_,
    new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_,
    new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_,
    new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_,
    new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_,
    new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_,
    new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_,
    new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_,
    new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_,
    new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_,
    new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_,
    new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_,
    new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_,
    new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_,
    new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_,
    new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_,
    new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_,
    new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_,
    new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_,
    new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_,
    new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_,
    new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_,
    new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_,
    new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_,
    new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_,
    new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_,
    new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_,
    new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_,
    new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_,
    new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_,
    new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_,
    new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_,
    new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_,
    new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_,
    new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_,
    new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_,
    new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_,
    new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_,
    new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_,
    new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_,
    new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_,
    new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_,
    new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_,
    new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_,
    new_n7398_, new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_,
    new_n7404_, new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_,
    new_n7410_, new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_,
    new_n7416_, new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_,
    new_n7422_, new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_,
    new_n7428_, new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_,
    new_n7434_, new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_,
    new_n7440_, new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_,
    new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_,
    new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_,
    new_n7458_, new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_,
    new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_,
    new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_,
    new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_,
    new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_,
    new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_,
    new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_,
    new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_,
    new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_,
    new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_,
    new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_,
    new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_,
    new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_,
    new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_,
    new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_,
    new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_,
    new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_,
    new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_,
    new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_,
    new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_, new_n7577_,
    new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_, new_n7583_,
    new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_, new_n7589_,
    new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_, new_n7595_,
    new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_, new_n7601_,
    new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_,
    new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_, new_n7613_,
    new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_,
    new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_,
    new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_,
    new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_,
    new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_,
    new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_,
    new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_,
    new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_,
    new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_,
    new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_,
    new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_,
    new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_,
    new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_, new_n7691_,
    new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_,
    new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_,
    new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_,
    new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_,
    new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_,
    new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_,
    new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_,
    new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_,
    new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_,
    new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_,
    new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_,
    new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_,
    new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_,
    new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_,
    new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_,
    new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_,
    new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_,
    new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_,
    new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_,
    new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_,
    new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_,
    new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_,
    new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_,
    new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_,
    new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_,
    new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_,
    new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_,
    new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_,
    new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_,
    new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_,
    new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_,
    new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_,
    new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_,
    new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_,
    new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_,
    new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_,
    new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_,
    new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_,
    new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_,
    new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_,
    new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_,
    new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_,
    new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_,
    new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_,
    new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_,
    new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_,
    new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_,
    new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_,
    new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_,
    new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_,
    new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_,
    new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_,
    new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_,
    new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_,
    new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_,
    new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_,
    new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_,
    new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_,
    new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_,
    new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_,
    new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_,
    new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_,
    new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_,
    new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_,
    new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_,
    new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_,
    new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_,
    new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_,
    new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_,
    new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_,
    new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_,
    new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_,
    new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_,
    new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_,
    new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_,
    new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_,
    new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_,
    new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_,
    new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_,
    new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_,
    new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_,
    new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_,
    new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_,
    new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_,
    new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_,
    new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_,
    new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_,
    new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_,
    new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_,
    new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_,
    new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_,
    new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_,
    new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_,
    new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_,
    new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_,
    new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_,
    new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_,
    new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_,
    new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_,
    new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_,
    new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_,
    new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_,
    new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_,
    new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_,
    new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_,
    new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_,
    new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_,
    new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_,
    new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_,
    new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_,
    new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_,
    new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_,
    new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_,
    new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_,
    new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_,
    new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_,
    new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_,
    new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_,
    new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_,
    new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_,
    new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_,
    new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_,
    new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_,
    new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_,
    new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_,
    new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_,
    new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_,
    new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_,
    new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_,
    new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_,
    new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_,
    new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_,
    new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_,
    new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_,
    new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_,
    new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_,
    new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_,
    new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_,
    new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_,
    new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12001_, new_n12002_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12015_,
    new_n12016_, new_n12017_, new_n12018_, new_n12019_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12079_, new_n12080_,
    new_n12081_, new_n12082_, new_n12083_, new_n12084_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12091_, new_n12092_, new_n12093_, new_n12094_, new_n12095_,
    new_n12096_, new_n12097_, new_n12098_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12137_, new_n12138_, new_n12139_, new_n12140_,
    new_n12141_, new_n12142_, new_n12143_, new_n12144_, new_n12145_,
    new_n12146_, new_n12147_, new_n12148_, new_n12149_, new_n12150_,
    new_n12151_, new_n12152_, new_n12153_, new_n12154_, new_n12155_,
    new_n12156_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12331_, new_n12332_, new_n12333_, new_n12334_, new_n12335_,
    new_n12336_, new_n12337_, new_n12338_, new_n12339_, new_n12340_,
    new_n12341_, new_n12342_, new_n12343_, new_n12344_, new_n12345_,
    new_n12346_, new_n12347_, new_n12348_, new_n12349_, new_n12350_,
    new_n12351_, new_n12352_, new_n12353_, new_n12354_, new_n12355_,
    new_n12356_, new_n12357_, new_n12358_, new_n12359_, new_n12360_,
    new_n12361_, new_n12362_, new_n12363_, new_n12364_, new_n12365_,
    new_n12366_, new_n12367_, new_n12368_, new_n12369_, new_n12370_,
    new_n12371_, new_n12372_, new_n12373_, new_n12374_, new_n12375_,
    new_n12376_, new_n12377_, new_n12378_, new_n12379_, new_n12380_,
    new_n12381_, new_n12382_, new_n12383_, new_n12384_, new_n12385_,
    new_n12386_, new_n12387_, new_n12388_, new_n12389_, new_n12390_,
    new_n12391_, new_n12392_, new_n12393_, new_n12394_, new_n12395_,
    new_n12396_, new_n12397_, new_n12398_, new_n12399_, new_n12400_,
    new_n12401_, new_n12402_, new_n12403_, new_n12404_, new_n12405_,
    new_n12406_, new_n12407_, new_n12408_, new_n12409_, new_n12410_,
    new_n12411_, new_n12412_, new_n12413_, new_n12414_, new_n12415_,
    new_n12416_, new_n12417_, new_n12418_, new_n12419_, new_n12420_,
    new_n12421_, new_n12422_, new_n12423_, new_n12424_, new_n12425_,
    new_n12426_, new_n12427_, new_n12428_, new_n12429_, new_n12430_,
    new_n12431_, new_n12432_, new_n12433_, new_n12434_, new_n12435_,
    new_n12436_, new_n12437_, new_n12438_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12454_, new_n12455_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13954_, new_n13955_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14025_,
    new_n14026_, new_n14027_, new_n14028_, new_n14029_, new_n14030_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14051_, new_n14052_, new_n14053_, new_n14054_, new_n14055_,
    new_n14056_, new_n14057_, new_n14058_, new_n14059_, new_n14060_,
    new_n14061_, new_n14062_, new_n14063_, new_n14064_, new_n14065_,
    new_n14066_, new_n14067_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14073_, new_n14074_, new_n14075_,
    new_n14076_, new_n14077_, new_n14078_, new_n14079_, new_n14080_,
    new_n14081_, new_n14082_, new_n14083_, new_n14084_, new_n14085_,
    new_n14086_, new_n14087_, new_n14088_, new_n14089_, new_n14090_,
    new_n14091_, new_n14092_, new_n14093_, new_n14094_, new_n14095_,
    new_n14096_, new_n14097_, new_n14098_, new_n14099_, new_n14100_,
    new_n14101_, new_n14102_, new_n14103_, new_n14104_, new_n14105_,
    new_n14106_, new_n14107_, new_n14108_, new_n14109_, new_n14110_,
    new_n14111_, new_n14112_, new_n14113_, new_n14114_, new_n14115_,
    new_n14116_, new_n14117_, new_n14118_, new_n14119_, new_n14120_,
    new_n14121_, new_n14122_, new_n14123_, new_n14124_, new_n14125_,
    new_n14126_, new_n14127_, new_n14128_, new_n14129_, new_n14130_,
    new_n14131_, new_n14132_, new_n14133_, new_n14134_, new_n14135_,
    new_n14136_, new_n14137_, new_n14138_, new_n14139_, new_n14140_,
    new_n14141_, new_n14142_, new_n14143_, new_n14144_, new_n14145_,
    new_n14146_, new_n14147_, new_n14148_, new_n14149_, new_n14150_,
    new_n14151_, new_n14152_, new_n14153_, new_n14154_, new_n14155_,
    new_n14156_, new_n14157_, new_n14158_, new_n14159_, new_n14160_,
    new_n14161_, new_n14162_, new_n14163_, new_n14164_, new_n14165_,
    new_n14166_, new_n14167_, new_n14168_, new_n14169_, new_n14170_,
    new_n14171_, new_n14172_, new_n14173_, new_n14174_, new_n14175_,
    new_n14176_, new_n14177_, new_n14178_, new_n14179_, new_n14180_,
    new_n14181_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14187_, new_n14188_, new_n14189_, new_n14190_,
    new_n14191_, new_n14192_, new_n14193_, new_n14194_, new_n14195_,
    new_n14196_, new_n14197_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14205_,
    new_n14206_, new_n14207_, new_n14208_, new_n14209_, new_n14210_,
    new_n14211_, new_n14212_, new_n14213_, new_n14214_, new_n14215_,
    new_n14216_, new_n14217_, new_n14218_, new_n14219_, new_n14220_,
    new_n14221_, new_n14222_, new_n14223_, new_n14224_, new_n14225_,
    new_n14226_, new_n14227_, new_n14228_, new_n14229_, new_n14230_,
    new_n14231_, new_n14232_, new_n14233_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14240_,
    new_n14241_, new_n14242_, new_n14243_, new_n14244_, new_n14245_,
    new_n14246_, new_n14247_, new_n14248_, new_n14249_, new_n14250_,
    new_n14251_, new_n14252_, new_n14253_, new_n14254_, new_n14255_,
    new_n14256_, new_n14257_, new_n14258_, new_n14259_, new_n14260_,
    new_n14261_, new_n14262_, new_n14263_, new_n14264_, new_n14265_,
    new_n14266_, new_n14267_, new_n14268_, new_n14269_, new_n14270_,
    new_n14271_, new_n14272_, new_n14273_, new_n14274_, new_n14275_,
    new_n14276_, new_n14277_, new_n14278_, new_n14279_, new_n14280_,
    new_n14281_, new_n14282_, new_n14283_, new_n14284_, new_n14285_,
    new_n14286_, new_n14287_, new_n14288_, new_n14289_, new_n14290_,
    new_n14291_, new_n14292_, new_n14293_, new_n14294_, new_n14295_,
    new_n14296_, new_n14297_, new_n14298_, new_n14299_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14306_, new_n14307_, new_n14308_, new_n14309_, new_n14310_,
    new_n14311_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14318_, new_n14319_, new_n14320_,
    new_n14321_, new_n14322_, new_n14323_, new_n14324_, new_n14325_,
    new_n14326_, new_n14327_, new_n14328_, new_n14329_, new_n14330_,
    new_n14331_, new_n14332_, new_n14333_, new_n14334_, new_n14335_,
    new_n14336_, new_n14337_, new_n14338_, new_n14339_, new_n14340_,
    new_n14341_, new_n14342_, new_n14343_, new_n14344_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14350_,
    new_n14351_, new_n14352_, new_n14353_, new_n14354_, new_n14355_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14366_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14372_, new_n14373_, new_n14374_, new_n14375_,
    new_n14376_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14382_, new_n14383_, new_n14384_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14400_,
    new_n14401_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14410_,
    new_n14411_, new_n14412_, new_n14413_, new_n14414_, new_n14415_,
    new_n14416_, new_n14417_, new_n14418_, new_n14419_, new_n14420_,
    new_n14421_, new_n14422_, new_n14423_, new_n14424_, new_n14425_,
    new_n14426_, new_n14427_, new_n14428_, new_n14429_, new_n14430_,
    new_n14431_, new_n14432_, new_n14433_, new_n14434_, new_n14435_,
    new_n14436_, new_n14437_, new_n14438_, new_n14439_, new_n14440_,
    new_n14441_, new_n14442_, new_n14443_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14449_, new_n14450_,
    new_n14451_, new_n14452_, new_n14453_, new_n14454_, new_n14455_,
    new_n14456_, new_n14457_, new_n14458_, new_n14459_, new_n14460_,
    new_n14461_, new_n14462_, new_n14463_, new_n14464_, new_n14465_,
    new_n14466_, new_n14467_, new_n14468_, new_n14469_, new_n14470_,
    new_n14471_, new_n14472_, new_n14473_, new_n14474_, new_n14475_,
    new_n14476_, new_n14477_, new_n14478_, new_n14479_, new_n14480_,
    new_n14481_, new_n14482_, new_n14483_, new_n14484_, new_n14485_,
    new_n14486_, new_n14487_, new_n14488_, new_n14489_, new_n14490_,
    new_n14491_, new_n14492_, new_n14493_, new_n14494_, new_n14495_,
    new_n14496_, new_n14497_, new_n14498_, new_n14499_, new_n14500_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14530_,
    new_n14531_, new_n14532_, new_n14533_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14540_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14581_, new_n14582_, new_n14583_, new_n14584_, new_n14585_,
    new_n14586_, new_n14587_, new_n14588_, new_n14589_, new_n14590_,
    new_n14591_, new_n14592_, new_n14593_, new_n14594_, new_n14595_,
    new_n14596_, new_n14597_, new_n14598_, new_n14599_, new_n14600_,
    new_n14601_, new_n14602_, new_n14603_, new_n14604_, new_n14605_,
    new_n14606_, new_n14607_, new_n14608_, new_n14609_, new_n14610_,
    new_n14611_, new_n14612_, new_n14613_, new_n14614_, new_n14615_,
    new_n14616_, new_n14617_, new_n14618_, new_n14619_, new_n14620_,
    new_n14621_, new_n14622_, new_n14623_, new_n14624_, new_n14625_,
    new_n14626_, new_n14627_, new_n14628_, new_n14629_, new_n14630_,
    new_n14631_, new_n14632_, new_n14633_, new_n14634_, new_n14635_,
    new_n14636_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14655_,
    new_n14656_, new_n14657_, new_n14658_, new_n14659_, new_n14660_,
    new_n14661_, new_n14662_, new_n14663_, new_n14664_, new_n14665_,
    new_n14666_, new_n14667_, new_n14668_, new_n14669_, new_n14670_,
    new_n14671_, new_n14672_, new_n14673_, new_n14674_, new_n14675_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14790_,
    new_n14791_, new_n14792_, new_n14793_, new_n14794_, new_n14795_,
    new_n14796_, new_n14797_, new_n14798_, new_n14799_, new_n14800_,
    new_n14801_, new_n14802_, new_n14803_, new_n14804_, new_n14805_,
    new_n14806_, new_n14807_, new_n14808_, new_n14809_, new_n14810_,
    new_n14811_, new_n14812_, new_n14813_, new_n14814_, new_n14815_,
    new_n14816_, new_n14817_, new_n14818_, new_n14819_, new_n14820_,
    new_n14821_, new_n14822_, new_n14823_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14838_, new_n14839_, new_n14840_,
    new_n14841_, new_n14842_, new_n14843_, new_n14844_, new_n14845_,
    new_n14846_, new_n14847_, new_n14848_, new_n14849_, new_n14850_,
    new_n14851_, new_n14852_, new_n14853_, new_n14854_, new_n14855_,
    new_n14856_, new_n14857_, new_n14858_, new_n14859_, new_n14860_,
    new_n14861_, new_n14862_, new_n14863_, new_n14864_, new_n14865_,
    new_n14866_, new_n14867_, new_n14868_, new_n14869_, new_n14870_,
    new_n14871_, new_n14872_, new_n14873_, new_n14874_, new_n14875_,
    new_n14876_, new_n14877_, new_n14878_, new_n14879_, new_n14880_,
    new_n14881_, new_n14882_, new_n14883_, new_n14884_, new_n14885_,
    new_n14886_, new_n14887_, new_n14888_, new_n14889_, new_n14890_,
    new_n14891_, new_n14892_, new_n14893_, new_n14894_, new_n14895_,
    new_n14896_, new_n14897_, new_n14898_, new_n14899_, new_n14900_,
    new_n14901_, new_n14902_, new_n14903_, new_n14904_, new_n14905_,
    new_n14906_, new_n14907_, new_n14908_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15031_, new_n15032_, new_n15033_, new_n15034_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15044_, new_n15045_,
    new_n15046_, new_n15047_, new_n15048_, new_n15049_, new_n15050_,
    new_n15051_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15146_, new_n15147_, new_n15148_, new_n15149_, new_n15150_,
    new_n15151_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15192_, new_n15193_, new_n15194_, new_n15195_,
    new_n15196_, new_n15197_, new_n15198_, new_n15199_, new_n15200_,
    new_n15201_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15231_, new_n15232_, new_n15233_, new_n15234_, new_n15235_,
    new_n15236_, new_n15237_, new_n15238_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15244_, new_n15245_,
    new_n15246_, new_n15247_, new_n15248_, new_n15249_, new_n15250_,
    new_n15251_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15281_, new_n15282_, new_n15283_, new_n15284_, new_n15285_,
    new_n15286_, new_n15287_, new_n15288_, new_n15289_, new_n15290_,
    new_n15291_, new_n15292_, new_n15293_, new_n15294_, new_n15295_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15314_, new_n15315_,
    new_n15316_, new_n15317_, new_n15318_, new_n15319_, new_n15320_,
    new_n15321_, new_n15322_, new_n15323_, new_n15324_, new_n15325_,
    new_n15326_, new_n15327_, new_n15328_, new_n15329_, new_n15330_,
    new_n15331_, new_n15332_, new_n15333_, new_n15334_, new_n15335_,
    new_n15336_, new_n15337_, new_n15338_, new_n15339_, new_n15340_,
    new_n15341_, new_n15342_, new_n15343_, new_n15344_, new_n15345_,
    new_n15346_, new_n15347_, new_n15348_, new_n15349_, new_n15350_,
    new_n15351_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15359_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15366_, new_n15367_, new_n15368_, new_n15369_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15377_, new_n15378_, new_n15379_, new_n15380_,
    new_n15381_, new_n15382_, new_n15383_, new_n15384_, new_n15385_,
    new_n15386_, new_n15387_, new_n15388_, new_n15389_, new_n15390_,
    new_n15391_, new_n15392_, new_n15393_, new_n15394_, new_n15395_,
    new_n15396_, new_n15397_, new_n15398_, new_n15399_, new_n15400_,
    new_n15401_, new_n15402_, new_n15403_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15431_, new_n15432_, new_n15433_, new_n15434_, new_n15435_,
    new_n15436_, new_n15437_, new_n15438_, new_n15439_, new_n15440_,
    new_n15441_, new_n15442_, new_n15443_, new_n15444_, new_n15445_,
    new_n15446_, new_n15447_, new_n15448_, new_n15449_, new_n15450_,
    new_n15451_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15456_, new_n15457_, new_n15458_, new_n15459_, new_n15460_,
    new_n15461_, new_n15462_, new_n15463_, new_n15464_, new_n15465_,
    new_n15466_, new_n15467_, new_n15468_, new_n15469_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15481_, new_n15482_, new_n15483_, new_n15484_, new_n15485_,
    new_n15486_, new_n15487_, new_n15488_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15494_, new_n15495_,
    new_n15496_, new_n15497_, new_n15498_, new_n15499_, new_n15500_,
    new_n15501_, new_n15502_, new_n15503_, new_n15504_, new_n15505_,
    new_n15506_, new_n15507_, new_n15508_, new_n15509_, new_n15510_,
    new_n15511_, new_n15512_, new_n15513_, new_n15514_, new_n15515_,
    new_n15516_, new_n15517_, new_n15518_, new_n15519_, new_n15520_,
    new_n15521_, new_n15522_, new_n15523_, new_n15524_, new_n15525_,
    new_n15526_, new_n15527_, new_n15528_, new_n15529_, new_n15530_,
    new_n15531_, new_n15532_, new_n15533_, new_n15534_, new_n15535_,
    new_n15536_, new_n15537_, new_n15538_, new_n15539_, new_n15540_,
    new_n15541_, new_n15542_, new_n15543_, new_n15544_, new_n15545_,
    new_n15546_, new_n15547_, new_n15548_, new_n15549_, new_n15550_,
    new_n15551_, new_n15552_, new_n15553_, new_n15554_, new_n15555_,
    new_n15556_, new_n15557_, new_n15558_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_;
  INV_X1     g00000(.I(\A[200] ), .ZN(new_n1003_));
  NAND2_X1   g00001(.A1(new_n1003_), .A2(\A[201] ), .ZN(new_n1004_));
  INV_X1     g00002(.I(new_n1004_), .ZN(new_n1005_));
  NOR2_X1    g00003(.A1(new_n1003_), .A2(\A[201] ), .ZN(new_n1006_));
  OAI21_X1   g00004(.A1(new_n1005_), .A2(new_n1006_), .B(\A[199] ), .ZN(new_n1007_));
  INV_X1     g00005(.I(\A[199] ), .ZN(new_n1008_));
  NAND2_X1   g00006(.A1(\A[200] ), .A2(\A[201] ), .ZN(new_n1009_));
  INV_X1     g00007(.I(new_n1009_), .ZN(new_n1010_));
  NOR2_X1    g00008(.A1(\A[200] ), .A2(\A[201] ), .ZN(new_n1011_));
  OAI21_X1   g00009(.A1(new_n1010_), .A2(new_n1011_), .B(new_n1008_), .ZN(new_n1012_));
  INV_X1     g00010(.I(\A[204] ), .ZN(new_n1013_));
  NOR2_X1    g00011(.A1(new_n1013_), .A2(\A[203] ), .ZN(new_n1014_));
  INV_X1     g00012(.I(\A[203] ), .ZN(new_n1015_));
  NOR2_X1    g00013(.A1(new_n1015_), .A2(\A[204] ), .ZN(new_n1016_));
  OAI21_X1   g00014(.A1(new_n1014_), .A2(new_n1016_), .B(\A[202] ), .ZN(new_n1017_));
  INV_X1     g00015(.I(\A[202] ), .ZN(new_n1018_));
  NAND2_X1   g00016(.A1(\A[203] ), .A2(\A[204] ), .ZN(new_n1019_));
  INV_X1     g00017(.I(new_n1019_), .ZN(new_n1020_));
  NOR2_X1    g00018(.A1(\A[203] ), .A2(\A[204] ), .ZN(new_n1021_));
  OAI21_X1   g00019(.A1(new_n1020_), .A2(new_n1021_), .B(new_n1018_), .ZN(new_n1022_));
  NAND4_X1   g00020(.A1(new_n1007_), .A2(new_n1012_), .A3(new_n1022_), .A4(new_n1017_), .ZN(new_n1023_));
  AOI21_X1   g00021(.A1(\A[203] ), .A2(\A[204] ), .B(\A[202] ), .ZN(new_n1024_));
  NOR2_X1    g00022(.A1(new_n1024_), .A2(new_n1021_), .ZN(new_n1025_));
  AOI21_X1   g00023(.A1(\A[200] ), .A2(\A[201] ), .B(\A[199] ), .ZN(new_n1026_));
  NOR2_X1    g00024(.A1(new_n1026_), .A2(new_n1011_), .ZN(new_n1027_));
  NOR2_X1    g00025(.A1(new_n1025_), .A2(new_n1027_), .ZN(new_n1028_));
  NOR4_X1    g00026(.A1(new_n1024_), .A2(new_n1026_), .A3(new_n1011_), .A4(new_n1021_), .ZN(new_n1029_));
  NOR2_X1    g00027(.A1(new_n1028_), .A2(new_n1029_), .ZN(new_n1030_));
  NAND2_X1   g00028(.A1(new_n1023_), .A2(new_n1030_), .ZN(new_n1031_));
  INV_X1     g00029(.I(\A[201] ), .ZN(new_n1032_));
  NAND2_X1   g00030(.A1(new_n1032_), .A2(\A[200] ), .ZN(new_n1033_));
  AOI21_X1   g00031(.A1(new_n1004_), .A2(new_n1033_), .B(new_n1008_), .ZN(new_n1034_));
  INV_X1     g00032(.I(new_n1011_), .ZN(new_n1035_));
  AOI21_X1   g00033(.A1(new_n1035_), .A2(new_n1009_), .B(\A[199] ), .ZN(new_n1036_));
  NAND2_X1   g00034(.A1(new_n1015_), .A2(\A[204] ), .ZN(new_n1037_));
  NAND2_X1   g00035(.A1(new_n1013_), .A2(\A[203] ), .ZN(new_n1038_));
  AOI21_X1   g00036(.A1(new_n1037_), .A2(new_n1038_), .B(new_n1018_), .ZN(new_n1039_));
  INV_X1     g00037(.I(new_n1021_), .ZN(new_n1040_));
  AOI21_X1   g00038(.A1(new_n1040_), .A2(new_n1019_), .B(\A[202] ), .ZN(new_n1041_));
  NOR4_X1    g00039(.A1(new_n1034_), .A2(new_n1036_), .A3(new_n1041_), .A4(new_n1039_), .ZN(new_n1042_));
  OAI22_X1   g00040(.A1(new_n1011_), .A2(new_n1026_), .B1(new_n1024_), .B2(new_n1021_), .ZN(new_n1043_));
  INV_X1     g00041(.I(new_n1029_), .ZN(new_n1044_));
  NAND2_X1   g00042(.A1(new_n1044_), .A2(new_n1043_), .ZN(new_n1045_));
  NAND2_X1   g00043(.A1(new_n1042_), .A2(new_n1045_), .ZN(new_n1046_));
  NAND2_X1   g00044(.A1(new_n1031_), .A2(new_n1046_), .ZN(new_n1047_));
  INV_X1     g00045(.I(\A[207] ), .ZN(new_n1048_));
  NOR2_X1    g00046(.A1(new_n1048_), .A2(\A[206] ), .ZN(new_n1049_));
  INV_X1     g00047(.I(\A[206] ), .ZN(new_n1050_));
  NOR2_X1    g00048(.A1(new_n1050_), .A2(\A[207] ), .ZN(new_n1051_));
  OAI21_X1   g00049(.A1(new_n1049_), .A2(new_n1051_), .B(\A[205] ), .ZN(new_n1052_));
  INV_X1     g00050(.I(\A[205] ), .ZN(new_n1053_));
  NAND2_X1   g00051(.A1(\A[206] ), .A2(\A[207] ), .ZN(new_n1054_));
  INV_X1     g00052(.I(new_n1054_), .ZN(new_n1055_));
  NOR2_X1    g00053(.A1(\A[206] ), .A2(\A[207] ), .ZN(new_n1056_));
  OAI21_X1   g00054(.A1(new_n1055_), .A2(new_n1056_), .B(new_n1053_), .ZN(new_n1057_));
  INV_X1     g00055(.I(\A[210] ), .ZN(new_n1058_));
  NOR2_X1    g00056(.A1(new_n1058_), .A2(\A[209] ), .ZN(new_n1059_));
  INV_X1     g00057(.I(\A[209] ), .ZN(new_n1060_));
  NOR2_X1    g00058(.A1(new_n1060_), .A2(\A[210] ), .ZN(new_n1061_));
  OAI21_X1   g00059(.A1(new_n1059_), .A2(new_n1061_), .B(\A[208] ), .ZN(new_n1062_));
  INV_X1     g00060(.I(\A[208] ), .ZN(new_n1063_));
  NAND2_X1   g00061(.A1(\A[209] ), .A2(\A[210] ), .ZN(new_n1064_));
  INV_X1     g00062(.I(new_n1064_), .ZN(new_n1065_));
  NOR2_X1    g00063(.A1(\A[209] ), .A2(\A[210] ), .ZN(new_n1066_));
  OAI21_X1   g00064(.A1(new_n1065_), .A2(new_n1066_), .B(new_n1063_), .ZN(new_n1067_));
  NAND4_X1   g00065(.A1(new_n1052_), .A2(new_n1057_), .A3(new_n1062_), .A4(new_n1067_), .ZN(new_n1068_));
  AOI21_X1   g00066(.A1(new_n1063_), .A2(new_n1064_), .B(new_n1066_), .ZN(new_n1069_));
  AOI21_X1   g00067(.A1(\A[206] ), .A2(\A[207] ), .B(\A[205] ), .ZN(new_n1070_));
  NOR2_X1    g00068(.A1(new_n1070_), .A2(new_n1056_), .ZN(new_n1071_));
  XNOR2_X1   g00069(.A1(new_n1069_), .A2(new_n1071_), .ZN(new_n1072_));
  NOR2_X1    g00070(.A1(new_n1072_), .A2(new_n1068_), .ZN(new_n1073_));
  NAND2_X1   g00071(.A1(new_n1050_), .A2(\A[207] ), .ZN(new_n1074_));
  NAND2_X1   g00072(.A1(new_n1048_), .A2(\A[206] ), .ZN(new_n1075_));
  AOI21_X1   g00073(.A1(new_n1074_), .A2(new_n1075_), .B(new_n1053_), .ZN(new_n1076_));
  INV_X1     g00074(.I(new_n1056_), .ZN(new_n1077_));
  AOI21_X1   g00075(.A1(new_n1077_), .A2(new_n1054_), .B(\A[205] ), .ZN(new_n1078_));
  NAND2_X1   g00076(.A1(new_n1060_), .A2(\A[210] ), .ZN(new_n1079_));
  NAND2_X1   g00077(.A1(new_n1058_), .A2(\A[209] ), .ZN(new_n1080_));
  AOI21_X1   g00078(.A1(new_n1079_), .A2(new_n1080_), .B(new_n1063_), .ZN(new_n1081_));
  INV_X1     g00079(.I(new_n1066_), .ZN(new_n1082_));
  AOI21_X1   g00080(.A1(new_n1082_), .A2(new_n1064_), .B(\A[208] ), .ZN(new_n1083_));
  NOR4_X1    g00081(.A1(new_n1076_), .A2(new_n1078_), .A3(new_n1083_), .A4(new_n1081_), .ZN(new_n1084_));
  XOR2_X1    g00082(.A1(new_n1069_), .A2(new_n1071_), .Z(new_n1085_));
  NOR2_X1    g00083(.A1(new_n1085_), .A2(new_n1084_), .ZN(new_n1086_));
  OAI22_X1   g00084(.A1(new_n1034_), .A2(new_n1036_), .B1(new_n1041_), .B2(new_n1039_), .ZN(new_n1087_));
  NAND2_X1   g00085(.A1(new_n1023_), .A2(new_n1087_), .ZN(new_n1088_));
  OAI22_X1   g00086(.A1(new_n1076_), .A2(new_n1078_), .B1(new_n1083_), .B2(new_n1081_), .ZN(new_n1089_));
  NAND2_X1   g00087(.A1(new_n1089_), .A2(new_n1068_), .ZN(new_n1090_));
  OAI22_X1   g00088(.A1(new_n1073_), .A2(new_n1086_), .B1(new_n1088_), .B2(new_n1090_), .ZN(new_n1091_));
  AOI22_X1   g00089(.A1(new_n1007_), .A2(new_n1012_), .B1(new_n1022_), .B2(new_n1017_), .ZN(new_n1092_));
  NOR2_X1    g00090(.A1(new_n1092_), .A2(new_n1042_), .ZN(new_n1093_));
  NAND3_X1   g00091(.A1(new_n1089_), .A2(new_n1069_), .A3(new_n1071_), .ZN(new_n1094_));
  AOI22_X1   g00092(.A1(new_n1052_), .A2(new_n1057_), .B1(new_n1062_), .B2(new_n1067_), .ZN(new_n1095_));
  NOR3_X1    g00093(.A1(new_n1072_), .A2(new_n1095_), .A3(new_n1084_), .ZN(new_n1096_));
  NAND3_X1   g00094(.A1(new_n1096_), .A2(new_n1093_), .A3(new_n1094_), .ZN(new_n1097_));
  NAND3_X1   g00095(.A1(new_n1091_), .A2(new_n1097_), .A3(new_n1047_), .ZN(new_n1098_));
  INV_X1     g00096(.I(new_n1047_), .ZN(new_n1099_));
  NAND2_X1   g00097(.A1(new_n1085_), .A2(new_n1084_), .ZN(new_n1100_));
  NAND2_X1   g00098(.A1(new_n1072_), .A2(new_n1068_), .ZN(new_n1101_));
  NOR2_X1    g00099(.A1(new_n1095_), .A2(new_n1084_), .ZN(new_n1102_));
  AOI22_X1   g00100(.A1(new_n1100_), .A2(new_n1101_), .B1(new_n1093_), .B2(new_n1102_), .ZN(new_n1103_));
  NOR4_X1    g00101(.A1(new_n1088_), .A2(new_n1084_), .A3(new_n1072_), .A4(new_n1095_), .ZN(new_n1104_));
  OAI21_X1   g00102(.A1(new_n1103_), .A2(new_n1104_), .B(new_n1099_), .ZN(new_n1105_));
  NAND2_X1   g00103(.A1(new_n1105_), .A2(new_n1098_), .ZN(new_n1106_));
  INV_X1     g00104(.I(\A[211] ), .ZN(new_n1107_));
  INV_X1     g00105(.I(\A[212] ), .ZN(new_n1108_));
  NAND2_X1   g00106(.A1(new_n1108_), .A2(\A[213] ), .ZN(new_n1109_));
  INV_X1     g00107(.I(\A[213] ), .ZN(new_n1110_));
  NAND2_X1   g00108(.A1(new_n1110_), .A2(\A[212] ), .ZN(new_n1111_));
  AOI21_X1   g00109(.A1(new_n1109_), .A2(new_n1111_), .B(new_n1107_), .ZN(new_n1112_));
  NAND2_X1   g00110(.A1(\A[212] ), .A2(\A[213] ), .ZN(new_n1113_));
  NOR2_X1    g00111(.A1(\A[212] ), .A2(\A[213] ), .ZN(new_n1114_));
  INV_X1     g00112(.I(new_n1114_), .ZN(new_n1115_));
  AOI21_X1   g00113(.A1(new_n1115_), .A2(new_n1113_), .B(\A[211] ), .ZN(new_n1116_));
  INV_X1     g00114(.I(\A[214] ), .ZN(new_n1117_));
  INV_X1     g00115(.I(\A[215] ), .ZN(new_n1118_));
  NAND2_X1   g00116(.A1(new_n1118_), .A2(\A[216] ), .ZN(new_n1119_));
  INV_X1     g00117(.I(\A[216] ), .ZN(new_n1120_));
  NAND2_X1   g00118(.A1(new_n1120_), .A2(\A[215] ), .ZN(new_n1121_));
  AOI21_X1   g00119(.A1(new_n1119_), .A2(new_n1121_), .B(new_n1117_), .ZN(new_n1122_));
  NAND2_X1   g00120(.A1(\A[215] ), .A2(\A[216] ), .ZN(new_n1123_));
  OR2_X2     g00121(.A1(\A[215] ), .A2(\A[216] ), .Z(new_n1124_));
  AOI21_X1   g00122(.A1(new_n1124_), .A2(new_n1123_), .B(\A[214] ), .ZN(new_n1125_));
  NOR4_X1    g00123(.A1(new_n1112_), .A2(new_n1116_), .A3(new_n1122_), .A4(new_n1125_), .ZN(new_n1126_));
  NOR2_X1    g00124(.A1(\A[215] ), .A2(\A[216] ), .ZN(new_n1127_));
  AOI21_X1   g00125(.A1(\A[215] ), .A2(\A[216] ), .B(\A[214] ), .ZN(new_n1128_));
  AOI21_X1   g00126(.A1(\A[212] ), .A2(\A[213] ), .B(\A[211] ), .ZN(new_n1129_));
  OAI22_X1   g00127(.A1(new_n1114_), .A2(new_n1129_), .B1(new_n1128_), .B2(new_n1127_), .ZN(new_n1130_));
  NOR4_X1    g00128(.A1(new_n1128_), .A2(new_n1129_), .A3(new_n1114_), .A4(new_n1127_), .ZN(new_n1131_));
  INV_X1     g00129(.I(new_n1131_), .ZN(new_n1132_));
  NAND2_X1   g00130(.A1(new_n1132_), .A2(new_n1130_), .ZN(new_n1133_));
  XOR2_X1    g00131(.A1(new_n1126_), .A2(new_n1133_), .Z(new_n1134_));
  INV_X1     g00132(.I(\A[219] ), .ZN(new_n1135_));
  NOR2_X1    g00133(.A1(new_n1135_), .A2(\A[218] ), .ZN(new_n1136_));
  INV_X1     g00134(.I(\A[218] ), .ZN(new_n1137_));
  NOR2_X1    g00135(.A1(new_n1137_), .A2(\A[219] ), .ZN(new_n1138_));
  OAI21_X1   g00136(.A1(new_n1136_), .A2(new_n1138_), .B(\A[217] ), .ZN(new_n1139_));
  INV_X1     g00137(.I(\A[217] ), .ZN(new_n1140_));
  AND2_X2    g00138(.A1(\A[218] ), .A2(\A[219] ), .Z(new_n1141_));
  NOR2_X1    g00139(.A1(\A[218] ), .A2(\A[219] ), .ZN(new_n1142_));
  OAI21_X1   g00140(.A1(new_n1141_), .A2(new_n1142_), .B(new_n1140_), .ZN(new_n1143_));
  INV_X1     g00141(.I(\A[222] ), .ZN(new_n1144_));
  NOR2_X1    g00142(.A1(new_n1144_), .A2(\A[221] ), .ZN(new_n1145_));
  INV_X1     g00143(.I(\A[221] ), .ZN(new_n1146_));
  NOR2_X1    g00144(.A1(new_n1146_), .A2(\A[222] ), .ZN(new_n1147_));
  OAI21_X1   g00145(.A1(new_n1145_), .A2(new_n1147_), .B(\A[220] ), .ZN(new_n1148_));
  INV_X1     g00146(.I(\A[220] ), .ZN(new_n1149_));
  AND2_X2    g00147(.A1(\A[221] ), .A2(\A[222] ), .Z(new_n1150_));
  NOR2_X1    g00148(.A1(\A[221] ), .A2(\A[222] ), .ZN(new_n1151_));
  OAI21_X1   g00149(.A1(new_n1150_), .A2(new_n1151_), .B(new_n1149_), .ZN(new_n1152_));
  NAND4_X1   g00150(.A1(new_n1139_), .A2(new_n1148_), .A3(new_n1143_), .A4(new_n1152_), .ZN(new_n1153_));
  AOI21_X1   g00151(.A1(\A[221] ), .A2(\A[222] ), .B(\A[220] ), .ZN(new_n1154_));
  AOI21_X1   g00152(.A1(\A[218] ), .A2(\A[219] ), .B(\A[217] ), .ZN(new_n1155_));
  NOR2_X1    g00153(.A1(new_n1155_), .A2(new_n1142_), .ZN(new_n1156_));
  NOR3_X1    g00154(.A1(new_n1156_), .A2(new_n1151_), .A3(new_n1154_), .ZN(new_n1157_));
  NOR2_X1    g00155(.A1(new_n1154_), .A2(new_n1151_), .ZN(new_n1158_));
  NOR3_X1    g00156(.A1(new_n1158_), .A2(new_n1142_), .A3(new_n1155_), .ZN(new_n1159_));
  NOR2_X1    g00157(.A1(new_n1159_), .A2(new_n1157_), .ZN(new_n1160_));
  NOR2_X1    g00158(.A1(new_n1160_), .A2(new_n1153_), .ZN(new_n1161_));
  NAND2_X1   g00159(.A1(new_n1137_), .A2(\A[219] ), .ZN(new_n1162_));
  NAND2_X1   g00160(.A1(new_n1135_), .A2(\A[218] ), .ZN(new_n1163_));
  AOI21_X1   g00161(.A1(new_n1162_), .A2(new_n1163_), .B(new_n1140_), .ZN(new_n1164_));
  NAND2_X1   g00162(.A1(\A[218] ), .A2(\A[219] ), .ZN(new_n1165_));
  INV_X1     g00163(.I(new_n1142_), .ZN(new_n1166_));
  AOI21_X1   g00164(.A1(new_n1166_), .A2(new_n1165_), .B(\A[217] ), .ZN(new_n1167_));
  NAND2_X1   g00165(.A1(new_n1146_), .A2(\A[222] ), .ZN(new_n1168_));
  NAND2_X1   g00166(.A1(new_n1144_), .A2(\A[221] ), .ZN(new_n1169_));
  AOI21_X1   g00167(.A1(new_n1168_), .A2(new_n1169_), .B(new_n1149_), .ZN(new_n1170_));
  NAND2_X1   g00168(.A1(\A[221] ), .A2(\A[222] ), .ZN(new_n1171_));
  OR2_X2     g00169(.A1(\A[221] ), .A2(\A[222] ), .Z(new_n1172_));
  AOI21_X1   g00170(.A1(new_n1172_), .A2(new_n1171_), .B(\A[220] ), .ZN(new_n1173_));
  NOR4_X1    g00171(.A1(new_n1164_), .A2(new_n1167_), .A3(new_n1170_), .A4(new_n1173_), .ZN(new_n1174_));
  XOR2_X1    g00172(.A1(new_n1158_), .A2(new_n1156_), .Z(new_n1175_));
  NOR2_X1    g00173(.A1(new_n1175_), .A2(new_n1174_), .ZN(new_n1176_));
  NOR2_X1    g00174(.A1(new_n1110_), .A2(\A[212] ), .ZN(new_n1177_));
  NOR2_X1    g00175(.A1(new_n1108_), .A2(\A[213] ), .ZN(new_n1178_));
  OAI21_X1   g00176(.A1(new_n1177_), .A2(new_n1178_), .B(\A[211] ), .ZN(new_n1179_));
  INV_X1     g00177(.I(new_n1113_), .ZN(new_n1180_));
  OAI21_X1   g00178(.A1(new_n1180_), .A2(new_n1114_), .B(new_n1107_), .ZN(new_n1181_));
  NOR2_X1    g00179(.A1(new_n1120_), .A2(\A[215] ), .ZN(new_n1182_));
  NOR2_X1    g00180(.A1(new_n1118_), .A2(\A[216] ), .ZN(new_n1183_));
  OAI21_X1   g00181(.A1(new_n1182_), .A2(new_n1183_), .B(\A[214] ), .ZN(new_n1184_));
  INV_X1     g00182(.I(new_n1123_), .ZN(new_n1185_));
  OAI21_X1   g00183(.A1(new_n1185_), .A2(new_n1127_), .B(new_n1117_), .ZN(new_n1186_));
  NAND4_X1   g00184(.A1(new_n1179_), .A2(new_n1181_), .A3(new_n1184_), .A4(new_n1186_), .ZN(new_n1187_));
  OAI22_X1   g00185(.A1(new_n1112_), .A2(new_n1116_), .B1(new_n1122_), .B2(new_n1125_), .ZN(new_n1188_));
  NAND2_X1   g00186(.A1(new_n1187_), .A2(new_n1188_), .ZN(new_n1189_));
  OAI22_X1   g00187(.A1(new_n1164_), .A2(new_n1167_), .B1(new_n1170_), .B2(new_n1173_), .ZN(new_n1190_));
  NAND2_X1   g00188(.A1(new_n1190_), .A2(new_n1153_), .ZN(new_n1191_));
  OAI22_X1   g00189(.A1(new_n1176_), .A2(new_n1161_), .B1(new_n1189_), .B2(new_n1191_), .ZN(new_n1192_));
  AOI22_X1   g00190(.A1(new_n1179_), .A2(new_n1181_), .B1(new_n1184_), .B2(new_n1186_), .ZN(new_n1193_));
  NOR2_X1    g00191(.A1(new_n1193_), .A2(new_n1126_), .ZN(new_n1194_));
  NAND3_X1   g00192(.A1(new_n1190_), .A2(new_n1158_), .A3(new_n1156_), .ZN(new_n1195_));
  AOI22_X1   g00193(.A1(new_n1139_), .A2(new_n1143_), .B1(new_n1148_), .B2(new_n1152_), .ZN(new_n1196_));
  NOR3_X1    g00194(.A1(new_n1160_), .A2(new_n1196_), .A3(new_n1174_), .ZN(new_n1197_));
  NAND3_X1   g00195(.A1(new_n1197_), .A2(new_n1194_), .A3(new_n1195_), .ZN(new_n1198_));
  AOI21_X1   g00196(.A1(new_n1192_), .A2(new_n1198_), .B(new_n1134_), .ZN(new_n1199_));
  XOR2_X1    g00197(.A1(new_n1187_), .A2(new_n1133_), .Z(new_n1200_));
  NAND2_X1   g00198(.A1(new_n1175_), .A2(new_n1174_), .ZN(new_n1201_));
  NAND2_X1   g00199(.A1(new_n1160_), .A2(new_n1153_), .ZN(new_n1202_));
  NOR2_X1    g00200(.A1(new_n1196_), .A2(new_n1174_), .ZN(new_n1203_));
  AOI22_X1   g00201(.A1(new_n1201_), .A2(new_n1202_), .B1(new_n1194_), .B2(new_n1203_), .ZN(new_n1204_));
  NOR4_X1    g00202(.A1(new_n1189_), .A2(new_n1174_), .A3(new_n1160_), .A4(new_n1196_), .ZN(new_n1205_));
  NOR3_X1    g00203(.A1(new_n1204_), .A2(new_n1200_), .A3(new_n1205_), .ZN(new_n1206_));
  NAND2_X1   g00204(.A1(new_n1093_), .A2(new_n1090_), .ZN(new_n1207_));
  NAND2_X1   g00205(.A1(new_n1102_), .A2(new_n1088_), .ZN(new_n1208_));
  NAND4_X1   g00206(.A1(new_n1187_), .A2(new_n1188_), .A3(new_n1190_), .A4(new_n1153_), .ZN(new_n1209_));
  OAI22_X1   g00207(.A1(new_n1126_), .A2(new_n1193_), .B1(new_n1196_), .B2(new_n1174_), .ZN(new_n1210_));
  NAND2_X1   g00208(.A1(new_n1210_), .A2(new_n1209_), .ZN(new_n1211_));
  AOI21_X1   g00209(.A1(new_n1207_), .A2(new_n1208_), .B(new_n1211_), .ZN(new_n1212_));
  OAI21_X1   g00210(.A1(new_n1199_), .A2(new_n1206_), .B(new_n1212_), .ZN(new_n1213_));
  INV_X1     g00211(.I(new_n1158_), .ZN(new_n1214_));
  INV_X1     g00212(.I(new_n1156_), .ZN(new_n1215_));
  NOR3_X1    g00213(.A1(new_n1196_), .A2(new_n1214_), .A3(new_n1215_), .ZN(new_n1216_));
  NAND3_X1   g00214(.A1(new_n1175_), .A2(new_n1153_), .A3(new_n1190_), .ZN(new_n1217_));
  NOR3_X1    g00215(.A1(new_n1217_), .A2(new_n1216_), .A3(new_n1189_), .ZN(new_n1218_));
  OAI21_X1   g00216(.A1(new_n1204_), .A2(new_n1218_), .B(new_n1200_), .ZN(new_n1219_));
  NAND4_X1   g00217(.A1(new_n1194_), .A2(new_n1153_), .A3(new_n1175_), .A4(new_n1190_), .ZN(new_n1220_));
  NAND3_X1   g00218(.A1(new_n1192_), .A2(new_n1134_), .A3(new_n1220_), .ZN(new_n1221_));
  NOR2_X1    g00219(.A1(new_n1102_), .A2(new_n1088_), .ZN(new_n1222_));
  NOR2_X1    g00220(.A1(new_n1093_), .A2(new_n1090_), .ZN(new_n1223_));
  NOR4_X1    g00221(.A1(new_n1126_), .A2(new_n1193_), .A3(new_n1196_), .A4(new_n1174_), .ZN(new_n1224_));
  AOI22_X1   g00222(.A1(new_n1187_), .A2(new_n1188_), .B1(new_n1190_), .B2(new_n1153_), .ZN(new_n1225_));
  NOR2_X1    g00223(.A1(new_n1224_), .A2(new_n1225_), .ZN(new_n1226_));
  OAI21_X1   g00224(.A1(new_n1222_), .A2(new_n1223_), .B(new_n1226_), .ZN(new_n1227_));
  NAND3_X1   g00225(.A1(new_n1227_), .A2(new_n1219_), .A3(new_n1221_), .ZN(new_n1228_));
  AOI21_X1   g00226(.A1(new_n1213_), .A2(new_n1228_), .B(new_n1106_), .ZN(new_n1229_));
  INV_X1     g00227(.I(new_n1069_), .ZN(new_n1230_));
  INV_X1     g00228(.I(new_n1071_), .ZN(new_n1231_));
  NOR3_X1    g00229(.A1(new_n1095_), .A2(new_n1230_), .A3(new_n1231_), .ZN(new_n1232_));
  NAND3_X1   g00230(.A1(new_n1085_), .A2(new_n1089_), .A3(new_n1068_), .ZN(new_n1233_));
  NOR3_X1    g00231(.A1(new_n1233_), .A2(new_n1232_), .A3(new_n1088_), .ZN(new_n1234_));
  NOR3_X1    g00232(.A1(new_n1103_), .A2(new_n1099_), .A3(new_n1234_), .ZN(new_n1235_));
  NAND4_X1   g00233(.A1(new_n1093_), .A2(new_n1068_), .A3(new_n1085_), .A4(new_n1089_), .ZN(new_n1236_));
  AOI21_X1   g00234(.A1(new_n1091_), .A2(new_n1236_), .B(new_n1047_), .ZN(new_n1237_));
  NOR2_X1    g00235(.A1(new_n1235_), .A2(new_n1237_), .ZN(new_n1238_));
  AOI21_X1   g00236(.A1(new_n1219_), .A2(new_n1221_), .B(new_n1227_), .ZN(new_n1239_));
  NOR3_X1    g00237(.A1(new_n1212_), .A2(new_n1206_), .A3(new_n1199_), .ZN(new_n1240_));
  NOR3_X1    g00238(.A1(new_n1239_), .A2(new_n1240_), .A3(new_n1238_), .ZN(new_n1241_));
  OR2_X2     g00239(.A1(new_n1241_), .A2(new_n1229_), .Z(new_n1242_));
  INV_X1     g00240(.I(\A[193] ), .ZN(new_n1243_));
  INV_X1     g00241(.I(\A[194] ), .ZN(new_n1244_));
  NAND2_X1   g00242(.A1(new_n1244_), .A2(\A[195] ), .ZN(new_n1245_));
  INV_X1     g00243(.I(\A[195] ), .ZN(new_n1246_));
  NAND2_X1   g00244(.A1(new_n1246_), .A2(\A[194] ), .ZN(new_n1247_));
  AOI21_X1   g00245(.A1(new_n1245_), .A2(new_n1247_), .B(new_n1243_), .ZN(new_n1248_));
  NOR2_X1    g00246(.A1(\A[194] ), .A2(\A[195] ), .ZN(new_n1249_));
  INV_X1     g00247(.I(new_n1249_), .ZN(new_n1250_));
  NAND2_X1   g00248(.A1(\A[194] ), .A2(\A[195] ), .ZN(new_n1251_));
  AOI21_X1   g00249(.A1(new_n1250_), .A2(new_n1251_), .B(\A[193] ), .ZN(new_n1252_));
  INV_X1     g00250(.I(\A[196] ), .ZN(new_n1253_));
  INV_X1     g00251(.I(\A[197] ), .ZN(new_n1254_));
  NAND2_X1   g00252(.A1(new_n1254_), .A2(\A[198] ), .ZN(new_n1255_));
  INV_X1     g00253(.I(\A[198] ), .ZN(new_n1256_));
  NAND2_X1   g00254(.A1(new_n1256_), .A2(\A[197] ), .ZN(new_n1257_));
  AOI21_X1   g00255(.A1(new_n1255_), .A2(new_n1257_), .B(new_n1253_), .ZN(new_n1258_));
  NOR2_X1    g00256(.A1(\A[197] ), .A2(\A[198] ), .ZN(new_n1259_));
  INV_X1     g00257(.I(new_n1259_), .ZN(new_n1260_));
  NAND2_X1   g00258(.A1(\A[197] ), .A2(\A[198] ), .ZN(new_n1261_));
  AOI21_X1   g00259(.A1(new_n1260_), .A2(new_n1261_), .B(\A[196] ), .ZN(new_n1262_));
  NOR4_X1    g00260(.A1(new_n1248_), .A2(new_n1252_), .A3(new_n1262_), .A4(new_n1258_), .ZN(new_n1263_));
  NOR2_X1    g00261(.A1(new_n1246_), .A2(\A[194] ), .ZN(new_n1264_));
  NOR2_X1    g00262(.A1(new_n1244_), .A2(\A[195] ), .ZN(new_n1265_));
  OAI21_X1   g00263(.A1(new_n1264_), .A2(new_n1265_), .B(\A[193] ), .ZN(new_n1266_));
  INV_X1     g00264(.I(new_n1251_), .ZN(new_n1267_));
  OAI21_X1   g00265(.A1(new_n1267_), .A2(new_n1249_), .B(new_n1243_), .ZN(new_n1268_));
  NOR2_X1    g00266(.A1(new_n1256_), .A2(\A[197] ), .ZN(new_n1269_));
  NOR2_X1    g00267(.A1(new_n1254_), .A2(\A[198] ), .ZN(new_n1270_));
  OAI21_X1   g00268(.A1(new_n1269_), .A2(new_n1270_), .B(\A[196] ), .ZN(new_n1271_));
  AND2_X2    g00269(.A1(\A[197] ), .A2(\A[198] ), .Z(new_n1272_));
  OAI21_X1   g00270(.A1(new_n1272_), .A2(new_n1259_), .B(new_n1253_), .ZN(new_n1273_));
  AOI22_X1   g00271(.A1(new_n1266_), .A2(new_n1268_), .B1(new_n1271_), .B2(new_n1273_), .ZN(new_n1274_));
  NOR2_X1    g00272(.A1(new_n1263_), .A2(new_n1274_), .ZN(new_n1275_));
  INV_X1     g00273(.I(\A[189] ), .ZN(new_n1276_));
  NOR2_X1    g00274(.A1(new_n1276_), .A2(\A[188] ), .ZN(new_n1277_));
  INV_X1     g00275(.I(\A[188] ), .ZN(new_n1278_));
  NOR2_X1    g00276(.A1(new_n1278_), .A2(\A[189] ), .ZN(new_n1279_));
  OAI21_X1   g00277(.A1(new_n1277_), .A2(new_n1279_), .B(\A[187] ), .ZN(new_n1280_));
  INV_X1     g00278(.I(\A[187] ), .ZN(new_n1281_));
  NAND2_X1   g00279(.A1(\A[188] ), .A2(\A[189] ), .ZN(new_n1282_));
  INV_X1     g00280(.I(new_n1282_), .ZN(new_n1283_));
  NOR2_X1    g00281(.A1(\A[188] ), .A2(\A[189] ), .ZN(new_n1284_));
  OAI21_X1   g00282(.A1(new_n1283_), .A2(new_n1284_), .B(new_n1281_), .ZN(new_n1285_));
  INV_X1     g00283(.I(\A[192] ), .ZN(new_n1286_));
  NOR2_X1    g00284(.A1(new_n1286_), .A2(\A[191] ), .ZN(new_n1287_));
  INV_X1     g00285(.I(\A[191] ), .ZN(new_n1288_));
  NOR2_X1    g00286(.A1(new_n1288_), .A2(\A[192] ), .ZN(new_n1289_));
  OAI21_X1   g00287(.A1(new_n1287_), .A2(new_n1289_), .B(\A[190] ), .ZN(new_n1290_));
  INV_X1     g00288(.I(\A[190] ), .ZN(new_n1291_));
  AND2_X2    g00289(.A1(\A[191] ), .A2(\A[192] ), .Z(new_n1292_));
  NOR2_X1    g00290(.A1(\A[191] ), .A2(\A[192] ), .ZN(new_n1293_));
  OAI21_X1   g00291(.A1(new_n1292_), .A2(new_n1293_), .B(new_n1291_), .ZN(new_n1294_));
  NAND4_X1   g00292(.A1(new_n1280_), .A2(new_n1290_), .A3(new_n1285_), .A4(new_n1294_), .ZN(new_n1295_));
  NAND2_X1   g00293(.A1(new_n1280_), .A2(new_n1285_), .ZN(new_n1296_));
  NAND2_X1   g00294(.A1(new_n1290_), .A2(new_n1294_), .ZN(new_n1297_));
  NAND2_X1   g00295(.A1(new_n1296_), .A2(new_n1297_), .ZN(new_n1298_));
  NAND2_X1   g00296(.A1(new_n1298_), .A2(new_n1295_), .ZN(new_n1299_));
  NAND2_X1   g00297(.A1(new_n1299_), .A2(new_n1275_), .ZN(new_n1300_));
  NAND4_X1   g00298(.A1(new_n1266_), .A2(new_n1271_), .A3(new_n1268_), .A4(new_n1273_), .ZN(new_n1301_));
  OAI22_X1   g00299(.A1(new_n1248_), .A2(new_n1252_), .B1(new_n1262_), .B2(new_n1258_), .ZN(new_n1302_));
  NAND2_X1   g00300(.A1(new_n1302_), .A2(new_n1301_), .ZN(new_n1303_));
  NAND2_X1   g00301(.A1(new_n1278_), .A2(\A[189] ), .ZN(new_n1304_));
  NAND2_X1   g00302(.A1(new_n1276_), .A2(\A[188] ), .ZN(new_n1305_));
  AOI21_X1   g00303(.A1(new_n1304_), .A2(new_n1305_), .B(new_n1281_), .ZN(new_n1306_));
  INV_X1     g00304(.I(new_n1284_), .ZN(new_n1307_));
  AOI21_X1   g00305(.A1(new_n1307_), .A2(new_n1282_), .B(\A[187] ), .ZN(new_n1308_));
  NAND2_X1   g00306(.A1(new_n1288_), .A2(\A[192] ), .ZN(new_n1309_));
  NAND2_X1   g00307(.A1(new_n1286_), .A2(\A[191] ), .ZN(new_n1310_));
  AOI21_X1   g00308(.A1(new_n1309_), .A2(new_n1310_), .B(new_n1291_), .ZN(new_n1311_));
  NAND2_X1   g00309(.A1(\A[191] ), .A2(\A[192] ), .ZN(new_n1312_));
  OR2_X2     g00310(.A1(\A[191] ), .A2(\A[192] ), .Z(new_n1313_));
  AOI21_X1   g00311(.A1(new_n1313_), .A2(new_n1312_), .B(\A[190] ), .ZN(new_n1314_));
  NOR4_X1    g00312(.A1(new_n1306_), .A2(new_n1308_), .A3(new_n1311_), .A4(new_n1314_), .ZN(new_n1315_));
  NOR2_X1    g00313(.A1(new_n1308_), .A2(new_n1306_), .ZN(new_n1316_));
  NOR2_X1    g00314(.A1(new_n1311_), .A2(new_n1314_), .ZN(new_n1317_));
  NOR2_X1    g00315(.A1(new_n1316_), .A2(new_n1317_), .ZN(new_n1318_));
  NOR2_X1    g00316(.A1(new_n1318_), .A2(new_n1315_), .ZN(new_n1319_));
  NAND2_X1   g00317(.A1(new_n1319_), .A2(new_n1303_), .ZN(new_n1320_));
  INV_X1     g00318(.I(\A[181] ), .ZN(new_n1321_));
  INV_X1     g00319(.I(\A[182] ), .ZN(new_n1322_));
  NAND2_X1   g00320(.A1(new_n1322_), .A2(\A[183] ), .ZN(new_n1323_));
  INV_X1     g00321(.I(\A[183] ), .ZN(new_n1324_));
  NAND2_X1   g00322(.A1(new_n1324_), .A2(\A[182] ), .ZN(new_n1325_));
  AOI21_X1   g00323(.A1(new_n1323_), .A2(new_n1325_), .B(new_n1321_), .ZN(new_n1326_));
  NOR2_X1    g00324(.A1(\A[182] ), .A2(\A[183] ), .ZN(new_n1327_));
  INV_X1     g00325(.I(new_n1327_), .ZN(new_n1328_));
  NAND2_X1   g00326(.A1(\A[182] ), .A2(\A[183] ), .ZN(new_n1329_));
  AOI21_X1   g00327(.A1(new_n1328_), .A2(new_n1329_), .B(\A[181] ), .ZN(new_n1330_));
  INV_X1     g00328(.I(\A[184] ), .ZN(new_n1331_));
  INV_X1     g00329(.I(\A[185] ), .ZN(new_n1332_));
  NAND2_X1   g00330(.A1(new_n1332_), .A2(\A[186] ), .ZN(new_n1333_));
  INV_X1     g00331(.I(\A[186] ), .ZN(new_n1334_));
  NAND2_X1   g00332(.A1(new_n1334_), .A2(\A[185] ), .ZN(new_n1335_));
  AOI21_X1   g00333(.A1(new_n1333_), .A2(new_n1335_), .B(new_n1331_), .ZN(new_n1336_));
  NOR2_X1    g00334(.A1(\A[185] ), .A2(\A[186] ), .ZN(new_n1337_));
  INV_X1     g00335(.I(new_n1337_), .ZN(new_n1338_));
  NAND2_X1   g00336(.A1(\A[185] ), .A2(\A[186] ), .ZN(new_n1339_));
  AOI21_X1   g00337(.A1(new_n1338_), .A2(new_n1339_), .B(\A[184] ), .ZN(new_n1340_));
  NOR4_X1    g00338(.A1(new_n1326_), .A2(new_n1330_), .A3(new_n1340_), .A4(new_n1336_), .ZN(new_n1341_));
  NOR2_X1    g00339(.A1(new_n1324_), .A2(\A[182] ), .ZN(new_n1342_));
  NOR2_X1    g00340(.A1(new_n1322_), .A2(\A[183] ), .ZN(new_n1343_));
  OAI21_X1   g00341(.A1(new_n1342_), .A2(new_n1343_), .B(\A[181] ), .ZN(new_n1344_));
  INV_X1     g00342(.I(new_n1329_), .ZN(new_n1345_));
  OAI21_X1   g00343(.A1(new_n1345_), .A2(new_n1327_), .B(new_n1321_), .ZN(new_n1346_));
  NOR2_X1    g00344(.A1(new_n1334_), .A2(\A[185] ), .ZN(new_n1347_));
  NOR2_X1    g00345(.A1(new_n1332_), .A2(\A[186] ), .ZN(new_n1348_));
  OAI21_X1   g00346(.A1(new_n1347_), .A2(new_n1348_), .B(\A[184] ), .ZN(new_n1349_));
  AND2_X2    g00347(.A1(\A[185] ), .A2(\A[186] ), .Z(new_n1350_));
  OAI21_X1   g00348(.A1(new_n1350_), .A2(new_n1337_), .B(new_n1331_), .ZN(new_n1351_));
  AOI22_X1   g00349(.A1(new_n1344_), .A2(new_n1346_), .B1(new_n1349_), .B2(new_n1351_), .ZN(new_n1352_));
  NOR2_X1    g00350(.A1(new_n1341_), .A2(new_n1352_), .ZN(new_n1353_));
  INV_X1     g00351(.I(\A[177] ), .ZN(new_n1354_));
  NOR2_X1    g00352(.A1(new_n1354_), .A2(\A[176] ), .ZN(new_n1355_));
  INV_X1     g00353(.I(\A[176] ), .ZN(new_n1356_));
  NOR2_X1    g00354(.A1(new_n1356_), .A2(\A[177] ), .ZN(new_n1357_));
  OAI21_X1   g00355(.A1(new_n1355_), .A2(new_n1357_), .B(\A[175] ), .ZN(new_n1358_));
  INV_X1     g00356(.I(\A[175] ), .ZN(new_n1359_));
  NAND2_X1   g00357(.A1(\A[176] ), .A2(\A[177] ), .ZN(new_n1360_));
  INV_X1     g00358(.I(new_n1360_), .ZN(new_n1361_));
  NOR2_X1    g00359(.A1(\A[176] ), .A2(\A[177] ), .ZN(new_n1362_));
  OAI21_X1   g00360(.A1(new_n1361_), .A2(new_n1362_), .B(new_n1359_), .ZN(new_n1363_));
  INV_X1     g00361(.I(\A[180] ), .ZN(new_n1364_));
  NOR2_X1    g00362(.A1(new_n1364_), .A2(\A[179] ), .ZN(new_n1365_));
  INV_X1     g00363(.I(\A[179] ), .ZN(new_n1366_));
  NOR2_X1    g00364(.A1(new_n1366_), .A2(\A[180] ), .ZN(new_n1367_));
  OAI21_X1   g00365(.A1(new_n1365_), .A2(new_n1367_), .B(\A[178] ), .ZN(new_n1368_));
  INV_X1     g00366(.I(\A[178] ), .ZN(new_n1369_));
  NAND2_X1   g00367(.A1(\A[179] ), .A2(\A[180] ), .ZN(new_n1370_));
  INV_X1     g00368(.I(new_n1370_), .ZN(new_n1371_));
  NOR2_X1    g00369(.A1(\A[179] ), .A2(\A[180] ), .ZN(new_n1372_));
  OAI21_X1   g00370(.A1(new_n1371_), .A2(new_n1372_), .B(new_n1369_), .ZN(new_n1373_));
  NAND4_X1   g00371(.A1(new_n1358_), .A2(new_n1363_), .A3(new_n1368_), .A4(new_n1373_), .ZN(new_n1374_));
  NAND2_X1   g00372(.A1(new_n1356_), .A2(\A[177] ), .ZN(new_n1375_));
  NAND2_X1   g00373(.A1(new_n1354_), .A2(\A[176] ), .ZN(new_n1376_));
  AOI21_X1   g00374(.A1(new_n1375_), .A2(new_n1376_), .B(new_n1359_), .ZN(new_n1377_));
  INV_X1     g00375(.I(new_n1362_), .ZN(new_n1378_));
  AOI21_X1   g00376(.A1(new_n1378_), .A2(new_n1360_), .B(\A[175] ), .ZN(new_n1379_));
  NAND2_X1   g00377(.A1(new_n1366_), .A2(\A[180] ), .ZN(new_n1380_));
  NAND2_X1   g00378(.A1(new_n1364_), .A2(\A[179] ), .ZN(new_n1381_));
  AOI21_X1   g00379(.A1(new_n1380_), .A2(new_n1381_), .B(new_n1369_), .ZN(new_n1382_));
  OR2_X2     g00380(.A1(\A[179] ), .A2(\A[180] ), .Z(new_n1383_));
  AOI21_X1   g00381(.A1(new_n1383_), .A2(new_n1370_), .B(\A[178] ), .ZN(new_n1384_));
  OAI22_X1   g00382(.A1(new_n1377_), .A2(new_n1379_), .B1(new_n1382_), .B2(new_n1384_), .ZN(new_n1385_));
  NAND2_X1   g00383(.A1(new_n1374_), .A2(new_n1385_), .ZN(new_n1386_));
  NAND2_X1   g00384(.A1(new_n1353_), .A2(new_n1386_), .ZN(new_n1387_));
  NAND4_X1   g00385(.A1(new_n1344_), .A2(new_n1349_), .A3(new_n1346_), .A4(new_n1351_), .ZN(new_n1388_));
  OAI22_X1   g00386(.A1(new_n1326_), .A2(new_n1330_), .B1(new_n1340_), .B2(new_n1336_), .ZN(new_n1389_));
  NAND2_X1   g00387(.A1(new_n1389_), .A2(new_n1388_), .ZN(new_n1390_));
  NOR4_X1    g00388(.A1(new_n1377_), .A2(new_n1379_), .A3(new_n1382_), .A4(new_n1384_), .ZN(new_n1391_));
  AOI22_X1   g00389(.A1(new_n1358_), .A2(new_n1363_), .B1(new_n1368_), .B2(new_n1373_), .ZN(new_n1392_));
  NOR2_X1    g00390(.A1(new_n1392_), .A2(new_n1391_), .ZN(new_n1393_));
  NAND2_X1   g00391(.A1(new_n1393_), .A2(new_n1390_), .ZN(new_n1394_));
  AOI22_X1   g00392(.A1(new_n1320_), .A2(new_n1300_), .B1(new_n1387_), .B2(new_n1394_), .ZN(new_n1395_));
  NOR2_X1    g00393(.A1(new_n1319_), .A2(new_n1303_), .ZN(new_n1396_));
  NOR2_X1    g00394(.A1(new_n1299_), .A2(new_n1275_), .ZN(new_n1397_));
  NOR2_X1    g00395(.A1(new_n1393_), .A2(new_n1390_), .ZN(new_n1398_));
  NOR2_X1    g00396(.A1(new_n1353_), .A2(new_n1386_), .ZN(new_n1399_));
  NOR4_X1    g00397(.A1(new_n1396_), .A2(new_n1397_), .A3(new_n1399_), .A4(new_n1398_), .ZN(new_n1400_));
  NOR2_X1    g00398(.A1(new_n1400_), .A2(new_n1395_), .ZN(new_n1401_));
  NOR2_X1    g00399(.A1(new_n1222_), .A2(new_n1223_), .ZN(new_n1402_));
  XOR2_X1    g00400(.A1(new_n1189_), .A2(new_n1191_), .Z(new_n1403_));
  NAND2_X1   g00401(.A1(new_n1403_), .A2(new_n1402_), .ZN(new_n1404_));
  NAND2_X1   g00402(.A1(new_n1208_), .A2(new_n1207_), .ZN(new_n1405_));
  XOR2_X1    g00403(.A1(new_n1194_), .A2(new_n1191_), .Z(new_n1406_));
  NAND2_X1   g00404(.A1(new_n1406_), .A2(new_n1405_), .ZN(new_n1407_));
  NAND2_X1   g00405(.A1(new_n1404_), .A2(new_n1407_), .ZN(new_n1408_));
  NAND2_X1   g00406(.A1(new_n1408_), .A2(new_n1401_), .ZN(new_n1409_));
  AOI21_X1   g00407(.A1(\A[191] ), .A2(\A[192] ), .B(\A[190] ), .ZN(new_n1410_));
  NOR2_X1    g00408(.A1(new_n1410_), .A2(new_n1293_), .ZN(new_n1411_));
  AOI21_X1   g00409(.A1(\A[188] ), .A2(\A[189] ), .B(\A[187] ), .ZN(new_n1412_));
  NOR2_X1    g00410(.A1(new_n1412_), .A2(new_n1284_), .ZN(new_n1413_));
  NOR2_X1    g00411(.A1(new_n1411_), .A2(new_n1413_), .ZN(new_n1414_));
  NOR4_X1    g00412(.A1(new_n1410_), .A2(new_n1412_), .A3(new_n1284_), .A4(new_n1293_), .ZN(new_n1415_));
  NOR2_X1    g00413(.A1(new_n1414_), .A2(new_n1415_), .ZN(new_n1416_));
  NAND2_X1   g00414(.A1(new_n1295_), .A2(new_n1416_), .ZN(new_n1417_));
  OAI22_X1   g00415(.A1(new_n1284_), .A2(new_n1412_), .B1(new_n1410_), .B2(new_n1293_), .ZN(new_n1418_));
  NAND2_X1   g00416(.A1(new_n1411_), .A2(new_n1413_), .ZN(new_n1419_));
  NAND2_X1   g00417(.A1(new_n1419_), .A2(new_n1418_), .ZN(new_n1420_));
  NAND2_X1   g00418(.A1(new_n1315_), .A2(new_n1420_), .ZN(new_n1421_));
  NAND2_X1   g00419(.A1(new_n1417_), .A2(new_n1421_), .ZN(new_n1422_));
  AOI21_X1   g00420(.A1(\A[197] ), .A2(\A[198] ), .B(\A[196] ), .ZN(new_n1423_));
  NOR2_X1    g00421(.A1(new_n1423_), .A2(new_n1259_), .ZN(new_n1424_));
  AOI21_X1   g00422(.A1(\A[194] ), .A2(\A[195] ), .B(\A[193] ), .ZN(new_n1425_));
  NOR2_X1    g00423(.A1(new_n1425_), .A2(new_n1249_), .ZN(new_n1426_));
  XOR2_X1    g00424(.A1(new_n1424_), .A2(new_n1426_), .Z(new_n1427_));
  NOR2_X1    g00425(.A1(new_n1427_), .A2(new_n1263_), .ZN(new_n1428_));
  NOR3_X1    g00426(.A1(new_n1426_), .A2(new_n1259_), .A3(new_n1423_), .ZN(new_n1429_));
  NOR3_X1    g00427(.A1(new_n1424_), .A2(new_n1249_), .A3(new_n1425_), .ZN(new_n1430_));
  NOR2_X1    g00428(.A1(new_n1429_), .A2(new_n1430_), .ZN(new_n1431_));
  NOR2_X1    g00429(.A1(new_n1431_), .A2(new_n1301_), .ZN(new_n1432_));
  NOR2_X1    g00430(.A1(new_n1428_), .A2(new_n1432_), .ZN(new_n1433_));
  NOR4_X1    g00431(.A1(new_n1318_), .A2(new_n1263_), .A3(new_n1274_), .A4(new_n1315_), .ZN(new_n1434_));
  NOR2_X1    g00432(.A1(new_n1433_), .A2(new_n1434_), .ZN(new_n1435_));
  NOR4_X1    g00433(.A1(new_n1299_), .A2(new_n1263_), .A3(new_n1274_), .A4(new_n1431_), .ZN(new_n1436_));
  NOR3_X1    g00434(.A1(new_n1435_), .A2(new_n1422_), .A3(new_n1436_), .ZN(new_n1437_));
  NOR2_X1    g00435(.A1(new_n1315_), .A2(new_n1420_), .ZN(new_n1438_));
  NOR2_X1    g00436(.A1(new_n1295_), .A2(new_n1416_), .ZN(new_n1439_));
  NOR2_X1    g00437(.A1(new_n1439_), .A2(new_n1438_), .ZN(new_n1440_));
  OAI22_X1   g00438(.A1(new_n1299_), .A2(new_n1303_), .B1(new_n1428_), .B2(new_n1432_), .ZN(new_n1441_));
  NAND2_X1   g00439(.A1(new_n1431_), .A2(new_n1301_), .ZN(new_n1442_));
  NAND2_X1   g00440(.A1(new_n1427_), .A2(new_n1263_), .ZN(new_n1443_));
  NAND3_X1   g00441(.A1(new_n1434_), .A2(new_n1442_), .A3(new_n1443_), .ZN(new_n1444_));
  AOI21_X1   g00442(.A1(new_n1444_), .A2(new_n1441_), .B(new_n1440_), .ZN(new_n1445_));
  NOR2_X1    g00443(.A1(new_n1437_), .A2(new_n1445_), .ZN(new_n1446_));
  OAI22_X1   g00444(.A1(new_n1396_), .A2(new_n1397_), .B1(new_n1399_), .B2(new_n1398_), .ZN(new_n1447_));
  AOI21_X1   g00445(.A1(\A[179] ), .A2(\A[180] ), .B(\A[178] ), .ZN(new_n1448_));
  NOR2_X1    g00446(.A1(new_n1448_), .A2(new_n1372_), .ZN(new_n1449_));
  AOI21_X1   g00447(.A1(\A[176] ), .A2(\A[177] ), .B(\A[175] ), .ZN(new_n1450_));
  NOR2_X1    g00448(.A1(new_n1450_), .A2(new_n1362_), .ZN(new_n1451_));
  NOR2_X1    g00449(.A1(new_n1449_), .A2(new_n1451_), .ZN(new_n1452_));
  NOR4_X1    g00450(.A1(new_n1448_), .A2(new_n1450_), .A3(new_n1362_), .A4(new_n1372_), .ZN(new_n1453_));
  NOR2_X1    g00451(.A1(new_n1452_), .A2(new_n1453_), .ZN(new_n1454_));
  NAND2_X1   g00452(.A1(new_n1374_), .A2(new_n1454_), .ZN(new_n1455_));
  NOR2_X1    g00453(.A1(new_n1379_), .A2(new_n1377_), .ZN(new_n1456_));
  NOR2_X1    g00454(.A1(new_n1382_), .A2(new_n1384_), .ZN(new_n1457_));
  OAI22_X1   g00455(.A1(new_n1362_), .A2(new_n1450_), .B1(new_n1448_), .B2(new_n1372_), .ZN(new_n1458_));
  NAND2_X1   g00456(.A1(new_n1370_), .A2(new_n1369_), .ZN(new_n1459_));
  NAND2_X1   g00457(.A1(new_n1360_), .A2(new_n1359_), .ZN(new_n1460_));
  NAND4_X1   g00458(.A1(new_n1459_), .A2(new_n1460_), .A3(new_n1378_), .A4(new_n1383_), .ZN(new_n1461_));
  NAND2_X1   g00459(.A1(new_n1461_), .A2(new_n1458_), .ZN(new_n1462_));
  NAND3_X1   g00460(.A1(new_n1462_), .A2(new_n1456_), .A3(new_n1457_), .ZN(new_n1463_));
  NAND2_X1   g00461(.A1(new_n1455_), .A2(new_n1463_), .ZN(new_n1464_));
  AOI21_X1   g00462(.A1(\A[185] ), .A2(\A[186] ), .B(\A[184] ), .ZN(new_n1465_));
  AOI21_X1   g00463(.A1(\A[182] ), .A2(\A[183] ), .B(\A[181] ), .ZN(new_n1466_));
  NOR2_X1    g00464(.A1(new_n1466_), .A2(new_n1327_), .ZN(new_n1467_));
  NOR3_X1    g00465(.A1(new_n1467_), .A2(new_n1337_), .A3(new_n1465_), .ZN(new_n1468_));
  NOR2_X1    g00466(.A1(new_n1465_), .A2(new_n1337_), .ZN(new_n1469_));
  NOR3_X1    g00467(.A1(new_n1469_), .A2(new_n1327_), .A3(new_n1466_), .ZN(new_n1470_));
  NOR3_X1    g00468(.A1(new_n1341_), .A2(new_n1468_), .A3(new_n1470_), .ZN(new_n1471_));
  NOR2_X1    g00469(.A1(new_n1468_), .A2(new_n1470_), .ZN(new_n1472_));
  NOR2_X1    g00470(.A1(new_n1472_), .A2(new_n1388_), .ZN(new_n1473_));
  NOR2_X1    g00471(.A1(new_n1471_), .A2(new_n1473_), .ZN(new_n1474_));
  NOR4_X1    g00472(.A1(new_n1341_), .A2(new_n1392_), .A3(new_n1352_), .A4(new_n1391_), .ZN(new_n1475_));
  OAI21_X1   g00473(.A1(new_n1474_), .A2(new_n1475_), .B(new_n1464_), .ZN(new_n1476_));
  NAND4_X1   g00474(.A1(new_n1389_), .A2(new_n1374_), .A3(new_n1385_), .A4(new_n1388_), .ZN(new_n1477_));
  NOR3_X1    g00475(.A1(new_n1477_), .A2(new_n1471_), .A3(new_n1473_), .ZN(new_n1478_));
  NOR2_X1    g00476(.A1(new_n1476_), .A2(new_n1478_), .ZN(new_n1479_));
  OAI21_X1   g00477(.A1(new_n1471_), .A2(new_n1473_), .B(new_n1477_), .ZN(new_n1480_));
  NAND2_X1   g00478(.A1(new_n1472_), .A2(new_n1388_), .ZN(new_n1481_));
  XOR2_X1    g00479(.A1(new_n1469_), .A2(new_n1467_), .Z(new_n1482_));
  NAND2_X1   g00480(.A1(new_n1482_), .A2(new_n1341_), .ZN(new_n1483_));
  NAND3_X1   g00481(.A1(new_n1475_), .A2(new_n1481_), .A3(new_n1483_), .ZN(new_n1484_));
  AOI21_X1   g00482(.A1(new_n1480_), .A2(new_n1484_), .B(new_n1464_), .ZN(new_n1485_));
  NOR3_X1    g00483(.A1(new_n1479_), .A2(new_n1485_), .A3(new_n1447_), .ZN(new_n1486_));
  NAND3_X1   g00484(.A1(new_n1480_), .A2(new_n1484_), .A3(new_n1464_), .ZN(new_n1487_));
  NOR2_X1    g00485(.A1(new_n1391_), .A2(new_n1462_), .ZN(new_n1488_));
  NOR2_X1    g00486(.A1(new_n1374_), .A2(new_n1454_), .ZN(new_n1489_));
  NOR2_X1    g00487(.A1(new_n1489_), .A2(new_n1488_), .ZN(new_n1490_));
  NOR2_X1    g00488(.A1(new_n1474_), .A2(new_n1475_), .ZN(new_n1491_));
  OAI21_X1   g00489(.A1(new_n1491_), .A2(new_n1478_), .B(new_n1490_), .ZN(new_n1492_));
  AOI21_X1   g00490(.A1(new_n1492_), .A2(new_n1487_), .B(new_n1395_), .ZN(new_n1493_));
  NOR3_X1    g00491(.A1(new_n1486_), .A2(new_n1493_), .A3(new_n1446_), .ZN(new_n1494_));
  NAND3_X1   g00492(.A1(new_n1444_), .A2(new_n1441_), .A3(new_n1440_), .ZN(new_n1495_));
  OAI21_X1   g00493(.A1(new_n1435_), .A2(new_n1436_), .B(new_n1422_), .ZN(new_n1496_));
  NAND2_X1   g00494(.A1(new_n1496_), .A2(new_n1495_), .ZN(new_n1497_));
  NAND3_X1   g00495(.A1(new_n1492_), .A2(new_n1487_), .A3(new_n1395_), .ZN(new_n1498_));
  OAI21_X1   g00496(.A1(new_n1479_), .A2(new_n1485_), .B(new_n1447_), .ZN(new_n1499_));
  AOI21_X1   g00497(.A1(new_n1499_), .A2(new_n1498_), .B(new_n1497_), .ZN(new_n1500_));
  OAI21_X1   g00498(.A1(new_n1494_), .A2(new_n1500_), .B(new_n1409_), .ZN(new_n1501_));
  INV_X1     g00499(.I(new_n1401_), .ZN(new_n1502_));
  NOR2_X1    g00500(.A1(new_n1406_), .A2(new_n1405_), .ZN(new_n1503_));
  NOR2_X1    g00501(.A1(new_n1403_), .A2(new_n1402_), .ZN(new_n1504_));
  NOR2_X1    g00502(.A1(new_n1504_), .A2(new_n1503_), .ZN(new_n1505_));
  NOR2_X1    g00503(.A1(new_n1502_), .A2(new_n1505_), .ZN(new_n1506_));
  NAND3_X1   g00504(.A1(new_n1499_), .A2(new_n1498_), .A3(new_n1497_), .ZN(new_n1507_));
  OAI21_X1   g00505(.A1(new_n1486_), .A2(new_n1493_), .B(new_n1446_), .ZN(new_n1508_));
  NAND3_X1   g00506(.A1(new_n1506_), .A2(new_n1508_), .A3(new_n1507_), .ZN(new_n1509_));
  NAND3_X1   g00507(.A1(new_n1242_), .A2(new_n1501_), .A3(new_n1509_), .ZN(new_n1510_));
  NOR2_X1    g00508(.A1(new_n1241_), .A2(new_n1229_), .ZN(new_n1511_));
  AOI21_X1   g00509(.A1(new_n1508_), .A2(new_n1507_), .B(new_n1506_), .ZN(new_n1512_));
  NOR3_X1    g00510(.A1(new_n1494_), .A2(new_n1500_), .A3(new_n1409_), .ZN(new_n1513_));
  OAI21_X1   g00511(.A1(new_n1512_), .A2(new_n1513_), .B(new_n1511_), .ZN(new_n1514_));
  NAND2_X1   g00512(.A1(new_n1510_), .A2(new_n1514_), .ZN(new_n1515_));
  NOR2_X1    g00513(.A1(new_n1408_), .A2(new_n1401_), .ZN(new_n1516_));
  NOR2_X1    g00514(.A1(new_n1506_), .A2(new_n1516_), .ZN(new_n1517_));
  INV_X1     g00515(.I(new_n1517_), .ZN(new_n1518_));
  INV_X1     g00516(.I(\A[265] ), .ZN(new_n1519_));
  INV_X1     g00517(.I(\A[266] ), .ZN(new_n1520_));
  NAND2_X1   g00518(.A1(new_n1520_), .A2(\A[267] ), .ZN(new_n1521_));
  INV_X1     g00519(.I(\A[267] ), .ZN(new_n1522_));
  NAND2_X1   g00520(.A1(new_n1522_), .A2(\A[266] ), .ZN(new_n1523_));
  AOI21_X1   g00521(.A1(new_n1521_), .A2(new_n1523_), .B(new_n1519_), .ZN(new_n1524_));
  NAND2_X1   g00522(.A1(\A[266] ), .A2(\A[267] ), .ZN(new_n1525_));
  NOR2_X1    g00523(.A1(\A[266] ), .A2(\A[267] ), .ZN(new_n1526_));
  INV_X1     g00524(.I(new_n1526_), .ZN(new_n1527_));
  AOI21_X1   g00525(.A1(new_n1527_), .A2(new_n1525_), .B(\A[265] ), .ZN(new_n1528_));
  NOR2_X1    g00526(.A1(new_n1528_), .A2(new_n1524_), .ZN(new_n1529_));
  INV_X1     g00527(.I(\A[270] ), .ZN(new_n1530_));
  NOR2_X1    g00528(.A1(new_n1530_), .A2(\A[269] ), .ZN(new_n1531_));
  INV_X1     g00529(.I(\A[269] ), .ZN(new_n1532_));
  NOR2_X1    g00530(.A1(new_n1532_), .A2(\A[270] ), .ZN(new_n1533_));
  OAI21_X1   g00531(.A1(new_n1531_), .A2(new_n1533_), .B(\A[268] ), .ZN(new_n1534_));
  INV_X1     g00532(.I(\A[268] ), .ZN(new_n1535_));
  AND2_X2    g00533(.A1(\A[269] ), .A2(\A[270] ), .Z(new_n1536_));
  NOR2_X1    g00534(.A1(\A[269] ), .A2(\A[270] ), .ZN(new_n1537_));
  OAI21_X1   g00535(.A1(new_n1536_), .A2(new_n1537_), .B(new_n1535_), .ZN(new_n1538_));
  NAND2_X1   g00536(.A1(new_n1534_), .A2(new_n1538_), .ZN(new_n1539_));
  NAND2_X1   g00537(.A1(new_n1529_), .A2(new_n1539_), .ZN(new_n1540_));
  NOR2_X1    g00538(.A1(new_n1522_), .A2(\A[266] ), .ZN(new_n1541_));
  NOR2_X1    g00539(.A1(new_n1520_), .A2(\A[267] ), .ZN(new_n1542_));
  OAI21_X1   g00540(.A1(new_n1541_), .A2(new_n1542_), .B(\A[265] ), .ZN(new_n1543_));
  INV_X1     g00541(.I(new_n1525_), .ZN(new_n1544_));
  OAI21_X1   g00542(.A1(new_n1544_), .A2(new_n1526_), .B(new_n1519_), .ZN(new_n1545_));
  NAND2_X1   g00543(.A1(new_n1543_), .A2(new_n1545_), .ZN(new_n1546_));
  NAND2_X1   g00544(.A1(new_n1532_), .A2(\A[270] ), .ZN(new_n1547_));
  NAND2_X1   g00545(.A1(new_n1530_), .A2(\A[269] ), .ZN(new_n1548_));
  AOI21_X1   g00546(.A1(new_n1547_), .A2(new_n1548_), .B(new_n1535_), .ZN(new_n1549_));
  NAND2_X1   g00547(.A1(\A[269] ), .A2(\A[270] ), .ZN(new_n1550_));
  INV_X1     g00548(.I(new_n1537_), .ZN(new_n1551_));
  AOI21_X1   g00549(.A1(new_n1551_), .A2(new_n1550_), .B(\A[268] ), .ZN(new_n1552_));
  NOR2_X1    g00550(.A1(new_n1552_), .A2(new_n1549_), .ZN(new_n1553_));
  NAND2_X1   g00551(.A1(new_n1553_), .A2(new_n1546_), .ZN(new_n1554_));
  NAND2_X1   g00552(.A1(new_n1554_), .A2(new_n1540_), .ZN(new_n1555_));
  INV_X1     g00553(.I(\A[259] ), .ZN(new_n1556_));
  INV_X1     g00554(.I(\A[260] ), .ZN(new_n1557_));
  NAND2_X1   g00555(.A1(new_n1557_), .A2(\A[261] ), .ZN(new_n1558_));
  INV_X1     g00556(.I(\A[261] ), .ZN(new_n1559_));
  NAND2_X1   g00557(.A1(new_n1559_), .A2(\A[260] ), .ZN(new_n1560_));
  AOI21_X1   g00558(.A1(new_n1558_), .A2(new_n1560_), .B(new_n1556_), .ZN(new_n1561_));
  NAND2_X1   g00559(.A1(\A[260] ), .A2(\A[261] ), .ZN(new_n1562_));
  NOR2_X1    g00560(.A1(\A[260] ), .A2(\A[261] ), .ZN(new_n1563_));
  INV_X1     g00561(.I(new_n1563_), .ZN(new_n1564_));
  AOI21_X1   g00562(.A1(new_n1564_), .A2(new_n1562_), .B(\A[259] ), .ZN(new_n1565_));
  NOR2_X1    g00563(.A1(new_n1565_), .A2(new_n1561_), .ZN(new_n1566_));
  INV_X1     g00564(.I(\A[264] ), .ZN(new_n1567_));
  NOR2_X1    g00565(.A1(new_n1567_), .A2(\A[263] ), .ZN(new_n1568_));
  INV_X1     g00566(.I(\A[263] ), .ZN(new_n1569_));
  NOR2_X1    g00567(.A1(new_n1569_), .A2(\A[264] ), .ZN(new_n1570_));
  OAI21_X1   g00568(.A1(new_n1568_), .A2(new_n1570_), .B(\A[262] ), .ZN(new_n1571_));
  INV_X1     g00569(.I(\A[262] ), .ZN(new_n1572_));
  NAND2_X1   g00570(.A1(\A[263] ), .A2(\A[264] ), .ZN(new_n1573_));
  INV_X1     g00571(.I(new_n1573_), .ZN(new_n1574_));
  NOR2_X1    g00572(.A1(\A[263] ), .A2(\A[264] ), .ZN(new_n1575_));
  OAI21_X1   g00573(.A1(new_n1574_), .A2(new_n1575_), .B(new_n1572_), .ZN(new_n1576_));
  NAND2_X1   g00574(.A1(new_n1571_), .A2(new_n1576_), .ZN(new_n1577_));
  NAND2_X1   g00575(.A1(new_n1566_), .A2(new_n1577_), .ZN(new_n1578_));
  NOR2_X1    g00576(.A1(new_n1559_), .A2(\A[260] ), .ZN(new_n1579_));
  NOR2_X1    g00577(.A1(new_n1557_), .A2(\A[261] ), .ZN(new_n1580_));
  OAI21_X1   g00578(.A1(new_n1579_), .A2(new_n1580_), .B(\A[259] ), .ZN(new_n1581_));
  AND2_X2    g00579(.A1(\A[260] ), .A2(\A[261] ), .Z(new_n1582_));
  OAI21_X1   g00580(.A1(new_n1582_), .A2(new_n1563_), .B(new_n1556_), .ZN(new_n1583_));
  NAND2_X1   g00581(.A1(new_n1581_), .A2(new_n1583_), .ZN(new_n1584_));
  NAND2_X1   g00582(.A1(new_n1569_), .A2(\A[264] ), .ZN(new_n1585_));
  NAND2_X1   g00583(.A1(new_n1567_), .A2(\A[263] ), .ZN(new_n1586_));
  AOI21_X1   g00584(.A1(new_n1585_), .A2(new_n1586_), .B(new_n1572_), .ZN(new_n1587_));
  INV_X1     g00585(.I(new_n1575_), .ZN(new_n1588_));
  AOI21_X1   g00586(.A1(new_n1588_), .A2(new_n1573_), .B(\A[262] ), .ZN(new_n1589_));
  NOR2_X1    g00587(.A1(new_n1589_), .A2(new_n1587_), .ZN(new_n1590_));
  NAND2_X1   g00588(.A1(new_n1590_), .A2(new_n1584_), .ZN(new_n1591_));
  NAND2_X1   g00589(.A1(new_n1578_), .A2(new_n1591_), .ZN(new_n1592_));
  NOR2_X1    g00590(.A1(new_n1555_), .A2(new_n1592_), .ZN(new_n1593_));
  XOR2_X1    g00591(.A1(new_n1529_), .A2(new_n1539_), .Z(new_n1594_));
  NOR2_X1    g00592(.A1(new_n1590_), .A2(new_n1584_), .ZN(new_n1595_));
  NOR2_X1    g00593(.A1(new_n1566_), .A2(new_n1577_), .ZN(new_n1596_));
  NOR2_X1    g00594(.A1(new_n1596_), .A2(new_n1595_), .ZN(new_n1597_));
  NOR2_X1    g00595(.A1(new_n1594_), .A2(new_n1597_), .ZN(new_n1598_));
  INV_X1     g00596(.I(\A[253] ), .ZN(new_n1599_));
  INV_X1     g00597(.I(\A[254] ), .ZN(new_n1600_));
  NAND2_X1   g00598(.A1(new_n1600_), .A2(\A[255] ), .ZN(new_n1601_));
  INV_X1     g00599(.I(\A[255] ), .ZN(new_n1602_));
  NAND2_X1   g00600(.A1(new_n1602_), .A2(\A[254] ), .ZN(new_n1603_));
  AOI21_X1   g00601(.A1(new_n1601_), .A2(new_n1603_), .B(new_n1599_), .ZN(new_n1604_));
  NAND2_X1   g00602(.A1(\A[254] ), .A2(\A[255] ), .ZN(new_n1605_));
  NOR2_X1    g00603(.A1(\A[254] ), .A2(\A[255] ), .ZN(new_n1606_));
  INV_X1     g00604(.I(new_n1606_), .ZN(new_n1607_));
  AOI21_X1   g00605(.A1(new_n1607_), .A2(new_n1605_), .B(\A[253] ), .ZN(new_n1608_));
  NOR2_X1    g00606(.A1(new_n1608_), .A2(new_n1604_), .ZN(new_n1609_));
  INV_X1     g00607(.I(\A[258] ), .ZN(new_n1610_));
  NOR2_X1    g00608(.A1(new_n1610_), .A2(\A[257] ), .ZN(new_n1611_));
  INV_X1     g00609(.I(\A[257] ), .ZN(new_n1612_));
  NOR2_X1    g00610(.A1(new_n1612_), .A2(\A[258] ), .ZN(new_n1613_));
  OAI21_X1   g00611(.A1(new_n1611_), .A2(new_n1613_), .B(\A[256] ), .ZN(new_n1614_));
  INV_X1     g00612(.I(\A[256] ), .ZN(new_n1615_));
  NAND2_X1   g00613(.A1(\A[257] ), .A2(\A[258] ), .ZN(new_n1616_));
  INV_X1     g00614(.I(new_n1616_), .ZN(new_n1617_));
  NOR2_X1    g00615(.A1(\A[257] ), .A2(\A[258] ), .ZN(new_n1618_));
  OAI21_X1   g00616(.A1(new_n1617_), .A2(new_n1618_), .B(new_n1615_), .ZN(new_n1619_));
  NAND2_X1   g00617(.A1(new_n1614_), .A2(new_n1619_), .ZN(new_n1620_));
  NAND2_X1   g00618(.A1(new_n1609_), .A2(new_n1620_), .ZN(new_n1621_));
  NOR2_X1    g00619(.A1(new_n1602_), .A2(\A[254] ), .ZN(new_n1622_));
  NOR2_X1    g00620(.A1(new_n1600_), .A2(\A[255] ), .ZN(new_n1623_));
  OAI21_X1   g00621(.A1(new_n1622_), .A2(new_n1623_), .B(\A[253] ), .ZN(new_n1624_));
  INV_X1     g00622(.I(new_n1605_), .ZN(new_n1625_));
  OAI21_X1   g00623(.A1(new_n1625_), .A2(new_n1606_), .B(new_n1599_), .ZN(new_n1626_));
  NAND2_X1   g00624(.A1(new_n1624_), .A2(new_n1626_), .ZN(new_n1627_));
  NAND2_X1   g00625(.A1(new_n1612_), .A2(\A[258] ), .ZN(new_n1628_));
  NAND2_X1   g00626(.A1(new_n1610_), .A2(\A[257] ), .ZN(new_n1629_));
  AOI21_X1   g00627(.A1(new_n1628_), .A2(new_n1629_), .B(new_n1615_), .ZN(new_n1630_));
  INV_X1     g00628(.I(new_n1618_), .ZN(new_n1631_));
  AOI21_X1   g00629(.A1(new_n1631_), .A2(new_n1616_), .B(\A[256] ), .ZN(new_n1632_));
  NOR2_X1    g00630(.A1(new_n1632_), .A2(new_n1630_), .ZN(new_n1633_));
  NAND2_X1   g00631(.A1(new_n1633_), .A2(new_n1627_), .ZN(new_n1634_));
  INV_X1     g00632(.I(\A[247] ), .ZN(new_n1635_));
  INV_X1     g00633(.I(\A[248] ), .ZN(new_n1636_));
  NAND2_X1   g00634(.A1(new_n1636_), .A2(\A[249] ), .ZN(new_n1637_));
  INV_X1     g00635(.I(\A[249] ), .ZN(new_n1638_));
  NAND2_X1   g00636(.A1(new_n1638_), .A2(\A[248] ), .ZN(new_n1639_));
  AOI21_X1   g00637(.A1(new_n1637_), .A2(new_n1639_), .B(new_n1635_), .ZN(new_n1640_));
  NAND2_X1   g00638(.A1(\A[248] ), .A2(\A[249] ), .ZN(new_n1641_));
  NOR2_X1    g00639(.A1(\A[248] ), .A2(\A[249] ), .ZN(new_n1642_));
  INV_X1     g00640(.I(new_n1642_), .ZN(new_n1643_));
  AOI21_X1   g00641(.A1(new_n1643_), .A2(new_n1641_), .B(\A[247] ), .ZN(new_n1644_));
  NOR2_X1    g00642(.A1(new_n1644_), .A2(new_n1640_), .ZN(new_n1645_));
  INV_X1     g00643(.I(\A[252] ), .ZN(new_n1646_));
  NOR2_X1    g00644(.A1(new_n1646_), .A2(\A[251] ), .ZN(new_n1647_));
  INV_X1     g00645(.I(\A[251] ), .ZN(new_n1648_));
  NOR2_X1    g00646(.A1(new_n1648_), .A2(\A[252] ), .ZN(new_n1649_));
  OAI21_X1   g00647(.A1(new_n1647_), .A2(new_n1649_), .B(\A[250] ), .ZN(new_n1650_));
  INV_X1     g00648(.I(\A[250] ), .ZN(new_n1651_));
  NAND2_X1   g00649(.A1(\A[251] ), .A2(\A[252] ), .ZN(new_n1652_));
  INV_X1     g00650(.I(new_n1652_), .ZN(new_n1653_));
  NOR2_X1    g00651(.A1(\A[251] ), .A2(\A[252] ), .ZN(new_n1654_));
  OAI21_X1   g00652(.A1(new_n1653_), .A2(new_n1654_), .B(new_n1651_), .ZN(new_n1655_));
  NAND2_X1   g00653(.A1(new_n1650_), .A2(new_n1655_), .ZN(new_n1656_));
  NAND2_X1   g00654(.A1(new_n1645_), .A2(new_n1656_), .ZN(new_n1657_));
  NOR2_X1    g00655(.A1(new_n1638_), .A2(\A[248] ), .ZN(new_n1658_));
  NOR2_X1    g00656(.A1(new_n1636_), .A2(\A[249] ), .ZN(new_n1659_));
  OAI21_X1   g00657(.A1(new_n1658_), .A2(new_n1659_), .B(\A[247] ), .ZN(new_n1660_));
  AND2_X2    g00658(.A1(\A[248] ), .A2(\A[249] ), .Z(new_n1661_));
  OAI21_X1   g00659(.A1(new_n1661_), .A2(new_n1642_), .B(new_n1635_), .ZN(new_n1662_));
  NAND2_X1   g00660(.A1(new_n1660_), .A2(new_n1662_), .ZN(new_n1663_));
  NAND2_X1   g00661(.A1(new_n1648_), .A2(\A[252] ), .ZN(new_n1664_));
  NAND2_X1   g00662(.A1(new_n1646_), .A2(\A[251] ), .ZN(new_n1665_));
  AOI21_X1   g00663(.A1(new_n1664_), .A2(new_n1665_), .B(new_n1651_), .ZN(new_n1666_));
  INV_X1     g00664(.I(new_n1654_), .ZN(new_n1667_));
  AOI21_X1   g00665(.A1(new_n1667_), .A2(new_n1652_), .B(\A[250] ), .ZN(new_n1668_));
  NOR2_X1    g00666(.A1(new_n1668_), .A2(new_n1666_), .ZN(new_n1669_));
  NAND2_X1   g00667(.A1(new_n1669_), .A2(new_n1663_), .ZN(new_n1670_));
  AOI22_X1   g00668(.A1(new_n1621_), .A2(new_n1634_), .B1(new_n1657_), .B2(new_n1670_), .ZN(new_n1671_));
  NAND2_X1   g00669(.A1(new_n1634_), .A2(new_n1621_), .ZN(new_n1672_));
  NAND2_X1   g00670(.A1(new_n1657_), .A2(new_n1670_), .ZN(new_n1673_));
  NOR2_X1    g00671(.A1(new_n1672_), .A2(new_n1673_), .ZN(new_n1674_));
  NOR4_X1    g00672(.A1(new_n1598_), .A2(new_n1593_), .A3(new_n1674_), .A4(new_n1671_), .ZN(new_n1675_));
  NAND2_X1   g00673(.A1(new_n1594_), .A2(new_n1597_), .ZN(new_n1676_));
  NAND2_X1   g00674(.A1(new_n1555_), .A2(new_n1592_), .ZN(new_n1677_));
  NAND2_X1   g00675(.A1(new_n1672_), .A2(new_n1673_), .ZN(new_n1678_));
  NOR2_X1    g00676(.A1(new_n1633_), .A2(new_n1627_), .ZN(new_n1679_));
  NOR2_X1    g00677(.A1(new_n1609_), .A2(new_n1620_), .ZN(new_n1680_));
  NOR2_X1    g00678(.A1(new_n1679_), .A2(new_n1680_), .ZN(new_n1681_));
  NOR2_X1    g00679(.A1(new_n1669_), .A2(new_n1663_), .ZN(new_n1682_));
  NOR2_X1    g00680(.A1(new_n1645_), .A2(new_n1656_), .ZN(new_n1683_));
  NOR2_X1    g00681(.A1(new_n1683_), .A2(new_n1682_), .ZN(new_n1684_));
  NAND2_X1   g00682(.A1(new_n1681_), .A2(new_n1684_), .ZN(new_n1685_));
  AOI22_X1   g00683(.A1(new_n1676_), .A2(new_n1677_), .B1(new_n1685_), .B2(new_n1678_), .ZN(new_n1686_));
  NOR2_X1    g00684(.A1(new_n1686_), .A2(new_n1675_), .ZN(new_n1687_));
  INV_X1     g00685(.I(\A[231] ), .ZN(new_n1688_));
  NOR2_X1    g00686(.A1(new_n1688_), .A2(\A[230] ), .ZN(new_n1689_));
  INV_X1     g00687(.I(\A[230] ), .ZN(new_n1690_));
  NOR2_X1    g00688(.A1(new_n1690_), .A2(\A[231] ), .ZN(new_n1691_));
  OAI21_X1   g00689(.A1(new_n1689_), .A2(new_n1691_), .B(\A[229] ), .ZN(new_n1692_));
  INV_X1     g00690(.I(\A[229] ), .ZN(new_n1693_));
  NOR2_X1    g00691(.A1(\A[230] ), .A2(\A[231] ), .ZN(new_n1694_));
  NAND2_X1   g00692(.A1(\A[230] ), .A2(\A[231] ), .ZN(new_n1695_));
  INV_X1     g00693(.I(new_n1695_), .ZN(new_n1696_));
  OAI21_X1   g00694(.A1(new_n1696_), .A2(new_n1694_), .B(new_n1693_), .ZN(new_n1697_));
  INV_X1     g00695(.I(\A[234] ), .ZN(new_n1698_));
  NOR2_X1    g00696(.A1(new_n1698_), .A2(\A[233] ), .ZN(new_n1699_));
  INV_X1     g00697(.I(\A[233] ), .ZN(new_n1700_));
  NOR2_X1    g00698(.A1(new_n1700_), .A2(\A[234] ), .ZN(new_n1701_));
  OAI21_X1   g00699(.A1(new_n1699_), .A2(new_n1701_), .B(\A[232] ), .ZN(new_n1702_));
  INV_X1     g00700(.I(\A[232] ), .ZN(new_n1703_));
  NOR2_X1    g00701(.A1(\A[233] ), .A2(\A[234] ), .ZN(new_n1704_));
  AND2_X2    g00702(.A1(\A[233] ), .A2(\A[234] ), .Z(new_n1705_));
  OAI21_X1   g00703(.A1(new_n1705_), .A2(new_n1704_), .B(new_n1703_), .ZN(new_n1706_));
  NAND4_X1   g00704(.A1(new_n1692_), .A2(new_n1702_), .A3(new_n1697_), .A4(new_n1706_), .ZN(new_n1707_));
  NAND2_X1   g00705(.A1(new_n1690_), .A2(\A[231] ), .ZN(new_n1708_));
  NAND2_X1   g00706(.A1(new_n1688_), .A2(\A[230] ), .ZN(new_n1709_));
  AOI21_X1   g00707(.A1(new_n1708_), .A2(new_n1709_), .B(new_n1693_), .ZN(new_n1710_));
  INV_X1     g00708(.I(new_n1694_), .ZN(new_n1711_));
  AOI21_X1   g00709(.A1(new_n1711_), .A2(new_n1695_), .B(\A[229] ), .ZN(new_n1712_));
  NAND2_X1   g00710(.A1(new_n1700_), .A2(\A[234] ), .ZN(new_n1713_));
  NAND2_X1   g00711(.A1(new_n1698_), .A2(\A[233] ), .ZN(new_n1714_));
  AOI21_X1   g00712(.A1(new_n1713_), .A2(new_n1714_), .B(new_n1703_), .ZN(new_n1715_));
  INV_X1     g00713(.I(new_n1704_), .ZN(new_n1716_));
  NAND2_X1   g00714(.A1(\A[233] ), .A2(\A[234] ), .ZN(new_n1717_));
  AOI21_X1   g00715(.A1(new_n1716_), .A2(new_n1717_), .B(\A[232] ), .ZN(new_n1718_));
  OAI22_X1   g00716(.A1(new_n1710_), .A2(new_n1712_), .B1(new_n1718_), .B2(new_n1715_), .ZN(new_n1719_));
  NAND2_X1   g00717(.A1(new_n1719_), .A2(new_n1707_), .ZN(new_n1720_));
  INV_X1     g00718(.I(\A[223] ), .ZN(new_n1721_));
  INV_X1     g00719(.I(\A[224] ), .ZN(new_n1722_));
  NAND2_X1   g00720(.A1(new_n1722_), .A2(\A[225] ), .ZN(new_n1723_));
  INV_X1     g00721(.I(\A[225] ), .ZN(new_n1724_));
  NAND2_X1   g00722(.A1(new_n1724_), .A2(\A[224] ), .ZN(new_n1725_));
  AOI21_X1   g00723(.A1(new_n1723_), .A2(new_n1725_), .B(new_n1721_), .ZN(new_n1726_));
  NAND2_X1   g00724(.A1(\A[224] ), .A2(\A[225] ), .ZN(new_n1727_));
  NOR2_X1    g00725(.A1(\A[224] ), .A2(\A[225] ), .ZN(new_n1728_));
  INV_X1     g00726(.I(new_n1728_), .ZN(new_n1729_));
  AOI21_X1   g00727(.A1(new_n1729_), .A2(new_n1727_), .B(\A[223] ), .ZN(new_n1730_));
  INV_X1     g00728(.I(\A[226] ), .ZN(new_n1731_));
  INV_X1     g00729(.I(\A[227] ), .ZN(new_n1732_));
  NAND2_X1   g00730(.A1(new_n1732_), .A2(\A[228] ), .ZN(new_n1733_));
  INV_X1     g00731(.I(\A[228] ), .ZN(new_n1734_));
  NAND2_X1   g00732(.A1(new_n1734_), .A2(\A[227] ), .ZN(new_n1735_));
  AOI21_X1   g00733(.A1(new_n1733_), .A2(new_n1735_), .B(new_n1731_), .ZN(new_n1736_));
  NAND2_X1   g00734(.A1(\A[227] ), .A2(\A[228] ), .ZN(new_n1737_));
  OR2_X2     g00735(.A1(\A[227] ), .A2(\A[228] ), .Z(new_n1738_));
  AOI21_X1   g00736(.A1(new_n1738_), .A2(new_n1737_), .B(\A[226] ), .ZN(new_n1739_));
  NOR4_X1    g00737(.A1(new_n1726_), .A2(new_n1730_), .A3(new_n1736_), .A4(new_n1739_), .ZN(new_n1740_));
  NOR2_X1    g00738(.A1(new_n1724_), .A2(\A[224] ), .ZN(new_n1741_));
  NOR2_X1    g00739(.A1(new_n1722_), .A2(\A[225] ), .ZN(new_n1742_));
  OAI21_X1   g00740(.A1(new_n1741_), .A2(new_n1742_), .B(\A[223] ), .ZN(new_n1743_));
  INV_X1     g00741(.I(new_n1727_), .ZN(new_n1744_));
  OAI21_X1   g00742(.A1(new_n1744_), .A2(new_n1728_), .B(new_n1721_), .ZN(new_n1745_));
  NOR2_X1    g00743(.A1(new_n1734_), .A2(\A[227] ), .ZN(new_n1746_));
  NOR2_X1    g00744(.A1(new_n1732_), .A2(\A[228] ), .ZN(new_n1747_));
  OAI21_X1   g00745(.A1(new_n1746_), .A2(new_n1747_), .B(\A[226] ), .ZN(new_n1748_));
  INV_X1     g00746(.I(new_n1737_), .ZN(new_n1749_));
  NOR2_X1    g00747(.A1(\A[227] ), .A2(\A[228] ), .ZN(new_n1750_));
  OAI21_X1   g00748(.A1(new_n1749_), .A2(new_n1750_), .B(new_n1731_), .ZN(new_n1751_));
  AOI22_X1   g00749(.A1(new_n1743_), .A2(new_n1745_), .B1(new_n1748_), .B2(new_n1751_), .ZN(new_n1752_));
  NOR2_X1    g00750(.A1(new_n1752_), .A2(new_n1740_), .ZN(new_n1753_));
  NAND2_X1   g00751(.A1(new_n1753_), .A2(new_n1720_), .ZN(new_n1754_));
  NOR4_X1    g00752(.A1(new_n1710_), .A2(new_n1712_), .A3(new_n1718_), .A4(new_n1715_), .ZN(new_n1755_));
  AOI22_X1   g00753(.A1(new_n1692_), .A2(new_n1697_), .B1(new_n1702_), .B2(new_n1706_), .ZN(new_n1756_));
  NOR2_X1    g00754(.A1(new_n1755_), .A2(new_n1756_), .ZN(new_n1757_));
  NAND4_X1   g00755(.A1(new_n1743_), .A2(new_n1745_), .A3(new_n1748_), .A4(new_n1751_), .ZN(new_n1758_));
  OAI22_X1   g00756(.A1(new_n1726_), .A2(new_n1730_), .B1(new_n1736_), .B2(new_n1739_), .ZN(new_n1759_));
  NAND2_X1   g00757(.A1(new_n1758_), .A2(new_n1759_), .ZN(new_n1760_));
  NAND2_X1   g00758(.A1(new_n1757_), .A2(new_n1760_), .ZN(new_n1761_));
  NAND2_X1   g00759(.A1(new_n1761_), .A2(new_n1754_), .ZN(new_n1762_));
  INV_X1     g00760(.I(\A[235] ), .ZN(new_n1763_));
  INV_X1     g00761(.I(\A[236] ), .ZN(new_n1764_));
  NAND2_X1   g00762(.A1(new_n1764_), .A2(\A[237] ), .ZN(new_n1765_));
  INV_X1     g00763(.I(\A[237] ), .ZN(new_n1766_));
  NAND2_X1   g00764(.A1(new_n1766_), .A2(\A[236] ), .ZN(new_n1767_));
  AOI21_X1   g00765(.A1(new_n1765_), .A2(new_n1767_), .B(new_n1763_), .ZN(new_n1768_));
  NAND2_X1   g00766(.A1(\A[236] ), .A2(\A[237] ), .ZN(new_n1769_));
  NOR2_X1    g00767(.A1(\A[236] ), .A2(\A[237] ), .ZN(new_n1770_));
  INV_X1     g00768(.I(new_n1770_), .ZN(new_n1771_));
  AOI21_X1   g00769(.A1(new_n1771_), .A2(new_n1769_), .B(\A[235] ), .ZN(new_n1772_));
  INV_X1     g00770(.I(\A[238] ), .ZN(new_n1773_));
  INV_X1     g00771(.I(\A[239] ), .ZN(new_n1774_));
  NAND2_X1   g00772(.A1(new_n1774_), .A2(\A[240] ), .ZN(new_n1775_));
  INV_X1     g00773(.I(\A[240] ), .ZN(new_n1776_));
  NAND2_X1   g00774(.A1(new_n1776_), .A2(\A[239] ), .ZN(new_n1777_));
  AOI21_X1   g00775(.A1(new_n1775_), .A2(new_n1777_), .B(new_n1773_), .ZN(new_n1778_));
  NAND2_X1   g00776(.A1(\A[239] ), .A2(\A[240] ), .ZN(new_n1779_));
  NOR2_X1    g00777(.A1(\A[239] ), .A2(\A[240] ), .ZN(new_n1780_));
  INV_X1     g00778(.I(new_n1780_), .ZN(new_n1781_));
  AOI21_X1   g00779(.A1(new_n1781_), .A2(new_n1779_), .B(\A[238] ), .ZN(new_n1782_));
  NOR4_X1    g00780(.A1(new_n1768_), .A2(new_n1772_), .A3(new_n1782_), .A4(new_n1778_), .ZN(new_n1783_));
  NOR2_X1    g00781(.A1(new_n1766_), .A2(\A[236] ), .ZN(new_n1784_));
  NOR2_X1    g00782(.A1(new_n1764_), .A2(\A[237] ), .ZN(new_n1785_));
  OAI21_X1   g00783(.A1(new_n1784_), .A2(new_n1785_), .B(\A[235] ), .ZN(new_n1786_));
  INV_X1     g00784(.I(new_n1769_), .ZN(new_n1787_));
  OAI21_X1   g00785(.A1(new_n1787_), .A2(new_n1770_), .B(new_n1763_), .ZN(new_n1788_));
  NOR2_X1    g00786(.A1(new_n1776_), .A2(\A[239] ), .ZN(new_n1789_));
  NOR2_X1    g00787(.A1(new_n1774_), .A2(\A[240] ), .ZN(new_n1790_));
  OAI21_X1   g00788(.A1(new_n1789_), .A2(new_n1790_), .B(\A[238] ), .ZN(new_n1791_));
  AND2_X2    g00789(.A1(\A[239] ), .A2(\A[240] ), .Z(new_n1792_));
  OAI21_X1   g00790(.A1(new_n1792_), .A2(new_n1780_), .B(new_n1773_), .ZN(new_n1793_));
  AOI22_X1   g00791(.A1(new_n1786_), .A2(new_n1788_), .B1(new_n1791_), .B2(new_n1793_), .ZN(new_n1794_));
  INV_X1     g00792(.I(\A[241] ), .ZN(new_n1795_));
  INV_X1     g00793(.I(\A[242] ), .ZN(new_n1796_));
  NAND2_X1   g00794(.A1(new_n1796_), .A2(\A[243] ), .ZN(new_n1797_));
  INV_X1     g00795(.I(\A[243] ), .ZN(new_n1798_));
  NAND2_X1   g00796(.A1(new_n1798_), .A2(\A[242] ), .ZN(new_n1799_));
  AOI21_X1   g00797(.A1(new_n1797_), .A2(new_n1799_), .B(new_n1795_), .ZN(new_n1800_));
  NAND2_X1   g00798(.A1(\A[242] ), .A2(\A[243] ), .ZN(new_n1801_));
  NOR2_X1    g00799(.A1(\A[242] ), .A2(\A[243] ), .ZN(new_n1802_));
  INV_X1     g00800(.I(new_n1802_), .ZN(new_n1803_));
  AOI21_X1   g00801(.A1(new_n1803_), .A2(new_n1801_), .B(\A[241] ), .ZN(new_n1804_));
  INV_X1     g00802(.I(\A[244] ), .ZN(new_n1805_));
  INV_X1     g00803(.I(\A[245] ), .ZN(new_n1806_));
  NAND2_X1   g00804(.A1(new_n1806_), .A2(\A[246] ), .ZN(new_n1807_));
  INV_X1     g00805(.I(\A[246] ), .ZN(new_n1808_));
  NAND2_X1   g00806(.A1(new_n1808_), .A2(\A[245] ), .ZN(new_n1809_));
  AOI21_X1   g00807(.A1(new_n1807_), .A2(new_n1809_), .B(new_n1805_), .ZN(new_n1810_));
  NAND2_X1   g00808(.A1(\A[245] ), .A2(\A[246] ), .ZN(new_n1811_));
  NOR2_X1    g00809(.A1(\A[245] ), .A2(\A[246] ), .ZN(new_n1812_));
  INV_X1     g00810(.I(new_n1812_), .ZN(new_n1813_));
  AOI21_X1   g00811(.A1(new_n1813_), .A2(new_n1811_), .B(\A[244] ), .ZN(new_n1814_));
  NOR4_X1    g00812(.A1(new_n1800_), .A2(new_n1804_), .A3(new_n1814_), .A4(new_n1810_), .ZN(new_n1815_));
  NOR2_X1    g00813(.A1(new_n1798_), .A2(\A[242] ), .ZN(new_n1816_));
  NOR2_X1    g00814(.A1(new_n1796_), .A2(\A[243] ), .ZN(new_n1817_));
  OAI21_X1   g00815(.A1(new_n1816_), .A2(new_n1817_), .B(\A[241] ), .ZN(new_n1818_));
  INV_X1     g00816(.I(new_n1801_), .ZN(new_n1819_));
  OAI21_X1   g00817(.A1(new_n1819_), .A2(new_n1802_), .B(new_n1795_), .ZN(new_n1820_));
  NOR2_X1    g00818(.A1(new_n1808_), .A2(\A[245] ), .ZN(new_n1821_));
  NOR2_X1    g00819(.A1(new_n1806_), .A2(\A[246] ), .ZN(new_n1822_));
  OAI21_X1   g00820(.A1(new_n1821_), .A2(new_n1822_), .B(\A[244] ), .ZN(new_n1823_));
  AND2_X2    g00821(.A1(\A[245] ), .A2(\A[246] ), .Z(new_n1824_));
  OAI21_X1   g00822(.A1(new_n1824_), .A2(new_n1812_), .B(new_n1805_), .ZN(new_n1825_));
  AOI22_X1   g00823(.A1(new_n1818_), .A2(new_n1820_), .B1(new_n1823_), .B2(new_n1825_), .ZN(new_n1826_));
  OAI22_X1   g00824(.A1(new_n1783_), .A2(new_n1794_), .B1(new_n1815_), .B2(new_n1826_), .ZN(new_n1827_));
  NAND4_X1   g00825(.A1(new_n1786_), .A2(new_n1791_), .A3(new_n1788_), .A4(new_n1793_), .ZN(new_n1828_));
  OAI22_X1   g00826(.A1(new_n1768_), .A2(new_n1772_), .B1(new_n1782_), .B2(new_n1778_), .ZN(new_n1829_));
  NAND4_X1   g00827(.A1(new_n1818_), .A2(new_n1823_), .A3(new_n1820_), .A4(new_n1825_), .ZN(new_n1830_));
  OAI22_X1   g00828(.A1(new_n1800_), .A2(new_n1804_), .B1(new_n1814_), .B2(new_n1810_), .ZN(new_n1831_));
  NAND4_X1   g00829(.A1(new_n1829_), .A2(new_n1831_), .A3(new_n1828_), .A4(new_n1830_), .ZN(new_n1832_));
  NAND2_X1   g00830(.A1(new_n1827_), .A2(new_n1832_), .ZN(new_n1833_));
  INV_X1     g00831(.I(new_n1833_), .ZN(new_n1834_));
  NOR2_X1    g00832(.A1(new_n1834_), .A2(new_n1762_), .ZN(new_n1835_));
  AOI21_X1   g00833(.A1(new_n1754_), .A2(new_n1761_), .B(new_n1833_), .ZN(new_n1836_));
  NOR2_X1    g00834(.A1(new_n1835_), .A2(new_n1836_), .ZN(new_n1837_));
  NAND2_X1   g00835(.A1(new_n1687_), .A2(new_n1837_), .ZN(new_n1838_));
  NOR2_X1    g00836(.A1(new_n1687_), .A2(new_n1837_), .ZN(new_n1839_));
  INV_X1     g00837(.I(new_n1839_), .ZN(new_n1840_));
  NAND2_X1   g00838(.A1(new_n1840_), .A2(new_n1838_), .ZN(new_n1841_));
  NOR2_X1    g00839(.A1(new_n1518_), .A2(new_n1841_), .ZN(new_n1842_));
  AOI21_X1   g00840(.A1(\A[239] ), .A2(\A[240] ), .B(\A[238] ), .ZN(new_n1843_));
  NOR2_X1    g00841(.A1(new_n1843_), .A2(new_n1780_), .ZN(new_n1844_));
  AOI21_X1   g00842(.A1(\A[236] ), .A2(\A[237] ), .B(\A[235] ), .ZN(new_n1845_));
  NOR2_X1    g00843(.A1(new_n1845_), .A2(new_n1770_), .ZN(new_n1846_));
  NOR2_X1    g00844(.A1(new_n1844_), .A2(new_n1846_), .ZN(new_n1847_));
  NOR4_X1    g00845(.A1(new_n1843_), .A2(new_n1845_), .A3(new_n1770_), .A4(new_n1780_), .ZN(new_n1848_));
  NOR2_X1    g00846(.A1(new_n1847_), .A2(new_n1848_), .ZN(new_n1849_));
  NAND2_X1   g00847(.A1(new_n1828_), .A2(new_n1849_), .ZN(new_n1850_));
  OAI22_X1   g00848(.A1(new_n1770_), .A2(new_n1845_), .B1(new_n1843_), .B2(new_n1780_), .ZN(new_n1851_));
  INV_X1     g00849(.I(new_n1848_), .ZN(new_n1852_));
  NAND2_X1   g00850(.A1(new_n1852_), .A2(new_n1851_), .ZN(new_n1853_));
  NAND2_X1   g00851(.A1(new_n1783_), .A2(new_n1853_), .ZN(new_n1854_));
  NAND2_X1   g00852(.A1(new_n1854_), .A2(new_n1850_), .ZN(new_n1855_));
  NOR4_X1    g00853(.A1(new_n1783_), .A2(new_n1794_), .A3(new_n1815_), .A4(new_n1826_), .ZN(new_n1856_));
  NAND2_X1   g00854(.A1(new_n1818_), .A2(new_n1820_), .ZN(new_n1857_));
  NAND2_X1   g00855(.A1(new_n1823_), .A2(new_n1825_), .ZN(new_n1858_));
  AOI21_X1   g00856(.A1(\A[245] ), .A2(\A[246] ), .B(\A[244] ), .ZN(new_n1859_));
  AOI21_X1   g00857(.A1(\A[242] ), .A2(\A[243] ), .B(\A[241] ), .ZN(new_n1860_));
  NOR2_X1    g00858(.A1(new_n1860_), .A2(new_n1802_), .ZN(new_n1861_));
  NOR3_X1    g00859(.A1(new_n1861_), .A2(new_n1812_), .A3(new_n1859_), .ZN(new_n1862_));
  NOR2_X1    g00860(.A1(new_n1859_), .A2(new_n1812_), .ZN(new_n1863_));
  NOR3_X1    g00861(.A1(new_n1863_), .A2(new_n1802_), .A3(new_n1860_), .ZN(new_n1864_));
  OAI22_X1   g00862(.A1(new_n1857_), .A2(new_n1858_), .B1(new_n1862_), .B2(new_n1864_), .ZN(new_n1865_));
  NOR2_X1    g00863(.A1(new_n1862_), .A2(new_n1864_), .ZN(new_n1866_));
  NAND2_X1   g00864(.A1(new_n1815_), .A2(new_n1866_), .ZN(new_n1867_));
  NAND2_X1   g00865(.A1(new_n1867_), .A2(new_n1865_), .ZN(new_n1868_));
  NOR2_X1    g00866(.A1(new_n1868_), .A2(new_n1856_), .ZN(new_n1869_));
  NOR2_X1    g00867(.A1(new_n1804_), .A2(new_n1800_), .ZN(new_n1870_));
  NOR2_X1    g00868(.A1(new_n1814_), .A2(new_n1810_), .ZN(new_n1871_));
  OAI21_X1   g00869(.A1(new_n1802_), .A2(new_n1860_), .B(new_n1863_), .ZN(new_n1872_));
  OAI21_X1   g00870(.A1(new_n1812_), .A2(new_n1859_), .B(new_n1861_), .ZN(new_n1873_));
  AOI22_X1   g00871(.A1(new_n1870_), .A2(new_n1871_), .B1(new_n1872_), .B2(new_n1873_), .ZN(new_n1874_));
  NOR4_X1    g00872(.A1(new_n1857_), .A2(new_n1858_), .A3(new_n1862_), .A4(new_n1864_), .ZN(new_n1875_));
  NOR2_X1    g00873(.A1(new_n1874_), .A2(new_n1875_), .ZN(new_n1876_));
  NOR2_X1    g00874(.A1(new_n1876_), .A2(new_n1832_), .ZN(new_n1877_));
  OR3_X2     g00875(.A1(new_n1869_), .A2(new_n1877_), .A3(new_n1855_), .Z(new_n1878_));
  NOR2_X1    g00876(.A1(new_n1783_), .A2(new_n1794_), .ZN(new_n1879_));
  NAND2_X1   g00877(.A1(new_n1863_), .A2(new_n1861_), .ZN(new_n1880_));
  INV_X1     g00878(.I(new_n1880_), .ZN(new_n1881_));
  NAND2_X1   g00879(.A1(new_n1831_), .A2(new_n1881_), .ZN(new_n1882_));
  NOR3_X1    g00880(.A1(new_n1866_), .A2(new_n1815_), .A3(new_n1826_), .ZN(new_n1883_));
  AND3_X2    g00881(.A1(new_n1883_), .A2(new_n1879_), .A3(new_n1882_), .Z(new_n1884_));
  OAI21_X1   g00882(.A1(new_n1884_), .A2(new_n1869_), .B(new_n1855_), .ZN(new_n1885_));
  NAND2_X1   g00883(.A1(new_n1878_), .A2(new_n1885_), .ZN(new_n1886_));
  AOI21_X1   g00884(.A1(\A[227] ), .A2(\A[228] ), .B(\A[226] ), .ZN(new_n1887_));
  NOR2_X1    g00885(.A1(new_n1887_), .A2(new_n1750_), .ZN(new_n1888_));
  AOI21_X1   g00886(.A1(\A[224] ), .A2(\A[225] ), .B(\A[223] ), .ZN(new_n1889_));
  NOR2_X1    g00887(.A1(new_n1889_), .A2(new_n1728_), .ZN(new_n1890_));
  NOR2_X1    g00888(.A1(new_n1888_), .A2(new_n1890_), .ZN(new_n1891_));
  NOR4_X1    g00889(.A1(new_n1887_), .A2(new_n1889_), .A3(new_n1728_), .A4(new_n1750_), .ZN(new_n1892_));
  NOR2_X1    g00890(.A1(new_n1891_), .A2(new_n1892_), .ZN(new_n1893_));
  NAND2_X1   g00891(.A1(new_n1758_), .A2(new_n1893_), .ZN(new_n1894_));
  NOR2_X1    g00892(.A1(new_n1730_), .A2(new_n1726_), .ZN(new_n1895_));
  NOR2_X1    g00893(.A1(new_n1736_), .A2(new_n1739_), .ZN(new_n1896_));
  OAI22_X1   g00894(.A1(new_n1728_), .A2(new_n1889_), .B1(new_n1887_), .B2(new_n1750_), .ZN(new_n1897_));
  NAND2_X1   g00895(.A1(new_n1888_), .A2(new_n1890_), .ZN(new_n1898_));
  NAND2_X1   g00896(.A1(new_n1898_), .A2(new_n1897_), .ZN(new_n1899_));
  NAND3_X1   g00897(.A1(new_n1899_), .A2(new_n1895_), .A3(new_n1896_), .ZN(new_n1900_));
  NAND2_X1   g00898(.A1(new_n1894_), .A2(new_n1900_), .ZN(new_n1901_));
  AOI21_X1   g00899(.A1(\A[233] ), .A2(\A[234] ), .B(\A[232] ), .ZN(new_n1902_));
  NOR2_X1    g00900(.A1(new_n1902_), .A2(new_n1704_), .ZN(new_n1903_));
  AOI21_X1   g00901(.A1(\A[230] ), .A2(\A[231] ), .B(\A[229] ), .ZN(new_n1904_));
  NOR2_X1    g00902(.A1(new_n1904_), .A2(new_n1694_), .ZN(new_n1905_));
  XOR2_X1    g00903(.A1(new_n1903_), .A2(new_n1905_), .Z(new_n1906_));
  NOR2_X1    g00904(.A1(new_n1906_), .A2(new_n1755_), .ZN(new_n1907_));
  NOR3_X1    g00905(.A1(new_n1905_), .A2(new_n1704_), .A3(new_n1902_), .ZN(new_n1908_));
  NOR3_X1    g00906(.A1(new_n1903_), .A2(new_n1694_), .A3(new_n1904_), .ZN(new_n1909_));
  NOR2_X1    g00907(.A1(new_n1908_), .A2(new_n1909_), .ZN(new_n1910_));
  NOR2_X1    g00908(.A1(new_n1910_), .A2(new_n1707_), .ZN(new_n1911_));
  OAI22_X1   g00909(.A1(new_n1907_), .A2(new_n1911_), .B1(new_n1760_), .B2(new_n1720_), .ZN(new_n1912_));
  NOR3_X1    g00910(.A1(new_n1755_), .A2(new_n1910_), .A3(new_n1756_), .ZN(new_n1913_));
  NOR2_X1    g00911(.A1(new_n1903_), .A2(new_n1905_), .ZN(new_n1914_));
  INV_X1     g00912(.I(new_n1914_), .ZN(new_n1915_));
  NAND2_X1   g00913(.A1(new_n1903_), .A2(new_n1905_), .ZN(new_n1916_));
  NAND2_X1   g00914(.A1(new_n1707_), .A2(new_n1916_), .ZN(new_n1917_));
  NAND2_X1   g00915(.A1(new_n1917_), .A2(new_n1915_), .ZN(new_n1918_));
  NAND3_X1   g00916(.A1(new_n1918_), .A2(new_n1753_), .A3(new_n1913_), .ZN(new_n1919_));
  NAND3_X1   g00917(.A1(new_n1919_), .A2(new_n1912_), .A3(new_n1901_), .ZN(new_n1920_));
  NOR2_X1    g00918(.A1(new_n1740_), .A2(new_n1899_), .ZN(new_n1921_));
  NOR2_X1    g00919(.A1(new_n1758_), .A2(new_n1893_), .ZN(new_n1922_));
  NOR2_X1    g00920(.A1(new_n1922_), .A2(new_n1921_), .ZN(new_n1923_));
  NAND2_X1   g00921(.A1(new_n1910_), .A2(new_n1707_), .ZN(new_n1924_));
  NAND2_X1   g00922(.A1(new_n1906_), .A2(new_n1755_), .ZN(new_n1925_));
  AOI22_X1   g00923(.A1(new_n1924_), .A2(new_n1925_), .B1(new_n1757_), .B2(new_n1753_), .ZN(new_n1926_));
  NOR4_X1    g00924(.A1(new_n1760_), .A2(new_n1755_), .A3(new_n1756_), .A4(new_n1910_), .ZN(new_n1927_));
  OAI21_X1   g00925(.A1(new_n1926_), .A2(new_n1927_), .B(new_n1923_), .ZN(new_n1928_));
  NAND3_X1   g00926(.A1(new_n1836_), .A2(new_n1920_), .A3(new_n1928_), .ZN(new_n1929_));
  AND2_X2    g00927(.A1(new_n1761_), .A2(new_n1754_), .Z(new_n1930_));
  NAND3_X1   g00928(.A1(new_n1906_), .A2(new_n1719_), .A3(new_n1707_), .ZN(new_n1931_));
  AOI21_X1   g00929(.A1(new_n1707_), .A2(new_n1916_), .B(new_n1914_), .ZN(new_n1932_));
  NOR3_X1    g00930(.A1(new_n1931_), .A2(new_n1760_), .A3(new_n1932_), .ZN(new_n1933_));
  NOR3_X1    g00931(.A1(new_n1926_), .A2(new_n1923_), .A3(new_n1933_), .ZN(new_n1934_));
  NOR4_X1    g00932(.A1(new_n1755_), .A2(new_n1752_), .A3(new_n1756_), .A4(new_n1740_), .ZN(new_n1935_));
  NAND3_X1   g00933(.A1(new_n1935_), .A2(new_n1924_), .A3(new_n1925_), .ZN(new_n1936_));
  AOI21_X1   g00934(.A1(new_n1936_), .A2(new_n1912_), .B(new_n1901_), .ZN(new_n1937_));
  OAI22_X1   g00935(.A1(new_n1937_), .A2(new_n1934_), .B1(new_n1930_), .B2(new_n1833_), .ZN(new_n1938_));
  NAND3_X1   g00936(.A1(new_n1886_), .A2(new_n1929_), .A3(new_n1938_), .ZN(new_n1939_));
  NOR3_X1    g00937(.A1(new_n1869_), .A2(new_n1877_), .A3(new_n1855_), .ZN(new_n1940_));
  INV_X1     g00938(.I(new_n1855_), .ZN(new_n1941_));
  NAND2_X1   g00939(.A1(new_n1876_), .A2(new_n1832_), .ZN(new_n1942_));
  NAND4_X1   g00940(.A1(new_n1883_), .A2(new_n1828_), .A3(new_n1882_), .A4(new_n1829_), .ZN(new_n1943_));
  AOI21_X1   g00941(.A1(new_n1942_), .A2(new_n1943_), .B(new_n1941_), .ZN(new_n1944_));
  NOR2_X1    g00942(.A1(new_n1940_), .A2(new_n1944_), .ZN(new_n1945_));
  NOR4_X1    g00943(.A1(new_n1937_), .A2(new_n1934_), .A3(new_n1930_), .A4(new_n1833_), .ZN(new_n1946_));
  AOI21_X1   g00944(.A1(new_n1920_), .A2(new_n1928_), .B(new_n1836_), .ZN(new_n1947_));
  OAI21_X1   g00945(.A1(new_n1947_), .A2(new_n1946_), .B(new_n1945_), .ZN(new_n1948_));
  NAND2_X1   g00946(.A1(new_n1939_), .A2(new_n1948_), .ZN(new_n1949_));
  INV_X1     g00947(.I(new_n1838_), .ZN(new_n1950_));
  NAND4_X1   g00948(.A1(new_n1660_), .A2(new_n1650_), .A3(new_n1655_), .A4(new_n1662_), .ZN(new_n1951_));
  AOI21_X1   g00949(.A1(\A[251] ), .A2(\A[252] ), .B(\A[250] ), .ZN(new_n1952_));
  AOI21_X1   g00950(.A1(\A[248] ), .A2(\A[249] ), .B(\A[247] ), .ZN(new_n1953_));
  OAI22_X1   g00951(.A1(new_n1642_), .A2(new_n1953_), .B1(new_n1952_), .B2(new_n1654_), .ZN(new_n1954_));
  NOR4_X1    g00952(.A1(new_n1952_), .A2(new_n1953_), .A3(new_n1642_), .A4(new_n1654_), .ZN(new_n1955_));
  INV_X1     g00953(.I(new_n1955_), .ZN(new_n1956_));
  NAND2_X1   g00954(.A1(new_n1956_), .A2(new_n1954_), .ZN(new_n1957_));
  XOR2_X1    g00955(.A1(new_n1957_), .A2(new_n1951_), .Z(new_n1958_));
  NOR4_X1    g00956(.A1(new_n1604_), .A2(new_n1608_), .A3(new_n1632_), .A4(new_n1630_), .ZN(new_n1959_));
  AOI21_X1   g00957(.A1(\A[257] ), .A2(\A[258] ), .B(\A[256] ), .ZN(new_n1960_));
  NOR2_X1    g00958(.A1(new_n1960_), .A2(new_n1618_), .ZN(new_n1961_));
  AOI21_X1   g00959(.A1(\A[254] ), .A2(\A[255] ), .B(\A[253] ), .ZN(new_n1962_));
  NOR2_X1    g00960(.A1(new_n1962_), .A2(new_n1606_), .ZN(new_n1963_));
  XOR2_X1    g00961(.A1(new_n1963_), .A2(new_n1961_), .Z(new_n1964_));
  NOR2_X1    g00962(.A1(new_n1964_), .A2(new_n1959_), .ZN(new_n1965_));
  NAND4_X1   g00963(.A1(new_n1624_), .A2(new_n1626_), .A3(new_n1614_), .A4(new_n1619_), .ZN(new_n1966_));
  NOR3_X1    g00964(.A1(new_n1963_), .A2(new_n1618_), .A3(new_n1960_), .ZN(new_n1967_));
  NOR3_X1    g00965(.A1(new_n1961_), .A2(new_n1606_), .A3(new_n1962_), .ZN(new_n1968_));
  NOR2_X1    g00966(.A1(new_n1967_), .A2(new_n1968_), .ZN(new_n1969_));
  NOR2_X1    g00967(.A1(new_n1966_), .A2(new_n1969_), .ZN(new_n1970_));
  NOR2_X1    g00968(.A1(new_n1965_), .A2(new_n1970_), .ZN(new_n1971_));
  OAI21_X1   g00969(.A1(new_n1671_), .A2(new_n1971_), .B(new_n1958_), .ZN(new_n1972_));
  NAND2_X1   g00970(.A1(new_n1966_), .A2(new_n1969_), .ZN(new_n1973_));
  NAND2_X1   g00971(.A1(new_n1964_), .A2(new_n1959_), .ZN(new_n1974_));
  NAND2_X1   g00972(.A1(new_n1974_), .A2(new_n1973_), .ZN(new_n1975_));
  INV_X1     g00973(.I(new_n1961_), .ZN(new_n1976_));
  INV_X1     g00974(.I(new_n1963_), .ZN(new_n1977_));
  NOR2_X1    g00975(.A1(new_n1609_), .A2(new_n1633_), .ZN(new_n1978_));
  NOR3_X1    g00976(.A1(new_n1978_), .A2(new_n1976_), .A3(new_n1977_), .ZN(new_n1979_));
  NOR4_X1    g00977(.A1(new_n1975_), .A2(new_n1681_), .A3(new_n1684_), .A4(new_n1979_), .ZN(new_n1980_));
  NOR2_X1    g00978(.A1(new_n1971_), .A2(new_n1671_), .ZN(new_n1981_));
  NOR4_X1    g00979(.A1(new_n1681_), .A2(new_n1684_), .A3(new_n1965_), .A4(new_n1970_), .ZN(new_n1982_));
  NOR2_X1    g00980(.A1(new_n1981_), .A2(new_n1982_), .ZN(new_n1983_));
  OAI22_X1   g00981(.A1(new_n1983_), .A2(new_n1958_), .B1(new_n1972_), .B2(new_n1980_), .ZN(new_n1984_));
  NAND4_X1   g00982(.A1(new_n1581_), .A2(new_n1571_), .A3(new_n1576_), .A4(new_n1583_), .ZN(new_n1985_));
  AOI21_X1   g00983(.A1(\A[263] ), .A2(\A[264] ), .B(\A[262] ), .ZN(new_n1986_));
  NOR2_X1    g00984(.A1(new_n1986_), .A2(new_n1575_), .ZN(new_n1987_));
  AOI21_X1   g00985(.A1(\A[260] ), .A2(\A[261] ), .B(\A[259] ), .ZN(new_n1988_));
  NOR2_X1    g00986(.A1(new_n1988_), .A2(new_n1563_), .ZN(new_n1989_));
  NOR2_X1    g00987(.A1(new_n1987_), .A2(new_n1989_), .ZN(new_n1990_));
  NOR4_X1    g00988(.A1(new_n1986_), .A2(new_n1988_), .A3(new_n1563_), .A4(new_n1575_), .ZN(new_n1991_));
  NOR2_X1    g00989(.A1(new_n1990_), .A2(new_n1991_), .ZN(new_n1992_));
  XOR2_X1    g00990(.A1(new_n1985_), .A2(new_n1992_), .Z(new_n1993_));
  NOR4_X1    g00991(.A1(new_n1524_), .A2(new_n1528_), .A3(new_n1552_), .A4(new_n1549_), .ZN(new_n1994_));
  AOI21_X1   g00992(.A1(\A[269] ), .A2(\A[270] ), .B(\A[268] ), .ZN(new_n1995_));
  NOR2_X1    g00993(.A1(new_n1995_), .A2(new_n1537_), .ZN(new_n1996_));
  AOI21_X1   g00994(.A1(\A[266] ), .A2(\A[267] ), .B(\A[265] ), .ZN(new_n1997_));
  NOR2_X1    g00995(.A1(new_n1997_), .A2(new_n1526_), .ZN(new_n1998_));
  XOR2_X1    g00996(.A1(new_n1996_), .A2(new_n1998_), .Z(new_n1999_));
  NOR2_X1    g00997(.A1(new_n1999_), .A2(new_n1994_), .ZN(new_n2000_));
  NAND4_X1   g00998(.A1(new_n1543_), .A2(new_n1534_), .A3(new_n1545_), .A4(new_n1538_), .ZN(new_n2001_));
  NOR3_X1    g00999(.A1(new_n1998_), .A2(new_n1537_), .A3(new_n1995_), .ZN(new_n2002_));
  NOR3_X1    g01000(.A1(new_n1996_), .A2(new_n1526_), .A3(new_n1997_), .ZN(new_n2003_));
  NOR2_X1    g01001(.A1(new_n2002_), .A2(new_n2003_), .ZN(new_n2004_));
  NOR2_X1    g01002(.A1(new_n2004_), .A2(new_n2001_), .ZN(new_n2005_));
  OAI22_X1   g01003(.A1(new_n1594_), .A2(new_n1597_), .B1(new_n2000_), .B2(new_n2005_), .ZN(new_n2006_));
  NOR2_X1    g01004(.A1(new_n2000_), .A2(new_n2005_), .ZN(new_n2007_));
  NAND2_X1   g01005(.A1(new_n1546_), .A2(new_n1539_), .ZN(new_n2008_));
  NAND3_X1   g01006(.A1(new_n2008_), .A2(new_n1996_), .A3(new_n1998_), .ZN(new_n2009_));
  NAND4_X1   g01007(.A1(new_n2007_), .A2(new_n1555_), .A3(new_n1592_), .A4(new_n2009_), .ZN(new_n2010_));
  AOI21_X1   g01008(.A1(new_n2010_), .A2(new_n2006_), .B(new_n1993_), .ZN(new_n2011_));
  NOR4_X1    g01009(.A1(new_n1561_), .A2(new_n1565_), .A3(new_n1589_), .A4(new_n1587_), .ZN(new_n2012_));
  XOR2_X1    g01010(.A1(new_n2012_), .A2(new_n1992_), .Z(new_n2013_));
  NAND2_X1   g01011(.A1(new_n2004_), .A2(new_n2001_), .ZN(new_n2014_));
  NAND2_X1   g01012(.A1(new_n1999_), .A2(new_n1994_), .ZN(new_n2015_));
  AOI22_X1   g01013(.A1(new_n1555_), .A2(new_n1592_), .B1(new_n2014_), .B2(new_n2015_), .ZN(new_n2016_));
  NAND2_X1   g01014(.A1(new_n2015_), .A2(new_n2014_), .ZN(new_n2017_));
  NOR3_X1    g01015(.A1(new_n2017_), .A2(new_n1594_), .A3(new_n1597_), .ZN(new_n2018_));
  NOR3_X1    g01016(.A1(new_n2018_), .A2(new_n2016_), .A3(new_n2013_), .ZN(new_n2019_));
  OAI21_X1   g01017(.A1(new_n2011_), .A2(new_n2019_), .B(new_n1675_), .ZN(new_n2020_));
  NAND4_X1   g01018(.A1(new_n1676_), .A2(new_n1677_), .A3(new_n1685_), .A4(new_n1678_), .ZN(new_n2021_));
  INV_X1     g01019(.I(new_n1996_), .ZN(new_n2022_));
  INV_X1     g01020(.I(new_n1998_), .ZN(new_n2023_));
  NOR2_X1    g01021(.A1(new_n1529_), .A2(new_n1553_), .ZN(new_n2024_));
  NOR3_X1    g01022(.A1(new_n2024_), .A2(new_n2022_), .A3(new_n2023_), .ZN(new_n2025_));
  NOR4_X1    g01023(.A1(new_n2017_), .A2(new_n1594_), .A3(new_n1597_), .A4(new_n2025_), .ZN(new_n2026_));
  OAI21_X1   g01024(.A1(new_n2026_), .A2(new_n2016_), .B(new_n2013_), .ZN(new_n2027_));
  NAND4_X1   g01025(.A1(new_n1555_), .A2(new_n1592_), .A3(new_n2014_), .A4(new_n2015_), .ZN(new_n2028_));
  NAND3_X1   g01026(.A1(new_n2006_), .A2(new_n2028_), .A3(new_n1993_), .ZN(new_n2029_));
  NAND3_X1   g01027(.A1(new_n2027_), .A2(new_n2021_), .A3(new_n2029_), .ZN(new_n2030_));
  AOI21_X1   g01028(.A1(new_n2020_), .A2(new_n2030_), .B(new_n1984_), .ZN(new_n2031_));
  NOR4_X1    g01029(.A1(new_n1640_), .A2(new_n1644_), .A3(new_n1668_), .A4(new_n1666_), .ZN(new_n2032_));
  XOR2_X1    g01030(.A1(new_n2032_), .A2(new_n1957_), .Z(new_n2033_));
  AOI21_X1   g01031(.A1(new_n1678_), .A2(new_n1975_), .B(new_n2033_), .ZN(new_n2034_));
  NAND2_X1   g01032(.A1(new_n1627_), .A2(new_n1620_), .ZN(new_n2035_));
  NAND3_X1   g01033(.A1(new_n2035_), .A2(new_n1961_), .A3(new_n1963_), .ZN(new_n2036_));
  NAND4_X1   g01034(.A1(new_n1971_), .A2(new_n1672_), .A3(new_n1673_), .A4(new_n2036_), .ZN(new_n2037_));
  OAI22_X1   g01035(.A1(new_n1681_), .A2(new_n1684_), .B1(new_n1965_), .B2(new_n1970_), .ZN(new_n2038_));
  NAND2_X1   g01036(.A1(new_n1971_), .A2(new_n1671_), .ZN(new_n2039_));
  NAND2_X1   g01037(.A1(new_n2039_), .A2(new_n2038_), .ZN(new_n2040_));
  AOI22_X1   g01038(.A1(new_n2040_), .A2(new_n2033_), .B1(new_n2034_), .B2(new_n2037_), .ZN(new_n2041_));
  AOI21_X1   g01039(.A1(new_n2027_), .A2(new_n2029_), .B(new_n2021_), .ZN(new_n2042_));
  NOR3_X1    g01040(.A1(new_n2011_), .A2(new_n2019_), .A3(new_n1675_), .ZN(new_n2043_));
  NOR3_X1    g01041(.A1(new_n2042_), .A2(new_n2043_), .A3(new_n2041_), .ZN(new_n2044_));
  OAI21_X1   g01042(.A1(new_n2031_), .A2(new_n2044_), .B(new_n1950_), .ZN(new_n2045_));
  OAI21_X1   g01043(.A1(new_n2042_), .A2(new_n2043_), .B(new_n2041_), .ZN(new_n2046_));
  NAND3_X1   g01044(.A1(new_n2020_), .A2(new_n2030_), .A3(new_n1984_), .ZN(new_n2047_));
  NAND3_X1   g01045(.A1(new_n2046_), .A2(new_n2047_), .A3(new_n1838_), .ZN(new_n2048_));
  AOI21_X1   g01046(.A1(new_n2045_), .A2(new_n2048_), .B(new_n1949_), .ZN(new_n2049_));
  AND2_X2    g01047(.A1(new_n1939_), .A2(new_n1948_), .Z(new_n2050_));
  AOI21_X1   g01048(.A1(new_n2046_), .A2(new_n2047_), .B(new_n1838_), .ZN(new_n2051_));
  NOR3_X1    g01049(.A1(new_n1950_), .A2(new_n2044_), .A3(new_n2031_), .ZN(new_n2052_));
  NOR3_X1    g01050(.A1(new_n2050_), .A2(new_n2052_), .A3(new_n2051_), .ZN(new_n2053_));
  OAI21_X1   g01051(.A1(new_n2053_), .A2(new_n2049_), .B(new_n1842_), .ZN(new_n2054_));
  NOR2_X1    g01052(.A1(new_n1950_), .A2(new_n1839_), .ZN(new_n2055_));
  NAND2_X1   g01053(.A1(new_n2055_), .A2(new_n1517_), .ZN(new_n2056_));
  OAI21_X1   g01054(.A1(new_n2052_), .A2(new_n2051_), .B(new_n2050_), .ZN(new_n2057_));
  NAND3_X1   g01055(.A1(new_n2045_), .A2(new_n2048_), .A3(new_n1949_), .ZN(new_n2058_));
  NAND3_X1   g01056(.A1(new_n2057_), .A2(new_n2058_), .A3(new_n2056_), .ZN(new_n2059_));
  AOI21_X1   g01057(.A1(new_n2054_), .A2(new_n2059_), .B(new_n1515_), .ZN(new_n2060_));
  INV_X1     g01058(.I(new_n1515_), .ZN(new_n2061_));
  AOI21_X1   g01059(.A1(new_n2057_), .A2(new_n2058_), .B(new_n2056_), .ZN(new_n2062_));
  NOR3_X1    g01060(.A1(new_n2053_), .A2(new_n2049_), .A3(new_n1842_), .ZN(new_n2063_));
  NOR3_X1    g01061(.A1(new_n2061_), .A2(new_n2062_), .A3(new_n2063_), .ZN(new_n2064_));
  NOR2_X1    g01062(.A1(new_n2064_), .A2(new_n2060_), .ZN(new_n2065_));
  NOR2_X1    g01063(.A1(new_n2055_), .A2(new_n1517_), .ZN(new_n2066_));
  NOR2_X1    g01064(.A1(new_n1842_), .A2(new_n2066_), .ZN(new_n2067_));
  INV_X1     g01065(.I(new_n2067_), .ZN(new_n2068_));
  INV_X1     g01066(.I(\A[169] ), .ZN(new_n2069_));
  INV_X1     g01067(.I(\A[170] ), .ZN(new_n2070_));
  NAND2_X1   g01068(.A1(new_n2070_), .A2(\A[171] ), .ZN(new_n2071_));
  INV_X1     g01069(.I(\A[171] ), .ZN(new_n2072_));
  NAND2_X1   g01070(.A1(new_n2072_), .A2(\A[170] ), .ZN(new_n2073_));
  AOI21_X1   g01071(.A1(new_n2071_), .A2(new_n2073_), .B(new_n2069_), .ZN(new_n2074_));
  NOR2_X1    g01072(.A1(\A[170] ), .A2(\A[171] ), .ZN(new_n2075_));
  INV_X1     g01073(.I(new_n2075_), .ZN(new_n2076_));
  NAND2_X1   g01074(.A1(\A[170] ), .A2(\A[171] ), .ZN(new_n2077_));
  AOI21_X1   g01075(.A1(new_n2076_), .A2(new_n2077_), .B(\A[169] ), .ZN(new_n2078_));
  INV_X1     g01076(.I(\A[172] ), .ZN(new_n2079_));
  INV_X1     g01077(.I(\A[173] ), .ZN(new_n2080_));
  NAND2_X1   g01078(.A1(new_n2080_), .A2(\A[174] ), .ZN(new_n2081_));
  INV_X1     g01079(.I(\A[174] ), .ZN(new_n2082_));
  NAND2_X1   g01080(.A1(new_n2082_), .A2(\A[173] ), .ZN(new_n2083_));
  AOI21_X1   g01081(.A1(new_n2081_), .A2(new_n2083_), .B(new_n2079_), .ZN(new_n2084_));
  NOR2_X1    g01082(.A1(\A[173] ), .A2(\A[174] ), .ZN(new_n2085_));
  INV_X1     g01083(.I(new_n2085_), .ZN(new_n2086_));
  NAND2_X1   g01084(.A1(\A[173] ), .A2(\A[174] ), .ZN(new_n2087_));
  AOI21_X1   g01085(.A1(new_n2086_), .A2(new_n2087_), .B(\A[172] ), .ZN(new_n2088_));
  NOR4_X1    g01086(.A1(new_n2074_), .A2(new_n2078_), .A3(new_n2088_), .A4(new_n2084_), .ZN(new_n2089_));
  OAI22_X1   g01087(.A1(new_n2074_), .A2(new_n2078_), .B1(new_n2088_), .B2(new_n2084_), .ZN(new_n2090_));
  INV_X1     g01088(.I(new_n2090_), .ZN(new_n2091_));
  NOR2_X1    g01089(.A1(new_n2091_), .A2(new_n2089_), .ZN(new_n2092_));
  INV_X1     g01090(.I(\A[165] ), .ZN(new_n2093_));
  NOR2_X1    g01091(.A1(new_n2093_), .A2(\A[164] ), .ZN(new_n2094_));
  INV_X1     g01092(.I(\A[164] ), .ZN(new_n2095_));
  NOR2_X1    g01093(.A1(new_n2095_), .A2(\A[165] ), .ZN(new_n2096_));
  OAI21_X1   g01094(.A1(new_n2094_), .A2(new_n2096_), .B(\A[163] ), .ZN(new_n2097_));
  INV_X1     g01095(.I(\A[163] ), .ZN(new_n2098_));
  NAND2_X1   g01096(.A1(\A[164] ), .A2(\A[165] ), .ZN(new_n2099_));
  INV_X1     g01097(.I(new_n2099_), .ZN(new_n2100_));
  NOR2_X1    g01098(.A1(\A[164] ), .A2(\A[165] ), .ZN(new_n2101_));
  OAI21_X1   g01099(.A1(new_n2100_), .A2(new_n2101_), .B(new_n2098_), .ZN(new_n2102_));
  INV_X1     g01100(.I(\A[168] ), .ZN(new_n2103_));
  NOR2_X1    g01101(.A1(new_n2103_), .A2(\A[167] ), .ZN(new_n2104_));
  INV_X1     g01102(.I(\A[167] ), .ZN(new_n2105_));
  NOR2_X1    g01103(.A1(new_n2105_), .A2(\A[168] ), .ZN(new_n2106_));
  OAI21_X1   g01104(.A1(new_n2104_), .A2(new_n2106_), .B(\A[166] ), .ZN(new_n2107_));
  INV_X1     g01105(.I(\A[166] ), .ZN(new_n2108_));
  AND2_X2    g01106(.A1(\A[167] ), .A2(\A[168] ), .Z(new_n2109_));
  NOR2_X1    g01107(.A1(\A[167] ), .A2(\A[168] ), .ZN(new_n2110_));
  OAI21_X1   g01108(.A1(new_n2109_), .A2(new_n2110_), .B(new_n2108_), .ZN(new_n2111_));
  NAND4_X1   g01109(.A1(new_n2097_), .A2(new_n2107_), .A3(new_n2102_), .A4(new_n2111_), .ZN(new_n2112_));
  NAND2_X1   g01110(.A1(new_n2095_), .A2(\A[165] ), .ZN(new_n2113_));
  NAND2_X1   g01111(.A1(new_n2093_), .A2(\A[164] ), .ZN(new_n2114_));
  AOI21_X1   g01112(.A1(new_n2113_), .A2(new_n2114_), .B(new_n2098_), .ZN(new_n2115_));
  INV_X1     g01113(.I(new_n2101_), .ZN(new_n2116_));
  AOI21_X1   g01114(.A1(new_n2116_), .A2(new_n2099_), .B(\A[163] ), .ZN(new_n2117_));
  NAND2_X1   g01115(.A1(new_n2105_), .A2(\A[168] ), .ZN(new_n2118_));
  NAND2_X1   g01116(.A1(new_n2103_), .A2(\A[167] ), .ZN(new_n2119_));
  AOI21_X1   g01117(.A1(new_n2118_), .A2(new_n2119_), .B(new_n2108_), .ZN(new_n2120_));
  NAND2_X1   g01118(.A1(\A[167] ), .A2(\A[168] ), .ZN(new_n2121_));
  OR2_X2     g01119(.A1(\A[167] ), .A2(\A[168] ), .Z(new_n2122_));
  AOI21_X1   g01120(.A1(new_n2122_), .A2(new_n2121_), .B(\A[166] ), .ZN(new_n2123_));
  OAI22_X1   g01121(.A1(new_n2115_), .A2(new_n2117_), .B1(new_n2120_), .B2(new_n2123_), .ZN(new_n2124_));
  NAND2_X1   g01122(.A1(new_n2124_), .A2(new_n2112_), .ZN(new_n2125_));
  NAND2_X1   g01123(.A1(new_n2092_), .A2(new_n2125_), .ZN(new_n2126_));
  NOR2_X1    g01124(.A1(new_n2072_), .A2(\A[170] ), .ZN(new_n2127_));
  NOR2_X1    g01125(.A1(new_n2070_), .A2(\A[171] ), .ZN(new_n2128_));
  OAI21_X1   g01126(.A1(new_n2127_), .A2(new_n2128_), .B(\A[169] ), .ZN(new_n2129_));
  INV_X1     g01127(.I(new_n2077_), .ZN(new_n2130_));
  OAI21_X1   g01128(.A1(new_n2130_), .A2(new_n2075_), .B(new_n2069_), .ZN(new_n2131_));
  NOR2_X1    g01129(.A1(new_n2082_), .A2(\A[173] ), .ZN(new_n2132_));
  NOR2_X1    g01130(.A1(new_n2080_), .A2(\A[174] ), .ZN(new_n2133_));
  OAI21_X1   g01131(.A1(new_n2132_), .A2(new_n2133_), .B(\A[172] ), .ZN(new_n2134_));
  INV_X1     g01132(.I(new_n2087_), .ZN(new_n2135_));
  OAI21_X1   g01133(.A1(new_n2135_), .A2(new_n2085_), .B(new_n2079_), .ZN(new_n2136_));
  NAND4_X1   g01134(.A1(new_n2129_), .A2(new_n2131_), .A3(new_n2134_), .A4(new_n2136_), .ZN(new_n2137_));
  NAND2_X1   g01135(.A1(new_n2090_), .A2(new_n2137_), .ZN(new_n2138_));
  NOR4_X1    g01136(.A1(new_n2115_), .A2(new_n2117_), .A3(new_n2120_), .A4(new_n2123_), .ZN(new_n2139_));
  AOI22_X1   g01137(.A1(new_n2097_), .A2(new_n2102_), .B1(new_n2107_), .B2(new_n2111_), .ZN(new_n2140_));
  NOR2_X1    g01138(.A1(new_n2140_), .A2(new_n2139_), .ZN(new_n2141_));
  NAND2_X1   g01139(.A1(new_n2138_), .A2(new_n2141_), .ZN(new_n2142_));
  INV_X1     g01140(.I(\A[157] ), .ZN(new_n2143_));
  INV_X1     g01141(.I(\A[158] ), .ZN(new_n2144_));
  NAND2_X1   g01142(.A1(new_n2144_), .A2(\A[159] ), .ZN(new_n2145_));
  INV_X1     g01143(.I(\A[159] ), .ZN(new_n2146_));
  NAND2_X1   g01144(.A1(new_n2146_), .A2(\A[158] ), .ZN(new_n2147_));
  AOI21_X1   g01145(.A1(new_n2145_), .A2(new_n2147_), .B(new_n2143_), .ZN(new_n2148_));
  NOR2_X1    g01146(.A1(\A[158] ), .A2(\A[159] ), .ZN(new_n2149_));
  INV_X1     g01147(.I(new_n2149_), .ZN(new_n2150_));
  NAND2_X1   g01148(.A1(\A[158] ), .A2(\A[159] ), .ZN(new_n2151_));
  AOI21_X1   g01149(.A1(new_n2150_), .A2(new_n2151_), .B(\A[157] ), .ZN(new_n2152_));
  INV_X1     g01150(.I(\A[160] ), .ZN(new_n2153_));
  INV_X1     g01151(.I(\A[161] ), .ZN(new_n2154_));
  NAND2_X1   g01152(.A1(new_n2154_), .A2(\A[162] ), .ZN(new_n2155_));
  INV_X1     g01153(.I(\A[162] ), .ZN(new_n2156_));
  NAND2_X1   g01154(.A1(new_n2156_), .A2(\A[161] ), .ZN(new_n2157_));
  AOI21_X1   g01155(.A1(new_n2155_), .A2(new_n2157_), .B(new_n2153_), .ZN(new_n2158_));
  NOR2_X1    g01156(.A1(\A[161] ), .A2(\A[162] ), .ZN(new_n2159_));
  INV_X1     g01157(.I(new_n2159_), .ZN(new_n2160_));
  NAND2_X1   g01158(.A1(\A[161] ), .A2(\A[162] ), .ZN(new_n2161_));
  AOI21_X1   g01159(.A1(new_n2160_), .A2(new_n2161_), .B(\A[160] ), .ZN(new_n2162_));
  NOR4_X1    g01160(.A1(new_n2148_), .A2(new_n2152_), .A3(new_n2162_), .A4(new_n2158_), .ZN(new_n2163_));
  NOR2_X1    g01161(.A1(new_n2146_), .A2(\A[158] ), .ZN(new_n2164_));
  NOR2_X1    g01162(.A1(new_n2144_), .A2(\A[159] ), .ZN(new_n2165_));
  OAI21_X1   g01163(.A1(new_n2164_), .A2(new_n2165_), .B(\A[157] ), .ZN(new_n2166_));
  INV_X1     g01164(.I(new_n2151_), .ZN(new_n2167_));
  OAI21_X1   g01165(.A1(new_n2167_), .A2(new_n2149_), .B(new_n2143_), .ZN(new_n2168_));
  NOR2_X1    g01166(.A1(new_n2156_), .A2(\A[161] ), .ZN(new_n2169_));
  NOR2_X1    g01167(.A1(new_n2154_), .A2(\A[162] ), .ZN(new_n2170_));
  OAI21_X1   g01168(.A1(new_n2169_), .A2(new_n2170_), .B(\A[160] ), .ZN(new_n2171_));
  AND2_X2    g01169(.A1(\A[161] ), .A2(\A[162] ), .Z(new_n2172_));
  OAI21_X1   g01170(.A1(new_n2172_), .A2(new_n2159_), .B(new_n2153_), .ZN(new_n2173_));
  AOI22_X1   g01171(.A1(new_n2166_), .A2(new_n2168_), .B1(new_n2171_), .B2(new_n2173_), .ZN(new_n2174_));
  NOR2_X1    g01172(.A1(new_n2163_), .A2(new_n2174_), .ZN(new_n2175_));
  INV_X1     g01173(.I(\A[153] ), .ZN(new_n2176_));
  NOR2_X1    g01174(.A1(new_n2176_), .A2(\A[152] ), .ZN(new_n2177_));
  INV_X1     g01175(.I(\A[152] ), .ZN(new_n2178_));
  NOR2_X1    g01176(.A1(new_n2178_), .A2(\A[153] ), .ZN(new_n2179_));
  OAI21_X1   g01177(.A1(new_n2177_), .A2(new_n2179_), .B(\A[151] ), .ZN(new_n2180_));
  INV_X1     g01178(.I(\A[151] ), .ZN(new_n2181_));
  NAND2_X1   g01179(.A1(\A[152] ), .A2(\A[153] ), .ZN(new_n2182_));
  INV_X1     g01180(.I(new_n2182_), .ZN(new_n2183_));
  NOR2_X1    g01181(.A1(\A[152] ), .A2(\A[153] ), .ZN(new_n2184_));
  OAI21_X1   g01182(.A1(new_n2183_), .A2(new_n2184_), .B(new_n2181_), .ZN(new_n2185_));
  INV_X1     g01183(.I(\A[156] ), .ZN(new_n2186_));
  NOR2_X1    g01184(.A1(new_n2186_), .A2(\A[155] ), .ZN(new_n2187_));
  INV_X1     g01185(.I(\A[155] ), .ZN(new_n2188_));
  NOR2_X1    g01186(.A1(new_n2188_), .A2(\A[156] ), .ZN(new_n2189_));
  OAI21_X1   g01187(.A1(new_n2187_), .A2(new_n2189_), .B(\A[154] ), .ZN(new_n2190_));
  INV_X1     g01188(.I(\A[154] ), .ZN(new_n2191_));
  NAND2_X1   g01189(.A1(\A[155] ), .A2(\A[156] ), .ZN(new_n2192_));
  INV_X1     g01190(.I(new_n2192_), .ZN(new_n2193_));
  NOR2_X1    g01191(.A1(\A[155] ), .A2(\A[156] ), .ZN(new_n2194_));
  OAI21_X1   g01192(.A1(new_n2193_), .A2(new_n2194_), .B(new_n2191_), .ZN(new_n2195_));
  NAND4_X1   g01193(.A1(new_n2180_), .A2(new_n2185_), .A3(new_n2190_), .A4(new_n2195_), .ZN(new_n2196_));
  NAND2_X1   g01194(.A1(new_n2178_), .A2(\A[153] ), .ZN(new_n2197_));
  NAND2_X1   g01195(.A1(new_n2176_), .A2(\A[152] ), .ZN(new_n2198_));
  AOI21_X1   g01196(.A1(new_n2197_), .A2(new_n2198_), .B(new_n2181_), .ZN(new_n2199_));
  INV_X1     g01197(.I(new_n2184_), .ZN(new_n2200_));
  AOI21_X1   g01198(.A1(new_n2200_), .A2(new_n2182_), .B(\A[151] ), .ZN(new_n2201_));
  NAND2_X1   g01199(.A1(new_n2188_), .A2(\A[156] ), .ZN(new_n2202_));
  NAND2_X1   g01200(.A1(new_n2186_), .A2(\A[155] ), .ZN(new_n2203_));
  AOI21_X1   g01201(.A1(new_n2202_), .A2(new_n2203_), .B(new_n2191_), .ZN(new_n2204_));
  OR2_X2     g01202(.A1(\A[155] ), .A2(\A[156] ), .Z(new_n2205_));
  AOI21_X1   g01203(.A1(new_n2205_), .A2(new_n2192_), .B(\A[154] ), .ZN(new_n2206_));
  OAI22_X1   g01204(.A1(new_n2199_), .A2(new_n2201_), .B1(new_n2204_), .B2(new_n2206_), .ZN(new_n2207_));
  NAND2_X1   g01205(.A1(new_n2196_), .A2(new_n2207_), .ZN(new_n2208_));
  NAND2_X1   g01206(.A1(new_n2175_), .A2(new_n2208_), .ZN(new_n2209_));
  NAND4_X1   g01207(.A1(new_n2166_), .A2(new_n2171_), .A3(new_n2168_), .A4(new_n2173_), .ZN(new_n2210_));
  OAI22_X1   g01208(.A1(new_n2148_), .A2(new_n2152_), .B1(new_n2162_), .B2(new_n2158_), .ZN(new_n2211_));
  NAND2_X1   g01209(.A1(new_n2211_), .A2(new_n2210_), .ZN(new_n2212_));
  NOR4_X1    g01210(.A1(new_n2199_), .A2(new_n2201_), .A3(new_n2204_), .A4(new_n2206_), .ZN(new_n2213_));
  AOI22_X1   g01211(.A1(new_n2180_), .A2(new_n2185_), .B1(new_n2190_), .B2(new_n2195_), .ZN(new_n2214_));
  NOR2_X1    g01212(.A1(new_n2214_), .A2(new_n2213_), .ZN(new_n2215_));
  NAND2_X1   g01213(.A1(new_n2215_), .A2(new_n2212_), .ZN(new_n2216_));
  AOI22_X1   g01214(.A1(new_n2126_), .A2(new_n2142_), .B1(new_n2209_), .B2(new_n2216_), .ZN(new_n2217_));
  NOR2_X1    g01215(.A1(new_n2138_), .A2(new_n2141_), .ZN(new_n2218_));
  NOR2_X1    g01216(.A1(new_n2092_), .A2(new_n2125_), .ZN(new_n2219_));
  NOR2_X1    g01217(.A1(new_n2215_), .A2(new_n2212_), .ZN(new_n2220_));
  NOR2_X1    g01218(.A1(new_n2175_), .A2(new_n2208_), .ZN(new_n2221_));
  NOR4_X1    g01219(.A1(new_n2219_), .A2(new_n2218_), .A3(new_n2221_), .A4(new_n2220_), .ZN(new_n2222_));
  NOR2_X1    g01220(.A1(new_n2222_), .A2(new_n2217_), .ZN(new_n2223_));
  INV_X1     g01221(.I(\A[145] ), .ZN(new_n2224_));
  INV_X1     g01222(.I(\A[146] ), .ZN(new_n2225_));
  NAND2_X1   g01223(.A1(new_n2225_), .A2(\A[147] ), .ZN(new_n2226_));
  INV_X1     g01224(.I(\A[147] ), .ZN(new_n2227_));
  NAND2_X1   g01225(.A1(new_n2227_), .A2(\A[146] ), .ZN(new_n2228_));
  AOI21_X1   g01226(.A1(new_n2226_), .A2(new_n2228_), .B(new_n2224_), .ZN(new_n2229_));
  NOR2_X1    g01227(.A1(\A[146] ), .A2(\A[147] ), .ZN(new_n2230_));
  INV_X1     g01228(.I(new_n2230_), .ZN(new_n2231_));
  NAND2_X1   g01229(.A1(\A[146] ), .A2(\A[147] ), .ZN(new_n2232_));
  AOI21_X1   g01230(.A1(new_n2231_), .A2(new_n2232_), .B(\A[145] ), .ZN(new_n2233_));
  INV_X1     g01231(.I(\A[148] ), .ZN(new_n2234_));
  INV_X1     g01232(.I(\A[149] ), .ZN(new_n2235_));
  NAND2_X1   g01233(.A1(new_n2235_), .A2(\A[150] ), .ZN(new_n2236_));
  INV_X1     g01234(.I(\A[150] ), .ZN(new_n2237_));
  NAND2_X1   g01235(.A1(new_n2237_), .A2(\A[149] ), .ZN(new_n2238_));
  AOI21_X1   g01236(.A1(new_n2236_), .A2(new_n2238_), .B(new_n2234_), .ZN(new_n2239_));
  NOR2_X1    g01237(.A1(\A[149] ), .A2(\A[150] ), .ZN(new_n2240_));
  INV_X1     g01238(.I(new_n2240_), .ZN(new_n2241_));
  NAND2_X1   g01239(.A1(\A[149] ), .A2(\A[150] ), .ZN(new_n2242_));
  AOI21_X1   g01240(.A1(new_n2241_), .A2(new_n2242_), .B(\A[148] ), .ZN(new_n2243_));
  NOR4_X1    g01241(.A1(new_n2229_), .A2(new_n2233_), .A3(new_n2243_), .A4(new_n2239_), .ZN(new_n2244_));
  OAI22_X1   g01242(.A1(new_n2229_), .A2(new_n2233_), .B1(new_n2243_), .B2(new_n2239_), .ZN(new_n2245_));
  INV_X1     g01243(.I(new_n2245_), .ZN(new_n2246_));
  NOR2_X1    g01244(.A1(new_n2246_), .A2(new_n2244_), .ZN(new_n2247_));
  INV_X1     g01245(.I(\A[141] ), .ZN(new_n2248_));
  NOR2_X1    g01246(.A1(new_n2248_), .A2(\A[140] ), .ZN(new_n2249_));
  INV_X1     g01247(.I(\A[140] ), .ZN(new_n2250_));
  NOR2_X1    g01248(.A1(new_n2250_), .A2(\A[141] ), .ZN(new_n2251_));
  OAI21_X1   g01249(.A1(new_n2249_), .A2(new_n2251_), .B(\A[139] ), .ZN(new_n2252_));
  INV_X1     g01250(.I(\A[139] ), .ZN(new_n2253_));
  NAND2_X1   g01251(.A1(\A[140] ), .A2(\A[141] ), .ZN(new_n2254_));
  INV_X1     g01252(.I(new_n2254_), .ZN(new_n2255_));
  NOR2_X1    g01253(.A1(\A[140] ), .A2(\A[141] ), .ZN(new_n2256_));
  OAI21_X1   g01254(.A1(new_n2255_), .A2(new_n2256_), .B(new_n2253_), .ZN(new_n2257_));
  INV_X1     g01255(.I(\A[144] ), .ZN(new_n2258_));
  NOR2_X1    g01256(.A1(new_n2258_), .A2(\A[143] ), .ZN(new_n2259_));
  INV_X1     g01257(.I(\A[143] ), .ZN(new_n2260_));
  NOR2_X1    g01258(.A1(new_n2260_), .A2(\A[144] ), .ZN(new_n2261_));
  OAI21_X1   g01259(.A1(new_n2259_), .A2(new_n2261_), .B(\A[142] ), .ZN(new_n2262_));
  INV_X1     g01260(.I(\A[142] ), .ZN(new_n2263_));
  NAND2_X1   g01261(.A1(\A[143] ), .A2(\A[144] ), .ZN(new_n2264_));
  INV_X1     g01262(.I(new_n2264_), .ZN(new_n2265_));
  NOR2_X1    g01263(.A1(\A[143] ), .A2(\A[144] ), .ZN(new_n2266_));
  OAI21_X1   g01264(.A1(new_n2265_), .A2(new_n2266_), .B(new_n2263_), .ZN(new_n2267_));
  NAND4_X1   g01265(.A1(new_n2252_), .A2(new_n2257_), .A3(new_n2262_), .A4(new_n2267_), .ZN(new_n2268_));
  NAND2_X1   g01266(.A1(new_n2250_), .A2(\A[141] ), .ZN(new_n2269_));
  NAND2_X1   g01267(.A1(new_n2248_), .A2(\A[140] ), .ZN(new_n2270_));
  AOI21_X1   g01268(.A1(new_n2269_), .A2(new_n2270_), .B(new_n2253_), .ZN(new_n2271_));
  INV_X1     g01269(.I(new_n2256_), .ZN(new_n2272_));
  AOI21_X1   g01270(.A1(new_n2272_), .A2(new_n2254_), .B(\A[139] ), .ZN(new_n2273_));
  NAND2_X1   g01271(.A1(new_n2260_), .A2(\A[144] ), .ZN(new_n2274_));
  NAND2_X1   g01272(.A1(new_n2258_), .A2(\A[143] ), .ZN(new_n2275_));
  AOI21_X1   g01273(.A1(new_n2274_), .A2(new_n2275_), .B(new_n2263_), .ZN(new_n2276_));
  INV_X1     g01274(.I(new_n2266_), .ZN(new_n2277_));
  AOI21_X1   g01275(.A1(new_n2277_), .A2(new_n2264_), .B(\A[142] ), .ZN(new_n2278_));
  OAI22_X1   g01276(.A1(new_n2271_), .A2(new_n2273_), .B1(new_n2278_), .B2(new_n2276_), .ZN(new_n2279_));
  NAND2_X1   g01277(.A1(new_n2279_), .A2(new_n2268_), .ZN(new_n2280_));
  NAND2_X1   g01278(.A1(new_n2247_), .A2(new_n2280_), .ZN(new_n2281_));
  INV_X1     g01279(.I(new_n2226_), .ZN(new_n2282_));
  NOR2_X1    g01280(.A1(new_n2225_), .A2(\A[147] ), .ZN(new_n2283_));
  OAI21_X1   g01281(.A1(new_n2282_), .A2(new_n2283_), .B(\A[145] ), .ZN(new_n2284_));
  INV_X1     g01282(.I(new_n2232_), .ZN(new_n2285_));
  OAI21_X1   g01283(.A1(new_n2285_), .A2(new_n2230_), .B(new_n2224_), .ZN(new_n2286_));
  NOR2_X1    g01284(.A1(new_n2237_), .A2(\A[149] ), .ZN(new_n2287_));
  NOR2_X1    g01285(.A1(new_n2235_), .A2(\A[150] ), .ZN(new_n2288_));
  OAI21_X1   g01286(.A1(new_n2287_), .A2(new_n2288_), .B(\A[148] ), .ZN(new_n2289_));
  INV_X1     g01287(.I(new_n2242_), .ZN(new_n2290_));
  OAI21_X1   g01288(.A1(new_n2290_), .A2(new_n2240_), .B(new_n2234_), .ZN(new_n2291_));
  NAND4_X1   g01289(.A1(new_n2284_), .A2(new_n2286_), .A3(new_n2291_), .A4(new_n2289_), .ZN(new_n2292_));
  NAND2_X1   g01290(.A1(new_n2292_), .A2(new_n2245_), .ZN(new_n2293_));
  NOR4_X1    g01291(.A1(new_n2271_), .A2(new_n2273_), .A3(new_n2278_), .A4(new_n2276_), .ZN(new_n2294_));
  NOR2_X1    g01292(.A1(new_n2273_), .A2(new_n2271_), .ZN(new_n2295_));
  NOR2_X1    g01293(.A1(new_n2278_), .A2(new_n2276_), .ZN(new_n2296_));
  NOR2_X1    g01294(.A1(new_n2295_), .A2(new_n2296_), .ZN(new_n2297_));
  NOR2_X1    g01295(.A1(new_n2297_), .A2(new_n2294_), .ZN(new_n2298_));
  NAND2_X1   g01296(.A1(new_n2298_), .A2(new_n2293_), .ZN(new_n2299_));
  INV_X1     g01297(.I(\A[133] ), .ZN(new_n2300_));
  INV_X1     g01298(.I(\A[134] ), .ZN(new_n2301_));
  NAND2_X1   g01299(.A1(new_n2301_), .A2(\A[135] ), .ZN(new_n2302_));
  INV_X1     g01300(.I(\A[135] ), .ZN(new_n2303_));
  NAND2_X1   g01301(.A1(new_n2303_), .A2(\A[134] ), .ZN(new_n2304_));
  AOI21_X1   g01302(.A1(new_n2302_), .A2(new_n2304_), .B(new_n2300_), .ZN(new_n2305_));
  NOR2_X1    g01303(.A1(\A[134] ), .A2(\A[135] ), .ZN(new_n2306_));
  INV_X1     g01304(.I(new_n2306_), .ZN(new_n2307_));
  NAND2_X1   g01305(.A1(\A[134] ), .A2(\A[135] ), .ZN(new_n2308_));
  AOI21_X1   g01306(.A1(new_n2307_), .A2(new_n2308_), .B(\A[133] ), .ZN(new_n2309_));
  INV_X1     g01307(.I(\A[136] ), .ZN(new_n2310_));
  INV_X1     g01308(.I(\A[137] ), .ZN(new_n2311_));
  NAND2_X1   g01309(.A1(new_n2311_), .A2(\A[138] ), .ZN(new_n2312_));
  INV_X1     g01310(.I(\A[138] ), .ZN(new_n2313_));
  NAND2_X1   g01311(.A1(new_n2313_), .A2(\A[137] ), .ZN(new_n2314_));
  AOI21_X1   g01312(.A1(new_n2312_), .A2(new_n2314_), .B(new_n2310_), .ZN(new_n2315_));
  NOR2_X1    g01313(.A1(\A[137] ), .A2(\A[138] ), .ZN(new_n2316_));
  INV_X1     g01314(.I(new_n2316_), .ZN(new_n2317_));
  NAND2_X1   g01315(.A1(\A[137] ), .A2(\A[138] ), .ZN(new_n2318_));
  AOI21_X1   g01316(.A1(new_n2317_), .A2(new_n2318_), .B(\A[136] ), .ZN(new_n2319_));
  NOR4_X1    g01317(.A1(new_n2305_), .A2(new_n2309_), .A3(new_n2319_), .A4(new_n2315_), .ZN(new_n2320_));
  INV_X1     g01318(.I(new_n2302_), .ZN(new_n2321_));
  NOR2_X1    g01319(.A1(new_n2301_), .A2(\A[135] ), .ZN(new_n2322_));
  OAI21_X1   g01320(.A1(new_n2321_), .A2(new_n2322_), .B(\A[133] ), .ZN(new_n2323_));
  INV_X1     g01321(.I(new_n2308_), .ZN(new_n2324_));
  OAI21_X1   g01322(.A1(new_n2324_), .A2(new_n2306_), .B(new_n2300_), .ZN(new_n2325_));
  NOR2_X1    g01323(.A1(new_n2313_), .A2(\A[137] ), .ZN(new_n2326_));
  NOR2_X1    g01324(.A1(new_n2311_), .A2(\A[138] ), .ZN(new_n2327_));
  OAI21_X1   g01325(.A1(new_n2326_), .A2(new_n2327_), .B(\A[136] ), .ZN(new_n2328_));
  INV_X1     g01326(.I(new_n2318_), .ZN(new_n2329_));
  OAI21_X1   g01327(.A1(new_n2329_), .A2(new_n2316_), .B(new_n2310_), .ZN(new_n2330_));
  AOI22_X1   g01328(.A1(new_n2323_), .A2(new_n2325_), .B1(new_n2330_), .B2(new_n2328_), .ZN(new_n2331_));
  NOR2_X1    g01329(.A1(new_n2331_), .A2(new_n2320_), .ZN(new_n2332_));
  INV_X1     g01330(.I(\A[129] ), .ZN(new_n2333_));
  NOR2_X1    g01331(.A1(new_n2333_), .A2(\A[128] ), .ZN(new_n2334_));
  INV_X1     g01332(.I(\A[128] ), .ZN(new_n2335_));
  NOR2_X1    g01333(.A1(new_n2335_), .A2(\A[129] ), .ZN(new_n2336_));
  OAI21_X1   g01334(.A1(new_n2334_), .A2(new_n2336_), .B(\A[127] ), .ZN(new_n2337_));
  INV_X1     g01335(.I(\A[127] ), .ZN(new_n2338_));
  NAND2_X1   g01336(.A1(\A[128] ), .A2(\A[129] ), .ZN(new_n2339_));
  INV_X1     g01337(.I(new_n2339_), .ZN(new_n2340_));
  NOR2_X1    g01338(.A1(\A[128] ), .A2(\A[129] ), .ZN(new_n2341_));
  OAI21_X1   g01339(.A1(new_n2340_), .A2(new_n2341_), .B(new_n2338_), .ZN(new_n2342_));
  INV_X1     g01340(.I(\A[132] ), .ZN(new_n2343_));
  NOR2_X1    g01341(.A1(new_n2343_), .A2(\A[131] ), .ZN(new_n2344_));
  INV_X1     g01342(.I(\A[131] ), .ZN(new_n2345_));
  NOR2_X1    g01343(.A1(new_n2345_), .A2(\A[132] ), .ZN(new_n2346_));
  OAI21_X1   g01344(.A1(new_n2344_), .A2(new_n2346_), .B(\A[130] ), .ZN(new_n2347_));
  INV_X1     g01345(.I(\A[130] ), .ZN(new_n2348_));
  NAND2_X1   g01346(.A1(\A[131] ), .A2(\A[132] ), .ZN(new_n2349_));
  INV_X1     g01347(.I(new_n2349_), .ZN(new_n2350_));
  NOR2_X1    g01348(.A1(\A[131] ), .A2(\A[132] ), .ZN(new_n2351_));
  OAI21_X1   g01349(.A1(new_n2350_), .A2(new_n2351_), .B(new_n2348_), .ZN(new_n2352_));
  NAND4_X1   g01350(.A1(new_n2337_), .A2(new_n2342_), .A3(new_n2347_), .A4(new_n2352_), .ZN(new_n2353_));
  NAND2_X1   g01351(.A1(new_n2335_), .A2(\A[129] ), .ZN(new_n2354_));
  NAND2_X1   g01352(.A1(new_n2333_), .A2(\A[128] ), .ZN(new_n2355_));
  AOI21_X1   g01353(.A1(new_n2354_), .A2(new_n2355_), .B(new_n2338_), .ZN(new_n2356_));
  INV_X1     g01354(.I(new_n2341_), .ZN(new_n2357_));
  AOI21_X1   g01355(.A1(new_n2357_), .A2(new_n2339_), .B(\A[127] ), .ZN(new_n2358_));
  NAND2_X1   g01356(.A1(new_n2345_), .A2(\A[132] ), .ZN(new_n2359_));
  NAND2_X1   g01357(.A1(new_n2343_), .A2(\A[131] ), .ZN(new_n2360_));
  AOI21_X1   g01358(.A1(new_n2359_), .A2(new_n2360_), .B(new_n2348_), .ZN(new_n2361_));
  INV_X1     g01359(.I(new_n2351_), .ZN(new_n2362_));
  AOI21_X1   g01360(.A1(new_n2362_), .A2(new_n2349_), .B(\A[130] ), .ZN(new_n2363_));
  OAI22_X1   g01361(.A1(new_n2356_), .A2(new_n2358_), .B1(new_n2363_), .B2(new_n2361_), .ZN(new_n2364_));
  NAND2_X1   g01362(.A1(new_n2364_), .A2(new_n2353_), .ZN(new_n2365_));
  NAND2_X1   g01363(.A1(new_n2332_), .A2(new_n2365_), .ZN(new_n2366_));
  NAND4_X1   g01364(.A1(new_n2323_), .A2(new_n2325_), .A3(new_n2330_), .A4(new_n2328_), .ZN(new_n2367_));
  OAI22_X1   g01365(.A1(new_n2305_), .A2(new_n2309_), .B1(new_n2319_), .B2(new_n2315_), .ZN(new_n2368_));
  NAND2_X1   g01366(.A1(new_n2367_), .A2(new_n2368_), .ZN(new_n2369_));
  NOR4_X1    g01367(.A1(new_n2356_), .A2(new_n2358_), .A3(new_n2363_), .A4(new_n2361_), .ZN(new_n2370_));
  AOI22_X1   g01368(.A1(new_n2337_), .A2(new_n2342_), .B1(new_n2347_), .B2(new_n2352_), .ZN(new_n2371_));
  NOR2_X1    g01369(.A1(new_n2371_), .A2(new_n2370_), .ZN(new_n2372_));
  NAND2_X1   g01370(.A1(new_n2372_), .A2(new_n2369_), .ZN(new_n2373_));
  AOI22_X1   g01371(.A1(new_n2281_), .A2(new_n2299_), .B1(new_n2366_), .B2(new_n2373_), .ZN(new_n2374_));
  NOR2_X1    g01372(.A1(new_n2298_), .A2(new_n2293_), .ZN(new_n2375_));
  NOR2_X1    g01373(.A1(new_n2247_), .A2(new_n2280_), .ZN(new_n2376_));
  NOR2_X1    g01374(.A1(new_n2372_), .A2(new_n2369_), .ZN(new_n2377_));
  NOR2_X1    g01375(.A1(new_n2332_), .A2(new_n2365_), .ZN(new_n2378_));
  NOR4_X1    g01376(.A1(new_n2375_), .A2(new_n2376_), .A3(new_n2377_), .A4(new_n2378_), .ZN(new_n2379_));
  NOR2_X1    g01377(.A1(new_n2379_), .A2(new_n2374_), .ZN(new_n2380_));
  NAND2_X1   g01378(.A1(new_n2380_), .A2(new_n2223_), .ZN(new_n2381_));
  INV_X1     g01379(.I(new_n2381_), .ZN(new_n2382_));
  NOR2_X1    g01380(.A1(new_n2380_), .A2(new_n2223_), .ZN(new_n2383_));
  NOR2_X1    g01381(.A1(new_n2382_), .A2(new_n2383_), .ZN(new_n2384_));
  INV_X1     g01382(.I(\A[123] ), .ZN(new_n2385_));
  NOR2_X1    g01383(.A1(new_n2385_), .A2(\A[122] ), .ZN(new_n2386_));
  INV_X1     g01384(.I(\A[122] ), .ZN(new_n2387_));
  NOR2_X1    g01385(.A1(new_n2387_), .A2(\A[123] ), .ZN(new_n2388_));
  OAI21_X1   g01386(.A1(new_n2386_), .A2(new_n2388_), .B(\A[121] ), .ZN(new_n2389_));
  INV_X1     g01387(.I(\A[121] ), .ZN(new_n2390_));
  NOR2_X1    g01388(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n2391_));
  NAND2_X1   g01389(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n2392_));
  INV_X1     g01390(.I(new_n2392_), .ZN(new_n2393_));
  OAI21_X1   g01391(.A1(new_n2393_), .A2(new_n2391_), .B(new_n2390_), .ZN(new_n2394_));
  INV_X1     g01392(.I(\A[126] ), .ZN(new_n2395_));
  NOR2_X1    g01393(.A1(new_n2395_), .A2(\A[125] ), .ZN(new_n2396_));
  INV_X1     g01394(.I(\A[125] ), .ZN(new_n2397_));
  NOR2_X1    g01395(.A1(new_n2397_), .A2(\A[126] ), .ZN(new_n2398_));
  OAI21_X1   g01396(.A1(new_n2396_), .A2(new_n2398_), .B(\A[124] ), .ZN(new_n2399_));
  INV_X1     g01397(.I(\A[124] ), .ZN(new_n2400_));
  NOR2_X1    g01398(.A1(\A[125] ), .A2(\A[126] ), .ZN(new_n2401_));
  NAND2_X1   g01399(.A1(\A[125] ), .A2(\A[126] ), .ZN(new_n2402_));
  INV_X1     g01400(.I(new_n2402_), .ZN(new_n2403_));
  OAI21_X1   g01401(.A1(new_n2403_), .A2(new_n2401_), .B(new_n2400_), .ZN(new_n2404_));
  NAND4_X1   g01402(.A1(new_n2389_), .A2(new_n2394_), .A3(new_n2399_), .A4(new_n2404_), .ZN(new_n2405_));
  NAND2_X1   g01403(.A1(new_n2387_), .A2(\A[123] ), .ZN(new_n2406_));
  NAND2_X1   g01404(.A1(new_n2385_), .A2(\A[122] ), .ZN(new_n2407_));
  AOI21_X1   g01405(.A1(new_n2406_), .A2(new_n2407_), .B(new_n2390_), .ZN(new_n2408_));
  INV_X1     g01406(.I(new_n2391_), .ZN(new_n2409_));
  AOI21_X1   g01407(.A1(new_n2409_), .A2(new_n2392_), .B(\A[121] ), .ZN(new_n2410_));
  NAND2_X1   g01408(.A1(new_n2397_), .A2(\A[126] ), .ZN(new_n2411_));
  NAND2_X1   g01409(.A1(new_n2395_), .A2(\A[125] ), .ZN(new_n2412_));
  AOI21_X1   g01410(.A1(new_n2411_), .A2(new_n2412_), .B(new_n2400_), .ZN(new_n2413_));
  INV_X1     g01411(.I(new_n2401_), .ZN(new_n2414_));
  AOI21_X1   g01412(.A1(new_n2414_), .A2(new_n2402_), .B(\A[124] ), .ZN(new_n2415_));
  OAI22_X1   g01413(.A1(new_n2408_), .A2(new_n2410_), .B1(new_n2415_), .B2(new_n2413_), .ZN(new_n2416_));
  NAND2_X1   g01414(.A1(new_n2416_), .A2(new_n2405_), .ZN(new_n2417_));
  INV_X1     g01415(.I(\A[115] ), .ZN(new_n2418_));
  INV_X1     g01416(.I(\A[116] ), .ZN(new_n2419_));
  NAND2_X1   g01417(.A1(new_n2419_), .A2(\A[117] ), .ZN(new_n2420_));
  INV_X1     g01418(.I(\A[117] ), .ZN(new_n2421_));
  NAND2_X1   g01419(.A1(new_n2421_), .A2(\A[116] ), .ZN(new_n2422_));
  AOI21_X1   g01420(.A1(new_n2420_), .A2(new_n2422_), .B(new_n2418_), .ZN(new_n2423_));
  NAND2_X1   g01421(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n2424_));
  NOR2_X1    g01422(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n2425_));
  INV_X1     g01423(.I(new_n2425_), .ZN(new_n2426_));
  AOI21_X1   g01424(.A1(new_n2426_), .A2(new_n2424_), .B(\A[115] ), .ZN(new_n2427_));
  INV_X1     g01425(.I(\A[118] ), .ZN(new_n2428_));
  INV_X1     g01426(.I(\A[119] ), .ZN(new_n2429_));
  NAND2_X1   g01427(.A1(new_n2429_), .A2(\A[120] ), .ZN(new_n2430_));
  INV_X1     g01428(.I(\A[120] ), .ZN(new_n2431_));
  NAND2_X1   g01429(.A1(new_n2431_), .A2(\A[119] ), .ZN(new_n2432_));
  AOI21_X1   g01430(.A1(new_n2430_), .A2(new_n2432_), .B(new_n2428_), .ZN(new_n2433_));
  NAND2_X1   g01431(.A1(\A[119] ), .A2(\A[120] ), .ZN(new_n2434_));
  OR2_X2     g01432(.A1(\A[119] ), .A2(\A[120] ), .Z(new_n2435_));
  AOI21_X1   g01433(.A1(new_n2435_), .A2(new_n2434_), .B(\A[118] ), .ZN(new_n2436_));
  NOR4_X1    g01434(.A1(new_n2423_), .A2(new_n2427_), .A3(new_n2433_), .A4(new_n2436_), .ZN(new_n2437_));
  NOR2_X1    g01435(.A1(new_n2421_), .A2(\A[116] ), .ZN(new_n2438_));
  NOR2_X1    g01436(.A1(new_n2419_), .A2(\A[117] ), .ZN(new_n2439_));
  OAI21_X1   g01437(.A1(new_n2438_), .A2(new_n2439_), .B(\A[115] ), .ZN(new_n2440_));
  INV_X1     g01438(.I(new_n2424_), .ZN(new_n2441_));
  OAI21_X1   g01439(.A1(new_n2441_), .A2(new_n2425_), .B(new_n2418_), .ZN(new_n2442_));
  NOR2_X1    g01440(.A1(new_n2431_), .A2(\A[119] ), .ZN(new_n2443_));
  NOR2_X1    g01441(.A1(new_n2429_), .A2(\A[120] ), .ZN(new_n2444_));
  OAI21_X1   g01442(.A1(new_n2443_), .A2(new_n2444_), .B(\A[118] ), .ZN(new_n2445_));
  AND2_X2    g01443(.A1(\A[119] ), .A2(\A[120] ), .Z(new_n2446_));
  NOR2_X1    g01444(.A1(\A[119] ), .A2(\A[120] ), .ZN(new_n2447_));
  OAI21_X1   g01445(.A1(new_n2446_), .A2(new_n2447_), .B(new_n2428_), .ZN(new_n2448_));
  AOI22_X1   g01446(.A1(new_n2440_), .A2(new_n2442_), .B1(new_n2445_), .B2(new_n2448_), .ZN(new_n2449_));
  NOR2_X1    g01447(.A1(new_n2449_), .A2(new_n2437_), .ZN(new_n2450_));
  NOR2_X1    g01448(.A1(new_n2417_), .A2(new_n2450_), .ZN(new_n2451_));
  NOR4_X1    g01449(.A1(new_n2408_), .A2(new_n2410_), .A3(new_n2415_), .A4(new_n2413_), .ZN(new_n2452_));
  AOI22_X1   g01450(.A1(new_n2389_), .A2(new_n2394_), .B1(new_n2399_), .B2(new_n2404_), .ZN(new_n2453_));
  NOR2_X1    g01451(.A1(new_n2453_), .A2(new_n2452_), .ZN(new_n2454_));
  NAND4_X1   g01452(.A1(new_n2440_), .A2(new_n2445_), .A3(new_n2442_), .A4(new_n2448_), .ZN(new_n2455_));
  OAI22_X1   g01453(.A1(new_n2423_), .A2(new_n2427_), .B1(new_n2433_), .B2(new_n2436_), .ZN(new_n2456_));
  NAND2_X1   g01454(.A1(new_n2456_), .A2(new_n2455_), .ZN(new_n2457_));
  NOR2_X1    g01455(.A1(new_n2454_), .A2(new_n2457_), .ZN(new_n2458_));
  INV_X1     g01456(.I(\A[111] ), .ZN(new_n2459_));
  NOR2_X1    g01457(.A1(new_n2459_), .A2(\A[110] ), .ZN(new_n2460_));
  INV_X1     g01458(.I(\A[110] ), .ZN(new_n2461_));
  NOR2_X1    g01459(.A1(new_n2461_), .A2(\A[111] ), .ZN(new_n2462_));
  OAI21_X1   g01460(.A1(new_n2460_), .A2(new_n2462_), .B(\A[109] ), .ZN(new_n2463_));
  INV_X1     g01461(.I(\A[109] ), .ZN(new_n2464_));
  NOR2_X1    g01462(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n2465_));
  NAND2_X1   g01463(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n2466_));
  INV_X1     g01464(.I(new_n2466_), .ZN(new_n2467_));
  OAI21_X1   g01465(.A1(new_n2467_), .A2(new_n2465_), .B(new_n2464_), .ZN(new_n2468_));
  INV_X1     g01466(.I(\A[114] ), .ZN(new_n2469_));
  NOR2_X1    g01467(.A1(new_n2469_), .A2(\A[113] ), .ZN(new_n2470_));
  INV_X1     g01468(.I(\A[113] ), .ZN(new_n2471_));
  NOR2_X1    g01469(.A1(new_n2471_), .A2(\A[114] ), .ZN(new_n2472_));
  OAI21_X1   g01470(.A1(new_n2470_), .A2(new_n2472_), .B(\A[112] ), .ZN(new_n2473_));
  INV_X1     g01471(.I(\A[112] ), .ZN(new_n2474_));
  NOR2_X1    g01472(.A1(\A[113] ), .A2(\A[114] ), .ZN(new_n2475_));
  NAND2_X1   g01473(.A1(\A[113] ), .A2(\A[114] ), .ZN(new_n2476_));
  INV_X1     g01474(.I(new_n2476_), .ZN(new_n2477_));
  OAI21_X1   g01475(.A1(new_n2477_), .A2(new_n2475_), .B(new_n2474_), .ZN(new_n2478_));
  NAND4_X1   g01476(.A1(new_n2463_), .A2(new_n2468_), .A3(new_n2473_), .A4(new_n2478_), .ZN(new_n2479_));
  NAND2_X1   g01477(.A1(new_n2461_), .A2(\A[111] ), .ZN(new_n2480_));
  NAND2_X1   g01478(.A1(new_n2459_), .A2(\A[110] ), .ZN(new_n2481_));
  AOI21_X1   g01479(.A1(new_n2480_), .A2(new_n2481_), .B(new_n2464_), .ZN(new_n2482_));
  INV_X1     g01480(.I(new_n2465_), .ZN(new_n2483_));
  AOI21_X1   g01481(.A1(new_n2483_), .A2(new_n2466_), .B(\A[109] ), .ZN(new_n2484_));
  NAND2_X1   g01482(.A1(new_n2471_), .A2(\A[114] ), .ZN(new_n2485_));
  NAND2_X1   g01483(.A1(new_n2469_), .A2(\A[113] ), .ZN(new_n2486_));
  AOI21_X1   g01484(.A1(new_n2485_), .A2(new_n2486_), .B(new_n2474_), .ZN(new_n2487_));
  INV_X1     g01485(.I(new_n2475_), .ZN(new_n2488_));
  AOI21_X1   g01486(.A1(new_n2488_), .A2(new_n2476_), .B(\A[112] ), .ZN(new_n2489_));
  OAI22_X1   g01487(.A1(new_n2482_), .A2(new_n2484_), .B1(new_n2489_), .B2(new_n2487_), .ZN(new_n2490_));
  NAND2_X1   g01488(.A1(new_n2490_), .A2(new_n2479_), .ZN(new_n2491_));
  INV_X1     g01489(.I(\A[103] ), .ZN(new_n2492_));
  INV_X1     g01490(.I(\A[104] ), .ZN(new_n2493_));
  NAND2_X1   g01491(.A1(new_n2493_), .A2(\A[105] ), .ZN(new_n2494_));
  INV_X1     g01492(.I(\A[105] ), .ZN(new_n2495_));
  NAND2_X1   g01493(.A1(new_n2495_), .A2(\A[104] ), .ZN(new_n2496_));
  AOI21_X1   g01494(.A1(new_n2494_), .A2(new_n2496_), .B(new_n2492_), .ZN(new_n2497_));
  NAND2_X1   g01495(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n2498_));
  NOR2_X1    g01496(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n2499_));
  INV_X1     g01497(.I(new_n2499_), .ZN(new_n2500_));
  AOI21_X1   g01498(.A1(new_n2500_), .A2(new_n2498_), .B(\A[103] ), .ZN(new_n2501_));
  INV_X1     g01499(.I(\A[106] ), .ZN(new_n2502_));
  INV_X1     g01500(.I(\A[107] ), .ZN(new_n2503_));
  NAND2_X1   g01501(.A1(new_n2503_), .A2(\A[108] ), .ZN(new_n2504_));
  INV_X1     g01502(.I(\A[108] ), .ZN(new_n2505_));
  NAND2_X1   g01503(.A1(new_n2505_), .A2(\A[107] ), .ZN(new_n2506_));
  AOI21_X1   g01504(.A1(new_n2504_), .A2(new_n2506_), .B(new_n2502_), .ZN(new_n2507_));
  NAND2_X1   g01505(.A1(\A[107] ), .A2(\A[108] ), .ZN(new_n2508_));
  OR2_X2     g01506(.A1(\A[107] ), .A2(\A[108] ), .Z(new_n2509_));
  AOI21_X1   g01507(.A1(new_n2509_), .A2(new_n2508_), .B(\A[106] ), .ZN(new_n2510_));
  NOR4_X1    g01508(.A1(new_n2497_), .A2(new_n2501_), .A3(new_n2507_), .A4(new_n2510_), .ZN(new_n2511_));
  NOR2_X1    g01509(.A1(new_n2495_), .A2(\A[104] ), .ZN(new_n2512_));
  NOR2_X1    g01510(.A1(new_n2493_), .A2(\A[105] ), .ZN(new_n2513_));
  OAI21_X1   g01511(.A1(new_n2512_), .A2(new_n2513_), .B(\A[103] ), .ZN(new_n2514_));
  INV_X1     g01512(.I(new_n2498_), .ZN(new_n2515_));
  OAI21_X1   g01513(.A1(new_n2515_), .A2(new_n2499_), .B(new_n2492_), .ZN(new_n2516_));
  NOR2_X1    g01514(.A1(new_n2505_), .A2(\A[107] ), .ZN(new_n2517_));
  NOR2_X1    g01515(.A1(new_n2503_), .A2(\A[108] ), .ZN(new_n2518_));
  OAI21_X1   g01516(.A1(new_n2517_), .A2(new_n2518_), .B(\A[106] ), .ZN(new_n2519_));
  INV_X1     g01517(.I(new_n2508_), .ZN(new_n2520_));
  NOR2_X1    g01518(.A1(\A[107] ), .A2(\A[108] ), .ZN(new_n2521_));
  OAI21_X1   g01519(.A1(new_n2520_), .A2(new_n2521_), .B(new_n2502_), .ZN(new_n2522_));
  AOI22_X1   g01520(.A1(new_n2514_), .A2(new_n2516_), .B1(new_n2519_), .B2(new_n2522_), .ZN(new_n2523_));
  NOR2_X1    g01521(.A1(new_n2523_), .A2(new_n2511_), .ZN(new_n2524_));
  NOR2_X1    g01522(.A1(new_n2491_), .A2(new_n2524_), .ZN(new_n2525_));
  NOR4_X1    g01523(.A1(new_n2482_), .A2(new_n2484_), .A3(new_n2489_), .A4(new_n2487_), .ZN(new_n2526_));
  AOI22_X1   g01524(.A1(new_n2463_), .A2(new_n2468_), .B1(new_n2473_), .B2(new_n2478_), .ZN(new_n2527_));
  NOR2_X1    g01525(.A1(new_n2527_), .A2(new_n2526_), .ZN(new_n2528_));
  NAND4_X1   g01526(.A1(new_n2514_), .A2(new_n2516_), .A3(new_n2519_), .A4(new_n2522_), .ZN(new_n2529_));
  OAI22_X1   g01527(.A1(new_n2497_), .A2(new_n2501_), .B1(new_n2507_), .B2(new_n2510_), .ZN(new_n2530_));
  NAND2_X1   g01528(.A1(new_n2529_), .A2(new_n2530_), .ZN(new_n2531_));
  NOR2_X1    g01529(.A1(new_n2528_), .A2(new_n2531_), .ZN(new_n2532_));
  OAI22_X1   g01530(.A1(new_n2525_), .A2(new_n2532_), .B1(new_n2451_), .B2(new_n2458_), .ZN(new_n2533_));
  NAND2_X1   g01531(.A1(new_n2454_), .A2(new_n2457_), .ZN(new_n2534_));
  NAND2_X1   g01532(.A1(new_n2417_), .A2(new_n2450_), .ZN(new_n2535_));
  NOR2_X1    g01533(.A1(new_n2532_), .A2(new_n2525_), .ZN(new_n2536_));
  NAND3_X1   g01534(.A1(new_n2536_), .A2(new_n2534_), .A3(new_n2535_), .ZN(new_n2537_));
  NAND2_X1   g01535(.A1(new_n2537_), .A2(new_n2533_), .ZN(new_n2538_));
  INV_X1     g01536(.I(\A[98] ), .ZN(new_n2539_));
  NAND2_X1   g01537(.A1(new_n2539_), .A2(\A[99] ), .ZN(new_n2540_));
  INV_X1     g01538(.I(\A[99] ), .ZN(new_n2541_));
  NAND2_X1   g01539(.A1(new_n2541_), .A2(\A[98] ), .ZN(new_n2542_));
  NAND2_X1   g01540(.A1(new_n2540_), .A2(new_n2542_), .ZN(new_n2543_));
  NAND2_X1   g01541(.A1(new_n2543_), .A2(\A[97] ), .ZN(new_n2544_));
  INV_X1     g01542(.I(\A[97] ), .ZN(new_n2545_));
  NOR2_X1    g01543(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n2546_));
  NAND2_X1   g01544(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n2547_));
  INV_X1     g01545(.I(new_n2547_), .ZN(new_n2548_));
  OAI21_X1   g01546(.A1(new_n2548_), .A2(new_n2546_), .B(new_n2545_), .ZN(new_n2549_));
  INV_X1     g01547(.I(\A[102] ), .ZN(new_n2550_));
  NOR2_X1    g01548(.A1(new_n2550_), .A2(\A[101] ), .ZN(new_n2551_));
  INV_X1     g01549(.I(\A[101] ), .ZN(new_n2552_));
  NOR2_X1    g01550(.A1(new_n2552_), .A2(\A[102] ), .ZN(new_n2553_));
  OAI21_X1   g01551(.A1(new_n2551_), .A2(new_n2553_), .B(\A[100] ), .ZN(new_n2554_));
  INV_X1     g01552(.I(\A[100] ), .ZN(new_n2555_));
  NOR2_X1    g01553(.A1(\A[101] ), .A2(\A[102] ), .ZN(new_n2556_));
  NAND2_X1   g01554(.A1(\A[101] ), .A2(\A[102] ), .ZN(new_n2557_));
  INV_X1     g01555(.I(new_n2557_), .ZN(new_n2558_));
  OAI21_X1   g01556(.A1(new_n2558_), .A2(new_n2556_), .B(new_n2555_), .ZN(new_n2559_));
  NAND4_X1   g01557(.A1(new_n2544_), .A2(new_n2549_), .A3(new_n2559_), .A4(new_n2554_), .ZN(new_n2560_));
  AOI21_X1   g01558(.A1(new_n2540_), .A2(new_n2542_), .B(new_n2545_), .ZN(new_n2561_));
  INV_X1     g01559(.I(new_n2546_), .ZN(new_n2562_));
  AOI21_X1   g01560(.A1(new_n2562_), .A2(new_n2547_), .B(\A[97] ), .ZN(new_n2563_));
  NAND2_X1   g01561(.A1(new_n2552_), .A2(\A[102] ), .ZN(new_n2564_));
  NAND2_X1   g01562(.A1(new_n2550_), .A2(\A[101] ), .ZN(new_n2565_));
  AOI21_X1   g01563(.A1(new_n2564_), .A2(new_n2565_), .B(new_n2555_), .ZN(new_n2566_));
  INV_X1     g01564(.I(new_n2556_), .ZN(new_n2567_));
  AOI21_X1   g01565(.A1(new_n2567_), .A2(new_n2557_), .B(\A[100] ), .ZN(new_n2568_));
  OAI22_X1   g01566(.A1(new_n2561_), .A2(new_n2563_), .B1(new_n2568_), .B2(new_n2566_), .ZN(new_n2569_));
  NAND2_X1   g01567(.A1(new_n2560_), .A2(new_n2569_), .ZN(new_n2570_));
  INV_X1     g01568(.I(\A[93] ), .ZN(new_n2571_));
  NOR2_X1    g01569(.A1(new_n2571_), .A2(\A[92] ), .ZN(new_n2572_));
  INV_X1     g01570(.I(\A[92] ), .ZN(new_n2573_));
  NOR2_X1    g01571(.A1(new_n2573_), .A2(\A[93] ), .ZN(new_n2574_));
  OAI21_X1   g01572(.A1(new_n2572_), .A2(new_n2574_), .B(\A[91] ), .ZN(new_n2575_));
  INV_X1     g01573(.I(\A[91] ), .ZN(new_n2576_));
  NAND2_X1   g01574(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n2577_));
  INV_X1     g01575(.I(new_n2577_), .ZN(new_n2578_));
  NOR2_X1    g01576(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n2579_));
  OAI21_X1   g01577(.A1(new_n2578_), .A2(new_n2579_), .B(new_n2576_), .ZN(new_n2580_));
  INV_X1     g01578(.I(\A[96] ), .ZN(new_n2581_));
  NOR2_X1    g01579(.A1(new_n2581_), .A2(\A[95] ), .ZN(new_n2582_));
  INV_X1     g01580(.I(\A[95] ), .ZN(new_n2583_));
  NOR2_X1    g01581(.A1(new_n2583_), .A2(\A[96] ), .ZN(new_n2584_));
  OAI21_X1   g01582(.A1(new_n2582_), .A2(new_n2584_), .B(\A[94] ), .ZN(new_n2585_));
  INV_X1     g01583(.I(\A[94] ), .ZN(new_n2586_));
  NAND2_X1   g01584(.A1(\A[95] ), .A2(\A[96] ), .ZN(new_n2587_));
  INV_X1     g01585(.I(new_n2587_), .ZN(new_n2588_));
  NOR2_X1    g01586(.A1(\A[95] ), .A2(\A[96] ), .ZN(new_n2589_));
  OAI21_X1   g01587(.A1(new_n2588_), .A2(new_n2589_), .B(new_n2586_), .ZN(new_n2590_));
  NAND4_X1   g01588(.A1(new_n2575_), .A2(new_n2580_), .A3(new_n2585_), .A4(new_n2590_), .ZN(new_n2591_));
  INV_X1     g01589(.I(new_n2572_), .ZN(new_n2592_));
  NAND2_X1   g01590(.A1(new_n2571_), .A2(\A[92] ), .ZN(new_n2593_));
  AOI21_X1   g01591(.A1(new_n2592_), .A2(new_n2593_), .B(new_n2576_), .ZN(new_n2594_));
  INV_X1     g01592(.I(new_n2579_), .ZN(new_n2595_));
  AOI21_X1   g01593(.A1(new_n2595_), .A2(new_n2577_), .B(\A[91] ), .ZN(new_n2596_));
  NAND2_X1   g01594(.A1(new_n2583_), .A2(\A[96] ), .ZN(new_n2597_));
  NAND2_X1   g01595(.A1(new_n2581_), .A2(\A[95] ), .ZN(new_n2598_));
  AOI21_X1   g01596(.A1(new_n2597_), .A2(new_n2598_), .B(new_n2586_), .ZN(new_n2599_));
  INV_X1     g01597(.I(new_n2589_), .ZN(new_n2600_));
  AOI21_X1   g01598(.A1(new_n2600_), .A2(new_n2587_), .B(\A[94] ), .ZN(new_n2601_));
  OAI22_X1   g01599(.A1(new_n2594_), .A2(new_n2596_), .B1(new_n2601_), .B2(new_n2599_), .ZN(new_n2602_));
  NAND2_X1   g01600(.A1(new_n2602_), .A2(new_n2591_), .ZN(new_n2603_));
  INV_X1     g01601(.I(new_n2603_), .ZN(new_n2604_));
  NOR2_X1    g01602(.A1(new_n2604_), .A2(new_n2570_), .ZN(new_n2605_));
  NOR4_X1    g01603(.A1(new_n2561_), .A2(new_n2563_), .A3(new_n2568_), .A4(new_n2566_), .ZN(new_n2606_));
  AOI22_X1   g01604(.A1(new_n2544_), .A2(new_n2549_), .B1(new_n2559_), .B2(new_n2554_), .ZN(new_n2607_));
  NOR2_X1    g01605(.A1(new_n2607_), .A2(new_n2606_), .ZN(new_n2608_));
  NOR2_X1    g01606(.A1(new_n2608_), .A2(new_n2603_), .ZN(new_n2609_));
  INV_X1     g01607(.I(\A[86] ), .ZN(new_n2610_));
  NAND2_X1   g01608(.A1(new_n2610_), .A2(\A[87] ), .ZN(new_n2611_));
  INV_X1     g01609(.I(new_n2611_), .ZN(new_n2612_));
  NOR2_X1    g01610(.A1(new_n2610_), .A2(\A[87] ), .ZN(new_n2613_));
  OAI21_X1   g01611(.A1(new_n2612_), .A2(new_n2613_), .B(\A[85] ), .ZN(new_n2614_));
  INV_X1     g01612(.I(\A[85] ), .ZN(new_n2615_));
  NOR2_X1    g01613(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n2616_));
  NAND2_X1   g01614(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n2617_));
  INV_X1     g01615(.I(new_n2617_), .ZN(new_n2618_));
  OAI21_X1   g01616(.A1(new_n2618_), .A2(new_n2616_), .B(new_n2615_), .ZN(new_n2619_));
  INV_X1     g01617(.I(\A[90] ), .ZN(new_n2620_));
  NOR2_X1    g01618(.A1(new_n2620_), .A2(\A[89] ), .ZN(new_n2621_));
  INV_X1     g01619(.I(\A[89] ), .ZN(new_n2622_));
  NOR2_X1    g01620(.A1(new_n2622_), .A2(\A[90] ), .ZN(new_n2623_));
  OAI21_X1   g01621(.A1(new_n2621_), .A2(new_n2623_), .B(\A[88] ), .ZN(new_n2624_));
  INV_X1     g01622(.I(\A[88] ), .ZN(new_n2625_));
  NOR2_X1    g01623(.A1(\A[89] ), .A2(\A[90] ), .ZN(new_n2626_));
  NAND2_X1   g01624(.A1(\A[89] ), .A2(\A[90] ), .ZN(new_n2627_));
  INV_X1     g01625(.I(new_n2627_), .ZN(new_n2628_));
  OAI21_X1   g01626(.A1(new_n2628_), .A2(new_n2626_), .B(new_n2625_), .ZN(new_n2629_));
  NAND4_X1   g01627(.A1(new_n2614_), .A2(new_n2619_), .A3(new_n2629_), .A4(new_n2624_), .ZN(new_n2630_));
  INV_X1     g01628(.I(\A[87] ), .ZN(new_n2631_));
  NAND2_X1   g01629(.A1(new_n2631_), .A2(\A[86] ), .ZN(new_n2632_));
  AOI21_X1   g01630(.A1(new_n2611_), .A2(new_n2632_), .B(new_n2615_), .ZN(new_n2633_));
  INV_X1     g01631(.I(new_n2616_), .ZN(new_n2634_));
  AOI21_X1   g01632(.A1(new_n2634_), .A2(new_n2617_), .B(\A[85] ), .ZN(new_n2635_));
  NAND2_X1   g01633(.A1(new_n2622_), .A2(\A[90] ), .ZN(new_n2636_));
  NAND2_X1   g01634(.A1(new_n2620_), .A2(\A[89] ), .ZN(new_n2637_));
  AOI21_X1   g01635(.A1(new_n2636_), .A2(new_n2637_), .B(new_n2625_), .ZN(new_n2638_));
  INV_X1     g01636(.I(new_n2626_), .ZN(new_n2639_));
  AOI21_X1   g01637(.A1(new_n2639_), .A2(new_n2627_), .B(\A[88] ), .ZN(new_n2640_));
  OAI22_X1   g01638(.A1(new_n2633_), .A2(new_n2635_), .B1(new_n2640_), .B2(new_n2638_), .ZN(new_n2641_));
  NAND2_X1   g01639(.A1(new_n2630_), .A2(new_n2641_), .ZN(new_n2642_));
  INV_X1     g01640(.I(\A[79] ), .ZN(new_n2643_));
  INV_X1     g01641(.I(\A[80] ), .ZN(new_n2644_));
  NAND2_X1   g01642(.A1(new_n2644_), .A2(\A[81] ), .ZN(new_n2645_));
  INV_X1     g01643(.I(\A[81] ), .ZN(new_n2646_));
  NAND2_X1   g01644(.A1(new_n2646_), .A2(\A[80] ), .ZN(new_n2647_));
  AOI21_X1   g01645(.A1(new_n2645_), .A2(new_n2647_), .B(new_n2643_), .ZN(new_n2648_));
  NAND2_X1   g01646(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n2649_));
  NOR2_X1    g01647(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n2650_));
  INV_X1     g01648(.I(new_n2650_), .ZN(new_n2651_));
  AOI21_X1   g01649(.A1(new_n2651_), .A2(new_n2649_), .B(\A[79] ), .ZN(new_n2652_));
  INV_X1     g01650(.I(\A[82] ), .ZN(new_n2653_));
  INV_X1     g01651(.I(\A[83] ), .ZN(new_n2654_));
  NAND2_X1   g01652(.A1(new_n2654_), .A2(\A[84] ), .ZN(new_n2655_));
  INV_X1     g01653(.I(\A[84] ), .ZN(new_n2656_));
  NAND2_X1   g01654(.A1(new_n2656_), .A2(\A[83] ), .ZN(new_n2657_));
  AOI21_X1   g01655(.A1(new_n2655_), .A2(new_n2657_), .B(new_n2653_), .ZN(new_n2658_));
  NAND2_X1   g01656(.A1(\A[83] ), .A2(\A[84] ), .ZN(new_n2659_));
  NOR2_X1    g01657(.A1(\A[83] ), .A2(\A[84] ), .ZN(new_n2660_));
  INV_X1     g01658(.I(new_n2660_), .ZN(new_n2661_));
  AOI21_X1   g01659(.A1(new_n2661_), .A2(new_n2659_), .B(\A[82] ), .ZN(new_n2662_));
  NOR4_X1    g01660(.A1(new_n2648_), .A2(new_n2652_), .A3(new_n2662_), .A4(new_n2658_), .ZN(new_n2663_));
  NOR2_X1    g01661(.A1(new_n2646_), .A2(\A[80] ), .ZN(new_n2664_));
  NOR2_X1    g01662(.A1(new_n2644_), .A2(\A[81] ), .ZN(new_n2665_));
  OAI21_X1   g01663(.A1(new_n2664_), .A2(new_n2665_), .B(\A[79] ), .ZN(new_n2666_));
  INV_X1     g01664(.I(new_n2649_), .ZN(new_n2667_));
  OAI21_X1   g01665(.A1(new_n2667_), .A2(new_n2650_), .B(new_n2643_), .ZN(new_n2668_));
  NOR2_X1    g01666(.A1(new_n2656_), .A2(\A[83] ), .ZN(new_n2669_));
  NOR2_X1    g01667(.A1(new_n2654_), .A2(\A[84] ), .ZN(new_n2670_));
  OAI21_X1   g01668(.A1(new_n2669_), .A2(new_n2670_), .B(\A[82] ), .ZN(new_n2671_));
  INV_X1     g01669(.I(new_n2659_), .ZN(new_n2672_));
  OAI21_X1   g01670(.A1(new_n2672_), .A2(new_n2660_), .B(new_n2653_), .ZN(new_n2673_));
  AOI22_X1   g01671(.A1(new_n2666_), .A2(new_n2668_), .B1(new_n2671_), .B2(new_n2673_), .ZN(new_n2674_));
  NOR2_X1    g01672(.A1(new_n2674_), .A2(new_n2663_), .ZN(new_n2675_));
  NOR2_X1    g01673(.A1(new_n2675_), .A2(new_n2642_), .ZN(new_n2676_));
  NOR4_X1    g01674(.A1(new_n2633_), .A2(new_n2635_), .A3(new_n2640_), .A4(new_n2638_), .ZN(new_n2677_));
  AOI22_X1   g01675(.A1(new_n2614_), .A2(new_n2619_), .B1(new_n2629_), .B2(new_n2624_), .ZN(new_n2678_));
  NOR2_X1    g01676(.A1(new_n2678_), .A2(new_n2677_), .ZN(new_n2679_));
  NAND4_X1   g01677(.A1(new_n2666_), .A2(new_n2668_), .A3(new_n2671_), .A4(new_n2673_), .ZN(new_n2680_));
  OAI22_X1   g01678(.A1(new_n2648_), .A2(new_n2652_), .B1(new_n2662_), .B2(new_n2658_), .ZN(new_n2681_));
  NAND2_X1   g01679(.A1(new_n2681_), .A2(new_n2680_), .ZN(new_n2682_));
  NOR2_X1    g01680(.A1(new_n2679_), .A2(new_n2682_), .ZN(new_n2683_));
  OAI22_X1   g01681(.A1(new_n2605_), .A2(new_n2609_), .B1(new_n2676_), .B2(new_n2683_), .ZN(new_n2684_));
  NAND2_X1   g01682(.A1(new_n2608_), .A2(new_n2603_), .ZN(new_n2685_));
  INV_X1     g01683(.I(new_n2609_), .ZN(new_n2686_));
  NOR2_X1    g01684(.A1(new_n2676_), .A2(new_n2683_), .ZN(new_n2687_));
  NAND3_X1   g01685(.A1(new_n2687_), .A2(new_n2686_), .A3(new_n2685_), .ZN(new_n2688_));
  NAND2_X1   g01686(.A1(new_n2688_), .A2(new_n2684_), .ZN(new_n2689_));
  NOR2_X1    g01687(.A1(new_n2689_), .A2(new_n2538_), .ZN(new_n2690_));
  NAND2_X1   g01688(.A1(new_n2689_), .A2(new_n2538_), .ZN(new_n2691_));
  INV_X1     g01689(.I(new_n2691_), .ZN(new_n2692_));
  NOR2_X1    g01690(.A1(new_n2692_), .A2(new_n2690_), .ZN(new_n2693_));
  NAND2_X1   g01691(.A1(new_n2693_), .A2(new_n2384_), .ZN(new_n2694_));
  NOR2_X1    g01692(.A1(new_n2693_), .A2(new_n2384_), .ZN(new_n2695_));
  INV_X1     g01693(.I(new_n2695_), .ZN(new_n2696_));
  NAND2_X1   g01694(.A1(new_n2696_), .A2(new_n2694_), .ZN(new_n2697_));
  NOR2_X1    g01695(.A1(new_n2068_), .A2(new_n2697_), .ZN(new_n2698_));
  AOI21_X1   g01696(.A1(\A[143] ), .A2(\A[144] ), .B(\A[142] ), .ZN(new_n2699_));
  NOR2_X1    g01697(.A1(new_n2699_), .A2(new_n2266_), .ZN(new_n2700_));
  AOI21_X1   g01698(.A1(\A[140] ), .A2(\A[141] ), .B(\A[139] ), .ZN(new_n2701_));
  NOR2_X1    g01699(.A1(new_n2701_), .A2(new_n2256_), .ZN(new_n2702_));
  NOR2_X1    g01700(.A1(new_n2700_), .A2(new_n2702_), .ZN(new_n2703_));
  NOR4_X1    g01701(.A1(new_n2699_), .A2(new_n2701_), .A3(new_n2256_), .A4(new_n2266_), .ZN(new_n2704_));
  NOR2_X1    g01702(.A1(new_n2703_), .A2(new_n2704_), .ZN(new_n2705_));
  NAND2_X1   g01703(.A1(new_n2268_), .A2(new_n2705_), .ZN(new_n2706_));
  OAI22_X1   g01704(.A1(new_n2256_), .A2(new_n2701_), .B1(new_n2699_), .B2(new_n2266_), .ZN(new_n2707_));
  INV_X1     g01705(.I(new_n2704_), .ZN(new_n2708_));
  NAND2_X1   g01706(.A1(new_n2708_), .A2(new_n2707_), .ZN(new_n2709_));
  NAND2_X1   g01707(.A1(new_n2294_), .A2(new_n2709_), .ZN(new_n2710_));
  NAND2_X1   g01708(.A1(new_n2710_), .A2(new_n2706_), .ZN(new_n2711_));
  AOI21_X1   g01709(.A1(\A[149] ), .A2(\A[150] ), .B(\A[148] ), .ZN(new_n2712_));
  NOR2_X1    g01710(.A1(new_n2712_), .A2(new_n2240_), .ZN(new_n2713_));
  AOI21_X1   g01711(.A1(\A[146] ), .A2(\A[147] ), .B(\A[145] ), .ZN(new_n2714_));
  NOR2_X1    g01712(.A1(new_n2714_), .A2(new_n2230_), .ZN(new_n2715_));
  XOR2_X1    g01713(.A1(new_n2713_), .A2(new_n2715_), .Z(new_n2716_));
  NOR2_X1    g01714(.A1(new_n2716_), .A2(new_n2244_), .ZN(new_n2717_));
  NOR3_X1    g01715(.A1(new_n2715_), .A2(new_n2240_), .A3(new_n2712_), .ZN(new_n2718_));
  NOR3_X1    g01716(.A1(new_n2713_), .A2(new_n2230_), .A3(new_n2714_), .ZN(new_n2719_));
  NOR2_X1    g01717(.A1(new_n2718_), .A2(new_n2719_), .ZN(new_n2720_));
  NOR2_X1    g01718(.A1(new_n2292_), .A2(new_n2720_), .ZN(new_n2721_));
  NOR2_X1    g01719(.A1(new_n2717_), .A2(new_n2721_), .ZN(new_n2722_));
  NOR2_X1    g01720(.A1(new_n2293_), .A2(new_n2280_), .ZN(new_n2723_));
  NOR2_X1    g01721(.A1(new_n2722_), .A2(new_n2723_), .ZN(new_n2724_));
  NAND4_X1   g01722(.A1(new_n2292_), .A2(new_n2245_), .A3(new_n2279_), .A4(new_n2268_), .ZN(new_n2725_));
  NOR3_X1    g01723(.A1(new_n2725_), .A2(new_n2717_), .A3(new_n2721_), .ZN(new_n2726_));
  NOR3_X1    g01724(.A1(new_n2724_), .A2(new_n2711_), .A3(new_n2726_), .ZN(new_n2727_));
  NOR2_X1    g01725(.A1(new_n2294_), .A2(new_n2709_), .ZN(new_n2728_));
  NOR2_X1    g01726(.A1(new_n2268_), .A2(new_n2705_), .ZN(new_n2729_));
  NOR2_X1    g01727(.A1(new_n2728_), .A2(new_n2729_), .ZN(new_n2730_));
  OAI21_X1   g01728(.A1(new_n2717_), .A2(new_n2721_), .B(new_n2725_), .ZN(new_n2731_));
  NAND4_X1   g01729(.A1(new_n2298_), .A2(new_n2292_), .A3(new_n2245_), .A4(new_n2716_), .ZN(new_n2732_));
  AOI21_X1   g01730(.A1(new_n2731_), .A2(new_n2732_), .B(new_n2730_), .ZN(new_n2733_));
  NOR2_X1    g01731(.A1(new_n2727_), .A2(new_n2733_), .ZN(new_n2734_));
  OAI22_X1   g01732(.A1(new_n2376_), .A2(new_n2375_), .B1(new_n2377_), .B2(new_n2378_), .ZN(new_n2735_));
  AOI21_X1   g01733(.A1(\A[131] ), .A2(\A[132] ), .B(\A[130] ), .ZN(new_n2736_));
  NOR2_X1    g01734(.A1(new_n2736_), .A2(new_n2351_), .ZN(new_n2737_));
  AOI21_X1   g01735(.A1(\A[128] ), .A2(\A[129] ), .B(\A[127] ), .ZN(new_n2738_));
  NOR2_X1    g01736(.A1(new_n2738_), .A2(new_n2341_), .ZN(new_n2739_));
  NOR2_X1    g01737(.A1(new_n2737_), .A2(new_n2739_), .ZN(new_n2740_));
  NOR4_X1    g01738(.A1(new_n2736_), .A2(new_n2738_), .A3(new_n2341_), .A4(new_n2351_), .ZN(new_n2741_));
  NOR2_X1    g01739(.A1(new_n2740_), .A2(new_n2741_), .ZN(new_n2742_));
  NAND2_X1   g01740(.A1(new_n2353_), .A2(new_n2742_), .ZN(new_n2743_));
  OAI22_X1   g01741(.A1(new_n2341_), .A2(new_n2738_), .B1(new_n2736_), .B2(new_n2351_), .ZN(new_n2744_));
  INV_X1     g01742(.I(new_n2741_), .ZN(new_n2745_));
  NAND2_X1   g01743(.A1(new_n2745_), .A2(new_n2744_), .ZN(new_n2746_));
  NAND2_X1   g01744(.A1(new_n2370_), .A2(new_n2746_), .ZN(new_n2747_));
  NAND2_X1   g01745(.A1(new_n2747_), .A2(new_n2743_), .ZN(new_n2748_));
  AOI21_X1   g01746(.A1(\A[137] ), .A2(\A[138] ), .B(\A[136] ), .ZN(new_n2749_));
  NOR2_X1    g01747(.A1(new_n2749_), .A2(new_n2316_), .ZN(new_n2750_));
  AOI21_X1   g01748(.A1(\A[134] ), .A2(\A[135] ), .B(\A[133] ), .ZN(new_n2751_));
  NOR2_X1    g01749(.A1(new_n2751_), .A2(new_n2306_), .ZN(new_n2752_));
  XOR2_X1    g01750(.A1(new_n2750_), .A2(new_n2752_), .Z(new_n2753_));
  NOR2_X1    g01751(.A1(new_n2753_), .A2(new_n2320_), .ZN(new_n2754_));
  NOR3_X1    g01752(.A1(new_n2752_), .A2(new_n2316_), .A3(new_n2749_), .ZN(new_n2755_));
  NOR3_X1    g01753(.A1(new_n2750_), .A2(new_n2306_), .A3(new_n2751_), .ZN(new_n2756_));
  NOR2_X1    g01754(.A1(new_n2755_), .A2(new_n2756_), .ZN(new_n2757_));
  NOR2_X1    g01755(.A1(new_n2367_), .A2(new_n2757_), .ZN(new_n2758_));
  NOR2_X1    g01756(.A1(new_n2754_), .A2(new_n2758_), .ZN(new_n2759_));
  NOR4_X1    g01757(.A1(new_n2320_), .A2(new_n2331_), .A3(new_n2371_), .A4(new_n2370_), .ZN(new_n2760_));
  OAI21_X1   g01758(.A1(new_n2759_), .A2(new_n2760_), .B(new_n2748_), .ZN(new_n2761_));
  NOR4_X1    g01759(.A1(new_n2365_), .A2(new_n2320_), .A3(new_n2331_), .A4(new_n2757_), .ZN(new_n2762_));
  NOR2_X1    g01760(.A1(new_n2761_), .A2(new_n2762_), .ZN(new_n2763_));
  OAI22_X1   g01761(.A1(new_n2754_), .A2(new_n2758_), .B1(new_n2369_), .B2(new_n2365_), .ZN(new_n2764_));
  NAND2_X1   g01762(.A1(new_n2759_), .A2(new_n2760_), .ZN(new_n2765_));
  AOI21_X1   g01763(.A1(new_n2765_), .A2(new_n2764_), .B(new_n2748_), .ZN(new_n2766_));
  NOR3_X1    g01764(.A1(new_n2763_), .A2(new_n2766_), .A3(new_n2735_), .ZN(new_n2767_));
  NAND3_X1   g01765(.A1(new_n2765_), .A2(new_n2764_), .A3(new_n2748_), .ZN(new_n2768_));
  NOR2_X1    g01766(.A1(new_n2370_), .A2(new_n2746_), .ZN(new_n2769_));
  NOR2_X1    g01767(.A1(new_n2353_), .A2(new_n2742_), .ZN(new_n2770_));
  NOR2_X1    g01768(.A1(new_n2769_), .A2(new_n2770_), .ZN(new_n2771_));
  NOR2_X1    g01769(.A1(new_n2759_), .A2(new_n2760_), .ZN(new_n2772_));
  OAI21_X1   g01770(.A1(new_n2772_), .A2(new_n2762_), .B(new_n2771_), .ZN(new_n2773_));
  AOI21_X1   g01771(.A1(new_n2773_), .A2(new_n2768_), .B(new_n2374_), .ZN(new_n2774_));
  NOR3_X1    g01772(.A1(new_n2767_), .A2(new_n2774_), .A3(new_n2734_), .ZN(new_n2775_));
  NAND3_X1   g01773(.A1(new_n2731_), .A2(new_n2732_), .A3(new_n2730_), .ZN(new_n2776_));
  OAI21_X1   g01774(.A1(new_n2724_), .A2(new_n2726_), .B(new_n2711_), .ZN(new_n2777_));
  NAND2_X1   g01775(.A1(new_n2777_), .A2(new_n2776_), .ZN(new_n2778_));
  NAND3_X1   g01776(.A1(new_n2773_), .A2(new_n2768_), .A3(new_n2374_), .ZN(new_n2779_));
  OAI21_X1   g01777(.A1(new_n2763_), .A2(new_n2766_), .B(new_n2735_), .ZN(new_n2780_));
  AOI21_X1   g01778(.A1(new_n2780_), .A2(new_n2779_), .B(new_n2778_), .ZN(new_n2781_));
  NOR2_X1    g01779(.A1(new_n2775_), .A2(new_n2781_), .ZN(new_n2782_));
  AOI21_X1   g01780(.A1(\A[155] ), .A2(\A[156] ), .B(\A[154] ), .ZN(new_n2783_));
  NOR2_X1    g01781(.A1(new_n2783_), .A2(new_n2194_), .ZN(new_n2784_));
  AOI21_X1   g01782(.A1(\A[152] ), .A2(\A[153] ), .B(\A[151] ), .ZN(new_n2785_));
  NOR2_X1    g01783(.A1(new_n2785_), .A2(new_n2184_), .ZN(new_n2786_));
  NOR2_X1    g01784(.A1(new_n2784_), .A2(new_n2786_), .ZN(new_n2787_));
  NOR4_X1    g01785(.A1(new_n2783_), .A2(new_n2785_), .A3(new_n2184_), .A4(new_n2194_), .ZN(new_n2788_));
  NOR2_X1    g01786(.A1(new_n2787_), .A2(new_n2788_), .ZN(new_n2789_));
  NAND2_X1   g01787(.A1(new_n2196_), .A2(new_n2789_), .ZN(new_n2790_));
  NOR2_X1    g01788(.A1(new_n2201_), .A2(new_n2199_), .ZN(new_n2791_));
  NOR2_X1    g01789(.A1(new_n2204_), .A2(new_n2206_), .ZN(new_n2792_));
  OAI22_X1   g01790(.A1(new_n2184_), .A2(new_n2785_), .B1(new_n2783_), .B2(new_n2194_), .ZN(new_n2793_));
  NAND2_X1   g01791(.A1(new_n2192_), .A2(new_n2191_), .ZN(new_n2794_));
  NAND2_X1   g01792(.A1(new_n2182_), .A2(new_n2181_), .ZN(new_n2795_));
  NAND4_X1   g01793(.A1(new_n2794_), .A2(new_n2795_), .A3(new_n2200_), .A4(new_n2205_), .ZN(new_n2796_));
  NAND2_X1   g01794(.A1(new_n2796_), .A2(new_n2793_), .ZN(new_n2797_));
  NAND3_X1   g01795(.A1(new_n2797_), .A2(new_n2791_), .A3(new_n2792_), .ZN(new_n2798_));
  NAND2_X1   g01796(.A1(new_n2790_), .A2(new_n2798_), .ZN(new_n2799_));
  AOI21_X1   g01797(.A1(\A[161] ), .A2(\A[162] ), .B(\A[160] ), .ZN(new_n2800_));
  AOI21_X1   g01798(.A1(\A[158] ), .A2(\A[159] ), .B(\A[157] ), .ZN(new_n2801_));
  NOR2_X1    g01799(.A1(new_n2801_), .A2(new_n2149_), .ZN(new_n2802_));
  NOR3_X1    g01800(.A1(new_n2802_), .A2(new_n2159_), .A3(new_n2800_), .ZN(new_n2803_));
  NOR2_X1    g01801(.A1(new_n2800_), .A2(new_n2159_), .ZN(new_n2804_));
  NOR3_X1    g01802(.A1(new_n2804_), .A2(new_n2149_), .A3(new_n2801_), .ZN(new_n2805_));
  NOR3_X1    g01803(.A1(new_n2163_), .A2(new_n2803_), .A3(new_n2805_), .ZN(new_n2806_));
  NOR2_X1    g01804(.A1(new_n2803_), .A2(new_n2805_), .ZN(new_n2807_));
  NOR2_X1    g01805(.A1(new_n2807_), .A2(new_n2210_), .ZN(new_n2808_));
  NOR2_X1    g01806(.A1(new_n2806_), .A2(new_n2808_), .ZN(new_n2809_));
  NOR4_X1    g01807(.A1(new_n2163_), .A2(new_n2214_), .A3(new_n2174_), .A4(new_n2213_), .ZN(new_n2810_));
  OAI21_X1   g01808(.A1(new_n2809_), .A2(new_n2810_), .B(new_n2799_), .ZN(new_n2811_));
  NAND2_X1   g01809(.A1(new_n2807_), .A2(new_n2210_), .ZN(new_n2812_));
  XOR2_X1    g01810(.A1(new_n2804_), .A2(new_n2802_), .Z(new_n2813_));
  NAND2_X1   g01811(.A1(new_n2813_), .A2(new_n2163_), .ZN(new_n2814_));
  NAND2_X1   g01812(.A1(new_n2814_), .A2(new_n2812_), .ZN(new_n2815_));
  NAND4_X1   g01813(.A1(new_n2211_), .A2(new_n2196_), .A3(new_n2207_), .A4(new_n2210_), .ZN(new_n2816_));
  NOR2_X1    g01814(.A1(new_n2815_), .A2(new_n2816_), .ZN(new_n2817_));
  NOR2_X1    g01815(.A1(new_n2809_), .A2(new_n2810_), .ZN(new_n2818_));
  NOR2_X1    g01816(.A1(new_n2818_), .A2(new_n2817_), .ZN(new_n2819_));
  OAI22_X1   g01817(.A1(new_n2819_), .A2(new_n2799_), .B1(new_n2811_), .B2(new_n2817_), .ZN(new_n2820_));
  AOI21_X1   g01818(.A1(\A[167] ), .A2(\A[168] ), .B(\A[166] ), .ZN(new_n2821_));
  NOR2_X1    g01819(.A1(new_n2821_), .A2(new_n2110_), .ZN(new_n2822_));
  AOI21_X1   g01820(.A1(\A[164] ), .A2(\A[165] ), .B(\A[163] ), .ZN(new_n2823_));
  NOR2_X1    g01821(.A1(new_n2823_), .A2(new_n2101_), .ZN(new_n2824_));
  NOR2_X1    g01822(.A1(new_n2822_), .A2(new_n2824_), .ZN(new_n2825_));
  NOR4_X1    g01823(.A1(new_n2821_), .A2(new_n2823_), .A3(new_n2101_), .A4(new_n2110_), .ZN(new_n2826_));
  NOR2_X1    g01824(.A1(new_n2825_), .A2(new_n2826_), .ZN(new_n2827_));
  NAND2_X1   g01825(.A1(new_n2112_), .A2(new_n2827_), .ZN(new_n2828_));
  OAI22_X1   g01826(.A1(new_n2101_), .A2(new_n2823_), .B1(new_n2821_), .B2(new_n2110_), .ZN(new_n2829_));
  NAND2_X1   g01827(.A1(new_n2822_), .A2(new_n2824_), .ZN(new_n2830_));
  NAND2_X1   g01828(.A1(new_n2830_), .A2(new_n2829_), .ZN(new_n2831_));
  NAND2_X1   g01829(.A1(new_n2139_), .A2(new_n2831_), .ZN(new_n2832_));
  NAND2_X1   g01830(.A1(new_n2828_), .A2(new_n2832_), .ZN(new_n2833_));
  AOI21_X1   g01831(.A1(\A[173] ), .A2(\A[174] ), .B(\A[172] ), .ZN(new_n2834_));
  AOI21_X1   g01832(.A1(\A[170] ), .A2(\A[171] ), .B(\A[169] ), .ZN(new_n2835_));
  NOR2_X1    g01833(.A1(new_n2835_), .A2(new_n2075_), .ZN(new_n2836_));
  NOR3_X1    g01834(.A1(new_n2836_), .A2(new_n2085_), .A3(new_n2834_), .ZN(new_n2837_));
  NOR2_X1    g01835(.A1(new_n2834_), .A2(new_n2085_), .ZN(new_n2838_));
  NOR3_X1    g01836(.A1(new_n2838_), .A2(new_n2075_), .A3(new_n2835_), .ZN(new_n2839_));
  NOR2_X1    g01837(.A1(new_n2837_), .A2(new_n2839_), .ZN(new_n2840_));
  NAND2_X1   g01838(.A1(new_n2137_), .A2(new_n2840_), .ZN(new_n2841_));
  XOR2_X1    g01839(.A1(new_n2838_), .A2(new_n2836_), .Z(new_n2842_));
  NAND2_X1   g01840(.A1(new_n2842_), .A2(new_n2089_), .ZN(new_n2843_));
  AOI22_X1   g01841(.A1(new_n2092_), .A2(new_n2141_), .B1(new_n2841_), .B2(new_n2843_), .ZN(new_n2844_));
  NOR4_X1    g01842(.A1(new_n2125_), .A2(new_n2091_), .A3(new_n2089_), .A4(new_n2840_), .ZN(new_n2845_));
  NOR3_X1    g01843(.A1(new_n2844_), .A2(new_n2833_), .A3(new_n2845_), .ZN(new_n2846_));
  NOR2_X1    g01844(.A1(new_n2139_), .A2(new_n2831_), .ZN(new_n2847_));
  NOR2_X1    g01845(.A1(new_n2112_), .A2(new_n2827_), .ZN(new_n2848_));
  NOR2_X1    g01846(.A1(new_n2848_), .A2(new_n2847_), .ZN(new_n2849_));
  NOR2_X1    g01847(.A1(new_n2842_), .A2(new_n2089_), .ZN(new_n2850_));
  NOR2_X1    g01848(.A1(new_n2137_), .A2(new_n2840_), .ZN(new_n2851_));
  OAI22_X1   g01849(.A1(new_n2850_), .A2(new_n2851_), .B1(new_n2138_), .B2(new_n2125_), .ZN(new_n2852_));
  NAND4_X1   g01850(.A1(new_n2141_), .A2(new_n2137_), .A3(new_n2090_), .A4(new_n2842_), .ZN(new_n2853_));
  AOI21_X1   g01851(.A1(new_n2852_), .A2(new_n2853_), .B(new_n2849_), .ZN(new_n2854_));
  OAI21_X1   g01852(.A1(new_n2846_), .A2(new_n2854_), .B(new_n2217_), .ZN(new_n2855_));
  OAI22_X1   g01853(.A1(new_n2219_), .A2(new_n2218_), .B1(new_n2221_), .B2(new_n2220_), .ZN(new_n2856_));
  NAND3_X1   g01854(.A1(new_n2852_), .A2(new_n2849_), .A3(new_n2853_), .ZN(new_n2857_));
  OAI21_X1   g01855(.A1(new_n2844_), .A2(new_n2845_), .B(new_n2833_), .ZN(new_n2858_));
  NAND3_X1   g01856(.A1(new_n2858_), .A2(new_n2856_), .A3(new_n2857_), .ZN(new_n2859_));
  AOI21_X1   g01857(.A1(new_n2855_), .A2(new_n2859_), .B(new_n2820_), .ZN(new_n2860_));
  NOR2_X1    g01858(.A1(new_n2213_), .A2(new_n2797_), .ZN(new_n2861_));
  NOR2_X1    g01859(.A1(new_n2196_), .A2(new_n2789_), .ZN(new_n2862_));
  NOR2_X1    g01860(.A1(new_n2862_), .A2(new_n2861_), .ZN(new_n2863_));
  AOI21_X1   g01861(.A1(new_n2815_), .A2(new_n2816_), .B(new_n2863_), .ZN(new_n2864_));
  NAND2_X1   g01862(.A1(new_n2809_), .A2(new_n2810_), .ZN(new_n2865_));
  NAND2_X1   g01863(.A1(new_n2815_), .A2(new_n2816_), .ZN(new_n2866_));
  NAND2_X1   g01864(.A1(new_n2865_), .A2(new_n2866_), .ZN(new_n2867_));
  AOI22_X1   g01865(.A1(new_n2867_), .A2(new_n2863_), .B1(new_n2864_), .B2(new_n2865_), .ZN(new_n2868_));
  AOI21_X1   g01866(.A1(new_n2858_), .A2(new_n2857_), .B(new_n2856_), .ZN(new_n2869_));
  NOR3_X1    g01867(.A1(new_n2846_), .A2(new_n2217_), .A3(new_n2854_), .ZN(new_n2870_));
  NOR3_X1    g01868(.A1(new_n2868_), .A2(new_n2869_), .A3(new_n2870_), .ZN(new_n2871_));
  OAI21_X1   g01869(.A1(new_n2860_), .A2(new_n2871_), .B(new_n2382_), .ZN(new_n2872_));
  OAI21_X1   g01870(.A1(new_n2869_), .A2(new_n2870_), .B(new_n2868_), .ZN(new_n2873_));
  NAND3_X1   g01871(.A1(new_n2820_), .A2(new_n2855_), .A3(new_n2859_), .ZN(new_n2874_));
  NAND3_X1   g01872(.A1(new_n2873_), .A2(new_n2874_), .A3(new_n2381_), .ZN(new_n2875_));
  NAND2_X1   g01873(.A1(new_n2872_), .A2(new_n2875_), .ZN(new_n2876_));
  NAND2_X1   g01874(.A1(new_n2876_), .A2(new_n2782_), .ZN(new_n2877_));
  AOI21_X1   g01875(.A1(new_n2873_), .A2(new_n2874_), .B(new_n2381_), .ZN(new_n2878_));
  NOR2_X1    g01876(.A1(new_n2878_), .A2(new_n2782_), .ZN(new_n2879_));
  NAND2_X1   g01877(.A1(new_n2879_), .A2(new_n2875_), .ZN(new_n2880_));
  NAND2_X1   g01878(.A1(new_n2877_), .A2(new_n2880_), .ZN(new_n2881_));
  INV_X1     g01879(.I(new_n2694_), .ZN(new_n2882_));
  AOI21_X1   g01880(.A1(\A[107] ), .A2(\A[108] ), .B(\A[106] ), .ZN(new_n2883_));
  NOR2_X1    g01881(.A1(new_n2883_), .A2(new_n2521_), .ZN(new_n2884_));
  AOI21_X1   g01882(.A1(\A[104] ), .A2(\A[105] ), .B(\A[103] ), .ZN(new_n2885_));
  NOR2_X1    g01883(.A1(new_n2885_), .A2(new_n2499_), .ZN(new_n2886_));
  NOR2_X1    g01884(.A1(new_n2884_), .A2(new_n2886_), .ZN(new_n2887_));
  NOR4_X1    g01885(.A1(new_n2883_), .A2(new_n2885_), .A3(new_n2499_), .A4(new_n2521_), .ZN(new_n2888_));
  NOR2_X1    g01886(.A1(new_n2887_), .A2(new_n2888_), .ZN(new_n2889_));
  NAND2_X1   g01887(.A1(new_n2529_), .A2(new_n2889_), .ZN(new_n2890_));
  OAI22_X1   g01888(.A1(new_n2499_), .A2(new_n2885_), .B1(new_n2883_), .B2(new_n2521_), .ZN(new_n2891_));
  NAND2_X1   g01889(.A1(new_n2884_), .A2(new_n2886_), .ZN(new_n2892_));
  NAND2_X1   g01890(.A1(new_n2892_), .A2(new_n2891_), .ZN(new_n2893_));
  NAND2_X1   g01891(.A1(new_n2511_), .A2(new_n2893_), .ZN(new_n2894_));
  NAND2_X1   g01892(.A1(new_n2890_), .A2(new_n2894_), .ZN(new_n2895_));
  AOI21_X1   g01893(.A1(\A[113] ), .A2(\A[114] ), .B(\A[112] ), .ZN(new_n2896_));
  NOR2_X1    g01894(.A1(new_n2896_), .A2(new_n2475_), .ZN(new_n2897_));
  AOI21_X1   g01895(.A1(\A[110] ), .A2(\A[111] ), .B(\A[109] ), .ZN(new_n2898_));
  NOR2_X1    g01896(.A1(new_n2898_), .A2(new_n2465_), .ZN(new_n2899_));
  XOR2_X1    g01897(.A1(new_n2897_), .A2(new_n2899_), .Z(new_n2900_));
  NOR2_X1    g01898(.A1(new_n2900_), .A2(new_n2526_), .ZN(new_n2901_));
  NOR3_X1    g01899(.A1(new_n2899_), .A2(new_n2475_), .A3(new_n2896_), .ZN(new_n2902_));
  NOR3_X1    g01900(.A1(new_n2897_), .A2(new_n2465_), .A3(new_n2898_), .ZN(new_n2903_));
  NOR2_X1    g01901(.A1(new_n2902_), .A2(new_n2903_), .ZN(new_n2904_));
  NOR2_X1    g01902(.A1(new_n2479_), .A2(new_n2904_), .ZN(new_n2905_));
  NOR2_X1    g01903(.A1(new_n2901_), .A2(new_n2905_), .ZN(new_n2906_));
  NOR4_X1    g01904(.A1(new_n2527_), .A2(new_n2523_), .A3(new_n2526_), .A4(new_n2511_), .ZN(new_n2907_));
  OAI21_X1   g01905(.A1(new_n2906_), .A2(new_n2907_), .B(new_n2895_), .ZN(new_n2908_));
  NAND2_X1   g01906(.A1(new_n2479_), .A2(new_n2904_), .ZN(new_n2909_));
  NAND2_X1   g01907(.A1(new_n2900_), .A2(new_n2526_), .ZN(new_n2910_));
  NAND2_X1   g01908(.A1(new_n2910_), .A2(new_n2909_), .ZN(new_n2911_));
  NOR3_X1    g01909(.A1(new_n2911_), .A2(new_n2491_), .A3(new_n2531_), .ZN(new_n2912_));
  OAI22_X1   g01910(.A1(new_n2901_), .A2(new_n2905_), .B1(new_n2491_), .B2(new_n2531_), .ZN(new_n2913_));
  INV_X1     g01911(.I(new_n2913_), .ZN(new_n2914_));
  NOR2_X1    g01912(.A1(new_n2914_), .A2(new_n2912_), .ZN(new_n2915_));
  OAI22_X1   g01913(.A1(new_n2915_), .A2(new_n2895_), .B1(new_n2908_), .B2(new_n2912_), .ZN(new_n2916_));
  NAND2_X1   g01914(.A1(new_n2528_), .A2(new_n2531_), .ZN(new_n2917_));
  NAND2_X1   g01915(.A1(new_n2491_), .A2(new_n2524_), .ZN(new_n2918_));
  AOI22_X1   g01916(.A1(new_n2917_), .A2(new_n2918_), .B1(new_n2535_), .B2(new_n2534_), .ZN(new_n2919_));
  AOI21_X1   g01917(.A1(\A[119] ), .A2(\A[120] ), .B(\A[118] ), .ZN(new_n2920_));
  AOI21_X1   g01918(.A1(\A[116] ), .A2(\A[117] ), .B(\A[115] ), .ZN(new_n2921_));
  OAI22_X1   g01919(.A1(new_n2425_), .A2(new_n2921_), .B1(new_n2920_), .B2(new_n2447_), .ZN(new_n2922_));
  INV_X1     g01920(.I(new_n2922_), .ZN(new_n2923_));
  NOR4_X1    g01921(.A1(new_n2920_), .A2(new_n2921_), .A3(new_n2425_), .A4(new_n2447_), .ZN(new_n2924_));
  NOR2_X1    g01922(.A1(new_n2923_), .A2(new_n2924_), .ZN(new_n2925_));
  NAND2_X1   g01923(.A1(new_n2925_), .A2(new_n2455_), .ZN(new_n2926_));
  OR4_X2     g01924(.A1(new_n2425_), .A2(new_n2920_), .A3(new_n2921_), .A4(new_n2447_), .Z(new_n2927_));
  NAND2_X1   g01925(.A1(new_n2927_), .A2(new_n2922_), .ZN(new_n2928_));
  NAND2_X1   g01926(.A1(new_n2437_), .A2(new_n2928_), .ZN(new_n2929_));
  NAND2_X1   g01927(.A1(new_n2926_), .A2(new_n2929_), .ZN(new_n2930_));
  AOI21_X1   g01928(.A1(\A[125] ), .A2(\A[126] ), .B(\A[124] ), .ZN(new_n2931_));
  AOI21_X1   g01929(.A1(\A[122] ), .A2(\A[123] ), .B(\A[121] ), .ZN(new_n2932_));
  NOR2_X1    g01930(.A1(new_n2932_), .A2(new_n2391_), .ZN(new_n2933_));
  NOR3_X1    g01931(.A1(new_n2933_), .A2(new_n2401_), .A3(new_n2931_), .ZN(new_n2934_));
  NOR2_X1    g01932(.A1(new_n2931_), .A2(new_n2401_), .ZN(new_n2935_));
  NOR3_X1    g01933(.A1(new_n2935_), .A2(new_n2391_), .A3(new_n2932_), .ZN(new_n2936_));
  NOR2_X1    g01934(.A1(new_n2934_), .A2(new_n2936_), .ZN(new_n2937_));
  NAND2_X1   g01935(.A1(new_n2405_), .A2(new_n2937_), .ZN(new_n2938_));
  XOR2_X1    g01936(.A1(new_n2935_), .A2(new_n2933_), .Z(new_n2939_));
  NAND2_X1   g01937(.A1(new_n2939_), .A2(new_n2452_), .ZN(new_n2940_));
  AOI22_X1   g01938(.A1(new_n2938_), .A2(new_n2940_), .B1(new_n2454_), .B2(new_n2450_), .ZN(new_n2941_));
  NOR4_X1    g01939(.A1(new_n2457_), .A2(new_n2452_), .A3(new_n2453_), .A4(new_n2937_), .ZN(new_n2942_));
  NOR3_X1    g01940(.A1(new_n2941_), .A2(new_n2942_), .A3(new_n2930_), .ZN(new_n2943_));
  NOR2_X1    g01941(.A1(new_n2437_), .A2(new_n2928_), .ZN(new_n2944_));
  NOR2_X1    g01942(.A1(new_n2925_), .A2(new_n2455_), .ZN(new_n2945_));
  NOR2_X1    g01943(.A1(new_n2945_), .A2(new_n2944_), .ZN(new_n2946_));
  NOR2_X1    g01944(.A1(new_n2939_), .A2(new_n2452_), .ZN(new_n2947_));
  NOR2_X1    g01945(.A1(new_n2405_), .A2(new_n2937_), .ZN(new_n2948_));
  OAI22_X1   g01946(.A1(new_n2947_), .A2(new_n2948_), .B1(new_n2417_), .B2(new_n2457_), .ZN(new_n2949_));
  NAND4_X1   g01947(.A1(new_n2450_), .A2(new_n2405_), .A3(new_n2416_), .A4(new_n2939_), .ZN(new_n2950_));
  AOI21_X1   g01948(.A1(new_n2949_), .A2(new_n2950_), .B(new_n2946_), .ZN(new_n2951_));
  OAI21_X1   g01949(.A1(new_n2943_), .A2(new_n2951_), .B(new_n2919_), .ZN(new_n2952_));
  NAND3_X1   g01950(.A1(new_n2949_), .A2(new_n2946_), .A3(new_n2950_), .ZN(new_n2953_));
  OAI21_X1   g01951(.A1(new_n2941_), .A2(new_n2942_), .B(new_n2930_), .ZN(new_n2954_));
  NAND3_X1   g01952(.A1(new_n2954_), .A2(new_n2533_), .A3(new_n2953_), .ZN(new_n2955_));
  NAND3_X1   g01953(.A1(new_n2916_), .A2(new_n2955_), .A3(new_n2952_), .ZN(new_n2956_));
  NOR2_X1    g01954(.A1(new_n2511_), .A2(new_n2893_), .ZN(new_n2957_));
  NOR2_X1    g01955(.A1(new_n2529_), .A2(new_n2889_), .ZN(new_n2958_));
  NOR2_X1    g01956(.A1(new_n2958_), .A2(new_n2957_), .ZN(new_n2959_));
  INV_X1     g01957(.I(new_n2907_), .ZN(new_n2960_));
  AOI21_X1   g01958(.A1(new_n2960_), .A2(new_n2911_), .B(new_n2959_), .ZN(new_n2961_));
  NAND2_X1   g01959(.A1(new_n2906_), .A2(new_n2907_), .ZN(new_n2962_));
  NAND2_X1   g01960(.A1(new_n2962_), .A2(new_n2913_), .ZN(new_n2963_));
  AOI22_X1   g01961(.A1(new_n2963_), .A2(new_n2959_), .B1(new_n2961_), .B2(new_n2962_), .ZN(new_n2964_));
  AOI21_X1   g01962(.A1(new_n2954_), .A2(new_n2953_), .B(new_n2533_), .ZN(new_n2965_));
  NOR3_X1    g01963(.A1(new_n2943_), .A2(new_n2951_), .A3(new_n2919_), .ZN(new_n2966_));
  OAI21_X1   g01964(.A1(new_n2965_), .A2(new_n2966_), .B(new_n2964_), .ZN(new_n2967_));
  NAND2_X1   g01965(.A1(new_n2956_), .A2(new_n2967_), .ZN(new_n2968_));
  NOR4_X1    g01966(.A1(new_n2594_), .A2(new_n2596_), .A3(new_n2601_), .A4(new_n2599_), .ZN(new_n2969_));
  AOI21_X1   g01967(.A1(\A[95] ), .A2(\A[96] ), .B(\A[94] ), .ZN(new_n2970_));
  AOI21_X1   g01968(.A1(\A[92] ), .A2(\A[93] ), .B(\A[91] ), .ZN(new_n2971_));
  OAI22_X1   g01969(.A1(new_n2579_), .A2(new_n2971_), .B1(new_n2970_), .B2(new_n2589_), .ZN(new_n2972_));
  NOR4_X1    g01970(.A1(new_n2970_), .A2(new_n2971_), .A3(new_n2579_), .A4(new_n2589_), .ZN(new_n2973_));
  INV_X1     g01971(.I(new_n2973_), .ZN(new_n2974_));
  NAND2_X1   g01972(.A1(new_n2974_), .A2(new_n2972_), .ZN(new_n2975_));
  NOR2_X1    g01973(.A1(new_n2969_), .A2(new_n2975_), .ZN(new_n2976_));
  INV_X1     g01974(.I(new_n2972_), .ZN(new_n2977_));
  NOR2_X1    g01975(.A1(new_n2977_), .A2(new_n2973_), .ZN(new_n2978_));
  NOR2_X1    g01976(.A1(new_n2978_), .A2(new_n2591_), .ZN(new_n2979_));
  NOR2_X1    g01977(.A1(new_n2976_), .A2(new_n2979_), .ZN(new_n2980_));
  AOI21_X1   g01978(.A1(new_n2555_), .A2(new_n2557_), .B(new_n2556_), .ZN(new_n2981_));
  AOI21_X1   g01979(.A1(new_n2545_), .A2(new_n2547_), .B(new_n2546_), .ZN(new_n2982_));
  XNOR2_X1   g01980(.A1(new_n2981_), .A2(new_n2982_), .ZN(new_n2983_));
  NAND2_X1   g01981(.A1(new_n2983_), .A2(new_n2560_), .ZN(new_n2984_));
  XOR2_X1    g01982(.A1(new_n2981_), .A2(new_n2982_), .Z(new_n2985_));
  NAND2_X1   g01983(.A1(new_n2985_), .A2(new_n2606_), .ZN(new_n2986_));
  NAND2_X1   g01984(.A1(new_n2984_), .A2(new_n2986_), .ZN(new_n2987_));
  NAND3_X1   g01985(.A1(new_n2608_), .A2(new_n2591_), .A3(new_n2602_), .ZN(new_n2988_));
  NAND2_X1   g01986(.A1(new_n2987_), .A2(new_n2988_), .ZN(new_n2989_));
  NOR4_X1    g01987(.A1(new_n2603_), .A2(new_n2606_), .A3(new_n2607_), .A4(new_n2983_), .ZN(new_n2990_));
  INV_X1     g01988(.I(new_n2990_), .ZN(new_n2991_));
  NAND3_X1   g01989(.A1(new_n2989_), .A2(new_n2991_), .A3(new_n2980_), .ZN(new_n2992_));
  NAND2_X1   g01990(.A1(new_n2978_), .A2(new_n2591_), .ZN(new_n2993_));
  NAND2_X1   g01991(.A1(new_n2969_), .A2(new_n2975_), .ZN(new_n2994_));
  NAND2_X1   g01992(.A1(new_n2994_), .A2(new_n2993_), .ZN(new_n2995_));
  NOR2_X1    g01993(.A1(new_n2985_), .A2(new_n2606_), .ZN(new_n2996_));
  NOR2_X1    g01994(.A1(new_n2983_), .A2(new_n2560_), .ZN(new_n2997_));
  NOR2_X1    g01995(.A1(new_n2997_), .A2(new_n2996_), .ZN(new_n2998_));
  NOR2_X1    g01996(.A1(new_n2570_), .A2(new_n2603_), .ZN(new_n2999_));
  NOR2_X1    g01997(.A1(new_n2998_), .A2(new_n2999_), .ZN(new_n3000_));
  OAI21_X1   g01998(.A1(new_n3000_), .A2(new_n2990_), .B(new_n2995_), .ZN(new_n3001_));
  NAND2_X1   g01999(.A1(new_n2992_), .A2(new_n3001_), .ZN(new_n3002_));
  NAND2_X1   g02000(.A1(new_n2679_), .A2(new_n2682_), .ZN(new_n3003_));
  NAND2_X1   g02001(.A1(new_n2675_), .A2(new_n2642_), .ZN(new_n3004_));
  AOI22_X1   g02002(.A1(new_n2686_), .A2(new_n2685_), .B1(new_n3003_), .B2(new_n3004_), .ZN(new_n3005_));
  AOI21_X1   g02003(.A1(\A[83] ), .A2(\A[84] ), .B(\A[82] ), .ZN(new_n3006_));
  AOI21_X1   g02004(.A1(\A[80] ), .A2(\A[81] ), .B(\A[79] ), .ZN(new_n3007_));
  OAI22_X1   g02005(.A1(new_n2650_), .A2(new_n3007_), .B1(new_n3006_), .B2(new_n2660_), .ZN(new_n3008_));
  NOR4_X1    g02006(.A1(new_n3006_), .A2(new_n3007_), .A3(new_n2650_), .A4(new_n2660_), .ZN(new_n3009_));
  INV_X1     g02007(.I(new_n3009_), .ZN(new_n3010_));
  NAND2_X1   g02008(.A1(new_n3010_), .A2(new_n3008_), .ZN(new_n3011_));
  NOR2_X1    g02009(.A1(new_n2663_), .A2(new_n3011_), .ZN(new_n3012_));
  NOR2_X1    g02010(.A1(new_n3006_), .A2(new_n2660_), .ZN(new_n3013_));
  NOR2_X1    g02011(.A1(new_n3007_), .A2(new_n2650_), .ZN(new_n3014_));
  NOR2_X1    g02012(.A1(new_n3013_), .A2(new_n3014_), .ZN(new_n3015_));
  NOR2_X1    g02013(.A1(new_n3015_), .A2(new_n3009_), .ZN(new_n3016_));
  NOR2_X1    g02014(.A1(new_n2680_), .A2(new_n3016_), .ZN(new_n3017_));
  NOR2_X1    g02015(.A1(new_n3012_), .A2(new_n3017_), .ZN(new_n3018_));
  AOI21_X1   g02016(.A1(\A[89] ), .A2(\A[90] ), .B(\A[88] ), .ZN(new_n3019_));
  AOI21_X1   g02017(.A1(\A[86] ), .A2(\A[87] ), .B(\A[85] ), .ZN(new_n3020_));
  NOR2_X1    g02018(.A1(new_n3020_), .A2(new_n2616_), .ZN(new_n3021_));
  NOR3_X1    g02019(.A1(new_n3021_), .A2(new_n2626_), .A3(new_n3019_), .ZN(new_n3022_));
  NOR2_X1    g02020(.A1(new_n3019_), .A2(new_n2626_), .ZN(new_n3023_));
  NOR3_X1    g02021(.A1(new_n3023_), .A2(new_n2616_), .A3(new_n3020_), .ZN(new_n3024_));
  NOR2_X1    g02022(.A1(new_n3022_), .A2(new_n3024_), .ZN(new_n3025_));
  NAND2_X1   g02023(.A1(new_n2630_), .A2(new_n3025_), .ZN(new_n3026_));
  XOR2_X1    g02024(.A1(new_n3023_), .A2(new_n3021_), .Z(new_n3027_));
  NAND2_X1   g02025(.A1(new_n3027_), .A2(new_n2677_), .ZN(new_n3028_));
  NAND2_X1   g02026(.A1(new_n3028_), .A2(new_n3026_), .ZN(new_n3029_));
  NAND2_X1   g02027(.A1(new_n2679_), .A2(new_n2675_), .ZN(new_n3030_));
  AOI21_X1   g02028(.A1(new_n3030_), .A2(new_n3029_), .B(new_n3018_), .ZN(new_n3031_));
  NAND4_X1   g02029(.A1(new_n2675_), .A2(new_n2630_), .A3(new_n2641_), .A4(new_n3027_), .ZN(new_n3032_));
  NAND2_X1   g02030(.A1(new_n3031_), .A2(new_n3032_), .ZN(new_n3033_));
  NOR2_X1    g02031(.A1(new_n3027_), .A2(new_n2677_), .ZN(new_n3034_));
  NOR2_X1    g02032(.A1(new_n2630_), .A2(new_n3025_), .ZN(new_n3035_));
  NOR2_X1    g02033(.A1(new_n3034_), .A2(new_n3035_), .ZN(new_n3036_));
  NOR2_X1    g02034(.A1(new_n2642_), .A2(new_n2682_), .ZN(new_n3037_));
  NOR2_X1    g02035(.A1(new_n3036_), .A2(new_n3037_), .ZN(new_n3038_));
  INV_X1     g02036(.I(new_n3032_), .ZN(new_n3039_));
  OAI21_X1   g02037(.A1(new_n3038_), .A2(new_n3039_), .B(new_n3018_), .ZN(new_n3040_));
  NAND3_X1   g02038(.A1(new_n3033_), .A2(new_n3040_), .A3(new_n3005_), .ZN(new_n3041_));
  NAND2_X1   g02039(.A1(new_n2680_), .A2(new_n3016_), .ZN(new_n3042_));
  NAND2_X1   g02040(.A1(new_n2663_), .A2(new_n3011_), .ZN(new_n3043_));
  NAND2_X1   g02041(.A1(new_n3043_), .A2(new_n3042_), .ZN(new_n3044_));
  OAI21_X1   g02042(.A1(new_n3036_), .A2(new_n3037_), .B(new_n3044_), .ZN(new_n3045_));
  NOR2_X1    g02043(.A1(new_n3045_), .A2(new_n3039_), .ZN(new_n3046_));
  NAND2_X1   g02044(.A1(new_n3030_), .A2(new_n3029_), .ZN(new_n3047_));
  AOI21_X1   g02045(.A1(new_n3047_), .A2(new_n3032_), .B(new_n3044_), .ZN(new_n3048_));
  OAI21_X1   g02046(.A1(new_n3046_), .A2(new_n3048_), .B(new_n2684_), .ZN(new_n3049_));
  NAND3_X1   g02047(.A1(new_n3049_), .A2(new_n3041_), .A3(new_n3002_), .ZN(new_n3050_));
  NOR3_X1    g02048(.A1(new_n3000_), .A2(new_n2995_), .A3(new_n2990_), .ZN(new_n3051_));
  AOI21_X1   g02049(.A1(new_n2989_), .A2(new_n2991_), .B(new_n2980_), .ZN(new_n3052_));
  NOR2_X1    g02050(.A1(new_n3052_), .A2(new_n3051_), .ZN(new_n3053_));
  NOR3_X1    g02051(.A1(new_n3046_), .A2(new_n3048_), .A3(new_n2684_), .ZN(new_n3054_));
  AOI21_X1   g02052(.A1(new_n3033_), .A2(new_n3040_), .B(new_n3005_), .ZN(new_n3055_));
  OAI21_X1   g02053(.A1(new_n3055_), .A2(new_n3054_), .B(new_n3053_), .ZN(new_n3056_));
  NAND3_X1   g02054(.A1(new_n3056_), .A2(new_n3050_), .A3(new_n2690_), .ZN(new_n3057_));
  INV_X1     g02055(.I(new_n2690_), .ZN(new_n3058_));
  NOR3_X1    g02056(.A1(new_n3054_), .A2(new_n3055_), .A3(new_n3053_), .ZN(new_n3059_));
  AOI21_X1   g02057(.A1(new_n3041_), .A2(new_n3049_), .B(new_n3002_), .ZN(new_n3060_));
  OAI21_X1   g02058(.A1(new_n3059_), .A2(new_n3060_), .B(new_n3058_), .ZN(new_n3061_));
  NAND3_X1   g02059(.A1(new_n3061_), .A2(new_n3057_), .A3(new_n2968_), .ZN(new_n3062_));
  INV_X1     g02060(.I(new_n2968_), .ZN(new_n3063_));
  NOR3_X1    g02061(.A1(new_n3058_), .A2(new_n3059_), .A3(new_n3060_), .ZN(new_n3064_));
  AOI21_X1   g02062(.A1(new_n3056_), .A2(new_n3050_), .B(new_n2690_), .ZN(new_n3065_));
  OAI21_X1   g02063(.A1(new_n3064_), .A2(new_n3065_), .B(new_n3063_), .ZN(new_n3066_));
  NAND3_X1   g02064(.A1(new_n3066_), .A2(new_n2882_), .A3(new_n3062_), .ZN(new_n3067_));
  NOR3_X1    g02065(.A1(new_n3063_), .A2(new_n3064_), .A3(new_n3065_), .ZN(new_n3068_));
  AOI21_X1   g02066(.A1(new_n3061_), .A2(new_n3057_), .B(new_n2968_), .ZN(new_n3069_));
  OAI21_X1   g02067(.A1(new_n3068_), .A2(new_n3069_), .B(new_n2694_), .ZN(new_n3070_));
  NAND3_X1   g02068(.A1(new_n2881_), .A2(new_n3067_), .A3(new_n3070_), .ZN(new_n3071_));
  AOI22_X1   g02069(.A1(new_n2876_), .A2(new_n2782_), .B1(new_n2879_), .B2(new_n2875_), .ZN(new_n3072_));
  NOR3_X1    g02070(.A1(new_n3068_), .A2(new_n3069_), .A3(new_n2694_), .ZN(new_n3073_));
  AOI21_X1   g02071(.A1(new_n3066_), .A2(new_n3062_), .B(new_n2882_), .ZN(new_n3074_));
  OAI21_X1   g02072(.A1(new_n3074_), .A2(new_n3073_), .B(new_n3072_), .ZN(new_n3075_));
  AOI21_X1   g02073(.A1(new_n3071_), .A2(new_n3075_), .B(new_n2698_), .ZN(new_n3076_));
  NOR2_X1    g02074(.A1(new_n2882_), .A2(new_n2695_), .ZN(new_n3077_));
  NAND2_X1   g02075(.A1(new_n3077_), .A2(new_n2067_), .ZN(new_n3078_));
  NOR3_X1    g02076(.A1(new_n3074_), .A2(new_n3073_), .A3(new_n3072_), .ZN(new_n3079_));
  AOI21_X1   g02077(.A1(new_n3067_), .A2(new_n3070_), .B(new_n2881_), .ZN(new_n3080_));
  NOR3_X1    g02078(.A1(new_n3080_), .A2(new_n3079_), .A3(new_n3078_), .ZN(new_n3081_));
  NOR3_X1    g02079(.A1(new_n3081_), .A2(new_n3076_), .A3(new_n2065_), .ZN(new_n3082_));
  INV_X1     g02080(.I(new_n2060_), .ZN(new_n3083_));
  NAND3_X1   g02081(.A1(new_n2054_), .A2(new_n2059_), .A3(new_n1515_), .ZN(new_n3084_));
  NAND2_X1   g02082(.A1(new_n3083_), .A2(new_n3084_), .ZN(new_n3085_));
  OAI21_X1   g02083(.A1(new_n3080_), .A2(new_n3079_), .B(new_n3078_), .ZN(new_n3086_));
  NAND3_X1   g02084(.A1(new_n3071_), .A2(new_n3075_), .A3(new_n2698_), .ZN(new_n3087_));
  AOI21_X1   g02085(.A1(new_n3086_), .A2(new_n3087_), .B(new_n3085_), .ZN(new_n3088_));
  NOR2_X1    g02086(.A1(new_n3088_), .A2(new_n3082_), .ZN(new_n3089_));
  INV_X1     g02087(.I(\A[385] ), .ZN(new_n3090_));
  INV_X1     g02088(.I(\A[386] ), .ZN(new_n3091_));
  NAND2_X1   g02089(.A1(new_n3091_), .A2(\A[387] ), .ZN(new_n3092_));
  INV_X1     g02090(.I(\A[387] ), .ZN(new_n3093_));
  NAND2_X1   g02091(.A1(new_n3093_), .A2(\A[386] ), .ZN(new_n3094_));
  AOI21_X1   g02092(.A1(new_n3092_), .A2(new_n3094_), .B(new_n3090_), .ZN(new_n3095_));
  NOR2_X1    g02093(.A1(\A[386] ), .A2(\A[387] ), .ZN(new_n3096_));
  INV_X1     g02094(.I(new_n3096_), .ZN(new_n3097_));
  NAND2_X1   g02095(.A1(\A[386] ), .A2(\A[387] ), .ZN(new_n3098_));
  AOI21_X1   g02096(.A1(new_n3097_), .A2(new_n3098_), .B(\A[385] ), .ZN(new_n3099_));
  INV_X1     g02097(.I(\A[388] ), .ZN(new_n3100_));
  INV_X1     g02098(.I(\A[389] ), .ZN(new_n3101_));
  NAND2_X1   g02099(.A1(new_n3101_), .A2(\A[390] ), .ZN(new_n3102_));
  INV_X1     g02100(.I(\A[390] ), .ZN(new_n3103_));
  NAND2_X1   g02101(.A1(new_n3103_), .A2(\A[389] ), .ZN(new_n3104_));
  AOI21_X1   g02102(.A1(new_n3102_), .A2(new_n3104_), .B(new_n3100_), .ZN(new_n3105_));
  NOR2_X1    g02103(.A1(\A[389] ), .A2(\A[390] ), .ZN(new_n3106_));
  INV_X1     g02104(.I(new_n3106_), .ZN(new_n3107_));
  NAND2_X1   g02105(.A1(\A[389] ), .A2(\A[390] ), .ZN(new_n3108_));
  AOI21_X1   g02106(.A1(new_n3107_), .A2(new_n3108_), .B(\A[388] ), .ZN(new_n3109_));
  NOR4_X1    g02107(.A1(new_n3095_), .A2(new_n3099_), .A3(new_n3109_), .A4(new_n3105_), .ZN(new_n3110_));
  NOR2_X1    g02108(.A1(new_n3093_), .A2(\A[386] ), .ZN(new_n3111_));
  NOR2_X1    g02109(.A1(new_n3091_), .A2(\A[387] ), .ZN(new_n3112_));
  OAI21_X1   g02110(.A1(new_n3111_), .A2(new_n3112_), .B(\A[385] ), .ZN(new_n3113_));
  INV_X1     g02111(.I(new_n3098_), .ZN(new_n3114_));
  OAI21_X1   g02112(.A1(new_n3114_), .A2(new_n3096_), .B(new_n3090_), .ZN(new_n3115_));
  NOR2_X1    g02113(.A1(new_n3103_), .A2(\A[389] ), .ZN(new_n3116_));
  NOR2_X1    g02114(.A1(new_n3101_), .A2(\A[390] ), .ZN(new_n3117_));
  OAI21_X1   g02115(.A1(new_n3116_), .A2(new_n3117_), .B(\A[388] ), .ZN(new_n3118_));
  AND2_X2    g02116(.A1(\A[389] ), .A2(\A[390] ), .Z(new_n3119_));
  OAI21_X1   g02117(.A1(new_n3119_), .A2(new_n3106_), .B(new_n3100_), .ZN(new_n3120_));
  AOI22_X1   g02118(.A1(new_n3113_), .A2(new_n3115_), .B1(new_n3118_), .B2(new_n3120_), .ZN(new_n3121_));
  NOR2_X1    g02119(.A1(new_n3110_), .A2(new_n3121_), .ZN(new_n3122_));
  INV_X1     g02120(.I(\A[381] ), .ZN(new_n3123_));
  NOR2_X1    g02121(.A1(new_n3123_), .A2(\A[380] ), .ZN(new_n3124_));
  INV_X1     g02122(.I(\A[380] ), .ZN(new_n3125_));
  NOR2_X1    g02123(.A1(new_n3125_), .A2(\A[381] ), .ZN(new_n3126_));
  OAI21_X1   g02124(.A1(new_n3124_), .A2(new_n3126_), .B(\A[379] ), .ZN(new_n3127_));
  INV_X1     g02125(.I(\A[379] ), .ZN(new_n3128_));
  NAND2_X1   g02126(.A1(\A[380] ), .A2(\A[381] ), .ZN(new_n3129_));
  INV_X1     g02127(.I(new_n3129_), .ZN(new_n3130_));
  NOR2_X1    g02128(.A1(\A[380] ), .A2(\A[381] ), .ZN(new_n3131_));
  OAI21_X1   g02129(.A1(new_n3130_), .A2(new_n3131_), .B(new_n3128_), .ZN(new_n3132_));
  INV_X1     g02130(.I(\A[384] ), .ZN(new_n3133_));
  NOR2_X1    g02131(.A1(new_n3133_), .A2(\A[383] ), .ZN(new_n3134_));
  INV_X1     g02132(.I(\A[383] ), .ZN(new_n3135_));
  NOR2_X1    g02133(.A1(new_n3135_), .A2(\A[384] ), .ZN(new_n3136_));
  OAI21_X1   g02134(.A1(new_n3134_), .A2(new_n3136_), .B(\A[382] ), .ZN(new_n3137_));
  INV_X1     g02135(.I(\A[382] ), .ZN(new_n3138_));
  AND2_X2    g02136(.A1(\A[383] ), .A2(\A[384] ), .Z(new_n3139_));
  NOR2_X1    g02137(.A1(\A[383] ), .A2(\A[384] ), .ZN(new_n3140_));
  OAI21_X1   g02138(.A1(new_n3139_), .A2(new_n3140_), .B(new_n3138_), .ZN(new_n3141_));
  NAND4_X1   g02139(.A1(new_n3127_), .A2(new_n3137_), .A3(new_n3132_), .A4(new_n3141_), .ZN(new_n3142_));
  NAND2_X1   g02140(.A1(new_n3127_), .A2(new_n3132_), .ZN(new_n3143_));
  NAND2_X1   g02141(.A1(new_n3137_), .A2(new_n3141_), .ZN(new_n3144_));
  NAND2_X1   g02142(.A1(new_n3143_), .A2(new_n3144_), .ZN(new_n3145_));
  NAND2_X1   g02143(.A1(new_n3145_), .A2(new_n3142_), .ZN(new_n3146_));
  NAND2_X1   g02144(.A1(new_n3146_), .A2(new_n3122_), .ZN(new_n3147_));
  NAND4_X1   g02145(.A1(new_n3113_), .A2(new_n3118_), .A3(new_n3115_), .A4(new_n3120_), .ZN(new_n3148_));
  OAI22_X1   g02146(.A1(new_n3095_), .A2(new_n3099_), .B1(new_n3109_), .B2(new_n3105_), .ZN(new_n3149_));
  NAND2_X1   g02147(.A1(new_n3149_), .A2(new_n3148_), .ZN(new_n3150_));
  NAND2_X1   g02148(.A1(new_n3125_), .A2(\A[381] ), .ZN(new_n3151_));
  NAND2_X1   g02149(.A1(new_n3123_), .A2(\A[380] ), .ZN(new_n3152_));
  AOI21_X1   g02150(.A1(new_n3151_), .A2(new_n3152_), .B(new_n3128_), .ZN(new_n3153_));
  INV_X1     g02151(.I(new_n3131_), .ZN(new_n3154_));
  AOI21_X1   g02152(.A1(new_n3154_), .A2(new_n3129_), .B(\A[379] ), .ZN(new_n3155_));
  NAND2_X1   g02153(.A1(new_n3135_), .A2(\A[384] ), .ZN(new_n3156_));
  NAND2_X1   g02154(.A1(new_n3133_), .A2(\A[383] ), .ZN(new_n3157_));
  AOI21_X1   g02155(.A1(new_n3156_), .A2(new_n3157_), .B(new_n3138_), .ZN(new_n3158_));
  NAND2_X1   g02156(.A1(\A[383] ), .A2(\A[384] ), .ZN(new_n3159_));
  OR2_X2     g02157(.A1(\A[383] ), .A2(\A[384] ), .Z(new_n3160_));
  AOI21_X1   g02158(.A1(new_n3160_), .A2(new_n3159_), .B(\A[382] ), .ZN(new_n3161_));
  NOR4_X1    g02159(.A1(new_n3153_), .A2(new_n3155_), .A3(new_n3158_), .A4(new_n3161_), .ZN(new_n3162_));
  NOR2_X1    g02160(.A1(new_n3155_), .A2(new_n3153_), .ZN(new_n3163_));
  NOR2_X1    g02161(.A1(new_n3158_), .A2(new_n3161_), .ZN(new_n3164_));
  NOR2_X1    g02162(.A1(new_n3163_), .A2(new_n3164_), .ZN(new_n3165_));
  NOR2_X1    g02163(.A1(new_n3165_), .A2(new_n3162_), .ZN(new_n3166_));
  NAND2_X1   g02164(.A1(new_n3166_), .A2(new_n3150_), .ZN(new_n3167_));
  INV_X1     g02165(.I(\A[373] ), .ZN(new_n3168_));
  INV_X1     g02166(.I(\A[374] ), .ZN(new_n3169_));
  NAND2_X1   g02167(.A1(new_n3169_), .A2(\A[375] ), .ZN(new_n3170_));
  INV_X1     g02168(.I(\A[375] ), .ZN(new_n3171_));
  NAND2_X1   g02169(.A1(new_n3171_), .A2(\A[374] ), .ZN(new_n3172_));
  AOI21_X1   g02170(.A1(new_n3170_), .A2(new_n3172_), .B(new_n3168_), .ZN(new_n3173_));
  NOR2_X1    g02171(.A1(\A[374] ), .A2(\A[375] ), .ZN(new_n3174_));
  INV_X1     g02172(.I(new_n3174_), .ZN(new_n3175_));
  NAND2_X1   g02173(.A1(\A[374] ), .A2(\A[375] ), .ZN(new_n3176_));
  AOI21_X1   g02174(.A1(new_n3175_), .A2(new_n3176_), .B(\A[373] ), .ZN(new_n3177_));
  INV_X1     g02175(.I(\A[376] ), .ZN(new_n3178_));
  INV_X1     g02176(.I(\A[377] ), .ZN(new_n3179_));
  NAND2_X1   g02177(.A1(new_n3179_), .A2(\A[378] ), .ZN(new_n3180_));
  INV_X1     g02178(.I(\A[378] ), .ZN(new_n3181_));
  NAND2_X1   g02179(.A1(new_n3181_), .A2(\A[377] ), .ZN(new_n3182_));
  AOI21_X1   g02180(.A1(new_n3180_), .A2(new_n3182_), .B(new_n3178_), .ZN(new_n3183_));
  NOR2_X1    g02181(.A1(\A[377] ), .A2(\A[378] ), .ZN(new_n3184_));
  INV_X1     g02182(.I(new_n3184_), .ZN(new_n3185_));
  NAND2_X1   g02183(.A1(\A[377] ), .A2(\A[378] ), .ZN(new_n3186_));
  AOI21_X1   g02184(.A1(new_n3185_), .A2(new_n3186_), .B(\A[376] ), .ZN(new_n3187_));
  NOR4_X1    g02185(.A1(new_n3173_), .A2(new_n3177_), .A3(new_n3187_), .A4(new_n3183_), .ZN(new_n3188_));
  NOR2_X1    g02186(.A1(new_n3171_), .A2(\A[374] ), .ZN(new_n3189_));
  NOR2_X1    g02187(.A1(new_n3169_), .A2(\A[375] ), .ZN(new_n3190_));
  OAI21_X1   g02188(.A1(new_n3189_), .A2(new_n3190_), .B(\A[373] ), .ZN(new_n3191_));
  INV_X1     g02189(.I(new_n3176_), .ZN(new_n3192_));
  OAI21_X1   g02190(.A1(new_n3192_), .A2(new_n3174_), .B(new_n3168_), .ZN(new_n3193_));
  NOR2_X1    g02191(.A1(new_n3181_), .A2(\A[377] ), .ZN(new_n3194_));
  NOR2_X1    g02192(.A1(new_n3179_), .A2(\A[378] ), .ZN(new_n3195_));
  OAI21_X1   g02193(.A1(new_n3194_), .A2(new_n3195_), .B(\A[376] ), .ZN(new_n3196_));
  AND2_X2    g02194(.A1(\A[377] ), .A2(\A[378] ), .Z(new_n3197_));
  OAI21_X1   g02195(.A1(new_n3197_), .A2(new_n3184_), .B(new_n3178_), .ZN(new_n3198_));
  AOI22_X1   g02196(.A1(new_n3191_), .A2(new_n3193_), .B1(new_n3196_), .B2(new_n3198_), .ZN(new_n3199_));
  NOR2_X1    g02197(.A1(new_n3188_), .A2(new_n3199_), .ZN(new_n3200_));
  INV_X1     g02198(.I(\A[369] ), .ZN(new_n3201_));
  NOR2_X1    g02199(.A1(new_n3201_), .A2(\A[368] ), .ZN(new_n3202_));
  INV_X1     g02200(.I(\A[368] ), .ZN(new_n3203_));
  NOR2_X1    g02201(.A1(new_n3203_), .A2(\A[369] ), .ZN(new_n3204_));
  OAI21_X1   g02202(.A1(new_n3202_), .A2(new_n3204_), .B(\A[367] ), .ZN(new_n3205_));
  INV_X1     g02203(.I(\A[367] ), .ZN(new_n3206_));
  NAND2_X1   g02204(.A1(\A[368] ), .A2(\A[369] ), .ZN(new_n3207_));
  INV_X1     g02205(.I(new_n3207_), .ZN(new_n3208_));
  NOR2_X1    g02206(.A1(\A[368] ), .A2(\A[369] ), .ZN(new_n3209_));
  OAI21_X1   g02207(.A1(new_n3208_), .A2(new_n3209_), .B(new_n3206_), .ZN(new_n3210_));
  INV_X1     g02208(.I(\A[372] ), .ZN(new_n3211_));
  NOR2_X1    g02209(.A1(new_n3211_), .A2(\A[371] ), .ZN(new_n3212_));
  INV_X1     g02210(.I(\A[371] ), .ZN(new_n3213_));
  NOR2_X1    g02211(.A1(new_n3213_), .A2(\A[372] ), .ZN(new_n3214_));
  OAI21_X1   g02212(.A1(new_n3212_), .A2(new_n3214_), .B(\A[370] ), .ZN(new_n3215_));
  INV_X1     g02213(.I(\A[370] ), .ZN(new_n3216_));
  NAND2_X1   g02214(.A1(\A[371] ), .A2(\A[372] ), .ZN(new_n3217_));
  INV_X1     g02215(.I(new_n3217_), .ZN(new_n3218_));
  NOR2_X1    g02216(.A1(\A[371] ), .A2(\A[372] ), .ZN(new_n3219_));
  OAI21_X1   g02217(.A1(new_n3218_), .A2(new_n3219_), .B(new_n3216_), .ZN(new_n3220_));
  NAND4_X1   g02218(.A1(new_n3205_), .A2(new_n3210_), .A3(new_n3215_), .A4(new_n3220_), .ZN(new_n3221_));
  NAND2_X1   g02219(.A1(new_n3203_), .A2(\A[369] ), .ZN(new_n3222_));
  NAND2_X1   g02220(.A1(new_n3201_), .A2(\A[368] ), .ZN(new_n3223_));
  AOI21_X1   g02221(.A1(new_n3222_), .A2(new_n3223_), .B(new_n3206_), .ZN(new_n3224_));
  INV_X1     g02222(.I(new_n3209_), .ZN(new_n3225_));
  AOI21_X1   g02223(.A1(new_n3225_), .A2(new_n3207_), .B(\A[367] ), .ZN(new_n3226_));
  NAND2_X1   g02224(.A1(new_n3213_), .A2(\A[372] ), .ZN(new_n3227_));
  NAND2_X1   g02225(.A1(new_n3211_), .A2(\A[371] ), .ZN(new_n3228_));
  AOI21_X1   g02226(.A1(new_n3227_), .A2(new_n3228_), .B(new_n3216_), .ZN(new_n3229_));
  OR2_X2     g02227(.A1(\A[371] ), .A2(\A[372] ), .Z(new_n3230_));
  AOI21_X1   g02228(.A1(new_n3230_), .A2(new_n3217_), .B(\A[370] ), .ZN(new_n3231_));
  OAI22_X1   g02229(.A1(new_n3224_), .A2(new_n3226_), .B1(new_n3229_), .B2(new_n3231_), .ZN(new_n3232_));
  NAND2_X1   g02230(.A1(new_n3221_), .A2(new_n3232_), .ZN(new_n3233_));
  NAND2_X1   g02231(.A1(new_n3200_), .A2(new_n3233_), .ZN(new_n3234_));
  NAND4_X1   g02232(.A1(new_n3191_), .A2(new_n3196_), .A3(new_n3193_), .A4(new_n3198_), .ZN(new_n3235_));
  OAI22_X1   g02233(.A1(new_n3173_), .A2(new_n3177_), .B1(new_n3187_), .B2(new_n3183_), .ZN(new_n3236_));
  NAND2_X1   g02234(.A1(new_n3236_), .A2(new_n3235_), .ZN(new_n3237_));
  NOR4_X1    g02235(.A1(new_n3224_), .A2(new_n3226_), .A3(new_n3229_), .A4(new_n3231_), .ZN(new_n3238_));
  AOI22_X1   g02236(.A1(new_n3205_), .A2(new_n3210_), .B1(new_n3215_), .B2(new_n3220_), .ZN(new_n3239_));
  NOR2_X1    g02237(.A1(new_n3239_), .A2(new_n3238_), .ZN(new_n3240_));
  NAND2_X1   g02238(.A1(new_n3240_), .A2(new_n3237_), .ZN(new_n3241_));
  AOI22_X1   g02239(.A1(new_n3167_), .A2(new_n3147_), .B1(new_n3234_), .B2(new_n3241_), .ZN(new_n3242_));
  NOR2_X1    g02240(.A1(new_n3166_), .A2(new_n3150_), .ZN(new_n3243_));
  NOR2_X1    g02241(.A1(new_n3146_), .A2(new_n3122_), .ZN(new_n3244_));
  NOR2_X1    g02242(.A1(new_n3240_), .A2(new_n3237_), .ZN(new_n3245_));
  NOR2_X1    g02243(.A1(new_n3200_), .A2(new_n3233_), .ZN(new_n3246_));
  NOR4_X1    g02244(.A1(new_n3243_), .A2(new_n3244_), .A3(new_n3246_), .A4(new_n3245_), .ZN(new_n3247_));
  NOR2_X1    g02245(.A1(new_n3247_), .A2(new_n3242_), .ZN(new_n3248_));
  INV_X1     g02246(.I(new_n3248_), .ZN(new_n3249_));
  INV_X1     g02247(.I(\A[391] ), .ZN(new_n3250_));
  INV_X1     g02248(.I(\A[393] ), .ZN(new_n3251_));
  NOR2_X1    g02249(.A1(new_n3251_), .A2(\A[392] ), .ZN(new_n3252_));
  INV_X1     g02250(.I(new_n3252_), .ZN(new_n3253_));
  NAND2_X1   g02251(.A1(new_n3251_), .A2(\A[392] ), .ZN(new_n3254_));
  AOI21_X1   g02252(.A1(new_n3253_), .A2(new_n3254_), .B(new_n3250_), .ZN(new_n3255_));
  NAND2_X1   g02253(.A1(\A[392] ), .A2(\A[393] ), .ZN(new_n3256_));
  NOR2_X1    g02254(.A1(\A[392] ), .A2(\A[393] ), .ZN(new_n3257_));
  INV_X1     g02255(.I(new_n3257_), .ZN(new_n3258_));
  AOI21_X1   g02256(.A1(new_n3258_), .A2(new_n3256_), .B(\A[391] ), .ZN(new_n3259_));
  INV_X1     g02257(.I(\A[394] ), .ZN(new_n3260_));
  INV_X1     g02258(.I(\A[395] ), .ZN(new_n3261_));
  NAND2_X1   g02259(.A1(new_n3261_), .A2(\A[396] ), .ZN(new_n3262_));
  INV_X1     g02260(.I(\A[396] ), .ZN(new_n3263_));
  NAND2_X1   g02261(.A1(new_n3263_), .A2(\A[395] ), .ZN(new_n3264_));
  AOI21_X1   g02262(.A1(new_n3262_), .A2(new_n3264_), .B(new_n3260_), .ZN(new_n3265_));
  NAND2_X1   g02263(.A1(\A[395] ), .A2(\A[396] ), .ZN(new_n3266_));
  NOR2_X1    g02264(.A1(\A[395] ), .A2(\A[396] ), .ZN(new_n3267_));
  INV_X1     g02265(.I(new_n3267_), .ZN(new_n3268_));
  AOI21_X1   g02266(.A1(new_n3268_), .A2(new_n3266_), .B(\A[394] ), .ZN(new_n3269_));
  NOR4_X1    g02267(.A1(new_n3255_), .A2(new_n3259_), .A3(new_n3269_), .A4(new_n3265_), .ZN(new_n3270_));
  INV_X1     g02268(.I(\A[392] ), .ZN(new_n3271_));
  NOR2_X1    g02269(.A1(new_n3271_), .A2(\A[393] ), .ZN(new_n3272_));
  OAI21_X1   g02270(.A1(new_n3252_), .A2(new_n3272_), .B(\A[391] ), .ZN(new_n3273_));
  INV_X1     g02271(.I(new_n3256_), .ZN(new_n3274_));
  OAI21_X1   g02272(.A1(new_n3274_), .A2(new_n3257_), .B(new_n3250_), .ZN(new_n3275_));
  NOR2_X1    g02273(.A1(new_n3263_), .A2(\A[395] ), .ZN(new_n3276_));
  NOR2_X1    g02274(.A1(new_n3261_), .A2(\A[396] ), .ZN(new_n3277_));
  OAI21_X1   g02275(.A1(new_n3276_), .A2(new_n3277_), .B(\A[394] ), .ZN(new_n3278_));
  INV_X1     g02276(.I(new_n3266_), .ZN(new_n3279_));
  OAI21_X1   g02277(.A1(new_n3279_), .A2(new_n3267_), .B(new_n3260_), .ZN(new_n3280_));
  AOI22_X1   g02278(.A1(new_n3273_), .A2(new_n3275_), .B1(new_n3278_), .B2(new_n3280_), .ZN(new_n3281_));
  NOR2_X1    g02279(.A1(new_n3270_), .A2(new_n3281_), .ZN(new_n3282_));
  INV_X1     g02280(.I(\A[398] ), .ZN(new_n3283_));
  NAND2_X1   g02281(.A1(new_n3283_), .A2(\A[399] ), .ZN(new_n3284_));
  INV_X1     g02282(.I(new_n3284_), .ZN(new_n3285_));
  NOR2_X1    g02283(.A1(new_n3283_), .A2(\A[399] ), .ZN(new_n3286_));
  OAI21_X1   g02284(.A1(new_n3285_), .A2(new_n3286_), .B(\A[397] ), .ZN(new_n3287_));
  INV_X1     g02285(.I(\A[397] ), .ZN(new_n3288_));
  NAND2_X1   g02286(.A1(\A[398] ), .A2(\A[399] ), .ZN(new_n3289_));
  INV_X1     g02287(.I(new_n3289_), .ZN(new_n3290_));
  NOR2_X1    g02288(.A1(\A[398] ), .A2(\A[399] ), .ZN(new_n3291_));
  OAI21_X1   g02289(.A1(new_n3290_), .A2(new_n3291_), .B(new_n3288_), .ZN(new_n3292_));
  INV_X1     g02290(.I(\A[402] ), .ZN(new_n3293_));
  NOR2_X1    g02291(.A1(new_n3293_), .A2(\A[401] ), .ZN(new_n3294_));
  INV_X1     g02292(.I(\A[401] ), .ZN(new_n3295_));
  NOR2_X1    g02293(.A1(new_n3295_), .A2(\A[402] ), .ZN(new_n3296_));
  OAI21_X1   g02294(.A1(new_n3294_), .A2(new_n3296_), .B(\A[400] ), .ZN(new_n3297_));
  INV_X1     g02295(.I(\A[400] ), .ZN(new_n3298_));
  NAND2_X1   g02296(.A1(\A[401] ), .A2(\A[402] ), .ZN(new_n3299_));
  INV_X1     g02297(.I(new_n3299_), .ZN(new_n3300_));
  NOR2_X1    g02298(.A1(\A[401] ), .A2(\A[402] ), .ZN(new_n3301_));
  OAI21_X1   g02299(.A1(new_n3300_), .A2(new_n3301_), .B(new_n3298_), .ZN(new_n3302_));
  NAND4_X1   g02300(.A1(new_n3287_), .A2(new_n3292_), .A3(new_n3302_), .A4(new_n3297_), .ZN(new_n3303_));
  INV_X1     g02301(.I(\A[399] ), .ZN(new_n3304_));
  NAND2_X1   g02302(.A1(new_n3304_), .A2(\A[398] ), .ZN(new_n3305_));
  AOI21_X1   g02303(.A1(new_n3284_), .A2(new_n3305_), .B(new_n3288_), .ZN(new_n3306_));
  INV_X1     g02304(.I(new_n3291_), .ZN(new_n3307_));
  AOI21_X1   g02305(.A1(new_n3307_), .A2(new_n3289_), .B(\A[397] ), .ZN(new_n3308_));
  NAND2_X1   g02306(.A1(new_n3295_), .A2(\A[402] ), .ZN(new_n3309_));
  NAND2_X1   g02307(.A1(new_n3293_), .A2(\A[401] ), .ZN(new_n3310_));
  AOI21_X1   g02308(.A1(new_n3309_), .A2(new_n3310_), .B(new_n3298_), .ZN(new_n3311_));
  INV_X1     g02309(.I(new_n3301_), .ZN(new_n3312_));
  AOI21_X1   g02310(.A1(new_n3312_), .A2(new_n3299_), .B(\A[400] ), .ZN(new_n3313_));
  OAI22_X1   g02311(.A1(new_n3306_), .A2(new_n3308_), .B1(new_n3313_), .B2(new_n3311_), .ZN(new_n3314_));
  NAND2_X1   g02312(.A1(new_n3303_), .A2(new_n3314_), .ZN(new_n3315_));
  NAND2_X1   g02313(.A1(new_n3282_), .A2(new_n3315_), .ZN(new_n3316_));
  NAND4_X1   g02314(.A1(new_n3273_), .A2(new_n3275_), .A3(new_n3278_), .A4(new_n3280_), .ZN(new_n3317_));
  OAI22_X1   g02315(.A1(new_n3255_), .A2(new_n3259_), .B1(new_n3269_), .B2(new_n3265_), .ZN(new_n3318_));
  NAND2_X1   g02316(.A1(new_n3318_), .A2(new_n3317_), .ZN(new_n3319_));
  NOR4_X1    g02317(.A1(new_n3306_), .A2(new_n3308_), .A3(new_n3313_), .A4(new_n3311_), .ZN(new_n3320_));
  AOI22_X1   g02318(.A1(new_n3287_), .A2(new_n3292_), .B1(new_n3302_), .B2(new_n3297_), .ZN(new_n3321_));
  NOR2_X1    g02319(.A1(new_n3321_), .A2(new_n3320_), .ZN(new_n3322_));
  NAND2_X1   g02320(.A1(new_n3322_), .A2(new_n3319_), .ZN(new_n3323_));
  NAND2_X1   g02321(.A1(new_n3323_), .A2(new_n3316_), .ZN(new_n3324_));
  INV_X1     g02322(.I(\A[403] ), .ZN(new_n3325_));
  INV_X1     g02323(.I(\A[404] ), .ZN(new_n3326_));
  NAND2_X1   g02324(.A1(new_n3326_), .A2(\A[405] ), .ZN(new_n3327_));
  INV_X1     g02325(.I(\A[405] ), .ZN(new_n3328_));
  NAND2_X1   g02326(.A1(new_n3328_), .A2(\A[404] ), .ZN(new_n3329_));
  AOI21_X1   g02327(.A1(new_n3327_), .A2(new_n3329_), .B(new_n3325_), .ZN(new_n3330_));
  NAND2_X1   g02328(.A1(\A[404] ), .A2(\A[405] ), .ZN(new_n3331_));
  NOR2_X1    g02329(.A1(\A[404] ), .A2(\A[405] ), .ZN(new_n3332_));
  INV_X1     g02330(.I(new_n3332_), .ZN(new_n3333_));
  AOI21_X1   g02331(.A1(new_n3333_), .A2(new_n3331_), .B(\A[403] ), .ZN(new_n3334_));
  INV_X1     g02332(.I(\A[406] ), .ZN(new_n3335_));
  INV_X1     g02333(.I(\A[407] ), .ZN(new_n3336_));
  NAND2_X1   g02334(.A1(new_n3336_), .A2(\A[408] ), .ZN(new_n3337_));
  INV_X1     g02335(.I(\A[408] ), .ZN(new_n3338_));
  NAND2_X1   g02336(.A1(new_n3338_), .A2(\A[407] ), .ZN(new_n3339_));
  AOI21_X1   g02337(.A1(new_n3337_), .A2(new_n3339_), .B(new_n3335_), .ZN(new_n3340_));
  NAND2_X1   g02338(.A1(\A[407] ), .A2(\A[408] ), .ZN(new_n3341_));
  OR2_X2     g02339(.A1(\A[407] ), .A2(\A[408] ), .Z(new_n3342_));
  AOI21_X1   g02340(.A1(new_n3342_), .A2(new_n3341_), .B(\A[406] ), .ZN(new_n3343_));
  NOR4_X1    g02341(.A1(new_n3330_), .A2(new_n3334_), .A3(new_n3340_), .A4(new_n3343_), .ZN(new_n3344_));
  NOR2_X1    g02342(.A1(new_n3328_), .A2(\A[404] ), .ZN(new_n3345_));
  NOR2_X1    g02343(.A1(new_n3326_), .A2(\A[405] ), .ZN(new_n3346_));
  OAI21_X1   g02344(.A1(new_n3345_), .A2(new_n3346_), .B(\A[403] ), .ZN(new_n3347_));
  INV_X1     g02345(.I(new_n3331_), .ZN(new_n3348_));
  OAI21_X1   g02346(.A1(new_n3348_), .A2(new_n3332_), .B(new_n3325_), .ZN(new_n3349_));
  NOR2_X1    g02347(.A1(new_n3338_), .A2(\A[407] ), .ZN(new_n3350_));
  NOR2_X1    g02348(.A1(new_n3336_), .A2(\A[408] ), .ZN(new_n3351_));
  OAI21_X1   g02349(.A1(new_n3350_), .A2(new_n3351_), .B(\A[406] ), .ZN(new_n3352_));
  INV_X1     g02350(.I(new_n3341_), .ZN(new_n3353_));
  NOR2_X1    g02351(.A1(\A[407] ), .A2(\A[408] ), .ZN(new_n3354_));
  OAI21_X1   g02352(.A1(new_n3353_), .A2(new_n3354_), .B(new_n3335_), .ZN(new_n3355_));
  AOI22_X1   g02353(.A1(new_n3347_), .A2(new_n3349_), .B1(new_n3352_), .B2(new_n3355_), .ZN(new_n3356_));
  NOR2_X1    g02354(.A1(new_n3356_), .A2(new_n3344_), .ZN(new_n3357_));
  INV_X1     g02355(.I(\A[411] ), .ZN(new_n3358_));
  NOR2_X1    g02356(.A1(new_n3358_), .A2(\A[410] ), .ZN(new_n3359_));
  INV_X1     g02357(.I(\A[410] ), .ZN(new_n3360_));
  NOR2_X1    g02358(.A1(new_n3360_), .A2(\A[411] ), .ZN(new_n3361_));
  OAI21_X1   g02359(.A1(new_n3359_), .A2(new_n3361_), .B(\A[409] ), .ZN(new_n3362_));
  INV_X1     g02360(.I(\A[409] ), .ZN(new_n3363_));
  AND2_X2    g02361(.A1(\A[410] ), .A2(\A[411] ), .Z(new_n3364_));
  NOR2_X1    g02362(.A1(\A[410] ), .A2(\A[411] ), .ZN(new_n3365_));
  OAI21_X1   g02363(.A1(new_n3364_), .A2(new_n3365_), .B(new_n3363_), .ZN(new_n3366_));
  INV_X1     g02364(.I(\A[414] ), .ZN(new_n3367_));
  NOR2_X1    g02365(.A1(new_n3367_), .A2(\A[413] ), .ZN(new_n3368_));
  INV_X1     g02366(.I(\A[413] ), .ZN(new_n3369_));
  NOR2_X1    g02367(.A1(new_n3369_), .A2(\A[414] ), .ZN(new_n3370_));
  OAI21_X1   g02368(.A1(new_n3368_), .A2(new_n3370_), .B(\A[412] ), .ZN(new_n3371_));
  INV_X1     g02369(.I(\A[412] ), .ZN(new_n3372_));
  AND2_X2    g02370(.A1(\A[413] ), .A2(\A[414] ), .Z(new_n3373_));
  NOR2_X1    g02371(.A1(\A[413] ), .A2(\A[414] ), .ZN(new_n3374_));
  OAI21_X1   g02372(.A1(new_n3373_), .A2(new_n3374_), .B(new_n3372_), .ZN(new_n3375_));
  NAND4_X1   g02373(.A1(new_n3362_), .A2(new_n3371_), .A3(new_n3366_), .A4(new_n3375_), .ZN(new_n3376_));
  NAND2_X1   g02374(.A1(new_n3360_), .A2(\A[411] ), .ZN(new_n3377_));
  NAND2_X1   g02375(.A1(new_n3358_), .A2(\A[410] ), .ZN(new_n3378_));
  AOI21_X1   g02376(.A1(new_n3377_), .A2(new_n3378_), .B(new_n3363_), .ZN(new_n3379_));
  NAND2_X1   g02377(.A1(\A[410] ), .A2(\A[411] ), .ZN(new_n3380_));
  INV_X1     g02378(.I(new_n3365_), .ZN(new_n3381_));
  AOI21_X1   g02379(.A1(new_n3381_), .A2(new_n3380_), .B(\A[409] ), .ZN(new_n3382_));
  NAND2_X1   g02380(.A1(new_n3369_), .A2(\A[414] ), .ZN(new_n3383_));
  NAND2_X1   g02381(.A1(new_n3367_), .A2(\A[413] ), .ZN(new_n3384_));
  AOI21_X1   g02382(.A1(new_n3383_), .A2(new_n3384_), .B(new_n3372_), .ZN(new_n3385_));
  NAND2_X1   g02383(.A1(\A[413] ), .A2(\A[414] ), .ZN(new_n3386_));
  OR2_X2     g02384(.A1(\A[413] ), .A2(\A[414] ), .Z(new_n3387_));
  AOI21_X1   g02385(.A1(new_n3387_), .A2(new_n3386_), .B(\A[412] ), .ZN(new_n3388_));
  OAI22_X1   g02386(.A1(new_n3379_), .A2(new_n3382_), .B1(new_n3385_), .B2(new_n3388_), .ZN(new_n3389_));
  NAND2_X1   g02387(.A1(new_n3389_), .A2(new_n3376_), .ZN(new_n3390_));
  XOR2_X1    g02388(.A1(new_n3357_), .A2(new_n3390_), .Z(new_n3391_));
  NOR2_X1    g02389(.A1(new_n3391_), .A2(new_n3324_), .ZN(new_n3392_));
  NOR2_X1    g02390(.A1(new_n3322_), .A2(new_n3319_), .ZN(new_n3393_));
  NOR2_X1    g02391(.A1(new_n3282_), .A2(new_n3315_), .ZN(new_n3394_));
  NOR2_X1    g02392(.A1(new_n3393_), .A2(new_n3394_), .ZN(new_n3395_));
  NAND4_X1   g02393(.A1(new_n3347_), .A2(new_n3349_), .A3(new_n3352_), .A4(new_n3355_), .ZN(new_n3396_));
  OAI22_X1   g02394(.A1(new_n3330_), .A2(new_n3334_), .B1(new_n3340_), .B2(new_n3343_), .ZN(new_n3397_));
  NAND2_X1   g02395(.A1(new_n3396_), .A2(new_n3397_), .ZN(new_n3398_));
  XOR2_X1    g02396(.A1(new_n3398_), .A2(new_n3390_), .Z(new_n3399_));
  NOR2_X1    g02397(.A1(new_n3399_), .A2(new_n3395_), .ZN(new_n3400_));
  NOR2_X1    g02398(.A1(new_n3400_), .A2(new_n3392_), .ZN(new_n3401_));
  NOR2_X1    g02399(.A1(new_n3249_), .A2(new_n3401_), .ZN(new_n3402_));
  NAND2_X1   g02400(.A1(new_n3399_), .A2(new_n3395_), .ZN(new_n3403_));
  NAND2_X1   g02401(.A1(new_n3391_), .A2(new_n3324_), .ZN(new_n3404_));
  NAND2_X1   g02402(.A1(new_n3403_), .A2(new_n3404_), .ZN(new_n3405_));
  NOR2_X1    g02403(.A1(new_n3405_), .A2(new_n3248_), .ZN(new_n3406_));
  NOR2_X1    g02404(.A1(new_n3402_), .A2(new_n3406_), .ZN(new_n3407_));
  INV_X1     g02405(.I(\A[457] ), .ZN(new_n3408_));
  INV_X1     g02406(.I(\A[458] ), .ZN(new_n3409_));
  NAND2_X1   g02407(.A1(new_n3409_), .A2(\A[459] ), .ZN(new_n3410_));
  INV_X1     g02408(.I(\A[459] ), .ZN(new_n3411_));
  NAND2_X1   g02409(.A1(new_n3411_), .A2(\A[458] ), .ZN(new_n3412_));
  AOI21_X1   g02410(.A1(new_n3410_), .A2(new_n3412_), .B(new_n3408_), .ZN(new_n3413_));
  NAND2_X1   g02411(.A1(\A[458] ), .A2(\A[459] ), .ZN(new_n3414_));
  NOR2_X1    g02412(.A1(\A[458] ), .A2(\A[459] ), .ZN(new_n3415_));
  INV_X1     g02413(.I(new_n3415_), .ZN(new_n3416_));
  AOI21_X1   g02414(.A1(new_n3416_), .A2(new_n3414_), .B(\A[457] ), .ZN(new_n3417_));
  NOR2_X1    g02415(.A1(new_n3417_), .A2(new_n3413_), .ZN(new_n3418_));
  INV_X1     g02416(.I(\A[462] ), .ZN(new_n3419_));
  NOR2_X1    g02417(.A1(new_n3419_), .A2(\A[461] ), .ZN(new_n3420_));
  INV_X1     g02418(.I(\A[461] ), .ZN(new_n3421_));
  NOR2_X1    g02419(.A1(new_n3421_), .A2(\A[462] ), .ZN(new_n3422_));
  OAI21_X1   g02420(.A1(new_n3420_), .A2(new_n3422_), .B(\A[460] ), .ZN(new_n3423_));
  INV_X1     g02421(.I(\A[460] ), .ZN(new_n3424_));
  AND2_X2    g02422(.A1(\A[461] ), .A2(\A[462] ), .Z(new_n3425_));
  NOR2_X1    g02423(.A1(\A[461] ), .A2(\A[462] ), .ZN(new_n3426_));
  OAI21_X1   g02424(.A1(new_n3425_), .A2(new_n3426_), .B(new_n3424_), .ZN(new_n3427_));
  NAND2_X1   g02425(.A1(new_n3423_), .A2(new_n3427_), .ZN(new_n3428_));
  NAND2_X1   g02426(.A1(new_n3418_), .A2(new_n3428_), .ZN(new_n3429_));
  NOR2_X1    g02427(.A1(new_n3411_), .A2(\A[458] ), .ZN(new_n3430_));
  NOR2_X1    g02428(.A1(new_n3409_), .A2(\A[459] ), .ZN(new_n3431_));
  OAI21_X1   g02429(.A1(new_n3430_), .A2(new_n3431_), .B(\A[457] ), .ZN(new_n3432_));
  INV_X1     g02430(.I(new_n3414_), .ZN(new_n3433_));
  OAI21_X1   g02431(.A1(new_n3433_), .A2(new_n3415_), .B(new_n3408_), .ZN(new_n3434_));
  NAND2_X1   g02432(.A1(new_n3432_), .A2(new_n3434_), .ZN(new_n3435_));
  NAND2_X1   g02433(.A1(new_n3421_), .A2(\A[462] ), .ZN(new_n3436_));
  NAND2_X1   g02434(.A1(new_n3419_), .A2(\A[461] ), .ZN(new_n3437_));
  AOI21_X1   g02435(.A1(new_n3436_), .A2(new_n3437_), .B(new_n3424_), .ZN(new_n3438_));
  NAND2_X1   g02436(.A1(\A[461] ), .A2(\A[462] ), .ZN(new_n3439_));
  INV_X1     g02437(.I(new_n3426_), .ZN(new_n3440_));
  AOI21_X1   g02438(.A1(new_n3440_), .A2(new_n3439_), .B(\A[460] ), .ZN(new_n3441_));
  NOR2_X1    g02439(.A1(new_n3441_), .A2(new_n3438_), .ZN(new_n3442_));
  NAND2_X1   g02440(.A1(new_n3442_), .A2(new_n3435_), .ZN(new_n3443_));
  NAND2_X1   g02441(.A1(new_n3443_), .A2(new_n3429_), .ZN(new_n3444_));
  INV_X1     g02442(.I(\A[451] ), .ZN(new_n3445_));
  INV_X1     g02443(.I(\A[452] ), .ZN(new_n3446_));
  NAND2_X1   g02444(.A1(new_n3446_), .A2(\A[453] ), .ZN(new_n3447_));
  INV_X1     g02445(.I(\A[453] ), .ZN(new_n3448_));
  NAND2_X1   g02446(.A1(new_n3448_), .A2(\A[452] ), .ZN(new_n3449_));
  AOI21_X1   g02447(.A1(new_n3447_), .A2(new_n3449_), .B(new_n3445_), .ZN(new_n3450_));
  NAND2_X1   g02448(.A1(\A[452] ), .A2(\A[453] ), .ZN(new_n3451_));
  NOR2_X1    g02449(.A1(\A[452] ), .A2(\A[453] ), .ZN(new_n3452_));
  INV_X1     g02450(.I(new_n3452_), .ZN(new_n3453_));
  AOI21_X1   g02451(.A1(new_n3453_), .A2(new_n3451_), .B(\A[451] ), .ZN(new_n3454_));
  NOR2_X1    g02452(.A1(new_n3454_), .A2(new_n3450_), .ZN(new_n3455_));
  INV_X1     g02453(.I(\A[456] ), .ZN(new_n3456_));
  NOR2_X1    g02454(.A1(new_n3456_), .A2(\A[455] ), .ZN(new_n3457_));
  INV_X1     g02455(.I(\A[455] ), .ZN(new_n3458_));
  NOR2_X1    g02456(.A1(new_n3458_), .A2(\A[456] ), .ZN(new_n3459_));
  OAI21_X1   g02457(.A1(new_n3457_), .A2(new_n3459_), .B(\A[454] ), .ZN(new_n3460_));
  INV_X1     g02458(.I(\A[454] ), .ZN(new_n3461_));
  NAND2_X1   g02459(.A1(\A[455] ), .A2(\A[456] ), .ZN(new_n3462_));
  INV_X1     g02460(.I(new_n3462_), .ZN(new_n3463_));
  NOR2_X1    g02461(.A1(\A[455] ), .A2(\A[456] ), .ZN(new_n3464_));
  OAI21_X1   g02462(.A1(new_n3463_), .A2(new_n3464_), .B(new_n3461_), .ZN(new_n3465_));
  NAND2_X1   g02463(.A1(new_n3460_), .A2(new_n3465_), .ZN(new_n3466_));
  NAND2_X1   g02464(.A1(new_n3455_), .A2(new_n3466_), .ZN(new_n3467_));
  NOR2_X1    g02465(.A1(new_n3448_), .A2(\A[452] ), .ZN(new_n3468_));
  NOR2_X1    g02466(.A1(new_n3446_), .A2(\A[453] ), .ZN(new_n3469_));
  OAI21_X1   g02467(.A1(new_n3468_), .A2(new_n3469_), .B(\A[451] ), .ZN(new_n3470_));
  AND2_X2    g02468(.A1(\A[452] ), .A2(\A[453] ), .Z(new_n3471_));
  OAI21_X1   g02469(.A1(new_n3471_), .A2(new_n3452_), .B(new_n3445_), .ZN(new_n3472_));
  NAND2_X1   g02470(.A1(new_n3470_), .A2(new_n3472_), .ZN(new_n3473_));
  NAND2_X1   g02471(.A1(new_n3458_), .A2(\A[456] ), .ZN(new_n3474_));
  NAND2_X1   g02472(.A1(new_n3456_), .A2(\A[455] ), .ZN(new_n3475_));
  AOI21_X1   g02473(.A1(new_n3474_), .A2(new_n3475_), .B(new_n3461_), .ZN(new_n3476_));
  INV_X1     g02474(.I(new_n3464_), .ZN(new_n3477_));
  AOI21_X1   g02475(.A1(new_n3477_), .A2(new_n3462_), .B(\A[454] ), .ZN(new_n3478_));
  NOR2_X1    g02476(.A1(new_n3478_), .A2(new_n3476_), .ZN(new_n3479_));
  NAND2_X1   g02477(.A1(new_n3479_), .A2(new_n3473_), .ZN(new_n3480_));
  NAND2_X1   g02478(.A1(new_n3467_), .A2(new_n3480_), .ZN(new_n3481_));
  NOR2_X1    g02479(.A1(new_n3444_), .A2(new_n3481_), .ZN(new_n3482_));
  XOR2_X1    g02480(.A1(new_n3418_), .A2(new_n3428_), .Z(new_n3483_));
  NOR2_X1    g02481(.A1(new_n3479_), .A2(new_n3473_), .ZN(new_n3484_));
  NOR2_X1    g02482(.A1(new_n3455_), .A2(new_n3466_), .ZN(new_n3485_));
  NOR2_X1    g02483(.A1(new_n3485_), .A2(new_n3484_), .ZN(new_n3486_));
  NOR2_X1    g02484(.A1(new_n3483_), .A2(new_n3486_), .ZN(new_n3487_));
  INV_X1     g02485(.I(\A[445] ), .ZN(new_n3488_));
  INV_X1     g02486(.I(\A[446] ), .ZN(new_n3489_));
  NAND2_X1   g02487(.A1(new_n3489_), .A2(\A[447] ), .ZN(new_n3490_));
  INV_X1     g02488(.I(\A[447] ), .ZN(new_n3491_));
  NAND2_X1   g02489(.A1(new_n3491_), .A2(\A[446] ), .ZN(new_n3492_));
  AOI21_X1   g02490(.A1(new_n3490_), .A2(new_n3492_), .B(new_n3488_), .ZN(new_n3493_));
  NAND2_X1   g02491(.A1(\A[446] ), .A2(\A[447] ), .ZN(new_n3494_));
  NOR2_X1    g02492(.A1(\A[446] ), .A2(\A[447] ), .ZN(new_n3495_));
  INV_X1     g02493(.I(new_n3495_), .ZN(new_n3496_));
  AOI21_X1   g02494(.A1(new_n3496_), .A2(new_n3494_), .B(\A[445] ), .ZN(new_n3497_));
  NOR2_X1    g02495(.A1(new_n3497_), .A2(new_n3493_), .ZN(new_n3498_));
  INV_X1     g02496(.I(\A[450] ), .ZN(new_n3499_));
  NOR2_X1    g02497(.A1(new_n3499_), .A2(\A[449] ), .ZN(new_n3500_));
  INV_X1     g02498(.I(\A[449] ), .ZN(new_n3501_));
  NOR2_X1    g02499(.A1(new_n3501_), .A2(\A[450] ), .ZN(new_n3502_));
  OAI21_X1   g02500(.A1(new_n3500_), .A2(new_n3502_), .B(\A[448] ), .ZN(new_n3503_));
  INV_X1     g02501(.I(\A[448] ), .ZN(new_n3504_));
  NAND2_X1   g02502(.A1(\A[449] ), .A2(\A[450] ), .ZN(new_n3505_));
  INV_X1     g02503(.I(new_n3505_), .ZN(new_n3506_));
  NOR2_X1    g02504(.A1(\A[449] ), .A2(\A[450] ), .ZN(new_n3507_));
  OAI21_X1   g02505(.A1(new_n3506_), .A2(new_n3507_), .B(new_n3504_), .ZN(new_n3508_));
  NAND2_X1   g02506(.A1(new_n3503_), .A2(new_n3508_), .ZN(new_n3509_));
  NAND2_X1   g02507(.A1(new_n3498_), .A2(new_n3509_), .ZN(new_n3510_));
  NOR2_X1    g02508(.A1(new_n3491_), .A2(\A[446] ), .ZN(new_n3511_));
  NOR2_X1    g02509(.A1(new_n3489_), .A2(\A[447] ), .ZN(new_n3512_));
  OAI21_X1   g02510(.A1(new_n3511_), .A2(new_n3512_), .B(\A[445] ), .ZN(new_n3513_));
  INV_X1     g02511(.I(new_n3494_), .ZN(new_n3514_));
  OAI21_X1   g02512(.A1(new_n3514_), .A2(new_n3495_), .B(new_n3488_), .ZN(new_n3515_));
  NAND2_X1   g02513(.A1(new_n3513_), .A2(new_n3515_), .ZN(new_n3516_));
  NAND2_X1   g02514(.A1(new_n3501_), .A2(\A[450] ), .ZN(new_n3517_));
  NAND2_X1   g02515(.A1(new_n3499_), .A2(\A[449] ), .ZN(new_n3518_));
  AOI21_X1   g02516(.A1(new_n3517_), .A2(new_n3518_), .B(new_n3504_), .ZN(new_n3519_));
  INV_X1     g02517(.I(new_n3507_), .ZN(new_n3520_));
  AOI21_X1   g02518(.A1(new_n3520_), .A2(new_n3505_), .B(\A[448] ), .ZN(new_n3521_));
  NOR2_X1    g02519(.A1(new_n3521_), .A2(new_n3519_), .ZN(new_n3522_));
  NAND2_X1   g02520(.A1(new_n3522_), .A2(new_n3516_), .ZN(new_n3523_));
  INV_X1     g02521(.I(\A[439] ), .ZN(new_n3524_));
  INV_X1     g02522(.I(\A[440] ), .ZN(new_n3525_));
  NAND2_X1   g02523(.A1(new_n3525_), .A2(\A[441] ), .ZN(new_n3526_));
  INV_X1     g02524(.I(\A[441] ), .ZN(new_n3527_));
  NAND2_X1   g02525(.A1(new_n3527_), .A2(\A[440] ), .ZN(new_n3528_));
  AOI21_X1   g02526(.A1(new_n3526_), .A2(new_n3528_), .B(new_n3524_), .ZN(new_n3529_));
  NAND2_X1   g02527(.A1(\A[440] ), .A2(\A[441] ), .ZN(new_n3530_));
  NOR2_X1    g02528(.A1(\A[440] ), .A2(\A[441] ), .ZN(new_n3531_));
  INV_X1     g02529(.I(new_n3531_), .ZN(new_n3532_));
  AOI21_X1   g02530(.A1(new_n3532_), .A2(new_n3530_), .B(\A[439] ), .ZN(new_n3533_));
  NOR2_X1    g02531(.A1(new_n3533_), .A2(new_n3529_), .ZN(new_n3534_));
  INV_X1     g02532(.I(\A[444] ), .ZN(new_n3535_));
  NOR2_X1    g02533(.A1(new_n3535_), .A2(\A[443] ), .ZN(new_n3536_));
  INV_X1     g02534(.I(\A[443] ), .ZN(new_n3537_));
  NOR2_X1    g02535(.A1(new_n3537_), .A2(\A[444] ), .ZN(new_n3538_));
  OAI21_X1   g02536(.A1(new_n3536_), .A2(new_n3538_), .B(\A[442] ), .ZN(new_n3539_));
  INV_X1     g02537(.I(\A[442] ), .ZN(new_n3540_));
  NAND2_X1   g02538(.A1(\A[443] ), .A2(\A[444] ), .ZN(new_n3541_));
  INV_X1     g02539(.I(new_n3541_), .ZN(new_n3542_));
  NOR2_X1    g02540(.A1(\A[443] ), .A2(\A[444] ), .ZN(new_n3543_));
  OAI21_X1   g02541(.A1(new_n3542_), .A2(new_n3543_), .B(new_n3540_), .ZN(new_n3544_));
  NAND2_X1   g02542(.A1(new_n3539_), .A2(new_n3544_), .ZN(new_n3545_));
  NAND2_X1   g02543(.A1(new_n3534_), .A2(new_n3545_), .ZN(new_n3546_));
  NOR2_X1    g02544(.A1(new_n3527_), .A2(\A[440] ), .ZN(new_n3547_));
  NOR2_X1    g02545(.A1(new_n3525_), .A2(\A[441] ), .ZN(new_n3548_));
  OAI21_X1   g02546(.A1(new_n3547_), .A2(new_n3548_), .B(\A[439] ), .ZN(new_n3549_));
  AND2_X2    g02547(.A1(\A[440] ), .A2(\A[441] ), .Z(new_n3550_));
  OAI21_X1   g02548(.A1(new_n3550_), .A2(new_n3531_), .B(new_n3524_), .ZN(new_n3551_));
  NAND2_X1   g02549(.A1(new_n3549_), .A2(new_n3551_), .ZN(new_n3552_));
  NAND2_X1   g02550(.A1(new_n3537_), .A2(\A[444] ), .ZN(new_n3553_));
  NAND2_X1   g02551(.A1(new_n3535_), .A2(\A[443] ), .ZN(new_n3554_));
  AOI21_X1   g02552(.A1(new_n3553_), .A2(new_n3554_), .B(new_n3540_), .ZN(new_n3555_));
  INV_X1     g02553(.I(new_n3543_), .ZN(new_n3556_));
  AOI21_X1   g02554(.A1(new_n3556_), .A2(new_n3541_), .B(\A[442] ), .ZN(new_n3557_));
  NOR2_X1    g02555(.A1(new_n3557_), .A2(new_n3555_), .ZN(new_n3558_));
  NAND2_X1   g02556(.A1(new_n3558_), .A2(new_n3552_), .ZN(new_n3559_));
  AOI22_X1   g02557(.A1(new_n3510_), .A2(new_n3523_), .B1(new_n3546_), .B2(new_n3559_), .ZN(new_n3560_));
  NAND2_X1   g02558(.A1(new_n3523_), .A2(new_n3510_), .ZN(new_n3561_));
  NAND2_X1   g02559(.A1(new_n3546_), .A2(new_n3559_), .ZN(new_n3562_));
  NOR2_X1    g02560(.A1(new_n3561_), .A2(new_n3562_), .ZN(new_n3563_));
  NOR4_X1    g02561(.A1(new_n3487_), .A2(new_n3482_), .A3(new_n3563_), .A4(new_n3560_), .ZN(new_n3564_));
  NAND2_X1   g02562(.A1(new_n3483_), .A2(new_n3486_), .ZN(new_n3565_));
  NAND2_X1   g02563(.A1(new_n3444_), .A2(new_n3481_), .ZN(new_n3566_));
  NAND2_X1   g02564(.A1(new_n3561_), .A2(new_n3562_), .ZN(new_n3567_));
  NOR2_X1    g02565(.A1(new_n3522_), .A2(new_n3516_), .ZN(new_n3568_));
  NOR2_X1    g02566(.A1(new_n3498_), .A2(new_n3509_), .ZN(new_n3569_));
  NOR2_X1    g02567(.A1(new_n3568_), .A2(new_n3569_), .ZN(new_n3570_));
  NOR2_X1    g02568(.A1(new_n3558_), .A2(new_n3552_), .ZN(new_n3571_));
  NOR2_X1    g02569(.A1(new_n3534_), .A2(new_n3545_), .ZN(new_n3572_));
  NOR2_X1    g02570(.A1(new_n3572_), .A2(new_n3571_), .ZN(new_n3573_));
  NAND2_X1   g02571(.A1(new_n3570_), .A2(new_n3573_), .ZN(new_n3574_));
  AOI22_X1   g02572(.A1(new_n3565_), .A2(new_n3566_), .B1(new_n3574_), .B2(new_n3567_), .ZN(new_n3575_));
  NOR2_X1    g02573(.A1(new_n3575_), .A2(new_n3564_), .ZN(new_n3576_));
  INV_X1     g02574(.I(new_n3576_), .ZN(new_n3577_));
  INV_X1     g02575(.I(\A[423] ), .ZN(new_n3578_));
  NOR2_X1    g02576(.A1(new_n3578_), .A2(\A[422] ), .ZN(new_n3579_));
  INV_X1     g02577(.I(\A[422] ), .ZN(new_n3580_));
  NOR2_X1    g02578(.A1(new_n3580_), .A2(\A[423] ), .ZN(new_n3581_));
  OAI21_X1   g02579(.A1(new_n3579_), .A2(new_n3581_), .B(\A[421] ), .ZN(new_n3582_));
  INV_X1     g02580(.I(\A[421] ), .ZN(new_n3583_));
  NOR2_X1    g02581(.A1(\A[422] ), .A2(\A[423] ), .ZN(new_n3584_));
  NAND2_X1   g02582(.A1(\A[422] ), .A2(\A[423] ), .ZN(new_n3585_));
  INV_X1     g02583(.I(new_n3585_), .ZN(new_n3586_));
  OAI21_X1   g02584(.A1(new_n3586_), .A2(new_n3584_), .B(new_n3583_), .ZN(new_n3587_));
  INV_X1     g02585(.I(\A[426] ), .ZN(new_n3588_));
  NOR2_X1    g02586(.A1(new_n3588_), .A2(\A[425] ), .ZN(new_n3589_));
  INV_X1     g02587(.I(\A[425] ), .ZN(new_n3590_));
  NOR2_X1    g02588(.A1(new_n3590_), .A2(\A[426] ), .ZN(new_n3591_));
  OAI21_X1   g02589(.A1(new_n3589_), .A2(new_n3591_), .B(\A[424] ), .ZN(new_n3592_));
  INV_X1     g02590(.I(\A[424] ), .ZN(new_n3593_));
  NOR2_X1    g02591(.A1(\A[425] ), .A2(\A[426] ), .ZN(new_n3594_));
  AND2_X2    g02592(.A1(\A[425] ), .A2(\A[426] ), .Z(new_n3595_));
  OAI21_X1   g02593(.A1(new_n3595_), .A2(new_n3594_), .B(new_n3593_), .ZN(new_n3596_));
  NAND4_X1   g02594(.A1(new_n3582_), .A2(new_n3592_), .A3(new_n3587_), .A4(new_n3596_), .ZN(new_n3597_));
  NAND2_X1   g02595(.A1(new_n3580_), .A2(\A[423] ), .ZN(new_n3598_));
  NAND2_X1   g02596(.A1(new_n3578_), .A2(\A[422] ), .ZN(new_n3599_));
  AOI21_X1   g02597(.A1(new_n3598_), .A2(new_n3599_), .B(new_n3583_), .ZN(new_n3600_));
  INV_X1     g02598(.I(new_n3584_), .ZN(new_n3601_));
  AOI21_X1   g02599(.A1(new_n3601_), .A2(new_n3585_), .B(\A[421] ), .ZN(new_n3602_));
  NAND2_X1   g02600(.A1(new_n3590_), .A2(\A[426] ), .ZN(new_n3603_));
  NAND2_X1   g02601(.A1(new_n3588_), .A2(\A[425] ), .ZN(new_n3604_));
  AOI21_X1   g02602(.A1(new_n3603_), .A2(new_n3604_), .B(new_n3593_), .ZN(new_n3605_));
  INV_X1     g02603(.I(new_n3594_), .ZN(new_n3606_));
  NAND2_X1   g02604(.A1(\A[425] ), .A2(\A[426] ), .ZN(new_n3607_));
  AOI21_X1   g02605(.A1(new_n3606_), .A2(new_n3607_), .B(\A[424] ), .ZN(new_n3608_));
  OAI22_X1   g02606(.A1(new_n3600_), .A2(new_n3602_), .B1(new_n3608_), .B2(new_n3605_), .ZN(new_n3609_));
  NAND2_X1   g02607(.A1(new_n3609_), .A2(new_n3597_), .ZN(new_n3610_));
  INV_X1     g02608(.I(\A[415] ), .ZN(new_n3611_));
  INV_X1     g02609(.I(\A[416] ), .ZN(new_n3612_));
  NAND2_X1   g02610(.A1(new_n3612_), .A2(\A[417] ), .ZN(new_n3613_));
  INV_X1     g02611(.I(\A[417] ), .ZN(new_n3614_));
  NAND2_X1   g02612(.A1(new_n3614_), .A2(\A[416] ), .ZN(new_n3615_));
  AOI21_X1   g02613(.A1(new_n3613_), .A2(new_n3615_), .B(new_n3611_), .ZN(new_n3616_));
  NAND2_X1   g02614(.A1(\A[416] ), .A2(\A[417] ), .ZN(new_n3617_));
  NOR2_X1    g02615(.A1(\A[416] ), .A2(\A[417] ), .ZN(new_n3618_));
  INV_X1     g02616(.I(new_n3618_), .ZN(new_n3619_));
  AOI21_X1   g02617(.A1(new_n3619_), .A2(new_n3617_), .B(\A[415] ), .ZN(new_n3620_));
  INV_X1     g02618(.I(\A[418] ), .ZN(new_n3621_));
  INV_X1     g02619(.I(\A[419] ), .ZN(new_n3622_));
  NAND2_X1   g02620(.A1(new_n3622_), .A2(\A[420] ), .ZN(new_n3623_));
  INV_X1     g02621(.I(\A[420] ), .ZN(new_n3624_));
  NAND2_X1   g02622(.A1(new_n3624_), .A2(\A[419] ), .ZN(new_n3625_));
  AOI21_X1   g02623(.A1(new_n3623_), .A2(new_n3625_), .B(new_n3621_), .ZN(new_n3626_));
  NAND2_X1   g02624(.A1(\A[419] ), .A2(\A[420] ), .ZN(new_n3627_));
  OR2_X2     g02625(.A1(\A[419] ), .A2(\A[420] ), .Z(new_n3628_));
  AOI21_X1   g02626(.A1(new_n3628_), .A2(new_n3627_), .B(\A[418] ), .ZN(new_n3629_));
  NOR4_X1    g02627(.A1(new_n3616_), .A2(new_n3620_), .A3(new_n3626_), .A4(new_n3629_), .ZN(new_n3630_));
  NOR2_X1    g02628(.A1(new_n3614_), .A2(\A[416] ), .ZN(new_n3631_));
  NOR2_X1    g02629(.A1(new_n3612_), .A2(\A[417] ), .ZN(new_n3632_));
  OAI21_X1   g02630(.A1(new_n3631_), .A2(new_n3632_), .B(\A[415] ), .ZN(new_n3633_));
  INV_X1     g02631(.I(new_n3617_), .ZN(new_n3634_));
  OAI21_X1   g02632(.A1(new_n3634_), .A2(new_n3618_), .B(new_n3611_), .ZN(new_n3635_));
  NOR2_X1    g02633(.A1(new_n3624_), .A2(\A[419] ), .ZN(new_n3636_));
  NOR2_X1    g02634(.A1(new_n3622_), .A2(\A[420] ), .ZN(new_n3637_));
  OAI21_X1   g02635(.A1(new_n3636_), .A2(new_n3637_), .B(\A[418] ), .ZN(new_n3638_));
  INV_X1     g02636(.I(new_n3627_), .ZN(new_n3639_));
  NOR2_X1    g02637(.A1(\A[419] ), .A2(\A[420] ), .ZN(new_n3640_));
  OAI21_X1   g02638(.A1(new_n3639_), .A2(new_n3640_), .B(new_n3621_), .ZN(new_n3641_));
  AOI22_X1   g02639(.A1(new_n3633_), .A2(new_n3635_), .B1(new_n3638_), .B2(new_n3641_), .ZN(new_n3642_));
  NOR2_X1    g02640(.A1(new_n3642_), .A2(new_n3630_), .ZN(new_n3643_));
  NAND2_X1   g02641(.A1(new_n3643_), .A2(new_n3610_), .ZN(new_n3644_));
  NOR4_X1    g02642(.A1(new_n3600_), .A2(new_n3602_), .A3(new_n3608_), .A4(new_n3605_), .ZN(new_n3645_));
  AOI22_X1   g02643(.A1(new_n3582_), .A2(new_n3587_), .B1(new_n3592_), .B2(new_n3596_), .ZN(new_n3646_));
  NOR2_X1    g02644(.A1(new_n3645_), .A2(new_n3646_), .ZN(new_n3647_));
  NAND4_X1   g02645(.A1(new_n3633_), .A2(new_n3635_), .A3(new_n3638_), .A4(new_n3641_), .ZN(new_n3648_));
  OAI22_X1   g02646(.A1(new_n3616_), .A2(new_n3620_), .B1(new_n3626_), .B2(new_n3629_), .ZN(new_n3649_));
  NAND2_X1   g02647(.A1(new_n3648_), .A2(new_n3649_), .ZN(new_n3650_));
  NAND2_X1   g02648(.A1(new_n3647_), .A2(new_n3650_), .ZN(new_n3651_));
  NAND2_X1   g02649(.A1(new_n3651_), .A2(new_n3644_), .ZN(new_n3652_));
  INV_X1     g02650(.I(new_n3652_), .ZN(new_n3653_));
  INV_X1     g02651(.I(\A[427] ), .ZN(new_n3654_));
  INV_X1     g02652(.I(\A[428] ), .ZN(new_n3655_));
  NAND2_X1   g02653(.A1(new_n3655_), .A2(\A[429] ), .ZN(new_n3656_));
  INV_X1     g02654(.I(\A[429] ), .ZN(new_n3657_));
  NAND2_X1   g02655(.A1(new_n3657_), .A2(\A[428] ), .ZN(new_n3658_));
  AOI21_X1   g02656(.A1(new_n3656_), .A2(new_n3658_), .B(new_n3654_), .ZN(new_n3659_));
  NAND2_X1   g02657(.A1(\A[428] ), .A2(\A[429] ), .ZN(new_n3660_));
  NOR2_X1    g02658(.A1(\A[428] ), .A2(\A[429] ), .ZN(new_n3661_));
  INV_X1     g02659(.I(new_n3661_), .ZN(new_n3662_));
  AOI21_X1   g02660(.A1(new_n3662_), .A2(new_n3660_), .B(\A[427] ), .ZN(new_n3663_));
  INV_X1     g02661(.I(\A[430] ), .ZN(new_n3664_));
  INV_X1     g02662(.I(\A[431] ), .ZN(new_n3665_));
  NAND2_X1   g02663(.A1(new_n3665_), .A2(\A[432] ), .ZN(new_n3666_));
  INV_X1     g02664(.I(\A[432] ), .ZN(new_n3667_));
  NAND2_X1   g02665(.A1(new_n3667_), .A2(\A[431] ), .ZN(new_n3668_));
  AOI21_X1   g02666(.A1(new_n3666_), .A2(new_n3668_), .B(new_n3664_), .ZN(new_n3669_));
  NAND2_X1   g02667(.A1(\A[431] ), .A2(\A[432] ), .ZN(new_n3670_));
  NOR2_X1    g02668(.A1(\A[431] ), .A2(\A[432] ), .ZN(new_n3671_));
  INV_X1     g02669(.I(new_n3671_), .ZN(new_n3672_));
  AOI21_X1   g02670(.A1(new_n3672_), .A2(new_n3670_), .B(\A[430] ), .ZN(new_n3673_));
  NOR4_X1    g02671(.A1(new_n3659_), .A2(new_n3663_), .A3(new_n3673_), .A4(new_n3669_), .ZN(new_n3674_));
  NOR2_X1    g02672(.A1(new_n3657_), .A2(\A[428] ), .ZN(new_n3675_));
  NOR2_X1    g02673(.A1(new_n3655_), .A2(\A[429] ), .ZN(new_n3676_));
  OAI21_X1   g02674(.A1(new_n3675_), .A2(new_n3676_), .B(\A[427] ), .ZN(new_n3677_));
  INV_X1     g02675(.I(new_n3660_), .ZN(new_n3678_));
  OAI21_X1   g02676(.A1(new_n3678_), .A2(new_n3661_), .B(new_n3654_), .ZN(new_n3679_));
  NOR2_X1    g02677(.A1(new_n3667_), .A2(\A[431] ), .ZN(new_n3680_));
  NOR2_X1    g02678(.A1(new_n3665_), .A2(\A[432] ), .ZN(new_n3681_));
  OAI21_X1   g02679(.A1(new_n3680_), .A2(new_n3681_), .B(\A[430] ), .ZN(new_n3682_));
  AND2_X2    g02680(.A1(\A[431] ), .A2(\A[432] ), .Z(new_n3683_));
  OAI21_X1   g02681(.A1(new_n3683_), .A2(new_n3671_), .B(new_n3664_), .ZN(new_n3684_));
  AOI22_X1   g02682(.A1(new_n3677_), .A2(new_n3679_), .B1(new_n3682_), .B2(new_n3684_), .ZN(new_n3685_));
  INV_X1     g02683(.I(\A[433] ), .ZN(new_n3686_));
  INV_X1     g02684(.I(\A[434] ), .ZN(new_n3687_));
  NAND2_X1   g02685(.A1(new_n3687_), .A2(\A[435] ), .ZN(new_n3688_));
  INV_X1     g02686(.I(\A[435] ), .ZN(new_n3689_));
  NAND2_X1   g02687(.A1(new_n3689_), .A2(\A[434] ), .ZN(new_n3690_));
  AOI21_X1   g02688(.A1(new_n3688_), .A2(new_n3690_), .B(new_n3686_), .ZN(new_n3691_));
  NAND2_X1   g02689(.A1(\A[434] ), .A2(\A[435] ), .ZN(new_n3692_));
  NOR2_X1    g02690(.A1(\A[434] ), .A2(\A[435] ), .ZN(new_n3693_));
  INV_X1     g02691(.I(new_n3693_), .ZN(new_n3694_));
  AOI21_X1   g02692(.A1(new_n3694_), .A2(new_n3692_), .B(\A[433] ), .ZN(new_n3695_));
  INV_X1     g02693(.I(\A[436] ), .ZN(new_n3696_));
  INV_X1     g02694(.I(\A[437] ), .ZN(new_n3697_));
  NAND2_X1   g02695(.A1(new_n3697_), .A2(\A[438] ), .ZN(new_n3698_));
  INV_X1     g02696(.I(\A[438] ), .ZN(new_n3699_));
  NAND2_X1   g02697(.A1(new_n3699_), .A2(\A[437] ), .ZN(new_n3700_));
  AOI21_X1   g02698(.A1(new_n3698_), .A2(new_n3700_), .B(new_n3696_), .ZN(new_n3701_));
  NAND2_X1   g02699(.A1(\A[437] ), .A2(\A[438] ), .ZN(new_n3702_));
  NOR2_X1    g02700(.A1(\A[437] ), .A2(\A[438] ), .ZN(new_n3703_));
  INV_X1     g02701(.I(new_n3703_), .ZN(new_n3704_));
  AOI21_X1   g02702(.A1(new_n3704_), .A2(new_n3702_), .B(\A[436] ), .ZN(new_n3705_));
  NOR4_X1    g02703(.A1(new_n3691_), .A2(new_n3695_), .A3(new_n3705_), .A4(new_n3701_), .ZN(new_n3706_));
  NOR2_X1    g02704(.A1(new_n3689_), .A2(\A[434] ), .ZN(new_n3707_));
  NOR2_X1    g02705(.A1(new_n3687_), .A2(\A[435] ), .ZN(new_n3708_));
  OAI21_X1   g02706(.A1(new_n3707_), .A2(new_n3708_), .B(\A[433] ), .ZN(new_n3709_));
  INV_X1     g02707(.I(new_n3692_), .ZN(new_n3710_));
  OAI21_X1   g02708(.A1(new_n3710_), .A2(new_n3693_), .B(new_n3686_), .ZN(new_n3711_));
  NOR2_X1    g02709(.A1(new_n3699_), .A2(\A[437] ), .ZN(new_n3712_));
  NOR2_X1    g02710(.A1(new_n3697_), .A2(\A[438] ), .ZN(new_n3713_));
  OAI21_X1   g02711(.A1(new_n3712_), .A2(new_n3713_), .B(\A[436] ), .ZN(new_n3714_));
  AND2_X2    g02712(.A1(\A[437] ), .A2(\A[438] ), .Z(new_n3715_));
  OAI21_X1   g02713(.A1(new_n3715_), .A2(new_n3703_), .B(new_n3696_), .ZN(new_n3716_));
  AOI22_X1   g02714(.A1(new_n3709_), .A2(new_n3711_), .B1(new_n3714_), .B2(new_n3716_), .ZN(new_n3717_));
  OAI22_X1   g02715(.A1(new_n3674_), .A2(new_n3685_), .B1(new_n3706_), .B2(new_n3717_), .ZN(new_n3718_));
  NAND4_X1   g02716(.A1(new_n3677_), .A2(new_n3682_), .A3(new_n3679_), .A4(new_n3684_), .ZN(new_n3719_));
  OAI22_X1   g02717(.A1(new_n3659_), .A2(new_n3663_), .B1(new_n3673_), .B2(new_n3669_), .ZN(new_n3720_));
  NAND4_X1   g02718(.A1(new_n3709_), .A2(new_n3714_), .A3(new_n3711_), .A4(new_n3716_), .ZN(new_n3721_));
  OAI22_X1   g02719(.A1(new_n3691_), .A2(new_n3695_), .B1(new_n3705_), .B2(new_n3701_), .ZN(new_n3722_));
  NAND4_X1   g02720(.A1(new_n3720_), .A2(new_n3722_), .A3(new_n3719_), .A4(new_n3721_), .ZN(new_n3723_));
  NAND2_X1   g02721(.A1(new_n3718_), .A2(new_n3723_), .ZN(new_n3724_));
  NAND2_X1   g02722(.A1(new_n3653_), .A2(new_n3724_), .ZN(new_n3725_));
  INV_X1     g02723(.I(new_n3724_), .ZN(new_n3726_));
  NAND2_X1   g02724(.A1(new_n3726_), .A2(new_n3652_), .ZN(new_n3727_));
  NAND2_X1   g02725(.A1(new_n3725_), .A2(new_n3727_), .ZN(new_n3728_));
  NOR2_X1    g02726(.A1(new_n3577_), .A2(new_n3728_), .ZN(new_n3729_));
  NOR2_X1    g02727(.A1(new_n3726_), .A2(new_n3652_), .ZN(new_n3730_));
  AOI21_X1   g02728(.A1(new_n3644_), .A2(new_n3651_), .B(new_n3724_), .ZN(new_n3731_));
  NOR2_X1    g02729(.A1(new_n3730_), .A2(new_n3731_), .ZN(new_n3732_));
  NOR2_X1    g02730(.A1(new_n3576_), .A2(new_n3732_), .ZN(new_n3733_));
  NOR2_X1    g02731(.A1(new_n3729_), .A2(new_n3733_), .ZN(new_n3734_));
  NAND2_X1   g02732(.A1(new_n3734_), .A2(new_n3407_), .ZN(new_n3735_));
  OAI22_X1   g02733(.A1(new_n3729_), .A2(new_n3733_), .B1(new_n3402_), .B2(new_n3406_), .ZN(new_n3736_));
  NAND2_X1   g02734(.A1(new_n3735_), .A2(new_n3736_), .ZN(new_n3737_));
  INV_X1     g02735(.I(\A[361] ), .ZN(new_n3738_));
  INV_X1     g02736(.I(\A[362] ), .ZN(new_n3739_));
  NAND2_X1   g02737(.A1(new_n3739_), .A2(\A[363] ), .ZN(new_n3740_));
  INV_X1     g02738(.I(\A[363] ), .ZN(new_n3741_));
  NAND2_X1   g02739(.A1(new_n3741_), .A2(\A[362] ), .ZN(new_n3742_));
  AOI21_X1   g02740(.A1(new_n3740_), .A2(new_n3742_), .B(new_n3738_), .ZN(new_n3743_));
  NAND2_X1   g02741(.A1(\A[362] ), .A2(\A[363] ), .ZN(new_n3744_));
  NOR2_X1    g02742(.A1(\A[362] ), .A2(\A[363] ), .ZN(new_n3745_));
  INV_X1     g02743(.I(new_n3745_), .ZN(new_n3746_));
  AOI21_X1   g02744(.A1(new_n3746_), .A2(new_n3744_), .B(\A[361] ), .ZN(new_n3747_));
  NOR2_X1    g02745(.A1(new_n3747_), .A2(new_n3743_), .ZN(new_n3748_));
  INV_X1     g02746(.I(\A[366] ), .ZN(new_n3749_));
  NOR2_X1    g02747(.A1(new_n3749_), .A2(\A[365] ), .ZN(new_n3750_));
  INV_X1     g02748(.I(\A[365] ), .ZN(new_n3751_));
  NOR2_X1    g02749(.A1(new_n3751_), .A2(\A[366] ), .ZN(new_n3752_));
  OAI21_X1   g02750(.A1(new_n3750_), .A2(new_n3752_), .B(\A[364] ), .ZN(new_n3753_));
  INV_X1     g02751(.I(\A[364] ), .ZN(new_n3754_));
  AND2_X2    g02752(.A1(\A[365] ), .A2(\A[366] ), .Z(new_n3755_));
  NOR2_X1    g02753(.A1(\A[365] ), .A2(\A[366] ), .ZN(new_n3756_));
  OAI21_X1   g02754(.A1(new_n3755_), .A2(new_n3756_), .B(new_n3754_), .ZN(new_n3757_));
  NAND2_X1   g02755(.A1(new_n3753_), .A2(new_n3757_), .ZN(new_n3758_));
  NAND2_X1   g02756(.A1(new_n3748_), .A2(new_n3758_), .ZN(new_n3759_));
  NOR2_X1    g02757(.A1(new_n3741_), .A2(\A[362] ), .ZN(new_n3760_));
  NOR2_X1    g02758(.A1(new_n3739_), .A2(\A[363] ), .ZN(new_n3761_));
  OAI21_X1   g02759(.A1(new_n3760_), .A2(new_n3761_), .B(\A[361] ), .ZN(new_n3762_));
  INV_X1     g02760(.I(new_n3744_), .ZN(new_n3763_));
  OAI21_X1   g02761(.A1(new_n3763_), .A2(new_n3745_), .B(new_n3738_), .ZN(new_n3764_));
  NAND2_X1   g02762(.A1(new_n3762_), .A2(new_n3764_), .ZN(new_n3765_));
  NAND2_X1   g02763(.A1(new_n3751_), .A2(\A[366] ), .ZN(new_n3766_));
  NAND2_X1   g02764(.A1(new_n3749_), .A2(\A[365] ), .ZN(new_n3767_));
  AOI21_X1   g02765(.A1(new_n3766_), .A2(new_n3767_), .B(new_n3754_), .ZN(new_n3768_));
  NAND2_X1   g02766(.A1(\A[365] ), .A2(\A[366] ), .ZN(new_n3769_));
  INV_X1     g02767(.I(new_n3756_), .ZN(new_n3770_));
  AOI21_X1   g02768(.A1(new_n3770_), .A2(new_n3769_), .B(\A[364] ), .ZN(new_n3771_));
  NOR2_X1    g02769(.A1(new_n3771_), .A2(new_n3768_), .ZN(new_n3772_));
  NAND2_X1   g02770(.A1(new_n3772_), .A2(new_n3765_), .ZN(new_n3773_));
  NAND2_X1   g02771(.A1(new_n3773_), .A2(new_n3759_), .ZN(new_n3774_));
  INV_X1     g02772(.I(\A[355] ), .ZN(new_n3775_));
  INV_X1     g02773(.I(\A[356] ), .ZN(new_n3776_));
  NAND2_X1   g02774(.A1(new_n3776_), .A2(\A[357] ), .ZN(new_n3777_));
  INV_X1     g02775(.I(\A[357] ), .ZN(new_n3778_));
  NAND2_X1   g02776(.A1(new_n3778_), .A2(\A[356] ), .ZN(new_n3779_));
  AOI21_X1   g02777(.A1(new_n3777_), .A2(new_n3779_), .B(new_n3775_), .ZN(new_n3780_));
  NAND2_X1   g02778(.A1(\A[356] ), .A2(\A[357] ), .ZN(new_n3781_));
  NOR2_X1    g02779(.A1(\A[356] ), .A2(\A[357] ), .ZN(new_n3782_));
  INV_X1     g02780(.I(new_n3782_), .ZN(new_n3783_));
  AOI21_X1   g02781(.A1(new_n3783_), .A2(new_n3781_), .B(\A[355] ), .ZN(new_n3784_));
  NOR2_X1    g02782(.A1(new_n3784_), .A2(new_n3780_), .ZN(new_n3785_));
  INV_X1     g02783(.I(\A[360] ), .ZN(new_n3786_));
  NOR2_X1    g02784(.A1(new_n3786_), .A2(\A[359] ), .ZN(new_n3787_));
  INV_X1     g02785(.I(\A[359] ), .ZN(new_n3788_));
  NOR2_X1    g02786(.A1(new_n3788_), .A2(\A[360] ), .ZN(new_n3789_));
  OAI21_X1   g02787(.A1(new_n3787_), .A2(new_n3789_), .B(\A[358] ), .ZN(new_n3790_));
  INV_X1     g02788(.I(\A[358] ), .ZN(new_n3791_));
  NAND2_X1   g02789(.A1(\A[359] ), .A2(\A[360] ), .ZN(new_n3792_));
  INV_X1     g02790(.I(new_n3792_), .ZN(new_n3793_));
  NOR2_X1    g02791(.A1(\A[359] ), .A2(\A[360] ), .ZN(new_n3794_));
  OAI21_X1   g02792(.A1(new_n3793_), .A2(new_n3794_), .B(new_n3791_), .ZN(new_n3795_));
  NAND2_X1   g02793(.A1(new_n3790_), .A2(new_n3795_), .ZN(new_n3796_));
  NAND2_X1   g02794(.A1(new_n3785_), .A2(new_n3796_), .ZN(new_n3797_));
  NOR2_X1    g02795(.A1(new_n3778_), .A2(\A[356] ), .ZN(new_n3798_));
  NOR2_X1    g02796(.A1(new_n3776_), .A2(\A[357] ), .ZN(new_n3799_));
  OAI21_X1   g02797(.A1(new_n3798_), .A2(new_n3799_), .B(\A[355] ), .ZN(new_n3800_));
  AND2_X2    g02798(.A1(\A[356] ), .A2(\A[357] ), .Z(new_n3801_));
  OAI21_X1   g02799(.A1(new_n3801_), .A2(new_n3782_), .B(new_n3775_), .ZN(new_n3802_));
  NAND2_X1   g02800(.A1(new_n3800_), .A2(new_n3802_), .ZN(new_n3803_));
  NAND2_X1   g02801(.A1(new_n3788_), .A2(\A[360] ), .ZN(new_n3804_));
  NAND2_X1   g02802(.A1(new_n3786_), .A2(\A[359] ), .ZN(new_n3805_));
  AOI21_X1   g02803(.A1(new_n3804_), .A2(new_n3805_), .B(new_n3791_), .ZN(new_n3806_));
  INV_X1     g02804(.I(new_n3794_), .ZN(new_n3807_));
  AOI21_X1   g02805(.A1(new_n3807_), .A2(new_n3792_), .B(\A[358] ), .ZN(new_n3808_));
  NOR2_X1    g02806(.A1(new_n3808_), .A2(new_n3806_), .ZN(new_n3809_));
  NAND2_X1   g02807(.A1(new_n3809_), .A2(new_n3803_), .ZN(new_n3810_));
  NAND2_X1   g02808(.A1(new_n3797_), .A2(new_n3810_), .ZN(new_n3811_));
  NOR2_X1    g02809(.A1(new_n3774_), .A2(new_n3811_), .ZN(new_n3812_));
  XOR2_X1    g02810(.A1(new_n3748_), .A2(new_n3758_), .Z(new_n3813_));
  NOR2_X1    g02811(.A1(new_n3809_), .A2(new_n3803_), .ZN(new_n3814_));
  NOR2_X1    g02812(.A1(new_n3785_), .A2(new_n3796_), .ZN(new_n3815_));
  NOR2_X1    g02813(.A1(new_n3815_), .A2(new_n3814_), .ZN(new_n3816_));
  NOR2_X1    g02814(.A1(new_n3813_), .A2(new_n3816_), .ZN(new_n3817_));
  INV_X1     g02815(.I(\A[349] ), .ZN(new_n3818_));
  INV_X1     g02816(.I(\A[350] ), .ZN(new_n3819_));
  NAND2_X1   g02817(.A1(new_n3819_), .A2(\A[351] ), .ZN(new_n3820_));
  INV_X1     g02818(.I(\A[351] ), .ZN(new_n3821_));
  NAND2_X1   g02819(.A1(new_n3821_), .A2(\A[350] ), .ZN(new_n3822_));
  AOI21_X1   g02820(.A1(new_n3820_), .A2(new_n3822_), .B(new_n3818_), .ZN(new_n3823_));
  NAND2_X1   g02821(.A1(\A[350] ), .A2(\A[351] ), .ZN(new_n3824_));
  NOR2_X1    g02822(.A1(\A[350] ), .A2(\A[351] ), .ZN(new_n3825_));
  INV_X1     g02823(.I(new_n3825_), .ZN(new_n3826_));
  AOI21_X1   g02824(.A1(new_n3826_), .A2(new_n3824_), .B(\A[349] ), .ZN(new_n3827_));
  NOR2_X1    g02825(.A1(new_n3827_), .A2(new_n3823_), .ZN(new_n3828_));
  INV_X1     g02826(.I(\A[354] ), .ZN(new_n3829_));
  NOR2_X1    g02827(.A1(new_n3829_), .A2(\A[353] ), .ZN(new_n3830_));
  INV_X1     g02828(.I(\A[353] ), .ZN(new_n3831_));
  NOR2_X1    g02829(.A1(new_n3831_), .A2(\A[354] ), .ZN(new_n3832_));
  OAI21_X1   g02830(.A1(new_n3830_), .A2(new_n3832_), .B(\A[352] ), .ZN(new_n3833_));
  INV_X1     g02831(.I(\A[352] ), .ZN(new_n3834_));
  AND2_X2    g02832(.A1(\A[353] ), .A2(\A[354] ), .Z(new_n3835_));
  NOR2_X1    g02833(.A1(\A[353] ), .A2(\A[354] ), .ZN(new_n3836_));
  OAI21_X1   g02834(.A1(new_n3835_), .A2(new_n3836_), .B(new_n3834_), .ZN(new_n3837_));
  NAND2_X1   g02835(.A1(new_n3833_), .A2(new_n3837_), .ZN(new_n3838_));
  NAND2_X1   g02836(.A1(new_n3828_), .A2(new_n3838_), .ZN(new_n3839_));
  NOR2_X1    g02837(.A1(new_n3821_), .A2(\A[350] ), .ZN(new_n3840_));
  NOR2_X1    g02838(.A1(new_n3819_), .A2(\A[351] ), .ZN(new_n3841_));
  OAI21_X1   g02839(.A1(new_n3840_), .A2(new_n3841_), .B(\A[349] ), .ZN(new_n3842_));
  INV_X1     g02840(.I(new_n3824_), .ZN(new_n3843_));
  OAI21_X1   g02841(.A1(new_n3843_), .A2(new_n3825_), .B(new_n3818_), .ZN(new_n3844_));
  NAND2_X1   g02842(.A1(new_n3842_), .A2(new_n3844_), .ZN(new_n3845_));
  NAND2_X1   g02843(.A1(new_n3831_), .A2(\A[354] ), .ZN(new_n3846_));
  NAND2_X1   g02844(.A1(new_n3829_), .A2(\A[353] ), .ZN(new_n3847_));
  AOI21_X1   g02845(.A1(new_n3846_), .A2(new_n3847_), .B(new_n3834_), .ZN(new_n3848_));
  NAND2_X1   g02846(.A1(\A[353] ), .A2(\A[354] ), .ZN(new_n3849_));
  INV_X1     g02847(.I(new_n3836_), .ZN(new_n3850_));
  AOI21_X1   g02848(.A1(new_n3850_), .A2(new_n3849_), .B(\A[352] ), .ZN(new_n3851_));
  NOR2_X1    g02849(.A1(new_n3851_), .A2(new_n3848_), .ZN(new_n3852_));
  NAND2_X1   g02850(.A1(new_n3852_), .A2(new_n3845_), .ZN(new_n3853_));
  INV_X1     g02851(.I(\A[343] ), .ZN(new_n3854_));
  INV_X1     g02852(.I(\A[344] ), .ZN(new_n3855_));
  NAND2_X1   g02853(.A1(new_n3855_), .A2(\A[345] ), .ZN(new_n3856_));
  INV_X1     g02854(.I(\A[345] ), .ZN(new_n3857_));
  NAND2_X1   g02855(.A1(new_n3857_), .A2(\A[344] ), .ZN(new_n3858_));
  AOI21_X1   g02856(.A1(new_n3856_), .A2(new_n3858_), .B(new_n3854_), .ZN(new_n3859_));
  NAND2_X1   g02857(.A1(\A[344] ), .A2(\A[345] ), .ZN(new_n3860_));
  NOR2_X1    g02858(.A1(\A[344] ), .A2(\A[345] ), .ZN(new_n3861_));
  INV_X1     g02859(.I(new_n3861_), .ZN(new_n3862_));
  AOI21_X1   g02860(.A1(new_n3862_), .A2(new_n3860_), .B(\A[343] ), .ZN(new_n3863_));
  NOR2_X1    g02861(.A1(new_n3863_), .A2(new_n3859_), .ZN(new_n3864_));
  INV_X1     g02862(.I(\A[348] ), .ZN(new_n3865_));
  NOR2_X1    g02863(.A1(new_n3865_), .A2(\A[347] ), .ZN(new_n3866_));
  INV_X1     g02864(.I(\A[347] ), .ZN(new_n3867_));
  NOR2_X1    g02865(.A1(new_n3867_), .A2(\A[348] ), .ZN(new_n3868_));
  OAI21_X1   g02866(.A1(new_n3866_), .A2(new_n3868_), .B(\A[346] ), .ZN(new_n3869_));
  INV_X1     g02867(.I(\A[346] ), .ZN(new_n3870_));
  AND2_X2    g02868(.A1(\A[347] ), .A2(\A[348] ), .Z(new_n3871_));
  NOR2_X1    g02869(.A1(\A[347] ), .A2(\A[348] ), .ZN(new_n3872_));
  OAI21_X1   g02870(.A1(new_n3871_), .A2(new_n3872_), .B(new_n3870_), .ZN(new_n3873_));
  NAND2_X1   g02871(.A1(new_n3869_), .A2(new_n3873_), .ZN(new_n3874_));
  NAND2_X1   g02872(.A1(new_n3864_), .A2(new_n3874_), .ZN(new_n3875_));
  NOR2_X1    g02873(.A1(new_n3857_), .A2(\A[344] ), .ZN(new_n3876_));
  NOR2_X1    g02874(.A1(new_n3855_), .A2(\A[345] ), .ZN(new_n3877_));
  OAI21_X1   g02875(.A1(new_n3876_), .A2(new_n3877_), .B(\A[343] ), .ZN(new_n3878_));
  AND2_X2    g02876(.A1(\A[344] ), .A2(\A[345] ), .Z(new_n3879_));
  OAI21_X1   g02877(.A1(new_n3879_), .A2(new_n3861_), .B(new_n3854_), .ZN(new_n3880_));
  NAND2_X1   g02878(.A1(new_n3878_), .A2(new_n3880_), .ZN(new_n3881_));
  NAND2_X1   g02879(.A1(new_n3867_), .A2(\A[348] ), .ZN(new_n3882_));
  NAND2_X1   g02880(.A1(new_n3865_), .A2(\A[347] ), .ZN(new_n3883_));
  AOI21_X1   g02881(.A1(new_n3882_), .A2(new_n3883_), .B(new_n3870_), .ZN(new_n3884_));
  NAND2_X1   g02882(.A1(\A[347] ), .A2(\A[348] ), .ZN(new_n3885_));
  INV_X1     g02883(.I(new_n3872_), .ZN(new_n3886_));
  AOI21_X1   g02884(.A1(new_n3886_), .A2(new_n3885_), .B(\A[346] ), .ZN(new_n3887_));
  NOR2_X1    g02885(.A1(new_n3887_), .A2(new_n3884_), .ZN(new_n3888_));
  NAND2_X1   g02886(.A1(new_n3888_), .A2(new_n3881_), .ZN(new_n3889_));
  AOI22_X1   g02887(.A1(new_n3839_), .A2(new_n3853_), .B1(new_n3875_), .B2(new_n3889_), .ZN(new_n3890_));
  NAND2_X1   g02888(.A1(new_n3853_), .A2(new_n3839_), .ZN(new_n3891_));
  NAND2_X1   g02889(.A1(new_n3875_), .A2(new_n3889_), .ZN(new_n3892_));
  NOR2_X1    g02890(.A1(new_n3891_), .A2(new_n3892_), .ZN(new_n3893_));
  NOR4_X1    g02891(.A1(new_n3817_), .A2(new_n3812_), .A3(new_n3893_), .A4(new_n3890_), .ZN(new_n3894_));
  NAND2_X1   g02892(.A1(new_n3813_), .A2(new_n3816_), .ZN(new_n3895_));
  NAND2_X1   g02893(.A1(new_n3774_), .A2(new_n3811_), .ZN(new_n3896_));
  NAND2_X1   g02894(.A1(new_n3891_), .A2(new_n3892_), .ZN(new_n3897_));
  XOR2_X1    g02895(.A1(new_n3828_), .A2(new_n3838_), .Z(new_n3898_));
  NOR2_X1    g02896(.A1(new_n3888_), .A2(new_n3881_), .ZN(new_n3899_));
  NOR2_X1    g02897(.A1(new_n3864_), .A2(new_n3874_), .ZN(new_n3900_));
  NOR2_X1    g02898(.A1(new_n3899_), .A2(new_n3900_), .ZN(new_n3901_));
  NAND2_X1   g02899(.A1(new_n3898_), .A2(new_n3901_), .ZN(new_n3902_));
  AOI22_X1   g02900(.A1(new_n3895_), .A2(new_n3896_), .B1(new_n3902_), .B2(new_n3897_), .ZN(new_n3903_));
  NOR2_X1    g02901(.A1(new_n3903_), .A2(new_n3894_), .ZN(new_n3904_));
  INV_X1     g02902(.I(\A[327] ), .ZN(new_n3905_));
  NOR2_X1    g02903(.A1(new_n3905_), .A2(\A[326] ), .ZN(new_n3906_));
  INV_X1     g02904(.I(\A[326] ), .ZN(new_n3907_));
  NOR2_X1    g02905(.A1(new_n3907_), .A2(\A[327] ), .ZN(new_n3908_));
  OAI21_X1   g02906(.A1(new_n3906_), .A2(new_n3908_), .B(\A[325] ), .ZN(new_n3909_));
  INV_X1     g02907(.I(\A[325] ), .ZN(new_n3910_));
  NOR2_X1    g02908(.A1(\A[326] ), .A2(\A[327] ), .ZN(new_n3911_));
  NAND2_X1   g02909(.A1(\A[326] ), .A2(\A[327] ), .ZN(new_n3912_));
  INV_X1     g02910(.I(new_n3912_), .ZN(new_n3913_));
  OAI21_X1   g02911(.A1(new_n3913_), .A2(new_n3911_), .B(new_n3910_), .ZN(new_n3914_));
  INV_X1     g02912(.I(\A[330] ), .ZN(new_n3915_));
  NOR2_X1    g02913(.A1(new_n3915_), .A2(\A[329] ), .ZN(new_n3916_));
  INV_X1     g02914(.I(\A[329] ), .ZN(new_n3917_));
  NOR2_X1    g02915(.A1(new_n3917_), .A2(\A[330] ), .ZN(new_n3918_));
  OAI21_X1   g02916(.A1(new_n3916_), .A2(new_n3918_), .B(\A[328] ), .ZN(new_n3919_));
  INV_X1     g02917(.I(\A[328] ), .ZN(new_n3920_));
  NOR2_X1    g02918(.A1(\A[329] ), .A2(\A[330] ), .ZN(new_n3921_));
  AND2_X2    g02919(.A1(\A[329] ), .A2(\A[330] ), .Z(new_n3922_));
  OAI21_X1   g02920(.A1(new_n3922_), .A2(new_n3921_), .B(new_n3920_), .ZN(new_n3923_));
  NAND4_X1   g02921(.A1(new_n3909_), .A2(new_n3919_), .A3(new_n3914_), .A4(new_n3923_), .ZN(new_n3924_));
  NAND2_X1   g02922(.A1(new_n3907_), .A2(\A[327] ), .ZN(new_n3925_));
  NAND2_X1   g02923(.A1(new_n3905_), .A2(\A[326] ), .ZN(new_n3926_));
  AOI21_X1   g02924(.A1(new_n3925_), .A2(new_n3926_), .B(new_n3910_), .ZN(new_n3927_));
  INV_X1     g02925(.I(new_n3911_), .ZN(new_n3928_));
  AOI21_X1   g02926(.A1(new_n3928_), .A2(new_n3912_), .B(\A[325] ), .ZN(new_n3929_));
  NAND2_X1   g02927(.A1(new_n3917_), .A2(\A[330] ), .ZN(new_n3930_));
  NAND2_X1   g02928(.A1(new_n3915_), .A2(\A[329] ), .ZN(new_n3931_));
  AOI21_X1   g02929(.A1(new_n3930_), .A2(new_n3931_), .B(new_n3920_), .ZN(new_n3932_));
  INV_X1     g02930(.I(new_n3921_), .ZN(new_n3933_));
  NAND2_X1   g02931(.A1(\A[329] ), .A2(\A[330] ), .ZN(new_n3934_));
  AOI21_X1   g02932(.A1(new_n3933_), .A2(new_n3934_), .B(\A[328] ), .ZN(new_n3935_));
  OAI22_X1   g02933(.A1(new_n3927_), .A2(new_n3929_), .B1(new_n3935_), .B2(new_n3932_), .ZN(new_n3936_));
  NAND2_X1   g02934(.A1(new_n3936_), .A2(new_n3924_), .ZN(new_n3937_));
  INV_X1     g02935(.I(\A[319] ), .ZN(new_n3938_));
  INV_X1     g02936(.I(\A[320] ), .ZN(new_n3939_));
  NAND2_X1   g02937(.A1(new_n3939_), .A2(\A[321] ), .ZN(new_n3940_));
  INV_X1     g02938(.I(\A[321] ), .ZN(new_n3941_));
  NAND2_X1   g02939(.A1(new_n3941_), .A2(\A[320] ), .ZN(new_n3942_));
  AOI21_X1   g02940(.A1(new_n3940_), .A2(new_n3942_), .B(new_n3938_), .ZN(new_n3943_));
  NAND2_X1   g02941(.A1(\A[320] ), .A2(\A[321] ), .ZN(new_n3944_));
  NOR2_X1    g02942(.A1(\A[320] ), .A2(\A[321] ), .ZN(new_n3945_));
  INV_X1     g02943(.I(new_n3945_), .ZN(new_n3946_));
  AOI21_X1   g02944(.A1(new_n3946_), .A2(new_n3944_), .B(\A[319] ), .ZN(new_n3947_));
  INV_X1     g02945(.I(\A[322] ), .ZN(new_n3948_));
  INV_X1     g02946(.I(\A[323] ), .ZN(new_n3949_));
  NAND2_X1   g02947(.A1(new_n3949_), .A2(\A[324] ), .ZN(new_n3950_));
  INV_X1     g02948(.I(\A[324] ), .ZN(new_n3951_));
  NAND2_X1   g02949(.A1(new_n3951_), .A2(\A[323] ), .ZN(new_n3952_));
  AOI21_X1   g02950(.A1(new_n3950_), .A2(new_n3952_), .B(new_n3948_), .ZN(new_n3953_));
  NAND2_X1   g02951(.A1(\A[323] ), .A2(\A[324] ), .ZN(new_n3954_));
  OR2_X2     g02952(.A1(\A[323] ), .A2(\A[324] ), .Z(new_n3955_));
  AOI21_X1   g02953(.A1(new_n3955_), .A2(new_n3954_), .B(\A[322] ), .ZN(new_n3956_));
  NOR4_X1    g02954(.A1(new_n3943_), .A2(new_n3947_), .A3(new_n3953_), .A4(new_n3956_), .ZN(new_n3957_));
  NOR2_X1    g02955(.A1(new_n3941_), .A2(\A[320] ), .ZN(new_n3958_));
  NOR2_X1    g02956(.A1(new_n3939_), .A2(\A[321] ), .ZN(new_n3959_));
  OAI21_X1   g02957(.A1(new_n3958_), .A2(new_n3959_), .B(\A[319] ), .ZN(new_n3960_));
  INV_X1     g02958(.I(new_n3944_), .ZN(new_n3961_));
  OAI21_X1   g02959(.A1(new_n3961_), .A2(new_n3945_), .B(new_n3938_), .ZN(new_n3962_));
  NOR2_X1    g02960(.A1(new_n3951_), .A2(\A[323] ), .ZN(new_n3963_));
  NOR2_X1    g02961(.A1(new_n3949_), .A2(\A[324] ), .ZN(new_n3964_));
  OAI21_X1   g02962(.A1(new_n3963_), .A2(new_n3964_), .B(\A[322] ), .ZN(new_n3965_));
  INV_X1     g02963(.I(new_n3954_), .ZN(new_n3966_));
  NOR2_X1    g02964(.A1(\A[323] ), .A2(\A[324] ), .ZN(new_n3967_));
  OAI21_X1   g02965(.A1(new_n3966_), .A2(new_n3967_), .B(new_n3948_), .ZN(new_n3968_));
  AOI22_X1   g02966(.A1(new_n3960_), .A2(new_n3962_), .B1(new_n3965_), .B2(new_n3968_), .ZN(new_n3969_));
  NOR2_X1    g02967(.A1(new_n3969_), .A2(new_n3957_), .ZN(new_n3970_));
  NAND2_X1   g02968(.A1(new_n3970_), .A2(new_n3937_), .ZN(new_n3971_));
  NOR4_X1    g02969(.A1(new_n3927_), .A2(new_n3929_), .A3(new_n3935_), .A4(new_n3932_), .ZN(new_n3972_));
  AOI22_X1   g02970(.A1(new_n3909_), .A2(new_n3914_), .B1(new_n3919_), .B2(new_n3923_), .ZN(new_n3973_));
  NOR2_X1    g02971(.A1(new_n3972_), .A2(new_n3973_), .ZN(new_n3974_));
  NAND4_X1   g02972(.A1(new_n3960_), .A2(new_n3962_), .A3(new_n3965_), .A4(new_n3968_), .ZN(new_n3975_));
  OAI22_X1   g02973(.A1(new_n3943_), .A2(new_n3947_), .B1(new_n3953_), .B2(new_n3956_), .ZN(new_n3976_));
  NAND2_X1   g02974(.A1(new_n3975_), .A2(new_n3976_), .ZN(new_n3977_));
  NAND2_X1   g02975(.A1(new_n3974_), .A2(new_n3977_), .ZN(new_n3978_));
  NAND2_X1   g02976(.A1(new_n3978_), .A2(new_n3971_), .ZN(new_n3979_));
  INV_X1     g02977(.I(\A[331] ), .ZN(new_n3980_));
  INV_X1     g02978(.I(\A[332] ), .ZN(new_n3981_));
  NAND2_X1   g02979(.A1(new_n3981_), .A2(\A[333] ), .ZN(new_n3982_));
  INV_X1     g02980(.I(\A[333] ), .ZN(new_n3983_));
  NAND2_X1   g02981(.A1(new_n3983_), .A2(\A[332] ), .ZN(new_n3984_));
  AOI21_X1   g02982(.A1(new_n3982_), .A2(new_n3984_), .B(new_n3980_), .ZN(new_n3985_));
  NAND2_X1   g02983(.A1(\A[332] ), .A2(\A[333] ), .ZN(new_n3986_));
  NOR2_X1    g02984(.A1(\A[332] ), .A2(\A[333] ), .ZN(new_n3987_));
  INV_X1     g02985(.I(new_n3987_), .ZN(new_n3988_));
  AOI21_X1   g02986(.A1(new_n3988_), .A2(new_n3986_), .B(\A[331] ), .ZN(new_n3989_));
  INV_X1     g02987(.I(\A[334] ), .ZN(new_n3990_));
  INV_X1     g02988(.I(\A[335] ), .ZN(new_n3991_));
  NAND2_X1   g02989(.A1(new_n3991_), .A2(\A[336] ), .ZN(new_n3992_));
  INV_X1     g02990(.I(\A[336] ), .ZN(new_n3993_));
  NAND2_X1   g02991(.A1(new_n3993_), .A2(\A[335] ), .ZN(new_n3994_));
  AOI21_X1   g02992(.A1(new_n3992_), .A2(new_n3994_), .B(new_n3990_), .ZN(new_n3995_));
  NAND2_X1   g02993(.A1(\A[335] ), .A2(\A[336] ), .ZN(new_n3996_));
  NOR2_X1    g02994(.A1(\A[335] ), .A2(\A[336] ), .ZN(new_n3997_));
  INV_X1     g02995(.I(new_n3997_), .ZN(new_n3998_));
  AOI21_X1   g02996(.A1(new_n3998_), .A2(new_n3996_), .B(\A[334] ), .ZN(new_n3999_));
  NOR4_X1    g02997(.A1(new_n3985_), .A2(new_n3989_), .A3(new_n3999_), .A4(new_n3995_), .ZN(new_n4000_));
  NOR2_X1    g02998(.A1(new_n3983_), .A2(\A[332] ), .ZN(new_n4001_));
  NOR2_X1    g02999(.A1(new_n3981_), .A2(\A[333] ), .ZN(new_n4002_));
  OAI21_X1   g03000(.A1(new_n4001_), .A2(new_n4002_), .B(\A[331] ), .ZN(new_n4003_));
  INV_X1     g03001(.I(new_n3986_), .ZN(new_n4004_));
  OAI21_X1   g03002(.A1(new_n4004_), .A2(new_n3987_), .B(new_n3980_), .ZN(new_n4005_));
  NOR2_X1    g03003(.A1(new_n3993_), .A2(\A[335] ), .ZN(new_n4006_));
  NOR2_X1    g03004(.A1(new_n3991_), .A2(\A[336] ), .ZN(new_n4007_));
  OAI21_X1   g03005(.A1(new_n4006_), .A2(new_n4007_), .B(\A[334] ), .ZN(new_n4008_));
  AND2_X2    g03006(.A1(\A[335] ), .A2(\A[336] ), .Z(new_n4009_));
  OAI21_X1   g03007(.A1(new_n4009_), .A2(new_n3997_), .B(new_n3990_), .ZN(new_n4010_));
  AOI22_X1   g03008(.A1(new_n4003_), .A2(new_n4005_), .B1(new_n4008_), .B2(new_n4010_), .ZN(new_n4011_));
  INV_X1     g03009(.I(\A[337] ), .ZN(new_n4012_));
  INV_X1     g03010(.I(\A[338] ), .ZN(new_n4013_));
  NAND2_X1   g03011(.A1(new_n4013_), .A2(\A[339] ), .ZN(new_n4014_));
  INV_X1     g03012(.I(\A[339] ), .ZN(new_n4015_));
  NAND2_X1   g03013(.A1(new_n4015_), .A2(\A[338] ), .ZN(new_n4016_));
  AOI21_X1   g03014(.A1(new_n4014_), .A2(new_n4016_), .B(new_n4012_), .ZN(new_n4017_));
  NAND2_X1   g03015(.A1(\A[338] ), .A2(\A[339] ), .ZN(new_n4018_));
  NOR2_X1    g03016(.A1(\A[338] ), .A2(\A[339] ), .ZN(new_n4019_));
  INV_X1     g03017(.I(new_n4019_), .ZN(new_n4020_));
  AOI21_X1   g03018(.A1(new_n4020_), .A2(new_n4018_), .B(\A[337] ), .ZN(new_n4021_));
  INV_X1     g03019(.I(\A[340] ), .ZN(new_n4022_));
  INV_X1     g03020(.I(\A[341] ), .ZN(new_n4023_));
  NAND2_X1   g03021(.A1(new_n4023_), .A2(\A[342] ), .ZN(new_n4024_));
  INV_X1     g03022(.I(\A[342] ), .ZN(new_n4025_));
  NAND2_X1   g03023(.A1(new_n4025_), .A2(\A[341] ), .ZN(new_n4026_));
  AOI21_X1   g03024(.A1(new_n4024_), .A2(new_n4026_), .B(new_n4022_), .ZN(new_n4027_));
  NAND2_X1   g03025(.A1(\A[341] ), .A2(\A[342] ), .ZN(new_n4028_));
  NOR2_X1    g03026(.A1(\A[341] ), .A2(\A[342] ), .ZN(new_n4029_));
  INV_X1     g03027(.I(new_n4029_), .ZN(new_n4030_));
  AOI21_X1   g03028(.A1(new_n4030_), .A2(new_n4028_), .B(\A[340] ), .ZN(new_n4031_));
  NOR4_X1    g03029(.A1(new_n4017_), .A2(new_n4021_), .A3(new_n4031_), .A4(new_n4027_), .ZN(new_n4032_));
  NOR2_X1    g03030(.A1(new_n4015_), .A2(\A[338] ), .ZN(new_n4033_));
  NOR2_X1    g03031(.A1(new_n4013_), .A2(\A[339] ), .ZN(new_n4034_));
  OAI21_X1   g03032(.A1(new_n4033_), .A2(new_n4034_), .B(\A[337] ), .ZN(new_n4035_));
  INV_X1     g03033(.I(new_n4018_), .ZN(new_n4036_));
  OAI21_X1   g03034(.A1(new_n4036_), .A2(new_n4019_), .B(new_n4012_), .ZN(new_n4037_));
  NOR2_X1    g03035(.A1(new_n4025_), .A2(\A[341] ), .ZN(new_n4038_));
  NOR2_X1    g03036(.A1(new_n4023_), .A2(\A[342] ), .ZN(new_n4039_));
  OAI21_X1   g03037(.A1(new_n4038_), .A2(new_n4039_), .B(\A[340] ), .ZN(new_n4040_));
  AND2_X2    g03038(.A1(\A[341] ), .A2(\A[342] ), .Z(new_n4041_));
  OAI21_X1   g03039(.A1(new_n4041_), .A2(new_n4029_), .B(new_n4022_), .ZN(new_n4042_));
  AOI22_X1   g03040(.A1(new_n4035_), .A2(new_n4037_), .B1(new_n4040_), .B2(new_n4042_), .ZN(new_n4043_));
  OAI22_X1   g03041(.A1(new_n4000_), .A2(new_n4011_), .B1(new_n4032_), .B2(new_n4043_), .ZN(new_n4044_));
  NAND4_X1   g03042(.A1(new_n4003_), .A2(new_n4008_), .A3(new_n4005_), .A4(new_n4010_), .ZN(new_n4045_));
  OAI22_X1   g03043(.A1(new_n3985_), .A2(new_n3989_), .B1(new_n3999_), .B2(new_n3995_), .ZN(new_n4046_));
  NAND4_X1   g03044(.A1(new_n4035_), .A2(new_n4040_), .A3(new_n4037_), .A4(new_n4042_), .ZN(new_n4047_));
  OAI22_X1   g03045(.A1(new_n4017_), .A2(new_n4021_), .B1(new_n4031_), .B2(new_n4027_), .ZN(new_n4048_));
  NAND4_X1   g03046(.A1(new_n4046_), .A2(new_n4048_), .A3(new_n4045_), .A4(new_n4047_), .ZN(new_n4049_));
  NAND2_X1   g03047(.A1(new_n4044_), .A2(new_n4049_), .ZN(new_n4050_));
  INV_X1     g03048(.I(new_n4050_), .ZN(new_n4051_));
  NOR2_X1    g03049(.A1(new_n4051_), .A2(new_n3979_), .ZN(new_n4052_));
  AOI21_X1   g03050(.A1(new_n3971_), .A2(new_n3978_), .B(new_n4050_), .ZN(new_n4053_));
  NOR2_X1    g03051(.A1(new_n4052_), .A2(new_n4053_), .ZN(new_n4054_));
  NAND2_X1   g03052(.A1(new_n3904_), .A2(new_n4054_), .ZN(new_n4055_));
  NOR2_X1    g03053(.A1(new_n3904_), .A2(new_n4054_), .ZN(new_n4056_));
  INV_X1     g03054(.I(new_n4056_), .ZN(new_n4057_));
  INV_X1     g03055(.I(\A[315] ), .ZN(new_n4058_));
  NOR2_X1    g03056(.A1(new_n4058_), .A2(\A[314] ), .ZN(new_n4059_));
  INV_X1     g03057(.I(\A[314] ), .ZN(new_n4060_));
  NOR2_X1    g03058(.A1(new_n4060_), .A2(\A[315] ), .ZN(new_n4061_));
  OAI21_X1   g03059(.A1(new_n4059_), .A2(new_n4061_), .B(\A[313] ), .ZN(new_n4062_));
  INV_X1     g03060(.I(\A[313] ), .ZN(new_n4063_));
  NOR2_X1    g03061(.A1(\A[314] ), .A2(\A[315] ), .ZN(new_n4064_));
  NAND2_X1   g03062(.A1(\A[314] ), .A2(\A[315] ), .ZN(new_n4065_));
  INV_X1     g03063(.I(new_n4065_), .ZN(new_n4066_));
  OAI21_X1   g03064(.A1(new_n4066_), .A2(new_n4064_), .B(new_n4063_), .ZN(new_n4067_));
  INV_X1     g03065(.I(\A[318] ), .ZN(new_n4068_));
  NOR2_X1    g03066(.A1(new_n4068_), .A2(\A[317] ), .ZN(new_n4069_));
  INV_X1     g03067(.I(\A[317] ), .ZN(new_n4070_));
  NOR2_X1    g03068(.A1(new_n4070_), .A2(\A[318] ), .ZN(new_n4071_));
  OAI21_X1   g03069(.A1(new_n4069_), .A2(new_n4071_), .B(\A[316] ), .ZN(new_n4072_));
  INV_X1     g03070(.I(\A[316] ), .ZN(new_n4073_));
  NOR2_X1    g03071(.A1(\A[317] ), .A2(\A[318] ), .ZN(new_n4074_));
  NAND2_X1   g03072(.A1(\A[317] ), .A2(\A[318] ), .ZN(new_n4075_));
  INV_X1     g03073(.I(new_n4075_), .ZN(new_n4076_));
  OAI21_X1   g03074(.A1(new_n4076_), .A2(new_n4074_), .B(new_n4073_), .ZN(new_n4077_));
  NAND4_X1   g03075(.A1(new_n4062_), .A2(new_n4067_), .A3(new_n4072_), .A4(new_n4077_), .ZN(new_n4078_));
  NAND2_X1   g03076(.A1(new_n4060_), .A2(\A[315] ), .ZN(new_n4079_));
  NAND2_X1   g03077(.A1(new_n4058_), .A2(\A[314] ), .ZN(new_n4080_));
  AOI21_X1   g03078(.A1(new_n4079_), .A2(new_n4080_), .B(new_n4063_), .ZN(new_n4081_));
  INV_X1     g03079(.I(new_n4064_), .ZN(new_n4082_));
  AOI21_X1   g03080(.A1(new_n4082_), .A2(new_n4065_), .B(\A[313] ), .ZN(new_n4083_));
  NAND2_X1   g03081(.A1(new_n4070_), .A2(\A[318] ), .ZN(new_n4084_));
  NAND2_X1   g03082(.A1(new_n4068_), .A2(\A[317] ), .ZN(new_n4085_));
  AOI21_X1   g03083(.A1(new_n4084_), .A2(new_n4085_), .B(new_n4073_), .ZN(new_n4086_));
  INV_X1     g03084(.I(new_n4074_), .ZN(new_n4087_));
  AOI21_X1   g03085(.A1(new_n4087_), .A2(new_n4075_), .B(\A[316] ), .ZN(new_n4088_));
  OAI22_X1   g03086(.A1(new_n4081_), .A2(new_n4083_), .B1(new_n4088_), .B2(new_n4086_), .ZN(new_n4089_));
  NAND2_X1   g03087(.A1(new_n4089_), .A2(new_n4078_), .ZN(new_n4090_));
  INV_X1     g03088(.I(\A[307] ), .ZN(new_n4091_));
  INV_X1     g03089(.I(\A[308] ), .ZN(new_n4092_));
  NAND2_X1   g03090(.A1(new_n4092_), .A2(\A[309] ), .ZN(new_n4093_));
  INV_X1     g03091(.I(\A[309] ), .ZN(new_n4094_));
  NAND2_X1   g03092(.A1(new_n4094_), .A2(\A[308] ), .ZN(new_n4095_));
  AOI21_X1   g03093(.A1(new_n4093_), .A2(new_n4095_), .B(new_n4091_), .ZN(new_n4096_));
  NAND2_X1   g03094(.A1(\A[308] ), .A2(\A[309] ), .ZN(new_n4097_));
  NOR2_X1    g03095(.A1(\A[308] ), .A2(\A[309] ), .ZN(new_n4098_));
  INV_X1     g03096(.I(new_n4098_), .ZN(new_n4099_));
  AOI21_X1   g03097(.A1(new_n4099_), .A2(new_n4097_), .B(\A[307] ), .ZN(new_n4100_));
  INV_X1     g03098(.I(\A[310] ), .ZN(new_n4101_));
  INV_X1     g03099(.I(\A[311] ), .ZN(new_n4102_));
  NAND2_X1   g03100(.A1(new_n4102_), .A2(\A[312] ), .ZN(new_n4103_));
  INV_X1     g03101(.I(\A[312] ), .ZN(new_n4104_));
  NAND2_X1   g03102(.A1(new_n4104_), .A2(\A[311] ), .ZN(new_n4105_));
  AOI21_X1   g03103(.A1(new_n4103_), .A2(new_n4105_), .B(new_n4101_), .ZN(new_n4106_));
  NAND2_X1   g03104(.A1(\A[311] ), .A2(\A[312] ), .ZN(new_n4107_));
  OR2_X2     g03105(.A1(\A[311] ), .A2(\A[312] ), .Z(new_n4108_));
  AOI21_X1   g03106(.A1(new_n4108_), .A2(new_n4107_), .B(\A[310] ), .ZN(new_n4109_));
  NOR4_X1    g03107(.A1(new_n4096_), .A2(new_n4100_), .A3(new_n4106_), .A4(new_n4109_), .ZN(new_n4110_));
  NOR2_X1    g03108(.A1(new_n4094_), .A2(\A[308] ), .ZN(new_n4111_));
  NOR2_X1    g03109(.A1(new_n4092_), .A2(\A[309] ), .ZN(new_n4112_));
  OAI21_X1   g03110(.A1(new_n4111_), .A2(new_n4112_), .B(\A[307] ), .ZN(new_n4113_));
  INV_X1     g03111(.I(new_n4097_), .ZN(new_n4114_));
  OAI21_X1   g03112(.A1(new_n4114_), .A2(new_n4098_), .B(new_n4091_), .ZN(new_n4115_));
  NOR2_X1    g03113(.A1(new_n4104_), .A2(\A[311] ), .ZN(new_n4116_));
  NOR2_X1    g03114(.A1(new_n4102_), .A2(\A[312] ), .ZN(new_n4117_));
  OAI21_X1   g03115(.A1(new_n4116_), .A2(new_n4117_), .B(\A[310] ), .ZN(new_n4118_));
  INV_X1     g03116(.I(new_n4107_), .ZN(new_n4119_));
  NOR2_X1    g03117(.A1(\A[311] ), .A2(\A[312] ), .ZN(new_n4120_));
  OAI21_X1   g03118(.A1(new_n4119_), .A2(new_n4120_), .B(new_n4101_), .ZN(new_n4121_));
  AOI22_X1   g03119(.A1(new_n4113_), .A2(new_n4115_), .B1(new_n4118_), .B2(new_n4121_), .ZN(new_n4122_));
  NOR2_X1    g03120(.A1(new_n4122_), .A2(new_n4110_), .ZN(new_n4123_));
  NOR2_X1    g03121(.A1(new_n4090_), .A2(new_n4123_), .ZN(new_n4124_));
  NOR4_X1    g03122(.A1(new_n4081_), .A2(new_n4083_), .A3(new_n4088_), .A4(new_n4086_), .ZN(new_n4125_));
  AOI22_X1   g03123(.A1(new_n4062_), .A2(new_n4067_), .B1(new_n4072_), .B2(new_n4077_), .ZN(new_n4126_));
  NOR2_X1    g03124(.A1(new_n4126_), .A2(new_n4125_), .ZN(new_n4127_));
  NAND4_X1   g03125(.A1(new_n4113_), .A2(new_n4115_), .A3(new_n4118_), .A4(new_n4121_), .ZN(new_n4128_));
  OAI22_X1   g03126(.A1(new_n4096_), .A2(new_n4100_), .B1(new_n4106_), .B2(new_n4109_), .ZN(new_n4129_));
  NAND2_X1   g03127(.A1(new_n4128_), .A2(new_n4129_), .ZN(new_n4130_));
  NOR2_X1    g03128(.A1(new_n4127_), .A2(new_n4130_), .ZN(new_n4131_));
  INV_X1     g03129(.I(\A[303] ), .ZN(new_n4132_));
  NOR2_X1    g03130(.A1(new_n4132_), .A2(\A[302] ), .ZN(new_n4133_));
  INV_X1     g03131(.I(\A[302] ), .ZN(new_n4134_));
  NOR2_X1    g03132(.A1(new_n4134_), .A2(\A[303] ), .ZN(new_n4135_));
  OAI21_X1   g03133(.A1(new_n4133_), .A2(new_n4135_), .B(\A[301] ), .ZN(new_n4136_));
  INV_X1     g03134(.I(\A[301] ), .ZN(new_n4137_));
  NOR2_X1    g03135(.A1(\A[302] ), .A2(\A[303] ), .ZN(new_n4138_));
  NAND2_X1   g03136(.A1(\A[302] ), .A2(\A[303] ), .ZN(new_n4139_));
  INV_X1     g03137(.I(new_n4139_), .ZN(new_n4140_));
  OAI21_X1   g03138(.A1(new_n4140_), .A2(new_n4138_), .B(new_n4137_), .ZN(new_n4141_));
  INV_X1     g03139(.I(\A[306] ), .ZN(new_n4142_));
  NOR2_X1    g03140(.A1(new_n4142_), .A2(\A[305] ), .ZN(new_n4143_));
  INV_X1     g03141(.I(\A[305] ), .ZN(new_n4144_));
  NOR2_X1    g03142(.A1(new_n4144_), .A2(\A[306] ), .ZN(new_n4145_));
  OAI21_X1   g03143(.A1(new_n4143_), .A2(new_n4145_), .B(\A[304] ), .ZN(new_n4146_));
  INV_X1     g03144(.I(\A[304] ), .ZN(new_n4147_));
  NOR2_X1    g03145(.A1(\A[305] ), .A2(\A[306] ), .ZN(new_n4148_));
  AND2_X2    g03146(.A1(\A[305] ), .A2(\A[306] ), .Z(new_n4149_));
  OAI21_X1   g03147(.A1(new_n4149_), .A2(new_n4148_), .B(new_n4147_), .ZN(new_n4150_));
  NAND4_X1   g03148(.A1(new_n4136_), .A2(new_n4146_), .A3(new_n4141_), .A4(new_n4150_), .ZN(new_n4151_));
  NAND2_X1   g03149(.A1(new_n4134_), .A2(\A[303] ), .ZN(new_n4152_));
  NAND2_X1   g03150(.A1(new_n4132_), .A2(\A[302] ), .ZN(new_n4153_));
  AOI21_X1   g03151(.A1(new_n4152_), .A2(new_n4153_), .B(new_n4137_), .ZN(new_n4154_));
  INV_X1     g03152(.I(new_n4138_), .ZN(new_n4155_));
  AOI21_X1   g03153(.A1(new_n4155_), .A2(new_n4139_), .B(\A[301] ), .ZN(new_n4156_));
  NAND2_X1   g03154(.A1(new_n4144_), .A2(\A[306] ), .ZN(new_n4157_));
  NAND2_X1   g03155(.A1(new_n4142_), .A2(\A[305] ), .ZN(new_n4158_));
  AOI21_X1   g03156(.A1(new_n4157_), .A2(new_n4158_), .B(new_n4147_), .ZN(new_n4159_));
  INV_X1     g03157(.I(new_n4148_), .ZN(new_n4160_));
  NAND2_X1   g03158(.A1(\A[305] ), .A2(\A[306] ), .ZN(new_n4161_));
  AOI21_X1   g03159(.A1(new_n4160_), .A2(new_n4161_), .B(\A[304] ), .ZN(new_n4162_));
  OAI22_X1   g03160(.A1(new_n4154_), .A2(new_n4156_), .B1(new_n4162_), .B2(new_n4159_), .ZN(new_n4163_));
  NAND2_X1   g03161(.A1(new_n4163_), .A2(new_n4151_), .ZN(new_n4164_));
  INV_X1     g03162(.I(\A[295] ), .ZN(new_n4165_));
  INV_X1     g03163(.I(\A[296] ), .ZN(new_n4166_));
  NAND2_X1   g03164(.A1(new_n4166_), .A2(\A[297] ), .ZN(new_n4167_));
  INV_X1     g03165(.I(\A[297] ), .ZN(new_n4168_));
  NAND2_X1   g03166(.A1(new_n4168_), .A2(\A[296] ), .ZN(new_n4169_));
  AOI21_X1   g03167(.A1(new_n4167_), .A2(new_n4169_), .B(new_n4165_), .ZN(new_n4170_));
  NAND2_X1   g03168(.A1(\A[296] ), .A2(\A[297] ), .ZN(new_n4171_));
  NOR2_X1    g03169(.A1(\A[296] ), .A2(\A[297] ), .ZN(new_n4172_));
  INV_X1     g03170(.I(new_n4172_), .ZN(new_n4173_));
  AOI21_X1   g03171(.A1(new_n4173_), .A2(new_n4171_), .B(\A[295] ), .ZN(new_n4174_));
  INV_X1     g03172(.I(\A[298] ), .ZN(new_n4175_));
  INV_X1     g03173(.I(\A[299] ), .ZN(new_n4176_));
  NAND2_X1   g03174(.A1(new_n4176_), .A2(\A[300] ), .ZN(new_n4177_));
  INV_X1     g03175(.I(\A[300] ), .ZN(new_n4178_));
  NAND2_X1   g03176(.A1(new_n4178_), .A2(\A[299] ), .ZN(new_n4179_));
  AOI21_X1   g03177(.A1(new_n4177_), .A2(new_n4179_), .B(new_n4175_), .ZN(new_n4180_));
  NAND2_X1   g03178(.A1(\A[299] ), .A2(\A[300] ), .ZN(new_n4181_));
  OR2_X2     g03179(.A1(\A[299] ), .A2(\A[300] ), .Z(new_n4182_));
  AOI21_X1   g03180(.A1(new_n4182_), .A2(new_n4181_), .B(\A[298] ), .ZN(new_n4183_));
  NOR4_X1    g03181(.A1(new_n4170_), .A2(new_n4174_), .A3(new_n4180_), .A4(new_n4183_), .ZN(new_n4184_));
  NOR2_X1    g03182(.A1(new_n4168_), .A2(\A[296] ), .ZN(new_n4185_));
  NOR2_X1    g03183(.A1(new_n4166_), .A2(\A[297] ), .ZN(new_n4186_));
  OAI21_X1   g03184(.A1(new_n4185_), .A2(new_n4186_), .B(\A[295] ), .ZN(new_n4187_));
  INV_X1     g03185(.I(new_n4171_), .ZN(new_n4188_));
  OAI21_X1   g03186(.A1(new_n4188_), .A2(new_n4172_), .B(new_n4165_), .ZN(new_n4189_));
  NOR2_X1    g03187(.A1(new_n4178_), .A2(\A[299] ), .ZN(new_n4190_));
  NOR2_X1    g03188(.A1(new_n4176_), .A2(\A[300] ), .ZN(new_n4191_));
  OAI21_X1   g03189(.A1(new_n4190_), .A2(new_n4191_), .B(\A[298] ), .ZN(new_n4192_));
  INV_X1     g03190(.I(new_n4181_), .ZN(new_n4193_));
  NOR2_X1    g03191(.A1(\A[299] ), .A2(\A[300] ), .ZN(new_n4194_));
  OAI21_X1   g03192(.A1(new_n4193_), .A2(new_n4194_), .B(new_n4175_), .ZN(new_n4195_));
  AOI22_X1   g03193(.A1(new_n4187_), .A2(new_n4189_), .B1(new_n4192_), .B2(new_n4195_), .ZN(new_n4196_));
  NOR2_X1    g03194(.A1(new_n4196_), .A2(new_n4184_), .ZN(new_n4197_));
  NOR2_X1    g03195(.A1(new_n4197_), .A2(new_n4164_), .ZN(new_n4198_));
  NOR4_X1    g03196(.A1(new_n4154_), .A2(new_n4156_), .A3(new_n4162_), .A4(new_n4159_), .ZN(new_n4199_));
  AOI22_X1   g03197(.A1(new_n4136_), .A2(new_n4141_), .B1(new_n4146_), .B2(new_n4150_), .ZN(new_n4200_));
  NOR2_X1    g03198(.A1(new_n4199_), .A2(new_n4200_), .ZN(new_n4201_));
  NAND4_X1   g03199(.A1(new_n4187_), .A2(new_n4189_), .A3(new_n4192_), .A4(new_n4195_), .ZN(new_n4202_));
  OAI22_X1   g03200(.A1(new_n4170_), .A2(new_n4174_), .B1(new_n4180_), .B2(new_n4183_), .ZN(new_n4203_));
  NAND2_X1   g03201(.A1(new_n4202_), .A2(new_n4203_), .ZN(new_n4204_));
  NOR2_X1    g03202(.A1(new_n4201_), .A2(new_n4204_), .ZN(new_n4205_));
  OAI22_X1   g03203(.A1(new_n4124_), .A2(new_n4131_), .B1(new_n4205_), .B2(new_n4198_), .ZN(new_n4206_));
  NOR2_X1    g03204(.A1(new_n4124_), .A2(new_n4131_), .ZN(new_n4207_));
  NAND2_X1   g03205(.A1(new_n4201_), .A2(new_n4204_), .ZN(new_n4208_));
  NAND2_X1   g03206(.A1(new_n4197_), .A2(new_n4164_), .ZN(new_n4209_));
  NAND3_X1   g03207(.A1(new_n4207_), .A2(new_n4208_), .A3(new_n4209_), .ZN(new_n4210_));
  NAND2_X1   g03208(.A1(new_n4210_), .A2(new_n4206_), .ZN(new_n4211_));
  INV_X1     g03209(.I(\A[291] ), .ZN(new_n4212_));
  NOR2_X1    g03210(.A1(new_n4212_), .A2(\A[290] ), .ZN(new_n4213_));
  NAND2_X1   g03211(.A1(new_n4212_), .A2(\A[290] ), .ZN(new_n4214_));
  INV_X1     g03212(.I(new_n4214_), .ZN(new_n4215_));
  OAI21_X1   g03213(.A1(new_n4215_), .A2(new_n4213_), .B(\A[289] ), .ZN(new_n4216_));
  INV_X1     g03214(.I(\A[289] ), .ZN(new_n4217_));
  NOR2_X1    g03215(.A1(\A[290] ), .A2(\A[291] ), .ZN(new_n4218_));
  NAND2_X1   g03216(.A1(\A[290] ), .A2(\A[291] ), .ZN(new_n4219_));
  INV_X1     g03217(.I(new_n4219_), .ZN(new_n4220_));
  OAI21_X1   g03218(.A1(new_n4220_), .A2(new_n4218_), .B(new_n4217_), .ZN(new_n4221_));
  INV_X1     g03219(.I(\A[294] ), .ZN(new_n4222_));
  NOR2_X1    g03220(.A1(new_n4222_), .A2(\A[293] ), .ZN(new_n4223_));
  INV_X1     g03221(.I(\A[293] ), .ZN(new_n4224_));
  NOR2_X1    g03222(.A1(new_n4224_), .A2(\A[294] ), .ZN(new_n4225_));
  OAI21_X1   g03223(.A1(new_n4223_), .A2(new_n4225_), .B(\A[292] ), .ZN(new_n4226_));
  INV_X1     g03224(.I(\A[292] ), .ZN(new_n4227_));
  NOR2_X1    g03225(.A1(\A[293] ), .A2(\A[294] ), .ZN(new_n4228_));
  NAND2_X1   g03226(.A1(\A[293] ), .A2(\A[294] ), .ZN(new_n4229_));
  INV_X1     g03227(.I(new_n4229_), .ZN(new_n4230_));
  OAI21_X1   g03228(.A1(new_n4230_), .A2(new_n4228_), .B(new_n4227_), .ZN(new_n4231_));
  NAND4_X1   g03229(.A1(new_n4216_), .A2(new_n4221_), .A3(new_n4231_), .A4(new_n4226_), .ZN(new_n4232_));
  INV_X1     g03230(.I(new_n4213_), .ZN(new_n4233_));
  AOI21_X1   g03231(.A1(new_n4233_), .A2(new_n4214_), .B(new_n4217_), .ZN(new_n4234_));
  INV_X1     g03232(.I(new_n4218_), .ZN(new_n4235_));
  AOI21_X1   g03233(.A1(new_n4235_), .A2(new_n4219_), .B(\A[289] ), .ZN(new_n4236_));
  NAND2_X1   g03234(.A1(new_n4224_), .A2(\A[294] ), .ZN(new_n4237_));
  NAND2_X1   g03235(.A1(new_n4222_), .A2(\A[293] ), .ZN(new_n4238_));
  AOI21_X1   g03236(.A1(new_n4237_), .A2(new_n4238_), .B(new_n4227_), .ZN(new_n4239_));
  INV_X1     g03237(.I(new_n4228_), .ZN(new_n4240_));
  AOI21_X1   g03238(.A1(new_n4240_), .A2(new_n4229_), .B(\A[292] ), .ZN(new_n4241_));
  OAI22_X1   g03239(.A1(new_n4234_), .A2(new_n4236_), .B1(new_n4241_), .B2(new_n4239_), .ZN(new_n4242_));
  NAND2_X1   g03240(.A1(new_n4242_), .A2(new_n4232_), .ZN(new_n4243_));
  INV_X1     g03241(.I(\A[283] ), .ZN(new_n4244_));
  INV_X1     g03242(.I(\A[284] ), .ZN(new_n4245_));
  NAND2_X1   g03243(.A1(new_n4245_), .A2(\A[285] ), .ZN(new_n4246_));
  INV_X1     g03244(.I(\A[285] ), .ZN(new_n4247_));
  NAND2_X1   g03245(.A1(new_n4247_), .A2(\A[284] ), .ZN(new_n4248_));
  AOI21_X1   g03246(.A1(new_n4246_), .A2(new_n4248_), .B(new_n4244_), .ZN(new_n4249_));
  NAND2_X1   g03247(.A1(\A[284] ), .A2(\A[285] ), .ZN(new_n4250_));
  NOR2_X1    g03248(.A1(\A[284] ), .A2(\A[285] ), .ZN(new_n4251_));
  INV_X1     g03249(.I(new_n4251_), .ZN(new_n4252_));
  AOI21_X1   g03250(.A1(new_n4252_), .A2(new_n4250_), .B(\A[283] ), .ZN(new_n4253_));
  INV_X1     g03251(.I(\A[286] ), .ZN(new_n4254_));
  INV_X1     g03252(.I(\A[287] ), .ZN(new_n4255_));
  NAND2_X1   g03253(.A1(new_n4255_), .A2(\A[288] ), .ZN(new_n4256_));
  INV_X1     g03254(.I(\A[288] ), .ZN(new_n4257_));
  NAND2_X1   g03255(.A1(new_n4257_), .A2(\A[287] ), .ZN(new_n4258_));
  AOI21_X1   g03256(.A1(new_n4256_), .A2(new_n4258_), .B(new_n4254_), .ZN(new_n4259_));
  NAND2_X1   g03257(.A1(\A[287] ), .A2(\A[288] ), .ZN(new_n4260_));
  NOR2_X1    g03258(.A1(\A[287] ), .A2(\A[288] ), .ZN(new_n4261_));
  INV_X1     g03259(.I(new_n4261_), .ZN(new_n4262_));
  AOI21_X1   g03260(.A1(new_n4262_), .A2(new_n4260_), .B(\A[286] ), .ZN(new_n4263_));
  NOR4_X1    g03261(.A1(new_n4249_), .A2(new_n4253_), .A3(new_n4263_), .A4(new_n4259_), .ZN(new_n4264_));
  INV_X1     g03262(.I(new_n4246_), .ZN(new_n4265_));
  NOR2_X1    g03263(.A1(new_n4245_), .A2(\A[285] ), .ZN(new_n4266_));
  OAI21_X1   g03264(.A1(new_n4265_), .A2(new_n4266_), .B(\A[283] ), .ZN(new_n4267_));
  INV_X1     g03265(.I(new_n4250_), .ZN(new_n4268_));
  OAI21_X1   g03266(.A1(new_n4268_), .A2(new_n4251_), .B(new_n4244_), .ZN(new_n4269_));
  NOR2_X1    g03267(.A1(new_n4257_), .A2(\A[287] ), .ZN(new_n4270_));
  NOR2_X1    g03268(.A1(new_n4255_), .A2(\A[288] ), .ZN(new_n4271_));
  OAI21_X1   g03269(.A1(new_n4270_), .A2(new_n4271_), .B(\A[286] ), .ZN(new_n4272_));
  INV_X1     g03270(.I(new_n4260_), .ZN(new_n4273_));
  OAI21_X1   g03271(.A1(new_n4273_), .A2(new_n4261_), .B(new_n4254_), .ZN(new_n4274_));
  AOI22_X1   g03272(.A1(new_n4267_), .A2(new_n4269_), .B1(new_n4274_), .B2(new_n4272_), .ZN(new_n4275_));
  NOR2_X1    g03273(.A1(new_n4275_), .A2(new_n4264_), .ZN(new_n4276_));
  NOR2_X1    g03274(.A1(new_n4243_), .A2(new_n4276_), .ZN(new_n4277_));
  NOR4_X1    g03275(.A1(new_n4234_), .A2(new_n4236_), .A3(new_n4241_), .A4(new_n4239_), .ZN(new_n4278_));
  AOI22_X1   g03276(.A1(new_n4216_), .A2(new_n4221_), .B1(new_n4231_), .B2(new_n4226_), .ZN(new_n4279_));
  NOR2_X1    g03277(.A1(new_n4278_), .A2(new_n4279_), .ZN(new_n4280_));
  NAND4_X1   g03278(.A1(new_n4267_), .A2(new_n4269_), .A3(new_n4274_), .A4(new_n4272_), .ZN(new_n4281_));
  OAI22_X1   g03279(.A1(new_n4249_), .A2(new_n4253_), .B1(new_n4263_), .B2(new_n4259_), .ZN(new_n4282_));
  NAND2_X1   g03280(.A1(new_n4281_), .A2(new_n4282_), .ZN(new_n4283_));
  NOR2_X1    g03281(.A1(new_n4280_), .A2(new_n4283_), .ZN(new_n4284_));
  INV_X1     g03282(.I(\A[277] ), .ZN(new_n4285_));
  INV_X1     g03283(.I(\A[278] ), .ZN(new_n4286_));
  NAND2_X1   g03284(.A1(new_n4286_), .A2(\A[279] ), .ZN(new_n4287_));
  INV_X1     g03285(.I(\A[279] ), .ZN(new_n4288_));
  NAND2_X1   g03286(.A1(new_n4288_), .A2(\A[278] ), .ZN(new_n4289_));
  AOI21_X1   g03287(.A1(new_n4287_), .A2(new_n4289_), .B(new_n4285_), .ZN(new_n4290_));
  NOR2_X1    g03288(.A1(\A[278] ), .A2(\A[279] ), .ZN(new_n4291_));
  INV_X1     g03289(.I(new_n4291_), .ZN(new_n4292_));
  NAND2_X1   g03290(.A1(\A[278] ), .A2(\A[279] ), .ZN(new_n4293_));
  AOI21_X1   g03291(.A1(new_n4292_), .A2(new_n4293_), .B(\A[277] ), .ZN(new_n4294_));
  INV_X1     g03292(.I(\A[280] ), .ZN(new_n4295_));
  INV_X1     g03293(.I(\A[281] ), .ZN(new_n4296_));
  NAND2_X1   g03294(.A1(new_n4296_), .A2(\A[282] ), .ZN(new_n4297_));
  INV_X1     g03295(.I(\A[282] ), .ZN(new_n4298_));
  NAND2_X1   g03296(.A1(new_n4298_), .A2(\A[281] ), .ZN(new_n4299_));
  AOI21_X1   g03297(.A1(new_n4297_), .A2(new_n4299_), .B(new_n4295_), .ZN(new_n4300_));
  NOR2_X1    g03298(.A1(\A[281] ), .A2(\A[282] ), .ZN(new_n4301_));
  INV_X1     g03299(.I(new_n4301_), .ZN(new_n4302_));
  NAND2_X1   g03300(.A1(\A[281] ), .A2(\A[282] ), .ZN(new_n4303_));
  AOI21_X1   g03301(.A1(new_n4302_), .A2(new_n4303_), .B(\A[280] ), .ZN(new_n4304_));
  NOR4_X1    g03302(.A1(new_n4290_), .A2(new_n4294_), .A3(new_n4304_), .A4(new_n4300_), .ZN(new_n4305_));
  INV_X1     g03303(.I(new_n4287_), .ZN(new_n4306_));
  NOR2_X1    g03304(.A1(new_n4286_), .A2(\A[279] ), .ZN(new_n4307_));
  OAI21_X1   g03305(.A1(new_n4306_), .A2(new_n4307_), .B(\A[277] ), .ZN(new_n4308_));
  INV_X1     g03306(.I(new_n4293_), .ZN(new_n4309_));
  OAI21_X1   g03307(.A1(new_n4309_), .A2(new_n4291_), .B(new_n4285_), .ZN(new_n4310_));
  NOR2_X1    g03308(.A1(new_n4298_), .A2(\A[281] ), .ZN(new_n4311_));
  NOR2_X1    g03309(.A1(new_n4296_), .A2(\A[282] ), .ZN(new_n4312_));
  OAI21_X1   g03310(.A1(new_n4311_), .A2(new_n4312_), .B(\A[280] ), .ZN(new_n4313_));
  INV_X1     g03311(.I(new_n4303_), .ZN(new_n4314_));
  OAI21_X1   g03312(.A1(new_n4314_), .A2(new_n4301_), .B(new_n4295_), .ZN(new_n4315_));
  AOI22_X1   g03313(.A1(new_n4308_), .A2(new_n4310_), .B1(new_n4315_), .B2(new_n4313_), .ZN(new_n4316_));
  NOR2_X1    g03314(.A1(new_n4316_), .A2(new_n4305_), .ZN(new_n4317_));
  INV_X1     g03315(.I(\A[273] ), .ZN(new_n4318_));
  NOR2_X1    g03316(.A1(new_n4318_), .A2(\A[272] ), .ZN(new_n4319_));
  INV_X1     g03317(.I(\A[272] ), .ZN(new_n4320_));
  NOR2_X1    g03318(.A1(new_n4320_), .A2(\A[273] ), .ZN(new_n4321_));
  OAI21_X1   g03319(.A1(new_n4319_), .A2(new_n4321_), .B(\A[271] ), .ZN(new_n4322_));
  INV_X1     g03320(.I(\A[271] ), .ZN(new_n4323_));
  NAND2_X1   g03321(.A1(\A[272] ), .A2(\A[273] ), .ZN(new_n4324_));
  INV_X1     g03322(.I(new_n4324_), .ZN(new_n4325_));
  NOR2_X1    g03323(.A1(\A[272] ), .A2(\A[273] ), .ZN(new_n4326_));
  OAI21_X1   g03324(.A1(new_n4325_), .A2(new_n4326_), .B(new_n4323_), .ZN(new_n4327_));
  INV_X1     g03325(.I(\A[276] ), .ZN(new_n4328_));
  NOR2_X1    g03326(.A1(new_n4328_), .A2(\A[275] ), .ZN(new_n4329_));
  INV_X1     g03327(.I(\A[275] ), .ZN(new_n4330_));
  NOR2_X1    g03328(.A1(new_n4330_), .A2(\A[276] ), .ZN(new_n4331_));
  OAI21_X1   g03329(.A1(new_n4329_), .A2(new_n4331_), .B(\A[274] ), .ZN(new_n4332_));
  INV_X1     g03330(.I(\A[274] ), .ZN(new_n4333_));
  NAND2_X1   g03331(.A1(\A[275] ), .A2(\A[276] ), .ZN(new_n4334_));
  INV_X1     g03332(.I(new_n4334_), .ZN(new_n4335_));
  NOR2_X1    g03333(.A1(\A[275] ), .A2(\A[276] ), .ZN(new_n4336_));
  OAI21_X1   g03334(.A1(new_n4335_), .A2(new_n4336_), .B(new_n4333_), .ZN(new_n4337_));
  NAND4_X1   g03335(.A1(new_n4322_), .A2(new_n4327_), .A3(new_n4332_), .A4(new_n4337_), .ZN(new_n4338_));
  NAND2_X1   g03336(.A1(new_n4320_), .A2(\A[273] ), .ZN(new_n4339_));
  NAND2_X1   g03337(.A1(new_n4318_), .A2(\A[272] ), .ZN(new_n4340_));
  AOI21_X1   g03338(.A1(new_n4339_), .A2(new_n4340_), .B(new_n4323_), .ZN(new_n4341_));
  INV_X1     g03339(.I(new_n4326_), .ZN(new_n4342_));
  AOI21_X1   g03340(.A1(new_n4342_), .A2(new_n4324_), .B(\A[271] ), .ZN(new_n4343_));
  NAND2_X1   g03341(.A1(new_n4330_), .A2(\A[276] ), .ZN(new_n4344_));
  NAND2_X1   g03342(.A1(new_n4328_), .A2(\A[275] ), .ZN(new_n4345_));
  AOI21_X1   g03343(.A1(new_n4344_), .A2(new_n4345_), .B(new_n4333_), .ZN(new_n4346_));
  INV_X1     g03344(.I(new_n4336_), .ZN(new_n4347_));
  AOI21_X1   g03345(.A1(new_n4347_), .A2(new_n4334_), .B(\A[274] ), .ZN(new_n4348_));
  OAI22_X1   g03346(.A1(new_n4341_), .A2(new_n4343_), .B1(new_n4348_), .B2(new_n4346_), .ZN(new_n4349_));
  NAND2_X1   g03347(.A1(new_n4349_), .A2(new_n4338_), .ZN(new_n4350_));
  NAND2_X1   g03348(.A1(new_n4317_), .A2(new_n4350_), .ZN(new_n4351_));
  INV_X1     g03349(.I(new_n4351_), .ZN(new_n4352_));
  NOR2_X1    g03350(.A1(new_n4317_), .A2(new_n4350_), .ZN(new_n4353_));
  OAI22_X1   g03351(.A1(new_n4352_), .A2(new_n4353_), .B1(new_n4277_), .B2(new_n4284_), .ZN(new_n4354_));
  NOR2_X1    g03352(.A1(new_n4277_), .A2(new_n4284_), .ZN(new_n4355_));
  INV_X1     g03353(.I(new_n4353_), .ZN(new_n4356_));
  NAND3_X1   g03354(.A1(new_n4355_), .A2(new_n4351_), .A3(new_n4356_), .ZN(new_n4357_));
  NAND2_X1   g03355(.A1(new_n4357_), .A2(new_n4354_), .ZN(new_n4358_));
  NOR2_X1    g03356(.A1(new_n4358_), .A2(new_n4211_), .ZN(new_n4359_));
  INV_X1     g03357(.I(new_n4359_), .ZN(new_n4360_));
  NAND2_X1   g03358(.A1(new_n4358_), .A2(new_n4211_), .ZN(new_n4361_));
  NAND4_X1   g03359(.A1(new_n4057_), .A2(new_n4361_), .A3(new_n4055_), .A4(new_n4360_), .ZN(new_n4362_));
  INV_X1     g03360(.I(new_n4055_), .ZN(new_n4363_));
  INV_X1     g03361(.I(new_n4361_), .ZN(new_n4364_));
  OAI22_X1   g03362(.A1(new_n4363_), .A2(new_n4056_), .B1(new_n4359_), .B2(new_n4364_), .ZN(new_n4365_));
  NAND2_X1   g03363(.A1(new_n4365_), .A2(new_n4362_), .ZN(new_n4366_));
  NOR2_X1    g03364(.A1(new_n4366_), .A2(new_n3737_), .ZN(new_n4367_));
  INV_X1     g03365(.I(new_n4367_), .ZN(new_n4368_));
  NAND2_X1   g03366(.A1(new_n4366_), .A2(new_n3737_), .ZN(new_n4369_));
  NOR2_X1    g03367(.A1(new_n3077_), .A2(new_n2067_), .ZN(new_n4370_));
  NOR2_X1    g03368(.A1(new_n2698_), .A2(new_n4370_), .ZN(new_n4371_));
  NAND3_X1   g03369(.A1(new_n4371_), .A2(new_n4368_), .A3(new_n4369_), .ZN(new_n4372_));
  AOI21_X1   g03370(.A1(\A[335] ), .A2(\A[336] ), .B(\A[334] ), .ZN(new_n4373_));
  NOR2_X1    g03371(.A1(new_n4373_), .A2(new_n3997_), .ZN(new_n4374_));
  AOI21_X1   g03372(.A1(\A[332] ), .A2(\A[333] ), .B(\A[331] ), .ZN(new_n4375_));
  NOR2_X1    g03373(.A1(new_n4375_), .A2(new_n3987_), .ZN(new_n4376_));
  NOR2_X1    g03374(.A1(new_n4374_), .A2(new_n4376_), .ZN(new_n4377_));
  NOR4_X1    g03375(.A1(new_n4373_), .A2(new_n4375_), .A3(new_n3987_), .A4(new_n3997_), .ZN(new_n4378_));
  NOR2_X1    g03376(.A1(new_n4377_), .A2(new_n4378_), .ZN(new_n4379_));
  NAND2_X1   g03377(.A1(new_n4045_), .A2(new_n4379_), .ZN(new_n4380_));
  OAI22_X1   g03378(.A1(new_n3987_), .A2(new_n4375_), .B1(new_n4373_), .B2(new_n3997_), .ZN(new_n4381_));
  INV_X1     g03379(.I(new_n4378_), .ZN(new_n4382_));
  NAND2_X1   g03380(.A1(new_n4382_), .A2(new_n4381_), .ZN(new_n4383_));
  NAND2_X1   g03381(.A1(new_n4000_), .A2(new_n4383_), .ZN(new_n4384_));
  NAND2_X1   g03382(.A1(new_n4384_), .A2(new_n4380_), .ZN(new_n4385_));
  NOR4_X1    g03383(.A1(new_n4000_), .A2(new_n4011_), .A3(new_n4032_), .A4(new_n4043_), .ZN(new_n4386_));
  NAND2_X1   g03384(.A1(new_n4035_), .A2(new_n4037_), .ZN(new_n4387_));
  NAND2_X1   g03385(.A1(new_n4040_), .A2(new_n4042_), .ZN(new_n4388_));
  AOI21_X1   g03386(.A1(\A[341] ), .A2(\A[342] ), .B(\A[340] ), .ZN(new_n4389_));
  AOI21_X1   g03387(.A1(\A[338] ), .A2(\A[339] ), .B(\A[337] ), .ZN(new_n4390_));
  NOR2_X1    g03388(.A1(new_n4390_), .A2(new_n4019_), .ZN(new_n4391_));
  NOR3_X1    g03389(.A1(new_n4391_), .A2(new_n4029_), .A3(new_n4389_), .ZN(new_n4392_));
  NOR2_X1    g03390(.A1(new_n4389_), .A2(new_n4029_), .ZN(new_n4393_));
  NOR3_X1    g03391(.A1(new_n4393_), .A2(new_n4019_), .A3(new_n4390_), .ZN(new_n4394_));
  OAI22_X1   g03392(.A1(new_n4387_), .A2(new_n4388_), .B1(new_n4392_), .B2(new_n4394_), .ZN(new_n4395_));
  NOR2_X1    g03393(.A1(new_n4392_), .A2(new_n4394_), .ZN(new_n4396_));
  NAND2_X1   g03394(.A1(new_n4032_), .A2(new_n4396_), .ZN(new_n4397_));
  NAND2_X1   g03395(.A1(new_n4397_), .A2(new_n4395_), .ZN(new_n4398_));
  NOR2_X1    g03396(.A1(new_n4398_), .A2(new_n4386_), .ZN(new_n4399_));
  NOR2_X1    g03397(.A1(new_n4021_), .A2(new_n4017_), .ZN(new_n4400_));
  NOR2_X1    g03398(.A1(new_n4031_), .A2(new_n4027_), .ZN(new_n4401_));
  OAI21_X1   g03399(.A1(new_n4019_), .A2(new_n4390_), .B(new_n4393_), .ZN(new_n4402_));
  OAI21_X1   g03400(.A1(new_n4029_), .A2(new_n4389_), .B(new_n4391_), .ZN(new_n4403_));
  AOI22_X1   g03401(.A1(new_n4400_), .A2(new_n4401_), .B1(new_n4402_), .B2(new_n4403_), .ZN(new_n4404_));
  NOR4_X1    g03402(.A1(new_n4387_), .A2(new_n4388_), .A3(new_n4392_), .A4(new_n4394_), .ZN(new_n4405_));
  NOR2_X1    g03403(.A1(new_n4404_), .A2(new_n4405_), .ZN(new_n4406_));
  NOR2_X1    g03404(.A1(new_n4406_), .A2(new_n4049_), .ZN(new_n4407_));
  NOR3_X1    g03405(.A1(new_n4399_), .A2(new_n4407_), .A3(new_n4385_), .ZN(new_n4408_));
  AND2_X2    g03406(.A1(new_n4384_), .A2(new_n4380_), .Z(new_n4409_));
  NAND2_X1   g03407(.A1(new_n4406_), .A2(new_n4049_), .ZN(new_n4410_));
  NAND2_X1   g03408(.A1(new_n4393_), .A2(new_n4391_), .ZN(new_n4411_));
  INV_X1     g03409(.I(new_n4411_), .ZN(new_n4412_));
  NAND2_X1   g03410(.A1(new_n4048_), .A2(new_n4412_), .ZN(new_n4413_));
  NOR3_X1    g03411(.A1(new_n4396_), .A2(new_n4032_), .A3(new_n4043_), .ZN(new_n4414_));
  NAND4_X1   g03412(.A1(new_n4414_), .A2(new_n4045_), .A3(new_n4413_), .A4(new_n4046_), .ZN(new_n4415_));
  AOI21_X1   g03413(.A1(new_n4410_), .A2(new_n4415_), .B(new_n4409_), .ZN(new_n4416_));
  NOR2_X1    g03414(.A1(new_n4408_), .A2(new_n4416_), .ZN(new_n4417_));
  INV_X1     g03415(.I(new_n3979_), .ZN(new_n4418_));
  AOI21_X1   g03416(.A1(\A[323] ), .A2(\A[324] ), .B(\A[322] ), .ZN(new_n4419_));
  AOI21_X1   g03417(.A1(\A[320] ), .A2(\A[321] ), .B(\A[319] ), .ZN(new_n4420_));
  OAI22_X1   g03418(.A1(new_n3945_), .A2(new_n4420_), .B1(new_n4419_), .B2(new_n3967_), .ZN(new_n4421_));
  NOR2_X1    g03419(.A1(new_n4419_), .A2(new_n3967_), .ZN(new_n4422_));
  NOR2_X1    g03420(.A1(new_n4420_), .A2(new_n3945_), .ZN(new_n4423_));
  NAND2_X1   g03421(.A1(new_n4422_), .A2(new_n4423_), .ZN(new_n4424_));
  NAND2_X1   g03422(.A1(new_n4424_), .A2(new_n4421_), .ZN(new_n4425_));
  NOR2_X1    g03423(.A1(new_n3957_), .A2(new_n4425_), .ZN(new_n4426_));
  NOR2_X1    g03424(.A1(new_n4422_), .A2(new_n4423_), .ZN(new_n4427_));
  NOR4_X1    g03425(.A1(new_n4419_), .A2(new_n4420_), .A3(new_n3945_), .A4(new_n3967_), .ZN(new_n4428_));
  NOR2_X1    g03426(.A1(new_n4427_), .A2(new_n4428_), .ZN(new_n4429_));
  NOR2_X1    g03427(.A1(new_n3975_), .A2(new_n4429_), .ZN(new_n4430_));
  NOR2_X1    g03428(.A1(new_n4430_), .A2(new_n4426_), .ZN(new_n4431_));
  AOI21_X1   g03429(.A1(\A[329] ), .A2(\A[330] ), .B(\A[328] ), .ZN(new_n4432_));
  AOI21_X1   g03430(.A1(\A[326] ), .A2(\A[327] ), .B(\A[325] ), .ZN(new_n4433_));
  NOR2_X1    g03431(.A1(new_n4433_), .A2(new_n3911_), .ZN(new_n4434_));
  NOR3_X1    g03432(.A1(new_n4434_), .A2(new_n3921_), .A3(new_n4432_), .ZN(new_n4435_));
  NOR2_X1    g03433(.A1(new_n4432_), .A2(new_n3921_), .ZN(new_n4436_));
  NOR3_X1    g03434(.A1(new_n4436_), .A2(new_n3911_), .A3(new_n4433_), .ZN(new_n4437_));
  NOR2_X1    g03435(.A1(new_n4435_), .A2(new_n4437_), .ZN(new_n4438_));
  NAND2_X1   g03436(.A1(new_n4438_), .A2(new_n3924_), .ZN(new_n4439_));
  XOR2_X1    g03437(.A1(new_n4436_), .A2(new_n4434_), .Z(new_n4440_));
  NAND2_X1   g03438(.A1(new_n4440_), .A2(new_n3972_), .ZN(new_n4441_));
  AOI22_X1   g03439(.A1(new_n4439_), .A2(new_n4441_), .B1(new_n3974_), .B2(new_n3970_), .ZN(new_n4442_));
  NAND3_X1   g03440(.A1(new_n4440_), .A2(new_n3936_), .A3(new_n3924_), .ZN(new_n4443_));
  NOR2_X1    g03441(.A1(new_n4436_), .A2(new_n4434_), .ZN(new_n4444_));
  NAND2_X1   g03442(.A1(new_n4436_), .A2(new_n4434_), .ZN(new_n4445_));
  AOI21_X1   g03443(.A1(new_n3924_), .A2(new_n4445_), .B(new_n4444_), .ZN(new_n4446_));
  NOR3_X1    g03444(.A1(new_n4443_), .A2(new_n3977_), .A3(new_n4446_), .ZN(new_n4447_));
  NOR3_X1    g03445(.A1(new_n4442_), .A2(new_n4431_), .A3(new_n4447_), .ZN(new_n4448_));
  NAND2_X1   g03446(.A1(new_n3975_), .A2(new_n4429_), .ZN(new_n4449_));
  NOR2_X1    g03447(.A1(new_n3947_), .A2(new_n3943_), .ZN(new_n4450_));
  NOR2_X1    g03448(.A1(new_n3953_), .A2(new_n3956_), .ZN(new_n4451_));
  NAND3_X1   g03449(.A1(new_n4425_), .A2(new_n4450_), .A3(new_n4451_), .ZN(new_n4452_));
  NAND2_X1   g03450(.A1(new_n4449_), .A2(new_n4452_), .ZN(new_n4453_));
  NOR2_X1    g03451(.A1(new_n4440_), .A2(new_n3972_), .ZN(new_n4454_));
  NOR2_X1    g03452(.A1(new_n4438_), .A2(new_n3924_), .ZN(new_n4455_));
  OAI22_X1   g03453(.A1(new_n4454_), .A2(new_n4455_), .B1(new_n3977_), .B2(new_n3937_), .ZN(new_n4456_));
  NOR4_X1    g03454(.A1(new_n3977_), .A2(new_n3972_), .A3(new_n3973_), .A4(new_n4438_), .ZN(new_n4457_));
  INV_X1     g03455(.I(new_n4457_), .ZN(new_n4458_));
  AOI21_X1   g03456(.A1(new_n4458_), .A2(new_n4456_), .B(new_n4453_), .ZN(new_n4459_));
  NOR4_X1    g03457(.A1(new_n4459_), .A2(new_n4448_), .A3(new_n4418_), .A4(new_n4050_), .ZN(new_n4460_));
  NOR3_X1    g03458(.A1(new_n3972_), .A2(new_n4438_), .A3(new_n3973_), .ZN(new_n4461_));
  INV_X1     g03459(.I(new_n4444_), .ZN(new_n4462_));
  NAND2_X1   g03460(.A1(new_n3924_), .A2(new_n4445_), .ZN(new_n4463_));
  NAND2_X1   g03461(.A1(new_n4463_), .A2(new_n4462_), .ZN(new_n4464_));
  NAND3_X1   g03462(.A1(new_n4464_), .A2(new_n3970_), .A3(new_n4461_), .ZN(new_n4465_));
  NAND3_X1   g03463(.A1(new_n4465_), .A2(new_n4456_), .A3(new_n4453_), .ZN(new_n4466_));
  OAI21_X1   g03464(.A1(new_n4442_), .A2(new_n4457_), .B(new_n4431_), .ZN(new_n4467_));
  AOI21_X1   g03465(.A1(new_n4466_), .A2(new_n4467_), .B(new_n4053_), .ZN(new_n4468_));
  NOR3_X1    g03466(.A1(new_n4460_), .A2(new_n4468_), .A3(new_n4417_), .ZN(new_n4469_));
  INV_X1     g03467(.I(new_n4469_), .ZN(new_n4470_));
  OAI21_X1   g03468(.A1(new_n4460_), .A2(new_n4468_), .B(new_n4417_), .ZN(new_n4471_));
  NAND2_X1   g03469(.A1(new_n4470_), .A2(new_n4471_), .ZN(new_n4472_));
  NOR4_X1    g03470(.A1(new_n3859_), .A2(new_n3863_), .A3(new_n3887_), .A4(new_n3884_), .ZN(new_n4473_));
  AOI21_X1   g03471(.A1(\A[347] ), .A2(\A[348] ), .B(\A[346] ), .ZN(new_n4474_));
  AOI21_X1   g03472(.A1(\A[344] ), .A2(\A[345] ), .B(\A[343] ), .ZN(new_n4475_));
  OAI22_X1   g03473(.A1(new_n3861_), .A2(new_n4475_), .B1(new_n4474_), .B2(new_n3872_), .ZN(new_n4476_));
  OR4_X2     g03474(.A1(new_n3861_), .A2(new_n4474_), .A3(new_n4475_), .A4(new_n3872_), .Z(new_n4477_));
  NAND2_X1   g03475(.A1(new_n4477_), .A2(new_n4476_), .ZN(new_n4478_));
  XOR2_X1    g03476(.A1(new_n4473_), .A2(new_n4478_), .Z(new_n4479_));
  NAND4_X1   g03477(.A1(new_n3842_), .A2(new_n3833_), .A3(new_n3844_), .A4(new_n3837_), .ZN(new_n4480_));
  AOI21_X1   g03478(.A1(\A[353] ), .A2(\A[354] ), .B(\A[352] ), .ZN(new_n4481_));
  AOI21_X1   g03479(.A1(\A[350] ), .A2(\A[351] ), .B(\A[349] ), .ZN(new_n4482_));
  NOR2_X1    g03480(.A1(new_n4482_), .A2(new_n3825_), .ZN(new_n4483_));
  NOR3_X1    g03481(.A1(new_n4483_), .A2(new_n3836_), .A3(new_n4481_), .ZN(new_n4484_));
  NOR2_X1    g03482(.A1(new_n4481_), .A2(new_n3836_), .ZN(new_n4485_));
  NOR3_X1    g03483(.A1(new_n4485_), .A2(new_n3825_), .A3(new_n4482_), .ZN(new_n4486_));
  NOR2_X1    g03484(.A1(new_n4484_), .A2(new_n4486_), .ZN(new_n4487_));
  NAND2_X1   g03485(.A1(new_n4487_), .A2(new_n4480_), .ZN(new_n4488_));
  NOR4_X1    g03486(.A1(new_n3823_), .A2(new_n3827_), .A3(new_n3851_), .A4(new_n3848_), .ZN(new_n4489_));
  XOR2_X1    g03487(.A1(new_n4483_), .A2(new_n4485_), .Z(new_n4490_));
  NAND2_X1   g03488(.A1(new_n4490_), .A2(new_n4489_), .ZN(new_n4491_));
  NAND2_X1   g03489(.A1(new_n4491_), .A2(new_n4488_), .ZN(new_n4492_));
  AOI21_X1   g03490(.A1(new_n3897_), .A2(new_n4492_), .B(new_n4479_), .ZN(new_n4493_));
  NOR2_X1    g03491(.A1(new_n4490_), .A2(new_n4489_), .ZN(new_n4494_));
  NOR2_X1    g03492(.A1(new_n4487_), .A2(new_n4480_), .ZN(new_n4495_));
  NOR2_X1    g03493(.A1(new_n4494_), .A2(new_n4495_), .ZN(new_n4496_));
  NAND2_X1   g03494(.A1(new_n3845_), .A2(new_n3838_), .ZN(new_n4497_));
  NAND3_X1   g03495(.A1(new_n4497_), .A2(new_n4485_), .A3(new_n4483_), .ZN(new_n4498_));
  NAND4_X1   g03496(.A1(new_n4496_), .A2(new_n3891_), .A3(new_n3892_), .A4(new_n4498_), .ZN(new_n4499_));
  OAI22_X1   g03497(.A1(new_n3898_), .A2(new_n3901_), .B1(new_n4494_), .B2(new_n4495_), .ZN(new_n4500_));
  NAND2_X1   g03498(.A1(new_n4496_), .A2(new_n3890_), .ZN(new_n4501_));
  NAND2_X1   g03499(.A1(new_n4501_), .A2(new_n4500_), .ZN(new_n4502_));
  AOI22_X1   g03500(.A1(new_n4502_), .A2(new_n4479_), .B1(new_n4493_), .B2(new_n4499_), .ZN(new_n4503_));
  NAND4_X1   g03501(.A1(new_n3895_), .A2(new_n3902_), .A3(new_n3896_), .A4(new_n3897_), .ZN(new_n4504_));
  NAND4_X1   g03502(.A1(new_n3800_), .A2(new_n3790_), .A3(new_n3795_), .A4(new_n3802_), .ZN(new_n4505_));
  AOI21_X1   g03503(.A1(\A[359] ), .A2(\A[360] ), .B(\A[358] ), .ZN(new_n4506_));
  NOR2_X1    g03504(.A1(new_n4506_), .A2(new_n3794_), .ZN(new_n4507_));
  AOI21_X1   g03505(.A1(\A[356] ), .A2(\A[357] ), .B(\A[355] ), .ZN(new_n4508_));
  NOR2_X1    g03506(.A1(new_n4508_), .A2(new_n3782_), .ZN(new_n4509_));
  NOR2_X1    g03507(.A1(new_n4507_), .A2(new_n4509_), .ZN(new_n4510_));
  NOR4_X1    g03508(.A1(new_n4506_), .A2(new_n4508_), .A3(new_n3782_), .A4(new_n3794_), .ZN(new_n4511_));
  NOR2_X1    g03509(.A1(new_n4510_), .A2(new_n4511_), .ZN(new_n4512_));
  XNOR2_X1   g03510(.A1(new_n4505_), .A2(new_n4512_), .ZN(new_n4513_));
  NAND4_X1   g03511(.A1(new_n3762_), .A2(new_n3753_), .A3(new_n3764_), .A4(new_n3757_), .ZN(new_n4514_));
  AOI21_X1   g03512(.A1(\A[365] ), .A2(\A[366] ), .B(\A[364] ), .ZN(new_n4515_));
  AOI21_X1   g03513(.A1(\A[362] ), .A2(\A[363] ), .B(\A[361] ), .ZN(new_n4516_));
  NOR2_X1    g03514(.A1(new_n4516_), .A2(new_n3745_), .ZN(new_n4517_));
  NOR3_X1    g03515(.A1(new_n4517_), .A2(new_n3756_), .A3(new_n4515_), .ZN(new_n4518_));
  NOR2_X1    g03516(.A1(new_n4515_), .A2(new_n3756_), .ZN(new_n4519_));
  NOR3_X1    g03517(.A1(new_n4519_), .A2(new_n3745_), .A3(new_n4516_), .ZN(new_n4520_));
  NOR2_X1    g03518(.A1(new_n4518_), .A2(new_n4520_), .ZN(new_n4521_));
  NAND2_X1   g03519(.A1(new_n4521_), .A2(new_n4514_), .ZN(new_n4522_));
  NOR4_X1    g03520(.A1(new_n3743_), .A2(new_n3747_), .A3(new_n3771_), .A4(new_n3768_), .ZN(new_n4523_));
  XOR2_X1    g03521(.A1(new_n4519_), .A2(new_n4517_), .Z(new_n4524_));
  NAND2_X1   g03522(.A1(new_n4524_), .A2(new_n4523_), .ZN(new_n4525_));
  AOI22_X1   g03523(.A1(new_n3774_), .A2(new_n3811_), .B1(new_n4522_), .B2(new_n4525_), .ZN(new_n4526_));
  NAND2_X1   g03524(.A1(new_n4525_), .A2(new_n4522_), .ZN(new_n4527_));
  INV_X1     g03525(.I(new_n4519_), .ZN(new_n4528_));
  INV_X1     g03526(.I(new_n4517_), .ZN(new_n4529_));
  NOR2_X1    g03527(.A1(new_n3748_), .A2(new_n3772_), .ZN(new_n4530_));
  NOR3_X1    g03528(.A1(new_n4530_), .A2(new_n4528_), .A3(new_n4529_), .ZN(new_n4531_));
  NOR4_X1    g03529(.A1(new_n4527_), .A2(new_n3813_), .A3(new_n3816_), .A4(new_n4531_), .ZN(new_n4532_));
  OAI21_X1   g03530(.A1(new_n4532_), .A2(new_n4526_), .B(new_n4513_), .ZN(new_n4533_));
  XOR2_X1    g03531(.A1(new_n4505_), .A2(new_n4512_), .Z(new_n4534_));
  NOR3_X1    g03532(.A1(new_n4523_), .A2(new_n4518_), .A3(new_n4520_), .ZN(new_n4535_));
  NOR2_X1    g03533(.A1(new_n4521_), .A2(new_n4514_), .ZN(new_n4536_));
  OAI22_X1   g03534(.A1(new_n3813_), .A2(new_n3816_), .B1(new_n4535_), .B2(new_n4536_), .ZN(new_n4537_));
  NAND4_X1   g03535(.A1(new_n3774_), .A2(new_n3811_), .A3(new_n4522_), .A4(new_n4525_), .ZN(new_n4538_));
  NAND3_X1   g03536(.A1(new_n4537_), .A2(new_n4538_), .A3(new_n4534_), .ZN(new_n4539_));
  AOI21_X1   g03537(.A1(new_n4533_), .A2(new_n4539_), .B(new_n4504_), .ZN(new_n4540_));
  NOR2_X1    g03538(.A1(new_n4535_), .A2(new_n4536_), .ZN(new_n4541_));
  NAND2_X1   g03539(.A1(new_n3765_), .A2(new_n3758_), .ZN(new_n4542_));
  NAND3_X1   g03540(.A1(new_n4542_), .A2(new_n4519_), .A3(new_n4517_), .ZN(new_n4543_));
  NAND4_X1   g03541(.A1(new_n4541_), .A2(new_n3774_), .A3(new_n3811_), .A4(new_n4543_), .ZN(new_n4544_));
  AOI21_X1   g03542(.A1(new_n4544_), .A2(new_n4537_), .B(new_n4534_), .ZN(new_n4545_));
  NOR3_X1    g03543(.A1(new_n4527_), .A2(new_n3813_), .A3(new_n3816_), .ZN(new_n4546_));
  NOR3_X1    g03544(.A1(new_n4546_), .A2(new_n4526_), .A3(new_n4513_), .ZN(new_n4547_));
  NOR3_X1    g03545(.A1(new_n4545_), .A2(new_n4547_), .A3(new_n3894_), .ZN(new_n4548_));
  OAI21_X1   g03546(.A1(new_n4540_), .A2(new_n4548_), .B(new_n4503_), .ZN(new_n4549_));
  NAND4_X1   g03547(.A1(new_n3878_), .A2(new_n3869_), .A3(new_n3880_), .A4(new_n3873_), .ZN(new_n4550_));
  XOR2_X1    g03548(.A1(new_n4550_), .A2(new_n4478_), .Z(new_n4551_));
  OAI21_X1   g03549(.A1(new_n4496_), .A2(new_n3890_), .B(new_n4551_), .ZN(new_n4552_));
  INV_X1     g03550(.I(new_n4485_), .ZN(new_n4553_));
  INV_X1     g03551(.I(new_n4483_), .ZN(new_n4554_));
  NOR2_X1    g03552(.A1(new_n3828_), .A2(new_n3852_), .ZN(new_n4555_));
  NOR3_X1    g03553(.A1(new_n4555_), .A2(new_n4553_), .A3(new_n4554_), .ZN(new_n4556_));
  NOR4_X1    g03554(.A1(new_n4492_), .A2(new_n3898_), .A3(new_n3901_), .A4(new_n4556_), .ZN(new_n4557_));
  AOI22_X1   g03555(.A1(new_n3891_), .A2(new_n3892_), .B1(new_n4488_), .B2(new_n4491_), .ZN(new_n4558_));
  NOR3_X1    g03556(.A1(new_n4492_), .A2(new_n3898_), .A3(new_n3901_), .ZN(new_n4559_));
  NOR2_X1    g03557(.A1(new_n4559_), .A2(new_n4558_), .ZN(new_n4560_));
  OAI22_X1   g03558(.A1(new_n4560_), .A2(new_n4551_), .B1(new_n4552_), .B2(new_n4557_), .ZN(new_n4561_));
  OAI21_X1   g03559(.A1(new_n4545_), .A2(new_n4547_), .B(new_n3894_), .ZN(new_n4562_));
  NAND3_X1   g03560(.A1(new_n4533_), .A2(new_n4504_), .A3(new_n4539_), .ZN(new_n4563_));
  NAND3_X1   g03561(.A1(new_n4562_), .A2(new_n4563_), .A3(new_n4561_), .ZN(new_n4564_));
  AOI21_X1   g03562(.A1(new_n4549_), .A2(new_n4564_), .B(new_n4055_), .ZN(new_n4565_));
  AOI21_X1   g03563(.A1(new_n4562_), .A2(new_n4563_), .B(new_n4561_), .ZN(new_n4566_));
  NOR3_X1    g03564(.A1(new_n4540_), .A2(new_n4548_), .A3(new_n4503_), .ZN(new_n4567_));
  NOR3_X1    g03565(.A1(new_n4363_), .A2(new_n4567_), .A3(new_n4566_), .ZN(new_n4568_));
  NOR2_X1    g03566(.A1(new_n4568_), .A2(new_n4565_), .ZN(new_n4569_));
  NOR2_X1    g03567(.A1(new_n4569_), .A2(new_n4472_), .ZN(new_n4570_));
  OAI21_X1   g03568(.A1(new_n4567_), .A2(new_n4566_), .B(new_n4363_), .ZN(new_n4571_));
  NAND2_X1   g03569(.A1(new_n4571_), .A2(new_n4472_), .ZN(new_n4572_));
  NOR2_X1    g03570(.A1(new_n4572_), .A2(new_n4568_), .ZN(new_n4573_));
  NOR2_X1    g03571(.A1(new_n4573_), .A2(new_n4570_), .ZN(new_n4574_));
  AOI21_X1   g03572(.A1(\A[299] ), .A2(\A[300] ), .B(\A[298] ), .ZN(new_n4575_));
  NOR2_X1    g03573(.A1(new_n4575_), .A2(new_n4194_), .ZN(new_n4576_));
  AOI21_X1   g03574(.A1(\A[296] ), .A2(\A[297] ), .B(\A[295] ), .ZN(new_n4577_));
  NOR2_X1    g03575(.A1(new_n4577_), .A2(new_n4172_), .ZN(new_n4578_));
  NOR2_X1    g03576(.A1(new_n4576_), .A2(new_n4578_), .ZN(new_n4579_));
  NOR4_X1    g03577(.A1(new_n4575_), .A2(new_n4577_), .A3(new_n4172_), .A4(new_n4194_), .ZN(new_n4580_));
  NOR2_X1    g03578(.A1(new_n4579_), .A2(new_n4580_), .ZN(new_n4581_));
  NAND2_X1   g03579(.A1(new_n4202_), .A2(new_n4581_), .ZN(new_n4582_));
  OAI22_X1   g03580(.A1(new_n4172_), .A2(new_n4577_), .B1(new_n4575_), .B2(new_n4194_), .ZN(new_n4583_));
  NAND2_X1   g03581(.A1(new_n4576_), .A2(new_n4578_), .ZN(new_n4584_));
  NAND2_X1   g03582(.A1(new_n4584_), .A2(new_n4583_), .ZN(new_n4585_));
  NAND2_X1   g03583(.A1(new_n4184_), .A2(new_n4585_), .ZN(new_n4586_));
  NAND2_X1   g03584(.A1(new_n4582_), .A2(new_n4586_), .ZN(new_n4587_));
  AOI21_X1   g03585(.A1(\A[305] ), .A2(\A[306] ), .B(\A[304] ), .ZN(new_n4588_));
  NOR2_X1    g03586(.A1(new_n4588_), .A2(new_n4148_), .ZN(new_n4589_));
  AOI21_X1   g03587(.A1(\A[302] ), .A2(\A[303] ), .B(\A[301] ), .ZN(new_n4590_));
  NOR2_X1    g03588(.A1(new_n4590_), .A2(new_n4138_), .ZN(new_n4591_));
  XOR2_X1    g03589(.A1(new_n4589_), .A2(new_n4591_), .Z(new_n4592_));
  NOR2_X1    g03590(.A1(new_n4592_), .A2(new_n4199_), .ZN(new_n4593_));
  NOR3_X1    g03591(.A1(new_n4591_), .A2(new_n4148_), .A3(new_n4588_), .ZN(new_n4594_));
  NOR3_X1    g03592(.A1(new_n4589_), .A2(new_n4138_), .A3(new_n4590_), .ZN(new_n4595_));
  NOR2_X1    g03593(.A1(new_n4594_), .A2(new_n4595_), .ZN(new_n4596_));
  NOR2_X1    g03594(.A1(new_n4596_), .A2(new_n4151_), .ZN(new_n4597_));
  NOR2_X1    g03595(.A1(new_n4593_), .A2(new_n4597_), .ZN(new_n4598_));
  NOR4_X1    g03596(.A1(new_n4196_), .A2(new_n4199_), .A3(new_n4200_), .A4(new_n4184_), .ZN(new_n4599_));
  OAI21_X1   g03597(.A1(new_n4598_), .A2(new_n4599_), .B(new_n4587_), .ZN(new_n4600_));
  NOR4_X1    g03598(.A1(new_n4204_), .A2(new_n4199_), .A3(new_n4200_), .A4(new_n4596_), .ZN(new_n4601_));
  OAI22_X1   g03599(.A1(new_n4593_), .A2(new_n4597_), .B1(new_n4204_), .B2(new_n4164_), .ZN(new_n4602_));
  INV_X1     g03600(.I(new_n4602_), .ZN(new_n4603_));
  NOR2_X1    g03601(.A1(new_n4603_), .A2(new_n4601_), .ZN(new_n4604_));
  OAI22_X1   g03602(.A1(new_n4604_), .A2(new_n4587_), .B1(new_n4600_), .B2(new_n4601_), .ZN(new_n4605_));
  NAND2_X1   g03603(.A1(new_n4127_), .A2(new_n4130_), .ZN(new_n4606_));
  NAND2_X1   g03604(.A1(new_n4090_), .A2(new_n4123_), .ZN(new_n4607_));
  AOI22_X1   g03605(.A1(new_n4606_), .A2(new_n4607_), .B1(new_n4208_), .B2(new_n4209_), .ZN(new_n4608_));
  AOI21_X1   g03606(.A1(\A[311] ), .A2(\A[312] ), .B(\A[310] ), .ZN(new_n4609_));
  AOI21_X1   g03607(.A1(\A[308] ), .A2(\A[309] ), .B(\A[307] ), .ZN(new_n4610_));
  OAI22_X1   g03608(.A1(new_n4098_), .A2(new_n4610_), .B1(new_n4609_), .B2(new_n4120_), .ZN(new_n4611_));
  INV_X1     g03609(.I(new_n4611_), .ZN(new_n4612_));
  NOR4_X1    g03610(.A1(new_n4609_), .A2(new_n4610_), .A3(new_n4098_), .A4(new_n4120_), .ZN(new_n4613_));
  NOR2_X1    g03611(.A1(new_n4612_), .A2(new_n4613_), .ZN(new_n4614_));
  NAND2_X1   g03612(.A1(new_n4614_), .A2(new_n4128_), .ZN(new_n4615_));
  INV_X1     g03613(.I(new_n4613_), .ZN(new_n4616_));
  NAND2_X1   g03614(.A1(new_n4616_), .A2(new_n4611_), .ZN(new_n4617_));
  NAND2_X1   g03615(.A1(new_n4110_), .A2(new_n4617_), .ZN(new_n4618_));
  NAND2_X1   g03616(.A1(new_n4615_), .A2(new_n4618_), .ZN(new_n4619_));
  AOI21_X1   g03617(.A1(\A[317] ), .A2(\A[318] ), .B(\A[316] ), .ZN(new_n4620_));
  AOI21_X1   g03618(.A1(\A[314] ), .A2(\A[315] ), .B(\A[313] ), .ZN(new_n4621_));
  NOR2_X1    g03619(.A1(new_n4621_), .A2(new_n4064_), .ZN(new_n4622_));
  NOR3_X1    g03620(.A1(new_n4622_), .A2(new_n4074_), .A3(new_n4620_), .ZN(new_n4623_));
  NOR2_X1    g03621(.A1(new_n4620_), .A2(new_n4074_), .ZN(new_n4624_));
  NOR3_X1    g03622(.A1(new_n4624_), .A2(new_n4064_), .A3(new_n4621_), .ZN(new_n4625_));
  NOR2_X1    g03623(.A1(new_n4623_), .A2(new_n4625_), .ZN(new_n4626_));
  NAND2_X1   g03624(.A1(new_n4078_), .A2(new_n4626_), .ZN(new_n4627_));
  XOR2_X1    g03625(.A1(new_n4624_), .A2(new_n4622_), .Z(new_n4628_));
  NAND2_X1   g03626(.A1(new_n4628_), .A2(new_n4125_), .ZN(new_n4629_));
  AOI22_X1   g03627(.A1(new_n4627_), .A2(new_n4629_), .B1(new_n4127_), .B2(new_n4123_), .ZN(new_n4630_));
  NOR4_X1    g03628(.A1(new_n4130_), .A2(new_n4125_), .A3(new_n4126_), .A4(new_n4626_), .ZN(new_n4631_));
  NOR3_X1    g03629(.A1(new_n4630_), .A2(new_n4619_), .A3(new_n4631_), .ZN(new_n4632_));
  NOR2_X1    g03630(.A1(new_n4110_), .A2(new_n4617_), .ZN(new_n4633_));
  NOR2_X1    g03631(.A1(new_n4614_), .A2(new_n4128_), .ZN(new_n4634_));
  NOR2_X1    g03632(.A1(new_n4634_), .A2(new_n4633_), .ZN(new_n4635_));
  NOR2_X1    g03633(.A1(new_n4628_), .A2(new_n4125_), .ZN(new_n4636_));
  NOR2_X1    g03634(.A1(new_n4078_), .A2(new_n4626_), .ZN(new_n4637_));
  OAI22_X1   g03635(.A1(new_n4636_), .A2(new_n4637_), .B1(new_n4090_), .B2(new_n4130_), .ZN(new_n4638_));
  NAND4_X1   g03636(.A1(new_n4123_), .A2(new_n4078_), .A3(new_n4089_), .A4(new_n4628_), .ZN(new_n4639_));
  AOI21_X1   g03637(.A1(new_n4638_), .A2(new_n4639_), .B(new_n4635_), .ZN(new_n4640_));
  OAI21_X1   g03638(.A1(new_n4632_), .A2(new_n4640_), .B(new_n4608_), .ZN(new_n4641_));
  NAND3_X1   g03639(.A1(new_n4638_), .A2(new_n4635_), .A3(new_n4639_), .ZN(new_n4642_));
  OAI21_X1   g03640(.A1(new_n4630_), .A2(new_n4631_), .B(new_n4619_), .ZN(new_n4643_));
  NAND3_X1   g03641(.A1(new_n4642_), .A2(new_n4643_), .A3(new_n4206_), .ZN(new_n4644_));
  NAND3_X1   g03642(.A1(new_n4605_), .A2(new_n4644_), .A3(new_n4641_), .ZN(new_n4645_));
  NOR2_X1    g03643(.A1(new_n4184_), .A2(new_n4585_), .ZN(new_n4646_));
  NOR2_X1    g03644(.A1(new_n4202_), .A2(new_n4581_), .ZN(new_n4647_));
  NOR2_X1    g03645(.A1(new_n4647_), .A2(new_n4646_), .ZN(new_n4648_));
  NAND2_X1   g03646(.A1(new_n4596_), .A2(new_n4151_), .ZN(new_n4649_));
  NAND2_X1   g03647(.A1(new_n4592_), .A2(new_n4199_), .ZN(new_n4650_));
  NAND2_X1   g03648(.A1(new_n4650_), .A2(new_n4649_), .ZN(new_n4651_));
  NAND2_X1   g03649(.A1(new_n4201_), .A2(new_n4197_), .ZN(new_n4652_));
  AOI21_X1   g03650(.A1(new_n4652_), .A2(new_n4651_), .B(new_n4648_), .ZN(new_n4653_));
  INV_X1     g03651(.I(new_n4601_), .ZN(new_n4654_));
  NAND2_X1   g03652(.A1(new_n4654_), .A2(new_n4602_), .ZN(new_n4655_));
  AOI22_X1   g03653(.A1(new_n4655_), .A2(new_n4648_), .B1(new_n4653_), .B2(new_n4654_), .ZN(new_n4656_));
  AOI21_X1   g03654(.A1(new_n4642_), .A2(new_n4643_), .B(new_n4206_), .ZN(new_n4657_));
  NOR3_X1    g03655(.A1(new_n4632_), .A2(new_n4640_), .A3(new_n4608_), .ZN(new_n4658_));
  OAI21_X1   g03656(.A1(new_n4657_), .A2(new_n4658_), .B(new_n4656_), .ZN(new_n4659_));
  NAND2_X1   g03657(.A1(new_n4645_), .A2(new_n4659_), .ZN(new_n4660_));
  INV_X1     g03658(.I(new_n4660_), .ZN(new_n4661_));
  AOI21_X1   g03659(.A1(\A[287] ), .A2(\A[288] ), .B(\A[286] ), .ZN(new_n4662_));
  AOI21_X1   g03660(.A1(\A[284] ), .A2(\A[285] ), .B(\A[283] ), .ZN(new_n4663_));
  OAI22_X1   g03661(.A1(new_n4251_), .A2(new_n4663_), .B1(new_n4662_), .B2(new_n4261_), .ZN(new_n4664_));
  INV_X1     g03662(.I(new_n4664_), .ZN(new_n4665_));
  NOR4_X1    g03663(.A1(new_n4662_), .A2(new_n4663_), .A3(new_n4251_), .A4(new_n4261_), .ZN(new_n4666_));
  NOR2_X1    g03664(.A1(new_n4665_), .A2(new_n4666_), .ZN(new_n4667_));
  NAND2_X1   g03665(.A1(new_n4281_), .A2(new_n4667_), .ZN(new_n4668_));
  INV_X1     g03666(.I(new_n4666_), .ZN(new_n4669_));
  NAND2_X1   g03667(.A1(new_n4669_), .A2(new_n4664_), .ZN(new_n4670_));
  NAND2_X1   g03668(.A1(new_n4264_), .A2(new_n4670_), .ZN(new_n4671_));
  NAND2_X1   g03669(.A1(new_n4668_), .A2(new_n4671_), .ZN(new_n4672_));
  AOI21_X1   g03670(.A1(new_n4227_), .A2(new_n4229_), .B(new_n4228_), .ZN(new_n4673_));
  AOI21_X1   g03671(.A1(new_n4217_), .A2(new_n4219_), .B(new_n4218_), .ZN(new_n4674_));
  XOR2_X1    g03672(.A1(new_n4673_), .A2(new_n4674_), .Z(new_n4675_));
  NOR2_X1    g03673(.A1(new_n4675_), .A2(new_n4278_), .ZN(new_n4676_));
  XNOR2_X1   g03674(.A1(new_n4673_), .A2(new_n4674_), .ZN(new_n4677_));
  NOR2_X1    g03675(.A1(new_n4677_), .A2(new_n4232_), .ZN(new_n4678_));
  NOR2_X1    g03676(.A1(new_n4678_), .A2(new_n4676_), .ZN(new_n4679_));
  NOR2_X1    g03677(.A1(new_n4243_), .A2(new_n4283_), .ZN(new_n4680_));
  NOR2_X1    g03678(.A1(new_n4679_), .A2(new_n4680_), .ZN(new_n4681_));
  NOR4_X1    g03679(.A1(new_n4283_), .A2(new_n4278_), .A3(new_n4279_), .A4(new_n4677_), .ZN(new_n4682_));
  NOR3_X1    g03680(.A1(new_n4681_), .A2(new_n4672_), .A3(new_n4682_), .ZN(new_n4683_));
  NOR2_X1    g03681(.A1(new_n4264_), .A2(new_n4670_), .ZN(new_n4684_));
  NOR2_X1    g03682(.A1(new_n4281_), .A2(new_n4667_), .ZN(new_n4685_));
  NOR2_X1    g03683(.A1(new_n4685_), .A2(new_n4684_), .ZN(new_n4686_));
  NAND2_X1   g03684(.A1(new_n4677_), .A2(new_n4232_), .ZN(new_n4687_));
  NAND2_X1   g03685(.A1(new_n4675_), .A2(new_n4278_), .ZN(new_n4688_));
  NAND2_X1   g03686(.A1(new_n4687_), .A2(new_n4688_), .ZN(new_n4689_));
  NAND2_X1   g03687(.A1(new_n4280_), .A2(new_n4276_), .ZN(new_n4690_));
  NAND2_X1   g03688(.A1(new_n4689_), .A2(new_n4690_), .ZN(new_n4691_));
  INV_X1     g03689(.I(new_n4682_), .ZN(new_n4692_));
  AOI21_X1   g03690(.A1(new_n4691_), .A2(new_n4692_), .B(new_n4686_), .ZN(new_n4693_));
  NOR2_X1    g03691(.A1(new_n4683_), .A2(new_n4693_), .ZN(new_n4694_));
  AOI21_X1   g03692(.A1(\A[275] ), .A2(\A[276] ), .B(\A[274] ), .ZN(new_n4695_));
  NOR2_X1    g03693(.A1(new_n4695_), .A2(new_n4336_), .ZN(new_n4696_));
  AOI21_X1   g03694(.A1(\A[272] ), .A2(\A[273] ), .B(\A[271] ), .ZN(new_n4697_));
  NOR2_X1    g03695(.A1(new_n4697_), .A2(new_n4326_), .ZN(new_n4698_));
  NOR2_X1    g03696(.A1(new_n4696_), .A2(new_n4698_), .ZN(new_n4699_));
  NOR4_X1    g03697(.A1(new_n4695_), .A2(new_n4697_), .A3(new_n4326_), .A4(new_n4336_), .ZN(new_n4700_));
  NOR2_X1    g03698(.A1(new_n4699_), .A2(new_n4700_), .ZN(new_n4701_));
  NAND2_X1   g03699(.A1(new_n4338_), .A2(new_n4701_), .ZN(new_n4702_));
  NOR4_X1    g03700(.A1(new_n4341_), .A2(new_n4343_), .A3(new_n4348_), .A4(new_n4346_), .ZN(new_n4703_));
  OAI22_X1   g03701(.A1(new_n4326_), .A2(new_n4697_), .B1(new_n4695_), .B2(new_n4336_), .ZN(new_n4704_));
  INV_X1     g03702(.I(new_n4700_), .ZN(new_n4705_));
  NAND2_X1   g03703(.A1(new_n4705_), .A2(new_n4704_), .ZN(new_n4706_));
  NAND2_X1   g03704(.A1(new_n4703_), .A2(new_n4706_), .ZN(new_n4707_));
  NAND2_X1   g03705(.A1(new_n4707_), .A2(new_n4702_), .ZN(new_n4708_));
  AOI21_X1   g03706(.A1(\A[281] ), .A2(\A[282] ), .B(\A[280] ), .ZN(new_n4709_));
  NOR2_X1    g03707(.A1(new_n4709_), .A2(new_n4301_), .ZN(new_n4710_));
  AOI21_X1   g03708(.A1(\A[278] ), .A2(\A[279] ), .B(\A[277] ), .ZN(new_n4711_));
  NOR2_X1    g03709(.A1(new_n4711_), .A2(new_n4291_), .ZN(new_n4712_));
  XOR2_X1    g03710(.A1(new_n4710_), .A2(new_n4712_), .Z(new_n4713_));
  NOR2_X1    g03711(.A1(new_n4713_), .A2(new_n4305_), .ZN(new_n4714_));
  NAND4_X1   g03712(.A1(new_n4308_), .A2(new_n4310_), .A3(new_n4315_), .A4(new_n4313_), .ZN(new_n4715_));
  NOR3_X1    g03713(.A1(new_n4712_), .A2(new_n4301_), .A3(new_n4709_), .ZN(new_n4716_));
  NOR3_X1    g03714(.A1(new_n4710_), .A2(new_n4291_), .A3(new_n4711_), .ZN(new_n4717_));
  NOR2_X1    g03715(.A1(new_n4716_), .A2(new_n4717_), .ZN(new_n4718_));
  NOR2_X1    g03716(.A1(new_n4715_), .A2(new_n4718_), .ZN(new_n4719_));
  NOR2_X1    g03717(.A1(new_n4714_), .A2(new_n4719_), .ZN(new_n4720_));
  OAI22_X1   g03718(.A1(new_n4290_), .A2(new_n4294_), .B1(new_n4304_), .B2(new_n4300_), .ZN(new_n4721_));
  NAND2_X1   g03719(.A1(new_n4715_), .A2(new_n4721_), .ZN(new_n4722_));
  NOR2_X1    g03720(.A1(new_n4722_), .A2(new_n4350_), .ZN(new_n4723_));
  OAI21_X1   g03721(.A1(new_n4720_), .A2(new_n4723_), .B(new_n4708_), .ZN(new_n4724_));
  NOR4_X1    g03722(.A1(new_n4350_), .A2(new_n4305_), .A3(new_n4316_), .A4(new_n4718_), .ZN(new_n4725_));
  NOR2_X1    g03723(.A1(new_n4724_), .A2(new_n4725_), .ZN(new_n4726_));
  OAI22_X1   g03724(.A1(new_n4714_), .A2(new_n4719_), .B1(new_n4722_), .B2(new_n4350_), .ZN(new_n4727_));
  INV_X1     g03725(.I(new_n4725_), .ZN(new_n4728_));
  AOI21_X1   g03726(.A1(new_n4728_), .A2(new_n4727_), .B(new_n4708_), .ZN(new_n4729_));
  NOR3_X1    g03727(.A1(new_n4726_), .A2(new_n4729_), .A3(new_n4354_), .ZN(new_n4730_));
  NAND2_X1   g03728(.A1(new_n4280_), .A2(new_n4283_), .ZN(new_n4731_));
  NAND2_X1   g03729(.A1(new_n4243_), .A2(new_n4276_), .ZN(new_n4732_));
  AOI22_X1   g03730(.A1(new_n4356_), .A2(new_n4351_), .B1(new_n4731_), .B2(new_n4732_), .ZN(new_n4733_));
  NOR2_X1    g03731(.A1(new_n4703_), .A2(new_n4706_), .ZN(new_n4734_));
  NOR2_X1    g03732(.A1(new_n4338_), .A2(new_n4701_), .ZN(new_n4735_));
  NOR2_X1    g03733(.A1(new_n4734_), .A2(new_n4735_), .ZN(new_n4736_));
  NAND2_X1   g03734(.A1(new_n4715_), .A2(new_n4718_), .ZN(new_n4737_));
  NAND2_X1   g03735(.A1(new_n4713_), .A2(new_n4305_), .ZN(new_n4738_));
  NAND2_X1   g03736(.A1(new_n4738_), .A2(new_n4737_), .ZN(new_n4739_));
  NAND3_X1   g03737(.A1(new_n4317_), .A2(new_n4338_), .A3(new_n4349_), .ZN(new_n4740_));
  AOI21_X1   g03738(.A1(new_n4740_), .A2(new_n4739_), .B(new_n4736_), .ZN(new_n4741_));
  NAND2_X1   g03739(.A1(new_n4741_), .A2(new_n4728_), .ZN(new_n4742_));
  NOR2_X1    g03740(.A1(new_n4720_), .A2(new_n4723_), .ZN(new_n4743_));
  OAI21_X1   g03741(.A1(new_n4743_), .A2(new_n4725_), .B(new_n4736_), .ZN(new_n4744_));
  AOI21_X1   g03742(.A1(new_n4744_), .A2(new_n4742_), .B(new_n4733_), .ZN(new_n4745_));
  NOR3_X1    g03743(.A1(new_n4730_), .A2(new_n4745_), .A3(new_n4694_), .ZN(new_n4746_));
  NAND3_X1   g03744(.A1(new_n4691_), .A2(new_n4692_), .A3(new_n4686_), .ZN(new_n4747_));
  OAI21_X1   g03745(.A1(new_n4681_), .A2(new_n4682_), .B(new_n4672_), .ZN(new_n4748_));
  NAND2_X1   g03746(.A1(new_n4748_), .A2(new_n4747_), .ZN(new_n4749_));
  NAND3_X1   g03747(.A1(new_n4744_), .A2(new_n4742_), .A3(new_n4733_), .ZN(new_n4750_));
  OAI21_X1   g03748(.A1(new_n4726_), .A2(new_n4729_), .B(new_n4354_), .ZN(new_n4751_));
  AOI21_X1   g03749(.A1(new_n4751_), .A2(new_n4750_), .B(new_n4749_), .ZN(new_n4752_));
  NOR3_X1    g03750(.A1(new_n4360_), .A2(new_n4746_), .A3(new_n4752_), .ZN(new_n4753_));
  NAND3_X1   g03751(.A1(new_n4750_), .A2(new_n4751_), .A3(new_n4749_), .ZN(new_n4754_));
  OAI21_X1   g03752(.A1(new_n4745_), .A2(new_n4730_), .B(new_n4694_), .ZN(new_n4755_));
  AOI21_X1   g03753(.A1(new_n4755_), .A2(new_n4754_), .B(new_n4359_), .ZN(new_n4756_));
  NOR3_X1    g03754(.A1(new_n4661_), .A2(new_n4753_), .A3(new_n4756_), .ZN(new_n4757_));
  NAND3_X1   g03755(.A1(new_n4755_), .A2(new_n4754_), .A3(new_n4359_), .ZN(new_n4758_));
  OAI21_X1   g03756(.A1(new_n4752_), .A2(new_n4746_), .B(new_n4360_), .ZN(new_n4759_));
  AOI21_X1   g03757(.A1(new_n4759_), .A2(new_n4758_), .B(new_n4660_), .ZN(new_n4760_));
  NOR3_X1    g03758(.A1(new_n4757_), .A2(new_n4760_), .A3(new_n4362_), .ZN(new_n4761_));
  INV_X1     g03759(.I(new_n4362_), .ZN(new_n4762_));
  NAND3_X1   g03760(.A1(new_n4759_), .A2(new_n4758_), .A3(new_n4660_), .ZN(new_n4763_));
  OAI21_X1   g03761(.A1(new_n4756_), .A2(new_n4753_), .B(new_n4661_), .ZN(new_n4764_));
  AOI21_X1   g03762(.A1(new_n4764_), .A2(new_n4763_), .B(new_n4762_), .ZN(new_n4765_));
  NOR3_X1    g03763(.A1(new_n4574_), .A2(new_n4765_), .A3(new_n4761_), .ZN(new_n4766_));
  OAI22_X1   g03764(.A1(new_n4572_), .A2(new_n4568_), .B1(new_n4569_), .B2(new_n4472_), .ZN(new_n4767_));
  NAND3_X1   g03765(.A1(new_n4764_), .A2(new_n4763_), .A3(new_n4762_), .ZN(new_n4768_));
  OAI21_X1   g03766(.A1(new_n4757_), .A2(new_n4760_), .B(new_n4362_), .ZN(new_n4769_));
  AOI21_X1   g03767(.A1(new_n4768_), .A2(new_n4769_), .B(new_n4767_), .ZN(new_n4770_));
  NOR2_X1    g03768(.A1(new_n4766_), .A2(new_n4770_), .ZN(new_n4771_));
  AOI21_X1   g03769(.A1(\A[395] ), .A2(\A[396] ), .B(\A[394] ), .ZN(new_n4772_));
  AOI21_X1   g03770(.A1(\A[392] ), .A2(\A[393] ), .B(\A[391] ), .ZN(new_n4773_));
  OAI22_X1   g03771(.A1(new_n3257_), .A2(new_n4773_), .B1(new_n4772_), .B2(new_n3267_), .ZN(new_n4774_));
  NOR4_X1    g03772(.A1(new_n4772_), .A2(new_n4773_), .A3(new_n3257_), .A4(new_n3267_), .ZN(new_n4775_));
  INV_X1     g03773(.I(new_n4775_), .ZN(new_n4776_));
  NAND3_X1   g03774(.A1(new_n3317_), .A2(new_n4774_), .A3(new_n4776_), .ZN(new_n4777_));
  NAND2_X1   g03775(.A1(new_n4776_), .A2(new_n4774_), .ZN(new_n4778_));
  NAND2_X1   g03776(.A1(new_n3270_), .A2(new_n4778_), .ZN(new_n4779_));
  NAND2_X1   g03777(.A1(new_n4779_), .A2(new_n4777_), .ZN(new_n4780_));
  AOI21_X1   g03778(.A1(\A[401] ), .A2(\A[402] ), .B(\A[400] ), .ZN(new_n4781_));
  AOI21_X1   g03779(.A1(\A[398] ), .A2(\A[399] ), .B(\A[397] ), .ZN(new_n4782_));
  NOR2_X1    g03780(.A1(new_n4782_), .A2(new_n3291_), .ZN(new_n4783_));
  NOR3_X1    g03781(.A1(new_n4783_), .A2(new_n3301_), .A3(new_n4781_), .ZN(new_n4784_));
  NOR2_X1    g03782(.A1(new_n4781_), .A2(new_n3301_), .ZN(new_n4785_));
  NOR3_X1    g03783(.A1(new_n4785_), .A2(new_n3291_), .A3(new_n4782_), .ZN(new_n4786_));
  NOR2_X1    g03784(.A1(new_n4784_), .A2(new_n4786_), .ZN(new_n4787_));
  NOR2_X1    g03785(.A1(new_n3303_), .A2(new_n4787_), .ZN(new_n4788_));
  XOR2_X1    g03786(.A1(new_n4785_), .A2(new_n4783_), .Z(new_n4789_));
  NOR2_X1    g03787(.A1(new_n4789_), .A2(new_n3320_), .ZN(new_n4790_));
  OAI22_X1   g03788(.A1(new_n3319_), .A2(new_n3315_), .B1(new_n4790_), .B2(new_n4788_), .ZN(new_n4791_));
  NAND3_X1   g03789(.A1(new_n3314_), .A2(new_n4785_), .A3(new_n4783_), .ZN(new_n4792_));
  NOR3_X1    g03790(.A1(new_n3321_), .A2(new_n3320_), .A3(new_n4787_), .ZN(new_n4793_));
  NAND3_X1   g03791(.A1(new_n4793_), .A2(new_n3282_), .A3(new_n4792_), .ZN(new_n4794_));
  NAND3_X1   g03792(.A1(new_n4791_), .A2(new_n4794_), .A3(new_n4780_), .ZN(new_n4795_));
  AND2_X2    g03793(.A1(new_n4779_), .A2(new_n4777_), .Z(new_n4796_));
  NAND2_X1   g03794(.A1(new_n4789_), .A2(new_n3320_), .ZN(new_n4797_));
  NAND2_X1   g03795(.A1(new_n3303_), .A2(new_n4787_), .ZN(new_n4798_));
  AOI22_X1   g03796(.A1(new_n3282_), .A2(new_n3322_), .B1(new_n4797_), .B2(new_n4798_), .ZN(new_n4799_));
  NOR4_X1    g03797(.A1(new_n3319_), .A2(new_n3320_), .A3(new_n3321_), .A4(new_n4787_), .ZN(new_n4800_));
  OAI21_X1   g03798(.A1(new_n4799_), .A2(new_n4800_), .B(new_n4796_), .ZN(new_n4801_));
  NAND2_X1   g03799(.A1(new_n4801_), .A2(new_n4795_), .ZN(new_n4802_));
  AOI21_X1   g03800(.A1(\A[407] ), .A2(\A[408] ), .B(\A[406] ), .ZN(new_n4803_));
  AOI21_X1   g03801(.A1(\A[404] ), .A2(\A[405] ), .B(\A[403] ), .ZN(new_n4804_));
  OAI22_X1   g03802(.A1(new_n3332_), .A2(new_n4804_), .B1(new_n4803_), .B2(new_n3354_), .ZN(new_n4805_));
  NOR4_X1    g03803(.A1(new_n4803_), .A2(new_n4804_), .A3(new_n3332_), .A4(new_n3354_), .ZN(new_n4806_));
  INV_X1     g03804(.I(new_n4806_), .ZN(new_n4807_));
  NAND2_X1   g03805(.A1(new_n4807_), .A2(new_n4805_), .ZN(new_n4808_));
  XOR2_X1    g03806(.A1(new_n3344_), .A2(new_n4808_), .Z(new_n4809_));
  AOI21_X1   g03807(.A1(\A[413] ), .A2(\A[414] ), .B(\A[412] ), .ZN(new_n4810_));
  AOI21_X1   g03808(.A1(\A[410] ), .A2(\A[411] ), .B(\A[409] ), .ZN(new_n4811_));
  NOR2_X1    g03809(.A1(new_n4811_), .A2(new_n3365_), .ZN(new_n4812_));
  NOR3_X1    g03810(.A1(new_n4812_), .A2(new_n3374_), .A3(new_n4810_), .ZN(new_n4813_));
  NOR2_X1    g03811(.A1(new_n4810_), .A2(new_n3374_), .ZN(new_n4814_));
  NOR3_X1    g03812(.A1(new_n4814_), .A2(new_n3365_), .A3(new_n4811_), .ZN(new_n4815_));
  NOR2_X1    g03813(.A1(new_n4815_), .A2(new_n4813_), .ZN(new_n4816_));
  NOR2_X1    g03814(.A1(new_n4816_), .A2(new_n3376_), .ZN(new_n4817_));
  NOR4_X1    g03815(.A1(new_n3379_), .A2(new_n3382_), .A3(new_n3385_), .A4(new_n3388_), .ZN(new_n4818_));
  XOR2_X1    g03816(.A1(new_n4814_), .A2(new_n4812_), .Z(new_n4819_));
  NOR2_X1    g03817(.A1(new_n4819_), .A2(new_n4818_), .ZN(new_n4820_));
  OAI22_X1   g03818(.A1(new_n4820_), .A2(new_n4817_), .B1(new_n3398_), .B2(new_n3390_), .ZN(new_n4821_));
  NAND3_X1   g03819(.A1(new_n3389_), .A2(new_n4814_), .A3(new_n4812_), .ZN(new_n4822_));
  AOI22_X1   g03820(.A1(new_n3362_), .A2(new_n3366_), .B1(new_n3371_), .B2(new_n3375_), .ZN(new_n4823_));
  NOR3_X1    g03821(.A1(new_n4823_), .A2(new_n4816_), .A3(new_n4818_), .ZN(new_n4824_));
  NAND3_X1   g03822(.A1(new_n4824_), .A2(new_n3357_), .A3(new_n4822_), .ZN(new_n4825_));
  AOI21_X1   g03823(.A1(new_n4821_), .A2(new_n4825_), .B(new_n4809_), .ZN(new_n4826_));
  XOR2_X1    g03824(.A1(new_n3396_), .A2(new_n4808_), .Z(new_n4827_));
  NOR2_X1    g03825(.A1(new_n4823_), .A2(new_n4818_), .ZN(new_n4828_));
  NAND2_X1   g03826(.A1(new_n4819_), .A2(new_n4818_), .ZN(new_n4829_));
  NAND2_X1   g03827(.A1(new_n4816_), .A2(new_n3376_), .ZN(new_n4830_));
  AOI22_X1   g03828(.A1(new_n4829_), .A2(new_n4830_), .B1(new_n3357_), .B2(new_n4828_), .ZN(new_n4831_));
  NAND4_X1   g03829(.A1(new_n3396_), .A2(new_n3397_), .A3(new_n3389_), .A4(new_n3376_), .ZN(new_n4832_));
  NOR3_X1    g03830(.A1(new_n4832_), .A2(new_n4817_), .A3(new_n4820_), .ZN(new_n4833_));
  NOR3_X1    g03831(.A1(new_n4831_), .A2(new_n4833_), .A3(new_n4827_), .ZN(new_n4834_));
  OAI22_X1   g03832(.A1(new_n3344_), .A2(new_n3356_), .B1(new_n4823_), .B2(new_n4818_), .ZN(new_n4835_));
  NAND2_X1   g03833(.A1(new_n4835_), .A2(new_n4832_), .ZN(new_n4836_));
  AOI21_X1   g03834(.A1(new_n3316_), .A2(new_n3323_), .B(new_n4836_), .ZN(new_n4837_));
  OAI21_X1   g03835(.A1(new_n4826_), .A2(new_n4834_), .B(new_n4837_), .ZN(new_n4838_));
  INV_X1     g03836(.I(new_n4814_), .ZN(new_n4839_));
  INV_X1     g03837(.I(new_n4812_), .ZN(new_n4840_));
  NOR3_X1    g03838(.A1(new_n4823_), .A2(new_n4839_), .A3(new_n4840_), .ZN(new_n4841_));
  NAND3_X1   g03839(.A1(new_n4819_), .A2(new_n3376_), .A3(new_n3389_), .ZN(new_n4842_));
  NOR3_X1    g03840(.A1(new_n4842_), .A2(new_n4841_), .A3(new_n3398_), .ZN(new_n4843_));
  OAI21_X1   g03841(.A1(new_n4831_), .A2(new_n4843_), .B(new_n4827_), .ZN(new_n4844_));
  NAND4_X1   g03842(.A1(new_n3357_), .A2(new_n3376_), .A3(new_n3389_), .A4(new_n4819_), .ZN(new_n4845_));
  NAND3_X1   g03843(.A1(new_n4821_), .A2(new_n4809_), .A3(new_n4845_), .ZN(new_n4846_));
  NOR4_X1    g03844(.A1(new_n3344_), .A2(new_n3356_), .A3(new_n4823_), .A4(new_n4818_), .ZN(new_n4847_));
  AOI22_X1   g03845(.A1(new_n3396_), .A2(new_n3397_), .B1(new_n3389_), .B2(new_n3376_), .ZN(new_n4848_));
  NOR2_X1    g03846(.A1(new_n4847_), .A2(new_n4848_), .ZN(new_n4849_));
  OAI21_X1   g03847(.A1(new_n3393_), .A2(new_n3394_), .B(new_n4849_), .ZN(new_n4850_));
  NAND3_X1   g03848(.A1(new_n4850_), .A2(new_n4844_), .A3(new_n4846_), .ZN(new_n4851_));
  AOI21_X1   g03849(.A1(new_n4838_), .A2(new_n4851_), .B(new_n4802_), .ZN(new_n4852_));
  INV_X1     g03850(.I(new_n4785_), .ZN(new_n4853_));
  INV_X1     g03851(.I(new_n4783_), .ZN(new_n4854_));
  NOR3_X1    g03852(.A1(new_n3321_), .A2(new_n4853_), .A3(new_n4854_), .ZN(new_n4855_));
  NAND3_X1   g03853(.A1(new_n4789_), .A2(new_n3303_), .A3(new_n3314_), .ZN(new_n4856_));
  NOR3_X1    g03854(.A1(new_n4856_), .A2(new_n4855_), .A3(new_n3319_), .ZN(new_n4857_));
  NOR3_X1    g03855(.A1(new_n4796_), .A2(new_n4799_), .A3(new_n4857_), .ZN(new_n4858_));
  NAND4_X1   g03856(.A1(new_n3282_), .A2(new_n3303_), .A3(new_n3314_), .A4(new_n4789_), .ZN(new_n4859_));
  AOI21_X1   g03857(.A1(new_n4791_), .A2(new_n4859_), .B(new_n4780_), .ZN(new_n4860_));
  NOR2_X1    g03858(.A1(new_n4858_), .A2(new_n4860_), .ZN(new_n4861_));
  AOI21_X1   g03859(.A1(new_n4844_), .A2(new_n4846_), .B(new_n4850_), .ZN(new_n4862_));
  NOR3_X1    g03860(.A1(new_n4837_), .A2(new_n4834_), .A3(new_n4826_), .ZN(new_n4863_));
  NOR3_X1    g03861(.A1(new_n4862_), .A2(new_n4863_), .A3(new_n4861_), .ZN(new_n4864_));
  NOR2_X1    g03862(.A1(new_n4864_), .A2(new_n4852_), .ZN(new_n4865_));
  AOI21_X1   g03863(.A1(\A[383] ), .A2(\A[384] ), .B(\A[382] ), .ZN(new_n4866_));
  AOI21_X1   g03864(.A1(\A[380] ), .A2(\A[381] ), .B(\A[379] ), .ZN(new_n4867_));
  OAI22_X1   g03865(.A1(new_n3131_), .A2(new_n4867_), .B1(new_n4866_), .B2(new_n3140_), .ZN(new_n4868_));
  NOR2_X1    g03866(.A1(new_n4866_), .A2(new_n3140_), .ZN(new_n4869_));
  NOR2_X1    g03867(.A1(new_n4867_), .A2(new_n3131_), .ZN(new_n4870_));
  NAND2_X1   g03868(.A1(new_n4869_), .A2(new_n4870_), .ZN(new_n4871_));
  NAND2_X1   g03869(.A1(new_n4871_), .A2(new_n4868_), .ZN(new_n4872_));
  NOR2_X1    g03870(.A1(new_n3162_), .A2(new_n4872_), .ZN(new_n4873_));
  NOR2_X1    g03871(.A1(new_n4869_), .A2(new_n4870_), .ZN(new_n4874_));
  NOR4_X1    g03872(.A1(new_n4866_), .A2(new_n4867_), .A3(new_n3131_), .A4(new_n3140_), .ZN(new_n4875_));
  NOR2_X1    g03873(.A1(new_n4874_), .A2(new_n4875_), .ZN(new_n4876_));
  NOR2_X1    g03874(.A1(new_n3142_), .A2(new_n4876_), .ZN(new_n4877_));
  NOR2_X1    g03875(.A1(new_n4877_), .A2(new_n4873_), .ZN(new_n4878_));
  AOI21_X1   g03876(.A1(\A[389] ), .A2(\A[390] ), .B(\A[388] ), .ZN(new_n4879_));
  NOR2_X1    g03877(.A1(new_n4879_), .A2(new_n3106_), .ZN(new_n4880_));
  AOI21_X1   g03878(.A1(\A[386] ), .A2(\A[387] ), .B(\A[385] ), .ZN(new_n4881_));
  NOR2_X1    g03879(.A1(new_n4881_), .A2(new_n3096_), .ZN(new_n4882_));
  XOR2_X1    g03880(.A1(new_n4880_), .A2(new_n4882_), .Z(new_n4883_));
  NOR2_X1    g03881(.A1(new_n4883_), .A2(new_n3110_), .ZN(new_n4884_));
  NOR3_X1    g03882(.A1(new_n4882_), .A2(new_n3106_), .A3(new_n4879_), .ZN(new_n4885_));
  NOR3_X1    g03883(.A1(new_n4880_), .A2(new_n3096_), .A3(new_n4881_), .ZN(new_n4886_));
  NOR2_X1    g03884(.A1(new_n4885_), .A2(new_n4886_), .ZN(new_n4887_));
  NOR2_X1    g03885(.A1(new_n4887_), .A2(new_n3148_), .ZN(new_n4888_));
  OAI22_X1   g03886(.A1(new_n3146_), .A2(new_n3150_), .B1(new_n4884_), .B2(new_n4888_), .ZN(new_n4889_));
  NAND2_X1   g03887(.A1(new_n4887_), .A2(new_n3148_), .ZN(new_n4890_));
  NAND2_X1   g03888(.A1(new_n4883_), .A2(new_n3110_), .ZN(new_n4891_));
  NOR4_X1    g03889(.A1(new_n3165_), .A2(new_n3110_), .A3(new_n3121_), .A4(new_n3162_), .ZN(new_n4892_));
  NAND3_X1   g03890(.A1(new_n4892_), .A2(new_n4890_), .A3(new_n4891_), .ZN(new_n4893_));
  NAND3_X1   g03891(.A1(new_n4893_), .A2(new_n4889_), .A3(new_n4878_), .ZN(new_n4894_));
  NAND2_X1   g03892(.A1(new_n3142_), .A2(new_n4876_), .ZN(new_n4895_));
  NAND2_X1   g03893(.A1(new_n3162_), .A2(new_n4872_), .ZN(new_n4896_));
  NAND2_X1   g03894(.A1(new_n4895_), .A2(new_n4896_), .ZN(new_n4897_));
  NOR2_X1    g03895(.A1(new_n4884_), .A2(new_n4888_), .ZN(new_n4898_));
  NOR2_X1    g03896(.A1(new_n4898_), .A2(new_n4892_), .ZN(new_n4899_));
  NOR4_X1    g03897(.A1(new_n3146_), .A2(new_n3110_), .A3(new_n3121_), .A4(new_n4887_), .ZN(new_n4900_));
  OAI21_X1   g03898(.A1(new_n4899_), .A2(new_n4900_), .B(new_n4897_), .ZN(new_n4901_));
  NAND2_X1   g03899(.A1(new_n4901_), .A2(new_n4894_), .ZN(new_n4902_));
  AOI21_X1   g03900(.A1(\A[371] ), .A2(\A[372] ), .B(\A[370] ), .ZN(new_n4903_));
  NOR2_X1    g03901(.A1(new_n4903_), .A2(new_n3219_), .ZN(new_n4904_));
  AOI21_X1   g03902(.A1(\A[368] ), .A2(\A[369] ), .B(\A[367] ), .ZN(new_n4905_));
  NOR2_X1    g03903(.A1(new_n4905_), .A2(new_n3209_), .ZN(new_n4906_));
  NOR2_X1    g03904(.A1(new_n4904_), .A2(new_n4906_), .ZN(new_n4907_));
  NOR4_X1    g03905(.A1(new_n4903_), .A2(new_n4905_), .A3(new_n3209_), .A4(new_n3219_), .ZN(new_n4908_));
  NOR2_X1    g03906(.A1(new_n4907_), .A2(new_n4908_), .ZN(new_n4909_));
  NAND2_X1   g03907(.A1(new_n3221_), .A2(new_n4909_), .ZN(new_n4910_));
  NOR2_X1    g03908(.A1(new_n3226_), .A2(new_n3224_), .ZN(new_n4911_));
  NOR2_X1    g03909(.A1(new_n3229_), .A2(new_n3231_), .ZN(new_n4912_));
  OAI22_X1   g03910(.A1(new_n3209_), .A2(new_n4905_), .B1(new_n4903_), .B2(new_n3219_), .ZN(new_n4913_));
  NAND2_X1   g03911(.A1(new_n3217_), .A2(new_n3216_), .ZN(new_n4914_));
  NAND2_X1   g03912(.A1(new_n3207_), .A2(new_n3206_), .ZN(new_n4915_));
  NAND4_X1   g03913(.A1(new_n4914_), .A2(new_n4915_), .A3(new_n3225_), .A4(new_n3230_), .ZN(new_n4916_));
  NAND2_X1   g03914(.A1(new_n4916_), .A2(new_n4913_), .ZN(new_n4917_));
  NAND3_X1   g03915(.A1(new_n4917_), .A2(new_n4911_), .A3(new_n4912_), .ZN(new_n4918_));
  NAND2_X1   g03916(.A1(new_n4910_), .A2(new_n4918_), .ZN(new_n4919_));
  AOI21_X1   g03917(.A1(\A[377] ), .A2(\A[378] ), .B(\A[376] ), .ZN(new_n4920_));
  AOI21_X1   g03918(.A1(\A[374] ), .A2(\A[375] ), .B(\A[373] ), .ZN(new_n4921_));
  NOR2_X1    g03919(.A1(new_n4921_), .A2(new_n3174_), .ZN(new_n4922_));
  NOR3_X1    g03920(.A1(new_n4922_), .A2(new_n3184_), .A3(new_n4920_), .ZN(new_n4923_));
  NOR2_X1    g03921(.A1(new_n4920_), .A2(new_n3184_), .ZN(new_n4924_));
  NOR3_X1    g03922(.A1(new_n4924_), .A2(new_n3174_), .A3(new_n4921_), .ZN(new_n4925_));
  NOR3_X1    g03923(.A1(new_n3188_), .A2(new_n4923_), .A3(new_n4925_), .ZN(new_n4926_));
  NOR2_X1    g03924(.A1(new_n4923_), .A2(new_n4925_), .ZN(new_n4927_));
  NOR2_X1    g03925(.A1(new_n4927_), .A2(new_n3235_), .ZN(new_n4928_));
  NAND4_X1   g03926(.A1(new_n3236_), .A2(new_n3221_), .A3(new_n3232_), .A4(new_n3235_), .ZN(new_n4929_));
  OAI21_X1   g03927(.A1(new_n4926_), .A2(new_n4928_), .B(new_n4929_), .ZN(new_n4930_));
  NAND2_X1   g03928(.A1(new_n4927_), .A2(new_n3235_), .ZN(new_n4931_));
  XOR2_X1    g03929(.A1(new_n4924_), .A2(new_n4922_), .Z(new_n4932_));
  NAND2_X1   g03930(.A1(new_n4932_), .A2(new_n3188_), .ZN(new_n4933_));
  NOR4_X1    g03931(.A1(new_n3188_), .A2(new_n3239_), .A3(new_n3199_), .A4(new_n3238_), .ZN(new_n4934_));
  NAND3_X1   g03932(.A1(new_n4934_), .A2(new_n4931_), .A3(new_n4933_), .ZN(new_n4935_));
  NAND3_X1   g03933(.A1(new_n4930_), .A2(new_n4935_), .A3(new_n4919_), .ZN(new_n4936_));
  NOR2_X1    g03934(.A1(new_n3238_), .A2(new_n4917_), .ZN(new_n4937_));
  NOR2_X1    g03935(.A1(new_n3221_), .A2(new_n4909_), .ZN(new_n4938_));
  NOR2_X1    g03936(.A1(new_n4938_), .A2(new_n4937_), .ZN(new_n4939_));
  NOR2_X1    g03937(.A1(new_n4926_), .A2(new_n4928_), .ZN(new_n4940_));
  NOR2_X1    g03938(.A1(new_n4940_), .A2(new_n4934_), .ZN(new_n4941_));
  NOR3_X1    g03939(.A1(new_n4929_), .A2(new_n4926_), .A3(new_n4928_), .ZN(new_n4942_));
  OAI21_X1   g03940(.A1(new_n4941_), .A2(new_n4942_), .B(new_n4939_), .ZN(new_n4943_));
  NAND3_X1   g03941(.A1(new_n4943_), .A2(new_n4936_), .A3(new_n3242_), .ZN(new_n4944_));
  OAI22_X1   g03942(.A1(new_n3243_), .A2(new_n3244_), .B1(new_n3246_), .B2(new_n3245_), .ZN(new_n4945_));
  OAI21_X1   g03943(.A1(new_n4940_), .A2(new_n4934_), .B(new_n4919_), .ZN(new_n4946_));
  NOR2_X1    g03944(.A1(new_n4946_), .A2(new_n4942_), .ZN(new_n4947_));
  AOI21_X1   g03945(.A1(new_n4930_), .A2(new_n4935_), .B(new_n4919_), .ZN(new_n4948_));
  OAI21_X1   g03946(.A1(new_n4947_), .A2(new_n4948_), .B(new_n4945_), .ZN(new_n4949_));
  NAND3_X1   g03947(.A1(new_n4949_), .A2(new_n4944_), .A3(new_n4902_), .ZN(new_n4950_));
  NOR3_X1    g03948(.A1(new_n4899_), .A2(new_n4897_), .A3(new_n4900_), .ZN(new_n4951_));
  AOI21_X1   g03949(.A1(new_n4893_), .A2(new_n4889_), .B(new_n4878_), .ZN(new_n4952_));
  NOR2_X1    g03950(.A1(new_n4951_), .A2(new_n4952_), .ZN(new_n4953_));
  NOR3_X1    g03951(.A1(new_n4947_), .A2(new_n4948_), .A3(new_n4945_), .ZN(new_n4954_));
  AOI21_X1   g03952(.A1(new_n4943_), .A2(new_n4936_), .B(new_n3242_), .ZN(new_n4955_));
  OAI21_X1   g03953(.A1(new_n4954_), .A2(new_n4955_), .B(new_n4953_), .ZN(new_n4956_));
  AOI21_X1   g03954(.A1(new_n4956_), .A2(new_n4950_), .B(new_n3402_), .ZN(new_n4957_));
  NAND2_X1   g03955(.A1(new_n3405_), .A2(new_n3248_), .ZN(new_n4958_));
  NOR3_X1    g03956(.A1(new_n4954_), .A2(new_n4955_), .A3(new_n4953_), .ZN(new_n4959_));
  AOI21_X1   g03957(.A1(new_n4949_), .A2(new_n4944_), .B(new_n4902_), .ZN(new_n4960_));
  NOR3_X1    g03958(.A1(new_n4959_), .A2(new_n4960_), .A3(new_n4958_), .ZN(new_n4961_));
  NOR3_X1    g03959(.A1(new_n4957_), .A2(new_n4961_), .A3(new_n4865_), .ZN(new_n4962_));
  OAI21_X1   g03960(.A1(new_n4957_), .A2(new_n4961_), .B(new_n4865_), .ZN(new_n4963_));
  INV_X1     g03961(.I(new_n4963_), .ZN(new_n4964_));
  NOR2_X1    g03962(.A1(new_n4964_), .A2(new_n4962_), .ZN(new_n4965_));
  AOI21_X1   g03963(.A1(\A[431] ), .A2(\A[432] ), .B(\A[430] ), .ZN(new_n4966_));
  NOR2_X1    g03964(.A1(new_n4966_), .A2(new_n3671_), .ZN(new_n4967_));
  AOI21_X1   g03965(.A1(\A[428] ), .A2(\A[429] ), .B(\A[427] ), .ZN(new_n4968_));
  NOR2_X1    g03966(.A1(new_n4968_), .A2(new_n3661_), .ZN(new_n4969_));
  NOR2_X1    g03967(.A1(new_n4967_), .A2(new_n4969_), .ZN(new_n4970_));
  NOR4_X1    g03968(.A1(new_n4966_), .A2(new_n4968_), .A3(new_n3661_), .A4(new_n3671_), .ZN(new_n4971_));
  NOR2_X1    g03969(.A1(new_n4970_), .A2(new_n4971_), .ZN(new_n4972_));
  NAND2_X1   g03970(.A1(new_n3719_), .A2(new_n4972_), .ZN(new_n4973_));
  OAI22_X1   g03971(.A1(new_n3661_), .A2(new_n4968_), .B1(new_n4966_), .B2(new_n3671_), .ZN(new_n4974_));
  INV_X1     g03972(.I(new_n4971_), .ZN(new_n4975_));
  NAND2_X1   g03973(.A1(new_n4975_), .A2(new_n4974_), .ZN(new_n4976_));
  NAND2_X1   g03974(.A1(new_n3674_), .A2(new_n4976_), .ZN(new_n4977_));
  NAND2_X1   g03975(.A1(new_n4977_), .A2(new_n4973_), .ZN(new_n4978_));
  NOR4_X1    g03976(.A1(new_n3674_), .A2(new_n3685_), .A3(new_n3706_), .A4(new_n3717_), .ZN(new_n4979_));
  NAND2_X1   g03977(.A1(new_n3709_), .A2(new_n3711_), .ZN(new_n4980_));
  NAND2_X1   g03978(.A1(new_n3714_), .A2(new_n3716_), .ZN(new_n4981_));
  AOI21_X1   g03979(.A1(\A[437] ), .A2(\A[438] ), .B(\A[436] ), .ZN(new_n4982_));
  AOI21_X1   g03980(.A1(\A[434] ), .A2(\A[435] ), .B(\A[433] ), .ZN(new_n4983_));
  NOR2_X1    g03981(.A1(new_n4983_), .A2(new_n3693_), .ZN(new_n4984_));
  NOR3_X1    g03982(.A1(new_n4984_), .A2(new_n3703_), .A3(new_n4982_), .ZN(new_n4985_));
  NOR2_X1    g03983(.A1(new_n4982_), .A2(new_n3703_), .ZN(new_n4986_));
  NOR3_X1    g03984(.A1(new_n4986_), .A2(new_n3693_), .A3(new_n4983_), .ZN(new_n4987_));
  OAI22_X1   g03985(.A1(new_n4980_), .A2(new_n4981_), .B1(new_n4985_), .B2(new_n4987_), .ZN(new_n4988_));
  NOR2_X1    g03986(.A1(new_n4985_), .A2(new_n4987_), .ZN(new_n4989_));
  NAND2_X1   g03987(.A1(new_n3706_), .A2(new_n4989_), .ZN(new_n4990_));
  NAND2_X1   g03988(.A1(new_n4990_), .A2(new_n4988_), .ZN(new_n4991_));
  NOR2_X1    g03989(.A1(new_n4991_), .A2(new_n4979_), .ZN(new_n4992_));
  NOR2_X1    g03990(.A1(new_n3695_), .A2(new_n3691_), .ZN(new_n4993_));
  NOR2_X1    g03991(.A1(new_n3705_), .A2(new_n3701_), .ZN(new_n4994_));
  OAI21_X1   g03992(.A1(new_n3693_), .A2(new_n4983_), .B(new_n4986_), .ZN(new_n4995_));
  OAI21_X1   g03993(.A1(new_n3703_), .A2(new_n4982_), .B(new_n4984_), .ZN(new_n4996_));
  AOI22_X1   g03994(.A1(new_n4993_), .A2(new_n4994_), .B1(new_n4995_), .B2(new_n4996_), .ZN(new_n4997_));
  NOR4_X1    g03995(.A1(new_n4980_), .A2(new_n4981_), .A3(new_n4985_), .A4(new_n4987_), .ZN(new_n4998_));
  NOR2_X1    g03996(.A1(new_n4997_), .A2(new_n4998_), .ZN(new_n4999_));
  NOR2_X1    g03997(.A1(new_n4999_), .A2(new_n3723_), .ZN(new_n5000_));
  NOR3_X1    g03998(.A1(new_n4992_), .A2(new_n5000_), .A3(new_n4978_), .ZN(new_n5001_));
  AND2_X2    g03999(.A1(new_n4977_), .A2(new_n4973_), .Z(new_n5002_));
  NAND2_X1   g04000(.A1(new_n4999_), .A2(new_n3723_), .ZN(new_n5003_));
  NAND2_X1   g04001(.A1(new_n4986_), .A2(new_n4984_), .ZN(new_n5004_));
  INV_X1     g04002(.I(new_n5004_), .ZN(new_n5005_));
  NAND2_X1   g04003(.A1(new_n3722_), .A2(new_n5005_), .ZN(new_n5006_));
  NOR3_X1    g04004(.A1(new_n4989_), .A2(new_n3706_), .A3(new_n3717_), .ZN(new_n5007_));
  NAND4_X1   g04005(.A1(new_n5007_), .A2(new_n3719_), .A3(new_n5006_), .A4(new_n3720_), .ZN(new_n5008_));
  AOI21_X1   g04006(.A1(new_n5003_), .A2(new_n5008_), .B(new_n5002_), .ZN(new_n5009_));
  NOR2_X1    g04007(.A1(new_n5001_), .A2(new_n5009_), .ZN(new_n5010_));
  AOI21_X1   g04008(.A1(\A[419] ), .A2(\A[420] ), .B(\A[418] ), .ZN(new_n5011_));
  AOI21_X1   g04009(.A1(\A[416] ), .A2(\A[417] ), .B(\A[415] ), .ZN(new_n5012_));
  OAI22_X1   g04010(.A1(new_n3618_), .A2(new_n5012_), .B1(new_n5011_), .B2(new_n3640_), .ZN(new_n5013_));
  NOR2_X1    g04011(.A1(new_n5011_), .A2(new_n3640_), .ZN(new_n5014_));
  NOR2_X1    g04012(.A1(new_n5012_), .A2(new_n3618_), .ZN(new_n5015_));
  NAND2_X1   g04013(.A1(new_n5014_), .A2(new_n5015_), .ZN(new_n5016_));
  NAND2_X1   g04014(.A1(new_n5016_), .A2(new_n5013_), .ZN(new_n5017_));
  NOR2_X1    g04015(.A1(new_n3630_), .A2(new_n5017_), .ZN(new_n5018_));
  NOR2_X1    g04016(.A1(new_n5014_), .A2(new_n5015_), .ZN(new_n5019_));
  NOR4_X1    g04017(.A1(new_n5011_), .A2(new_n5012_), .A3(new_n3618_), .A4(new_n3640_), .ZN(new_n5020_));
  NOR2_X1    g04018(.A1(new_n5019_), .A2(new_n5020_), .ZN(new_n5021_));
  NOR2_X1    g04019(.A1(new_n3648_), .A2(new_n5021_), .ZN(new_n5022_));
  NOR2_X1    g04020(.A1(new_n5022_), .A2(new_n5018_), .ZN(new_n5023_));
  AOI21_X1   g04021(.A1(\A[425] ), .A2(\A[426] ), .B(\A[424] ), .ZN(new_n5024_));
  AOI21_X1   g04022(.A1(\A[422] ), .A2(\A[423] ), .B(\A[421] ), .ZN(new_n5025_));
  NOR2_X1    g04023(.A1(new_n5025_), .A2(new_n3584_), .ZN(new_n5026_));
  NOR3_X1    g04024(.A1(new_n5026_), .A2(new_n3594_), .A3(new_n5024_), .ZN(new_n5027_));
  NOR2_X1    g04025(.A1(new_n5024_), .A2(new_n3594_), .ZN(new_n5028_));
  NOR3_X1    g04026(.A1(new_n5028_), .A2(new_n3584_), .A3(new_n5025_), .ZN(new_n5029_));
  NOR2_X1    g04027(.A1(new_n5027_), .A2(new_n5029_), .ZN(new_n5030_));
  NAND2_X1   g04028(.A1(new_n5030_), .A2(new_n3597_), .ZN(new_n5031_));
  XOR2_X1    g04029(.A1(new_n5028_), .A2(new_n5026_), .Z(new_n5032_));
  NAND2_X1   g04030(.A1(new_n5032_), .A2(new_n3645_), .ZN(new_n5033_));
  AOI22_X1   g04031(.A1(new_n5031_), .A2(new_n5033_), .B1(new_n3647_), .B2(new_n3643_), .ZN(new_n5034_));
  NAND3_X1   g04032(.A1(new_n5032_), .A2(new_n3609_), .A3(new_n3597_), .ZN(new_n5035_));
  NOR2_X1    g04033(.A1(new_n5028_), .A2(new_n5026_), .ZN(new_n5036_));
  NAND2_X1   g04034(.A1(new_n5028_), .A2(new_n5026_), .ZN(new_n5037_));
  AOI21_X1   g04035(.A1(new_n3597_), .A2(new_n5037_), .B(new_n5036_), .ZN(new_n5038_));
  NOR3_X1    g04036(.A1(new_n5035_), .A2(new_n3650_), .A3(new_n5038_), .ZN(new_n5039_));
  NOR3_X1    g04037(.A1(new_n5034_), .A2(new_n5023_), .A3(new_n5039_), .ZN(new_n5040_));
  NAND2_X1   g04038(.A1(new_n3648_), .A2(new_n5021_), .ZN(new_n5041_));
  NOR2_X1    g04039(.A1(new_n3620_), .A2(new_n3616_), .ZN(new_n5042_));
  NOR2_X1    g04040(.A1(new_n3626_), .A2(new_n3629_), .ZN(new_n5043_));
  NAND3_X1   g04041(.A1(new_n5017_), .A2(new_n5042_), .A3(new_n5043_), .ZN(new_n5044_));
  NAND2_X1   g04042(.A1(new_n5041_), .A2(new_n5044_), .ZN(new_n5045_));
  NOR2_X1    g04043(.A1(new_n5032_), .A2(new_n3645_), .ZN(new_n5046_));
  NOR2_X1    g04044(.A1(new_n5030_), .A2(new_n3597_), .ZN(new_n5047_));
  OAI22_X1   g04045(.A1(new_n5046_), .A2(new_n5047_), .B1(new_n3650_), .B2(new_n3610_), .ZN(new_n5048_));
  NOR4_X1    g04046(.A1(new_n3650_), .A2(new_n3645_), .A3(new_n3646_), .A4(new_n5030_), .ZN(new_n5049_));
  INV_X1     g04047(.I(new_n5049_), .ZN(new_n5050_));
  AOI21_X1   g04048(.A1(new_n5050_), .A2(new_n5048_), .B(new_n5045_), .ZN(new_n5051_));
  NOR3_X1    g04049(.A1(new_n3727_), .A2(new_n5051_), .A3(new_n5040_), .ZN(new_n5052_));
  NOR3_X1    g04050(.A1(new_n3645_), .A2(new_n5030_), .A3(new_n3646_), .ZN(new_n5053_));
  INV_X1     g04051(.I(new_n5036_), .ZN(new_n5054_));
  NAND2_X1   g04052(.A1(new_n3597_), .A2(new_n5037_), .ZN(new_n5055_));
  NAND2_X1   g04053(.A1(new_n5055_), .A2(new_n5054_), .ZN(new_n5056_));
  NAND3_X1   g04054(.A1(new_n5056_), .A2(new_n3643_), .A3(new_n5053_), .ZN(new_n5057_));
  NAND3_X1   g04055(.A1(new_n5057_), .A2(new_n5048_), .A3(new_n5045_), .ZN(new_n5058_));
  OAI21_X1   g04056(.A1(new_n5034_), .A2(new_n5049_), .B(new_n5023_), .ZN(new_n5059_));
  AOI21_X1   g04057(.A1(new_n5058_), .A2(new_n5059_), .B(new_n3731_), .ZN(new_n5060_));
  NOR3_X1    g04058(.A1(new_n5052_), .A2(new_n5060_), .A3(new_n5010_), .ZN(new_n5061_));
  OAI21_X1   g04059(.A1(new_n5052_), .A2(new_n5060_), .B(new_n5010_), .ZN(new_n5062_));
  INV_X1     g04060(.I(new_n5062_), .ZN(new_n5063_));
  NOR2_X1    g04061(.A1(new_n5063_), .A2(new_n5061_), .ZN(new_n5064_));
  NAND2_X1   g04062(.A1(new_n3576_), .A2(new_n3732_), .ZN(new_n5065_));
  NOR4_X1    g04063(.A1(new_n3529_), .A2(new_n3533_), .A3(new_n3557_), .A4(new_n3555_), .ZN(new_n5066_));
  AOI21_X1   g04064(.A1(\A[443] ), .A2(\A[444] ), .B(\A[442] ), .ZN(new_n5067_));
  AOI21_X1   g04065(.A1(\A[440] ), .A2(\A[441] ), .B(\A[439] ), .ZN(new_n5068_));
  OAI22_X1   g04066(.A1(new_n3531_), .A2(new_n5068_), .B1(new_n5067_), .B2(new_n3543_), .ZN(new_n5069_));
  NOR4_X1    g04067(.A1(new_n5067_), .A2(new_n5068_), .A3(new_n3531_), .A4(new_n3543_), .ZN(new_n5070_));
  INV_X1     g04068(.I(new_n5070_), .ZN(new_n5071_));
  NAND2_X1   g04069(.A1(new_n5071_), .A2(new_n5069_), .ZN(new_n5072_));
  XOR2_X1    g04070(.A1(new_n5066_), .A2(new_n5072_), .Z(new_n5073_));
  NOR4_X1    g04071(.A1(new_n3493_), .A2(new_n3497_), .A3(new_n3521_), .A4(new_n3519_), .ZN(new_n5074_));
  AOI21_X1   g04072(.A1(\A[449] ), .A2(\A[450] ), .B(\A[448] ), .ZN(new_n5075_));
  AOI21_X1   g04073(.A1(\A[446] ), .A2(\A[447] ), .B(\A[445] ), .ZN(new_n5076_));
  NOR2_X1    g04074(.A1(new_n5076_), .A2(new_n3495_), .ZN(new_n5077_));
  NOR3_X1    g04075(.A1(new_n5077_), .A2(new_n3507_), .A3(new_n5075_), .ZN(new_n5078_));
  NOR2_X1    g04076(.A1(new_n5075_), .A2(new_n3507_), .ZN(new_n5079_));
  NOR3_X1    g04077(.A1(new_n5079_), .A2(new_n3495_), .A3(new_n5076_), .ZN(new_n5080_));
  NOR2_X1    g04078(.A1(new_n5078_), .A2(new_n5080_), .ZN(new_n5081_));
  XOR2_X1    g04079(.A1(new_n5074_), .A2(new_n5081_), .Z(new_n5082_));
  AOI21_X1   g04080(.A1(new_n3567_), .A2(new_n5082_), .B(new_n5073_), .ZN(new_n5083_));
  NOR3_X1    g04081(.A1(new_n5074_), .A2(new_n5078_), .A3(new_n5080_), .ZN(new_n5084_));
  NAND4_X1   g04082(.A1(new_n3513_), .A2(new_n3515_), .A3(new_n3503_), .A4(new_n3508_), .ZN(new_n5085_));
  NOR2_X1    g04083(.A1(new_n5085_), .A2(new_n5081_), .ZN(new_n5086_));
  NOR2_X1    g04084(.A1(new_n5084_), .A2(new_n5086_), .ZN(new_n5087_));
  NAND2_X1   g04085(.A1(new_n3516_), .A2(new_n3509_), .ZN(new_n5088_));
  NAND3_X1   g04086(.A1(new_n5088_), .A2(new_n5079_), .A3(new_n5077_), .ZN(new_n5089_));
  NAND4_X1   g04087(.A1(new_n5087_), .A2(new_n3561_), .A3(new_n3562_), .A4(new_n5089_), .ZN(new_n5090_));
  OAI22_X1   g04088(.A1(new_n3570_), .A2(new_n3573_), .B1(new_n5084_), .B2(new_n5086_), .ZN(new_n5091_));
  NAND2_X1   g04089(.A1(new_n5087_), .A2(new_n3560_), .ZN(new_n5092_));
  NAND2_X1   g04090(.A1(new_n5092_), .A2(new_n5091_), .ZN(new_n5093_));
  AOI22_X1   g04091(.A1(new_n5093_), .A2(new_n5073_), .B1(new_n5083_), .B2(new_n5090_), .ZN(new_n5094_));
  NAND4_X1   g04092(.A1(new_n3565_), .A2(new_n3566_), .A3(new_n3574_), .A4(new_n3567_), .ZN(new_n5095_));
  NAND4_X1   g04093(.A1(new_n3470_), .A2(new_n3460_), .A3(new_n3465_), .A4(new_n3472_), .ZN(new_n5096_));
  AOI21_X1   g04094(.A1(\A[455] ), .A2(\A[456] ), .B(\A[454] ), .ZN(new_n5097_));
  NOR2_X1    g04095(.A1(new_n5097_), .A2(new_n3464_), .ZN(new_n5098_));
  AOI21_X1   g04096(.A1(\A[452] ), .A2(\A[453] ), .B(\A[451] ), .ZN(new_n5099_));
  NOR2_X1    g04097(.A1(new_n5099_), .A2(new_n3452_), .ZN(new_n5100_));
  NOR2_X1    g04098(.A1(new_n5098_), .A2(new_n5100_), .ZN(new_n5101_));
  NOR4_X1    g04099(.A1(new_n5097_), .A2(new_n5099_), .A3(new_n3452_), .A4(new_n3464_), .ZN(new_n5102_));
  NOR2_X1    g04100(.A1(new_n5101_), .A2(new_n5102_), .ZN(new_n5103_));
  XNOR2_X1   g04101(.A1(new_n5096_), .A2(new_n5103_), .ZN(new_n5104_));
  NAND4_X1   g04102(.A1(new_n3432_), .A2(new_n3423_), .A3(new_n3434_), .A4(new_n3427_), .ZN(new_n5105_));
  AOI21_X1   g04103(.A1(\A[461] ), .A2(\A[462] ), .B(\A[460] ), .ZN(new_n5106_));
  AOI21_X1   g04104(.A1(\A[458] ), .A2(\A[459] ), .B(\A[457] ), .ZN(new_n5107_));
  NOR2_X1    g04105(.A1(new_n5107_), .A2(new_n3415_), .ZN(new_n5108_));
  NOR3_X1    g04106(.A1(new_n5108_), .A2(new_n3426_), .A3(new_n5106_), .ZN(new_n5109_));
  NOR2_X1    g04107(.A1(new_n5106_), .A2(new_n3426_), .ZN(new_n5110_));
  NOR3_X1    g04108(.A1(new_n5110_), .A2(new_n3415_), .A3(new_n5107_), .ZN(new_n5111_));
  NOR2_X1    g04109(.A1(new_n5109_), .A2(new_n5111_), .ZN(new_n5112_));
  NAND2_X1   g04110(.A1(new_n5112_), .A2(new_n5105_), .ZN(new_n5113_));
  NOR4_X1    g04111(.A1(new_n3413_), .A2(new_n3417_), .A3(new_n3441_), .A4(new_n3438_), .ZN(new_n5114_));
  XOR2_X1    g04112(.A1(new_n5110_), .A2(new_n5108_), .Z(new_n5115_));
  NAND2_X1   g04113(.A1(new_n5115_), .A2(new_n5114_), .ZN(new_n5116_));
  AOI22_X1   g04114(.A1(new_n3444_), .A2(new_n3481_), .B1(new_n5113_), .B2(new_n5116_), .ZN(new_n5117_));
  NAND2_X1   g04115(.A1(new_n5116_), .A2(new_n5113_), .ZN(new_n5118_));
  INV_X1     g04116(.I(new_n5110_), .ZN(new_n5119_));
  INV_X1     g04117(.I(new_n5108_), .ZN(new_n5120_));
  NOR2_X1    g04118(.A1(new_n3418_), .A2(new_n3442_), .ZN(new_n5121_));
  NOR3_X1    g04119(.A1(new_n5121_), .A2(new_n5119_), .A3(new_n5120_), .ZN(new_n5122_));
  NOR4_X1    g04120(.A1(new_n5118_), .A2(new_n3483_), .A3(new_n3486_), .A4(new_n5122_), .ZN(new_n5123_));
  OAI21_X1   g04121(.A1(new_n5123_), .A2(new_n5117_), .B(new_n5104_), .ZN(new_n5124_));
  XOR2_X1    g04122(.A1(new_n5096_), .A2(new_n5103_), .Z(new_n5125_));
  NOR2_X1    g04123(.A1(new_n5115_), .A2(new_n5114_), .ZN(new_n5126_));
  NOR2_X1    g04124(.A1(new_n5112_), .A2(new_n5105_), .ZN(new_n5127_));
  OAI22_X1   g04125(.A1(new_n3483_), .A2(new_n3486_), .B1(new_n5126_), .B2(new_n5127_), .ZN(new_n5128_));
  NAND4_X1   g04126(.A1(new_n3444_), .A2(new_n3481_), .A3(new_n5113_), .A4(new_n5116_), .ZN(new_n5129_));
  NAND3_X1   g04127(.A1(new_n5128_), .A2(new_n5129_), .A3(new_n5125_), .ZN(new_n5130_));
  AOI21_X1   g04128(.A1(new_n5124_), .A2(new_n5130_), .B(new_n5095_), .ZN(new_n5131_));
  NOR2_X1    g04129(.A1(new_n5126_), .A2(new_n5127_), .ZN(new_n5132_));
  NAND2_X1   g04130(.A1(new_n3435_), .A2(new_n3428_), .ZN(new_n5133_));
  NAND3_X1   g04131(.A1(new_n5133_), .A2(new_n5110_), .A3(new_n5108_), .ZN(new_n5134_));
  NAND4_X1   g04132(.A1(new_n5132_), .A2(new_n3444_), .A3(new_n3481_), .A4(new_n5134_), .ZN(new_n5135_));
  AOI21_X1   g04133(.A1(new_n5135_), .A2(new_n5128_), .B(new_n5125_), .ZN(new_n5136_));
  NOR3_X1    g04134(.A1(new_n5118_), .A2(new_n3483_), .A3(new_n3486_), .ZN(new_n5137_));
  NOR3_X1    g04135(.A1(new_n5137_), .A2(new_n5117_), .A3(new_n5104_), .ZN(new_n5138_));
  NOR3_X1    g04136(.A1(new_n5136_), .A2(new_n5138_), .A3(new_n3564_), .ZN(new_n5139_));
  OAI21_X1   g04137(.A1(new_n5131_), .A2(new_n5139_), .B(new_n5094_), .ZN(new_n5140_));
  NAND4_X1   g04138(.A1(new_n3549_), .A2(new_n3539_), .A3(new_n3544_), .A4(new_n3551_), .ZN(new_n5141_));
  XOR2_X1    g04139(.A1(new_n5072_), .A2(new_n5141_), .Z(new_n5142_));
  NAND2_X1   g04140(.A1(new_n5091_), .A2(new_n5142_), .ZN(new_n5143_));
  INV_X1     g04141(.I(new_n5079_), .ZN(new_n5144_));
  INV_X1     g04142(.I(new_n5077_), .ZN(new_n5145_));
  NOR2_X1    g04143(.A1(new_n3498_), .A2(new_n3522_), .ZN(new_n5146_));
  NOR3_X1    g04144(.A1(new_n5146_), .A2(new_n5144_), .A3(new_n5145_), .ZN(new_n5147_));
  NOR4_X1    g04145(.A1(new_n5082_), .A2(new_n3570_), .A3(new_n3573_), .A4(new_n5147_), .ZN(new_n5148_));
  NOR2_X1    g04146(.A1(new_n5087_), .A2(new_n3560_), .ZN(new_n5149_));
  NOR4_X1    g04147(.A1(new_n3570_), .A2(new_n3573_), .A3(new_n5084_), .A4(new_n5086_), .ZN(new_n5150_));
  NOR2_X1    g04148(.A1(new_n5149_), .A2(new_n5150_), .ZN(new_n5151_));
  OAI22_X1   g04149(.A1(new_n5151_), .A2(new_n5142_), .B1(new_n5143_), .B2(new_n5148_), .ZN(new_n5152_));
  OAI21_X1   g04150(.A1(new_n5136_), .A2(new_n5138_), .B(new_n3564_), .ZN(new_n5153_));
  NAND3_X1   g04151(.A1(new_n5124_), .A2(new_n5095_), .A3(new_n5130_), .ZN(new_n5154_));
  NAND3_X1   g04152(.A1(new_n5154_), .A2(new_n5153_), .A3(new_n5152_), .ZN(new_n5155_));
  AOI21_X1   g04153(.A1(new_n5140_), .A2(new_n5155_), .B(new_n5065_), .ZN(new_n5156_));
  AOI21_X1   g04154(.A1(new_n5153_), .A2(new_n5154_), .B(new_n5152_), .ZN(new_n5157_));
  NOR3_X1    g04155(.A1(new_n5131_), .A2(new_n5139_), .A3(new_n5094_), .ZN(new_n5158_));
  NOR3_X1    g04156(.A1(new_n3729_), .A2(new_n5158_), .A3(new_n5157_), .ZN(new_n5159_));
  OAI21_X1   g04157(.A1(new_n5159_), .A2(new_n5156_), .B(new_n5064_), .ZN(new_n5160_));
  OR2_X2     g04158(.A1(new_n5001_), .A2(new_n5009_), .Z(new_n5161_));
  NAND3_X1   g04159(.A1(new_n3731_), .A2(new_n5058_), .A3(new_n5059_), .ZN(new_n5162_));
  OAI22_X1   g04160(.A1(new_n5051_), .A2(new_n5040_), .B1(new_n3653_), .B2(new_n3724_), .ZN(new_n5163_));
  NAND3_X1   g04161(.A1(new_n5161_), .A2(new_n5163_), .A3(new_n5162_), .ZN(new_n5164_));
  NAND2_X1   g04162(.A1(new_n5164_), .A2(new_n5062_), .ZN(new_n5165_));
  OAI21_X1   g04163(.A1(new_n5157_), .A2(new_n5158_), .B(new_n3729_), .ZN(new_n5166_));
  NAND3_X1   g04164(.A1(new_n5140_), .A2(new_n5155_), .A3(new_n5065_), .ZN(new_n5167_));
  NAND3_X1   g04165(.A1(new_n5166_), .A2(new_n5167_), .A3(new_n5165_), .ZN(new_n5168_));
  AOI21_X1   g04166(.A1(new_n5160_), .A2(new_n5168_), .B(new_n3735_), .ZN(new_n5169_));
  INV_X1     g04167(.I(new_n3735_), .ZN(new_n5170_));
  AOI21_X1   g04168(.A1(new_n5166_), .A2(new_n5167_), .B(new_n5165_), .ZN(new_n5171_));
  NOR3_X1    g04169(.A1(new_n5064_), .A2(new_n5159_), .A3(new_n5156_), .ZN(new_n5172_));
  NOR3_X1    g04170(.A1(new_n5170_), .A2(new_n5172_), .A3(new_n5171_), .ZN(new_n5173_));
  OAI21_X1   g04171(.A1(new_n5173_), .A2(new_n5169_), .B(new_n4965_), .ZN(new_n5174_));
  INV_X1     g04172(.I(new_n4962_), .ZN(new_n5175_));
  NAND2_X1   g04173(.A1(new_n5175_), .A2(new_n4963_), .ZN(new_n5176_));
  OAI21_X1   g04174(.A1(new_n5172_), .A2(new_n5171_), .B(new_n5170_), .ZN(new_n5177_));
  NAND3_X1   g04175(.A1(new_n5160_), .A2(new_n5168_), .A3(new_n3735_), .ZN(new_n5178_));
  NAND3_X1   g04176(.A1(new_n5177_), .A2(new_n5176_), .A3(new_n5178_), .ZN(new_n5179_));
  AOI21_X1   g04177(.A1(new_n5174_), .A2(new_n5179_), .B(new_n4368_), .ZN(new_n5180_));
  AOI21_X1   g04178(.A1(new_n5177_), .A2(new_n5178_), .B(new_n5176_), .ZN(new_n5181_));
  NOR3_X1    g04179(.A1(new_n4965_), .A2(new_n5173_), .A3(new_n5169_), .ZN(new_n5182_));
  NOR3_X1    g04180(.A1(new_n5181_), .A2(new_n5182_), .A3(new_n4367_), .ZN(new_n5183_));
  OAI21_X1   g04181(.A1(new_n5183_), .A2(new_n5180_), .B(new_n4771_), .ZN(new_n5184_));
  NAND3_X1   g04182(.A1(new_n4768_), .A2(new_n4769_), .A3(new_n4767_), .ZN(new_n5185_));
  OAI21_X1   g04183(.A1(new_n4761_), .A2(new_n4765_), .B(new_n4574_), .ZN(new_n5186_));
  NAND2_X1   g04184(.A1(new_n5186_), .A2(new_n5185_), .ZN(new_n5187_));
  OAI21_X1   g04185(.A1(new_n5181_), .A2(new_n5182_), .B(new_n4367_), .ZN(new_n5188_));
  NAND3_X1   g04186(.A1(new_n5174_), .A2(new_n5179_), .A3(new_n4368_), .ZN(new_n5189_));
  NAND3_X1   g04187(.A1(new_n5187_), .A2(new_n5188_), .A3(new_n5189_), .ZN(new_n5190_));
  AOI21_X1   g04188(.A1(new_n5184_), .A2(new_n5190_), .B(new_n4372_), .ZN(new_n5191_));
  NAND3_X1   g04189(.A1(new_n5184_), .A2(new_n5190_), .A3(new_n4372_), .ZN(new_n5192_));
  OAI21_X1   g04190(.A1(new_n3089_), .A2(new_n5191_), .B(new_n5192_), .ZN(new_n5193_));
  INV_X1     g04191(.I(new_n5193_), .ZN(new_n5194_));
  AOI21_X1   g04192(.A1(new_n2987_), .A2(new_n2988_), .B(new_n2980_), .ZN(new_n5195_));
  NAND2_X1   g04193(.A1(new_n2981_), .A2(new_n2982_), .ZN(new_n5196_));
  NOR2_X1    g04194(.A1(new_n2981_), .A2(new_n2982_), .ZN(new_n5197_));
  AOI21_X1   g04195(.A1(new_n2560_), .A2(new_n5196_), .B(new_n5197_), .ZN(new_n5198_));
  AOI21_X1   g04196(.A1(new_n2591_), .A2(new_n2974_), .B(new_n2977_), .ZN(new_n5199_));
  NOR2_X1    g04197(.A1(new_n5198_), .A2(new_n5199_), .ZN(new_n5200_));
  INV_X1     g04198(.I(new_n5196_), .ZN(new_n5201_));
  INV_X1     g04199(.I(new_n5197_), .ZN(new_n5202_));
  OAI21_X1   g04200(.A1(new_n2606_), .A2(new_n5201_), .B(new_n5202_), .ZN(new_n5203_));
  OAI21_X1   g04201(.A1(new_n2969_), .A2(new_n2973_), .B(new_n2972_), .ZN(new_n5204_));
  NOR2_X1    g04202(.A1(new_n5204_), .A2(new_n5203_), .ZN(new_n5205_));
  NOR2_X1    g04203(.A1(new_n5200_), .A2(new_n5205_), .ZN(new_n5206_));
  OAI21_X1   g04204(.A1(new_n5195_), .A2(new_n2990_), .B(new_n5206_), .ZN(new_n5207_));
  OAI21_X1   g04205(.A1(new_n2998_), .A2(new_n2999_), .B(new_n2995_), .ZN(new_n5208_));
  NAND2_X1   g04206(.A1(new_n5204_), .A2(new_n5203_), .ZN(new_n5209_));
  NAND2_X1   g04207(.A1(new_n5198_), .A2(new_n5199_), .ZN(new_n5210_));
  NAND2_X1   g04208(.A1(new_n5210_), .A2(new_n5209_), .ZN(new_n5211_));
  NAND3_X1   g04209(.A1(new_n5208_), .A2(new_n5211_), .A3(new_n2991_), .ZN(new_n5212_));
  NAND2_X1   g04210(.A1(new_n5207_), .A2(new_n5212_), .ZN(new_n5213_));
  NOR4_X1    g04211(.A1(new_n3019_), .A2(new_n3020_), .A3(new_n2616_), .A4(new_n2626_), .ZN(new_n5214_));
  NOR2_X1    g04212(.A1(new_n3023_), .A2(new_n3021_), .ZN(new_n5215_));
  INV_X1     g04213(.I(new_n5215_), .ZN(new_n5216_));
  OAI21_X1   g04214(.A1(new_n2677_), .A2(new_n5214_), .B(new_n5216_), .ZN(new_n5217_));
  AOI21_X1   g04215(.A1(new_n2680_), .A2(new_n3010_), .B(new_n3015_), .ZN(new_n5218_));
  NOR3_X1    g04216(.A1(new_n3031_), .A2(new_n3039_), .A3(new_n5218_), .ZN(new_n5219_));
  INV_X1     g04217(.I(new_n5218_), .ZN(new_n5220_));
  AOI21_X1   g04218(.A1(new_n3045_), .A2(new_n3032_), .B(new_n5220_), .ZN(new_n5221_));
  NOR3_X1    g04219(.A1(new_n5219_), .A2(new_n5221_), .A3(new_n5217_), .ZN(new_n5222_));
  INV_X1     g04220(.I(new_n5217_), .ZN(new_n5223_));
  NAND3_X1   g04221(.A1(new_n3045_), .A2(new_n3032_), .A3(new_n5220_), .ZN(new_n5224_));
  OAI21_X1   g04222(.A1(new_n3031_), .A2(new_n3039_), .B(new_n5218_), .ZN(new_n5225_));
  AOI21_X1   g04223(.A1(new_n5225_), .A2(new_n5224_), .B(new_n5223_), .ZN(new_n5226_));
  OAI21_X1   g04224(.A1(new_n5222_), .A2(new_n5226_), .B(new_n5213_), .ZN(new_n5227_));
  AOI21_X1   g04225(.A1(new_n5208_), .A2(new_n2991_), .B(new_n5211_), .ZN(new_n5228_));
  NOR3_X1    g04226(.A1(new_n5195_), .A2(new_n5206_), .A3(new_n2990_), .ZN(new_n5229_));
  NOR2_X1    g04227(.A1(new_n5229_), .A2(new_n5228_), .ZN(new_n5230_));
  NAND3_X1   g04228(.A1(new_n5225_), .A2(new_n5224_), .A3(new_n5223_), .ZN(new_n5231_));
  OAI21_X1   g04229(.A1(new_n5219_), .A2(new_n5221_), .B(new_n5217_), .ZN(new_n5232_));
  NAND3_X1   g04230(.A1(new_n5230_), .A2(new_n5232_), .A3(new_n5231_), .ZN(new_n5233_));
  OAI21_X1   g04231(.A1(new_n3002_), .A2(new_n3054_), .B(new_n3049_), .ZN(new_n5234_));
  NAND3_X1   g04232(.A1(new_n5227_), .A2(new_n5233_), .A3(new_n5234_), .ZN(new_n5235_));
  AOI21_X1   g04233(.A1(new_n5232_), .A2(new_n5231_), .B(new_n5230_), .ZN(new_n5236_));
  NOR3_X1    g04234(.A1(new_n5222_), .A2(new_n5226_), .A3(new_n5213_), .ZN(new_n5237_));
  AOI21_X1   g04235(.A1(new_n3053_), .A2(new_n3041_), .B(new_n3055_), .ZN(new_n5238_));
  OAI21_X1   g04236(.A1(new_n5236_), .A2(new_n5237_), .B(new_n5238_), .ZN(new_n5239_));
  OAI21_X1   g04237(.A1(new_n2964_), .A2(new_n2965_), .B(new_n2955_), .ZN(new_n5240_));
  NAND2_X1   g04238(.A1(new_n2940_), .A2(new_n2938_), .ZN(new_n5241_));
  NAND2_X1   g04239(.A1(new_n2454_), .A2(new_n2450_), .ZN(new_n5242_));
  AOI21_X1   g04240(.A1(new_n5241_), .A2(new_n5242_), .B(new_n2946_), .ZN(new_n5243_));
  NAND2_X1   g04241(.A1(new_n2935_), .A2(new_n2933_), .ZN(new_n5244_));
  NOR2_X1    g04242(.A1(new_n2935_), .A2(new_n2933_), .ZN(new_n5245_));
  AOI21_X1   g04243(.A1(new_n2405_), .A2(new_n5244_), .B(new_n5245_), .ZN(new_n5246_));
  AOI21_X1   g04244(.A1(new_n2455_), .A2(new_n2927_), .B(new_n2923_), .ZN(new_n5247_));
  NOR2_X1    g04245(.A1(new_n5246_), .A2(new_n5247_), .ZN(new_n5248_));
  INV_X1     g04246(.I(new_n5244_), .ZN(new_n5249_));
  INV_X1     g04247(.I(new_n5245_), .ZN(new_n5250_));
  OAI21_X1   g04248(.A1(new_n2452_), .A2(new_n5249_), .B(new_n5250_), .ZN(new_n5251_));
  OAI21_X1   g04249(.A1(new_n2437_), .A2(new_n2924_), .B(new_n2922_), .ZN(new_n5252_));
  NOR2_X1    g04250(.A1(new_n5251_), .A2(new_n5252_), .ZN(new_n5253_));
  NOR2_X1    g04251(.A1(new_n5253_), .A2(new_n5248_), .ZN(new_n5254_));
  OAI21_X1   g04252(.A1(new_n5243_), .A2(new_n2942_), .B(new_n5254_), .ZN(new_n5255_));
  NOR2_X1    g04253(.A1(new_n2947_), .A2(new_n2948_), .ZN(new_n5256_));
  NOR2_X1    g04254(.A1(new_n2417_), .A2(new_n2457_), .ZN(new_n5257_));
  OAI21_X1   g04255(.A1(new_n5256_), .A2(new_n5257_), .B(new_n2930_), .ZN(new_n5258_));
  NAND2_X1   g04256(.A1(new_n5251_), .A2(new_n5252_), .ZN(new_n5259_));
  NAND2_X1   g04257(.A1(new_n5246_), .A2(new_n5247_), .ZN(new_n5260_));
  NAND2_X1   g04258(.A1(new_n5259_), .A2(new_n5260_), .ZN(new_n5261_));
  NAND3_X1   g04259(.A1(new_n5258_), .A2(new_n5261_), .A3(new_n2950_), .ZN(new_n5262_));
  NAND2_X1   g04260(.A1(new_n5255_), .A2(new_n5262_), .ZN(new_n5263_));
  NOR4_X1    g04261(.A1(new_n2896_), .A2(new_n2898_), .A3(new_n2465_), .A4(new_n2475_), .ZN(new_n5264_));
  NOR2_X1    g04262(.A1(new_n2897_), .A2(new_n2899_), .ZN(new_n5265_));
  INV_X1     g04263(.I(new_n5265_), .ZN(new_n5266_));
  OAI21_X1   g04264(.A1(new_n2526_), .A2(new_n5264_), .B(new_n5266_), .ZN(new_n5267_));
  AOI21_X1   g04265(.A1(new_n2529_), .A2(new_n2892_), .B(new_n2887_), .ZN(new_n5268_));
  NOR3_X1    g04266(.A1(new_n2961_), .A2(new_n2912_), .A3(new_n5268_), .ZN(new_n5269_));
  INV_X1     g04267(.I(new_n5268_), .ZN(new_n5270_));
  AOI21_X1   g04268(.A1(new_n2908_), .A2(new_n2962_), .B(new_n5270_), .ZN(new_n5271_));
  NOR3_X1    g04269(.A1(new_n5269_), .A2(new_n5271_), .A3(new_n5267_), .ZN(new_n5272_));
  INV_X1     g04270(.I(new_n5267_), .ZN(new_n5273_));
  NAND3_X1   g04271(.A1(new_n2908_), .A2(new_n2962_), .A3(new_n5270_), .ZN(new_n5274_));
  OAI21_X1   g04272(.A1(new_n2961_), .A2(new_n2912_), .B(new_n5268_), .ZN(new_n5275_));
  AOI21_X1   g04273(.A1(new_n5275_), .A2(new_n5274_), .B(new_n5273_), .ZN(new_n5276_));
  OAI21_X1   g04274(.A1(new_n5272_), .A2(new_n5276_), .B(new_n5263_), .ZN(new_n5277_));
  AOI21_X1   g04275(.A1(new_n5258_), .A2(new_n2950_), .B(new_n5261_), .ZN(new_n5278_));
  OAI21_X1   g04276(.A1(new_n2941_), .A2(new_n2946_), .B(new_n2950_), .ZN(new_n5279_));
  NOR2_X1    g04277(.A1(new_n5279_), .A2(new_n5254_), .ZN(new_n5280_));
  NOR2_X1    g04278(.A1(new_n5280_), .A2(new_n5278_), .ZN(new_n5281_));
  NAND3_X1   g04279(.A1(new_n5275_), .A2(new_n5274_), .A3(new_n5273_), .ZN(new_n5282_));
  OAI21_X1   g04280(.A1(new_n5269_), .A2(new_n5271_), .B(new_n5267_), .ZN(new_n5283_));
  NAND3_X1   g04281(.A1(new_n5281_), .A2(new_n5283_), .A3(new_n5282_), .ZN(new_n5284_));
  NAND3_X1   g04282(.A1(new_n5284_), .A2(new_n5277_), .A3(new_n5240_), .ZN(new_n5285_));
  AOI21_X1   g04283(.A1(new_n2916_), .A2(new_n2952_), .B(new_n2966_), .ZN(new_n5286_));
  AOI21_X1   g04284(.A1(new_n5282_), .A2(new_n5283_), .B(new_n5281_), .ZN(new_n5287_));
  NOR3_X1    g04285(.A1(new_n5272_), .A2(new_n5276_), .A3(new_n5263_), .ZN(new_n5288_));
  OAI21_X1   g04286(.A1(new_n5287_), .A2(new_n5288_), .B(new_n5286_), .ZN(new_n5289_));
  NAND4_X1   g04287(.A1(new_n5239_), .A2(new_n5235_), .A3(new_n5289_), .A4(new_n5285_), .ZN(new_n5290_));
  NOR3_X1    g04288(.A1(new_n5236_), .A2(new_n5237_), .A3(new_n5238_), .ZN(new_n5291_));
  AOI21_X1   g04289(.A1(new_n5233_), .A2(new_n5227_), .B(new_n5234_), .ZN(new_n5292_));
  NOR3_X1    g04290(.A1(new_n5287_), .A2(new_n5288_), .A3(new_n5286_), .ZN(new_n5293_));
  AOI21_X1   g04291(.A1(new_n5284_), .A2(new_n5277_), .B(new_n5240_), .ZN(new_n5294_));
  OAI22_X1   g04292(.A1(new_n5291_), .A2(new_n5292_), .B1(new_n5294_), .B2(new_n5293_), .ZN(new_n5295_));
  OAI21_X1   g04293(.A1(new_n2968_), .A2(new_n3064_), .B(new_n3061_), .ZN(new_n5296_));
  NAND3_X1   g04294(.A1(new_n5295_), .A2(new_n5290_), .A3(new_n5296_), .ZN(new_n5297_));
  NOR4_X1    g04295(.A1(new_n5291_), .A2(new_n5292_), .A3(new_n5294_), .A4(new_n5293_), .ZN(new_n5298_));
  AOI22_X1   g04296(.A1(new_n5239_), .A2(new_n5235_), .B1(new_n5289_), .B2(new_n5285_), .ZN(new_n5299_));
  AOI21_X1   g04297(.A1(new_n3063_), .A2(new_n3057_), .B(new_n3065_), .ZN(new_n5300_));
  OAI21_X1   g04298(.A1(new_n5298_), .A2(new_n5299_), .B(new_n5300_), .ZN(new_n5301_));
  OAI21_X1   g04299(.A1(new_n2782_), .A2(new_n2878_), .B(new_n2875_), .ZN(new_n5302_));
  XOR2_X1    g04300(.A1(new_n2244_), .A2(new_n2720_), .Z(new_n5303_));
  AOI21_X1   g04301(.A1(new_n5303_), .A2(new_n2725_), .B(new_n2730_), .ZN(new_n5304_));
  NAND2_X1   g04302(.A1(new_n2713_), .A2(new_n2715_), .ZN(new_n5305_));
  NOR2_X1    g04303(.A1(new_n2713_), .A2(new_n2715_), .ZN(new_n5306_));
  AOI21_X1   g04304(.A1(new_n2292_), .A2(new_n5305_), .B(new_n5306_), .ZN(new_n5307_));
  AOI21_X1   g04305(.A1(new_n2268_), .A2(new_n2708_), .B(new_n2703_), .ZN(new_n5308_));
  NOR2_X1    g04306(.A1(new_n5307_), .A2(new_n5308_), .ZN(new_n5309_));
  INV_X1     g04307(.I(new_n5305_), .ZN(new_n5310_));
  NOR2_X1    g04308(.A1(new_n2244_), .A2(new_n5310_), .ZN(new_n5311_));
  AOI21_X1   g04309(.A1(new_n2295_), .A2(new_n2296_), .B(new_n2704_), .ZN(new_n5312_));
  NOR4_X1    g04310(.A1(new_n5311_), .A2(new_n5312_), .A3(new_n2703_), .A4(new_n5306_), .ZN(new_n5313_));
  NOR2_X1    g04311(.A1(new_n5313_), .A2(new_n5309_), .ZN(new_n5314_));
  OAI21_X1   g04312(.A1(new_n5304_), .A2(new_n2726_), .B(new_n5314_), .ZN(new_n5315_));
  OAI21_X1   g04313(.A1(new_n2722_), .A2(new_n2723_), .B(new_n2711_), .ZN(new_n5316_));
  OAI22_X1   g04314(.A1(new_n5311_), .A2(new_n5306_), .B1(new_n5312_), .B2(new_n2703_), .ZN(new_n5317_));
  NAND2_X1   g04315(.A1(new_n5307_), .A2(new_n5308_), .ZN(new_n5318_));
  NAND2_X1   g04316(.A1(new_n5317_), .A2(new_n5318_), .ZN(new_n5319_));
  NAND3_X1   g04317(.A1(new_n5316_), .A2(new_n5319_), .A3(new_n2732_), .ZN(new_n5320_));
  NAND2_X1   g04318(.A1(new_n5315_), .A2(new_n5320_), .ZN(new_n5321_));
  NOR4_X1    g04319(.A1(new_n2749_), .A2(new_n2751_), .A3(new_n2306_), .A4(new_n2316_), .ZN(new_n5322_));
  NOR2_X1    g04320(.A1(new_n2750_), .A2(new_n2752_), .ZN(new_n5323_));
  INV_X1     g04321(.I(new_n5323_), .ZN(new_n5324_));
  OAI21_X1   g04322(.A1(new_n2320_), .A2(new_n5322_), .B(new_n5324_), .ZN(new_n5325_));
  NAND2_X1   g04323(.A1(new_n2367_), .A2(new_n2757_), .ZN(new_n5326_));
  NAND2_X1   g04324(.A1(new_n2753_), .A2(new_n2320_), .ZN(new_n5327_));
  NAND2_X1   g04325(.A1(new_n5327_), .A2(new_n5326_), .ZN(new_n5328_));
  NAND2_X1   g04326(.A1(new_n2332_), .A2(new_n2372_), .ZN(new_n5329_));
  AOI21_X1   g04327(.A1(new_n5329_), .A2(new_n5328_), .B(new_n2771_), .ZN(new_n5330_));
  AOI21_X1   g04328(.A1(new_n2353_), .A2(new_n2745_), .B(new_n2740_), .ZN(new_n5331_));
  NOR3_X1    g04329(.A1(new_n5330_), .A2(new_n2762_), .A3(new_n5331_), .ZN(new_n5332_));
  INV_X1     g04330(.I(new_n5331_), .ZN(new_n5333_));
  AOI21_X1   g04331(.A1(new_n2761_), .A2(new_n2765_), .B(new_n5333_), .ZN(new_n5334_));
  NOR3_X1    g04332(.A1(new_n5332_), .A2(new_n5334_), .A3(new_n5325_), .ZN(new_n5335_));
  INV_X1     g04333(.I(new_n5325_), .ZN(new_n5336_));
  NAND3_X1   g04334(.A1(new_n2761_), .A2(new_n2765_), .A3(new_n5333_), .ZN(new_n5337_));
  OAI21_X1   g04335(.A1(new_n5330_), .A2(new_n2762_), .B(new_n5331_), .ZN(new_n5338_));
  AOI21_X1   g04336(.A1(new_n5338_), .A2(new_n5337_), .B(new_n5336_), .ZN(new_n5339_));
  OAI21_X1   g04337(.A1(new_n5335_), .A2(new_n5339_), .B(new_n5321_), .ZN(new_n5340_));
  AOI21_X1   g04338(.A1(new_n5316_), .A2(new_n2732_), .B(new_n5319_), .ZN(new_n5341_));
  NOR3_X1    g04339(.A1(new_n5304_), .A2(new_n5314_), .A3(new_n2726_), .ZN(new_n5342_));
  NOR2_X1    g04340(.A1(new_n5342_), .A2(new_n5341_), .ZN(new_n5343_));
  NAND3_X1   g04341(.A1(new_n5338_), .A2(new_n5337_), .A3(new_n5336_), .ZN(new_n5344_));
  OAI21_X1   g04342(.A1(new_n5332_), .A2(new_n5334_), .B(new_n5325_), .ZN(new_n5345_));
  NAND3_X1   g04343(.A1(new_n5343_), .A2(new_n5345_), .A3(new_n5344_), .ZN(new_n5346_));
  OAI21_X1   g04344(.A1(new_n2778_), .A2(new_n2767_), .B(new_n2780_), .ZN(new_n5347_));
  NAND3_X1   g04345(.A1(new_n5346_), .A2(new_n5340_), .A3(new_n5347_), .ZN(new_n5348_));
  AOI21_X1   g04346(.A1(new_n5344_), .A2(new_n5345_), .B(new_n5343_), .ZN(new_n5349_));
  NOR3_X1    g04347(.A1(new_n5335_), .A2(new_n5339_), .A3(new_n5321_), .ZN(new_n5350_));
  AOI21_X1   g04348(.A1(new_n2734_), .A2(new_n2779_), .B(new_n2774_), .ZN(new_n5351_));
  OAI21_X1   g04349(.A1(new_n5349_), .A2(new_n5350_), .B(new_n5351_), .ZN(new_n5352_));
  OAI21_X1   g04350(.A1(new_n2868_), .A2(new_n2869_), .B(new_n2859_), .ZN(new_n5353_));
  NAND2_X1   g04351(.A1(new_n2843_), .A2(new_n2841_), .ZN(new_n5354_));
  NAND3_X1   g04352(.A1(new_n2141_), .A2(new_n2137_), .A3(new_n2090_), .ZN(new_n5355_));
  AOI21_X1   g04353(.A1(new_n5354_), .A2(new_n5355_), .B(new_n2849_), .ZN(new_n5356_));
  NAND2_X1   g04354(.A1(new_n2838_), .A2(new_n2836_), .ZN(new_n5357_));
  NOR2_X1    g04355(.A1(new_n2838_), .A2(new_n2836_), .ZN(new_n5358_));
  AOI21_X1   g04356(.A1(new_n2137_), .A2(new_n5357_), .B(new_n5358_), .ZN(new_n5359_));
  AOI21_X1   g04357(.A1(new_n2112_), .A2(new_n2830_), .B(new_n2825_), .ZN(new_n5360_));
  NOR2_X1    g04358(.A1(new_n5359_), .A2(new_n5360_), .ZN(new_n5361_));
  INV_X1     g04359(.I(new_n5357_), .ZN(new_n5362_));
  NOR2_X1    g04360(.A1(new_n2089_), .A2(new_n5362_), .ZN(new_n5363_));
  NOR2_X1    g04361(.A1(new_n2117_), .A2(new_n2115_), .ZN(new_n5364_));
  NOR2_X1    g04362(.A1(new_n2120_), .A2(new_n2123_), .ZN(new_n5365_));
  AOI21_X1   g04363(.A1(new_n5364_), .A2(new_n5365_), .B(new_n2826_), .ZN(new_n5366_));
  NOR4_X1    g04364(.A1(new_n5363_), .A2(new_n5366_), .A3(new_n2825_), .A4(new_n5358_), .ZN(new_n5367_));
  NOR2_X1    g04365(.A1(new_n5367_), .A2(new_n5361_), .ZN(new_n5368_));
  OAI21_X1   g04366(.A1(new_n5356_), .A2(new_n2845_), .B(new_n5368_), .ZN(new_n5369_));
  NOR2_X1    g04367(.A1(new_n2850_), .A2(new_n2851_), .ZN(new_n5370_));
  NOR2_X1    g04368(.A1(new_n2138_), .A2(new_n2125_), .ZN(new_n5371_));
  OAI21_X1   g04369(.A1(new_n5370_), .A2(new_n5371_), .B(new_n2833_), .ZN(new_n5372_));
  OAI22_X1   g04370(.A1(new_n5363_), .A2(new_n5358_), .B1(new_n5366_), .B2(new_n2825_), .ZN(new_n5373_));
  NAND2_X1   g04371(.A1(new_n5359_), .A2(new_n5360_), .ZN(new_n5374_));
  NAND2_X1   g04372(.A1(new_n5373_), .A2(new_n5374_), .ZN(new_n5375_));
  NAND3_X1   g04373(.A1(new_n5372_), .A2(new_n5375_), .A3(new_n2853_), .ZN(new_n5376_));
  NAND2_X1   g04374(.A1(new_n5369_), .A2(new_n5376_), .ZN(new_n5377_));
  NOR4_X1    g04375(.A1(new_n2800_), .A2(new_n2801_), .A3(new_n2149_), .A4(new_n2159_), .ZN(new_n5378_));
  NOR2_X1    g04376(.A1(new_n2804_), .A2(new_n2802_), .ZN(new_n5379_));
  INV_X1     g04377(.I(new_n5379_), .ZN(new_n5380_));
  OAI21_X1   g04378(.A1(new_n2163_), .A2(new_n5378_), .B(new_n5380_), .ZN(new_n5381_));
  AOI21_X1   g04379(.A1(new_n2196_), .A2(new_n2796_), .B(new_n2787_), .ZN(new_n5382_));
  NOR3_X1    g04380(.A1(new_n2864_), .A2(new_n2817_), .A3(new_n5382_), .ZN(new_n5383_));
  INV_X1     g04381(.I(new_n5382_), .ZN(new_n5384_));
  AOI21_X1   g04382(.A1(new_n2811_), .A2(new_n2865_), .B(new_n5384_), .ZN(new_n5385_));
  NOR3_X1    g04383(.A1(new_n5383_), .A2(new_n5385_), .A3(new_n5381_), .ZN(new_n5386_));
  INV_X1     g04384(.I(new_n5381_), .ZN(new_n5387_));
  NAND3_X1   g04385(.A1(new_n2811_), .A2(new_n2865_), .A3(new_n5384_), .ZN(new_n5388_));
  OAI21_X1   g04386(.A1(new_n2864_), .A2(new_n2817_), .B(new_n5382_), .ZN(new_n5389_));
  AOI21_X1   g04387(.A1(new_n5389_), .A2(new_n5388_), .B(new_n5387_), .ZN(new_n5390_));
  OAI21_X1   g04388(.A1(new_n5386_), .A2(new_n5390_), .B(new_n5377_), .ZN(new_n5391_));
  AOI21_X1   g04389(.A1(new_n2852_), .A2(new_n2833_), .B(new_n2845_), .ZN(new_n5392_));
  NOR2_X1    g04390(.A1(new_n5392_), .A2(new_n5375_), .ZN(new_n5393_));
  NOR3_X1    g04391(.A1(new_n5356_), .A2(new_n5368_), .A3(new_n2845_), .ZN(new_n5394_));
  NOR2_X1    g04392(.A1(new_n5393_), .A2(new_n5394_), .ZN(new_n5395_));
  NAND3_X1   g04393(.A1(new_n5389_), .A2(new_n5388_), .A3(new_n5387_), .ZN(new_n5396_));
  OAI21_X1   g04394(.A1(new_n5383_), .A2(new_n5385_), .B(new_n5381_), .ZN(new_n5397_));
  NAND3_X1   g04395(.A1(new_n5395_), .A2(new_n5397_), .A3(new_n5396_), .ZN(new_n5398_));
  NAND3_X1   g04396(.A1(new_n5398_), .A2(new_n5391_), .A3(new_n5353_), .ZN(new_n5399_));
  AOI21_X1   g04397(.A1(new_n2820_), .A2(new_n2855_), .B(new_n2870_), .ZN(new_n5400_));
  AOI21_X1   g04398(.A1(new_n5396_), .A2(new_n5397_), .B(new_n5395_), .ZN(new_n5401_));
  NOR3_X1    g04399(.A1(new_n5386_), .A2(new_n5390_), .A3(new_n5377_), .ZN(new_n5402_));
  OAI21_X1   g04400(.A1(new_n5401_), .A2(new_n5402_), .B(new_n5400_), .ZN(new_n5403_));
  NAND4_X1   g04401(.A1(new_n5348_), .A2(new_n5352_), .A3(new_n5403_), .A4(new_n5399_), .ZN(new_n5404_));
  NOR3_X1    g04402(.A1(new_n5349_), .A2(new_n5350_), .A3(new_n5351_), .ZN(new_n5405_));
  AOI21_X1   g04403(.A1(new_n5346_), .A2(new_n5340_), .B(new_n5347_), .ZN(new_n5406_));
  NOR3_X1    g04404(.A1(new_n5401_), .A2(new_n5402_), .A3(new_n5400_), .ZN(new_n5407_));
  AOI21_X1   g04405(.A1(new_n5398_), .A2(new_n5391_), .B(new_n5353_), .ZN(new_n5408_));
  OAI22_X1   g04406(.A1(new_n5405_), .A2(new_n5406_), .B1(new_n5408_), .B2(new_n5407_), .ZN(new_n5409_));
  NAND3_X1   g04407(.A1(new_n5409_), .A2(new_n5404_), .A3(new_n5302_), .ZN(new_n5410_));
  INV_X1     g04408(.I(new_n2782_), .ZN(new_n5411_));
  NOR3_X1    g04409(.A1(new_n2382_), .A2(new_n2860_), .A3(new_n2871_), .ZN(new_n5412_));
  AOI21_X1   g04410(.A1(new_n5411_), .A2(new_n2872_), .B(new_n5412_), .ZN(new_n5413_));
  NOR4_X1    g04411(.A1(new_n5405_), .A2(new_n5406_), .A3(new_n5408_), .A4(new_n5407_), .ZN(new_n5414_));
  AOI22_X1   g04412(.A1(new_n5352_), .A2(new_n5348_), .B1(new_n5403_), .B2(new_n5399_), .ZN(new_n5415_));
  OAI21_X1   g04413(.A1(new_n5414_), .A2(new_n5415_), .B(new_n5413_), .ZN(new_n5416_));
  NAND4_X1   g04414(.A1(new_n5297_), .A2(new_n5301_), .A3(new_n5416_), .A4(new_n5410_), .ZN(new_n5417_));
  NOR3_X1    g04415(.A1(new_n5298_), .A2(new_n5299_), .A3(new_n5300_), .ZN(new_n5418_));
  AOI21_X1   g04416(.A1(new_n5295_), .A2(new_n5290_), .B(new_n5296_), .ZN(new_n5419_));
  NOR3_X1    g04417(.A1(new_n5414_), .A2(new_n5415_), .A3(new_n5413_), .ZN(new_n5420_));
  AOI21_X1   g04418(.A1(new_n5409_), .A2(new_n5404_), .B(new_n5302_), .ZN(new_n5421_));
  OAI22_X1   g04419(.A1(new_n5418_), .A2(new_n5419_), .B1(new_n5420_), .B2(new_n5421_), .ZN(new_n5422_));
  OAI21_X1   g04420(.A1(new_n2881_), .A2(new_n3073_), .B(new_n3070_), .ZN(new_n5423_));
  NAND3_X1   g04421(.A1(new_n5422_), .A2(new_n5417_), .A3(new_n5423_), .ZN(new_n5424_));
  NOR4_X1    g04422(.A1(new_n5418_), .A2(new_n5419_), .A3(new_n5420_), .A4(new_n5421_), .ZN(new_n5425_));
  AOI22_X1   g04423(.A1(new_n5297_), .A2(new_n5301_), .B1(new_n5416_), .B2(new_n5410_), .ZN(new_n5426_));
  AOI21_X1   g04424(.A1(new_n3072_), .A2(new_n3067_), .B(new_n3074_), .ZN(new_n5427_));
  OAI21_X1   g04425(.A1(new_n5425_), .A2(new_n5426_), .B(new_n5427_), .ZN(new_n5428_));
  OAI21_X1   g04426(.A1(new_n2061_), .A2(new_n2062_), .B(new_n2059_), .ZN(new_n5429_));
  NAND2_X1   g04427(.A1(new_n1443_), .A2(new_n1442_), .ZN(new_n5430_));
  NAND3_X1   g04428(.A1(new_n1275_), .A2(new_n1295_), .A3(new_n1298_), .ZN(new_n5431_));
  AOI21_X1   g04429(.A1(new_n5431_), .A2(new_n5430_), .B(new_n1440_), .ZN(new_n5432_));
  NOR4_X1    g04430(.A1(new_n1423_), .A2(new_n1425_), .A3(new_n1249_), .A4(new_n1259_), .ZN(new_n5433_));
  INV_X1     g04431(.I(new_n5433_), .ZN(new_n5434_));
  NAND2_X1   g04432(.A1(new_n1301_), .A2(new_n5434_), .ZN(new_n5435_));
  NOR2_X1    g04433(.A1(new_n1424_), .A2(new_n1426_), .ZN(new_n5436_));
  INV_X1     g04434(.I(new_n5436_), .ZN(new_n5437_));
  OAI21_X1   g04435(.A1(new_n1296_), .A2(new_n1297_), .B(new_n1419_), .ZN(new_n5438_));
  AOI22_X1   g04436(.A1(new_n5435_), .A2(new_n5437_), .B1(new_n5438_), .B2(new_n1418_), .ZN(new_n5439_));
  NOR2_X1    g04437(.A1(new_n1252_), .A2(new_n1248_), .ZN(new_n5440_));
  NOR2_X1    g04438(.A1(new_n1262_), .A2(new_n1258_), .ZN(new_n5441_));
  AOI21_X1   g04439(.A1(new_n5440_), .A2(new_n5441_), .B(new_n5433_), .ZN(new_n5442_));
  AOI21_X1   g04440(.A1(new_n1316_), .A2(new_n1317_), .B(new_n1415_), .ZN(new_n5443_));
  NOR4_X1    g04441(.A1(new_n5442_), .A2(new_n5443_), .A3(new_n1414_), .A4(new_n5436_), .ZN(new_n5444_));
  NOR2_X1    g04442(.A1(new_n5439_), .A2(new_n5444_), .ZN(new_n5445_));
  OAI21_X1   g04443(.A1(new_n5432_), .A2(new_n1436_), .B(new_n5445_), .ZN(new_n5446_));
  OAI21_X1   g04444(.A1(new_n1433_), .A2(new_n1434_), .B(new_n1422_), .ZN(new_n5447_));
  OAI22_X1   g04445(.A1(new_n5442_), .A2(new_n5436_), .B1(new_n5443_), .B2(new_n1414_), .ZN(new_n5448_));
  NAND4_X1   g04446(.A1(new_n5435_), .A2(new_n5438_), .A3(new_n1418_), .A4(new_n5437_), .ZN(new_n5449_));
  NAND2_X1   g04447(.A1(new_n5448_), .A2(new_n5449_), .ZN(new_n5450_));
  NAND3_X1   g04448(.A1(new_n5447_), .A2(new_n5450_), .A3(new_n1444_), .ZN(new_n5451_));
  NAND2_X1   g04449(.A1(new_n5446_), .A2(new_n5451_), .ZN(new_n5452_));
  NOR4_X1    g04450(.A1(new_n1465_), .A2(new_n1466_), .A3(new_n1327_), .A4(new_n1337_), .ZN(new_n5453_));
  NOR2_X1    g04451(.A1(new_n1469_), .A2(new_n1467_), .ZN(new_n5454_));
  INV_X1     g04452(.I(new_n5454_), .ZN(new_n5455_));
  OAI21_X1   g04453(.A1(new_n1341_), .A2(new_n5453_), .B(new_n5455_), .ZN(new_n5456_));
  NAND2_X1   g04454(.A1(new_n1483_), .A2(new_n1481_), .ZN(new_n5457_));
  AOI21_X1   g04455(.A1(new_n5457_), .A2(new_n1477_), .B(new_n1490_), .ZN(new_n5458_));
  AOI21_X1   g04456(.A1(new_n1374_), .A2(new_n1461_), .B(new_n1452_), .ZN(new_n5459_));
  NOR3_X1    g04457(.A1(new_n5458_), .A2(new_n1478_), .A3(new_n5459_), .ZN(new_n5460_));
  INV_X1     g04458(.I(new_n5459_), .ZN(new_n5461_));
  AOI21_X1   g04459(.A1(new_n1476_), .A2(new_n1484_), .B(new_n5461_), .ZN(new_n5462_));
  NOR3_X1    g04460(.A1(new_n5460_), .A2(new_n5462_), .A3(new_n5456_), .ZN(new_n5463_));
  INV_X1     g04461(.I(new_n5456_), .ZN(new_n5464_));
  NAND3_X1   g04462(.A1(new_n1476_), .A2(new_n1484_), .A3(new_n5461_), .ZN(new_n5465_));
  OAI21_X1   g04463(.A1(new_n5458_), .A2(new_n1478_), .B(new_n5459_), .ZN(new_n5466_));
  AOI21_X1   g04464(.A1(new_n5466_), .A2(new_n5465_), .B(new_n5464_), .ZN(new_n5467_));
  OAI21_X1   g04465(.A1(new_n5463_), .A2(new_n5467_), .B(new_n5452_), .ZN(new_n5468_));
  AOI21_X1   g04466(.A1(new_n5447_), .A2(new_n1444_), .B(new_n5450_), .ZN(new_n5469_));
  NOR3_X1    g04467(.A1(new_n5432_), .A2(new_n5445_), .A3(new_n1436_), .ZN(new_n5470_));
  NOR2_X1    g04468(.A1(new_n5469_), .A2(new_n5470_), .ZN(new_n5471_));
  NAND3_X1   g04469(.A1(new_n5466_), .A2(new_n5465_), .A3(new_n5464_), .ZN(new_n5472_));
  OAI21_X1   g04470(.A1(new_n5460_), .A2(new_n5462_), .B(new_n5456_), .ZN(new_n5473_));
  NAND3_X1   g04471(.A1(new_n5471_), .A2(new_n5473_), .A3(new_n5472_), .ZN(new_n5474_));
  OAI21_X1   g04472(.A1(new_n1497_), .A2(new_n1486_), .B(new_n1499_), .ZN(new_n5475_));
  NAND3_X1   g04473(.A1(new_n5474_), .A2(new_n5468_), .A3(new_n5475_), .ZN(new_n5476_));
  AOI21_X1   g04474(.A1(new_n5472_), .A2(new_n5473_), .B(new_n5471_), .ZN(new_n5477_));
  NOR3_X1    g04475(.A1(new_n5463_), .A2(new_n5467_), .A3(new_n5452_), .ZN(new_n5478_));
  AOI21_X1   g04476(.A1(new_n1446_), .A2(new_n1498_), .B(new_n1493_), .ZN(new_n5479_));
  OAI21_X1   g04477(.A1(new_n5477_), .A2(new_n5478_), .B(new_n5479_), .ZN(new_n5480_));
  OAI21_X1   g04478(.A1(new_n1239_), .A2(new_n1238_), .B(new_n1228_), .ZN(new_n5481_));
  OAI21_X1   g04479(.A1(new_n1204_), .A2(new_n1134_), .B(new_n1198_), .ZN(new_n5482_));
  NOR2_X1    g04480(.A1(new_n1153_), .A2(new_n1215_), .ZN(new_n5483_));
  AOI21_X1   g04481(.A1(new_n1153_), .A2(new_n1215_), .B(new_n1214_), .ZN(new_n5484_));
  INV_X1     g04482(.I(new_n1130_), .ZN(new_n5485_));
  AOI21_X1   g04483(.A1(new_n1187_), .A2(new_n1132_), .B(new_n5485_), .ZN(new_n5486_));
  OAI21_X1   g04484(.A1(new_n5483_), .A2(new_n5484_), .B(new_n5486_), .ZN(new_n5487_));
  NAND2_X1   g04485(.A1(new_n1174_), .A2(new_n1156_), .ZN(new_n5488_));
  OAI21_X1   g04486(.A1(new_n1174_), .A2(new_n1156_), .B(new_n1158_), .ZN(new_n5489_));
  OAI21_X1   g04487(.A1(new_n1126_), .A2(new_n1131_), .B(new_n1130_), .ZN(new_n5490_));
  NAND3_X1   g04488(.A1(new_n5489_), .A2(new_n5490_), .A3(new_n5488_), .ZN(new_n5491_));
  NAND2_X1   g04489(.A1(new_n5487_), .A2(new_n5491_), .ZN(new_n5492_));
  NAND2_X1   g04490(.A1(new_n5482_), .A2(new_n5492_), .ZN(new_n5493_));
  AOI21_X1   g04491(.A1(new_n1192_), .A2(new_n1200_), .B(new_n1218_), .ZN(new_n5494_));
  AOI21_X1   g04492(.A1(new_n5488_), .A2(new_n5489_), .B(new_n5490_), .ZN(new_n5495_));
  NOR3_X1    g04493(.A1(new_n5486_), .A2(new_n5484_), .A3(new_n5483_), .ZN(new_n5496_));
  NOR2_X1    g04494(.A1(new_n5495_), .A2(new_n5496_), .ZN(new_n5497_));
  NAND2_X1   g04495(.A1(new_n5494_), .A2(new_n5497_), .ZN(new_n5498_));
  OAI21_X1   g04496(.A1(new_n1103_), .A2(new_n1099_), .B(new_n1097_), .ZN(new_n5499_));
  NOR2_X1    g04497(.A1(new_n1068_), .A2(new_n1231_), .ZN(new_n5500_));
  AOI21_X1   g04498(.A1(new_n1068_), .A2(new_n1231_), .B(new_n1230_), .ZN(new_n5501_));
  AOI21_X1   g04499(.A1(new_n1023_), .A2(new_n1044_), .B(new_n1028_), .ZN(new_n5502_));
  OAI21_X1   g04500(.A1(new_n5500_), .A2(new_n5501_), .B(new_n5502_), .ZN(new_n5503_));
  NAND2_X1   g04501(.A1(new_n1084_), .A2(new_n1071_), .ZN(new_n5504_));
  OAI21_X1   g04502(.A1(new_n1084_), .A2(new_n1071_), .B(new_n1069_), .ZN(new_n5505_));
  OAI21_X1   g04503(.A1(new_n1042_), .A2(new_n1029_), .B(new_n1043_), .ZN(new_n5506_));
  NAND3_X1   g04504(.A1(new_n5505_), .A2(new_n5506_), .A3(new_n5504_), .ZN(new_n5507_));
  NAND2_X1   g04505(.A1(new_n5503_), .A2(new_n5507_), .ZN(new_n5508_));
  NAND2_X1   g04506(.A1(new_n5499_), .A2(new_n5508_), .ZN(new_n5509_));
  AOI21_X1   g04507(.A1(new_n1091_), .A2(new_n1047_), .B(new_n1234_), .ZN(new_n5510_));
  AOI21_X1   g04508(.A1(new_n5504_), .A2(new_n5505_), .B(new_n5506_), .ZN(new_n5511_));
  NOR3_X1    g04509(.A1(new_n5502_), .A2(new_n5501_), .A3(new_n5500_), .ZN(new_n5512_));
  NOR2_X1    g04510(.A1(new_n5511_), .A2(new_n5512_), .ZN(new_n5513_));
  NAND2_X1   g04511(.A1(new_n5510_), .A2(new_n5513_), .ZN(new_n5514_));
  NAND4_X1   g04512(.A1(new_n5509_), .A2(new_n5493_), .A3(new_n5514_), .A4(new_n5498_), .ZN(new_n5515_));
  NOR2_X1    g04513(.A1(new_n5494_), .A2(new_n5497_), .ZN(new_n5516_));
  NOR2_X1    g04514(.A1(new_n5482_), .A2(new_n5492_), .ZN(new_n5517_));
  NOR2_X1    g04515(.A1(new_n5510_), .A2(new_n5513_), .ZN(new_n5518_));
  NOR2_X1    g04516(.A1(new_n5499_), .A2(new_n5508_), .ZN(new_n5519_));
  OAI22_X1   g04517(.A1(new_n5519_), .A2(new_n5518_), .B1(new_n5517_), .B2(new_n5516_), .ZN(new_n5520_));
  NAND3_X1   g04518(.A1(new_n5520_), .A2(new_n5481_), .A3(new_n5515_), .ZN(new_n5521_));
  AOI21_X1   g04519(.A1(new_n1213_), .A2(new_n1106_), .B(new_n1240_), .ZN(new_n5522_));
  NOR4_X1    g04520(.A1(new_n5519_), .A2(new_n5517_), .A3(new_n5518_), .A4(new_n5516_), .ZN(new_n5523_));
  AOI22_X1   g04521(.A1(new_n5509_), .A2(new_n5514_), .B1(new_n5493_), .B2(new_n5498_), .ZN(new_n5524_));
  OAI21_X1   g04522(.A1(new_n5523_), .A2(new_n5524_), .B(new_n5522_), .ZN(new_n5525_));
  NAND4_X1   g04523(.A1(new_n5480_), .A2(new_n5476_), .A3(new_n5525_), .A4(new_n5521_), .ZN(new_n5526_));
  NOR3_X1    g04524(.A1(new_n5477_), .A2(new_n5478_), .A3(new_n5479_), .ZN(new_n5527_));
  AOI21_X1   g04525(.A1(new_n5474_), .A2(new_n5468_), .B(new_n5475_), .ZN(new_n5528_));
  NOR3_X1    g04526(.A1(new_n5522_), .A2(new_n5523_), .A3(new_n5524_), .ZN(new_n5529_));
  AOI21_X1   g04527(.A1(new_n5515_), .A2(new_n5520_), .B(new_n5481_), .ZN(new_n5530_));
  OAI22_X1   g04528(.A1(new_n5528_), .A2(new_n5527_), .B1(new_n5529_), .B2(new_n5530_), .ZN(new_n5531_));
  OAI21_X1   g04529(.A1(new_n1242_), .A2(new_n1513_), .B(new_n1501_), .ZN(new_n5532_));
  NAND3_X1   g04530(.A1(new_n5531_), .A2(new_n5526_), .A3(new_n5532_), .ZN(new_n5533_));
  NOR4_X1    g04531(.A1(new_n5528_), .A2(new_n5527_), .A3(new_n5529_), .A4(new_n5530_), .ZN(new_n5534_));
  AOI22_X1   g04532(.A1(new_n5480_), .A2(new_n5476_), .B1(new_n5525_), .B2(new_n5521_), .ZN(new_n5535_));
  AOI21_X1   g04533(.A1(new_n1511_), .A2(new_n1509_), .B(new_n1512_), .ZN(new_n5536_));
  OAI21_X1   g04534(.A1(new_n5535_), .A2(new_n5534_), .B(new_n5536_), .ZN(new_n5537_));
  OAI21_X1   g04535(.A1(new_n2050_), .A2(new_n2051_), .B(new_n2048_), .ZN(new_n5538_));
  AOI22_X1   g04536(.A1(new_n1876_), .A2(new_n1832_), .B1(new_n1850_), .B2(new_n1854_), .ZN(new_n5539_));
  NOR2_X1    g04537(.A1(new_n1863_), .A2(new_n1861_), .ZN(new_n5540_));
  AOI21_X1   g04538(.A1(new_n1830_), .A2(new_n1880_), .B(new_n5540_), .ZN(new_n5541_));
  AOI21_X1   g04539(.A1(new_n1828_), .A2(new_n1852_), .B(new_n1847_), .ZN(new_n5542_));
  NOR2_X1    g04540(.A1(new_n5541_), .A2(new_n5542_), .ZN(new_n5543_));
  INV_X1     g04541(.I(new_n5540_), .ZN(new_n5544_));
  OAI21_X1   g04542(.A1(new_n1815_), .A2(new_n1881_), .B(new_n5544_), .ZN(new_n5545_));
  OAI21_X1   g04543(.A1(new_n1783_), .A2(new_n1848_), .B(new_n1851_), .ZN(new_n5546_));
  NOR2_X1    g04544(.A1(new_n5545_), .A2(new_n5546_), .ZN(new_n5547_));
  NOR2_X1    g04545(.A1(new_n5547_), .A2(new_n5543_), .ZN(new_n5548_));
  OAI21_X1   g04546(.A1(new_n1884_), .A2(new_n5539_), .B(new_n5548_), .ZN(new_n5549_));
  OAI21_X1   g04547(.A1(new_n1856_), .A2(new_n1868_), .B(new_n1855_), .ZN(new_n5550_));
  NAND2_X1   g04548(.A1(new_n5545_), .A2(new_n5546_), .ZN(new_n5551_));
  NAND2_X1   g04549(.A1(new_n5541_), .A2(new_n5542_), .ZN(new_n5552_));
  NAND2_X1   g04550(.A1(new_n5551_), .A2(new_n5552_), .ZN(new_n5553_));
  NAND3_X1   g04551(.A1(new_n5550_), .A2(new_n5553_), .A3(new_n1943_), .ZN(new_n5554_));
  NAND2_X1   g04552(.A1(new_n5549_), .A2(new_n5554_), .ZN(new_n5555_));
  NAND2_X1   g04553(.A1(new_n1925_), .A2(new_n1924_), .ZN(new_n5556_));
  NAND2_X1   g04554(.A1(new_n1757_), .A2(new_n1753_), .ZN(new_n5557_));
  AOI21_X1   g04555(.A1(new_n5557_), .A2(new_n5556_), .B(new_n1923_), .ZN(new_n5558_));
  AOI21_X1   g04556(.A1(new_n1758_), .A2(new_n1898_), .B(new_n1891_), .ZN(new_n5559_));
  NOR3_X1    g04557(.A1(new_n5558_), .A2(new_n1933_), .A3(new_n5559_), .ZN(new_n5560_));
  NOR2_X1    g04558(.A1(new_n1907_), .A2(new_n1911_), .ZN(new_n5561_));
  OAI21_X1   g04559(.A1(new_n5561_), .A2(new_n1935_), .B(new_n1901_), .ZN(new_n5562_));
  INV_X1     g04560(.I(new_n5559_), .ZN(new_n5563_));
  AOI21_X1   g04561(.A1(new_n5562_), .A2(new_n1919_), .B(new_n5563_), .ZN(new_n5564_));
  NOR3_X1    g04562(.A1(new_n5560_), .A2(new_n5564_), .A3(new_n1918_), .ZN(new_n5565_));
  NAND3_X1   g04563(.A1(new_n5562_), .A2(new_n1919_), .A3(new_n5563_), .ZN(new_n5566_));
  OAI21_X1   g04564(.A1(new_n5558_), .A2(new_n1933_), .B(new_n5559_), .ZN(new_n5567_));
  AOI21_X1   g04565(.A1(new_n5567_), .A2(new_n5566_), .B(new_n1932_), .ZN(new_n5568_));
  OAI21_X1   g04566(.A1(new_n5565_), .A2(new_n5568_), .B(new_n5555_), .ZN(new_n5569_));
  AOI21_X1   g04567(.A1(new_n5550_), .A2(new_n1943_), .B(new_n5553_), .ZN(new_n5570_));
  NOR3_X1    g04568(.A1(new_n5539_), .A2(new_n5548_), .A3(new_n1884_), .ZN(new_n5571_));
  NOR2_X1    g04569(.A1(new_n5570_), .A2(new_n5571_), .ZN(new_n5572_));
  NAND3_X1   g04570(.A1(new_n5567_), .A2(new_n5566_), .A3(new_n1932_), .ZN(new_n5573_));
  OAI21_X1   g04571(.A1(new_n5560_), .A2(new_n5564_), .B(new_n1918_), .ZN(new_n5574_));
  NAND3_X1   g04572(.A1(new_n5572_), .A2(new_n5574_), .A3(new_n5573_), .ZN(new_n5575_));
  OAI21_X1   g04573(.A1(new_n1886_), .A2(new_n1946_), .B(new_n1938_), .ZN(new_n5576_));
  NAND3_X1   g04574(.A1(new_n5575_), .A2(new_n5569_), .A3(new_n5576_), .ZN(new_n5577_));
  AOI21_X1   g04575(.A1(new_n5574_), .A2(new_n5573_), .B(new_n5572_), .ZN(new_n5578_));
  NOR3_X1    g04576(.A1(new_n5565_), .A2(new_n5568_), .A3(new_n5555_), .ZN(new_n5579_));
  AOI21_X1   g04577(.A1(new_n1945_), .A2(new_n1929_), .B(new_n1947_), .ZN(new_n5580_));
  OAI21_X1   g04578(.A1(new_n5578_), .A2(new_n5579_), .B(new_n5580_), .ZN(new_n5581_));
  OAI21_X1   g04579(.A1(new_n2041_), .A2(new_n2042_), .B(new_n2030_), .ZN(new_n5582_));
  NOR2_X1    g04580(.A1(new_n2016_), .A2(new_n1993_), .ZN(new_n5583_));
  NOR2_X1    g04581(.A1(new_n2001_), .A2(new_n2023_), .ZN(new_n5584_));
  AOI21_X1   g04582(.A1(new_n2001_), .A2(new_n2023_), .B(new_n2022_), .ZN(new_n5585_));
  INV_X1     g04583(.I(new_n1991_), .ZN(new_n5586_));
  AOI21_X1   g04584(.A1(new_n1985_), .A2(new_n5586_), .B(new_n1990_), .ZN(new_n5587_));
  OAI21_X1   g04585(.A1(new_n5584_), .A2(new_n5585_), .B(new_n5587_), .ZN(new_n5588_));
  INV_X1     g04586(.I(new_n5584_), .ZN(new_n5589_));
  OAI21_X1   g04587(.A1(new_n1994_), .A2(new_n1998_), .B(new_n1996_), .ZN(new_n5590_));
  INV_X1     g04588(.I(new_n1990_), .ZN(new_n5591_));
  OAI21_X1   g04589(.A1(new_n2012_), .A2(new_n1991_), .B(new_n5591_), .ZN(new_n5592_));
  NAND3_X1   g04590(.A1(new_n5589_), .A2(new_n5590_), .A3(new_n5592_), .ZN(new_n5593_));
  NAND2_X1   g04591(.A1(new_n5593_), .A2(new_n5588_), .ZN(new_n5594_));
  OAI21_X1   g04592(.A1(new_n5583_), .A2(new_n2026_), .B(new_n5594_), .ZN(new_n5595_));
  NAND2_X1   g04593(.A1(new_n2006_), .A2(new_n2013_), .ZN(new_n5596_));
  AOI21_X1   g04594(.A1(new_n5589_), .A2(new_n5590_), .B(new_n5592_), .ZN(new_n5597_));
  NOR3_X1    g04595(.A1(new_n5585_), .A2(new_n5587_), .A3(new_n5584_), .ZN(new_n5598_));
  NOR2_X1    g04596(.A1(new_n5597_), .A2(new_n5598_), .ZN(new_n5599_));
  NAND3_X1   g04597(.A1(new_n5596_), .A2(new_n2010_), .A3(new_n5599_), .ZN(new_n5600_));
  NOR2_X1    g04598(.A1(new_n1966_), .A2(new_n1977_), .ZN(new_n5601_));
  AOI21_X1   g04599(.A1(new_n1966_), .A2(new_n1977_), .B(new_n1976_), .ZN(new_n5602_));
  INV_X1     g04600(.I(new_n1954_), .ZN(new_n5603_));
  AOI21_X1   g04601(.A1(new_n1951_), .A2(new_n1956_), .B(new_n5603_), .ZN(new_n5604_));
  OAI21_X1   g04602(.A1(new_n5602_), .A2(new_n5601_), .B(new_n5604_), .ZN(new_n5605_));
  NAND2_X1   g04603(.A1(new_n1959_), .A2(new_n1963_), .ZN(new_n5606_));
  OAI21_X1   g04604(.A1(new_n1959_), .A2(new_n1963_), .B(new_n1961_), .ZN(new_n5607_));
  OAI21_X1   g04605(.A1(new_n2032_), .A2(new_n1955_), .B(new_n1954_), .ZN(new_n5608_));
  NAND3_X1   g04606(.A1(new_n5607_), .A2(new_n5608_), .A3(new_n5606_), .ZN(new_n5609_));
  NAND2_X1   g04607(.A1(new_n5609_), .A2(new_n5605_), .ZN(new_n5610_));
  OAI21_X1   g04608(.A1(new_n2034_), .A2(new_n1980_), .B(new_n5610_), .ZN(new_n5611_));
  AOI21_X1   g04609(.A1(new_n5607_), .A2(new_n5606_), .B(new_n5608_), .ZN(new_n5612_));
  NOR3_X1    g04610(.A1(new_n5602_), .A2(new_n5604_), .A3(new_n5601_), .ZN(new_n5613_));
  NOR2_X1    g04611(.A1(new_n5612_), .A2(new_n5613_), .ZN(new_n5614_));
  NAND3_X1   g04612(.A1(new_n1972_), .A2(new_n5614_), .A3(new_n2037_), .ZN(new_n5615_));
  NAND4_X1   g04613(.A1(new_n5600_), .A2(new_n5595_), .A3(new_n5611_), .A4(new_n5615_), .ZN(new_n5616_));
  AOI21_X1   g04614(.A1(new_n5596_), .A2(new_n2010_), .B(new_n5599_), .ZN(new_n5617_));
  NOR3_X1    g04615(.A1(new_n5583_), .A2(new_n2026_), .A3(new_n5594_), .ZN(new_n5618_));
  AOI21_X1   g04616(.A1(new_n1972_), .A2(new_n2037_), .B(new_n5614_), .ZN(new_n5619_));
  NOR3_X1    g04617(.A1(new_n2034_), .A2(new_n1980_), .A3(new_n5610_), .ZN(new_n5620_));
  OAI22_X1   g04618(.A1(new_n5617_), .A2(new_n5618_), .B1(new_n5620_), .B2(new_n5619_), .ZN(new_n5621_));
  NAND3_X1   g04619(.A1(new_n5582_), .A2(new_n5616_), .A3(new_n5621_), .ZN(new_n5622_));
  AOI21_X1   g04620(.A1(new_n1984_), .A2(new_n2020_), .B(new_n2043_), .ZN(new_n5623_));
  NOR4_X1    g04621(.A1(new_n5617_), .A2(new_n5618_), .A3(new_n5620_), .A4(new_n5619_), .ZN(new_n5624_));
  AOI22_X1   g04622(.A1(new_n5600_), .A2(new_n5595_), .B1(new_n5611_), .B2(new_n5615_), .ZN(new_n5625_));
  OAI21_X1   g04623(.A1(new_n5624_), .A2(new_n5625_), .B(new_n5623_), .ZN(new_n5626_));
  NAND4_X1   g04624(.A1(new_n5626_), .A2(new_n5581_), .A3(new_n5577_), .A4(new_n5622_), .ZN(new_n5627_));
  NOR3_X1    g04625(.A1(new_n5578_), .A2(new_n5579_), .A3(new_n5580_), .ZN(new_n5628_));
  AOI21_X1   g04626(.A1(new_n5575_), .A2(new_n5569_), .B(new_n5576_), .ZN(new_n5629_));
  NOR3_X1    g04627(.A1(new_n5623_), .A2(new_n5624_), .A3(new_n5625_), .ZN(new_n5630_));
  AOI21_X1   g04628(.A1(new_n5616_), .A2(new_n5621_), .B(new_n5582_), .ZN(new_n5631_));
  OAI22_X1   g04629(.A1(new_n5630_), .A2(new_n5631_), .B1(new_n5629_), .B2(new_n5628_), .ZN(new_n5632_));
  NAND3_X1   g04630(.A1(new_n5632_), .A2(new_n5627_), .A3(new_n5538_), .ZN(new_n5633_));
  AOI21_X1   g04631(.A1(new_n2045_), .A2(new_n1949_), .B(new_n2052_), .ZN(new_n5634_));
  NOR4_X1    g04632(.A1(new_n5631_), .A2(new_n5629_), .A3(new_n5628_), .A4(new_n5630_), .ZN(new_n5635_));
  AOI22_X1   g04633(.A1(new_n5626_), .A2(new_n5622_), .B1(new_n5581_), .B2(new_n5577_), .ZN(new_n5636_));
  OAI21_X1   g04634(.A1(new_n5636_), .A2(new_n5635_), .B(new_n5634_), .ZN(new_n5637_));
  NAND4_X1   g04635(.A1(new_n5637_), .A2(new_n5633_), .A3(new_n5537_), .A4(new_n5533_), .ZN(new_n5638_));
  NOR3_X1    g04636(.A1(new_n5535_), .A2(new_n5534_), .A3(new_n5536_), .ZN(new_n5639_));
  AOI21_X1   g04637(.A1(new_n5531_), .A2(new_n5526_), .B(new_n5532_), .ZN(new_n5640_));
  NOR3_X1    g04638(.A1(new_n5636_), .A2(new_n5635_), .A3(new_n5634_), .ZN(new_n5641_));
  AOI21_X1   g04639(.A1(new_n5632_), .A2(new_n5627_), .B(new_n5538_), .ZN(new_n5642_));
  OAI22_X1   g04640(.A1(new_n5641_), .A2(new_n5642_), .B1(new_n5639_), .B2(new_n5640_), .ZN(new_n5643_));
  NAND3_X1   g04641(.A1(new_n5643_), .A2(new_n5638_), .A3(new_n5429_), .ZN(new_n5644_));
  AOI21_X1   g04642(.A1(new_n1515_), .A2(new_n2054_), .B(new_n2063_), .ZN(new_n5645_));
  NOR4_X1    g04643(.A1(new_n5641_), .A2(new_n5642_), .A3(new_n5639_), .A4(new_n5640_), .ZN(new_n5646_));
  AOI22_X1   g04644(.A1(new_n5637_), .A2(new_n5633_), .B1(new_n5537_), .B2(new_n5533_), .ZN(new_n5647_));
  OAI21_X1   g04645(.A1(new_n5646_), .A2(new_n5647_), .B(new_n5645_), .ZN(new_n5648_));
  NAND4_X1   g04646(.A1(new_n5428_), .A2(new_n5424_), .A3(new_n5648_), .A4(new_n5644_), .ZN(new_n5649_));
  NOR3_X1    g04647(.A1(new_n5425_), .A2(new_n5426_), .A3(new_n5427_), .ZN(new_n5650_));
  AOI21_X1   g04648(.A1(new_n5422_), .A2(new_n5417_), .B(new_n5423_), .ZN(new_n5651_));
  NOR3_X1    g04649(.A1(new_n5646_), .A2(new_n5647_), .A3(new_n5645_), .ZN(new_n5652_));
  AOI21_X1   g04650(.A1(new_n5643_), .A2(new_n5638_), .B(new_n5429_), .ZN(new_n5653_));
  OAI22_X1   g04651(.A1(new_n5650_), .A2(new_n5651_), .B1(new_n5652_), .B2(new_n5653_), .ZN(new_n5654_));
  OAI21_X1   g04652(.A1(new_n3085_), .A2(new_n3081_), .B(new_n3086_), .ZN(new_n5655_));
  NAND3_X1   g04653(.A1(new_n5654_), .A2(new_n5649_), .A3(new_n5655_), .ZN(new_n5656_));
  NOR4_X1    g04654(.A1(new_n5650_), .A2(new_n5651_), .A3(new_n5652_), .A4(new_n5653_), .ZN(new_n5657_));
  AOI22_X1   g04655(.A1(new_n5428_), .A2(new_n5424_), .B1(new_n5648_), .B2(new_n5644_), .ZN(new_n5658_));
  AOI21_X1   g04656(.A1(new_n2065_), .A2(new_n3087_), .B(new_n3076_), .ZN(new_n5659_));
  OAI21_X1   g04657(.A1(new_n5657_), .A2(new_n5658_), .B(new_n5659_), .ZN(new_n5660_));
  OAI21_X1   g04658(.A1(new_n4771_), .A2(new_n5180_), .B(new_n5189_), .ZN(new_n5661_));
  AOI21_X1   g04659(.A1(new_n4689_), .A2(new_n4690_), .B(new_n4686_), .ZN(new_n5662_));
  NAND2_X1   g04660(.A1(new_n4673_), .A2(new_n4674_), .ZN(new_n5663_));
  NOR2_X1    g04661(.A1(new_n4673_), .A2(new_n4674_), .ZN(new_n5664_));
  AOI21_X1   g04662(.A1(new_n4232_), .A2(new_n5663_), .B(new_n5664_), .ZN(new_n5665_));
  AOI21_X1   g04663(.A1(new_n4281_), .A2(new_n4669_), .B(new_n4665_), .ZN(new_n5666_));
  NOR2_X1    g04664(.A1(new_n5665_), .A2(new_n5666_), .ZN(new_n5667_));
  INV_X1     g04665(.I(new_n5663_), .ZN(new_n5668_));
  INV_X1     g04666(.I(new_n5664_), .ZN(new_n5669_));
  OAI21_X1   g04667(.A1(new_n4278_), .A2(new_n5668_), .B(new_n5669_), .ZN(new_n5670_));
  OAI21_X1   g04668(.A1(new_n4264_), .A2(new_n4666_), .B(new_n4664_), .ZN(new_n5671_));
  NOR2_X1    g04669(.A1(new_n5670_), .A2(new_n5671_), .ZN(new_n5672_));
  NOR2_X1    g04670(.A1(new_n5667_), .A2(new_n5672_), .ZN(new_n5673_));
  OAI21_X1   g04671(.A1(new_n5662_), .A2(new_n4682_), .B(new_n5673_), .ZN(new_n5674_));
  OAI21_X1   g04672(.A1(new_n4679_), .A2(new_n4680_), .B(new_n4672_), .ZN(new_n5675_));
  NAND2_X1   g04673(.A1(new_n5670_), .A2(new_n5671_), .ZN(new_n5676_));
  NAND2_X1   g04674(.A1(new_n5665_), .A2(new_n5666_), .ZN(new_n5677_));
  NAND2_X1   g04675(.A1(new_n5677_), .A2(new_n5676_), .ZN(new_n5678_));
  NAND3_X1   g04676(.A1(new_n5675_), .A2(new_n5678_), .A3(new_n4692_), .ZN(new_n5679_));
  NAND2_X1   g04677(.A1(new_n5674_), .A2(new_n5679_), .ZN(new_n5680_));
  NOR4_X1    g04678(.A1(new_n4709_), .A2(new_n4711_), .A3(new_n4291_), .A4(new_n4301_), .ZN(new_n5681_));
  NOR2_X1    g04679(.A1(new_n4710_), .A2(new_n4712_), .ZN(new_n5682_));
  INV_X1     g04680(.I(new_n5682_), .ZN(new_n5683_));
  OAI21_X1   g04681(.A1(new_n4305_), .A2(new_n5681_), .B(new_n5683_), .ZN(new_n5684_));
  AOI21_X1   g04682(.A1(new_n4338_), .A2(new_n4705_), .B(new_n4699_), .ZN(new_n5685_));
  NOR3_X1    g04683(.A1(new_n4741_), .A2(new_n4725_), .A3(new_n5685_), .ZN(new_n5686_));
  INV_X1     g04684(.I(new_n5685_), .ZN(new_n5687_));
  AOI21_X1   g04685(.A1(new_n4724_), .A2(new_n4728_), .B(new_n5687_), .ZN(new_n5688_));
  NOR3_X1    g04686(.A1(new_n5686_), .A2(new_n5688_), .A3(new_n5684_), .ZN(new_n5689_));
  INV_X1     g04687(.I(new_n5684_), .ZN(new_n5690_));
  NAND3_X1   g04688(.A1(new_n4724_), .A2(new_n4728_), .A3(new_n5687_), .ZN(new_n5691_));
  OAI21_X1   g04689(.A1(new_n4741_), .A2(new_n4725_), .B(new_n5685_), .ZN(new_n5692_));
  AOI21_X1   g04690(.A1(new_n5692_), .A2(new_n5691_), .B(new_n5690_), .ZN(new_n5693_));
  OAI21_X1   g04691(.A1(new_n5689_), .A2(new_n5693_), .B(new_n5680_), .ZN(new_n5694_));
  AOI21_X1   g04692(.A1(new_n5675_), .A2(new_n4692_), .B(new_n5678_), .ZN(new_n5695_));
  NOR3_X1    g04693(.A1(new_n5662_), .A2(new_n5673_), .A3(new_n4682_), .ZN(new_n5696_));
  NOR2_X1    g04694(.A1(new_n5695_), .A2(new_n5696_), .ZN(new_n5697_));
  NAND3_X1   g04695(.A1(new_n5692_), .A2(new_n5691_), .A3(new_n5690_), .ZN(new_n5698_));
  OAI21_X1   g04696(.A1(new_n5686_), .A2(new_n5688_), .B(new_n5684_), .ZN(new_n5699_));
  NAND3_X1   g04697(.A1(new_n5697_), .A2(new_n5699_), .A3(new_n5698_), .ZN(new_n5700_));
  OAI21_X1   g04698(.A1(new_n4749_), .A2(new_n4730_), .B(new_n4751_), .ZN(new_n5701_));
  NAND3_X1   g04699(.A1(new_n5694_), .A2(new_n5700_), .A3(new_n5701_), .ZN(new_n5702_));
  AOI21_X1   g04700(.A1(new_n5699_), .A2(new_n5698_), .B(new_n5697_), .ZN(new_n5703_));
  NOR3_X1    g04701(.A1(new_n5693_), .A2(new_n5689_), .A3(new_n5680_), .ZN(new_n5704_));
  AOI21_X1   g04702(.A1(new_n4694_), .A2(new_n4750_), .B(new_n4745_), .ZN(new_n5705_));
  OAI21_X1   g04703(.A1(new_n5703_), .A2(new_n5704_), .B(new_n5705_), .ZN(new_n5706_));
  OAI21_X1   g04704(.A1(new_n4656_), .A2(new_n4657_), .B(new_n4644_), .ZN(new_n5707_));
  NAND2_X1   g04705(.A1(new_n4629_), .A2(new_n4627_), .ZN(new_n5708_));
  NAND2_X1   g04706(.A1(new_n4127_), .A2(new_n4123_), .ZN(new_n5709_));
  AOI21_X1   g04707(.A1(new_n5708_), .A2(new_n5709_), .B(new_n4635_), .ZN(new_n5710_));
  NAND2_X1   g04708(.A1(new_n4624_), .A2(new_n4622_), .ZN(new_n5711_));
  NOR2_X1    g04709(.A1(new_n4624_), .A2(new_n4622_), .ZN(new_n5712_));
  AOI21_X1   g04710(.A1(new_n4078_), .A2(new_n5711_), .B(new_n5712_), .ZN(new_n5713_));
  AOI21_X1   g04711(.A1(new_n4128_), .A2(new_n4616_), .B(new_n4612_), .ZN(new_n5714_));
  NOR2_X1    g04712(.A1(new_n5713_), .A2(new_n5714_), .ZN(new_n5715_));
  INV_X1     g04713(.I(new_n5711_), .ZN(new_n5716_));
  INV_X1     g04714(.I(new_n5712_), .ZN(new_n5717_));
  OAI21_X1   g04715(.A1(new_n4125_), .A2(new_n5716_), .B(new_n5717_), .ZN(new_n5718_));
  OAI21_X1   g04716(.A1(new_n4110_), .A2(new_n4613_), .B(new_n4611_), .ZN(new_n5719_));
  NOR2_X1    g04717(.A1(new_n5718_), .A2(new_n5719_), .ZN(new_n5720_));
  NOR2_X1    g04718(.A1(new_n5715_), .A2(new_n5720_), .ZN(new_n5721_));
  OAI21_X1   g04719(.A1(new_n5710_), .A2(new_n4631_), .B(new_n5721_), .ZN(new_n5722_));
  NOR2_X1    g04720(.A1(new_n4636_), .A2(new_n4637_), .ZN(new_n5723_));
  NOR2_X1    g04721(.A1(new_n4090_), .A2(new_n4130_), .ZN(new_n5724_));
  OAI21_X1   g04722(.A1(new_n5723_), .A2(new_n5724_), .B(new_n4619_), .ZN(new_n5725_));
  NAND2_X1   g04723(.A1(new_n5718_), .A2(new_n5719_), .ZN(new_n5726_));
  NAND2_X1   g04724(.A1(new_n5713_), .A2(new_n5714_), .ZN(new_n5727_));
  NAND2_X1   g04725(.A1(new_n5727_), .A2(new_n5726_), .ZN(new_n5728_));
  NAND3_X1   g04726(.A1(new_n5725_), .A2(new_n5728_), .A3(new_n4639_), .ZN(new_n5729_));
  NAND2_X1   g04727(.A1(new_n5722_), .A2(new_n5729_), .ZN(new_n5730_));
  NOR4_X1    g04728(.A1(new_n4588_), .A2(new_n4590_), .A3(new_n4138_), .A4(new_n4148_), .ZN(new_n5731_));
  NOR2_X1    g04729(.A1(new_n4589_), .A2(new_n4591_), .ZN(new_n5732_));
  INV_X1     g04730(.I(new_n5732_), .ZN(new_n5733_));
  OAI21_X1   g04731(.A1(new_n4199_), .A2(new_n5731_), .B(new_n5733_), .ZN(new_n5734_));
  AOI21_X1   g04732(.A1(new_n4202_), .A2(new_n4584_), .B(new_n4579_), .ZN(new_n5735_));
  NOR3_X1    g04733(.A1(new_n4653_), .A2(new_n4601_), .A3(new_n5735_), .ZN(new_n5736_));
  INV_X1     g04734(.I(new_n5735_), .ZN(new_n5737_));
  AOI21_X1   g04735(.A1(new_n4600_), .A2(new_n4654_), .B(new_n5737_), .ZN(new_n5738_));
  NOR3_X1    g04736(.A1(new_n5736_), .A2(new_n5738_), .A3(new_n5734_), .ZN(new_n5739_));
  INV_X1     g04737(.I(new_n5734_), .ZN(new_n5740_));
  NAND3_X1   g04738(.A1(new_n4600_), .A2(new_n4654_), .A3(new_n5737_), .ZN(new_n5741_));
  OAI21_X1   g04739(.A1(new_n4653_), .A2(new_n4601_), .B(new_n5735_), .ZN(new_n5742_));
  AOI21_X1   g04740(.A1(new_n5742_), .A2(new_n5741_), .B(new_n5740_), .ZN(new_n5743_));
  OAI21_X1   g04741(.A1(new_n5739_), .A2(new_n5743_), .B(new_n5730_), .ZN(new_n5744_));
  AOI21_X1   g04742(.A1(new_n5725_), .A2(new_n4639_), .B(new_n5728_), .ZN(new_n5745_));
  NOR3_X1    g04743(.A1(new_n5710_), .A2(new_n5721_), .A3(new_n4631_), .ZN(new_n5746_));
  NOR2_X1    g04744(.A1(new_n5746_), .A2(new_n5745_), .ZN(new_n5747_));
  NAND3_X1   g04745(.A1(new_n5742_), .A2(new_n5741_), .A3(new_n5740_), .ZN(new_n5748_));
  OAI21_X1   g04746(.A1(new_n5736_), .A2(new_n5738_), .B(new_n5734_), .ZN(new_n5749_));
  NAND3_X1   g04747(.A1(new_n5747_), .A2(new_n5749_), .A3(new_n5748_), .ZN(new_n5750_));
  NAND3_X1   g04748(.A1(new_n5744_), .A2(new_n5750_), .A3(new_n5707_), .ZN(new_n5751_));
  AOI21_X1   g04749(.A1(new_n4605_), .A2(new_n4641_), .B(new_n4658_), .ZN(new_n5752_));
  AOI21_X1   g04750(.A1(new_n5748_), .A2(new_n5749_), .B(new_n5747_), .ZN(new_n5753_));
  NOR3_X1    g04751(.A1(new_n5739_), .A2(new_n5743_), .A3(new_n5730_), .ZN(new_n5754_));
  OAI21_X1   g04752(.A1(new_n5753_), .A2(new_n5754_), .B(new_n5752_), .ZN(new_n5755_));
  NAND4_X1   g04753(.A1(new_n5706_), .A2(new_n5702_), .A3(new_n5755_), .A4(new_n5751_), .ZN(new_n5756_));
  NOR3_X1    g04754(.A1(new_n5703_), .A2(new_n5704_), .A3(new_n5705_), .ZN(new_n5757_));
  AOI21_X1   g04755(.A1(new_n5694_), .A2(new_n5700_), .B(new_n5701_), .ZN(new_n5758_));
  NOR3_X1    g04756(.A1(new_n5753_), .A2(new_n5754_), .A3(new_n5752_), .ZN(new_n5759_));
  AOI21_X1   g04757(.A1(new_n5744_), .A2(new_n5750_), .B(new_n5707_), .ZN(new_n5760_));
  OAI22_X1   g04758(.A1(new_n5757_), .A2(new_n5758_), .B1(new_n5759_), .B2(new_n5760_), .ZN(new_n5761_));
  OAI21_X1   g04759(.A1(new_n4660_), .A2(new_n4753_), .B(new_n4759_), .ZN(new_n5762_));
  NAND3_X1   g04760(.A1(new_n5761_), .A2(new_n5762_), .A3(new_n5756_), .ZN(new_n5763_));
  NOR4_X1    g04761(.A1(new_n5757_), .A2(new_n5758_), .A3(new_n5759_), .A4(new_n5760_), .ZN(new_n5764_));
  AOI22_X1   g04762(.A1(new_n5706_), .A2(new_n5702_), .B1(new_n5755_), .B2(new_n5751_), .ZN(new_n5765_));
  AOI21_X1   g04763(.A1(new_n4661_), .A2(new_n4758_), .B(new_n4756_), .ZN(new_n5766_));
  OAI21_X1   g04764(.A1(new_n5764_), .A2(new_n5765_), .B(new_n5766_), .ZN(new_n5767_));
  INV_X1     g04765(.I(new_n4471_), .ZN(new_n5768_));
  NOR2_X1    g04766(.A1(new_n5768_), .A2(new_n4469_), .ZN(new_n5769_));
  NAND3_X1   g04767(.A1(new_n4549_), .A2(new_n4564_), .A3(new_n4055_), .ZN(new_n5770_));
  OAI21_X1   g04768(.A1(new_n5769_), .A2(new_n4565_), .B(new_n5770_), .ZN(new_n5771_));
  NOR2_X1    g04769(.A1(new_n4000_), .A2(new_n4011_), .ZN(new_n5772_));
  AND3_X2    g04770(.A1(new_n4414_), .A2(new_n5772_), .A3(new_n4413_), .Z(new_n5773_));
  AOI22_X1   g04771(.A1(new_n4406_), .A2(new_n4049_), .B1(new_n4380_), .B2(new_n4384_), .ZN(new_n5774_));
  NOR2_X1    g04772(.A1(new_n4393_), .A2(new_n4391_), .ZN(new_n5775_));
  AOI21_X1   g04773(.A1(new_n4047_), .A2(new_n4411_), .B(new_n5775_), .ZN(new_n5776_));
  AOI21_X1   g04774(.A1(new_n4045_), .A2(new_n4382_), .B(new_n4377_), .ZN(new_n5777_));
  NOR2_X1    g04775(.A1(new_n5776_), .A2(new_n5777_), .ZN(new_n5778_));
  INV_X1     g04776(.I(new_n5775_), .ZN(new_n5779_));
  OAI21_X1   g04777(.A1(new_n4032_), .A2(new_n4412_), .B(new_n5779_), .ZN(new_n5780_));
  OAI21_X1   g04778(.A1(new_n4000_), .A2(new_n4378_), .B(new_n4381_), .ZN(new_n5781_));
  NOR2_X1    g04779(.A1(new_n5780_), .A2(new_n5781_), .ZN(new_n5782_));
  NOR2_X1    g04780(.A1(new_n5782_), .A2(new_n5778_), .ZN(new_n5783_));
  OAI21_X1   g04781(.A1(new_n5773_), .A2(new_n5774_), .B(new_n5783_), .ZN(new_n5784_));
  OAI21_X1   g04782(.A1(new_n4386_), .A2(new_n4398_), .B(new_n4385_), .ZN(new_n5785_));
  NAND2_X1   g04783(.A1(new_n5780_), .A2(new_n5781_), .ZN(new_n5786_));
  NAND2_X1   g04784(.A1(new_n5776_), .A2(new_n5777_), .ZN(new_n5787_));
  NAND2_X1   g04785(.A1(new_n5786_), .A2(new_n5787_), .ZN(new_n5788_));
  NAND3_X1   g04786(.A1(new_n5785_), .A2(new_n5788_), .A3(new_n4415_), .ZN(new_n5789_));
  NAND2_X1   g04787(.A1(new_n5784_), .A2(new_n5789_), .ZN(new_n5790_));
  NAND2_X1   g04788(.A1(new_n4441_), .A2(new_n4439_), .ZN(new_n5791_));
  NAND2_X1   g04789(.A1(new_n3974_), .A2(new_n3970_), .ZN(new_n5792_));
  AOI21_X1   g04790(.A1(new_n5792_), .A2(new_n5791_), .B(new_n4431_), .ZN(new_n5793_));
  AOI21_X1   g04791(.A1(new_n3975_), .A2(new_n4424_), .B(new_n4427_), .ZN(new_n5794_));
  NOR3_X1    g04792(.A1(new_n5793_), .A2(new_n4447_), .A3(new_n5794_), .ZN(new_n5795_));
  NOR2_X1    g04793(.A1(new_n4454_), .A2(new_n4455_), .ZN(new_n5796_));
  NOR4_X1    g04794(.A1(new_n3972_), .A2(new_n3969_), .A3(new_n3973_), .A4(new_n3957_), .ZN(new_n5797_));
  OAI21_X1   g04795(.A1(new_n5796_), .A2(new_n5797_), .B(new_n4453_), .ZN(new_n5798_));
  INV_X1     g04796(.I(new_n5794_), .ZN(new_n5799_));
  AOI21_X1   g04797(.A1(new_n5798_), .A2(new_n4465_), .B(new_n5799_), .ZN(new_n5800_));
  NOR3_X1    g04798(.A1(new_n5795_), .A2(new_n5800_), .A3(new_n4464_), .ZN(new_n5801_));
  NAND3_X1   g04799(.A1(new_n5798_), .A2(new_n4465_), .A3(new_n5799_), .ZN(new_n5802_));
  OAI21_X1   g04800(.A1(new_n5793_), .A2(new_n4447_), .B(new_n5794_), .ZN(new_n5803_));
  AOI21_X1   g04801(.A1(new_n5803_), .A2(new_n5802_), .B(new_n4446_), .ZN(new_n5804_));
  OAI21_X1   g04802(.A1(new_n5801_), .A2(new_n5804_), .B(new_n5790_), .ZN(new_n5805_));
  AOI21_X1   g04803(.A1(new_n5785_), .A2(new_n4415_), .B(new_n5788_), .ZN(new_n5806_));
  NOR3_X1    g04804(.A1(new_n5774_), .A2(new_n5783_), .A3(new_n5773_), .ZN(new_n5807_));
  NOR2_X1    g04805(.A1(new_n5806_), .A2(new_n5807_), .ZN(new_n5808_));
  NAND3_X1   g04806(.A1(new_n5803_), .A2(new_n5802_), .A3(new_n4446_), .ZN(new_n5809_));
  OAI21_X1   g04807(.A1(new_n5795_), .A2(new_n5800_), .B(new_n4464_), .ZN(new_n5810_));
  NAND3_X1   g04808(.A1(new_n5808_), .A2(new_n5810_), .A3(new_n5809_), .ZN(new_n5811_));
  OR2_X2     g04809(.A1(new_n4408_), .A2(new_n4416_), .Z(new_n5812_));
  OAI22_X1   g04810(.A1(new_n4459_), .A2(new_n4448_), .B1(new_n4418_), .B2(new_n4050_), .ZN(new_n5813_));
  OAI21_X1   g04811(.A1(new_n5812_), .A2(new_n4460_), .B(new_n5813_), .ZN(new_n5814_));
  NAND3_X1   g04812(.A1(new_n5805_), .A2(new_n5811_), .A3(new_n5814_), .ZN(new_n5815_));
  AOI21_X1   g04813(.A1(new_n5810_), .A2(new_n5809_), .B(new_n5808_), .ZN(new_n5816_));
  NOR3_X1    g04814(.A1(new_n5801_), .A2(new_n5804_), .A3(new_n5790_), .ZN(new_n5817_));
  NAND3_X1   g04815(.A1(new_n4053_), .A2(new_n4466_), .A3(new_n4467_), .ZN(new_n5818_));
  AOI21_X1   g04816(.A1(new_n4417_), .A2(new_n5818_), .B(new_n4468_), .ZN(new_n5819_));
  OAI21_X1   g04817(.A1(new_n5816_), .A2(new_n5817_), .B(new_n5819_), .ZN(new_n5820_));
  OAI21_X1   g04818(.A1(new_n4503_), .A2(new_n4540_), .B(new_n4563_), .ZN(new_n5821_));
  NOR2_X1    g04819(.A1(new_n4526_), .A2(new_n4534_), .ZN(new_n5822_));
  NOR2_X1    g04820(.A1(new_n4514_), .A2(new_n4529_), .ZN(new_n5823_));
  AOI21_X1   g04821(.A1(new_n4514_), .A2(new_n4529_), .B(new_n4528_), .ZN(new_n5824_));
  INV_X1     g04822(.I(new_n4511_), .ZN(new_n5825_));
  AOI21_X1   g04823(.A1(new_n4505_), .A2(new_n5825_), .B(new_n4510_), .ZN(new_n5826_));
  OAI21_X1   g04824(.A1(new_n5823_), .A2(new_n5824_), .B(new_n5826_), .ZN(new_n5827_));
  NOR2_X1    g04825(.A1(new_n5824_), .A2(new_n5823_), .ZN(new_n5828_));
  INV_X1     g04826(.I(new_n5826_), .ZN(new_n5829_));
  NAND2_X1   g04827(.A1(new_n5828_), .A2(new_n5829_), .ZN(new_n5830_));
  NAND2_X1   g04828(.A1(new_n5830_), .A2(new_n5827_), .ZN(new_n5831_));
  OAI21_X1   g04829(.A1(new_n5822_), .A2(new_n4532_), .B(new_n5831_), .ZN(new_n5832_));
  OAI21_X1   g04830(.A1(new_n3817_), .A2(new_n4541_), .B(new_n4513_), .ZN(new_n5833_));
  NOR2_X1    g04831(.A1(new_n5828_), .A2(new_n5829_), .ZN(new_n5834_));
  NOR3_X1    g04832(.A1(new_n5824_), .A2(new_n5826_), .A3(new_n5823_), .ZN(new_n5835_));
  NOR2_X1    g04833(.A1(new_n5834_), .A2(new_n5835_), .ZN(new_n5836_));
  NAND3_X1   g04834(.A1(new_n5833_), .A2(new_n5836_), .A3(new_n4544_), .ZN(new_n5837_));
  NOR2_X1    g04835(.A1(new_n4480_), .A2(new_n4554_), .ZN(new_n5838_));
  AOI21_X1   g04836(.A1(new_n4480_), .A2(new_n4554_), .B(new_n4553_), .ZN(new_n5839_));
  INV_X1     g04837(.I(new_n4476_), .ZN(new_n5840_));
  AOI21_X1   g04838(.A1(new_n4550_), .A2(new_n4477_), .B(new_n5840_), .ZN(new_n5841_));
  OAI21_X1   g04839(.A1(new_n5838_), .A2(new_n5839_), .B(new_n5841_), .ZN(new_n5842_));
  NAND2_X1   g04840(.A1(new_n4489_), .A2(new_n4483_), .ZN(new_n5843_));
  OAI21_X1   g04841(.A1(new_n4489_), .A2(new_n4483_), .B(new_n4485_), .ZN(new_n5844_));
  INV_X1     g04842(.I(new_n4477_), .ZN(new_n5845_));
  OAI21_X1   g04843(.A1(new_n4473_), .A2(new_n5845_), .B(new_n4476_), .ZN(new_n5846_));
  NAND3_X1   g04844(.A1(new_n5844_), .A2(new_n5846_), .A3(new_n5843_), .ZN(new_n5847_));
  NAND2_X1   g04845(.A1(new_n5847_), .A2(new_n5842_), .ZN(new_n5848_));
  OAI21_X1   g04846(.A1(new_n4493_), .A2(new_n4557_), .B(new_n5848_), .ZN(new_n5849_));
  AOI21_X1   g04847(.A1(new_n5843_), .A2(new_n5844_), .B(new_n5846_), .ZN(new_n5850_));
  NOR3_X1    g04848(.A1(new_n5839_), .A2(new_n5841_), .A3(new_n5838_), .ZN(new_n5851_));
  NOR2_X1    g04849(.A1(new_n5850_), .A2(new_n5851_), .ZN(new_n5852_));
  NAND3_X1   g04850(.A1(new_n4552_), .A2(new_n5852_), .A3(new_n4499_), .ZN(new_n5853_));
  NAND4_X1   g04851(.A1(new_n5832_), .A2(new_n5837_), .A3(new_n5849_), .A4(new_n5853_), .ZN(new_n5854_));
  AOI21_X1   g04852(.A1(new_n4544_), .A2(new_n5833_), .B(new_n5836_), .ZN(new_n5855_));
  NOR3_X1    g04853(.A1(new_n5822_), .A2(new_n5831_), .A3(new_n4532_), .ZN(new_n5856_));
  AOI21_X1   g04854(.A1(new_n4552_), .A2(new_n4499_), .B(new_n5852_), .ZN(new_n5857_));
  NOR3_X1    g04855(.A1(new_n4493_), .A2(new_n4557_), .A3(new_n5848_), .ZN(new_n5858_));
  OAI22_X1   g04856(.A1(new_n5855_), .A2(new_n5856_), .B1(new_n5858_), .B2(new_n5857_), .ZN(new_n5859_));
  NAND3_X1   g04857(.A1(new_n5821_), .A2(new_n5854_), .A3(new_n5859_), .ZN(new_n5860_));
  AOI21_X1   g04858(.A1(new_n4561_), .A2(new_n4562_), .B(new_n4548_), .ZN(new_n5861_));
  NOR4_X1    g04859(.A1(new_n5855_), .A2(new_n5856_), .A3(new_n5858_), .A4(new_n5857_), .ZN(new_n5862_));
  AOI22_X1   g04860(.A1(new_n5832_), .A2(new_n5837_), .B1(new_n5849_), .B2(new_n5853_), .ZN(new_n5863_));
  OAI21_X1   g04861(.A1(new_n5862_), .A2(new_n5863_), .B(new_n5861_), .ZN(new_n5864_));
  NAND4_X1   g04862(.A1(new_n5864_), .A2(new_n5815_), .A3(new_n5820_), .A4(new_n5860_), .ZN(new_n5865_));
  NOR3_X1    g04863(.A1(new_n5816_), .A2(new_n5817_), .A3(new_n5819_), .ZN(new_n5866_));
  AOI21_X1   g04864(.A1(new_n5811_), .A2(new_n5805_), .B(new_n5814_), .ZN(new_n5867_));
  NOR3_X1    g04865(.A1(new_n5861_), .A2(new_n5862_), .A3(new_n5863_), .ZN(new_n5868_));
  AOI21_X1   g04866(.A1(new_n5854_), .A2(new_n5859_), .B(new_n5821_), .ZN(new_n5869_));
  OAI22_X1   g04867(.A1(new_n5868_), .A2(new_n5869_), .B1(new_n5867_), .B2(new_n5866_), .ZN(new_n5870_));
  NAND3_X1   g04868(.A1(new_n5870_), .A2(new_n5865_), .A3(new_n5771_), .ZN(new_n5871_));
  AOI21_X1   g04869(.A1(new_n4571_), .A2(new_n4472_), .B(new_n4568_), .ZN(new_n5872_));
  NOR4_X1    g04870(.A1(new_n5867_), .A2(new_n5869_), .A3(new_n5866_), .A4(new_n5868_), .ZN(new_n5873_));
  AOI22_X1   g04871(.A1(new_n5860_), .A2(new_n5864_), .B1(new_n5815_), .B2(new_n5820_), .ZN(new_n5874_));
  OAI21_X1   g04872(.A1(new_n5874_), .A2(new_n5873_), .B(new_n5872_), .ZN(new_n5875_));
  NAND4_X1   g04873(.A1(new_n5763_), .A2(new_n5767_), .A3(new_n5875_), .A4(new_n5871_), .ZN(new_n5876_));
  NOR3_X1    g04874(.A1(new_n5764_), .A2(new_n5765_), .A3(new_n5766_), .ZN(new_n5877_));
  AOI21_X1   g04875(.A1(new_n5761_), .A2(new_n5756_), .B(new_n5762_), .ZN(new_n5878_));
  NOR3_X1    g04876(.A1(new_n5874_), .A2(new_n5873_), .A3(new_n5872_), .ZN(new_n5879_));
  AOI21_X1   g04877(.A1(new_n5870_), .A2(new_n5865_), .B(new_n5771_), .ZN(new_n5880_));
  OAI22_X1   g04878(.A1(new_n5878_), .A2(new_n5877_), .B1(new_n5879_), .B2(new_n5880_), .ZN(new_n5881_));
  OAI21_X1   g04879(.A1(new_n4767_), .A2(new_n4761_), .B(new_n4769_), .ZN(new_n5882_));
  NAND3_X1   g04880(.A1(new_n5881_), .A2(new_n5876_), .A3(new_n5882_), .ZN(new_n5883_));
  NOR4_X1    g04881(.A1(new_n5878_), .A2(new_n5877_), .A3(new_n5879_), .A4(new_n5880_), .ZN(new_n5884_));
  AOI22_X1   g04882(.A1(new_n5763_), .A2(new_n5767_), .B1(new_n5875_), .B2(new_n5871_), .ZN(new_n5885_));
  AOI21_X1   g04883(.A1(new_n4574_), .A2(new_n4768_), .B(new_n4765_), .ZN(new_n5886_));
  OAI21_X1   g04884(.A1(new_n5884_), .A2(new_n5885_), .B(new_n5886_), .ZN(new_n5887_));
  OAI21_X1   g04885(.A1(new_n4965_), .A2(new_n5169_), .B(new_n5178_), .ZN(new_n5888_));
  NAND2_X1   g04886(.A1(new_n4891_), .A2(new_n4890_), .ZN(new_n5889_));
  NAND3_X1   g04887(.A1(new_n3122_), .A2(new_n3142_), .A3(new_n3145_), .ZN(new_n5890_));
  AOI21_X1   g04888(.A1(new_n5890_), .A2(new_n5889_), .B(new_n4878_), .ZN(new_n5891_));
  NOR4_X1    g04889(.A1(new_n4879_), .A2(new_n4881_), .A3(new_n3096_), .A4(new_n3106_), .ZN(new_n5892_));
  INV_X1     g04890(.I(new_n5892_), .ZN(new_n5893_));
  NAND2_X1   g04891(.A1(new_n3148_), .A2(new_n5893_), .ZN(new_n5894_));
  NOR2_X1    g04892(.A1(new_n4880_), .A2(new_n4882_), .ZN(new_n5895_));
  INV_X1     g04893(.I(new_n5895_), .ZN(new_n5896_));
  OAI21_X1   g04894(.A1(new_n3143_), .A2(new_n3144_), .B(new_n4871_), .ZN(new_n5897_));
  AOI22_X1   g04895(.A1(new_n5894_), .A2(new_n5896_), .B1(new_n5897_), .B2(new_n4868_), .ZN(new_n5898_));
  NOR2_X1    g04896(.A1(new_n3099_), .A2(new_n3095_), .ZN(new_n5899_));
  NOR2_X1    g04897(.A1(new_n3109_), .A2(new_n3105_), .ZN(new_n5900_));
  AOI21_X1   g04898(.A1(new_n5899_), .A2(new_n5900_), .B(new_n5892_), .ZN(new_n5901_));
  AOI21_X1   g04899(.A1(new_n3163_), .A2(new_n3164_), .B(new_n4875_), .ZN(new_n5902_));
  NOR4_X1    g04900(.A1(new_n5901_), .A2(new_n5902_), .A3(new_n4874_), .A4(new_n5895_), .ZN(new_n5903_));
  NOR2_X1    g04901(.A1(new_n5898_), .A2(new_n5903_), .ZN(new_n5904_));
  OAI21_X1   g04902(.A1(new_n5891_), .A2(new_n4900_), .B(new_n5904_), .ZN(new_n5905_));
  OAI21_X1   g04903(.A1(new_n4898_), .A2(new_n4892_), .B(new_n4897_), .ZN(new_n5906_));
  OAI22_X1   g04904(.A1(new_n5901_), .A2(new_n5895_), .B1(new_n5902_), .B2(new_n4874_), .ZN(new_n5907_));
  NAND4_X1   g04905(.A1(new_n5894_), .A2(new_n5897_), .A3(new_n4868_), .A4(new_n5896_), .ZN(new_n5908_));
  NAND2_X1   g04906(.A1(new_n5907_), .A2(new_n5908_), .ZN(new_n5909_));
  NAND3_X1   g04907(.A1(new_n5906_), .A2(new_n5909_), .A3(new_n4893_), .ZN(new_n5910_));
  NAND2_X1   g04908(.A1(new_n5905_), .A2(new_n5910_), .ZN(new_n5911_));
  NOR4_X1    g04909(.A1(new_n4920_), .A2(new_n4921_), .A3(new_n3174_), .A4(new_n3184_), .ZN(new_n5912_));
  NOR2_X1    g04910(.A1(new_n4924_), .A2(new_n4922_), .ZN(new_n5913_));
  INV_X1     g04911(.I(new_n5913_), .ZN(new_n5914_));
  OAI21_X1   g04912(.A1(new_n3188_), .A2(new_n5912_), .B(new_n5914_), .ZN(new_n5915_));
  NAND2_X1   g04913(.A1(new_n4933_), .A2(new_n4931_), .ZN(new_n5916_));
  AOI21_X1   g04914(.A1(new_n5916_), .A2(new_n4929_), .B(new_n4939_), .ZN(new_n5917_));
  AOI21_X1   g04915(.A1(new_n3221_), .A2(new_n4916_), .B(new_n4907_), .ZN(new_n5918_));
  NOR3_X1    g04916(.A1(new_n5917_), .A2(new_n4942_), .A3(new_n5918_), .ZN(new_n5919_));
  INV_X1     g04917(.I(new_n5918_), .ZN(new_n5920_));
  AOI21_X1   g04918(.A1(new_n4946_), .A2(new_n4935_), .B(new_n5920_), .ZN(new_n5921_));
  NOR3_X1    g04919(.A1(new_n5919_), .A2(new_n5921_), .A3(new_n5915_), .ZN(new_n5922_));
  INV_X1     g04920(.I(new_n5915_), .ZN(new_n5923_));
  NAND3_X1   g04921(.A1(new_n4946_), .A2(new_n4935_), .A3(new_n5920_), .ZN(new_n5924_));
  OAI21_X1   g04922(.A1(new_n5917_), .A2(new_n4942_), .B(new_n5918_), .ZN(new_n5925_));
  AOI21_X1   g04923(.A1(new_n5925_), .A2(new_n5924_), .B(new_n5923_), .ZN(new_n5926_));
  OAI21_X1   g04924(.A1(new_n5922_), .A2(new_n5926_), .B(new_n5911_), .ZN(new_n5927_));
  AOI21_X1   g04925(.A1(new_n5906_), .A2(new_n4893_), .B(new_n5909_), .ZN(new_n5928_));
  NOR3_X1    g04926(.A1(new_n5891_), .A2(new_n5904_), .A3(new_n4900_), .ZN(new_n5929_));
  NOR2_X1    g04927(.A1(new_n5928_), .A2(new_n5929_), .ZN(new_n5930_));
  NAND3_X1   g04928(.A1(new_n5925_), .A2(new_n5924_), .A3(new_n5923_), .ZN(new_n5931_));
  OAI21_X1   g04929(.A1(new_n5919_), .A2(new_n5921_), .B(new_n5915_), .ZN(new_n5932_));
  NAND3_X1   g04930(.A1(new_n5930_), .A2(new_n5932_), .A3(new_n5931_), .ZN(new_n5933_));
  OAI21_X1   g04931(.A1(new_n4902_), .A2(new_n4954_), .B(new_n4949_), .ZN(new_n5934_));
  NAND3_X1   g04932(.A1(new_n5933_), .A2(new_n5927_), .A3(new_n5934_), .ZN(new_n5935_));
  AOI21_X1   g04933(.A1(new_n5931_), .A2(new_n5932_), .B(new_n5930_), .ZN(new_n5936_));
  NOR3_X1    g04934(.A1(new_n5922_), .A2(new_n5926_), .A3(new_n5911_), .ZN(new_n5937_));
  AOI21_X1   g04935(.A1(new_n4953_), .A2(new_n4944_), .B(new_n4955_), .ZN(new_n5938_));
  OAI21_X1   g04936(.A1(new_n5936_), .A2(new_n5937_), .B(new_n5938_), .ZN(new_n5939_));
  OAI21_X1   g04937(.A1(new_n4862_), .A2(new_n4861_), .B(new_n4851_), .ZN(new_n5940_));
  OAI21_X1   g04938(.A1(new_n4831_), .A2(new_n4809_), .B(new_n4825_), .ZN(new_n5941_));
  NOR2_X1    g04939(.A1(new_n3376_), .A2(new_n4840_), .ZN(new_n5942_));
  AOI21_X1   g04940(.A1(new_n3376_), .A2(new_n4840_), .B(new_n4839_), .ZN(new_n5943_));
  INV_X1     g04941(.I(new_n4805_), .ZN(new_n5944_));
  AOI21_X1   g04942(.A1(new_n3396_), .A2(new_n4807_), .B(new_n5944_), .ZN(new_n5945_));
  OAI21_X1   g04943(.A1(new_n5942_), .A2(new_n5943_), .B(new_n5945_), .ZN(new_n5946_));
  NAND2_X1   g04944(.A1(new_n4818_), .A2(new_n4812_), .ZN(new_n5947_));
  OAI21_X1   g04945(.A1(new_n4818_), .A2(new_n4812_), .B(new_n4814_), .ZN(new_n5948_));
  OAI21_X1   g04946(.A1(new_n3344_), .A2(new_n4806_), .B(new_n4805_), .ZN(new_n5949_));
  NAND3_X1   g04947(.A1(new_n5948_), .A2(new_n5949_), .A3(new_n5947_), .ZN(new_n5950_));
  NAND2_X1   g04948(.A1(new_n5946_), .A2(new_n5950_), .ZN(new_n5951_));
  NAND2_X1   g04949(.A1(new_n5941_), .A2(new_n5951_), .ZN(new_n5952_));
  AOI21_X1   g04950(.A1(new_n4821_), .A2(new_n4827_), .B(new_n4843_), .ZN(new_n5953_));
  AOI21_X1   g04951(.A1(new_n5947_), .A2(new_n5948_), .B(new_n5949_), .ZN(new_n5954_));
  NOR3_X1    g04952(.A1(new_n5945_), .A2(new_n5943_), .A3(new_n5942_), .ZN(new_n5955_));
  NOR2_X1    g04953(.A1(new_n5954_), .A2(new_n5955_), .ZN(new_n5956_));
  NAND2_X1   g04954(.A1(new_n5953_), .A2(new_n5956_), .ZN(new_n5957_));
  OAI21_X1   g04955(.A1(new_n4796_), .A2(new_n4799_), .B(new_n4794_), .ZN(new_n5958_));
  NOR2_X1    g04956(.A1(new_n3303_), .A2(new_n4854_), .ZN(new_n5959_));
  AOI21_X1   g04957(.A1(new_n3303_), .A2(new_n4854_), .B(new_n4853_), .ZN(new_n5960_));
  NOR2_X1    g04958(.A1(new_n4772_), .A2(new_n3267_), .ZN(new_n5961_));
  NOR2_X1    g04959(.A1(new_n4773_), .A2(new_n3257_), .ZN(new_n5962_));
  NOR2_X1    g04960(.A1(new_n5961_), .A2(new_n5962_), .ZN(new_n5963_));
  AOI21_X1   g04961(.A1(new_n3317_), .A2(new_n4776_), .B(new_n5963_), .ZN(new_n5964_));
  OAI21_X1   g04962(.A1(new_n5960_), .A2(new_n5959_), .B(new_n5964_), .ZN(new_n5965_));
  NAND2_X1   g04963(.A1(new_n3320_), .A2(new_n4783_), .ZN(new_n5966_));
  OAI21_X1   g04964(.A1(new_n3320_), .A2(new_n4783_), .B(new_n4785_), .ZN(new_n5967_));
  OAI21_X1   g04965(.A1(new_n3270_), .A2(new_n4775_), .B(new_n4774_), .ZN(new_n5968_));
  NAND3_X1   g04966(.A1(new_n5968_), .A2(new_n5967_), .A3(new_n5966_), .ZN(new_n5969_));
  NAND2_X1   g04967(.A1(new_n5965_), .A2(new_n5969_), .ZN(new_n5970_));
  NAND2_X1   g04968(.A1(new_n5958_), .A2(new_n5970_), .ZN(new_n5971_));
  AOI21_X1   g04969(.A1(new_n4791_), .A2(new_n4780_), .B(new_n4857_), .ZN(new_n5972_));
  AOI21_X1   g04970(.A1(new_n5966_), .A2(new_n5967_), .B(new_n5968_), .ZN(new_n5973_));
  NOR3_X1    g04971(.A1(new_n5960_), .A2(new_n5964_), .A3(new_n5959_), .ZN(new_n5974_));
  NOR2_X1    g04972(.A1(new_n5973_), .A2(new_n5974_), .ZN(new_n5975_));
  NAND2_X1   g04973(.A1(new_n5972_), .A2(new_n5975_), .ZN(new_n5976_));
  NAND4_X1   g04974(.A1(new_n5971_), .A2(new_n5976_), .A3(new_n5952_), .A4(new_n5957_), .ZN(new_n5977_));
  NOR2_X1    g04975(.A1(new_n5953_), .A2(new_n5956_), .ZN(new_n5978_));
  NOR2_X1    g04976(.A1(new_n5941_), .A2(new_n5951_), .ZN(new_n5979_));
  NOR2_X1    g04977(.A1(new_n5972_), .A2(new_n5975_), .ZN(new_n5980_));
  NOR2_X1    g04978(.A1(new_n5958_), .A2(new_n5970_), .ZN(new_n5981_));
  OAI22_X1   g04979(.A1(new_n5981_), .A2(new_n5980_), .B1(new_n5979_), .B2(new_n5978_), .ZN(new_n5982_));
  NAND3_X1   g04980(.A1(new_n5982_), .A2(new_n5940_), .A3(new_n5977_), .ZN(new_n5983_));
  AOI21_X1   g04981(.A1(new_n4838_), .A2(new_n4802_), .B(new_n4863_), .ZN(new_n5984_));
  NOR4_X1    g04982(.A1(new_n5980_), .A2(new_n5981_), .A3(new_n5979_), .A4(new_n5978_), .ZN(new_n5985_));
  AOI22_X1   g04983(.A1(new_n5971_), .A2(new_n5976_), .B1(new_n5952_), .B2(new_n5957_), .ZN(new_n5986_));
  OAI21_X1   g04984(.A1(new_n5985_), .A2(new_n5986_), .B(new_n5984_), .ZN(new_n5987_));
  NAND4_X1   g04985(.A1(new_n5939_), .A2(new_n5935_), .A3(new_n5987_), .A4(new_n5983_), .ZN(new_n5988_));
  NOR3_X1    g04986(.A1(new_n5936_), .A2(new_n5937_), .A3(new_n5938_), .ZN(new_n5989_));
  AOI21_X1   g04987(.A1(new_n5933_), .A2(new_n5927_), .B(new_n5934_), .ZN(new_n5990_));
  NOR3_X1    g04988(.A1(new_n5984_), .A2(new_n5985_), .A3(new_n5986_), .ZN(new_n5991_));
  AOI21_X1   g04989(.A1(new_n5977_), .A2(new_n5982_), .B(new_n5940_), .ZN(new_n5992_));
  OAI22_X1   g04990(.A1(new_n5990_), .A2(new_n5989_), .B1(new_n5991_), .B2(new_n5992_), .ZN(new_n5993_));
  OR2_X2     g04991(.A1(new_n4864_), .A2(new_n4852_), .Z(new_n5994_));
  OAI21_X1   g04992(.A1(new_n4959_), .A2(new_n4960_), .B(new_n4958_), .ZN(new_n5995_));
  OAI21_X1   g04993(.A1(new_n5994_), .A2(new_n4961_), .B(new_n5995_), .ZN(new_n5996_));
  NAND3_X1   g04994(.A1(new_n5993_), .A2(new_n5988_), .A3(new_n5996_), .ZN(new_n5997_));
  NOR4_X1    g04995(.A1(new_n5990_), .A2(new_n5989_), .A3(new_n5991_), .A4(new_n5992_), .ZN(new_n5998_));
  AOI22_X1   g04996(.A1(new_n5939_), .A2(new_n5935_), .B1(new_n5987_), .B2(new_n5983_), .ZN(new_n5999_));
  NAND3_X1   g04997(.A1(new_n3402_), .A2(new_n4956_), .A3(new_n4950_), .ZN(new_n6000_));
  AOI21_X1   g04998(.A1(new_n4865_), .A2(new_n6000_), .B(new_n4957_), .ZN(new_n6001_));
  OAI21_X1   g04999(.A1(new_n5999_), .A2(new_n5998_), .B(new_n6001_), .ZN(new_n6002_));
  OAI21_X1   g05000(.A1(new_n5064_), .A2(new_n5156_), .B(new_n5167_), .ZN(new_n6003_));
  NOR2_X1    g05001(.A1(new_n3674_), .A2(new_n3685_), .ZN(new_n6004_));
  AND3_X2    g05002(.A1(new_n5007_), .A2(new_n6004_), .A3(new_n5006_), .Z(new_n6005_));
  AOI22_X1   g05003(.A1(new_n4999_), .A2(new_n3723_), .B1(new_n4973_), .B2(new_n4977_), .ZN(new_n6006_));
  NOR2_X1    g05004(.A1(new_n4986_), .A2(new_n4984_), .ZN(new_n6007_));
  AOI21_X1   g05005(.A1(new_n3721_), .A2(new_n5004_), .B(new_n6007_), .ZN(new_n6008_));
  AOI21_X1   g05006(.A1(new_n3719_), .A2(new_n4975_), .B(new_n4970_), .ZN(new_n6009_));
  NOR2_X1    g05007(.A1(new_n6008_), .A2(new_n6009_), .ZN(new_n6010_));
  INV_X1     g05008(.I(new_n6007_), .ZN(new_n6011_));
  OAI21_X1   g05009(.A1(new_n3706_), .A2(new_n5005_), .B(new_n6011_), .ZN(new_n6012_));
  OAI21_X1   g05010(.A1(new_n3674_), .A2(new_n4971_), .B(new_n4974_), .ZN(new_n6013_));
  NOR2_X1    g05011(.A1(new_n6012_), .A2(new_n6013_), .ZN(new_n6014_));
  NOR2_X1    g05012(.A1(new_n6014_), .A2(new_n6010_), .ZN(new_n6015_));
  OAI21_X1   g05013(.A1(new_n6005_), .A2(new_n6006_), .B(new_n6015_), .ZN(new_n6016_));
  OAI21_X1   g05014(.A1(new_n4979_), .A2(new_n4991_), .B(new_n4978_), .ZN(new_n6017_));
  NAND2_X1   g05015(.A1(new_n6012_), .A2(new_n6013_), .ZN(new_n6018_));
  NAND2_X1   g05016(.A1(new_n6008_), .A2(new_n6009_), .ZN(new_n6019_));
  NAND2_X1   g05017(.A1(new_n6018_), .A2(new_n6019_), .ZN(new_n6020_));
  NAND3_X1   g05018(.A1(new_n6017_), .A2(new_n6020_), .A3(new_n5008_), .ZN(new_n6021_));
  NAND2_X1   g05019(.A1(new_n6016_), .A2(new_n6021_), .ZN(new_n6022_));
  NAND2_X1   g05020(.A1(new_n5033_), .A2(new_n5031_), .ZN(new_n6023_));
  NAND2_X1   g05021(.A1(new_n3647_), .A2(new_n3643_), .ZN(new_n6024_));
  AOI21_X1   g05022(.A1(new_n6024_), .A2(new_n6023_), .B(new_n5023_), .ZN(new_n6025_));
  AOI21_X1   g05023(.A1(new_n3648_), .A2(new_n5016_), .B(new_n5019_), .ZN(new_n6026_));
  NOR3_X1    g05024(.A1(new_n6025_), .A2(new_n5039_), .A3(new_n6026_), .ZN(new_n6027_));
  NOR2_X1    g05025(.A1(new_n5046_), .A2(new_n5047_), .ZN(new_n6028_));
  NOR4_X1    g05026(.A1(new_n3645_), .A2(new_n3642_), .A3(new_n3646_), .A4(new_n3630_), .ZN(new_n6029_));
  OAI21_X1   g05027(.A1(new_n6028_), .A2(new_n6029_), .B(new_n5045_), .ZN(new_n6030_));
  INV_X1     g05028(.I(new_n6026_), .ZN(new_n6031_));
  AOI21_X1   g05029(.A1(new_n6030_), .A2(new_n5057_), .B(new_n6031_), .ZN(new_n6032_));
  NOR3_X1    g05030(.A1(new_n6027_), .A2(new_n6032_), .A3(new_n5056_), .ZN(new_n6033_));
  NAND3_X1   g05031(.A1(new_n6030_), .A2(new_n5057_), .A3(new_n6031_), .ZN(new_n6034_));
  OAI21_X1   g05032(.A1(new_n6025_), .A2(new_n5039_), .B(new_n6026_), .ZN(new_n6035_));
  AOI21_X1   g05033(.A1(new_n6035_), .A2(new_n6034_), .B(new_n5038_), .ZN(new_n6036_));
  OAI21_X1   g05034(.A1(new_n6033_), .A2(new_n6036_), .B(new_n6022_), .ZN(new_n6037_));
  AOI21_X1   g05035(.A1(new_n6017_), .A2(new_n5008_), .B(new_n6020_), .ZN(new_n6038_));
  NOR3_X1    g05036(.A1(new_n6006_), .A2(new_n6015_), .A3(new_n6005_), .ZN(new_n6039_));
  NOR2_X1    g05037(.A1(new_n6038_), .A2(new_n6039_), .ZN(new_n6040_));
  NAND3_X1   g05038(.A1(new_n6035_), .A2(new_n6034_), .A3(new_n5038_), .ZN(new_n6041_));
  OAI21_X1   g05039(.A1(new_n6027_), .A2(new_n6032_), .B(new_n5056_), .ZN(new_n6042_));
  NAND3_X1   g05040(.A1(new_n6040_), .A2(new_n6042_), .A3(new_n6041_), .ZN(new_n6043_));
  OAI21_X1   g05041(.A1(new_n5161_), .A2(new_n5052_), .B(new_n5163_), .ZN(new_n6044_));
  NAND3_X1   g05042(.A1(new_n6037_), .A2(new_n6043_), .A3(new_n6044_), .ZN(new_n6045_));
  AOI21_X1   g05043(.A1(new_n6042_), .A2(new_n6041_), .B(new_n6040_), .ZN(new_n6046_));
  NOR3_X1    g05044(.A1(new_n6033_), .A2(new_n6036_), .A3(new_n6022_), .ZN(new_n6047_));
  AOI21_X1   g05045(.A1(new_n5010_), .A2(new_n5162_), .B(new_n5060_), .ZN(new_n6048_));
  OAI21_X1   g05046(.A1(new_n6046_), .A2(new_n6047_), .B(new_n6048_), .ZN(new_n6049_));
  OAI21_X1   g05047(.A1(new_n5094_), .A2(new_n5131_), .B(new_n5154_), .ZN(new_n6050_));
  NOR2_X1    g05048(.A1(new_n5117_), .A2(new_n5125_), .ZN(new_n6051_));
  NOR2_X1    g05049(.A1(new_n5105_), .A2(new_n5120_), .ZN(new_n6052_));
  AOI21_X1   g05050(.A1(new_n5105_), .A2(new_n5120_), .B(new_n5119_), .ZN(new_n6053_));
  INV_X1     g05051(.I(new_n5102_), .ZN(new_n6054_));
  AOI21_X1   g05052(.A1(new_n5096_), .A2(new_n6054_), .B(new_n5101_), .ZN(new_n6055_));
  OAI21_X1   g05053(.A1(new_n6052_), .A2(new_n6053_), .B(new_n6055_), .ZN(new_n6056_));
  OR3_X2     g05054(.A1(new_n6053_), .A2(new_n6055_), .A3(new_n6052_), .Z(new_n6057_));
  NAND2_X1   g05055(.A1(new_n6057_), .A2(new_n6056_), .ZN(new_n6058_));
  OAI21_X1   g05056(.A1(new_n6051_), .A2(new_n5123_), .B(new_n6058_), .ZN(new_n6059_));
  NAND2_X1   g05057(.A1(new_n5128_), .A2(new_n5104_), .ZN(new_n6060_));
  INV_X1     g05058(.I(new_n6056_), .ZN(new_n6061_));
  NOR3_X1    g05059(.A1(new_n6053_), .A2(new_n6055_), .A3(new_n6052_), .ZN(new_n6062_));
  NOR2_X1    g05060(.A1(new_n6061_), .A2(new_n6062_), .ZN(new_n6063_));
  NAND3_X1   g05061(.A1(new_n6060_), .A2(new_n6063_), .A3(new_n5135_), .ZN(new_n6064_));
  NOR2_X1    g05062(.A1(new_n5085_), .A2(new_n5145_), .ZN(new_n6065_));
  AOI21_X1   g05063(.A1(new_n5085_), .A2(new_n5145_), .B(new_n5144_), .ZN(new_n6066_));
  INV_X1     g05064(.I(new_n5069_), .ZN(new_n6067_));
  AOI21_X1   g05065(.A1(new_n5141_), .A2(new_n5071_), .B(new_n6067_), .ZN(new_n6068_));
  OAI21_X1   g05066(.A1(new_n6066_), .A2(new_n6065_), .B(new_n6068_), .ZN(new_n6069_));
  NAND2_X1   g05067(.A1(new_n5074_), .A2(new_n5077_), .ZN(new_n6070_));
  OAI21_X1   g05068(.A1(new_n5074_), .A2(new_n5077_), .B(new_n5079_), .ZN(new_n6071_));
  OAI21_X1   g05069(.A1(new_n5066_), .A2(new_n5070_), .B(new_n5069_), .ZN(new_n6072_));
  NAND3_X1   g05070(.A1(new_n6071_), .A2(new_n6072_), .A3(new_n6070_), .ZN(new_n6073_));
  NAND2_X1   g05071(.A1(new_n6073_), .A2(new_n6069_), .ZN(new_n6074_));
  OAI21_X1   g05072(.A1(new_n5148_), .A2(new_n5083_), .B(new_n6074_), .ZN(new_n6075_));
  AOI21_X1   g05073(.A1(new_n6071_), .A2(new_n6070_), .B(new_n6072_), .ZN(new_n6076_));
  NOR3_X1    g05074(.A1(new_n6066_), .A2(new_n6068_), .A3(new_n6065_), .ZN(new_n6077_));
  NOR2_X1    g05075(.A1(new_n6076_), .A2(new_n6077_), .ZN(new_n6078_));
  NAND3_X1   g05076(.A1(new_n5143_), .A2(new_n6078_), .A3(new_n5090_), .ZN(new_n6079_));
  NAND4_X1   g05077(.A1(new_n6064_), .A2(new_n6059_), .A3(new_n6075_), .A4(new_n6079_), .ZN(new_n6080_));
  AOI21_X1   g05078(.A1(new_n6060_), .A2(new_n5135_), .B(new_n6063_), .ZN(new_n6081_));
  NOR3_X1    g05079(.A1(new_n6051_), .A2(new_n6058_), .A3(new_n5123_), .ZN(new_n6082_));
  AOI21_X1   g05080(.A1(new_n5143_), .A2(new_n5090_), .B(new_n6078_), .ZN(new_n6083_));
  NOR3_X1    g05081(.A1(new_n5148_), .A2(new_n5083_), .A3(new_n6074_), .ZN(new_n6084_));
  OAI22_X1   g05082(.A1(new_n6081_), .A2(new_n6082_), .B1(new_n6084_), .B2(new_n6083_), .ZN(new_n6085_));
  NAND3_X1   g05083(.A1(new_n6050_), .A2(new_n6085_), .A3(new_n6080_), .ZN(new_n6086_));
  AOI21_X1   g05084(.A1(new_n5152_), .A2(new_n5153_), .B(new_n5139_), .ZN(new_n6087_));
  NOR4_X1    g05085(.A1(new_n6081_), .A2(new_n6082_), .A3(new_n6084_), .A4(new_n6083_), .ZN(new_n6088_));
  AOI22_X1   g05086(.A1(new_n6064_), .A2(new_n6059_), .B1(new_n6075_), .B2(new_n6079_), .ZN(new_n6089_));
  OAI21_X1   g05087(.A1(new_n6088_), .A2(new_n6089_), .B(new_n6087_), .ZN(new_n6090_));
  NAND4_X1   g05088(.A1(new_n6090_), .A2(new_n6045_), .A3(new_n6049_), .A4(new_n6086_), .ZN(new_n6091_));
  NOR3_X1    g05089(.A1(new_n6046_), .A2(new_n6047_), .A3(new_n6048_), .ZN(new_n6092_));
  AOI21_X1   g05090(.A1(new_n6043_), .A2(new_n6037_), .B(new_n6044_), .ZN(new_n6093_));
  NOR3_X1    g05091(.A1(new_n6087_), .A2(new_n6088_), .A3(new_n6089_), .ZN(new_n6094_));
  AOI21_X1   g05092(.A1(new_n6080_), .A2(new_n6085_), .B(new_n6050_), .ZN(new_n6095_));
  OAI22_X1   g05093(.A1(new_n6094_), .A2(new_n6095_), .B1(new_n6093_), .B2(new_n6092_), .ZN(new_n6096_));
  NAND3_X1   g05094(.A1(new_n6096_), .A2(new_n6091_), .A3(new_n6003_), .ZN(new_n6097_));
  AOI21_X1   g05095(.A1(new_n5165_), .A2(new_n5166_), .B(new_n5159_), .ZN(new_n6098_));
  NOR4_X1    g05096(.A1(new_n6095_), .A2(new_n6093_), .A3(new_n6092_), .A4(new_n6094_), .ZN(new_n6099_));
  AOI22_X1   g05097(.A1(new_n6086_), .A2(new_n6090_), .B1(new_n6045_), .B2(new_n6049_), .ZN(new_n6100_));
  OAI21_X1   g05098(.A1(new_n6100_), .A2(new_n6099_), .B(new_n6098_), .ZN(new_n6101_));
  NAND4_X1   g05099(.A1(new_n6101_), .A2(new_n6097_), .A3(new_n6002_), .A4(new_n5997_), .ZN(new_n6102_));
  NOR3_X1    g05100(.A1(new_n5999_), .A2(new_n5998_), .A3(new_n6001_), .ZN(new_n6103_));
  AOI21_X1   g05101(.A1(new_n5993_), .A2(new_n5988_), .B(new_n5996_), .ZN(new_n6104_));
  NOR3_X1    g05102(.A1(new_n6100_), .A2(new_n6099_), .A3(new_n6098_), .ZN(new_n6105_));
  AOI21_X1   g05103(.A1(new_n6096_), .A2(new_n6091_), .B(new_n6003_), .ZN(new_n6106_));
  OAI22_X1   g05104(.A1(new_n6105_), .A2(new_n6106_), .B1(new_n6103_), .B2(new_n6104_), .ZN(new_n6107_));
  NAND3_X1   g05105(.A1(new_n6107_), .A2(new_n6102_), .A3(new_n5888_), .ZN(new_n6108_));
  AOI21_X1   g05106(.A1(new_n5176_), .A2(new_n5177_), .B(new_n5173_), .ZN(new_n6109_));
  NOR4_X1    g05107(.A1(new_n6105_), .A2(new_n6106_), .A3(new_n6103_), .A4(new_n6104_), .ZN(new_n6110_));
  AOI22_X1   g05108(.A1(new_n6101_), .A2(new_n6097_), .B1(new_n6002_), .B2(new_n5997_), .ZN(new_n6111_));
  OAI21_X1   g05109(.A1(new_n6110_), .A2(new_n6111_), .B(new_n6109_), .ZN(new_n6112_));
  NAND4_X1   g05110(.A1(new_n5887_), .A2(new_n5883_), .A3(new_n6112_), .A4(new_n6108_), .ZN(new_n6113_));
  NOR3_X1    g05111(.A1(new_n5884_), .A2(new_n5885_), .A3(new_n5886_), .ZN(new_n6114_));
  AOI21_X1   g05112(.A1(new_n5881_), .A2(new_n5876_), .B(new_n5882_), .ZN(new_n6115_));
  NOR3_X1    g05113(.A1(new_n6110_), .A2(new_n6111_), .A3(new_n6109_), .ZN(new_n6116_));
  AOI21_X1   g05114(.A1(new_n6107_), .A2(new_n6102_), .B(new_n5888_), .ZN(new_n6117_));
  OAI22_X1   g05115(.A1(new_n6114_), .A2(new_n6115_), .B1(new_n6116_), .B2(new_n6117_), .ZN(new_n6118_));
  NAND3_X1   g05116(.A1(new_n6118_), .A2(new_n6113_), .A3(new_n5661_), .ZN(new_n6119_));
  AOI21_X1   g05117(.A1(new_n5187_), .A2(new_n5188_), .B(new_n5183_), .ZN(new_n6120_));
  NOR4_X1    g05118(.A1(new_n6114_), .A2(new_n6115_), .A3(new_n6116_), .A4(new_n6117_), .ZN(new_n6121_));
  AOI22_X1   g05119(.A1(new_n5887_), .A2(new_n5883_), .B1(new_n6112_), .B2(new_n6108_), .ZN(new_n6122_));
  OAI21_X1   g05120(.A1(new_n6121_), .A2(new_n6122_), .B(new_n6120_), .ZN(new_n6123_));
  NAND4_X1   g05121(.A1(new_n5660_), .A2(new_n6123_), .A3(new_n5656_), .A4(new_n6119_), .ZN(new_n6124_));
  AOI22_X1   g05122(.A1(new_n5656_), .A2(new_n5660_), .B1(new_n6123_), .B2(new_n6119_), .ZN(new_n6125_));
  OAI21_X1   g05123(.A1(new_n6125_), .A2(new_n5194_), .B(new_n6124_), .ZN(new_n6126_));
  AOI21_X1   g05124(.A1(new_n5661_), .A2(new_n6118_), .B(new_n6121_), .ZN(new_n6127_));
  AOI21_X1   g05125(.A1(new_n5888_), .A2(new_n6107_), .B(new_n6110_), .ZN(new_n6128_));
  AOI21_X1   g05126(.A1(new_n6003_), .A2(new_n6096_), .B(new_n6099_), .ZN(new_n6129_));
  OAI21_X1   g05127(.A1(new_n6050_), .A2(new_n6088_), .B(new_n6085_), .ZN(new_n6130_));
  OAI21_X1   g05128(.A1(new_n6051_), .A2(new_n5123_), .B(new_n6057_), .ZN(new_n6131_));
  NAND2_X1   g05129(.A1(new_n6131_), .A2(new_n6056_), .ZN(new_n6132_));
  OAI21_X1   g05130(.A1(new_n5148_), .A2(new_n5083_), .B(new_n6073_), .ZN(new_n6133_));
  NAND3_X1   g05131(.A1(new_n6132_), .A2(new_n6069_), .A3(new_n6133_), .ZN(new_n6134_));
  NAND2_X1   g05132(.A1(new_n6133_), .A2(new_n6069_), .ZN(new_n6135_));
  NAND3_X1   g05133(.A1(new_n6135_), .A2(new_n6056_), .A3(new_n6131_), .ZN(new_n6136_));
  NAND2_X1   g05134(.A1(new_n6136_), .A2(new_n6134_), .ZN(new_n6137_));
  NAND2_X1   g05135(.A1(new_n6137_), .A2(new_n6130_), .ZN(new_n6138_));
  NAND2_X1   g05136(.A1(new_n6087_), .A2(new_n6080_), .ZN(new_n6139_));
  NAND4_X1   g05137(.A1(new_n6139_), .A2(new_n6085_), .A3(new_n6134_), .A4(new_n6136_), .ZN(new_n6140_));
  NOR2_X1    g05138(.A1(new_n6046_), .A2(new_n6044_), .ZN(new_n6141_));
  NOR2_X1    g05139(.A1(new_n6032_), .A2(new_n5038_), .ZN(new_n6142_));
  NOR2_X1    g05140(.A1(new_n6006_), .A2(new_n6005_), .ZN(new_n6143_));
  AOI21_X1   g05141(.A1(new_n6143_), .A2(new_n6019_), .B(new_n6010_), .ZN(new_n6144_));
  OAI21_X1   g05142(.A1(new_n6142_), .A2(new_n6027_), .B(new_n6144_), .ZN(new_n6145_));
  NAND2_X1   g05143(.A1(new_n6035_), .A2(new_n5056_), .ZN(new_n6146_));
  NAND2_X1   g05144(.A1(new_n6017_), .A2(new_n5008_), .ZN(new_n6147_));
  OAI21_X1   g05145(.A1(new_n6147_), .A2(new_n6014_), .B(new_n6018_), .ZN(new_n6148_));
  NAND3_X1   g05146(.A1(new_n6146_), .A2(new_n6148_), .A3(new_n6034_), .ZN(new_n6149_));
  NAND2_X1   g05147(.A1(new_n6145_), .A2(new_n6149_), .ZN(new_n6150_));
  OAI21_X1   g05148(.A1(new_n6141_), .A2(new_n6047_), .B(new_n6150_), .ZN(new_n6151_));
  NAND2_X1   g05149(.A1(new_n6037_), .A2(new_n6048_), .ZN(new_n6152_));
  AOI21_X1   g05150(.A1(new_n6034_), .A2(new_n6146_), .B(new_n6148_), .ZN(new_n6153_));
  NOR3_X1    g05151(.A1(new_n6144_), .A2(new_n6142_), .A3(new_n6027_), .ZN(new_n6154_));
  NOR2_X1    g05152(.A1(new_n6153_), .A2(new_n6154_), .ZN(new_n6155_));
  NAND3_X1   g05153(.A1(new_n6152_), .A2(new_n6155_), .A3(new_n6043_), .ZN(new_n6156_));
  AOI22_X1   g05154(.A1(new_n6138_), .A2(new_n6140_), .B1(new_n6151_), .B2(new_n6156_), .ZN(new_n6157_));
  AOI22_X1   g05155(.A1(new_n6139_), .A2(new_n6085_), .B1(new_n6134_), .B2(new_n6136_), .ZN(new_n6158_));
  NOR2_X1    g05156(.A1(new_n6137_), .A2(new_n6130_), .ZN(new_n6159_));
  AOI21_X1   g05157(.A1(new_n6152_), .A2(new_n6043_), .B(new_n6155_), .ZN(new_n6160_));
  NOR3_X1    g05158(.A1(new_n6141_), .A2(new_n6047_), .A3(new_n6150_), .ZN(new_n6161_));
  NOR4_X1    g05159(.A1(new_n6158_), .A2(new_n6159_), .A3(new_n6161_), .A4(new_n6160_), .ZN(new_n6162_));
  NOR3_X1    g05160(.A1(new_n6129_), .A2(new_n6157_), .A3(new_n6162_), .ZN(new_n6163_));
  OAI21_X1   g05161(.A1(new_n6100_), .A2(new_n6098_), .B(new_n6091_), .ZN(new_n6164_));
  OAI22_X1   g05162(.A1(new_n6158_), .A2(new_n6159_), .B1(new_n6161_), .B2(new_n6160_), .ZN(new_n6165_));
  NAND4_X1   g05163(.A1(new_n6138_), .A2(new_n6140_), .A3(new_n6151_), .A4(new_n6156_), .ZN(new_n6166_));
  AOI21_X1   g05164(.A1(new_n6165_), .A2(new_n6166_), .B(new_n6164_), .ZN(new_n6167_));
  AOI21_X1   g05165(.A1(new_n5993_), .A2(new_n5996_), .B(new_n5998_), .ZN(new_n6168_));
  NAND2_X1   g05166(.A1(new_n5927_), .A2(new_n5938_), .ZN(new_n6169_));
  NOR2_X1    g05167(.A1(new_n5921_), .A2(new_n5923_), .ZN(new_n6170_));
  NOR2_X1    g05168(.A1(new_n5891_), .A2(new_n4900_), .ZN(new_n6171_));
  AOI21_X1   g05169(.A1(new_n6171_), .A2(new_n5908_), .B(new_n5898_), .ZN(new_n6172_));
  OAI21_X1   g05170(.A1(new_n6170_), .A2(new_n5919_), .B(new_n6172_), .ZN(new_n6173_));
  NAND2_X1   g05171(.A1(new_n5925_), .A2(new_n5915_), .ZN(new_n6174_));
  NAND2_X1   g05172(.A1(new_n5906_), .A2(new_n4893_), .ZN(new_n6175_));
  OAI21_X1   g05173(.A1(new_n6175_), .A2(new_n5903_), .B(new_n5907_), .ZN(new_n6176_));
  NAND3_X1   g05174(.A1(new_n6174_), .A2(new_n6176_), .A3(new_n5924_), .ZN(new_n6177_));
  NAND2_X1   g05175(.A1(new_n6173_), .A2(new_n6177_), .ZN(new_n6178_));
  AOI21_X1   g05176(.A1(new_n6169_), .A2(new_n5933_), .B(new_n6178_), .ZN(new_n6179_));
  NOR2_X1    g05177(.A1(new_n5936_), .A2(new_n5934_), .ZN(new_n6180_));
  AOI21_X1   g05178(.A1(new_n5924_), .A2(new_n6174_), .B(new_n6176_), .ZN(new_n6181_));
  NOR3_X1    g05179(.A1(new_n6172_), .A2(new_n6170_), .A3(new_n5919_), .ZN(new_n6182_));
  NOR2_X1    g05180(.A1(new_n6181_), .A2(new_n6182_), .ZN(new_n6183_));
  NOR3_X1    g05181(.A1(new_n6180_), .A2(new_n6183_), .A3(new_n5937_), .ZN(new_n6184_));
  AOI21_X1   g05182(.A1(new_n5984_), .A2(new_n5977_), .B(new_n5986_), .ZN(new_n6185_));
  OAI21_X1   g05183(.A1(new_n5953_), .A2(new_n5955_), .B(new_n5946_), .ZN(new_n6186_));
  OAI21_X1   g05184(.A1(new_n5972_), .A2(new_n5974_), .B(new_n5965_), .ZN(new_n6187_));
  XOR2_X1    g05185(.A1(new_n6187_), .A2(new_n6186_), .Z(new_n6188_));
  NOR2_X1    g05186(.A1(new_n6185_), .A2(new_n6188_), .ZN(new_n6189_));
  OAI21_X1   g05187(.A1(new_n5940_), .A2(new_n5985_), .B(new_n5982_), .ZN(new_n6190_));
  AOI21_X1   g05188(.A1(new_n5958_), .A2(new_n5969_), .B(new_n5973_), .ZN(new_n6191_));
  XOR2_X1    g05189(.A1(new_n6191_), .A2(new_n6186_), .Z(new_n6192_));
  NOR2_X1    g05190(.A1(new_n6190_), .A2(new_n6192_), .ZN(new_n6193_));
  NOR4_X1    g05191(.A1(new_n6179_), .A2(new_n6184_), .A3(new_n6189_), .A4(new_n6193_), .ZN(new_n6194_));
  OAI21_X1   g05192(.A1(new_n6180_), .A2(new_n5937_), .B(new_n6183_), .ZN(new_n6195_));
  NAND3_X1   g05193(.A1(new_n6169_), .A2(new_n6178_), .A3(new_n5933_), .ZN(new_n6196_));
  NAND2_X1   g05194(.A1(new_n6190_), .A2(new_n6192_), .ZN(new_n6197_));
  NAND2_X1   g05195(.A1(new_n6185_), .A2(new_n6188_), .ZN(new_n6198_));
  AOI22_X1   g05196(.A1(new_n6195_), .A2(new_n6196_), .B1(new_n6197_), .B2(new_n6198_), .ZN(new_n6199_));
  NOR3_X1    g05197(.A1(new_n6168_), .A2(new_n6194_), .A3(new_n6199_), .ZN(new_n6200_));
  OAI21_X1   g05198(.A1(new_n5999_), .A2(new_n6001_), .B(new_n5988_), .ZN(new_n6201_));
  NAND4_X1   g05199(.A1(new_n6195_), .A2(new_n6196_), .A3(new_n6197_), .A4(new_n6198_), .ZN(new_n6202_));
  OAI22_X1   g05200(.A1(new_n6179_), .A2(new_n6184_), .B1(new_n6189_), .B2(new_n6193_), .ZN(new_n6203_));
  AOI21_X1   g05201(.A1(new_n6202_), .A2(new_n6203_), .B(new_n6201_), .ZN(new_n6204_));
  NOR4_X1    g05202(.A1(new_n6167_), .A2(new_n6163_), .A3(new_n6204_), .A4(new_n6200_), .ZN(new_n6205_));
  NAND3_X1   g05203(.A1(new_n6164_), .A2(new_n6165_), .A3(new_n6166_), .ZN(new_n6206_));
  OAI21_X1   g05204(.A1(new_n6157_), .A2(new_n6162_), .B(new_n6129_), .ZN(new_n6207_));
  NAND3_X1   g05205(.A1(new_n6201_), .A2(new_n6202_), .A3(new_n6203_), .ZN(new_n6208_));
  OAI21_X1   g05206(.A1(new_n6194_), .A2(new_n6199_), .B(new_n6168_), .ZN(new_n6209_));
  AOI22_X1   g05207(.A1(new_n6207_), .A2(new_n6206_), .B1(new_n6209_), .B2(new_n6208_), .ZN(new_n6210_));
  NOR3_X1    g05208(.A1(new_n6210_), .A2(new_n6128_), .A3(new_n6205_), .ZN(new_n6211_));
  OAI21_X1   g05209(.A1(new_n6109_), .A2(new_n6111_), .B(new_n6102_), .ZN(new_n6212_));
  NAND4_X1   g05210(.A1(new_n6207_), .A2(new_n6209_), .A3(new_n6206_), .A4(new_n6208_), .ZN(new_n6213_));
  OAI22_X1   g05211(.A1(new_n6167_), .A2(new_n6163_), .B1(new_n6204_), .B2(new_n6200_), .ZN(new_n6214_));
  AOI21_X1   g05212(.A1(new_n6213_), .A2(new_n6214_), .B(new_n6212_), .ZN(new_n6215_));
  AOI21_X1   g05213(.A1(new_n5881_), .A2(new_n5882_), .B(new_n5884_), .ZN(new_n6216_));
  AOI21_X1   g05214(.A1(new_n5771_), .A2(new_n5870_), .B(new_n5873_), .ZN(new_n6217_));
  OAI21_X1   g05215(.A1(new_n5821_), .A2(new_n5862_), .B(new_n5859_), .ZN(new_n6218_));
  OAI21_X1   g05216(.A1(new_n5822_), .A2(new_n4532_), .B(new_n5830_), .ZN(new_n6219_));
  NAND2_X1   g05217(.A1(new_n6219_), .A2(new_n5827_), .ZN(new_n6220_));
  OAI21_X1   g05218(.A1(new_n4493_), .A2(new_n4557_), .B(new_n5847_), .ZN(new_n6221_));
  NAND3_X1   g05219(.A1(new_n6220_), .A2(new_n5842_), .A3(new_n6221_), .ZN(new_n6222_));
  NAND2_X1   g05220(.A1(new_n6221_), .A2(new_n5842_), .ZN(new_n6223_));
  NAND3_X1   g05221(.A1(new_n6223_), .A2(new_n5827_), .A3(new_n6219_), .ZN(new_n6224_));
  NAND2_X1   g05222(.A1(new_n6222_), .A2(new_n6224_), .ZN(new_n6225_));
  NAND2_X1   g05223(.A1(new_n6218_), .A2(new_n6225_), .ZN(new_n6226_));
  NAND2_X1   g05224(.A1(new_n4562_), .A2(new_n4561_), .ZN(new_n6227_));
  NAND3_X1   g05225(.A1(new_n6227_), .A2(new_n5854_), .A3(new_n4563_), .ZN(new_n6228_));
  NAND4_X1   g05226(.A1(new_n6228_), .A2(new_n5859_), .A3(new_n6222_), .A4(new_n6224_), .ZN(new_n6229_));
  OAI21_X1   g05227(.A1(new_n5816_), .A2(new_n5814_), .B(new_n5811_), .ZN(new_n6230_));
  NOR2_X1    g05228(.A1(new_n5800_), .A2(new_n4446_), .ZN(new_n6231_));
  NOR2_X1    g05229(.A1(new_n5774_), .A2(new_n5773_), .ZN(new_n6232_));
  AOI21_X1   g05230(.A1(new_n6232_), .A2(new_n5787_), .B(new_n5778_), .ZN(new_n6233_));
  OAI21_X1   g05231(.A1(new_n6231_), .A2(new_n5795_), .B(new_n6233_), .ZN(new_n6234_));
  NAND2_X1   g05232(.A1(new_n5803_), .A2(new_n4464_), .ZN(new_n6235_));
  NAND2_X1   g05233(.A1(new_n5785_), .A2(new_n4415_), .ZN(new_n6236_));
  OAI21_X1   g05234(.A1(new_n6236_), .A2(new_n5782_), .B(new_n5786_), .ZN(new_n6237_));
  NAND3_X1   g05235(.A1(new_n6235_), .A2(new_n6237_), .A3(new_n5802_), .ZN(new_n6238_));
  NAND2_X1   g05236(.A1(new_n6234_), .A2(new_n6238_), .ZN(new_n6239_));
  NAND2_X1   g05237(.A1(new_n6230_), .A2(new_n6239_), .ZN(new_n6240_));
  NAND2_X1   g05238(.A1(new_n5805_), .A2(new_n5819_), .ZN(new_n6241_));
  AOI21_X1   g05239(.A1(new_n6235_), .A2(new_n5802_), .B(new_n6237_), .ZN(new_n6242_));
  NOR3_X1    g05240(.A1(new_n6233_), .A2(new_n6231_), .A3(new_n5795_), .ZN(new_n6243_));
  NOR2_X1    g05241(.A1(new_n6242_), .A2(new_n6243_), .ZN(new_n6244_));
  NAND3_X1   g05242(.A1(new_n6241_), .A2(new_n6244_), .A3(new_n5811_), .ZN(new_n6245_));
  AOI22_X1   g05243(.A1(new_n6240_), .A2(new_n6245_), .B1(new_n6226_), .B2(new_n6229_), .ZN(new_n6246_));
  AOI22_X1   g05244(.A1(new_n6228_), .A2(new_n5859_), .B1(new_n6222_), .B2(new_n6224_), .ZN(new_n6247_));
  NOR2_X1    g05245(.A1(new_n6218_), .A2(new_n6225_), .ZN(new_n6248_));
  AOI21_X1   g05246(.A1(new_n6241_), .A2(new_n5811_), .B(new_n6244_), .ZN(new_n6249_));
  NOR2_X1    g05247(.A1(new_n6230_), .A2(new_n6239_), .ZN(new_n6250_));
  NOR4_X1    g05248(.A1(new_n6250_), .A2(new_n6249_), .A3(new_n6248_), .A4(new_n6247_), .ZN(new_n6251_));
  NOR3_X1    g05249(.A1(new_n6217_), .A2(new_n6246_), .A3(new_n6251_), .ZN(new_n6252_));
  OAI21_X1   g05250(.A1(new_n5874_), .A2(new_n5872_), .B(new_n5865_), .ZN(new_n6253_));
  OAI22_X1   g05251(.A1(new_n6250_), .A2(new_n6249_), .B1(new_n6248_), .B2(new_n6247_), .ZN(new_n6254_));
  NAND4_X1   g05252(.A1(new_n6240_), .A2(new_n6226_), .A3(new_n6245_), .A4(new_n6229_), .ZN(new_n6255_));
  AOI21_X1   g05253(.A1(new_n6254_), .A2(new_n6255_), .B(new_n6253_), .ZN(new_n6256_));
  AOI21_X1   g05254(.A1(new_n5761_), .A2(new_n5762_), .B(new_n5764_), .ZN(new_n6257_));
  AOI21_X1   g05255(.A1(new_n5694_), .A2(new_n5705_), .B(new_n5704_), .ZN(new_n6258_));
  NOR2_X1    g05256(.A1(new_n5688_), .A2(new_n5690_), .ZN(new_n6259_));
  NOR2_X1    g05257(.A1(new_n5662_), .A2(new_n4682_), .ZN(new_n6260_));
  AOI21_X1   g05258(.A1(new_n6260_), .A2(new_n5677_), .B(new_n5667_), .ZN(new_n6261_));
  OAI21_X1   g05259(.A1(new_n6259_), .A2(new_n5686_), .B(new_n6261_), .ZN(new_n6262_));
  NAND2_X1   g05260(.A1(new_n5692_), .A2(new_n5684_), .ZN(new_n6263_));
  NAND2_X1   g05261(.A1(new_n5675_), .A2(new_n4692_), .ZN(new_n6264_));
  OAI21_X1   g05262(.A1(new_n6264_), .A2(new_n5672_), .B(new_n5676_), .ZN(new_n6265_));
  NAND3_X1   g05263(.A1(new_n6265_), .A2(new_n6263_), .A3(new_n5691_), .ZN(new_n6266_));
  NAND2_X1   g05264(.A1(new_n6262_), .A2(new_n6266_), .ZN(new_n6267_));
  NOR2_X1    g05265(.A1(new_n6258_), .A2(new_n6267_), .ZN(new_n6268_));
  NOR2_X1    g05266(.A1(new_n5703_), .A2(new_n5701_), .ZN(new_n6269_));
  AOI21_X1   g05267(.A1(new_n5691_), .A2(new_n6263_), .B(new_n6265_), .ZN(new_n6270_));
  NOR3_X1    g05268(.A1(new_n6261_), .A2(new_n6259_), .A3(new_n5686_), .ZN(new_n6271_));
  NOR2_X1    g05269(.A1(new_n6270_), .A2(new_n6271_), .ZN(new_n6272_));
  NOR3_X1    g05270(.A1(new_n6269_), .A2(new_n6272_), .A3(new_n5704_), .ZN(new_n6273_));
  NAND2_X1   g05271(.A1(new_n5744_), .A2(new_n5752_), .ZN(new_n6274_));
  AOI21_X1   g05272(.A1(new_n4602_), .A2(new_n4587_), .B(new_n4601_), .ZN(new_n6275_));
  OAI21_X1   g05273(.A1(new_n6275_), .A2(new_n5737_), .B(new_n5734_), .ZN(new_n6276_));
  NAND2_X1   g05274(.A1(new_n6276_), .A2(new_n5741_), .ZN(new_n6277_));
  OAI21_X1   g05275(.A1(new_n4630_), .A2(new_n4635_), .B(new_n4639_), .ZN(new_n6278_));
  OAI21_X1   g05276(.A1(new_n6278_), .A2(new_n5720_), .B(new_n5726_), .ZN(new_n6279_));
  INV_X1     g05277(.I(new_n6279_), .ZN(new_n6280_));
  NAND2_X1   g05278(.A1(new_n6277_), .A2(new_n6280_), .ZN(new_n6281_));
  NAND3_X1   g05279(.A1(new_n6279_), .A2(new_n6276_), .A3(new_n5741_), .ZN(new_n6282_));
  NAND2_X1   g05280(.A1(new_n6281_), .A2(new_n6282_), .ZN(new_n6283_));
  AOI21_X1   g05281(.A1(new_n6274_), .A2(new_n5750_), .B(new_n6283_), .ZN(new_n6284_));
  NOR2_X1    g05282(.A1(new_n5753_), .A2(new_n5707_), .ZN(new_n6285_));
  AOI21_X1   g05283(.A1(new_n5741_), .A2(new_n6276_), .B(new_n6279_), .ZN(new_n6286_));
  INV_X1     g05284(.I(new_n6282_), .ZN(new_n6287_));
  NOR2_X1    g05285(.A1(new_n6287_), .A2(new_n6286_), .ZN(new_n6288_));
  NOR3_X1    g05286(.A1(new_n6285_), .A2(new_n6288_), .A3(new_n5754_), .ZN(new_n6289_));
  NOR4_X1    g05287(.A1(new_n6268_), .A2(new_n6273_), .A3(new_n6289_), .A4(new_n6284_), .ZN(new_n6290_));
  OAI21_X1   g05288(.A1(new_n5703_), .A2(new_n5701_), .B(new_n5700_), .ZN(new_n6291_));
  NAND2_X1   g05289(.A1(new_n6291_), .A2(new_n6272_), .ZN(new_n6292_));
  NAND2_X1   g05290(.A1(new_n5694_), .A2(new_n5705_), .ZN(new_n6293_));
  NAND3_X1   g05291(.A1(new_n6293_), .A2(new_n6267_), .A3(new_n5700_), .ZN(new_n6294_));
  OAI21_X1   g05292(.A1(new_n6285_), .A2(new_n5754_), .B(new_n6288_), .ZN(new_n6295_));
  NAND3_X1   g05293(.A1(new_n6274_), .A2(new_n6283_), .A3(new_n5750_), .ZN(new_n6296_));
  AOI22_X1   g05294(.A1(new_n6292_), .A2(new_n6294_), .B1(new_n6295_), .B2(new_n6296_), .ZN(new_n6297_));
  NOR3_X1    g05295(.A1(new_n6257_), .A2(new_n6290_), .A3(new_n6297_), .ZN(new_n6298_));
  OAI21_X1   g05296(.A1(new_n5765_), .A2(new_n5766_), .B(new_n5756_), .ZN(new_n6299_));
  NAND4_X1   g05297(.A1(new_n6292_), .A2(new_n6294_), .A3(new_n6295_), .A4(new_n6296_), .ZN(new_n6300_));
  OAI22_X1   g05298(.A1(new_n6268_), .A2(new_n6273_), .B1(new_n6289_), .B2(new_n6284_), .ZN(new_n6301_));
  AOI21_X1   g05299(.A1(new_n6300_), .A2(new_n6301_), .B(new_n6299_), .ZN(new_n6302_));
  NOR4_X1    g05300(.A1(new_n6298_), .A2(new_n6302_), .A3(new_n6256_), .A4(new_n6252_), .ZN(new_n6303_));
  NAND3_X1   g05301(.A1(new_n6253_), .A2(new_n6254_), .A3(new_n6255_), .ZN(new_n6304_));
  OAI21_X1   g05302(.A1(new_n6246_), .A2(new_n6251_), .B(new_n6217_), .ZN(new_n6305_));
  NAND3_X1   g05303(.A1(new_n6299_), .A2(new_n6300_), .A3(new_n6301_), .ZN(new_n6306_));
  OAI21_X1   g05304(.A1(new_n6290_), .A2(new_n6297_), .B(new_n6257_), .ZN(new_n6307_));
  AOI22_X1   g05305(.A1(new_n6307_), .A2(new_n6306_), .B1(new_n6305_), .B2(new_n6304_), .ZN(new_n6308_));
  NOR3_X1    g05306(.A1(new_n6216_), .A2(new_n6308_), .A3(new_n6303_), .ZN(new_n6309_));
  OAI21_X1   g05307(.A1(new_n5885_), .A2(new_n5886_), .B(new_n5876_), .ZN(new_n6310_));
  NAND4_X1   g05308(.A1(new_n6307_), .A2(new_n6305_), .A3(new_n6306_), .A4(new_n6304_), .ZN(new_n6311_));
  OAI22_X1   g05309(.A1(new_n6302_), .A2(new_n6298_), .B1(new_n6256_), .B2(new_n6252_), .ZN(new_n6312_));
  AOI21_X1   g05310(.A1(new_n6311_), .A2(new_n6312_), .B(new_n6310_), .ZN(new_n6313_));
  NOR4_X1    g05311(.A1(new_n6309_), .A2(new_n6313_), .A3(new_n6211_), .A4(new_n6215_), .ZN(new_n6314_));
  NAND3_X1   g05312(.A1(new_n6213_), .A2(new_n6214_), .A3(new_n6212_), .ZN(new_n6315_));
  OAI21_X1   g05313(.A1(new_n6210_), .A2(new_n6205_), .B(new_n6128_), .ZN(new_n6316_));
  NAND3_X1   g05314(.A1(new_n6310_), .A2(new_n6312_), .A3(new_n6311_), .ZN(new_n6317_));
  OAI21_X1   g05315(.A1(new_n6303_), .A2(new_n6308_), .B(new_n6216_), .ZN(new_n6318_));
  AOI22_X1   g05316(.A1(new_n6318_), .A2(new_n6317_), .B1(new_n6316_), .B2(new_n6315_), .ZN(new_n6319_));
  NOR3_X1    g05317(.A1(new_n6314_), .A2(new_n6319_), .A3(new_n6127_), .ZN(new_n6320_));
  OAI21_X1   g05318(.A1(new_n6120_), .A2(new_n6122_), .B(new_n6113_), .ZN(new_n6321_));
  NAND4_X1   g05319(.A1(new_n6318_), .A2(new_n6317_), .A3(new_n6316_), .A4(new_n6315_), .ZN(new_n6322_));
  OAI22_X1   g05320(.A1(new_n6309_), .A2(new_n6313_), .B1(new_n6211_), .B2(new_n6215_), .ZN(new_n6323_));
  AOI21_X1   g05321(.A1(new_n6323_), .A2(new_n6322_), .B(new_n6321_), .ZN(new_n6324_));
  AOI21_X1   g05322(.A1(new_n5654_), .A2(new_n5655_), .B(new_n5657_), .ZN(new_n6325_));
  AOI21_X1   g05323(.A1(new_n5429_), .A2(new_n5643_), .B(new_n5646_), .ZN(new_n6326_));
  AOI21_X1   g05324(.A1(new_n5538_), .A2(new_n5632_), .B(new_n5635_), .ZN(new_n6327_));
  OAI21_X1   g05325(.A1(new_n5582_), .A2(new_n5624_), .B(new_n5621_), .ZN(new_n6328_));
  OAI21_X1   g05326(.A1(new_n5583_), .A2(new_n2026_), .B(new_n5593_), .ZN(new_n6329_));
  NAND2_X1   g05327(.A1(new_n6329_), .A2(new_n5588_), .ZN(new_n6330_));
  OAI21_X1   g05328(.A1(new_n2034_), .A2(new_n1980_), .B(new_n5609_), .ZN(new_n6331_));
  NAND3_X1   g05329(.A1(new_n6330_), .A2(new_n5605_), .A3(new_n6331_), .ZN(new_n6332_));
  NAND2_X1   g05330(.A1(new_n6331_), .A2(new_n5605_), .ZN(new_n6333_));
  NAND3_X1   g05331(.A1(new_n6333_), .A2(new_n5588_), .A3(new_n6329_), .ZN(new_n6334_));
  NAND2_X1   g05332(.A1(new_n6332_), .A2(new_n6334_), .ZN(new_n6335_));
  NAND2_X1   g05333(.A1(new_n6328_), .A2(new_n6335_), .ZN(new_n6336_));
  NAND2_X1   g05334(.A1(new_n2020_), .A2(new_n1984_), .ZN(new_n6337_));
  NAND3_X1   g05335(.A1(new_n6337_), .A2(new_n5616_), .A3(new_n2030_), .ZN(new_n6338_));
  NAND4_X1   g05336(.A1(new_n6338_), .A2(new_n5621_), .A3(new_n6332_), .A4(new_n6334_), .ZN(new_n6339_));
  NOR2_X1    g05337(.A1(new_n5578_), .A2(new_n5576_), .ZN(new_n6340_));
  NOR2_X1    g05338(.A1(new_n5564_), .A2(new_n1932_), .ZN(new_n6341_));
  NOR2_X1    g05339(.A1(new_n5539_), .A2(new_n1884_), .ZN(new_n6342_));
  AOI21_X1   g05340(.A1(new_n6342_), .A2(new_n5552_), .B(new_n5543_), .ZN(new_n6343_));
  OAI21_X1   g05341(.A1(new_n6341_), .A2(new_n5560_), .B(new_n6343_), .ZN(new_n6344_));
  NAND2_X1   g05342(.A1(new_n5567_), .A2(new_n1918_), .ZN(new_n6345_));
  NAND2_X1   g05343(.A1(new_n5550_), .A2(new_n1943_), .ZN(new_n6346_));
  OAI21_X1   g05344(.A1(new_n6346_), .A2(new_n5547_), .B(new_n5551_), .ZN(new_n6347_));
  NAND3_X1   g05345(.A1(new_n6345_), .A2(new_n6347_), .A3(new_n5566_), .ZN(new_n6348_));
  NAND2_X1   g05346(.A1(new_n6344_), .A2(new_n6348_), .ZN(new_n6349_));
  OAI21_X1   g05347(.A1(new_n6340_), .A2(new_n5579_), .B(new_n6349_), .ZN(new_n6350_));
  NAND2_X1   g05348(.A1(new_n5569_), .A2(new_n5580_), .ZN(new_n6351_));
  AOI21_X1   g05349(.A1(new_n5566_), .A2(new_n6345_), .B(new_n6347_), .ZN(new_n6352_));
  NOR3_X1    g05350(.A1(new_n6343_), .A2(new_n6341_), .A3(new_n5560_), .ZN(new_n6353_));
  NOR2_X1    g05351(.A1(new_n6352_), .A2(new_n6353_), .ZN(new_n6354_));
  NAND3_X1   g05352(.A1(new_n6351_), .A2(new_n6354_), .A3(new_n5575_), .ZN(new_n6355_));
  AOI22_X1   g05353(.A1(new_n6336_), .A2(new_n6339_), .B1(new_n6350_), .B2(new_n6355_), .ZN(new_n6356_));
  AOI22_X1   g05354(.A1(new_n6338_), .A2(new_n5621_), .B1(new_n6332_), .B2(new_n6334_), .ZN(new_n6357_));
  NOR2_X1    g05355(.A1(new_n6328_), .A2(new_n6335_), .ZN(new_n6358_));
  AOI21_X1   g05356(.A1(new_n6351_), .A2(new_n5575_), .B(new_n6354_), .ZN(new_n6359_));
  NOR3_X1    g05357(.A1(new_n6340_), .A2(new_n5579_), .A3(new_n6349_), .ZN(new_n6360_));
  NOR4_X1    g05358(.A1(new_n6358_), .A2(new_n6360_), .A3(new_n6359_), .A4(new_n6357_), .ZN(new_n6361_));
  NOR3_X1    g05359(.A1(new_n6327_), .A2(new_n6356_), .A3(new_n6361_), .ZN(new_n6362_));
  OAI21_X1   g05360(.A1(new_n5636_), .A2(new_n5634_), .B(new_n5627_), .ZN(new_n6363_));
  OAI22_X1   g05361(.A1(new_n6359_), .A2(new_n6360_), .B1(new_n6358_), .B2(new_n6357_), .ZN(new_n6364_));
  NAND4_X1   g05362(.A1(new_n6336_), .A2(new_n6350_), .A3(new_n6355_), .A4(new_n6339_), .ZN(new_n6365_));
  AOI21_X1   g05363(.A1(new_n6364_), .A2(new_n6365_), .B(new_n6363_), .ZN(new_n6366_));
  AOI21_X1   g05364(.A1(new_n5531_), .A2(new_n5532_), .B(new_n5534_), .ZN(new_n6367_));
  NAND2_X1   g05365(.A1(new_n5468_), .A2(new_n5479_), .ZN(new_n6368_));
  NOR2_X1    g05366(.A1(new_n5462_), .A2(new_n5464_), .ZN(new_n6369_));
  NOR2_X1    g05367(.A1(new_n5432_), .A2(new_n1436_), .ZN(new_n6370_));
  AOI21_X1   g05368(.A1(new_n6370_), .A2(new_n5449_), .B(new_n5439_), .ZN(new_n6371_));
  OAI21_X1   g05369(.A1(new_n6369_), .A2(new_n5460_), .B(new_n6371_), .ZN(new_n6372_));
  NAND2_X1   g05370(.A1(new_n5466_), .A2(new_n5456_), .ZN(new_n6373_));
  NAND2_X1   g05371(.A1(new_n5447_), .A2(new_n1444_), .ZN(new_n6374_));
  OAI21_X1   g05372(.A1(new_n6374_), .A2(new_n5444_), .B(new_n5448_), .ZN(new_n6375_));
  NAND3_X1   g05373(.A1(new_n6373_), .A2(new_n6375_), .A3(new_n5465_), .ZN(new_n6376_));
  NAND2_X1   g05374(.A1(new_n6372_), .A2(new_n6376_), .ZN(new_n6377_));
  AOI21_X1   g05375(.A1(new_n6368_), .A2(new_n5474_), .B(new_n6377_), .ZN(new_n6378_));
  NOR2_X1    g05376(.A1(new_n5477_), .A2(new_n5475_), .ZN(new_n6379_));
  AOI21_X1   g05377(.A1(new_n5465_), .A2(new_n6373_), .B(new_n6375_), .ZN(new_n6380_));
  NOR3_X1    g05378(.A1(new_n6371_), .A2(new_n6369_), .A3(new_n5460_), .ZN(new_n6381_));
  NOR2_X1    g05379(.A1(new_n6380_), .A2(new_n6381_), .ZN(new_n6382_));
  NOR3_X1    g05380(.A1(new_n6379_), .A2(new_n6382_), .A3(new_n5478_), .ZN(new_n6383_));
  AOI21_X1   g05381(.A1(new_n5522_), .A2(new_n5515_), .B(new_n5524_), .ZN(new_n6384_));
  OAI21_X1   g05382(.A1(new_n5494_), .A2(new_n5496_), .B(new_n5487_), .ZN(new_n6385_));
  OAI21_X1   g05383(.A1(new_n5510_), .A2(new_n5512_), .B(new_n5503_), .ZN(new_n6386_));
  XOR2_X1    g05384(.A1(new_n6386_), .A2(new_n6385_), .Z(new_n6387_));
  NOR2_X1    g05385(.A1(new_n6384_), .A2(new_n6387_), .ZN(new_n6388_));
  OAI21_X1   g05386(.A1(new_n5481_), .A2(new_n5523_), .B(new_n5520_), .ZN(new_n6389_));
  XNOR2_X1   g05387(.A1(new_n6386_), .A2(new_n6385_), .ZN(new_n6390_));
  NOR2_X1    g05388(.A1(new_n6389_), .A2(new_n6390_), .ZN(new_n6391_));
  NOR4_X1    g05389(.A1(new_n6378_), .A2(new_n6383_), .A3(new_n6388_), .A4(new_n6391_), .ZN(new_n6392_));
  OAI21_X1   g05390(.A1(new_n6379_), .A2(new_n5478_), .B(new_n6382_), .ZN(new_n6393_));
  NAND3_X1   g05391(.A1(new_n6368_), .A2(new_n6377_), .A3(new_n5474_), .ZN(new_n6394_));
  NAND2_X1   g05392(.A1(new_n6389_), .A2(new_n6390_), .ZN(new_n6395_));
  NAND2_X1   g05393(.A1(new_n6384_), .A2(new_n6387_), .ZN(new_n6396_));
  AOI22_X1   g05394(.A1(new_n6393_), .A2(new_n6394_), .B1(new_n6395_), .B2(new_n6396_), .ZN(new_n6397_));
  NOR3_X1    g05395(.A1(new_n6367_), .A2(new_n6392_), .A3(new_n6397_), .ZN(new_n6398_));
  OAI21_X1   g05396(.A1(new_n5535_), .A2(new_n5536_), .B(new_n5526_), .ZN(new_n6399_));
  NAND4_X1   g05397(.A1(new_n6393_), .A2(new_n6394_), .A3(new_n6395_), .A4(new_n6396_), .ZN(new_n6400_));
  OAI22_X1   g05398(.A1(new_n6378_), .A2(new_n6383_), .B1(new_n6388_), .B2(new_n6391_), .ZN(new_n6401_));
  AOI21_X1   g05399(.A1(new_n6400_), .A2(new_n6401_), .B(new_n6399_), .ZN(new_n6402_));
  NOR4_X1    g05400(.A1(new_n6366_), .A2(new_n6362_), .A3(new_n6402_), .A4(new_n6398_), .ZN(new_n6403_));
  NAND3_X1   g05401(.A1(new_n6363_), .A2(new_n6364_), .A3(new_n6365_), .ZN(new_n6404_));
  OAI21_X1   g05402(.A1(new_n6356_), .A2(new_n6361_), .B(new_n6327_), .ZN(new_n6405_));
  NAND3_X1   g05403(.A1(new_n6399_), .A2(new_n6400_), .A3(new_n6401_), .ZN(new_n6406_));
  OAI21_X1   g05404(.A1(new_n6392_), .A2(new_n6397_), .B(new_n6367_), .ZN(new_n6407_));
  AOI22_X1   g05405(.A1(new_n6405_), .A2(new_n6404_), .B1(new_n6407_), .B2(new_n6406_), .ZN(new_n6408_));
  NOR3_X1    g05406(.A1(new_n6408_), .A2(new_n6326_), .A3(new_n6403_), .ZN(new_n6409_));
  OAI21_X1   g05407(.A1(new_n5645_), .A2(new_n5647_), .B(new_n5638_), .ZN(new_n6410_));
  NAND4_X1   g05408(.A1(new_n6405_), .A2(new_n6407_), .A3(new_n6404_), .A4(new_n6406_), .ZN(new_n6411_));
  OAI22_X1   g05409(.A1(new_n6366_), .A2(new_n6362_), .B1(new_n6402_), .B2(new_n6398_), .ZN(new_n6412_));
  AOI21_X1   g05410(.A1(new_n6411_), .A2(new_n6412_), .B(new_n6410_), .ZN(new_n6413_));
  AOI21_X1   g05411(.A1(new_n5422_), .A2(new_n5423_), .B(new_n5425_), .ZN(new_n6414_));
  AOI21_X1   g05412(.A1(new_n5302_), .A2(new_n5409_), .B(new_n5414_), .ZN(new_n6415_));
  NOR2_X1    g05413(.A1(new_n5349_), .A2(new_n5347_), .ZN(new_n6416_));
  NAND2_X1   g05414(.A1(new_n5338_), .A2(new_n5325_), .ZN(new_n6417_));
  NAND2_X1   g05415(.A1(new_n5316_), .A2(new_n2732_), .ZN(new_n6418_));
  OAI21_X1   g05416(.A1(new_n6418_), .A2(new_n5313_), .B(new_n5317_), .ZN(new_n6419_));
  AOI21_X1   g05417(.A1(new_n6417_), .A2(new_n5337_), .B(new_n6419_), .ZN(new_n6420_));
  NOR2_X1    g05418(.A1(new_n5334_), .A2(new_n5336_), .ZN(new_n6421_));
  AOI21_X1   g05419(.A1(new_n2731_), .A2(new_n2711_), .B(new_n2726_), .ZN(new_n6422_));
  AOI21_X1   g05420(.A1(new_n6422_), .A2(new_n5318_), .B(new_n5309_), .ZN(new_n6423_));
  NOR3_X1    g05421(.A1(new_n6421_), .A2(new_n6423_), .A3(new_n5332_), .ZN(new_n6424_));
  NOR2_X1    g05422(.A1(new_n6420_), .A2(new_n6424_), .ZN(new_n6425_));
  OAI21_X1   g05423(.A1(new_n6416_), .A2(new_n5350_), .B(new_n6425_), .ZN(new_n6426_));
  NAND2_X1   g05424(.A1(new_n5340_), .A2(new_n5351_), .ZN(new_n6427_));
  OAI21_X1   g05425(.A1(new_n6421_), .A2(new_n5332_), .B(new_n6423_), .ZN(new_n6428_));
  NAND3_X1   g05426(.A1(new_n6419_), .A2(new_n6417_), .A3(new_n5337_), .ZN(new_n6429_));
  NAND2_X1   g05427(.A1(new_n6429_), .A2(new_n6428_), .ZN(new_n6430_));
  NAND3_X1   g05428(.A1(new_n6427_), .A2(new_n6430_), .A3(new_n5346_), .ZN(new_n6431_));
  NOR2_X1    g05429(.A1(new_n5401_), .A2(new_n5353_), .ZN(new_n6432_));
  NAND2_X1   g05430(.A1(new_n5389_), .A2(new_n5381_), .ZN(new_n6433_));
  NAND2_X1   g05431(.A1(new_n5372_), .A2(new_n2853_), .ZN(new_n6434_));
  OAI21_X1   g05432(.A1(new_n6434_), .A2(new_n5367_), .B(new_n5373_), .ZN(new_n6435_));
  AOI21_X1   g05433(.A1(new_n5388_), .A2(new_n6433_), .B(new_n6435_), .ZN(new_n6436_));
  NOR2_X1    g05434(.A1(new_n5385_), .A2(new_n5387_), .ZN(new_n6437_));
  AOI21_X1   g05435(.A1(new_n5392_), .A2(new_n5374_), .B(new_n5361_), .ZN(new_n6438_));
  NOR3_X1    g05436(.A1(new_n6437_), .A2(new_n5383_), .A3(new_n6438_), .ZN(new_n6439_));
  NOR2_X1    g05437(.A1(new_n6436_), .A2(new_n6439_), .ZN(new_n6440_));
  OAI21_X1   g05438(.A1(new_n6432_), .A2(new_n5402_), .B(new_n6440_), .ZN(new_n6441_));
  NAND2_X1   g05439(.A1(new_n5391_), .A2(new_n5400_), .ZN(new_n6442_));
  OAI21_X1   g05440(.A1(new_n6437_), .A2(new_n5383_), .B(new_n6438_), .ZN(new_n6443_));
  NAND3_X1   g05441(.A1(new_n6433_), .A2(new_n6435_), .A3(new_n5388_), .ZN(new_n6444_));
  NAND2_X1   g05442(.A1(new_n6444_), .A2(new_n6443_), .ZN(new_n6445_));
  NAND3_X1   g05443(.A1(new_n6442_), .A2(new_n5398_), .A3(new_n6445_), .ZN(new_n6446_));
  NAND4_X1   g05444(.A1(new_n6426_), .A2(new_n6441_), .A3(new_n6431_), .A4(new_n6446_), .ZN(new_n6447_));
  AOI21_X1   g05445(.A1(new_n6427_), .A2(new_n5346_), .B(new_n6430_), .ZN(new_n6448_));
  NOR3_X1    g05446(.A1(new_n6416_), .A2(new_n5350_), .A3(new_n6425_), .ZN(new_n6449_));
  AOI21_X1   g05447(.A1(new_n6442_), .A2(new_n5398_), .B(new_n6445_), .ZN(new_n6450_));
  NOR3_X1    g05448(.A1(new_n6432_), .A2(new_n5402_), .A3(new_n6440_), .ZN(new_n6451_));
  OAI22_X1   g05449(.A1(new_n6449_), .A2(new_n6448_), .B1(new_n6451_), .B2(new_n6450_), .ZN(new_n6452_));
  NAND2_X1   g05450(.A1(new_n6452_), .A2(new_n6447_), .ZN(new_n6453_));
  NOR2_X1    g05451(.A1(new_n6453_), .A2(new_n6415_), .ZN(new_n6454_));
  OAI21_X1   g05452(.A1(new_n5413_), .A2(new_n5415_), .B(new_n5404_), .ZN(new_n6455_));
  AOI21_X1   g05453(.A1(new_n6447_), .A2(new_n6452_), .B(new_n6455_), .ZN(new_n6456_));
  AOI21_X1   g05454(.A1(new_n5295_), .A2(new_n5296_), .B(new_n5298_), .ZN(new_n6457_));
  NAND2_X1   g05455(.A1(new_n5238_), .A2(new_n5227_), .ZN(new_n6458_));
  NOR2_X1    g05456(.A1(new_n5221_), .A2(new_n5223_), .ZN(new_n6459_));
  NOR2_X1    g05457(.A1(new_n5195_), .A2(new_n2990_), .ZN(new_n6460_));
  AOI21_X1   g05458(.A1(new_n6460_), .A2(new_n5210_), .B(new_n5200_), .ZN(new_n6461_));
  OAI21_X1   g05459(.A1(new_n6459_), .A2(new_n5219_), .B(new_n6461_), .ZN(new_n6462_));
  NAND2_X1   g05460(.A1(new_n5225_), .A2(new_n5217_), .ZN(new_n6463_));
  NAND2_X1   g05461(.A1(new_n5208_), .A2(new_n2991_), .ZN(new_n6464_));
  OAI21_X1   g05462(.A1(new_n6464_), .A2(new_n5205_), .B(new_n5209_), .ZN(new_n6465_));
  NAND3_X1   g05463(.A1(new_n6465_), .A2(new_n6463_), .A3(new_n5224_), .ZN(new_n6466_));
  NAND2_X1   g05464(.A1(new_n6462_), .A2(new_n6466_), .ZN(new_n6467_));
  AOI21_X1   g05465(.A1(new_n6458_), .A2(new_n5233_), .B(new_n6467_), .ZN(new_n6468_));
  NOR2_X1    g05466(.A1(new_n5236_), .A2(new_n5234_), .ZN(new_n6469_));
  AOI21_X1   g05467(.A1(new_n5224_), .A2(new_n6463_), .B(new_n6465_), .ZN(new_n6470_));
  NOR3_X1    g05468(.A1(new_n6461_), .A2(new_n6459_), .A3(new_n5219_), .ZN(new_n6471_));
  NOR2_X1    g05469(.A1(new_n6470_), .A2(new_n6471_), .ZN(new_n6472_));
  NOR3_X1    g05470(.A1(new_n6469_), .A2(new_n6472_), .A3(new_n5237_), .ZN(new_n6473_));
  NOR2_X1    g05471(.A1(new_n5287_), .A2(new_n5240_), .ZN(new_n6474_));
  NAND2_X1   g05472(.A1(new_n5275_), .A2(new_n5267_), .ZN(new_n6475_));
  OAI21_X1   g05473(.A1(new_n5279_), .A2(new_n5253_), .B(new_n5259_), .ZN(new_n6476_));
  AOI21_X1   g05474(.A1(new_n6475_), .A2(new_n5274_), .B(new_n6476_), .ZN(new_n6477_));
  NOR2_X1    g05475(.A1(new_n5271_), .A2(new_n5273_), .ZN(new_n6478_));
  AOI21_X1   g05476(.A1(new_n2949_), .A2(new_n2930_), .B(new_n2942_), .ZN(new_n6479_));
  AOI21_X1   g05477(.A1(new_n6479_), .A2(new_n5260_), .B(new_n5248_), .ZN(new_n6480_));
  NOR3_X1    g05478(.A1(new_n6478_), .A2(new_n6480_), .A3(new_n5269_), .ZN(new_n6481_));
  NOR2_X1    g05479(.A1(new_n6477_), .A2(new_n6481_), .ZN(new_n6482_));
  OAI21_X1   g05480(.A1(new_n6474_), .A2(new_n5288_), .B(new_n6482_), .ZN(new_n6483_));
  NAND2_X1   g05481(.A1(new_n5277_), .A2(new_n5286_), .ZN(new_n6484_));
  OAI21_X1   g05482(.A1(new_n6478_), .A2(new_n5269_), .B(new_n6480_), .ZN(new_n6485_));
  NAND3_X1   g05483(.A1(new_n6475_), .A2(new_n6476_), .A3(new_n5274_), .ZN(new_n6486_));
  NAND2_X1   g05484(.A1(new_n6486_), .A2(new_n6485_), .ZN(new_n6487_));
  NAND3_X1   g05485(.A1(new_n6484_), .A2(new_n5284_), .A3(new_n6487_), .ZN(new_n6488_));
  NAND2_X1   g05486(.A1(new_n6483_), .A2(new_n6488_), .ZN(new_n6489_));
  NOR3_X1    g05487(.A1(new_n6489_), .A2(new_n6468_), .A3(new_n6473_), .ZN(new_n6490_));
  OAI21_X1   g05488(.A1(new_n6469_), .A2(new_n5237_), .B(new_n6472_), .ZN(new_n6491_));
  NAND3_X1   g05489(.A1(new_n6458_), .A2(new_n6467_), .A3(new_n5233_), .ZN(new_n6492_));
  AOI22_X1   g05490(.A1(new_n6491_), .A2(new_n6492_), .B1(new_n6483_), .B2(new_n6488_), .ZN(new_n6493_));
  NOR3_X1    g05491(.A1(new_n6457_), .A2(new_n6490_), .A3(new_n6493_), .ZN(new_n6494_));
  OAI21_X1   g05492(.A1(new_n5299_), .A2(new_n5300_), .B(new_n5290_), .ZN(new_n6495_));
  NAND4_X1   g05493(.A1(new_n6491_), .A2(new_n6492_), .A3(new_n6483_), .A4(new_n6488_), .ZN(new_n6496_));
  AOI21_X1   g05494(.A1(new_n6484_), .A2(new_n5284_), .B(new_n6487_), .ZN(new_n6497_));
  NOR3_X1    g05495(.A1(new_n6474_), .A2(new_n5288_), .A3(new_n6482_), .ZN(new_n6498_));
  OAI22_X1   g05496(.A1(new_n6468_), .A2(new_n6473_), .B1(new_n6498_), .B2(new_n6497_), .ZN(new_n6499_));
  AOI21_X1   g05497(.A1(new_n6496_), .A2(new_n6499_), .B(new_n6495_), .ZN(new_n6500_));
  NOR4_X1    g05498(.A1(new_n6454_), .A2(new_n6494_), .A3(new_n6500_), .A4(new_n6456_), .ZN(new_n6501_));
  NAND3_X1   g05499(.A1(new_n6455_), .A2(new_n6447_), .A3(new_n6452_), .ZN(new_n6502_));
  NAND2_X1   g05500(.A1(new_n6453_), .A2(new_n6415_), .ZN(new_n6503_));
  NAND3_X1   g05501(.A1(new_n6495_), .A2(new_n6496_), .A3(new_n6499_), .ZN(new_n6504_));
  OAI21_X1   g05502(.A1(new_n6490_), .A2(new_n6493_), .B(new_n6457_), .ZN(new_n6505_));
  AOI22_X1   g05503(.A1(new_n6505_), .A2(new_n6504_), .B1(new_n6503_), .B2(new_n6502_), .ZN(new_n6506_));
  NOR3_X1    g05504(.A1(new_n6501_), .A2(new_n6506_), .A3(new_n6414_), .ZN(new_n6507_));
  OAI21_X1   g05505(.A1(new_n5426_), .A2(new_n5427_), .B(new_n5417_), .ZN(new_n6508_));
  NAND4_X1   g05506(.A1(new_n6505_), .A2(new_n6503_), .A3(new_n6502_), .A4(new_n6504_), .ZN(new_n6509_));
  OAI22_X1   g05507(.A1(new_n6494_), .A2(new_n6500_), .B1(new_n6454_), .B2(new_n6456_), .ZN(new_n6510_));
  AOI21_X1   g05508(.A1(new_n6510_), .A2(new_n6509_), .B(new_n6508_), .ZN(new_n6511_));
  NOR4_X1    g05509(.A1(new_n6507_), .A2(new_n6511_), .A3(new_n6409_), .A4(new_n6413_), .ZN(new_n6512_));
  NAND3_X1   g05510(.A1(new_n6411_), .A2(new_n6412_), .A3(new_n6410_), .ZN(new_n6513_));
  OAI21_X1   g05511(.A1(new_n6408_), .A2(new_n6403_), .B(new_n6326_), .ZN(new_n6514_));
  NAND3_X1   g05512(.A1(new_n6510_), .A2(new_n6508_), .A3(new_n6509_), .ZN(new_n6515_));
  OAI21_X1   g05513(.A1(new_n6501_), .A2(new_n6506_), .B(new_n6414_), .ZN(new_n6516_));
  AOI22_X1   g05514(.A1(new_n6516_), .A2(new_n6515_), .B1(new_n6514_), .B2(new_n6513_), .ZN(new_n6517_));
  NOR3_X1    g05515(.A1(new_n6512_), .A2(new_n6517_), .A3(new_n6325_), .ZN(new_n6518_));
  OAI21_X1   g05516(.A1(new_n5658_), .A2(new_n5659_), .B(new_n5649_), .ZN(new_n6519_));
  NAND4_X1   g05517(.A1(new_n6516_), .A2(new_n6515_), .A3(new_n6514_), .A4(new_n6513_), .ZN(new_n6520_));
  OAI22_X1   g05518(.A1(new_n6507_), .A2(new_n6511_), .B1(new_n6409_), .B2(new_n6413_), .ZN(new_n6521_));
  AOI21_X1   g05519(.A1(new_n6521_), .A2(new_n6520_), .B(new_n6519_), .ZN(new_n6522_));
  NOR4_X1    g05520(.A1(new_n6320_), .A2(new_n6324_), .A3(new_n6518_), .A4(new_n6522_), .ZN(new_n6523_));
  OAI22_X1   g05521(.A1(new_n6320_), .A2(new_n6324_), .B1(new_n6518_), .B2(new_n6522_), .ZN(new_n6524_));
  AOI21_X1   g05522(.A1(new_n6126_), .A2(new_n6524_), .B(new_n6523_), .ZN(new_n6525_));
  AOI21_X1   g05523(.A1(new_n6519_), .A2(new_n6521_), .B(new_n6512_), .ZN(new_n6526_));
  OAI21_X1   g05524(.A1(new_n6506_), .A2(new_n6414_), .B(new_n6509_), .ZN(new_n6527_));
  NAND2_X1   g05525(.A1(new_n6442_), .A2(new_n5398_), .ZN(new_n6528_));
  AOI21_X1   g05526(.A1(new_n6433_), .A2(new_n5388_), .B(new_n6438_), .ZN(new_n6529_));
  INV_X1     g05527(.I(new_n6529_), .ZN(new_n6530_));
  NOR3_X1    g05528(.A1(new_n6435_), .A2(new_n6437_), .A3(new_n5383_), .ZN(new_n6531_));
  OAI21_X1   g05529(.A1(new_n6528_), .A2(new_n6531_), .B(new_n6530_), .ZN(new_n6532_));
  NOR2_X1    g05530(.A1(new_n6421_), .A2(new_n5332_), .ZN(new_n6533_));
  NOR2_X1    g05531(.A1(new_n6533_), .A2(new_n6423_), .ZN(new_n6534_));
  AOI21_X1   g05532(.A1(new_n6427_), .A2(new_n5346_), .B(new_n6534_), .ZN(new_n6535_));
  AOI21_X1   g05533(.A1(new_n6533_), .A2(new_n6423_), .B(new_n6535_), .ZN(new_n6536_));
  NOR2_X1    g05534(.A1(new_n6536_), .A2(new_n6532_), .ZN(new_n6537_));
  NOR2_X1    g05535(.A1(new_n6416_), .A2(new_n5350_), .ZN(new_n6538_));
  NAND2_X1   g05536(.A1(new_n6538_), .A2(new_n6425_), .ZN(new_n6539_));
  NAND2_X1   g05537(.A1(new_n6533_), .A2(new_n6423_), .ZN(new_n6540_));
  AOI22_X1   g05538(.A1(new_n6441_), .A2(new_n6446_), .B1(new_n6535_), .B2(new_n6540_), .ZN(new_n6541_));
  AOI22_X1   g05539(.A1(new_n6415_), .A2(new_n6447_), .B1(new_n6539_), .B2(new_n6541_), .ZN(new_n6542_));
  INV_X1     g05540(.I(new_n6532_), .ZN(new_n6543_));
  OAI21_X1   g05541(.A1(new_n6538_), .A2(new_n6534_), .B(new_n6540_), .ZN(new_n6544_));
  NOR2_X1    g05542(.A1(new_n6543_), .A2(new_n6544_), .ZN(new_n6545_));
  NOR3_X1    g05543(.A1(new_n6542_), .A2(new_n6537_), .A3(new_n6545_), .ZN(new_n6546_));
  INV_X1     g05544(.I(new_n6447_), .ZN(new_n6547_));
  NAND2_X1   g05545(.A1(new_n6541_), .A2(new_n6539_), .ZN(new_n6548_));
  OAI21_X1   g05546(.A1(new_n6455_), .A2(new_n6547_), .B(new_n6548_), .ZN(new_n6549_));
  NOR2_X1    g05547(.A1(new_n6545_), .A2(new_n6537_), .ZN(new_n6550_));
  NOR2_X1    g05548(.A1(new_n6549_), .A2(new_n6550_), .ZN(new_n6551_));
  NAND2_X1   g05549(.A1(new_n6484_), .A2(new_n5284_), .ZN(new_n6552_));
  NOR2_X1    g05550(.A1(new_n6478_), .A2(new_n5269_), .ZN(new_n6553_));
  NOR2_X1    g05551(.A1(new_n6553_), .A2(new_n6480_), .ZN(new_n6554_));
  INV_X1     g05552(.I(new_n6554_), .ZN(new_n6555_));
  NAND2_X1   g05553(.A1(new_n6553_), .A2(new_n6480_), .ZN(new_n6556_));
  INV_X1     g05554(.I(new_n6556_), .ZN(new_n6557_));
  OAI21_X1   g05555(.A1(new_n6552_), .A2(new_n6557_), .B(new_n6555_), .ZN(new_n6558_));
  NOR2_X1    g05556(.A1(new_n6459_), .A2(new_n5219_), .ZN(new_n6559_));
  NOR2_X1    g05557(.A1(new_n6559_), .A2(new_n6461_), .ZN(new_n6560_));
  AOI21_X1   g05558(.A1(new_n6458_), .A2(new_n5233_), .B(new_n6560_), .ZN(new_n6561_));
  AOI21_X1   g05559(.A1(new_n6559_), .A2(new_n6461_), .B(new_n6561_), .ZN(new_n6562_));
  NOR2_X1    g05560(.A1(new_n6562_), .A2(new_n6558_), .ZN(new_n6563_));
  NOR2_X1    g05561(.A1(new_n6469_), .A2(new_n5237_), .ZN(new_n6564_));
  NAND2_X1   g05562(.A1(new_n6564_), .A2(new_n6472_), .ZN(new_n6565_));
  NAND2_X1   g05563(.A1(new_n6559_), .A2(new_n6461_), .ZN(new_n6566_));
  AOI22_X1   g05564(.A1(new_n6561_), .A2(new_n6566_), .B1(new_n6483_), .B2(new_n6488_), .ZN(new_n6567_));
  AOI22_X1   g05565(.A1(new_n6457_), .A2(new_n6496_), .B1(new_n6565_), .B2(new_n6567_), .ZN(new_n6568_));
  INV_X1     g05566(.I(new_n6558_), .ZN(new_n6569_));
  OAI21_X1   g05567(.A1(new_n6564_), .A2(new_n6560_), .B(new_n6566_), .ZN(new_n6570_));
  NOR2_X1    g05568(.A1(new_n6569_), .A2(new_n6570_), .ZN(new_n6571_));
  NOR3_X1    g05569(.A1(new_n6568_), .A2(new_n6563_), .A3(new_n6571_), .ZN(new_n6572_));
  NAND2_X1   g05570(.A1(new_n6561_), .A2(new_n6566_), .ZN(new_n6573_));
  NAND3_X1   g05571(.A1(new_n6573_), .A2(new_n6489_), .A3(new_n6565_), .ZN(new_n6574_));
  OAI21_X1   g05572(.A1(new_n6495_), .A2(new_n6490_), .B(new_n6574_), .ZN(new_n6575_));
  NOR2_X1    g05573(.A1(new_n6563_), .A2(new_n6571_), .ZN(new_n6576_));
  NOR2_X1    g05574(.A1(new_n6575_), .A2(new_n6576_), .ZN(new_n6577_));
  OAI22_X1   g05575(.A1(new_n6546_), .A2(new_n6551_), .B1(new_n6577_), .B2(new_n6572_), .ZN(new_n6578_));
  NAND2_X1   g05576(.A1(new_n6543_), .A2(new_n6544_), .ZN(new_n6579_));
  NAND2_X1   g05577(.A1(new_n6536_), .A2(new_n6532_), .ZN(new_n6580_));
  NAND3_X1   g05578(.A1(new_n6549_), .A2(new_n6579_), .A3(new_n6580_), .ZN(new_n6581_));
  NAND2_X1   g05579(.A1(new_n6579_), .A2(new_n6580_), .ZN(new_n6582_));
  NAND2_X1   g05580(.A1(new_n6542_), .A2(new_n6582_), .ZN(new_n6583_));
  NAND2_X1   g05581(.A1(new_n6569_), .A2(new_n6570_), .ZN(new_n6584_));
  NAND2_X1   g05582(.A1(new_n6562_), .A2(new_n6558_), .ZN(new_n6585_));
  NAND3_X1   g05583(.A1(new_n6575_), .A2(new_n6584_), .A3(new_n6585_), .ZN(new_n6586_));
  NAND2_X1   g05584(.A1(new_n6585_), .A2(new_n6584_), .ZN(new_n6587_));
  NAND2_X1   g05585(.A1(new_n6587_), .A2(new_n6568_), .ZN(new_n6588_));
  NAND4_X1   g05586(.A1(new_n6581_), .A2(new_n6586_), .A3(new_n6588_), .A4(new_n6583_), .ZN(new_n6589_));
  AOI21_X1   g05587(.A1(new_n6578_), .A2(new_n6589_), .B(new_n6527_), .ZN(new_n6590_));
  AOI21_X1   g05588(.A1(new_n6508_), .A2(new_n6510_), .B(new_n6501_), .ZN(new_n6591_));
  AOI22_X1   g05589(.A1(new_n6581_), .A2(new_n6583_), .B1(new_n6586_), .B2(new_n6588_), .ZN(new_n6592_));
  NOR4_X1    g05590(.A1(new_n6551_), .A2(new_n6577_), .A3(new_n6572_), .A4(new_n6546_), .ZN(new_n6593_));
  NOR3_X1    g05591(.A1(new_n6591_), .A2(new_n6592_), .A3(new_n6593_), .ZN(new_n6594_));
  OAI21_X1   g05592(.A1(new_n6408_), .A2(new_n6326_), .B(new_n6411_), .ZN(new_n6595_));
  NAND2_X1   g05593(.A1(new_n6367_), .A2(new_n6400_), .ZN(new_n6596_));
  NOR2_X1    g05594(.A1(new_n6369_), .A2(new_n5460_), .ZN(new_n6597_));
  NAND2_X1   g05595(.A1(new_n6597_), .A2(new_n6371_), .ZN(new_n6598_));
  NOR2_X1    g05596(.A1(new_n6597_), .A2(new_n6371_), .ZN(new_n6599_));
  AOI21_X1   g05597(.A1(new_n6368_), .A2(new_n5474_), .B(new_n6599_), .ZN(new_n6600_));
  NAND2_X1   g05598(.A1(new_n6600_), .A2(new_n6598_), .ZN(new_n6601_));
  INV_X1     g05599(.I(new_n6385_), .ZN(new_n6602_));
  AOI21_X1   g05600(.A1(new_n5499_), .A2(new_n5507_), .B(new_n5511_), .ZN(new_n6603_));
  NOR2_X1    g05601(.A1(new_n6602_), .A2(new_n6603_), .ZN(new_n6604_));
  INV_X1     g05602(.I(new_n6604_), .ZN(new_n6605_));
  NOR2_X1    g05603(.A1(new_n6386_), .A2(new_n6385_), .ZN(new_n6606_));
  NOR2_X1    g05604(.A1(new_n6384_), .A2(new_n6606_), .ZN(new_n6607_));
  AOI22_X1   g05605(.A1(new_n6607_), .A2(new_n6605_), .B1(new_n6384_), .B2(new_n6390_), .ZN(new_n6608_));
  NAND3_X1   g05606(.A1(new_n6368_), .A2(new_n6382_), .A3(new_n5474_), .ZN(new_n6609_));
  NAND3_X1   g05607(.A1(new_n6608_), .A2(new_n6601_), .A3(new_n6609_), .ZN(new_n6610_));
  INV_X1     g05608(.I(new_n6598_), .ZN(new_n6611_));
  INV_X1     g05609(.I(new_n6606_), .ZN(new_n6612_));
  AOI21_X1   g05610(.A1(new_n6389_), .A2(new_n6612_), .B(new_n6604_), .ZN(new_n6613_));
  NOR3_X1    g05611(.A1(new_n6613_), .A2(new_n6600_), .A3(new_n6611_), .ZN(new_n6614_));
  INV_X1     g05612(.I(new_n6614_), .ZN(new_n6615_));
  OAI21_X1   g05613(.A1(new_n6611_), .A2(new_n6600_), .B(new_n6613_), .ZN(new_n6616_));
  NAND2_X1   g05614(.A1(new_n6615_), .A2(new_n6616_), .ZN(new_n6617_));
  AOI21_X1   g05615(.A1(new_n6596_), .A2(new_n6610_), .B(new_n6617_), .ZN(new_n6618_));
  NOR2_X1    g05616(.A1(new_n6399_), .A2(new_n6392_), .ZN(new_n6619_));
  INV_X1     g05617(.I(new_n6610_), .ZN(new_n6620_));
  INV_X1     g05618(.I(new_n6616_), .ZN(new_n6621_));
  NOR2_X1    g05619(.A1(new_n6621_), .A2(new_n6614_), .ZN(new_n6622_));
  NOR3_X1    g05620(.A1(new_n6622_), .A2(new_n6620_), .A3(new_n6619_), .ZN(new_n6623_));
  NOR2_X1    g05621(.A1(new_n6618_), .A2(new_n6623_), .ZN(new_n6624_));
  NOR2_X1    g05622(.A1(new_n6340_), .A2(new_n5579_), .ZN(new_n6625_));
  NOR2_X1    g05623(.A1(new_n6341_), .A2(new_n5560_), .ZN(new_n6626_));
  NAND2_X1   g05624(.A1(new_n6626_), .A2(new_n6343_), .ZN(new_n6627_));
  NOR2_X1    g05625(.A1(new_n6626_), .A2(new_n6343_), .ZN(new_n6628_));
  OAI21_X1   g05626(.A1(new_n6625_), .A2(new_n6628_), .B(new_n6627_), .ZN(new_n6629_));
  AOI21_X1   g05627(.A1(new_n5623_), .A2(new_n5616_), .B(new_n5625_), .ZN(new_n6630_));
  NAND2_X1   g05628(.A1(new_n6330_), .A2(new_n6333_), .ZN(new_n6631_));
  NOR2_X1    g05629(.A1(new_n6330_), .A2(new_n6333_), .ZN(new_n6632_));
  OAI21_X1   g05630(.A1(new_n6630_), .A2(new_n6632_), .B(new_n6631_), .ZN(new_n6633_));
  INV_X1     g05631(.I(new_n6633_), .ZN(new_n6634_));
  NAND2_X1   g05632(.A1(new_n6629_), .A2(new_n6634_), .ZN(new_n6635_));
  NAND2_X1   g05633(.A1(new_n6351_), .A2(new_n5575_), .ZN(new_n6636_));
  INV_X1     g05634(.I(new_n6627_), .ZN(new_n6637_));
  INV_X1     g05635(.I(new_n6628_), .ZN(new_n6638_));
  AOI21_X1   g05636(.A1(new_n6636_), .A2(new_n6638_), .B(new_n6637_), .ZN(new_n6639_));
  NAND2_X1   g05637(.A1(new_n6639_), .A2(new_n6633_), .ZN(new_n6640_));
  NAND2_X1   g05638(.A1(new_n6635_), .A2(new_n6640_), .ZN(new_n6641_));
  NOR2_X1    g05639(.A1(new_n6363_), .A2(new_n6356_), .ZN(new_n6642_));
  OAI21_X1   g05640(.A1(new_n6642_), .A2(new_n6361_), .B(new_n6641_), .ZN(new_n6643_));
  NOR2_X1    g05641(.A1(new_n6639_), .A2(new_n6633_), .ZN(new_n6644_));
  NOR2_X1    g05642(.A1(new_n6629_), .A2(new_n6634_), .ZN(new_n6645_));
  NOR2_X1    g05643(.A1(new_n6645_), .A2(new_n6644_), .ZN(new_n6646_));
  NAND2_X1   g05644(.A1(new_n6327_), .A2(new_n6364_), .ZN(new_n6647_));
  NAND3_X1   g05645(.A1(new_n6647_), .A2(new_n6646_), .A3(new_n6365_), .ZN(new_n6648_));
  NAND2_X1   g05646(.A1(new_n6643_), .A2(new_n6648_), .ZN(new_n6649_));
  NAND2_X1   g05647(.A1(new_n6649_), .A2(new_n6624_), .ZN(new_n6650_));
  OAI21_X1   g05648(.A1(new_n6619_), .A2(new_n6620_), .B(new_n6622_), .ZN(new_n6651_));
  NAND3_X1   g05649(.A1(new_n6596_), .A2(new_n6617_), .A3(new_n6610_), .ZN(new_n6652_));
  NAND2_X1   g05650(.A1(new_n6651_), .A2(new_n6652_), .ZN(new_n6653_));
  AOI21_X1   g05651(.A1(new_n6647_), .A2(new_n6365_), .B(new_n6646_), .ZN(new_n6654_));
  NOR3_X1    g05652(.A1(new_n6641_), .A2(new_n6642_), .A3(new_n6361_), .ZN(new_n6655_));
  NOR2_X1    g05653(.A1(new_n6654_), .A2(new_n6655_), .ZN(new_n6656_));
  NAND2_X1   g05654(.A1(new_n6656_), .A2(new_n6653_), .ZN(new_n6657_));
  AOI21_X1   g05655(.A1(new_n6650_), .A2(new_n6657_), .B(new_n6595_), .ZN(new_n6658_));
  AOI21_X1   g05656(.A1(new_n6410_), .A2(new_n6412_), .B(new_n6403_), .ZN(new_n6659_));
  NOR2_X1    g05657(.A1(new_n6656_), .A2(new_n6653_), .ZN(new_n6660_));
  NOR2_X1    g05658(.A1(new_n6649_), .A2(new_n6624_), .ZN(new_n6661_));
  NOR3_X1    g05659(.A1(new_n6661_), .A2(new_n6660_), .A3(new_n6659_), .ZN(new_n6662_));
  NOR4_X1    g05660(.A1(new_n6590_), .A2(new_n6594_), .A3(new_n6658_), .A4(new_n6662_), .ZN(new_n6663_));
  OAI21_X1   g05661(.A1(new_n6592_), .A2(new_n6593_), .B(new_n6591_), .ZN(new_n6664_));
  NAND3_X1   g05662(.A1(new_n6578_), .A2(new_n6527_), .A3(new_n6589_), .ZN(new_n6665_));
  OAI21_X1   g05663(.A1(new_n6661_), .A2(new_n6660_), .B(new_n6659_), .ZN(new_n6666_));
  NAND3_X1   g05664(.A1(new_n6650_), .A2(new_n6657_), .A3(new_n6595_), .ZN(new_n6667_));
  AOI22_X1   g05665(.A1(new_n6664_), .A2(new_n6665_), .B1(new_n6666_), .B2(new_n6667_), .ZN(new_n6668_));
  NOR3_X1    g05666(.A1(new_n6663_), .A2(new_n6668_), .A3(new_n6526_), .ZN(new_n6669_));
  OAI21_X1   g05667(.A1(new_n6325_), .A2(new_n6517_), .B(new_n6520_), .ZN(new_n6670_));
  NAND4_X1   g05668(.A1(new_n6664_), .A2(new_n6665_), .A3(new_n6666_), .A4(new_n6667_), .ZN(new_n6671_));
  OAI22_X1   g05669(.A1(new_n6590_), .A2(new_n6594_), .B1(new_n6658_), .B2(new_n6662_), .ZN(new_n6672_));
  AOI21_X1   g05670(.A1(new_n6672_), .A2(new_n6671_), .B(new_n6670_), .ZN(new_n6673_));
  AOI21_X1   g05671(.A1(new_n6321_), .A2(new_n6323_), .B(new_n6314_), .ZN(new_n6674_));
  OAI21_X1   g05672(.A1(new_n6308_), .A2(new_n6216_), .B(new_n6311_), .ZN(new_n6675_));
  NAND2_X1   g05673(.A1(new_n5761_), .A2(new_n5762_), .ZN(new_n6676_));
  NAND3_X1   g05674(.A1(new_n6676_), .A2(new_n6300_), .A3(new_n5756_), .ZN(new_n6677_));
  NOR2_X1    g05675(.A1(new_n6259_), .A2(new_n5686_), .ZN(new_n6678_));
  NAND2_X1   g05676(.A1(new_n6678_), .A2(new_n6261_), .ZN(new_n6679_));
  INV_X1     g05677(.I(new_n6679_), .ZN(new_n6680_));
  NOR2_X1    g05678(.A1(new_n6678_), .A2(new_n6261_), .ZN(new_n6681_));
  NOR3_X1    g05679(.A1(new_n6258_), .A2(new_n6680_), .A3(new_n6681_), .ZN(new_n6682_));
  AOI21_X1   g05680(.A1(new_n5752_), .A2(new_n5744_), .B(new_n5754_), .ZN(new_n6683_));
  NOR2_X1    g05681(.A1(new_n6277_), .A2(new_n6279_), .ZN(new_n6684_));
  NAND2_X1   g05682(.A1(new_n6277_), .A2(new_n6279_), .ZN(new_n6685_));
  INV_X1     g05683(.I(new_n6685_), .ZN(new_n6686_));
  NOR3_X1    g05684(.A1(new_n6683_), .A2(new_n6684_), .A3(new_n6686_), .ZN(new_n6687_));
  NAND2_X1   g05685(.A1(new_n6274_), .A2(new_n5750_), .ZN(new_n6688_));
  NOR2_X1    g05686(.A1(new_n6688_), .A2(new_n6283_), .ZN(new_n6689_));
  NOR2_X1    g05687(.A1(new_n6291_), .A2(new_n6267_), .ZN(new_n6690_));
  NOR4_X1    g05688(.A1(new_n6689_), .A2(new_n6682_), .A3(new_n6687_), .A4(new_n6690_), .ZN(new_n6691_));
  INV_X1     g05689(.I(new_n6691_), .ZN(new_n6692_));
  INV_X1     g05690(.I(new_n6684_), .ZN(new_n6693_));
  OAI21_X1   g05691(.A1(new_n6683_), .A2(new_n6686_), .B(new_n6693_), .ZN(new_n6694_));
  INV_X1     g05692(.I(new_n6681_), .ZN(new_n6695_));
  AOI21_X1   g05693(.A1(new_n6291_), .A2(new_n6695_), .B(new_n6680_), .ZN(new_n6696_));
  NAND2_X1   g05694(.A1(new_n6696_), .A2(new_n6694_), .ZN(new_n6697_));
  AOI21_X1   g05695(.A1(new_n6688_), .A2(new_n6685_), .B(new_n6684_), .ZN(new_n6698_));
  OAI21_X1   g05696(.A1(new_n6258_), .A2(new_n6681_), .B(new_n6679_), .ZN(new_n6699_));
  NAND2_X1   g05697(.A1(new_n6698_), .A2(new_n6699_), .ZN(new_n6700_));
  NAND2_X1   g05698(.A1(new_n6700_), .A2(new_n6697_), .ZN(new_n6701_));
  AOI21_X1   g05699(.A1(new_n6677_), .A2(new_n6692_), .B(new_n6701_), .ZN(new_n6702_));
  NOR2_X1    g05700(.A1(new_n6299_), .A2(new_n6290_), .ZN(new_n6703_));
  XOR2_X1    g05701(.A1(new_n6696_), .A2(new_n6694_), .Z(new_n6704_));
  NOR3_X1    g05702(.A1(new_n6703_), .A2(new_n6704_), .A3(new_n6691_), .ZN(new_n6705_));
  NOR2_X1    g05703(.A1(new_n6705_), .A2(new_n6702_), .ZN(new_n6706_));
  NAND2_X1   g05704(.A1(new_n6235_), .A2(new_n5802_), .ZN(new_n6707_));
  NOR2_X1    g05705(.A1(new_n6707_), .A2(new_n6237_), .ZN(new_n6708_));
  NAND2_X1   g05706(.A1(new_n6707_), .A2(new_n6237_), .ZN(new_n6709_));
  AOI21_X1   g05707(.A1(new_n6230_), .A2(new_n6709_), .B(new_n6708_), .ZN(new_n6710_));
  INV_X1     g05708(.I(new_n6220_), .ZN(new_n6711_));
  INV_X1     g05709(.I(new_n6223_), .ZN(new_n6712_));
  NOR2_X1    g05710(.A1(new_n6711_), .A2(new_n6712_), .ZN(new_n6713_));
  NOR2_X1    g05711(.A1(new_n6220_), .A2(new_n6223_), .ZN(new_n6714_));
  INV_X1     g05712(.I(new_n6714_), .ZN(new_n6715_));
  AOI21_X1   g05713(.A1(new_n6218_), .A2(new_n6715_), .B(new_n6713_), .ZN(new_n6716_));
  XOR2_X1    g05714(.A1(new_n6710_), .A2(new_n6716_), .Z(new_n6717_));
  NOR2_X1    g05715(.A1(new_n6253_), .A2(new_n6246_), .ZN(new_n6718_));
  OAI21_X1   g05716(.A1(new_n6718_), .A2(new_n6251_), .B(new_n6717_), .ZN(new_n6719_));
  AOI21_X1   g05717(.A1(new_n6228_), .A2(new_n5859_), .B(new_n6714_), .ZN(new_n6720_));
  NOR3_X1    g05718(.A1(new_n6710_), .A2(new_n6713_), .A3(new_n6720_), .ZN(new_n6721_));
  AOI22_X1   g05719(.A1(new_n6241_), .A2(new_n5811_), .B1(new_n6707_), .B2(new_n6237_), .ZN(new_n6722_));
  NOR3_X1    g05720(.A1(new_n6716_), .A2(new_n6722_), .A3(new_n6708_), .ZN(new_n6723_));
  NOR2_X1    g05721(.A1(new_n6721_), .A2(new_n6723_), .ZN(new_n6724_));
  NAND2_X1   g05722(.A1(new_n5870_), .A2(new_n5771_), .ZN(new_n6725_));
  NAND3_X1   g05723(.A1(new_n6725_), .A2(new_n6254_), .A3(new_n5865_), .ZN(new_n6726_));
  NAND3_X1   g05724(.A1(new_n6726_), .A2(new_n6255_), .A3(new_n6724_), .ZN(new_n6727_));
  NAND2_X1   g05725(.A1(new_n6719_), .A2(new_n6727_), .ZN(new_n6728_));
  NAND2_X1   g05726(.A1(new_n6706_), .A2(new_n6728_), .ZN(new_n6729_));
  OAI21_X1   g05727(.A1(new_n6703_), .A2(new_n6691_), .B(new_n6704_), .ZN(new_n6730_));
  NAND3_X1   g05728(.A1(new_n6677_), .A2(new_n6692_), .A3(new_n6701_), .ZN(new_n6731_));
  NAND2_X1   g05729(.A1(new_n6730_), .A2(new_n6731_), .ZN(new_n6732_));
  AOI21_X1   g05730(.A1(new_n6726_), .A2(new_n6255_), .B(new_n6724_), .ZN(new_n6733_));
  NOR3_X1    g05731(.A1(new_n6718_), .A2(new_n6717_), .A3(new_n6251_), .ZN(new_n6734_));
  NOR2_X1    g05732(.A1(new_n6734_), .A2(new_n6733_), .ZN(new_n6735_));
  NAND2_X1   g05733(.A1(new_n6732_), .A2(new_n6735_), .ZN(new_n6736_));
  AOI21_X1   g05734(.A1(new_n6729_), .A2(new_n6736_), .B(new_n6675_), .ZN(new_n6737_));
  AOI21_X1   g05735(.A1(new_n6310_), .A2(new_n6312_), .B(new_n6303_), .ZN(new_n6738_));
  NOR2_X1    g05736(.A1(new_n6732_), .A2(new_n6735_), .ZN(new_n6739_));
  NOR2_X1    g05737(.A1(new_n6706_), .A2(new_n6728_), .ZN(new_n6740_));
  NOR3_X1    g05738(.A1(new_n6738_), .A2(new_n6739_), .A3(new_n6740_), .ZN(new_n6741_));
  OAI21_X1   g05739(.A1(new_n6210_), .A2(new_n6128_), .B(new_n6213_), .ZN(new_n6742_));
  NAND2_X1   g05740(.A1(new_n5993_), .A2(new_n5996_), .ZN(new_n6743_));
  NAND3_X1   g05741(.A1(new_n6743_), .A2(new_n6202_), .A3(new_n5988_), .ZN(new_n6744_));
  NOR2_X1    g05742(.A1(new_n6170_), .A2(new_n5919_), .ZN(new_n6745_));
  NAND2_X1   g05743(.A1(new_n6745_), .A2(new_n6172_), .ZN(new_n6746_));
  NOR2_X1    g05744(.A1(new_n6745_), .A2(new_n6172_), .ZN(new_n6747_));
  AOI21_X1   g05745(.A1(new_n6169_), .A2(new_n5933_), .B(new_n6747_), .ZN(new_n6748_));
  NAND2_X1   g05746(.A1(new_n6748_), .A2(new_n6746_), .ZN(new_n6749_));
  INV_X1     g05747(.I(new_n6186_), .ZN(new_n6750_));
  NOR2_X1    g05748(.A1(new_n6750_), .A2(new_n6191_), .ZN(new_n6751_));
  NOR2_X1    g05749(.A1(new_n6187_), .A2(new_n6186_), .ZN(new_n6752_));
  NOR3_X1    g05750(.A1(new_n6185_), .A2(new_n6751_), .A3(new_n6752_), .ZN(new_n6753_));
  NOR2_X1    g05751(.A1(new_n6190_), .A2(new_n6188_), .ZN(new_n6754_));
  NOR2_X1    g05752(.A1(new_n6753_), .A2(new_n6754_), .ZN(new_n6755_));
  NAND3_X1   g05753(.A1(new_n6169_), .A2(new_n6183_), .A3(new_n5933_), .ZN(new_n6756_));
  NAND3_X1   g05754(.A1(new_n6755_), .A2(new_n6749_), .A3(new_n6756_), .ZN(new_n6757_));
  OAI22_X1   g05755(.A1(new_n6180_), .A2(new_n5937_), .B1(new_n6745_), .B2(new_n6172_), .ZN(new_n6758_));
  INV_X1     g05756(.I(new_n6751_), .ZN(new_n6759_));
  OAI21_X1   g05757(.A1(new_n6185_), .A2(new_n6752_), .B(new_n6759_), .ZN(new_n6760_));
  NAND3_X1   g05758(.A1(new_n6758_), .A2(new_n6760_), .A3(new_n6746_), .ZN(new_n6761_));
  INV_X1     g05759(.I(new_n6746_), .ZN(new_n6762_));
  INV_X1     g05760(.I(new_n6752_), .ZN(new_n6763_));
  AOI21_X1   g05761(.A1(new_n6190_), .A2(new_n6763_), .B(new_n6751_), .ZN(new_n6764_));
  OAI21_X1   g05762(.A1(new_n6762_), .A2(new_n6748_), .B(new_n6764_), .ZN(new_n6765_));
  NAND2_X1   g05763(.A1(new_n6761_), .A2(new_n6765_), .ZN(new_n6766_));
  AOI21_X1   g05764(.A1(new_n6744_), .A2(new_n6757_), .B(new_n6766_), .ZN(new_n6767_));
  NOR2_X1    g05765(.A1(new_n6201_), .A2(new_n6194_), .ZN(new_n6768_));
  INV_X1     g05766(.I(new_n6757_), .ZN(new_n6769_));
  NOR3_X1    g05767(.A1(new_n6764_), .A2(new_n6748_), .A3(new_n6762_), .ZN(new_n6770_));
  NOR2_X1    g05768(.A1(new_n6748_), .A2(new_n6762_), .ZN(new_n6771_));
  NOR2_X1    g05769(.A1(new_n6771_), .A2(new_n6760_), .ZN(new_n6772_));
  NOR2_X1    g05770(.A1(new_n6772_), .A2(new_n6770_), .ZN(new_n6773_));
  NOR3_X1    g05771(.A1(new_n6768_), .A2(new_n6769_), .A3(new_n6773_), .ZN(new_n6774_));
  NOR2_X1    g05772(.A1(new_n6774_), .A2(new_n6767_), .ZN(new_n6775_));
  NOR3_X1    g05773(.A1(new_n6148_), .A2(new_n6142_), .A3(new_n6027_), .ZN(new_n6776_));
  NAND2_X1   g05774(.A1(new_n6146_), .A2(new_n6034_), .ZN(new_n6777_));
  AOI22_X1   g05775(.A1(new_n6152_), .A2(new_n6043_), .B1(new_n6777_), .B2(new_n6148_), .ZN(new_n6778_));
  NAND2_X1   g05776(.A1(new_n6135_), .A2(new_n6132_), .ZN(new_n6779_));
  INV_X1     g05777(.I(new_n6779_), .ZN(new_n6780_));
  NAND4_X1   g05778(.A1(new_n6133_), .A2(new_n6131_), .A3(new_n6056_), .A4(new_n6069_), .ZN(new_n6781_));
  AOI21_X1   g05779(.A1(new_n6130_), .A2(new_n6781_), .B(new_n6780_), .ZN(new_n6782_));
  OAI21_X1   g05780(.A1(new_n6776_), .A2(new_n6778_), .B(new_n6782_), .ZN(new_n6783_));
  NOR3_X1    g05781(.A1(new_n6782_), .A2(new_n6778_), .A3(new_n6776_), .ZN(new_n6784_));
  INV_X1     g05782(.I(new_n6784_), .ZN(new_n6785_));
  NAND2_X1   g05783(.A1(new_n6785_), .A2(new_n6783_), .ZN(new_n6786_));
  NOR2_X1    g05784(.A1(new_n6164_), .A2(new_n6157_), .ZN(new_n6787_));
  OAI21_X1   g05785(.A1(new_n6787_), .A2(new_n6162_), .B(new_n6786_), .ZN(new_n6788_));
  NOR2_X1    g05786(.A1(new_n6778_), .A2(new_n6776_), .ZN(new_n6789_));
  INV_X1     g05787(.I(new_n6782_), .ZN(new_n6790_));
  NOR2_X1    g05788(.A1(new_n6789_), .A2(new_n6790_), .ZN(new_n6791_));
  NOR2_X1    g05789(.A1(new_n6791_), .A2(new_n6784_), .ZN(new_n6792_));
  NAND2_X1   g05790(.A1(new_n6129_), .A2(new_n6165_), .ZN(new_n6793_));
  NAND3_X1   g05791(.A1(new_n6793_), .A2(new_n6792_), .A3(new_n6166_), .ZN(new_n6794_));
  NAND2_X1   g05792(.A1(new_n6788_), .A2(new_n6794_), .ZN(new_n6795_));
  NAND2_X1   g05793(.A1(new_n6795_), .A2(new_n6775_), .ZN(new_n6796_));
  OAI21_X1   g05794(.A1(new_n6768_), .A2(new_n6769_), .B(new_n6773_), .ZN(new_n6797_));
  NAND3_X1   g05795(.A1(new_n6744_), .A2(new_n6766_), .A3(new_n6757_), .ZN(new_n6798_));
  NAND2_X1   g05796(.A1(new_n6797_), .A2(new_n6798_), .ZN(new_n6799_));
  NAND3_X1   g05797(.A1(new_n6799_), .A2(new_n6788_), .A3(new_n6794_), .ZN(new_n6800_));
  AOI21_X1   g05798(.A1(new_n6796_), .A2(new_n6800_), .B(new_n6742_), .ZN(new_n6801_));
  AOI21_X1   g05799(.A1(new_n6212_), .A2(new_n6214_), .B(new_n6205_), .ZN(new_n6802_));
  AOI21_X1   g05800(.A1(new_n6793_), .A2(new_n6166_), .B(new_n6792_), .ZN(new_n6803_));
  NOR3_X1    g05801(.A1(new_n6786_), .A2(new_n6787_), .A3(new_n6162_), .ZN(new_n6804_));
  NOR2_X1    g05802(.A1(new_n6803_), .A2(new_n6804_), .ZN(new_n6805_));
  NOR2_X1    g05803(.A1(new_n6805_), .A2(new_n6799_), .ZN(new_n6806_));
  NOR3_X1    g05804(.A1(new_n6775_), .A2(new_n6803_), .A3(new_n6804_), .ZN(new_n6807_));
  NOR3_X1    g05805(.A1(new_n6806_), .A2(new_n6807_), .A3(new_n6802_), .ZN(new_n6808_));
  NOR4_X1    g05806(.A1(new_n6737_), .A2(new_n6741_), .A3(new_n6801_), .A4(new_n6808_), .ZN(new_n6809_));
  OAI21_X1   g05807(.A1(new_n6739_), .A2(new_n6740_), .B(new_n6738_), .ZN(new_n6810_));
  NAND3_X1   g05808(.A1(new_n6675_), .A2(new_n6736_), .A3(new_n6729_), .ZN(new_n6811_));
  OAI21_X1   g05809(.A1(new_n6806_), .A2(new_n6807_), .B(new_n6802_), .ZN(new_n6812_));
  NAND3_X1   g05810(.A1(new_n6796_), .A2(new_n6742_), .A3(new_n6800_), .ZN(new_n6813_));
  AOI22_X1   g05811(.A1(new_n6810_), .A2(new_n6811_), .B1(new_n6812_), .B2(new_n6813_), .ZN(new_n6814_));
  NOR3_X1    g05812(.A1(new_n6674_), .A2(new_n6809_), .A3(new_n6814_), .ZN(new_n6815_));
  OAI21_X1   g05813(.A1(new_n6127_), .A2(new_n6319_), .B(new_n6322_), .ZN(new_n6816_));
  NAND4_X1   g05814(.A1(new_n6810_), .A2(new_n6812_), .A3(new_n6811_), .A4(new_n6813_), .ZN(new_n6817_));
  OAI22_X1   g05815(.A1(new_n6737_), .A2(new_n6741_), .B1(new_n6801_), .B2(new_n6808_), .ZN(new_n6818_));
  AOI21_X1   g05816(.A1(new_n6818_), .A2(new_n6817_), .B(new_n6816_), .ZN(new_n6819_));
  NOR4_X1    g05817(.A1(new_n6669_), .A2(new_n6673_), .A3(new_n6815_), .A4(new_n6819_), .ZN(new_n6820_));
  NAND3_X1   g05818(.A1(new_n6672_), .A2(new_n6671_), .A3(new_n6670_), .ZN(new_n6821_));
  OAI21_X1   g05819(.A1(new_n6663_), .A2(new_n6668_), .B(new_n6526_), .ZN(new_n6822_));
  NAND3_X1   g05820(.A1(new_n6818_), .A2(new_n6817_), .A3(new_n6816_), .ZN(new_n6823_));
  OAI21_X1   g05821(.A1(new_n6809_), .A2(new_n6814_), .B(new_n6674_), .ZN(new_n6824_));
  AOI22_X1   g05822(.A1(new_n6821_), .A2(new_n6822_), .B1(new_n6824_), .B2(new_n6823_), .ZN(new_n6825_));
  NOR3_X1    g05823(.A1(new_n6820_), .A2(new_n6825_), .A3(new_n6525_), .ZN(new_n6826_));
  NOR3_X1    g05824(.A1(new_n5657_), .A2(new_n5658_), .A3(new_n5659_), .ZN(new_n6827_));
  AOI21_X1   g05825(.A1(new_n5654_), .A2(new_n5649_), .B(new_n5655_), .ZN(new_n6828_));
  NOR3_X1    g05826(.A1(new_n6121_), .A2(new_n6122_), .A3(new_n6120_), .ZN(new_n6829_));
  AOI21_X1   g05827(.A1(new_n6118_), .A2(new_n6113_), .B(new_n5661_), .ZN(new_n6830_));
  NOR4_X1    g05828(.A1(new_n6827_), .A2(new_n6828_), .A3(new_n6829_), .A4(new_n6830_), .ZN(new_n6831_));
  OAI22_X1   g05829(.A1(new_n6827_), .A2(new_n6828_), .B1(new_n6829_), .B2(new_n6830_), .ZN(new_n6832_));
  AOI21_X1   g05830(.A1(new_n5193_), .A2(new_n6832_), .B(new_n6831_), .ZN(new_n6833_));
  NAND3_X1   g05831(.A1(new_n6323_), .A2(new_n6322_), .A3(new_n6321_), .ZN(new_n6834_));
  OAI21_X1   g05832(.A1(new_n6314_), .A2(new_n6319_), .B(new_n6127_), .ZN(new_n6835_));
  NAND3_X1   g05833(.A1(new_n6521_), .A2(new_n6520_), .A3(new_n6519_), .ZN(new_n6836_));
  OAI21_X1   g05834(.A1(new_n6512_), .A2(new_n6517_), .B(new_n6325_), .ZN(new_n6837_));
  NAND4_X1   g05835(.A1(new_n6834_), .A2(new_n6835_), .A3(new_n6837_), .A4(new_n6836_), .ZN(new_n6838_));
  AOI22_X1   g05836(.A1(new_n6836_), .A2(new_n6837_), .B1(new_n6835_), .B2(new_n6834_), .ZN(new_n6839_));
  OAI21_X1   g05837(.A1(new_n6833_), .A2(new_n6839_), .B(new_n6838_), .ZN(new_n6840_));
  NAND4_X1   g05838(.A1(new_n6822_), .A2(new_n6824_), .A3(new_n6821_), .A4(new_n6823_), .ZN(new_n6841_));
  OAI22_X1   g05839(.A1(new_n6669_), .A2(new_n6673_), .B1(new_n6815_), .B2(new_n6819_), .ZN(new_n6842_));
  AOI21_X1   g05840(.A1(new_n6842_), .A2(new_n6841_), .B(new_n6840_), .ZN(new_n6843_));
  NOR2_X1    g05841(.A1(new_n6826_), .A2(new_n6843_), .ZN(new_n6844_));
  INV_X1     g05842(.I(\A[957] ), .ZN(new_n6845_));
  NOR2_X1    g05843(.A1(new_n6845_), .A2(\A[956] ), .ZN(new_n6846_));
  INV_X1     g05844(.I(\A[956] ), .ZN(new_n6847_));
  NOR2_X1    g05845(.A1(new_n6847_), .A2(\A[957] ), .ZN(new_n6848_));
  OAI21_X1   g05846(.A1(new_n6846_), .A2(new_n6848_), .B(\A[955] ), .ZN(new_n6849_));
  INV_X1     g05847(.I(\A[955] ), .ZN(new_n6850_));
  NOR2_X1    g05848(.A1(new_n6847_), .A2(new_n6845_), .ZN(new_n6851_));
  NOR2_X1    g05849(.A1(\A[956] ), .A2(\A[957] ), .ZN(new_n6852_));
  OAI21_X1   g05850(.A1(new_n6851_), .A2(new_n6852_), .B(new_n6850_), .ZN(new_n6853_));
  INV_X1     g05851(.I(\A[960] ), .ZN(new_n6854_));
  NOR2_X1    g05852(.A1(new_n6854_), .A2(\A[959] ), .ZN(new_n6855_));
  INV_X1     g05853(.I(\A[959] ), .ZN(new_n6856_));
  NOR2_X1    g05854(.A1(new_n6856_), .A2(\A[960] ), .ZN(new_n6857_));
  OAI21_X1   g05855(.A1(new_n6855_), .A2(new_n6857_), .B(\A[958] ), .ZN(new_n6858_));
  INV_X1     g05856(.I(\A[958] ), .ZN(new_n6859_));
  NAND2_X1   g05857(.A1(\A[959] ), .A2(\A[960] ), .ZN(new_n6860_));
  INV_X1     g05858(.I(new_n6860_), .ZN(new_n6861_));
  NOR2_X1    g05859(.A1(\A[959] ), .A2(\A[960] ), .ZN(new_n6862_));
  OAI21_X1   g05860(.A1(new_n6861_), .A2(new_n6862_), .B(new_n6859_), .ZN(new_n6863_));
  NAND4_X1   g05861(.A1(new_n6849_), .A2(new_n6853_), .A3(new_n6858_), .A4(new_n6863_), .ZN(new_n6864_));
  NAND2_X1   g05862(.A1(new_n6853_), .A2(new_n6849_), .ZN(new_n6865_));
  NAND2_X1   g05863(.A1(new_n6858_), .A2(new_n6863_), .ZN(new_n6866_));
  NAND2_X1   g05864(.A1(new_n6865_), .A2(new_n6866_), .ZN(new_n6867_));
  NAND2_X1   g05865(.A1(new_n6867_), .A2(new_n6864_), .ZN(new_n6868_));
  INV_X1     g05866(.I(\A[961] ), .ZN(new_n6869_));
  INV_X1     g05867(.I(\A[962] ), .ZN(new_n6870_));
  NAND2_X1   g05868(.A1(new_n6870_), .A2(\A[963] ), .ZN(new_n6871_));
  INV_X1     g05869(.I(\A[963] ), .ZN(new_n6872_));
  NAND2_X1   g05870(.A1(new_n6872_), .A2(\A[962] ), .ZN(new_n6873_));
  AOI21_X1   g05871(.A1(new_n6871_), .A2(new_n6873_), .B(new_n6869_), .ZN(new_n6874_));
  NAND2_X1   g05872(.A1(\A[962] ), .A2(\A[963] ), .ZN(new_n6875_));
  NOR2_X1    g05873(.A1(\A[962] ), .A2(\A[963] ), .ZN(new_n6876_));
  INV_X1     g05874(.I(new_n6876_), .ZN(new_n6877_));
  AOI21_X1   g05875(.A1(new_n6877_), .A2(new_n6875_), .B(\A[961] ), .ZN(new_n6878_));
  NOR2_X1    g05876(.A1(new_n6878_), .A2(new_n6874_), .ZN(new_n6879_));
  INV_X1     g05877(.I(\A[966] ), .ZN(new_n6880_));
  NOR2_X1    g05878(.A1(new_n6880_), .A2(\A[965] ), .ZN(new_n6881_));
  INV_X1     g05879(.I(\A[965] ), .ZN(new_n6882_));
  NOR2_X1    g05880(.A1(new_n6882_), .A2(\A[966] ), .ZN(new_n6883_));
  OAI21_X1   g05881(.A1(new_n6881_), .A2(new_n6883_), .B(\A[964] ), .ZN(new_n6884_));
  INV_X1     g05882(.I(\A[964] ), .ZN(new_n6885_));
  NAND2_X1   g05883(.A1(\A[965] ), .A2(\A[966] ), .ZN(new_n6886_));
  INV_X1     g05884(.I(new_n6886_), .ZN(new_n6887_));
  NOR2_X1    g05885(.A1(\A[965] ), .A2(\A[966] ), .ZN(new_n6888_));
  OAI21_X1   g05886(.A1(new_n6887_), .A2(new_n6888_), .B(new_n6885_), .ZN(new_n6889_));
  NAND2_X1   g05887(.A1(new_n6884_), .A2(new_n6889_), .ZN(new_n6890_));
  XOR2_X1    g05888(.A1(new_n6879_), .A2(new_n6890_), .Z(new_n6891_));
  NOR2_X1    g05889(.A1(new_n6891_), .A2(new_n6868_), .ZN(new_n6892_));
  NAND2_X1   g05890(.A1(new_n6879_), .A2(new_n6890_), .ZN(new_n6893_));
  NOR2_X1    g05891(.A1(new_n6872_), .A2(\A[962] ), .ZN(new_n6894_));
  NOR2_X1    g05892(.A1(new_n6870_), .A2(\A[963] ), .ZN(new_n6895_));
  OAI21_X1   g05893(.A1(new_n6894_), .A2(new_n6895_), .B(\A[961] ), .ZN(new_n6896_));
  INV_X1     g05894(.I(new_n6875_), .ZN(new_n6897_));
  OAI21_X1   g05895(.A1(new_n6897_), .A2(new_n6876_), .B(new_n6869_), .ZN(new_n6898_));
  NAND2_X1   g05896(.A1(new_n6896_), .A2(new_n6898_), .ZN(new_n6899_));
  NAND3_X1   g05897(.A1(new_n6899_), .A2(new_n6884_), .A3(new_n6889_), .ZN(new_n6900_));
  NAND2_X1   g05898(.A1(new_n6893_), .A2(new_n6900_), .ZN(new_n6901_));
  AOI21_X1   g05899(.A1(new_n6859_), .A2(new_n6860_), .B(new_n6862_), .ZN(new_n6902_));
  INV_X1     g05900(.I(new_n6852_), .ZN(new_n6903_));
  OAI21_X1   g05901(.A1(\A[955] ), .A2(new_n6851_), .B(new_n6903_), .ZN(new_n6904_));
  INV_X1     g05902(.I(new_n6904_), .ZN(new_n6905_));
  AOI21_X1   g05903(.A1(new_n6864_), .A2(new_n6867_), .B(new_n6901_), .ZN(new_n6906_));
  NOR2_X1    g05904(.A1(new_n6906_), .A2(new_n6892_), .ZN(new_n6907_));
  INV_X1     g05905(.I(\A[945] ), .ZN(new_n6908_));
  NOR2_X1    g05906(.A1(new_n6908_), .A2(\A[944] ), .ZN(new_n6909_));
  INV_X1     g05907(.I(\A[944] ), .ZN(new_n6910_));
  NOR2_X1    g05908(.A1(new_n6910_), .A2(\A[945] ), .ZN(new_n6911_));
  OAI21_X1   g05909(.A1(new_n6909_), .A2(new_n6911_), .B(\A[943] ), .ZN(new_n6912_));
  INV_X1     g05910(.I(\A[943] ), .ZN(new_n6913_));
  NAND2_X1   g05911(.A1(\A[944] ), .A2(\A[945] ), .ZN(new_n6914_));
  INV_X1     g05912(.I(new_n6914_), .ZN(new_n6915_));
  NOR2_X1    g05913(.A1(\A[944] ), .A2(\A[945] ), .ZN(new_n6916_));
  OAI21_X1   g05914(.A1(new_n6915_), .A2(new_n6916_), .B(new_n6913_), .ZN(new_n6917_));
  INV_X1     g05915(.I(\A[948] ), .ZN(new_n6918_));
  NOR2_X1    g05916(.A1(new_n6918_), .A2(\A[947] ), .ZN(new_n6919_));
  INV_X1     g05917(.I(\A[947] ), .ZN(new_n6920_));
  NOR2_X1    g05918(.A1(new_n6920_), .A2(\A[948] ), .ZN(new_n6921_));
  OAI21_X1   g05919(.A1(new_n6919_), .A2(new_n6921_), .B(\A[946] ), .ZN(new_n6922_));
  INV_X1     g05920(.I(\A[946] ), .ZN(new_n6923_));
  NAND2_X1   g05921(.A1(\A[947] ), .A2(\A[948] ), .ZN(new_n6924_));
  INV_X1     g05922(.I(new_n6924_), .ZN(new_n6925_));
  NOR2_X1    g05923(.A1(\A[947] ), .A2(\A[948] ), .ZN(new_n6926_));
  OAI21_X1   g05924(.A1(new_n6925_), .A2(new_n6926_), .B(new_n6923_), .ZN(new_n6927_));
  NAND4_X1   g05925(.A1(new_n6912_), .A2(new_n6917_), .A3(new_n6922_), .A4(new_n6927_), .ZN(new_n6928_));
  AOI22_X1   g05926(.A1(new_n6912_), .A2(new_n6917_), .B1(new_n6922_), .B2(new_n6927_), .ZN(new_n6929_));
  INV_X1     g05927(.I(new_n6929_), .ZN(new_n6930_));
  INV_X1     g05928(.I(\A[951] ), .ZN(new_n6931_));
  NOR2_X1    g05929(.A1(new_n6931_), .A2(\A[950] ), .ZN(new_n6932_));
  INV_X1     g05930(.I(\A[950] ), .ZN(new_n6933_));
  NOR2_X1    g05931(.A1(new_n6933_), .A2(\A[951] ), .ZN(new_n6934_));
  OAI21_X1   g05932(.A1(new_n6932_), .A2(new_n6934_), .B(\A[949] ), .ZN(new_n6935_));
  INV_X1     g05933(.I(\A[949] ), .ZN(new_n6936_));
  NAND2_X1   g05934(.A1(\A[950] ), .A2(\A[951] ), .ZN(new_n6937_));
  INV_X1     g05935(.I(new_n6937_), .ZN(new_n6938_));
  NOR2_X1    g05936(.A1(\A[950] ), .A2(\A[951] ), .ZN(new_n6939_));
  OAI21_X1   g05937(.A1(new_n6938_), .A2(new_n6939_), .B(new_n6936_), .ZN(new_n6940_));
  NAND2_X1   g05938(.A1(new_n6935_), .A2(new_n6940_), .ZN(new_n6941_));
  INV_X1     g05939(.I(\A[954] ), .ZN(new_n6942_));
  NOR2_X1    g05940(.A1(new_n6942_), .A2(\A[953] ), .ZN(new_n6943_));
  INV_X1     g05941(.I(\A[953] ), .ZN(new_n6944_));
  NOR2_X1    g05942(.A1(new_n6944_), .A2(\A[954] ), .ZN(new_n6945_));
  OAI21_X1   g05943(.A1(new_n6943_), .A2(new_n6945_), .B(\A[952] ), .ZN(new_n6946_));
  INV_X1     g05944(.I(\A[952] ), .ZN(new_n6947_));
  NOR2_X1    g05945(.A1(new_n6944_), .A2(new_n6942_), .ZN(new_n6948_));
  NOR2_X1    g05946(.A1(\A[953] ), .A2(\A[954] ), .ZN(new_n6949_));
  OAI21_X1   g05947(.A1(new_n6948_), .A2(new_n6949_), .B(new_n6947_), .ZN(new_n6950_));
  NAND2_X1   g05948(.A1(new_n6950_), .A2(new_n6946_), .ZN(new_n6951_));
  XOR2_X1    g05949(.A1(new_n6951_), .A2(new_n6941_), .Z(new_n6952_));
  NAND3_X1   g05950(.A1(new_n6952_), .A2(new_n6928_), .A3(new_n6930_), .ZN(new_n6953_));
  NAND2_X1   g05951(.A1(new_n6930_), .A2(new_n6928_), .ZN(new_n6954_));
  AOI21_X1   g05952(.A1(new_n6946_), .A2(new_n6950_), .B(new_n6941_), .ZN(new_n6955_));
  NAND2_X1   g05953(.A1(new_n6933_), .A2(\A[951] ), .ZN(new_n6956_));
  NAND2_X1   g05954(.A1(new_n6931_), .A2(\A[950] ), .ZN(new_n6957_));
  AOI21_X1   g05955(.A1(new_n6956_), .A2(new_n6957_), .B(new_n6936_), .ZN(new_n6958_));
  INV_X1     g05956(.I(new_n6939_), .ZN(new_n6959_));
  AOI21_X1   g05957(.A1(new_n6959_), .A2(new_n6937_), .B(\A[949] ), .ZN(new_n6960_));
  NOR2_X1    g05958(.A1(new_n6960_), .A2(new_n6958_), .ZN(new_n6961_));
  NOR2_X1    g05959(.A1(new_n6961_), .A2(new_n6951_), .ZN(new_n6962_));
  NOR2_X1    g05960(.A1(new_n6955_), .A2(new_n6962_), .ZN(new_n6963_));
  AOI21_X1   g05961(.A1(new_n6923_), .A2(new_n6924_), .B(new_n6926_), .ZN(new_n6964_));
  INV_X1     g05962(.I(new_n6964_), .ZN(new_n6965_));
  AOI21_X1   g05963(.A1(new_n6913_), .A2(new_n6914_), .B(new_n6916_), .ZN(new_n6966_));
  INV_X1     g05964(.I(new_n6966_), .ZN(new_n6967_));
  NOR3_X1    g05965(.A1(new_n6928_), .A2(new_n6965_), .A3(new_n6967_), .ZN(new_n6968_));
  OAI21_X1   g05966(.A1(new_n6954_), .A2(new_n6968_), .B(new_n6963_), .ZN(new_n6969_));
  NAND2_X1   g05967(.A1(new_n6969_), .A2(new_n6953_), .ZN(new_n6970_));
  XNOR2_X1   g05968(.A1(new_n6970_), .A2(new_n6907_), .ZN(new_n6971_));
  INV_X1     g05969(.I(\A[975] ), .ZN(new_n6972_));
  NOR2_X1    g05970(.A1(new_n6972_), .A2(\A[974] ), .ZN(new_n6973_));
  INV_X1     g05971(.I(\A[974] ), .ZN(new_n6974_));
  NOR2_X1    g05972(.A1(new_n6974_), .A2(\A[975] ), .ZN(new_n6975_));
  OAI21_X1   g05973(.A1(new_n6973_), .A2(new_n6975_), .B(\A[973] ), .ZN(new_n6976_));
  INV_X1     g05974(.I(\A[973] ), .ZN(new_n6977_));
  NOR2_X1    g05975(.A1(\A[974] ), .A2(\A[975] ), .ZN(new_n6978_));
  NAND2_X1   g05976(.A1(\A[974] ), .A2(\A[975] ), .ZN(new_n6979_));
  INV_X1     g05977(.I(new_n6979_), .ZN(new_n6980_));
  OAI21_X1   g05978(.A1(new_n6980_), .A2(new_n6978_), .B(new_n6977_), .ZN(new_n6981_));
  NAND2_X1   g05979(.A1(new_n6976_), .A2(new_n6981_), .ZN(new_n6982_));
  INV_X1     g05980(.I(\A[978] ), .ZN(new_n6983_));
  NOR2_X1    g05981(.A1(new_n6983_), .A2(\A[977] ), .ZN(new_n6984_));
  INV_X1     g05982(.I(\A[977] ), .ZN(new_n6985_));
  NOR2_X1    g05983(.A1(new_n6985_), .A2(\A[978] ), .ZN(new_n6986_));
  OAI21_X1   g05984(.A1(new_n6984_), .A2(new_n6986_), .B(\A[976] ), .ZN(new_n6987_));
  INV_X1     g05985(.I(\A[976] ), .ZN(new_n6988_));
  NOR2_X1    g05986(.A1(\A[977] ), .A2(\A[978] ), .ZN(new_n6989_));
  NAND2_X1   g05987(.A1(\A[977] ), .A2(\A[978] ), .ZN(new_n6990_));
  INV_X1     g05988(.I(new_n6990_), .ZN(new_n6991_));
  OAI21_X1   g05989(.A1(new_n6991_), .A2(new_n6989_), .B(new_n6988_), .ZN(new_n6992_));
  NAND2_X1   g05990(.A1(new_n6987_), .A2(new_n6992_), .ZN(new_n6993_));
  NOR2_X1    g05991(.A1(new_n6982_), .A2(new_n6993_), .ZN(new_n6994_));
  NAND2_X1   g05992(.A1(new_n6974_), .A2(\A[975] ), .ZN(new_n6995_));
  NAND2_X1   g05993(.A1(new_n6972_), .A2(\A[974] ), .ZN(new_n6996_));
  AOI21_X1   g05994(.A1(new_n6995_), .A2(new_n6996_), .B(new_n6977_), .ZN(new_n6997_));
  INV_X1     g05995(.I(new_n6978_), .ZN(new_n6998_));
  AOI21_X1   g05996(.A1(new_n6998_), .A2(new_n6979_), .B(\A[973] ), .ZN(new_n6999_));
  NOR2_X1    g05997(.A1(new_n6999_), .A2(new_n6997_), .ZN(new_n7000_));
  NAND2_X1   g05998(.A1(new_n6985_), .A2(\A[978] ), .ZN(new_n7001_));
  NAND2_X1   g05999(.A1(new_n6983_), .A2(\A[977] ), .ZN(new_n7002_));
  AOI21_X1   g06000(.A1(new_n7001_), .A2(new_n7002_), .B(new_n6988_), .ZN(new_n7003_));
  INV_X1     g06001(.I(new_n6989_), .ZN(new_n7004_));
  AOI21_X1   g06002(.A1(new_n7004_), .A2(new_n6990_), .B(\A[976] ), .ZN(new_n7005_));
  NOR2_X1    g06003(.A1(new_n7005_), .A2(new_n7003_), .ZN(new_n7006_));
  NOR2_X1    g06004(.A1(new_n7000_), .A2(new_n7006_), .ZN(new_n7007_));
  INV_X1     g06005(.I(\A[967] ), .ZN(new_n7008_));
  INV_X1     g06006(.I(\A[968] ), .ZN(new_n7009_));
  NAND2_X1   g06007(.A1(new_n7009_), .A2(\A[969] ), .ZN(new_n7010_));
  INV_X1     g06008(.I(\A[969] ), .ZN(new_n7011_));
  NAND2_X1   g06009(.A1(new_n7011_), .A2(\A[968] ), .ZN(new_n7012_));
  AOI21_X1   g06010(.A1(new_n7010_), .A2(new_n7012_), .B(new_n7008_), .ZN(new_n7013_));
  NAND2_X1   g06011(.A1(\A[968] ), .A2(\A[969] ), .ZN(new_n7014_));
  NOR2_X1    g06012(.A1(\A[968] ), .A2(\A[969] ), .ZN(new_n7015_));
  INV_X1     g06013(.I(new_n7015_), .ZN(new_n7016_));
  AOI21_X1   g06014(.A1(new_n7016_), .A2(new_n7014_), .B(\A[967] ), .ZN(new_n7017_));
  INV_X1     g06015(.I(\A[970] ), .ZN(new_n7018_));
  INV_X1     g06016(.I(\A[971] ), .ZN(new_n7019_));
  NAND2_X1   g06017(.A1(new_n7019_), .A2(\A[972] ), .ZN(new_n7020_));
  INV_X1     g06018(.I(\A[972] ), .ZN(new_n7021_));
  NAND2_X1   g06019(.A1(new_n7021_), .A2(\A[971] ), .ZN(new_n7022_));
  AOI21_X1   g06020(.A1(new_n7020_), .A2(new_n7022_), .B(new_n7018_), .ZN(new_n7023_));
  NAND2_X1   g06021(.A1(\A[971] ), .A2(\A[972] ), .ZN(new_n7024_));
  NOR2_X1    g06022(.A1(\A[971] ), .A2(\A[972] ), .ZN(new_n7025_));
  INV_X1     g06023(.I(new_n7025_), .ZN(new_n7026_));
  AOI21_X1   g06024(.A1(new_n7026_), .A2(new_n7024_), .B(\A[970] ), .ZN(new_n7027_));
  NOR4_X1    g06025(.A1(new_n7013_), .A2(new_n7017_), .A3(new_n7027_), .A4(new_n7023_), .ZN(new_n7028_));
  NOR2_X1    g06026(.A1(new_n7011_), .A2(\A[968] ), .ZN(new_n7029_));
  NOR2_X1    g06027(.A1(new_n7009_), .A2(\A[969] ), .ZN(new_n7030_));
  OAI21_X1   g06028(.A1(new_n7029_), .A2(new_n7030_), .B(\A[967] ), .ZN(new_n7031_));
  INV_X1     g06029(.I(new_n7014_), .ZN(new_n7032_));
  OAI21_X1   g06030(.A1(new_n7032_), .A2(new_n7015_), .B(new_n7008_), .ZN(new_n7033_));
  NOR2_X1    g06031(.A1(new_n7021_), .A2(\A[971] ), .ZN(new_n7034_));
  NOR2_X1    g06032(.A1(new_n7019_), .A2(\A[972] ), .ZN(new_n7035_));
  OAI21_X1   g06033(.A1(new_n7034_), .A2(new_n7035_), .B(\A[970] ), .ZN(new_n7036_));
  INV_X1     g06034(.I(new_n7024_), .ZN(new_n7037_));
  OAI21_X1   g06035(.A1(new_n7037_), .A2(new_n7025_), .B(new_n7018_), .ZN(new_n7038_));
  AOI22_X1   g06036(.A1(new_n7031_), .A2(new_n7033_), .B1(new_n7036_), .B2(new_n7038_), .ZN(new_n7039_));
  NOR2_X1    g06037(.A1(new_n7039_), .A2(new_n7028_), .ZN(new_n7040_));
  OAI21_X1   g06038(.A1(new_n6994_), .A2(new_n7007_), .B(new_n7040_), .ZN(new_n7041_));
  NAND4_X1   g06039(.A1(new_n6976_), .A2(new_n6981_), .A3(new_n6987_), .A4(new_n6992_), .ZN(new_n7042_));
  NAND2_X1   g06040(.A1(new_n6982_), .A2(new_n6993_), .ZN(new_n7043_));
  NAND4_X1   g06041(.A1(new_n7031_), .A2(new_n7033_), .A3(new_n7036_), .A4(new_n7038_), .ZN(new_n7044_));
  OAI22_X1   g06042(.A1(new_n7013_), .A2(new_n7017_), .B1(new_n7027_), .B2(new_n7023_), .ZN(new_n7045_));
  NAND2_X1   g06043(.A1(new_n7045_), .A2(new_n7044_), .ZN(new_n7046_));
  NAND3_X1   g06044(.A1(new_n7046_), .A2(new_n7042_), .A3(new_n7043_), .ZN(new_n7047_));
  NAND2_X1   g06045(.A1(new_n7041_), .A2(new_n7047_), .ZN(new_n7048_));
  INV_X1     g06046(.I(\A[987] ), .ZN(new_n7049_));
  NOR2_X1    g06047(.A1(new_n7049_), .A2(\A[986] ), .ZN(new_n7050_));
  INV_X1     g06048(.I(\A[986] ), .ZN(new_n7051_));
  NOR2_X1    g06049(.A1(new_n7051_), .A2(\A[987] ), .ZN(new_n7052_));
  OAI21_X1   g06050(.A1(new_n7050_), .A2(new_n7052_), .B(\A[985] ), .ZN(new_n7053_));
  INV_X1     g06051(.I(\A[985] ), .ZN(new_n7054_));
  NOR2_X1    g06052(.A1(\A[986] ), .A2(\A[987] ), .ZN(new_n7055_));
  NAND2_X1   g06053(.A1(\A[986] ), .A2(\A[987] ), .ZN(new_n7056_));
  INV_X1     g06054(.I(new_n7056_), .ZN(new_n7057_));
  OAI21_X1   g06055(.A1(new_n7057_), .A2(new_n7055_), .B(new_n7054_), .ZN(new_n7058_));
  INV_X1     g06056(.I(\A[990] ), .ZN(new_n7059_));
  NOR2_X1    g06057(.A1(new_n7059_), .A2(\A[989] ), .ZN(new_n7060_));
  INV_X1     g06058(.I(\A[989] ), .ZN(new_n7061_));
  NOR2_X1    g06059(.A1(new_n7061_), .A2(\A[990] ), .ZN(new_n7062_));
  OAI21_X1   g06060(.A1(new_n7060_), .A2(new_n7062_), .B(\A[988] ), .ZN(new_n7063_));
  INV_X1     g06061(.I(\A[988] ), .ZN(new_n7064_));
  NOR2_X1    g06062(.A1(\A[989] ), .A2(\A[990] ), .ZN(new_n7065_));
  NAND2_X1   g06063(.A1(\A[989] ), .A2(\A[990] ), .ZN(new_n7066_));
  INV_X1     g06064(.I(new_n7066_), .ZN(new_n7067_));
  OAI21_X1   g06065(.A1(new_n7067_), .A2(new_n7065_), .B(new_n7064_), .ZN(new_n7068_));
  NAND4_X1   g06066(.A1(new_n7053_), .A2(new_n7058_), .A3(new_n7063_), .A4(new_n7068_), .ZN(new_n7069_));
  NAND2_X1   g06067(.A1(new_n7051_), .A2(\A[987] ), .ZN(new_n7070_));
  NAND2_X1   g06068(.A1(new_n7049_), .A2(\A[986] ), .ZN(new_n7071_));
  AOI21_X1   g06069(.A1(new_n7070_), .A2(new_n7071_), .B(new_n7054_), .ZN(new_n7072_));
  INV_X1     g06070(.I(new_n7055_), .ZN(new_n7073_));
  AOI21_X1   g06071(.A1(new_n7073_), .A2(new_n7056_), .B(\A[985] ), .ZN(new_n7074_));
  NAND2_X1   g06072(.A1(new_n7061_), .A2(\A[990] ), .ZN(new_n7075_));
  NAND2_X1   g06073(.A1(new_n7059_), .A2(\A[989] ), .ZN(new_n7076_));
  AOI21_X1   g06074(.A1(new_n7075_), .A2(new_n7076_), .B(new_n7064_), .ZN(new_n7077_));
  INV_X1     g06075(.I(new_n7065_), .ZN(new_n7078_));
  AOI21_X1   g06076(.A1(new_n7078_), .A2(new_n7066_), .B(\A[988] ), .ZN(new_n7079_));
  OAI22_X1   g06077(.A1(new_n7072_), .A2(new_n7074_), .B1(new_n7079_), .B2(new_n7077_), .ZN(new_n7080_));
  NAND2_X1   g06078(.A1(new_n7080_), .A2(new_n7069_), .ZN(new_n7081_));
  INV_X1     g06079(.I(\A[981] ), .ZN(new_n7082_));
  NOR2_X1    g06080(.A1(new_n7082_), .A2(\A[980] ), .ZN(new_n7083_));
  INV_X1     g06081(.I(\A[980] ), .ZN(new_n7084_));
  NOR2_X1    g06082(.A1(new_n7084_), .A2(\A[981] ), .ZN(new_n7085_));
  OAI21_X1   g06083(.A1(new_n7083_), .A2(new_n7085_), .B(\A[979] ), .ZN(new_n7086_));
  INV_X1     g06084(.I(\A[979] ), .ZN(new_n7087_));
  NAND2_X1   g06085(.A1(\A[980] ), .A2(\A[981] ), .ZN(new_n7088_));
  INV_X1     g06086(.I(new_n7088_), .ZN(new_n7089_));
  NOR2_X1    g06087(.A1(\A[980] ), .A2(\A[981] ), .ZN(new_n7090_));
  OAI21_X1   g06088(.A1(new_n7089_), .A2(new_n7090_), .B(new_n7087_), .ZN(new_n7091_));
  INV_X1     g06089(.I(\A[984] ), .ZN(new_n7092_));
  NOR2_X1    g06090(.A1(new_n7092_), .A2(\A[983] ), .ZN(new_n7093_));
  INV_X1     g06091(.I(\A[983] ), .ZN(new_n7094_));
  NOR2_X1    g06092(.A1(new_n7094_), .A2(\A[984] ), .ZN(new_n7095_));
  OAI21_X1   g06093(.A1(new_n7093_), .A2(new_n7095_), .B(\A[982] ), .ZN(new_n7096_));
  INV_X1     g06094(.I(\A[982] ), .ZN(new_n7097_));
  NAND2_X1   g06095(.A1(\A[983] ), .A2(\A[984] ), .ZN(new_n7098_));
  INV_X1     g06096(.I(new_n7098_), .ZN(new_n7099_));
  NOR2_X1    g06097(.A1(\A[983] ), .A2(\A[984] ), .ZN(new_n7100_));
  OAI21_X1   g06098(.A1(new_n7099_), .A2(new_n7100_), .B(new_n7097_), .ZN(new_n7101_));
  NAND4_X1   g06099(.A1(new_n7086_), .A2(new_n7091_), .A3(new_n7096_), .A4(new_n7101_), .ZN(new_n7102_));
  NAND2_X1   g06100(.A1(new_n7084_), .A2(\A[981] ), .ZN(new_n7103_));
  NAND2_X1   g06101(.A1(new_n7082_), .A2(\A[980] ), .ZN(new_n7104_));
  AOI21_X1   g06102(.A1(new_n7103_), .A2(new_n7104_), .B(new_n7087_), .ZN(new_n7105_));
  INV_X1     g06103(.I(new_n7090_), .ZN(new_n7106_));
  AOI21_X1   g06104(.A1(new_n7106_), .A2(new_n7088_), .B(\A[979] ), .ZN(new_n7107_));
  NAND2_X1   g06105(.A1(new_n7094_), .A2(\A[984] ), .ZN(new_n7108_));
  NAND2_X1   g06106(.A1(new_n7092_), .A2(\A[983] ), .ZN(new_n7109_));
  AOI21_X1   g06107(.A1(new_n7108_), .A2(new_n7109_), .B(new_n7097_), .ZN(new_n7110_));
  INV_X1     g06108(.I(new_n7100_), .ZN(new_n7111_));
  AOI21_X1   g06109(.A1(new_n7111_), .A2(new_n7098_), .B(\A[982] ), .ZN(new_n7112_));
  OAI22_X1   g06110(.A1(new_n7105_), .A2(new_n7107_), .B1(new_n7112_), .B2(new_n7110_), .ZN(new_n7113_));
  NAND3_X1   g06111(.A1(new_n7081_), .A2(new_n7102_), .A3(new_n7113_), .ZN(new_n7114_));
  NAND2_X1   g06112(.A1(new_n7113_), .A2(new_n7102_), .ZN(new_n7115_));
  NAND3_X1   g06113(.A1(new_n7115_), .A2(new_n7069_), .A3(new_n7080_), .ZN(new_n7116_));
  NAND2_X1   g06114(.A1(new_n7114_), .A2(new_n7116_), .ZN(new_n7117_));
  XOR2_X1    g06115(.A1(new_n7048_), .A2(new_n7117_), .Z(new_n7118_));
  NAND2_X1   g06116(.A1(new_n6971_), .A2(new_n7118_), .ZN(new_n7119_));
  INV_X1     g06117(.I(new_n7119_), .ZN(new_n7120_));
  NOR2_X1    g06118(.A1(new_n6971_), .A2(new_n7118_), .ZN(new_n7121_));
  OR2_X2     g06119(.A1(new_n7120_), .A2(new_n7121_), .Z(new_n7122_));
  INV_X1     g06120(.I(\A[61] ), .ZN(new_n7123_));
  INV_X1     g06121(.I(\A[62] ), .ZN(new_n7124_));
  NAND2_X1   g06122(.A1(new_n7124_), .A2(\A[63] ), .ZN(new_n7125_));
  INV_X1     g06123(.I(\A[63] ), .ZN(new_n7126_));
  NAND2_X1   g06124(.A1(new_n7126_), .A2(\A[62] ), .ZN(new_n7127_));
  AOI21_X1   g06125(.A1(new_n7125_), .A2(new_n7127_), .B(new_n7123_), .ZN(new_n7128_));
  NOR2_X1    g06126(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n7129_));
  INV_X1     g06127(.I(new_n7129_), .ZN(new_n7130_));
  NAND2_X1   g06128(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n7131_));
  AOI21_X1   g06129(.A1(new_n7130_), .A2(new_n7131_), .B(\A[61] ), .ZN(new_n7132_));
  NOR2_X1    g06130(.A1(new_n7132_), .A2(new_n7128_), .ZN(new_n7133_));
  INV_X1     g06131(.I(\A[66] ), .ZN(new_n7134_));
  NOR2_X1    g06132(.A1(new_n7134_), .A2(\A[65] ), .ZN(new_n7135_));
  INV_X1     g06133(.I(\A[65] ), .ZN(new_n7136_));
  NOR2_X1    g06134(.A1(new_n7136_), .A2(\A[66] ), .ZN(new_n7137_));
  OAI21_X1   g06135(.A1(new_n7135_), .A2(new_n7137_), .B(\A[64] ), .ZN(new_n7138_));
  INV_X1     g06136(.I(\A[64] ), .ZN(new_n7139_));
  NOR2_X1    g06137(.A1(\A[65] ), .A2(\A[66] ), .ZN(new_n7140_));
  NAND2_X1   g06138(.A1(\A[65] ), .A2(\A[66] ), .ZN(new_n7141_));
  INV_X1     g06139(.I(new_n7141_), .ZN(new_n7142_));
  OAI21_X1   g06140(.A1(new_n7142_), .A2(new_n7140_), .B(new_n7139_), .ZN(new_n7143_));
  NAND2_X1   g06141(.A1(new_n7138_), .A2(new_n7143_), .ZN(new_n7144_));
  NAND2_X1   g06142(.A1(new_n7133_), .A2(new_n7144_), .ZN(new_n7145_));
  NOR2_X1    g06143(.A1(new_n7126_), .A2(\A[62] ), .ZN(new_n7146_));
  NOR2_X1    g06144(.A1(new_n7124_), .A2(\A[63] ), .ZN(new_n7147_));
  OAI21_X1   g06145(.A1(new_n7146_), .A2(new_n7147_), .B(\A[61] ), .ZN(new_n7148_));
  INV_X1     g06146(.I(new_n7131_), .ZN(new_n7149_));
  OAI21_X1   g06147(.A1(new_n7149_), .A2(new_n7129_), .B(new_n7123_), .ZN(new_n7150_));
  NAND2_X1   g06148(.A1(new_n7148_), .A2(new_n7150_), .ZN(new_n7151_));
  NAND2_X1   g06149(.A1(new_n7136_), .A2(\A[66] ), .ZN(new_n7152_));
  NAND2_X1   g06150(.A1(new_n7134_), .A2(\A[65] ), .ZN(new_n7153_));
  AOI21_X1   g06151(.A1(new_n7152_), .A2(new_n7153_), .B(new_n7139_), .ZN(new_n7154_));
  INV_X1     g06152(.I(new_n7140_), .ZN(new_n7155_));
  AOI21_X1   g06153(.A1(new_n7155_), .A2(new_n7141_), .B(\A[64] ), .ZN(new_n7156_));
  NOR2_X1    g06154(.A1(new_n7156_), .A2(new_n7154_), .ZN(new_n7157_));
  NAND2_X1   g06155(.A1(new_n7157_), .A2(new_n7151_), .ZN(new_n7158_));
  INV_X1     g06156(.I(\A[55] ), .ZN(new_n7159_));
  INV_X1     g06157(.I(\A[56] ), .ZN(new_n7160_));
  NAND2_X1   g06158(.A1(new_n7160_), .A2(\A[57] ), .ZN(new_n7161_));
  INV_X1     g06159(.I(\A[57] ), .ZN(new_n7162_));
  NAND2_X1   g06160(.A1(new_n7162_), .A2(\A[56] ), .ZN(new_n7163_));
  AOI21_X1   g06161(.A1(new_n7161_), .A2(new_n7163_), .B(new_n7159_), .ZN(new_n7164_));
  NAND2_X1   g06162(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n7165_));
  NOR2_X1    g06163(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n7166_));
  INV_X1     g06164(.I(new_n7166_), .ZN(new_n7167_));
  AOI21_X1   g06165(.A1(new_n7167_), .A2(new_n7165_), .B(\A[55] ), .ZN(new_n7168_));
  NOR2_X1    g06166(.A1(new_n7168_), .A2(new_n7164_), .ZN(new_n7169_));
  INV_X1     g06167(.I(\A[60] ), .ZN(new_n7170_));
  NOR2_X1    g06168(.A1(new_n7170_), .A2(\A[59] ), .ZN(new_n7171_));
  INV_X1     g06169(.I(\A[59] ), .ZN(new_n7172_));
  NOR2_X1    g06170(.A1(new_n7172_), .A2(\A[60] ), .ZN(new_n7173_));
  OAI21_X1   g06171(.A1(new_n7171_), .A2(new_n7173_), .B(\A[58] ), .ZN(new_n7174_));
  INV_X1     g06172(.I(\A[58] ), .ZN(new_n7175_));
  NAND2_X1   g06173(.A1(\A[59] ), .A2(\A[60] ), .ZN(new_n7176_));
  INV_X1     g06174(.I(new_n7176_), .ZN(new_n7177_));
  NOR2_X1    g06175(.A1(\A[59] ), .A2(\A[60] ), .ZN(new_n7178_));
  OAI21_X1   g06176(.A1(new_n7177_), .A2(new_n7178_), .B(new_n7175_), .ZN(new_n7179_));
  NAND2_X1   g06177(.A1(new_n7174_), .A2(new_n7179_), .ZN(new_n7180_));
  NAND2_X1   g06178(.A1(new_n7169_), .A2(new_n7180_), .ZN(new_n7181_));
  NOR2_X1    g06179(.A1(new_n7162_), .A2(\A[56] ), .ZN(new_n7182_));
  NOR2_X1    g06180(.A1(new_n7160_), .A2(\A[57] ), .ZN(new_n7183_));
  OAI21_X1   g06181(.A1(new_n7182_), .A2(new_n7183_), .B(\A[55] ), .ZN(new_n7184_));
  INV_X1     g06182(.I(new_n7165_), .ZN(new_n7185_));
  OAI21_X1   g06183(.A1(new_n7185_), .A2(new_n7166_), .B(new_n7159_), .ZN(new_n7186_));
  NAND2_X1   g06184(.A1(new_n7184_), .A2(new_n7186_), .ZN(new_n7187_));
  NAND2_X1   g06185(.A1(new_n7172_), .A2(\A[60] ), .ZN(new_n7188_));
  NAND2_X1   g06186(.A1(new_n7170_), .A2(\A[59] ), .ZN(new_n7189_));
  AOI21_X1   g06187(.A1(new_n7188_), .A2(new_n7189_), .B(new_n7175_), .ZN(new_n7190_));
  INV_X1     g06188(.I(new_n7178_), .ZN(new_n7191_));
  AOI21_X1   g06189(.A1(new_n7191_), .A2(new_n7176_), .B(\A[58] ), .ZN(new_n7192_));
  NOR2_X1    g06190(.A1(new_n7192_), .A2(new_n7190_), .ZN(new_n7193_));
  NAND2_X1   g06191(.A1(new_n7193_), .A2(new_n7187_), .ZN(new_n7194_));
  AOI22_X1   g06192(.A1(new_n7145_), .A2(new_n7158_), .B1(new_n7181_), .B2(new_n7194_), .ZN(new_n7195_));
  NOR2_X1    g06193(.A1(new_n7157_), .A2(new_n7151_), .ZN(new_n7196_));
  NOR2_X1    g06194(.A1(new_n7133_), .A2(new_n7144_), .ZN(new_n7197_));
  NOR2_X1    g06195(.A1(new_n7193_), .A2(new_n7187_), .ZN(new_n7198_));
  NOR2_X1    g06196(.A1(new_n7169_), .A2(new_n7180_), .ZN(new_n7199_));
  NOR4_X1    g06197(.A1(new_n7196_), .A2(new_n7197_), .A3(new_n7198_), .A4(new_n7199_), .ZN(new_n7200_));
  INV_X1     g06198(.I(\A[73] ), .ZN(new_n7201_));
  INV_X1     g06199(.I(\A[74] ), .ZN(new_n7202_));
  NAND2_X1   g06200(.A1(new_n7202_), .A2(\A[75] ), .ZN(new_n7203_));
  INV_X1     g06201(.I(\A[75] ), .ZN(new_n7204_));
  NAND2_X1   g06202(.A1(new_n7204_), .A2(\A[74] ), .ZN(new_n7205_));
  AOI21_X1   g06203(.A1(new_n7203_), .A2(new_n7205_), .B(new_n7201_), .ZN(new_n7206_));
  NOR2_X1    g06204(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n7207_));
  INV_X1     g06205(.I(new_n7207_), .ZN(new_n7208_));
  NAND2_X1   g06206(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n7209_));
  AOI21_X1   g06207(.A1(new_n7208_), .A2(new_n7209_), .B(\A[73] ), .ZN(new_n7210_));
  NOR2_X1    g06208(.A1(new_n7210_), .A2(new_n7206_), .ZN(new_n7211_));
  INV_X1     g06209(.I(\A[78] ), .ZN(new_n7212_));
  NOR2_X1    g06210(.A1(new_n7212_), .A2(\A[77] ), .ZN(new_n7213_));
  INV_X1     g06211(.I(\A[77] ), .ZN(new_n7214_));
  NOR2_X1    g06212(.A1(new_n7214_), .A2(\A[78] ), .ZN(new_n7215_));
  OAI21_X1   g06213(.A1(new_n7213_), .A2(new_n7215_), .B(\A[76] ), .ZN(new_n7216_));
  INV_X1     g06214(.I(\A[76] ), .ZN(new_n7217_));
  NOR2_X1    g06215(.A1(\A[77] ), .A2(\A[78] ), .ZN(new_n7218_));
  AND2_X2    g06216(.A1(\A[77] ), .A2(\A[78] ), .Z(new_n7219_));
  OAI21_X1   g06217(.A1(new_n7219_), .A2(new_n7218_), .B(new_n7217_), .ZN(new_n7220_));
  NAND2_X1   g06218(.A1(new_n7216_), .A2(new_n7220_), .ZN(new_n7221_));
  NAND2_X1   g06219(.A1(new_n7211_), .A2(new_n7221_), .ZN(new_n7222_));
  NOR2_X1    g06220(.A1(new_n7204_), .A2(\A[74] ), .ZN(new_n7223_));
  NOR2_X1    g06221(.A1(new_n7202_), .A2(\A[75] ), .ZN(new_n7224_));
  OAI21_X1   g06222(.A1(new_n7223_), .A2(new_n7224_), .B(\A[73] ), .ZN(new_n7225_));
  INV_X1     g06223(.I(new_n7209_), .ZN(new_n7226_));
  OAI21_X1   g06224(.A1(new_n7226_), .A2(new_n7207_), .B(new_n7201_), .ZN(new_n7227_));
  NAND2_X1   g06225(.A1(new_n7225_), .A2(new_n7227_), .ZN(new_n7228_));
  NAND2_X1   g06226(.A1(new_n7214_), .A2(\A[78] ), .ZN(new_n7229_));
  NAND2_X1   g06227(.A1(new_n7212_), .A2(\A[77] ), .ZN(new_n7230_));
  AOI21_X1   g06228(.A1(new_n7229_), .A2(new_n7230_), .B(new_n7217_), .ZN(new_n7231_));
  INV_X1     g06229(.I(new_n7218_), .ZN(new_n7232_));
  NAND2_X1   g06230(.A1(\A[77] ), .A2(\A[78] ), .ZN(new_n7233_));
  AOI21_X1   g06231(.A1(new_n7232_), .A2(new_n7233_), .B(\A[76] ), .ZN(new_n7234_));
  NOR2_X1    g06232(.A1(new_n7234_), .A2(new_n7231_), .ZN(new_n7235_));
  NAND2_X1   g06233(.A1(new_n7235_), .A2(new_n7228_), .ZN(new_n7236_));
  INV_X1     g06234(.I(\A[67] ), .ZN(new_n7237_));
  INV_X1     g06235(.I(\A[68] ), .ZN(new_n7238_));
  NAND2_X1   g06236(.A1(new_n7238_), .A2(\A[69] ), .ZN(new_n7239_));
  INV_X1     g06237(.I(\A[69] ), .ZN(new_n7240_));
  NAND2_X1   g06238(.A1(new_n7240_), .A2(\A[68] ), .ZN(new_n7241_));
  AOI21_X1   g06239(.A1(new_n7239_), .A2(new_n7241_), .B(new_n7237_), .ZN(new_n7242_));
  NAND2_X1   g06240(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n7243_));
  NOR2_X1    g06241(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n7244_));
  INV_X1     g06242(.I(new_n7244_), .ZN(new_n7245_));
  AOI21_X1   g06243(.A1(new_n7245_), .A2(new_n7243_), .B(\A[67] ), .ZN(new_n7246_));
  NOR2_X1    g06244(.A1(new_n7246_), .A2(new_n7242_), .ZN(new_n7247_));
  INV_X1     g06245(.I(\A[72] ), .ZN(new_n7248_));
  NOR2_X1    g06246(.A1(new_n7248_), .A2(\A[71] ), .ZN(new_n7249_));
  INV_X1     g06247(.I(\A[71] ), .ZN(new_n7250_));
  NOR2_X1    g06248(.A1(new_n7250_), .A2(\A[72] ), .ZN(new_n7251_));
  OAI21_X1   g06249(.A1(new_n7249_), .A2(new_n7251_), .B(\A[70] ), .ZN(new_n7252_));
  INV_X1     g06250(.I(\A[70] ), .ZN(new_n7253_));
  AND2_X2    g06251(.A1(\A[71] ), .A2(\A[72] ), .Z(new_n7254_));
  NOR2_X1    g06252(.A1(\A[71] ), .A2(\A[72] ), .ZN(new_n7255_));
  OAI21_X1   g06253(.A1(new_n7254_), .A2(new_n7255_), .B(new_n7253_), .ZN(new_n7256_));
  NAND2_X1   g06254(.A1(new_n7252_), .A2(new_n7256_), .ZN(new_n7257_));
  NAND2_X1   g06255(.A1(new_n7247_), .A2(new_n7257_), .ZN(new_n7258_));
  NOR2_X1    g06256(.A1(new_n7240_), .A2(\A[68] ), .ZN(new_n7259_));
  NOR2_X1    g06257(.A1(new_n7238_), .A2(\A[69] ), .ZN(new_n7260_));
  OAI21_X1   g06258(.A1(new_n7259_), .A2(new_n7260_), .B(\A[67] ), .ZN(new_n7261_));
  AND2_X2    g06259(.A1(\A[68] ), .A2(\A[69] ), .Z(new_n7262_));
  OAI21_X1   g06260(.A1(new_n7262_), .A2(new_n7244_), .B(new_n7237_), .ZN(new_n7263_));
  NAND2_X1   g06261(.A1(new_n7261_), .A2(new_n7263_), .ZN(new_n7264_));
  NAND2_X1   g06262(.A1(new_n7250_), .A2(\A[72] ), .ZN(new_n7265_));
  NAND2_X1   g06263(.A1(new_n7248_), .A2(\A[71] ), .ZN(new_n7266_));
  AOI21_X1   g06264(.A1(new_n7265_), .A2(new_n7266_), .B(new_n7253_), .ZN(new_n7267_));
  NAND2_X1   g06265(.A1(\A[71] ), .A2(\A[72] ), .ZN(new_n7268_));
  INV_X1     g06266(.I(new_n7255_), .ZN(new_n7269_));
  AOI21_X1   g06267(.A1(new_n7269_), .A2(new_n7268_), .B(\A[70] ), .ZN(new_n7270_));
  NOR2_X1    g06268(.A1(new_n7270_), .A2(new_n7267_), .ZN(new_n7271_));
  NAND2_X1   g06269(.A1(new_n7271_), .A2(new_n7264_), .ZN(new_n7272_));
  AOI22_X1   g06270(.A1(new_n7222_), .A2(new_n7236_), .B1(new_n7258_), .B2(new_n7272_), .ZN(new_n7273_));
  NOR2_X1    g06271(.A1(new_n7235_), .A2(new_n7228_), .ZN(new_n7274_));
  NOR2_X1    g06272(.A1(new_n7211_), .A2(new_n7221_), .ZN(new_n7275_));
  NOR2_X1    g06273(.A1(new_n7271_), .A2(new_n7264_), .ZN(new_n7276_));
  NOR2_X1    g06274(.A1(new_n7247_), .A2(new_n7257_), .ZN(new_n7277_));
  NOR4_X1    g06275(.A1(new_n7274_), .A2(new_n7275_), .A3(new_n7276_), .A4(new_n7277_), .ZN(new_n7278_));
  OAI22_X1   g06276(.A1(new_n7200_), .A2(new_n7195_), .B1(new_n7278_), .B2(new_n7273_), .ZN(new_n7279_));
  INV_X1     g06277(.I(new_n7279_), .ZN(new_n7280_));
  NOR4_X1    g06278(.A1(new_n7195_), .A2(new_n7200_), .A3(new_n7278_), .A4(new_n7273_), .ZN(new_n7281_));
  INV_X1     g06279(.I(\A[39] ), .ZN(new_n7282_));
  NOR2_X1    g06280(.A1(new_n7282_), .A2(\A[38] ), .ZN(new_n7283_));
  INV_X1     g06281(.I(\A[38] ), .ZN(new_n7284_));
  NOR2_X1    g06282(.A1(new_n7284_), .A2(\A[39] ), .ZN(new_n7285_));
  OAI21_X1   g06283(.A1(new_n7283_), .A2(new_n7285_), .B(\A[37] ), .ZN(new_n7286_));
  INV_X1     g06284(.I(\A[37] ), .ZN(new_n7287_));
  NOR2_X1    g06285(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n7288_));
  NAND2_X1   g06286(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n7289_));
  INV_X1     g06287(.I(new_n7289_), .ZN(new_n7290_));
  OAI21_X1   g06288(.A1(new_n7290_), .A2(new_n7288_), .B(new_n7287_), .ZN(new_n7291_));
  NAND2_X1   g06289(.A1(new_n7286_), .A2(new_n7291_), .ZN(new_n7292_));
  INV_X1     g06290(.I(\A[40] ), .ZN(new_n7293_));
  INV_X1     g06291(.I(\A[41] ), .ZN(new_n7294_));
  NAND2_X1   g06292(.A1(new_n7294_), .A2(\A[42] ), .ZN(new_n7295_));
  INV_X1     g06293(.I(\A[42] ), .ZN(new_n7296_));
  NAND2_X1   g06294(.A1(new_n7296_), .A2(\A[41] ), .ZN(new_n7297_));
  AOI21_X1   g06295(.A1(new_n7295_), .A2(new_n7297_), .B(new_n7293_), .ZN(new_n7298_));
  NOR2_X1    g06296(.A1(\A[41] ), .A2(\A[42] ), .ZN(new_n7299_));
  INV_X1     g06297(.I(new_n7299_), .ZN(new_n7300_));
  NAND2_X1   g06298(.A1(\A[41] ), .A2(\A[42] ), .ZN(new_n7301_));
  AOI21_X1   g06299(.A1(new_n7300_), .A2(new_n7301_), .B(\A[40] ), .ZN(new_n7302_));
  NOR2_X1    g06300(.A1(new_n7302_), .A2(new_n7298_), .ZN(new_n7303_));
  NOR2_X1    g06301(.A1(new_n7303_), .A2(new_n7292_), .ZN(new_n7304_));
  NAND2_X1   g06302(.A1(new_n7284_), .A2(\A[39] ), .ZN(new_n7305_));
  NAND2_X1   g06303(.A1(new_n7282_), .A2(\A[38] ), .ZN(new_n7306_));
  AOI21_X1   g06304(.A1(new_n7305_), .A2(new_n7306_), .B(new_n7287_), .ZN(new_n7307_));
  INV_X1     g06305(.I(new_n7288_), .ZN(new_n7308_));
  AOI21_X1   g06306(.A1(new_n7308_), .A2(new_n7289_), .B(\A[37] ), .ZN(new_n7309_));
  NOR2_X1    g06307(.A1(new_n7309_), .A2(new_n7307_), .ZN(new_n7310_));
  NOR2_X1    g06308(.A1(new_n7296_), .A2(\A[41] ), .ZN(new_n7311_));
  NOR2_X1    g06309(.A1(new_n7294_), .A2(\A[42] ), .ZN(new_n7312_));
  OAI21_X1   g06310(.A1(new_n7311_), .A2(new_n7312_), .B(\A[40] ), .ZN(new_n7313_));
  INV_X1     g06311(.I(new_n7301_), .ZN(new_n7314_));
  OAI21_X1   g06312(.A1(new_n7314_), .A2(new_n7299_), .B(new_n7293_), .ZN(new_n7315_));
  NAND2_X1   g06313(.A1(new_n7313_), .A2(new_n7315_), .ZN(new_n7316_));
  NOR2_X1    g06314(.A1(new_n7310_), .A2(new_n7316_), .ZN(new_n7317_));
  INV_X1     g06315(.I(\A[33] ), .ZN(new_n7318_));
  NOR2_X1    g06316(.A1(new_n7318_), .A2(\A[32] ), .ZN(new_n7319_));
  INV_X1     g06317(.I(\A[32] ), .ZN(new_n7320_));
  NOR2_X1    g06318(.A1(new_n7320_), .A2(\A[33] ), .ZN(new_n7321_));
  OAI21_X1   g06319(.A1(new_n7319_), .A2(new_n7321_), .B(\A[31] ), .ZN(new_n7322_));
  INV_X1     g06320(.I(\A[31] ), .ZN(new_n7323_));
  NOR2_X1    g06321(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n7324_));
  NAND2_X1   g06322(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n7325_));
  INV_X1     g06323(.I(new_n7325_), .ZN(new_n7326_));
  OAI21_X1   g06324(.A1(new_n7326_), .A2(new_n7324_), .B(new_n7323_), .ZN(new_n7327_));
  NAND2_X1   g06325(.A1(new_n7322_), .A2(new_n7327_), .ZN(new_n7328_));
  INV_X1     g06326(.I(\A[34] ), .ZN(new_n7329_));
  INV_X1     g06327(.I(\A[35] ), .ZN(new_n7330_));
  NAND2_X1   g06328(.A1(new_n7330_), .A2(\A[36] ), .ZN(new_n7331_));
  INV_X1     g06329(.I(\A[36] ), .ZN(new_n7332_));
  NAND2_X1   g06330(.A1(new_n7332_), .A2(\A[35] ), .ZN(new_n7333_));
  AOI21_X1   g06331(.A1(new_n7331_), .A2(new_n7333_), .B(new_n7329_), .ZN(new_n7334_));
  NOR2_X1    g06332(.A1(\A[35] ), .A2(\A[36] ), .ZN(new_n7335_));
  INV_X1     g06333(.I(new_n7335_), .ZN(new_n7336_));
  NAND2_X1   g06334(.A1(\A[35] ), .A2(\A[36] ), .ZN(new_n7337_));
  AOI21_X1   g06335(.A1(new_n7336_), .A2(new_n7337_), .B(\A[34] ), .ZN(new_n7338_));
  NOR2_X1    g06336(.A1(new_n7338_), .A2(new_n7334_), .ZN(new_n7339_));
  NOR2_X1    g06337(.A1(new_n7339_), .A2(new_n7328_), .ZN(new_n7340_));
  NAND2_X1   g06338(.A1(new_n7320_), .A2(\A[33] ), .ZN(new_n7341_));
  NAND2_X1   g06339(.A1(new_n7318_), .A2(\A[32] ), .ZN(new_n7342_));
  AOI21_X1   g06340(.A1(new_n7341_), .A2(new_n7342_), .B(new_n7323_), .ZN(new_n7343_));
  INV_X1     g06341(.I(new_n7324_), .ZN(new_n7344_));
  AOI21_X1   g06342(.A1(new_n7344_), .A2(new_n7325_), .B(\A[31] ), .ZN(new_n7345_));
  NOR2_X1    g06343(.A1(new_n7345_), .A2(new_n7343_), .ZN(new_n7346_));
  NOR2_X1    g06344(.A1(new_n7332_), .A2(\A[35] ), .ZN(new_n7347_));
  NOR2_X1    g06345(.A1(new_n7330_), .A2(\A[36] ), .ZN(new_n7348_));
  OAI21_X1   g06346(.A1(new_n7347_), .A2(new_n7348_), .B(\A[34] ), .ZN(new_n7349_));
  INV_X1     g06347(.I(new_n7337_), .ZN(new_n7350_));
  OAI21_X1   g06348(.A1(new_n7350_), .A2(new_n7335_), .B(new_n7329_), .ZN(new_n7351_));
  NAND2_X1   g06349(.A1(new_n7349_), .A2(new_n7351_), .ZN(new_n7352_));
  NOR2_X1    g06350(.A1(new_n7346_), .A2(new_n7352_), .ZN(new_n7353_));
  OAI22_X1   g06351(.A1(new_n7304_), .A2(new_n7317_), .B1(new_n7340_), .B2(new_n7353_), .ZN(new_n7354_));
  NOR2_X1    g06352(.A1(new_n7304_), .A2(new_n7317_), .ZN(new_n7355_));
  NOR2_X1    g06353(.A1(new_n7340_), .A2(new_n7353_), .ZN(new_n7356_));
  NAND2_X1   g06354(.A1(new_n7355_), .A2(new_n7356_), .ZN(new_n7357_));
  INV_X1     g06355(.I(\A[51] ), .ZN(new_n7358_));
  NOR2_X1    g06356(.A1(new_n7358_), .A2(\A[50] ), .ZN(new_n7359_));
  INV_X1     g06357(.I(\A[50] ), .ZN(new_n7360_));
  NOR2_X1    g06358(.A1(new_n7360_), .A2(\A[51] ), .ZN(new_n7361_));
  OAI21_X1   g06359(.A1(new_n7359_), .A2(new_n7361_), .B(\A[49] ), .ZN(new_n7362_));
  INV_X1     g06360(.I(\A[49] ), .ZN(new_n7363_));
  NOR2_X1    g06361(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n7364_));
  NAND2_X1   g06362(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n7365_));
  INV_X1     g06363(.I(new_n7365_), .ZN(new_n7366_));
  OAI21_X1   g06364(.A1(new_n7366_), .A2(new_n7364_), .B(new_n7363_), .ZN(new_n7367_));
  NAND2_X1   g06365(.A1(new_n7362_), .A2(new_n7367_), .ZN(new_n7368_));
  INV_X1     g06366(.I(\A[52] ), .ZN(new_n7369_));
  INV_X1     g06367(.I(\A[53] ), .ZN(new_n7370_));
  NAND2_X1   g06368(.A1(new_n7370_), .A2(\A[54] ), .ZN(new_n7371_));
  INV_X1     g06369(.I(\A[54] ), .ZN(new_n7372_));
  NAND2_X1   g06370(.A1(new_n7372_), .A2(\A[53] ), .ZN(new_n7373_));
  AOI21_X1   g06371(.A1(new_n7371_), .A2(new_n7373_), .B(new_n7369_), .ZN(new_n7374_));
  NOR2_X1    g06372(.A1(\A[53] ), .A2(\A[54] ), .ZN(new_n7375_));
  INV_X1     g06373(.I(new_n7375_), .ZN(new_n7376_));
  NAND2_X1   g06374(.A1(\A[53] ), .A2(\A[54] ), .ZN(new_n7377_));
  AOI21_X1   g06375(.A1(new_n7376_), .A2(new_n7377_), .B(\A[52] ), .ZN(new_n7378_));
  NOR2_X1    g06376(.A1(new_n7378_), .A2(new_n7374_), .ZN(new_n7379_));
  NOR2_X1    g06377(.A1(new_n7379_), .A2(new_n7368_), .ZN(new_n7380_));
  NAND2_X1   g06378(.A1(new_n7360_), .A2(\A[51] ), .ZN(new_n7381_));
  NAND2_X1   g06379(.A1(new_n7358_), .A2(\A[50] ), .ZN(new_n7382_));
  AOI21_X1   g06380(.A1(new_n7381_), .A2(new_n7382_), .B(new_n7363_), .ZN(new_n7383_));
  INV_X1     g06381(.I(new_n7364_), .ZN(new_n7384_));
  AOI21_X1   g06382(.A1(new_n7384_), .A2(new_n7365_), .B(\A[49] ), .ZN(new_n7385_));
  NOR2_X1    g06383(.A1(new_n7385_), .A2(new_n7383_), .ZN(new_n7386_));
  NOR2_X1    g06384(.A1(new_n7372_), .A2(\A[53] ), .ZN(new_n7387_));
  NOR2_X1    g06385(.A1(new_n7370_), .A2(\A[54] ), .ZN(new_n7388_));
  OAI21_X1   g06386(.A1(new_n7387_), .A2(new_n7388_), .B(\A[52] ), .ZN(new_n7389_));
  INV_X1     g06387(.I(new_n7377_), .ZN(new_n7390_));
  OAI21_X1   g06388(.A1(new_n7390_), .A2(new_n7375_), .B(new_n7369_), .ZN(new_n7391_));
  NAND2_X1   g06389(.A1(new_n7389_), .A2(new_n7391_), .ZN(new_n7392_));
  NOR2_X1    g06390(.A1(new_n7386_), .A2(new_n7392_), .ZN(new_n7393_));
  INV_X1     g06391(.I(\A[45] ), .ZN(new_n7394_));
  NOR2_X1    g06392(.A1(new_n7394_), .A2(\A[44] ), .ZN(new_n7395_));
  INV_X1     g06393(.I(\A[44] ), .ZN(new_n7396_));
  NOR2_X1    g06394(.A1(new_n7396_), .A2(\A[45] ), .ZN(new_n7397_));
  OAI21_X1   g06395(.A1(new_n7395_), .A2(new_n7397_), .B(\A[43] ), .ZN(new_n7398_));
  INV_X1     g06396(.I(\A[43] ), .ZN(new_n7399_));
  NOR2_X1    g06397(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n7400_));
  NAND2_X1   g06398(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n7401_));
  INV_X1     g06399(.I(new_n7401_), .ZN(new_n7402_));
  OAI21_X1   g06400(.A1(new_n7402_), .A2(new_n7400_), .B(new_n7399_), .ZN(new_n7403_));
  NAND2_X1   g06401(.A1(new_n7398_), .A2(new_n7403_), .ZN(new_n7404_));
  INV_X1     g06402(.I(\A[46] ), .ZN(new_n7405_));
  INV_X1     g06403(.I(\A[47] ), .ZN(new_n7406_));
  NAND2_X1   g06404(.A1(new_n7406_), .A2(\A[48] ), .ZN(new_n7407_));
  INV_X1     g06405(.I(\A[48] ), .ZN(new_n7408_));
  NAND2_X1   g06406(.A1(new_n7408_), .A2(\A[47] ), .ZN(new_n7409_));
  AOI21_X1   g06407(.A1(new_n7407_), .A2(new_n7409_), .B(new_n7405_), .ZN(new_n7410_));
  NOR2_X1    g06408(.A1(\A[47] ), .A2(\A[48] ), .ZN(new_n7411_));
  INV_X1     g06409(.I(new_n7411_), .ZN(new_n7412_));
  NAND2_X1   g06410(.A1(\A[47] ), .A2(\A[48] ), .ZN(new_n7413_));
  AOI21_X1   g06411(.A1(new_n7412_), .A2(new_n7413_), .B(\A[46] ), .ZN(new_n7414_));
  NOR2_X1    g06412(.A1(new_n7414_), .A2(new_n7410_), .ZN(new_n7415_));
  NOR2_X1    g06413(.A1(new_n7415_), .A2(new_n7404_), .ZN(new_n7416_));
  NAND2_X1   g06414(.A1(new_n7396_), .A2(\A[45] ), .ZN(new_n7417_));
  NAND2_X1   g06415(.A1(new_n7394_), .A2(\A[44] ), .ZN(new_n7418_));
  AOI21_X1   g06416(.A1(new_n7417_), .A2(new_n7418_), .B(new_n7399_), .ZN(new_n7419_));
  INV_X1     g06417(.I(new_n7400_), .ZN(new_n7420_));
  AOI21_X1   g06418(.A1(new_n7420_), .A2(new_n7401_), .B(\A[43] ), .ZN(new_n7421_));
  NOR2_X1    g06419(.A1(new_n7421_), .A2(new_n7419_), .ZN(new_n7422_));
  NOR2_X1    g06420(.A1(new_n7408_), .A2(\A[47] ), .ZN(new_n7423_));
  NOR2_X1    g06421(.A1(new_n7406_), .A2(\A[48] ), .ZN(new_n7424_));
  OAI21_X1   g06422(.A1(new_n7423_), .A2(new_n7424_), .B(\A[46] ), .ZN(new_n7425_));
  INV_X1     g06423(.I(new_n7413_), .ZN(new_n7426_));
  OAI21_X1   g06424(.A1(new_n7426_), .A2(new_n7411_), .B(new_n7405_), .ZN(new_n7427_));
  NAND2_X1   g06425(.A1(new_n7425_), .A2(new_n7427_), .ZN(new_n7428_));
  NOR2_X1    g06426(.A1(new_n7422_), .A2(new_n7428_), .ZN(new_n7429_));
  OAI22_X1   g06427(.A1(new_n7380_), .A2(new_n7393_), .B1(new_n7416_), .B2(new_n7429_), .ZN(new_n7430_));
  NOR4_X1    g06428(.A1(new_n7380_), .A2(new_n7393_), .A3(new_n7416_), .A4(new_n7429_), .ZN(new_n7431_));
  INV_X1     g06429(.I(new_n7431_), .ZN(new_n7432_));
  AOI22_X1   g06430(.A1(new_n7432_), .A2(new_n7430_), .B1(new_n7357_), .B2(new_n7354_), .ZN(new_n7433_));
  NAND2_X1   g06431(.A1(new_n7310_), .A2(new_n7316_), .ZN(new_n7434_));
  NAND2_X1   g06432(.A1(new_n7303_), .A2(new_n7292_), .ZN(new_n7435_));
  NAND2_X1   g06433(.A1(new_n7346_), .A2(new_n7352_), .ZN(new_n7436_));
  NAND2_X1   g06434(.A1(new_n7339_), .A2(new_n7328_), .ZN(new_n7437_));
  AOI22_X1   g06435(.A1(new_n7434_), .A2(new_n7435_), .B1(new_n7436_), .B2(new_n7437_), .ZN(new_n7438_));
  NAND2_X1   g06436(.A1(new_n7434_), .A2(new_n7435_), .ZN(new_n7439_));
  NAND2_X1   g06437(.A1(new_n7436_), .A2(new_n7437_), .ZN(new_n7440_));
  NOR2_X1    g06438(.A1(new_n7439_), .A2(new_n7440_), .ZN(new_n7441_));
  NAND2_X1   g06439(.A1(new_n7386_), .A2(new_n7392_), .ZN(new_n7442_));
  NAND2_X1   g06440(.A1(new_n7379_), .A2(new_n7368_), .ZN(new_n7443_));
  NAND2_X1   g06441(.A1(new_n7422_), .A2(new_n7428_), .ZN(new_n7444_));
  NAND2_X1   g06442(.A1(new_n7415_), .A2(new_n7404_), .ZN(new_n7445_));
  AOI22_X1   g06443(.A1(new_n7444_), .A2(new_n7445_), .B1(new_n7442_), .B2(new_n7443_), .ZN(new_n7446_));
  NOR4_X1    g06444(.A1(new_n7441_), .A2(new_n7438_), .A3(new_n7446_), .A4(new_n7431_), .ZN(new_n7447_));
  NOR4_X1    g06445(.A1(new_n7280_), .A2(new_n7433_), .A3(new_n7281_), .A4(new_n7447_), .ZN(new_n7448_));
  OR4_X2     g06446(.A1(new_n7195_), .A2(new_n7200_), .A3(new_n7273_), .A4(new_n7278_), .Z(new_n7449_));
  INV_X1     g06447(.I(new_n7433_), .ZN(new_n7450_));
  NAND4_X1   g06448(.A1(new_n7432_), .A2(new_n7357_), .A3(new_n7354_), .A4(new_n7430_), .ZN(new_n7451_));
  AOI22_X1   g06449(.A1(new_n7450_), .A2(new_n7451_), .B1(new_n7279_), .B2(new_n7449_), .ZN(new_n7452_));
  NOR2_X1    g06450(.A1(new_n7452_), .A2(new_n7448_), .ZN(new_n7453_));
  INV_X1     g06451(.I(\A[993] ), .ZN(new_n7454_));
  NOR2_X1    g06452(.A1(new_n7454_), .A2(\A[992] ), .ZN(new_n7455_));
  INV_X1     g06453(.I(\A[992] ), .ZN(new_n7456_));
  NOR2_X1    g06454(.A1(new_n7456_), .A2(\A[993] ), .ZN(new_n7457_));
  OAI21_X1   g06455(.A1(new_n7455_), .A2(new_n7457_), .B(\A[991] ), .ZN(new_n7458_));
  NOR2_X1    g06456(.A1(\A[992] ), .A2(\A[993] ), .ZN(new_n7459_));
  NOR2_X1    g06457(.A1(new_n7456_), .A2(new_n7454_), .ZN(new_n7460_));
  NOR2_X1    g06458(.A1(new_n7460_), .A2(new_n7459_), .ZN(new_n7461_));
  OAI21_X1   g06459(.A1(\A[991] ), .A2(new_n7461_), .B(new_n7458_), .ZN(new_n7462_));
  INV_X1     g06460(.I(\A[996] ), .ZN(new_n7463_));
  NOR2_X1    g06461(.A1(new_n7463_), .A2(\A[995] ), .ZN(new_n7464_));
  INV_X1     g06462(.I(\A[995] ), .ZN(new_n7465_));
  NOR2_X1    g06463(.A1(new_n7465_), .A2(\A[996] ), .ZN(new_n7466_));
  OAI21_X1   g06464(.A1(new_n7464_), .A2(new_n7466_), .B(\A[994] ), .ZN(new_n7467_));
  NOR2_X1    g06465(.A1(\A[995] ), .A2(\A[996] ), .ZN(new_n7468_));
  NOR2_X1    g06466(.A1(new_n7465_), .A2(new_n7463_), .ZN(new_n7469_));
  NOR2_X1    g06467(.A1(new_n7469_), .A2(new_n7468_), .ZN(new_n7470_));
  OAI21_X1   g06468(.A1(\A[994] ), .A2(new_n7470_), .B(new_n7467_), .ZN(new_n7471_));
  XNOR2_X1   g06469(.A1(new_n7462_), .A2(new_n7471_), .ZN(new_n7472_));
  XOR2_X1    g06470(.A1(\A[998] ), .A2(\A[999] ), .Z(new_n7473_));
  NAND2_X1   g06471(.A1(new_n7473_), .A2(\A[997] ), .ZN(new_n7474_));
  INV_X1     g06472(.I(\A[997] ), .ZN(new_n7475_));
  AND2_X2    g06473(.A1(\A[998] ), .A2(\A[999] ), .Z(new_n7476_));
  NOR2_X1    g06474(.A1(\A[998] ), .A2(\A[999] ), .ZN(new_n7477_));
  OAI21_X1   g06475(.A1(new_n7476_), .A2(new_n7477_), .B(new_n7475_), .ZN(new_n7478_));
  NAND2_X1   g06476(.A1(new_n7474_), .A2(new_n7478_), .ZN(new_n7479_));
  INV_X1     g06477(.I(\A[5] ), .ZN(new_n7480_));
  NOR2_X1    g06478(.A1(new_n7480_), .A2(\A[4] ), .ZN(new_n7481_));
  INV_X1     g06479(.I(\A[4] ), .ZN(new_n7482_));
  NOR2_X1    g06480(.A1(new_n7482_), .A2(\A[5] ), .ZN(new_n7483_));
  OAI21_X1   g06481(.A1(new_n7481_), .A2(new_n7483_), .B(\A[3] ), .ZN(new_n7484_));
  INV_X1     g06482(.I(\A[3] ), .ZN(new_n7485_));
  NAND2_X1   g06483(.A1(\A[4] ), .A2(\A[5] ), .ZN(new_n7486_));
  INV_X1     g06484(.I(new_n7486_), .ZN(new_n7487_));
  NOR2_X1    g06485(.A1(\A[4] ), .A2(\A[5] ), .ZN(new_n7488_));
  OAI21_X1   g06486(.A1(new_n7487_), .A2(new_n7488_), .B(new_n7485_), .ZN(new_n7489_));
  NAND2_X1   g06487(.A1(new_n7484_), .A2(new_n7489_), .ZN(new_n7490_));
  INV_X1     g06488(.I(\A[6] ), .ZN(new_n7491_));
  INV_X1     g06489(.I(\A[1] ), .ZN(new_n7492_));
  NAND2_X1   g06490(.A1(new_n7492_), .A2(\A[2] ), .ZN(new_n7493_));
  INV_X1     g06491(.I(\A[2] ), .ZN(new_n7494_));
  NAND2_X1   g06492(.A1(new_n7494_), .A2(\A[1] ), .ZN(new_n7495_));
  AOI21_X1   g06493(.A1(new_n7493_), .A2(new_n7495_), .B(\A[0] ), .ZN(new_n7496_));
  INV_X1     g06494(.I(\A[0] ), .ZN(new_n7497_));
  NAND2_X1   g06495(.A1(\A[1] ), .A2(\A[2] ), .ZN(new_n7498_));
  NOR2_X1    g06496(.A1(\A[1] ), .A2(\A[2] ), .ZN(new_n7499_));
  INV_X1     g06497(.I(new_n7499_), .ZN(new_n7500_));
  AOI21_X1   g06498(.A1(new_n7500_), .A2(new_n7498_), .B(new_n7497_), .ZN(new_n7501_));
  OAI21_X1   g06499(.A1(new_n7501_), .A2(new_n7496_), .B(new_n7491_), .ZN(new_n7502_));
  NOR2_X1    g06500(.A1(new_n7494_), .A2(\A[1] ), .ZN(new_n7503_));
  NOR2_X1    g06501(.A1(new_n7492_), .A2(\A[2] ), .ZN(new_n7504_));
  OAI21_X1   g06502(.A1(new_n7503_), .A2(new_n7504_), .B(new_n7497_), .ZN(new_n7505_));
  NAND3_X1   g06503(.A1(new_n7493_), .A2(new_n7495_), .A3(\A[0] ), .ZN(new_n7506_));
  NAND3_X1   g06504(.A1(new_n7505_), .A2(new_n7506_), .A3(\A[6] ), .ZN(new_n7507_));
  AOI21_X1   g06505(.A1(new_n7502_), .A2(new_n7507_), .B(new_n7490_), .ZN(new_n7508_));
  NAND2_X1   g06506(.A1(new_n7482_), .A2(\A[5] ), .ZN(new_n7509_));
  NAND2_X1   g06507(.A1(new_n7480_), .A2(\A[4] ), .ZN(new_n7510_));
  AOI21_X1   g06508(.A1(new_n7509_), .A2(new_n7510_), .B(new_n7485_), .ZN(new_n7511_));
  INV_X1     g06509(.I(new_n7488_), .ZN(new_n7512_));
  AOI21_X1   g06510(.A1(new_n7512_), .A2(new_n7486_), .B(\A[3] ), .ZN(new_n7513_));
  NOR2_X1    g06511(.A1(new_n7513_), .A2(new_n7511_), .ZN(new_n7514_));
  AND2_X2    g06512(.A1(\A[1] ), .A2(\A[2] ), .Z(new_n7515_));
  OAI21_X1   g06513(.A1(new_n7515_), .A2(new_n7499_), .B(\A[0] ), .ZN(new_n7516_));
  AOI21_X1   g06514(.A1(new_n7505_), .A2(new_n7516_), .B(\A[6] ), .ZN(new_n7517_));
  NOR3_X1    g06515(.A1(new_n7503_), .A2(new_n7504_), .A3(new_n7497_), .ZN(new_n7518_));
  NOR3_X1    g06516(.A1(new_n7496_), .A2(new_n7518_), .A3(new_n7491_), .ZN(new_n7519_));
  NOR3_X1    g06517(.A1(new_n7519_), .A2(new_n7517_), .A3(new_n7514_), .ZN(new_n7520_));
  NOR3_X1    g06518(.A1(new_n7520_), .A2(new_n7508_), .A3(new_n7479_), .ZN(new_n7521_));
  INV_X1     g06519(.I(new_n7479_), .ZN(new_n7522_));
  OAI21_X1   g06520(.A1(new_n7519_), .A2(new_n7517_), .B(new_n7514_), .ZN(new_n7523_));
  NAND3_X1   g06521(.A1(new_n7502_), .A2(new_n7507_), .A3(new_n7490_), .ZN(new_n7524_));
  AOI21_X1   g06522(.A1(new_n7523_), .A2(new_n7524_), .B(new_n7522_), .ZN(new_n7525_));
  OAI21_X1   g06523(.A1(new_n7521_), .A2(new_n7525_), .B(new_n7472_), .ZN(new_n7526_));
  NOR3_X1    g06524(.A1(new_n7472_), .A2(new_n7525_), .A3(new_n7521_), .ZN(new_n7527_));
  INV_X1     g06525(.I(new_n7527_), .ZN(new_n7528_));
  NAND2_X1   g06526(.A1(new_n7528_), .A2(new_n7526_), .ZN(new_n7529_));
  INV_X1     g06527(.I(\A[13] ), .ZN(new_n7530_));
  INV_X1     g06528(.I(\A[14] ), .ZN(new_n7531_));
  NAND2_X1   g06529(.A1(new_n7531_), .A2(\A[15] ), .ZN(new_n7532_));
  INV_X1     g06530(.I(\A[15] ), .ZN(new_n7533_));
  NAND2_X1   g06531(.A1(new_n7533_), .A2(\A[14] ), .ZN(new_n7534_));
  AOI21_X1   g06532(.A1(new_n7532_), .A2(new_n7534_), .B(new_n7530_), .ZN(new_n7535_));
  NOR2_X1    g06533(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n7536_));
  INV_X1     g06534(.I(new_n7536_), .ZN(new_n7537_));
  NAND2_X1   g06535(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n7538_));
  AOI21_X1   g06536(.A1(new_n7537_), .A2(new_n7538_), .B(\A[13] ), .ZN(new_n7539_));
  NOR2_X1    g06537(.A1(new_n7539_), .A2(new_n7535_), .ZN(new_n7540_));
  INV_X1     g06538(.I(\A[18] ), .ZN(new_n7541_));
  NOR2_X1    g06539(.A1(new_n7541_), .A2(\A[17] ), .ZN(new_n7542_));
  INV_X1     g06540(.I(\A[17] ), .ZN(new_n7543_));
  NOR2_X1    g06541(.A1(new_n7543_), .A2(\A[18] ), .ZN(new_n7544_));
  OAI21_X1   g06542(.A1(new_n7542_), .A2(new_n7544_), .B(\A[16] ), .ZN(new_n7545_));
  INV_X1     g06543(.I(\A[16] ), .ZN(new_n7546_));
  NOR2_X1    g06544(.A1(\A[17] ), .A2(\A[18] ), .ZN(new_n7547_));
  AND2_X2    g06545(.A1(\A[17] ), .A2(\A[18] ), .Z(new_n7548_));
  OAI21_X1   g06546(.A1(new_n7548_), .A2(new_n7547_), .B(new_n7546_), .ZN(new_n7549_));
  NAND2_X1   g06547(.A1(new_n7545_), .A2(new_n7549_), .ZN(new_n7550_));
  NAND2_X1   g06548(.A1(new_n7540_), .A2(new_n7550_), .ZN(new_n7551_));
  NOR2_X1    g06549(.A1(new_n7533_), .A2(\A[14] ), .ZN(new_n7552_));
  NOR2_X1    g06550(.A1(new_n7531_), .A2(\A[15] ), .ZN(new_n7553_));
  OAI21_X1   g06551(.A1(new_n7552_), .A2(new_n7553_), .B(\A[13] ), .ZN(new_n7554_));
  INV_X1     g06552(.I(new_n7538_), .ZN(new_n7555_));
  OAI21_X1   g06553(.A1(new_n7555_), .A2(new_n7536_), .B(new_n7530_), .ZN(new_n7556_));
  NAND2_X1   g06554(.A1(new_n7554_), .A2(new_n7556_), .ZN(new_n7557_));
  NAND2_X1   g06555(.A1(new_n7543_), .A2(\A[18] ), .ZN(new_n7558_));
  NAND2_X1   g06556(.A1(new_n7541_), .A2(\A[17] ), .ZN(new_n7559_));
  AOI21_X1   g06557(.A1(new_n7558_), .A2(new_n7559_), .B(new_n7546_), .ZN(new_n7560_));
  INV_X1     g06558(.I(new_n7547_), .ZN(new_n7561_));
  NAND2_X1   g06559(.A1(\A[17] ), .A2(\A[18] ), .ZN(new_n7562_));
  AOI21_X1   g06560(.A1(new_n7561_), .A2(new_n7562_), .B(\A[16] ), .ZN(new_n7563_));
  NOR2_X1    g06561(.A1(new_n7563_), .A2(new_n7560_), .ZN(new_n7564_));
  NAND2_X1   g06562(.A1(new_n7564_), .A2(new_n7557_), .ZN(new_n7565_));
  INV_X1     g06563(.I(\A[7] ), .ZN(new_n7566_));
  INV_X1     g06564(.I(\A[8] ), .ZN(new_n7567_));
  NAND2_X1   g06565(.A1(new_n7567_), .A2(\A[9] ), .ZN(new_n7568_));
  INV_X1     g06566(.I(\A[9] ), .ZN(new_n7569_));
  NAND2_X1   g06567(.A1(new_n7569_), .A2(\A[8] ), .ZN(new_n7570_));
  AOI21_X1   g06568(.A1(new_n7568_), .A2(new_n7570_), .B(new_n7566_), .ZN(new_n7571_));
  NAND2_X1   g06569(.A1(\A[8] ), .A2(\A[9] ), .ZN(new_n7572_));
  NOR2_X1    g06570(.A1(\A[8] ), .A2(\A[9] ), .ZN(new_n7573_));
  INV_X1     g06571(.I(new_n7573_), .ZN(new_n7574_));
  AOI21_X1   g06572(.A1(new_n7574_), .A2(new_n7572_), .B(\A[7] ), .ZN(new_n7575_));
  NOR2_X1    g06573(.A1(new_n7575_), .A2(new_n7571_), .ZN(new_n7576_));
  INV_X1     g06574(.I(\A[12] ), .ZN(new_n7577_));
  NOR2_X1    g06575(.A1(new_n7577_), .A2(\A[11] ), .ZN(new_n7578_));
  INV_X1     g06576(.I(\A[11] ), .ZN(new_n7579_));
  NOR2_X1    g06577(.A1(new_n7579_), .A2(\A[12] ), .ZN(new_n7580_));
  OAI21_X1   g06578(.A1(new_n7578_), .A2(new_n7580_), .B(\A[10] ), .ZN(new_n7581_));
  INV_X1     g06579(.I(\A[10] ), .ZN(new_n7582_));
  NAND2_X1   g06580(.A1(\A[11] ), .A2(\A[12] ), .ZN(new_n7583_));
  INV_X1     g06581(.I(new_n7583_), .ZN(new_n7584_));
  NOR2_X1    g06582(.A1(\A[11] ), .A2(\A[12] ), .ZN(new_n7585_));
  OAI21_X1   g06583(.A1(new_n7584_), .A2(new_n7585_), .B(new_n7582_), .ZN(new_n7586_));
  NAND2_X1   g06584(.A1(new_n7581_), .A2(new_n7586_), .ZN(new_n7587_));
  NAND2_X1   g06585(.A1(new_n7576_), .A2(new_n7587_), .ZN(new_n7588_));
  NOR2_X1    g06586(.A1(new_n7569_), .A2(\A[8] ), .ZN(new_n7589_));
  NOR2_X1    g06587(.A1(new_n7567_), .A2(\A[9] ), .ZN(new_n7590_));
  OAI21_X1   g06588(.A1(new_n7589_), .A2(new_n7590_), .B(\A[7] ), .ZN(new_n7591_));
  INV_X1     g06589(.I(new_n7572_), .ZN(new_n7592_));
  OAI21_X1   g06590(.A1(new_n7592_), .A2(new_n7573_), .B(new_n7566_), .ZN(new_n7593_));
  NAND2_X1   g06591(.A1(new_n7591_), .A2(new_n7593_), .ZN(new_n7594_));
  NAND2_X1   g06592(.A1(new_n7579_), .A2(\A[12] ), .ZN(new_n7595_));
  NAND2_X1   g06593(.A1(new_n7577_), .A2(\A[11] ), .ZN(new_n7596_));
  AOI21_X1   g06594(.A1(new_n7595_), .A2(new_n7596_), .B(new_n7582_), .ZN(new_n7597_));
  INV_X1     g06595(.I(new_n7585_), .ZN(new_n7598_));
  AOI21_X1   g06596(.A1(new_n7598_), .A2(new_n7583_), .B(\A[10] ), .ZN(new_n7599_));
  NOR2_X1    g06597(.A1(new_n7599_), .A2(new_n7597_), .ZN(new_n7600_));
  NAND2_X1   g06598(.A1(new_n7600_), .A2(new_n7594_), .ZN(new_n7601_));
  AOI22_X1   g06599(.A1(new_n7588_), .A2(new_n7601_), .B1(new_n7565_), .B2(new_n7551_), .ZN(new_n7602_));
  NOR2_X1    g06600(.A1(new_n7564_), .A2(new_n7557_), .ZN(new_n7603_));
  NOR2_X1    g06601(.A1(new_n7540_), .A2(new_n7550_), .ZN(new_n7604_));
  NOR2_X1    g06602(.A1(new_n7600_), .A2(new_n7594_), .ZN(new_n7605_));
  NOR2_X1    g06603(.A1(new_n7576_), .A2(new_n7587_), .ZN(new_n7606_));
  NOR4_X1    g06604(.A1(new_n7603_), .A2(new_n7605_), .A3(new_n7606_), .A4(new_n7604_), .ZN(new_n7607_));
  NOR2_X1    g06605(.A1(new_n7607_), .A2(new_n7602_), .ZN(new_n7608_));
  INV_X1     g06606(.I(\A[27] ), .ZN(new_n7609_));
  NOR2_X1    g06607(.A1(new_n7609_), .A2(\A[26] ), .ZN(new_n7610_));
  INV_X1     g06608(.I(\A[26] ), .ZN(new_n7611_));
  NOR2_X1    g06609(.A1(new_n7611_), .A2(\A[27] ), .ZN(new_n7612_));
  OAI21_X1   g06610(.A1(new_n7610_), .A2(new_n7612_), .B(\A[25] ), .ZN(new_n7613_));
  INV_X1     g06611(.I(\A[25] ), .ZN(new_n7614_));
  NOR2_X1    g06612(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n7615_));
  NAND2_X1   g06613(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n7616_));
  INV_X1     g06614(.I(new_n7616_), .ZN(new_n7617_));
  OAI21_X1   g06615(.A1(new_n7617_), .A2(new_n7615_), .B(new_n7614_), .ZN(new_n7618_));
  NAND2_X1   g06616(.A1(new_n7613_), .A2(new_n7618_), .ZN(new_n7619_));
  INV_X1     g06617(.I(\A[28] ), .ZN(new_n7620_));
  INV_X1     g06618(.I(\A[29] ), .ZN(new_n7621_));
  NAND2_X1   g06619(.A1(new_n7621_), .A2(\A[30] ), .ZN(new_n7622_));
  INV_X1     g06620(.I(\A[30] ), .ZN(new_n7623_));
  NAND2_X1   g06621(.A1(new_n7623_), .A2(\A[29] ), .ZN(new_n7624_));
  AOI21_X1   g06622(.A1(new_n7622_), .A2(new_n7624_), .B(new_n7620_), .ZN(new_n7625_));
  NOR2_X1    g06623(.A1(\A[29] ), .A2(\A[30] ), .ZN(new_n7626_));
  INV_X1     g06624(.I(new_n7626_), .ZN(new_n7627_));
  NAND2_X1   g06625(.A1(\A[29] ), .A2(\A[30] ), .ZN(new_n7628_));
  AOI21_X1   g06626(.A1(new_n7627_), .A2(new_n7628_), .B(\A[28] ), .ZN(new_n7629_));
  NOR2_X1    g06627(.A1(new_n7629_), .A2(new_n7625_), .ZN(new_n7630_));
  NOR2_X1    g06628(.A1(new_n7630_), .A2(new_n7619_), .ZN(new_n7631_));
  NAND2_X1   g06629(.A1(new_n7611_), .A2(\A[27] ), .ZN(new_n7632_));
  NAND2_X1   g06630(.A1(new_n7609_), .A2(\A[26] ), .ZN(new_n7633_));
  AOI21_X1   g06631(.A1(new_n7632_), .A2(new_n7633_), .B(new_n7614_), .ZN(new_n7634_));
  INV_X1     g06632(.I(new_n7615_), .ZN(new_n7635_));
  AOI21_X1   g06633(.A1(new_n7635_), .A2(new_n7616_), .B(\A[25] ), .ZN(new_n7636_));
  NOR2_X1    g06634(.A1(new_n7636_), .A2(new_n7634_), .ZN(new_n7637_));
  NOR2_X1    g06635(.A1(new_n7623_), .A2(\A[29] ), .ZN(new_n7638_));
  NOR2_X1    g06636(.A1(new_n7621_), .A2(\A[30] ), .ZN(new_n7639_));
  OAI21_X1   g06637(.A1(new_n7638_), .A2(new_n7639_), .B(\A[28] ), .ZN(new_n7640_));
  AND2_X2    g06638(.A1(\A[29] ), .A2(\A[30] ), .Z(new_n7641_));
  OAI21_X1   g06639(.A1(new_n7641_), .A2(new_n7626_), .B(new_n7620_), .ZN(new_n7642_));
  NAND2_X1   g06640(.A1(new_n7640_), .A2(new_n7642_), .ZN(new_n7643_));
  NOR2_X1    g06641(.A1(new_n7637_), .A2(new_n7643_), .ZN(new_n7644_));
  INV_X1     g06642(.I(\A[21] ), .ZN(new_n7645_));
  NOR2_X1    g06643(.A1(new_n7645_), .A2(\A[20] ), .ZN(new_n7646_));
  INV_X1     g06644(.I(\A[20] ), .ZN(new_n7647_));
  NOR2_X1    g06645(.A1(new_n7647_), .A2(\A[21] ), .ZN(new_n7648_));
  OAI21_X1   g06646(.A1(new_n7646_), .A2(new_n7648_), .B(\A[19] ), .ZN(new_n7649_));
  INV_X1     g06647(.I(\A[19] ), .ZN(new_n7650_));
  AND2_X2    g06648(.A1(\A[20] ), .A2(\A[21] ), .Z(new_n7651_));
  NOR2_X1    g06649(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n7652_));
  OAI21_X1   g06650(.A1(new_n7651_), .A2(new_n7652_), .B(new_n7650_), .ZN(new_n7653_));
  NAND2_X1   g06651(.A1(new_n7649_), .A2(new_n7653_), .ZN(new_n7654_));
  INV_X1     g06652(.I(\A[22] ), .ZN(new_n7655_));
  INV_X1     g06653(.I(\A[23] ), .ZN(new_n7656_));
  NAND2_X1   g06654(.A1(new_n7656_), .A2(\A[24] ), .ZN(new_n7657_));
  INV_X1     g06655(.I(\A[24] ), .ZN(new_n7658_));
  NAND2_X1   g06656(.A1(new_n7658_), .A2(\A[23] ), .ZN(new_n7659_));
  AOI21_X1   g06657(.A1(new_n7657_), .A2(new_n7659_), .B(new_n7655_), .ZN(new_n7660_));
  NAND2_X1   g06658(.A1(\A[23] ), .A2(\A[24] ), .ZN(new_n7661_));
  NOR2_X1    g06659(.A1(\A[23] ), .A2(\A[24] ), .ZN(new_n7662_));
  INV_X1     g06660(.I(new_n7662_), .ZN(new_n7663_));
  AOI21_X1   g06661(.A1(new_n7663_), .A2(new_n7661_), .B(\A[22] ), .ZN(new_n7664_));
  NOR2_X1    g06662(.A1(new_n7664_), .A2(new_n7660_), .ZN(new_n7665_));
  NOR2_X1    g06663(.A1(new_n7665_), .A2(new_n7654_), .ZN(new_n7666_));
  NAND2_X1   g06664(.A1(new_n7647_), .A2(\A[21] ), .ZN(new_n7667_));
  NAND2_X1   g06665(.A1(new_n7645_), .A2(\A[20] ), .ZN(new_n7668_));
  AOI21_X1   g06666(.A1(new_n7667_), .A2(new_n7668_), .B(new_n7650_), .ZN(new_n7669_));
  NAND2_X1   g06667(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n7670_));
  INV_X1     g06668(.I(new_n7652_), .ZN(new_n7671_));
  AOI21_X1   g06669(.A1(new_n7671_), .A2(new_n7670_), .B(\A[19] ), .ZN(new_n7672_));
  NOR2_X1    g06670(.A1(new_n7672_), .A2(new_n7669_), .ZN(new_n7673_));
  NOR2_X1    g06671(.A1(new_n7658_), .A2(\A[23] ), .ZN(new_n7674_));
  NOR2_X1    g06672(.A1(new_n7656_), .A2(\A[24] ), .ZN(new_n7675_));
  OAI21_X1   g06673(.A1(new_n7674_), .A2(new_n7675_), .B(\A[22] ), .ZN(new_n7676_));
  AND2_X2    g06674(.A1(\A[23] ), .A2(\A[24] ), .Z(new_n7677_));
  OAI21_X1   g06675(.A1(new_n7677_), .A2(new_n7662_), .B(new_n7655_), .ZN(new_n7678_));
  NAND2_X1   g06676(.A1(new_n7676_), .A2(new_n7678_), .ZN(new_n7679_));
  NOR2_X1    g06677(.A1(new_n7673_), .A2(new_n7679_), .ZN(new_n7680_));
  OAI22_X1   g06678(.A1(new_n7631_), .A2(new_n7644_), .B1(new_n7666_), .B2(new_n7680_), .ZN(new_n7681_));
  NAND2_X1   g06679(.A1(new_n7637_), .A2(new_n7643_), .ZN(new_n7682_));
  NAND2_X1   g06680(.A1(new_n7630_), .A2(new_n7619_), .ZN(new_n7683_));
  NAND2_X1   g06681(.A1(new_n7673_), .A2(new_n7679_), .ZN(new_n7684_));
  NAND2_X1   g06682(.A1(new_n7665_), .A2(new_n7654_), .ZN(new_n7685_));
  NAND4_X1   g06683(.A1(new_n7682_), .A2(new_n7683_), .A3(new_n7684_), .A4(new_n7685_), .ZN(new_n7686_));
  NAND2_X1   g06684(.A1(new_n7681_), .A2(new_n7686_), .ZN(new_n7687_));
  NOR2_X1    g06685(.A1(new_n7608_), .A2(new_n7687_), .ZN(new_n7688_));
  NAND2_X1   g06686(.A1(new_n7608_), .A2(new_n7687_), .ZN(new_n7689_));
  INV_X1     g06687(.I(new_n7689_), .ZN(new_n7690_));
  NOR3_X1    g06688(.A1(new_n7529_), .A2(new_n7690_), .A3(new_n7688_), .ZN(new_n7691_));
  INV_X1     g06689(.I(new_n7526_), .ZN(new_n7692_));
  NOR2_X1    g06690(.A1(new_n7692_), .A2(new_n7527_), .ZN(new_n7693_));
  INV_X1     g06691(.I(new_n7688_), .ZN(new_n7694_));
  AOI21_X1   g06692(.A1(new_n7689_), .A2(new_n7694_), .B(new_n7693_), .ZN(new_n7695_));
  NOR2_X1    g06693(.A1(new_n7695_), .A2(new_n7691_), .ZN(new_n7696_));
  XOR2_X1    g06694(.A1(new_n7696_), .A2(new_n7453_), .Z(new_n7697_));
  NOR2_X1    g06695(.A1(new_n7697_), .A2(new_n7122_), .ZN(new_n7698_));
  NOR2_X1    g06696(.A1(new_n7594_), .A2(new_n7587_), .ZN(new_n7699_));
  AOI21_X1   g06697(.A1(\A[11] ), .A2(\A[12] ), .B(\A[10] ), .ZN(new_n7700_));
  AOI21_X1   g06698(.A1(\A[8] ), .A2(\A[9] ), .B(\A[7] ), .ZN(new_n7701_));
  NOR4_X1    g06699(.A1(new_n7700_), .A2(new_n7701_), .A3(new_n7573_), .A4(new_n7585_), .ZN(new_n7702_));
  NAND2_X1   g06700(.A1(new_n7699_), .A2(new_n7702_), .ZN(new_n7703_));
  AOI21_X1   g06701(.A1(\A[17] ), .A2(\A[18] ), .B(\A[16] ), .ZN(new_n7704_));
  AOI21_X1   g06702(.A1(\A[14] ), .A2(\A[15] ), .B(\A[13] ), .ZN(new_n7705_));
  NOR2_X1    g06703(.A1(new_n7705_), .A2(new_n7536_), .ZN(new_n7706_));
  NOR3_X1    g06704(.A1(new_n7706_), .A2(new_n7547_), .A3(new_n7704_), .ZN(new_n7707_));
  NOR2_X1    g06705(.A1(new_n7704_), .A2(new_n7547_), .ZN(new_n7708_));
  NOR3_X1    g06706(.A1(new_n7708_), .A2(new_n7536_), .A3(new_n7705_), .ZN(new_n7709_));
  OAI22_X1   g06707(.A1(new_n7557_), .A2(new_n7550_), .B1(new_n7707_), .B2(new_n7709_), .ZN(new_n7710_));
  INV_X1     g06708(.I(new_n7706_), .ZN(new_n7711_));
  NAND2_X1   g06709(.A1(new_n7711_), .A2(new_n7708_), .ZN(new_n7712_));
  INV_X1     g06710(.I(new_n7708_), .ZN(new_n7713_));
  NAND2_X1   g06711(.A1(new_n7713_), .A2(new_n7706_), .ZN(new_n7714_));
  NAND4_X1   g06712(.A1(new_n7540_), .A2(new_n7564_), .A3(new_n7714_), .A4(new_n7712_), .ZN(new_n7715_));
  NAND2_X1   g06713(.A1(new_n7715_), .A2(new_n7710_), .ZN(new_n7716_));
  NOR2_X1    g06714(.A1(new_n7711_), .A2(new_n7713_), .ZN(new_n7717_));
  OAI21_X1   g06715(.A1(new_n7540_), .A2(new_n7564_), .B(new_n7717_), .ZN(new_n7718_));
  NAND4_X1   g06716(.A1(new_n7602_), .A2(new_n7716_), .A3(new_n7703_), .A4(new_n7718_), .ZN(new_n7719_));
  INV_X1     g06717(.I(new_n7702_), .ZN(new_n7720_));
  OAI22_X1   g06718(.A1(new_n7573_), .A2(new_n7701_), .B1(new_n7700_), .B2(new_n7585_), .ZN(new_n7721_));
  NAND2_X1   g06719(.A1(new_n7720_), .A2(new_n7721_), .ZN(new_n7722_));
  XOR2_X1    g06720(.A1(new_n7699_), .A2(new_n7722_), .Z(new_n7723_));
  NOR2_X1    g06721(.A1(new_n7557_), .A2(new_n7550_), .ZN(new_n7724_));
  AOI22_X1   g06722(.A1(new_n7699_), .A2(new_n7702_), .B1(new_n7724_), .B2(new_n7717_), .ZN(new_n7725_));
  AOI21_X1   g06723(.A1(new_n7602_), .A2(new_n7725_), .B(new_n7716_), .ZN(new_n7726_));
  NOR2_X1    g06724(.A1(new_n7726_), .A2(new_n7723_), .ZN(new_n7727_));
  OAI22_X1   g06725(.A1(new_n7605_), .A2(new_n7606_), .B1(new_n7603_), .B2(new_n7604_), .ZN(new_n7728_));
  AOI22_X1   g06726(.A1(new_n7540_), .A2(new_n7564_), .B1(new_n7714_), .B2(new_n7712_), .ZN(new_n7729_));
  NOR4_X1    g06727(.A1(new_n7557_), .A2(new_n7550_), .A3(new_n7707_), .A4(new_n7709_), .ZN(new_n7730_));
  NOR2_X1    g06728(.A1(new_n7729_), .A2(new_n7730_), .ZN(new_n7731_));
  NAND2_X1   g06729(.A1(new_n7576_), .A2(new_n7600_), .ZN(new_n7732_));
  NAND4_X1   g06730(.A1(new_n7554_), .A2(new_n7545_), .A3(new_n7556_), .A4(new_n7549_), .ZN(new_n7733_));
  INV_X1     g06731(.I(new_n7717_), .ZN(new_n7734_));
  OAI22_X1   g06732(.A1(new_n7732_), .A2(new_n7720_), .B1(new_n7734_), .B2(new_n7733_), .ZN(new_n7735_));
  OAI21_X1   g06733(.A1(new_n7728_), .A2(new_n7735_), .B(new_n7731_), .ZN(new_n7736_));
  NAND3_X1   g06734(.A1(new_n7602_), .A2(new_n7725_), .A3(new_n7716_), .ZN(new_n7737_));
  NAND2_X1   g06735(.A1(new_n7736_), .A2(new_n7737_), .ZN(new_n7738_));
  AOI22_X1   g06736(.A1(new_n7738_), .A2(new_n7723_), .B1(new_n7727_), .B2(new_n7719_), .ZN(new_n7739_));
  NAND3_X1   g06737(.A1(new_n7608_), .A2(new_n7681_), .A3(new_n7686_), .ZN(new_n7740_));
  NAND4_X1   g06738(.A1(new_n7649_), .A2(new_n7676_), .A3(new_n7653_), .A4(new_n7678_), .ZN(new_n7741_));
  AOI21_X1   g06739(.A1(\A[23] ), .A2(\A[24] ), .B(\A[22] ), .ZN(new_n7742_));
  AOI21_X1   g06740(.A1(\A[20] ), .A2(\A[21] ), .B(\A[19] ), .ZN(new_n7743_));
  OAI22_X1   g06741(.A1(new_n7652_), .A2(new_n7743_), .B1(new_n7742_), .B2(new_n7662_), .ZN(new_n7744_));
  NOR4_X1    g06742(.A1(new_n7742_), .A2(new_n7743_), .A3(new_n7652_), .A4(new_n7662_), .ZN(new_n7745_));
  INV_X1     g06743(.I(new_n7745_), .ZN(new_n7746_));
  NAND2_X1   g06744(.A1(new_n7746_), .A2(new_n7744_), .ZN(new_n7747_));
  XNOR2_X1   g06745(.A1(new_n7747_), .A2(new_n7741_), .ZN(new_n7748_));
  AOI21_X1   g06746(.A1(\A[29] ), .A2(\A[30] ), .B(\A[28] ), .ZN(new_n7749_));
  NOR2_X1    g06747(.A1(new_n7749_), .A2(new_n7626_), .ZN(new_n7750_));
  AOI21_X1   g06748(.A1(\A[26] ), .A2(\A[27] ), .B(\A[25] ), .ZN(new_n7751_));
  NOR2_X1    g06749(.A1(new_n7751_), .A2(new_n7615_), .ZN(new_n7752_));
  NAND2_X1   g06750(.A1(new_n7750_), .A2(new_n7752_), .ZN(new_n7753_));
  NAND4_X1   g06751(.A1(new_n7613_), .A2(new_n7640_), .A3(new_n7618_), .A4(new_n7642_), .ZN(new_n7754_));
  OAI22_X1   g06752(.A1(new_n7753_), .A2(new_n7754_), .B1(new_n7741_), .B2(new_n7746_), .ZN(new_n7755_));
  NOR3_X1    g06753(.A1(new_n7752_), .A2(new_n7626_), .A3(new_n7749_), .ZN(new_n7756_));
  NOR3_X1    g06754(.A1(new_n7750_), .A2(new_n7615_), .A3(new_n7751_), .ZN(new_n7757_));
  NOR2_X1    g06755(.A1(new_n7756_), .A2(new_n7757_), .ZN(new_n7758_));
  NAND2_X1   g06756(.A1(new_n7758_), .A2(new_n7754_), .ZN(new_n7759_));
  NOR4_X1    g06757(.A1(new_n7634_), .A2(new_n7636_), .A3(new_n7629_), .A4(new_n7625_), .ZN(new_n7760_));
  XOR2_X1    g06758(.A1(new_n7750_), .A2(new_n7752_), .Z(new_n7761_));
  NAND2_X1   g06759(.A1(new_n7761_), .A2(new_n7760_), .ZN(new_n7762_));
  NAND2_X1   g06760(.A1(new_n7762_), .A2(new_n7759_), .ZN(new_n7763_));
  OAI21_X1   g06761(.A1(new_n7681_), .A2(new_n7755_), .B(new_n7763_), .ZN(new_n7764_));
  AOI22_X1   g06762(.A1(new_n7682_), .A2(new_n7683_), .B1(new_n7684_), .B2(new_n7685_), .ZN(new_n7765_));
  INV_X1     g06763(.I(new_n7741_), .ZN(new_n7766_));
  INV_X1     g06764(.I(new_n7753_), .ZN(new_n7767_));
  AOI22_X1   g06765(.A1(new_n7766_), .A2(new_n7745_), .B1(new_n7767_), .B2(new_n7760_), .ZN(new_n7768_));
  NOR2_X1    g06766(.A1(new_n7761_), .A2(new_n7760_), .ZN(new_n7769_));
  NOR2_X1    g06767(.A1(new_n7758_), .A2(new_n7754_), .ZN(new_n7770_));
  NOR2_X1    g06768(.A1(new_n7769_), .A2(new_n7770_), .ZN(new_n7771_));
  NAND3_X1   g06769(.A1(new_n7771_), .A2(new_n7765_), .A3(new_n7768_), .ZN(new_n7772_));
  NAND3_X1   g06770(.A1(new_n7764_), .A2(new_n7772_), .A3(new_n7748_), .ZN(new_n7773_));
  XOR2_X1    g06771(.A1(new_n7747_), .A2(new_n7741_), .Z(new_n7774_));
  AOI21_X1   g06772(.A1(new_n7765_), .A2(new_n7768_), .B(new_n7771_), .ZN(new_n7775_));
  NAND3_X1   g06773(.A1(new_n7673_), .A2(new_n7665_), .A3(new_n7745_), .ZN(new_n7776_));
  NAND3_X1   g06774(.A1(new_n7762_), .A2(new_n7759_), .A3(new_n7776_), .ZN(new_n7777_));
  AOI21_X1   g06775(.A1(new_n7619_), .A2(new_n7643_), .B(new_n7753_), .ZN(new_n7778_));
  NOR3_X1    g06776(.A1(new_n7777_), .A2(new_n7681_), .A3(new_n7778_), .ZN(new_n7779_));
  OAI21_X1   g06777(.A1(new_n7775_), .A2(new_n7779_), .B(new_n7774_), .ZN(new_n7780_));
  AOI21_X1   g06778(.A1(new_n7780_), .A2(new_n7773_), .B(new_n7740_), .ZN(new_n7781_));
  NOR3_X1    g06779(.A1(new_n7687_), .A2(new_n7602_), .A3(new_n7607_), .ZN(new_n7782_));
  NOR3_X1    g06780(.A1(new_n7681_), .A2(new_n7763_), .A3(new_n7755_), .ZN(new_n7783_));
  NOR3_X1    g06781(.A1(new_n7775_), .A2(new_n7783_), .A3(new_n7774_), .ZN(new_n7784_));
  INV_X1     g06782(.I(new_n7778_), .ZN(new_n7785_));
  NAND4_X1   g06783(.A1(new_n7771_), .A2(new_n7765_), .A3(new_n7776_), .A4(new_n7785_), .ZN(new_n7786_));
  AOI21_X1   g06784(.A1(new_n7786_), .A2(new_n7764_), .B(new_n7748_), .ZN(new_n7787_));
  NOR3_X1    g06785(.A1(new_n7787_), .A2(new_n7784_), .A3(new_n7782_), .ZN(new_n7788_));
  OAI21_X1   g06786(.A1(new_n7788_), .A2(new_n7781_), .B(new_n7739_), .ZN(new_n7789_));
  XOR2_X1    g06787(.A1(new_n7732_), .A2(new_n7722_), .Z(new_n7790_));
  NAND3_X1   g06788(.A1(new_n7736_), .A2(new_n7719_), .A3(new_n7790_), .ZN(new_n7791_));
  NOR3_X1    g06789(.A1(new_n7728_), .A2(new_n7731_), .A3(new_n7735_), .ZN(new_n7792_));
  OAI21_X1   g06790(.A1(new_n7726_), .A2(new_n7792_), .B(new_n7723_), .ZN(new_n7793_));
  NAND2_X1   g06791(.A1(new_n7793_), .A2(new_n7791_), .ZN(new_n7794_));
  OAI21_X1   g06792(.A1(new_n7787_), .A2(new_n7784_), .B(new_n7782_), .ZN(new_n7795_));
  NAND3_X1   g06793(.A1(new_n7780_), .A2(new_n7773_), .A3(new_n7740_), .ZN(new_n7796_));
  NAND3_X1   g06794(.A1(new_n7795_), .A2(new_n7796_), .A3(new_n7794_), .ZN(new_n7797_));
  NAND2_X1   g06795(.A1(new_n7789_), .A2(new_n7797_), .ZN(new_n7798_));
  OAI21_X1   g06796(.A1(new_n7688_), .A2(new_n7690_), .B(new_n7693_), .ZN(new_n7799_));
  NOR2_X1    g06797(.A1(new_n7462_), .A2(new_n7471_), .ZN(new_n7800_));
  NOR2_X1    g06798(.A1(new_n7469_), .A2(\A[994] ), .ZN(new_n7801_));
  NOR2_X1    g06799(.A1(new_n7801_), .A2(new_n7468_), .ZN(new_n7802_));
  NOR2_X1    g06800(.A1(new_n7460_), .A2(\A[991] ), .ZN(new_n7803_));
  NOR2_X1    g06801(.A1(new_n7803_), .A2(new_n7459_), .ZN(new_n7804_));
  NOR2_X1    g06802(.A1(new_n7802_), .A2(new_n7804_), .ZN(new_n7805_));
  INV_X1     g06803(.I(new_n7805_), .ZN(new_n7806_));
  NAND2_X1   g06804(.A1(new_n7802_), .A2(new_n7804_), .ZN(new_n7807_));
  NAND2_X1   g06805(.A1(new_n7806_), .A2(new_n7807_), .ZN(new_n7808_));
  XOR2_X1    g06806(.A1(new_n7808_), .A2(new_n7800_), .Z(new_n7809_));
  NOR2_X1    g06807(.A1(new_n7476_), .A2(\A[997] ), .ZN(new_n7810_));
  NOR2_X1    g06808(.A1(new_n7810_), .A2(new_n7477_), .ZN(new_n7811_));
  INV_X1     g06809(.I(new_n7811_), .ZN(new_n7812_));
  AOI21_X1   g06810(.A1(new_n7485_), .A2(new_n7486_), .B(new_n7488_), .ZN(new_n7813_));
  AOI21_X1   g06811(.A1(new_n7497_), .A2(new_n7498_), .B(new_n7499_), .ZN(new_n7814_));
  XOR2_X1    g06812(.A1(new_n7814_), .A2(new_n7813_), .Z(new_n7815_));
  AOI21_X1   g06813(.A1(new_n7505_), .A2(new_n7516_), .B(new_n7491_), .ZN(new_n7816_));
  INV_X1     g06814(.I(new_n7816_), .ZN(new_n7817_));
  AOI21_X1   g06815(.A1(new_n7523_), .A2(new_n7817_), .B(new_n7815_), .ZN(new_n7818_));
  NAND2_X1   g06816(.A1(new_n7814_), .A2(new_n7813_), .ZN(new_n7819_));
  OR2_X2     g06817(.A1(new_n7814_), .A2(new_n7813_), .Z(new_n7820_));
  NAND2_X1   g06818(.A1(new_n7820_), .A2(new_n7819_), .ZN(new_n7821_));
  NOR3_X1    g06819(.A1(new_n7508_), .A2(new_n7821_), .A3(new_n7816_), .ZN(new_n7822_));
  OAI21_X1   g06820(.A1(new_n7818_), .A2(new_n7822_), .B(new_n7521_), .ZN(new_n7823_));
  NAND3_X1   g06821(.A1(new_n7523_), .A2(new_n7524_), .A3(new_n7522_), .ZN(new_n7824_));
  OAI21_X1   g06822(.A1(new_n7508_), .A2(new_n7816_), .B(new_n7821_), .ZN(new_n7825_));
  NAND3_X1   g06823(.A1(new_n7523_), .A2(new_n7815_), .A3(new_n7817_), .ZN(new_n7826_));
  NAND3_X1   g06824(.A1(new_n7824_), .A2(new_n7825_), .A3(new_n7826_), .ZN(new_n7827_));
  AOI21_X1   g06825(.A1(new_n7823_), .A2(new_n7827_), .B(new_n7812_), .ZN(new_n7828_));
  AOI21_X1   g06826(.A1(new_n7825_), .A2(new_n7826_), .B(new_n7824_), .ZN(new_n7829_));
  NOR3_X1    g06827(.A1(new_n7521_), .A2(new_n7822_), .A3(new_n7818_), .ZN(new_n7830_));
  NOR3_X1    g06828(.A1(new_n7829_), .A2(new_n7830_), .A3(new_n7811_), .ZN(new_n7831_));
  OAI21_X1   g06829(.A1(new_n7831_), .A2(new_n7828_), .B(new_n7527_), .ZN(new_n7832_));
  OAI21_X1   g06830(.A1(new_n7829_), .A2(new_n7830_), .B(new_n7811_), .ZN(new_n7833_));
  NAND3_X1   g06831(.A1(new_n7823_), .A2(new_n7827_), .A3(new_n7812_), .ZN(new_n7834_));
  NAND3_X1   g06832(.A1(new_n7833_), .A2(new_n7834_), .A3(new_n7528_), .ZN(new_n7835_));
  NAND3_X1   g06833(.A1(new_n7832_), .A2(new_n7835_), .A3(new_n7809_), .ZN(new_n7836_));
  INV_X1     g06834(.I(new_n7809_), .ZN(new_n7837_));
  AOI21_X1   g06835(.A1(new_n7833_), .A2(new_n7834_), .B(new_n7528_), .ZN(new_n7838_));
  NOR3_X1    g06836(.A1(new_n7831_), .A2(new_n7828_), .A3(new_n7527_), .ZN(new_n7839_));
  OAI21_X1   g06837(.A1(new_n7839_), .A2(new_n7838_), .B(new_n7837_), .ZN(new_n7840_));
  NAND3_X1   g06838(.A1(new_n7840_), .A2(new_n7836_), .A3(new_n7799_), .ZN(new_n7841_));
  AOI21_X1   g06839(.A1(new_n7689_), .A2(new_n7694_), .B(new_n7529_), .ZN(new_n7842_));
  NOR3_X1    g06840(.A1(new_n7839_), .A2(new_n7838_), .A3(new_n7837_), .ZN(new_n7843_));
  AOI21_X1   g06841(.A1(new_n7832_), .A2(new_n7835_), .B(new_n7809_), .ZN(new_n7844_));
  OAI21_X1   g06842(.A1(new_n7843_), .A2(new_n7844_), .B(new_n7842_), .ZN(new_n7845_));
  NAND3_X1   g06843(.A1(new_n7845_), .A2(new_n7841_), .A3(new_n7798_), .ZN(new_n7846_));
  AOI21_X1   g06844(.A1(new_n7795_), .A2(new_n7796_), .B(new_n7794_), .ZN(new_n7847_));
  NOR3_X1    g06845(.A1(new_n7739_), .A2(new_n7788_), .A3(new_n7781_), .ZN(new_n7848_));
  NOR2_X1    g06846(.A1(new_n7848_), .A2(new_n7847_), .ZN(new_n7849_));
  NOR3_X1    g06847(.A1(new_n7843_), .A2(new_n7844_), .A3(new_n7842_), .ZN(new_n7850_));
  AOI21_X1   g06848(.A1(new_n7840_), .A2(new_n7836_), .B(new_n7799_), .ZN(new_n7851_));
  OAI21_X1   g06849(.A1(new_n7850_), .A2(new_n7851_), .B(new_n7849_), .ZN(new_n7852_));
  NAND2_X1   g06850(.A1(new_n7852_), .A2(new_n7846_), .ZN(new_n7853_));
  OAI21_X1   g06851(.A1(new_n7691_), .A2(new_n7695_), .B(new_n7453_), .ZN(new_n7854_));
  INV_X1     g06852(.I(new_n7854_), .ZN(new_n7855_));
  NOR2_X1    g06853(.A1(new_n7187_), .A2(new_n7180_), .ZN(new_n7856_));
  AOI21_X1   g06854(.A1(new_n7175_), .A2(new_n7176_), .B(new_n7178_), .ZN(new_n7857_));
  INV_X1     g06855(.I(new_n7857_), .ZN(new_n7858_));
  AOI21_X1   g06856(.A1(new_n7159_), .A2(new_n7165_), .B(new_n7166_), .ZN(new_n7859_));
  INV_X1     g06857(.I(new_n7859_), .ZN(new_n7860_));
  NOR2_X1    g06858(.A1(new_n7858_), .A2(new_n7860_), .ZN(new_n7861_));
  NAND2_X1   g06859(.A1(new_n7856_), .A2(new_n7861_), .ZN(new_n7862_));
  AOI21_X1   g06860(.A1(\A[65] ), .A2(\A[66] ), .B(\A[64] ), .ZN(new_n7863_));
  AOI21_X1   g06861(.A1(\A[62] ), .A2(\A[63] ), .B(\A[61] ), .ZN(new_n7864_));
  NOR2_X1    g06862(.A1(new_n7864_), .A2(new_n7129_), .ZN(new_n7865_));
  NOR3_X1    g06863(.A1(new_n7865_), .A2(new_n7140_), .A3(new_n7863_), .ZN(new_n7866_));
  NOR2_X1    g06864(.A1(new_n7863_), .A2(new_n7140_), .ZN(new_n7867_));
  NOR3_X1    g06865(.A1(new_n7867_), .A2(new_n7129_), .A3(new_n7864_), .ZN(new_n7868_));
  OAI22_X1   g06866(.A1(new_n7151_), .A2(new_n7144_), .B1(new_n7866_), .B2(new_n7868_), .ZN(new_n7869_));
  NOR4_X1    g06867(.A1(new_n7128_), .A2(new_n7132_), .A3(new_n7156_), .A4(new_n7154_), .ZN(new_n7870_));
  INV_X1     g06868(.I(new_n7865_), .ZN(new_n7871_));
  NAND2_X1   g06869(.A1(new_n7871_), .A2(new_n7867_), .ZN(new_n7872_));
  INV_X1     g06870(.I(new_n7867_), .ZN(new_n7873_));
  NAND2_X1   g06871(.A1(new_n7873_), .A2(new_n7865_), .ZN(new_n7874_));
  NAND3_X1   g06872(.A1(new_n7870_), .A2(new_n7872_), .A3(new_n7874_), .ZN(new_n7875_));
  NAND2_X1   g06873(.A1(new_n7875_), .A2(new_n7869_), .ZN(new_n7876_));
  NOR2_X1    g06874(.A1(new_n7873_), .A2(new_n7871_), .ZN(new_n7877_));
  OAI21_X1   g06875(.A1(new_n7133_), .A2(new_n7157_), .B(new_n7877_), .ZN(new_n7878_));
  NAND4_X1   g06876(.A1(new_n7195_), .A2(new_n7876_), .A3(new_n7862_), .A4(new_n7878_), .ZN(new_n7879_));
  NOR2_X1    g06877(.A1(new_n7857_), .A2(new_n7859_), .ZN(new_n7880_));
  NOR2_X1    g06878(.A1(new_n7861_), .A2(new_n7880_), .ZN(new_n7881_));
  XOR2_X1    g06879(.A1(new_n7881_), .A2(new_n7856_), .Z(new_n7882_));
  OAI22_X1   g06880(.A1(new_n7196_), .A2(new_n7197_), .B1(new_n7198_), .B2(new_n7199_), .ZN(new_n7883_));
  AOI22_X1   g06881(.A1(new_n7133_), .A2(new_n7157_), .B1(new_n7872_), .B2(new_n7874_), .ZN(new_n7884_));
  NOR4_X1    g06882(.A1(new_n7151_), .A2(new_n7144_), .A3(new_n7866_), .A4(new_n7868_), .ZN(new_n7885_));
  NOR2_X1    g06883(.A1(new_n7884_), .A2(new_n7885_), .ZN(new_n7886_));
  NAND2_X1   g06884(.A1(new_n7169_), .A2(new_n7193_), .ZN(new_n7887_));
  INV_X1     g06885(.I(new_n7861_), .ZN(new_n7888_));
  NAND4_X1   g06886(.A1(new_n7148_), .A2(new_n7150_), .A3(new_n7138_), .A4(new_n7143_), .ZN(new_n7889_));
  INV_X1     g06887(.I(new_n7877_), .ZN(new_n7890_));
  OAI22_X1   g06888(.A1(new_n7887_), .A2(new_n7888_), .B1(new_n7890_), .B2(new_n7889_), .ZN(new_n7891_));
  OAI21_X1   g06889(.A1(new_n7883_), .A2(new_n7891_), .B(new_n7886_), .ZN(new_n7892_));
  NAND3_X1   g06890(.A1(new_n7879_), .A2(new_n7892_), .A3(new_n7882_), .ZN(new_n7893_));
  XOR2_X1    g06891(.A1(new_n7881_), .A2(new_n7887_), .Z(new_n7894_));
  AOI22_X1   g06892(.A1(new_n7856_), .A2(new_n7861_), .B1(new_n7870_), .B2(new_n7877_), .ZN(new_n7895_));
  AOI21_X1   g06893(.A1(new_n7195_), .A2(new_n7895_), .B(new_n7876_), .ZN(new_n7896_));
  NOR3_X1    g06894(.A1(new_n7883_), .A2(new_n7886_), .A3(new_n7891_), .ZN(new_n7897_));
  OAI21_X1   g06895(.A1(new_n7896_), .A2(new_n7897_), .B(new_n7894_), .ZN(new_n7898_));
  NAND2_X1   g06896(.A1(new_n7898_), .A2(new_n7893_), .ZN(new_n7899_));
  NAND4_X1   g06897(.A1(new_n7261_), .A2(new_n7252_), .A3(new_n7263_), .A4(new_n7256_), .ZN(new_n7900_));
  AOI21_X1   g06898(.A1(\A[71] ), .A2(\A[72] ), .B(\A[70] ), .ZN(new_n7901_));
  NOR2_X1    g06899(.A1(new_n7901_), .A2(new_n7255_), .ZN(new_n7902_));
  AOI21_X1   g06900(.A1(\A[68] ), .A2(\A[69] ), .B(\A[67] ), .ZN(new_n7903_));
  NOR2_X1    g06901(.A1(new_n7903_), .A2(new_n7244_), .ZN(new_n7904_));
  NOR2_X1    g06902(.A1(new_n7902_), .A2(new_n7904_), .ZN(new_n7905_));
  NOR4_X1    g06903(.A1(new_n7901_), .A2(new_n7903_), .A3(new_n7244_), .A4(new_n7255_), .ZN(new_n7906_));
  NOR2_X1    g06904(.A1(new_n7905_), .A2(new_n7906_), .ZN(new_n7907_));
  XNOR2_X1   g06905(.A1(new_n7900_), .A2(new_n7907_), .ZN(new_n7908_));
  INV_X1     g06906(.I(new_n7900_), .ZN(new_n7909_));
  AOI21_X1   g06907(.A1(\A[77] ), .A2(\A[78] ), .B(\A[76] ), .ZN(new_n7910_));
  NOR2_X1    g06908(.A1(new_n7910_), .A2(new_n7218_), .ZN(new_n7911_));
  AOI21_X1   g06909(.A1(\A[74] ), .A2(\A[75] ), .B(\A[73] ), .ZN(new_n7912_));
  NOR2_X1    g06910(.A1(new_n7912_), .A2(new_n7207_), .ZN(new_n7913_));
  NAND2_X1   g06911(.A1(new_n7911_), .A2(new_n7913_), .ZN(new_n7914_));
  INV_X1     g06912(.I(new_n7914_), .ZN(new_n7915_));
  NOR4_X1    g06913(.A1(new_n7206_), .A2(new_n7210_), .A3(new_n7234_), .A4(new_n7231_), .ZN(new_n7916_));
  AOI22_X1   g06914(.A1(new_n7909_), .A2(new_n7906_), .B1(new_n7915_), .B2(new_n7916_), .ZN(new_n7917_));
  NAND4_X1   g06915(.A1(new_n7225_), .A2(new_n7216_), .A3(new_n7227_), .A4(new_n7220_), .ZN(new_n7918_));
  NOR3_X1    g06916(.A1(new_n7913_), .A2(new_n7218_), .A3(new_n7910_), .ZN(new_n7919_));
  NOR3_X1    g06917(.A1(new_n7911_), .A2(new_n7207_), .A3(new_n7912_), .ZN(new_n7920_));
  NOR2_X1    g06918(.A1(new_n7919_), .A2(new_n7920_), .ZN(new_n7921_));
  NAND2_X1   g06919(.A1(new_n7921_), .A2(new_n7918_), .ZN(new_n7922_));
  XOR2_X1    g06920(.A1(new_n7911_), .A2(new_n7913_), .Z(new_n7923_));
  NAND2_X1   g06921(.A1(new_n7923_), .A2(new_n7916_), .ZN(new_n7924_));
  AOI22_X1   g06922(.A1(new_n7273_), .A2(new_n7917_), .B1(new_n7922_), .B2(new_n7924_), .ZN(new_n7925_));
  OAI22_X1   g06923(.A1(new_n7274_), .A2(new_n7275_), .B1(new_n7276_), .B2(new_n7277_), .ZN(new_n7926_));
  INV_X1     g06924(.I(new_n7906_), .ZN(new_n7927_));
  OAI22_X1   g06925(.A1(new_n7914_), .A2(new_n7918_), .B1(new_n7900_), .B2(new_n7927_), .ZN(new_n7928_));
  NAND2_X1   g06926(.A1(new_n7924_), .A2(new_n7922_), .ZN(new_n7929_));
  NOR3_X1    g06927(.A1(new_n7926_), .A2(new_n7929_), .A3(new_n7928_), .ZN(new_n7930_));
  NOR3_X1    g06928(.A1(new_n7925_), .A2(new_n7930_), .A3(new_n7908_), .ZN(new_n7931_));
  XOR2_X1    g06929(.A1(new_n7900_), .A2(new_n7907_), .Z(new_n7932_));
  OAI21_X1   g06930(.A1(new_n7926_), .A2(new_n7928_), .B(new_n7929_), .ZN(new_n7933_));
  NAND3_X1   g06931(.A1(new_n7247_), .A2(new_n7271_), .A3(new_n7906_), .ZN(new_n7934_));
  NOR2_X1    g06932(.A1(new_n7923_), .A2(new_n7916_), .ZN(new_n7935_));
  NOR2_X1    g06933(.A1(new_n7921_), .A2(new_n7918_), .ZN(new_n7936_));
  NOR2_X1    g06934(.A1(new_n7935_), .A2(new_n7936_), .ZN(new_n7937_));
  AOI21_X1   g06935(.A1(new_n7228_), .A2(new_n7221_), .B(new_n7914_), .ZN(new_n7938_));
  INV_X1     g06936(.I(new_n7938_), .ZN(new_n7939_));
  NAND4_X1   g06937(.A1(new_n7937_), .A2(new_n7273_), .A3(new_n7934_), .A4(new_n7939_), .ZN(new_n7940_));
  AOI21_X1   g06938(.A1(new_n7940_), .A2(new_n7933_), .B(new_n7932_), .ZN(new_n7941_));
  OAI21_X1   g06939(.A1(new_n7941_), .A2(new_n7931_), .B(new_n7281_), .ZN(new_n7942_));
  NAND3_X1   g06940(.A1(new_n7937_), .A2(new_n7273_), .A3(new_n7917_), .ZN(new_n7943_));
  NAND3_X1   g06941(.A1(new_n7933_), .A2(new_n7943_), .A3(new_n7932_), .ZN(new_n7944_));
  NAND3_X1   g06942(.A1(new_n7924_), .A2(new_n7922_), .A3(new_n7934_), .ZN(new_n7945_));
  NOR3_X1    g06943(.A1(new_n7945_), .A2(new_n7926_), .A3(new_n7938_), .ZN(new_n7946_));
  OAI21_X1   g06944(.A1(new_n7925_), .A2(new_n7946_), .B(new_n7908_), .ZN(new_n7947_));
  NAND3_X1   g06945(.A1(new_n7947_), .A2(new_n7944_), .A3(new_n7449_), .ZN(new_n7948_));
  AOI21_X1   g06946(.A1(new_n7942_), .A2(new_n7948_), .B(new_n7899_), .ZN(new_n7949_));
  INV_X1     g06947(.I(new_n7862_), .ZN(new_n7950_));
  INV_X1     g06948(.I(new_n7878_), .ZN(new_n7951_));
  NOR4_X1    g06949(.A1(new_n7883_), .A2(new_n7950_), .A3(new_n7886_), .A4(new_n7951_), .ZN(new_n7952_));
  NOR3_X1    g06950(.A1(new_n7952_), .A2(new_n7896_), .A3(new_n7894_), .ZN(new_n7953_));
  NAND3_X1   g06951(.A1(new_n7195_), .A2(new_n7876_), .A3(new_n7895_), .ZN(new_n7954_));
  AOI21_X1   g06952(.A1(new_n7892_), .A2(new_n7954_), .B(new_n7882_), .ZN(new_n7955_));
  NOR2_X1    g06953(.A1(new_n7953_), .A2(new_n7955_), .ZN(new_n7956_));
  AOI21_X1   g06954(.A1(new_n7947_), .A2(new_n7944_), .B(new_n7449_), .ZN(new_n7957_));
  NOR3_X1    g06955(.A1(new_n7941_), .A2(new_n7931_), .A3(new_n7281_), .ZN(new_n7958_));
  NOR3_X1    g06956(.A1(new_n7958_), .A2(new_n7957_), .A3(new_n7956_), .ZN(new_n7959_));
  OAI21_X1   g06957(.A1(new_n7959_), .A2(new_n7949_), .B(new_n7448_), .ZN(new_n7960_));
  INV_X1     g06958(.I(new_n7448_), .ZN(new_n7961_));
  OAI21_X1   g06959(.A1(new_n7958_), .A2(new_n7957_), .B(new_n7956_), .ZN(new_n7962_));
  NAND3_X1   g06960(.A1(new_n7942_), .A2(new_n7948_), .A3(new_n7899_), .ZN(new_n7963_));
  NAND3_X1   g06961(.A1(new_n7962_), .A2(new_n7963_), .A3(new_n7961_), .ZN(new_n7964_));
  NOR4_X1    g06962(.A1(new_n7343_), .A2(new_n7345_), .A3(new_n7338_), .A4(new_n7334_), .ZN(new_n7965_));
  AOI21_X1   g06963(.A1(\A[35] ), .A2(\A[36] ), .B(\A[34] ), .ZN(new_n7966_));
  NOR2_X1    g06964(.A1(new_n7966_), .A2(new_n7335_), .ZN(new_n7967_));
  AOI21_X1   g06965(.A1(\A[32] ), .A2(\A[33] ), .B(\A[31] ), .ZN(new_n7968_));
  NOR2_X1    g06966(.A1(new_n7968_), .A2(new_n7324_), .ZN(new_n7969_));
  NOR2_X1    g06967(.A1(new_n7967_), .A2(new_n7969_), .ZN(new_n7970_));
  NOR4_X1    g06968(.A1(new_n7966_), .A2(new_n7968_), .A3(new_n7324_), .A4(new_n7335_), .ZN(new_n7971_));
  NOR2_X1    g06969(.A1(new_n7970_), .A2(new_n7971_), .ZN(new_n7972_));
  XNOR2_X1   g06970(.A1(new_n7965_), .A2(new_n7972_), .ZN(new_n7973_));
  NAND4_X1   g06971(.A1(new_n7286_), .A2(new_n7291_), .A3(new_n7313_), .A4(new_n7315_), .ZN(new_n7974_));
  AOI21_X1   g06972(.A1(new_n7293_), .A2(new_n7301_), .B(new_n7299_), .ZN(new_n7975_));
  AOI21_X1   g06973(.A1(\A[38] ), .A2(\A[39] ), .B(\A[37] ), .ZN(new_n7976_));
  NOR2_X1    g06974(.A1(new_n7976_), .A2(new_n7288_), .ZN(new_n7977_));
  XNOR2_X1   g06975(.A1(new_n7975_), .A2(new_n7977_), .ZN(new_n7978_));
  NAND2_X1   g06976(.A1(new_n7978_), .A2(new_n7974_), .ZN(new_n7979_));
  NOR4_X1    g06977(.A1(new_n7307_), .A2(new_n7309_), .A3(new_n7302_), .A4(new_n7298_), .ZN(new_n7980_));
  XOR2_X1    g06978(.A1(new_n7975_), .A2(new_n7977_), .Z(new_n7981_));
  NAND2_X1   g06979(.A1(new_n7981_), .A2(new_n7980_), .ZN(new_n7982_));
  NAND2_X1   g06980(.A1(new_n7979_), .A2(new_n7982_), .ZN(new_n7983_));
  AOI21_X1   g06981(.A1(new_n7354_), .A2(new_n7983_), .B(new_n7973_), .ZN(new_n7984_));
  NOR2_X1    g06982(.A1(new_n7981_), .A2(new_n7980_), .ZN(new_n7985_));
  NOR2_X1    g06983(.A1(new_n7978_), .A2(new_n7974_), .ZN(new_n7986_));
  NOR2_X1    g06984(.A1(new_n7986_), .A2(new_n7985_), .ZN(new_n7987_));
  NAND2_X1   g06985(.A1(new_n7975_), .A2(new_n7977_), .ZN(new_n7988_));
  INV_X1     g06986(.I(new_n7988_), .ZN(new_n7989_));
  NOR2_X1    g06987(.A1(new_n7975_), .A2(new_n7977_), .ZN(new_n7990_));
  INV_X1     g06988(.I(new_n7990_), .ZN(new_n7991_));
  OAI21_X1   g06989(.A1(new_n7980_), .A2(new_n7989_), .B(new_n7991_), .ZN(new_n7992_));
  AOI21_X1   g06990(.A1(new_n7974_), .A2(new_n7988_), .B(new_n7990_), .ZN(new_n7993_));
  AND3_X2    g06991(.A1(new_n7346_), .A2(new_n7339_), .A3(new_n7971_), .Z(new_n7994_));
  AOI21_X1   g06992(.A1(new_n7439_), .A2(new_n7993_), .B(new_n7994_), .ZN(new_n7995_));
  NAND4_X1   g06993(.A1(new_n7995_), .A2(new_n7438_), .A3(new_n7987_), .A4(new_n7992_), .ZN(new_n7996_));
  NAND2_X1   g06994(.A1(new_n7983_), .A2(new_n7354_), .ZN(new_n7997_));
  NAND4_X1   g06995(.A1(new_n7439_), .A2(new_n7440_), .A3(new_n7979_), .A4(new_n7982_), .ZN(new_n7998_));
  NAND2_X1   g06996(.A1(new_n7997_), .A2(new_n7998_), .ZN(new_n7999_));
  AOI22_X1   g06997(.A1(new_n7999_), .A2(new_n7973_), .B1(new_n7996_), .B2(new_n7984_), .ZN(new_n8000_));
  NAND4_X1   g06998(.A1(new_n7398_), .A2(new_n7403_), .A3(new_n7425_), .A4(new_n7427_), .ZN(new_n8001_));
  AOI21_X1   g06999(.A1(\A[47] ), .A2(\A[48] ), .B(\A[46] ), .ZN(new_n8002_));
  AOI21_X1   g07000(.A1(\A[44] ), .A2(\A[45] ), .B(\A[43] ), .ZN(new_n8003_));
  OAI22_X1   g07001(.A1(new_n7400_), .A2(new_n8003_), .B1(new_n8002_), .B2(new_n7411_), .ZN(new_n8004_));
  NOR4_X1    g07002(.A1(new_n8002_), .A2(new_n8003_), .A3(new_n7400_), .A4(new_n7411_), .ZN(new_n8005_));
  INV_X1     g07003(.I(new_n8005_), .ZN(new_n8006_));
  NAND2_X1   g07004(.A1(new_n8006_), .A2(new_n8004_), .ZN(new_n8007_));
  XOR2_X1    g07005(.A1(new_n8001_), .A2(new_n8007_), .Z(new_n8008_));
  NOR4_X1    g07006(.A1(new_n7383_), .A2(new_n7385_), .A3(new_n7378_), .A4(new_n7374_), .ZN(new_n8009_));
  AOI21_X1   g07007(.A1(new_n7369_), .A2(new_n7377_), .B(new_n7375_), .ZN(new_n8010_));
  AOI21_X1   g07008(.A1(\A[50] ), .A2(\A[51] ), .B(\A[49] ), .ZN(new_n8011_));
  NOR2_X1    g07009(.A1(new_n8011_), .A2(new_n7364_), .ZN(new_n8012_));
  XOR2_X1    g07010(.A1(new_n8010_), .A2(new_n8012_), .Z(new_n8013_));
  NOR2_X1    g07011(.A1(new_n8013_), .A2(new_n8009_), .ZN(new_n8014_));
  NAND4_X1   g07012(.A1(new_n7362_), .A2(new_n7367_), .A3(new_n7389_), .A4(new_n7391_), .ZN(new_n8015_));
  XNOR2_X1   g07013(.A1(new_n8010_), .A2(new_n8012_), .ZN(new_n8016_));
  NOR2_X1    g07014(.A1(new_n8016_), .A2(new_n8015_), .ZN(new_n8017_));
  NOR2_X1    g07015(.A1(new_n8017_), .A2(new_n8014_), .ZN(new_n8018_));
  NOR2_X1    g07016(.A1(new_n8018_), .A2(new_n7446_), .ZN(new_n8019_));
  NAND2_X1   g07017(.A1(new_n8016_), .A2(new_n8015_), .ZN(new_n8020_));
  NAND2_X1   g07018(.A1(new_n8013_), .A2(new_n8009_), .ZN(new_n8021_));
  NAND2_X1   g07019(.A1(new_n8020_), .A2(new_n8021_), .ZN(new_n8022_));
  NOR2_X1    g07020(.A1(new_n8022_), .A2(new_n7430_), .ZN(new_n8023_));
  NOR3_X1    g07021(.A1(new_n8023_), .A2(new_n8019_), .A3(new_n8008_), .ZN(new_n8024_));
  NOR4_X1    g07022(.A1(new_n7419_), .A2(new_n7421_), .A3(new_n7414_), .A4(new_n7410_), .ZN(new_n8025_));
  XOR2_X1    g07023(.A1(new_n8025_), .A2(new_n8007_), .Z(new_n8026_));
  NAND2_X1   g07024(.A1(new_n8022_), .A2(new_n7430_), .ZN(new_n8027_));
  NAND2_X1   g07025(.A1(new_n8025_), .A2(new_n8005_), .ZN(new_n8028_));
  NAND2_X1   g07026(.A1(new_n8010_), .A2(new_n8012_), .ZN(new_n8029_));
  AOI21_X1   g07027(.A1(new_n7368_), .A2(new_n7392_), .B(new_n8029_), .ZN(new_n8030_));
  INV_X1     g07028(.I(new_n8030_), .ZN(new_n8031_));
  NAND4_X1   g07029(.A1(new_n8018_), .A2(new_n7446_), .A3(new_n8028_), .A4(new_n8031_), .ZN(new_n8032_));
  AOI21_X1   g07030(.A1(new_n8032_), .A2(new_n8027_), .B(new_n8026_), .ZN(new_n8033_));
  OAI21_X1   g07031(.A1(new_n8033_), .A2(new_n8024_), .B(new_n7447_), .ZN(new_n8034_));
  NAND2_X1   g07032(.A1(new_n8018_), .A2(new_n7446_), .ZN(new_n8035_));
  NAND3_X1   g07033(.A1(new_n8027_), .A2(new_n8035_), .A3(new_n8026_), .ZN(new_n8036_));
  NAND3_X1   g07034(.A1(new_n8020_), .A2(new_n8021_), .A3(new_n8028_), .ZN(new_n8037_));
  NOR3_X1    g07035(.A1(new_n8037_), .A2(new_n7430_), .A3(new_n8030_), .ZN(new_n8038_));
  OAI21_X1   g07036(.A1(new_n8038_), .A2(new_n8019_), .B(new_n8008_), .ZN(new_n8039_));
  NAND3_X1   g07037(.A1(new_n8039_), .A2(new_n8036_), .A3(new_n7451_), .ZN(new_n8040_));
  NAND3_X1   g07038(.A1(new_n8034_), .A2(new_n8040_), .A3(new_n8000_), .ZN(new_n8041_));
  XOR2_X1    g07039(.A1(new_n7965_), .A2(new_n7972_), .Z(new_n8042_));
  OAI21_X1   g07040(.A1(new_n7438_), .A2(new_n7987_), .B(new_n8042_), .ZN(new_n8043_));
  NAND2_X1   g07041(.A1(new_n7965_), .A2(new_n7971_), .ZN(new_n8044_));
  OAI21_X1   g07042(.A1(new_n7355_), .A2(new_n7992_), .B(new_n8044_), .ZN(new_n8045_));
  NOR3_X1    g07043(.A1(new_n7998_), .A2(new_n8045_), .A3(new_n7993_), .ZN(new_n8046_));
  AOI22_X1   g07044(.A1(new_n7439_), .A2(new_n7440_), .B1(new_n7979_), .B2(new_n7982_), .ZN(new_n8047_));
  NOR4_X1    g07045(.A1(new_n7355_), .A2(new_n7356_), .A3(new_n7985_), .A4(new_n7986_), .ZN(new_n8048_));
  NOR2_X1    g07046(.A1(new_n8047_), .A2(new_n8048_), .ZN(new_n8049_));
  OAI22_X1   g07047(.A1(new_n8042_), .A2(new_n8049_), .B1(new_n8046_), .B2(new_n8043_), .ZN(new_n8050_));
  AOI21_X1   g07048(.A1(new_n8039_), .A2(new_n8036_), .B(new_n7451_), .ZN(new_n8051_));
  NOR3_X1    g07049(.A1(new_n8033_), .A2(new_n8024_), .A3(new_n7447_), .ZN(new_n8052_));
  OAI21_X1   g07050(.A1(new_n8052_), .A2(new_n8051_), .B(new_n8050_), .ZN(new_n8053_));
  NAND2_X1   g07051(.A1(new_n8053_), .A2(new_n8041_), .ZN(new_n8054_));
  AOI21_X1   g07052(.A1(new_n7960_), .A2(new_n7964_), .B(new_n8054_), .ZN(new_n8055_));
  AOI21_X1   g07053(.A1(new_n7962_), .A2(new_n7963_), .B(new_n7961_), .ZN(new_n8056_));
  NOR3_X1    g07054(.A1(new_n7959_), .A2(new_n7949_), .A3(new_n7448_), .ZN(new_n8057_));
  NOR3_X1    g07055(.A1(new_n8052_), .A2(new_n8051_), .A3(new_n8050_), .ZN(new_n8058_));
  AOI21_X1   g07056(.A1(new_n8034_), .A2(new_n8040_), .B(new_n8000_), .ZN(new_n8059_));
  NOR2_X1    g07057(.A1(new_n8058_), .A2(new_n8059_), .ZN(new_n8060_));
  NOR3_X1    g07058(.A1(new_n8056_), .A2(new_n8057_), .A3(new_n8060_), .ZN(new_n8061_));
  OAI21_X1   g07059(.A1(new_n8061_), .A2(new_n8055_), .B(new_n7855_), .ZN(new_n8062_));
  OAI21_X1   g07060(.A1(new_n8056_), .A2(new_n8057_), .B(new_n8060_), .ZN(new_n8063_));
  NAND3_X1   g07061(.A1(new_n7960_), .A2(new_n7964_), .A3(new_n8054_), .ZN(new_n8064_));
  NAND3_X1   g07062(.A1(new_n8063_), .A2(new_n8064_), .A3(new_n7854_), .ZN(new_n8065_));
  AOI21_X1   g07063(.A1(new_n8062_), .A2(new_n8065_), .B(new_n7853_), .ZN(new_n8066_));
  NOR3_X1    g07064(.A1(new_n7850_), .A2(new_n7851_), .A3(new_n7849_), .ZN(new_n8067_));
  AOI21_X1   g07065(.A1(new_n7845_), .A2(new_n7841_), .B(new_n7798_), .ZN(new_n8068_));
  NOR2_X1    g07066(.A1(new_n8067_), .A2(new_n8068_), .ZN(new_n8069_));
  AOI21_X1   g07067(.A1(new_n8063_), .A2(new_n8064_), .B(new_n7854_), .ZN(new_n8070_));
  NOR3_X1    g07068(.A1(new_n8061_), .A2(new_n8055_), .A3(new_n7855_), .ZN(new_n8071_));
  NOR3_X1    g07069(.A1(new_n8071_), .A2(new_n8070_), .A3(new_n8069_), .ZN(new_n8072_));
  OAI21_X1   g07070(.A1(new_n8072_), .A2(new_n8066_), .B(new_n7698_), .ZN(new_n8073_));
  NOR3_X1    g07071(.A1(new_n8072_), .A2(new_n8066_), .A3(new_n7698_), .ZN(new_n8074_));
  NOR3_X1    g07072(.A1(new_n7046_), .A2(new_n6994_), .A3(new_n7007_), .ZN(new_n8075_));
  AOI21_X1   g07073(.A1(\A[971] ), .A2(\A[972] ), .B(\A[970] ), .ZN(new_n8076_));
  NOR2_X1    g07074(.A1(new_n8076_), .A2(new_n7025_), .ZN(new_n8077_));
  AOI21_X1   g07075(.A1(\A[968] ), .A2(\A[969] ), .B(\A[967] ), .ZN(new_n8078_));
  NOR2_X1    g07076(.A1(new_n8078_), .A2(new_n7015_), .ZN(new_n8079_));
  NAND3_X1   g07077(.A1(new_n7028_), .A2(new_n8077_), .A3(new_n8079_), .ZN(new_n8080_));
  AOI21_X1   g07078(.A1(new_n6988_), .A2(new_n6990_), .B(new_n6989_), .ZN(new_n8081_));
  AOI21_X1   g07079(.A1(new_n6977_), .A2(new_n6979_), .B(new_n6978_), .ZN(new_n8082_));
  XOR2_X1    g07080(.A1(new_n8081_), .A2(new_n8082_), .Z(new_n8083_));
  NAND2_X1   g07081(.A1(new_n8083_), .A2(new_n7042_), .ZN(new_n8084_));
  INV_X1     g07082(.I(new_n8082_), .ZN(new_n8085_));
  NAND2_X1   g07083(.A1(new_n8085_), .A2(new_n8081_), .ZN(new_n8086_));
  INV_X1     g07084(.I(new_n8081_), .ZN(new_n8087_));
  NAND2_X1   g07085(.A1(new_n8087_), .A2(new_n8082_), .ZN(new_n8088_));
  NAND4_X1   g07086(.A1(new_n7000_), .A2(new_n8086_), .A3(new_n8088_), .A4(new_n7006_), .ZN(new_n8089_));
  NAND2_X1   g07087(.A1(new_n8084_), .A2(new_n8089_), .ZN(new_n8090_));
  NAND2_X1   g07088(.A1(new_n8081_), .A2(new_n8082_), .ZN(new_n8091_));
  INV_X1     g07089(.I(new_n8091_), .ZN(new_n8092_));
  NAND2_X1   g07090(.A1(new_n7043_), .A2(new_n8092_), .ZN(new_n8093_));
  NAND4_X1   g07091(.A1(new_n8090_), .A2(new_n8075_), .A3(new_n8080_), .A4(new_n8093_), .ZN(new_n8094_));
  OAI22_X1   g07092(.A1(new_n7015_), .A2(new_n8078_), .B1(new_n8076_), .B2(new_n7025_), .ZN(new_n8095_));
  NAND2_X1   g07093(.A1(new_n8077_), .A2(new_n8079_), .ZN(new_n8096_));
  NAND2_X1   g07094(.A1(new_n8096_), .A2(new_n8095_), .ZN(new_n8097_));
  XOR2_X1    g07095(.A1(new_n7028_), .A2(new_n8097_), .Z(new_n8098_));
  AOI22_X1   g07096(.A1(new_n8086_), .A2(new_n8088_), .B1(new_n7000_), .B2(new_n7006_), .ZN(new_n8099_));
  NOR2_X1    g07097(.A1(new_n8083_), .A2(new_n7042_), .ZN(new_n8100_));
  NOR2_X1    g07098(.A1(new_n8100_), .A2(new_n8099_), .ZN(new_n8101_));
  NAND4_X1   g07099(.A1(new_n7040_), .A2(new_n8080_), .A3(new_n7042_), .A4(new_n7043_), .ZN(new_n8102_));
  AOI21_X1   g07100(.A1(new_n8102_), .A2(new_n8101_), .B(new_n8098_), .ZN(new_n8103_));
  NAND2_X1   g07101(.A1(new_n8102_), .A2(new_n8101_), .ZN(new_n8104_));
  INV_X1     g07102(.I(new_n8077_), .ZN(new_n8105_));
  NOR4_X1    g07103(.A1(new_n7044_), .A2(new_n7015_), .A3(new_n8105_), .A4(new_n8078_), .ZN(new_n8106_));
  NOR4_X1    g07104(.A1(new_n8106_), .A2(new_n7046_), .A3(new_n6994_), .A4(new_n7007_), .ZN(new_n8107_));
  NAND2_X1   g07105(.A1(new_n8107_), .A2(new_n8090_), .ZN(new_n8108_));
  NAND2_X1   g07106(.A1(new_n8108_), .A2(new_n8104_), .ZN(new_n8109_));
  AOI22_X1   g07107(.A1(new_n8109_), .A2(new_n8098_), .B1(new_n8094_), .B2(new_n8103_), .ZN(new_n8110_));
  NAND2_X1   g07108(.A1(new_n7048_), .A2(new_n7117_), .ZN(new_n8111_));
  AOI21_X1   g07109(.A1(new_n7097_), .A2(new_n7098_), .B(new_n7100_), .ZN(new_n8112_));
  AOI21_X1   g07110(.A1(new_n7087_), .A2(new_n7088_), .B(new_n7090_), .ZN(new_n8113_));
  XOR2_X1    g07111(.A1(new_n8112_), .A2(new_n8113_), .Z(new_n8114_));
  XOR2_X1    g07112(.A1(new_n8114_), .A2(new_n7102_), .Z(new_n8115_));
  NAND4_X1   g07113(.A1(new_n7080_), .A2(new_n7113_), .A3(new_n7069_), .A4(new_n7102_), .ZN(new_n8116_));
  NOR4_X1    g07114(.A1(new_n7072_), .A2(new_n7074_), .A3(new_n7079_), .A4(new_n7077_), .ZN(new_n8117_));
  AOI21_X1   g07115(.A1(new_n7064_), .A2(new_n7066_), .B(new_n7065_), .ZN(new_n8118_));
  AOI21_X1   g07116(.A1(\A[986] ), .A2(\A[987] ), .B(\A[985] ), .ZN(new_n8119_));
  NOR2_X1    g07117(.A1(new_n8119_), .A2(new_n7055_), .ZN(new_n8120_));
  NAND2_X1   g07118(.A1(new_n8118_), .A2(new_n8120_), .ZN(new_n8121_));
  INV_X1     g07119(.I(new_n8121_), .ZN(new_n8122_));
  NAND2_X1   g07120(.A1(new_n8117_), .A2(new_n8122_), .ZN(new_n8123_));
  NOR4_X1    g07121(.A1(new_n7105_), .A2(new_n7107_), .A3(new_n7112_), .A4(new_n7110_), .ZN(new_n8124_));
  NAND3_X1   g07122(.A1(new_n8124_), .A2(new_n8112_), .A3(new_n8113_), .ZN(new_n8125_));
  NAND2_X1   g07123(.A1(new_n8125_), .A2(new_n8123_), .ZN(new_n8126_));
  XNOR2_X1   g07124(.A1(new_n8118_), .A2(new_n8120_), .ZN(new_n8127_));
  NOR2_X1    g07125(.A1(new_n8127_), .A2(new_n7069_), .ZN(new_n8128_));
  XOR2_X1    g07126(.A1(new_n8118_), .A2(new_n8120_), .Z(new_n8129_));
  NOR2_X1    g07127(.A1(new_n8129_), .A2(new_n8117_), .ZN(new_n8130_));
  OAI22_X1   g07128(.A1(new_n8126_), .A2(new_n8116_), .B1(new_n8128_), .B2(new_n8130_), .ZN(new_n8131_));
  AOI22_X1   g07129(.A1(new_n7053_), .A2(new_n7058_), .B1(new_n7063_), .B2(new_n7068_), .ZN(new_n8132_));
  AOI22_X1   g07130(.A1(new_n7086_), .A2(new_n7091_), .B1(new_n7096_), .B2(new_n7101_), .ZN(new_n8133_));
  NOR4_X1    g07131(.A1(new_n8117_), .A2(new_n8132_), .A3(new_n8133_), .A4(new_n8124_), .ZN(new_n8134_));
  NOR2_X1    g07132(.A1(new_n7069_), .A2(new_n8121_), .ZN(new_n8135_));
  INV_X1     g07133(.I(new_n8112_), .ZN(new_n8136_));
  INV_X1     g07134(.I(new_n8113_), .ZN(new_n8137_));
  NOR3_X1    g07135(.A1(new_n7102_), .A2(new_n8136_), .A3(new_n8137_), .ZN(new_n8138_));
  NOR2_X1    g07136(.A1(new_n8138_), .A2(new_n8135_), .ZN(new_n8139_));
  NOR2_X1    g07137(.A1(new_n8128_), .A2(new_n8130_), .ZN(new_n8140_));
  NAND3_X1   g07138(.A1(new_n8140_), .A2(new_n8139_), .A3(new_n8134_), .ZN(new_n8141_));
  NAND3_X1   g07139(.A1(new_n8141_), .A2(new_n8131_), .A3(new_n8115_), .ZN(new_n8142_));
  XOR2_X1    g07140(.A1(new_n8114_), .A2(new_n8124_), .Z(new_n8143_));
  NAND2_X1   g07141(.A1(new_n8129_), .A2(new_n8117_), .ZN(new_n8144_));
  NAND2_X1   g07142(.A1(new_n8127_), .A2(new_n7069_), .ZN(new_n8145_));
  AOI22_X1   g07143(.A1(new_n8139_), .A2(new_n8134_), .B1(new_n8144_), .B2(new_n8145_), .ZN(new_n8146_));
  NAND2_X1   g07144(.A1(new_n8145_), .A2(new_n8144_), .ZN(new_n8147_));
  NOR2_X1    g07145(.A1(new_n8132_), .A2(new_n8121_), .ZN(new_n8148_));
  NOR4_X1    g07146(.A1(new_n8147_), .A2(new_n8116_), .A3(new_n8138_), .A4(new_n8148_), .ZN(new_n8149_));
  OAI21_X1   g07147(.A1(new_n8149_), .A2(new_n8146_), .B(new_n8143_), .ZN(new_n8150_));
  AOI21_X1   g07148(.A1(new_n8150_), .A2(new_n8142_), .B(new_n8111_), .ZN(new_n8151_));
  AOI22_X1   g07149(.A1(new_n7041_), .A2(new_n7047_), .B1(new_n7114_), .B2(new_n7116_), .ZN(new_n8152_));
  NOR3_X1    g07150(.A1(new_n8147_), .A2(new_n8126_), .A3(new_n8116_), .ZN(new_n8153_));
  NOR3_X1    g07151(.A1(new_n8146_), .A2(new_n8153_), .A3(new_n8143_), .ZN(new_n8154_));
  INV_X1     g07152(.I(new_n8148_), .ZN(new_n8155_));
  NAND4_X1   g07153(.A1(new_n8140_), .A2(new_n8134_), .A3(new_n8125_), .A4(new_n8155_), .ZN(new_n8156_));
  AOI21_X1   g07154(.A1(new_n8156_), .A2(new_n8131_), .B(new_n8115_), .ZN(new_n8157_));
  NOR3_X1    g07155(.A1(new_n8157_), .A2(new_n8154_), .A3(new_n8152_), .ZN(new_n8158_));
  OAI21_X1   g07156(.A1(new_n8158_), .A2(new_n8151_), .B(new_n8110_), .ZN(new_n8159_));
  NAND2_X1   g07157(.A1(new_n8103_), .A2(new_n8094_), .ZN(new_n8160_));
  NOR2_X1    g07158(.A1(new_n8107_), .A2(new_n8090_), .ZN(new_n8161_));
  NOR2_X1    g07159(.A1(new_n8102_), .A2(new_n8101_), .ZN(new_n8162_));
  OAI21_X1   g07160(.A1(new_n8161_), .A2(new_n8162_), .B(new_n8098_), .ZN(new_n8163_));
  NAND2_X1   g07161(.A1(new_n8163_), .A2(new_n8160_), .ZN(new_n8164_));
  OAI21_X1   g07162(.A1(new_n8157_), .A2(new_n8154_), .B(new_n8152_), .ZN(new_n8165_));
  NAND3_X1   g07163(.A1(new_n8150_), .A2(new_n8142_), .A3(new_n8111_), .ZN(new_n8166_));
  NAND3_X1   g07164(.A1(new_n8165_), .A2(new_n8166_), .A3(new_n8164_), .ZN(new_n8167_));
  NAND2_X1   g07165(.A1(new_n8159_), .A2(new_n8167_), .ZN(new_n8168_));
  XNOR2_X1   g07166(.A1(new_n6964_), .A2(new_n6966_), .ZN(new_n8169_));
  XNOR2_X1   g07167(.A1(new_n8169_), .A2(new_n6928_), .ZN(new_n8170_));
  NAND3_X1   g07168(.A1(new_n6952_), .A2(new_n6928_), .A3(new_n6930_), .ZN(new_n8171_));
  NOR2_X1    g07169(.A1(new_n6951_), .A2(new_n6941_), .ZN(new_n8172_));
  AOI21_X1   g07170(.A1(\A[953] ), .A2(\A[954] ), .B(\A[952] ), .ZN(new_n8173_));
  NOR2_X1    g07171(.A1(new_n8173_), .A2(new_n6949_), .ZN(new_n8174_));
  AOI21_X1   g07172(.A1(new_n6936_), .A2(new_n6937_), .B(new_n6939_), .ZN(new_n8175_));
  XOR2_X1    g07173(.A1(new_n8175_), .A2(new_n8174_), .Z(new_n8176_));
  XNOR2_X1   g07174(.A1(new_n8172_), .A2(new_n8176_), .ZN(new_n8177_));
  AOI21_X1   g07175(.A1(new_n8177_), .A2(new_n8171_), .B(new_n8170_), .ZN(new_n8178_));
  INV_X1     g07176(.I(new_n6928_), .ZN(new_n8179_));
  NOR3_X1    g07177(.A1(new_n6963_), .A2(new_n8179_), .A3(new_n6929_), .ZN(new_n8180_));
  AND2_X2    g07178(.A1(new_n8175_), .A2(new_n8174_), .Z(new_n8181_));
  OAI21_X1   g07179(.A1(new_n6955_), .A2(new_n6962_), .B(new_n8181_), .ZN(new_n8182_));
  NAND3_X1   g07180(.A1(new_n8180_), .A2(new_n8176_), .A3(new_n8182_), .ZN(new_n8183_));
  NAND2_X1   g07181(.A1(new_n8177_), .A2(new_n8171_), .ZN(new_n8184_));
  XOR2_X1    g07182(.A1(new_n8172_), .A2(new_n8176_), .Z(new_n8185_));
  NAND2_X1   g07183(.A1(new_n8185_), .A2(new_n8180_), .ZN(new_n8186_));
  NAND2_X1   g07184(.A1(new_n8184_), .A2(new_n8186_), .ZN(new_n8187_));
  AOI22_X1   g07185(.A1(new_n8187_), .A2(new_n8170_), .B1(new_n8178_), .B2(new_n8183_), .ZN(new_n8188_));
  NOR3_X1    g07186(.A1(new_n6970_), .A2(new_n6892_), .A3(new_n6906_), .ZN(new_n8189_));
  INV_X1     g07187(.I(new_n6902_), .ZN(new_n8190_));
  NAND2_X1   g07188(.A1(new_n8190_), .A2(new_n6904_), .ZN(new_n8191_));
  NAND2_X1   g07189(.A1(new_n6905_), .A2(new_n6902_), .ZN(new_n8192_));
  NAND2_X1   g07190(.A1(new_n8192_), .A2(new_n8191_), .ZN(new_n8193_));
  XNOR2_X1   g07191(.A1(new_n8193_), .A2(new_n6864_), .ZN(new_n8194_));
  NAND3_X1   g07192(.A1(new_n6901_), .A2(new_n6864_), .A3(new_n6867_), .ZN(new_n8195_));
  NAND3_X1   g07193(.A1(new_n6879_), .A2(new_n6884_), .A3(new_n6889_), .ZN(new_n8196_));
  AOI21_X1   g07194(.A1(new_n6885_), .A2(new_n6886_), .B(new_n6888_), .ZN(new_n8197_));
  AOI21_X1   g07195(.A1(new_n6869_), .A2(new_n6875_), .B(new_n6876_), .ZN(new_n8198_));
  XOR2_X1    g07196(.A1(new_n8197_), .A2(new_n8198_), .Z(new_n8199_));
  XOR2_X1    g07197(.A1(new_n8196_), .A2(new_n8199_), .Z(new_n8200_));
  INV_X1     g07198(.I(new_n8197_), .ZN(new_n8201_));
  INV_X1     g07199(.I(new_n8198_), .ZN(new_n8202_));
  NOR3_X1    g07200(.A1(new_n6891_), .A2(new_n8201_), .A3(new_n8202_), .ZN(new_n8203_));
  OAI21_X1   g07201(.A1(new_n8203_), .A2(new_n8200_), .B(new_n8195_), .ZN(new_n8204_));
  NOR3_X1    g07202(.A1(new_n6864_), .A2(new_n8190_), .A3(new_n6904_), .ZN(new_n8205_));
  NOR3_X1    g07203(.A1(new_n6891_), .A2(new_n6868_), .A3(new_n8205_), .ZN(new_n8206_));
  NAND3_X1   g07204(.A1(new_n6901_), .A2(new_n8197_), .A3(new_n8198_), .ZN(new_n8207_));
  NAND3_X1   g07205(.A1(new_n8206_), .A2(new_n8199_), .A3(new_n8207_), .ZN(new_n8208_));
  AOI21_X1   g07206(.A1(new_n8204_), .A2(new_n8208_), .B(new_n8194_), .ZN(new_n8209_));
  XOR2_X1    g07207(.A1(new_n8193_), .A2(new_n6864_), .Z(new_n8210_));
  NOR2_X1    g07208(.A1(new_n6899_), .A2(new_n6890_), .ZN(new_n8211_));
  XOR2_X1    g07209(.A1(new_n8211_), .A2(new_n8199_), .Z(new_n8212_));
  AOI21_X1   g07210(.A1(new_n8212_), .A2(new_n8207_), .B(new_n8206_), .ZN(new_n8213_));
  NOR3_X1    g07211(.A1(new_n8203_), .A2(new_n8200_), .A3(new_n8195_), .ZN(new_n8214_));
  NOR3_X1    g07212(.A1(new_n8213_), .A2(new_n8214_), .A3(new_n8210_), .ZN(new_n8215_));
  OAI21_X1   g07213(.A1(new_n8215_), .A2(new_n8209_), .B(new_n8189_), .ZN(new_n8216_));
  NAND3_X1   g07214(.A1(new_n6907_), .A2(new_n6953_), .A3(new_n6969_), .ZN(new_n8217_));
  XNOR2_X1   g07215(.A1(new_n8197_), .A2(new_n8198_), .ZN(new_n8218_));
  NOR3_X1    g07216(.A1(new_n8203_), .A2(new_n8195_), .A3(new_n8218_), .ZN(new_n8219_));
  OAI21_X1   g07217(.A1(new_n8213_), .A2(new_n8219_), .B(new_n8210_), .ZN(new_n8220_));
  NAND3_X1   g07218(.A1(new_n8206_), .A2(new_n8212_), .A3(new_n8207_), .ZN(new_n8221_));
  NAND3_X1   g07219(.A1(new_n8204_), .A2(new_n8221_), .A3(new_n8194_), .ZN(new_n8222_));
  NAND3_X1   g07220(.A1(new_n8220_), .A2(new_n8222_), .A3(new_n8217_), .ZN(new_n8223_));
  NAND3_X1   g07221(.A1(new_n8216_), .A2(new_n8223_), .A3(new_n8188_), .ZN(new_n8224_));
  XOR2_X1    g07222(.A1(new_n8169_), .A2(new_n6928_), .Z(new_n8225_));
  OAI21_X1   g07223(.A1(new_n8180_), .A2(new_n8185_), .B(new_n8225_), .ZN(new_n8226_));
  NAND2_X1   g07224(.A1(new_n8182_), .A2(new_n8176_), .ZN(new_n8227_));
  NOR2_X1    g07225(.A1(new_n8171_), .A2(new_n8227_), .ZN(new_n8228_));
  NOR2_X1    g07226(.A1(new_n8185_), .A2(new_n8180_), .ZN(new_n8229_));
  NOR2_X1    g07227(.A1(new_n8177_), .A2(new_n8171_), .ZN(new_n8230_));
  NOR2_X1    g07228(.A1(new_n8230_), .A2(new_n8229_), .ZN(new_n8231_));
  OAI22_X1   g07229(.A1(new_n8231_), .A2(new_n8225_), .B1(new_n8226_), .B2(new_n8228_), .ZN(new_n8232_));
  AOI21_X1   g07230(.A1(new_n8220_), .A2(new_n8222_), .B(new_n8217_), .ZN(new_n8233_));
  NOR3_X1    g07231(.A1(new_n8215_), .A2(new_n8209_), .A3(new_n8189_), .ZN(new_n8234_));
  OAI21_X1   g07232(.A1(new_n8234_), .A2(new_n8233_), .B(new_n8232_), .ZN(new_n8235_));
  NAND3_X1   g07233(.A1(new_n8168_), .A2(new_n8235_), .A3(new_n8224_), .ZN(new_n8236_));
  AND2_X2    g07234(.A1(new_n8159_), .A2(new_n8167_), .Z(new_n8237_));
  NAND2_X1   g07235(.A1(new_n8235_), .A2(new_n8224_), .ZN(new_n8238_));
  NAND2_X1   g07236(.A1(new_n8238_), .A2(new_n8237_), .ZN(new_n8239_));
  NAND3_X1   g07237(.A1(new_n8239_), .A2(new_n7120_), .A3(new_n8236_), .ZN(new_n8240_));
  NAND2_X1   g07238(.A1(new_n8239_), .A2(new_n8236_), .ZN(new_n8241_));
  NAND2_X1   g07239(.A1(new_n8241_), .A2(new_n7119_), .ZN(new_n8242_));
  NAND2_X1   g07240(.A1(new_n8242_), .A2(new_n8240_), .ZN(new_n8243_));
  AOI21_X1   g07241(.A1(new_n8073_), .A2(new_n8243_), .B(new_n8074_), .ZN(new_n8244_));
  AOI21_X1   g07242(.A1(new_n8224_), .A2(new_n8235_), .B(new_n8168_), .ZN(new_n8245_));
  AOI21_X1   g07243(.A1(new_n7119_), .A2(new_n8236_), .B(new_n8245_), .ZN(new_n8246_));
  OAI21_X1   g07244(.A1(new_n8188_), .A2(new_n8233_), .B(new_n8223_), .ZN(new_n8247_));
  AOI21_X1   g07245(.A1(new_n8204_), .A2(new_n8210_), .B(new_n8219_), .ZN(new_n8248_));
  NAND2_X1   g07246(.A1(new_n8211_), .A2(new_n8198_), .ZN(new_n8249_));
  OAI21_X1   g07247(.A1(new_n8211_), .A2(new_n8198_), .B(new_n8197_), .ZN(new_n8250_));
  INV_X1     g07248(.I(new_n8191_), .ZN(new_n8251_));
  AOI21_X1   g07249(.A1(new_n6864_), .A2(new_n8192_), .B(new_n8251_), .ZN(new_n8252_));
  INV_X1     g07250(.I(new_n8252_), .ZN(new_n8253_));
  NAND3_X1   g07251(.A1(new_n8253_), .A2(new_n8249_), .A3(new_n8250_), .ZN(new_n8254_));
  NAND2_X1   g07252(.A1(new_n8250_), .A2(new_n8249_), .ZN(new_n8255_));
  NAND2_X1   g07253(.A1(new_n8255_), .A2(new_n8252_), .ZN(new_n8256_));
  NAND2_X1   g07254(.A1(new_n8254_), .A2(new_n8256_), .ZN(new_n8257_));
  NOR2_X1    g07255(.A1(new_n8248_), .A2(new_n8257_), .ZN(new_n8258_));
  NAND2_X1   g07256(.A1(new_n8212_), .A2(new_n8207_), .ZN(new_n8259_));
  AOI21_X1   g07257(.A1(new_n8259_), .A2(new_n8195_), .B(new_n8194_), .ZN(new_n8260_));
  NOR2_X1    g07258(.A1(new_n8255_), .A2(new_n8252_), .ZN(new_n8261_));
  AOI21_X1   g07259(.A1(new_n8249_), .A2(new_n8250_), .B(new_n8253_), .ZN(new_n8262_));
  NOR2_X1    g07260(.A1(new_n8262_), .A2(new_n8261_), .ZN(new_n8263_));
  NOR3_X1    g07261(.A1(new_n8260_), .A2(new_n8263_), .A3(new_n8219_), .ZN(new_n8264_));
  NOR2_X1    g07262(.A1(new_n8175_), .A2(new_n8174_), .ZN(new_n8265_));
  INV_X1     g07263(.I(new_n8265_), .ZN(new_n8266_));
  OAI21_X1   g07264(.A1(new_n8172_), .A2(new_n8181_), .B(new_n8266_), .ZN(new_n8267_));
  NOR2_X1    g07265(.A1(new_n6964_), .A2(new_n6966_), .ZN(new_n8268_));
  NOR2_X1    g07266(.A1(new_n6965_), .A2(new_n6967_), .ZN(new_n8269_));
  NOR2_X1    g07267(.A1(new_n8179_), .A2(new_n8269_), .ZN(new_n8270_));
  NOR2_X1    g07268(.A1(new_n8270_), .A2(new_n8268_), .ZN(new_n8271_));
  NOR3_X1    g07269(.A1(new_n8178_), .A2(new_n8228_), .A3(new_n8271_), .ZN(new_n8272_));
  INV_X1     g07270(.I(new_n8271_), .ZN(new_n8273_));
  AOI21_X1   g07271(.A1(new_n8226_), .A2(new_n8183_), .B(new_n8273_), .ZN(new_n8274_));
  NOR3_X1    g07272(.A1(new_n8272_), .A2(new_n8274_), .A3(new_n8267_), .ZN(new_n8275_));
  INV_X1     g07273(.I(new_n8267_), .ZN(new_n8276_));
  NAND3_X1   g07274(.A1(new_n8226_), .A2(new_n8183_), .A3(new_n8273_), .ZN(new_n8277_));
  OAI21_X1   g07275(.A1(new_n8178_), .A2(new_n8228_), .B(new_n8271_), .ZN(new_n8278_));
  AOI21_X1   g07276(.A1(new_n8278_), .A2(new_n8277_), .B(new_n8276_), .ZN(new_n8279_));
  OAI22_X1   g07277(.A1(new_n8275_), .A2(new_n8279_), .B1(new_n8258_), .B2(new_n8264_), .ZN(new_n8280_));
  OAI21_X1   g07278(.A1(new_n8260_), .A2(new_n8219_), .B(new_n8263_), .ZN(new_n8281_));
  NAND2_X1   g07279(.A1(new_n8248_), .A2(new_n8257_), .ZN(new_n8282_));
  NAND3_X1   g07280(.A1(new_n8278_), .A2(new_n8277_), .A3(new_n8276_), .ZN(new_n8283_));
  OAI21_X1   g07281(.A1(new_n8272_), .A2(new_n8274_), .B(new_n8267_), .ZN(new_n8284_));
  NAND4_X1   g07282(.A1(new_n8284_), .A2(new_n8283_), .A3(new_n8282_), .A4(new_n8281_), .ZN(new_n8285_));
  NAND3_X1   g07283(.A1(new_n8280_), .A2(new_n8247_), .A3(new_n8285_), .ZN(new_n8286_));
  AOI21_X1   g07284(.A1(new_n8232_), .A2(new_n8216_), .B(new_n8234_), .ZN(new_n8287_));
  AOI22_X1   g07285(.A1(new_n8284_), .A2(new_n8283_), .B1(new_n8282_), .B2(new_n8281_), .ZN(new_n8288_));
  NOR4_X1    g07286(.A1(new_n8275_), .A2(new_n8279_), .A3(new_n8258_), .A4(new_n8264_), .ZN(new_n8289_));
  OAI21_X1   g07287(.A1(new_n8288_), .A2(new_n8289_), .B(new_n8287_), .ZN(new_n8290_));
  OAI21_X1   g07288(.A1(new_n8110_), .A2(new_n8151_), .B(new_n8166_), .ZN(new_n8291_));
  XOR2_X1    g07289(.A1(new_n7044_), .A2(new_n8097_), .Z(new_n8292_));
  OAI21_X1   g07290(.A1(new_n8107_), .A2(new_n8090_), .B(new_n8292_), .ZN(new_n8293_));
  NOR2_X1    g07291(.A1(new_n8081_), .A2(new_n8082_), .ZN(new_n8294_));
  AOI21_X1   g07292(.A1(new_n7042_), .A2(new_n8091_), .B(new_n8294_), .ZN(new_n8295_));
  INV_X1     g07293(.I(new_n8095_), .ZN(new_n8296_));
  AOI21_X1   g07294(.A1(new_n7044_), .A2(new_n8096_), .B(new_n8296_), .ZN(new_n8297_));
  XOR2_X1    g07295(.A1(new_n8295_), .A2(new_n8297_), .Z(new_n8298_));
  AOI21_X1   g07296(.A1(new_n8293_), .A2(new_n8094_), .B(new_n8298_), .ZN(new_n8299_));
  NAND3_X1   g07297(.A1(new_n7040_), .A2(new_n7042_), .A3(new_n7043_), .ZN(new_n8300_));
  NOR2_X1    g07298(.A1(new_n7007_), .A2(new_n8091_), .ZN(new_n8301_));
  NOR4_X1    g07299(.A1(new_n8101_), .A2(new_n8300_), .A3(new_n8106_), .A4(new_n8301_), .ZN(new_n8302_));
  XNOR2_X1   g07300(.A1(new_n8295_), .A2(new_n8297_), .ZN(new_n8303_));
  NOR3_X1    g07301(.A1(new_n8103_), .A2(new_n8303_), .A3(new_n8302_), .ZN(new_n8304_));
  NOR2_X1    g07302(.A1(new_n8126_), .A2(new_n8116_), .ZN(new_n8305_));
  OAI21_X1   g07303(.A1(new_n8305_), .A2(new_n8140_), .B(new_n8143_), .ZN(new_n8306_));
  NOR2_X1    g07304(.A1(new_n8118_), .A2(new_n8120_), .ZN(new_n8307_));
  AOI21_X1   g07305(.A1(new_n7069_), .A2(new_n8121_), .B(new_n8307_), .ZN(new_n8308_));
  NOR2_X1    g07306(.A1(new_n8112_), .A2(new_n8113_), .ZN(new_n8309_));
  NAND2_X1   g07307(.A1(new_n8112_), .A2(new_n8113_), .ZN(new_n8310_));
  AOI21_X1   g07308(.A1(new_n7102_), .A2(new_n8310_), .B(new_n8309_), .ZN(new_n8311_));
  XOR2_X1    g07309(.A1(new_n8308_), .A2(new_n8311_), .Z(new_n8312_));
  AOI21_X1   g07310(.A1(new_n8306_), .A2(new_n8156_), .B(new_n8312_), .ZN(new_n8313_));
  NAND2_X1   g07311(.A1(new_n8139_), .A2(new_n8134_), .ZN(new_n8314_));
  AOI21_X1   g07312(.A1(new_n8314_), .A2(new_n8147_), .B(new_n8115_), .ZN(new_n8315_));
  XNOR2_X1   g07313(.A1(new_n8308_), .A2(new_n8311_), .ZN(new_n8316_));
  NOR3_X1    g07314(.A1(new_n8315_), .A2(new_n8149_), .A3(new_n8316_), .ZN(new_n8317_));
  OAI22_X1   g07315(.A1(new_n8317_), .A2(new_n8313_), .B1(new_n8304_), .B2(new_n8299_), .ZN(new_n8318_));
  OAI21_X1   g07316(.A1(new_n8103_), .A2(new_n8302_), .B(new_n8303_), .ZN(new_n8319_));
  NAND3_X1   g07317(.A1(new_n8293_), .A2(new_n8298_), .A3(new_n8094_), .ZN(new_n8320_));
  OAI21_X1   g07318(.A1(new_n8315_), .A2(new_n8149_), .B(new_n8316_), .ZN(new_n8321_));
  NAND3_X1   g07319(.A1(new_n8306_), .A2(new_n8156_), .A3(new_n8312_), .ZN(new_n8322_));
  NAND4_X1   g07320(.A1(new_n8321_), .A2(new_n8322_), .A3(new_n8319_), .A4(new_n8320_), .ZN(new_n8323_));
  NAND3_X1   g07321(.A1(new_n8291_), .A2(new_n8318_), .A3(new_n8323_), .ZN(new_n8324_));
  AOI21_X1   g07322(.A1(new_n8164_), .A2(new_n8165_), .B(new_n8158_), .ZN(new_n8325_));
  NAND2_X1   g07323(.A1(new_n8318_), .A2(new_n8323_), .ZN(new_n8326_));
  NAND2_X1   g07324(.A1(new_n8326_), .A2(new_n8325_), .ZN(new_n8327_));
  AOI22_X1   g07325(.A1(new_n8290_), .A2(new_n8286_), .B1(new_n8324_), .B2(new_n8327_), .ZN(new_n8328_));
  NOR3_X1    g07326(.A1(new_n8287_), .A2(new_n8289_), .A3(new_n8288_), .ZN(new_n8329_));
  AOI21_X1   g07327(.A1(new_n8280_), .A2(new_n8285_), .B(new_n8247_), .ZN(new_n8330_));
  NAND2_X1   g07328(.A1(new_n8327_), .A2(new_n8324_), .ZN(new_n8331_));
  NOR3_X1    g07329(.A1(new_n8329_), .A2(new_n8331_), .A3(new_n8330_), .ZN(new_n8332_));
  NOR3_X1    g07330(.A1(new_n8246_), .A2(new_n8328_), .A3(new_n8332_), .ZN(new_n8333_));
  NAND2_X1   g07331(.A1(new_n8236_), .A2(new_n7119_), .ZN(new_n8334_));
  NAND2_X1   g07332(.A1(new_n8334_), .A2(new_n8239_), .ZN(new_n8335_));
  OAI21_X1   g07333(.A1(new_n8329_), .A2(new_n8330_), .B(new_n8331_), .ZN(new_n8336_));
  NAND4_X1   g07334(.A1(new_n8290_), .A2(new_n8286_), .A3(new_n8324_), .A4(new_n8327_), .ZN(new_n8337_));
  AOI21_X1   g07335(.A1(new_n8336_), .A2(new_n8337_), .B(new_n8335_), .ZN(new_n8338_));
  NOR2_X1    g07336(.A1(new_n8338_), .A2(new_n8333_), .ZN(new_n8339_));
  AOI21_X1   g07337(.A1(new_n7853_), .A2(new_n8062_), .B(new_n8071_), .ZN(new_n8340_));
  INV_X1     g07338(.I(new_n8340_), .ZN(new_n8341_));
  OAI21_X1   g07339(.A1(new_n8056_), .A2(new_n8060_), .B(new_n7964_), .ZN(new_n8342_));
  NAND2_X1   g07340(.A1(new_n8040_), .A2(new_n8000_), .ZN(new_n8343_));
  INV_X1     g07341(.I(new_n7970_), .ZN(new_n8344_));
  OAI21_X1   g07342(.A1(new_n7965_), .A2(new_n7971_), .B(new_n8344_), .ZN(new_n8345_));
  XOR2_X1    g07343(.A1(new_n8345_), .A2(new_n7993_), .Z(new_n8346_));
  OAI21_X1   g07344(.A1(new_n8046_), .A2(new_n7984_), .B(new_n8346_), .ZN(new_n8347_));
  XOR2_X1    g07345(.A1(new_n7992_), .A2(new_n8345_), .Z(new_n8348_));
  NAND3_X1   g07346(.A1(new_n7996_), .A2(new_n8043_), .A3(new_n8348_), .ZN(new_n8349_));
  AOI21_X1   g07347(.A1(new_n8022_), .A2(new_n7430_), .B(new_n8026_), .ZN(new_n8350_));
  NOR2_X1    g07348(.A1(new_n8010_), .A2(new_n8012_), .ZN(new_n8351_));
  AOI21_X1   g07349(.A1(new_n8015_), .A2(new_n8029_), .B(new_n8351_), .ZN(new_n8352_));
  OAI21_X1   g07350(.A1(new_n8025_), .A2(new_n8005_), .B(new_n8004_), .ZN(new_n8353_));
  NOR2_X1    g07351(.A1(new_n8353_), .A2(new_n8352_), .ZN(new_n8354_));
  INV_X1     g07352(.I(new_n8029_), .ZN(new_n8355_));
  INV_X1     g07353(.I(new_n8351_), .ZN(new_n8356_));
  OAI21_X1   g07354(.A1(new_n8009_), .A2(new_n8355_), .B(new_n8356_), .ZN(new_n8357_));
  INV_X1     g07355(.I(new_n8004_), .ZN(new_n8358_));
  AOI21_X1   g07356(.A1(new_n8001_), .A2(new_n8006_), .B(new_n8358_), .ZN(new_n8359_));
  NOR2_X1    g07357(.A1(new_n8357_), .A2(new_n8359_), .ZN(new_n8360_));
  NOR2_X1    g07358(.A1(new_n8354_), .A2(new_n8360_), .ZN(new_n8361_));
  OAI21_X1   g07359(.A1(new_n8350_), .A2(new_n8038_), .B(new_n8361_), .ZN(new_n8362_));
  OAI21_X1   g07360(.A1(new_n8018_), .A2(new_n7446_), .B(new_n8008_), .ZN(new_n8363_));
  NAND2_X1   g07361(.A1(new_n8357_), .A2(new_n8359_), .ZN(new_n8364_));
  NAND2_X1   g07362(.A1(new_n8353_), .A2(new_n8352_), .ZN(new_n8365_));
  NAND2_X1   g07363(.A1(new_n8364_), .A2(new_n8365_), .ZN(new_n8366_));
  NAND3_X1   g07364(.A1(new_n8363_), .A2(new_n8032_), .A3(new_n8366_), .ZN(new_n8367_));
  NAND4_X1   g07365(.A1(new_n8347_), .A2(new_n8349_), .A3(new_n8362_), .A4(new_n8367_), .ZN(new_n8368_));
  AOI21_X1   g07366(.A1(new_n7996_), .A2(new_n8043_), .B(new_n8348_), .ZN(new_n8369_));
  NOR3_X1    g07367(.A1(new_n8046_), .A2(new_n7984_), .A3(new_n8346_), .ZN(new_n8370_));
  AOI21_X1   g07368(.A1(new_n8363_), .A2(new_n8032_), .B(new_n8366_), .ZN(new_n8371_));
  NOR3_X1    g07369(.A1(new_n8350_), .A2(new_n8038_), .A3(new_n8361_), .ZN(new_n8372_));
  OAI22_X1   g07370(.A1(new_n8370_), .A2(new_n8369_), .B1(new_n8372_), .B2(new_n8371_), .ZN(new_n8373_));
  AOI22_X1   g07371(.A1(new_n8343_), .A2(new_n8034_), .B1(new_n8373_), .B2(new_n8368_), .ZN(new_n8374_));
  NOR2_X1    g07372(.A1(new_n8052_), .A2(new_n8050_), .ZN(new_n8375_));
  NOR4_X1    g07373(.A1(new_n8370_), .A2(new_n8369_), .A3(new_n8372_), .A4(new_n8371_), .ZN(new_n8376_));
  AOI22_X1   g07374(.A1(new_n8347_), .A2(new_n8349_), .B1(new_n8362_), .B2(new_n8367_), .ZN(new_n8377_));
  NOR4_X1    g07375(.A1(new_n8375_), .A2(new_n8377_), .A3(new_n8376_), .A4(new_n8051_), .ZN(new_n8378_));
  AOI21_X1   g07376(.A1(new_n7899_), .A2(new_n7942_), .B(new_n7958_), .ZN(new_n8379_));
  NOR2_X1    g07377(.A1(new_n7896_), .A2(new_n7894_), .ZN(new_n8380_));
  NOR2_X1    g07378(.A1(new_n7867_), .A2(new_n7865_), .ZN(new_n8381_));
  AOI21_X1   g07379(.A1(new_n7890_), .A2(new_n7889_), .B(new_n8381_), .ZN(new_n8382_));
  INV_X1     g07380(.I(new_n7880_), .ZN(new_n8383_));
  OAI21_X1   g07381(.A1(new_n7856_), .A2(new_n7861_), .B(new_n8383_), .ZN(new_n8384_));
  XOR2_X1    g07382(.A1(new_n8384_), .A2(new_n8382_), .Z(new_n8385_));
  OAI21_X1   g07383(.A1(new_n8380_), .A2(new_n7952_), .B(new_n8385_), .ZN(new_n8386_));
  NAND2_X1   g07384(.A1(new_n7892_), .A2(new_n7882_), .ZN(new_n8387_));
  AOI21_X1   g07385(.A1(new_n7887_), .A2(new_n7888_), .B(new_n7880_), .ZN(new_n8388_));
  XOR2_X1    g07386(.A1(new_n8388_), .A2(new_n8382_), .Z(new_n8389_));
  NAND3_X1   g07387(.A1(new_n8387_), .A2(new_n8389_), .A3(new_n7879_), .ZN(new_n8390_));
  NAND2_X1   g07388(.A1(new_n7273_), .A2(new_n7917_), .ZN(new_n8391_));
  AOI21_X1   g07389(.A1(new_n8391_), .A2(new_n7929_), .B(new_n7932_), .ZN(new_n8392_));
  NOR2_X1    g07390(.A1(new_n7911_), .A2(new_n7913_), .ZN(new_n8393_));
  AOI21_X1   g07391(.A1(new_n7918_), .A2(new_n7914_), .B(new_n8393_), .ZN(new_n8394_));
  AOI21_X1   g07392(.A1(new_n7900_), .A2(new_n7927_), .B(new_n7905_), .ZN(new_n8395_));
  XNOR2_X1   g07393(.A1(new_n8394_), .A2(new_n8395_), .ZN(new_n8396_));
  OAI21_X1   g07394(.A1(new_n8392_), .A2(new_n7946_), .B(new_n8396_), .ZN(new_n8397_));
  NOR2_X1    g07395(.A1(new_n7926_), .A2(new_n7928_), .ZN(new_n8398_));
  OAI21_X1   g07396(.A1(new_n8398_), .A2(new_n7937_), .B(new_n7908_), .ZN(new_n8399_));
  XOR2_X1    g07397(.A1(new_n8394_), .A2(new_n8395_), .Z(new_n8400_));
  NAND3_X1   g07398(.A1(new_n8399_), .A2(new_n7940_), .A3(new_n8400_), .ZN(new_n8401_));
  AOI22_X1   g07399(.A1(new_n8386_), .A2(new_n8390_), .B1(new_n8397_), .B2(new_n8401_), .ZN(new_n8402_));
  AOI21_X1   g07400(.A1(new_n8387_), .A2(new_n7879_), .B(new_n8389_), .ZN(new_n8403_));
  NOR3_X1    g07401(.A1(new_n8380_), .A2(new_n7952_), .A3(new_n8385_), .ZN(new_n8404_));
  AOI21_X1   g07402(.A1(new_n8399_), .A2(new_n7940_), .B(new_n8400_), .ZN(new_n8405_));
  NOR3_X1    g07403(.A1(new_n8392_), .A2(new_n7946_), .A3(new_n8396_), .ZN(new_n8406_));
  NOR4_X1    g07404(.A1(new_n8403_), .A2(new_n8404_), .A3(new_n8405_), .A4(new_n8406_), .ZN(new_n8407_));
  NOR3_X1    g07405(.A1(new_n8379_), .A2(new_n8402_), .A3(new_n8407_), .ZN(new_n8408_));
  OAI21_X1   g07406(.A1(new_n7956_), .A2(new_n7957_), .B(new_n7948_), .ZN(new_n8409_));
  OAI22_X1   g07407(.A1(new_n8403_), .A2(new_n8404_), .B1(new_n8405_), .B2(new_n8406_), .ZN(new_n8410_));
  NAND4_X1   g07408(.A1(new_n8386_), .A2(new_n8390_), .A3(new_n8397_), .A4(new_n8401_), .ZN(new_n8411_));
  AOI21_X1   g07409(.A1(new_n8410_), .A2(new_n8411_), .B(new_n8409_), .ZN(new_n8412_));
  OAI22_X1   g07410(.A1(new_n8412_), .A2(new_n8408_), .B1(new_n8374_), .B2(new_n8378_), .ZN(new_n8413_));
  OAI22_X1   g07411(.A1(new_n8375_), .A2(new_n8051_), .B1(new_n8377_), .B2(new_n8376_), .ZN(new_n8414_));
  AOI21_X1   g07412(.A1(new_n8000_), .A2(new_n8040_), .B(new_n8051_), .ZN(new_n8415_));
  NAND3_X1   g07413(.A1(new_n8415_), .A2(new_n8368_), .A3(new_n8373_), .ZN(new_n8416_));
  NAND3_X1   g07414(.A1(new_n8409_), .A2(new_n8410_), .A3(new_n8411_), .ZN(new_n8417_));
  OAI21_X1   g07415(.A1(new_n8402_), .A2(new_n8407_), .B(new_n8379_), .ZN(new_n8418_));
  NAND4_X1   g07416(.A1(new_n8418_), .A2(new_n8414_), .A3(new_n8416_), .A4(new_n8417_), .ZN(new_n8419_));
  NAND3_X1   g07417(.A1(new_n8419_), .A2(new_n8413_), .A3(new_n8342_), .ZN(new_n8420_));
  AOI21_X1   g07418(.A1(new_n7960_), .A2(new_n8054_), .B(new_n8057_), .ZN(new_n8421_));
  AOI22_X1   g07419(.A1(new_n8418_), .A2(new_n8417_), .B1(new_n8416_), .B2(new_n8414_), .ZN(new_n8422_));
  NOR4_X1    g07420(.A1(new_n8412_), .A2(new_n8408_), .A3(new_n8374_), .A4(new_n8378_), .ZN(new_n8423_));
  OAI21_X1   g07421(.A1(new_n8422_), .A2(new_n8423_), .B(new_n8421_), .ZN(new_n8424_));
  NAND2_X1   g07422(.A1(new_n8424_), .A2(new_n8420_), .ZN(new_n8425_));
  NAND2_X1   g07423(.A1(new_n7736_), .A2(new_n7790_), .ZN(new_n8426_));
  NOR2_X1    g07424(.A1(new_n7708_), .A2(new_n7706_), .ZN(new_n8427_));
  AOI21_X1   g07425(.A1(new_n7734_), .A2(new_n7733_), .B(new_n8427_), .ZN(new_n8428_));
  INV_X1     g07426(.I(new_n7721_), .ZN(new_n8429_));
  AOI21_X1   g07427(.A1(new_n7732_), .A2(new_n7720_), .B(new_n8429_), .ZN(new_n8430_));
  XOR2_X1    g07428(.A1(new_n8430_), .A2(new_n8428_), .Z(new_n8431_));
  AOI21_X1   g07429(.A1(new_n8426_), .A2(new_n7719_), .B(new_n8431_), .ZN(new_n8432_));
  INV_X1     g07430(.I(new_n7719_), .ZN(new_n8433_));
  OAI21_X1   g07431(.A1(new_n7699_), .A2(new_n7702_), .B(new_n7721_), .ZN(new_n8434_));
  XOR2_X1    g07432(.A1(new_n8434_), .A2(new_n8428_), .Z(new_n8435_));
  NOR3_X1    g07433(.A1(new_n7727_), .A2(new_n8433_), .A3(new_n8435_), .ZN(new_n8436_));
  NOR2_X1    g07434(.A1(new_n7681_), .A2(new_n7755_), .ZN(new_n8437_));
  OAI21_X1   g07435(.A1(new_n8437_), .A2(new_n7771_), .B(new_n7774_), .ZN(new_n8438_));
  NOR2_X1    g07436(.A1(new_n7750_), .A2(new_n7752_), .ZN(new_n8439_));
  AOI21_X1   g07437(.A1(new_n7754_), .A2(new_n7753_), .B(new_n8439_), .ZN(new_n8440_));
  INV_X1     g07438(.I(new_n7744_), .ZN(new_n8441_));
  AOI21_X1   g07439(.A1(new_n7741_), .A2(new_n7746_), .B(new_n8441_), .ZN(new_n8442_));
  XOR2_X1    g07440(.A1(new_n8440_), .A2(new_n8442_), .Z(new_n8443_));
  AOI21_X1   g07441(.A1(new_n8438_), .A2(new_n7786_), .B(new_n8443_), .ZN(new_n8444_));
  NAND2_X1   g07442(.A1(new_n7765_), .A2(new_n7768_), .ZN(new_n8445_));
  AOI21_X1   g07443(.A1(new_n8445_), .A2(new_n7763_), .B(new_n7748_), .ZN(new_n8446_));
  XNOR2_X1   g07444(.A1(new_n8440_), .A2(new_n8442_), .ZN(new_n8447_));
  NOR3_X1    g07445(.A1(new_n8446_), .A2(new_n7779_), .A3(new_n8447_), .ZN(new_n8448_));
  NOR4_X1    g07446(.A1(new_n8432_), .A2(new_n8436_), .A3(new_n8444_), .A4(new_n8448_), .ZN(new_n8449_));
  OAI21_X1   g07447(.A1(new_n7727_), .A2(new_n8433_), .B(new_n8435_), .ZN(new_n8450_));
  NAND3_X1   g07448(.A1(new_n8426_), .A2(new_n8431_), .A3(new_n7719_), .ZN(new_n8451_));
  OAI21_X1   g07449(.A1(new_n8446_), .A2(new_n7779_), .B(new_n8447_), .ZN(new_n8452_));
  NAND3_X1   g07450(.A1(new_n8438_), .A2(new_n7786_), .A3(new_n8443_), .ZN(new_n8453_));
  AOI22_X1   g07451(.A1(new_n8450_), .A2(new_n8451_), .B1(new_n8452_), .B2(new_n8453_), .ZN(new_n8454_));
  AOI21_X1   g07452(.A1(new_n7794_), .A2(new_n7795_), .B(new_n7788_), .ZN(new_n8455_));
  NOR3_X1    g07453(.A1(new_n8455_), .A2(new_n8449_), .A3(new_n8454_), .ZN(new_n8456_));
  NAND4_X1   g07454(.A1(new_n8450_), .A2(new_n8451_), .A3(new_n8452_), .A4(new_n8453_), .ZN(new_n8457_));
  OAI22_X1   g07455(.A1(new_n8432_), .A2(new_n8436_), .B1(new_n8444_), .B2(new_n8448_), .ZN(new_n8458_));
  OAI21_X1   g07456(.A1(new_n7739_), .A2(new_n7781_), .B(new_n7796_), .ZN(new_n8459_));
  AOI21_X1   g07457(.A1(new_n8457_), .A2(new_n8458_), .B(new_n8459_), .ZN(new_n8460_));
  NOR2_X1    g07458(.A1(new_n8460_), .A2(new_n8456_), .ZN(new_n8461_));
  INV_X1     g07459(.I(new_n8461_), .ZN(new_n8462_));
  NOR2_X1    g07460(.A1(new_n7851_), .A2(new_n7798_), .ZN(new_n8463_));
  NAND2_X1   g07461(.A1(new_n7827_), .A2(new_n7811_), .ZN(new_n8464_));
  NAND3_X1   g07462(.A1(new_n7523_), .A2(new_n7819_), .A3(new_n7817_), .ZN(new_n8465_));
  NAND2_X1   g07463(.A1(new_n8465_), .A2(new_n7820_), .ZN(new_n8466_));
  AOI21_X1   g07464(.A1(new_n8464_), .A2(new_n7823_), .B(new_n8466_), .ZN(new_n8467_));
  INV_X1     g07465(.I(new_n8467_), .ZN(new_n8468_));
  NAND3_X1   g07466(.A1(new_n8464_), .A2(new_n7823_), .A3(new_n8466_), .ZN(new_n8469_));
  NAND2_X1   g07467(.A1(new_n8468_), .A2(new_n8469_), .ZN(new_n8470_));
  NAND2_X1   g07468(.A1(new_n7835_), .A2(new_n7837_), .ZN(new_n8471_));
  INV_X1     g07469(.I(new_n7800_), .ZN(new_n8472_));
  AOI21_X1   g07470(.A1(new_n8472_), .A2(new_n7807_), .B(new_n7805_), .ZN(new_n8473_));
  INV_X1     g07471(.I(new_n8473_), .ZN(new_n8474_));
  AOI21_X1   g07472(.A1(new_n8471_), .A2(new_n7832_), .B(new_n8474_), .ZN(new_n8475_));
  NOR2_X1    g07473(.A1(new_n7839_), .A2(new_n7809_), .ZN(new_n8476_));
  NOR3_X1    g07474(.A1(new_n8476_), .A2(new_n7838_), .A3(new_n8473_), .ZN(new_n8477_));
  NOR3_X1    g07475(.A1(new_n8477_), .A2(new_n8475_), .A3(new_n8470_), .ZN(new_n8478_));
  INV_X1     g07476(.I(new_n8469_), .ZN(new_n8479_));
  NOR2_X1    g07477(.A1(new_n8479_), .A2(new_n8467_), .ZN(new_n8480_));
  OAI21_X1   g07478(.A1(new_n8476_), .A2(new_n7838_), .B(new_n8473_), .ZN(new_n8481_));
  NAND3_X1   g07479(.A1(new_n8471_), .A2(new_n7832_), .A3(new_n8474_), .ZN(new_n8482_));
  AOI21_X1   g07480(.A1(new_n8481_), .A2(new_n8482_), .B(new_n8480_), .ZN(new_n8483_));
  NOR4_X1    g07481(.A1(new_n8463_), .A2(new_n8478_), .A3(new_n8483_), .A4(new_n7850_), .ZN(new_n8484_));
  NAND2_X1   g07482(.A1(new_n7845_), .A2(new_n7849_), .ZN(new_n8485_));
  NAND3_X1   g07483(.A1(new_n8481_), .A2(new_n8482_), .A3(new_n8480_), .ZN(new_n8486_));
  OAI21_X1   g07484(.A1(new_n8477_), .A2(new_n8475_), .B(new_n8470_), .ZN(new_n8487_));
  AOI22_X1   g07485(.A1(new_n8485_), .A2(new_n7841_), .B1(new_n8487_), .B2(new_n8486_), .ZN(new_n8488_));
  NOR3_X1    g07486(.A1(new_n8488_), .A2(new_n8484_), .A3(new_n8462_), .ZN(new_n8489_));
  NAND4_X1   g07487(.A1(new_n8485_), .A2(new_n8487_), .A3(new_n8486_), .A4(new_n7841_), .ZN(new_n8490_));
  OAI22_X1   g07488(.A1(new_n7850_), .A2(new_n8463_), .B1(new_n8478_), .B2(new_n8483_), .ZN(new_n8491_));
  AOI21_X1   g07489(.A1(new_n8491_), .A2(new_n8490_), .B(new_n8461_), .ZN(new_n8492_));
  NOR3_X1    g07490(.A1(new_n8425_), .A2(new_n8489_), .A3(new_n8492_), .ZN(new_n8493_));
  NAND3_X1   g07491(.A1(new_n8491_), .A2(new_n8490_), .A3(new_n8461_), .ZN(new_n8494_));
  OAI21_X1   g07492(.A1(new_n8488_), .A2(new_n8484_), .B(new_n8462_), .ZN(new_n8495_));
  AOI22_X1   g07493(.A1(new_n8495_), .A2(new_n8494_), .B1(new_n8420_), .B2(new_n8424_), .ZN(new_n8496_));
  NOR3_X1    g07494(.A1(new_n8496_), .A2(new_n8493_), .A3(new_n8341_), .ZN(new_n8497_));
  NAND4_X1   g07495(.A1(new_n8495_), .A2(new_n8494_), .A3(new_n8420_), .A4(new_n8424_), .ZN(new_n8498_));
  NOR3_X1    g07496(.A1(new_n8422_), .A2(new_n8423_), .A3(new_n8421_), .ZN(new_n8499_));
  AOI21_X1   g07497(.A1(new_n8419_), .A2(new_n8413_), .B(new_n8342_), .ZN(new_n8500_));
  OAI22_X1   g07498(.A1(new_n8489_), .A2(new_n8492_), .B1(new_n8499_), .B2(new_n8500_), .ZN(new_n8501_));
  AOI21_X1   g07499(.A1(new_n8501_), .A2(new_n8498_), .B(new_n8340_), .ZN(new_n8502_));
  OAI21_X1   g07500(.A1(new_n8497_), .A2(new_n8502_), .B(new_n8339_), .ZN(new_n8503_));
  NOR3_X1    g07501(.A1(new_n8497_), .A2(new_n8502_), .A3(new_n8339_), .ZN(new_n8504_));
  AOI21_X1   g07502(.A1(new_n8244_), .A2(new_n8503_), .B(new_n8504_), .ZN(new_n8505_));
  AOI21_X1   g07503(.A1(new_n8335_), .A2(new_n8336_), .B(new_n8332_), .ZN(new_n8506_));
  NAND2_X1   g07504(.A1(new_n8325_), .A2(new_n8323_), .ZN(new_n8507_));
  NAND2_X1   g07505(.A1(new_n8507_), .A2(new_n8318_), .ZN(new_n8508_));
  INV_X1     g07506(.I(new_n8311_), .ZN(new_n8509_));
  NAND3_X1   g07507(.A1(new_n8306_), .A2(new_n8156_), .A3(new_n8509_), .ZN(new_n8510_));
  AOI21_X1   g07508(.A1(new_n8306_), .A2(new_n8156_), .B(new_n8509_), .ZN(new_n8511_));
  OAI21_X1   g07509(.A1(new_n8308_), .A2(new_n8511_), .B(new_n8510_), .ZN(new_n8512_));
  INV_X1     g07510(.I(new_n8295_), .ZN(new_n8513_));
  NAND2_X1   g07511(.A1(new_n8293_), .A2(new_n8094_), .ZN(new_n8514_));
  NOR2_X1    g07512(.A1(new_n8514_), .A2(new_n8297_), .ZN(new_n8515_));
  NAND2_X1   g07513(.A1(new_n8514_), .A2(new_n8297_), .ZN(new_n8516_));
  AOI21_X1   g07514(.A1(new_n8513_), .A2(new_n8516_), .B(new_n8515_), .ZN(new_n8517_));
  XOR2_X1    g07515(.A1(new_n8517_), .A2(new_n8512_), .Z(new_n8518_));
  NAND2_X1   g07516(.A1(new_n8518_), .A2(new_n8508_), .ZN(new_n8519_));
  INV_X1     g07517(.I(new_n8318_), .ZN(new_n8520_));
  AOI21_X1   g07518(.A1(new_n8325_), .A2(new_n8323_), .B(new_n8520_), .ZN(new_n8521_));
  NOR2_X1    g07519(.A1(new_n8103_), .A2(new_n8302_), .ZN(new_n8522_));
  INV_X1     g07520(.I(new_n8297_), .ZN(new_n8523_));
  NAND2_X1   g07521(.A1(new_n8522_), .A2(new_n8523_), .ZN(new_n8524_));
  NOR2_X1    g07522(.A1(new_n8522_), .A2(new_n8523_), .ZN(new_n8525_));
  OAI21_X1   g07523(.A1(new_n8525_), .A2(new_n8295_), .B(new_n8524_), .ZN(new_n8526_));
  XOR2_X1    g07524(.A1(new_n8526_), .A2(new_n8512_), .Z(new_n8527_));
  NAND2_X1   g07525(.A1(new_n8527_), .A2(new_n8521_), .ZN(new_n8528_));
  OAI21_X1   g07526(.A1(new_n8288_), .A2(new_n8247_), .B(new_n8285_), .ZN(new_n8529_));
  OAI21_X1   g07527(.A1(new_n8276_), .A2(new_n8274_), .B(new_n8277_), .ZN(new_n8530_));
  OAI21_X1   g07528(.A1(new_n8248_), .A2(new_n8261_), .B(new_n8256_), .ZN(new_n8531_));
  INV_X1     g07529(.I(new_n8531_), .ZN(new_n8532_));
  NAND2_X1   g07530(.A1(new_n8532_), .A2(new_n8530_), .ZN(new_n8533_));
  INV_X1     g07531(.I(new_n8530_), .ZN(new_n8534_));
  NAND2_X1   g07532(.A1(new_n8534_), .A2(new_n8531_), .ZN(new_n8535_));
  NAND2_X1   g07533(.A1(new_n8533_), .A2(new_n8535_), .ZN(new_n8536_));
  NAND2_X1   g07534(.A1(new_n8536_), .A2(new_n8529_), .ZN(new_n8537_));
  AOI21_X1   g07535(.A1(new_n8287_), .A2(new_n8280_), .B(new_n8289_), .ZN(new_n8538_));
  NOR2_X1    g07536(.A1(new_n8534_), .A2(new_n8531_), .ZN(new_n8539_));
  NOR2_X1    g07537(.A1(new_n8532_), .A2(new_n8530_), .ZN(new_n8540_));
  NOR2_X1    g07538(.A1(new_n8540_), .A2(new_n8539_), .ZN(new_n8541_));
  NAND2_X1   g07539(.A1(new_n8538_), .A2(new_n8541_), .ZN(new_n8542_));
  AOI22_X1   g07540(.A1(new_n8542_), .A2(new_n8537_), .B1(new_n8528_), .B2(new_n8519_), .ZN(new_n8543_));
  NOR2_X1    g07541(.A1(new_n8527_), .A2(new_n8521_), .ZN(new_n8544_));
  NOR2_X1    g07542(.A1(new_n8518_), .A2(new_n8508_), .ZN(new_n8545_));
  NOR2_X1    g07543(.A1(new_n8538_), .A2(new_n8541_), .ZN(new_n8546_));
  NOR2_X1    g07544(.A1(new_n8536_), .A2(new_n8529_), .ZN(new_n8547_));
  NOR4_X1    g07545(.A1(new_n8546_), .A2(new_n8547_), .A3(new_n8544_), .A4(new_n8545_), .ZN(new_n8548_));
  NOR3_X1    g07546(.A1(new_n8506_), .A2(new_n8543_), .A3(new_n8548_), .ZN(new_n8549_));
  OAI21_X1   g07547(.A1(new_n8246_), .A2(new_n8328_), .B(new_n8337_), .ZN(new_n8550_));
  OAI22_X1   g07548(.A1(new_n8546_), .A2(new_n8547_), .B1(new_n8544_), .B2(new_n8545_), .ZN(new_n8551_));
  NAND4_X1   g07549(.A1(new_n8542_), .A2(new_n8537_), .A3(new_n8528_), .A4(new_n8519_), .ZN(new_n8552_));
  AOI21_X1   g07550(.A1(new_n8551_), .A2(new_n8552_), .B(new_n8550_), .ZN(new_n8553_));
  NOR2_X1    g07551(.A1(new_n8553_), .A2(new_n8549_), .ZN(new_n8554_));
  NOR2_X1    g07552(.A1(new_n8505_), .A2(new_n8554_), .ZN(new_n8555_));
  AOI21_X1   g07553(.A1(new_n8342_), .A2(new_n8413_), .B(new_n8423_), .ZN(new_n8556_));
  OAI21_X1   g07554(.A1(new_n8409_), .A2(new_n8407_), .B(new_n8410_), .ZN(new_n8557_));
  INV_X1     g07555(.I(new_n8394_), .ZN(new_n8558_));
  NOR3_X1    g07556(.A1(new_n8392_), .A2(new_n7946_), .A3(new_n8395_), .ZN(new_n8559_));
  OAI21_X1   g07557(.A1(new_n8392_), .A2(new_n7946_), .B(new_n8395_), .ZN(new_n8560_));
  AOI21_X1   g07558(.A1(new_n8558_), .A2(new_n8560_), .B(new_n8559_), .ZN(new_n8561_));
  NAND3_X1   g07559(.A1(new_n8387_), .A2(new_n7879_), .A3(new_n8384_), .ZN(new_n8562_));
  AOI21_X1   g07560(.A1(new_n8387_), .A2(new_n7879_), .B(new_n8384_), .ZN(new_n8563_));
  OAI21_X1   g07561(.A1(new_n8382_), .A2(new_n8563_), .B(new_n8562_), .ZN(new_n8564_));
  XOR2_X1    g07562(.A1(new_n8564_), .A2(new_n8561_), .Z(new_n8565_));
  NAND2_X1   g07563(.A1(new_n8565_), .A2(new_n8557_), .ZN(new_n8566_));
  AOI21_X1   g07564(.A1(new_n8379_), .A2(new_n8411_), .B(new_n8402_), .ZN(new_n8567_));
  XNOR2_X1   g07565(.A1(new_n8564_), .A2(new_n8561_), .ZN(new_n8568_));
  NAND2_X1   g07566(.A1(new_n8568_), .A2(new_n8567_), .ZN(new_n8569_));
  OAI21_X1   g07567(.A1(new_n8415_), .A2(new_n8376_), .B(new_n8373_), .ZN(new_n8570_));
  NOR3_X1    g07568(.A1(new_n8350_), .A2(new_n8038_), .A3(new_n8359_), .ZN(new_n8571_));
  OAI21_X1   g07569(.A1(new_n8350_), .A2(new_n8038_), .B(new_n8359_), .ZN(new_n8572_));
  AOI21_X1   g07570(.A1(new_n8357_), .A2(new_n8572_), .B(new_n8571_), .ZN(new_n8573_));
  NAND3_X1   g07571(.A1(new_n7996_), .A2(new_n8043_), .A3(new_n8345_), .ZN(new_n8574_));
  AOI21_X1   g07572(.A1(new_n7996_), .A2(new_n8043_), .B(new_n8345_), .ZN(new_n8575_));
  OAI21_X1   g07573(.A1(new_n7993_), .A2(new_n8575_), .B(new_n8574_), .ZN(new_n8576_));
  XOR2_X1    g07574(.A1(new_n8576_), .A2(new_n8573_), .Z(new_n8577_));
  NAND2_X1   g07575(.A1(new_n8577_), .A2(new_n8570_), .ZN(new_n8578_));
  OAI21_X1   g07576(.A1(new_n8050_), .A2(new_n8052_), .B(new_n8034_), .ZN(new_n8579_));
  AOI21_X1   g07577(.A1(new_n8579_), .A2(new_n8368_), .B(new_n8377_), .ZN(new_n8580_));
  XNOR2_X1   g07578(.A1(new_n8576_), .A2(new_n8573_), .ZN(new_n8581_));
  NAND2_X1   g07579(.A1(new_n8581_), .A2(new_n8580_), .ZN(new_n8582_));
  AOI22_X1   g07580(.A1(new_n8569_), .A2(new_n8566_), .B1(new_n8578_), .B2(new_n8582_), .ZN(new_n8583_));
  NOR2_X1    g07581(.A1(new_n8568_), .A2(new_n8567_), .ZN(new_n8584_));
  NOR2_X1    g07582(.A1(new_n8565_), .A2(new_n8557_), .ZN(new_n8585_));
  NOR2_X1    g07583(.A1(new_n8581_), .A2(new_n8580_), .ZN(new_n8586_));
  NOR2_X1    g07584(.A1(new_n8577_), .A2(new_n8570_), .ZN(new_n8587_));
  NOR4_X1    g07585(.A1(new_n8584_), .A2(new_n8585_), .A3(new_n8586_), .A4(new_n8587_), .ZN(new_n8588_));
  NOR3_X1    g07586(.A1(new_n8583_), .A2(new_n8588_), .A3(new_n8556_), .ZN(new_n8589_));
  OAI21_X1   g07587(.A1(new_n8422_), .A2(new_n8421_), .B(new_n8419_), .ZN(new_n8590_));
  OAI22_X1   g07588(.A1(new_n8584_), .A2(new_n8585_), .B1(new_n8586_), .B2(new_n8587_), .ZN(new_n8591_));
  NAND4_X1   g07589(.A1(new_n8569_), .A2(new_n8566_), .A3(new_n8582_), .A4(new_n8578_), .ZN(new_n8592_));
  AOI21_X1   g07590(.A1(new_n8591_), .A2(new_n8592_), .B(new_n8590_), .ZN(new_n8593_));
  AOI21_X1   g07591(.A1(new_n8461_), .A2(new_n8490_), .B(new_n8488_), .ZN(new_n8594_));
  AOI21_X1   g07592(.A1(new_n7837_), .A2(new_n7835_), .B(new_n7838_), .ZN(new_n8595_));
  NAND2_X1   g07593(.A1(new_n8595_), .A2(new_n8470_), .ZN(new_n8596_));
  AOI21_X1   g07594(.A1(new_n8596_), .A2(new_n8473_), .B(new_n8468_), .ZN(new_n8597_));
  OAI21_X1   g07595(.A1(new_n7809_), .A2(new_n7839_), .B(new_n7832_), .ZN(new_n8598_));
  AOI21_X1   g07596(.A1(new_n8598_), .A2(new_n8473_), .B(new_n8480_), .ZN(new_n8599_));
  NOR3_X1    g07597(.A1(new_n8599_), .A2(new_n8467_), .A3(new_n8477_), .ZN(new_n8600_));
  AOI21_X1   g07598(.A1(new_n8455_), .A2(new_n8457_), .B(new_n8454_), .ZN(new_n8601_));
  INV_X1     g07599(.I(new_n8442_), .ZN(new_n8602_));
  NAND3_X1   g07600(.A1(new_n8438_), .A2(new_n7786_), .A3(new_n8602_), .ZN(new_n8603_));
  AOI21_X1   g07601(.A1(new_n8438_), .A2(new_n7786_), .B(new_n8602_), .ZN(new_n8604_));
  OAI21_X1   g07602(.A1(new_n8440_), .A2(new_n8604_), .B(new_n8603_), .ZN(new_n8605_));
  INV_X1     g07603(.I(new_n8428_), .ZN(new_n8606_));
  NOR3_X1    g07604(.A1(new_n7727_), .A2(new_n8433_), .A3(new_n8430_), .ZN(new_n8607_));
  OAI21_X1   g07605(.A1(new_n7727_), .A2(new_n8433_), .B(new_n8430_), .ZN(new_n8608_));
  AOI21_X1   g07606(.A1(new_n8606_), .A2(new_n8608_), .B(new_n8607_), .ZN(new_n8609_));
  NOR2_X1    g07607(.A1(new_n8609_), .A2(new_n8605_), .ZN(new_n8610_));
  INV_X1     g07608(.I(new_n8440_), .ZN(new_n8611_));
  NOR3_X1    g07609(.A1(new_n8446_), .A2(new_n7779_), .A3(new_n8442_), .ZN(new_n8612_));
  OAI21_X1   g07610(.A1(new_n8446_), .A2(new_n7779_), .B(new_n8442_), .ZN(new_n8613_));
  AOI21_X1   g07611(.A1(new_n8611_), .A2(new_n8613_), .B(new_n8612_), .ZN(new_n8614_));
  NAND3_X1   g07612(.A1(new_n8426_), .A2(new_n7719_), .A3(new_n8434_), .ZN(new_n8615_));
  AOI21_X1   g07613(.A1(new_n8426_), .A2(new_n7719_), .B(new_n8434_), .ZN(new_n8616_));
  OAI21_X1   g07614(.A1(new_n8428_), .A2(new_n8616_), .B(new_n8615_), .ZN(new_n8617_));
  NOR2_X1    g07615(.A1(new_n8617_), .A2(new_n8614_), .ZN(new_n8618_));
  NOR3_X1    g07616(.A1(new_n8601_), .A2(new_n8610_), .A3(new_n8618_), .ZN(new_n8619_));
  OAI21_X1   g07617(.A1(new_n8459_), .A2(new_n8449_), .B(new_n8458_), .ZN(new_n8620_));
  NAND2_X1   g07618(.A1(new_n8617_), .A2(new_n8614_), .ZN(new_n8621_));
  NAND2_X1   g07619(.A1(new_n8609_), .A2(new_n8605_), .ZN(new_n8622_));
  AOI21_X1   g07620(.A1(new_n8621_), .A2(new_n8622_), .B(new_n8620_), .ZN(new_n8623_));
  OAI22_X1   g07621(.A1(new_n8623_), .A2(new_n8619_), .B1(new_n8600_), .B2(new_n8597_), .ZN(new_n8624_));
  NOR2_X1    g07622(.A1(new_n8598_), .A2(new_n8480_), .ZN(new_n8625_));
  OAI21_X1   g07623(.A1(new_n8625_), .A2(new_n8474_), .B(new_n8467_), .ZN(new_n8626_));
  OAI21_X1   g07624(.A1(new_n8595_), .A2(new_n8474_), .B(new_n8470_), .ZN(new_n8627_));
  NAND3_X1   g07625(.A1(new_n8627_), .A2(new_n8468_), .A3(new_n8482_), .ZN(new_n8628_));
  NAND3_X1   g07626(.A1(new_n8620_), .A2(new_n8621_), .A3(new_n8622_), .ZN(new_n8629_));
  NAND2_X1   g07627(.A1(new_n8621_), .A2(new_n8622_), .ZN(new_n8630_));
  NAND2_X1   g07628(.A1(new_n8630_), .A2(new_n8601_), .ZN(new_n8631_));
  NAND4_X1   g07629(.A1(new_n8631_), .A2(new_n8628_), .A3(new_n8629_), .A4(new_n8626_), .ZN(new_n8632_));
  NAND2_X1   g07630(.A1(new_n8624_), .A2(new_n8632_), .ZN(new_n8633_));
  NOR2_X1    g07631(.A1(new_n8594_), .A2(new_n8633_), .ZN(new_n8634_));
  OAI21_X1   g07632(.A1(new_n8462_), .A2(new_n8484_), .B(new_n8491_), .ZN(new_n8635_));
  AOI22_X1   g07633(.A1(new_n8631_), .A2(new_n8629_), .B1(new_n8628_), .B2(new_n8626_), .ZN(new_n8636_));
  NOR4_X1    g07634(.A1(new_n8623_), .A2(new_n8619_), .A3(new_n8600_), .A4(new_n8597_), .ZN(new_n8637_));
  NOR2_X1    g07635(.A1(new_n8637_), .A2(new_n8636_), .ZN(new_n8638_));
  NOR2_X1    g07636(.A1(new_n8638_), .A2(new_n8635_), .ZN(new_n8639_));
  NOR4_X1    g07637(.A1(new_n8639_), .A2(new_n8634_), .A3(new_n8589_), .A4(new_n8593_), .ZN(new_n8640_));
  NAND3_X1   g07638(.A1(new_n8591_), .A2(new_n8592_), .A3(new_n8590_), .ZN(new_n8641_));
  OAI21_X1   g07639(.A1(new_n8583_), .A2(new_n8588_), .B(new_n8556_), .ZN(new_n8642_));
  NAND2_X1   g07640(.A1(new_n8638_), .A2(new_n8635_), .ZN(new_n8643_));
  NAND2_X1   g07641(.A1(new_n8594_), .A2(new_n8633_), .ZN(new_n8644_));
  AOI22_X1   g07642(.A1(new_n8643_), .A2(new_n8644_), .B1(new_n8641_), .B2(new_n8642_), .ZN(new_n8645_));
  NOR2_X1    g07643(.A1(new_n8645_), .A2(new_n8640_), .ZN(new_n8646_));
  AOI21_X1   g07644(.A1(new_n8341_), .A2(new_n8501_), .B(new_n8493_), .ZN(new_n8647_));
  NOR2_X1    g07645(.A1(new_n8646_), .A2(new_n8647_), .ZN(new_n8648_));
  NAND4_X1   g07646(.A1(new_n8643_), .A2(new_n8644_), .A3(new_n8641_), .A4(new_n8642_), .ZN(new_n8649_));
  OAI22_X1   g07647(.A1(new_n8639_), .A2(new_n8634_), .B1(new_n8589_), .B2(new_n8593_), .ZN(new_n8650_));
  NAND2_X1   g07648(.A1(new_n8650_), .A2(new_n8649_), .ZN(new_n8651_));
  OAI21_X1   g07649(.A1(new_n8496_), .A2(new_n8340_), .B(new_n8498_), .ZN(new_n8652_));
  NOR2_X1    g07650(.A1(new_n8651_), .A2(new_n8652_), .ZN(new_n8653_));
  NOR2_X1    g07651(.A1(new_n8648_), .A2(new_n8653_), .ZN(new_n8654_));
  INV_X1     g07652(.I(new_n8339_), .ZN(new_n8655_));
  NAND3_X1   g07653(.A1(new_n8501_), .A2(new_n8498_), .A3(new_n8340_), .ZN(new_n8656_));
  OAI21_X1   g07654(.A1(new_n8496_), .A2(new_n8493_), .B(new_n8341_), .ZN(new_n8657_));
  NAND3_X1   g07655(.A1(new_n8657_), .A2(new_n8656_), .A3(new_n8655_), .ZN(new_n8658_));
  NAND2_X1   g07656(.A1(new_n8503_), .A2(new_n8244_), .ZN(new_n8659_));
  NAND3_X1   g07657(.A1(new_n8659_), .A2(new_n8658_), .A3(new_n8554_), .ZN(new_n8660_));
  OAI21_X1   g07658(.A1(new_n8555_), .A2(new_n8654_), .B(new_n8660_), .ZN(new_n8661_));
  NAND3_X1   g07659(.A1(new_n8529_), .A2(new_n8533_), .A3(new_n8535_), .ZN(new_n8662_));
  NOR2_X1    g07660(.A1(new_n8526_), .A2(new_n8512_), .ZN(new_n8663_));
  INV_X1     g07661(.I(new_n8663_), .ZN(new_n8664_));
  AOI21_X1   g07662(.A1(new_n8512_), .A2(new_n8526_), .B(new_n8521_), .ZN(new_n8665_));
  NAND2_X1   g07663(.A1(new_n8665_), .A2(new_n8664_), .ZN(new_n8666_));
  NAND2_X1   g07664(.A1(new_n8518_), .A2(new_n8521_), .ZN(new_n8667_));
  NAND2_X1   g07665(.A1(new_n8538_), .A2(new_n8536_), .ZN(new_n8668_));
  NAND4_X1   g07666(.A1(new_n8666_), .A2(new_n8662_), .A3(new_n8667_), .A4(new_n8668_), .ZN(new_n8669_));
  OAI21_X1   g07667(.A1(new_n8550_), .A2(new_n8548_), .B(new_n8669_), .ZN(new_n8670_));
  NOR2_X1    g07668(.A1(new_n8665_), .A2(new_n8663_), .ZN(new_n8671_));
  OAI21_X1   g07669(.A1(new_n8538_), .A2(new_n8539_), .B(new_n8535_), .ZN(new_n8672_));
  XOR2_X1    g07670(.A1(new_n8671_), .A2(new_n8672_), .Z(new_n8673_));
  AND2_X2    g07671(.A1(new_n8670_), .A2(new_n8673_), .Z(new_n8674_));
  NOR2_X1    g07672(.A1(new_n8670_), .A2(new_n8673_), .ZN(new_n8675_));
  OR2_X2     g07673(.A1(new_n8674_), .A2(new_n8675_), .Z(new_n8676_));
  AOI21_X1   g07674(.A1(new_n8650_), .A2(new_n8652_), .B(new_n8640_), .ZN(new_n8677_));
  NOR2_X1    g07675(.A1(new_n8484_), .A2(new_n8462_), .ZN(new_n8678_));
  OAI21_X1   g07676(.A1(new_n8678_), .A2(new_n8488_), .B(new_n8624_), .ZN(new_n8679_));
  NAND3_X1   g07677(.A1(new_n8627_), .A2(new_n8467_), .A3(new_n8482_), .ZN(new_n8680_));
  NOR2_X1    g07678(.A1(new_n8617_), .A2(new_n8605_), .ZN(new_n8681_));
  INV_X1     g07679(.I(new_n8681_), .ZN(new_n8682_));
  OAI21_X1   g07680(.A1(new_n8614_), .A2(new_n8609_), .B(new_n8620_), .ZN(new_n8683_));
  AOI21_X1   g07681(.A1(new_n8683_), .A2(new_n8682_), .B(new_n8680_), .ZN(new_n8684_));
  NAND3_X1   g07682(.A1(new_n8683_), .A2(new_n8680_), .A3(new_n8682_), .ZN(new_n8685_));
  INV_X1     g07683(.I(new_n8685_), .ZN(new_n8686_));
  NOR2_X1    g07684(.A1(new_n8686_), .A2(new_n8684_), .ZN(new_n8687_));
  NAND3_X1   g07685(.A1(new_n8679_), .A2(new_n8687_), .A3(new_n8632_), .ZN(new_n8688_));
  NAND2_X1   g07686(.A1(new_n8490_), .A2(new_n8461_), .ZN(new_n8689_));
  AOI21_X1   g07687(.A1(new_n8689_), .A2(new_n8491_), .B(new_n8636_), .ZN(new_n8690_));
  NOR3_X1    g07688(.A1(new_n8599_), .A2(new_n8468_), .A3(new_n8477_), .ZN(new_n8691_));
  AOI21_X1   g07689(.A1(new_n8605_), .A2(new_n8617_), .B(new_n8601_), .ZN(new_n8692_));
  OAI21_X1   g07690(.A1(new_n8692_), .A2(new_n8681_), .B(new_n8691_), .ZN(new_n8693_));
  NAND2_X1   g07691(.A1(new_n8693_), .A2(new_n8685_), .ZN(new_n8694_));
  OAI21_X1   g07692(.A1(new_n8690_), .A2(new_n8637_), .B(new_n8694_), .ZN(new_n8695_));
  NAND2_X1   g07693(.A1(new_n8688_), .A2(new_n8695_), .ZN(new_n8696_));
  NAND2_X1   g07694(.A1(new_n8592_), .A2(new_n8556_), .ZN(new_n8697_));
  INV_X1     g07695(.I(new_n8574_), .ZN(new_n8698_));
  NOR2_X1    g07696(.A1(new_n8575_), .A2(new_n7993_), .ZN(new_n8699_));
  NOR2_X1    g07697(.A1(new_n8699_), .A2(new_n8698_), .ZN(new_n8700_));
  NAND2_X1   g07698(.A1(new_n8700_), .A2(new_n8573_), .ZN(new_n8701_));
  INV_X1     g07699(.I(new_n8701_), .ZN(new_n8702_));
  NOR2_X1    g07700(.A1(new_n8700_), .A2(new_n8573_), .ZN(new_n8703_));
  NOR3_X1    g07701(.A1(new_n8702_), .A2(new_n8580_), .A3(new_n8703_), .ZN(new_n8704_));
  INV_X1     g07702(.I(new_n8559_), .ZN(new_n8705_));
  NAND2_X1   g07703(.A1(new_n8560_), .A2(new_n8558_), .ZN(new_n8706_));
  NAND2_X1   g07704(.A1(new_n8706_), .A2(new_n8705_), .ZN(new_n8707_));
  NOR2_X1    g07705(.A1(new_n8707_), .A2(new_n8564_), .ZN(new_n8708_));
  AND2_X2    g07706(.A1(new_n8707_), .A2(new_n8564_), .Z(new_n8709_));
  NOR3_X1    g07707(.A1(new_n8709_), .A2(new_n8567_), .A3(new_n8708_), .ZN(new_n8710_));
  NOR2_X1    g07708(.A1(new_n8568_), .A2(new_n8557_), .ZN(new_n8711_));
  NOR2_X1    g07709(.A1(new_n8581_), .A2(new_n8570_), .ZN(new_n8712_));
  NOR4_X1    g07710(.A1(new_n8711_), .A2(new_n8710_), .A3(new_n8712_), .A4(new_n8704_), .ZN(new_n8713_));
  INV_X1     g07711(.I(new_n8713_), .ZN(new_n8714_));
  NAND2_X1   g07712(.A1(new_n8707_), .A2(new_n8564_), .ZN(new_n8715_));
  AOI21_X1   g07713(.A1(new_n8557_), .A2(new_n8715_), .B(new_n8708_), .ZN(new_n8716_));
  OAI21_X1   g07714(.A1(new_n8580_), .A2(new_n8703_), .B(new_n8701_), .ZN(new_n8717_));
  XNOR2_X1   g07715(.A1(new_n8717_), .A2(new_n8716_), .ZN(new_n8718_));
  AOI21_X1   g07716(.A1(new_n8697_), .A2(new_n8714_), .B(new_n8718_), .ZN(new_n8719_));
  NOR2_X1    g07717(.A1(new_n8588_), .A2(new_n8590_), .ZN(new_n8720_));
  XOR2_X1    g07718(.A1(new_n8717_), .A2(new_n8716_), .Z(new_n8721_));
  NOR3_X1    g07719(.A1(new_n8720_), .A2(new_n8713_), .A3(new_n8721_), .ZN(new_n8722_));
  NOR2_X1    g07720(.A1(new_n8722_), .A2(new_n8719_), .ZN(new_n8723_));
  NAND2_X1   g07721(.A1(new_n8696_), .A2(new_n8723_), .ZN(new_n8724_));
  NOR3_X1    g07722(.A1(new_n8690_), .A2(new_n8637_), .A3(new_n8694_), .ZN(new_n8725_));
  AOI21_X1   g07723(.A1(new_n8679_), .A2(new_n8632_), .B(new_n8687_), .ZN(new_n8726_));
  NOR2_X1    g07724(.A1(new_n8726_), .A2(new_n8725_), .ZN(new_n8727_));
  OAI21_X1   g07725(.A1(new_n8720_), .A2(new_n8713_), .B(new_n8721_), .ZN(new_n8728_));
  AOI21_X1   g07726(.A1(new_n8556_), .A2(new_n8592_), .B(new_n8713_), .ZN(new_n8729_));
  NAND2_X1   g07727(.A1(new_n8729_), .A2(new_n8718_), .ZN(new_n8730_));
  NAND2_X1   g07728(.A1(new_n8730_), .A2(new_n8728_), .ZN(new_n8731_));
  NAND2_X1   g07729(.A1(new_n8727_), .A2(new_n8731_), .ZN(new_n8732_));
  NAND3_X1   g07730(.A1(new_n8677_), .A2(new_n8732_), .A3(new_n8724_), .ZN(new_n8733_));
  OAI21_X1   g07731(.A1(new_n8647_), .A2(new_n8645_), .B(new_n8649_), .ZN(new_n8734_));
  NOR2_X1    g07732(.A1(new_n8727_), .A2(new_n8731_), .ZN(new_n8735_));
  NOR2_X1    g07733(.A1(new_n8696_), .A2(new_n8723_), .ZN(new_n8736_));
  OAI21_X1   g07734(.A1(new_n8735_), .A2(new_n8736_), .B(new_n8734_), .ZN(new_n8737_));
  AOI21_X1   g07735(.A1(new_n8737_), .A2(new_n8733_), .B(new_n8676_), .ZN(new_n8738_));
  NOR2_X1    g07736(.A1(new_n8674_), .A2(new_n8675_), .ZN(new_n8739_));
  NOR3_X1    g07737(.A1(new_n8734_), .A2(new_n8735_), .A3(new_n8736_), .ZN(new_n8740_));
  AOI21_X1   g07738(.A1(new_n8724_), .A2(new_n8732_), .B(new_n8677_), .ZN(new_n8741_));
  NOR3_X1    g07739(.A1(new_n8741_), .A2(new_n8740_), .A3(new_n8739_), .ZN(new_n8742_));
  NOR2_X1    g07740(.A1(new_n8742_), .A2(new_n8738_), .ZN(new_n8743_));
  NOR2_X1    g07741(.A1(new_n8743_), .A2(new_n8661_), .ZN(new_n8744_));
  INV_X1     g07742(.I(new_n8244_), .ZN(new_n8745_));
  AOI21_X1   g07743(.A1(new_n8657_), .A2(new_n8656_), .B(new_n8655_), .ZN(new_n8746_));
  OAI21_X1   g07744(.A1(new_n8745_), .A2(new_n8746_), .B(new_n8658_), .ZN(new_n8747_));
  NAND3_X1   g07745(.A1(new_n8550_), .A2(new_n8551_), .A3(new_n8552_), .ZN(new_n8748_));
  OAI21_X1   g07746(.A1(new_n8543_), .A2(new_n8548_), .B(new_n8506_), .ZN(new_n8749_));
  NAND2_X1   g07747(.A1(new_n8749_), .A2(new_n8748_), .ZN(new_n8750_));
  NAND2_X1   g07748(.A1(new_n8651_), .A2(new_n8652_), .ZN(new_n8751_));
  NAND2_X1   g07749(.A1(new_n8646_), .A2(new_n8647_), .ZN(new_n8752_));
  AOI22_X1   g07750(.A1(new_n8747_), .A2(new_n8750_), .B1(new_n8751_), .B2(new_n8752_), .ZN(new_n8753_));
  NOR2_X1    g07751(.A1(new_n8747_), .A2(new_n8750_), .ZN(new_n8754_));
  NOR2_X1    g07752(.A1(new_n8753_), .A2(new_n8754_), .ZN(new_n8755_));
  OAI21_X1   g07753(.A1(new_n8741_), .A2(new_n8740_), .B(new_n8739_), .ZN(new_n8756_));
  NAND3_X1   g07754(.A1(new_n8737_), .A2(new_n8733_), .A3(new_n8676_), .ZN(new_n8757_));
  NAND2_X1   g07755(.A1(new_n8756_), .A2(new_n8757_), .ZN(new_n8758_));
  NOR2_X1    g07756(.A1(new_n8758_), .A2(new_n8755_), .ZN(new_n8759_));
  NOR2_X1    g07757(.A1(new_n8744_), .A2(new_n8759_), .ZN(new_n8760_));
  INV_X1     g07758(.I(\A[847] ), .ZN(new_n8761_));
  INV_X1     g07759(.I(\A[848] ), .ZN(new_n8762_));
  NAND2_X1   g07760(.A1(new_n8762_), .A2(\A[849] ), .ZN(new_n8763_));
  INV_X1     g07761(.I(\A[849] ), .ZN(new_n8764_));
  NAND2_X1   g07762(.A1(new_n8764_), .A2(\A[848] ), .ZN(new_n8765_));
  AOI21_X1   g07763(.A1(new_n8763_), .A2(new_n8765_), .B(new_n8761_), .ZN(new_n8766_));
  NAND2_X1   g07764(.A1(\A[848] ), .A2(\A[849] ), .ZN(new_n8767_));
  NOR2_X1    g07765(.A1(\A[848] ), .A2(\A[849] ), .ZN(new_n8768_));
  INV_X1     g07766(.I(new_n8768_), .ZN(new_n8769_));
  AOI21_X1   g07767(.A1(new_n8769_), .A2(new_n8767_), .B(\A[847] ), .ZN(new_n8770_));
  INV_X1     g07768(.I(\A[850] ), .ZN(new_n8771_));
  INV_X1     g07769(.I(\A[851] ), .ZN(new_n8772_));
  NAND2_X1   g07770(.A1(new_n8772_), .A2(\A[852] ), .ZN(new_n8773_));
  INV_X1     g07771(.I(\A[852] ), .ZN(new_n8774_));
  NAND2_X1   g07772(.A1(new_n8774_), .A2(\A[851] ), .ZN(new_n8775_));
  AOI21_X1   g07773(.A1(new_n8773_), .A2(new_n8775_), .B(new_n8771_), .ZN(new_n8776_));
  NAND2_X1   g07774(.A1(\A[851] ), .A2(\A[852] ), .ZN(new_n8777_));
  NOR2_X1    g07775(.A1(\A[851] ), .A2(\A[852] ), .ZN(new_n8778_));
  INV_X1     g07776(.I(new_n8778_), .ZN(new_n8779_));
  AOI21_X1   g07777(.A1(new_n8779_), .A2(new_n8777_), .B(\A[850] ), .ZN(new_n8780_));
  OR4_X2     g07778(.A1(new_n8766_), .A2(new_n8770_), .A3(new_n8780_), .A4(new_n8776_), .Z(new_n8781_));
  AOI21_X1   g07779(.A1(\A[851] ), .A2(\A[852] ), .B(\A[850] ), .ZN(new_n8782_));
  AOI21_X1   g07780(.A1(\A[848] ), .A2(\A[849] ), .B(\A[847] ), .ZN(new_n8783_));
  OAI22_X1   g07781(.A1(new_n8768_), .A2(new_n8783_), .B1(new_n8782_), .B2(new_n8778_), .ZN(new_n8784_));
  INV_X1     g07782(.I(new_n8784_), .ZN(new_n8785_));
  NOR4_X1    g07783(.A1(new_n8782_), .A2(new_n8783_), .A3(new_n8768_), .A4(new_n8778_), .ZN(new_n8786_));
  NOR2_X1    g07784(.A1(new_n8785_), .A2(new_n8786_), .ZN(new_n8787_));
  NAND2_X1   g07785(.A1(new_n8781_), .A2(new_n8787_), .ZN(new_n8788_));
  NOR4_X1    g07786(.A1(new_n8766_), .A2(new_n8770_), .A3(new_n8780_), .A4(new_n8776_), .ZN(new_n8789_));
  INV_X1     g07787(.I(new_n8786_), .ZN(new_n8790_));
  NAND2_X1   g07788(.A1(new_n8790_), .A2(new_n8784_), .ZN(new_n8791_));
  NAND2_X1   g07789(.A1(new_n8789_), .A2(new_n8791_), .ZN(new_n8792_));
  NAND2_X1   g07790(.A1(new_n8788_), .A2(new_n8792_), .ZN(new_n8793_));
  INV_X1     g07791(.I(\A[854] ), .ZN(new_n8794_));
  NAND2_X1   g07792(.A1(new_n8794_), .A2(\A[855] ), .ZN(new_n8795_));
  INV_X1     g07793(.I(new_n8795_), .ZN(new_n8796_));
  NOR2_X1    g07794(.A1(new_n8794_), .A2(\A[855] ), .ZN(new_n8797_));
  OAI21_X1   g07795(.A1(new_n8796_), .A2(new_n8797_), .B(\A[853] ), .ZN(new_n8798_));
  INV_X1     g07796(.I(\A[853] ), .ZN(new_n8799_));
  NOR2_X1    g07797(.A1(\A[854] ), .A2(\A[855] ), .ZN(new_n8800_));
  NAND2_X1   g07798(.A1(\A[854] ), .A2(\A[855] ), .ZN(new_n8801_));
  INV_X1     g07799(.I(new_n8801_), .ZN(new_n8802_));
  OAI21_X1   g07800(.A1(new_n8802_), .A2(new_n8800_), .B(new_n8799_), .ZN(new_n8803_));
  INV_X1     g07801(.I(\A[858] ), .ZN(new_n8804_));
  NOR2_X1    g07802(.A1(new_n8804_), .A2(\A[857] ), .ZN(new_n8805_));
  INV_X1     g07803(.I(\A[857] ), .ZN(new_n8806_));
  NOR2_X1    g07804(.A1(new_n8806_), .A2(\A[858] ), .ZN(new_n8807_));
  OAI21_X1   g07805(.A1(new_n8805_), .A2(new_n8807_), .B(\A[856] ), .ZN(new_n8808_));
  INV_X1     g07806(.I(\A[856] ), .ZN(new_n8809_));
  NOR2_X1    g07807(.A1(\A[857] ), .A2(\A[858] ), .ZN(new_n8810_));
  NAND2_X1   g07808(.A1(\A[857] ), .A2(\A[858] ), .ZN(new_n8811_));
  INV_X1     g07809(.I(new_n8811_), .ZN(new_n8812_));
  OAI21_X1   g07810(.A1(new_n8812_), .A2(new_n8810_), .B(new_n8809_), .ZN(new_n8813_));
  NAND4_X1   g07811(.A1(new_n8798_), .A2(new_n8803_), .A3(new_n8813_), .A4(new_n8808_), .ZN(new_n8814_));
  AOI21_X1   g07812(.A1(\A[857] ), .A2(\A[858] ), .B(\A[856] ), .ZN(new_n8815_));
  AOI21_X1   g07813(.A1(\A[854] ), .A2(\A[855] ), .B(\A[853] ), .ZN(new_n8816_));
  NOR2_X1    g07814(.A1(new_n8816_), .A2(new_n8800_), .ZN(new_n8817_));
  NOR3_X1    g07815(.A1(new_n8817_), .A2(new_n8810_), .A3(new_n8815_), .ZN(new_n8818_));
  NOR2_X1    g07816(.A1(new_n8815_), .A2(new_n8810_), .ZN(new_n8819_));
  NOR3_X1    g07817(.A1(new_n8819_), .A2(new_n8800_), .A3(new_n8816_), .ZN(new_n8820_));
  NOR2_X1    g07818(.A1(new_n8818_), .A2(new_n8820_), .ZN(new_n8821_));
  XOR2_X1    g07819(.A1(new_n8814_), .A2(new_n8821_), .Z(new_n8822_));
  INV_X1     g07820(.I(\A[855] ), .ZN(new_n8823_));
  NAND2_X1   g07821(.A1(new_n8823_), .A2(\A[854] ), .ZN(new_n8824_));
  AOI21_X1   g07822(.A1(new_n8795_), .A2(new_n8824_), .B(new_n8799_), .ZN(new_n8825_));
  INV_X1     g07823(.I(new_n8800_), .ZN(new_n8826_));
  AOI21_X1   g07824(.A1(new_n8826_), .A2(new_n8801_), .B(\A[853] ), .ZN(new_n8827_));
  NAND2_X1   g07825(.A1(new_n8806_), .A2(\A[858] ), .ZN(new_n8828_));
  NAND2_X1   g07826(.A1(new_n8804_), .A2(\A[857] ), .ZN(new_n8829_));
  AOI21_X1   g07827(.A1(new_n8828_), .A2(new_n8829_), .B(new_n8809_), .ZN(new_n8830_));
  INV_X1     g07828(.I(new_n8810_), .ZN(new_n8831_));
  AOI21_X1   g07829(.A1(new_n8831_), .A2(new_n8811_), .B(\A[856] ), .ZN(new_n8832_));
  OAI22_X1   g07830(.A1(new_n8825_), .A2(new_n8827_), .B1(new_n8832_), .B2(new_n8830_), .ZN(new_n8833_));
  NAND2_X1   g07831(.A1(new_n8814_), .A2(new_n8833_), .ZN(new_n8834_));
  OAI22_X1   g07832(.A1(new_n8766_), .A2(new_n8770_), .B1(new_n8780_), .B2(new_n8776_), .ZN(new_n8835_));
  NAND2_X1   g07833(.A1(new_n8781_), .A2(new_n8835_), .ZN(new_n8836_));
  NOR2_X1    g07834(.A1(new_n8836_), .A2(new_n8834_), .ZN(new_n8837_));
  OAI21_X1   g07835(.A1(new_n8822_), .A2(new_n8837_), .B(new_n8793_), .ZN(new_n8838_));
  NOR4_X1    g07836(.A1(new_n8825_), .A2(new_n8827_), .A3(new_n8832_), .A4(new_n8830_), .ZN(new_n8839_));
  XOR2_X1    g07837(.A1(new_n8839_), .A2(new_n8821_), .Z(new_n8840_));
  NAND4_X1   g07838(.A1(new_n8781_), .A2(new_n8814_), .A3(new_n8833_), .A4(new_n8835_), .ZN(new_n8841_));
  NOR2_X1    g07839(.A1(new_n8840_), .A2(new_n8841_), .ZN(new_n8842_));
  NOR2_X1    g07840(.A1(new_n8838_), .A2(new_n8842_), .ZN(new_n8843_));
  NAND2_X1   g07841(.A1(new_n8840_), .A2(new_n8841_), .ZN(new_n8844_));
  NAND2_X1   g07842(.A1(new_n8822_), .A2(new_n8837_), .ZN(new_n8845_));
  AOI21_X1   g07843(.A1(new_n8845_), .A2(new_n8844_), .B(new_n8793_), .ZN(new_n8846_));
  NOR2_X1    g07844(.A1(new_n8846_), .A2(new_n8843_), .ZN(new_n8847_));
  INV_X1     g07845(.I(new_n8847_), .ZN(new_n8848_));
  INV_X1     g07846(.I(\A[865] ), .ZN(new_n8849_));
  INV_X1     g07847(.I(\A[866] ), .ZN(new_n8850_));
  NAND2_X1   g07848(.A1(new_n8850_), .A2(\A[867] ), .ZN(new_n8851_));
  INV_X1     g07849(.I(\A[867] ), .ZN(new_n8852_));
  NAND2_X1   g07850(.A1(new_n8852_), .A2(\A[866] ), .ZN(new_n8853_));
  AOI21_X1   g07851(.A1(new_n8851_), .A2(new_n8853_), .B(new_n8849_), .ZN(new_n8854_));
  NAND2_X1   g07852(.A1(\A[866] ), .A2(\A[867] ), .ZN(new_n8855_));
  NOR2_X1    g07853(.A1(\A[866] ), .A2(\A[867] ), .ZN(new_n8856_));
  INV_X1     g07854(.I(new_n8856_), .ZN(new_n8857_));
  AOI21_X1   g07855(.A1(new_n8857_), .A2(new_n8855_), .B(\A[865] ), .ZN(new_n8858_));
  NOR2_X1    g07856(.A1(new_n8858_), .A2(new_n8854_), .ZN(new_n8859_));
  INV_X1     g07857(.I(\A[870] ), .ZN(new_n8860_));
  NOR2_X1    g07858(.A1(new_n8860_), .A2(\A[869] ), .ZN(new_n8861_));
  INV_X1     g07859(.I(\A[869] ), .ZN(new_n8862_));
  NOR2_X1    g07860(.A1(new_n8862_), .A2(\A[870] ), .ZN(new_n8863_));
  OAI21_X1   g07861(.A1(new_n8861_), .A2(new_n8863_), .B(\A[868] ), .ZN(new_n8864_));
  INV_X1     g07862(.I(\A[868] ), .ZN(new_n8865_));
  NAND2_X1   g07863(.A1(\A[869] ), .A2(\A[870] ), .ZN(new_n8866_));
  INV_X1     g07864(.I(new_n8866_), .ZN(new_n8867_));
  NOR2_X1    g07865(.A1(\A[869] ), .A2(\A[870] ), .ZN(new_n8868_));
  OAI21_X1   g07866(.A1(new_n8867_), .A2(new_n8868_), .B(new_n8865_), .ZN(new_n8869_));
  NAND2_X1   g07867(.A1(new_n8864_), .A2(new_n8869_), .ZN(new_n8870_));
  NAND2_X1   g07868(.A1(new_n8859_), .A2(new_n8870_), .ZN(new_n8871_));
  NOR2_X1    g07869(.A1(new_n8852_), .A2(\A[866] ), .ZN(new_n8872_));
  NOR2_X1    g07870(.A1(new_n8850_), .A2(\A[867] ), .ZN(new_n8873_));
  OAI21_X1   g07871(.A1(new_n8872_), .A2(new_n8873_), .B(\A[865] ), .ZN(new_n8874_));
  INV_X1     g07872(.I(new_n8855_), .ZN(new_n8875_));
  OAI21_X1   g07873(.A1(new_n8875_), .A2(new_n8856_), .B(new_n8849_), .ZN(new_n8876_));
  NAND2_X1   g07874(.A1(new_n8874_), .A2(new_n8876_), .ZN(new_n8877_));
  NAND2_X1   g07875(.A1(new_n8862_), .A2(\A[870] ), .ZN(new_n8878_));
  NAND2_X1   g07876(.A1(new_n8860_), .A2(\A[869] ), .ZN(new_n8879_));
  AOI21_X1   g07877(.A1(new_n8878_), .A2(new_n8879_), .B(new_n8865_), .ZN(new_n8880_));
  INV_X1     g07878(.I(new_n8868_), .ZN(new_n8881_));
  AOI21_X1   g07879(.A1(new_n8881_), .A2(new_n8866_), .B(\A[868] ), .ZN(new_n8882_));
  NOR2_X1    g07880(.A1(new_n8882_), .A2(new_n8880_), .ZN(new_n8883_));
  NAND2_X1   g07881(.A1(new_n8883_), .A2(new_n8877_), .ZN(new_n8884_));
  NAND2_X1   g07882(.A1(new_n8871_), .A2(new_n8884_), .ZN(new_n8885_));
  INV_X1     g07883(.I(\A[859] ), .ZN(new_n8886_));
  INV_X1     g07884(.I(\A[860] ), .ZN(new_n8887_));
  NAND2_X1   g07885(.A1(new_n8887_), .A2(\A[861] ), .ZN(new_n8888_));
  INV_X1     g07886(.I(\A[861] ), .ZN(new_n8889_));
  NAND2_X1   g07887(.A1(new_n8889_), .A2(\A[860] ), .ZN(new_n8890_));
  AOI21_X1   g07888(.A1(new_n8888_), .A2(new_n8890_), .B(new_n8886_), .ZN(new_n8891_));
  NAND2_X1   g07889(.A1(\A[860] ), .A2(\A[861] ), .ZN(new_n8892_));
  NOR2_X1    g07890(.A1(\A[860] ), .A2(\A[861] ), .ZN(new_n8893_));
  INV_X1     g07891(.I(new_n8893_), .ZN(new_n8894_));
  AOI21_X1   g07892(.A1(new_n8894_), .A2(new_n8892_), .B(\A[859] ), .ZN(new_n8895_));
  NOR2_X1    g07893(.A1(new_n8895_), .A2(new_n8891_), .ZN(new_n8896_));
  INV_X1     g07894(.I(\A[862] ), .ZN(new_n8897_));
  INV_X1     g07895(.I(\A[863] ), .ZN(new_n8898_));
  NAND2_X1   g07896(.A1(new_n8898_), .A2(\A[864] ), .ZN(new_n8899_));
  INV_X1     g07897(.I(\A[864] ), .ZN(new_n8900_));
  NAND2_X1   g07898(.A1(new_n8900_), .A2(\A[863] ), .ZN(new_n8901_));
  AOI21_X1   g07899(.A1(new_n8899_), .A2(new_n8901_), .B(new_n8897_), .ZN(new_n8902_));
  NAND2_X1   g07900(.A1(\A[863] ), .A2(\A[864] ), .ZN(new_n8903_));
  NOR2_X1    g07901(.A1(\A[863] ), .A2(\A[864] ), .ZN(new_n8904_));
  INV_X1     g07902(.I(new_n8904_), .ZN(new_n8905_));
  AOI21_X1   g07903(.A1(new_n8905_), .A2(new_n8903_), .B(\A[862] ), .ZN(new_n8906_));
  NOR2_X1    g07904(.A1(new_n8906_), .A2(new_n8902_), .ZN(new_n8907_));
  NAND2_X1   g07905(.A1(new_n8896_), .A2(new_n8907_), .ZN(new_n8908_));
  NOR2_X1    g07906(.A1(new_n8889_), .A2(\A[860] ), .ZN(new_n8909_));
  NOR2_X1    g07907(.A1(new_n8887_), .A2(\A[861] ), .ZN(new_n8910_));
  OAI21_X1   g07908(.A1(new_n8909_), .A2(new_n8910_), .B(\A[859] ), .ZN(new_n8911_));
  INV_X1     g07909(.I(new_n8892_), .ZN(new_n8912_));
  OAI21_X1   g07910(.A1(new_n8912_), .A2(new_n8893_), .B(new_n8886_), .ZN(new_n8913_));
  NAND2_X1   g07911(.A1(new_n8911_), .A2(new_n8913_), .ZN(new_n8914_));
  NOR2_X1    g07912(.A1(new_n8900_), .A2(\A[863] ), .ZN(new_n8915_));
  NOR2_X1    g07913(.A1(new_n8898_), .A2(\A[864] ), .ZN(new_n8916_));
  OAI21_X1   g07914(.A1(new_n8915_), .A2(new_n8916_), .B(\A[862] ), .ZN(new_n8917_));
  INV_X1     g07915(.I(new_n8903_), .ZN(new_n8918_));
  OAI21_X1   g07916(.A1(new_n8918_), .A2(new_n8904_), .B(new_n8897_), .ZN(new_n8919_));
  NAND2_X1   g07917(.A1(new_n8917_), .A2(new_n8919_), .ZN(new_n8920_));
  NAND2_X1   g07918(.A1(new_n8914_), .A2(new_n8920_), .ZN(new_n8921_));
  NAND2_X1   g07919(.A1(new_n8908_), .A2(new_n8921_), .ZN(new_n8922_));
  AOI21_X1   g07920(.A1(new_n8865_), .A2(new_n8866_), .B(new_n8868_), .ZN(new_n8923_));
  NAND4_X1   g07921(.A1(new_n8874_), .A2(new_n8876_), .A3(new_n8864_), .A4(new_n8869_), .ZN(new_n8924_));
  AOI21_X1   g07922(.A1(new_n8849_), .A2(new_n8855_), .B(new_n8856_), .ZN(new_n8925_));
  INV_X1     g07923(.I(new_n8925_), .ZN(new_n8926_));
  NOR2_X1    g07924(.A1(new_n8924_), .A2(new_n8926_), .ZN(new_n8927_));
  NAND2_X1   g07925(.A1(new_n8927_), .A2(new_n8923_), .ZN(new_n8928_));
  NAND3_X1   g07926(.A1(new_n8928_), .A2(new_n8885_), .A3(new_n8922_), .ZN(new_n8929_));
  NOR2_X1    g07927(.A1(new_n8883_), .A2(new_n8877_), .ZN(new_n8930_));
  NOR2_X1    g07928(.A1(new_n8859_), .A2(new_n8870_), .ZN(new_n8931_));
  NOR2_X1    g07929(.A1(new_n8930_), .A2(new_n8931_), .ZN(new_n8932_));
  AOI21_X1   g07930(.A1(new_n8897_), .A2(new_n8903_), .B(new_n8904_), .ZN(new_n8933_));
  AOI21_X1   g07931(.A1(new_n8886_), .A2(new_n8892_), .B(new_n8893_), .ZN(new_n8934_));
  NAND3_X1   g07932(.A1(new_n8932_), .A2(new_n8908_), .A3(new_n8921_), .ZN(new_n8935_));
  NAND2_X1   g07933(.A1(new_n8929_), .A2(new_n8935_), .ZN(new_n8936_));
  NOR2_X1    g07934(.A1(new_n8827_), .A2(new_n8825_), .ZN(new_n8937_));
  NAND2_X1   g07935(.A1(new_n8808_), .A2(new_n8813_), .ZN(new_n8938_));
  XOR2_X1    g07936(.A1(new_n8937_), .A2(new_n8938_), .Z(new_n8939_));
  AOI21_X1   g07937(.A1(new_n8836_), .A2(new_n8939_), .B(new_n8837_), .ZN(new_n8940_));
  NAND2_X1   g07938(.A1(new_n8936_), .A2(new_n8940_), .ZN(new_n8941_));
  NOR2_X1    g07939(.A1(new_n8914_), .A2(new_n8920_), .ZN(new_n8942_));
  NOR2_X1    g07940(.A1(new_n8933_), .A2(new_n8934_), .ZN(new_n8943_));
  AND2_X2    g07941(.A1(new_n8933_), .A2(new_n8934_), .Z(new_n8944_));
  NOR2_X1    g07942(.A1(new_n8944_), .A2(new_n8943_), .ZN(new_n8945_));
  XOR2_X1    g07943(.A1(new_n8942_), .A2(new_n8945_), .Z(new_n8946_));
  XNOR2_X1   g07944(.A1(new_n8923_), .A2(new_n8925_), .ZN(new_n8947_));
  XOR2_X1    g07945(.A1(new_n8947_), .A2(new_n8924_), .Z(new_n8948_));
  NAND3_X1   g07946(.A1(new_n8885_), .A2(new_n8923_), .A3(new_n8925_), .ZN(new_n8949_));
  NOR2_X1    g07947(.A1(new_n8932_), .A2(new_n8922_), .ZN(new_n8950_));
  AOI21_X1   g07948(.A1(new_n8948_), .A2(new_n8949_), .B(new_n8950_), .ZN(new_n8951_));
  INV_X1     g07949(.I(new_n8923_), .ZN(new_n8952_));
  NOR3_X1    g07950(.A1(new_n8932_), .A2(new_n8952_), .A3(new_n8926_), .ZN(new_n8953_));
  NOR4_X1    g07951(.A1(new_n8953_), .A2(new_n8932_), .A3(new_n8922_), .A4(new_n8947_), .ZN(new_n8954_));
  OAI21_X1   g07952(.A1(new_n8951_), .A2(new_n8954_), .B(new_n8946_), .ZN(new_n8955_));
  INV_X1     g07953(.I(new_n8946_), .ZN(new_n8956_));
  NAND2_X1   g07954(.A1(new_n8947_), .A2(new_n8924_), .ZN(new_n8957_));
  INV_X1     g07955(.I(new_n8924_), .ZN(new_n8958_));
  NAND2_X1   g07956(.A1(new_n8926_), .A2(new_n8923_), .ZN(new_n8959_));
  NAND2_X1   g07957(.A1(new_n8952_), .A2(new_n8925_), .ZN(new_n8960_));
  NAND2_X1   g07958(.A1(new_n8959_), .A2(new_n8960_), .ZN(new_n8961_));
  NAND2_X1   g07959(.A1(new_n8958_), .A2(new_n8961_), .ZN(new_n8962_));
  NAND2_X1   g07960(.A1(new_n8962_), .A2(new_n8957_), .ZN(new_n8963_));
  NOR2_X1    g07961(.A1(new_n8896_), .A2(new_n8907_), .ZN(new_n8964_));
  NOR2_X1    g07962(.A1(new_n8964_), .A2(new_n8942_), .ZN(new_n8965_));
  NAND2_X1   g07963(.A1(new_n8965_), .A2(new_n8885_), .ZN(new_n8966_));
  OAI21_X1   g07964(.A1(new_n8953_), .A2(new_n8963_), .B(new_n8966_), .ZN(new_n8967_));
  NAND3_X1   g07965(.A1(new_n8948_), .A2(new_n8950_), .A3(new_n8949_), .ZN(new_n8968_));
  NAND3_X1   g07966(.A1(new_n8967_), .A2(new_n8968_), .A3(new_n8956_), .ZN(new_n8969_));
  AOI21_X1   g07967(.A1(new_n8955_), .A2(new_n8969_), .B(new_n8941_), .ZN(new_n8970_));
  AND2_X2    g07968(.A1(new_n8936_), .A2(new_n8940_), .Z(new_n8971_));
  NAND4_X1   g07969(.A1(new_n8949_), .A2(new_n8885_), .A3(new_n8965_), .A4(new_n8961_), .ZN(new_n8972_));
  AOI21_X1   g07970(.A1(new_n8967_), .A2(new_n8972_), .B(new_n8956_), .ZN(new_n8973_));
  NOR3_X1    g07971(.A1(new_n8953_), .A2(new_n8966_), .A3(new_n8963_), .ZN(new_n8974_));
  NOR3_X1    g07972(.A1(new_n8951_), .A2(new_n8974_), .A3(new_n8946_), .ZN(new_n8975_));
  NOR3_X1    g07973(.A1(new_n8971_), .A2(new_n8975_), .A3(new_n8973_), .ZN(new_n8976_));
  NOR3_X1    g07974(.A1(new_n8976_), .A2(new_n8970_), .A3(new_n8848_), .ZN(new_n8977_));
  OAI21_X1   g07975(.A1(new_n8975_), .A2(new_n8973_), .B(new_n8971_), .ZN(new_n8978_));
  NAND3_X1   g07976(.A1(new_n8955_), .A2(new_n8969_), .A3(new_n8941_), .ZN(new_n8979_));
  AOI21_X1   g07977(.A1(new_n8978_), .A2(new_n8979_), .B(new_n8847_), .ZN(new_n8980_));
  NOR2_X1    g07978(.A1(new_n8980_), .A2(new_n8977_), .ZN(new_n8981_));
  INV_X1     g07979(.I(\A[889] ), .ZN(new_n8982_));
  INV_X1     g07980(.I(\A[890] ), .ZN(new_n8983_));
  NAND2_X1   g07981(.A1(new_n8983_), .A2(\A[891] ), .ZN(new_n8984_));
  INV_X1     g07982(.I(\A[891] ), .ZN(new_n8985_));
  NAND2_X1   g07983(.A1(new_n8985_), .A2(\A[890] ), .ZN(new_n8986_));
  AOI21_X1   g07984(.A1(new_n8984_), .A2(new_n8986_), .B(new_n8982_), .ZN(new_n8987_));
  NAND2_X1   g07985(.A1(\A[890] ), .A2(\A[891] ), .ZN(new_n8988_));
  NOR2_X1    g07986(.A1(\A[890] ), .A2(\A[891] ), .ZN(new_n8989_));
  INV_X1     g07987(.I(new_n8989_), .ZN(new_n8990_));
  AOI21_X1   g07988(.A1(new_n8990_), .A2(new_n8988_), .B(\A[889] ), .ZN(new_n8991_));
  NOR2_X1    g07989(.A1(new_n8991_), .A2(new_n8987_), .ZN(new_n8992_));
  INV_X1     g07990(.I(\A[894] ), .ZN(new_n8993_));
  NOR2_X1    g07991(.A1(new_n8993_), .A2(\A[893] ), .ZN(new_n8994_));
  INV_X1     g07992(.I(\A[893] ), .ZN(new_n8995_));
  NOR2_X1    g07993(.A1(new_n8995_), .A2(\A[894] ), .ZN(new_n8996_));
  OAI21_X1   g07994(.A1(new_n8994_), .A2(new_n8996_), .B(\A[892] ), .ZN(new_n8997_));
  INV_X1     g07995(.I(\A[892] ), .ZN(new_n8998_));
  NAND2_X1   g07996(.A1(\A[893] ), .A2(\A[894] ), .ZN(new_n8999_));
  INV_X1     g07997(.I(new_n8999_), .ZN(new_n9000_));
  NOR2_X1    g07998(.A1(\A[893] ), .A2(\A[894] ), .ZN(new_n9001_));
  OAI21_X1   g07999(.A1(new_n9000_), .A2(new_n9001_), .B(new_n8998_), .ZN(new_n9002_));
  NAND2_X1   g08000(.A1(new_n8997_), .A2(new_n9002_), .ZN(new_n9003_));
  NAND2_X1   g08001(.A1(new_n8992_), .A2(new_n9003_), .ZN(new_n9004_));
  NOR2_X1    g08002(.A1(new_n8985_), .A2(\A[890] ), .ZN(new_n9005_));
  NOR2_X1    g08003(.A1(new_n8983_), .A2(\A[891] ), .ZN(new_n9006_));
  OAI21_X1   g08004(.A1(new_n9005_), .A2(new_n9006_), .B(\A[889] ), .ZN(new_n9007_));
  INV_X1     g08005(.I(new_n8988_), .ZN(new_n9008_));
  OAI21_X1   g08006(.A1(new_n9008_), .A2(new_n8989_), .B(new_n8982_), .ZN(new_n9009_));
  NAND2_X1   g08007(.A1(new_n9007_), .A2(new_n9009_), .ZN(new_n9010_));
  NAND2_X1   g08008(.A1(new_n8995_), .A2(\A[894] ), .ZN(new_n9011_));
  NAND2_X1   g08009(.A1(new_n8993_), .A2(\A[893] ), .ZN(new_n9012_));
  AOI21_X1   g08010(.A1(new_n9011_), .A2(new_n9012_), .B(new_n8998_), .ZN(new_n9013_));
  INV_X1     g08011(.I(new_n9001_), .ZN(new_n9014_));
  AOI21_X1   g08012(.A1(new_n9014_), .A2(new_n8999_), .B(\A[892] ), .ZN(new_n9015_));
  NOR2_X1    g08013(.A1(new_n9015_), .A2(new_n9013_), .ZN(new_n9016_));
  NAND2_X1   g08014(.A1(new_n9016_), .A2(new_n9010_), .ZN(new_n9017_));
  NAND2_X1   g08015(.A1(new_n9004_), .A2(new_n9017_), .ZN(new_n9018_));
  INV_X1     g08016(.I(\A[883] ), .ZN(new_n9019_));
  INV_X1     g08017(.I(\A[884] ), .ZN(new_n9020_));
  NAND2_X1   g08018(.A1(new_n9020_), .A2(\A[885] ), .ZN(new_n9021_));
  INV_X1     g08019(.I(\A[885] ), .ZN(new_n9022_));
  NAND2_X1   g08020(.A1(new_n9022_), .A2(\A[884] ), .ZN(new_n9023_));
  AOI21_X1   g08021(.A1(new_n9021_), .A2(new_n9023_), .B(new_n9019_), .ZN(new_n9024_));
  NAND2_X1   g08022(.A1(\A[884] ), .A2(\A[885] ), .ZN(new_n9025_));
  NOR2_X1    g08023(.A1(\A[884] ), .A2(\A[885] ), .ZN(new_n9026_));
  INV_X1     g08024(.I(new_n9026_), .ZN(new_n9027_));
  AOI21_X1   g08025(.A1(new_n9027_), .A2(new_n9025_), .B(\A[883] ), .ZN(new_n9028_));
  INV_X1     g08026(.I(\A[886] ), .ZN(new_n9029_));
  INV_X1     g08027(.I(\A[887] ), .ZN(new_n9030_));
  NAND2_X1   g08028(.A1(new_n9030_), .A2(\A[888] ), .ZN(new_n9031_));
  INV_X1     g08029(.I(\A[888] ), .ZN(new_n9032_));
  NAND2_X1   g08030(.A1(new_n9032_), .A2(\A[887] ), .ZN(new_n9033_));
  AOI21_X1   g08031(.A1(new_n9031_), .A2(new_n9033_), .B(new_n9029_), .ZN(new_n9034_));
  NAND2_X1   g08032(.A1(\A[887] ), .A2(\A[888] ), .ZN(new_n9035_));
  NOR2_X1    g08033(.A1(\A[887] ), .A2(\A[888] ), .ZN(new_n9036_));
  INV_X1     g08034(.I(new_n9036_), .ZN(new_n9037_));
  AOI21_X1   g08035(.A1(new_n9037_), .A2(new_n9035_), .B(\A[886] ), .ZN(new_n9038_));
  NOR4_X1    g08036(.A1(new_n9024_), .A2(new_n9028_), .A3(new_n9038_), .A4(new_n9034_), .ZN(new_n9039_));
  INV_X1     g08037(.I(new_n9021_), .ZN(new_n9040_));
  NOR2_X1    g08038(.A1(new_n9020_), .A2(\A[885] ), .ZN(new_n9041_));
  OAI21_X1   g08039(.A1(new_n9040_), .A2(new_n9041_), .B(\A[883] ), .ZN(new_n9042_));
  INV_X1     g08040(.I(new_n9025_), .ZN(new_n9043_));
  OAI21_X1   g08041(.A1(new_n9043_), .A2(new_n9026_), .B(new_n9019_), .ZN(new_n9044_));
  NOR2_X1    g08042(.A1(new_n9032_), .A2(\A[887] ), .ZN(new_n9045_));
  NOR2_X1    g08043(.A1(new_n9030_), .A2(\A[888] ), .ZN(new_n9046_));
  OAI21_X1   g08044(.A1(new_n9045_), .A2(new_n9046_), .B(\A[886] ), .ZN(new_n9047_));
  INV_X1     g08045(.I(new_n9035_), .ZN(new_n9048_));
  OAI21_X1   g08046(.A1(new_n9048_), .A2(new_n9036_), .B(new_n9029_), .ZN(new_n9049_));
  AOI22_X1   g08047(.A1(new_n9042_), .A2(new_n9044_), .B1(new_n9049_), .B2(new_n9047_), .ZN(new_n9050_));
  NOR2_X1    g08048(.A1(new_n9050_), .A2(new_n9039_), .ZN(new_n9051_));
  AOI21_X1   g08049(.A1(new_n8998_), .A2(new_n8999_), .B(new_n9001_), .ZN(new_n9052_));
  NAND4_X1   g08050(.A1(new_n9007_), .A2(new_n9009_), .A3(new_n8997_), .A4(new_n9002_), .ZN(new_n9053_));
  AOI21_X1   g08051(.A1(new_n8982_), .A2(new_n8988_), .B(new_n8989_), .ZN(new_n9054_));
  INV_X1     g08052(.I(new_n9054_), .ZN(new_n9055_));
  NOR2_X1    g08053(.A1(new_n9053_), .A2(new_n9055_), .ZN(new_n9056_));
  AOI21_X1   g08054(.A1(new_n9052_), .A2(new_n9056_), .B(new_n9051_), .ZN(new_n9057_));
  NAND4_X1   g08055(.A1(new_n9042_), .A2(new_n9044_), .A3(new_n9049_), .A4(new_n9047_), .ZN(new_n9058_));
  AOI21_X1   g08056(.A1(new_n9029_), .A2(new_n9035_), .B(new_n9036_), .ZN(new_n9059_));
  INV_X1     g08057(.I(new_n9059_), .ZN(new_n9060_));
  AOI21_X1   g08058(.A1(new_n9019_), .A2(new_n9025_), .B(new_n9026_), .ZN(new_n9061_));
  INV_X1     g08059(.I(new_n9061_), .ZN(new_n9062_));
  NOR3_X1    g08060(.A1(new_n9058_), .A2(new_n9060_), .A3(new_n9062_), .ZN(new_n9063_));
  NOR2_X1    g08061(.A1(new_n9018_), .A2(new_n9063_), .ZN(new_n9064_));
  AOI22_X1   g08062(.A1(new_n9018_), .A2(new_n9057_), .B1(new_n9064_), .B2(new_n9051_), .ZN(new_n9065_));
  INV_X1     g08063(.I(\A[873] ), .ZN(new_n9066_));
  NOR2_X1    g08064(.A1(new_n9066_), .A2(\A[872] ), .ZN(new_n9067_));
  INV_X1     g08065(.I(\A[872] ), .ZN(new_n9068_));
  NOR2_X1    g08066(.A1(new_n9068_), .A2(\A[873] ), .ZN(new_n9069_));
  OAI21_X1   g08067(.A1(new_n9067_), .A2(new_n9069_), .B(\A[871] ), .ZN(new_n9070_));
  INV_X1     g08068(.I(\A[871] ), .ZN(new_n9071_));
  NAND2_X1   g08069(.A1(\A[872] ), .A2(\A[873] ), .ZN(new_n9072_));
  INV_X1     g08070(.I(new_n9072_), .ZN(new_n9073_));
  NOR2_X1    g08071(.A1(\A[872] ), .A2(\A[873] ), .ZN(new_n9074_));
  OAI21_X1   g08072(.A1(new_n9073_), .A2(new_n9074_), .B(new_n9071_), .ZN(new_n9075_));
  INV_X1     g08073(.I(\A[876] ), .ZN(new_n9076_));
  NOR2_X1    g08074(.A1(new_n9076_), .A2(\A[875] ), .ZN(new_n9077_));
  INV_X1     g08075(.I(\A[875] ), .ZN(new_n9078_));
  NOR2_X1    g08076(.A1(new_n9078_), .A2(\A[876] ), .ZN(new_n9079_));
  OAI21_X1   g08077(.A1(new_n9077_), .A2(new_n9079_), .B(\A[874] ), .ZN(new_n9080_));
  INV_X1     g08078(.I(\A[874] ), .ZN(new_n9081_));
  NAND2_X1   g08079(.A1(\A[875] ), .A2(\A[876] ), .ZN(new_n9082_));
  INV_X1     g08080(.I(new_n9082_), .ZN(new_n9083_));
  NOR2_X1    g08081(.A1(\A[875] ), .A2(\A[876] ), .ZN(new_n9084_));
  OAI21_X1   g08082(.A1(new_n9083_), .A2(new_n9084_), .B(new_n9081_), .ZN(new_n9085_));
  NAND4_X1   g08083(.A1(new_n9070_), .A2(new_n9075_), .A3(new_n9080_), .A4(new_n9085_), .ZN(new_n9086_));
  INV_X1     g08084(.I(new_n9067_), .ZN(new_n9087_));
  NAND2_X1   g08085(.A1(new_n9066_), .A2(\A[872] ), .ZN(new_n9088_));
  AOI21_X1   g08086(.A1(new_n9087_), .A2(new_n9088_), .B(new_n9071_), .ZN(new_n9089_));
  INV_X1     g08087(.I(new_n9074_), .ZN(new_n9090_));
  AOI21_X1   g08088(.A1(new_n9090_), .A2(new_n9072_), .B(\A[871] ), .ZN(new_n9091_));
  NAND2_X1   g08089(.A1(new_n9078_), .A2(\A[876] ), .ZN(new_n9092_));
  NAND2_X1   g08090(.A1(new_n9076_), .A2(\A[875] ), .ZN(new_n9093_));
  AOI21_X1   g08091(.A1(new_n9092_), .A2(new_n9093_), .B(new_n9081_), .ZN(new_n9094_));
  INV_X1     g08092(.I(new_n9084_), .ZN(new_n9095_));
  AOI21_X1   g08093(.A1(new_n9095_), .A2(new_n9082_), .B(\A[874] ), .ZN(new_n9096_));
  OAI22_X1   g08094(.A1(new_n9089_), .A2(new_n9091_), .B1(new_n9096_), .B2(new_n9094_), .ZN(new_n9097_));
  NAND2_X1   g08095(.A1(new_n9097_), .A2(new_n9086_), .ZN(new_n9098_));
  INV_X1     g08096(.I(\A[879] ), .ZN(new_n9099_));
  NOR2_X1    g08097(.A1(new_n9099_), .A2(\A[878] ), .ZN(new_n9100_));
  INV_X1     g08098(.I(\A[878] ), .ZN(new_n9101_));
  NOR2_X1    g08099(.A1(new_n9101_), .A2(\A[879] ), .ZN(new_n9102_));
  OAI21_X1   g08100(.A1(new_n9100_), .A2(new_n9102_), .B(\A[877] ), .ZN(new_n9103_));
  INV_X1     g08101(.I(\A[877] ), .ZN(new_n9104_));
  NAND2_X1   g08102(.A1(\A[878] ), .A2(\A[879] ), .ZN(new_n9105_));
  INV_X1     g08103(.I(new_n9105_), .ZN(new_n9106_));
  NOR2_X1    g08104(.A1(\A[878] ), .A2(\A[879] ), .ZN(new_n9107_));
  OAI21_X1   g08105(.A1(new_n9106_), .A2(new_n9107_), .B(new_n9104_), .ZN(new_n9108_));
  NAND2_X1   g08106(.A1(new_n9103_), .A2(new_n9108_), .ZN(new_n9109_));
  INV_X1     g08107(.I(\A[880] ), .ZN(new_n9110_));
  INV_X1     g08108(.I(\A[881] ), .ZN(new_n9111_));
  NAND2_X1   g08109(.A1(new_n9111_), .A2(\A[882] ), .ZN(new_n9112_));
  INV_X1     g08110(.I(\A[882] ), .ZN(new_n9113_));
  NAND2_X1   g08111(.A1(new_n9113_), .A2(\A[881] ), .ZN(new_n9114_));
  AOI21_X1   g08112(.A1(new_n9112_), .A2(new_n9114_), .B(new_n9110_), .ZN(new_n9115_));
  NAND2_X1   g08113(.A1(\A[881] ), .A2(\A[882] ), .ZN(new_n9116_));
  NOR2_X1    g08114(.A1(\A[881] ), .A2(\A[882] ), .ZN(new_n9117_));
  INV_X1     g08115(.I(new_n9117_), .ZN(new_n9118_));
  AOI21_X1   g08116(.A1(new_n9118_), .A2(new_n9116_), .B(\A[880] ), .ZN(new_n9119_));
  NOR2_X1    g08117(.A1(new_n9119_), .A2(new_n9115_), .ZN(new_n9120_));
  NOR2_X1    g08118(.A1(new_n9120_), .A2(new_n9109_), .ZN(new_n9121_));
  NAND2_X1   g08119(.A1(new_n9101_), .A2(\A[879] ), .ZN(new_n9122_));
  NAND2_X1   g08120(.A1(new_n9099_), .A2(\A[878] ), .ZN(new_n9123_));
  AOI21_X1   g08121(.A1(new_n9122_), .A2(new_n9123_), .B(new_n9104_), .ZN(new_n9124_));
  INV_X1     g08122(.I(new_n9107_), .ZN(new_n9125_));
  AOI21_X1   g08123(.A1(new_n9125_), .A2(new_n9105_), .B(\A[877] ), .ZN(new_n9126_));
  NOR2_X1    g08124(.A1(new_n9126_), .A2(new_n9124_), .ZN(new_n9127_));
  NOR2_X1    g08125(.A1(new_n9113_), .A2(\A[881] ), .ZN(new_n9128_));
  NOR2_X1    g08126(.A1(new_n9111_), .A2(\A[882] ), .ZN(new_n9129_));
  OAI21_X1   g08127(.A1(new_n9128_), .A2(new_n9129_), .B(\A[880] ), .ZN(new_n9130_));
  INV_X1     g08128(.I(new_n9116_), .ZN(new_n9131_));
  OAI21_X1   g08129(.A1(new_n9131_), .A2(new_n9117_), .B(new_n9110_), .ZN(new_n9132_));
  NAND2_X1   g08130(.A1(new_n9130_), .A2(new_n9132_), .ZN(new_n9133_));
  NOR2_X1    g08131(.A1(new_n9127_), .A2(new_n9133_), .ZN(new_n9134_));
  NOR2_X1    g08132(.A1(new_n9121_), .A2(new_n9134_), .ZN(new_n9135_));
  AOI21_X1   g08133(.A1(new_n9081_), .A2(new_n9082_), .B(new_n9084_), .ZN(new_n9136_));
  AOI21_X1   g08134(.A1(new_n9071_), .A2(new_n9072_), .B(new_n9074_), .ZN(new_n9137_));
  NAND2_X1   g08135(.A1(new_n9097_), .A2(new_n9086_), .ZN(new_n9138_));
  NAND2_X1   g08136(.A1(new_n9135_), .A2(new_n9138_), .ZN(new_n9139_));
  OAI21_X1   g08137(.A1(new_n9098_), .A2(new_n9135_), .B(new_n9139_), .ZN(new_n9140_));
  NOR2_X1    g08138(.A1(new_n9065_), .A2(new_n9140_), .ZN(new_n9141_));
  NOR2_X1    g08139(.A1(new_n9016_), .A2(new_n9010_), .ZN(new_n9142_));
  NOR2_X1    g08140(.A1(new_n8992_), .A2(new_n9003_), .ZN(new_n9143_));
  NOR2_X1    g08141(.A1(new_n9142_), .A2(new_n9143_), .ZN(new_n9144_));
  OAI22_X1   g08142(.A1(new_n9024_), .A2(new_n9028_), .B1(new_n9038_), .B2(new_n9034_), .ZN(new_n9145_));
  NAND2_X1   g08143(.A1(new_n9058_), .A2(new_n9145_), .ZN(new_n9146_));
  NAND2_X1   g08144(.A1(new_n9056_), .A2(new_n9052_), .ZN(new_n9147_));
  NAND2_X1   g08145(.A1(new_n9147_), .A2(new_n9146_), .ZN(new_n9148_));
  NAND3_X1   g08146(.A1(new_n9039_), .A2(new_n9059_), .A3(new_n9061_), .ZN(new_n9149_));
  NAND2_X1   g08147(.A1(new_n9144_), .A2(new_n9149_), .ZN(new_n9150_));
  OAI22_X1   g08148(.A1(new_n9148_), .A2(new_n9144_), .B1(new_n9150_), .B2(new_n9146_), .ZN(new_n9151_));
  NOR2_X1    g08149(.A1(new_n9135_), .A2(new_n9098_), .ZN(new_n9152_));
  AOI21_X1   g08150(.A1(new_n9135_), .A2(new_n9138_), .B(new_n9152_), .ZN(new_n9153_));
  NOR2_X1    g08151(.A1(new_n9151_), .A2(new_n9153_), .ZN(new_n9154_));
  NOR2_X1    g08152(.A1(new_n8936_), .A2(new_n8940_), .ZN(new_n9155_));
  NOR4_X1    g08153(.A1(new_n8971_), .A2(new_n9141_), .A3(new_n9154_), .A4(new_n9155_), .ZN(new_n9156_));
  NOR4_X1    g08154(.A1(new_n9089_), .A2(new_n9091_), .A3(new_n9096_), .A4(new_n9094_), .ZN(new_n9157_));
  XOR2_X1    g08155(.A1(new_n9136_), .A2(new_n9137_), .Z(new_n9158_));
  XOR2_X1    g08156(.A1(new_n9158_), .A2(new_n9157_), .Z(new_n9159_));
  INV_X1     g08157(.I(new_n9097_), .ZN(new_n9160_));
  NOR3_X1    g08158(.A1(new_n9135_), .A2(new_n9157_), .A3(new_n9160_), .ZN(new_n9161_));
  NOR2_X1    g08159(.A1(new_n9109_), .A2(new_n9133_), .ZN(new_n9162_));
  AOI21_X1   g08160(.A1(new_n9110_), .A2(new_n9116_), .B(new_n9117_), .ZN(new_n9163_));
  AOI21_X1   g08161(.A1(new_n9104_), .A2(new_n9105_), .B(new_n9107_), .ZN(new_n9164_));
  XOR2_X1    g08162(.A1(new_n9163_), .A2(new_n9164_), .Z(new_n9165_));
  XOR2_X1    g08163(.A1(new_n9162_), .A2(new_n9165_), .Z(new_n9166_));
  OAI21_X1   g08164(.A1(new_n9166_), .A2(new_n9161_), .B(new_n9159_), .ZN(new_n9167_));
  NAND2_X1   g08165(.A1(new_n9127_), .A2(new_n9133_), .ZN(new_n9168_));
  NAND2_X1   g08166(.A1(new_n9120_), .A2(new_n9109_), .ZN(new_n9169_));
  NAND2_X1   g08167(.A1(new_n9168_), .A2(new_n9169_), .ZN(new_n9170_));
  NAND3_X1   g08168(.A1(new_n9170_), .A2(new_n9086_), .A3(new_n9097_), .ZN(new_n9171_));
  NAND2_X1   g08169(.A1(new_n9163_), .A2(new_n9164_), .ZN(new_n9172_));
  OAI21_X1   g08170(.A1(new_n9135_), .A2(new_n9172_), .B(new_n9165_), .ZN(new_n9173_));
  NOR2_X1    g08171(.A1(new_n9173_), .A2(new_n9171_), .ZN(new_n9174_));
  NOR3_X1    g08172(.A1(new_n9165_), .A2(new_n9109_), .A3(new_n9133_), .ZN(new_n9175_));
  XNOR2_X1   g08173(.A1(new_n9163_), .A2(new_n9164_), .ZN(new_n9176_));
  NOR2_X1    g08174(.A1(new_n9162_), .A2(new_n9176_), .ZN(new_n9177_));
  NOR2_X1    g08175(.A1(new_n9177_), .A2(new_n9175_), .ZN(new_n9178_));
  XOR2_X1    g08176(.A1(new_n9171_), .A2(new_n9178_), .Z(new_n9179_));
  OAI22_X1   g08177(.A1(new_n9179_), .A2(new_n9159_), .B1(new_n9167_), .B2(new_n9174_), .ZN(new_n9180_));
  NOR2_X1    g08178(.A1(new_n9059_), .A2(new_n9061_), .ZN(new_n9181_));
  NOR2_X1    g08179(.A1(new_n9060_), .A2(new_n9062_), .ZN(new_n9182_));
  NOR2_X1    g08180(.A1(new_n9182_), .A2(new_n9181_), .ZN(new_n9183_));
  XOR2_X1    g08181(.A1(new_n9183_), .A2(new_n9058_), .Z(new_n9184_));
  XOR2_X1    g08182(.A1(new_n9052_), .A2(new_n9054_), .Z(new_n9185_));
  XOR2_X1    g08183(.A1(new_n9185_), .A2(new_n9053_), .Z(new_n9186_));
  INV_X1     g08184(.I(new_n9052_), .ZN(new_n9187_));
  NOR3_X1    g08185(.A1(new_n9144_), .A2(new_n9187_), .A3(new_n9055_), .ZN(new_n9188_));
  NAND2_X1   g08186(.A1(new_n9018_), .A2(new_n9051_), .ZN(new_n9189_));
  OAI21_X1   g08187(.A1(new_n9188_), .A2(new_n9186_), .B(new_n9189_), .ZN(new_n9190_));
  NAND3_X1   g08188(.A1(new_n9018_), .A2(new_n9052_), .A3(new_n9054_), .ZN(new_n9191_));
  NAND4_X1   g08189(.A1(new_n9191_), .A2(new_n9018_), .A3(new_n9051_), .A4(new_n9185_), .ZN(new_n9192_));
  AOI21_X1   g08190(.A1(new_n9190_), .A2(new_n9192_), .B(new_n9184_), .ZN(new_n9193_));
  INV_X1     g08191(.I(new_n9184_), .ZN(new_n9194_));
  INV_X1     g08192(.I(new_n9053_), .ZN(new_n9195_));
  NOR2_X1    g08193(.A1(new_n9195_), .A2(new_n9185_), .ZN(new_n9196_));
  XNOR2_X1   g08194(.A1(new_n9052_), .A2(new_n9054_), .ZN(new_n9197_));
  NOR2_X1    g08195(.A1(new_n9197_), .A2(new_n9053_), .ZN(new_n9198_));
  NOR2_X1    g08196(.A1(new_n9196_), .A2(new_n9198_), .ZN(new_n9199_));
  NOR2_X1    g08197(.A1(new_n9144_), .A2(new_n9146_), .ZN(new_n9200_));
  AOI21_X1   g08198(.A1(new_n9191_), .A2(new_n9199_), .B(new_n9200_), .ZN(new_n9201_));
  NOR3_X1    g08199(.A1(new_n9188_), .A2(new_n9186_), .A3(new_n9189_), .ZN(new_n9202_));
  NOR3_X1    g08200(.A1(new_n9202_), .A2(new_n9201_), .A3(new_n9194_), .ZN(new_n9203_));
  OAI21_X1   g08201(.A1(new_n9203_), .A2(new_n9193_), .B(new_n9141_), .ZN(new_n9204_));
  NAND2_X1   g08202(.A1(new_n9151_), .A2(new_n9153_), .ZN(new_n9205_));
  NOR4_X1    g08203(.A1(new_n9188_), .A2(new_n9144_), .A3(new_n9146_), .A4(new_n9197_), .ZN(new_n9206_));
  OAI21_X1   g08204(.A1(new_n9206_), .A2(new_n9201_), .B(new_n9194_), .ZN(new_n9207_));
  NAND3_X1   g08205(.A1(new_n9191_), .A2(new_n9199_), .A3(new_n9200_), .ZN(new_n9208_));
  NAND3_X1   g08206(.A1(new_n9190_), .A2(new_n9208_), .A3(new_n9184_), .ZN(new_n9209_));
  NAND3_X1   g08207(.A1(new_n9207_), .A2(new_n9209_), .A3(new_n9205_), .ZN(new_n9210_));
  AOI21_X1   g08208(.A1(new_n9204_), .A2(new_n9210_), .B(new_n9180_), .ZN(new_n9211_));
  XOR2_X1    g08209(.A1(new_n9158_), .A2(new_n9086_), .Z(new_n9212_));
  AOI21_X1   g08210(.A1(new_n9171_), .A2(new_n9178_), .B(new_n9212_), .ZN(new_n9213_));
  INV_X1     g08211(.I(new_n9172_), .ZN(new_n9214_));
  AOI21_X1   g08212(.A1(new_n9170_), .A2(new_n9214_), .B(new_n9176_), .ZN(new_n9215_));
  NAND2_X1   g08213(.A1(new_n9161_), .A2(new_n9215_), .ZN(new_n9216_));
  XOR2_X1    g08214(.A1(new_n9161_), .A2(new_n9178_), .Z(new_n9217_));
  AOI22_X1   g08215(.A1(new_n9217_), .A2(new_n9212_), .B1(new_n9213_), .B2(new_n9216_), .ZN(new_n9218_));
  AOI21_X1   g08216(.A1(new_n9207_), .A2(new_n9209_), .B(new_n9205_), .ZN(new_n9219_));
  NOR3_X1    g08217(.A1(new_n9203_), .A2(new_n9193_), .A3(new_n9141_), .ZN(new_n9220_));
  NOR3_X1    g08218(.A1(new_n9218_), .A2(new_n9220_), .A3(new_n9219_), .ZN(new_n9221_));
  OAI21_X1   g08219(.A1(new_n9221_), .A2(new_n9211_), .B(new_n9156_), .ZN(new_n9222_));
  INV_X1     g08220(.I(new_n9156_), .ZN(new_n9223_));
  OAI21_X1   g08221(.A1(new_n9219_), .A2(new_n9220_), .B(new_n9218_), .ZN(new_n9224_));
  NAND3_X1   g08222(.A1(new_n9180_), .A2(new_n9204_), .A3(new_n9210_), .ZN(new_n9225_));
  NAND3_X1   g08223(.A1(new_n9224_), .A2(new_n9225_), .A3(new_n9223_), .ZN(new_n9226_));
  NAND3_X1   g08224(.A1(new_n9222_), .A2(new_n9226_), .A3(new_n8981_), .ZN(new_n9227_));
  NAND3_X1   g08225(.A1(new_n8978_), .A2(new_n8979_), .A3(new_n8847_), .ZN(new_n9228_));
  OAI21_X1   g08226(.A1(new_n8976_), .A2(new_n8970_), .B(new_n8848_), .ZN(new_n9229_));
  NAND2_X1   g08227(.A1(new_n9228_), .A2(new_n9229_), .ZN(new_n9230_));
  AOI21_X1   g08228(.A1(new_n9224_), .A2(new_n9225_), .B(new_n9223_), .ZN(new_n9231_));
  NOR3_X1    g08229(.A1(new_n9221_), .A2(new_n9211_), .A3(new_n9156_), .ZN(new_n9232_));
  OAI21_X1   g08230(.A1(new_n9232_), .A2(new_n9231_), .B(new_n9230_), .ZN(new_n9233_));
  NAND2_X1   g08231(.A1(new_n9233_), .A2(new_n9227_), .ZN(new_n9234_));
  INV_X1     g08232(.I(\A[939] ), .ZN(new_n9235_));
  NOR2_X1    g08233(.A1(new_n9235_), .A2(\A[938] ), .ZN(new_n9236_));
  INV_X1     g08234(.I(\A[938] ), .ZN(new_n9237_));
  NOR2_X1    g08235(.A1(new_n9237_), .A2(\A[939] ), .ZN(new_n9238_));
  OAI21_X1   g08236(.A1(new_n9236_), .A2(new_n9238_), .B(\A[937] ), .ZN(new_n9239_));
  INV_X1     g08237(.I(\A[937] ), .ZN(new_n9240_));
  NAND2_X1   g08238(.A1(\A[938] ), .A2(\A[939] ), .ZN(new_n9241_));
  INV_X1     g08239(.I(new_n9241_), .ZN(new_n9242_));
  NOR2_X1    g08240(.A1(\A[938] ), .A2(\A[939] ), .ZN(new_n9243_));
  OAI21_X1   g08241(.A1(new_n9242_), .A2(new_n9243_), .B(new_n9240_), .ZN(new_n9244_));
  NAND2_X1   g08242(.A1(new_n9239_), .A2(new_n9244_), .ZN(new_n9245_));
  INV_X1     g08243(.I(\A[940] ), .ZN(new_n9246_));
  INV_X1     g08244(.I(\A[941] ), .ZN(new_n9247_));
  NAND2_X1   g08245(.A1(new_n9247_), .A2(\A[942] ), .ZN(new_n9248_));
  INV_X1     g08246(.I(\A[942] ), .ZN(new_n9249_));
  NAND2_X1   g08247(.A1(new_n9249_), .A2(\A[941] ), .ZN(new_n9250_));
  AOI21_X1   g08248(.A1(new_n9248_), .A2(new_n9250_), .B(new_n9246_), .ZN(new_n9251_));
  NAND2_X1   g08249(.A1(\A[941] ), .A2(\A[942] ), .ZN(new_n9252_));
  NOR2_X1    g08250(.A1(\A[941] ), .A2(\A[942] ), .ZN(new_n9253_));
  INV_X1     g08251(.I(new_n9253_), .ZN(new_n9254_));
  AOI21_X1   g08252(.A1(new_n9254_), .A2(new_n9252_), .B(\A[940] ), .ZN(new_n9255_));
  NOR2_X1    g08253(.A1(new_n9255_), .A2(new_n9251_), .ZN(new_n9256_));
  NOR2_X1    g08254(.A1(new_n9256_), .A2(new_n9245_), .ZN(new_n9257_));
  NAND2_X1   g08255(.A1(new_n9237_), .A2(\A[939] ), .ZN(new_n9258_));
  NAND2_X1   g08256(.A1(new_n9235_), .A2(\A[938] ), .ZN(new_n9259_));
  AOI21_X1   g08257(.A1(new_n9258_), .A2(new_n9259_), .B(new_n9240_), .ZN(new_n9260_));
  INV_X1     g08258(.I(new_n9243_), .ZN(new_n9261_));
  AOI21_X1   g08259(.A1(new_n9261_), .A2(new_n9241_), .B(\A[937] ), .ZN(new_n9262_));
  NOR2_X1    g08260(.A1(new_n9262_), .A2(new_n9260_), .ZN(new_n9263_));
  NOR2_X1    g08261(.A1(new_n9249_), .A2(\A[941] ), .ZN(new_n9264_));
  NOR2_X1    g08262(.A1(new_n9247_), .A2(\A[942] ), .ZN(new_n9265_));
  OAI21_X1   g08263(.A1(new_n9264_), .A2(new_n9265_), .B(\A[940] ), .ZN(new_n9266_));
  INV_X1     g08264(.I(new_n9252_), .ZN(new_n9267_));
  OAI21_X1   g08265(.A1(new_n9267_), .A2(new_n9253_), .B(new_n9246_), .ZN(new_n9268_));
  NAND2_X1   g08266(.A1(new_n9266_), .A2(new_n9268_), .ZN(new_n9269_));
  NOR2_X1    g08267(.A1(new_n9263_), .A2(new_n9269_), .ZN(new_n9270_));
  NOR2_X1    g08268(.A1(new_n9257_), .A2(new_n9270_), .ZN(new_n9271_));
  INV_X1     g08269(.I(\A[933] ), .ZN(new_n9272_));
  NOR2_X1    g08270(.A1(new_n9272_), .A2(\A[932] ), .ZN(new_n9273_));
  INV_X1     g08271(.I(\A[932] ), .ZN(new_n9274_));
  NOR2_X1    g08272(.A1(new_n9274_), .A2(\A[933] ), .ZN(new_n9275_));
  OAI21_X1   g08273(.A1(new_n9273_), .A2(new_n9275_), .B(\A[931] ), .ZN(new_n9276_));
  INV_X1     g08274(.I(\A[931] ), .ZN(new_n9277_));
  NAND2_X1   g08275(.A1(\A[932] ), .A2(\A[933] ), .ZN(new_n9278_));
  INV_X1     g08276(.I(new_n9278_), .ZN(new_n9279_));
  NOR2_X1    g08277(.A1(\A[932] ), .A2(\A[933] ), .ZN(new_n9280_));
  OAI21_X1   g08278(.A1(new_n9279_), .A2(new_n9280_), .B(new_n9277_), .ZN(new_n9281_));
  INV_X1     g08279(.I(\A[936] ), .ZN(new_n9282_));
  NOR2_X1    g08280(.A1(new_n9282_), .A2(\A[935] ), .ZN(new_n9283_));
  INV_X1     g08281(.I(\A[935] ), .ZN(new_n9284_));
  NOR2_X1    g08282(.A1(new_n9284_), .A2(\A[936] ), .ZN(new_n9285_));
  OAI21_X1   g08283(.A1(new_n9283_), .A2(new_n9285_), .B(\A[934] ), .ZN(new_n9286_));
  INV_X1     g08284(.I(\A[934] ), .ZN(new_n9287_));
  NAND2_X1   g08285(.A1(\A[935] ), .A2(\A[936] ), .ZN(new_n9288_));
  INV_X1     g08286(.I(new_n9288_), .ZN(new_n9289_));
  NOR2_X1    g08287(.A1(\A[935] ), .A2(\A[936] ), .ZN(new_n9290_));
  OAI21_X1   g08288(.A1(new_n9289_), .A2(new_n9290_), .B(new_n9287_), .ZN(new_n9291_));
  NAND4_X1   g08289(.A1(new_n9276_), .A2(new_n9281_), .A3(new_n9286_), .A4(new_n9291_), .ZN(new_n9292_));
  NAND2_X1   g08290(.A1(new_n9274_), .A2(\A[933] ), .ZN(new_n9293_));
  NAND2_X1   g08291(.A1(new_n9272_), .A2(\A[932] ), .ZN(new_n9294_));
  AOI21_X1   g08292(.A1(new_n9293_), .A2(new_n9294_), .B(new_n9277_), .ZN(new_n9295_));
  INV_X1     g08293(.I(new_n9280_), .ZN(new_n9296_));
  AOI21_X1   g08294(.A1(new_n9296_), .A2(new_n9278_), .B(\A[931] ), .ZN(new_n9297_));
  NAND2_X1   g08295(.A1(new_n9284_), .A2(\A[936] ), .ZN(new_n9298_));
  NAND2_X1   g08296(.A1(new_n9282_), .A2(\A[935] ), .ZN(new_n9299_));
  AOI21_X1   g08297(.A1(new_n9298_), .A2(new_n9299_), .B(new_n9287_), .ZN(new_n9300_));
  INV_X1     g08298(.I(new_n9290_), .ZN(new_n9301_));
  AOI21_X1   g08299(.A1(new_n9301_), .A2(new_n9288_), .B(\A[934] ), .ZN(new_n9302_));
  OAI22_X1   g08300(.A1(new_n9295_), .A2(new_n9297_), .B1(new_n9302_), .B2(new_n9300_), .ZN(new_n9303_));
  NAND2_X1   g08301(.A1(new_n9303_), .A2(new_n9292_), .ZN(new_n9304_));
  AOI21_X1   g08302(.A1(\A[941] ), .A2(\A[942] ), .B(\A[940] ), .ZN(new_n9305_));
  NOR2_X1    g08303(.A1(new_n9305_), .A2(new_n9253_), .ZN(new_n9306_));
  INV_X1     g08304(.I(new_n9306_), .ZN(new_n9307_));
  NOR4_X1    g08305(.A1(new_n9260_), .A2(new_n9262_), .A3(new_n9255_), .A4(new_n9251_), .ZN(new_n9308_));
  AOI21_X1   g08306(.A1(\A[938] ), .A2(\A[939] ), .B(\A[937] ), .ZN(new_n9309_));
  NOR2_X1    g08307(.A1(new_n9309_), .A2(new_n9243_), .ZN(new_n9310_));
  NAND2_X1   g08308(.A1(new_n9308_), .A2(new_n9310_), .ZN(new_n9311_));
  OAI21_X1   g08309(.A1(new_n9307_), .A2(new_n9311_), .B(new_n9304_), .ZN(new_n9312_));
  NAND2_X1   g08310(.A1(new_n9263_), .A2(new_n9269_), .ZN(new_n9313_));
  NAND2_X1   g08311(.A1(new_n9256_), .A2(new_n9245_), .ZN(new_n9314_));
  NOR4_X1    g08312(.A1(new_n9295_), .A2(new_n9297_), .A3(new_n9302_), .A4(new_n9300_), .ZN(new_n9315_));
  AOI21_X1   g08313(.A1(new_n9287_), .A2(new_n9288_), .B(new_n9290_), .ZN(new_n9316_));
  AOI21_X1   g08314(.A1(new_n9277_), .A2(new_n9278_), .B(new_n9280_), .ZN(new_n9317_));
  NAND3_X1   g08315(.A1(new_n9315_), .A2(new_n9316_), .A3(new_n9317_), .ZN(new_n9318_));
  NAND3_X1   g08316(.A1(new_n9318_), .A2(new_n9313_), .A3(new_n9314_), .ZN(new_n9319_));
  OAI22_X1   g08317(.A1(new_n9312_), .A2(new_n9271_), .B1(new_n9319_), .B2(new_n9304_), .ZN(new_n9320_));
  INV_X1     g08318(.I(\A[921] ), .ZN(new_n9321_));
  NOR2_X1    g08319(.A1(new_n9321_), .A2(\A[920] ), .ZN(new_n9322_));
  INV_X1     g08320(.I(\A[920] ), .ZN(new_n9323_));
  NOR2_X1    g08321(.A1(new_n9323_), .A2(\A[921] ), .ZN(new_n9324_));
  OAI21_X1   g08322(.A1(new_n9322_), .A2(new_n9324_), .B(\A[919] ), .ZN(new_n9325_));
  INV_X1     g08323(.I(\A[919] ), .ZN(new_n9326_));
  NAND2_X1   g08324(.A1(\A[920] ), .A2(\A[921] ), .ZN(new_n9327_));
  INV_X1     g08325(.I(new_n9327_), .ZN(new_n9328_));
  NOR2_X1    g08326(.A1(\A[920] ), .A2(\A[921] ), .ZN(new_n9329_));
  OAI21_X1   g08327(.A1(new_n9328_), .A2(new_n9329_), .B(new_n9326_), .ZN(new_n9330_));
  INV_X1     g08328(.I(\A[924] ), .ZN(new_n9331_));
  NOR2_X1    g08329(.A1(new_n9331_), .A2(\A[923] ), .ZN(new_n9332_));
  INV_X1     g08330(.I(\A[923] ), .ZN(new_n9333_));
  NOR2_X1    g08331(.A1(new_n9333_), .A2(\A[924] ), .ZN(new_n9334_));
  OAI21_X1   g08332(.A1(new_n9332_), .A2(new_n9334_), .B(\A[922] ), .ZN(new_n9335_));
  INV_X1     g08333(.I(\A[922] ), .ZN(new_n9336_));
  NAND2_X1   g08334(.A1(\A[923] ), .A2(\A[924] ), .ZN(new_n9337_));
  INV_X1     g08335(.I(new_n9337_), .ZN(new_n9338_));
  NOR2_X1    g08336(.A1(\A[923] ), .A2(\A[924] ), .ZN(new_n9339_));
  OAI21_X1   g08337(.A1(new_n9338_), .A2(new_n9339_), .B(new_n9336_), .ZN(new_n9340_));
  NAND4_X1   g08338(.A1(new_n9325_), .A2(new_n9330_), .A3(new_n9335_), .A4(new_n9340_), .ZN(new_n9341_));
  NAND2_X1   g08339(.A1(new_n9323_), .A2(\A[921] ), .ZN(new_n9342_));
  NAND2_X1   g08340(.A1(new_n9321_), .A2(\A[920] ), .ZN(new_n9343_));
  AOI21_X1   g08341(.A1(new_n9342_), .A2(new_n9343_), .B(new_n9326_), .ZN(new_n9344_));
  INV_X1     g08342(.I(new_n9329_), .ZN(new_n9345_));
  AOI21_X1   g08343(.A1(new_n9345_), .A2(new_n9327_), .B(\A[919] ), .ZN(new_n9346_));
  NAND2_X1   g08344(.A1(new_n9333_), .A2(\A[924] ), .ZN(new_n9347_));
  NAND2_X1   g08345(.A1(new_n9331_), .A2(\A[923] ), .ZN(new_n9348_));
  AOI21_X1   g08346(.A1(new_n9347_), .A2(new_n9348_), .B(new_n9336_), .ZN(new_n9349_));
  INV_X1     g08347(.I(new_n9339_), .ZN(new_n9350_));
  AOI21_X1   g08348(.A1(new_n9350_), .A2(new_n9337_), .B(\A[922] ), .ZN(new_n9351_));
  OAI22_X1   g08349(.A1(new_n9344_), .A2(new_n9346_), .B1(new_n9351_), .B2(new_n9349_), .ZN(new_n9352_));
  NAND2_X1   g08350(.A1(new_n9352_), .A2(new_n9341_), .ZN(new_n9353_));
  INV_X1     g08351(.I(\A[925] ), .ZN(new_n9354_));
  INV_X1     g08352(.I(\A[926] ), .ZN(new_n9355_));
  NAND2_X1   g08353(.A1(new_n9355_), .A2(\A[927] ), .ZN(new_n9356_));
  INV_X1     g08354(.I(\A[927] ), .ZN(new_n9357_));
  NAND2_X1   g08355(.A1(new_n9357_), .A2(\A[926] ), .ZN(new_n9358_));
  AOI21_X1   g08356(.A1(new_n9356_), .A2(new_n9358_), .B(new_n9354_), .ZN(new_n9359_));
  NAND2_X1   g08357(.A1(\A[926] ), .A2(\A[927] ), .ZN(new_n9360_));
  NOR2_X1    g08358(.A1(\A[926] ), .A2(\A[927] ), .ZN(new_n9361_));
  INV_X1     g08359(.I(new_n9361_), .ZN(new_n9362_));
  AOI21_X1   g08360(.A1(new_n9362_), .A2(new_n9360_), .B(\A[925] ), .ZN(new_n9363_));
  NOR2_X1    g08361(.A1(new_n9363_), .A2(new_n9359_), .ZN(new_n9364_));
  INV_X1     g08362(.I(\A[930] ), .ZN(new_n9365_));
  NOR2_X1    g08363(.A1(new_n9365_), .A2(\A[929] ), .ZN(new_n9366_));
  INV_X1     g08364(.I(\A[929] ), .ZN(new_n9367_));
  NOR2_X1    g08365(.A1(new_n9367_), .A2(\A[930] ), .ZN(new_n9368_));
  OAI21_X1   g08366(.A1(new_n9366_), .A2(new_n9368_), .B(\A[928] ), .ZN(new_n9369_));
  INV_X1     g08367(.I(\A[928] ), .ZN(new_n9370_));
  NAND2_X1   g08368(.A1(\A[929] ), .A2(\A[930] ), .ZN(new_n9371_));
  INV_X1     g08369(.I(new_n9371_), .ZN(new_n9372_));
  NOR2_X1    g08370(.A1(\A[929] ), .A2(\A[930] ), .ZN(new_n9373_));
  OAI21_X1   g08371(.A1(new_n9372_), .A2(new_n9373_), .B(new_n9370_), .ZN(new_n9374_));
  NAND2_X1   g08372(.A1(new_n9369_), .A2(new_n9374_), .ZN(new_n9375_));
  NAND2_X1   g08373(.A1(new_n9364_), .A2(new_n9375_), .ZN(new_n9376_));
  NOR2_X1    g08374(.A1(new_n9357_), .A2(\A[926] ), .ZN(new_n9377_));
  NOR2_X1    g08375(.A1(new_n9355_), .A2(\A[927] ), .ZN(new_n9378_));
  OAI21_X1   g08376(.A1(new_n9377_), .A2(new_n9378_), .B(\A[925] ), .ZN(new_n9379_));
  INV_X1     g08377(.I(new_n9360_), .ZN(new_n9380_));
  OAI21_X1   g08378(.A1(new_n9380_), .A2(new_n9361_), .B(new_n9354_), .ZN(new_n9381_));
  NAND2_X1   g08379(.A1(new_n9379_), .A2(new_n9381_), .ZN(new_n9382_));
  NAND2_X1   g08380(.A1(new_n9367_), .A2(\A[930] ), .ZN(new_n9383_));
  NAND2_X1   g08381(.A1(new_n9365_), .A2(\A[929] ), .ZN(new_n9384_));
  AOI21_X1   g08382(.A1(new_n9383_), .A2(new_n9384_), .B(new_n9370_), .ZN(new_n9385_));
  INV_X1     g08383(.I(new_n9373_), .ZN(new_n9386_));
  AOI21_X1   g08384(.A1(new_n9386_), .A2(new_n9371_), .B(\A[928] ), .ZN(new_n9387_));
  NOR2_X1    g08385(.A1(new_n9387_), .A2(new_n9385_), .ZN(new_n9388_));
  NAND2_X1   g08386(.A1(new_n9388_), .A2(new_n9382_), .ZN(new_n9389_));
  AOI21_X1   g08387(.A1(new_n9376_), .A2(new_n9389_), .B(new_n9353_), .ZN(new_n9390_));
  NAND2_X1   g08388(.A1(new_n9376_), .A2(new_n9389_), .ZN(new_n9391_));
  NOR4_X1    g08389(.A1(new_n9344_), .A2(new_n9346_), .A3(new_n9351_), .A4(new_n9349_), .ZN(new_n9392_));
  AOI22_X1   g08390(.A1(new_n9325_), .A2(new_n9330_), .B1(new_n9335_), .B2(new_n9340_), .ZN(new_n9393_));
  AOI21_X1   g08391(.A1(\A[923] ), .A2(\A[924] ), .B(\A[922] ), .ZN(new_n9394_));
  NOR2_X1    g08392(.A1(new_n9394_), .A2(new_n9339_), .ZN(new_n9395_));
  AOI21_X1   g08393(.A1(\A[920] ), .A2(\A[921] ), .B(\A[919] ), .ZN(new_n9396_));
  NOR2_X1    g08394(.A1(new_n9396_), .A2(new_n9329_), .ZN(new_n9397_));
  NOR2_X1    g08395(.A1(new_n9393_), .A2(new_n9392_), .ZN(new_n9398_));
  NOR2_X1    g08396(.A1(new_n9391_), .A2(new_n9398_), .ZN(new_n9399_));
  NOR2_X1    g08397(.A1(new_n9399_), .A2(new_n9390_), .ZN(new_n9400_));
  NAND2_X1   g08398(.A1(new_n9320_), .A2(new_n9400_), .ZN(new_n9401_));
  NAND2_X1   g08399(.A1(new_n9313_), .A2(new_n9314_), .ZN(new_n9402_));
  AOI22_X1   g08400(.A1(new_n9276_), .A2(new_n9281_), .B1(new_n9286_), .B2(new_n9291_), .ZN(new_n9403_));
  NOR2_X1    g08401(.A1(new_n9403_), .A2(new_n9315_), .ZN(new_n9404_));
  NAND4_X1   g08402(.A1(new_n9239_), .A2(new_n9244_), .A3(new_n9266_), .A4(new_n9268_), .ZN(new_n9405_));
  INV_X1     g08403(.I(new_n9310_), .ZN(new_n9406_));
  NOR2_X1    g08404(.A1(new_n9405_), .A2(new_n9406_), .ZN(new_n9407_));
  AOI21_X1   g08405(.A1(new_n9306_), .A2(new_n9407_), .B(new_n9404_), .ZN(new_n9408_));
  INV_X1     g08406(.I(new_n9316_), .ZN(new_n9409_));
  INV_X1     g08407(.I(new_n9317_), .ZN(new_n9410_));
  NOR3_X1    g08408(.A1(new_n9292_), .A2(new_n9409_), .A3(new_n9410_), .ZN(new_n9411_));
  NOR2_X1    g08409(.A1(new_n9402_), .A2(new_n9411_), .ZN(new_n9412_));
  AOI22_X1   g08410(.A1(new_n9404_), .A2(new_n9412_), .B1(new_n9408_), .B2(new_n9402_), .ZN(new_n9413_));
  NOR2_X1    g08411(.A1(new_n9393_), .A2(new_n9392_), .ZN(new_n9414_));
  NAND2_X1   g08412(.A1(new_n9391_), .A2(new_n9414_), .ZN(new_n9415_));
  OAI21_X1   g08413(.A1(new_n9391_), .A2(new_n9398_), .B(new_n9415_), .ZN(new_n9416_));
  NAND2_X1   g08414(.A1(new_n9413_), .A2(new_n9416_), .ZN(new_n9417_));
  NAND2_X1   g08415(.A1(new_n9417_), .A2(new_n9401_), .ZN(new_n9418_));
  INV_X1     g08416(.I(\A[907] ), .ZN(new_n9419_));
  INV_X1     g08417(.I(\A[908] ), .ZN(new_n9420_));
  NAND2_X1   g08418(.A1(new_n9420_), .A2(\A[909] ), .ZN(new_n9421_));
  INV_X1     g08419(.I(\A[909] ), .ZN(new_n9422_));
  NAND2_X1   g08420(.A1(new_n9422_), .A2(\A[908] ), .ZN(new_n9423_));
  AOI21_X1   g08421(.A1(new_n9421_), .A2(new_n9423_), .B(new_n9419_), .ZN(new_n9424_));
  NAND2_X1   g08422(.A1(\A[908] ), .A2(\A[909] ), .ZN(new_n9425_));
  NOR2_X1    g08423(.A1(\A[908] ), .A2(\A[909] ), .ZN(new_n9426_));
  INV_X1     g08424(.I(new_n9426_), .ZN(new_n9427_));
  AOI21_X1   g08425(.A1(new_n9427_), .A2(new_n9425_), .B(\A[907] ), .ZN(new_n9428_));
  INV_X1     g08426(.I(\A[910] ), .ZN(new_n9429_));
  INV_X1     g08427(.I(\A[911] ), .ZN(new_n9430_));
  NAND2_X1   g08428(.A1(new_n9430_), .A2(\A[912] ), .ZN(new_n9431_));
  INV_X1     g08429(.I(\A[912] ), .ZN(new_n9432_));
  NAND2_X1   g08430(.A1(new_n9432_), .A2(\A[911] ), .ZN(new_n9433_));
  AOI21_X1   g08431(.A1(new_n9431_), .A2(new_n9433_), .B(new_n9429_), .ZN(new_n9434_));
  NAND2_X1   g08432(.A1(\A[911] ), .A2(\A[912] ), .ZN(new_n9435_));
  NAND2_X1   g08433(.A1(new_n9430_), .A2(new_n9432_), .ZN(new_n9436_));
  AOI21_X1   g08434(.A1(new_n9436_), .A2(new_n9435_), .B(\A[910] ), .ZN(new_n9437_));
  NOR4_X1    g08435(.A1(new_n9424_), .A2(new_n9428_), .A3(new_n9437_), .A4(new_n9434_), .ZN(new_n9438_));
  NOR2_X1    g08436(.A1(new_n9428_), .A2(new_n9424_), .ZN(new_n9439_));
  NOR2_X1    g08437(.A1(new_n9437_), .A2(new_n9434_), .ZN(new_n9440_));
  NOR2_X1    g08438(.A1(new_n9439_), .A2(new_n9440_), .ZN(new_n9441_));
  INV_X1     g08439(.I(\A[915] ), .ZN(new_n9442_));
  NOR2_X1    g08440(.A1(new_n9442_), .A2(\A[914] ), .ZN(new_n9443_));
  INV_X1     g08441(.I(\A[914] ), .ZN(new_n9444_));
  NOR2_X1    g08442(.A1(new_n9444_), .A2(\A[915] ), .ZN(new_n9445_));
  OAI21_X1   g08443(.A1(new_n9443_), .A2(new_n9445_), .B(\A[913] ), .ZN(new_n9446_));
  INV_X1     g08444(.I(\A[913] ), .ZN(new_n9447_));
  NAND2_X1   g08445(.A1(\A[914] ), .A2(\A[915] ), .ZN(new_n9448_));
  INV_X1     g08446(.I(new_n9448_), .ZN(new_n9449_));
  NOR2_X1    g08447(.A1(\A[914] ), .A2(\A[915] ), .ZN(new_n9450_));
  OAI21_X1   g08448(.A1(new_n9449_), .A2(new_n9450_), .B(new_n9447_), .ZN(new_n9451_));
  NAND2_X1   g08449(.A1(new_n9446_), .A2(new_n9451_), .ZN(new_n9452_));
  INV_X1     g08450(.I(\A[916] ), .ZN(new_n9453_));
  INV_X1     g08451(.I(\A[917] ), .ZN(new_n9454_));
  NAND2_X1   g08452(.A1(new_n9454_), .A2(\A[918] ), .ZN(new_n9455_));
  INV_X1     g08453(.I(\A[918] ), .ZN(new_n9456_));
  NAND2_X1   g08454(.A1(new_n9456_), .A2(\A[917] ), .ZN(new_n9457_));
  AOI21_X1   g08455(.A1(new_n9455_), .A2(new_n9457_), .B(new_n9453_), .ZN(new_n9458_));
  NAND2_X1   g08456(.A1(\A[917] ), .A2(\A[918] ), .ZN(new_n9459_));
  NOR2_X1    g08457(.A1(\A[917] ), .A2(\A[918] ), .ZN(new_n9460_));
  INV_X1     g08458(.I(new_n9460_), .ZN(new_n9461_));
  AOI21_X1   g08459(.A1(new_n9461_), .A2(new_n9459_), .B(\A[916] ), .ZN(new_n9462_));
  NOR2_X1    g08460(.A1(new_n9462_), .A2(new_n9458_), .ZN(new_n9463_));
  NOR2_X1    g08461(.A1(new_n9463_), .A2(new_n9452_), .ZN(new_n9464_));
  NAND2_X1   g08462(.A1(new_n9444_), .A2(\A[915] ), .ZN(new_n9465_));
  NAND2_X1   g08463(.A1(new_n9442_), .A2(\A[914] ), .ZN(new_n9466_));
  AOI21_X1   g08464(.A1(new_n9465_), .A2(new_n9466_), .B(new_n9447_), .ZN(new_n9467_));
  INV_X1     g08465(.I(new_n9450_), .ZN(new_n9468_));
  AOI21_X1   g08466(.A1(new_n9468_), .A2(new_n9448_), .B(\A[913] ), .ZN(new_n9469_));
  NOR2_X1    g08467(.A1(new_n9469_), .A2(new_n9467_), .ZN(new_n9470_));
  NOR2_X1    g08468(.A1(new_n9456_), .A2(\A[917] ), .ZN(new_n9471_));
  NOR2_X1    g08469(.A1(new_n9454_), .A2(\A[918] ), .ZN(new_n9472_));
  OAI21_X1   g08470(.A1(new_n9471_), .A2(new_n9472_), .B(\A[916] ), .ZN(new_n9473_));
  INV_X1     g08471(.I(new_n9459_), .ZN(new_n9474_));
  OAI21_X1   g08472(.A1(new_n9474_), .A2(new_n9460_), .B(new_n9453_), .ZN(new_n9475_));
  NAND2_X1   g08473(.A1(new_n9473_), .A2(new_n9475_), .ZN(new_n9476_));
  NOR2_X1    g08474(.A1(new_n9470_), .A2(new_n9476_), .ZN(new_n9477_));
  NOR2_X1    g08475(.A1(new_n9464_), .A2(new_n9477_), .ZN(new_n9478_));
  NOR3_X1    g08476(.A1(new_n9478_), .A2(new_n9438_), .A3(new_n9441_), .ZN(new_n9479_));
  NOR2_X1    g08477(.A1(new_n9441_), .A2(new_n9438_), .ZN(new_n9480_));
  NAND2_X1   g08478(.A1(new_n9470_), .A2(new_n9476_), .ZN(new_n9481_));
  NAND2_X1   g08479(.A1(new_n9463_), .A2(new_n9452_), .ZN(new_n9482_));
  NAND2_X1   g08480(.A1(new_n9481_), .A2(new_n9482_), .ZN(new_n9483_));
  NAND2_X1   g08481(.A1(new_n9435_), .A2(new_n9429_), .ZN(new_n9484_));
  NAND2_X1   g08482(.A1(new_n9484_), .A2(new_n9436_), .ZN(new_n9485_));
  INV_X1     g08483(.I(new_n9485_), .ZN(new_n9486_));
  AOI21_X1   g08484(.A1(new_n9419_), .A2(new_n9425_), .B(new_n9426_), .ZN(new_n9487_));
  NAND3_X1   g08485(.A1(new_n9438_), .A2(new_n9486_), .A3(new_n9487_), .ZN(new_n9488_));
  AOI21_X1   g08486(.A1(new_n9480_), .A2(new_n9488_), .B(new_n9483_), .ZN(new_n9489_));
  INV_X1     g08487(.I(\A[897] ), .ZN(new_n9490_));
  NOR2_X1    g08488(.A1(new_n9490_), .A2(\A[896] ), .ZN(new_n9491_));
  INV_X1     g08489(.I(\A[896] ), .ZN(new_n9492_));
  NOR2_X1    g08490(.A1(new_n9492_), .A2(\A[897] ), .ZN(new_n9493_));
  OAI21_X1   g08491(.A1(new_n9491_), .A2(new_n9493_), .B(\A[895] ), .ZN(new_n9494_));
  INV_X1     g08492(.I(\A[895] ), .ZN(new_n9495_));
  NAND2_X1   g08493(.A1(\A[896] ), .A2(\A[897] ), .ZN(new_n9496_));
  INV_X1     g08494(.I(new_n9496_), .ZN(new_n9497_));
  NOR2_X1    g08495(.A1(\A[896] ), .A2(\A[897] ), .ZN(new_n9498_));
  OAI21_X1   g08496(.A1(new_n9497_), .A2(new_n9498_), .B(new_n9495_), .ZN(new_n9499_));
  INV_X1     g08497(.I(\A[900] ), .ZN(new_n9500_));
  NOR2_X1    g08498(.A1(new_n9500_), .A2(\A[899] ), .ZN(new_n9501_));
  INV_X1     g08499(.I(\A[899] ), .ZN(new_n9502_));
  NOR2_X1    g08500(.A1(new_n9502_), .A2(\A[900] ), .ZN(new_n9503_));
  OAI21_X1   g08501(.A1(new_n9501_), .A2(new_n9503_), .B(\A[898] ), .ZN(new_n9504_));
  INV_X1     g08502(.I(\A[898] ), .ZN(new_n9505_));
  NAND2_X1   g08503(.A1(\A[899] ), .A2(\A[900] ), .ZN(new_n9506_));
  INV_X1     g08504(.I(new_n9506_), .ZN(new_n9507_));
  NOR2_X1    g08505(.A1(\A[899] ), .A2(\A[900] ), .ZN(new_n9508_));
  OAI21_X1   g08506(.A1(new_n9507_), .A2(new_n9508_), .B(new_n9505_), .ZN(new_n9509_));
  NAND4_X1   g08507(.A1(new_n9494_), .A2(new_n9499_), .A3(new_n9504_), .A4(new_n9509_), .ZN(new_n9510_));
  INV_X1     g08508(.I(new_n9491_), .ZN(new_n9511_));
  NAND2_X1   g08509(.A1(new_n9490_), .A2(\A[896] ), .ZN(new_n9512_));
  AOI21_X1   g08510(.A1(new_n9511_), .A2(new_n9512_), .B(new_n9495_), .ZN(new_n9513_));
  INV_X1     g08511(.I(new_n9498_), .ZN(new_n9514_));
  AOI21_X1   g08512(.A1(new_n9514_), .A2(new_n9496_), .B(\A[895] ), .ZN(new_n9515_));
  NAND2_X1   g08513(.A1(new_n9502_), .A2(\A[900] ), .ZN(new_n9516_));
  NAND2_X1   g08514(.A1(new_n9500_), .A2(\A[899] ), .ZN(new_n9517_));
  AOI21_X1   g08515(.A1(new_n9516_), .A2(new_n9517_), .B(new_n9505_), .ZN(new_n9518_));
  INV_X1     g08516(.I(new_n9508_), .ZN(new_n9519_));
  AOI21_X1   g08517(.A1(new_n9519_), .A2(new_n9506_), .B(\A[898] ), .ZN(new_n9520_));
  OAI22_X1   g08518(.A1(new_n9513_), .A2(new_n9515_), .B1(new_n9520_), .B2(new_n9518_), .ZN(new_n9521_));
  NAND2_X1   g08519(.A1(new_n9521_), .A2(new_n9510_), .ZN(new_n9522_));
  INV_X1     g08520(.I(\A[903] ), .ZN(new_n9523_));
  NOR2_X1    g08521(.A1(new_n9523_), .A2(\A[902] ), .ZN(new_n9524_));
  INV_X1     g08522(.I(\A[902] ), .ZN(new_n9525_));
  NOR2_X1    g08523(.A1(new_n9525_), .A2(\A[903] ), .ZN(new_n9526_));
  OAI21_X1   g08524(.A1(new_n9524_), .A2(new_n9526_), .B(\A[901] ), .ZN(new_n9527_));
  INV_X1     g08525(.I(\A[901] ), .ZN(new_n9528_));
  NAND2_X1   g08526(.A1(\A[902] ), .A2(\A[903] ), .ZN(new_n9529_));
  INV_X1     g08527(.I(new_n9529_), .ZN(new_n9530_));
  NOR2_X1    g08528(.A1(\A[902] ), .A2(\A[903] ), .ZN(new_n9531_));
  OAI21_X1   g08529(.A1(new_n9530_), .A2(new_n9531_), .B(new_n9528_), .ZN(new_n9532_));
  NAND2_X1   g08530(.A1(new_n9527_), .A2(new_n9532_), .ZN(new_n9533_));
  INV_X1     g08531(.I(\A[904] ), .ZN(new_n9534_));
  INV_X1     g08532(.I(\A[905] ), .ZN(new_n9535_));
  NAND2_X1   g08533(.A1(new_n9535_), .A2(\A[906] ), .ZN(new_n9536_));
  INV_X1     g08534(.I(\A[906] ), .ZN(new_n9537_));
  NAND2_X1   g08535(.A1(new_n9537_), .A2(\A[905] ), .ZN(new_n9538_));
  AOI21_X1   g08536(.A1(new_n9536_), .A2(new_n9538_), .B(new_n9534_), .ZN(new_n9539_));
  NAND2_X1   g08537(.A1(\A[905] ), .A2(\A[906] ), .ZN(new_n9540_));
  NOR2_X1    g08538(.A1(\A[905] ), .A2(\A[906] ), .ZN(new_n9541_));
  INV_X1     g08539(.I(new_n9541_), .ZN(new_n9542_));
  AOI21_X1   g08540(.A1(new_n9542_), .A2(new_n9540_), .B(\A[904] ), .ZN(new_n9543_));
  NOR2_X1    g08541(.A1(new_n9543_), .A2(new_n9539_), .ZN(new_n9544_));
  NOR2_X1    g08542(.A1(new_n9544_), .A2(new_n9533_), .ZN(new_n9545_));
  NAND2_X1   g08543(.A1(new_n9525_), .A2(\A[903] ), .ZN(new_n9546_));
  NAND2_X1   g08544(.A1(new_n9523_), .A2(\A[902] ), .ZN(new_n9547_));
  AOI21_X1   g08545(.A1(new_n9546_), .A2(new_n9547_), .B(new_n9528_), .ZN(new_n9548_));
  INV_X1     g08546(.I(new_n9531_), .ZN(new_n9549_));
  AOI21_X1   g08547(.A1(new_n9549_), .A2(new_n9529_), .B(\A[901] ), .ZN(new_n9550_));
  NOR2_X1    g08548(.A1(new_n9550_), .A2(new_n9548_), .ZN(new_n9551_));
  NOR2_X1    g08549(.A1(new_n9537_), .A2(\A[905] ), .ZN(new_n9552_));
  NOR2_X1    g08550(.A1(new_n9535_), .A2(\A[906] ), .ZN(new_n9553_));
  OAI21_X1   g08551(.A1(new_n9552_), .A2(new_n9553_), .B(\A[904] ), .ZN(new_n9554_));
  INV_X1     g08552(.I(new_n9540_), .ZN(new_n9555_));
  OAI21_X1   g08553(.A1(new_n9555_), .A2(new_n9541_), .B(new_n9534_), .ZN(new_n9556_));
  NAND2_X1   g08554(.A1(new_n9554_), .A2(new_n9556_), .ZN(new_n9557_));
  NOR2_X1    g08555(.A1(new_n9551_), .A2(new_n9557_), .ZN(new_n9558_));
  NOR2_X1    g08556(.A1(new_n9545_), .A2(new_n9558_), .ZN(new_n9559_));
  NOR2_X1    g08557(.A1(new_n9559_), .A2(new_n9522_), .ZN(new_n9560_));
  NAND2_X1   g08558(.A1(new_n9551_), .A2(new_n9557_), .ZN(new_n9561_));
  NAND2_X1   g08559(.A1(new_n9544_), .A2(new_n9533_), .ZN(new_n9562_));
  NAND2_X1   g08560(.A1(new_n9561_), .A2(new_n9562_), .ZN(new_n9563_));
  AOI21_X1   g08561(.A1(new_n9505_), .A2(new_n9506_), .B(new_n9508_), .ZN(new_n9564_));
  AOI21_X1   g08562(.A1(new_n9495_), .A2(new_n9496_), .B(new_n9498_), .ZN(new_n9565_));
  AOI21_X1   g08563(.A1(new_n9510_), .A2(new_n9521_), .B(new_n9563_), .ZN(new_n9566_));
  NOR4_X1    g08564(.A1(new_n9489_), .A2(new_n9566_), .A3(new_n9479_), .A4(new_n9560_), .ZN(new_n9567_));
  NOR2_X1    g08565(.A1(new_n9489_), .A2(new_n9479_), .ZN(new_n9568_));
  NOR2_X1    g08566(.A1(new_n9566_), .A2(new_n9560_), .ZN(new_n9569_));
  NOR2_X1    g08567(.A1(new_n9568_), .A2(new_n9569_), .ZN(new_n9570_));
  NOR3_X1    g08568(.A1(new_n9418_), .A2(new_n9567_), .A3(new_n9570_), .ZN(new_n9571_));
  NOR2_X1    g08569(.A1(new_n9413_), .A2(new_n9416_), .ZN(new_n9572_));
  NOR2_X1    g08570(.A1(new_n9320_), .A2(new_n9400_), .ZN(new_n9573_));
  NOR2_X1    g08571(.A1(new_n9572_), .A2(new_n9573_), .ZN(new_n9574_));
  NOR2_X1    g08572(.A1(new_n9570_), .A2(new_n9567_), .ZN(new_n9575_));
  NOR2_X1    g08573(.A1(new_n9575_), .A2(new_n9574_), .ZN(new_n9576_));
  NOR2_X1    g08574(.A1(new_n9576_), .A2(new_n9571_), .ZN(new_n9577_));
  NOR2_X1    g08575(.A1(new_n9154_), .A2(new_n9141_), .ZN(new_n9578_));
  NOR2_X1    g08576(.A1(new_n8971_), .A2(new_n9155_), .ZN(new_n9579_));
  NOR2_X1    g08577(.A1(new_n9579_), .A2(new_n9578_), .ZN(new_n9580_));
  NOR2_X1    g08578(.A1(new_n9580_), .A2(new_n9156_), .ZN(new_n9581_));
  NAND2_X1   g08579(.A1(new_n9581_), .A2(new_n9577_), .ZN(new_n9582_));
  NAND2_X1   g08580(.A1(new_n9575_), .A2(new_n9574_), .ZN(new_n9583_));
  OAI22_X1   g08581(.A1(new_n9329_), .A2(new_n9396_), .B1(new_n9394_), .B2(new_n9339_), .ZN(new_n9584_));
  NAND2_X1   g08582(.A1(new_n9395_), .A2(new_n9397_), .ZN(new_n9585_));
  NAND2_X1   g08583(.A1(new_n9585_), .A2(new_n9584_), .ZN(new_n9586_));
  XOR2_X1    g08584(.A1(new_n9392_), .A2(new_n9586_), .Z(new_n9587_));
  NAND3_X1   g08585(.A1(new_n9392_), .A2(new_n9395_), .A3(new_n9397_), .ZN(new_n9588_));
  NAND3_X1   g08586(.A1(new_n9391_), .A2(new_n9414_), .A3(new_n9588_), .ZN(new_n9589_));
  AOI21_X1   g08587(.A1(new_n9370_), .A2(new_n9371_), .B(new_n9373_), .ZN(new_n9590_));
  AOI21_X1   g08588(.A1(\A[926] ), .A2(\A[927] ), .B(\A[925] ), .ZN(new_n9591_));
  NOR2_X1    g08589(.A1(new_n9591_), .A2(new_n9361_), .ZN(new_n9592_));
  XOR2_X1    g08590(.A1(new_n9590_), .A2(new_n9592_), .Z(new_n9593_));
  NOR3_X1    g08591(.A1(new_n9593_), .A2(new_n9382_), .A3(new_n9375_), .ZN(new_n9594_));
  NOR2_X1    g08592(.A1(new_n9382_), .A2(new_n9375_), .ZN(new_n9595_));
  XNOR2_X1   g08593(.A1(new_n9590_), .A2(new_n9592_), .ZN(new_n9596_));
  NOR2_X1    g08594(.A1(new_n9595_), .A2(new_n9596_), .ZN(new_n9597_));
  NOR2_X1    g08595(.A1(new_n9597_), .A2(new_n9594_), .ZN(new_n9598_));
  AOI21_X1   g08596(.A1(new_n9589_), .A2(new_n9598_), .B(new_n9587_), .ZN(new_n9599_));
  NOR2_X1    g08597(.A1(new_n9388_), .A2(new_n9382_), .ZN(new_n9600_));
  NOR2_X1    g08598(.A1(new_n9364_), .A2(new_n9375_), .ZN(new_n9601_));
  AND2_X2    g08599(.A1(new_n9590_), .A2(new_n9592_), .Z(new_n9602_));
  OAI21_X1   g08600(.A1(new_n9600_), .A2(new_n9601_), .B(new_n9602_), .ZN(new_n9603_));
  NAND4_X1   g08601(.A1(new_n9390_), .A2(new_n9588_), .A3(new_n9593_), .A4(new_n9603_), .ZN(new_n9604_));
  NAND2_X1   g08602(.A1(new_n9595_), .A2(new_n9596_), .ZN(new_n9605_));
  OAI21_X1   g08603(.A1(new_n9382_), .A2(new_n9375_), .B(new_n9593_), .ZN(new_n9606_));
  NAND2_X1   g08604(.A1(new_n9606_), .A2(new_n9605_), .ZN(new_n9607_));
  XOR2_X1    g08605(.A1(new_n9589_), .A2(new_n9607_), .Z(new_n9608_));
  AOI22_X1   g08606(.A1(new_n9608_), .A2(new_n9587_), .B1(new_n9599_), .B2(new_n9604_), .ZN(new_n9609_));
  NOR2_X1    g08607(.A1(new_n9316_), .A2(new_n9317_), .ZN(new_n9610_));
  NOR2_X1    g08608(.A1(new_n9409_), .A2(new_n9410_), .ZN(new_n9611_));
  NOR2_X1    g08609(.A1(new_n9611_), .A2(new_n9610_), .ZN(new_n9612_));
  XOR2_X1    g08610(.A1(new_n9612_), .A2(new_n9292_), .Z(new_n9613_));
  INV_X1     g08611(.I(new_n9613_), .ZN(new_n9614_));
  NOR3_X1    g08612(.A1(new_n9310_), .A2(new_n9253_), .A3(new_n9305_), .ZN(new_n9615_));
  NOR3_X1    g08613(.A1(new_n9306_), .A2(new_n9243_), .A3(new_n9309_), .ZN(new_n9616_));
  OR2_X2     g08614(.A1(new_n9615_), .A2(new_n9616_), .Z(new_n9617_));
  NOR2_X1    g08615(.A1(new_n9617_), .A2(new_n9308_), .ZN(new_n9618_));
  NOR2_X1    g08616(.A1(new_n9615_), .A2(new_n9616_), .ZN(new_n9619_));
  NOR2_X1    g08617(.A1(new_n9405_), .A2(new_n9619_), .ZN(new_n9620_));
  NOR2_X1    g08618(.A1(new_n9618_), .A2(new_n9620_), .ZN(new_n9621_));
  NAND3_X1   g08619(.A1(new_n9402_), .A2(new_n9306_), .A3(new_n9310_), .ZN(new_n9622_));
  AOI21_X1   g08620(.A1(new_n9313_), .A2(new_n9314_), .B(new_n9304_), .ZN(new_n9623_));
  AOI21_X1   g08621(.A1(new_n9622_), .A2(new_n9621_), .B(new_n9623_), .ZN(new_n9624_));
  NOR3_X1    g08622(.A1(new_n9271_), .A2(new_n9307_), .A3(new_n9406_), .ZN(new_n9625_));
  AOI21_X1   g08623(.A1(new_n9313_), .A2(new_n9314_), .B(new_n9619_), .ZN(new_n9626_));
  INV_X1     g08624(.I(new_n9626_), .ZN(new_n9627_));
  NOR3_X1    g08625(.A1(new_n9625_), .A2(new_n9627_), .A3(new_n9304_), .ZN(new_n9628_));
  OAI21_X1   g08626(.A1(new_n9628_), .A2(new_n9624_), .B(new_n9614_), .ZN(new_n9629_));
  XOR2_X1    g08627(.A1(new_n9308_), .A2(new_n9619_), .Z(new_n9630_));
  NAND2_X1   g08628(.A1(new_n9402_), .A2(new_n9404_), .ZN(new_n9631_));
  OAI21_X1   g08629(.A1(new_n9625_), .A2(new_n9630_), .B(new_n9631_), .ZN(new_n9632_));
  NAND3_X1   g08630(.A1(new_n9622_), .A2(new_n9623_), .A3(new_n9621_), .ZN(new_n9633_));
  NAND3_X1   g08631(.A1(new_n9632_), .A2(new_n9633_), .A3(new_n9613_), .ZN(new_n9634_));
  AOI21_X1   g08632(.A1(new_n9629_), .A2(new_n9634_), .B(new_n9401_), .ZN(new_n9635_));
  NAND3_X1   g08633(.A1(new_n9622_), .A2(new_n9404_), .A3(new_n9626_), .ZN(new_n9636_));
  AOI21_X1   g08634(.A1(new_n9632_), .A2(new_n9636_), .B(new_n9613_), .ZN(new_n9637_));
  NOR3_X1    g08635(.A1(new_n9625_), .A2(new_n9631_), .A3(new_n9630_), .ZN(new_n9638_));
  NOR3_X1    g08636(.A1(new_n9638_), .A2(new_n9624_), .A3(new_n9614_), .ZN(new_n9639_));
  NOR3_X1    g08637(.A1(new_n9639_), .A2(new_n9637_), .A3(new_n9572_), .ZN(new_n9640_));
  OAI21_X1   g08638(.A1(new_n9635_), .A2(new_n9640_), .B(new_n9609_), .ZN(new_n9641_));
  XOR2_X1    g08639(.A1(new_n9341_), .A2(new_n9586_), .Z(new_n9642_));
  NOR2_X1    g08640(.A1(new_n9600_), .A2(new_n9601_), .ZN(new_n9643_));
  NOR3_X1    g08641(.A1(new_n9643_), .A2(new_n9392_), .A3(new_n9393_), .ZN(new_n9644_));
  OAI21_X1   g08642(.A1(new_n9644_), .A2(new_n9607_), .B(new_n9642_), .ZN(new_n9645_));
  NAND2_X1   g08643(.A1(new_n9603_), .A2(new_n9593_), .ZN(new_n9646_));
  NOR2_X1    g08644(.A1(new_n9646_), .A2(new_n9589_), .ZN(new_n9647_));
  XOR2_X1    g08645(.A1(new_n9589_), .A2(new_n9598_), .Z(new_n9648_));
  OAI22_X1   g08646(.A1(new_n9648_), .A2(new_n9642_), .B1(new_n9645_), .B2(new_n9647_), .ZN(new_n9649_));
  OAI21_X1   g08647(.A1(new_n9639_), .A2(new_n9637_), .B(new_n9572_), .ZN(new_n9650_));
  NAND3_X1   g08648(.A1(new_n9629_), .A2(new_n9634_), .A3(new_n9401_), .ZN(new_n9651_));
  NAND3_X1   g08649(.A1(new_n9650_), .A2(new_n9649_), .A3(new_n9651_), .ZN(new_n9652_));
  AOI21_X1   g08650(.A1(new_n9641_), .A2(new_n9652_), .B(new_n9583_), .ZN(new_n9653_));
  AOI21_X1   g08651(.A1(new_n9650_), .A2(new_n9651_), .B(new_n9649_), .ZN(new_n9654_));
  NOR3_X1    g08652(.A1(new_n9640_), .A2(new_n9609_), .A3(new_n9635_), .ZN(new_n9655_));
  NOR3_X1    g08653(.A1(new_n9654_), .A2(new_n9655_), .A3(new_n9571_), .ZN(new_n9656_));
  XOR2_X1    g08654(.A1(new_n9564_), .A2(new_n9565_), .Z(new_n9657_));
  XOR2_X1    g08655(.A1(new_n9657_), .A2(new_n9510_), .Z(new_n9658_));
  NAND3_X1   g08656(.A1(new_n9563_), .A2(new_n9510_), .A3(new_n9521_), .ZN(new_n9659_));
  NOR2_X1    g08657(.A1(new_n9533_), .A2(new_n9557_), .ZN(new_n9660_));
  AOI21_X1   g08658(.A1(new_n9534_), .A2(new_n9540_), .B(new_n9541_), .ZN(new_n9661_));
  AOI21_X1   g08659(.A1(new_n9528_), .A2(new_n9529_), .B(new_n9531_), .ZN(new_n9662_));
  XNOR2_X1   g08660(.A1(new_n9661_), .A2(new_n9662_), .ZN(new_n9663_));
  XOR2_X1    g08661(.A1(new_n9660_), .A2(new_n9663_), .Z(new_n9664_));
  AOI21_X1   g08662(.A1(new_n9664_), .A2(new_n9659_), .B(new_n9658_), .ZN(new_n9665_));
  NOR4_X1    g08663(.A1(new_n9513_), .A2(new_n9515_), .A3(new_n9520_), .A4(new_n9518_), .ZN(new_n9666_));
  INV_X1     g08664(.I(new_n9521_), .ZN(new_n9667_));
  NOR3_X1    g08665(.A1(new_n9559_), .A2(new_n9666_), .A3(new_n9667_), .ZN(new_n9668_));
  NAND2_X1   g08666(.A1(new_n9661_), .A2(new_n9662_), .ZN(new_n9669_));
  INV_X1     g08667(.I(new_n9669_), .ZN(new_n9670_));
  AOI21_X1   g08668(.A1(new_n9563_), .A2(new_n9670_), .B(new_n9663_), .ZN(new_n9671_));
  NAND2_X1   g08669(.A1(new_n9668_), .A2(new_n9671_), .ZN(new_n9672_));
  NAND2_X1   g08670(.A1(new_n9665_), .A2(new_n9672_), .ZN(new_n9673_));
  NAND2_X1   g08671(.A1(new_n9664_), .A2(new_n9659_), .ZN(new_n9674_));
  NAND2_X1   g08672(.A1(new_n9660_), .A2(new_n9663_), .ZN(new_n9675_));
  XOR2_X1    g08673(.A1(new_n9661_), .A2(new_n9662_), .Z(new_n9676_));
  OAI21_X1   g08674(.A1(new_n9533_), .A2(new_n9557_), .B(new_n9676_), .ZN(new_n9677_));
  NAND2_X1   g08675(.A1(new_n9677_), .A2(new_n9675_), .ZN(new_n9678_));
  NAND2_X1   g08676(.A1(new_n9668_), .A2(new_n9678_), .ZN(new_n9679_));
  NAND2_X1   g08677(.A1(new_n9674_), .A2(new_n9679_), .ZN(new_n9680_));
  NAND2_X1   g08678(.A1(new_n9680_), .A2(new_n9658_), .ZN(new_n9681_));
  NAND2_X1   g08679(.A1(new_n9681_), .A2(new_n9673_), .ZN(new_n9682_));
  NAND2_X1   g08680(.A1(new_n9568_), .A2(new_n9569_), .ZN(new_n9683_));
  NOR2_X1    g08681(.A1(new_n9486_), .A2(new_n9487_), .ZN(new_n9684_));
  INV_X1     g08682(.I(new_n9487_), .ZN(new_n9685_));
  NOR2_X1    g08683(.A1(new_n9685_), .A2(new_n9485_), .ZN(new_n9686_));
  NOR2_X1    g08684(.A1(new_n9684_), .A2(new_n9686_), .ZN(new_n9687_));
  XOR2_X1    g08685(.A1(new_n9687_), .A2(new_n9438_), .Z(new_n9688_));
  NOR3_X1    g08686(.A1(new_n9478_), .A2(new_n9438_), .A3(new_n9441_), .ZN(new_n9689_));
  NAND4_X1   g08687(.A1(new_n9446_), .A2(new_n9451_), .A3(new_n9473_), .A4(new_n9475_), .ZN(new_n9690_));
  INV_X1     g08688(.I(new_n9690_), .ZN(new_n9691_));
  AOI21_X1   g08689(.A1(new_n9453_), .A2(new_n9459_), .B(new_n9460_), .ZN(new_n9692_));
  AOI21_X1   g08690(.A1(new_n9447_), .A2(new_n9448_), .B(new_n9450_), .ZN(new_n9693_));
  XOR2_X1    g08691(.A1(new_n9692_), .A2(new_n9693_), .Z(new_n9694_));
  NOR2_X1    g08692(.A1(new_n9691_), .A2(new_n9694_), .ZN(new_n9695_));
  XNOR2_X1   g08693(.A1(new_n9692_), .A2(new_n9693_), .ZN(new_n9696_));
  NOR2_X1    g08694(.A1(new_n9696_), .A2(new_n9690_), .ZN(new_n9697_));
  NOR2_X1    g08695(.A1(new_n9695_), .A2(new_n9697_), .ZN(new_n9698_));
  NAND3_X1   g08696(.A1(new_n9483_), .A2(new_n9692_), .A3(new_n9693_), .ZN(new_n9699_));
  AOI21_X1   g08697(.A1(new_n9698_), .A2(new_n9699_), .B(new_n9689_), .ZN(new_n9700_));
  NAND3_X1   g08698(.A1(new_n9483_), .A2(new_n9480_), .A3(new_n9488_), .ZN(new_n9701_));
  INV_X1     g08699(.I(new_n9692_), .ZN(new_n9702_));
  INV_X1     g08700(.I(new_n9693_), .ZN(new_n9703_));
  NOR3_X1    g08701(.A1(new_n9478_), .A2(new_n9702_), .A3(new_n9703_), .ZN(new_n9704_));
  NOR3_X1    g08702(.A1(new_n9704_), .A2(new_n9701_), .A3(new_n9696_), .ZN(new_n9705_));
  OAI21_X1   g08703(.A1(new_n9700_), .A2(new_n9705_), .B(new_n9688_), .ZN(new_n9706_));
  XNOR2_X1   g08704(.A1(new_n9687_), .A2(new_n9438_), .ZN(new_n9707_));
  XOR2_X1    g08705(.A1(new_n9694_), .A2(new_n9690_), .Z(new_n9708_));
  OAI21_X1   g08706(.A1(new_n9708_), .A2(new_n9704_), .B(new_n9701_), .ZN(new_n9709_));
  NAND3_X1   g08707(.A1(new_n9689_), .A2(new_n9699_), .A3(new_n9698_), .ZN(new_n9710_));
  NAND3_X1   g08708(.A1(new_n9709_), .A2(new_n9710_), .A3(new_n9707_), .ZN(new_n9711_));
  AOI21_X1   g08709(.A1(new_n9706_), .A2(new_n9711_), .B(new_n9683_), .ZN(new_n9712_));
  NAND3_X1   g08710(.A1(new_n9689_), .A2(new_n9699_), .A3(new_n9694_), .ZN(new_n9713_));
  AOI21_X1   g08711(.A1(new_n9709_), .A2(new_n9713_), .B(new_n9707_), .ZN(new_n9714_));
  NOR3_X1    g08712(.A1(new_n9708_), .A2(new_n9704_), .A3(new_n9701_), .ZN(new_n9715_));
  NOR3_X1    g08713(.A1(new_n9700_), .A2(new_n9715_), .A3(new_n9688_), .ZN(new_n9716_));
  NOR3_X1    g08714(.A1(new_n9716_), .A2(new_n9714_), .A3(new_n9567_), .ZN(new_n9717_));
  NOR3_X1    g08715(.A1(new_n9682_), .A2(new_n9717_), .A3(new_n9712_), .ZN(new_n9718_));
  AOI22_X1   g08716(.A1(new_n9680_), .A2(new_n9658_), .B1(new_n9665_), .B2(new_n9672_), .ZN(new_n9719_));
  OAI21_X1   g08717(.A1(new_n9716_), .A2(new_n9714_), .B(new_n9567_), .ZN(new_n9720_));
  NAND3_X1   g08718(.A1(new_n9706_), .A2(new_n9711_), .A3(new_n9683_), .ZN(new_n9721_));
  AOI21_X1   g08719(.A1(new_n9720_), .A2(new_n9721_), .B(new_n9719_), .ZN(new_n9722_));
  NOR2_X1    g08720(.A1(new_n9718_), .A2(new_n9722_), .ZN(new_n9723_));
  OAI21_X1   g08721(.A1(new_n9656_), .A2(new_n9653_), .B(new_n9723_), .ZN(new_n9724_));
  OAI21_X1   g08722(.A1(new_n9654_), .A2(new_n9655_), .B(new_n9571_), .ZN(new_n9725_));
  NAND3_X1   g08723(.A1(new_n9641_), .A2(new_n9652_), .A3(new_n9583_), .ZN(new_n9726_));
  NAND3_X1   g08724(.A1(new_n9720_), .A2(new_n9721_), .A3(new_n9719_), .ZN(new_n9727_));
  OAI21_X1   g08725(.A1(new_n9717_), .A2(new_n9712_), .B(new_n9682_), .ZN(new_n9728_));
  NAND2_X1   g08726(.A1(new_n9728_), .A2(new_n9727_), .ZN(new_n9729_));
  NAND3_X1   g08727(.A1(new_n9725_), .A2(new_n9729_), .A3(new_n9726_), .ZN(new_n9730_));
  AOI21_X1   g08728(.A1(new_n9730_), .A2(new_n9724_), .B(new_n9582_), .ZN(new_n9731_));
  INV_X1     g08729(.I(new_n9582_), .ZN(new_n9732_));
  AOI21_X1   g08730(.A1(new_n9725_), .A2(new_n9726_), .B(new_n9729_), .ZN(new_n9733_));
  NOR3_X1    g08731(.A1(new_n9656_), .A2(new_n9653_), .A3(new_n9723_), .ZN(new_n9734_));
  NOR3_X1    g08732(.A1(new_n9733_), .A2(new_n9734_), .A3(new_n9732_), .ZN(new_n9735_));
  NOR3_X1    g08733(.A1(new_n9735_), .A2(new_n9731_), .A3(new_n9234_), .ZN(new_n9736_));
  NOR3_X1    g08734(.A1(new_n9232_), .A2(new_n9231_), .A3(new_n9230_), .ZN(new_n9737_));
  AOI21_X1   g08735(.A1(new_n9222_), .A2(new_n9226_), .B(new_n8981_), .ZN(new_n9738_));
  NOR2_X1    g08736(.A1(new_n9738_), .A2(new_n9737_), .ZN(new_n9739_));
  OAI21_X1   g08737(.A1(new_n9733_), .A2(new_n9734_), .B(new_n9732_), .ZN(new_n9740_));
  NAND3_X1   g08738(.A1(new_n9730_), .A2(new_n9724_), .A3(new_n9582_), .ZN(new_n9741_));
  AOI21_X1   g08739(.A1(new_n9740_), .A2(new_n9741_), .B(new_n9739_), .ZN(new_n9742_));
  XNOR2_X1   g08740(.A1(new_n9581_), .A2(new_n9577_), .ZN(new_n9743_));
  NOR2_X1    g08741(.A1(new_n7120_), .A2(new_n7121_), .ZN(new_n9744_));
  XNOR2_X1   g08742(.A1(new_n7696_), .A2(new_n7453_), .ZN(new_n9745_));
  NOR2_X1    g08743(.A1(new_n9745_), .A2(new_n9744_), .ZN(new_n9746_));
  OR3_X2     g08744(.A1(new_n9746_), .A2(new_n9743_), .A3(new_n7698_), .Z(new_n9747_));
  OAI21_X1   g08745(.A1(new_n9736_), .A2(new_n9742_), .B(new_n9747_), .ZN(new_n9748_));
  OAI21_X1   g08746(.A1(new_n9739_), .A2(new_n9731_), .B(new_n9741_), .ZN(new_n9749_));
  AOI21_X1   g08747(.A1(new_n9230_), .A2(new_n9222_), .B(new_n9232_), .ZN(new_n9750_));
  OAI21_X1   g08748(.A1(new_n8847_), .A2(new_n8970_), .B(new_n8979_), .ZN(new_n9751_));
  OAI21_X1   g08749(.A1(new_n8951_), .A2(new_n8956_), .B(new_n8972_), .ZN(new_n9752_));
  AOI21_X1   g08750(.A1(new_n8924_), .A2(new_n8926_), .B(new_n8952_), .ZN(new_n9753_));
  NOR2_X1    g08751(.A1(new_n9753_), .A2(new_n8927_), .ZN(new_n9754_));
  INV_X1     g08752(.I(new_n8943_), .ZN(new_n9755_));
  OAI21_X1   g08753(.A1(new_n8942_), .A2(new_n8944_), .B(new_n9755_), .ZN(new_n9756_));
  NAND2_X1   g08754(.A1(new_n9754_), .A2(new_n9756_), .ZN(new_n9757_));
  INV_X1     g08755(.I(new_n9757_), .ZN(new_n9758_));
  NOR2_X1    g08756(.A1(new_n9754_), .A2(new_n9756_), .ZN(new_n9759_));
  NOR2_X1    g08757(.A1(new_n9758_), .A2(new_n9759_), .ZN(new_n9760_));
  NAND2_X1   g08758(.A1(new_n9752_), .A2(new_n9760_), .ZN(new_n9761_));
  NAND2_X1   g08759(.A1(new_n8967_), .A2(new_n8946_), .ZN(new_n9762_));
  INV_X1     g08760(.I(new_n9759_), .ZN(new_n9763_));
  NAND2_X1   g08761(.A1(new_n9763_), .A2(new_n9757_), .ZN(new_n9764_));
  NAND3_X1   g08762(.A1(new_n9762_), .A2(new_n9764_), .A3(new_n8972_), .ZN(new_n9765_));
  NAND2_X1   g08763(.A1(new_n9761_), .A2(new_n9765_), .ZN(new_n9766_));
  NOR3_X1    g08764(.A1(new_n8814_), .A2(new_n8800_), .A3(new_n8816_), .ZN(new_n9767_));
  NOR2_X1    g08765(.A1(new_n8839_), .A2(new_n8817_), .ZN(new_n9768_));
  NOR3_X1    g08766(.A1(new_n9768_), .A2(new_n8810_), .A3(new_n8815_), .ZN(new_n9769_));
  NOR2_X1    g08767(.A1(new_n9769_), .A2(new_n9767_), .ZN(new_n9770_));
  INV_X1     g08768(.I(new_n9770_), .ZN(new_n9771_));
  AOI22_X1   g08769(.A1(new_n8840_), .A2(new_n8841_), .B1(new_n8788_), .B2(new_n8792_), .ZN(new_n9772_));
  AOI21_X1   g08770(.A1(new_n8781_), .A2(new_n8790_), .B(new_n8785_), .ZN(new_n9773_));
  NOR3_X1    g08771(.A1(new_n9772_), .A2(new_n8842_), .A3(new_n9773_), .ZN(new_n9774_));
  INV_X1     g08772(.I(new_n9773_), .ZN(new_n9775_));
  AOI21_X1   g08773(.A1(new_n8838_), .A2(new_n8845_), .B(new_n9775_), .ZN(new_n9776_));
  NOR3_X1    g08774(.A1(new_n9774_), .A2(new_n9776_), .A3(new_n9771_), .ZN(new_n9777_));
  NAND3_X1   g08775(.A1(new_n8838_), .A2(new_n8845_), .A3(new_n9775_), .ZN(new_n9778_));
  OAI21_X1   g08776(.A1(new_n9772_), .A2(new_n8842_), .B(new_n9773_), .ZN(new_n9779_));
  AOI21_X1   g08777(.A1(new_n9779_), .A2(new_n9778_), .B(new_n9770_), .ZN(new_n9780_));
  NOR2_X1    g08778(.A1(new_n9777_), .A2(new_n9780_), .ZN(new_n9781_));
  NAND2_X1   g08779(.A1(new_n9781_), .A2(new_n9766_), .ZN(new_n9782_));
  AOI21_X1   g08780(.A1(new_n9762_), .A2(new_n8972_), .B(new_n9764_), .ZN(new_n9783_));
  NOR2_X1    g08781(.A1(new_n9752_), .A2(new_n9760_), .ZN(new_n9784_));
  NOR2_X1    g08782(.A1(new_n9784_), .A2(new_n9783_), .ZN(new_n9785_));
  NAND3_X1   g08783(.A1(new_n9779_), .A2(new_n9778_), .A3(new_n9770_), .ZN(new_n9786_));
  OAI21_X1   g08784(.A1(new_n9774_), .A2(new_n9776_), .B(new_n9771_), .ZN(new_n9787_));
  NAND2_X1   g08785(.A1(new_n9787_), .A2(new_n9786_), .ZN(new_n9788_));
  NAND2_X1   g08786(.A1(new_n9785_), .A2(new_n9788_), .ZN(new_n9789_));
  NAND3_X1   g08787(.A1(new_n9782_), .A2(new_n9789_), .A3(new_n9751_), .ZN(new_n9790_));
  AOI21_X1   g08788(.A1(new_n8978_), .A2(new_n8848_), .B(new_n8976_), .ZN(new_n9791_));
  NOR2_X1    g08789(.A1(new_n9785_), .A2(new_n9788_), .ZN(new_n9792_));
  NOR2_X1    g08790(.A1(new_n9781_), .A2(new_n9766_), .ZN(new_n9793_));
  OAI21_X1   g08791(.A1(new_n9793_), .A2(new_n9792_), .B(new_n9791_), .ZN(new_n9794_));
  OAI21_X1   g08792(.A1(new_n9218_), .A2(new_n9219_), .B(new_n9210_), .ZN(new_n9795_));
  NAND2_X1   g08793(.A1(new_n9190_), .A2(new_n9194_), .ZN(new_n9796_));
  AOI21_X1   g08794(.A1(new_n9053_), .A2(new_n9055_), .B(new_n9187_), .ZN(new_n9797_));
  NOR2_X1    g08795(.A1(new_n9797_), .A2(new_n9056_), .ZN(new_n9798_));
  NOR2_X1    g08796(.A1(new_n9039_), .A2(new_n9182_), .ZN(new_n9799_));
  NOR2_X1    g08797(.A1(new_n9799_), .A2(new_n9181_), .ZN(new_n9800_));
  INV_X1     g08798(.I(new_n9800_), .ZN(new_n9801_));
  NAND2_X1   g08799(.A1(new_n9801_), .A2(new_n9798_), .ZN(new_n9802_));
  INV_X1     g08800(.I(new_n9798_), .ZN(new_n9803_));
  NAND2_X1   g08801(.A1(new_n9803_), .A2(new_n9800_), .ZN(new_n9804_));
  NAND2_X1   g08802(.A1(new_n9804_), .A2(new_n9802_), .ZN(new_n9805_));
  AOI21_X1   g08803(.A1(new_n9796_), .A2(new_n9192_), .B(new_n9805_), .ZN(new_n9806_));
  NOR2_X1    g08804(.A1(new_n9201_), .A2(new_n9184_), .ZN(new_n9807_));
  NOR2_X1    g08805(.A1(new_n9803_), .A2(new_n9800_), .ZN(new_n9808_));
  NOR2_X1    g08806(.A1(new_n9801_), .A2(new_n9798_), .ZN(new_n9809_));
  NOR2_X1    g08807(.A1(new_n9808_), .A2(new_n9809_), .ZN(new_n9810_));
  NOR3_X1    g08808(.A1(new_n9807_), .A2(new_n9810_), .A3(new_n9206_), .ZN(new_n9811_));
  NOR2_X1    g08809(.A1(new_n9163_), .A2(new_n9164_), .ZN(new_n9812_));
  INV_X1     g08810(.I(new_n9812_), .ZN(new_n9813_));
  OAI21_X1   g08811(.A1(new_n9162_), .A2(new_n9214_), .B(new_n9813_), .ZN(new_n9814_));
  NOR2_X1    g08812(.A1(new_n9136_), .A2(new_n9137_), .ZN(new_n9815_));
  NAND2_X1   g08813(.A1(new_n9136_), .A2(new_n9137_), .ZN(new_n9816_));
  AOI21_X1   g08814(.A1(new_n9086_), .A2(new_n9816_), .B(new_n9815_), .ZN(new_n9817_));
  NOR3_X1    g08815(.A1(new_n9213_), .A2(new_n9174_), .A3(new_n9817_), .ZN(new_n9818_));
  INV_X1     g08816(.I(new_n9817_), .ZN(new_n9819_));
  AOI21_X1   g08817(.A1(new_n9167_), .A2(new_n9216_), .B(new_n9819_), .ZN(new_n9820_));
  NOR3_X1    g08818(.A1(new_n9818_), .A2(new_n9820_), .A3(new_n9814_), .ZN(new_n9821_));
  INV_X1     g08819(.I(new_n9814_), .ZN(new_n9822_));
  NAND3_X1   g08820(.A1(new_n9167_), .A2(new_n9216_), .A3(new_n9819_), .ZN(new_n9823_));
  OAI21_X1   g08821(.A1(new_n9213_), .A2(new_n9174_), .B(new_n9817_), .ZN(new_n9824_));
  AOI21_X1   g08822(.A1(new_n9824_), .A2(new_n9823_), .B(new_n9822_), .ZN(new_n9825_));
  OAI22_X1   g08823(.A1(new_n9821_), .A2(new_n9825_), .B1(new_n9806_), .B2(new_n9811_), .ZN(new_n9826_));
  OAI21_X1   g08824(.A1(new_n9807_), .A2(new_n9206_), .B(new_n9810_), .ZN(new_n9827_));
  NAND3_X1   g08825(.A1(new_n9796_), .A2(new_n9805_), .A3(new_n9192_), .ZN(new_n9828_));
  NAND3_X1   g08826(.A1(new_n9824_), .A2(new_n9823_), .A3(new_n9822_), .ZN(new_n9829_));
  OAI21_X1   g08827(.A1(new_n9818_), .A2(new_n9820_), .B(new_n9814_), .ZN(new_n9830_));
  NAND4_X1   g08828(.A1(new_n9830_), .A2(new_n9829_), .A3(new_n9827_), .A4(new_n9828_), .ZN(new_n9831_));
  NAND3_X1   g08829(.A1(new_n9826_), .A2(new_n9795_), .A3(new_n9831_), .ZN(new_n9832_));
  AOI21_X1   g08830(.A1(new_n9180_), .A2(new_n9204_), .B(new_n9220_), .ZN(new_n9833_));
  AOI22_X1   g08831(.A1(new_n9830_), .A2(new_n9829_), .B1(new_n9827_), .B2(new_n9828_), .ZN(new_n9834_));
  NOR4_X1    g08832(.A1(new_n9821_), .A2(new_n9825_), .A3(new_n9806_), .A4(new_n9811_), .ZN(new_n9835_));
  OAI21_X1   g08833(.A1(new_n9835_), .A2(new_n9834_), .B(new_n9833_), .ZN(new_n9836_));
  AOI22_X1   g08834(.A1(new_n9794_), .A2(new_n9790_), .B1(new_n9836_), .B2(new_n9832_), .ZN(new_n9837_));
  NOR3_X1    g08835(.A1(new_n9793_), .A2(new_n9792_), .A3(new_n9791_), .ZN(new_n9838_));
  AOI21_X1   g08836(.A1(new_n9782_), .A2(new_n9789_), .B(new_n9751_), .ZN(new_n9839_));
  NOR3_X1    g08837(.A1(new_n9834_), .A2(new_n9835_), .A3(new_n9833_), .ZN(new_n9840_));
  AOI21_X1   g08838(.A1(new_n9826_), .A2(new_n9831_), .B(new_n9795_), .ZN(new_n9841_));
  NOR4_X1    g08839(.A1(new_n9839_), .A2(new_n9838_), .A3(new_n9840_), .A4(new_n9841_), .ZN(new_n9842_));
  NOR3_X1    g08840(.A1(new_n9842_), .A2(new_n9837_), .A3(new_n9750_), .ZN(new_n9843_));
  OAI21_X1   g08841(.A1(new_n8981_), .A2(new_n9231_), .B(new_n9226_), .ZN(new_n9844_));
  OAI22_X1   g08842(.A1(new_n9839_), .A2(new_n9838_), .B1(new_n9840_), .B2(new_n9841_), .ZN(new_n9845_));
  NAND4_X1   g08843(.A1(new_n9794_), .A2(new_n9790_), .A3(new_n9836_), .A4(new_n9832_), .ZN(new_n9846_));
  AOI21_X1   g08844(.A1(new_n9845_), .A2(new_n9846_), .B(new_n9844_), .ZN(new_n9847_));
  AOI21_X1   g08845(.A1(new_n9725_), .A2(new_n9729_), .B(new_n9656_), .ZN(new_n9848_));
  OAI21_X1   g08846(.A1(new_n9719_), .A2(new_n9712_), .B(new_n9721_), .ZN(new_n9849_));
  NAND2_X1   g08847(.A1(new_n9709_), .A2(new_n9688_), .ZN(new_n9850_));
  NAND2_X1   g08848(.A1(new_n9691_), .A2(new_n9693_), .ZN(new_n9851_));
  OAI21_X1   g08849(.A1(new_n9691_), .A2(new_n9693_), .B(new_n9692_), .ZN(new_n9852_));
  INV_X1     g08850(.I(new_n9684_), .ZN(new_n9853_));
  OAI21_X1   g08851(.A1(new_n9438_), .A2(new_n9686_), .B(new_n9853_), .ZN(new_n9854_));
  NAND3_X1   g08852(.A1(new_n9854_), .A2(new_n9852_), .A3(new_n9851_), .ZN(new_n9855_));
  NAND2_X1   g08853(.A1(new_n9852_), .A2(new_n9851_), .ZN(new_n9856_));
  NOR2_X1    g08854(.A1(new_n9438_), .A2(new_n9686_), .ZN(new_n9857_));
  NOR2_X1    g08855(.A1(new_n9857_), .A2(new_n9684_), .ZN(new_n9858_));
  NAND2_X1   g08856(.A1(new_n9856_), .A2(new_n9858_), .ZN(new_n9859_));
  NAND2_X1   g08857(.A1(new_n9859_), .A2(new_n9855_), .ZN(new_n9860_));
  AOI21_X1   g08858(.A1(new_n9850_), .A2(new_n9713_), .B(new_n9860_), .ZN(new_n9861_));
  NOR2_X1    g08859(.A1(new_n9700_), .A2(new_n9707_), .ZN(new_n9862_));
  INV_X1     g08860(.I(new_n9855_), .ZN(new_n9863_));
  AOI21_X1   g08861(.A1(new_n9852_), .A2(new_n9851_), .B(new_n9854_), .ZN(new_n9864_));
  NOR2_X1    g08862(.A1(new_n9863_), .A2(new_n9864_), .ZN(new_n9865_));
  NOR3_X1    g08863(.A1(new_n9862_), .A2(new_n9865_), .A3(new_n9705_), .ZN(new_n9866_));
  NOR2_X1    g08864(.A1(new_n9661_), .A2(new_n9662_), .ZN(new_n9867_));
  INV_X1     g08865(.I(new_n9867_), .ZN(new_n9868_));
  OAI21_X1   g08866(.A1(new_n9660_), .A2(new_n9670_), .B(new_n9868_), .ZN(new_n9869_));
  OAI21_X1   g08867(.A1(new_n9559_), .A2(new_n9669_), .B(new_n9676_), .ZN(new_n9870_));
  NOR2_X1    g08868(.A1(new_n9870_), .A2(new_n9659_), .ZN(new_n9871_));
  NOR2_X1    g08869(.A1(new_n9564_), .A2(new_n9565_), .ZN(new_n9872_));
  NAND2_X1   g08870(.A1(new_n9564_), .A2(new_n9565_), .ZN(new_n9873_));
  AOI21_X1   g08871(.A1(new_n9510_), .A2(new_n9873_), .B(new_n9872_), .ZN(new_n9874_));
  NOR3_X1    g08872(.A1(new_n9665_), .A2(new_n9871_), .A3(new_n9874_), .ZN(new_n9875_));
  NAND2_X1   g08873(.A1(new_n9657_), .A2(new_n9510_), .ZN(new_n9876_));
  INV_X1     g08874(.I(new_n9873_), .ZN(new_n9877_));
  OAI21_X1   g08875(.A1(new_n9872_), .A2(new_n9877_), .B(new_n9666_), .ZN(new_n9878_));
  NAND2_X1   g08876(.A1(new_n9878_), .A2(new_n9876_), .ZN(new_n9879_));
  OAI21_X1   g08877(.A1(new_n9668_), .A2(new_n9678_), .B(new_n9879_), .ZN(new_n9880_));
  INV_X1     g08878(.I(new_n9874_), .ZN(new_n9881_));
  AOI21_X1   g08879(.A1(new_n9880_), .A2(new_n9672_), .B(new_n9881_), .ZN(new_n9882_));
  NOR3_X1    g08880(.A1(new_n9875_), .A2(new_n9882_), .A3(new_n9869_), .ZN(new_n9883_));
  INV_X1     g08881(.I(new_n9869_), .ZN(new_n9884_));
  NAND3_X1   g08882(.A1(new_n9880_), .A2(new_n9672_), .A3(new_n9881_), .ZN(new_n9885_));
  OAI21_X1   g08883(.A1(new_n9665_), .A2(new_n9871_), .B(new_n9874_), .ZN(new_n9886_));
  AOI21_X1   g08884(.A1(new_n9886_), .A2(new_n9885_), .B(new_n9884_), .ZN(new_n9887_));
  OAI22_X1   g08885(.A1(new_n9883_), .A2(new_n9887_), .B1(new_n9866_), .B2(new_n9861_), .ZN(new_n9888_));
  OAI21_X1   g08886(.A1(new_n9862_), .A2(new_n9705_), .B(new_n9865_), .ZN(new_n9889_));
  NAND3_X1   g08887(.A1(new_n9850_), .A2(new_n9713_), .A3(new_n9860_), .ZN(new_n9890_));
  NAND3_X1   g08888(.A1(new_n9886_), .A2(new_n9885_), .A3(new_n9884_), .ZN(new_n9891_));
  OAI21_X1   g08889(.A1(new_n9875_), .A2(new_n9882_), .B(new_n9869_), .ZN(new_n9892_));
  NAND4_X1   g08890(.A1(new_n9892_), .A2(new_n9891_), .A3(new_n9889_), .A4(new_n9890_), .ZN(new_n9893_));
  NAND3_X1   g08891(.A1(new_n9849_), .A2(new_n9888_), .A3(new_n9893_), .ZN(new_n9894_));
  AOI21_X1   g08892(.A1(new_n9682_), .A2(new_n9720_), .B(new_n9717_), .ZN(new_n9895_));
  AOI22_X1   g08893(.A1(new_n9892_), .A2(new_n9891_), .B1(new_n9889_), .B2(new_n9890_), .ZN(new_n9896_));
  NOR4_X1    g08894(.A1(new_n9883_), .A2(new_n9887_), .A3(new_n9866_), .A4(new_n9861_), .ZN(new_n9897_));
  OAI21_X1   g08895(.A1(new_n9896_), .A2(new_n9897_), .B(new_n9895_), .ZN(new_n9898_));
  OAI21_X1   g08896(.A1(new_n9609_), .A2(new_n9635_), .B(new_n9651_), .ZN(new_n9899_));
  NAND2_X1   g08897(.A1(new_n9632_), .A2(new_n9614_), .ZN(new_n9900_));
  AOI21_X1   g08898(.A1(new_n9405_), .A2(new_n9406_), .B(new_n9307_), .ZN(new_n9901_));
  NOR2_X1    g08899(.A1(new_n9901_), .A2(new_n9407_), .ZN(new_n9902_));
  INV_X1     g08900(.I(new_n9610_), .ZN(new_n9903_));
  OAI21_X1   g08901(.A1(new_n9315_), .A2(new_n9611_), .B(new_n9903_), .ZN(new_n9904_));
  NAND2_X1   g08902(.A1(new_n9902_), .A2(new_n9904_), .ZN(new_n9905_));
  NOR2_X1    g08903(.A1(new_n9902_), .A2(new_n9904_), .ZN(new_n9906_));
  INV_X1     g08904(.I(new_n9906_), .ZN(new_n9907_));
  NAND2_X1   g08905(.A1(new_n9907_), .A2(new_n9905_), .ZN(new_n9908_));
  AOI21_X1   g08906(.A1(new_n9900_), .A2(new_n9636_), .B(new_n9908_), .ZN(new_n9909_));
  NOR2_X1    g08907(.A1(new_n9624_), .A2(new_n9613_), .ZN(new_n9910_));
  INV_X1     g08908(.I(new_n9905_), .ZN(new_n9911_));
  NOR2_X1    g08909(.A1(new_n9911_), .A2(new_n9906_), .ZN(new_n9912_));
  NOR3_X1    g08910(.A1(new_n9910_), .A2(new_n9912_), .A3(new_n9628_), .ZN(new_n9913_));
  NOR2_X1    g08911(.A1(new_n9590_), .A2(new_n9592_), .ZN(new_n9914_));
  INV_X1     g08912(.I(new_n9914_), .ZN(new_n9915_));
  OAI21_X1   g08913(.A1(new_n9595_), .A2(new_n9602_), .B(new_n9915_), .ZN(new_n9916_));
  NAND2_X1   g08914(.A1(new_n9341_), .A2(new_n9585_), .ZN(new_n9917_));
  NAND2_X1   g08915(.A1(new_n9917_), .A2(new_n9584_), .ZN(new_n9918_));
  INV_X1     g08916(.I(new_n9918_), .ZN(new_n9919_));
  NOR3_X1    g08917(.A1(new_n9599_), .A2(new_n9647_), .A3(new_n9919_), .ZN(new_n9920_));
  AOI21_X1   g08918(.A1(new_n9645_), .A2(new_n9604_), .B(new_n9918_), .ZN(new_n9921_));
  NOR3_X1    g08919(.A1(new_n9920_), .A2(new_n9921_), .A3(new_n9916_), .ZN(new_n9922_));
  INV_X1     g08920(.I(new_n9916_), .ZN(new_n9923_));
  NAND3_X1   g08921(.A1(new_n9645_), .A2(new_n9604_), .A3(new_n9918_), .ZN(new_n9924_));
  OAI21_X1   g08922(.A1(new_n9599_), .A2(new_n9647_), .B(new_n9919_), .ZN(new_n9925_));
  AOI21_X1   g08923(.A1(new_n9925_), .A2(new_n9924_), .B(new_n9923_), .ZN(new_n9926_));
  OAI22_X1   g08924(.A1(new_n9922_), .A2(new_n9926_), .B1(new_n9909_), .B2(new_n9913_), .ZN(new_n9927_));
  OAI21_X1   g08925(.A1(new_n9910_), .A2(new_n9628_), .B(new_n9912_), .ZN(new_n9928_));
  NAND3_X1   g08926(.A1(new_n9900_), .A2(new_n9908_), .A3(new_n9636_), .ZN(new_n9929_));
  NAND3_X1   g08927(.A1(new_n9925_), .A2(new_n9924_), .A3(new_n9923_), .ZN(new_n9930_));
  OAI21_X1   g08928(.A1(new_n9920_), .A2(new_n9921_), .B(new_n9916_), .ZN(new_n9931_));
  NAND4_X1   g08929(.A1(new_n9931_), .A2(new_n9930_), .A3(new_n9928_), .A4(new_n9929_), .ZN(new_n9932_));
  NAND3_X1   g08930(.A1(new_n9927_), .A2(new_n9899_), .A3(new_n9932_), .ZN(new_n9933_));
  AOI21_X1   g08931(.A1(new_n9649_), .A2(new_n9650_), .B(new_n9640_), .ZN(new_n9934_));
  AOI22_X1   g08932(.A1(new_n9931_), .A2(new_n9930_), .B1(new_n9928_), .B2(new_n9929_), .ZN(new_n9935_));
  NOR4_X1    g08933(.A1(new_n9922_), .A2(new_n9926_), .A3(new_n9909_), .A4(new_n9913_), .ZN(new_n9936_));
  OAI21_X1   g08934(.A1(new_n9935_), .A2(new_n9936_), .B(new_n9934_), .ZN(new_n9937_));
  AOI22_X1   g08935(.A1(new_n9898_), .A2(new_n9894_), .B1(new_n9937_), .B2(new_n9933_), .ZN(new_n9938_));
  NOR3_X1    g08936(.A1(new_n9895_), .A2(new_n9896_), .A3(new_n9897_), .ZN(new_n9939_));
  AOI21_X1   g08937(.A1(new_n9888_), .A2(new_n9893_), .B(new_n9849_), .ZN(new_n9940_));
  NOR3_X1    g08938(.A1(new_n9934_), .A2(new_n9936_), .A3(new_n9935_), .ZN(new_n9941_));
  AOI21_X1   g08939(.A1(new_n9927_), .A2(new_n9932_), .B(new_n9899_), .ZN(new_n9942_));
  NOR4_X1    g08940(.A1(new_n9939_), .A2(new_n9940_), .A3(new_n9941_), .A4(new_n9942_), .ZN(new_n9943_));
  NOR3_X1    g08941(.A1(new_n9938_), .A2(new_n9943_), .A3(new_n9848_), .ZN(new_n9944_));
  OAI21_X1   g08942(.A1(new_n9723_), .A2(new_n9653_), .B(new_n9726_), .ZN(new_n9945_));
  OAI22_X1   g08943(.A1(new_n9939_), .A2(new_n9940_), .B1(new_n9941_), .B2(new_n9942_), .ZN(new_n9946_));
  NAND4_X1   g08944(.A1(new_n9898_), .A2(new_n9937_), .A3(new_n9894_), .A4(new_n9933_), .ZN(new_n9947_));
  AOI21_X1   g08945(.A1(new_n9946_), .A2(new_n9947_), .B(new_n9945_), .ZN(new_n9948_));
  OAI22_X1   g08946(.A1(new_n9843_), .A2(new_n9847_), .B1(new_n9944_), .B2(new_n9948_), .ZN(new_n9949_));
  NAND3_X1   g08947(.A1(new_n9845_), .A2(new_n9846_), .A3(new_n9844_), .ZN(new_n9950_));
  OAI21_X1   g08948(.A1(new_n9842_), .A2(new_n9837_), .B(new_n9750_), .ZN(new_n9951_));
  NAND3_X1   g08949(.A1(new_n9946_), .A2(new_n9947_), .A3(new_n9945_), .ZN(new_n9952_));
  OAI21_X1   g08950(.A1(new_n9938_), .A2(new_n9943_), .B(new_n9848_), .ZN(new_n9953_));
  NAND4_X1   g08951(.A1(new_n9951_), .A2(new_n9950_), .A3(new_n9953_), .A4(new_n9952_), .ZN(new_n9954_));
  NAND3_X1   g08952(.A1(new_n9949_), .A2(new_n9954_), .A3(new_n9749_), .ZN(new_n9955_));
  INV_X1     g08953(.I(new_n9749_), .ZN(new_n9956_));
  AOI22_X1   g08954(.A1(new_n9951_), .A2(new_n9950_), .B1(new_n9953_), .B2(new_n9952_), .ZN(new_n9957_));
  NOR4_X1    g08955(.A1(new_n9843_), .A2(new_n9847_), .A3(new_n9944_), .A4(new_n9948_), .ZN(new_n9958_));
  OAI21_X1   g08956(.A1(new_n9958_), .A2(new_n9957_), .B(new_n9956_), .ZN(new_n9959_));
  NAND2_X1   g08957(.A1(new_n9959_), .A2(new_n9955_), .ZN(new_n9960_));
  NAND2_X1   g08958(.A1(new_n9745_), .A2(new_n9744_), .ZN(new_n9961_));
  OAI21_X1   g08959(.A1(new_n8071_), .A2(new_n8070_), .B(new_n8069_), .ZN(new_n9962_));
  NAND3_X1   g08960(.A1(new_n8062_), .A2(new_n8065_), .A3(new_n7853_), .ZN(new_n9963_));
  AOI21_X1   g08961(.A1(new_n9962_), .A2(new_n9963_), .B(new_n9961_), .ZN(new_n9964_));
  XOR2_X1    g08962(.A1(new_n8241_), .A2(new_n7119_), .Z(new_n9965_));
  OAI21_X1   g08963(.A1(new_n8074_), .A2(new_n9964_), .B(new_n9965_), .ZN(new_n9966_));
  NAND3_X1   g08964(.A1(new_n9962_), .A2(new_n9963_), .A3(new_n9961_), .ZN(new_n9967_));
  NAND3_X1   g08965(.A1(new_n8073_), .A2(new_n9967_), .A3(new_n8243_), .ZN(new_n9968_));
  NAND3_X1   g08966(.A1(new_n9739_), .A2(new_n9740_), .A3(new_n9741_), .ZN(new_n9969_));
  OAI21_X1   g08967(.A1(new_n9735_), .A2(new_n9731_), .B(new_n9234_), .ZN(new_n9970_));
  NAND2_X1   g08968(.A1(new_n7697_), .A2(new_n7122_), .ZN(new_n9971_));
  NAND2_X1   g08969(.A1(new_n9961_), .A2(new_n9971_), .ZN(new_n9972_));
  NOR2_X1    g08970(.A1(new_n9972_), .A2(new_n9743_), .ZN(new_n9973_));
  NAND3_X1   g08971(.A1(new_n9973_), .A2(new_n9970_), .A3(new_n9969_), .ZN(new_n9974_));
  NAND3_X1   g08972(.A1(new_n9966_), .A2(new_n9968_), .A3(new_n9974_), .ZN(new_n9975_));
  AOI21_X1   g08973(.A1(new_n9748_), .A2(new_n9975_), .B(new_n9960_), .ZN(new_n9976_));
  AOI21_X1   g08974(.A1(new_n9749_), .A2(new_n9949_), .B(new_n9958_), .ZN(new_n9977_));
  OAI21_X1   g08975(.A1(new_n9938_), .A2(new_n9848_), .B(new_n9947_), .ZN(new_n9978_));
  NOR2_X1    g08976(.A1(new_n9935_), .A2(new_n9899_), .ZN(new_n9979_));
  NOR2_X1    g08977(.A1(new_n9979_), .A2(new_n9936_), .ZN(new_n9980_));
  OAI21_X1   g08978(.A1(new_n9923_), .A2(new_n9921_), .B(new_n9924_), .ZN(new_n9981_));
  NAND2_X1   g08979(.A1(new_n9900_), .A2(new_n9636_), .ZN(new_n9982_));
  NAND2_X1   g08980(.A1(new_n9982_), .A2(new_n9905_), .ZN(new_n9983_));
  NAND3_X1   g08981(.A1(new_n9983_), .A2(new_n9907_), .A3(new_n9981_), .ZN(new_n9984_));
  AOI21_X1   g08982(.A1(new_n9916_), .A2(new_n9925_), .B(new_n9920_), .ZN(new_n9985_));
  NOR2_X1    g08983(.A1(new_n9910_), .A2(new_n9628_), .ZN(new_n9986_));
  OAI21_X1   g08984(.A1(new_n9986_), .A2(new_n9911_), .B(new_n9907_), .ZN(new_n9987_));
  NAND2_X1   g08985(.A1(new_n9987_), .A2(new_n9985_), .ZN(new_n9988_));
  AND2_X2    g08986(.A1(new_n9984_), .A2(new_n9988_), .Z(new_n9989_));
  NOR2_X1    g08987(.A1(new_n9980_), .A2(new_n9989_), .ZN(new_n9990_));
  NAND2_X1   g08988(.A1(new_n9984_), .A2(new_n9988_), .ZN(new_n9991_));
  NOR3_X1    g08989(.A1(new_n9991_), .A2(new_n9979_), .A3(new_n9936_), .ZN(new_n9992_));
  AOI21_X1   g08990(.A1(new_n9895_), .A2(new_n9888_), .B(new_n9897_), .ZN(new_n9993_));
  OAI21_X1   g08991(.A1(new_n9884_), .A2(new_n9882_), .B(new_n9885_), .ZN(new_n9994_));
  NAND2_X1   g08992(.A1(new_n9850_), .A2(new_n9713_), .ZN(new_n9995_));
  AOI21_X1   g08993(.A1(new_n9995_), .A2(new_n9855_), .B(new_n9864_), .ZN(new_n9996_));
  XOR2_X1    g08994(.A1(new_n9996_), .A2(new_n9994_), .Z(new_n9997_));
  NOR2_X1    g08995(.A1(new_n9997_), .A2(new_n9993_), .ZN(new_n9998_));
  OAI21_X1   g08996(.A1(new_n9896_), .A2(new_n9849_), .B(new_n9893_), .ZN(new_n9999_));
  NAND2_X1   g08997(.A1(new_n9996_), .A2(new_n9994_), .ZN(new_n10000_));
  INV_X1     g08998(.I(new_n9994_), .ZN(new_n10001_));
  NOR2_X1    g08999(.A1(new_n9862_), .A2(new_n9705_), .ZN(new_n10002_));
  OAI21_X1   g09000(.A1(new_n10002_), .A2(new_n9863_), .B(new_n9859_), .ZN(new_n10003_));
  NAND2_X1   g09001(.A1(new_n10003_), .A2(new_n10001_), .ZN(new_n10004_));
  NAND2_X1   g09002(.A1(new_n10004_), .A2(new_n10000_), .ZN(new_n10005_));
  NOR2_X1    g09003(.A1(new_n10005_), .A2(new_n9999_), .ZN(new_n10006_));
  OAI22_X1   g09004(.A1(new_n9990_), .A2(new_n9992_), .B1(new_n9998_), .B2(new_n10006_), .ZN(new_n10007_));
  OAI21_X1   g09005(.A1(new_n9936_), .A2(new_n9979_), .B(new_n9991_), .ZN(new_n10008_));
  NAND2_X1   g09006(.A1(new_n9980_), .A2(new_n9989_), .ZN(new_n10009_));
  NAND2_X1   g09007(.A1(new_n10005_), .A2(new_n9999_), .ZN(new_n10010_));
  NAND2_X1   g09008(.A1(new_n9997_), .A2(new_n9993_), .ZN(new_n10011_));
  NAND4_X1   g09009(.A1(new_n10009_), .A2(new_n10008_), .A3(new_n10011_), .A4(new_n10010_), .ZN(new_n10012_));
  NAND3_X1   g09010(.A1(new_n9978_), .A2(new_n10007_), .A3(new_n10012_), .ZN(new_n10013_));
  AOI21_X1   g09011(.A1(new_n9945_), .A2(new_n9946_), .B(new_n9943_), .ZN(new_n10014_));
  AOI22_X1   g09012(.A1(new_n10009_), .A2(new_n10008_), .B1(new_n10011_), .B2(new_n10010_), .ZN(new_n10015_));
  NOR4_X1    g09013(.A1(new_n9990_), .A2(new_n9998_), .A3(new_n9992_), .A4(new_n10006_), .ZN(new_n10016_));
  OAI21_X1   g09014(.A1(new_n10015_), .A2(new_n10016_), .B(new_n10014_), .ZN(new_n10017_));
  OAI21_X1   g09015(.A1(new_n9837_), .A2(new_n9750_), .B(new_n9846_), .ZN(new_n10018_));
  NAND2_X1   g09016(.A1(new_n9826_), .A2(new_n9833_), .ZN(new_n10019_));
  AOI21_X1   g09017(.A1(new_n9814_), .A2(new_n9824_), .B(new_n9818_), .ZN(new_n10020_));
  NOR2_X1    g09018(.A1(new_n9807_), .A2(new_n9206_), .ZN(new_n10021_));
  OAI21_X1   g09019(.A1(new_n10021_), .A2(new_n9808_), .B(new_n9804_), .ZN(new_n10022_));
  NOR2_X1    g09020(.A1(new_n10022_), .A2(new_n10020_), .ZN(new_n10023_));
  OAI21_X1   g09021(.A1(new_n9822_), .A2(new_n9820_), .B(new_n9823_), .ZN(new_n10024_));
  NAND2_X1   g09022(.A1(new_n9796_), .A2(new_n9192_), .ZN(new_n10025_));
  AOI21_X1   g09023(.A1(new_n10025_), .A2(new_n9802_), .B(new_n9809_), .ZN(new_n10026_));
  NOR2_X1    g09024(.A1(new_n10026_), .A2(new_n10024_), .ZN(new_n10027_));
  NOR2_X1    g09025(.A1(new_n10023_), .A2(new_n10027_), .ZN(new_n10028_));
  AOI21_X1   g09026(.A1(new_n9831_), .A2(new_n10019_), .B(new_n10028_), .ZN(new_n10029_));
  NOR2_X1    g09027(.A1(new_n9834_), .A2(new_n9795_), .ZN(new_n10030_));
  NAND2_X1   g09028(.A1(new_n10026_), .A2(new_n10024_), .ZN(new_n10031_));
  NAND2_X1   g09029(.A1(new_n10022_), .A2(new_n10020_), .ZN(new_n10032_));
  NAND2_X1   g09030(.A1(new_n10032_), .A2(new_n10031_), .ZN(new_n10033_));
  NOR3_X1    g09031(.A1(new_n10033_), .A2(new_n10030_), .A3(new_n9835_), .ZN(new_n10034_));
  NAND2_X1   g09032(.A1(new_n9782_), .A2(new_n9791_), .ZN(new_n10035_));
  AOI21_X1   g09033(.A1(new_n9770_), .A2(new_n9779_), .B(new_n9774_), .ZN(new_n10036_));
  AOI21_X1   g09034(.A1(new_n9752_), .A2(new_n9757_), .B(new_n9759_), .ZN(new_n10037_));
  INV_X1     g09035(.I(new_n10037_), .ZN(new_n10038_));
  NOR2_X1    g09036(.A1(new_n10038_), .A2(new_n10036_), .ZN(new_n10039_));
  INV_X1     g09037(.I(new_n10036_), .ZN(new_n10040_));
  NOR2_X1    g09038(.A1(new_n10040_), .A2(new_n10037_), .ZN(new_n10041_));
  NOR2_X1    g09039(.A1(new_n10039_), .A2(new_n10041_), .ZN(new_n10042_));
  AOI21_X1   g09040(.A1(new_n10035_), .A2(new_n9789_), .B(new_n10042_), .ZN(new_n10043_));
  NOR2_X1    g09041(.A1(new_n9792_), .A2(new_n9751_), .ZN(new_n10044_));
  NAND2_X1   g09042(.A1(new_n10040_), .A2(new_n10037_), .ZN(new_n10045_));
  NAND2_X1   g09043(.A1(new_n10038_), .A2(new_n10036_), .ZN(new_n10046_));
  NAND2_X1   g09044(.A1(new_n10046_), .A2(new_n10045_), .ZN(new_n10047_));
  NOR3_X1    g09045(.A1(new_n10044_), .A2(new_n10047_), .A3(new_n9793_), .ZN(new_n10048_));
  OAI22_X1   g09046(.A1(new_n10043_), .A2(new_n10048_), .B1(new_n10029_), .B2(new_n10034_), .ZN(new_n10049_));
  OAI21_X1   g09047(.A1(new_n9835_), .A2(new_n10030_), .B(new_n10033_), .ZN(new_n10050_));
  INV_X1     g09048(.I(new_n10034_), .ZN(new_n10051_));
  OAI21_X1   g09049(.A1(new_n10044_), .A2(new_n9793_), .B(new_n10047_), .ZN(new_n10052_));
  NAND3_X1   g09050(.A1(new_n10035_), .A2(new_n10042_), .A3(new_n9789_), .ZN(new_n10053_));
  NAND4_X1   g09051(.A1(new_n10051_), .A2(new_n10050_), .A3(new_n10052_), .A4(new_n10053_), .ZN(new_n10054_));
  NAND3_X1   g09052(.A1(new_n10054_), .A2(new_n10018_), .A3(new_n10049_), .ZN(new_n10055_));
  AOI21_X1   g09053(.A1(new_n9844_), .A2(new_n9845_), .B(new_n9842_), .ZN(new_n10056_));
  AOI22_X1   g09054(.A1(new_n10051_), .A2(new_n10050_), .B1(new_n10052_), .B2(new_n10053_), .ZN(new_n10057_));
  NOR4_X1    g09055(.A1(new_n10043_), .A2(new_n10029_), .A3(new_n10048_), .A4(new_n10034_), .ZN(new_n10058_));
  OAI21_X1   g09056(.A1(new_n10057_), .A2(new_n10058_), .B(new_n10056_), .ZN(new_n10059_));
  AOI22_X1   g09057(.A1(new_n10059_), .A2(new_n10055_), .B1(new_n10017_), .B2(new_n10013_), .ZN(new_n10060_));
  NOR3_X1    g09058(.A1(new_n10014_), .A2(new_n10016_), .A3(new_n10015_), .ZN(new_n10061_));
  AOI21_X1   g09059(.A1(new_n10007_), .A2(new_n10012_), .B(new_n9978_), .ZN(new_n10062_));
  NOR3_X1    g09060(.A1(new_n10056_), .A2(new_n10057_), .A3(new_n10058_), .ZN(new_n10063_));
  AOI21_X1   g09061(.A1(new_n10049_), .A2(new_n10054_), .B(new_n10018_), .ZN(new_n10064_));
  NOR4_X1    g09062(.A1(new_n10064_), .A2(new_n10063_), .A3(new_n10062_), .A4(new_n10061_), .ZN(new_n10065_));
  NOR3_X1    g09063(.A1(new_n10060_), .A2(new_n10065_), .A3(new_n9977_), .ZN(new_n10066_));
  OAI21_X1   g09064(.A1(new_n9956_), .A2(new_n9957_), .B(new_n9954_), .ZN(new_n10067_));
  OAI22_X1   g09065(.A1(new_n10064_), .A2(new_n10063_), .B1(new_n10062_), .B2(new_n10061_), .ZN(new_n10068_));
  NAND4_X1   g09066(.A1(new_n10059_), .A2(new_n10017_), .A3(new_n10055_), .A4(new_n10013_), .ZN(new_n10069_));
  AOI21_X1   g09067(.A1(new_n10068_), .A2(new_n10069_), .B(new_n10067_), .ZN(new_n10070_));
  NOR2_X1    g09068(.A1(new_n10066_), .A2(new_n10070_), .ZN(new_n10071_));
  INV_X1     g09069(.I(new_n9748_), .ZN(new_n10072_));
  NOR3_X1    g09070(.A1(new_n9958_), .A2(new_n9957_), .A3(new_n9956_), .ZN(new_n10073_));
  AOI21_X1   g09071(.A1(new_n9949_), .A2(new_n9954_), .B(new_n9749_), .ZN(new_n10074_));
  NOR2_X1    g09072(.A1(new_n10073_), .A2(new_n10074_), .ZN(new_n10075_));
  AOI21_X1   g09073(.A1(new_n8073_), .A2(new_n9967_), .B(new_n8243_), .ZN(new_n10076_));
  NOR3_X1    g09074(.A1(new_n9964_), .A2(new_n8074_), .A3(new_n9965_), .ZN(new_n10077_));
  NOR3_X1    g09075(.A1(new_n9742_), .A2(new_n9747_), .A3(new_n9736_), .ZN(new_n10078_));
  NOR3_X1    g09076(.A1(new_n10077_), .A2(new_n10076_), .A3(new_n10078_), .ZN(new_n10079_));
  NOR3_X1    g09077(.A1(new_n10075_), .A2(new_n10079_), .A3(new_n10072_), .ZN(new_n10080_));
  OAI21_X1   g09078(.A1(new_n8504_), .A2(new_n8746_), .B(new_n8745_), .ZN(new_n10081_));
  NAND3_X1   g09079(.A1(new_n8503_), .A2(new_n8658_), .A3(new_n8244_), .ZN(new_n10082_));
  AOI21_X1   g09080(.A1(new_n10081_), .A2(new_n10082_), .B(new_n10080_), .ZN(new_n10083_));
  NOR3_X1    g09081(.A1(new_n10083_), .A2(new_n9976_), .A3(new_n10071_), .ZN(new_n10084_));
  NAND2_X1   g09082(.A1(new_n8652_), .A2(new_n8750_), .ZN(new_n10085_));
  NAND2_X1   g09083(.A1(new_n8501_), .A2(new_n8341_), .ZN(new_n10086_));
  NAND3_X1   g09084(.A1(new_n8554_), .A2(new_n10086_), .A3(new_n8498_), .ZN(new_n10087_));
  NAND3_X1   g09085(.A1(new_n8651_), .A2(new_n10085_), .A3(new_n10087_), .ZN(new_n10088_));
  NOR2_X1    g09086(.A1(new_n8647_), .A2(new_n8554_), .ZN(new_n10089_));
  NOR2_X1    g09087(.A1(new_n8652_), .A2(new_n8750_), .ZN(new_n10090_));
  OAI21_X1   g09088(.A1(new_n10089_), .A2(new_n10090_), .B(new_n8646_), .ZN(new_n10091_));
  AOI21_X1   g09089(.A1(new_n10088_), .A2(new_n10091_), .B(new_n8747_), .ZN(new_n10092_));
  NOR3_X1    g09090(.A1(new_n8646_), .A2(new_n10090_), .A3(new_n10089_), .ZN(new_n10093_));
  AOI21_X1   g09091(.A1(new_n10085_), .A2(new_n10087_), .B(new_n8651_), .ZN(new_n10094_));
  NOR3_X1    g09092(.A1(new_n8505_), .A2(new_n10093_), .A3(new_n10094_), .ZN(new_n10095_));
  NOR2_X1    g09093(.A1(new_n10092_), .A2(new_n10095_), .ZN(new_n10096_));
  OAI21_X1   g09094(.A1(new_n10083_), .A2(new_n9976_), .B(new_n10071_), .ZN(new_n10097_));
  OAI21_X1   g09095(.A1(new_n10084_), .A2(new_n10096_), .B(new_n10097_), .ZN(new_n10098_));
  AOI21_X1   g09096(.A1(new_n10067_), .A2(new_n10068_), .B(new_n10065_), .ZN(new_n10099_));
  AOI21_X1   g09097(.A1(new_n10035_), .A2(new_n9789_), .B(new_n10039_), .ZN(new_n10100_));
  NAND2_X1   g09098(.A1(new_n10100_), .A2(new_n10046_), .ZN(new_n10101_));
  OAI21_X1   g09099(.A1(new_n10029_), .A2(new_n10034_), .B(new_n10101_), .ZN(new_n10102_));
  NOR3_X1    g09100(.A1(new_n10042_), .A2(new_n10044_), .A3(new_n9793_), .ZN(new_n10103_));
  OAI22_X1   g09101(.A1(new_n10102_), .A2(new_n10103_), .B1(new_n10018_), .B2(new_n10058_), .ZN(new_n10104_));
  NOR2_X1    g09102(.A1(new_n10030_), .A2(new_n9835_), .ZN(new_n10105_));
  OAI21_X1   g09103(.A1(new_n10105_), .A2(new_n10023_), .B(new_n10032_), .ZN(new_n10106_));
  NOR2_X1    g09104(.A1(new_n10100_), .A2(new_n10041_), .ZN(new_n10107_));
  XNOR2_X1   g09105(.A1(new_n10107_), .A2(new_n10106_), .ZN(new_n10108_));
  NAND2_X1   g09106(.A1(new_n10104_), .A2(new_n10108_), .ZN(new_n10109_));
  NOR2_X1    g09107(.A1(new_n10018_), .A2(new_n10058_), .ZN(new_n10110_));
  NOR2_X1    g09108(.A1(new_n10029_), .A2(new_n10034_), .ZN(new_n10111_));
  INV_X1     g09109(.I(new_n10101_), .ZN(new_n10112_));
  NOR3_X1    g09110(.A1(new_n10112_), .A2(new_n10111_), .A3(new_n10103_), .ZN(new_n10113_));
  NOR2_X1    g09111(.A1(new_n10110_), .A2(new_n10113_), .ZN(new_n10114_));
  INV_X1     g09112(.I(new_n10108_), .ZN(new_n10115_));
  NAND2_X1   g09113(.A1(new_n10115_), .A2(new_n10114_), .ZN(new_n10116_));
  NAND2_X1   g09114(.A1(new_n10014_), .A2(new_n10012_), .ZN(new_n10117_));
  NAND2_X1   g09115(.A1(new_n10009_), .A2(new_n10008_), .ZN(new_n10118_));
  NAND3_X1   g09116(.A1(new_n9999_), .A2(new_n10000_), .A3(new_n10004_), .ZN(new_n10119_));
  NAND2_X1   g09117(.A1(new_n9993_), .A2(new_n10005_), .ZN(new_n10120_));
  NAND3_X1   g09118(.A1(new_n10118_), .A2(new_n10119_), .A3(new_n10120_), .ZN(new_n10121_));
  NAND2_X1   g09119(.A1(new_n10117_), .A2(new_n10121_), .ZN(new_n10122_));
  OAI21_X1   g09120(.A1(new_n9979_), .A2(new_n9936_), .B(new_n9984_), .ZN(new_n10123_));
  NAND2_X1   g09121(.A1(new_n10123_), .A2(new_n9988_), .ZN(new_n10124_));
  NAND2_X1   g09122(.A1(new_n9999_), .A2(new_n10000_), .ZN(new_n10125_));
  NAND2_X1   g09123(.A1(new_n10125_), .A2(new_n10004_), .ZN(new_n10126_));
  XOR2_X1    g09124(.A1(new_n10126_), .A2(new_n10124_), .Z(new_n10127_));
  NAND2_X1   g09125(.A1(new_n10122_), .A2(new_n10127_), .ZN(new_n10128_));
  XNOR2_X1   g09126(.A1(new_n10126_), .A2(new_n10124_), .ZN(new_n10129_));
  NAND3_X1   g09127(.A1(new_n10129_), .A2(new_n10117_), .A3(new_n10121_), .ZN(new_n10130_));
  NAND4_X1   g09128(.A1(new_n10116_), .A2(new_n10109_), .A3(new_n10128_), .A4(new_n10130_), .ZN(new_n10131_));
  NOR2_X1    g09129(.A1(new_n10115_), .A2(new_n10114_), .ZN(new_n10132_));
  NOR2_X1    g09130(.A1(new_n10104_), .A2(new_n10108_), .ZN(new_n10133_));
  AOI21_X1   g09131(.A1(new_n10117_), .A2(new_n10121_), .B(new_n10129_), .ZN(new_n10134_));
  INV_X1     g09132(.I(new_n10130_), .ZN(new_n10135_));
  OAI22_X1   g09133(.A1(new_n10132_), .A2(new_n10133_), .B1(new_n10135_), .B2(new_n10134_), .ZN(new_n10136_));
  NAND2_X1   g09134(.A1(new_n10136_), .A2(new_n10131_), .ZN(new_n10137_));
  XOR2_X1    g09135(.A1(new_n10137_), .A2(new_n10099_), .Z(new_n10138_));
  NOR2_X1    g09136(.A1(new_n10098_), .A2(new_n10138_), .ZN(new_n10139_));
  OAI21_X1   g09137(.A1(new_n10072_), .A2(new_n10079_), .B(new_n10075_), .ZN(new_n10140_));
  NAND3_X1   g09138(.A1(new_n10068_), .A2(new_n10069_), .A3(new_n10067_), .ZN(new_n10141_));
  OAI21_X1   g09139(.A1(new_n10060_), .A2(new_n10065_), .B(new_n9977_), .ZN(new_n10142_));
  NAND2_X1   g09140(.A1(new_n10142_), .A2(new_n10141_), .ZN(new_n10143_));
  NAND3_X1   g09141(.A1(new_n9960_), .A2(new_n9975_), .A3(new_n9748_), .ZN(new_n10144_));
  AOI21_X1   g09142(.A1(new_n8503_), .A2(new_n8658_), .B(new_n8244_), .ZN(new_n10145_));
  NOR3_X1    g09143(.A1(new_n8504_), .A2(new_n8746_), .A3(new_n8745_), .ZN(new_n10146_));
  OAI21_X1   g09144(.A1(new_n10146_), .A2(new_n10145_), .B(new_n10144_), .ZN(new_n10147_));
  NAND3_X1   g09145(.A1(new_n10147_), .A2(new_n10140_), .A3(new_n10143_), .ZN(new_n10148_));
  OAI21_X1   g09146(.A1(new_n10093_), .A2(new_n10094_), .B(new_n8505_), .ZN(new_n10149_));
  NAND3_X1   g09147(.A1(new_n10091_), .A2(new_n8747_), .A3(new_n10088_), .ZN(new_n10150_));
  NAND2_X1   g09148(.A1(new_n10149_), .A2(new_n10150_), .ZN(new_n10151_));
  NAND2_X1   g09149(.A1(new_n10151_), .A2(new_n10148_), .ZN(new_n10152_));
  INV_X1     g09150(.I(new_n10099_), .ZN(new_n10153_));
  XOR2_X1    g09151(.A1(new_n10137_), .A2(new_n10153_), .Z(new_n10154_));
  AOI21_X1   g09152(.A1(new_n10152_), .A2(new_n10097_), .B(new_n10154_), .ZN(new_n10155_));
  OAI21_X1   g09153(.A1(new_n10139_), .A2(new_n10155_), .B(new_n8760_), .ZN(new_n10156_));
  NAND2_X1   g09154(.A1(new_n8758_), .A2(new_n8755_), .ZN(new_n10157_));
  NAND3_X1   g09155(.A1(new_n8661_), .A2(new_n8756_), .A3(new_n8757_), .ZN(new_n10158_));
  NAND2_X1   g09156(.A1(new_n10157_), .A2(new_n10158_), .ZN(new_n10159_));
  NAND3_X1   g09157(.A1(new_n10152_), .A2(new_n10097_), .A3(new_n10154_), .ZN(new_n10160_));
  NAND2_X1   g09158(.A1(new_n10081_), .A2(new_n10082_), .ZN(new_n10161_));
  AOI21_X1   g09159(.A1(new_n10161_), .A2(new_n10144_), .B(new_n9976_), .ZN(new_n10162_));
  AOI22_X1   g09160(.A1(new_n10162_), .A2(new_n10143_), .B1(new_n10149_), .B2(new_n10150_), .ZN(new_n10163_));
  AOI21_X1   g09161(.A1(new_n10147_), .A2(new_n10140_), .B(new_n10143_), .ZN(new_n10164_));
  OAI21_X1   g09162(.A1(new_n10163_), .A2(new_n10164_), .B(new_n10138_), .ZN(new_n10165_));
  NAND3_X1   g09163(.A1(new_n10165_), .A2(new_n10160_), .A3(new_n10159_), .ZN(new_n10166_));
  NAND2_X1   g09164(.A1(new_n10156_), .A2(new_n10166_), .ZN(new_n10167_));
  NAND2_X1   g09165(.A1(new_n10167_), .A2(new_n6844_), .ZN(new_n10168_));
  NAND3_X1   g09166(.A1(new_n6832_), .A2(new_n6124_), .A3(new_n5193_), .ZN(new_n10169_));
  OAI21_X1   g09167(.A1(new_n6831_), .A2(new_n6125_), .B(new_n5194_), .ZN(new_n10170_));
  NAND2_X1   g09168(.A1(new_n10170_), .A2(new_n10169_), .ZN(new_n10171_));
  NAND2_X1   g09169(.A1(new_n10140_), .A2(new_n10144_), .ZN(new_n10172_));
  AOI21_X1   g09170(.A1(new_n8503_), .A2(new_n8658_), .B(new_n8745_), .ZN(new_n10173_));
  NOR3_X1    g09171(.A1(new_n8504_), .A2(new_n8746_), .A3(new_n8244_), .ZN(new_n10174_));
  NOR2_X1    g09172(.A1(new_n10174_), .A2(new_n10173_), .ZN(new_n10175_));
  NOR2_X1    g09173(.A1(new_n10172_), .A2(new_n10175_), .ZN(new_n10176_));
  NOR2_X1    g09174(.A1(new_n9976_), .A2(new_n10080_), .ZN(new_n10177_));
  OAI21_X1   g09175(.A1(new_n8504_), .A2(new_n8746_), .B(new_n8244_), .ZN(new_n10178_));
  NAND3_X1   g09176(.A1(new_n8503_), .A2(new_n8658_), .A3(new_n8745_), .ZN(new_n10179_));
  NAND2_X1   g09177(.A1(new_n10178_), .A2(new_n10179_), .ZN(new_n10180_));
  NOR2_X1    g09178(.A1(new_n10177_), .A2(new_n10180_), .ZN(new_n10181_));
  NOR2_X1    g09179(.A1(new_n10176_), .A2(new_n10181_), .ZN(new_n10182_));
  NOR2_X1    g09180(.A1(new_n10171_), .A2(new_n10182_), .ZN(new_n10183_));
  NOR2_X1    g09181(.A1(new_n10077_), .A2(new_n10076_), .ZN(new_n10184_));
  NAND2_X1   g09182(.A1(new_n9748_), .A2(new_n9974_), .ZN(new_n10185_));
  XOR2_X1    g09183(.A1(new_n10184_), .A2(new_n10185_), .Z(new_n10186_));
  INV_X1     g09184(.I(new_n10186_), .ZN(new_n10187_));
  NAND2_X1   g09185(.A1(new_n4368_), .A2(new_n4369_), .ZN(new_n10188_));
  OAI21_X1   g09186(.A1(new_n2698_), .A2(new_n4370_), .B(new_n10188_), .ZN(new_n10189_));
  NAND2_X1   g09187(.A1(new_n4372_), .A2(new_n10189_), .ZN(new_n10190_));
  AND2_X2    g09188(.A1(new_n9972_), .A2(new_n9743_), .Z(new_n10191_));
  NOR3_X1    g09189(.A1(new_n10190_), .A2(new_n9973_), .A3(new_n10191_), .ZN(new_n10192_));
  NAND3_X1   g09190(.A1(new_n3085_), .A2(new_n3086_), .A3(new_n3087_), .ZN(new_n10193_));
  OAI21_X1   g09191(.A1(new_n3081_), .A2(new_n3076_), .B(new_n2065_), .ZN(new_n10194_));
  NAND2_X1   g09192(.A1(new_n10193_), .A2(new_n10194_), .ZN(new_n10195_));
  INV_X1     g09193(.I(new_n4372_), .ZN(new_n10196_));
  AOI21_X1   g09194(.A1(new_n5188_), .A2(new_n5189_), .B(new_n5187_), .ZN(new_n10197_));
  NOR3_X1    g09195(.A1(new_n5180_), .A2(new_n5183_), .A3(new_n4771_), .ZN(new_n10198_));
  OAI21_X1   g09196(.A1(new_n10197_), .A2(new_n10198_), .B(new_n10196_), .ZN(new_n10199_));
  AOI21_X1   g09197(.A1(new_n10199_), .A2(new_n5192_), .B(new_n10195_), .ZN(new_n10200_));
  NOR3_X1    g09198(.A1(new_n10197_), .A2(new_n10198_), .A3(new_n10196_), .ZN(new_n10201_));
  NOR3_X1    g09199(.A1(new_n3089_), .A2(new_n10201_), .A3(new_n5191_), .ZN(new_n10202_));
  OAI21_X1   g09200(.A1(new_n10202_), .A2(new_n10200_), .B(new_n10192_), .ZN(new_n10203_));
  NOR3_X1    g09201(.A1(new_n10202_), .A2(new_n10200_), .A3(new_n10192_), .ZN(new_n10204_));
  AOI21_X1   g09202(.A1(new_n10187_), .A2(new_n10203_), .B(new_n10204_), .ZN(new_n10205_));
  AOI21_X1   g09203(.A1(new_n10171_), .A2(new_n10182_), .B(new_n10205_), .ZN(new_n10206_));
  NOR2_X1    g09204(.A1(new_n10206_), .A2(new_n10183_), .ZN(new_n10207_));
  NAND3_X1   g09205(.A1(new_n6524_), .A2(new_n6838_), .A3(new_n6126_), .ZN(new_n10208_));
  OAI21_X1   g09206(.A1(new_n6523_), .A2(new_n6839_), .B(new_n6833_), .ZN(new_n10209_));
  NAND2_X1   g09207(.A1(new_n10143_), .A2(new_n8747_), .ZN(new_n10210_));
  NAND2_X1   g09208(.A1(new_n10071_), .A2(new_n8505_), .ZN(new_n10211_));
  NAND2_X1   g09209(.A1(new_n10211_), .A2(new_n10210_), .ZN(new_n10212_));
  NOR2_X1    g09210(.A1(new_n10093_), .A2(new_n10094_), .ZN(new_n10213_));
  NOR3_X1    g09211(.A1(new_n10083_), .A2(new_n9976_), .A3(new_n10213_), .ZN(new_n10214_));
  NAND2_X1   g09212(.A1(new_n10091_), .A2(new_n10088_), .ZN(new_n10215_));
  AOI21_X1   g09213(.A1(new_n10147_), .A2(new_n10140_), .B(new_n10215_), .ZN(new_n10216_));
  OAI21_X1   g09214(.A1(new_n10214_), .A2(new_n10216_), .B(new_n10212_), .ZN(new_n10217_));
  NOR2_X1    g09215(.A1(new_n10071_), .A2(new_n8505_), .ZN(new_n10218_));
  NOR2_X1    g09216(.A1(new_n8746_), .A2(new_n8745_), .ZN(new_n10219_));
  NOR4_X1    g09217(.A1(new_n10219_), .A2(new_n8504_), .A3(new_n10066_), .A4(new_n10070_), .ZN(new_n10220_));
  NOR2_X1    g09218(.A1(new_n10218_), .A2(new_n10220_), .ZN(new_n10221_));
  NAND3_X1   g09219(.A1(new_n10147_), .A2(new_n10215_), .A3(new_n10140_), .ZN(new_n10222_));
  OAI21_X1   g09220(.A1(new_n10083_), .A2(new_n9976_), .B(new_n10213_), .ZN(new_n10223_));
  NAND3_X1   g09221(.A1(new_n10223_), .A2(new_n10222_), .A3(new_n10221_), .ZN(new_n10224_));
  NAND4_X1   g09222(.A1(new_n10209_), .A2(new_n10208_), .A3(new_n10217_), .A4(new_n10224_), .ZN(new_n10225_));
  AOI22_X1   g09223(.A1(new_n10209_), .A2(new_n10208_), .B1(new_n10217_), .B2(new_n10224_), .ZN(new_n10226_));
  OAI21_X1   g09224(.A1(new_n10207_), .A2(new_n10226_), .B(new_n10225_), .ZN(new_n10227_));
  OAI21_X1   g09225(.A1(new_n10167_), .A2(new_n6844_), .B(new_n10227_), .ZN(new_n10228_));
  NAND2_X1   g09226(.A1(new_n10228_), .A2(new_n10168_), .ZN(new_n10229_));
  AOI21_X1   g09227(.A1(new_n6840_), .A2(new_n6842_), .B(new_n6820_), .ZN(new_n10230_));
  AOI21_X1   g09228(.A1(new_n6816_), .A2(new_n6818_), .B(new_n6809_), .ZN(new_n10231_));
  NOR2_X1    g09229(.A1(new_n6703_), .A2(new_n6691_), .ZN(new_n10232_));
  NOR2_X1    g09230(.A1(new_n6698_), .A2(new_n6696_), .ZN(new_n10233_));
  NOR2_X1    g09231(.A1(new_n6699_), .A2(new_n6694_), .ZN(new_n10234_));
  NOR3_X1    g09232(.A1(new_n10232_), .A2(new_n10233_), .A3(new_n10234_), .ZN(new_n10235_));
  NOR3_X1    g09233(.A1(new_n6703_), .A2(new_n6691_), .A3(new_n6701_), .ZN(new_n10236_));
  NOR3_X1    g09234(.A1(new_n10235_), .A2(new_n6728_), .A3(new_n10236_), .ZN(new_n10237_));
  AOI21_X1   g09235(.A1(new_n6738_), .A2(new_n6729_), .B(new_n10237_), .ZN(new_n10238_));
  NAND2_X1   g09236(.A1(new_n6726_), .A2(new_n6255_), .ZN(new_n10239_));
  NOR2_X1    g09237(.A1(new_n6710_), .A2(new_n6716_), .ZN(new_n10240_));
  NAND2_X1   g09238(.A1(new_n6710_), .A2(new_n6716_), .ZN(new_n10241_));
  AOI21_X1   g09239(.A1(new_n10239_), .A2(new_n10241_), .B(new_n10240_), .ZN(new_n10242_));
  INV_X1     g09240(.I(new_n10233_), .ZN(new_n10243_));
  OAI21_X1   g09241(.A1(new_n10232_), .A2(new_n10234_), .B(new_n10243_), .ZN(new_n10244_));
  XNOR2_X1   g09242(.A1(new_n10244_), .A2(new_n10242_), .ZN(new_n10245_));
  NOR2_X1    g09243(.A1(new_n10238_), .A2(new_n10245_), .ZN(new_n10246_));
  NAND2_X1   g09244(.A1(new_n6738_), .A2(new_n6729_), .ZN(new_n10247_));
  INV_X1     g09245(.I(new_n10237_), .ZN(new_n10248_));
  NAND2_X1   g09246(.A1(new_n10247_), .A2(new_n10248_), .ZN(new_n10249_));
  XOR2_X1    g09247(.A1(new_n10244_), .A2(new_n10242_), .Z(new_n10250_));
  NOR2_X1    g09248(.A1(new_n10249_), .A2(new_n10250_), .ZN(new_n10251_));
  NAND2_X1   g09249(.A1(new_n6796_), .A2(new_n6802_), .ZN(new_n10252_));
  NAND2_X1   g09250(.A1(new_n6744_), .A2(new_n6757_), .ZN(new_n10253_));
  NOR2_X1    g09251(.A1(new_n6771_), .A2(new_n6764_), .ZN(new_n10254_));
  INV_X1     g09252(.I(new_n10254_), .ZN(new_n10255_));
  NAND2_X1   g09253(.A1(new_n6771_), .A2(new_n6764_), .ZN(new_n10256_));
  NAND3_X1   g09254(.A1(new_n10253_), .A2(new_n10255_), .A3(new_n10256_), .ZN(new_n10257_));
  NAND3_X1   g09255(.A1(new_n6744_), .A2(new_n6757_), .A3(new_n6773_), .ZN(new_n10258_));
  NAND3_X1   g09256(.A1(new_n6805_), .A2(new_n10257_), .A3(new_n10258_), .ZN(new_n10259_));
  NOR2_X1    g09257(.A1(new_n6789_), .A2(new_n6782_), .ZN(new_n10260_));
  AOI22_X1   g09258(.A1(new_n6793_), .A2(new_n6166_), .B1(new_n6789_), .B2(new_n6782_), .ZN(new_n10261_));
  NOR2_X1    g09259(.A1(new_n10261_), .A2(new_n10260_), .ZN(new_n10262_));
  AOI21_X1   g09260(.A1(new_n10253_), .A2(new_n10256_), .B(new_n10254_), .ZN(new_n10263_));
  XOR2_X1    g09261(.A1(new_n10262_), .A2(new_n10263_), .Z(new_n10264_));
  AOI21_X1   g09262(.A1(new_n10252_), .A2(new_n10259_), .B(new_n10264_), .ZN(new_n10265_));
  OAI21_X1   g09263(.A1(new_n6742_), .A2(new_n6806_), .B(new_n10259_), .ZN(new_n10266_));
  XNOR2_X1   g09264(.A1(new_n10262_), .A2(new_n10263_), .ZN(new_n10267_));
  NOR2_X1    g09265(.A1(new_n10267_), .A2(new_n10266_), .ZN(new_n10268_));
  NOR4_X1    g09266(.A1(new_n10251_), .A2(new_n10265_), .A3(new_n10268_), .A4(new_n10246_), .ZN(new_n10269_));
  NAND2_X1   g09267(.A1(new_n10249_), .A2(new_n10250_), .ZN(new_n10270_));
  NAND2_X1   g09268(.A1(new_n10238_), .A2(new_n10245_), .ZN(new_n10271_));
  NAND2_X1   g09269(.A1(new_n10267_), .A2(new_n10266_), .ZN(new_n10272_));
  NAND3_X1   g09270(.A1(new_n10264_), .A2(new_n10252_), .A3(new_n10259_), .ZN(new_n10273_));
  AOI22_X1   g09271(.A1(new_n10270_), .A2(new_n10271_), .B1(new_n10272_), .B2(new_n10273_), .ZN(new_n10274_));
  NOR3_X1    g09272(.A1(new_n10269_), .A2(new_n10231_), .A3(new_n10274_), .ZN(new_n10275_));
  OAI21_X1   g09273(.A1(new_n6674_), .A2(new_n6814_), .B(new_n6817_), .ZN(new_n10276_));
  NAND4_X1   g09274(.A1(new_n10270_), .A2(new_n10272_), .A3(new_n10273_), .A4(new_n10271_), .ZN(new_n10277_));
  OAI22_X1   g09275(.A1(new_n10246_), .A2(new_n10251_), .B1(new_n10265_), .B2(new_n10268_), .ZN(new_n10278_));
  AOI21_X1   g09276(.A1(new_n10278_), .A2(new_n10277_), .B(new_n10276_), .ZN(new_n10279_));
  AOI21_X1   g09277(.A1(new_n6670_), .A2(new_n6672_), .B(new_n6663_), .ZN(new_n10280_));
  OAI21_X1   g09278(.A1(new_n6592_), .A2(new_n6527_), .B(new_n6589_), .ZN(new_n10281_));
  OAI21_X1   g09279(.A1(new_n6542_), .A2(new_n6545_), .B(new_n6579_), .ZN(new_n10282_));
  OAI21_X1   g09280(.A1(new_n6568_), .A2(new_n6571_), .B(new_n6584_), .ZN(new_n10283_));
  XNOR2_X1   g09281(.A1(new_n10283_), .A2(new_n10282_), .ZN(new_n10284_));
  NAND2_X1   g09282(.A1(new_n10281_), .A2(new_n10284_), .ZN(new_n10285_));
  AOI21_X1   g09283(.A1(new_n6591_), .A2(new_n6578_), .B(new_n6593_), .ZN(new_n10286_));
  XOR2_X1    g09284(.A1(new_n10283_), .A2(new_n10282_), .Z(new_n10287_));
  NAND2_X1   g09285(.A1(new_n10286_), .A2(new_n10287_), .ZN(new_n10288_));
  NAND2_X1   g09286(.A1(new_n6596_), .A2(new_n6610_), .ZN(new_n10289_));
  NOR2_X1    g09287(.A1(new_n6600_), .A2(new_n6611_), .ZN(new_n10290_));
  NOR2_X1    g09288(.A1(new_n10290_), .A2(new_n6613_), .ZN(new_n10291_));
  INV_X1     g09289(.I(new_n10291_), .ZN(new_n10292_));
  NAND2_X1   g09290(.A1(new_n10290_), .A2(new_n6613_), .ZN(new_n10293_));
  NAND3_X1   g09291(.A1(new_n10289_), .A2(new_n10292_), .A3(new_n10293_), .ZN(new_n10294_));
  NAND3_X1   g09292(.A1(new_n6596_), .A2(new_n6622_), .A3(new_n6610_), .ZN(new_n10295_));
  NAND3_X1   g09293(.A1(new_n6656_), .A2(new_n10294_), .A3(new_n10295_), .ZN(new_n10296_));
  OAI21_X1   g09294(.A1(new_n6595_), .A2(new_n6660_), .B(new_n10296_), .ZN(new_n10297_));
  NAND2_X1   g09295(.A1(new_n6629_), .A2(new_n6633_), .ZN(new_n10298_));
  INV_X1     g09296(.I(new_n10298_), .ZN(new_n10299_));
  AOI22_X1   g09297(.A1(new_n6647_), .A2(new_n6365_), .B1(new_n6639_), .B2(new_n6634_), .ZN(new_n10300_));
  NOR2_X1    g09298(.A1(new_n10300_), .A2(new_n10299_), .ZN(new_n10301_));
  AOI21_X1   g09299(.A1(new_n10289_), .A2(new_n10293_), .B(new_n10291_), .ZN(new_n10302_));
  XNOR2_X1   g09300(.A1(new_n10301_), .A2(new_n10302_), .ZN(new_n10303_));
  NAND2_X1   g09301(.A1(new_n10303_), .A2(new_n10297_), .ZN(new_n10304_));
  NAND2_X1   g09302(.A1(new_n6650_), .A2(new_n6659_), .ZN(new_n10305_));
  XOR2_X1    g09303(.A1(new_n10301_), .A2(new_n10302_), .Z(new_n10306_));
  NAND3_X1   g09304(.A1(new_n10306_), .A2(new_n10305_), .A3(new_n10296_), .ZN(new_n10307_));
  NAND4_X1   g09305(.A1(new_n10304_), .A2(new_n10307_), .A3(new_n10288_), .A4(new_n10285_), .ZN(new_n10308_));
  INV_X1     g09306(.I(new_n10308_), .ZN(new_n10309_));
  AOI22_X1   g09307(.A1(new_n10304_), .A2(new_n10307_), .B1(new_n10288_), .B2(new_n10285_), .ZN(new_n10310_));
  NOR3_X1    g09308(.A1(new_n10309_), .A2(new_n10280_), .A3(new_n10310_), .ZN(new_n10311_));
  OAI21_X1   g09309(.A1(new_n6526_), .A2(new_n6668_), .B(new_n6671_), .ZN(new_n10312_));
  NAND2_X1   g09310(.A1(new_n10288_), .A2(new_n10285_), .ZN(new_n10313_));
  NAND2_X1   g09311(.A1(new_n10304_), .A2(new_n10307_), .ZN(new_n10314_));
  NAND2_X1   g09312(.A1(new_n10314_), .A2(new_n10313_), .ZN(new_n10315_));
  AOI21_X1   g09313(.A1(new_n10315_), .A2(new_n10308_), .B(new_n10312_), .ZN(new_n10316_));
  NOR4_X1    g09314(.A1(new_n10311_), .A2(new_n10275_), .A3(new_n10316_), .A4(new_n10279_), .ZN(new_n10317_));
  NAND3_X1   g09315(.A1(new_n10278_), .A2(new_n10276_), .A3(new_n10277_), .ZN(new_n10318_));
  OAI21_X1   g09316(.A1(new_n10269_), .A2(new_n10274_), .B(new_n10231_), .ZN(new_n10319_));
  NAND3_X1   g09317(.A1(new_n10315_), .A2(new_n10312_), .A3(new_n10308_), .ZN(new_n10320_));
  OAI21_X1   g09318(.A1(new_n10309_), .A2(new_n10310_), .B(new_n10280_), .ZN(new_n10321_));
  AOI22_X1   g09319(.A1(new_n10320_), .A2(new_n10321_), .B1(new_n10319_), .B2(new_n10318_), .ZN(new_n10322_));
  NOR3_X1    g09320(.A1(new_n10230_), .A2(new_n10322_), .A3(new_n10317_), .ZN(new_n10323_));
  OAI21_X1   g09321(.A1(new_n6825_), .A2(new_n6525_), .B(new_n6841_), .ZN(new_n10324_));
  NAND4_X1   g09322(.A1(new_n10321_), .A2(new_n10319_), .A3(new_n10320_), .A4(new_n10318_), .ZN(new_n10325_));
  OAI22_X1   g09323(.A1(new_n10311_), .A2(new_n10316_), .B1(new_n10275_), .B2(new_n10279_), .ZN(new_n10326_));
  AOI21_X1   g09324(.A1(new_n10325_), .A2(new_n10326_), .B(new_n10324_), .ZN(new_n10327_));
  AOI21_X1   g09325(.A1(new_n10148_), .A2(new_n10151_), .B(new_n10164_), .ZN(new_n10328_));
  NAND2_X1   g09326(.A1(new_n8758_), .A2(new_n8661_), .ZN(new_n10329_));
  NAND2_X1   g09327(.A1(new_n8743_), .A2(new_n8755_), .ZN(new_n10330_));
  AOI22_X1   g09328(.A1(new_n10328_), .A2(new_n10154_), .B1(new_n10330_), .B2(new_n10329_), .ZN(new_n10331_));
  NOR2_X1    g09329(.A1(new_n10331_), .A2(new_n10155_), .ZN(new_n10332_));
  NOR4_X1    g09330(.A1(new_n10132_), .A2(new_n10135_), .A3(new_n10133_), .A4(new_n10134_), .ZN(new_n10333_));
  AOI21_X1   g09331(.A1(new_n10136_), .A2(new_n10099_), .B(new_n10333_), .ZN(new_n10334_));
  NAND2_X1   g09332(.A1(new_n10126_), .A2(new_n10124_), .ZN(new_n10335_));
  NAND4_X1   g09333(.A1(new_n10125_), .A2(new_n10123_), .A3(new_n9988_), .A4(new_n10004_), .ZN(new_n10336_));
  NAND2_X1   g09334(.A1(new_n10122_), .A2(new_n10336_), .ZN(new_n10337_));
  NAND2_X1   g09335(.A1(new_n10337_), .A2(new_n10335_), .ZN(new_n10338_));
  INV_X1     g09336(.I(new_n10107_), .ZN(new_n10339_));
  NAND2_X1   g09337(.A1(new_n10339_), .A2(new_n10106_), .ZN(new_n10340_));
  NOR2_X1    g09338(.A1(new_n10339_), .A2(new_n10106_), .ZN(new_n10341_));
  OAI21_X1   g09339(.A1(new_n10114_), .A2(new_n10341_), .B(new_n10340_), .ZN(new_n10342_));
  XNOR2_X1   g09340(.A1(new_n10338_), .A2(new_n10342_), .ZN(new_n10343_));
  XNOR2_X1   g09341(.A1(new_n10343_), .A2(new_n10334_), .ZN(new_n10344_));
  NAND2_X1   g09342(.A1(new_n8677_), .A2(new_n8724_), .ZN(new_n10345_));
  INV_X1     g09343(.I(new_n8729_), .ZN(new_n10346_));
  INV_X1     g09344(.I(new_n8717_), .ZN(new_n10347_));
  NOR2_X1    g09345(.A1(new_n10347_), .A2(new_n8716_), .ZN(new_n10348_));
  INV_X1     g09346(.I(new_n10348_), .ZN(new_n10349_));
  NAND2_X1   g09347(.A1(new_n10347_), .A2(new_n8716_), .ZN(new_n10350_));
  NAND3_X1   g09348(.A1(new_n10346_), .A2(new_n10349_), .A3(new_n10350_), .ZN(new_n10351_));
  NAND2_X1   g09349(.A1(new_n8729_), .A2(new_n8721_), .ZN(new_n10352_));
  NAND3_X1   g09350(.A1(new_n8727_), .A2(new_n10351_), .A3(new_n10352_), .ZN(new_n10353_));
  INV_X1     g09351(.I(new_n10350_), .ZN(new_n10354_));
  OAI21_X1   g09352(.A1(new_n8729_), .A2(new_n10354_), .B(new_n10349_), .ZN(new_n10355_));
  NOR2_X1    g09353(.A1(new_n8690_), .A2(new_n8637_), .ZN(new_n10356_));
  AOI21_X1   g09354(.A1(new_n10356_), .A2(new_n8685_), .B(new_n8684_), .ZN(new_n10357_));
  NAND2_X1   g09355(.A1(new_n10357_), .A2(new_n10355_), .ZN(new_n10358_));
  INV_X1     g09356(.I(new_n10355_), .ZN(new_n10359_));
  NAND3_X1   g09357(.A1(new_n8679_), .A2(new_n8632_), .A3(new_n8685_), .ZN(new_n10360_));
  NAND2_X1   g09358(.A1(new_n10360_), .A2(new_n8693_), .ZN(new_n10361_));
  NAND2_X1   g09359(.A1(new_n10359_), .A2(new_n10361_), .ZN(new_n10362_));
  NAND2_X1   g09360(.A1(new_n10362_), .A2(new_n10358_), .ZN(new_n10363_));
  AOI21_X1   g09361(.A1(new_n10345_), .A2(new_n10353_), .B(new_n10363_), .ZN(new_n10364_));
  OAI21_X1   g09362(.A1(new_n8734_), .A2(new_n8735_), .B(new_n10353_), .ZN(new_n10365_));
  XOR2_X1    g09363(.A1(new_n10357_), .A2(new_n10355_), .Z(new_n10366_));
  NOR2_X1    g09364(.A1(new_n10365_), .A2(new_n10366_), .ZN(new_n10367_));
  INV_X1     g09365(.I(new_n8672_), .ZN(new_n10368_));
  NOR2_X1    g09366(.A1(new_n10368_), .A2(new_n8671_), .ZN(new_n10369_));
  NAND2_X1   g09367(.A1(new_n10368_), .A2(new_n8671_), .ZN(new_n10370_));
  AOI21_X1   g09368(.A1(new_n8670_), .A2(new_n10370_), .B(new_n10369_), .ZN(new_n10371_));
  NOR3_X1    g09369(.A1(new_n10367_), .A2(new_n10364_), .A3(new_n10371_), .ZN(new_n10372_));
  NOR3_X1    g09370(.A1(new_n8738_), .A2(new_n8753_), .A3(new_n8754_), .ZN(new_n10373_));
  INV_X1     g09371(.I(new_n10371_), .ZN(new_n10374_));
  INV_X1     g09372(.I(new_n10352_), .ZN(new_n10375_));
  NOR2_X1    g09373(.A1(new_n8696_), .A2(new_n10375_), .ZN(new_n10376_));
  AOI22_X1   g09374(.A1(new_n8677_), .A2(new_n8724_), .B1(new_n10376_), .B2(new_n10351_), .ZN(new_n10377_));
  NOR2_X1    g09375(.A1(new_n10359_), .A2(new_n10357_), .ZN(new_n10378_));
  NOR2_X1    g09376(.A1(new_n10361_), .A2(new_n10355_), .ZN(new_n10379_));
  NOR3_X1    g09377(.A1(new_n10377_), .A2(new_n10378_), .A3(new_n10379_), .ZN(new_n10380_));
  NOR2_X1    g09378(.A1(new_n10365_), .A2(new_n10363_), .ZN(new_n10381_));
  NOR3_X1    g09379(.A1(new_n10380_), .A2(new_n10381_), .A3(new_n10374_), .ZN(new_n10382_));
  NOR4_X1    g09380(.A1(new_n10373_), .A2(new_n10382_), .A3(new_n10372_), .A4(new_n8742_), .ZN(new_n10383_));
  OAI22_X1   g09381(.A1(new_n8505_), .A2(new_n8554_), .B1(new_n8648_), .B2(new_n8653_), .ZN(new_n10384_));
  NAND3_X1   g09382(.A1(new_n8756_), .A2(new_n10384_), .A3(new_n8660_), .ZN(new_n10385_));
  INV_X1     g09383(.I(new_n10378_), .ZN(new_n10386_));
  INV_X1     g09384(.I(new_n10379_), .ZN(new_n10387_));
  NAND3_X1   g09385(.A1(new_n10365_), .A2(new_n10386_), .A3(new_n10387_), .ZN(new_n10388_));
  NAND2_X1   g09386(.A1(new_n10377_), .A2(new_n10366_), .ZN(new_n10389_));
  NAND3_X1   g09387(.A1(new_n10388_), .A2(new_n10389_), .A3(new_n10371_), .ZN(new_n10390_));
  OAI21_X1   g09388(.A1(new_n10380_), .A2(new_n10381_), .B(new_n10374_), .ZN(new_n10391_));
  AOI22_X1   g09389(.A1(new_n10385_), .A2(new_n8757_), .B1(new_n10391_), .B2(new_n10390_), .ZN(new_n10392_));
  OAI21_X1   g09390(.A1(new_n10392_), .A2(new_n10383_), .B(new_n10344_), .ZN(new_n10393_));
  XOR2_X1    g09391(.A1(new_n10343_), .A2(new_n10334_), .Z(new_n10394_));
  NAND2_X1   g09392(.A1(new_n10365_), .A2(new_n10366_), .ZN(new_n10395_));
  NAND2_X1   g09393(.A1(new_n10377_), .A2(new_n10363_), .ZN(new_n10396_));
  NAND3_X1   g09394(.A1(new_n10396_), .A2(new_n10395_), .A3(new_n10374_), .ZN(new_n10397_));
  NAND4_X1   g09395(.A1(new_n10385_), .A2(new_n10390_), .A3(new_n10397_), .A4(new_n8757_), .ZN(new_n10398_));
  AOI21_X1   g09396(.A1(new_n10388_), .A2(new_n10389_), .B(new_n10371_), .ZN(new_n10399_));
  OAI22_X1   g09397(.A1(new_n10382_), .A2(new_n10399_), .B1(new_n10373_), .B2(new_n8742_), .ZN(new_n10400_));
  NAND3_X1   g09398(.A1(new_n10400_), .A2(new_n10398_), .A3(new_n10394_), .ZN(new_n10401_));
  NAND2_X1   g09399(.A1(new_n10393_), .A2(new_n10401_), .ZN(new_n10402_));
  NOR2_X1    g09400(.A1(new_n10402_), .A2(new_n10332_), .ZN(new_n10403_));
  NOR2_X1    g09401(.A1(new_n8743_), .A2(new_n8755_), .ZN(new_n10404_));
  NOR2_X1    g09402(.A1(new_n8758_), .A2(new_n8661_), .ZN(new_n10405_));
  OAI22_X1   g09403(.A1(new_n10098_), .A2(new_n10138_), .B1(new_n10404_), .B2(new_n10405_), .ZN(new_n10406_));
  NAND2_X1   g09404(.A1(new_n10406_), .A2(new_n10165_), .ZN(new_n10407_));
  AOI21_X1   g09405(.A1(new_n10400_), .A2(new_n10398_), .B(new_n10394_), .ZN(new_n10408_));
  NOR3_X1    g09406(.A1(new_n10392_), .A2(new_n10383_), .A3(new_n10344_), .ZN(new_n10409_));
  NOR2_X1    g09407(.A1(new_n10408_), .A2(new_n10409_), .ZN(new_n10410_));
  NOR2_X1    g09408(.A1(new_n10410_), .A2(new_n10407_), .ZN(new_n10411_));
  OAI22_X1   g09409(.A1(new_n10411_), .A2(new_n10403_), .B1(new_n10323_), .B2(new_n10327_), .ZN(new_n10412_));
  NOR4_X1    g09410(.A1(new_n10411_), .A2(new_n10403_), .A3(new_n10323_), .A4(new_n10327_), .ZN(new_n10413_));
  OAI21_X1   g09411(.A1(new_n10229_), .A2(new_n10413_), .B(new_n10412_), .ZN(new_n10414_));
  OAI21_X1   g09412(.A1(new_n10322_), .A2(new_n10230_), .B(new_n10325_), .ZN(new_n10415_));
  INV_X1     g09413(.I(new_n10242_), .ZN(new_n10416_));
  NAND2_X1   g09414(.A1(new_n10416_), .A2(new_n10244_), .ZN(new_n10417_));
  INV_X1     g09415(.I(new_n10417_), .ZN(new_n10418_));
  NOR2_X1    g09416(.A1(new_n10416_), .A2(new_n10244_), .ZN(new_n10419_));
  NOR3_X1    g09417(.A1(new_n10238_), .A2(new_n10418_), .A3(new_n10419_), .ZN(new_n10420_));
  INV_X1     g09418(.I(new_n10420_), .ZN(new_n10421_));
  OR2_X2     g09419(.A1(new_n10262_), .A2(new_n10263_), .Z(new_n10422_));
  NAND2_X1   g09420(.A1(new_n10262_), .A2(new_n10263_), .ZN(new_n10423_));
  NAND3_X1   g09421(.A1(new_n10266_), .A2(new_n10422_), .A3(new_n10423_), .ZN(new_n10424_));
  NAND3_X1   g09422(.A1(new_n10267_), .A2(new_n10252_), .A3(new_n10259_), .ZN(new_n10425_));
  NAND3_X1   g09423(.A1(new_n10421_), .A2(new_n10424_), .A3(new_n10425_), .ZN(new_n10426_));
  NOR2_X1    g09424(.A1(new_n10249_), .A2(new_n10245_), .ZN(new_n10427_));
  OAI22_X1   g09425(.A1(new_n10426_), .A2(new_n10427_), .B1(new_n10269_), .B2(new_n10276_), .ZN(new_n10428_));
  NAND2_X1   g09426(.A1(new_n10266_), .A2(new_n10423_), .ZN(new_n10429_));
  NAND2_X1   g09427(.A1(new_n10429_), .A2(new_n10422_), .ZN(new_n10430_));
  OAI21_X1   g09428(.A1(new_n10238_), .A2(new_n10419_), .B(new_n10417_), .ZN(new_n10431_));
  XNOR2_X1   g09429(.A1(new_n10430_), .A2(new_n10431_), .ZN(new_n10432_));
  NAND2_X1   g09430(.A1(new_n10428_), .A2(new_n10432_), .ZN(new_n10433_));
  NAND2_X1   g09431(.A1(new_n10425_), .A2(new_n10424_), .ZN(new_n10434_));
  NOR3_X1    g09432(.A1(new_n10434_), .A2(new_n10420_), .A3(new_n10427_), .ZN(new_n10435_));
  AOI21_X1   g09433(.A1(new_n10231_), .A2(new_n10277_), .B(new_n10435_), .ZN(new_n10436_));
  XOR2_X1    g09434(.A1(new_n10430_), .A2(new_n10431_), .Z(new_n10437_));
  NAND2_X1   g09435(.A1(new_n10436_), .A2(new_n10437_), .ZN(new_n10438_));
  NAND2_X1   g09436(.A1(new_n10283_), .A2(new_n10282_), .ZN(new_n10439_));
  OR2_X2     g09437(.A1(new_n10283_), .A2(new_n10282_), .Z(new_n10440_));
  NAND3_X1   g09438(.A1(new_n10281_), .A2(new_n10439_), .A3(new_n10440_), .ZN(new_n10441_));
  OR2_X2     g09439(.A1(new_n10301_), .A2(new_n10302_), .Z(new_n10442_));
  NAND2_X1   g09440(.A1(new_n10301_), .A2(new_n10302_), .ZN(new_n10443_));
  NAND3_X1   g09441(.A1(new_n10297_), .A2(new_n10442_), .A3(new_n10443_), .ZN(new_n10444_));
  NAND3_X1   g09442(.A1(new_n10303_), .A2(new_n10305_), .A3(new_n10296_), .ZN(new_n10445_));
  NAND2_X1   g09443(.A1(new_n10286_), .A2(new_n10284_), .ZN(new_n10446_));
  NAND4_X1   g09444(.A1(new_n10444_), .A2(new_n10445_), .A3(new_n10441_), .A4(new_n10446_), .ZN(new_n10447_));
  OAI21_X1   g09445(.A1(new_n10309_), .A2(new_n10312_), .B(new_n10447_), .ZN(new_n10448_));
  NAND2_X1   g09446(.A1(new_n10297_), .A2(new_n10443_), .ZN(new_n10449_));
  NAND2_X1   g09447(.A1(new_n10449_), .A2(new_n10442_), .ZN(new_n10450_));
  NAND2_X1   g09448(.A1(new_n10281_), .A2(new_n10440_), .ZN(new_n10451_));
  NAND2_X1   g09449(.A1(new_n10451_), .A2(new_n10439_), .ZN(new_n10452_));
  XNOR2_X1   g09450(.A1(new_n10450_), .A2(new_n10452_), .ZN(new_n10453_));
  NAND2_X1   g09451(.A1(new_n10453_), .A2(new_n10448_), .ZN(new_n10454_));
  INV_X1     g09452(.I(new_n10447_), .ZN(new_n10455_));
  AOI21_X1   g09453(.A1(new_n10280_), .A2(new_n10308_), .B(new_n10455_), .ZN(new_n10456_));
  XOR2_X1    g09454(.A1(new_n10450_), .A2(new_n10452_), .Z(new_n10457_));
  NAND2_X1   g09455(.A1(new_n10456_), .A2(new_n10457_), .ZN(new_n10458_));
  NAND4_X1   g09456(.A1(new_n10438_), .A2(new_n10458_), .A3(new_n10433_), .A4(new_n10454_), .ZN(new_n10459_));
  NOR2_X1    g09457(.A1(new_n10436_), .A2(new_n10437_), .ZN(new_n10460_));
  NOR2_X1    g09458(.A1(new_n10428_), .A2(new_n10432_), .ZN(new_n10461_));
  NOR2_X1    g09459(.A1(new_n10456_), .A2(new_n10457_), .ZN(new_n10462_));
  NOR2_X1    g09460(.A1(new_n10453_), .A2(new_n10448_), .ZN(new_n10463_));
  OAI22_X1   g09461(.A1(new_n10460_), .A2(new_n10461_), .B1(new_n10462_), .B2(new_n10463_), .ZN(new_n10464_));
  NAND3_X1   g09462(.A1(new_n10464_), .A2(new_n10415_), .A3(new_n10459_), .ZN(new_n10465_));
  AOI21_X1   g09463(.A1(new_n10464_), .A2(new_n10459_), .B(new_n10415_), .ZN(new_n10466_));
  INV_X1     g09464(.I(new_n10466_), .ZN(new_n10467_));
  NAND2_X1   g09465(.A1(new_n10467_), .A2(new_n10465_), .ZN(new_n10468_));
  NOR2_X1    g09466(.A1(new_n10414_), .A2(new_n10468_), .ZN(new_n10469_));
  NOR3_X1    g09467(.A1(new_n10408_), .A2(new_n10331_), .A3(new_n10155_), .ZN(new_n10470_));
  NOR2_X1    g09468(.A1(new_n10470_), .A2(new_n10409_), .ZN(new_n10471_));
  NAND3_X1   g09469(.A1(new_n10396_), .A2(new_n10395_), .A3(new_n10371_), .ZN(new_n10472_));
  OAI21_X1   g09470(.A1(new_n10373_), .A2(new_n8742_), .B(new_n10472_), .ZN(new_n10473_));
  NOR3_X1    g09471(.A1(new_n10380_), .A2(new_n10381_), .A3(new_n10371_), .ZN(new_n10474_));
  INV_X1     g09472(.I(new_n10474_), .ZN(new_n10475_));
  NAND2_X1   g09473(.A1(new_n10473_), .A2(new_n10475_), .ZN(new_n10476_));
  AOI21_X1   g09474(.A1(new_n10365_), .A2(new_n10387_), .B(new_n10378_), .ZN(new_n10477_));
  INV_X1     g09475(.I(new_n10477_), .ZN(new_n10478_));
  NAND2_X1   g09476(.A1(new_n10338_), .A2(new_n10342_), .ZN(new_n10479_));
  NOR2_X1    g09477(.A1(new_n10338_), .A2(new_n10342_), .ZN(new_n10480_));
  OAI21_X1   g09478(.A1(new_n10334_), .A2(new_n10480_), .B(new_n10479_), .ZN(new_n10481_));
  XOR2_X1    g09479(.A1(new_n10481_), .A2(new_n10478_), .Z(new_n10482_));
  XNOR2_X1   g09480(.A1(new_n10476_), .A2(new_n10482_), .ZN(new_n10483_));
  NOR2_X1    g09481(.A1(new_n10471_), .A2(new_n10483_), .ZN(new_n10484_));
  NAND3_X1   g09482(.A1(new_n10393_), .A2(new_n10406_), .A3(new_n10165_), .ZN(new_n10485_));
  NAND2_X1   g09483(.A1(new_n10485_), .A2(new_n10401_), .ZN(new_n10486_));
  XOR2_X1    g09484(.A1(new_n10476_), .A2(new_n10482_), .Z(new_n10487_));
  NOR2_X1    g09485(.A1(new_n10486_), .A2(new_n10487_), .ZN(new_n10488_));
  NOR2_X1    g09486(.A1(new_n10484_), .A2(new_n10488_), .ZN(new_n10489_));
  AOI21_X1   g09487(.A1(new_n10414_), .A2(new_n10468_), .B(new_n10489_), .ZN(new_n10490_));
  AOI21_X1   g09488(.A1(new_n10324_), .A2(new_n10326_), .B(new_n10317_), .ZN(new_n10491_));
  NAND2_X1   g09489(.A1(new_n10491_), .A2(new_n10459_), .ZN(new_n10492_));
  NAND2_X1   g09490(.A1(new_n10430_), .A2(new_n10431_), .ZN(new_n10493_));
  NOR2_X1    g09491(.A1(new_n10430_), .A2(new_n10431_), .ZN(new_n10494_));
  INV_X1     g09492(.I(new_n10494_), .ZN(new_n10495_));
  NAND3_X1   g09493(.A1(new_n10428_), .A2(new_n10493_), .A3(new_n10495_), .ZN(new_n10496_));
  NAND2_X1   g09494(.A1(new_n10450_), .A2(new_n10452_), .ZN(new_n10497_));
  NAND4_X1   g09495(.A1(new_n10449_), .A2(new_n10451_), .A3(new_n10439_), .A4(new_n10442_), .ZN(new_n10498_));
  NAND3_X1   g09496(.A1(new_n10448_), .A2(new_n10497_), .A3(new_n10498_), .ZN(new_n10499_));
  NAND2_X1   g09497(.A1(new_n10456_), .A2(new_n10453_), .ZN(new_n10500_));
  NAND2_X1   g09498(.A1(new_n10436_), .A2(new_n10432_), .ZN(new_n10501_));
  NAND4_X1   g09499(.A1(new_n10501_), .A2(new_n10500_), .A3(new_n10496_), .A4(new_n10499_), .ZN(new_n10502_));
  INV_X1     g09500(.I(new_n10493_), .ZN(new_n10503_));
  AOI21_X1   g09501(.A1(new_n10428_), .A2(new_n10495_), .B(new_n10503_), .ZN(new_n10504_));
  INV_X1     g09502(.I(new_n10497_), .ZN(new_n10505_));
  AOI21_X1   g09503(.A1(new_n10448_), .A2(new_n10498_), .B(new_n10505_), .ZN(new_n10506_));
  XNOR2_X1   g09504(.A1(new_n10504_), .A2(new_n10506_), .ZN(new_n10507_));
  NAND3_X1   g09505(.A1(new_n10492_), .A2(new_n10507_), .A3(new_n10502_), .ZN(new_n10508_));
  AOI21_X1   g09506(.A1(new_n10473_), .A2(new_n10475_), .B(new_n10477_), .ZN(new_n10509_));
  INV_X1     g09507(.I(new_n10481_), .ZN(new_n10510_));
  NOR2_X1    g09508(.A1(new_n10367_), .A2(new_n10364_), .ZN(new_n10511_));
  AOI22_X1   g09509(.A1(new_n10385_), .A2(new_n8757_), .B1(new_n10511_), .B2(new_n10371_), .ZN(new_n10512_));
  OAI21_X1   g09510(.A1(new_n10512_), .A2(new_n10474_), .B(new_n10478_), .ZN(new_n10513_));
  NAND3_X1   g09511(.A1(new_n10473_), .A2(new_n10475_), .A3(new_n10477_), .ZN(new_n10514_));
  NAND2_X1   g09512(.A1(new_n10513_), .A2(new_n10514_), .ZN(new_n10515_));
  AOI22_X1   g09513(.A1(new_n10485_), .A2(new_n10401_), .B1(new_n10510_), .B2(new_n10515_), .ZN(new_n10516_));
  NAND3_X1   g09514(.A1(new_n10513_), .A2(new_n10514_), .A3(new_n10481_), .ZN(new_n10517_));
  INV_X1     g09515(.I(new_n10517_), .ZN(new_n10518_));
  NOR3_X1    g09516(.A1(new_n10516_), .A2(new_n10509_), .A3(new_n10518_), .ZN(new_n10519_));
  NOR3_X1    g09517(.A1(new_n10512_), .A2(new_n10474_), .A3(new_n10478_), .ZN(new_n10520_));
  OAI21_X1   g09518(.A1(new_n10520_), .A2(new_n10509_), .B(new_n10510_), .ZN(new_n10521_));
  OAI21_X1   g09519(.A1(new_n10470_), .A2(new_n10409_), .B(new_n10521_), .ZN(new_n10522_));
  NOR2_X1    g09520(.A1(new_n10522_), .A2(new_n10513_), .ZN(new_n10523_));
  NOR2_X1    g09521(.A1(new_n10519_), .A2(new_n10523_), .ZN(new_n10524_));
  NOR4_X1    g09522(.A1(new_n10460_), .A2(new_n10462_), .A3(new_n10461_), .A4(new_n10463_), .ZN(new_n10525_));
  OAI21_X1   g09523(.A1(new_n10415_), .A2(new_n10525_), .B(new_n10502_), .ZN(new_n10526_));
  XOR2_X1    g09524(.A1(new_n10504_), .A2(new_n10506_), .Z(new_n10527_));
  NAND2_X1   g09525(.A1(new_n10526_), .A2(new_n10527_), .ZN(new_n10528_));
  AOI21_X1   g09526(.A1(new_n10508_), .A2(new_n10528_), .B(new_n10524_), .ZN(new_n10529_));
  NOR3_X1    g09527(.A1(new_n10490_), .A2(new_n10529_), .A3(new_n10469_), .ZN(new_n10530_));
  NOR2_X1    g09528(.A1(new_n10504_), .A2(new_n10506_), .ZN(new_n10531_));
  INV_X1     g09529(.I(new_n10531_), .ZN(new_n10532_));
  NAND2_X1   g09530(.A1(new_n10504_), .A2(new_n10506_), .ZN(new_n10533_));
  NAND3_X1   g09531(.A1(new_n10526_), .A2(new_n10532_), .A3(new_n10533_), .ZN(new_n10534_));
  NAND2_X1   g09532(.A1(new_n10534_), .A2(new_n10508_), .ZN(new_n10535_));
  NAND3_X1   g09533(.A1(new_n10522_), .A2(new_n10513_), .A3(new_n10517_), .ZN(new_n10536_));
  NAND3_X1   g09534(.A1(new_n10486_), .A2(new_n10509_), .A3(new_n10521_), .ZN(new_n10537_));
  NAND2_X1   g09535(.A1(new_n10536_), .A2(new_n10537_), .ZN(new_n10538_));
  NOR2_X1    g09536(.A1(new_n10535_), .A2(new_n10538_), .ZN(new_n10539_));
  NOR2_X1    g09537(.A1(new_n10530_), .A2(new_n10539_), .ZN(new_n10540_));
  NAND2_X1   g09538(.A1(new_n10526_), .A2(new_n10533_), .ZN(new_n10541_));
  AOI21_X1   g09539(.A1(new_n10541_), .A2(new_n10532_), .B(new_n10537_), .ZN(new_n10542_));
  INV_X1     g09540(.I(new_n10542_), .ZN(new_n10543_));
  NAND3_X1   g09541(.A1(new_n10541_), .A2(new_n10532_), .A3(new_n10537_), .ZN(new_n10544_));
  INV_X1     g09542(.I(new_n10544_), .ZN(new_n10545_));
  AOI21_X1   g09543(.A1(new_n10540_), .A2(new_n10543_), .B(new_n10545_), .ZN(new_n10546_));
  INV_X1     g09544(.I(new_n10546_), .ZN(new_n10547_));
  INV_X1     g09545(.I(\A[795] ), .ZN(new_n10548_));
  NOR2_X1    g09546(.A1(new_n10548_), .A2(\A[794] ), .ZN(new_n10549_));
  INV_X1     g09547(.I(\A[794] ), .ZN(new_n10550_));
  NOR2_X1    g09548(.A1(new_n10550_), .A2(\A[795] ), .ZN(new_n10551_));
  OAI21_X1   g09549(.A1(new_n10549_), .A2(new_n10551_), .B(\A[793] ), .ZN(new_n10552_));
  INV_X1     g09550(.I(\A[793] ), .ZN(new_n10553_));
  NAND2_X1   g09551(.A1(\A[794] ), .A2(\A[795] ), .ZN(new_n10554_));
  INV_X1     g09552(.I(new_n10554_), .ZN(new_n10555_));
  NOR2_X1    g09553(.A1(\A[794] ), .A2(\A[795] ), .ZN(new_n10556_));
  OAI21_X1   g09554(.A1(new_n10555_), .A2(new_n10556_), .B(new_n10553_), .ZN(new_n10557_));
  NAND2_X1   g09555(.A1(new_n10552_), .A2(new_n10557_), .ZN(new_n10558_));
  INV_X1     g09556(.I(\A[798] ), .ZN(new_n10559_));
  NOR2_X1    g09557(.A1(new_n10559_), .A2(\A[797] ), .ZN(new_n10560_));
  INV_X1     g09558(.I(\A[797] ), .ZN(new_n10561_));
  NOR2_X1    g09559(.A1(new_n10561_), .A2(\A[798] ), .ZN(new_n10562_));
  OAI21_X1   g09560(.A1(new_n10560_), .A2(new_n10562_), .B(\A[796] ), .ZN(new_n10563_));
  INV_X1     g09561(.I(\A[796] ), .ZN(new_n10564_));
  NAND2_X1   g09562(.A1(\A[797] ), .A2(\A[798] ), .ZN(new_n10565_));
  INV_X1     g09563(.I(new_n10565_), .ZN(new_n10566_));
  NOR2_X1    g09564(.A1(\A[797] ), .A2(\A[798] ), .ZN(new_n10567_));
  OAI21_X1   g09565(.A1(new_n10566_), .A2(new_n10567_), .B(new_n10564_), .ZN(new_n10568_));
  NAND2_X1   g09566(.A1(new_n10563_), .A2(new_n10568_), .ZN(new_n10569_));
  NOR2_X1    g09567(.A1(new_n10558_), .A2(new_n10569_), .ZN(new_n10570_));
  AOI21_X1   g09568(.A1(new_n10553_), .A2(new_n10554_), .B(new_n10556_), .ZN(new_n10571_));
  NAND2_X1   g09569(.A1(new_n10570_), .A2(new_n10571_), .ZN(new_n10572_));
  AOI21_X1   g09570(.A1(new_n10564_), .A2(new_n10565_), .B(new_n10567_), .ZN(new_n10573_));
  OAI21_X1   g09571(.A1(new_n10570_), .A2(new_n10571_), .B(new_n10573_), .ZN(new_n10574_));
  INV_X1     g09572(.I(\A[787] ), .ZN(new_n10575_));
  INV_X1     g09573(.I(\A[788] ), .ZN(new_n10576_));
  NAND2_X1   g09574(.A1(new_n10576_), .A2(\A[789] ), .ZN(new_n10577_));
  INV_X1     g09575(.I(\A[789] ), .ZN(new_n10578_));
  NAND2_X1   g09576(.A1(new_n10578_), .A2(\A[788] ), .ZN(new_n10579_));
  AOI21_X1   g09577(.A1(new_n10577_), .A2(new_n10579_), .B(new_n10575_), .ZN(new_n10580_));
  NAND2_X1   g09578(.A1(\A[788] ), .A2(\A[789] ), .ZN(new_n10581_));
  NOR2_X1    g09579(.A1(\A[788] ), .A2(\A[789] ), .ZN(new_n10582_));
  INV_X1     g09580(.I(new_n10582_), .ZN(new_n10583_));
  AOI21_X1   g09581(.A1(new_n10583_), .A2(new_n10581_), .B(\A[787] ), .ZN(new_n10584_));
  INV_X1     g09582(.I(\A[790] ), .ZN(new_n10585_));
  INV_X1     g09583(.I(\A[791] ), .ZN(new_n10586_));
  NAND2_X1   g09584(.A1(new_n10586_), .A2(\A[792] ), .ZN(new_n10587_));
  INV_X1     g09585(.I(\A[792] ), .ZN(new_n10588_));
  NAND2_X1   g09586(.A1(new_n10588_), .A2(\A[791] ), .ZN(new_n10589_));
  AOI21_X1   g09587(.A1(new_n10587_), .A2(new_n10589_), .B(new_n10585_), .ZN(new_n10590_));
  NAND2_X1   g09588(.A1(\A[791] ), .A2(\A[792] ), .ZN(new_n10591_));
  NOR2_X1    g09589(.A1(\A[791] ), .A2(\A[792] ), .ZN(new_n10592_));
  INV_X1     g09590(.I(new_n10592_), .ZN(new_n10593_));
  AOI21_X1   g09591(.A1(new_n10593_), .A2(new_n10591_), .B(\A[790] ), .ZN(new_n10594_));
  NOR4_X1    g09592(.A1(new_n10580_), .A2(new_n10584_), .A3(new_n10594_), .A4(new_n10590_), .ZN(new_n10595_));
  AOI21_X1   g09593(.A1(new_n10585_), .A2(new_n10591_), .B(new_n10592_), .ZN(new_n10596_));
  AOI21_X1   g09594(.A1(new_n10575_), .A2(new_n10581_), .B(new_n10582_), .ZN(new_n10597_));
  NOR2_X1    g09595(.A1(new_n10596_), .A2(new_n10597_), .ZN(new_n10598_));
  INV_X1     g09596(.I(new_n10598_), .ZN(new_n10599_));
  AND2_X2    g09597(.A1(new_n10596_), .A2(new_n10597_), .Z(new_n10600_));
  OAI21_X1   g09598(.A1(new_n10595_), .A2(new_n10600_), .B(new_n10599_), .ZN(new_n10601_));
  AOI21_X1   g09599(.A1(new_n10574_), .A2(new_n10572_), .B(new_n10601_), .ZN(new_n10602_));
  NOR2_X1    g09600(.A1(new_n10600_), .A2(new_n10598_), .ZN(new_n10603_));
  XOR2_X1    g09601(.A1(new_n10603_), .A2(new_n10595_), .Z(new_n10604_));
  NAND2_X1   g09602(.A1(new_n10550_), .A2(\A[795] ), .ZN(new_n10605_));
  NAND2_X1   g09603(.A1(new_n10548_), .A2(\A[794] ), .ZN(new_n10606_));
  AOI21_X1   g09604(.A1(new_n10605_), .A2(new_n10606_), .B(new_n10553_), .ZN(new_n10607_));
  INV_X1     g09605(.I(new_n10556_), .ZN(new_n10608_));
  AOI21_X1   g09606(.A1(new_n10608_), .A2(new_n10554_), .B(\A[793] ), .ZN(new_n10609_));
  NOR2_X1    g09607(.A1(new_n10609_), .A2(new_n10607_), .ZN(new_n10610_));
  NAND2_X1   g09608(.A1(new_n10561_), .A2(\A[798] ), .ZN(new_n10611_));
  NAND2_X1   g09609(.A1(new_n10559_), .A2(\A[797] ), .ZN(new_n10612_));
  AOI21_X1   g09610(.A1(new_n10611_), .A2(new_n10612_), .B(new_n10564_), .ZN(new_n10613_));
  INV_X1     g09611(.I(new_n10567_), .ZN(new_n10614_));
  AOI21_X1   g09612(.A1(new_n10614_), .A2(new_n10565_), .B(\A[796] ), .ZN(new_n10615_));
  NOR2_X1    g09613(.A1(new_n10615_), .A2(new_n10613_), .ZN(new_n10616_));
  NAND2_X1   g09614(.A1(new_n10610_), .A2(new_n10616_), .ZN(new_n10617_));
  XNOR2_X1   g09615(.A1(new_n10573_), .A2(new_n10571_), .ZN(new_n10618_));
  NOR2_X1    g09616(.A1(new_n10617_), .A2(new_n10618_), .ZN(new_n10619_));
  XOR2_X1    g09617(.A1(new_n10573_), .A2(new_n10571_), .Z(new_n10620_));
  NOR2_X1    g09618(.A1(new_n10570_), .A2(new_n10620_), .ZN(new_n10621_));
  INV_X1     g09619(.I(new_n10595_), .ZN(new_n10622_));
  OAI22_X1   g09620(.A1(new_n10580_), .A2(new_n10584_), .B1(new_n10594_), .B2(new_n10590_), .ZN(new_n10623_));
  NAND2_X1   g09621(.A1(new_n10558_), .A2(new_n10569_), .ZN(new_n10624_));
  NAND4_X1   g09622(.A1(new_n10622_), .A2(new_n10617_), .A3(new_n10624_), .A4(new_n10623_), .ZN(new_n10625_));
  OAI21_X1   g09623(.A1(new_n10619_), .A2(new_n10621_), .B(new_n10625_), .ZN(new_n10626_));
  NAND2_X1   g09624(.A1(new_n10622_), .A2(new_n10623_), .ZN(new_n10627_));
  NOR2_X1    g09625(.A1(new_n10610_), .A2(new_n10616_), .ZN(new_n10628_));
  INV_X1     g09626(.I(new_n10573_), .ZN(new_n10629_));
  INV_X1     g09627(.I(new_n10571_), .ZN(new_n10630_));
  NOR3_X1    g09628(.A1(new_n10628_), .A2(new_n10629_), .A3(new_n10630_), .ZN(new_n10631_));
  NAND3_X1   g09629(.A1(new_n10617_), .A2(new_n10624_), .A3(new_n10620_), .ZN(new_n10632_));
  NOR3_X1    g09630(.A1(new_n10632_), .A2(new_n10631_), .A3(new_n10627_), .ZN(new_n10633_));
  AOI21_X1   g09631(.A1(new_n10626_), .A2(new_n10604_), .B(new_n10633_), .ZN(new_n10634_));
  NAND2_X1   g09632(.A1(new_n10574_), .A2(new_n10572_), .ZN(new_n10635_));
  INV_X1     g09633(.I(new_n10601_), .ZN(new_n10636_));
  NOR2_X1    g09634(.A1(new_n10635_), .A2(new_n10636_), .ZN(new_n10637_));
  NOR2_X1    g09635(.A1(new_n10634_), .A2(new_n10637_), .ZN(new_n10638_));
  NOR2_X1    g09636(.A1(new_n10638_), .A2(new_n10602_), .ZN(new_n10639_));
  INV_X1     g09637(.I(\A[784] ), .ZN(new_n10640_));
  NAND2_X1   g09638(.A1(\A[785] ), .A2(\A[786] ), .ZN(new_n10641_));
  NOR2_X1    g09639(.A1(\A[785] ), .A2(\A[786] ), .ZN(new_n10642_));
  AOI21_X1   g09640(.A1(new_n10640_), .A2(new_n10641_), .B(new_n10642_), .ZN(new_n10643_));
  INV_X1     g09641(.I(\A[781] ), .ZN(new_n10644_));
  INV_X1     g09642(.I(\A[782] ), .ZN(new_n10645_));
  NAND2_X1   g09643(.A1(new_n10645_), .A2(\A[783] ), .ZN(new_n10646_));
  INV_X1     g09644(.I(\A[783] ), .ZN(new_n10647_));
  NAND2_X1   g09645(.A1(new_n10647_), .A2(\A[782] ), .ZN(new_n10648_));
  AOI21_X1   g09646(.A1(new_n10646_), .A2(new_n10648_), .B(new_n10644_), .ZN(new_n10649_));
  NAND2_X1   g09647(.A1(\A[782] ), .A2(\A[783] ), .ZN(new_n10650_));
  NOR2_X1    g09648(.A1(\A[782] ), .A2(\A[783] ), .ZN(new_n10651_));
  INV_X1     g09649(.I(new_n10651_), .ZN(new_n10652_));
  AOI21_X1   g09650(.A1(new_n10652_), .A2(new_n10650_), .B(\A[781] ), .ZN(new_n10653_));
  NOR2_X1    g09651(.A1(new_n10653_), .A2(new_n10649_), .ZN(new_n10654_));
  INV_X1     g09652(.I(\A[785] ), .ZN(new_n10655_));
  NAND2_X1   g09653(.A1(new_n10655_), .A2(\A[786] ), .ZN(new_n10656_));
  INV_X1     g09654(.I(\A[786] ), .ZN(new_n10657_));
  NAND2_X1   g09655(.A1(new_n10657_), .A2(\A[785] ), .ZN(new_n10658_));
  AOI21_X1   g09656(.A1(new_n10656_), .A2(new_n10658_), .B(new_n10640_), .ZN(new_n10659_));
  INV_X1     g09657(.I(new_n10642_), .ZN(new_n10660_));
  AOI21_X1   g09658(.A1(new_n10660_), .A2(new_n10641_), .B(\A[784] ), .ZN(new_n10661_));
  NOR2_X1    g09659(.A1(new_n10661_), .A2(new_n10659_), .ZN(new_n10662_));
  NAND2_X1   g09660(.A1(new_n10654_), .A2(new_n10662_), .ZN(new_n10663_));
  AOI21_X1   g09661(.A1(new_n10644_), .A2(new_n10650_), .B(new_n10651_), .ZN(new_n10664_));
  INV_X1     g09662(.I(new_n10664_), .ZN(new_n10665_));
  NOR2_X1    g09663(.A1(new_n10663_), .A2(new_n10665_), .ZN(new_n10666_));
  NAND2_X1   g09664(.A1(new_n10663_), .A2(new_n10665_), .ZN(new_n10667_));
  AOI21_X1   g09665(.A1(new_n10643_), .A2(new_n10667_), .B(new_n10666_), .ZN(new_n10668_));
  INV_X1     g09666(.I(\A[778] ), .ZN(new_n10669_));
  NAND2_X1   g09667(.A1(\A[779] ), .A2(\A[780] ), .ZN(new_n10670_));
  NOR2_X1    g09668(.A1(\A[779] ), .A2(\A[780] ), .ZN(new_n10671_));
  AOI21_X1   g09669(.A1(new_n10669_), .A2(new_n10670_), .B(new_n10671_), .ZN(new_n10672_));
  INV_X1     g09670(.I(\A[775] ), .ZN(new_n10673_));
  NAND2_X1   g09671(.A1(\A[776] ), .A2(\A[777] ), .ZN(new_n10674_));
  NOR2_X1    g09672(.A1(\A[776] ), .A2(\A[777] ), .ZN(new_n10675_));
  AOI21_X1   g09673(.A1(new_n10673_), .A2(new_n10674_), .B(new_n10675_), .ZN(new_n10676_));
  NOR2_X1    g09674(.A1(new_n10672_), .A2(new_n10676_), .ZN(new_n10677_));
  INV_X1     g09675(.I(\A[776] ), .ZN(new_n10678_));
  NAND2_X1   g09676(.A1(new_n10678_), .A2(\A[777] ), .ZN(new_n10679_));
  INV_X1     g09677(.I(\A[777] ), .ZN(new_n10680_));
  NAND2_X1   g09678(.A1(new_n10680_), .A2(\A[776] ), .ZN(new_n10681_));
  AOI21_X1   g09679(.A1(new_n10679_), .A2(new_n10681_), .B(new_n10673_), .ZN(new_n10682_));
  INV_X1     g09680(.I(new_n10675_), .ZN(new_n10683_));
  AOI21_X1   g09681(.A1(new_n10683_), .A2(new_n10674_), .B(\A[775] ), .ZN(new_n10684_));
  INV_X1     g09682(.I(\A[779] ), .ZN(new_n10685_));
  NAND2_X1   g09683(.A1(new_n10685_), .A2(\A[780] ), .ZN(new_n10686_));
  INV_X1     g09684(.I(\A[780] ), .ZN(new_n10687_));
  NAND2_X1   g09685(.A1(new_n10687_), .A2(\A[779] ), .ZN(new_n10688_));
  AOI21_X1   g09686(.A1(new_n10686_), .A2(new_n10688_), .B(new_n10669_), .ZN(new_n10689_));
  INV_X1     g09687(.I(new_n10671_), .ZN(new_n10690_));
  AOI21_X1   g09688(.A1(new_n10690_), .A2(new_n10670_), .B(\A[778] ), .ZN(new_n10691_));
  NOR4_X1    g09689(.A1(new_n10682_), .A2(new_n10684_), .A3(new_n10691_), .A4(new_n10689_), .ZN(new_n10692_));
  AND2_X2    g09690(.A1(new_n10672_), .A2(new_n10676_), .Z(new_n10693_));
  NOR2_X1    g09691(.A1(new_n10692_), .A2(new_n10693_), .ZN(new_n10694_));
  NOR2_X1    g09692(.A1(new_n10694_), .A2(new_n10677_), .ZN(new_n10695_));
  INV_X1     g09693(.I(new_n10695_), .ZN(new_n10696_));
  NOR2_X1    g09694(.A1(new_n10668_), .A2(new_n10696_), .ZN(new_n10697_));
  NOR2_X1    g09695(.A1(new_n10693_), .A2(new_n10677_), .ZN(new_n10698_));
  XOR2_X1    g09696(.A1(new_n10698_), .A2(new_n10692_), .Z(new_n10699_));
  NOR2_X1    g09697(.A1(new_n10684_), .A2(new_n10682_), .ZN(new_n10700_));
  NOR2_X1    g09698(.A1(new_n10691_), .A2(new_n10689_), .ZN(new_n10701_));
  XNOR2_X1   g09699(.A1(new_n10700_), .A2(new_n10701_), .ZN(new_n10702_));
  NOR2_X1    g09700(.A1(new_n10647_), .A2(\A[782] ), .ZN(new_n10703_));
  NOR2_X1    g09701(.A1(new_n10645_), .A2(\A[783] ), .ZN(new_n10704_));
  OAI21_X1   g09702(.A1(new_n10703_), .A2(new_n10704_), .B(\A[781] ), .ZN(new_n10705_));
  INV_X1     g09703(.I(new_n10650_), .ZN(new_n10706_));
  OAI21_X1   g09704(.A1(new_n10706_), .A2(new_n10651_), .B(new_n10644_), .ZN(new_n10707_));
  NAND2_X1   g09705(.A1(new_n10705_), .A2(new_n10707_), .ZN(new_n10708_));
  NOR2_X1    g09706(.A1(new_n10657_), .A2(\A[785] ), .ZN(new_n10709_));
  NOR2_X1    g09707(.A1(new_n10655_), .A2(\A[786] ), .ZN(new_n10710_));
  OAI21_X1   g09708(.A1(new_n10709_), .A2(new_n10710_), .B(\A[784] ), .ZN(new_n10711_));
  INV_X1     g09709(.I(new_n10641_), .ZN(new_n10712_));
  OAI21_X1   g09710(.A1(new_n10712_), .A2(new_n10642_), .B(new_n10640_), .ZN(new_n10713_));
  NAND2_X1   g09711(.A1(new_n10711_), .A2(new_n10713_), .ZN(new_n10714_));
  NAND2_X1   g09712(.A1(new_n10708_), .A2(new_n10714_), .ZN(new_n10715_));
  NAND2_X1   g09713(.A1(new_n10663_), .A2(new_n10715_), .ZN(new_n10716_));
  XNOR2_X1   g09714(.A1(new_n10643_), .A2(new_n10664_), .ZN(new_n10717_));
  NOR2_X1    g09715(.A1(new_n10663_), .A2(new_n10717_), .ZN(new_n10718_));
  NOR2_X1    g09716(.A1(new_n10708_), .A2(new_n10714_), .ZN(new_n10719_));
  XOR2_X1    g09717(.A1(new_n10643_), .A2(new_n10664_), .Z(new_n10720_));
  NOR2_X1    g09718(.A1(new_n10719_), .A2(new_n10720_), .ZN(new_n10721_));
  OAI22_X1   g09719(.A1(new_n10702_), .A2(new_n10716_), .B1(new_n10718_), .B2(new_n10721_), .ZN(new_n10722_));
  NAND2_X1   g09720(.A1(new_n10722_), .A2(new_n10699_), .ZN(new_n10723_));
  NOR2_X1    g09721(.A1(new_n10700_), .A2(new_n10701_), .ZN(new_n10724_));
  NOR2_X1    g09722(.A1(new_n10724_), .A2(new_n10692_), .ZN(new_n10725_));
  NAND3_X1   g09723(.A1(new_n10715_), .A2(new_n10643_), .A3(new_n10664_), .ZN(new_n10726_));
  NOR2_X1    g09724(.A1(new_n10654_), .A2(new_n10662_), .ZN(new_n10727_));
  NOR3_X1    g09725(.A1(new_n10719_), .A2(new_n10727_), .A3(new_n10717_), .ZN(new_n10728_));
  NAND3_X1   g09726(.A1(new_n10728_), .A2(new_n10726_), .A3(new_n10725_), .ZN(new_n10729_));
  NAND2_X1   g09727(.A1(new_n10719_), .A2(new_n10664_), .ZN(new_n10730_));
  OAI21_X1   g09728(.A1(new_n10719_), .A2(new_n10664_), .B(new_n10643_), .ZN(new_n10731_));
  NAND2_X1   g09729(.A1(new_n10731_), .A2(new_n10730_), .ZN(new_n10732_));
  NOR2_X1    g09730(.A1(new_n10732_), .A2(new_n10695_), .ZN(new_n10733_));
  AOI21_X1   g09731(.A1(new_n10723_), .A2(new_n10729_), .B(new_n10733_), .ZN(new_n10734_));
  NOR2_X1    g09732(.A1(new_n10734_), .A2(new_n10697_), .ZN(new_n10735_));
  NOR2_X1    g09733(.A1(new_n10639_), .A2(new_n10735_), .ZN(new_n10736_));
  INV_X1     g09734(.I(new_n10729_), .ZN(new_n10737_));
  NOR2_X1    g09735(.A1(new_n10727_), .A2(new_n10719_), .ZN(new_n10738_));
  NAND2_X1   g09736(.A1(new_n10719_), .A2(new_n10720_), .ZN(new_n10739_));
  NAND2_X1   g09737(.A1(new_n10663_), .A2(new_n10717_), .ZN(new_n10740_));
  AOI22_X1   g09738(.A1(new_n10725_), .A2(new_n10738_), .B1(new_n10740_), .B2(new_n10739_), .ZN(new_n10741_));
  NAND4_X1   g09739(.A1(new_n10725_), .A2(new_n10663_), .A3(new_n10715_), .A4(new_n10720_), .ZN(new_n10742_));
  INV_X1     g09740(.I(new_n10742_), .ZN(new_n10743_));
  NOR2_X1    g09741(.A1(new_n10743_), .A2(new_n10741_), .ZN(new_n10744_));
  OAI22_X1   g09742(.A1(new_n10744_), .A2(new_n10699_), .B1(new_n10723_), .B2(new_n10737_), .ZN(new_n10745_));
  XNOR2_X1   g09743(.A1(new_n10603_), .A2(new_n10595_), .ZN(new_n10746_));
  OR3_X2     g09744(.A1(new_n10632_), .A2(new_n10631_), .A3(new_n10627_), .Z(new_n10747_));
  AOI21_X1   g09745(.A1(new_n10747_), .A2(new_n10626_), .B(new_n10746_), .ZN(new_n10748_));
  INV_X1     g09746(.I(new_n10623_), .ZN(new_n10749_));
  NOR2_X1    g09747(.A1(new_n10749_), .A2(new_n10595_), .ZN(new_n10750_));
  NOR2_X1    g09748(.A1(new_n10628_), .A2(new_n10570_), .ZN(new_n10751_));
  NAND2_X1   g09749(.A1(new_n10570_), .A2(new_n10620_), .ZN(new_n10752_));
  NAND2_X1   g09750(.A1(new_n10617_), .A2(new_n10618_), .ZN(new_n10753_));
  AOI22_X1   g09751(.A1(new_n10750_), .A2(new_n10751_), .B1(new_n10753_), .B2(new_n10752_), .ZN(new_n10754_));
  NOR3_X1    g09752(.A1(new_n10625_), .A2(new_n10619_), .A3(new_n10621_), .ZN(new_n10755_));
  NOR3_X1    g09753(.A1(new_n10754_), .A2(new_n10755_), .A3(new_n10604_), .ZN(new_n10756_));
  XOR2_X1    g09754(.A1(new_n10716_), .A2(new_n10725_), .Z(new_n10757_));
  NAND2_X1   g09755(.A1(new_n10617_), .A2(new_n10624_), .ZN(new_n10758_));
  NAND2_X1   g09756(.A1(new_n10627_), .A2(new_n10758_), .ZN(new_n10759_));
  NAND2_X1   g09757(.A1(new_n10759_), .A2(new_n10625_), .ZN(new_n10760_));
  NOR2_X1    g09758(.A1(new_n10757_), .A2(new_n10760_), .ZN(new_n10761_));
  OAI21_X1   g09759(.A1(new_n10748_), .A2(new_n10756_), .B(new_n10761_), .ZN(new_n10762_));
  NOR3_X1    g09760(.A1(new_n10761_), .A2(new_n10748_), .A3(new_n10756_), .ZN(new_n10763_));
  AOI21_X1   g09761(.A1(new_n10762_), .A2(new_n10745_), .B(new_n10763_), .ZN(new_n10764_));
  OAI21_X1   g09762(.A1(new_n10754_), .A2(new_n10746_), .B(new_n10747_), .ZN(new_n10765_));
  XOR2_X1    g09763(.A1(new_n10635_), .A2(new_n10601_), .Z(new_n10766_));
  NAND2_X1   g09764(.A1(new_n10765_), .A2(new_n10766_), .ZN(new_n10767_));
  NOR2_X1    g09765(.A1(new_n10637_), .A2(new_n10602_), .ZN(new_n10768_));
  NAND2_X1   g09766(.A1(new_n10634_), .A2(new_n10768_), .ZN(new_n10769_));
  XNOR2_X1   g09767(.A1(new_n10698_), .A2(new_n10692_), .ZN(new_n10770_));
  NOR2_X1    g09768(.A1(new_n10741_), .A2(new_n10770_), .ZN(new_n10771_));
  OAI22_X1   g09769(.A1(new_n10771_), .A2(new_n10737_), .B1(new_n10697_), .B2(new_n10733_), .ZN(new_n10772_));
  NAND2_X1   g09770(.A1(new_n10732_), .A2(new_n10695_), .ZN(new_n10773_));
  NAND2_X1   g09771(.A1(new_n10668_), .A2(new_n10696_), .ZN(new_n10774_));
  NAND4_X1   g09772(.A1(new_n10723_), .A2(new_n10729_), .A3(new_n10773_), .A4(new_n10774_), .ZN(new_n10775_));
  NAND4_X1   g09773(.A1(new_n10767_), .A2(new_n10775_), .A3(new_n10769_), .A4(new_n10772_), .ZN(new_n10776_));
  AOI22_X1   g09774(.A1(new_n10767_), .A2(new_n10769_), .B1(new_n10775_), .B2(new_n10772_), .ZN(new_n10777_));
  AOI21_X1   g09775(.A1(new_n10764_), .A2(new_n10776_), .B(new_n10777_), .ZN(new_n10778_));
  NAND2_X1   g09776(.A1(new_n10639_), .A2(new_n10735_), .ZN(new_n10779_));
  INV_X1     g09777(.I(new_n10779_), .ZN(new_n10780_));
  NOR3_X1    g09778(.A1(new_n10778_), .A2(new_n10736_), .A3(new_n10780_), .ZN(new_n10781_));
  INV_X1     g09779(.I(new_n10781_), .ZN(new_n10782_));
  OAI21_X1   g09780(.A1(new_n10736_), .A2(new_n10780_), .B(new_n10778_), .ZN(new_n10783_));
  NAND2_X1   g09781(.A1(new_n10782_), .A2(new_n10783_), .ZN(new_n10784_));
  INV_X1     g09782(.I(new_n10784_), .ZN(new_n10785_));
  INV_X1     g09783(.I(\A[769] ), .ZN(new_n10786_));
  INV_X1     g09784(.I(\A[770] ), .ZN(new_n10787_));
  NAND2_X1   g09785(.A1(new_n10787_), .A2(\A[771] ), .ZN(new_n10788_));
  INV_X1     g09786(.I(\A[771] ), .ZN(new_n10789_));
  NAND2_X1   g09787(.A1(new_n10789_), .A2(\A[770] ), .ZN(new_n10790_));
  AOI21_X1   g09788(.A1(new_n10788_), .A2(new_n10790_), .B(new_n10786_), .ZN(new_n10791_));
  NOR2_X1    g09789(.A1(\A[770] ), .A2(\A[771] ), .ZN(new_n10792_));
  INV_X1     g09790(.I(new_n10792_), .ZN(new_n10793_));
  NAND2_X1   g09791(.A1(\A[770] ), .A2(\A[771] ), .ZN(new_n10794_));
  AOI21_X1   g09792(.A1(new_n10793_), .A2(new_n10794_), .B(\A[769] ), .ZN(new_n10795_));
  NOR2_X1    g09793(.A1(new_n10795_), .A2(new_n10791_), .ZN(new_n10796_));
  INV_X1     g09794(.I(\A[772] ), .ZN(new_n10797_));
  INV_X1     g09795(.I(\A[773] ), .ZN(new_n10798_));
  NAND2_X1   g09796(.A1(new_n10798_), .A2(\A[774] ), .ZN(new_n10799_));
  INV_X1     g09797(.I(\A[774] ), .ZN(new_n10800_));
  NAND2_X1   g09798(.A1(new_n10800_), .A2(\A[773] ), .ZN(new_n10801_));
  AOI21_X1   g09799(.A1(new_n10799_), .A2(new_n10801_), .B(new_n10797_), .ZN(new_n10802_));
  NOR2_X1    g09800(.A1(\A[773] ), .A2(\A[774] ), .ZN(new_n10803_));
  INV_X1     g09801(.I(new_n10803_), .ZN(new_n10804_));
  NAND2_X1   g09802(.A1(\A[773] ), .A2(\A[774] ), .ZN(new_n10805_));
  AOI21_X1   g09803(.A1(new_n10804_), .A2(new_n10805_), .B(\A[772] ), .ZN(new_n10806_));
  NOR2_X1    g09804(.A1(new_n10806_), .A2(new_n10802_), .ZN(new_n10807_));
  NAND2_X1   g09805(.A1(new_n10796_), .A2(new_n10807_), .ZN(new_n10808_));
  NOR2_X1    g09806(.A1(new_n10789_), .A2(\A[770] ), .ZN(new_n10809_));
  NOR2_X1    g09807(.A1(new_n10787_), .A2(\A[771] ), .ZN(new_n10810_));
  OAI21_X1   g09808(.A1(new_n10809_), .A2(new_n10810_), .B(\A[769] ), .ZN(new_n10811_));
  INV_X1     g09809(.I(new_n10794_), .ZN(new_n10812_));
  OAI21_X1   g09810(.A1(new_n10812_), .A2(new_n10792_), .B(new_n10786_), .ZN(new_n10813_));
  NAND2_X1   g09811(.A1(new_n10811_), .A2(new_n10813_), .ZN(new_n10814_));
  NOR2_X1    g09812(.A1(new_n10800_), .A2(\A[773] ), .ZN(new_n10815_));
  NOR2_X1    g09813(.A1(new_n10798_), .A2(\A[774] ), .ZN(new_n10816_));
  OAI21_X1   g09814(.A1(new_n10815_), .A2(new_n10816_), .B(\A[772] ), .ZN(new_n10817_));
  INV_X1     g09815(.I(new_n10805_), .ZN(new_n10818_));
  OAI21_X1   g09816(.A1(new_n10818_), .A2(new_n10803_), .B(new_n10797_), .ZN(new_n10819_));
  NAND2_X1   g09817(.A1(new_n10817_), .A2(new_n10819_), .ZN(new_n10820_));
  NAND2_X1   g09818(.A1(new_n10814_), .A2(new_n10820_), .ZN(new_n10821_));
  INV_X1     g09819(.I(\A[765] ), .ZN(new_n10822_));
  NOR2_X1    g09820(.A1(new_n10822_), .A2(\A[764] ), .ZN(new_n10823_));
  INV_X1     g09821(.I(\A[764] ), .ZN(new_n10824_));
  NOR2_X1    g09822(.A1(new_n10824_), .A2(\A[765] ), .ZN(new_n10825_));
  OAI21_X1   g09823(.A1(new_n10823_), .A2(new_n10825_), .B(\A[763] ), .ZN(new_n10826_));
  INV_X1     g09824(.I(\A[763] ), .ZN(new_n10827_));
  NAND2_X1   g09825(.A1(\A[764] ), .A2(\A[765] ), .ZN(new_n10828_));
  INV_X1     g09826(.I(new_n10828_), .ZN(new_n10829_));
  NOR2_X1    g09827(.A1(\A[764] ), .A2(\A[765] ), .ZN(new_n10830_));
  OAI21_X1   g09828(.A1(new_n10829_), .A2(new_n10830_), .B(new_n10827_), .ZN(new_n10831_));
  NAND2_X1   g09829(.A1(new_n10826_), .A2(new_n10831_), .ZN(new_n10832_));
  INV_X1     g09830(.I(\A[768] ), .ZN(new_n10833_));
  NOR2_X1    g09831(.A1(new_n10833_), .A2(\A[767] ), .ZN(new_n10834_));
  INV_X1     g09832(.I(\A[767] ), .ZN(new_n10835_));
  NOR2_X1    g09833(.A1(new_n10835_), .A2(\A[768] ), .ZN(new_n10836_));
  OAI21_X1   g09834(.A1(new_n10834_), .A2(new_n10836_), .B(\A[766] ), .ZN(new_n10837_));
  INV_X1     g09835(.I(\A[766] ), .ZN(new_n10838_));
  NAND2_X1   g09836(.A1(\A[767] ), .A2(\A[768] ), .ZN(new_n10839_));
  INV_X1     g09837(.I(new_n10839_), .ZN(new_n10840_));
  NOR2_X1    g09838(.A1(\A[767] ), .A2(\A[768] ), .ZN(new_n10841_));
  OAI21_X1   g09839(.A1(new_n10840_), .A2(new_n10841_), .B(new_n10838_), .ZN(new_n10842_));
  NAND2_X1   g09840(.A1(new_n10837_), .A2(new_n10842_), .ZN(new_n10843_));
  NOR2_X1    g09841(.A1(new_n10832_), .A2(new_n10843_), .ZN(new_n10844_));
  NAND2_X1   g09842(.A1(new_n10824_), .A2(\A[765] ), .ZN(new_n10845_));
  NAND2_X1   g09843(.A1(new_n10822_), .A2(\A[764] ), .ZN(new_n10846_));
  AOI21_X1   g09844(.A1(new_n10845_), .A2(new_n10846_), .B(new_n10827_), .ZN(new_n10847_));
  INV_X1     g09845(.I(new_n10830_), .ZN(new_n10848_));
  AOI21_X1   g09846(.A1(new_n10848_), .A2(new_n10828_), .B(\A[763] ), .ZN(new_n10849_));
  NOR2_X1    g09847(.A1(new_n10849_), .A2(new_n10847_), .ZN(new_n10850_));
  NAND2_X1   g09848(.A1(new_n10835_), .A2(\A[768] ), .ZN(new_n10851_));
  NAND2_X1   g09849(.A1(new_n10833_), .A2(\A[767] ), .ZN(new_n10852_));
  AOI21_X1   g09850(.A1(new_n10851_), .A2(new_n10852_), .B(new_n10838_), .ZN(new_n10853_));
  INV_X1     g09851(.I(new_n10841_), .ZN(new_n10854_));
  AOI21_X1   g09852(.A1(new_n10854_), .A2(new_n10839_), .B(\A[766] ), .ZN(new_n10855_));
  NOR2_X1    g09853(.A1(new_n10855_), .A2(new_n10853_), .ZN(new_n10856_));
  NOR2_X1    g09854(.A1(new_n10850_), .A2(new_n10856_), .ZN(new_n10857_));
  NOR2_X1    g09855(.A1(new_n10857_), .A2(new_n10844_), .ZN(new_n10858_));
  AOI21_X1   g09856(.A1(new_n10797_), .A2(new_n10805_), .B(new_n10803_), .ZN(new_n10859_));
  AOI21_X1   g09857(.A1(new_n10786_), .A2(new_n10794_), .B(new_n10792_), .ZN(new_n10860_));
  XOR2_X1    g09858(.A1(new_n10859_), .A2(new_n10860_), .Z(new_n10861_));
  NAND4_X1   g09859(.A1(new_n10858_), .A2(new_n10808_), .A3(new_n10821_), .A4(new_n10861_), .ZN(new_n10862_));
  INV_X1     g09860(.I(new_n10862_), .ZN(new_n10863_));
  AOI21_X1   g09861(.A1(\A[767] ), .A2(\A[768] ), .B(\A[766] ), .ZN(new_n10864_));
  AOI21_X1   g09862(.A1(\A[764] ), .A2(\A[765] ), .B(\A[763] ), .ZN(new_n10865_));
  OAI22_X1   g09863(.A1(new_n10830_), .A2(new_n10865_), .B1(new_n10864_), .B2(new_n10841_), .ZN(new_n10866_));
  NOR4_X1    g09864(.A1(new_n10864_), .A2(new_n10865_), .A3(new_n10830_), .A4(new_n10841_), .ZN(new_n10867_));
  INV_X1     g09865(.I(new_n10867_), .ZN(new_n10868_));
  NAND2_X1   g09866(.A1(new_n10868_), .A2(new_n10866_), .ZN(new_n10869_));
  XOR2_X1    g09867(.A1(new_n10844_), .A2(new_n10869_), .Z(new_n10870_));
  NOR2_X1    g09868(.A1(new_n10814_), .A2(new_n10820_), .ZN(new_n10871_));
  NOR2_X1    g09869(.A1(new_n10871_), .A2(new_n10861_), .ZN(new_n10872_));
  XNOR2_X1   g09870(.A1(new_n10859_), .A2(new_n10860_), .ZN(new_n10873_));
  NOR2_X1    g09871(.A1(new_n10808_), .A2(new_n10873_), .ZN(new_n10874_));
  OR2_X2     g09872(.A1(new_n10874_), .A2(new_n10872_), .Z(new_n10875_));
  NOR2_X1    g09873(.A1(new_n10796_), .A2(new_n10807_), .ZN(new_n10876_));
  NOR2_X1    g09874(.A1(new_n10876_), .A2(new_n10871_), .ZN(new_n10877_));
  NAND2_X1   g09875(.A1(new_n10858_), .A2(new_n10877_), .ZN(new_n10878_));
  AOI21_X1   g09876(.A1(new_n10875_), .A2(new_n10878_), .B(new_n10870_), .ZN(new_n10879_));
  INV_X1     g09877(.I(new_n10859_), .ZN(new_n10880_));
  INV_X1     g09878(.I(new_n10860_), .ZN(new_n10881_));
  NOR2_X1    g09879(.A1(new_n10880_), .A2(new_n10881_), .ZN(new_n10882_));
  INV_X1     g09880(.I(new_n10882_), .ZN(new_n10883_));
  NOR2_X1    g09881(.A1(new_n10859_), .A2(new_n10860_), .ZN(new_n10884_));
  AOI21_X1   g09882(.A1(new_n10808_), .A2(new_n10883_), .B(new_n10884_), .ZN(new_n10885_));
  NAND2_X1   g09883(.A1(new_n10850_), .A2(new_n10856_), .ZN(new_n10886_));
  INV_X1     g09884(.I(new_n10866_), .ZN(new_n10887_));
  AOI21_X1   g09885(.A1(new_n10886_), .A2(new_n10868_), .B(new_n10887_), .ZN(new_n10888_));
  NOR2_X1    g09886(.A1(new_n10885_), .A2(new_n10888_), .ZN(new_n10889_));
  INV_X1     g09887(.I(new_n10884_), .ZN(new_n10890_));
  OAI21_X1   g09888(.A1(new_n10871_), .A2(new_n10882_), .B(new_n10890_), .ZN(new_n10891_));
  OAI21_X1   g09889(.A1(new_n10844_), .A2(new_n10867_), .B(new_n10866_), .ZN(new_n10892_));
  NOR2_X1    g09890(.A1(new_n10891_), .A2(new_n10892_), .ZN(new_n10893_));
  NOR2_X1    g09891(.A1(new_n10889_), .A2(new_n10893_), .ZN(new_n10894_));
  OAI21_X1   g09892(.A1(new_n10879_), .A2(new_n10863_), .B(new_n10894_), .ZN(new_n10895_));
  XOR2_X1    g09893(.A1(new_n10886_), .A2(new_n10869_), .Z(new_n10896_));
  NAND2_X1   g09894(.A1(new_n10808_), .A2(new_n10821_), .ZN(new_n10897_));
  NAND2_X1   g09895(.A1(new_n10832_), .A2(new_n10843_), .ZN(new_n10898_));
  NAND2_X1   g09896(.A1(new_n10886_), .A2(new_n10898_), .ZN(new_n10899_));
  OAI22_X1   g09897(.A1(new_n10897_), .A2(new_n10899_), .B1(new_n10874_), .B2(new_n10872_), .ZN(new_n10900_));
  NAND2_X1   g09898(.A1(new_n10900_), .A2(new_n10896_), .ZN(new_n10901_));
  NAND2_X1   g09899(.A1(new_n10891_), .A2(new_n10892_), .ZN(new_n10902_));
  NAND2_X1   g09900(.A1(new_n10885_), .A2(new_n10888_), .ZN(new_n10903_));
  NAND2_X1   g09901(.A1(new_n10903_), .A2(new_n10902_), .ZN(new_n10904_));
  NAND3_X1   g09902(.A1(new_n10901_), .A2(new_n10904_), .A3(new_n10862_), .ZN(new_n10905_));
  NAND2_X1   g09903(.A1(new_n10895_), .A2(new_n10905_), .ZN(new_n10906_));
  INV_X1     g09904(.I(\A[759] ), .ZN(new_n10907_));
  NOR2_X1    g09905(.A1(new_n10907_), .A2(\A[758] ), .ZN(new_n10908_));
  INV_X1     g09906(.I(\A[758] ), .ZN(new_n10909_));
  NOR2_X1    g09907(.A1(new_n10909_), .A2(\A[759] ), .ZN(new_n10910_));
  OAI21_X1   g09908(.A1(new_n10908_), .A2(new_n10910_), .B(\A[757] ), .ZN(new_n10911_));
  INV_X1     g09909(.I(\A[757] ), .ZN(new_n10912_));
  NOR2_X1    g09910(.A1(\A[758] ), .A2(\A[759] ), .ZN(new_n10913_));
  NAND2_X1   g09911(.A1(\A[758] ), .A2(\A[759] ), .ZN(new_n10914_));
  INV_X1     g09912(.I(new_n10914_), .ZN(new_n10915_));
  OAI21_X1   g09913(.A1(new_n10915_), .A2(new_n10913_), .B(new_n10912_), .ZN(new_n10916_));
  NAND2_X1   g09914(.A1(new_n10911_), .A2(new_n10916_), .ZN(new_n10917_));
  INV_X1     g09915(.I(\A[762] ), .ZN(new_n10918_));
  NOR2_X1    g09916(.A1(new_n10918_), .A2(\A[761] ), .ZN(new_n10919_));
  INV_X1     g09917(.I(\A[761] ), .ZN(new_n10920_));
  NOR2_X1    g09918(.A1(new_n10920_), .A2(\A[762] ), .ZN(new_n10921_));
  OAI21_X1   g09919(.A1(new_n10919_), .A2(new_n10921_), .B(\A[760] ), .ZN(new_n10922_));
  INV_X1     g09920(.I(\A[760] ), .ZN(new_n10923_));
  NOR2_X1    g09921(.A1(\A[761] ), .A2(\A[762] ), .ZN(new_n10924_));
  NAND2_X1   g09922(.A1(\A[761] ), .A2(\A[762] ), .ZN(new_n10925_));
  INV_X1     g09923(.I(new_n10925_), .ZN(new_n10926_));
  OAI21_X1   g09924(.A1(new_n10926_), .A2(new_n10924_), .B(new_n10923_), .ZN(new_n10927_));
  NAND2_X1   g09925(.A1(new_n10922_), .A2(new_n10927_), .ZN(new_n10928_));
  NOR2_X1    g09926(.A1(new_n10917_), .A2(new_n10928_), .ZN(new_n10929_));
  AOI21_X1   g09927(.A1(new_n10923_), .A2(new_n10925_), .B(new_n10924_), .ZN(new_n10930_));
  AOI21_X1   g09928(.A1(new_n10912_), .A2(new_n10914_), .B(new_n10913_), .ZN(new_n10931_));
  AND2_X2    g09929(.A1(new_n10930_), .A2(new_n10931_), .Z(new_n10932_));
  NOR2_X1    g09930(.A1(new_n10930_), .A2(new_n10931_), .ZN(new_n10933_));
  INV_X1     g09931(.I(new_n10933_), .ZN(new_n10934_));
  OAI21_X1   g09932(.A1(new_n10929_), .A2(new_n10932_), .B(new_n10934_), .ZN(new_n10935_));
  INV_X1     g09933(.I(\A[751] ), .ZN(new_n10936_));
  INV_X1     g09934(.I(\A[752] ), .ZN(new_n10937_));
  NAND2_X1   g09935(.A1(new_n10937_), .A2(\A[753] ), .ZN(new_n10938_));
  INV_X1     g09936(.I(\A[753] ), .ZN(new_n10939_));
  NAND2_X1   g09937(.A1(new_n10939_), .A2(\A[752] ), .ZN(new_n10940_));
  AOI21_X1   g09938(.A1(new_n10938_), .A2(new_n10940_), .B(new_n10936_), .ZN(new_n10941_));
  NAND2_X1   g09939(.A1(\A[752] ), .A2(\A[753] ), .ZN(new_n10942_));
  NOR2_X1    g09940(.A1(\A[752] ), .A2(\A[753] ), .ZN(new_n10943_));
  INV_X1     g09941(.I(new_n10943_), .ZN(new_n10944_));
  AOI21_X1   g09942(.A1(new_n10944_), .A2(new_n10942_), .B(\A[751] ), .ZN(new_n10945_));
  INV_X1     g09943(.I(\A[754] ), .ZN(new_n10946_));
  INV_X1     g09944(.I(\A[755] ), .ZN(new_n10947_));
  NAND2_X1   g09945(.A1(new_n10947_), .A2(\A[756] ), .ZN(new_n10948_));
  INV_X1     g09946(.I(\A[756] ), .ZN(new_n10949_));
  NAND2_X1   g09947(.A1(new_n10949_), .A2(\A[755] ), .ZN(new_n10950_));
  AOI21_X1   g09948(.A1(new_n10948_), .A2(new_n10950_), .B(new_n10946_), .ZN(new_n10951_));
  NAND2_X1   g09949(.A1(\A[755] ), .A2(\A[756] ), .ZN(new_n10952_));
  NOR2_X1    g09950(.A1(\A[755] ), .A2(\A[756] ), .ZN(new_n10953_));
  INV_X1     g09951(.I(new_n10953_), .ZN(new_n10954_));
  AOI21_X1   g09952(.A1(new_n10954_), .A2(new_n10952_), .B(\A[754] ), .ZN(new_n10955_));
  NOR4_X1    g09953(.A1(new_n10941_), .A2(new_n10945_), .A3(new_n10955_), .A4(new_n10951_), .ZN(new_n10956_));
  AOI21_X1   g09954(.A1(new_n10946_), .A2(new_n10952_), .B(new_n10953_), .ZN(new_n10957_));
  AOI21_X1   g09955(.A1(new_n10936_), .A2(new_n10942_), .B(new_n10943_), .ZN(new_n10958_));
  NOR2_X1    g09956(.A1(new_n10957_), .A2(new_n10958_), .ZN(new_n10959_));
  INV_X1     g09957(.I(new_n10959_), .ZN(new_n10960_));
  NAND2_X1   g09958(.A1(new_n10957_), .A2(new_n10958_), .ZN(new_n10961_));
  NAND2_X1   g09959(.A1(new_n10960_), .A2(new_n10961_), .ZN(new_n10962_));
  XOR2_X1    g09960(.A1(new_n10962_), .A2(new_n10956_), .Z(new_n10963_));
  NAND2_X1   g09961(.A1(new_n10909_), .A2(\A[759] ), .ZN(new_n10964_));
  NAND2_X1   g09962(.A1(new_n10907_), .A2(\A[758] ), .ZN(new_n10965_));
  AOI21_X1   g09963(.A1(new_n10964_), .A2(new_n10965_), .B(new_n10912_), .ZN(new_n10966_));
  INV_X1     g09964(.I(new_n10913_), .ZN(new_n10967_));
  AOI21_X1   g09965(.A1(new_n10967_), .A2(new_n10914_), .B(\A[757] ), .ZN(new_n10968_));
  NOR2_X1    g09966(.A1(new_n10968_), .A2(new_n10966_), .ZN(new_n10969_));
  NAND2_X1   g09967(.A1(new_n10920_), .A2(\A[762] ), .ZN(new_n10970_));
  NAND2_X1   g09968(.A1(new_n10918_), .A2(\A[761] ), .ZN(new_n10971_));
  AOI21_X1   g09969(.A1(new_n10970_), .A2(new_n10971_), .B(new_n10923_), .ZN(new_n10972_));
  INV_X1     g09970(.I(new_n10924_), .ZN(new_n10973_));
  AOI21_X1   g09971(.A1(new_n10973_), .A2(new_n10925_), .B(\A[760] ), .ZN(new_n10974_));
  NOR2_X1    g09972(.A1(new_n10974_), .A2(new_n10972_), .ZN(new_n10975_));
  NOR2_X1    g09973(.A1(new_n10969_), .A2(new_n10975_), .ZN(new_n10976_));
  NOR2_X1    g09974(.A1(new_n10976_), .A2(new_n10929_), .ZN(new_n10977_));
  OAI22_X1   g09975(.A1(new_n10941_), .A2(new_n10945_), .B1(new_n10955_), .B2(new_n10951_), .ZN(new_n10978_));
  INV_X1     g09976(.I(new_n10978_), .ZN(new_n10979_));
  NOR2_X1    g09977(.A1(new_n10979_), .A2(new_n10956_), .ZN(new_n10980_));
  NAND2_X1   g09978(.A1(new_n10969_), .A2(new_n10975_), .ZN(new_n10981_));
  XNOR2_X1   g09979(.A1(new_n10930_), .A2(new_n10931_), .ZN(new_n10982_));
  NAND2_X1   g09980(.A1(new_n10981_), .A2(new_n10982_), .ZN(new_n10983_));
  XOR2_X1    g09981(.A1(new_n10930_), .A2(new_n10931_), .Z(new_n10984_));
  NAND2_X1   g09982(.A1(new_n10929_), .A2(new_n10984_), .ZN(new_n10985_));
  AOI22_X1   g09983(.A1(new_n10980_), .A2(new_n10977_), .B1(new_n10983_), .B2(new_n10985_), .ZN(new_n10986_));
  NOR2_X1    g09984(.A1(new_n10986_), .A2(new_n10963_), .ZN(new_n10987_));
  NAND2_X1   g09985(.A1(new_n10983_), .A2(new_n10985_), .ZN(new_n10988_));
  NAND2_X1   g09986(.A1(new_n10980_), .A2(new_n10977_), .ZN(new_n10989_));
  NOR2_X1    g09987(.A1(new_n10989_), .A2(new_n10988_), .ZN(new_n10990_));
  NOR2_X1    g09988(.A1(new_n10945_), .A2(new_n10941_), .ZN(new_n10991_));
  NOR2_X1    g09989(.A1(new_n10955_), .A2(new_n10951_), .ZN(new_n10992_));
  NAND2_X1   g09990(.A1(new_n10991_), .A2(new_n10992_), .ZN(new_n10993_));
  AOI21_X1   g09991(.A1(new_n10993_), .A2(new_n10961_), .B(new_n10959_), .ZN(new_n10994_));
  NOR3_X1    g09992(.A1(new_n10987_), .A2(new_n10990_), .A3(new_n10994_), .ZN(new_n10995_));
  NAND3_X1   g09993(.A1(new_n10993_), .A2(new_n10960_), .A3(new_n10961_), .ZN(new_n10996_));
  NAND2_X1   g09994(.A1(new_n10962_), .A2(new_n10956_), .ZN(new_n10997_));
  NAND2_X1   g09995(.A1(new_n10996_), .A2(new_n10997_), .ZN(new_n10998_));
  XOR2_X1    g09996(.A1(new_n10929_), .A2(new_n10984_), .Z(new_n10999_));
  NAND2_X1   g09997(.A1(new_n10917_), .A2(new_n10928_), .ZN(new_n11000_));
  NAND2_X1   g09998(.A1(new_n10981_), .A2(new_n11000_), .ZN(new_n11001_));
  NAND2_X1   g09999(.A1(new_n10993_), .A2(new_n10978_), .ZN(new_n11002_));
  NOR2_X1    g10000(.A1(new_n11001_), .A2(new_n11002_), .ZN(new_n11003_));
  OAI21_X1   g10001(.A1(new_n10999_), .A2(new_n11003_), .B(new_n10998_), .ZN(new_n11004_));
  NAND3_X1   g10002(.A1(new_n11003_), .A2(new_n10983_), .A3(new_n10985_), .ZN(new_n11005_));
  INV_X1     g10003(.I(new_n10994_), .ZN(new_n11006_));
  AOI21_X1   g10004(.A1(new_n11004_), .A2(new_n11005_), .B(new_n11006_), .ZN(new_n11007_));
  NOR3_X1    g10005(.A1(new_n10995_), .A2(new_n11007_), .A3(new_n10935_), .ZN(new_n11008_));
  INV_X1     g10006(.I(new_n10935_), .ZN(new_n11009_));
  NAND3_X1   g10007(.A1(new_n11004_), .A2(new_n11005_), .A3(new_n11006_), .ZN(new_n11010_));
  OAI21_X1   g10008(.A1(new_n10987_), .A2(new_n10990_), .B(new_n10994_), .ZN(new_n11011_));
  AOI21_X1   g10009(.A1(new_n11011_), .A2(new_n11010_), .B(new_n11009_), .ZN(new_n11012_));
  OAI21_X1   g10010(.A1(new_n11008_), .A2(new_n11012_), .B(new_n10906_), .ZN(new_n11013_));
  AOI21_X1   g10011(.A1(new_n10901_), .A2(new_n10862_), .B(new_n10904_), .ZN(new_n11014_));
  NOR3_X1    g10012(.A1(new_n10879_), .A2(new_n10863_), .A3(new_n10894_), .ZN(new_n11015_));
  NOR2_X1    g10013(.A1(new_n11015_), .A2(new_n11014_), .ZN(new_n11016_));
  NAND3_X1   g10014(.A1(new_n11011_), .A2(new_n11010_), .A3(new_n11009_), .ZN(new_n11017_));
  OAI21_X1   g10015(.A1(new_n10995_), .A2(new_n11007_), .B(new_n10935_), .ZN(new_n11018_));
  NAND3_X1   g10016(.A1(new_n11016_), .A2(new_n11018_), .A3(new_n11017_), .ZN(new_n11019_));
  NAND3_X1   g10017(.A1(new_n10900_), .A2(new_n10870_), .A3(new_n10862_), .ZN(new_n11020_));
  AOI21_X1   g10018(.A1(new_n10900_), .A2(new_n10862_), .B(new_n10870_), .ZN(new_n11021_));
  INV_X1     g10019(.I(new_n11021_), .ZN(new_n11022_));
  NAND2_X1   g10020(.A1(new_n11022_), .A2(new_n11020_), .ZN(new_n11023_));
  NOR2_X1    g10021(.A1(new_n10858_), .A2(new_n10897_), .ZN(new_n11024_));
  NOR2_X1    g10022(.A1(new_n10877_), .A2(new_n10899_), .ZN(new_n11025_));
  NOR2_X1    g10023(.A1(new_n10980_), .A2(new_n11001_), .ZN(new_n11026_));
  NOR2_X1    g10024(.A1(new_n10977_), .A2(new_n11002_), .ZN(new_n11027_));
  OAI22_X1   g10025(.A1(new_n11024_), .A2(new_n11025_), .B1(new_n11026_), .B2(new_n11027_), .ZN(new_n11028_));
  NOR2_X1    g10026(.A1(new_n11004_), .A2(new_n10990_), .ZN(new_n11029_));
  NAND2_X1   g10027(.A1(new_n10989_), .A2(new_n10988_), .ZN(new_n11030_));
  AOI21_X1   g10028(.A1(new_n11030_), .A2(new_n11005_), .B(new_n10998_), .ZN(new_n11031_));
  NOR3_X1    g10029(.A1(new_n11029_), .A2(new_n11031_), .A3(new_n11028_), .ZN(new_n11032_));
  OAI21_X1   g10030(.A1(new_n11029_), .A2(new_n11031_), .B(new_n11028_), .ZN(new_n11033_));
  OAI21_X1   g10031(.A1(new_n11023_), .A2(new_n11032_), .B(new_n11033_), .ZN(new_n11034_));
  NAND3_X1   g10032(.A1(new_n11013_), .A2(new_n11019_), .A3(new_n11034_), .ZN(new_n11035_));
  AOI21_X1   g10033(.A1(new_n11018_), .A2(new_n11017_), .B(new_n11016_), .ZN(new_n11036_));
  NOR3_X1    g10034(.A1(new_n11008_), .A2(new_n11012_), .A3(new_n10906_), .ZN(new_n11037_));
  INV_X1     g10035(.I(new_n11020_), .ZN(new_n11038_));
  NOR2_X1    g10036(.A1(new_n11038_), .A2(new_n11021_), .ZN(new_n11039_));
  NAND2_X1   g10037(.A1(new_n10877_), .A2(new_n10899_), .ZN(new_n11040_));
  NAND2_X1   g10038(.A1(new_n10858_), .A2(new_n10897_), .ZN(new_n11041_));
  NAND2_X1   g10039(.A1(new_n10977_), .A2(new_n11002_), .ZN(new_n11042_));
  NAND2_X1   g10040(.A1(new_n10980_), .A2(new_n11001_), .ZN(new_n11043_));
  AOI22_X1   g10041(.A1(new_n11040_), .A2(new_n11041_), .B1(new_n11043_), .B2(new_n11042_), .ZN(new_n11044_));
  NAND2_X1   g10042(.A1(new_n10987_), .A2(new_n11005_), .ZN(new_n11045_));
  OAI21_X1   g10043(.A1(new_n10990_), .A2(new_n10986_), .B(new_n10963_), .ZN(new_n11046_));
  NAND3_X1   g10044(.A1(new_n11045_), .A2(new_n11046_), .A3(new_n11044_), .ZN(new_n11047_));
  AOI21_X1   g10045(.A1(new_n11045_), .A2(new_n11046_), .B(new_n11044_), .ZN(new_n11048_));
  AOI21_X1   g10046(.A1(new_n11039_), .A2(new_n11047_), .B(new_n11048_), .ZN(new_n11049_));
  OAI21_X1   g10047(.A1(new_n11036_), .A2(new_n11037_), .B(new_n11049_), .ZN(new_n11050_));
  NAND2_X1   g10048(.A1(new_n10722_), .A2(new_n10742_), .ZN(new_n11051_));
  AOI22_X1   g10049(.A1(new_n11051_), .A2(new_n10770_), .B1(new_n10771_), .B2(new_n10729_), .ZN(new_n11052_));
  OAI21_X1   g10050(.A1(new_n10754_), .A2(new_n10633_), .B(new_n10604_), .ZN(new_n11053_));
  NAND4_X1   g10051(.A1(new_n10750_), .A2(new_n10617_), .A3(new_n10624_), .A4(new_n10620_), .ZN(new_n11054_));
  NAND3_X1   g10052(.A1(new_n10626_), .A2(new_n10746_), .A3(new_n11054_), .ZN(new_n11055_));
  NAND2_X1   g10053(.A1(new_n10716_), .A2(new_n10725_), .ZN(new_n11056_));
  NAND2_X1   g10054(.A1(new_n10702_), .A2(new_n10738_), .ZN(new_n11057_));
  NAND2_X1   g10055(.A1(new_n11057_), .A2(new_n11056_), .ZN(new_n11058_));
  INV_X1     g10056(.I(new_n10625_), .ZN(new_n11059_));
  AOI22_X1   g10057(.A1(new_n10622_), .A2(new_n10623_), .B1(new_n10617_), .B2(new_n10624_), .ZN(new_n11060_));
  NOR2_X1    g10058(.A1(new_n11059_), .A2(new_n11060_), .ZN(new_n11061_));
  NAND2_X1   g10059(.A1(new_n11058_), .A2(new_n11061_), .ZN(new_n11062_));
  AOI21_X1   g10060(.A1(new_n11053_), .A2(new_n11055_), .B(new_n11062_), .ZN(new_n11063_));
  NAND3_X1   g10061(.A1(new_n11062_), .A2(new_n11053_), .A3(new_n11055_), .ZN(new_n11064_));
  OAI21_X1   g10062(.A1(new_n11063_), .A2(new_n11052_), .B(new_n11064_), .ZN(new_n11065_));
  NOR2_X1    g10063(.A1(new_n10634_), .A2(new_n10768_), .ZN(new_n11066_));
  NOR2_X1    g10064(.A1(new_n10765_), .A2(new_n10766_), .ZN(new_n11067_));
  AOI22_X1   g10065(.A1(new_n10723_), .A2(new_n10729_), .B1(new_n10773_), .B2(new_n10774_), .ZN(new_n11068_));
  NOR4_X1    g10066(.A1(new_n10771_), .A2(new_n10737_), .A3(new_n10697_), .A4(new_n10733_), .ZN(new_n11069_));
  OAI22_X1   g10067(.A1(new_n11067_), .A2(new_n11066_), .B1(new_n11068_), .B2(new_n11069_), .ZN(new_n11070_));
  NAND3_X1   g10068(.A1(new_n11070_), .A2(new_n11065_), .A3(new_n10776_), .ZN(new_n11071_));
  NOR4_X1    g10069(.A1(new_n11067_), .A2(new_n11066_), .A3(new_n11068_), .A4(new_n11069_), .ZN(new_n11072_));
  OAI21_X1   g10070(.A1(new_n11072_), .A2(new_n10777_), .B(new_n10764_), .ZN(new_n11073_));
  NAND4_X1   g10071(.A1(new_n11050_), .A2(new_n11035_), .A3(new_n11073_), .A4(new_n11071_), .ZN(new_n11074_));
  AOI22_X1   g10072(.A1(new_n11050_), .A2(new_n11035_), .B1(new_n11073_), .B2(new_n11071_), .ZN(new_n11075_));
  AOI21_X1   g10073(.A1(new_n10762_), .A2(new_n11064_), .B(new_n10745_), .ZN(new_n11076_));
  NOR3_X1    g10074(.A1(new_n11063_), .A2(new_n10763_), .A3(new_n11052_), .ZN(new_n11077_));
  NOR2_X1    g10075(.A1(new_n11076_), .A2(new_n11077_), .ZN(new_n11078_));
  NOR4_X1    g10076(.A1(new_n11024_), .A2(new_n11025_), .A3(new_n11026_), .A4(new_n11027_), .ZN(new_n11079_));
  NOR2_X1    g10077(.A1(new_n11079_), .A2(new_n11044_), .ZN(new_n11080_));
  INV_X1     g10078(.I(new_n11080_), .ZN(new_n11081_));
  XOR2_X1    g10079(.A1(new_n10627_), .A2(new_n10758_), .Z(new_n11082_));
  NAND2_X1   g10080(.A1(new_n11082_), .A2(new_n10757_), .ZN(new_n11083_));
  XOR2_X1    g10081(.A1(new_n10750_), .A2(new_n10758_), .Z(new_n11084_));
  NAND2_X1   g10082(.A1(new_n11084_), .A2(new_n11058_), .ZN(new_n11085_));
  AOI21_X1   g10083(.A1(new_n11083_), .A2(new_n11085_), .B(new_n11081_), .ZN(new_n11086_));
  NAND3_X1   g10084(.A1(new_n11033_), .A2(new_n11047_), .A3(new_n11023_), .ZN(new_n11087_));
  OAI21_X1   g10085(.A1(new_n11032_), .A2(new_n11048_), .B(new_n11039_), .ZN(new_n11088_));
  AOI21_X1   g10086(.A1(new_n11088_), .A2(new_n11087_), .B(new_n11086_), .ZN(new_n11089_));
  NAND3_X1   g10087(.A1(new_n11086_), .A2(new_n11088_), .A3(new_n11087_), .ZN(new_n11090_));
  AOI21_X1   g10088(.A1(new_n11078_), .A2(new_n11090_), .B(new_n11089_), .ZN(new_n11091_));
  OAI21_X1   g10089(.A1(new_n11075_), .A2(new_n11091_), .B(new_n11074_), .ZN(new_n11092_));
  AOI21_X1   g10090(.A1(new_n11013_), .A2(new_n11049_), .B(new_n11037_), .ZN(new_n11093_));
  AOI21_X1   g10091(.A1(new_n10935_), .A2(new_n11011_), .B(new_n10995_), .ZN(new_n11094_));
  NAND2_X1   g10092(.A1(new_n10901_), .A2(new_n10862_), .ZN(new_n11095_));
  OAI21_X1   g10093(.A1(new_n11095_), .A2(new_n10893_), .B(new_n10902_), .ZN(new_n11096_));
  XOR2_X1    g10094(.A1(new_n11094_), .A2(new_n11096_), .Z(new_n11097_));
  NOR2_X1    g10095(.A1(new_n11093_), .A2(new_n11097_), .ZN(new_n11098_));
  OAI21_X1   g10096(.A1(new_n11036_), .A2(new_n11034_), .B(new_n11019_), .ZN(new_n11099_));
  XNOR2_X1   g10097(.A1(new_n11094_), .A2(new_n11096_), .ZN(new_n11100_));
  NOR2_X1    g10098(.A1(new_n11100_), .A2(new_n11099_), .ZN(new_n11101_));
  NOR2_X1    g10099(.A1(new_n11101_), .A2(new_n11098_), .ZN(new_n11102_));
  NAND2_X1   g10100(.A1(new_n11092_), .A2(new_n11102_), .ZN(new_n11103_));
  NOR3_X1    g10101(.A1(new_n11036_), .A2(new_n11037_), .A3(new_n11049_), .ZN(new_n11104_));
  AOI21_X1   g10102(.A1(new_n11013_), .A2(new_n11019_), .B(new_n11034_), .ZN(new_n11105_));
  NOR3_X1    g10103(.A1(new_n10764_), .A2(new_n11072_), .A3(new_n10777_), .ZN(new_n11106_));
  AOI21_X1   g10104(.A1(new_n10776_), .A2(new_n11070_), .B(new_n11065_), .ZN(new_n11107_));
  NOR4_X1    g10105(.A1(new_n11104_), .A2(new_n11105_), .A3(new_n11106_), .A4(new_n11107_), .ZN(new_n11108_));
  OAI22_X1   g10106(.A1(new_n11104_), .A2(new_n11105_), .B1(new_n11106_), .B2(new_n11107_), .ZN(new_n11109_));
  OR2_X2     g10107(.A1(new_n11076_), .A2(new_n11077_), .Z(new_n11110_));
  NAND2_X1   g10108(.A1(new_n11083_), .A2(new_n11085_), .ZN(new_n11111_));
  NAND2_X1   g10109(.A1(new_n11111_), .A2(new_n11080_), .ZN(new_n11112_));
  NOR3_X1    g10110(.A1(new_n11032_), .A2(new_n11048_), .A3(new_n11039_), .ZN(new_n11113_));
  AOI21_X1   g10111(.A1(new_n11033_), .A2(new_n11047_), .B(new_n11023_), .ZN(new_n11114_));
  OAI21_X1   g10112(.A1(new_n11113_), .A2(new_n11114_), .B(new_n11112_), .ZN(new_n11115_));
  NOR3_X1    g10113(.A1(new_n11113_), .A2(new_n11114_), .A3(new_n11112_), .ZN(new_n11116_));
  OAI21_X1   g10114(.A1(new_n11110_), .A2(new_n11116_), .B(new_n11115_), .ZN(new_n11117_));
  AOI21_X1   g10115(.A1(new_n11109_), .A2(new_n11117_), .B(new_n11108_), .ZN(new_n11118_));
  INV_X1     g10116(.I(new_n11102_), .ZN(new_n11119_));
  NAND2_X1   g10117(.A1(new_n11119_), .A2(new_n11118_), .ZN(new_n11120_));
  AOI21_X1   g10118(.A1(new_n11120_), .A2(new_n11103_), .B(new_n10785_), .ZN(new_n11121_));
  NOR2_X1    g10119(.A1(new_n11119_), .A2(new_n11118_), .ZN(new_n11122_));
  NOR2_X1    g10120(.A1(new_n11092_), .A2(new_n11102_), .ZN(new_n11123_));
  NOR3_X1    g10121(.A1(new_n11122_), .A2(new_n11123_), .A3(new_n10784_), .ZN(new_n11124_));
  NOR2_X1    g10122(.A1(new_n11124_), .A2(new_n11121_), .ZN(new_n11125_));
  INV_X1     g10123(.I(new_n11125_), .ZN(new_n11126_));
  INV_X1     g10124(.I(\A[811] ), .ZN(new_n11127_));
  INV_X1     g10125(.I(\A[812] ), .ZN(new_n11128_));
  NAND2_X1   g10126(.A1(new_n11128_), .A2(\A[813] ), .ZN(new_n11129_));
  INV_X1     g10127(.I(\A[813] ), .ZN(new_n11130_));
  NAND2_X1   g10128(.A1(new_n11130_), .A2(\A[812] ), .ZN(new_n11131_));
  AOI21_X1   g10129(.A1(new_n11129_), .A2(new_n11131_), .B(new_n11127_), .ZN(new_n11132_));
  NAND2_X1   g10130(.A1(\A[812] ), .A2(\A[813] ), .ZN(new_n11133_));
  NOR2_X1    g10131(.A1(\A[812] ), .A2(\A[813] ), .ZN(new_n11134_));
  INV_X1     g10132(.I(new_n11134_), .ZN(new_n11135_));
  AOI21_X1   g10133(.A1(new_n11135_), .A2(new_n11133_), .B(\A[811] ), .ZN(new_n11136_));
  NOR2_X1    g10134(.A1(new_n11136_), .A2(new_n11132_), .ZN(new_n11137_));
  INV_X1     g10135(.I(\A[814] ), .ZN(new_n11138_));
  INV_X1     g10136(.I(\A[815] ), .ZN(new_n11139_));
  NAND2_X1   g10137(.A1(new_n11139_), .A2(\A[816] ), .ZN(new_n11140_));
  INV_X1     g10138(.I(\A[816] ), .ZN(new_n11141_));
  NAND2_X1   g10139(.A1(new_n11141_), .A2(\A[815] ), .ZN(new_n11142_));
  AOI21_X1   g10140(.A1(new_n11140_), .A2(new_n11142_), .B(new_n11138_), .ZN(new_n11143_));
  NAND2_X1   g10141(.A1(\A[815] ), .A2(\A[816] ), .ZN(new_n11144_));
  NOR2_X1    g10142(.A1(\A[815] ), .A2(\A[816] ), .ZN(new_n11145_));
  INV_X1     g10143(.I(new_n11145_), .ZN(new_n11146_));
  AOI21_X1   g10144(.A1(new_n11146_), .A2(new_n11144_), .B(\A[814] ), .ZN(new_n11147_));
  NOR2_X1    g10145(.A1(new_n11147_), .A2(new_n11143_), .ZN(new_n11148_));
  NAND2_X1   g10146(.A1(new_n11137_), .A2(new_n11148_), .ZN(new_n11149_));
  AOI21_X1   g10147(.A1(new_n11138_), .A2(new_n11144_), .B(new_n11145_), .ZN(new_n11150_));
  AOI21_X1   g10148(.A1(new_n11127_), .A2(new_n11133_), .B(new_n11134_), .ZN(new_n11151_));
  NOR2_X1    g10149(.A1(new_n11150_), .A2(new_n11151_), .ZN(new_n11152_));
  NAND2_X1   g10150(.A1(new_n11150_), .A2(new_n11151_), .ZN(new_n11153_));
  INV_X1     g10151(.I(new_n11153_), .ZN(new_n11154_));
  NOR2_X1    g10152(.A1(new_n11154_), .A2(new_n11152_), .ZN(new_n11155_));
  NAND2_X1   g10153(.A1(new_n11155_), .A2(new_n11149_), .ZN(new_n11156_));
  NOR2_X1    g10154(.A1(new_n11130_), .A2(\A[812] ), .ZN(new_n11157_));
  NOR2_X1    g10155(.A1(new_n11128_), .A2(\A[813] ), .ZN(new_n11158_));
  OAI21_X1   g10156(.A1(new_n11157_), .A2(new_n11158_), .B(\A[811] ), .ZN(new_n11159_));
  INV_X1     g10157(.I(new_n11133_), .ZN(new_n11160_));
  OAI21_X1   g10158(.A1(new_n11160_), .A2(new_n11134_), .B(new_n11127_), .ZN(new_n11161_));
  NAND2_X1   g10159(.A1(new_n11159_), .A2(new_n11161_), .ZN(new_n11162_));
  NOR2_X1    g10160(.A1(new_n11141_), .A2(\A[815] ), .ZN(new_n11163_));
  NOR2_X1    g10161(.A1(new_n11139_), .A2(\A[816] ), .ZN(new_n11164_));
  OAI21_X1   g10162(.A1(new_n11163_), .A2(new_n11164_), .B(\A[814] ), .ZN(new_n11165_));
  INV_X1     g10163(.I(new_n11144_), .ZN(new_n11166_));
  OAI21_X1   g10164(.A1(new_n11166_), .A2(new_n11145_), .B(new_n11138_), .ZN(new_n11167_));
  NAND2_X1   g10165(.A1(new_n11165_), .A2(new_n11167_), .ZN(new_n11168_));
  NOR2_X1    g10166(.A1(new_n11162_), .A2(new_n11168_), .ZN(new_n11169_));
  INV_X1     g10167(.I(new_n11152_), .ZN(new_n11170_));
  NAND2_X1   g10168(.A1(new_n11170_), .A2(new_n11153_), .ZN(new_n11171_));
  NAND2_X1   g10169(.A1(new_n11171_), .A2(new_n11169_), .ZN(new_n11172_));
  NAND2_X1   g10170(.A1(new_n11172_), .A2(new_n11156_), .ZN(new_n11173_));
  INV_X1     g10171(.I(\A[817] ), .ZN(new_n11174_));
  INV_X1     g10172(.I(\A[818] ), .ZN(new_n11175_));
  NAND2_X1   g10173(.A1(new_n11175_), .A2(\A[819] ), .ZN(new_n11176_));
  INV_X1     g10174(.I(\A[819] ), .ZN(new_n11177_));
  NAND2_X1   g10175(.A1(new_n11177_), .A2(\A[818] ), .ZN(new_n11178_));
  AOI21_X1   g10176(.A1(new_n11176_), .A2(new_n11178_), .B(new_n11174_), .ZN(new_n11179_));
  NAND2_X1   g10177(.A1(\A[818] ), .A2(\A[819] ), .ZN(new_n11180_));
  NOR2_X1    g10178(.A1(\A[818] ), .A2(\A[819] ), .ZN(new_n11181_));
  INV_X1     g10179(.I(new_n11181_), .ZN(new_n11182_));
  AOI21_X1   g10180(.A1(new_n11182_), .A2(new_n11180_), .B(\A[817] ), .ZN(new_n11183_));
  NOR2_X1    g10181(.A1(new_n11183_), .A2(new_n11179_), .ZN(new_n11184_));
  INV_X1     g10182(.I(\A[820] ), .ZN(new_n11185_));
  INV_X1     g10183(.I(\A[821] ), .ZN(new_n11186_));
  NAND2_X1   g10184(.A1(new_n11186_), .A2(\A[822] ), .ZN(new_n11187_));
  INV_X1     g10185(.I(\A[822] ), .ZN(new_n11188_));
  NAND2_X1   g10186(.A1(new_n11188_), .A2(\A[821] ), .ZN(new_n11189_));
  AOI21_X1   g10187(.A1(new_n11187_), .A2(new_n11189_), .B(new_n11185_), .ZN(new_n11190_));
  NAND2_X1   g10188(.A1(\A[821] ), .A2(\A[822] ), .ZN(new_n11191_));
  NOR2_X1    g10189(.A1(\A[821] ), .A2(\A[822] ), .ZN(new_n11192_));
  INV_X1     g10190(.I(new_n11192_), .ZN(new_n11193_));
  AOI21_X1   g10191(.A1(new_n11193_), .A2(new_n11191_), .B(\A[820] ), .ZN(new_n11194_));
  NOR2_X1    g10192(.A1(new_n11194_), .A2(new_n11190_), .ZN(new_n11195_));
  NAND2_X1   g10193(.A1(new_n11184_), .A2(new_n11195_), .ZN(new_n11196_));
  AOI21_X1   g10194(.A1(new_n11185_), .A2(new_n11191_), .B(new_n11192_), .ZN(new_n11197_));
  AOI21_X1   g10195(.A1(new_n11174_), .A2(new_n11180_), .B(new_n11181_), .ZN(new_n11198_));
  XOR2_X1    g10196(.A1(new_n11197_), .A2(new_n11198_), .Z(new_n11199_));
  NAND2_X1   g10197(.A1(new_n11196_), .A2(new_n11199_), .ZN(new_n11200_));
  NOR2_X1    g10198(.A1(new_n11177_), .A2(\A[818] ), .ZN(new_n11201_));
  NOR2_X1    g10199(.A1(new_n11175_), .A2(\A[819] ), .ZN(new_n11202_));
  OAI21_X1   g10200(.A1(new_n11201_), .A2(new_n11202_), .B(\A[817] ), .ZN(new_n11203_));
  INV_X1     g10201(.I(new_n11180_), .ZN(new_n11204_));
  OAI21_X1   g10202(.A1(new_n11204_), .A2(new_n11181_), .B(new_n11174_), .ZN(new_n11205_));
  NAND2_X1   g10203(.A1(new_n11203_), .A2(new_n11205_), .ZN(new_n11206_));
  NOR2_X1    g10204(.A1(new_n11188_), .A2(\A[821] ), .ZN(new_n11207_));
  NOR2_X1    g10205(.A1(new_n11186_), .A2(\A[822] ), .ZN(new_n11208_));
  OAI21_X1   g10206(.A1(new_n11207_), .A2(new_n11208_), .B(\A[820] ), .ZN(new_n11209_));
  INV_X1     g10207(.I(new_n11191_), .ZN(new_n11210_));
  OAI21_X1   g10208(.A1(new_n11210_), .A2(new_n11192_), .B(new_n11185_), .ZN(new_n11211_));
  NAND2_X1   g10209(.A1(new_n11209_), .A2(new_n11211_), .ZN(new_n11212_));
  NOR2_X1    g10210(.A1(new_n11206_), .A2(new_n11212_), .ZN(new_n11213_));
  XNOR2_X1   g10211(.A1(new_n11197_), .A2(new_n11198_), .ZN(new_n11214_));
  NAND2_X1   g10212(.A1(new_n11213_), .A2(new_n11214_), .ZN(new_n11215_));
  NAND2_X1   g10213(.A1(new_n11215_), .A2(new_n11200_), .ZN(new_n11216_));
  NAND2_X1   g10214(.A1(new_n11162_), .A2(new_n11168_), .ZN(new_n11217_));
  NAND2_X1   g10215(.A1(new_n11149_), .A2(new_n11217_), .ZN(new_n11218_));
  NAND2_X1   g10216(.A1(new_n11206_), .A2(new_n11212_), .ZN(new_n11219_));
  NAND2_X1   g10217(.A1(new_n11196_), .A2(new_n11219_), .ZN(new_n11220_));
  NOR2_X1    g10218(.A1(new_n11218_), .A2(new_n11220_), .ZN(new_n11221_));
  NOR2_X1    g10219(.A1(new_n11221_), .A2(new_n11216_), .ZN(new_n11222_));
  NOR2_X1    g10220(.A1(new_n11213_), .A2(new_n11214_), .ZN(new_n11223_));
  NOR2_X1    g10221(.A1(new_n11196_), .A2(new_n11199_), .ZN(new_n11224_));
  NOR2_X1    g10222(.A1(new_n11223_), .A2(new_n11224_), .ZN(new_n11225_));
  NOR2_X1    g10223(.A1(new_n11137_), .A2(new_n11148_), .ZN(new_n11226_));
  NOR2_X1    g10224(.A1(new_n11226_), .A2(new_n11169_), .ZN(new_n11227_));
  NOR2_X1    g10225(.A1(new_n11184_), .A2(new_n11195_), .ZN(new_n11228_));
  NOR2_X1    g10226(.A1(new_n11228_), .A2(new_n11213_), .ZN(new_n11229_));
  NAND2_X1   g10227(.A1(new_n11227_), .A2(new_n11229_), .ZN(new_n11230_));
  NOR2_X1    g10228(.A1(new_n11230_), .A2(new_n11225_), .ZN(new_n11231_));
  NOR3_X1    g10229(.A1(new_n11231_), .A2(new_n11222_), .A3(new_n11173_), .ZN(new_n11232_));
  INV_X1     g10230(.I(new_n11232_), .ZN(new_n11233_));
  INV_X1     g10231(.I(new_n11197_), .ZN(new_n11234_));
  INV_X1     g10232(.I(new_n11198_), .ZN(new_n11235_));
  NOR2_X1    g10233(.A1(new_n11234_), .A2(new_n11235_), .ZN(new_n11236_));
  NOR4_X1    g10234(.A1(new_n11218_), .A2(new_n11200_), .A3(new_n11228_), .A4(new_n11236_), .ZN(new_n11237_));
  OAI21_X1   g10235(.A1(new_n11222_), .A2(new_n11237_), .B(new_n11173_), .ZN(new_n11238_));
  NAND2_X1   g10236(.A1(new_n11233_), .A2(new_n11238_), .ZN(new_n11239_));
  NAND2_X1   g10237(.A1(new_n11229_), .A2(new_n11218_), .ZN(new_n11240_));
  NAND2_X1   g10238(.A1(new_n11227_), .A2(new_n11220_), .ZN(new_n11241_));
  INV_X1     g10239(.I(\A[807] ), .ZN(new_n11242_));
  NOR2_X1    g10240(.A1(new_n11242_), .A2(\A[806] ), .ZN(new_n11243_));
  INV_X1     g10241(.I(\A[806] ), .ZN(new_n11244_));
  NOR2_X1    g10242(.A1(new_n11244_), .A2(\A[807] ), .ZN(new_n11245_));
  OAI21_X1   g10243(.A1(new_n11243_), .A2(new_n11245_), .B(\A[805] ), .ZN(new_n11246_));
  INV_X1     g10244(.I(\A[805] ), .ZN(new_n11247_));
  NOR2_X1    g10245(.A1(\A[806] ), .A2(\A[807] ), .ZN(new_n11248_));
  NAND2_X1   g10246(.A1(\A[806] ), .A2(\A[807] ), .ZN(new_n11249_));
  INV_X1     g10247(.I(new_n11249_), .ZN(new_n11250_));
  OAI21_X1   g10248(.A1(new_n11250_), .A2(new_n11248_), .B(new_n11247_), .ZN(new_n11251_));
  NAND2_X1   g10249(.A1(new_n11246_), .A2(new_n11251_), .ZN(new_n11252_));
  INV_X1     g10250(.I(\A[810] ), .ZN(new_n11253_));
  NOR2_X1    g10251(.A1(new_n11253_), .A2(\A[809] ), .ZN(new_n11254_));
  INV_X1     g10252(.I(\A[809] ), .ZN(new_n11255_));
  NOR2_X1    g10253(.A1(new_n11255_), .A2(\A[810] ), .ZN(new_n11256_));
  OAI21_X1   g10254(.A1(new_n11254_), .A2(new_n11256_), .B(\A[808] ), .ZN(new_n11257_));
  INV_X1     g10255(.I(\A[808] ), .ZN(new_n11258_));
  NOR2_X1    g10256(.A1(\A[809] ), .A2(\A[810] ), .ZN(new_n11259_));
  NAND2_X1   g10257(.A1(\A[809] ), .A2(\A[810] ), .ZN(new_n11260_));
  INV_X1     g10258(.I(new_n11260_), .ZN(new_n11261_));
  OAI21_X1   g10259(.A1(new_n11261_), .A2(new_n11259_), .B(new_n11258_), .ZN(new_n11262_));
  NAND2_X1   g10260(.A1(new_n11257_), .A2(new_n11262_), .ZN(new_n11263_));
  NOR2_X1    g10261(.A1(new_n11252_), .A2(new_n11263_), .ZN(new_n11264_));
  NAND2_X1   g10262(.A1(new_n11244_), .A2(\A[807] ), .ZN(new_n11265_));
  NAND2_X1   g10263(.A1(new_n11242_), .A2(\A[806] ), .ZN(new_n11266_));
  AOI21_X1   g10264(.A1(new_n11265_), .A2(new_n11266_), .B(new_n11247_), .ZN(new_n11267_));
  INV_X1     g10265(.I(new_n11248_), .ZN(new_n11268_));
  AOI21_X1   g10266(.A1(new_n11268_), .A2(new_n11249_), .B(\A[805] ), .ZN(new_n11269_));
  NOR2_X1    g10267(.A1(new_n11269_), .A2(new_n11267_), .ZN(new_n11270_));
  NAND2_X1   g10268(.A1(new_n11255_), .A2(\A[810] ), .ZN(new_n11271_));
  NAND2_X1   g10269(.A1(new_n11253_), .A2(\A[809] ), .ZN(new_n11272_));
  AOI21_X1   g10270(.A1(new_n11271_), .A2(new_n11272_), .B(new_n11258_), .ZN(new_n11273_));
  INV_X1     g10271(.I(new_n11259_), .ZN(new_n11274_));
  AOI21_X1   g10272(.A1(new_n11274_), .A2(new_n11260_), .B(\A[808] ), .ZN(new_n11275_));
  NOR2_X1    g10273(.A1(new_n11275_), .A2(new_n11273_), .ZN(new_n11276_));
  NOR2_X1    g10274(.A1(new_n11270_), .A2(new_n11276_), .ZN(new_n11277_));
  NOR2_X1    g10275(.A1(new_n11277_), .A2(new_n11264_), .ZN(new_n11278_));
  INV_X1     g10276(.I(\A[799] ), .ZN(new_n11279_));
  INV_X1     g10277(.I(\A[800] ), .ZN(new_n11280_));
  NAND2_X1   g10278(.A1(new_n11280_), .A2(\A[801] ), .ZN(new_n11281_));
  INV_X1     g10279(.I(\A[801] ), .ZN(new_n11282_));
  NAND2_X1   g10280(.A1(new_n11282_), .A2(\A[800] ), .ZN(new_n11283_));
  AOI21_X1   g10281(.A1(new_n11281_), .A2(new_n11283_), .B(new_n11279_), .ZN(new_n11284_));
  NAND2_X1   g10282(.A1(\A[800] ), .A2(\A[801] ), .ZN(new_n11285_));
  NOR2_X1    g10283(.A1(\A[800] ), .A2(\A[801] ), .ZN(new_n11286_));
  INV_X1     g10284(.I(new_n11286_), .ZN(new_n11287_));
  AOI21_X1   g10285(.A1(new_n11287_), .A2(new_n11285_), .B(\A[799] ), .ZN(new_n11288_));
  INV_X1     g10286(.I(\A[802] ), .ZN(new_n11289_));
  INV_X1     g10287(.I(\A[803] ), .ZN(new_n11290_));
  NAND2_X1   g10288(.A1(new_n11290_), .A2(\A[804] ), .ZN(new_n11291_));
  INV_X1     g10289(.I(\A[804] ), .ZN(new_n11292_));
  NAND2_X1   g10290(.A1(new_n11292_), .A2(\A[803] ), .ZN(new_n11293_));
  AOI21_X1   g10291(.A1(new_n11291_), .A2(new_n11293_), .B(new_n11289_), .ZN(new_n11294_));
  NAND2_X1   g10292(.A1(\A[803] ), .A2(\A[804] ), .ZN(new_n11295_));
  NOR2_X1    g10293(.A1(\A[803] ), .A2(\A[804] ), .ZN(new_n11296_));
  INV_X1     g10294(.I(new_n11296_), .ZN(new_n11297_));
  AOI21_X1   g10295(.A1(new_n11297_), .A2(new_n11295_), .B(\A[802] ), .ZN(new_n11298_));
  NOR4_X1    g10296(.A1(new_n11284_), .A2(new_n11288_), .A3(new_n11298_), .A4(new_n11294_), .ZN(new_n11299_));
  NOR2_X1    g10297(.A1(new_n11288_), .A2(new_n11284_), .ZN(new_n11300_));
  NOR2_X1    g10298(.A1(new_n11298_), .A2(new_n11294_), .ZN(new_n11301_));
  NOR2_X1    g10299(.A1(new_n11300_), .A2(new_n11301_), .ZN(new_n11302_));
  OAI21_X1   g10300(.A1(new_n11299_), .A2(new_n11302_), .B(new_n11278_), .ZN(new_n11303_));
  NAND2_X1   g10301(.A1(new_n11270_), .A2(new_n11276_), .ZN(new_n11304_));
  NAND2_X1   g10302(.A1(new_n11252_), .A2(new_n11263_), .ZN(new_n11305_));
  NAND2_X1   g10303(.A1(new_n11304_), .A2(new_n11305_), .ZN(new_n11306_));
  NOR2_X1    g10304(.A1(new_n11302_), .A2(new_n11299_), .ZN(new_n11307_));
  NAND2_X1   g10305(.A1(new_n11306_), .A2(new_n11307_), .ZN(new_n11308_));
  AOI22_X1   g10306(.A1(new_n11303_), .A2(new_n11308_), .B1(new_n11240_), .B2(new_n11241_), .ZN(new_n11309_));
  AOI21_X1   g10307(.A1(new_n11289_), .A2(new_n11295_), .B(new_n11296_), .ZN(new_n11310_));
  AOI21_X1   g10308(.A1(new_n11279_), .A2(new_n11285_), .B(new_n11286_), .ZN(new_n11311_));
  XOR2_X1    g10309(.A1(new_n11310_), .A2(new_n11311_), .Z(new_n11312_));
  XNOR2_X1   g10310(.A1(new_n11312_), .A2(new_n11299_), .ZN(new_n11313_));
  AOI21_X1   g10311(.A1(new_n11258_), .A2(new_n11260_), .B(new_n11259_), .ZN(new_n11314_));
  AOI21_X1   g10312(.A1(new_n11247_), .A2(new_n11249_), .B(new_n11248_), .ZN(new_n11315_));
  XOR2_X1    g10313(.A1(new_n11314_), .A2(new_n11315_), .Z(new_n11316_));
  XOR2_X1    g10314(.A1(new_n11304_), .A2(new_n11316_), .Z(new_n11317_));
  NAND2_X1   g10315(.A1(new_n11278_), .A2(new_n11307_), .ZN(new_n11318_));
  AOI21_X1   g10316(.A1(new_n11318_), .A2(new_n11317_), .B(new_n11313_), .ZN(new_n11319_));
  XOR2_X1    g10317(.A1(new_n11264_), .A2(new_n11316_), .Z(new_n11320_));
  NOR3_X1    g10318(.A1(new_n11306_), .A2(new_n11299_), .A3(new_n11302_), .ZN(new_n11321_));
  NAND2_X1   g10319(.A1(new_n11320_), .A2(new_n11321_), .ZN(new_n11322_));
  NAND2_X1   g10320(.A1(new_n11319_), .A2(new_n11322_), .ZN(new_n11323_));
  NOR2_X1    g10321(.A1(new_n11320_), .A2(new_n11321_), .ZN(new_n11324_));
  NOR2_X1    g10322(.A1(new_n11317_), .A2(new_n11318_), .ZN(new_n11325_));
  OAI21_X1   g10323(.A1(new_n11324_), .A2(new_n11325_), .B(new_n11313_), .ZN(new_n11326_));
  NAND3_X1   g10324(.A1(new_n11323_), .A2(new_n11326_), .A3(new_n11309_), .ZN(new_n11327_));
  NAND2_X1   g10325(.A1(new_n11240_), .A2(new_n11241_), .ZN(new_n11328_));
  NAND2_X1   g10326(.A1(new_n11303_), .A2(new_n11308_), .ZN(new_n11329_));
  NAND2_X1   g10327(.A1(new_n11329_), .A2(new_n11328_), .ZN(new_n11330_));
  XOR2_X1    g10328(.A1(new_n11312_), .A2(new_n11299_), .Z(new_n11331_));
  OAI21_X1   g10329(.A1(new_n11320_), .A2(new_n11321_), .B(new_n11331_), .ZN(new_n11332_));
  NOR2_X1    g10330(.A1(new_n11332_), .A2(new_n11325_), .ZN(new_n11333_));
  NAND2_X1   g10331(.A1(new_n11317_), .A2(new_n11318_), .ZN(new_n11334_));
  AOI21_X1   g10332(.A1(new_n11322_), .A2(new_n11334_), .B(new_n11331_), .ZN(new_n11335_));
  OAI21_X1   g10333(.A1(new_n11335_), .A2(new_n11333_), .B(new_n11330_), .ZN(new_n11336_));
  NAND3_X1   g10334(.A1(new_n11239_), .A2(new_n11327_), .A3(new_n11336_), .ZN(new_n11337_));
  INV_X1     g10335(.I(new_n11238_), .ZN(new_n11338_));
  NOR2_X1    g10336(.A1(new_n11338_), .A2(new_n11232_), .ZN(new_n11339_));
  NOR3_X1    g10337(.A1(new_n11335_), .A2(new_n11333_), .A3(new_n11330_), .ZN(new_n11340_));
  AOI21_X1   g10338(.A1(new_n11323_), .A2(new_n11326_), .B(new_n11309_), .ZN(new_n11341_));
  OAI21_X1   g10339(.A1(new_n11340_), .A2(new_n11341_), .B(new_n11339_), .ZN(new_n11342_));
  NAND2_X1   g10340(.A1(new_n11342_), .A2(new_n11337_), .ZN(new_n11343_));
  INV_X1     g10341(.I(\A[837] ), .ZN(new_n11344_));
  NOR2_X1    g10342(.A1(new_n11344_), .A2(\A[836] ), .ZN(new_n11345_));
  INV_X1     g10343(.I(\A[836] ), .ZN(new_n11346_));
  NOR2_X1    g10344(.A1(new_n11346_), .A2(\A[837] ), .ZN(new_n11347_));
  OAI21_X1   g10345(.A1(new_n11345_), .A2(new_n11347_), .B(\A[835] ), .ZN(new_n11348_));
  INV_X1     g10346(.I(\A[835] ), .ZN(new_n11349_));
  NAND2_X1   g10347(.A1(\A[836] ), .A2(\A[837] ), .ZN(new_n11350_));
  INV_X1     g10348(.I(new_n11350_), .ZN(new_n11351_));
  NOR2_X1    g10349(.A1(\A[836] ), .A2(\A[837] ), .ZN(new_n11352_));
  OAI21_X1   g10350(.A1(new_n11351_), .A2(new_n11352_), .B(new_n11349_), .ZN(new_n11353_));
  NAND2_X1   g10351(.A1(new_n11348_), .A2(new_n11353_), .ZN(new_n11354_));
  INV_X1     g10352(.I(\A[840] ), .ZN(new_n11355_));
  NOR2_X1    g10353(.A1(new_n11355_), .A2(\A[839] ), .ZN(new_n11356_));
  INV_X1     g10354(.I(\A[839] ), .ZN(new_n11357_));
  NOR2_X1    g10355(.A1(new_n11357_), .A2(\A[840] ), .ZN(new_n11358_));
  OAI21_X1   g10356(.A1(new_n11356_), .A2(new_n11358_), .B(\A[838] ), .ZN(new_n11359_));
  INV_X1     g10357(.I(\A[838] ), .ZN(new_n11360_));
  NAND2_X1   g10358(.A1(\A[839] ), .A2(\A[840] ), .ZN(new_n11361_));
  INV_X1     g10359(.I(new_n11361_), .ZN(new_n11362_));
  NOR2_X1    g10360(.A1(\A[839] ), .A2(\A[840] ), .ZN(new_n11363_));
  OAI21_X1   g10361(.A1(new_n11362_), .A2(new_n11363_), .B(new_n11360_), .ZN(new_n11364_));
  NAND2_X1   g10362(.A1(new_n11359_), .A2(new_n11364_), .ZN(new_n11365_));
  NOR2_X1    g10363(.A1(new_n11354_), .A2(new_n11365_), .ZN(new_n11366_));
  NAND2_X1   g10364(.A1(new_n11346_), .A2(\A[837] ), .ZN(new_n11367_));
  NAND2_X1   g10365(.A1(new_n11344_), .A2(\A[836] ), .ZN(new_n11368_));
  AOI21_X1   g10366(.A1(new_n11367_), .A2(new_n11368_), .B(new_n11349_), .ZN(new_n11369_));
  INV_X1     g10367(.I(new_n11352_), .ZN(new_n11370_));
  AOI21_X1   g10368(.A1(new_n11370_), .A2(new_n11350_), .B(\A[835] ), .ZN(new_n11371_));
  NOR2_X1    g10369(.A1(new_n11371_), .A2(new_n11369_), .ZN(new_n11372_));
  NAND2_X1   g10370(.A1(new_n11357_), .A2(\A[840] ), .ZN(new_n11373_));
  NAND2_X1   g10371(.A1(new_n11355_), .A2(\A[839] ), .ZN(new_n11374_));
  AOI21_X1   g10372(.A1(new_n11373_), .A2(new_n11374_), .B(new_n11360_), .ZN(new_n11375_));
  INV_X1     g10373(.I(new_n11363_), .ZN(new_n11376_));
  AOI21_X1   g10374(.A1(new_n11376_), .A2(new_n11361_), .B(\A[838] ), .ZN(new_n11377_));
  NOR2_X1    g10375(.A1(new_n11377_), .A2(new_n11375_), .ZN(new_n11378_));
  NOR2_X1    g10376(.A1(new_n11372_), .A2(new_n11378_), .ZN(new_n11379_));
  NOR2_X1    g10377(.A1(new_n11379_), .A2(new_n11366_), .ZN(new_n11380_));
  INV_X1     g10378(.I(\A[841] ), .ZN(new_n11381_));
  INV_X1     g10379(.I(\A[842] ), .ZN(new_n11382_));
  NAND2_X1   g10380(.A1(new_n11382_), .A2(\A[843] ), .ZN(new_n11383_));
  INV_X1     g10381(.I(\A[843] ), .ZN(new_n11384_));
  NAND2_X1   g10382(.A1(new_n11384_), .A2(\A[842] ), .ZN(new_n11385_));
  AOI21_X1   g10383(.A1(new_n11383_), .A2(new_n11385_), .B(new_n11381_), .ZN(new_n11386_));
  NAND2_X1   g10384(.A1(\A[842] ), .A2(\A[843] ), .ZN(new_n11387_));
  NOR2_X1    g10385(.A1(\A[842] ), .A2(\A[843] ), .ZN(new_n11388_));
  INV_X1     g10386(.I(new_n11388_), .ZN(new_n11389_));
  AOI21_X1   g10387(.A1(new_n11389_), .A2(new_n11387_), .B(\A[841] ), .ZN(new_n11390_));
  NOR2_X1    g10388(.A1(new_n11390_), .A2(new_n11386_), .ZN(new_n11391_));
  INV_X1     g10389(.I(\A[844] ), .ZN(new_n11392_));
  INV_X1     g10390(.I(\A[845] ), .ZN(new_n11393_));
  NAND2_X1   g10391(.A1(new_n11393_), .A2(\A[846] ), .ZN(new_n11394_));
  INV_X1     g10392(.I(\A[846] ), .ZN(new_n11395_));
  NAND2_X1   g10393(.A1(new_n11395_), .A2(\A[845] ), .ZN(new_n11396_));
  AOI21_X1   g10394(.A1(new_n11394_), .A2(new_n11396_), .B(new_n11392_), .ZN(new_n11397_));
  NAND2_X1   g10395(.A1(\A[845] ), .A2(\A[846] ), .ZN(new_n11398_));
  NOR2_X1    g10396(.A1(\A[845] ), .A2(\A[846] ), .ZN(new_n11399_));
  INV_X1     g10397(.I(new_n11399_), .ZN(new_n11400_));
  AOI21_X1   g10398(.A1(new_n11400_), .A2(new_n11398_), .B(\A[844] ), .ZN(new_n11401_));
  NOR2_X1    g10399(.A1(new_n11401_), .A2(new_n11397_), .ZN(new_n11402_));
  NAND2_X1   g10400(.A1(new_n11391_), .A2(new_n11402_), .ZN(new_n11403_));
  NOR2_X1    g10401(.A1(new_n11384_), .A2(\A[842] ), .ZN(new_n11404_));
  NOR2_X1    g10402(.A1(new_n11382_), .A2(\A[843] ), .ZN(new_n11405_));
  OAI21_X1   g10403(.A1(new_n11404_), .A2(new_n11405_), .B(\A[841] ), .ZN(new_n11406_));
  INV_X1     g10404(.I(new_n11387_), .ZN(new_n11407_));
  OAI21_X1   g10405(.A1(new_n11407_), .A2(new_n11388_), .B(new_n11381_), .ZN(new_n11408_));
  NAND2_X1   g10406(.A1(new_n11406_), .A2(new_n11408_), .ZN(new_n11409_));
  NOR2_X1    g10407(.A1(new_n11395_), .A2(\A[845] ), .ZN(new_n11410_));
  NOR2_X1    g10408(.A1(new_n11393_), .A2(\A[846] ), .ZN(new_n11411_));
  OAI21_X1   g10409(.A1(new_n11410_), .A2(new_n11411_), .B(\A[844] ), .ZN(new_n11412_));
  INV_X1     g10410(.I(new_n11398_), .ZN(new_n11413_));
  OAI21_X1   g10411(.A1(new_n11413_), .A2(new_n11399_), .B(new_n11392_), .ZN(new_n11414_));
  NAND2_X1   g10412(.A1(new_n11412_), .A2(new_n11414_), .ZN(new_n11415_));
  NAND2_X1   g10413(.A1(new_n11409_), .A2(new_n11415_), .ZN(new_n11416_));
  NAND2_X1   g10414(.A1(new_n11403_), .A2(new_n11416_), .ZN(new_n11417_));
  XOR2_X1    g10415(.A1(new_n11380_), .A2(new_n11417_), .Z(new_n11418_));
  INV_X1     g10416(.I(\A[823] ), .ZN(new_n11419_));
  INV_X1     g10417(.I(\A[824] ), .ZN(new_n11420_));
  NAND2_X1   g10418(.A1(new_n11420_), .A2(\A[825] ), .ZN(new_n11421_));
  INV_X1     g10419(.I(\A[825] ), .ZN(new_n11422_));
  NAND2_X1   g10420(.A1(new_n11422_), .A2(\A[824] ), .ZN(new_n11423_));
  AOI21_X1   g10421(.A1(new_n11421_), .A2(new_n11423_), .B(new_n11419_), .ZN(new_n11424_));
  NAND2_X1   g10422(.A1(\A[824] ), .A2(\A[825] ), .ZN(new_n11425_));
  NOR2_X1    g10423(.A1(\A[824] ), .A2(\A[825] ), .ZN(new_n11426_));
  INV_X1     g10424(.I(new_n11426_), .ZN(new_n11427_));
  AOI21_X1   g10425(.A1(new_n11427_), .A2(new_n11425_), .B(\A[823] ), .ZN(new_n11428_));
  INV_X1     g10426(.I(\A[826] ), .ZN(new_n11429_));
  INV_X1     g10427(.I(\A[827] ), .ZN(new_n11430_));
  NAND2_X1   g10428(.A1(new_n11430_), .A2(\A[828] ), .ZN(new_n11431_));
  INV_X1     g10429(.I(\A[828] ), .ZN(new_n11432_));
  NAND2_X1   g10430(.A1(new_n11432_), .A2(\A[827] ), .ZN(new_n11433_));
  AOI21_X1   g10431(.A1(new_n11431_), .A2(new_n11433_), .B(new_n11429_), .ZN(new_n11434_));
  NAND2_X1   g10432(.A1(\A[827] ), .A2(\A[828] ), .ZN(new_n11435_));
  NOR2_X1    g10433(.A1(\A[827] ), .A2(\A[828] ), .ZN(new_n11436_));
  INV_X1     g10434(.I(new_n11436_), .ZN(new_n11437_));
  AOI21_X1   g10435(.A1(new_n11437_), .A2(new_n11435_), .B(\A[826] ), .ZN(new_n11438_));
  NOR4_X1    g10436(.A1(new_n11424_), .A2(new_n11428_), .A3(new_n11438_), .A4(new_n11434_), .ZN(new_n11439_));
  NOR2_X1    g10437(.A1(new_n11428_), .A2(new_n11424_), .ZN(new_n11440_));
  NOR2_X1    g10438(.A1(new_n11438_), .A2(new_n11434_), .ZN(new_n11441_));
  NOR2_X1    g10439(.A1(new_n11440_), .A2(new_n11441_), .ZN(new_n11442_));
  NOR2_X1    g10440(.A1(new_n11442_), .A2(new_n11439_), .ZN(new_n11443_));
  INV_X1     g10441(.I(\A[829] ), .ZN(new_n11444_));
  INV_X1     g10442(.I(\A[830] ), .ZN(new_n11445_));
  NAND2_X1   g10443(.A1(new_n11445_), .A2(\A[831] ), .ZN(new_n11446_));
  INV_X1     g10444(.I(\A[831] ), .ZN(new_n11447_));
  NAND2_X1   g10445(.A1(new_n11447_), .A2(\A[830] ), .ZN(new_n11448_));
  AOI21_X1   g10446(.A1(new_n11446_), .A2(new_n11448_), .B(new_n11444_), .ZN(new_n11449_));
  NAND2_X1   g10447(.A1(\A[830] ), .A2(\A[831] ), .ZN(new_n11450_));
  NOR2_X1    g10448(.A1(\A[830] ), .A2(\A[831] ), .ZN(new_n11451_));
  INV_X1     g10449(.I(new_n11451_), .ZN(new_n11452_));
  AOI21_X1   g10450(.A1(new_n11452_), .A2(new_n11450_), .B(\A[829] ), .ZN(new_n11453_));
  NOR2_X1    g10451(.A1(new_n11453_), .A2(new_n11449_), .ZN(new_n11454_));
  INV_X1     g10452(.I(\A[832] ), .ZN(new_n11455_));
  INV_X1     g10453(.I(\A[833] ), .ZN(new_n11456_));
  NAND2_X1   g10454(.A1(new_n11456_), .A2(\A[834] ), .ZN(new_n11457_));
  INV_X1     g10455(.I(\A[834] ), .ZN(new_n11458_));
  NAND2_X1   g10456(.A1(new_n11458_), .A2(\A[833] ), .ZN(new_n11459_));
  AOI21_X1   g10457(.A1(new_n11457_), .A2(new_n11459_), .B(new_n11455_), .ZN(new_n11460_));
  NAND2_X1   g10458(.A1(\A[833] ), .A2(\A[834] ), .ZN(new_n11461_));
  NOR2_X1    g10459(.A1(\A[833] ), .A2(\A[834] ), .ZN(new_n11462_));
  INV_X1     g10460(.I(new_n11462_), .ZN(new_n11463_));
  AOI21_X1   g10461(.A1(new_n11463_), .A2(new_n11461_), .B(\A[832] ), .ZN(new_n11464_));
  NOR2_X1    g10462(.A1(new_n11464_), .A2(new_n11460_), .ZN(new_n11465_));
  NAND2_X1   g10463(.A1(new_n11454_), .A2(new_n11465_), .ZN(new_n11466_));
  NOR2_X1    g10464(.A1(new_n11447_), .A2(\A[830] ), .ZN(new_n11467_));
  NOR2_X1    g10465(.A1(new_n11445_), .A2(\A[831] ), .ZN(new_n11468_));
  OAI21_X1   g10466(.A1(new_n11467_), .A2(new_n11468_), .B(\A[829] ), .ZN(new_n11469_));
  INV_X1     g10467(.I(new_n11450_), .ZN(new_n11470_));
  OAI21_X1   g10468(.A1(new_n11470_), .A2(new_n11451_), .B(new_n11444_), .ZN(new_n11471_));
  NAND2_X1   g10469(.A1(new_n11469_), .A2(new_n11471_), .ZN(new_n11472_));
  NOR2_X1    g10470(.A1(new_n11458_), .A2(\A[833] ), .ZN(new_n11473_));
  NOR2_X1    g10471(.A1(new_n11456_), .A2(\A[834] ), .ZN(new_n11474_));
  OAI21_X1   g10472(.A1(new_n11473_), .A2(new_n11474_), .B(\A[832] ), .ZN(new_n11475_));
  INV_X1     g10473(.I(new_n11461_), .ZN(new_n11476_));
  OAI21_X1   g10474(.A1(new_n11476_), .A2(new_n11462_), .B(new_n11455_), .ZN(new_n11477_));
  NAND2_X1   g10475(.A1(new_n11475_), .A2(new_n11477_), .ZN(new_n11478_));
  NAND2_X1   g10476(.A1(new_n11472_), .A2(new_n11478_), .ZN(new_n11479_));
  NAND2_X1   g10477(.A1(new_n11466_), .A2(new_n11479_), .ZN(new_n11480_));
  NOR2_X1    g10478(.A1(new_n11480_), .A2(new_n11443_), .ZN(new_n11481_));
  NAND2_X1   g10479(.A1(new_n11440_), .A2(new_n11441_), .ZN(new_n11482_));
  OAI22_X1   g10480(.A1(new_n11424_), .A2(new_n11428_), .B1(new_n11438_), .B2(new_n11434_), .ZN(new_n11483_));
  NAND2_X1   g10481(.A1(new_n11482_), .A2(new_n11483_), .ZN(new_n11484_));
  NOR2_X1    g10482(.A1(new_n11472_), .A2(new_n11478_), .ZN(new_n11485_));
  NOR2_X1    g10483(.A1(new_n11454_), .A2(new_n11465_), .ZN(new_n11486_));
  NOR2_X1    g10484(.A1(new_n11486_), .A2(new_n11485_), .ZN(new_n11487_));
  NOR2_X1    g10485(.A1(new_n11487_), .A2(new_n11484_), .ZN(new_n11488_));
  NOR2_X1    g10486(.A1(new_n11481_), .A2(new_n11488_), .ZN(new_n11489_));
  NOR2_X1    g10487(.A1(new_n11418_), .A2(new_n11489_), .ZN(new_n11490_));
  NAND2_X1   g10488(.A1(new_n11372_), .A2(new_n11378_), .ZN(new_n11491_));
  NAND2_X1   g10489(.A1(new_n11354_), .A2(new_n11365_), .ZN(new_n11492_));
  NAND2_X1   g10490(.A1(new_n11491_), .A2(new_n11492_), .ZN(new_n11493_));
  NOR2_X1    g10491(.A1(new_n11409_), .A2(new_n11415_), .ZN(new_n11494_));
  NOR2_X1    g10492(.A1(new_n11391_), .A2(new_n11402_), .ZN(new_n11495_));
  NOR2_X1    g10493(.A1(new_n11495_), .A2(new_n11494_), .ZN(new_n11496_));
  NAND2_X1   g10494(.A1(new_n11496_), .A2(new_n11493_), .ZN(new_n11497_));
  NAND2_X1   g10495(.A1(new_n11380_), .A2(new_n11417_), .ZN(new_n11498_));
  NAND2_X1   g10496(.A1(new_n11497_), .A2(new_n11498_), .ZN(new_n11499_));
  NAND2_X1   g10497(.A1(new_n11487_), .A2(new_n11484_), .ZN(new_n11500_));
  NAND2_X1   g10498(.A1(new_n11480_), .A2(new_n11443_), .ZN(new_n11501_));
  NAND2_X1   g10499(.A1(new_n11501_), .A2(new_n11500_), .ZN(new_n11502_));
  NOR2_X1    g10500(.A1(new_n11499_), .A2(new_n11502_), .ZN(new_n11503_));
  NOR2_X1    g10501(.A1(new_n11490_), .A2(new_n11503_), .ZN(new_n11504_));
  NOR2_X1    g10502(.A1(new_n11329_), .A2(new_n11328_), .ZN(new_n11505_));
  NOR2_X1    g10503(.A1(new_n11505_), .A2(new_n11309_), .ZN(new_n11506_));
  NAND2_X1   g10504(.A1(new_n11504_), .A2(new_n11506_), .ZN(new_n11507_));
  INV_X1     g10505(.I(new_n11507_), .ZN(new_n11508_));
  AOI21_X1   g10506(.A1(new_n11429_), .A2(new_n11435_), .B(new_n11436_), .ZN(new_n11509_));
  AOI21_X1   g10507(.A1(new_n11419_), .A2(new_n11425_), .B(new_n11426_), .ZN(new_n11510_));
  NOR2_X1    g10508(.A1(new_n11509_), .A2(new_n11510_), .ZN(new_n11511_));
  INV_X1     g10509(.I(new_n11511_), .ZN(new_n11512_));
  NAND2_X1   g10510(.A1(new_n11509_), .A2(new_n11510_), .ZN(new_n11513_));
  NAND2_X1   g10511(.A1(new_n11512_), .A2(new_n11513_), .ZN(new_n11514_));
  NOR2_X1    g10512(.A1(new_n11514_), .A2(new_n11439_), .ZN(new_n11515_));
  AOI21_X1   g10513(.A1(new_n11512_), .A2(new_n11513_), .B(new_n11482_), .ZN(new_n11516_));
  AOI21_X1   g10514(.A1(new_n11455_), .A2(new_n11461_), .B(new_n11462_), .ZN(new_n11517_));
  AOI21_X1   g10515(.A1(new_n11444_), .A2(new_n11450_), .B(new_n11451_), .ZN(new_n11518_));
  XOR2_X1    g10516(.A1(new_n11517_), .A2(new_n11518_), .Z(new_n11519_));
  NAND2_X1   g10517(.A1(new_n11466_), .A2(new_n11519_), .ZN(new_n11520_));
  XNOR2_X1   g10518(.A1(new_n11517_), .A2(new_n11518_), .ZN(new_n11521_));
  NAND2_X1   g10519(.A1(new_n11485_), .A2(new_n11521_), .ZN(new_n11522_));
  NAND2_X1   g10520(.A1(new_n11522_), .A2(new_n11520_), .ZN(new_n11523_));
  NOR4_X1    g10521(.A1(new_n11442_), .A2(new_n11486_), .A3(new_n11485_), .A4(new_n11439_), .ZN(new_n11524_));
  OAI22_X1   g10522(.A1(new_n11523_), .A2(new_n11524_), .B1(new_n11515_), .B2(new_n11516_), .ZN(new_n11525_));
  NOR2_X1    g10523(.A1(new_n11485_), .A2(new_n11521_), .ZN(new_n11526_));
  NAND2_X1   g10524(.A1(new_n11517_), .A2(new_n11518_), .ZN(new_n11527_));
  NAND4_X1   g10525(.A1(new_n11526_), .A2(new_n11443_), .A3(new_n11479_), .A4(new_n11527_), .ZN(new_n11528_));
  INV_X1     g10526(.I(new_n11528_), .ZN(new_n11529_));
  NOR2_X1    g10527(.A1(new_n11525_), .A2(new_n11529_), .ZN(new_n11530_));
  INV_X1     g10528(.I(new_n11515_), .ZN(new_n11531_));
  NAND2_X1   g10529(.A1(new_n11514_), .A2(new_n11439_), .ZN(new_n11532_));
  NAND2_X1   g10530(.A1(new_n11531_), .A2(new_n11532_), .ZN(new_n11533_));
  NOR2_X1    g10531(.A1(new_n11466_), .A2(new_n11519_), .ZN(new_n11534_));
  NOR2_X1    g10532(.A1(new_n11526_), .A2(new_n11534_), .ZN(new_n11535_));
  NAND2_X1   g10533(.A1(new_n11487_), .A2(new_n11443_), .ZN(new_n11536_));
  NAND2_X1   g10534(.A1(new_n11535_), .A2(new_n11536_), .ZN(new_n11537_));
  NAND2_X1   g10535(.A1(new_n11523_), .A2(new_n11524_), .ZN(new_n11538_));
  AOI21_X1   g10536(.A1(new_n11537_), .A2(new_n11538_), .B(new_n11533_), .ZN(new_n11539_));
  OR2_X2     g10537(.A1(new_n11530_), .A2(new_n11539_), .Z(new_n11540_));
  AOI21_X1   g10538(.A1(new_n11360_), .A2(new_n11361_), .B(new_n11363_), .ZN(new_n11541_));
  AOI21_X1   g10539(.A1(new_n11349_), .A2(new_n11350_), .B(new_n11352_), .ZN(new_n11542_));
  NOR2_X1    g10540(.A1(new_n11541_), .A2(new_n11542_), .ZN(new_n11543_));
  INV_X1     g10541(.I(new_n11543_), .ZN(new_n11544_));
  NAND2_X1   g10542(.A1(new_n11541_), .A2(new_n11542_), .ZN(new_n11545_));
  NAND3_X1   g10543(.A1(new_n11491_), .A2(new_n11544_), .A3(new_n11545_), .ZN(new_n11546_));
  NAND2_X1   g10544(.A1(new_n11544_), .A2(new_n11545_), .ZN(new_n11547_));
  NAND2_X1   g10545(.A1(new_n11547_), .A2(new_n11366_), .ZN(new_n11548_));
  NAND2_X1   g10546(.A1(new_n11548_), .A2(new_n11546_), .ZN(new_n11549_));
  INV_X1     g10547(.I(new_n11549_), .ZN(new_n11550_));
  AOI21_X1   g10548(.A1(new_n11392_), .A2(new_n11398_), .B(new_n11399_), .ZN(new_n11551_));
  AOI21_X1   g10549(.A1(new_n11381_), .A2(new_n11387_), .B(new_n11388_), .ZN(new_n11552_));
  XOR2_X1    g10550(.A1(new_n11551_), .A2(new_n11552_), .Z(new_n11553_));
  NAND2_X1   g10551(.A1(new_n11403_), .A2(new_n11553_), .ZN(new_n11554_));
  XNOR2_X1   g10552(.A1(new_n11551_), .A2(new_n11552_), .ZN(new_n11555_));
  NAND2_X1   g10553(.A1(new_n11494_), .A2(new_n11555_), .ZN(new_n11556_));
  NAND4_X1   g10554(.A1(new_n11491_), .A2(new_n11492_), .A3(new_n11403_), .A4(new_n11416_), .ZN(new_n11557_));
  NAND3_X1   g10555(.A1(new_n11557_), .A2(new_n11554_), .A3(new_n11556_), .ZN(new_n11558_));
  NAND4_X1   g10556(.A1(new_n11380_), .A2(new_n11403_), .A3(new_n11416_), .A4(new_n11553_), .ZN(new_n11559_));
  AND3_X2    g10557(.A1(new_n11550_), .A2(new_n11558_), .A3(new_n11559_), .Z(new_n11560_));
  INV_X1     g10558(.I(new_n11551_), .ZN(new_n11561_));
  INV_X1     g10559(.I(new_n11552_), .ZN(new_n11562_));
  NOR2_X1    g10560(.A1(new_n11561_), .A2(new_n11562_), .ZN(new_n11563_));
  NOR4_X1    g10561(.A1(new_n11493_), .A2(new_n11554_), .A3(new_n11495_), .A4(new_n11563_), .ZN(new_n11564_));
  INV_X1     g10562(.I(new_n11564_), .ZN(new_n11565_));
  AOI21_X1   g10563(.A1(new_n11565_), .A2(new_n11558_), .B(new_n11550_), .ZN(new_n11566_));
  OAI21_X1   g10564(.A1(new_n11560_), .A2(new_n11566_), .B(new_n11490_), .ZN(new_n11567_));
  NAND2_X1   g10565(.A1(new_n11499_), .A2(new_n11502_), .ZN(new_n11568_));
  NAND3_X1   g10566(.A1(new_n11550_), .A2(new_n11558_), .A3(new_n11559_), .ZN(new_n11569_));
  INV_X1     g10567(.I(new_n11558_), .ZN(new_n11570_));
  OAI21_X1   g10568(.A1(new_n11570_), .A2(new_n11564_), .B(new_n11549_), .ZN(new_n11571_));
  NAND3_X1   g10569(.A1(new_n11571_), .A2(new_n11568_), .A3(new_n11569_), .ZN(new_n11572_));
  AOI21_X1   g10570(.A1(new_n11567_), .A2(new_n11572_), .B(new_n11540_), .ZN(new_n11573_));
  NOR2_X1    g10571(.A1(new_n11530_), .A2(new_n11539_), .ZN(new_n11574_));
  AOI21_X1   g10572(.A1(new_n11571_), .A2(new_n11569_), .B(new_n11568_), .ZN(new_n11575_));
  NOR3_X1    g10573(.A1(new_n11560_), .A2(new_n11490_), .A3(new_n11566_), .ZN(new_n11576_));
  NOR3_X1    g10574(.A1(new_n11576_), .A2(new_n11575_), .A3(new_n11574_), .ZN(new_n11577_));
  OAI21_X1   g10575(.A1(new_n11573_), .A2(new_n11577_), .B(new_n11508_), .ZN(new_n11578_));
  NOR3_X1    g10576(.A1(new_n11573_), .A2(new_n11508_), .A3(new_n11577_), .ZN(new_n11579_));
  AOI21_X1   g10577(.A1(new_n11343_), .A2(new_n11578_), .B(new_n11579_), .ZN(new_n11580_));
  AOI22_X1   g10578(.A1(new_n11230_), .A2(new_n11225_), .B1(new_n11156_), .B2(new_n11172_), .ZN(new_n11581_));
  INV_X1     g10579(.I(new_n11236_), .ZN(new_n11582_));
  NOR2_X1    g10580(.A1(new_n11197_), .A2(new_n11198_), .ZN(new_n11583_));
  AOI21_X1   g10581(.A1(new_n11196_), .A2(new_n11582_), .B(new_n11583_), .ZN(new_n11584_));
  AOI21_X1   g10582(.A1(new_n11149_), .A2(new_n11153_), .B(new_n11152_), .ZN(new_n11585_));
  NOR2_X1    g10583(.A1(new_n11584_), .A2(new_n11585_), .ZN(new_n11586_));
  INV_X1     g10584(.I(new_n11583_), .ZN(new_n11587_));
  OAI21_X1   g10585(.A1(new_n11213_), .A2(new_n11236_), .B(new_n11587_), .ZN(new_n11588_));
  OAI21_X1   g10586(.A1(new_n11169_), .A2(new_n11154_), .B(new_n11170_), .ZN(new_n11589_));
  NOR2_X1    g10587(.A1(new_n11588_), .A2(new_n11589_), .ZN(new_n11590_));
  NOR2_X1    g10588(.A1(new_n11586_), .A2(new_n11590_), .ZN(new_n11591_));
  OAI21_X1   g10589(.A1(new_n11581_), .A2(new_n11237_), .B(new_n11591_), .ZN(new_n11592_));
  INV_X1     g10590(.I(new_n11237_), .ZN(new_n11593_));
  OAI21_X1   g10591(.A1(new_n11216_), .A2(new_n11221_), .B(new_n11173_), .ZN(new_n11594_));
  NAND2_X1   g10592(.A1(new_n11588_), .A2(new_n11589_), .ZN(new_n11595_));
  NAND2_X1   g10593(.A1(new_n11584_), .A2(new_n11585_), .ZN(new_n11596_));
  NAND2_X1   g10594(.A1(new_n11596_), .A2(new_n11595_), .ZN(new_n11597_));
  NAND3_X1   g10595(.A1(new_n11594_), .A2(new_n11597_), .A3(new_n11593_), .ZN(new_n11598_));
  NAND2_X1   g10596(.A1(new_n11592_), .A2(new_n11598_), .ZN(new_n11599_));
  AND2_X2    g10597(.A1(new_n11314_), .A2(new_n11315_), .Z(new_n11600_));
  NOR2_X1    g10598(.A1(new_n11314_), .A2(new_n11315_), .ZN(new_n11601_));
  INV_X1     g10599(.I(new_n11601_), .ZN(new_n11602_));
  OAI21_X1   g10600(.A1(new_n11264_), .A2(new_n11600_), .B(new_n11602_), .ZN(new_n11603_));
  INV_X1     g10601(.I(new_n11299_), .ZN(new_n11604_));
  NOR2_X1    g10602(.A1(new_n11310_), .A2(new_n11311_), .ZN(new_n11605_));
  NAND2_X1   g10603(.A1(new_n11310_), .A2(new_n11311_), .ZN(new_n11606_));
  AOI21_X1   g10604(.A1(new_n11604_), .A2(new_n11606_), .B(new_n11605_), .ZN(new_n11607_));
  NOR3_X1    g10605(.A1(new_n11319_), .A2(new_n11325_), .A3(new_n11607_), .ZN(new_n11608_));
  INV_X1     g10606(.I(new_n11607_), .ZN(new_n11609_));
  AOI21_X1   g10607(.A1(new_n11332_), .A2(new_n11322_), .B(new_n11609_), .ZN(new_n11610_));
  NOR3_X1    g10608(.A1(new_n11608_), .A2(new_n11610_), .A3(new_n11603_), .ZN(new_n11611_));
  INV_X1     g10609(.I(new_n11603_), .ZN(new_n11612_));
  NAND3_X1   g10610(.A1(new_n11332_), .A2(new_n11322_), .A3(new_n11609_), .ZN(new_n11613_));
  OAI21_X1   g10611(.A1(new_n11319_), .A2(new_n11325_), .B(new_n11607_), .ZN(new_n11614_));
  AOI21_X1   g10612(.A1(new_n11614_), .A2(new_n11613_), .B(new_n11612_), .ZN(new_n11615_));
  OAI21_X1   g10613(.A1(new_n11611_), .A2(new_n11615_), .B(new_n11599_), .ZN(new_n11616_));
  AOI21_X1   g10614(.A1(new_n11594_), .A2(new_n11593_), .B(new_n11597_), .ZN(new_n11617_));
  NOR3_X1    g10615(.A1(new_n11581_), .A2(new_n11591_), .A3(new_n11237_), .ZN(new_n11618_));
  NOR2_X1    g10616(.A1(new_n11618_), .A2(new_n11617_), .ZN(new_n11619_));
  NAND3_X1   g10617(.A1(new_n11614_), .A2(new_n11613_), .A3(new_n11612_), .ZN(new_n11620_));
  OAI21_X1   g10618(.A1(new_n11608_), .A2(new_n11610_), .B(new_n11603_), .ZN(new_n11621_));
  NAND3_X1   g10619(.A1(new_n11621_), .A2(new_n11620_), .A3(new_n11619_), .ZN(new_n11622_));
  OAI21_X1   g10620(.A1(new_n11239_), .A2(new_n11340_), .B(new_n11336_), .ZN(new_n11623_));
  NAND3_X1   g10621(.A1(new_n11616_), .A2(new_n11623_), .A3(new_n11622_), .ZN(new_n11624_));
  AOI21_X1   g10622(.A1(new_n11621_), .A2(new_n11620_), .B(new_n11619_), .ZN(new_n11625_));
  NOR3_X1    g10623(.A1(new_n11611_), .A2(new_n11615_), .A3(new_n11599_), .ZN(new_n11626_));
  AOI21_X1   g10624(.A1(new_n11339_), .A2(new_n11327_), .B(new_n11341_), .ZN(new_n11627_));
  OAI21_X1   g10625(.A1(new_n11625_), .A2(new_n11626_), .B(new_n11627_), .ZN(new_n11628_));
  OAI21_X1   g10626(.A1(new_n11574_), .A2(new_n11575_), .B(new_n11572_), .ZN(new_n11629_));
  NOR2_X1    g10627(.A1(new_n11494_), .A2(new_n11555_), .ZN(new_n11630_));
  NOR2_X1    g10628(.A1(new_n11403_), .A2(new_n11553_), .ZN(new_n11631_));
  NOR2_X1    g10629(.A1(new_n11630_), .A2(new_n11631_), .ZN(new_n11632_));
  AOI22_X1   g10630(.A1(new_n11632_), .A2(new_n11557_), .B1(new_n11546_), .B2(new_n11548_), .ZN(new_n11633_));
  INV_X1     g10631(.I(new_n11563_), .ZN(new_n11634_));
  NOR2_X1    g10632(.A1(new_n11551_), .A2(new_n11552_), .ZN(new_n11635_));
  AOI21_X1   g10633(.A1(new_n11403_), .A2(new_n11634_), .B(new_n11635_), .ZN(new_n11636_));
  AOI21_X1   g10634(.A1(new_n11491_), .A2(new_n11545_), .B(new_n11543_), .ZN(new_n11637_));
  NOR2_X1    g10635(.A1(new_n11636_), .A2(new_n11637_), .ZN(new_n11638_));
  INV_X1     g10636(.I(new_n11635_), .ZN(new_n11639_));
  OAI21_X1   g10637(.A1(new_n11494_), .A2(new_n11563_), .B(new_n11639_), .ZN(new_n11640_));
  INV_X1     g10638(.I(new_n11545_), .ZN(new_n11641_));
  OAI21_X1   g10639(.A1(new_n11366_), .A2(new_n11641_), .B(new_n11544_), .ZN(new_n11642_));
  NOR2_X1    g10640(.A1(new_n11640_), .A2(new_n11642_), .ZN(new_n11643_));
  NOR2_X1    g10641(.A1(new_n11638_), .A2(new_n11643_), .ZN(new_n11644_));
  OAI21_X1   g10642(.A1(new_n11633_), .A2(new_n11564_), .B(new_n11644_), .ZN(new_n11645_));
  AOI21_X1   g10643(.A1(new_n11558_), .A2(new_n11549_), .B(new_n11564_), .ZN(new_n11646_));
  NAND2_X1   g10644(.A1(new_n11640_), .A2(new_n11642_), .ZN(new_n11647_));
  NAND2_X1   g10645(.A1(new_n11636_), .A2(new_n11637_), .ZN(new_n11648_));
  NAND2_X1   g10646(.A1(new_n11648_), .A2(new_n11647_), .ZN(new_n11649_));
  NAND2_X1   g10647(.A1(new_n11646_), .A2(new_n11649_), .ZN(new_n11650_));
  NAND2_X1   g10648(.A1(new_n11650_), .A2(new_n11645_), .ZN(new_n11651_));
  NOR2_X1    g10649(.A1(new_n11517_), .A2(new_n11518_), .ZN(new_n11652_));
  AOI21_X1   g10650(.A1(new_n11466_), .A2(new_n11527_), .B(new_n11652_), .ZN(new_n11653_));
  INV_X1     g10651(.I(new_n11653_), .ZN(new_n11654_));
  AOI22_X1   g10652(.A1(new_n11535_), .A2(new_n11536_), .B1(new_n11531_), .B2(new_n11532_), .ZN(new_n11655_));
  AOI21_X1   g10653(.A1(new_n11482_), .A2(new_n11513_), .B(new_n11511_), .ZN(new_n11656_));
  NOR3_X1    g10654(.A1(new_n11655_), .A2(new_n11529_), .A3(new_n11656_), .ZN(new_n11657_));
  INV_X1     g10655(.I(new_n11656_), .ZN(new_n11658_));
  AOI21_X1   g10656(.A1(new_n11525_), .A2(new_n11528_), .B(new_n11658_), .ZN(new_n11659_));
  NOR3_X1    g10657(.A1(new_n11657_), .A2(new_n11659_), .A3(new_n11654_), .ZN(new_n11660_));
  NAND3_X1   g10658(.A1(new_n11525_), .A2(new_n11528_), .A3(new_n11658_), .ZN(new_n11661_));
  OAI21_X1   g10659(.A1(new_n11655_), .A2(new_n11529_), .B(new_n11656_), .ZN(new_n11662_));
  AOI21_X1   g10660(.A1(new_n11662_), .A2(new_n11661_), .B(new_n11653_), .ZN(new_n11663_));
  OAI21_X1   g10661(.A1(new_n11660_), .A2(new_n11663_), .B(new_n11651_), .ZN(new_n11664_));
  NOR2_X1    g10662(.A1(new_n11646_), .A2(new_n11649_), .ZN(new_n11665_));
  NOR3_X1    g10663(.A1(new_n11633_), .A2(new_n11644_), .A3(new_n11564_), .ZN(new_n11666_));
  NOR2_X1    g10664(.A1(new_n11665_), .A2(new_n11666_), .ZN(new_n11667_));
  NAND3_X1   g10665(.A1(new_n11662_), .A2(new_n11661_), .A3(new_n11653_), .ZN(new_n11668_));
  OAI21_X1   g10666(.A1(new_n11657_), .A2(new_n11659_), .B(new_n11654_), .ZN(new_n11669_));
  NAND3_X1   g10667(.A1(new_n11668_), .A2(new_n11669_), .A3(new_n11667_), .ZN(new_n11670_));
  NAND3_X1   g10668(.A1(new_n11664_), .A2(new_n11670_), .A3(new_n11629_), .ZN(new_n11671_));
  AOI21_X1   g10669(.A1(new_n11540_), .A2(new_n11567_), .B(new_n11576_), .ZN(new_n11672_));
  AOI21_X1   g10670(.A1(new_n11668_), .A2(new_n11669_), .B(new_n11667_), .ZN(new_n11673_));
  NOR3_X1    g10671(.A1(new_n11651_), .A2(new_n11660_), .A3(new_n11663_), .ZN(new_n11674_));
  OAI21_X1   g10672(.A1(new_n11674_), .A2(new_n11673_), .B(new_n11672_), .ZN(new_n11675_));
  NAND4_X1   g10673(.A1(new_n11628_), .A2(new_n11675_), .A3(new_n11624_), .A4(new_n11671_), .ZN(new_n11676_));
  AOI22_X1   g10674(.A1(new_n11628_), .A2(new_n11624_), .B1(new_n11675_), .B2(new_n11671_), .ZN(new_n11677_));
  OAI21_X1   g10675(.A1(new_n11677_), .A2(new_n11580_), .B(new_n11676_), .ZN(new_n11678_));
  NAND2_X1   g10676(.A1(new_n11627_), .A2(new_n11616_), .ZN(new_n11679_));
  NAND2_X1   g10677(.A1(new_n11679_), .A2(new_n11622_), .ZN(new_n11680_));
  AOI21_X1   g10678(.A1(new_n11603_), .A2(new_n11614_), .B(new_n11608_), .ZN(new_n11681_));
  NOR2_X1    g10679(.A1(new_n11581_), .A2(new_n11237_), .ZN(new_n11682_));
  AOI21_X1   g10680(.A1(new_n11682_), .A2(new_n11596_), .B(new_n11586_), .ZN(new_n11683_));
  INV_X1     g10681(.I(new_n11683_), .ZN(new_n11684_));
  NOR2_X1    g10682(.A1(new_n11684_), .A2(new_n11681_), .ZN(new_n11685_));
  OAI21_X1   g10683(.A1(new_n11612_), .A2(new_n11610_), .B(new_n11613_), .ZN(new_n11686_));
  NOR2_X1    g10684(.A1(new_n11686_), .A2(new_n11683_), .ZN(new_n11687_));
  NOR2_X1    g10685(.A1(new_n11685_), .A2(new_n11687_), .ZN(new_n11688_));
  NAND2_X1   g10686(.A1(new_n11680_), .A2(new_n11688_), .ZN(new_n11689_));
  INV_X1     g10687(.I(new_n11688_), .ZN(new_n11690_));
  NAND3_X1   g10688(.A1(new_n11690_), .A2(new_n11622_), .A3(new_n11679_), .ZN(new_n11691_));
  OAI21_X1   g10689(.A1(new_n11629_), .A2(new_n11673_), .B(new_n11670_), .ZN(new_n11692_));
  OAI21_X1   g10690(.A1(new_n11653_), .A2(new_n11659_), .B(new_n11661_), .ZN(new_n11693_));
  AOI21_X1   g10691(.A1(new_n11646_), .A2(new_n11648_), .B(new_n11638_), .ZN(new_n11694_));
  XOR2_X1    g10692(.A1(new_n11693_), .A2(new_n11694_), .Z(new_n11695_));
  NAND2_X1   g10693(.A1(new_n11692_), .A2(new_n11695_), .ZN(new_n11696_));
  AOI21_X1   g10694(.A1(new_n11672_), .A2(new_n11664_), .B(new_n11674_), .ZN(new_n11697_));
  INV_X1     g10695(.I(new_n11695_), .ZN(new_n11698_));
  NAND2_X1   g10696(.A1(new_n11698_), .A2(new_n11697_), .ZN(new_n11699_));
  NAND4_X1   g10697(.A1(new_n11689_), .A2(new_n11691_), .A3(new_n11696_), .A4(new_n11699_), .ZN(new_n11700_));
  AOI21_X1   g10698(.A1(new_n11622_), .A2(new_n11679_), .B(new_n11690_), .ZN(new_n11701_));
  NOR2_X1    g10699(.A1(new_n11680_), .A2(new_n11688_), .ZN(new_n11702_));
  INV_X1     g10700(.I(new_n11696_), .ZN(new_n11703_));
  NOR2_X1    g10701(.A1(new_n11692_), .A2(new_n11695_), .ZN(new_n11704_));
  OAI22_X1   g10702(.A1(new_n11701_), .A2(new_n11702_), .B1(new_n11703_), .B2(new_n11704_), .ZN(new_n11705_));
  NAND3_X1   g10703(.A1(new_n11705_), .A2(new_n11700_), .A3(new_n11678_), .ZN(new_n11706_));
  AOI21_X1   g10704(.A1(new_n11705_), .A2(new_n11700_), .B(new_n11678_), .ZN(new_n11707_));
  INV_X1     g10705(.I(new_n11707_), .ZN(new_n11708_));
  NAND2_X1   g10706(.A1(new_n11708_), .A2(new_n11706_), .ZN(new_n11709_));
  NOR3_X1    g10707(.A1(new_n11089_), .A2(new_n11116_), .A3(new_n11078_), .ZN(new_n11710_));
  AOI21_X1   g10708(.A1(new_n11115_), .A2(new_n11090_), .B(new_n11110_), .ZN(new_n11711_));
  NOR2_X1    g10709(.A1(new_n11711_), .A2(new_n11710_), .ZN(new_n11712_));
  NOR2_X1    g10710(.A1(new_n11111_), .A2(new_n11080_), .ZN(new_n11713_));
  NOR2_X1    g10711(.A1(new_n11086_), .A2(new_n11713_), .ZN(new_n11714_));
  NOR2_X1    g10712(.A1(new_n11504_), .A2(new_n11506_), .ZN(new_n11715_));
  NOR2_X1    g10713(.A1(new_n11508_), .A2(new_n11715_), .ZN(new_n11716_));
  NAND2_X1   g10714(.A1(new_n11716_), .A2(new_n11714_), .ZN(new_n11717_));
  NOR3_X1    g10715(.A1(new_n11339_), .A2(new_n11341_), .A3(new_n11340_), .ZN(new_n11718_));
  AOI21_X1   g10716(.A1(new_n11336_), .A2(new_n11327_), .B(new_n11239_), .ZN(new_n11719_));
  NOR2_X1    g10717(.A1(new_n11719_), .A2(new_n11718_), .ZN(new_n11720_));
  OAI21_X1   g10718(.A1(new_n11576_), .A2(new_n11575_), .B(new_n11574_), .ZN(new_n11721_));
  NAND3_X1   g10719(.A1(new_n11540_), .A2(new_n11567_), .A3(new_n11572_), .ZN(new_n11722_));
  AOI21_X1   g10720(.A1(new_n11722_), .A2(new_n11721_), .B(new_n11507_), .ZN(new_n11723_));
  OAI21_X1   g10721(.A1(new_n11579_), .A2(new_n11723_), .B(new_n11720_), .ZN(new_n11724_));
  NAND3_X1   g10722(.A1(new_n11722_), .A2(new_n11721_), .A3(new_n11507_), .ZN(new_n11725_));
  NAND3_X1   g10723(.A1(new_n11578_), .A2(new_n11343_), .A3(new_n11725_), .ZN(new_n11726_));
  AOI21_X1   g10724(.A1(new_n11724_), .A2(new_n11726_), .B(new_n11717_), .ZN(new_n11727_));
  NAND3_X1   g10725(.A1(new_n11724_), .A2(new_n11726_), .A3(new_n11717_), .ZN(new_n11728_));
  OAI21_X1   g10726(.A1(new_n11727_), .A2(new_n11712_), .B(new_n11728_), .ZN(new_n11729_));
  NOR3_X1    g10727(.A1(new_n11075_), .A2(new_n11108_), .A3(new_n11091_), .ZN(new_n11730_));
  AOI21_X1   g10728(.A1(new_n11109_), .A2(new_n11074_), .B(new_n11117_), .ZN(new_n11731_));
  NOR3_X1    g10729(.A1(new_n11626_), .A2(new_n11627_), .A3(new_n11625_), .ZN(new_n11732_));
  AOI21_X1   g10730(.A1(new_n11616_), .A2(new_n11622_), .B(new_n11623_), .ZN(new_n11733_));
  NOR3_X1    g10731(.A1(new_n11672_), .A2(new_n11674_), .A3(new_n11673_), .ZN(new_n11734_));
  AOI21_X1   g10732(.A1(new_n11664_), .A2(new_n11670_), .B(new_n11629_), .ZN(new_n11735_));
  NOR4_X1    g10733(.A1(new_n11732_), .A2(new_n11733_), .A3(new_n11734_), .A4(new_n11735_), .ZN(new_n11736_));
  NOR3_X1    g10734(.A1(new_n11677_), .A2(new_n11736_), .A3(new_n11580_), .ZN(new_n11737_));
  OAI21_X1   g10735(.A1(new_n11720_), .A2(new_n11723_), .B(new_n11725_), .ZN(new_n11738_));
  OAI22_X1   g10736(.A1(new_n11732_), .A2(new_n11733_), .B1(new_n11734_), .B2(new_n11735_), .ZN(new_n11739_));
  AOI21_X1   g10737(.A1(new_n11739_), .A2(new_n11676_), .B(new_n11738_), .ZN(new_n11740_));
  NOR4_X1    g10738(.A1(new_n11737_), .A2(new_n11740_), .A3(new_n11730_), .A4(new_n11731_), .ZN(new_n11741_));
  OAI22_X1   g10739(.A1(new_n11737_), .A2(new_n11740_), .B1(new_n11730_), .B2(new_n11731_), .ZN(new_n11742_));
  AOI21_X1   g10740(.A1(new_n11729_), .A2(new_n11742_), .B(new_n11741_), .ZN(new_n11743_));
  NOR2_X1    g10741(.A1(new_n11709_), .A2(new_n11743_), .ZN(new_n11744_));
  INV_X1     g10742(.I(new_n11706_), .ZN(new_n11745_));
  NOR2_X1    g10743(.A1(new_n11745_), .A2(new_n11707_), .ZN(new_n11746_));
  OR2_X2     g10744(.A1(new_n11711_), .A2(new_n11710_), .Z(new_n11747_));
  INV_X1     g10745(.I(new_n11717_), .ZN(new_n11748_));
  AOI21_X1   g10746(.A1(new_n11578_), .A2(new_n11725_), .B(new_n11343_), .ZN(new_n11749_));
  NOR3_X1    g10747(.A1(new_n11579_), .A2(new_n11720_), .A3(new_n11723_), .ZN(new_n11750_));
  OAI21_X1   g10748(.A1(new_n11750_), .A2(new_n11749_), .B(new_n11748_), .ZN(new_n11751_));
  NOR3_X1    g10749(.A1(new_n11748_), .A2(new_n11750_), .A3(new_n11749_), .ZN(new_n11752_));
  AOI21_X1   g10750(.A1(new_n11747_), .A2(new_n11751_), .B(new_n11752_), .ZN(new_n11753_));
  NAND3_X1   g10751(.A1(new_n11109_), .A2(new_n11074_), .A3(new_n11117_), .ZN(new_n11754_));
  OAI21_X1   g10752(.A1(new_n11075_), .A2(new_n11108_), .B(new_n11091_), .ZN(new_n11755_));
  NAND3_X1   g10753(.A1(new_n11739_), .A2(new_n11676_), .A3(new_n11738_), .ZN(new_n11756_));
  OAI21_X1   g10754(.A1(new_n11677_), .A2(new_n11736_), .B(new_n11580_), .ZN(new_n11757_));
  NAND4_X1   g10755(.A1(new_n11757_), .A2(new_n11756_), .A3(new_n11755_), .A4(new_n11754_), .ZN(new_n11758_));
  AOI22_X1   g10756(.A1(new_n11757_), .A2(new_n11756_), .B1(new_n11755_), .B2(new_n11754_), .ZN(new_n11759_));
  OAI21_X1   g10757(.A1(new_n11753_), .A2(new_n11759_), .B(new_n11758_), .ZN(new_n11760_));
  NOR2_X1    g10758(.A1(new_n11746_), .A2(new_n11760_), .ZN(new_n11761_));
  NOR3_X1    g10759(.A1(new_n11744_), .A2(new_n11761_), .A3(new_n11126_), .ZN(new_n11762_));
  NAND2_X1   g10760(.A1(new_n11746_), .A2(new_n11760_), .ZN(new_n11763_));
  NAND2_X1   g10761(.A1(new_n11709_), .A2(new_n11743_), .ZN(new_n11764_));
  AOI21_X1   g10762(.A1(new_n11764_), .A2(new_n11763_), .B(new_n11125_), .ZN(new_n11765_));
  NOR2_X1    g10763(.A1(new_n11762_), .A2(new_n11765_), .ZN(new_n11766_));
  INV_X1     g10764(.I(\A[673] ), .ZN(new_n11767_));
  INV_X1     g10765(.I(\A[674] ), .ZN(new_n11768_));
  NAND2_X1   g10766(.A1(new_n11768_), .A2(\A[675] ), .ZN(new_n11769_));
  INV_X1     g10767(.I(\A[675] ), .ZN(new_n11770_));
  NAND2_X1   g10768(.A1(new_n11770_), .A2(\A[674] ), .ZN(new_n11771_));
  AOI21_X1   g10769(.A1(new_n11769_), .A2(new_n11771_), .B(new_n11767_), .ZN(new_n11772_));
  NOR2_X1    g10770(.A1(\A[674] ), .A2(\A[675] ), .ZN(new_n11773_));
  INV_X1     g10771(.I(new_n11773_), .ZN(new_n11774_));
  NAND2_X1   g10772(.A1(\A[674] ), .A2(\A[675] ), .ZN(new_n11775_));
  AOI21_X1   g10773(.A1(new_n11774_), .A2(new_n11775_), .B(\A[673] ), .ZN(new_n11776_));
  NOR2_X1    g10774(.A1(new_n11776_), .A2(new_n11772_), .ZN(new_n11777_));
  INV_X1     g10775(.I(\A[676] ), .ZN(new_n11778_));
  INV_X1     g10776(.I(\A[677] ), .ZN(new_n11779_));
  NAND2_X1   g10777(.A1(new_n11779_), .A2(\A[678] ), .ZN(new_n11780_));
  INV_X1     g10778(.I(\A[678] ), .ZN(new_n11781_));
  NAND2_X1   g10779(.A1(new_n11781_), .A2(\A[677] ), .ZN(new_n11782_));
  AOI21_X1   g10780(.A1(new_n11780_), .A2(new_n11782_), .B(new_n11778_), .ZN(new_n11783_));
  NOR2_X1    g10781(.A1(\A[677] ), .A2(\A[678] ), .ZN(new_n11784_));
  INV_X1     g10782(.I(new_n11784_), .ZN(new_n11785_));
  NAND2_X1   g10783(.A1(\A[677] ), .A2(\A[678] ), .ZN(new_n11786_));
  AOI21_X1   g10784(.A1(new_n11785_), .A2(new_n11786_), .B(\A[676] ), .ZN(new_n11787_));
  NOR2_X1    g10785(.A1(new_n11787_), .A2(new_n11783_), .ZN(new_n11788_));
  NAND2_X1   g10786(.A1(new_n11777_), .A2(new_n11788_), .ZN(new_n11789_));
  AOI21_X1   g10787(.A1(new_n11778_), .A2(new_n11786_), .B(new_n11784_), .ZN(new_n11790_));
  AOI21_X1   g10788(.A1(new_n11767_), .A2(new_n11775_), .B(new_n11773_), .ZN(new_n11791_));
  XNOR2_X1   g10789(.A1(new_n11790_), .A2(new_n11791_), .ZN(new_n11792_));
  XNOR2_X1   g10790(.A1(new_n11789_), .A2(new_n11792_), .ZN(new_n11793_));
  INV_X1     g10791(.I(new_n11789_), .ZN(new_n11794_));
  NOR2_X1    g10792(.A1(new_n11777_), .A2(new_n11788_), .ZN(new_n11795_));
  NOR2_X1    g10793(.A1(new_n11794_), .A2(new_n11795_), .ZN(new_n11796_));
  INV_X1     g10794(.I(\A[669] ), .ZN(new_n11797_));
  NOR2_X1    g10795(.A1(new_n11797_), .A2(\A[668] ), .ZN(new_n11798_));
  INV_X1     g10796(.I(\A[668] ), .ZN(new_n11799_));
  NOR2_X1    g10797(.A1(new_n11799_), .A2(\A[669] ), .ZN(new_n11800_));
  OAI21_X1   g10798(.A1(new_n11798_), .A2(new_n11800_), .B(\A[667] ), .ZN(new_n11801_));
  INV_X1     g10799(.I(\A[667] ), .ZN(new_n11802_));
  NAND2_X1   g10800(.A1(\A[668] ), .A2(\A[669] ), .ZN(new_n11803_));
  INV_X1     g10801(.I(new_n11803_), .ZN(new_n11804_));
  NOR2_X1    g10802(.A1(\A[668] ), .A2(\A[669] ), .ZN(new_n11805_));
  OAI21_X1   g10803(.A1(new_n11804_), .A2(new_n11805_), .B(new_n11802_), .ZN(new_n11806_));
  INV_X1     g10804(.I(\A[672] ), .ZN(new_n11807_));
  NOR2_X1    g10805(.A1(new_n11807_), .A2(\A[671] ), .ZN(new_n11808_));
  INV_X1     g10806(.I(\A[671] ), .ZN(new_n11809_));
  NOR2_X1    g10807(.A1(new_n11809_), .A2(\A[672] ), .ZN(new_n11810_));
  OAI21_X1   g10808(.A1(new_n11808_), .A2(new_n11810_), .B(\A[670] ), .ZN(new_n11811_));
  INV_X1     g10809(.I(\A[670] ), .ZN(new_n11812_));
  NAND2_X1   g10810(.A1(\A[671] ), .A2(\A[672] ), .ZN(new_n11813_));
  INV_X1     g10811(.I(new_n11813_), .ZN(new_n11814_));
  NOR2_X1    g10812(.A1(\A[671] ), .A2(\A[672] ), .ZN(new_n11815_));
  OAI21_X1   g10813(.A1(new_n11814_), .A2(new_n11815_), .B(new_n11812_), .ZN(new_n11816_));
  NAND4_X1   g10814(.A1(new_n11801_), .A2(new_n11806_), .A3(new_n11811_), .A4(new_n11816_), .ZN(new_n11817_));
  NAND2_X1   g10815(.A1(new_n11801_), .A2(new_n11806_), .ZN(new_n11818_));
  NAND2_X1   g10816(.A1(new_n11811_), .A2(new_n11816_), .ZN(new_n11819_));
  NAND2_X1   g10817(.A1(new_n11818_), .A2(new_n11819_), .ZN(new_n11820_));
  NAND2_X1   g10818(.A1(new_n11820_), .A2(new_n11817_), .ZN(new_n11821_));
  INV_X1     g10819(.I(new_n11821_), .ZN(new_n11822_));
  NAND2_X1   g10820(.A1(new_n11796_), .A2(new_n11822_), .ZN(new_n11823_));
  NOR2_X1    g10821(.A1(new_n11823_), .A2(new_n11793_), .ZN(new_n11824_));
  AOI21_X1   g10822(.A1(new_n11812_), .A2(new_n11813_), .B(new_n11815_), .ZN(new_n11825_));
  AOI21_X1   g10823(.A1(new_n11802_), .A2(new_n11803_), .B(new_n11805_), .ZN(new_n11826_));
  NOR2_X1    g10824(.A1(new_n11825_), .A2(new_n11826_), .ZN(new_n11827_));
  INV_X1     g10825(.I(new_n11827_), .ZN(new_n11828_));
  NAND2_X1   g10826(.A1(new_n11825_), .A2(new_n11826_), .ZN(new_n11829_));
  NAND2_X1   g10827(.A1(new_n11828_), .A2(new_n11829_), .ZN(new_n11830_));
  XNOR2_X1   g10828(.A1(new_n11830_), .A2(new_n11817_), .ZN(new_n11831_));
  AOI21_X1   g10829(.A1(new_n11823_), .A2(new_n11793_), .B(new_n11831_), .ZN(new_n11832_));
  NAND2_X1   g10830(.A1(new_n11790_), .A2(new_n11791_), .ZN(new_n11833_));
  NOR2_X1    g10831(.A1(new_n11790_), .A2(new_n11791_), .ZN(new_n11834_));
  AOI21_X1   g10832(.A1(new_n11789_), .A2(new_n11833_), .B(new_n11834_), .ZN(new_n11835_));
  AOI21_X1   g10833(.A1(new_n11817_), .A2(new_n11829_), .B(new_n11827_), .ZN(new_n11836_));
  NOR2_X1    g10834(.A1(new_n11835_), .A2(new_n11836_), .ZN(new_n11837_));
  NAND2_X1   g10835(.A1(new_n11835_), .A2(new_n11836_), .ZN(new_n11838_));
  INV_X1     g10836(.I(new_n11838_), .ZN(new_n11839_));
  NOR2_X1    g10837(.A1(new_n11839_), .A2(new_n11837_), .ZN(new_n11840_));
  OAI21_X1   g10838(.A1(new_n11832_), .A2(new_n11824_), .B(new_n11840_), .ZN(new_n11841_));
  XOR2_X1    g10839(.A1(new_n11789_), .A2(new_n11792_), .Z(new_n11842_));
  INV_X1     g10840(.I(new_n11795_), .ZN(new_n11843_));
  NAND2_X1   g10841(.A1(new_n11843_), .A2(new_n11789_), .ZN(new_n11844_));
  NOR2_X1    g10842(.A1(new_n11844_), .A2(new_n11821_), .ZN(new_n11845_));
  NAND2_X1   g10843(.A1(new_n11845_), .A2(new_n11842_), .ZN(new_n11846_));
  XOR2_X1    g10844(.A1(new_n11830_), .A2(new_n11817_), .Z(new_n11847_));
  OAI21_X1   g10845(.A1(new_n11845_), .A2(new_n11842_), .B(new_n11847_), .ZN(new_n11848_));
  INV_X1     g10846(.I(new_n11837_), .ZN(new_n11849_));
  NAND2_X1   g10847(.A1(new_n11849_), .A2(new_n11838_), .ZN(new_n11850_));
  NAND3_X1   g10848(.A1(new_n11848_), .A2(new_n11850_), .A3(new_n11846_), .ZN(new_n11851_));
  NAND2_X1   g10849(.A1(new_n11841_), .A2(new_n11851_), .ZN(new_n11852_));
  INV_X1     g10850(.I(\A[663] ), .ZN(new_n11853_));
  NOR2_X1    g10851(.A1(new_n11853_), .A2(\A[662] ), .ZN(new_n11854_));
  INV_X1     g10852(.I(\A[662] ), .ZN(new_n11855_));
  NOR2_X1    g10853(.A1(new_n11855_), .A2(\A[663] ), .ZN(new_n11856_));
  OAI21_X1   g10854(.A1(new_n11854_), .A2(new_n11856_), .B(\A[661] ), .ZN(new_n11857_));
  INV_X1     g10855(.I(\A[661] ), .ZN(new_n11858_));
  NOR2_X1    g10856(.A1(\A[662] ), .A2(\A[663] ), .ZN(new_n11859_));
  NAND2_X1   g10857(.A1(\A[662] ), .A2(\A[663] ), .ZN(new_n11860_));
  INV_X1     g10858(.I(new_n11860_), .ZN(new_n11861_));
  OAI21_X1   g10859(.A1(new_n11861_), .A2(new_n11859_), .B(new_n11858_), .ZN(new_n11862_));
  NAND2_X1   g10860(.A1(new_n11857_), .A2(new_n11862_), .ZN(new_n11863_));
  INV_X1     g10861(.I(\A[666] ), .ZN(new_n11864_));
  NOR2_X1    g10862(.A1(new_n11864_), .A2(\A[665] ), .ZN(new_n11865_));
  INV_X1     g10863(.I(\A[665] ), .ZN(new_n11866_));
  NOR2_X1    g10864(.A1(new_n11866_), .A2(\A[666] ), .ZN(new_n11867_));
  OAI21_X1   g10865(.A1(new_n11865_), .A2(new_n11867_), .B(\A[664] ), .ZN(new_n11868_));
  INV_X1     g10866(.I(\A[664] ), .ZN(new_n11869_));
  NOR2_X1    g10867(.A1(\A[665] ), .A2(\A[666] ), .ZN(new_n11870_));
  NAND2_X1   g10868(.A1(\A[665] ), .A2(\A[666] ), .ZN(new_n11871_));
  INV_X1     g10869(.I(new_n11871_), .ZN(new_n11872_));
  OAI21_X1   g10870(.A1(new_n11872_), .A2(new_n11870_), .B(new_n11869_), .ZN(new_n11873_));
  NAND2_X1   g10871(.A1(new_n11868_), .A2(new_n11873_), .ZN(new_n11874_));
  NOR2_X1    g10872(.A1(new_n11863_), .A2(new_n11874_), .ZN(new_n11875_));
  AOI21_X1   g10873(.A1(new_n11869_), .A2(new_n11871_), .B(new_n11870_), .ZN(new_n11876_));
  AOI21_X1   g10874(.A1(new_n11858_), .A2(new_n11860_), .B(new_n11859_), .ZN(new_n11877_));
  AOI21_X1   g10875(.A1(new_n11876_), .A2(new_n11877_), .B(new_n11875_), .ZN(new_n11878_));
  NOR2_X1    g10876(.A1(new_n11876_), .A2(new_n11877_), .ZN(new_n11879_));
  NOR2_X1    g10877(.A1(new_n11878_), .A2(new_n11879_), .ZN(new_n11880_));
  INV_X1     g10878(.I(new_n11880_), .ZN(new_n11881_));
  INV_X1     g10879(.I(\A[655] ), .ZN(new_n11882_));
  INV_X1     g10880(.I(\A[656] ), .ZN(new_n11883_));
  NAND2_X1   g10881(.A1(new_n11883_), .A2(\A[657] ), .ZN(new_n11884_));
  INV_X1     g10882(.I(\A[657] ), .ZN(new_n11885_));
  NAND2_X1   g10883(.A1(new_n11885_), .A2(\A[656] ), .ZN(new_n11886_));
  AOI21_X1   g10884(.A1(new_n11884_), .A2(new_n11886_), .B(new_n11882_), .ZN(new_n11887_));
  NAND2_X1   g10885(.A1(\A[656] ), .A2(\A[657] ), .ZN(new_n11888_));
  NOR2_X1    g10886(.A1(\A[656] ), .A2(\A[657] ), .ZN(new_n11889_));
  INV_X1     g10887(.I(new_n11889_), .ZN(new_n11890_));
  AOI21_X1   g10888(.A1(new_n11890_), .A2(new_n11888_), .B(\A[655] ), .ZN(new_n11891_));
  INV_X1     g10889(.I(\A[658] ), .ZN(new_n11892_));
  INV_X1     g10890(.I(\A[659] ), .ZN(new_n11893_));
  NAND2_X1   g10891(.A1(new_n11893_), .A2(\A[660] ), .ZN(new_n11894_));
  INV_X1     g10892(.I(\A[660] ), .ZN(new_n11895_));
  NAND2_X1   g10893(.A1(new_n11895_), .A2(\A[659] ), .ZN(new_n11896_));
  AOI21_X1   g10894(.A1(new_n11894_), .A2(new_n11896_), .B(new_n11892_), .ZN(new_n11897_));
  NAND2_X1   g10895(.A1(\A[659] ), .A2(\A[660] ), .ZN(new_n11898_));
  NOR2_X1    g10896(.A1(\A[659] ), .A2(\A[660] ), .ZN(new_n11899_));
  INV_X1     g10897(.I(new_n11899_), .ZN(new_n11900_));
  AOI21_X1   g10898(.A1(new_n11900_), .A2(new_n11898_), .B(\A[658] ), .ZN(new_n11901_));
  NOR4_X1    g10899(.A1(new_n11887_), .A2(new_n11891_), .A3(new_n11901_), .A4(new_n11897_), .ZN(new_n11902_));
  AOI21_X1   g10900(.A1(new_n11892_), .A2(new_n11898_), .B(new_n11899_), .ZN(new_n11903_));
  AOI21_X1   g10901(.A1(new_n11882_), .A2(new_n11888_), .B(new_n11889_), .ZN(new_n11904_));
  NOR2_X1    g10902(.A1(new_n11903_), .A2(new_n11904_), .ZN(new_n11905_));
  NAND2_X1   g10903(.A1(new_n11903_), .A2(new_n11904_), .ZN(new_n11906_));
  INV_X1     g10904(.I(new_n11906_), .ZN(new_n11907_));
  NOR2_X1    g10905(.A1(new_n11907_), .A2(new_n11905_), .ZN(new_n11908_));
  XNOR2_X1   g10906(.A1(new_n11908_), .A2(new_n11902_), .ZN(new_n11909_));
  XOR2_X1    g10907(.A1(new_n11876_), .A2(new_n11877_), .Z(new_n11910_));
  NOR2_X1    g10908(.A1(new_n11875_), .A2(new_n11910_), .ZN(new_n11911_));
  NAND2_X1   g10909(.A1(new_n11855_), .A2(\A[663] ), .ZN(new_n11912_));
  NAND2_X1   g10910(.A1(new_n11853_), .A2(\A[662] ), .ZN(new_n11913_));
  AOI21_X1   g10911(.A1(new_n11912_), .A2(new_n11913_), .B(new_n11858_), .ZN(new_n11914_));
  INV_X1     g10912(.I(new_n11859_), .ZN(new_n11915_));
  AOI21_X1   g10913(.A1(new_n11915_), .A2(new_n11860_), .B(\A[661] ), .ZN(new_n11916_));
  NOR2_X1    g10914(.A1(new_n11916_), .A2(new_n11914_), .ZN(new_n11917_));
  NAND2_X1   g10915(.A1(new_n11866_), .A2(\A[666] ), .ZN(new_n11918_));
  NAND2_X1   g10916(.A1(new_n11864_), .A2(\A[665] ), .ZN(new_n11919_));
  AOI21_X1   g10917(.A1(new_n11918_), .A2(new_n11919_), .B(new_n11869_), .ZN(new_n11920_));
  INV_X1     g10918(.I(new_n11870_), .ZN(new_n11921_));
  AOI21_X1   g10919(.A1(new_n11921_), .A2(new_n11871_), .B(\A[664] ), .ZN(new_n11922_));
  NOR2_X1    g10920(.A1(new_n11922_), .A2(new_n11920_), .ZN(new_n11923_));
  NAND2_X1   g10921(.A1(new_n11917_), .A2(new_n11923_), .ZN(new_n11924_));
  XNOR2_X1   g10922(.A1(new_n11876_), .A2(new_n11877_), .ZN(new_n11925_));
  NOR2_X1    g10923(.A1(new_n11924_), .A2(new_n11925_), .ZN(new_n11926_));
  NOR2_X1    g10924(.A1(new_n11926_), .A2(new_n11911_), .ZN(new_n11927_));
  INV_X1     g10925(.I(new_n11927_), .ZN(new_n11928_));
  NOR2_X1    g10926(.A1(new_n11917_), .A2(new_n11923_), .ZN(new_n11929_));
  NOR2_X1    g10927(.A1(new_n11929_), .A2(new_n11875_), .ZN(new_n11930_));
  NOR2_X1    g10928(.A1(new_n11891_), .A2(new_n11887_), .ZN(new_n11931_));
  NOR2_X1    g10929(.A1(new_n11901_), .A2(new_n11897_), .ZN(new_n11932_));
  NOR2_X1    g10930(.A1(new_n11931_), .A2(new_n11932_), .ZN(new_n11933_));
  NOR2_X1    g10931(.A1(new_n11933_), .A2(new_n11902_), .ZN(new_n11934_));
  NAND2_X1   g10932(.A1(new_n11930_), .A2(new_n11934_), .ZN(new_n11935_));
  AOI21_X1   g10933(.A1(new_n11928_), .A2(new_n11935_), .B(new_n11909_), .ZN(new_n11936_));
  NOR2_X1    g10934(.A1(new_n11928_), .A2(new_n11935_), .ZN(new_n11937_));
  INV_X1     g10935(.I(new_n11905_), .ZN(new_n11938_));
  OAI21_X1   g10936(.A1(new_n11902_), .A2(new_n11907_), .B(new_n11938_), .ZN(new_n11939_));
  INV_X1     g10937(.I(new_n11939_), .ZN(new_n11940_));
  NOR3_X1    g10938(.A1(new_n11936_), .A2(new_n11937_), .A3(new_n11940_), .ZN(new_n11941_));
  XOR2_X1    g10939(.A1(new_n11908_), .A2(new_n11902_), .Z(new_n11942_));
  NAND2_X1   g10940(.A1(new_n11863_), .A2(new_n11874_), .ZN(new_n11943_));
  NAND2_X1   g10941(.A1(new_n11924_), .A2(new_n11943_), .ZN(new_n11944_));
  OR2_X2     g10942(.A1(new_n11933_), .A2(new_n11902_), .Z(new_n11945_));
  OAI22_X1   g10943(.A1(new_n11945_), .A2(new_n11944_), .B1(new_n11911_), .B2(new_n11926_), .ZN(new_n11946_));
  NAND2_X1   g10944(.A1(new_n11946_), .A2(new_n11942_), .ZN(new_n11947_));
  NAND3_X1   g10945(.A1(new_n11927_), .A2(new_n11930_), .A3(new_n11934_), .ZN(new_n11948_));
  AOI21_X1   g10946(.A1(new_n11947_), .A2(new_n11948_), .B(new_n11939_), .ZN(new_n11949_));
  NOR3_X1    g10947(.A1(new_n11941_), .A2(new_n11949_), .A3(new_n11881_), .ZN(new_n11950_));
  NAND3_X1   g10948(.A1(new_n11947_), .A2(new_n11948_), .A3(new_n11939_), .ZN(new_n11951_));
  OAI21_X1   g10949(.A1(new_n11936_), .A2(new_n11937_), .B(new_n11940_), .ZN(new_n11952_));
  AOI21_X1   g10950(.A1(new_n11952_), .A2(new_n11951_), .B(new_n11880_), .ZN(new_n11953_));
  OAI21_X1   g10951(.A1(new_n11950_), .A2(new_n11953_), .B(new_n11852_), .ZN(new_n11954_));
  AOI21_X1   g10952(.A1(new_n11848_), .A2(new_n11846_), .B(new_n11850_), .ZN(new_n11955_));
  NOR3_X1    g10953(.A1(new_n11832_), .A2(new_n11824_), .A3(new_n11840_), .ZN(new_n11956_));
  NOR2_X1    g10954(.A1(new_n11956_), .A2(new_n11955_), .ZN(new_n11957_));
  NAND3_X1   g10955(.A1(new_n11952_), .A2(new_n11951_), .A3(new_n11880_), .ZN(new_n11958_));
  OAI21_X1   g10956(.A1(new_n11941_), .A2(new_n11949_), .B(new_n11881_), .ZN(new_n11959_));
  NAND3_X1   g10957(.A1(new_n11957_), .A2(new_n11959_), .A3(new_n11958_), .ZN(new_n11960_));
  NAND2_X1   g10958(.A1(new_n11823_), .A2(new_n11793_), .ZN(new_n11961_));
  NAND3_X1   g10959(.A1(new_n11961_), .A2(new_n11846_), .A3(new_n11831_), .ZN(new_n11962_));
  NOR2_X1    g10960(.A1(new_n11845_), .A2(new_n11842_), .ZN(new_n11963_));
  OAI21_X1   g10961(.A1(new_n11824_), .A2(new_n11963_), .B(new_n11847_), .ZN(new_n11964_));
  NAND2_X1   g10962(.A1(new_n11964_), .A2(new_n11962_), .ZN(new_n11965_));
  NOR2_X1    g10963(.A1(new_n11947_), .A2(new_n11937_), .ZN(new_n11966_));
  AOI21_X1   g10964(.A1(new_n11948_), .A2(new_n11946_), .B(new_n11942_), .ZN(new_n11967_));
  NAND2_X1   g10965(.A1(new_n11796_), .A2(new_n11821_), .ZN(new_n11968_));
  NAND2_X1   g10966(.A1(new_n11844_), .A2(new_n11822_), .ZN(new_n11969_));
  NAND2_X1   g10967(.A1(new_n11969_), .A2(new_n11968_), .ZN(new_n11970_));
  NAND2_X1   g10968(.A1(new_n11945_), .A2(new_n11930_), .ZN(new_n11971_));
  NAND2_X1   g10969(.A1(new_n11944_), .A2(new_n11934_), .ZN(new_n11972_));
  NAND2_X1   g10970(.A1(new_n11971_), .A2(new_n11972_), .ZN(new_n11973_));
  NAND2_X1   g10971(.A1(new_n11970_), .A2(new_n11973_), .ZN(new_n11974_));
  NOR3_X1    g10972(.A1(new_n11966_), .A2(new_n11967_), .A3(new_n11974_), .ZN(new_n11975_));
  OAI21_X1   g10973(.A1(new_n11966_), .A2(new_n11967_), .B(new_n11974_), .ZN(new_n11976_));
  OAI21_X1   g10974(.A1(new_n11965_), .A2(new_n11975_), .B(new_n11976_), .ZN(new_n11977_));
  NAND3_X1   g10975(.A1(new_n11960_), .A2(new_n11954_), .A3(new_n11977_), .ZN(new_n11978_));
  AOI21_X1   g10976(.A1(new_n11958_), .A2(new_n11959_), .B(new_n11957_), .ZN(new_n11979_));
  NOR3_X1    g10977(.A1(new_n11950_), .A2(new_n11953_), .A3(new_n11852_), .ZN(new_n11980_));
  NOR3_X1    g10978(.A1(new_n11824_), .A2(new_n11963_), .A3(new_n11847_), .ZN(new_n11981_));
  AOI21_X1   g10979(.A1(new_n11961_), .A2(new_n11846_), .B(new_n11831_), .ZN(new_n11982_));
  NOR2_X1    g10980(.A1(new_n11982_), .A2(new_n11981_), .ZN(new_n11983_));
  NAND3_X1   g10981(.A1(new_n11948_), .A2(new_n11946_), .A3(new_n11942_), .ZN(new_n11984_));
  INV_X1     g10982(.I(new_n11967_), .ZN(new_n11985_));
  AOI22_X1   g10983(.A1(new_n11969_), .A2(new_n11968_), .B1(new_n11971_), .B2(new_n11972_), .ZN(new_n11986_));
  NAND3_X1   g10984(.A1(new_n11985_), .A2(new_n11984_), .A3(new_n11986_), .ZN(new_n11987_));
  AOI21_X1   g10985(.A1(new_n11985_), .A2(new_n11984_), .B(new_n11986_), .ZN(new_n11988_));
  AOI21_X1   g10986(.A1(new_n11983_), .A2(new_n11987_), .B(new_n11988_), .ZN(new_n11989_));
  OAI21_X1   g10987(.A1(new_n11979_), .A2(new_n11980_), .B(new_n11989_), .ZN(new_n11990_));
  INV_X1     g10988(.I(\A[679] ), .ZN(new_n11991_));
  INV_X1     g10989(.I(\A[680] ), .ZN(new_n11992_));
  NAND2_X1   g10990(.A1(new_n11992_), .A2(\A[681] ), .ZN(new_n11993_));
  INV_X1     g10991(.I(\A[681] ), .ZN(new_n11994_));
  NAND2_X1   g10992(.A1(new_n11994_), .A2(\A[680] ), .ZN(new_n11995_));
  AOI21_X1   g10993(.A1(new_n11993_), .A2(new_n11995_), .B(new_n11991_), .ZN(new_n11996_));
  NAND2_X1   g10994(.A1(\A[680] ), .A2(\A[681] ), .ZN(new_n11997_));
  NOR2_X1    g10995(.A1(\A[680] ), .A2(\A[681] ), .ZN(new_n11998_));
  INV_X1     g10996(.I(new_n11998_), .ZN(new_n11999_));
  AOI21_X1   g10997(.A1(new_n11999_), .A2(new_n11997_), .B(\A[679] ), .ZN(new_n12000_));
  INV_X1     g10998(.I(\A[682] ), .ZN(new_n12001_));
  INV_X1     g10999(.I(\A[683] ), .ZN(new_n12002_));
  NAND2_X1   g11000(.A1(new_n12002_), .A2(\A[684] ), .ZN(new_n12003_));
  INV_X1     g11001(.I(\A[684] ), .ZN(new_n12004_));
  NAND2_X1   g11002(.A1(new_n12004_), .A2(\A[683] ), .ZN(new_n12005_));
  AOI21_X1   g11003(.A1(new_n12003_), .A2(new_n12005_), .B(new_n12001_), .ZN(new_n12006_));
  NAND2_X1   g11004(.A1(\A[683] ), .A2(\A[684] ), .ZN(new_n12007_));
  NOR2_X1    g11005(.A1(\A[683] ), .A2(\A[684] ), .ZN(new_n12008_));
  INV_X1     g11006(.I(new_n12008_), .ZN(new_n12009_));
  AOI21_X1   g11007(.A1(new_n12009_), .A2(new_n12007_), .B(\A[682] ), .ZN(new_n12010_));
  NOR4_X1    g11008(.A1(new_n11996_), .A2(new_n12000_), .A3(new_n12010_), .A4(new_n12006_), .ZN(new_n12011_));
  AOI21_X1   g11009(.A1(new_n12001_), .A2(new_n12007_), .B(new_n12008_), .ZN(new_n12012_));
  AOI21_X1   g11010(.A1(\A[680] ), .A2(\A[681] ), .B(\A[679] ), .ZN(new_n12013_));
  NOR2_X1    g11011(.A1(new_n12013_), .A2(new_n11998_), .ZN(new_n12014_));
  NOR2_X1    g11012(.A1(new_n12012_), .A2(new_n12014_), .ZN(new_n12015_));
  NAND2_X1   g11013(.A1(new_n12012_), .A2(new_n12014_), .ZN(new_n12016_));
  INV_X1     g11014(.I(new_n12016_), .ZN(new_n12017_));
  NOR2_X1    g11015(.A1(new_n12017_), .A2(new_n12015_), .ZN(new_n12018_));
  XNOR2_X1   g11016(.A1(new_n12018_), .A2(new_n12011_), .ZN(new_n12019_));
  INV_X1     g11017(.I(\A[687] ), .ZN(new_n12020_));
  NOR2_X1    g11018(.A1(new_n12020_), .A2(\A[686] ), .ZN(new_n12021_));
  INV_X1     g11019(.I(\A[686] ), .ZN(new_n12022_));
  NOR2_X1    g11020(.A1(new_n12022_), .A2(\A[687] ), .ZN(new_n12023_));
  OAI21_X1   g11021(.A1(new_n12021_), .A2(new_n12023_), .B(\A[685] ), .ZN(new_n12024_));
  INV_X1     g11022(.I(\A[685] ), .ZN(new_n12025_));
  NOR2_X1    g11023(.A1(\A[686] ), .A2(\A[687] ), .ZN(new_n12026_));
  NOR2_X1    g11024(.A1(new_n12022_), .A2(new_n12020_), .ZN(new_n12027_));
  OAI21_X1   g11025(.A1(new_n12027_), .A2(new_n12026_), .B(new_n12025_), .ZN(new_n12028_));
  INV_X1     g11026(.I(\A[690] ), .ZN(new_n12029_));
  NOR2_X1    g11027(.A1(new_n12029_), .A2(\A[689] ), .ZN(new_n12030_));
  INV_X1     g11028(.I(\A[689] ), .ZN(new_n12031_));
  NOR2_X1    g11029(.A1(new_n12031_), .A2(\A[690] ), .ZN(new_n12032_));
  OAI21_X1   g11030(.A1(new_n12030_), .A2(new_n12032_), .B(\A[688] ), .ZN(new_n12033_));
  INV_X1     g11031(.I(\A[688] ), .ZN(new_n12034_));
  NOR2_X1    g11032(.A1(\A[689] ), .A2(\A[690] ), .ZN(new_n12035_));
  NOR2_X1    g11033(.A1(new_n12031_), .A2(new_n12029_), .ZN(new_n12036_));
  OAI21_X1   g11034(.A1(new_n12036_), .A2(new_n12035_), .B(new_n12034_), .ZN(new_n12037_));
  NAND4_X1   g11035(.A1(new_n12024_), .A2(new_n12028_), .A3(new_n12037_), .A4(new_n12033_), .ZN(new_n12038_));
  AOI21_X1   g11036(.A1(\A[689] ), .A2(\A[690] ), .B(\A[688] ), .ZN(new_n12039_));
  NOR2_X1    g11037(.A1(new_n12039_), .A2(new_n12035_), .ZN(new_n12040_));
  AOI21_X1   g11038(.A1(\A[686] ), .A2(\A[687] ), .B(\A[685] ), .ZN(new_n12041_));
  NOR2_X1    g11039(.A1(new_n12041_), .A2(new_n12026_), .ZN(new_n12042_));
  XNOR2_X1   g11040(.A1(new_n12040_), .A2(new_n12042_), .ZN(new_n12043_));
  XNOR2_X1   g11041(.A1(new_n12043_), .A2(new_n12038_), .ZN(new_n12044_));
  NAND2_X1   g11042(.A1(new_n12028_), .A2(new_n12024_), .ZN(new_n12045_));
  NAND2_X1   g11043(.A1(new_n12037_), .A2(new_n12033_), .ZN(new_n12046_));
  NAND2_X1   g11044(.A1(new_n12045_), .A2(new_n12046_), .ZN(new_n12047_));
  NAND2_X1   g11045(.A1(new_n12047_), .A2(new_n12038_), .ZN(new_n12048_));
  INV_X1     g11046(.I(new_n12048_), .ZN(new_n12049_));
  OAI22_X1   g11047(.A1(new_n11996_), .A2(new_n12000_), .B1(new_n12010_), .B2(new_n12006_), .ZN(new_n12050_));
  INV_X1     g11048(.I(new_n12050_), .ZN(new_n12051_));
  NOR2_X1    g11049(.A1(new_n12051_), .A2(new_n12011_), .ZN(new_n12052_));
  NAND2_X1   g11050(.A1(new_n12049_), .A2(new_n12052_), .ZN(new_n12053_));
  AOI21_X1   g11051(.A1(new_n12053_), .A2(new_n12044_), .B(new_n12019_), .ZN(new_n12054_));
  XOR2_X1    g11052(.A1(new_n12043_), .A2(new_n12038_), .Z(new_n12055_));
  INV_X1     g11053(.I(new_n12011_), .ZN(new_n12056_));
  NAND2_X1   g11054(.A1(new_n12056_), .A2(new_n12050_), .ZN(new_n12057_));
  NOR2_X1    g11055(.A1(new_n12057_), .A2(new_n12048_), .ZN(new_n12058_));
  NAND2_X1   g11056(.A1(new_n12055_), .A2(new_n12058_), .ZN(new_n12059_));
  NAND2_X1   g11057(.A1(new_n12053_), .A2(new_n12044_), .ZN(new_n12060_));
  NAND2_X1   g11058(.A1(new_n12060_), .A2(new_n12059_), .ZN(new_n12061_));
  AOI22_X1   g11059(.A1(new_n12061_), .A2(new_n12019_), .B1(new_n12054_), .B2(new_n12059_), .ZN(new_n12062_));
  INV_X1     g11060(.I(\A[699] ), .ZN(new_n12063_));
  NOR2_X1    g11061(.A1(new_n12063_), .A2(\A[698] ), .ZN(new_n12064_));
  INV_X1     g11062(.I(\A[698] ), .ZN(new_n12065_));
  NOR2_X1    g11063(.A1(new_n12065_), .A2(\A[699] ), .ZN(new_n12066_));
  OAI21_X1   g11064(.A1(new_n12064_), .A2(new_n12066_), .B(\A[697] ), .ZN(new_n12067_));
  INV_X1     g11065(.I(\A[697] ), .ZN(new_n12068_));
  NOR2_X1    g11066(.A1(\A[698] ), .A2(\A[699] ), .ZN(new_n12069_));
  NAND2_X1   g11067(.A1(\A[698] ), .A2(\A[699] ), .ZN(new_n12070_));
  INV_X1     g11068(.I(new_n12070_), .ZN(new_n12071_));
  OAI21_X1   g11069(.A1(new_n12071_), .A2(new_n12069_), .B(new_n12068_), .ZN(new_n12072_));
  NAND2_X1   g11070(.A1(new_n12067_), .A2(new_n12072_), .ZN(new_n12073_));
  INV_X1     g11071(.I(\A[702] ), .ZN(new_n12074_));
  NOR2_X1    g11072(.A1(new_n12074_), .A2(\A[701] ), .ZN(new_n12075_));
  INV_X1     g11073(.I(\A[701] ), .ZN(new_n12076_));
  NOR2_X1    g11074(.A1(new_n12076_), .A2(\A[702] ), .ZN(new_n12077_));
  OAI21_X1   g11075(.A1(new_n12075_), .A2(new_n12077_), .B(\A[700] ), .ZN(new_n12078_));
  INV_X1     g11076(.I(\A[700] ), .ZN(new_n12079_));
  NOR2_X1    g11077(.A1(\A[701] ), .A2(\A[702] ), .ZN(new_n12080_));
  NAND2_X1   g11078(.A1(\A[701] ), .A2(\A[702] ), .ZN(new_n12081_));
  INV_X1     g11079(.I(new_n12081_), .ZN(new_n12082_));
  OAI21_X1   g11080(.A1(new_n12082_), .A2(new_n12080_), .B(new_n12079_), .ZN(new_n12083_));
  NAND2_X1   g11081(.A1(new_n12078_), .A2(new_n12083_), .ZN(new_n12084_));
  NOR2_X1    g11082(.A1(new_n12073_), .A2(new_n12084_), .ZN(new_n12085_));
  NAND2_X1   g11083(.A1(new_n12065_), .A2(\A[699] ), .ZN(new_n12086_));
  NAND2_X1   g11084(.A1(new_n12063_), .A2(\A[698] ), .ZN(new_n12087_));
  AOI21_X1   g11085(.A1(new_n12086_), .A2(new_n12087_), .B(new_n12068_), .ZN(new_n12088_));
  INV_X1     g11086(.I(new_n12069_), .ZN(new_n12089_));
  AOI21_X1   g11087(.A1(new_n12089_), .A2(new_n12070_), .B(\A[697] ), .ZN(new_n12090_));
  NOR2_X1    g11088(.A1(new_n12090_), .A2(new_n12088_), .ZN(new_n12091_));
  NAND2_X1   g11089(.A1(new_n12076_), .A2(\A[702] ), .ZN(new_n12092_));
  NAND2_X1   g11090(.A1(new_n12074_), .A2(\A[701] ), .ZN(new_n12093_));
  AOI21_X1   g11091(.A1(new_n12092_), .A2(new_n12093_), .B(new_n12079_), .ZN(new_n12094_));
  INV_X1     g11092(.I(new_n12080_), .ZN(new_n12095_));
  AOI21_X1   g11093(.A1(new_n12095_), .A2(new_n12081_), .B(\A[700] ), .ZN(new_n12096_));
  NOR2_X1    g11094(.A1(new_n12096_), .A2(new_n12094_), .ZN(new_n12097_));
  NOR2_X1    g11095(.A1(new_n12091_), .A2(new_n12097_), .ZN(new_n12098_));
  NOR2_X1    g11096(.A1(new_n12098_), .A2(new_n12085_), .ZN(new_n12099_));
  INV_X1     g11097(.I(\A[691] ), .ZN(new_n12100_));
  INV_X1     g11098(.I(\A[692] ), .ZN(new_n12101_));
  NAND2_X1   g11099(.A1(new_n12101_), .A2(\A[693] ), .ZN(new_n12102_));
  INV_X1     g11100(.I(\A[693] ), .ZN(new_n12103_));
  NAND2_X1   g11101(.A1(new_n12103_), .A2(\A[692] ), .ZN(new_n12104_));
  AOI21_X1   g11102(.A1(new_n12102_), .A2(new_n12104_), .B(new_n12100_), .ZN(new_n12105_));
  NAND2_X1   g11103(.A1(\A[692] ), .A2(\A[693] ), .ZN(new_n12106_));
  NOR2_X1    g11104(.A1(\A[692] ), .A2(\A[693] ), .ZN(new_n12107_));
  INV_X1     g11105(.I(new_n12107_), .ZN(new_n12108_));
  AOI21_X1   g11106(.A1(new_n12108_), .A2(new_n12106_), .B(\A[691] ), .ZN(new_n12109_));
  NOR2_X1    g11107(.A1(new_n12109_), .A2(new_n12105_), .ZN(new_n12110_));
  INV_X1     g11108(.I(\A[694] ), .ZN(new_n12111_));
  INV_X1     g11109(.I(\A[695] ), .ZN(new_n12112_));
  NAND2_X1   g11110(.A1(new_n12112_), .A2(\A[696] ), .ZN(new_n12113_));
  INV_X1     g11111(.I(\A[696] ), .ZN(new_n12114_));
  NAND2_X1   g11112(.A1(new_n12114_), .A2(\A[695] ), .ZN(new_n12115_));
  AOI21_X1   g11113(.A1(new_n12113_), .A2(new_n12115_), .B(new_n12111_), .ZN(new_n12116_));
  NAND2_X1   g11114(.A1(\A[695] ), .A2(\A[696] ), .ZN(new_n12117_));
  NOR2_X1    g11115(.A1(\A[695] ), .A2(\A[696] ), .ZN(new_n12118_));
  INV_X1     g11116(.I(new_n12118_), .ZN(new_n12119_));
  AOI21_X1   g11117(.A1(new_n12119_), .A2(new_n12117_), .B(\A[694] ), .ZN(new_n12120_));
  NOR2_X1    g11118(.A1(new_n12120_), .A2(new_n12116_), .ZN(new_n12121_));
  NAND2_X1   g11119(.A1(new_n12110_), .A2(new_n12121_), .ZN(new_n12122_));
  NOR2_X1    g11120(.A1(new_n12103_), .A2(\A[692] ), .ZN(new_n12123_));
  NOR2_X1    g11121(.A1(new_n12101_), .A2(\A[693] ), .ZN(new_n12124_));
  OAI21_X1   g11122(.A1(new_n12123_), .A2(new_n12124_), .B(\A[691] ), .ZN(new_n12125_));
  INV_X1     g11123(.I(new_n12106_), .ZN(new_n12126_));
  OAI21_X1   g11124(.A1(new_n12126_), .A2(new_n12107_), .B(new_n12100_), .ZN(new_n12127_));
  NAND2_X1   g11125(.A1(new_n12125_), .A2(new_n12127_), .ZN(new_n12128_));
  NOR2_X1    g11126(.A1(new_n12114_), .A2(\A[695] ), .ZN(new_n12129_));
  NOR2_X1    g11127(.A1(new_n12112_), .A2(\A[696] ), .ZN(new_n12130_));
  OAI21_X1   g11128(.A1(new_n12129_), .A2(new_n12130_), .B(\A[694] ), .ZN(new_n12131_));
  INV_X1     g11129(.I(new_n12117_), .ZN(new_n12132_));
  OAI21_X1   g11130(.A1(new_n12132_), .A2(new_n12118_), .B(new_n12111_), .ZN(new_n12133_));
  NAND2_X1   g11131(.A1(new_n12131_), .A2(new_n12133_), .ZN(new_n12134_));
  NAND2_X1   g11132(.A1(new_n12128_), .A2(new_n12134_), .ZN(new_n12135_));
  NAND2_X1   g11133(.A1(new_n12122_), .A2(new_n12135_), .ZN(new_n12136_));
  NAND2_X1   g11134(.A1(new_n12099_), .A2(new_n12136_), .ZN(new_n12137_));
  NAND2_X1   g11135(.A1(new_n12091_), .A2(new_n12097_), .ZN(new_n12138_));
  NAND2_X1   g11136(.A1(new_n12073_), .A2(new_n12084_), .ZN(new_n12139_));
  NAND2_X1   g11137(.A1(new_n12138_), .A2(new_n12139_), .ZN(new_n12140_));
  NOR2_X1    g11138(.A1(new_n12128_), .A2(new_n12134_), .ZN(new_n12141_));
  NOR2_X1    g11139(.A1(new_n12110_), .A2(new_n12121_), .ZN(new_n12142_));
  NOR2_X1    g11140(.A1(new_n12142_), .A2(new_n12141_), .ZN(new_n12143_));
  NAND2_X1   g11141(.A1(new_n12143_), .A2(new_n12140_), .ZN(new_n12144_));
  NAND2_X1   g11142(.A1(new_n12049_), .A2(new_n12057_), .ZN(new_n12145_));
  NAND2_X1   g11143(.A1(new_n12052_), .A2(new_n12048_), .ZN(new_n12146_));
  AOI22_X1   g11144(.A1(new_n12145_), .A2(new_n12146_), .B1(new_n12144_), .B2(new_n12137_), .ZN(new_n12147_));
  INV_X1     g11145(.I(new_n12147_), .ZN(new_n12148_));
  AOI21_X1   g11146(.A1(\A[695] ), .A2(\A[696] ), .B(\A[694] ), .ZN(new_n12149_));
  AOI21_X1   g11147(.A1(\A[692] ), .A2(\A[693] ), .B(\A[691] ), .ZN(new_n12150_));
  OAI22_X1   g11148(.A1(new_n12107_), .A2(new_n12150_), .B1(new_n12149_), .B2(new_n12118_), .ZN(new_n12151_));
  NOR4_X1    g11149(.A1(new_n12149_), .A2(new_n12150_), .A3(new_n12107_), .A4(new_n12118_), .ZN(new_n12152_));
  INV_X1     g11150(.I(new_n12152_), .ZN(new_n12153_));
  NAND2_X1   g11151(.A1(new_n12153_), .A2(new_n12151_), .ZN(new_n12154_));
  XOR2_X1    g11152(.A1(new_n12141_), .A2(new_n12154_), .Z(new_n12155_));
  AOI21_X1   g11153(.A1(new_n12079_), .A2(new_n12081_), .B(new_n12080_), .ZN(new_n12156_));
  AOI21_X1   g11154(.A1(new_n12068_), .A2(new_n12070_), .B(new_n12069_), .ZN(new_n12157_));
  XOR2_X1    g11155(.A1(new_n12156_), .A2(new_n12157_), .Z(new_n12158_));
  NOR2_X1    g11156(.A1(new_n12085_), .A2(new_n12158_), .ZN(new_n12159_));
  XNOR2_X1   g11157(.A1(new_n12156_), .A2(new_n12157_), .ZN(new_n12160_));
  NOR2_X1    g11158(.A1(new_n12138_), .A2(new_n12160_), .ZN(new_n12161_));
  OAI22_X1   g11159(.A1(new_n12140_), .A2(new_n12136_), .B1(new_n12161_), .B2(new_n12159_), .ZN(new_n12162_));
  NOR2_X1    g11160(.A1(new_n12161_), .A2(new_n12159_), .ZN(new_n12163_));
  NAND3_X1   g11161(.A1(new_n12163_), .A2(new_n12099_), .A3(new_n12143_), .ZN(new_n12164_));
  NAND3_X1   g11162(.A1(new_n12164_), .A2(new_n12162_), .A3(new_n12155_), .ZN(new_n12165_));
  XOR2_X1    g11163(.A1(new_n12122_), .A2(new_n12154_), .Z(new_n12166_));
  INV_X1     g11164(.I(new_n12162_), .ZN(new_n12167_));
  NAND2_X1   g11165(.A1(new_n12143_), .A2(new_n12099_), .ZN(new_n12168_));
  NOR3_X1    g11166(.A1(new_n12168_), .A2(new_n12159_), .A3(new_n12161_), .ZN(new_n12169_));
  OAI21_X1   g11167(.A1(new_n12167_), .A2(new_n12169_), .B(new_n12166_), .ZN(new_n12170_));
  AOI21_X1   g11168(.A1(new_n12170_), .A2(new_n12165_), .B(new_n12148_), .ZN(new_n12171_));
  NAND3_X1   g11169(.A1(new_n12148_), .A2(new_n12170_), .A3(new_n12165_), .ZN(new_n12172_));
  OAI21_X1   g11170(.A1(new_n12171_), .A2(new_n12062_), .B(new_n12172_), .ZN(new_n12173_));
  INV_X1     g11171(.I(new_n12163_), .ZN(new_n12174_));
  AOI21_X1   g11172(.A1(new_n12174_), .A2(new_n12168_), .B(new_n12155_), .ZN(new_n12175_));
  INV_X1     g11173(.I(new_n12156_), .ZN(new_n12176_));
  INV_X1     g11174(.I(new_n12157_), .ZN(new_n12177_));
  NOR2_X1    g11175(.A1(new_n12176_), .A2(new_n12177_), .ZN(new_n12178_));
  INV_X1     g11176(.I(new_n12178_), .ZN(new_n12179_));
  NOR2_X1    g11177(.A1(new_n12156_), .A2(new_n12157_), .ZN(new_n12180_));
  AOI21_X1   g11178(.A1(new_n12138_), .A2(new_n12179_), .B(new_n12180_), .ZN(new_n12181_));
  INV_X1     g11179(.I(new_n12151_), .ZN(new_n12182_));
  AOI21_X1   g11180(.A1(new_n12122_), .A2(new_n12153_), .B(new_n12182_), .ZN(new_n12183_));
  NOR2_X1    g11181(.A1(new_n12181_), .A2(new_n12183_), .ZN(new_n12184_));
  INV_X1     g11182(.I(new_n12180_), .ZN(new_n12185_));
  OAI21_X1   g11183(.A1(new_n12085_), .A2(new_n12178_), .B(new_n12185_), .ZN(new_n12186_));
  OAI21_X1   g11184(.A1(new_n12141_), .A2(new_n12152_), .B(new_n12151_), .ZN(new_n12187_));
  NOR2_X1    g11185(.A1(new_n12186_), .A2(new_n12187_), .ZN(new_n12188_));
  NOR2_X1    g11186(.A1(new_n12184_), .A2(new_n12188_), .ZN(new_n12189_));
  OAI21_X1   g11187(.A1(new_n12175_), .A2(new_n12169_), .B(new_n12189_), .ZN(new_n12190_));
  NAND2_X1   g11188(.A1(new_n12162_), .A2(new_n12166_), .ZN(new_n12191_));
  NAND2_X1   g11189(.A1(new_n12186_), .A2(new_n12187_), .ZN(new_n12192_));
  NAND2_X1   g11190(.A1(new_n12181_), .A2(new_n12183_), .ZN(new_n12193_));
  NAND2_X1   g11191(.A1(new_n12193_), .A2(new_n12192_), .ZN(new_n12194_));
  NAND3_X1   g11192(.A1(new_n12191_), .A2(new_n12194_), .A3(new_n12164_), .ZN(new_n12195_));
  NAND2_X1   g11193(.A1(new_n12190_), .A2(new_n12195_), .ZN(new_n12196_));
  NOR4_X1    g11194(.A1(new_n12039_), .A2(new_n12041_), .A3(new_n12026_), .A4(new_n12035_), .ZN(new_n12197_));
  INV_X1     g11195(.I(new_n12197_), .ZN(new_n12198_));
  NOR2_X1    g11196(.A1(new_n12040_), .A2(new_n12042_), .ZN(new_n12199_));
  AOI21_X1   g11197(.A1(new_n12038_), .A2(new_n12198_), .B(new_n12199_), .ZN(new_n12200_));
  INV_X1     g11198(.I(new_n12200_), .ZN(new_n12201_));
  NOR2_X1    g11199(.A1(new_n12053_), .A2(new_n12044_), .ZN(new_n12202_));
  INV_X1     g11200(.I(new_n12015_), .ZN(new_n12203_));
  OAI21_X1   g11201(.A1(new_n12011_), .A2(new_n12017_), .B(new_n12203_), .ZN(new_n12204_));
  INV_X1     g11202(.I(new_n12204_), .ZN(new_n12205_));
  NOR3_X1    g11203(.A1(new_n12054_), .A2(new_n12202_), .A3(new_n12205_), .ZN(new_n12206_));
  XOR2_X1    g11204(.A1(new_n12018_), .A2(new_n12011_), .Z(new_n12207_));
  OAI21_X1   g11205(.A1(new_n12055_), .A2(new_n12058_), .B(new_n12207_), .ZN(new_n12208_));
  AOI21_X1   g11206(.A1(new_n12208_), .A2(new_n12059_), .B(new_n12204_), .ZN(new_n12209_));
  NOR3_X1    g11207(.A1(new_n12206_), .A2(new_n12209_), .A3(new_n12201_), .ZN(new_n12210_));
  NAND3_X1   g11208(.A1(new_n12208_), .A2(new_n12059_), .A3(new_n12204_), .ZN(new_n12211_));
  OAI21_X1   g11209(.A1(new_n12054_), .A2(new_n12202_), .B(new_n12205_), .ZN(new_n12212_));
  AOI21_X1   g11210(.A1(new_n12212_), .A2(new_n12211_), .B(new_n12200_), .ZN(new_n12213_));
  OAI21_X1   g11211(.A1(new_n12210_), .A2(new_n12213_), .B(new_n12196_), .ZN(new_n12214_));
  AOI21_X1   g11212(.A1(new_n12191_), .A2(new_n12164_), .B(new_n12194_), .ZN(new_n12215_));
  NOR3_X1    g11213(.A1(new_n12175_), .A2(new_n12169_), .A3(new_n12189_), .ZN(new_n12216_));
  NOR2_X1    g11214(.A1(new_n12216_), .A2(new_n12215_), .ZN(new_n12217_));
  NAND3_X1   g11215(.A1(new_n12212_), .A2(new_n12211_), .A3(new_n12200_), .ZN(new_n12218_));
  OAI21_X1   g11216(.A1(new_n12206_), .A2(new_n12209_), .B(new_n12201_), .ZN(new_n12219_));
  NAND3_X1   g11217(.A1(new_n12219_), .A2(new_n12218_), .A3(new_n12217_), .ZN(new_n12220_));
  NAND3_X1   g11218(.A1(new_n12220_), .A2(new_n12214_), .A3(new_n12173_), .ZN(new_n12221_));
  NOR2_X1    g11219(.A1(new_n12055_), .A2(new_n12058_), .ZN(new_n12222_));
  NOR2_X1    g11220(.A1(new_n12202_), .A2(new_n12222_), .ZN(new_n12223_));
  OAI22_X1   g11221(.A1(new_n12223_), .A2(new_n12207_), .B1(new_n12208_), .B2(new_n12202_), .ZN(new_n12224_));
  NOR3_X1    g11222(.A1(new_n12167_), .A2(new_n12169_), .A3(new_n12166_), .ZN(new_n12225_));
  AOI21_X1   g11223(.A1(new_n12164_), .A2(new_n12162_), .B(new_n12155_), .ZN(new_n12226_));
  OAI21_X1   g11224(.A1(new_n12225_), .A2(new_n12226_), .B(new_n12147_), .ZN(new_n12227_));
  NOR3_X1    g11225(.A1(new_n12225_), .A2(new_n12147_), .A3(new_n12226_), .ZN(new_n12228_));
  AOI21_X1   g11226(.A1(new_n12224_), .A2(new_n12227_), .B(new_n12228_), .ZN(new_n12229_));
  AOI21_X1   g11227(.A1(new_n12219_), .A2(new_n12218_), .B(new_n12217_), .ZN(new_n12230_));
  NOR3_X1    g11228(.A1(new_n12210_), .A2(new_n12213_), .A3(new_n12196_), .ZN(new_n12231_));
  OAI21_X1   g11229(.A1(new_n12230_), .A2(new_n12231_), .B(new_n12229_), .ZN(new_n12232_));
  NAND4_X1   g11230(.A1(new_n11990_), .A2(new_n11978_), .A3(new_n12232_), .A4(new_n12221_), .ZN(new_n12233_));
  NOR3_X1    g11231(.A1(new_n11979_), .A2(new_n11980_), .A3(new_n11989_), .ZN(new_n12234_));
  AOI21_X1   g11232(.A1(new_n11960_), .A2(new_n11954_), .B(new_n11977_), .ZN(new_n12235_));
  NOR3_X1    g11233(.A1(new_n12230_), .A2(new_n12231_), .A3(new_n12229_), .ZN(new_n12236_));
  AOI21_X1   g11234(.A1(new_n12220_), .A2(new_n12214_), .B(new_n12173_), .ZN(new_n12237_));
  OAI22_X1   g11235(.A1(new_n12234_), .A2(new_n12235_), .B1(new_n12237_), .B2(new_n12236_), .ZN(new_n12238_));
  NAND3_X1   g11236(.A1(new_n12224_), .A2(new_n12172_), .A3(new_n12227_), .ZN(new_n12239_));
  OAI21_X1   g11237(.A1(new_n12171_), .A2(new_n12228_), .B(new_n12062_), .ZN(new_n12240_));
  NAND2_X1   g11238(.A1(new_n12240_), .A2(new_n12239_), .ZN(new_n12241_));
  NOR3_X1    g11239(.A1(new_n11988_), .A2(new_n11975_), .A3(new_n11983_), .ZN(new_n12242_));
  AOI21_X1   g11240(.A1(new_n11987_), .A2(new_n11976_), .B(new_n11965_), .ZN(new_n12243_));
  AND4_X2    g11241(.A1(new_n12137_), .A2(new_n12145_), .A3(new_n12144_), .A4(new_n12146_), .Z(new_n12244_));
  NOR2_X1    g11242(.A1(new_n12244_), .A2(new_n12147_), .ZN(new_n12245_));
  NOR2_X1    g11243(.A1(new_n11970_), .A2(new_n11973_), .ZN(new_n12246_));
  NOR2_X1    g11244(.A1(new_n12246_), .A2(new_n11986_), .ZN(new_n12247_));
  NAND2_X1   g11245(.A1(new_n12247_), .A2(new_n12245_), .ZN(new_n12248_));
  NOR3_X1    g11246(.A1(new_n12242_), .A2(new_n12243_), .A3(new_n12248_), .ZN(new_n12249_));
  OAI21_X1   g11247(.A1(new_n12242_), .A2(new_n12243_), .B(new_n12248_), .ZN(new_n12250_));
  OAI21_X1   g11248(.A1(new_n12241_), .A2(new_n12249_), .B(new_n12250_), .ZN(new_n12251_));
  NAND3_X1   g11249(.A1(new_n12238_), .A2(new_n12233_), .A3(new_n12251_), .ZN(new_n12252_));
  NOR4_X1    g11250(.A1(new_n12234_), .A2(new_n12235_), .A3(new_n12237_), .A4(new_n12236_), .ZN(new_n12253_));
  AOI22_X1   g11251(.A1(new_n11990_), .A2(new_n11978_), .B1(new_n12232_), .B2(new_n12221_), .ZN(new_n12254_));
  INV_X1     g11252(.I(new_n12241_), .ZN(new_n12255_));
  NAND3_X1   g11253(.A1(new_n11987_), .A2(new_n11976_), .A3(new_n11965_), .ZN(new_n12256_));
  OAI21_X1   g11254(.A1(new_n11988_), .A2(new_n11975_), .B(new_n11983_), .ZN(new_n12257_));
  INV_X1     g11255(.I(new_n12248_), .ZN(new_n12258_));
  NAND3_X1   g11256(.A1(new_n12257_), .A2(new_n12258_), .A3(new_n12256_), .ZN(new_n12259_));
  AOI21_X1   g11257(.A1(new_n12257_), .A2(new_n12256_), .B(new_n12258_), .ZN(new_n12260_));
  AOI21_X1   g11258(.A1(new_n12255_), .A2(new_n12259_), .B(new_n12260_), .ZN(new_n12261_));
  OAI21_X1   g11259(.A1(new_n12253_), .A2(new_n12254_), .B(new_n12261_), .ZN(new_n12262_));
  INV_X1     g11260(.I(\A[717] ), .ZN(new_n12263_));
  NOR2_X1    g11261(.A1(new_n12263_), .A2(\A[716] ), .ZN(new_n12264_));
  INV_X1     g11262(.I(\A[716] ), .ZN(new_n12265_));
  NOR2_X1    g11263(.A1(new_n12265_), .A2(\A[717] ), .ZN(new_n12266_));
  OAI21_X1   g11264(.A1(new_n12264_), .A2(new_n12266_), .B(\A[715] ), .ZN(new_n12267_));
  INV_X1     g11265(.I(\A[715] ), .ZN(new_n12268_));
  NAND2_X1   g11266(.A1(\A[716] ), .A2(\A[717] ), .ZN(new_n12269_));
  INV_X1     g11267(.I(new_n12269_), .ZN(new_n12270_));
  NOR2_X1    g11268(.A1(\A[716] ), .A2(\A[717] ), .ZN(new_n12271_));
  OAI21_X1   g11269(.A1(new_n12270_), .A2(new_n12271_), .B(new_n12268_), .ZN(new_n12272_));
  INV_X1     g11270(.I(\A[720] ), .ZN(new_n12273_));
  NOR2_X1    g11271(.A1(new_n12273_), .A2(\A[719] ), .ZN(new_n12274_));
  INV_X1     g11272(.I(\A[719] ), .ZN(new_n12275_));
  NOR2_X1    g11273(.A1(new_n12275_), .A2(\A[720] ), .ZN(new_n12276_));
  OAI21_X1   g11274(.A1(new_n12274_), .A2(new_n12276_), .B(\A[718] ), .ZN(new_n12277_));
  INV_X1     g11275(.I(\A[718] ), .ZN(new_n12278_));
  NAND2_X1   g11276(.A1(\A[719] ), .A2(\A[720] ), .ZN(new_n12279_));
  INV_X1     g11277(.I(new_n12279_), .ZN(new_n12280_));
  NOR2_X1    g11278(.A1(\A[719] ), .A2(\A[720] ), .ZN(new_n12281_));
  OAI21_X1   g11279(.A1(new_n12280_), .A2(new_n12281_), .B(new_n12278_), .ZN(new_n12282_));
  NAND4_X1   g11280(.A1(new_n12267_), .A2(new_n12272_), .A3(new_n12277_), .A4(new_n12282_), .ZN(new_n12283_));
  AOI21_X1   g11281(.A1(new_n12278_), .A2(new_n12279_), .B(new_n12281_), .ZN(new_n12284_));
  AOI21_X1   g11282(.A1(new_n12268_), .A2(new_n12269_), .B(new_n12271_), .ZN(new_n12285_));
  NOR2_X1    g11283(.A1(new_n12284_), .A2(new_n12285_), .ZN(new_n12286_));
  NAND2_X1   g11284(.A1(new_n12284_), .A2(new_n12285_), .ZN(new_n12287_));
  INV_X1     g11285(.I(new_n12287_), .ZN(new_n12288_));
  NOR2_X1    g11286(.A1(new_n12288_), .A2(new_n12286_), .ZN(new_n12289_));
  NAND2_X1   g11287(.A1(new_n12289_), .A2(new_n12283_), .ZN(new_n12290_));
  INV_X1     g11288(.I(new_n12283_), .ZN(new_n12291_));
  INV_X1     g11289(.I(new_n12286_), .ZN(new_n12292_));
  NAND2_X1   g11290(.A1(new_n12292_), .A2(new_n12287_), .ZN(new_n12293_));
  NAND2_X1   g11291(.A1(new_n12291_), .A2(new_n12293_), .ZN(new_n12294_));
  NAND2_X1   g11292(.A1(new_n12294_), .A2(new_n12290_), .ZN(new_n12295_));
  INV_X1     g11293(.I(\A[721] ), .ZN(new_n12296_));
  INV_X1     g11294(.I(\A[722] ), .ZN(new_n12297_));
  NAND2_X1   g11295(.A1(new_n12297_), .A2(\A[723] ), .ZN(new_n12298_));
  INV_X1     g11296(.I(\A[723] ), .ZN(new_n12299_));
  NAND2_X1   g11297(.A1(new_n12299_), .A2(\A[722] ), .ZN(new_n12300_));
  AOI21_X1   g11298(.A1(new_n12298_), .A2(new_n12300_), .B(new_n12296_), .ZN(new_n12301_));
  NAND2_X1   g11299(.A1(\A[722] ), .A2(\A[723] ), .ZN(new_n12302_));
  NOR2_X1    g11300(.A1(\A[722] ), .A2(\A[723] ), .ZN(new_n12303_));
  INV_X1     g11301(.I(new_n12303_), .ZN(new_n12304_));
  AOI21_X1   g11302(.A1(new_n12304_), .A2(new_n12302_), .B(\A[721] ), .ZN(new_n12305_));
  NOR2_X1    g11303(.A1(new_n12305_), .A2(new_n12301_), .ZN(new_n12306_));
  INV_X1     g11304(.I(\A[724] ), .ZN(new_n12307_));
  INV_X1     g11305(.I(\A[725] ), .ZN(new_n12308_));
  NAND2_X1   g11306(.A1(new_n12308_), .A2(\A[726] ), .ZN(new_n12309_));
  INV_X1     g11307(.I(\A[726] ), .ZN(new_n12310_));
  NAND2_X1   g11308(.A1(new_n12310_), .A2(\A[725] ), .ZN(new_n12311_));
  AOI21_X1   g11309(.A1(new_n12309_), .A2(new_n12311_), .B(new_n12307_), .ZN(new_n12312_));
  NAND2_X1   g11310(.A1(\A[725] ), .A2(\A[726] ), .ZN(new_n12313_));
  NOR2_X1    g11311(.A1(\A[725] ), .A2(\A[726] ), .ZN(new_n12314_));
  INV_X1     g11312(.I(new_n12314_), .ZN(new_n12315_));
  AOI21_X1   g11313(.A1(new_n12315_), .A2(new_n12313_), .B(\A[724] ), .ZN(new_n12316_));
  NOR2_X1    g11314(.A1(new_n12316_), .A2(new_n12312_), .ZN(new_n12317_));
  NAND2_X1   g11315(.A1(new_n12306_), .A2(new_n12317_), .ZN(new_n12318_));
  AOI21_X1   g11316(.A1(new_n12307_), .A2(new_n12313_), .B(new_n12314_), .ZN(new_n12319_));
  AOI21_X1   g11317(.A1(new_n12296_), .A2(new_n12302_), .B(new_n12303_), .ZN(new_n12320_));
  XOR2_X1    g11318(.A1(new_n12319_), .A2(new_n12320_), .Z(new_n12321_));
  NAND2_X1   g11319(.A1(new_n12318_), .A2(new_n12321_), .ZN(new_n12322_));
  NOR2_X1    g11320(.A1(new_n12299_), .A2(\A[722] ), .ZN(new_n12323_));
  NOR2_X1    g11321(.A1(new_n12297_), .A2(\A[723] ), .ZN(new_n12324_));
  OAI21_X1   g11322(.A1(new_n12323_), .A2(new_n12324_), .B(\A[721] ), .ZN(new_n12325_));
  INV_X1     g11323(.I(new_n12302_), .ZN(new_n12326_));
  OAI21_X1   g11324(.A1(new_n12326_), .A2(new_n12303_), .B(new_n12296_), .ZN(new_n12327_));
  NAND2_X1   g11325(.A1(new_n12325_), .A2(new_n12327_), .ZN(new_n12328_));
  NOR2_X1    g11326(.A1(new_n12310_), .A2(\A[725] ), .ZN(new_n12329_));
  NOR2_X1    g11327(.A1(new_n12308_), .A2(\A[726] ), .ZN(new_n12330_));
  OAI21_X1   g11328(.A1(new_n12329_), .A2(new_n12330_), .B(\A[724] ), .ZN(new_n12331_));
  INV_X1     g11329(.I(new_n12313_), .ZN(new_n12332_));
  OAI21_X1   g11330(.A1(new_n12332_), .A2(new_n12314_), .B(new_n12307_), .ZN(new_n12333_));
  NAND2_X1   g11331(.A1(new_n12331_), .A2(new_n12333_), .ZN(new_n12334_));
  NOR2_X1    g11332(.A1(new_n12328_), .A2(new_n12334_), .ZN(new_n12335_));
  XNOR2_X1   g11333(.A1(new_n12319_), .A2(new_n12320_), .ZN(new_n12336_));
  NAND2_X1   g11334(.A1(new_n12335_), .A2(new_n12336_), .ZN(new_n12337_));
  NAND2_X1   g11335(.A1(new_n12337_), .A2(new_n12322_), .ZN(new_n12338_));
  NAND2_X1   g11336(.A1(new_n12267_), .A2(new_n12272_), .ZN(new_n12339_));
  NAND2_X1   g11337(.A1(new_n12277_), .A2(new_n12282_), .ZN(new_n12340_));
  NAND2_X1   g11338(.A1(new_n12339_), .A2(new_n12340_), .ZN(new_n12341_));
  NAND2_X1   g11339(.A1(new_n12341_), .A2(new_n12283_), .ZN(new_n12342_));
  NAND2_X1   g11340(.A1(new_n12328_), .A2(new_n12334_), .ZN(new_n12343_));
  NAND2_X1   g11341(.A1(new_n12318_), .A2(new_n12343_), .ZN(new_n12344_));
  NOR2_X1    g11342(.A1(new_n12344_), .A2(new_n12342_), .ZN(new_n12345_));
  NOR2_X1    g11343(.A1(new_n12338_), .A2(new_n12345_), .ZN(new_n12346_));
  NOR2_X1    g11344(.A1(new_n12335_), .A2(new_n12336_), .ZN(new_n12347_));
  NOR2_X1    g11345(.A1(new_n12318_), .A2(new_n12321_), .ZN(new_n12348_));
  NOR2_X1    g11346(.A1(new_n12347_), .A2(new_n12348_), .ZN(new_n12349_));
  NOR2_X1    g11347(.A1(new_n12306_), .A2(new_n12317_), .ZN(new_n12350_));
  NOR2_X1    g11348(.A1(new_n12350_), .A2(new_n12335_), .ZN(new_n12351_));
  NAND3_X1   g11349(.A1(new_n12351_), .A2(new_n12283_), .A3(new_n12341_), .ZN(new_n12352_));
  NOR2_X1    g11350(.A1(new_n12352_), .A2(new_n12349_), .ZN(new_n12353_));
  NOR3_X1    g11351(.A1(new_n12353_), .A2(new_n12346_), .A3(new_n12295_), .ZN(new_n12354_));
  XOR2_X1    g11352(.A1(new_n12289_), .A2(new_n12283_), .Z(new_n12355_));
  NAND2_X1   g11353(.A1(new_n12352_), .A2(new_n12349_), .ZN(new_n12356_));
  INV_X1     g11354(.I(new_n12319_), .ZN(new_n12357_));
  INV_X1     g11355(.I(new_n12320_), .ZN(new_n12358_));
  NOR2_X1    g11356(.A1(new_n12357_), .A2(new_n12358_), .ZN(new_n12359_));
  NOR4_X1    g11357(.A1(new_n12322_), .A2(new_n12342_), .A3(new_n12350_), .A4(new_n12359_), .ZN(new_n12360_));
  INV_X1     g11358(.I(new_n12360_), .ZN(new_n12361_));
  AOI21_X1   g11359(.A1(new_n12356_), .A2(new_n12361_), .B(new_n12355_), .ZN(new_n12362_));
  OR2_X2     g11360(.A1(new_n12354_), .A2(new_n12362_), .Z(new_n12363_));
  INV_X1     g11361(.I(\A[703] ), .ZN(new_n12364_));
  INV_X1     g11362(.I(\A[704] ), .ZN(new_n12365_));
  NAND2_X1   g11363(.A1(new_n12365_), .A2(\A[705] ), .ZN(new_n12366_));
  INV_X1     g11364(.I(\A[705] ), .ZN(new_n12367_));
  NAND2_X1   g11365(.A1(new_n12367_), .A2(\A[704] ), .ZN(new_n12368_));
  AOI21_X1   g11366(.A1(new_n12366_), .A2(new_n12368_), .B(new_n12364_), .ZN(new_n12369_));
  NAND2_X1   g11367(.A1(\A[704] ), .A2(\A[705] ), .ZN(new_n12370_));
  NOR2_X1    g11368(.A1(\A[704] ), .A2(\A[705] ), .ZN(new_n12371_));
  INV_X1     g11369(.I(new_n12371_), .ZN(new_n12372_));
  AOI21_X1   g11370(.A1(new_n12372_), .A2(new_n12370_), .B(\A[703] ), .ZN(new_n12373_));
  INV_X1     g11371(.I(\A[706] ), .ZN(new_n12374_));
  INV_X1     g11372(.I(\A[707] ), .ZN(new_n12375_));
  NAND2_X1   g11373(.A1(new_n12375_), .A2(\A[708] ), .ZN(new_n12376_));
  INV_X1     g11374(.I(\A[708] ), .ZN(new_n12377_));
  NAND2_X1   g11375(.A1(new_n12377_), .A2(\A[707] ), .ZN(new_n12378_));
  AOI21_X1   g11376(.A1(new_n12376_), .A2(new_n12378_), .B(new_n12374_), .ZN(new_n12379_));
  NAND2_X1   g11377(.A1(\A[707] ), .A2(\A[708] ), .ZN(new_n12380_));
  NOR2_X1    g11378(.A1(\A[707] ), .A2(\A[708] ), .ZN(new_n12381_));
  INV_X1     g11379(.I(new_n12381_), .ZN(new_n12382_));
  AOI21_X1   g11380(.A1(new_n12382_), .A2(new_n12380_), .B(\A[706] ), .ZN(new_n12383_));
  NOR4_X1    g11381(.A1(new_n12369_), .A2(new_n12373_), .A3(new_n12383_), .A4(new_n12379_), .ZN(new_n12384_));
  AOI21_X1   g11382(.A1(new_n12374_), .A2(new_n12380_), .B(new_n12381_), .ZN(new_n12385_));
  AOI21_X1   g11383(.A1(new_n12364_), .A2(new_n12370_), .B(new_n12371_), .ZN(new_n12386_));
  XOR2_X1    g11384(.A1(new_n12385_), .A2(new_n12386_), .Z(new_n12387_));
  XNOR2_X1   g11385(.A1(new_n12387_), .A2(new_n12384_), .ZN(new_n12388_));
  INV_X1     g11386(.I(\A[709] ), .ZN(new_n12389_));
  INV_X1     g11387(.I(\A[710] ), .ZN(new_n12390_));
  NAND2_X1   g11388(.A1(new_n12390_), .A2(\A[711] ), .ZN(new_n12391_));
  INV_X1     g11389(.I(\A[711] ), .ZN(new_n12392_));
  NAND2_X1   g11390(.A1(new_n12392_), .A2(\A[710] ), .ZN(new_n12393_));
  AOI21_X1   g11391(.A1(new_n12391_), .A2(new_n12393_), .B(new_n12389_), .ZN(new_n12394_));
  NOR2_X1    g11392(.A1(\A[710] ), .A2(\A[711] ), .ZN(new_n12395_));
  INV_X1     g11393(.I(new_n12395_), .ZN(new_n12396_));
  NAND2_X1   g11394(.A1(\A[710] ), .A2(\A[711] ), .ZN(new_n12397_));
  AOI21_X1   g11395(.A1(new_n12396_), .A2(new_n12397_), .B(\A[709] ), .ZN(new_n12398_));
  NOR2_X1    g11396(.A1(new_n12398_), .A2(new_n12394_), .ZN(new_n12399_));
  INV_X1     g11397(.I(\A[712] ), .ZN(new_n12400_));
  INV_X1     g11398(.I(\A[713] ), .ZN(new_n12401_));
  NAND2_X1   g11399(.A1(new_n12401_), .A2(\A[714] ), .ZN(new_n12402_));
  INV_X1     g11400(.I(\A[714] ), .ZN(new_n12403_));
  NAND2_X1   g11401(.A1(new_n12403_), .A2(\A[713] ), .ZN(new_n12404_));
  AOI21_X1   g11402(.A1(new_n12402_), .A2(new_n12404_), .B(new_n12400_), .ZN(new_n12405_));
  NOR2_X1    g11403(.A1(\A[713] ), .A2(\A[714] ), .ZN(new_n12406_));
  INV_X1     g11404(.I(new_n12406_), .ZN(new_n12407_));
  NAND2_X1   g11405(.A1(\A[713] ), .A2(\A[714] ), .ZN(new_n12408_));
  AOI21_X1   g11406(.A1(new_n12407_), .A2(new_n12408_), .B(\A[712] ), .ZN(new_n12409_));
  NOR2_X1    g11407(.A1(new_n12409_), .A2(new_n12405_), .ZN(new_n12410_));
  NAND2_X1   g11408(.A1(new_n12399_), .A2(new_n12410_), .ZN(new_n12411_));
  AOI21_X1   g11409(.A1(new_n12400_), .A2(new_n12408_), .B(new_n12406_), .ZN(new_n12412_));
  AOI21_X1   g11410(.A1(new_n12389_), .A2(new_n12397_), .B(new_n12395_), .ZN(new_n12413_));
  XOR2_X1    g11411(.A1(new_n12412_), .A2(new_n12413_), .Z(new_n12414_));
  XOR2_X1    g11412(.A1(new_n12411_), .A2(new_n12414_), .Z(new_n12415_));
  NOR2_X1    g11413(.A1(new_n12392_), .A2(\A[710] ), .ZN(new_n12416_));
  NOR2_X1    g11414(.A1(new_n12390_), .A2(\A[711] ), .ZN(new_n12417_));
  OAI21_X1   g11415(.A1(new_n12416_), .A2(new_n12417_), .B(\A[709] ), .ZN(new_n12418_));
  INV_X1     g11416(.I(new_n12397_), .ZN(new_n12419_));
  OAI21_X1   g11417(.A1(new_n12419_), .A2(new_n12395_), .B(new_n12389_), .ZN(new_n12420_));
  NAND2_X1   g11418(.A1(new_n12418_), .A2(new_n12420_), .ZN(new_n12421_));
  NOR2_X1    g11419(.A1(new_n12403_), .A2(\A[713] ), .ZN(new_n12422_));
  NOR2_X1    g11420(.A1(new_n12401_), .A2(\A[714] ), .ZN(new_n12423_));
  OAI21_X1   g11421(.A1(new_n12422_), .A2(new_n12423_), .B(\A[712] ), .ZN(new_n12424_));
  INV_X1     g11422(.I(new_n12408_), .ZN(new_n12425_));
  OAI21_X1   g11423(.A1(new_n12425_), .A2(new_n12406_), .B(new_n12400_), .ZN(new_n12426_));
  NAND2_X1   g11424(.A1(new_n12424_), .A2(new_n12426_), .ZN(new_n12427_));
  NOR2_X1    g11425(.A1(new_n12421_), .A2(new_n12427_), .ZN(new_n12428_));
  NOR2_X1    g11426(.A1(new_n12399_), .A2(new_n12410_), .ZN(new_n12429_));
  NOR2_X1    g11427(.A1(new_n12429_), .A2(new_n12428_), .ZN(new_n12430_));
  OAI22_X1   g11428(.A1(new_n12369_), .A2(new_n12373_), .B1(new_n12383_), .B2(new_n12379_), .ZN(new_n12431_));
  INV_X1     g11429(.I(new_n12431_), .ZN(new_n12432_));
  NOR2_X1    g11430(.A1(new_n12432_), .A2(new_n12384_), .ZN(new_n12433_));
  NAND2_X1   g11431(.A1(new_n12433_), .A2(new_n12430_), .ZN(new_n12434_));
  AOI21_X1   g11432(.A1(new_n12415_), .A2(new_n12434_), .B(new_n12388_), .ZN(new_n12435_));
  XOR2_X1    g11433(.A1(new_n12428_), .A2(new_n12414_), .Z(new_n12436_));
  NAND2_X1   g11434(.A1(new_n12421_), .A2(new_n12427_), .ZN(new_n12437_));
  NAND2_X1   g11435(.A1(new_n12411_), .A2(new_n12437_), .ZN(new_n12438_));
  INV_X1     g11436(.I(new_n12384_), .ZN(new_n12439_));
  NAND2_X1   g11437(.A1(new_n12439_), .A2(new_n12431_), .ZN(new_n12440_));
  NOR2_X1    g11438(.A1(new_n12440_), .A2(new_n12438_), .ZN(new_n12441_));
  NAND2_X1   g11439(.A1(new_n12436_), .A2(new_n12441_), .ZN(new_n12442_));
  NAND2_X1   g11440(.A1(new_n12435_), .A2(new_n12442_), .ZN(new_n12443_));
  NOR2_X1    g11441(.A1(new_n12436_), .A2(new_n12441_), .ZN(new_n12444_));
  NOR2_X1    g11442(.A1(new_n12415_), .A2(new_n12434_), .ZN(new_n12445_));
  OAI21_X1   g11443(.A1(new_n12445_), .A2(new_n12444_), .B(new_n12388_), .ZN(new_n12446_));
  NAND2_X1   g11444(.A1(new_n12351_), .A2(new_n12342_), .ZN(new_n12447_));
  INV_X1     g11445(.I(new_n12342_), .ZN(new_n12448_));
  NAND2_X1   g11446(.A1(new_n12448_), .A2(new_n12344_), .ZN(new_n12449_));
  NAND2_X1   g11447(.A1(new_n12440_), .A2(new_n12430_), .ZN(new_n12450_));
  NAND2_X1   g11448(.A1(new_n12433_), .A2(new_n12438_), .ZN(new_n12451_));
  AOI22_X1   g11449(.A1(new_n12449_), .A2(new_n12447_), .B1(new_n12450_), .B2(new_n12451_), .ZN(new_n12452_));
  NAND3_X1   g11450(.A1(new_n12443_), .A2(new_n12446_), .A3(new_n12452_), .ZN(new_n12453_));
  XOR2_X1    g11451(.A1(new_n12387_), .A2(new_n12384_), .Z(new_n12454_));
  OAI21_X1   g11452(.A1(new_n12436_), .A2(new_n12441_), .B(new_n12454_), .ZN(new_n12455_));
  NOR2_X1    g11453(.A1(new_n12455_), .A2(new_n12445_), .ZN(new_n12456_));
  NAND2_X1   g11454(.A1(new_n12415_), .A2(new_n12434_), .ZN(new_n12457_));
  AOI21_X1   g11455(.A1(new_n12457_), .A2(new_n12442_), .B(new_n12454_), .ZN(new_n12458_));
  XOR2_X1    g11456(.A1(new_n12344_), .A2(new_n12342_), .Z(new_n12459_));
  NAND2_X1   g11457(.A1(new_n12450_), .A2(new_n12451_), .ZN(new_n12460_));
  NAND2_X1   g11458(.A1(new_n12459_), .A2(new_n12460_), .ZN(new_n12461_));
  OAI21_X1   g11459(.A1(new_n12458_), .A2(new_n12456_), .B(new_n12461_), .ZN(new_n12462_));
  NAND3_X1   g11460(.A1(new_n12363_), .A2(new_n12453_), .A3(new_n12462_), .ZN(new_n12463_));
  NOR2_X1    g11461(.A1(new_n12354_), .A2(new_n12362_), .ZN(new_n12464_));
  NOR3_X1    g11462(.A1(new_n12458_), .A2(new_n12456_), .A3(new_n12461_), .ZN(new_n12465_));
  AOI21_X1   g11463(.A1(new_n12443_), .A2(new_n12446_), .B(new_n12452_), .ZN(new_n12466_));
  OAI21_X1   g11464(.A1(new_n12466_), .A2(new_n12465_), .B(new_n12464_), .ZN(new_n12467_));
  AND2_X2    g11465(.A1(new_n12463_), .A2(new_n12467_), .Z(new_n12468_));
  INV_X1     g11466(.I(\A[741] ), .ZN(new_n12469_));
  NOR2_X1    g11467(.A1(new_n12469_), .A2(\A[740] ), .ZN(new_n12470_));
  INV_X1     g11468(.I(\A[740] ), .ZN(new_n12471_));
  NOR2_X1    g11469(.A1(new_n12471_), .A2(\A[741] ), .ZN(new_n12472_));
  OAI21_X1   g11470(.A1(new_n12470_), .A2(new_n12472_), .B(\A[739] ), .ZN(new_n12473_));
  INV_X1     g11471(.I(\A[739] ), .ZN(new_n12474_));
  NAND2_X1   g11472(.A1(\A[740] ), .A2(\A[741] ), .ZN(new_n12475_));
  INV_X1     g11473(.I(new_n12475_), .ZN(new_n12476_));
  NOR2_X1    g11474(.A1(\A[740] ), .A2(\A[741] ), .ZN(new_n12477_));
  OAI21_X1   g11475(.A1(new_n12476_), .A2(new_n12477_), .B(new_n12474_), .ZN(new_n12478_));
  INV_X1     g11476(.I(\A[744] ), .ZN(new_n12479_));
  NOR2_X1    g11477(.A1(new_n12479_), .A2(\A[743] ), .ZN(new_n12480_));
  INV_X1     g11478(.I(\A[743] ), .ZN(new_n12481_));
  NOR2_X1    g11479(.A1(new_n12481_), .A2(\A[744] ), .ZN(new_n12482_));
  OAI21_X1   g11480(.A1(new_n12480_), .A2(new_n12482_), .B(\A[742] ), .ZN(new_n12483_));
  INV_X1     g11481(.I(\A[742] ), .ZN(new_n12484_));
  NAND2_X1   g11482(.A1(\A[743] ), .A2(\A[744] ), .ZN(new_n12485_));
  INV_X1     g11483(.I(new_n12485_), .ZN(new_n12486_));
  NOR2_X1    g11484(.A1(\A[743] ), .A2(\A[744] ), .ZN(new_n12487_));
  OAI21_X1   g11485(.A1(new_n12486_), .A2(new_n12487_), .B(new_n12484_), .ZN(new_n12488_));
  NAND4_X1   g11486(.A1(new_n12473_), .A2(new_n12478_), .A3(new_n12483_), .A4(new_n12488_), .ZN(new_n12489_));
  NAND2_X1   g11487(.A1(new_n12473_), .A2(new_n12478_), .ZN(new_n12490_));
  NAND2_X1   g11488(.A1(new_n12483_), .A2(new_n12488_), .ZN(new_n12491_));
  NAND2_X1   g11489(.A1(new_n12490_), .A2(new_n12491_), .ZN(new_n12492_));
  NAND2_X1   g11490(.A1(new_n12492_), .A2(new_n12489_), .ZN(new_n12493_));
  INV_X1     g11491(.I(new_n12493_), .ZN(new_n12494_));
  INV_X1     g11492(.I(\A[745] ), .ZN(new_n12495_));
  INV_X1     g11493(.I(\A[746] ), .ZN(new_n12496_));
  NAND2_X1   g11494(.A1(new_n12496_), .A2(\A[747] ), .ZN(new_n12497_));
  INV_X1     g11495(.I(\A[747] ), .ZN(new_n12498_));
  NAND2_X1   g11496(.A1(new_n12498_), .A2(\A[746] ), .ZN(new_n12499_));
  AOI21_X1   g11497(.A1(new_n12497_), .A2(new_n12499_), .B(new_n12495_), .ZN(new_n12500_));
  NAND2_X1   g11498(.A1(\A[746] ), .A2(\A[747] ), .ZN(new_n12501_));
  NOR2_X1    g11499(.A1(\A[746] ), .A2(\A[747] ), .ZN(new_n12502_));
  INV_X1     g11500(.I(new_n12502_), .ZN(new_n12503_));
  AOI21_X1   g11501(.A1(new_n12503_), .A2(new_n12501_), .B(\A[745] ), .ZN(new_n12504_));
  NOR2_X1    g11502(.A1(new_n12504_), .A2(new_n12500_), .ZN(new_n12505_));
  INV_X1     g11503(.I(\A[748] ), .ZN(new_n12506_));
  INV_X1     g11504(.I(\A[749] ), .ZN(new_n12507_));
  NAND2_X1   g11505(.A1(new_n12507_), .A2(\A[750] ), .ZN(new_n12508_));
  INV_X1     g11506(.I(\A[750] ), .ZN(new_n12509_));
  NAND2_X1   g11507(.A1(new_n12509_), .A2(\A[749] ), .ZN(new_n12510_));
  AOI21_X1   g11508(.A1(new_n12508_), .A2(new_n12510_), .B(new_n12506_), .ZN(new_n12511_));
  NAND2_X1   g11509(.A1(\A[749] ), .A2(\A[750] ), .ZN(new_n12512_));
  NOR2_X1    g11510(.A1(\A[749] ), .A2(\A[750] ), .ZN(new_n12513_));
  INV_X1     g11511(.I(new_n12513_), .ZN(new_n12514_));
  AOI21_X1   g11512(.A1(new_n12514_), .A2(new_n12512_), .B(\A[748] ), .ZN(new_n12515_));
  NOR2_X1    g11513(.A1(new_n12515_), .A2(new_n12511_), .ZN(new_n12516_));
  NAND2_X1   g11514(.A1(new_n12505_), .A2(new_n12516_), .ZN(new_n12517_));
  NOR2_X1    g11515(.A1(new_n12498_), .A2(\A[746] ), .ZN(new_n12518_));
  NOR2_X1    g11516(.A1(new_n12496_), .A2(\A[747] ), .ZN(new_n12519_));
  OAI21_X1   g11517(.A1(new_n12518_), .A2(new_n12519_), .B(\A[745] ), .ZN(new_n12520_));
  INV_X1     g11518(.I(new_n12501_), .ZN(new_n12521_));
  OAI21_X1   g11519(.A1(new_n12521_), .A2(new_n12502_), .B(new_n12495_), .ZN(new_n12522_));
  NAND2_X1   g11520(.A1(new_n12520_), .A2(new_n12522_), .ZN(new_n12523_));
  NOR2_X1    g11521(.A1(new_n12509_), .A2(\A[749] ), .ZN(new_n12524_));
  NOR2_X1    g11522(.A1(new_n12507_), .A2(\A[750] ), .ZN(new_n12525_));
  OAI21_X1   g11523(.A1(new_n12524_), .A2(new_n12525_), .B(\A[748] ), .ZN(new_n12526_));
  INV_X1     g11524(.I(new_n12512_), .ZN(new_n12527_));
  OAI21_X1   g11525(.A1(new_n12527_), .A2(new_n12513_), .B(new_n12506_), .ZN(new_n12528_));
  NAND2_X1   g11526(.A1(new_n12526_), .A2(new_n12528_), .ZN(new_n12529_));
  NAND2_X1   g11527(.A1(new_n12523_), .A2(new_n12529_), .ZN(new_n12530_));
  NAND2_X1   g11528(.A1(new_n12517_), .A2(new_n12530_), .ZN(new_n12531_));
  NOR2_X1    g11529(.A1(new_n12494_), .A2(new_n12531_), .ZN(new_n12532_));
  NOR2_X1    g11530(.A1(new_n12523_), .A2(new_n12529_), .ZN(new_n12533_));
  INV_X1     g11531(.I(new_n12530_), .ZN(new_n12534_));
  NOR2_X1    g11532(.A1(new_n12534_), .A2(new_n12533_), .ZN(new_n12535_));
  NOR2_X1    g11533(.A1(new_n12535_), .A2(new_n12493_), .ZN(new_n12536_));
  NOR2_X1    g11534(.A1(new_n12536_), .A2(new_n12532_), .ZN(new_n12537_));
  INV_X1     g11535(.I(\A[727] ), .ZN(new_n12538_));
  INV_X1     g11536(.I(\A[728] ), .ZN(new_n12539_));
  NAND2_X1   g11537(.A1(new_n12539_), .A2(\A[729] ), .ZN(new_n12540_));
  INV_X1     g11538(.I(\A[729] ), .ZN(new_n12541_));
  NAND2_X1   g11539(.A1(new_n12541_), .A2(\A[728] ), .ZN(new_n12542_));
  AOI21_X1   g11540(.A1(new_n12540_), .A2(new_n12542_), .B(new_n12538_), .ZN(new_n12543_));
  NAND2_X1   g11541(.A1(\A[728] ), .A2(\A[729] ), .ZN(new_n12544_));
  NOR2_X1    g11542(.A1(\A[728] ), .A2(\A[729] ), .ZN(new_n12545_));
  INV_X1     g11543(.I(new_n12545_), .ZN(new_n12546_));
  AOI21_X1   g11544(.A1(new_n12546_), .A2(new_n12544_), .B(\A[727] ), .ZN(new_n12547_));
  INV_X1     g11545(.I(\A[730] ), .ZN(new_n12548_));
  INV_X1     g11546(.I(\A[731] ), .ZN(new_n12549_));
  NAND2_X1   g11547(.A1(new_n12549_), .A2(\A[732] ), .ZN(new_n12550_));
  INV_X1     g11548(.I(\A[732] ), .ZN(new_n12551_));
  NAND2_X1   g11549(.A1(new_n12551_), .A2(\A[731] ), .ZN(new_n12552_));
  AOI21_X1   g11550(.A1(new_n12550_), .A2(new_n12552_), .B(new_n12548_), .ZN(new_n12553_));
  NAND2_X1   g11551(.A1(\A[731] ), .A2(\A[732] ), .ZN(new_n12554_));
  NOR2_X1    g11552(.A1(\A[731] ), .A2(\A[732] ), .ZN(new_n12555_));
  INV_X1     g11553(.I(new_n12555_), .ZN(new_n12556_));
  AOI21_X1   g11554(.A1(new_n12556_), .A2(new_n12554_), .B(\A[730] ), .ZN(new_n12557_));
  NOR4_X1    g11555(.A1(new_n12543_), .A2(new_n12547_), .A3(new_n12557_), .A4(new_n12553_), .ZN(new_n12558_));
  OAI22_X1   g11556(.A1(new_n12543_), .A2(new_n12547_), .B1(new_n12557_), .B2(new_n12553_), .ZN(new_n12559_));
  INV_X1     g11557(.I(new_n12559_), .ZN(new_n12560_));
  NOR2_X1    g11558(.A1(new_n12560_), .A2(new_n12558_), .ZN(new_n12561_));
  INV_X1     g11559(.I(\A[733] ), .ZN(new_n12562_));
  INV_X1     g11560(.I(\A[734] ), .ZN(new_n12563_));
  NAND2_X1   g11561(.A1(new_n12563_), .A2(\A[735] ), .ZN(new_n12564_));
  INV_X1     g11562(.I(\A[735] ), .ZN(new_n12565_));
  NAND2_X1   g11563(.A1(new_n12565_), .A2(\A[734] ), .ZN(new_n12566_));
  AOI21_X1   g11564(.A1(new_n12564_), .A2(new_n12566_), .B(new_n12562_), .ZN(new_n12567_));
  NAND2_X1   g11565(.A1(\A[734] ), .A2(\A[735] ), .ZN(new_n12568_));
  NOR2_X1    g11566(.A1(\A[734] ), .A2(\A[735] ), .ZN(new_n12569_));
  INV_X1     g11567(.I(new_n12569_), .ZN(new_n12570_));
  AOI21_X1   g11568(.A1(new_n12570_), .A2(new_n12568_), .B(\A[733] ), .ZN(new_n12571_));
  NOR2_X1    g11569(.A1(new_n12571_), .A2(new_n12567_), .ZN(new_n12572_));
  INV_X1     g11570(.I(\A[736] ), .ZN(new_n12573_));
  INV_X1     g11571(.I(\A[737] ), .ZN(new_n12574_));
  NAND2_X1   g11572(.A1(new_n12574_), .A2(\A[738] ), .ZN(new_n12575_));
  INV_X1     g11573(.I(\A[738] ), .ZN(new_n12576_));
  NAND2_X1   g11574(.A1(new_n12576_), .A2(\A[737] ), .ZN(new_n12577_));
  AOI21_X1   g11575(.A1(new_n12575_), .A2(new_n12577_), .B(new_n12573_), .ZN(new_n12578_));
  NAND2_X1   g11576(.A1(\A[737] ), .A2(\A[738] ), .ZN(new_n12579_));
  NOR2_X1    g11577(.A1(\A[737] ), .A2(\A[738] ), .ZN(new_n12580_));
  INV_X1     g11578(.I(new_n12580_), .ZN(new_n12581_));
  AOI21_X1   g11579(.A1(new_n12581_), .A2(new_n12579_), .B(\A[736] ), .ZN(new_n12582_));
  NOR2_X1    g11580(.A1(new_n12582_), .A2(new_n12578_), .ZN(new_n12583_));
  NAND2_X1   g11581(.A1(new_n12572_), .A2(new_n12583_), .ZN(new_n12584_));
  NOR2_X1    g11582(.A1(new_n12565_), .A2(\A[734] ), .ZN(new_n12585_));
  NOR2_X1    g11583(.A1(new_n12563_), .A2(\A[735] ), .ZN(new_n12586_));
  OAI21_X1   g11584(.A1(new_n12585_), .A2(new_n12586_), .B(\A[733] ), .ZN(new_n12587_));
  INV_X1     g11585(.I(new_n12568_), .ZN(new_n12588_));
  OAI21_X1   g11586(.A1(new_n12588_), .A2(new_n12569_), .B(new_n12562_), .ZN(new_n12589_));
  NAND2_X1   g11587(.A1(new_n12587_), .A2(new_n12589_), .ZN(new_n12590_));
  NOR2_X1    g11588(.A1(new_n12576_), .A2(\A[737] ), .ZN(new_n12591_));
  NOR2_X1    g11589(.A1(new_n12574_), .A2(\A[738] ), .ZN(new_n12592_));
  OAI21_X1   g11590(.A1(new_n12591_), .A2(new_n12592_), .B(\A[736] ), .ZN(new_n12593_));
  INV_X1     g11591(.I(new_n12579_), .ZN(new_n12594_));
  OAI21_X1   g11592(.A1(new_n12594_), .A2(new_n12580_), .B(new_n12573_), .ZN(new_n12595_));
  NAND2_X1   g11593(.A1(new_n12593_), .A2(new_n12595_), .ZN(new_n12596_));
  NAND2_X1   g11594(.A1(new_n12590_), .A2(new_n12596_), .ZN(new_n12597_));
  NAND2_X1   g11595(.A1(new_n12584_), .A2(new_n12597_), .ZN(new_n12598_));
  NOR2_X1    g11596(.A1(new_n12561_), .A2(new_n12598_), .ZN(new_n12599_));
  NOR2_X1    g11597(.A1(new_n12547_), .A2(new_n12543_), .ZN(new_n12600_));
  NOR2_X1    g11598(.A1(new_n12557_), .A2(new_n12553_), .ZN(new_n12601_));
  NAND2_X1   g11599(.A1(new_n12600_), .A2(new_n12601_), .ZN(new_n12602_));
  NAND2_X1   g11600(.A1(new_n12602_), .A2(new_n12559_), .ZN(new_n12603_));
  NOR2_X1    g11601(.A1(new_n12590_), .A2(new_n12596_), .ZN(new_n12604_));
  NOR2_X1    g11602(.A1(new_n12572_), .A2(new_n12583_), .ZN(new_n12605_));
  NOR2_X1    g11603(.A1(new_n12605_), .A2(new_n12604_), .ZN(new_n12606_));
  NOR2_X1    g11604(.A1(new_n12606_), .A2(new_n12603_), .ZN(new_n12607_));
  NOR2_X1    g11605(.A1(new_n12599_), .A2(new_n12607_), .ZN(new_n12608_));
  NOR2_X1    g11606(.A1(new_n12537_), .A2(new_n12608_), .ZN(new_n12609_));
  NOR4_X1    g11607(.A1(new_n12532_), .A2(new_n12536_), .A3(new_n12599_), .A4(new_n12607_), .ZN(new_n12610_));
  NOR2_X1    g11608(.A1(new_n12609_), .A2(new_n12610_), .ZN(new_n12611_));
  NOR2_X1    g11609(.A1(new_n12459_), .A2(new_n12460_), .ZN(new_n12612_));
  NOR2_X1    g11610(.A1(new_n12612_), .A2(new_n12452_), .ZN(new_n12613_));
  NAND2_X1   g11611(.A1(new_n12611_), .A2(new_n12613_), .ZN(new_n12614_));
  AOI21_X1   g11612(.A1(new_n12548_), .A2(new_n12554_), .B(new_n12555_), .ZN(new_n12615_));
  AOI21_X1   g11613(.A1(new_n12538_), .A2(new_n12544_), .B(new_n12545_), .ZN(new_n12616_));
  NOR2_X1    g11614(.A1(new_n12615_), .A2(new_n12616_), .ZN(new_n12617_));
  INV_X1     g11615(.I(new_n12617_), .ZN(new_n12618_));
  NAND2_X1   g11616(.A1(new_n12615_), .A2(new_n12616_), .ZN(new_n12619_));
  NAND2_X1   g11617(.A1(new_n12618_), .A2(new_n12619_), .ZN(new_n12620_));
  NOR2_X1    g11618(.A1(new_n12620_), .A2(new_n12558_), .ZN(new_n12621_));
  INV_X1     g11619(.I(new_n12619_), .ZN(new_n12622_));
  NOR2_X1    g11620(.A1(new_n12622_), .A2(new_n12617_), .ZN(new_n12623_));
  NOR2_X1    g11621(.A1(new_n12623_), .A2(new_n12602_), .ZN(new_n12624_));
  NOR2_X1    g11622(.A1(new_n12624_), .A2(new_n12621_), .ZN(new_n12625_));
  AOI21_X1   g11623(.A1(new_n12573_), .A2(new_n12579_), .B(new_n12580_), .ZN(new_n12626_));
  AOI21_X1   g11624(.A1(new_n12562_), .A2(new_n12568_), .B(new_n12569_), .ZN(new_n12627_));
  XNOR2_X1   g11625(.A1(new_n12626_), .A2(new_n12627_), .ZN(new_n12628_));
  NOR2_X1    g11626(.A1(new_n12604_), .A2(new_n12628_), .ZN(new_n12629_));
  XOR2_X1    g11627(.A1(new_n12626_), .A2(new_n12627_), .Z(new_n12630_));
  NOR2_X1    g11628(.A1(new_n12584_), .A2(new_n12630_), .ZN(new_n12631_));
  NOR2_X1    g11629(.A1(new_n12629_), .A2(new_n12631_), .ZN(new_n12632_));
  NAND2_X1   g11630(.A1(new_n12561_), .A2(new_n12606_), .ZN(new_n12633_));
  AOI21_X1   g11631(.A1(new_n12632_), .A2(new_n12633_), .B(new_n12625_), .ZN(new_n12634_));
  NAND2_X1   g11632(.A1(new_n12626_), .A2(new_n12627_), .ZN(new_n12635_));
  NAND4_X1   g11633(.A1(new_n12561_), .A2(new_n12629_), .A3(new_n12597_), .A4(new_n12635_), .ZN(new_n12636_));
  NOR2_X1    g11634(.A1(new_n12598_), .A2(new_n12603_), .ZN(new_n12637_));
  XOR2_X1    g11635(.A1(new_n12632_), .A2(new_n12637_), .Z(new_n12638_));
  AOI22_X1   g11636(.A1(new_n12638_), .A2(new_n12625_), .B1(new_n12634_), .B2(new_n12636_), .ZN(new_n12639_));
  OAI22_X1   g11637(.A1(new_n12536_), .A2(new_n12532_), .B1(new_n12599_), .B2(new_n12607_), .ZN(new_n12640_));
  INV_X1     g11638(.I(new_n12489_), .ZN(new_n12641_));
  AOI21_X1   g11639(.A1(new_n12484_), .A2(new_n12485_), .B(new_n12487_), .ZN(new_n12642_));
  AOI21_X1   g11640(.A1(new_n12474_), .A2(new_n12475_), .B(new_n12477_), .ZN(new_n12643_));
  NOR2_X1    g11641(.A1(new_n12642_), .A2(new_n12643_), .ZN(new_n12644_));
  INV_X1     g11642(.I(new_n12644_), .ZN(new_n12645_));
  NAND2_X1   g11643(.A1(new_n12642_), .A2(new_n12643_), .ZN(new_n12646_));
  NAND2_X1   g11644(.A1(new_n12645_), .A2(new_n12646_), .ZN(new_n12647_));
  NOR2_X1    g11645(.A1(new_n12641_), .A2(new_n12647_), .ZN(new_n12648_));
  INV_X1     g11646(.I(new_n12646_), .ZN(new_n12649_));
  NOR2_X1    g11647(.A1(new_n12649_), .A2(new_n12644_), .ZN(new_n12650_));
  NOR2_X1    g11648(.A1(new_n12650_), .A2(new_n12489_), .ZN(new_n12651_));
  NOR2_X1    g11649(.A1(new_n12648_), .A2(new_n12651_), .ZN(new_n12652_));
  AOI21_X1   g11650(.A1(new_n12506_), .A2(new_n12512_), .B(new_n12513_), .ZN(new_n12653_));
  AOI21_X1   g11651(.A1(new_n12495_), .A2(new_n12501_), .B(new_n12502_), .ZN(new_n12654_));
  XNOR2_X1   g11652(.A1(new_n12653_), .A2(new_n12654_), .ZN(new_n12655_));
  NOR2_X1    g11653(.A1(new_n12533_), .A2(new_n12655_), .ZN(new_n12656_));
  XOR2_X1    g11654(.A1(new_n12653_), .A2(new_n12654_), .Z(new_n12657_));
  NOR2_X1    g11655(.A1(new_n12517_), .A2(new_n12657_), .ZN(new_n12658_));
  NOR2_X1    g11656(.A1(new_n12656_), .A2(new_n12658_), .ZN(new_n12659_));
  NAND4_X1   g11657(.A1(new_n12492_), .A2(new_n12517_), .A3(new_n12530_), .A4(new_n12489_), .ZN(new_n12660_));
  NAND2_X1   g11658(.A1(new_n12659_), .A2(new_n12660_), .ZN(new_n12661_));
  NAND2_X1   g11659(.A1(new_n12517_), .A2(new_n12657_), .ZN(new_n12662_));
  NAND2_X1   g11660(.A1(new_n12533_), .A2(new_n12655_), .ZN(new_n12663_));
  NAND2_X1   g11661(.A1(new_n12663_), .A2(new_n12662_), .ZN(new_n12664_));
  INV_X1     g11662(.I(new_n12660_), .ZN(new_n12665_));
  NAND2_X1   g11663(.A1(new_n12665_), .A2(new_n12664_), .ZN(new_n12666_));
  NAND3_X1   g11664(.A1(new_n12666_), .A2(new_n12661_), .A3(new_n12652_), .ZN(new_n12667_));
  NAND2_X1   g11665(.A1(new_n12650_), .A2(new_n12489_), .ZN(new_n12668_));
  NAND2_X1   g11666(.A1(new_n12641_), .A2(new_n12647_), .ZN(new_n12669_));
  NAND2_X1   g11667(.A1(new_n12669_), .A2(new_n12668_), .ZN(new_n12670_));
  NOR2_X1    g11668(.A1(new_n12665_), .A2(new_n12664_), .ZN(new_n12671_));
  INV_X1     g11669(.I(new_n12653_), .ZN(new_n12672_));
  INV_X1     g11670(.I(new_n12654_), .ZN(new_n12673_));
  NOR2_X1    g11671(.A1(new_n12672_), .A2(new_n12673_), .ZN(new_n12674_));
  NOR4_X1    g11672(.A1(new_n12662_), .A2(new_n12493_), .A3(new_n12534_), .A4(new_n12674_), .ZN(new_n12675_));
  OAI21_X1   g11673(.A1(new_n12671_), .A2(new_n12675_), .B(new_n12670_), .ZN(new_n12676_));
  AOI21_X1   g11674(.A1(new_n12676_), .A2(new_n12667_), .B(new_n12640_), .ZN(new_n12677_));
  NOR2_X1    g11675(.A1(new_n12659_), .A2(new_n12660_), .ZN(new_n12678_));
  NOR3_X1    g11676(.A1(new_n12671_), .A2(new_n12678_), .A3(new_n12670_), .ZN(new_n12679_));
  INV_X1     g11677(.I(new_n12675_), .ZN(new_n12680_));
  AOI21_X1   g11678(.A1(new_n12680_), .A2(new_n12661_), .B(new_n12652_), .ZN(new_n12681_));
  NOR3_X1    g11679(.A1(new_n12609_), .A2(new_n12679_), .A3(new_n12681_), .ZN(new_n12682_));
  OAI21_X1   g11680(.A1(new_n12677_), .A2(new_n12682_), .B(new_n12639_), .ZN(new_n12683_));
  NAND2_X1   g11681(.A1(new_n12623_), .A2(new_n12602_), .ZN(new_n12684_));
  NAND2_X1   g11682(.A1(new_n12620_), .A2(new_n12558_), .ZN(new_n12685_));
  NAND2_X1   g11683(.A1(new_n12684_), .A2(new_n12685_), .ZN(new_n12686_));
  NAND2_X1   g11684(.A1(new_n12584_), .A2(new_n12630_), .ZN(new_n12687_));
  NAND2_X1   g11685(.A1(new_n12604_), .A2(new_n12628_), .ZN(new_n12688_));
  NAND2_X1   g11686(.A1(new_n12688_), .A2(new_n12687_), .ZN(new_n12689_));
  OAI21_X1   g11687(.A1(new_n12689_), .A2(new_n12637_), .B(new_n12686_), .ZN(new_n12690_));
  INV_X1     g11688(.I(new_n12636_), .ZN(new_n12691_));
  XOR2_X1    g11689(.A1(new_n12689_), .A2(new_n12637_), .Z(new_n12692_));
  OAI22_X1   g11690(.A1(new_n12692_), .A2(new_n12686_), .B1(new_n12690_), .B2(new_n12691_), .ZN(new_n12693_));
  OAI21_X1   g11691(.A1(new_n12679_), .A2(new_n12681_), .B(new_n12609_), .ZN(new_n12694_));
  NAND3_X1   g11692(.A1(new_n12676_), .A2(new_n12667_), .A3(new_n12640_), .ZN(new_n12695_));
  NAND3_X1   g11693(.A1(new_n12694_), .A2(new_n12693_), .A3(new_n12695_), .ZN(new_n12696_));
  AOI21_X1   g11694(.A1(new_n12683_), .A2(new_n12696_), .B(new_n12614_), .ZN(new_n12697_));
  NAND3_X1   g11695(.A1(new_n12683_), .A2(new_n12696_), .A3(new_n12614_), .ZN(new_n12698_));
  OAI21_X1   g11696(.A1(new_n12468_), .A2(new_n12697_), .B(new_n12698_), .ZN(new_n12699_));
  AOI21_X1   g11697(.A1(new_n12349_), .A2(new_n12352_), .B(new_n12355_), .ZN(new_n12700_));
  INV_X1     g11698(.I(new_n12359_), .ZN(new_n12701_));
  NOR2_X1    g11699(.A1(new_n12319_), .A2(new_n12320_), .ZN(new_n12702_));
  AOI21_X1   g11700(.A1(new_n12318_), .A2(new_n12701_), .B(new_n12702_), .ZN(new_n12703_));
  AOI21_X1   g11701(.A1(new_n12283_), .A2(new_n12287_), .B(new_n12286_), .ZN(new_n12704_));
  NOR2_X1    g11702(.A1(new_n12703_), .A2(new_n12704_), .ZN(new_n12705_));
  INV_X1     g11703(.I(new_n12702_), .ZN(new_n12706_));
  OAI21_X1   g11704(.A1(new_n12335_), .A2(new_n12359_), .B(new_n12706_), .ZN(new_n12707_));
  INV_X1     g11705(.I(new_n12704_), .ZN(new_n12708_));
  NOR2_X1    g11706(.A1(new_n12708_), .A2(new_n12707_), .ZN(new_n12709_));
  NOR2_X1    g11707(.A1(new_n12709_), .A2(new_n12705_), .ZN(new_n12710_));
  OAI21_X1   g11708(.A1(new_n12700_), .A2(new_n12360_), .B(new_n12710_), .ZN(new_n12711_));
  OAI21_X1   g11709(.A1(new_n12338_), .A2(new_n12345_), .B(new_n12295_), .ZN(new_n12712_));
  NAND2_X1   g11710(.A1(new_n12708_), .A2(new_n12707_), .ZN(new_n12713_));
  NAND2_X1   g11711(.A1(new_n12703_), .A2(new_n12704_), .ZN(new_n12714_));
  NAND2_X1   g11712(.A1(new_n12713_), .A2(new_n12714_), .ZN(new_n12715_));
  NAND3_X1   g11713(.A1(new_n12712_), .A2(new_n12715_), .A3(new_n12361_), .ZN(new_n12716_));
  NAND2_X1   g11714(.A1(new_n12711_), .A2(new_n12716_), .ZN(new_n12717_));
  AND2_X2    g11715(.A1(new_n12412_), .A2(new_n12413_), .Z(new_n12718_));
  NOR2_X1    g11716(.A1(new_n12412_), .A2(new_n12413_), .ZN(new_n12719_));
  INV_X1     g11717(.I(new_n12719_), .ZN(new_n12720_));
  OAI21_X1   g11718(.A1(new_n12428_), .A2(new_n12718_), .B(new_n12720_), .ZN(new_n12721_));
  NOR2_X1    g11719(.A1(new_n12385_), .A2(new_n12386_), .ZN(new_n12722_));
  NAND2_X1   g11720(.A1(new_n12385_), .A2(new_n12386_), .ZN(new_n12723_));
  AOI21_X1   g11721(.A1(new_n12439_), .A2(new_n12723_), .B(new_n12722_), .ZN(new_n12724_));
  NOR3_X1    g11722(.A1(new_n12435_), .A2(new_n12445_), .A3(new_n12724_), .ZN(new_n12725_));
  INV_X1     g11723(.I(new_n12724_), .ZN(new_n12726_));
  AOI21_X1   g11724(.A1(new_n12455_), .A2(new_n12442_), .B(new_n12726_), .ZN(new_n12727_));
  NOR3_X1    g11725(.A1(new_n12725_), .A2(new_n12727_), .A3(new_n12721_), .ZN(new_n12728_));
  INV_X1     g11726(.I(new_n12721_), .ZN(new_n12729_));
  NAND3_X1   g11727(.A1(new_n12455_), .A2(new_n12442_), .A3(new_n12726_), .ZN(new_n12730_));
  OAI21_X1   g11728(.A1(new_n12435_), .A2(new_n12445_), .B(new_n12724_), .ZN(new_n12731_));
  AOI21_X1   g11729(.A1(new_n12731_), .A2(new_n12730_), .B(new_n12729_), .ZN(new_n12732_));
  OAI21_X1   g11730(.A1(new_n12728_), .A2(new_n12732_), .B(new_n12717_), .ZN(new_n12733_));
  AOI21_X1   g11731(.A1(new_n12712_), .A2(new_n12361_), .B(new_n12715_), .ZN(new_n12734_));
  NOR3_X1    g11732(.A1(new_n12700_), .A2(new_n12360_), .A3(new_n12710_), .ZN(new_n12735_));
  NOR2_X1    g11733(.A1(new_n12735_), .A2(new_n12734_), .ZN(new_n12736_));
  NAND3_X1   g11734(.A1(new_n12731_), .A2(new_n12730_), .A3(new_n12729_), .ZN(new_n12737_));
  OAI21_X1   g11735(.A1(new_n12725_), .A2(new_n12727_), .B(new_n12721_), .ZN(new_n12738_));
  NAND3_X1   g11736(.A1(new_n12738_), .A2(new_n12737_), .A3(new_n12736_), .ZN(new_n12739_));
  OAI21_X1   g11737(.A1(new_n12363_), .A2(new_n12465_), .B(new_n12462_), .ZN(new_n12740_));
  NAND3_X1   g11738(.A1(new_n12733_), .A2(new_n12739_), .A3(new_n12740_), .ZN(new_n12741_));
  AOI21_X1   g11739(.A1(new_n12738_), .A2(new_n12737_), .B(new_n12736_), .ZN(new_n12742_));
  NOR3_X1    g11740(.A1(new_n12728_), .A2(new_n12732_), .A3(new_n12717_), .ZN(new_n12743_));
  AOI21_X1   g11741(.A1(new_n12464_), .A2(new_n12453_), .B(new_n12466_), .ZN(new_n12744_));
  OAI21_X1   g11742(.A1(new_n12742_), .A2(new_n12743_), .B(new_n12744_), .ZN(new_n12745_));
  OAI21_X1   g11743(.A1(new_n12639_), .A2(new_n12677_), .B(new_n12695_), .ZN(new_n12746_));
  AOI21_X1   g11744(.A1(new_n12659_), .A2(new_n12660_), .B(new_n12652_), .ZN(new_n12747_));
  INV_X1     g11745(.I(new_n12674_), .ZN(new_n12748_));
  NOR2_X1    g11746(.A1(new_n12653_), .A2(new_n12654_), .ZN(new_n12749_));
  AOI21_X1   g11747(.A1(new_n12517_), .A2(new_n12748_), .B(new_n12749_), .ZN(new_n12750_));
  AOI21_X1   g11748(.A1(new_n12489_), .A2(new_n12646_), .B(new_n12644_), .ZN(new_n12751_));
  NOR2_X1    g11749(.A1(new_n12750_), .A2(new_n12751_), .ZN(new_n12752_));
  INV_X1     g11750(.I(new_n12749_), .ZN(new_n12753_));
  OAI21_X1   g11751(.A1(new_n12533_), .A2(new_n12674_), .B(new_n12753_), .ZN(new_n12754_));
  INV_X1     g11752(.I(new_n12751_), .ZN(new_n12755_));
  NOR2_X1    g11753(.A1(new_n12755_), .A2(new_n12754_), .ZN(new_n12756_));
  NOR2_X1    g11754(.A1(new_n12756_), .A2(new_n12752_), .ZN(new_n12757_));
  OAI21_X1   g11755(.A1(new_n12747_), .A2(new_n12675_), .B(new_n12757_), .ZN(new_n12758_));
  OAI21_X1   g11756(.A1(new_n12665_), .A2(new_n12664_), .B(new_n12670_), .ZN(new_n12759_));
  NAND2_X1   g11757(.A1(new_n12755_), .A2(new_n12754_), .ZN(new_n12760_));
  NAND2_X1   g11758(.A1(new_n12750_), .A2(new_n12751_), .ZN(new_n12761_));
  NAND2_X1   g11759(.A1(new_n12760_), .A2(new_n12761_), .ZN(new_n12762_));
  NAND3_X1   g11760(.A1(new_n12759_), .A2(new_n12762_), .A3(new_n12680_), .ZN(new_n12763_));
  NAND2_X1   g11761(.A1(new_n12758_), .A2(new_n12763_), .ZN(new_n12764_));
  NOR2_X1    g11762(.A1(new_n12626_), .A2(new_n12627_), .ZN(new_n12765_));
  AOI21_X1   g11763(.A1(new_n12584_), .A2(new_n12635_), .B(new_n12765_), .ZN(new_n12766_));
  INV_X1     g11764(.I(new_n12766_), .ZN(new_n12767_));
  AOI21_X1   g11765(.A1(new_n12602_), .A2(new_n12619_), .B(new_n12617_), .ZN(new_n12768_));
  NOR3_X1    g11766(.A1(new_n12634_), .A2(new_n12691_), .A3(new_n12768_), .ZN(new_n12769_));
  INV_X1     g11767(.I(new_n12768_), .ZN(new_n12770_));
  AOI21_X1   g11768(.A1(new_n12690_), .A2(new_n12636_), .B(new_n12770_), .ZN(new_n12771_));
  NOR3_X1    g11769(.A1(new_n12769_), .A2(new_n12771_), .A3(new_n12767_), .ZN(new_n12772_));
  NAND3_X1   g11770(.A1(new_n12690_), .A2(new_n12636_), .A3(new_n12770_), .ZN(new_n12773_));
  OAI21_X1   g11771(.A1(new_n12634_), .A2(new_n12691_), .B(new_n12768_), .ZN(new_n12774_));
  AOI21_X1   g11772(.A1(new_n12774_), .A2(new_n12773_), .B(new_n12766_), .ZN(new_n12775_));
  OAI21_X1   g11773(.A1(new_n12772_), .A2(new_n12775_), .B(new_n12764_), .ZN(new_n12776_));
  AOI21_X1   g11774(.A1(new_n12661_), .A2(new_n12670_), .B(new_n12675_), .ZN(new_n12777_));
  NOR2_X1    g11775(.A1(new_n12777_), .A2(new_n12762_), .ZN(new_n12778_));
  NOR3_X1    g11776(.A1(new_n12747_), .A2(new_n12757_), .A3(new_n12675_), .ZN(new_n12779_));
  NOR2_X1    g11777(.A1(new_n12778_), .A2(new_n12779_), .ZN(new_n12780_));
  NAND3_X1   g11778(.A1(new_n12774_), .A2(new_n12773_), .A3(new_n12766_), .ZN(new_n12781_));
  OAI21_X1   g11779(.A1(new_n12769_), .A2(new_n12771_), .B(new_n12767_), .ZN(new_n12782_));
  NAND3_X1   g11780(.A1(new_n12780_), .A2(new_n12782_), .A3(new_n12781_), .ZN(new_n12783_));
  NAND3_X1   g11781(.A1(new_n12783_), .A2(new_n12776_), .A3(new_n12746_), .ZN(new_n12784_));
  AOI21_X1   g11782(.A1(new_n12694_), .A2(new_n12693_), .B(new_n12682_), .ZN(new_n12785_));
  AOI21_X1   g11783(.A1(new_n12781_), .A2(new_n12782_), .B(new_n12780_), .ZN(new_n12786_));
  NOR3_X1    g11784(.A1(new_n12772_), .A2(new_n12775_), .A3(new_n12764_), .ZN(new_n12787_));
  OAI21_X1   g11785(.A1(new_n12786_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n12788_));
  NAND4_X1   g11786(.A1(new_n12745_), .A2(new_n12741_), .A3(new_n12788_), .A4(new_n12784_), .ZN(new_n12789_));
  NOR3_X1    g11787(.A1(new_n12742_), .A2(new_n12743_), .A3(new_n12744_), .ZN(new_n12790_));
  AOI21_X1   g11788(.A1(new_n12733_), .A2(new_n12739_), .B(new_n12740_), .ZN(new_n12791_));
  NOR3_X1    g11789(.A1(new_n12786_), .A2(new_n12785_), .A3(new_n12787_), .ZN(new_n12792_));
  AOI21_X1   g11790(.A1(new_n12783_), .A2(new_n12776_), .B(new_n12746_), .ZN(new_n12793_));
  OAI22_X1   g11791(.A1(new_n12790_), .A2(new_n12791_), .B1(new_n12792_), .B2(new_n12793_), .ZN(new_n12794_));
  NAND3_X1   g11792(.A1(new_n12794_), .A2(new_n12789_), .A3(new_n12699_), .ZN(new_n12795_));
  NAND2_X1   g11793(.A1(new_n12463_), .A2(new_n12467_), .ZN(new_n12796_));
  INV_X1     g11794(.I(new_n12610_), .ZN(new_n12797_));
  NAND2_X1   g11795(.A1(new_n12797_), .A2(new_n12640_), .ZN(new_n12798_));
  NOR3_X1    g11796(.A1(new_n12798_), .A2(new_n12452_), .A3(new_n12612_), .ZN(new_n12799_));
  AOI21_X1   g11797(.A1(new_n12694_), .A2(new_n12695_), .B(new_n12693_), .ZN(new_n12800_));
  NOR3_X1    g11798(.A1(new_n12639_), .A2(new_n12682_), .A3(new_n12677_), .ZN(new_n12801_));
  OAI21_X1   g11799(.A1(new_n12800_), .A2(new_n12801_), .B(new_n12799_), .ZN(new_n12802_));
  NOR3_X1    g11800(.A1(new_n12800_), .A2(new_n12801_), .A3(new_n12799_), .ZN(new_n12803_));
  AOI21_X1   g11801(.A1(new_n12796_), .A2(new_n12802_), .B(new_n12803_), .ZN(new_n12804_));
  NOR4_X1    g11802(.A1(new_n12790_), .A2(new_n12791_), .A3(new_n12792_), .A4(new_n12793_), .ZN(new_n12805_));
  AOI22_X1   g11803(.A1(new_n12745_), .A2(new_n12741_), .B1(new_n12788_), .B2(new_n12784_), .ZN(new_n12806_));
  OAI21_X1   g11804(.A1(new_n12805_), .A2(new_n12806_), .B(new_n12804_), .ZN(new_n12807_));
  NAND4_X1   g11805(.A1(new_n12262_), .A2(new_n12252_), .A3(new_n12807_), .A4(new_n12795_), .ZN(new_n12808_));
  AOI22_X1   g11806(.A1(new_n12262_), .A2(new_n12252_), .B1(new_n12807_), .B2(new_n12795_), .ZN(new_n12809_));
  AOI21_X1   g11807(.A1(new_n12802_), .A2(new_n12698_), .B(new_n12796_), .ZN(new_n12810_));
  NOR3_X1    g11808(.A1(new_n12468_), .A2(new_n12697_), .A3(new_n12803_), .ZN(new_n12811_));
  NOR2_X1    g11809(.A1(new_n12811_), .A2(new_n12810_), .ZN(new_n12812_));
  NAND3_X1   g11810(.A1(new_n12259_), .A2(new_n12250_), .A3(new_n12241_), .ZN(new_n12813_));
  OAI21_X1   g11811(.A1(new_n12249_), .A2(new_n12260_), .B(new_n12255_), .ZN(new_n12814_));
  NOR2_X1    g11812(.A1(new_n12611_), .A2(new_n12613_), .ZN(new_n12815_));
  NOR2_X1    g11813(.A1(new_n12799_), .A2(new_n12815_), .ZN(new_n12816_));
  NOR2_X1    g11814(.A1(new_n12247_), .A2(new_n12245_), .ZN(new_n12817_));
  NOR2_X1    g11815(.A1(new_n12258_), .A2(new_n12817_), .ZN(new_n12818_));
  NAND2_X1   g11816(.A1(new_n12818_), .A2(new_n12816_), .ZN(new_n12819_));
  INV_X1     g11817(.I(new_n12819_), .ZN(new_n12820_));
  NAND3_X1   g11818(.A1(new_n12814_), .A2(new_n12813_), .A3(new_n12820_), .ZN(new_n12821_));
  AOI21_X1   g11819(.A1(new_n12814_), .A2(new_n12813_), .B(new_n12820_), .ZN(new_n12822_));
  AOI21_X1   g11820(.A1(new_n12812_), .A2(new_n12821_), .B(new_n12822_), .ZN(new_n12823_));
  OAI21_X1   g11821(.A1(new_n12809_), .A2(new_n12823_), .B(new_n12808_), .ZN(new_n12824_));
  OAI21_X1   g11822(.A1(new_n12804_), .A2(new_n12806_), .B(new_n12789_), .ZN(new_n12825_));
  NOR2_X1    g11823(.A1(new_n12742_), .A2(new_n12740_), .ZN(new_n12826_));
  NOR2_X1    g11824(.A1(new_n12727_), .A2(new_n12729_), .ZN(new_n12827_));
  NOR2_X1    g11825(.A1(new_n12827_), .A2(new_n12725_), .ZN(new_n12828_));
  NAND2_X1   g11826(.A1(new_n12712_), .A2(new_n12361_), .ZN(new_n12829_));
  OAI21_X1   g11827(.A1(new_n12829_), .A2(new_n12709_), .B(new_n12713_), .ZN(new_n12830_));
  NOR2_X1    g11828(.A1(new_n12828_), .A2(new_n12830_), .ZN(new_n12831_));
  NOR2_X1    g11829(.A1(new_n12700_), .A2(new_n12360_), .ZN(new_n12832_));
  AOI21_X1   g11830(.A1(new_n12832_), .A2(new_n12714_), .B(new_n12705_), .ZN(new_n12833_));
  NOR3_X1    g11831(.A1(new_n12833_), .A2(new_n12827_), .A3(new_n12725_), .ZN(new_n12834_));
  NOR2_X1    g11832(.A1(new_n12831_), .A2(new_n12834_), .ZN(new_n12835_));
  OAI21_X1   g11833(.A1(new_n12743_), .A2(new_n12826_), .B(new_n12835_), .ZN(new_n12836_));
  NAND2_X1   g11834(.A1(new_n12744_), .A2(new_n12733_), .ZN(new_n12837_));
  OAI21_X1   g11835(.A1(new_n12725_), .A2(new_n12827_), .B(new_n12833_), .ZN(new_n12838_));
  NAND2_X1   g11836(.A1(new_n12731_), .A2(new_n12721_), .ZN(new_n12839_));
  NAND3_X1   g11837(.A1(new_n12839_), .A2(new_n12830_), .A3(new_n12730_), .ZN(new_n12840_));
  NAND2_X1   g11838(.A1(new_n12838_), .A2(new_n12840_), .ZN(new_n12841_));
  NAND3_X1   g11839(.A1(new_n12837_), .A2(new_n12841_), .A3(new_n12739_), .ZN(new_n12842_));
  NAND2_X1   g11840(.A1(new_n12785_), .A2(new_n12776_), .ZN(new_n12843_));
  NAND2_X1   g11841(.A1(new_n12843_), .A2(new_n12783_), .ZN(new_n12844_));
  NOR2_X1    g11842(.A1(new_n12771_), .A2(new_n12766_), .ZN(new_n12845_));
  AOI21_X1   g11843(.A1(new_n12777_), .A2(new_n12761_), .B(new_n12752_), .ZN(new_n12846_));
  OAI21_X1   g11844(.A1(new_n12845_), .A2(new_n12769_), .B(new_n12846_), .ZN(new_n12847_));
  INV_X1     g11845(.I(new_n12847_), .ZN(new_n12848_));
  NOR3_X1    g11846(.A1(new_n12845_), .A2(new_n12846_), .A3(new_n12769_), .ZN(new_n12849_));
  NOR2_X1    g11847(.A1(new_n12848_), .A2(new_n12849_), .ZN(new_n12850_));
  NAND2_X1   g11848(.A1(new_n12844_), .A2(new_n12850_), .ZN(new_n12851_));
  INV_X1     g11849(.I(new_n12849_), .ZN(new_n12852_));
  NAND2_X1   g11850(.A1(new_n12852_), .A2(new_n12847_), .ZN(new_n12853_));
  NAND3_X1   g11851(.A1(new_n12853_), .A2(new_n12843_), .A3(new_n12783_), .ZN(new_n12854_));
  NAND4_X1   g11852(.A1(new_n12851_), .A2(new_n12836_), .A3(new_n12842_), .A4(new_n12854_), .ZN(new_n12855_));
  AOI21_X1   g11853(.A1(new_n12837_), .A2(new_n12739_), .B(new_n12841_), .ZN(new_n12856_));
  NOR3_X1    g11854(.A1(new_n12835_), .A2(new_n12826_), .A3(new_n12743_), .ZN(new_n12857_));
  AOI21_X1   g11855(.A1(new_n12843_), .A2(new_n12783_), .B(new_n12853_), .ZN(new_n12858_));
  NOR2_X1    g11856(.A1(new_n12786_), .A2(new_n12746_), .ZN(new_n12859_));
  NOR3_X1    g11857(.A1(new_n12850_), .A2(new_n12859_), .A3(new_n12787_), .ZN(new_n12860_));
  OAI22_X1   g11858(.A1(new_n12858_), .A2(new_n12860_), .B1(new_n12856_), .B2(new_n12857_), .ZN(new_n12861_));
  NAND3_X1   g11859(.A1(new_n12825_), .A2(new_n12855_), .A3(new_n12861_), .ZN(new_n12862_));
  AOI21_X1   g11860(.A1(new_n12699_), .A2(new_n12794_), .B(new_n12805_), .ZN(new_n12863_));
  NAND2_X1   g11861(.A1(new_n12855_), .A2(new_n12861_), .ZN(new_n12864_));
  NAND2_X1   g11862(.A1(new_n12864_), .A2(new_n12863_), .ZN(new_n12865_));
  OAI21_X1   g11863(.A1(new_n12254_), .A2(new_n12261_), .B(new_n12233_), .ZN(new_n12866_));
  NAND2_X1   g11864(.A1(new_n12214_), .A2(new_n12229_), .ZN(new_n12867_));
  NAND2_X1   g11865(.A1(new_n12867_), .A2(new_n12220_), .ZN(new_n12868_));
  AOI21_X1   g11866(.A1(new_n12201_), .A2(new_n12212_), .B(new_n12206_), .ZN(new_n12869_));
  NOR2_X1    g11867(.A1(new_n12175_), .A2(new_n12169_), .ZN(new_n12870_));
  AOI21_X1   g11868(.A1(new_n12870_), .A2(new_n12193_), .B(new_n12184_), .ZN(new_n12871_));
  XNOR2_X1   g11869(.A1(new_n12869_), .A2(new_n12871_), .ZN(new_n12872_));
  NAND2_X1   g11870(.A1(new_n12868_), .A2(new_n12872_), .ZN(new_n12873_));
  AOI21_X1   g11871(.A1(new_n12229_), .A2(new_n12214_), .B(new_n12231_), .ZN(new_n12874_));
  XOR2_X1    g11872(.A1(new_n12869_), .A2(new_n12871_), .Z(new_n12875_));
  NAND2_X1   g11873(.A1(new_n12874_), .A2(new_n12875_), .ZN(new_n12876_));
  NOR2_X1    g11874(.A1(new_n11979_), .A2(new_n11977_), .ZN(new_n12877_));
  NAND2_X1   g11875(.A1(new_n11952_), .A2(new_n11881_), .ZN(new_n12878_));
  NAND2_X1   g11876(.A1(new_n11848_), .A2(new_n11846_), .ZN(new_n12879_));
  OAI21_X1   g11877(.A1(new_n12879_), .A2(new_n11839_), .B(new_n11849_), .ZN(new_n12880_));
  AOI21_X1   g11878(.A1(new_n12878_), .A2(new_n11951_), .B(new_n12880_), .ZN(new_n12881_));
  NOR2_X1    g11879(.A1(new_n11949_), .A2(new_n11880_), .ZN(new_n12882_));
  NOR2_X1    g11880(.A1(new_n11832_), .A2(new_n11824_), .ZN(new_n12883_));
  AOI21_X1   g11881(.A1(new_n12883_), .A2(new_n11838_), .B(new_n11837_), .ZN(new_n12884_));
  NOR3_X1    g11882(.A1(new_n12884_), .A2(new_n12882_), .A3(new_n11941_), .ZN(new_n12885_));
  NOR2_X1    g11883(.A1(new_n12881_), .A2(new_n12885_), .ZN(new_n12886_));
  OAI21_X1   g11884(.A1(new_n12877_), .A2(new_n11980_), .B(new_n12886_), .ZN(new_n12887_));
  NAND2_X1   g11885(.A1(new_n11954_), .A2(new_n11989_), .ZN(new_n12888_));
  OAI21_X1   g11886(.A1(new_n11941_), .A2(new_n12882_), .B(new_n12884_), .ZN(new_n12889_));
  NAND3_X1   g11887(.A1(new_n12878_), .A2(new_n12880_), .A3(new_n11951_), .ZN(new_n12890_));
  NAND2_X1   g11888(.A1(new_n12889_), .A2(new_n12890_), .ZN(new_n12891_));
  NAND3_X1   g11889(.A1(new_n12888_), .A2(new_n12891_), .A3(new_n11960_), .ZN(new_n12892_));
  NAND4_X1   g11890(.A1(new_n12873_), .A2(new_n12876_), .A3(new_n12887_), .A4(new_n12892_), .ZN(new_n12893_));
  NOR2_X1    g11891(.A1(new_n12874_), .A2(new_n12875_), .ZN(new_n12894_));
  NOR2_X1    g11892(.A1(new_n12868_), .A2(new_n12872_), .ZN(new_n12895_));
  AOI21_X1   g11893(.A1(new_n12888_), .A2(new_n11960_), .B(new_n12891_), .ZN(new_n12896_));
  NOR3_X1    g11894(.A1(new_n12877_), .A2(new_n12886_), .A3(new_n11980_), .ZN(new_n12897_));
  OAI22_X1   g11895(.A1(new_n12895_), .A2(new_n12894_), .B1(new_n12896_), .B2(new_n12897_), .ZN(new_n12898_));
  NAND3_X1   g11896(.A1(new_n12866_), .A2(new_n12898_), .A3(new_n12893_), .ZN(new_n12899_));
  AOI21_X1   g11897(.A1(new_n12238_), .A2(new_n12251_), .B(new_n12253_), .ZN(new_n12900_));
  NAND2_X1   g11898(.A1(new_n12898_), .A2(new_n12893_), .ZN(new_n12901_));
  NAND2_X1   g11899(.A1(new_n12901_), .A2(new_n12900_), .ZN(new_n12902_));
  NAND4_X1   g11900(.A1(new_n12902_), .A2(new_n12865_), .A3(new_n12862_), .A4(new_n12899_), .ZN(new_n12903_));
  NOR2_X1    g11901(.A1(new_n12864_), .A2(new_n12863_), .ZN(new_n12904_));
  AOI21_X1   g11902(.A1(new_n12855_), .A2(new_n12861_), .B(new_n12825_), .ZN(new_n12905_));
  INV_X1     g11903(.I(new_n12899_), .ZN(new_n12906_));
  AOI21_X1   g11904(.A1(new_n12898_), .A2(new_n12893_), .B(new_n12866_), .ZN(new_n12907_));
  OAI22_X1   g11905(.A1(new_n12906_), .A2(new_n12907_), .B1(new_n12904_), .B2(new_n12905_), .ZN(new_n12908_));
  NAND3_X1   g11906(.A1(new_n12908_), .A2(new_n12903_), .A3(new_n12824_), .ZN(new_n12909_));
  NOR3_X1    g11907(.A1(new_n12253_), .A2(new_n12254_), .A3(new_n12261_), .ZN(new_n12910_));
  AOI21_X1   g11908(.A1(new_n12238_), .A2(new_n12233_), .B(new_n12251_), .ZN(new_n12911_));
  NOR3_X1    g11909(.A1(new_n12805_), .A2(new_n12806_), .A3(new_n12804_), .ZN(new_n12912_));
  AOI21_X1   g11910(.A1(new_n12794_), .A2(new_n12789_), .B(new_n12699_), .ZN(new_n12913_));
  NOR4_X1    g11911(.A1(new_n12910_), .A2(new_n12911_), .A3(new_n12912_), .A4(new_n12913_), .ZN(new_n12914_));
  OAI22_X1   g11912(.A1(new_n12910_), .A2(new_n12911_), .B1(new_n12912_), .B2(new_n12913_), .ZN(new_n12915_));
  INV_X1     g11913(.I(new_n12812_), .ZN(new_n12916_));
  NOR3_X1    g11914(.A1(new_n12255_), .A2(new_n12260_), .A3(new_n12249_), .ZN(new_n12917_));
  AOI21_X1   g11915(.A1(new_n12259_), .A2(new_n12250_), .B(new_n12241_), .ZN(new_n12918_));
  NOR3_X1    g11916(.A1(new_n12917_), .A2(new_n12918_), .A3(new_n12819_), .ZN(new_n12919_));
  OAI21_X1   g11917(.A1(new_n12917_), .A2(new_n12918_), .B(new_n12819_), .ZN(new_n12920_));
  OAI21_X1   g11918(.A1(new_n12916_), .A2(new_n12919_), .B(new_n12920_), .ZN(new_n12921_));
  AOI21_X1   g11919(.A1(new_n12915_), .A2(new_n12921_), .B(new_n12914_), .ZN(new_n12922_));
  NOR4_X1    g11920(.A1(new_n12906_), .A2(new_n12904_), .A3(new_n12905_), .A4(new_n12907_), .ZN(new_n12923_));
  AOI22_X1   g11921(.A1(new_n12902_), .A2(new_n12899_), .B1(new_n12865_), .B2(new_n12862_), .ZN(new_n12924_));
  OAI21_X1   g11922(.A1(new_n12924_), .A2(new_n12923_), .B(new_n12922_), .ZN(new_n12925_));
  NAND2_X1   g11923(.A1(new_n12925_), .A2(new_n12909_), .ZN(new_n12926_));
  NAND3_X1   g11924(.A1(new_n12916_), .A2(new_n12821_), .A3(new_n12920_), .ZN(new_n12927_));
  OAI21_X1   g11925(.A1(new_n12822_), .A2(new_n12919_), .B(new_n12812_), .ZN(new_n12928_));
  AND2_X2    g11926(.A1(new_n12927_), .A2(new_n12928_), .Z(new_n12929_));
  NOR2_X1    g11927(.A1(new_n11716_), .A2(new_n11714_), .ZN(new_n12930_));
  NOR2_X1    g11928(.A1(new_n11748_), .A2(new_n12930_), .ZN(new_n12931_));
  NOR2_X1    g11929(.A1(new_n12818_), .A2(new_n12816_), .ZN(new_n12932_));
  NOR2_X1    g11930(.A1(new_n12820_), .A2(new_n12932_), .ZN(new_n12933_));
  NAND2_X1   g11931(.A1(new_n12933_), .A2(new_n12931_), .ZN(new_n12934_));
  OAI21_X1   g11932(.A1(new_n11752_), .A2(new_n11727_), .B(new_n11712_), .ZN(new_n12935_));
  NAND3_X1   g11933(.A1(new_n11747_), .A2(new_n11751_), .A3(new_n11728_), .ZN(new_n12936_));
  AOI21_X1   g11934(.A1(new_n12936_), .A2(new_n12935_), .B(new_n12934_), .ZN(new_n12937_));
  NAND3_X1   g11935(.A1(new_n12936_), .A2(new_n12934_), .A3(new_n12935_), .ZN(new_n12938_));
  OAI21_X1   g11936(.A1(new_n12929_), .A2(new_n12937_), .B(new_n12938_), .ZN(new_n12939_));
  NOR3_X1    g11937(.A1(new_n12914_), .A2(new_n12809_), .A3(new_n12823_), .ZN(new_n12940_));
  AOI21_X1   g11938(.A1(new_n12915_), .A2(new_n12808_), .B(new_n12921_), .ZN(new_n12941_));
  NOR3_X1    g11939(.A1(new_n11741_), .A2(new_n11759_), .A3(new_n11753_), .ZN(new_n12942_));
  AOI21_X1   g11940(.A1(new_n11742_), .A2(new_n11758_), .B(new_n11729_), .ZN(new_n12943_));
  NOR4_X1    g11941(.A1(new_n12940_), .A2(new_n12941_), .A3(new_n12942_), .A4(new_n12943_), .ZN(new_n12944_));
  OAI22_X1   g11942(.A1(new_n12940_), .A2(new_n12941_), .B1(new_n12942_), .B2(new_n12943_), .ZN(new_n12945_));
  AOI21_X1   g11943(.A1(new_n12939_), .A2(new_n12945_), .B(new_n12944_), .ZN(new_n12946_));
  NOR2_X1    g11944(.A1(new_n12926_), .A2(new_n12946_), .ZN(new_n12947_));
  NAND2_X1   g11945(.A1(new_n12926_), .A2(new_n12946_), .ZN(new_n12948_));
  AOI21_X1   g11946(.A1(new_n11766_), .A2(new_n12948_), .B(new_n12947_), .ZN(new_n12949_));
  NOR2_X1    g11947(.A1(new_n11761_), .A2(new_n11126_), .ZN(new_n12950_));
  NOR2_X1    g11948(.A1(new_n12950_), .A2(new_n11744_), .ZN(new_n12951_));
  INV_X1     g11949(.I(new_n11694_), .ZN(new_n12952_));
  NOR2_X1    g11950(.A1(new_n11693_), .A2(new_n12952_), .ZN(new_n12953_));
  INV_X1     g11951(.I(new_n12953_), .ZN(new_n12954_));
  NAND2_X1   g11952(.A1(new_n11693_), .A2(new_n12952_), .ZN(new_n12955_));
  NAND2_X1   g11953(.A1(new_n11692_), .A2(new_n12955_), .ZN(new_n12956_));
  NAND2_X1   g11954(.A1(new_n11681_), .A2(new_n11683_), .ZN(new_n12957_));
  NAND2_X1   g11955(.A1(new_n11684_), .A2(new_n11686_), .ZN(new_n12958_));
  NAND2_X1   g11956(.A1(new_n11680_), .A2(new_n12958_), .ZN(new_n12959_));
  AOI22_X1   g11957(.A1(new_n12959_), .A2(new_n12957_), .B1(new_n12954_), .B2(new_n12956_), .ZN(new_n12960_));
  AOI21_X1   g11958(.A1(new_n11738_), .A2(new_n11739_), .B(new_n11736_), .ZN(new_n12961_));
  NAND2_X1   g11959(.A1(new_n11700_), .A2(new_n12961_), .ZN(new_n12962_));
  AOI22_X1   g11960(.A1(new_n11679_), .A2(new_n11622_), .B1(new_n11686_), .B2(new_n11684_), .ZN(new_n12963_));
  NAND2_X1   g11961(.A1(new_n12963_), .A2(new_n12957_), .ZN(new_n12964_));
  NOR2_X1    g11962(.A1(new_n12956_), .A2(new_n12953_), .ZN(new_n12965_));
  NOR2_X1    g11963(.A1(new_n11698_), .A2(new_n11692_), .ZN(new_n12966_));
  NOR2_X1    g11964(.A1(new_n12965_), .A2(new_n12966_), .ZN(new_n12967_));
  NOR2_X1    g11965(.A1(new_n11680_), .A2(new_n11690_), .ZN(new_n12968_));
  INV_X1     g11966(.I(new_n12968_), .ZN(new_n12969_));
  NAND3_X1   g11967(.A1(new_n12967_), .A2(new_n12964_), .A3(new_n12969_), .ZN(new_n12970_));
  NAND2_X1   g11968(.A1(new_n12962_), .A2(new_n12970_), .ZN(new_n12971_));
  NOR2_X1    g11969(.A1(new_n11701_), .A2(new_n11702_), .ZN(new_n12972_));
  NOR2_X1    g11970(.A1(new_n11703_), .A2(new_n11704_), .ZN(new_n12973_));
  AOI21_X1   g11971(.A1(new_n12972_), .A2(new_n12973_), .B(new_n11678_), .ZN(new_n12974_));
  INV_X1     g11972(.I(new_n12964_), .ZN(new_n12975_));
  NOR4_X1    g11973(.A1(new_n12975_), .A2(new_n12965_), .A3(new_n12966_), .A4(new_n12968_), .ZN(new_n12976_));
  NAND4_X1   g11974(.A1(new_n12959_), .A2(new_n12956_), .A3(new_n12954_), .A4(new_n12957_), .ZN(new_n12977_));
  OAI21_X1   g11975(.A1(new_n12974_), .A2(new_n12976_), .B(new_n12977_), .ZN(new_n12978_));
  INV_X1     g11976(.I(new_n12977_), .ZN(new_n12979_));
  NOR2_X1    g11977(.A1(new_n12979_), .A2(new_n12960_), .ZN(new_n12980_));
  OAI22_X1   g11978(.A1(new_n12978_), .A2(new_n12960_), .B1(new_n12971_), .B2(new_n12980_), .ZN(new_n12981_));
  AOI21_X1   g11979(.A1(new_n11119_), .A2(new_n10784_), .B(new_n11092_), .ZN(new_n12982_));
  NOR2_X1    g11980(.A1(new_n11119_), .A2(new_n10784_), .ZN(new_n12983_));
  INV_X1     g11981(.I(new_n11096_), .ZN(new_n12984_));
  NAND2_X1   g11982(.A1(new_n12984_), .A2(new_n11094_), .ZN(new_n12985_));
  INV_X1     g11983(.I(new_n12985_), .ZN(new_n12986_));
  NOR2_X1    g11984(.A1(new_n12984_), .A2(new_n11094_), .ZN(new_n12987_));
  NOR2_X1    g11985(.A1(new_n11093_), .A2(new_n12987_), .ZN(new_n12988_));
  NOR2_X1    g11986(.A1(new_n12988_), .A2(new_n12986_), .ZN(new_n12989_));
  NOR2_X1    g11987(.A1(new_n10778_), .A2(new_n10780_), .ZN(new_n12990_));
  NOR2_X1    g11988(.A1(new_n12990_), .A2(new_n10736_), .ZN(new_n12991_));
  XNOR2_X1   g11989(.A1(new_n12989_), .A2(new_n12991_), .ZN(new_n12992_));
  OAI21_X1   g11990(.A1(new_n12982_), .A2(new_n12983_), .B(new_n12992_), .ZN(new_n12993_));
  OAI21_X1   g11991(.A1(new_n10785_), .A2(new_n11102_), .B(new_n11118_), .ZN(new_n12994_));
  NAND2_X1   g11992(.A1(new_n10785_), .A2(new_n11102_), .ZN(new_n12995_));
  XOR2_X1    g11993(.A1(new_n12989_), .A2(new_n12991_), .Z(new_n12996_));
  NAND3_X1   g11994(.A1(new_n12996_), .A2(new_n12994_), .A3(new_n12995_), .ZN(new_n12997_));
  NAND3_X1   g11995(.A1(new_n12981_), .A2(new_n12993_), .A3(new_n12997_), .ZN(new_n12998_));
  INV_X1     g11996(.I(new_n12960_), .ZN(new_n12999_));
  INV_X1     g11997(.I(new_n12971_), .ZN(new_n13000_));
  AOI21_X1   g11998(.A1(new_n12962_), .A2(new_n12970_), .B(new_n12979_), .ZN(new_n13001_));
  INV_X1     g11999(.I(new_n12980_), .ZN(new_n13002_));
  AOI22_X1   g12000(.A1(new_n13000_), .A2(new_n13002_), .B1(new_n13001_), .B2(new_n12999_), .ZN(new_n13003_));
  NAND2_X1   g12001(.A1(new_n12993_), .A2(new_n12997_), .ZN(new_n13004_));
  NAND2_X1   g12002(.A1(new_n13003_), .A2(new_n13004_), .ZN(new_n13005_));
  NAND2_X1   g12003(.A1(new_n13005_), .A2(new_n12998_), .ZN(new_n13006_));
  NAND2_X1   g12004(.A1(new_n13006_), .A2(new_n12951_), .ZN(new_n13007_));
  NAND2_X1   g12005(.A1(new_n11764_), .A2(new_n11125_), .ZN(new_n13008_));
  NAND2_X1   g12006(.A1(new_n13008_), .A2(new_n11763_), .ZN(new_n13009_));
  NAND3_X1   g12007(.A1(new_n13009_), .A2(new_n12998_), .A3(new_n13005_), .ZN(new_n13010_));
  NAND2_X1   g12008(.A1(new_n12908_), .A2(new_n12824_), .ZN(new_n13011_));
  NOR2_X1    g12009(.A1(new_n12845_), .A2(new_n12769_), .ZN(new_n13012_));
  INV_X1     g12010(.I(new_n13012_), .ZN(new_n13013_));
  INV_X1     g12011(.I(new_n12846_), .ZN(new_n13014_));
  NOR2_X1    g12012(.A1(new_n13013_), .A2(new_n13014_), .ZN(new_n13015_));
  INV_X1     g12013(.I(new_n13015_), .ZN(new_n13016_));
  NAND2_X1   g12014(.A1(new_n13013_), .A2(new_n13014_), .ZN(new_n13017_));
  NAND2_X1   g12015(.A1(new_n12844_), .A2(new_n13017_), .ZN(new_n13018_));
  INV_X1     g12016(.I(new_n12828_), .ZN(new_n13019_));
  NOR2_X1    g12017(.A1(new_n13019_), .A2(new_n12830_), .ZN(new_n13020_));
  INV_X1     g12018(.I(new_n13020_), .ZN(new_n13021_));
  NAND2_X1   g12019(.A1(new_n12837_), .A2(new_n12739_), .ZN(new_n13022_));
  NAND2_X1   g12020(.A1(new_n13019_), .A2(new_n12830_), .ZN(new_n13023_));
  NAND2_X1   g12021(.A1(new_n13022_), .A2(new_n13023_), .ZN(new_n13024_));
  AOI22_X1   g12022(.A1(new_n13024_), .A2(new_n13021_), .B1(new_n13018_), .B2(new_n13016_), .ZN(new_n13025_));
  NAND2_X1   g12023(.A1(new_n12863_), .A2(new_n12855_), .ZN(new_n13026_));
  NAND3_X1   g12024(.A1(new_n13022_), .A2(new_n13021_), .A3(new_n13023_), .ZN(new_n13027_));
  NAND3_X1   g12025(.A1(new_n12844_), .A2(new_n13016_), .A3(new_n13017_), .ZN(new_n13028_));
  NAND3_X1   g12026(.A1(new_n12850_), .A2(new_n12843_), .A3(new_n12783_), .ZN(new_n13029_));
  NOR2_X1    g12027(.A1(new_n12826_), .A2(new_n12743_), .ZN(new_n13030_));
  NAND2_X1   g12028(.A1(new_n13030_), .A2(new_n12835_), .ZN(new_n13031_));
  NAND4_X1   g12029(.A1(new_n13027_), .A2(new_n13028_), .A3(new_n13031_), .A4(new_n13029_), .ZN(new_n13032_));
  NAND2_X1   g12030(.A1(new_n13026_), .A2(new_n13032_), .ZN(new_n13033_));
  NOR4_X1    g12031(.A1(new_n12860_), .A2(new_n12857_), .A3(new_n12856_), .A4(new_n12858_), .ZN(new_n13034_));
  NOR2_X1    g12032(.A1(new_n13034_), .A2(new_n12825_), .ZN(new_n13035_));
  INV_X1     g12033(.I(new_n13032_), .ZN(new_n13036_));
  NAND4_X1   g12034(.A1(new_n13024_), .A2(new_n13018_), .A3(new_n13016_), .A4(new_n13021_), .ZN(new_n13037_));
  OAI21_X1   g12035(.A1(new_n13035_), .A2(new_n13036_), .B(new_n13037_), .ZN(new_n13038_));
  INV_X1     g12036(.I(new_n13037_), .ZN(new_n13039_));
  NOR2_X1    g12037(.A1(new_n13039_), .A2(new_n13025_), .ZN(new_n13040_));
  OAI22_X1   g12038(.A1(new_n13038_), .A2(new_n13025_), .B1(new_n13033_), .B2(new_n13040_), .ZN(new_n13041_));
  NAND2_X1   g12039(.A1(new_n12900_), .A2(new_n12893_), .ZN(new_n13042_));
  INV_X1     g12040(.I(new_n12869_), .ZN(new_n13043_));
  INV_X1     g12041(.I(new_n12871_), .ZN(new_n13044_));
  NOR2_X1    g12042(.A1(new_n13043_), .A2(new_n13044_), .ZN(new_n13045_));
  INV_X1     g12043(.I(new_n13045_), .ZN(new_n13046_));
  NOR2_X1    g12044(.A1(new_n12869_), .A2(new_n12871_), .ZN(new_n13047_));
  OAI21_X1   g12045(.A1(new_n12874_), .A2(new_n13047_), .B(new_n13046_), .ZN(new_n13048_));
  NOR2_X1    g12046(.A1(new_n12877_), .A2(new_n11980_), .ZN(new_n13049_));
  NOR2_X1    g12047(.A1(new_n12882_), .A2(new_n11941_), .ZN(new_n13050_));
  NAND2_X1   g12048(.A1(new_n13050_), .A2(new_n12884_), .ZN(new_n13051_));
  NOR2_X1    g12049(.A1(new_n13050_), .A2(new_n12884_), .ZN(new_n13052_));
  OAI21_X1   g12050(.A1(new_n13049_), .A2(new_n13052_), .B(new_n13051_), .ZN(new_n13053_));
  XOR2_X1    g12051(.A1(new_n13053_), .A2(new_n13048_), .Z(new_n13054_));
  AOI21_X1   g12052(.A1(new_n12898_), .A2(new_n13042_), .B(new_n13054_), .ZN(new_n13055_));
  INV_X1     g12053(.I(new_n12898_), .ZN(new_n13056_));
  NOR4_X1    g12054(.A1(new_n12895_), .A2(new_n12894_), .A3(new_n12896_), .A4(new_n12897_), .ZN(new_n13057_));
  NOR2_X1    g12055(.A1(new_n12866_), .A2(new_n13057_), .ZN(new_n13058_));
  INV_X1     g12056(.I(new_n13047_), .ZN(new_n13059_));
  AOI21_X1   g12057(.A1(new_n12868_), .A2(new_n13059_), .B(new_n13045_), .ZN(new_n13060_));
  XOR2_X1    g12058(.A1(new_n13053_), .A2(new_n13060_), .Z(new_n13061_));
  NOR3_X1    g12059(.A1(new_n13061_), .A2(new_n13058_), .A3(new_n13056_), .ZN(new_n13062_));
  NOR2_X1    g12060(.A1(new_n13055_), .A2(new_n13062_), .ZN(new_n13063_));
  NAND2_X1   g12061(.A1(new_n13063_), .A2(new_n13041_), .ZN(new_n13064_));
  INV_X1     g12062(.I(new_n13025_), .ZN(new_n13065_));
  NOR2_X1    g12063(.A1(new_n13035_), .A2(new_n13036_), .ZN(new_n13066_));
  AOI21_X1   g12064(.A1(new_n13026_), .A2(new_n13032_), .B(new_n13039_), .ZN(new_n13067_));
  NAND2_X1   g12065(.A1(new_n13065_), .A2(new_n13037_), .ZN(new_n13068_));
  AOI22_X1   g12066(.A1(new_n13065_), .A2(new_n13067_), .B1(new_n13066_), .B2(new_n13068_), .ZN(new_n13069_));
  OAI21_X1   g12067(.A1(new_n13056_), .A2(new_n13058_), .B(new_n13061_), .ZN(new_n13070_));
  NAND3_X1   g12068(.A1(new_n13054_), .A2(new_n12898_), .A3(new_n13042_), .ZN(new_n13071_));
  NAND2_X1   g12069(.A1(new_n13070_), .A2(new_n13071_), .ZN(new_n13072_));
  NAND2_X1   g12070(.A1(new_n13072_), .A2(new_n13069_), .ZN(new_n13073_));
  NAND4_X1   g12071(.A1(new_n13064_), .A2(new_n13073_), .A3(new_n12903_), .A4(new_n13011_), .ZN(new_n13074_));
  OAI21_X1   g12072(.A1(new_n12924_), .A2(new_n12922_), .B(new_n12903_), .ZN(new_n13075_));
  NOR2_X1    g12073(.A1(new_n13072_), .A2(new_n13069_), .ZN(new_n13076_));
  NOR2_X1    g12074(.A1(new_n13063_), .A2(new_n13041_), .ZN(new_n13077_));
  OAI21_X1   g12075(.A1(new_n13077_), .A2(new_n13076_), .B(new_n13075_), .ZN(new_n13078_));
  NAND2_X1   g12076(.A1(new_n13074_), .A2(new_n13078_), .ZN(new_n13079_));
  NAND3_X1   g12077(.A1(new_n13079_), .A2(new_n13007_), .A3(new_n13010_), .ZN(new_n13080_));
  AOI21_X1   g12078(.A1(new_n13007_), .A2(new_n13010_), .B(new_n13079_), .ZN(new_n13081_));
  OAI21_X1   g12079(.A1(new_n13081_), .A2(new_n12949_), .B(new_n13080_), .ZN(new_n13082_));
  NAND3_X1   g12080(.A1(new_n13064_), .A2(new_n12903_), .A3(new_n13011_), .ZN(new_n13083_));
  AND2_X2    g12081(.A1(new_n13053_), .A2(new_n13048_), .Z(new_n13084_));
  NAND2_X1   g12082(.A1(new_n13042_), .A2(new_n12898_), .ZN(new_n13085_));
  NOR2_X1    g12083(.A1(new_n13053_), .A2(new_n13048_), .ZN(new_n13086_));
  INV_X1     g12084(.I(new_n13086_), .ZN(new_n13087_));
  NAND2_X1   g12085(.A1(new_n13085_), .A2(new_n13087_), .ZN(new_n13088_));
  NOR2_X1    g12086(.A1(new_n13088_), .A2(new_n13084_), .ZN(new_n13089_));
  NOR2_X1    g12087(.A1(new_n13085_), .A2(new_n13054_), .ZN(new_n13090_));
  NOR3_X1    g12088(.A1(new_n13089_), .A2(new_n13041_), .A3(new_n13090_), .ZN(new_n13091_));
  INV_X1     g12089(.I(new_n13091_), .ZN(new_n13092_));
  NOR2_X1    g12090(.A1(new_n13067_), .A2(new_n13025_), .ZN(new_n13093_));
  AOI21_X1   g12091(.A1(new_n13085_), .A2(new_n13087_), .B(new_n13084_), .ZN(new_n13094_));
  XOR2_X1    g12092(.A1(new_n13094_), .A2(new_n13093_), .Z(new_n13095_));
  AOI21_X1   g12093(.A1(new_n13083_), .A2(new_n13092_), .B(new_n13095_), .ZN(new_n13096_));
  NOR2_X1    g12094(.A1(new_n13076_), .A2(new_n13075_), .ZN(new_n13097_));
  XNOR2_X1   g12095(.A1(new_n13094_), .A2(new_n13093_), .ZN(new_n13098_));
  NOR3_X1    g12096(.A1(new_n13098_), .A2(new_n13097_), .A3(new_n13091_), .ZN(new_n13099_));
  NAND3_X1   g12097(.A1(new_n13008_), .A2(new_n12998_), .A3(new_n11763_), .ZN(new_n13100_));
  NOR2_X1    g12098(.A1(new_n12989_), .A2(new_n12991_), .ZN(new_n13101_));
  NAND2_X1   g12099(.A1(new_n12994_), .A2(new_n12995_), .ZN(new_n13102_));
  NAND2_X1   g12100(.A1(new_n12989_), .A2(new_n12991_), .ZN(new_n13103_));
  NAND2_X1   g12101(.A1(new_n13102_), .A2(new_n13103_), .ZN(new_n13104_));
  NOR2_X1    g12102(.A1(new_n13104_), .A2(new_n13101_), .ZN(new_n13105_));
  NOR2_X1    g12103(.A1(new_n13102_), .A2(new_n12996_), .ZN(new_n13106_));
  NOR3_X1    g12104(.A1(new_n13105_), .A2(new_n12981_), .A3(new_n13106_), .ZN(new_n13107_));
  INV_X1     g12105(.I(new_n13107_), .ZN(new_n13108_));
  NOR2_X1    g12106(.A1(new_n13001_), .A2(new_n12960_), .ZN(new_n13109_));
  AOI21_X1   g12107(.A1(new_n13102_), .A2(new_n13103_), .B(new_n13101_), .ZN(new_n13110_));
  XOR2_X1    g12108(.A1(new_n13110_), .A2(new_n13109_), .Z(new_n13111_));
  AOI21_X1   g12109(.A1(new_n13100_), .A2(new_n13108_), .B(new_n13111_), .ZN(new_n13112_));
  NOR2_X1    g12110(.A1(new_n13003_), .A2(new_n13004_), .ZN(new_n13113_));
  NOR3_X1    g12111(.A1(new_n13113_), .A2(new_n12950_), .A3(new_n11744_), .ZN(new_n13114_));
  XNOR2_X1   g12112(.A1(new_n13110_), .A2(new_n13109_), .ZN(new_n13115_));
  NOR3_X1    g12113(.A1(new_n13114_), .A2(new_n13115_), .A3(new_n13107_), .ZN(new_n13116_));
  NOR4_X1    g12114(.A1(new_n13116_), .A2(new_n13112_), .A3(new_n13096_), .A4(new_n13099_), .ZN(new_n13117_));
  OAI21_X1   g12115(.A1(new_n13097_), .A2(new_n13091_), .B(new_n13098_), .ZN(new_n13118_));
  NAND3_X1   g12116(.A1(new_n13083_), .A2(new_n13092_), .A3(new_n13095_), .ZN(new_n13119_));
  OAI21_X1   g12117(.A1(new_n13114_), .A2(new_n13107_), .B(new_n13115_), .ZN(new_n13120_));
  NAND3_X1   g12118(.A1(new_n13100_), .A2(new_n13108_), .A3(new_n13111_), .ZN(new_n13121_));
  AOI22_X1   g12119(.A1(new_n13120_), .A2(new_n13121_), .B1(new_n13118_), .B2(new_n13119_), .ZN(new_n13122_));
  NOR2_X1    g12120(.A1(new_n13117_), .A2(new_n13122_), .ZN(new_n13123_));
  NAND2_X1   g12121(.A1(new_n13123_), .A2(new_n13082_), .ZN(new_n13124_));
  NAND3_X1   g12122(.A1(new_n11764_), .A2(new_n11763_), .A3(new_n11125_), .ZN(new_n13125_));
  OAI21_X1   g12123(.A1(new_n11744_), .A2(new_n11761_), .B(new_n11126_), .ZN(new_n13126_));
  NAND2_X1   g12124(.A1(new_n13126_), .A2(new_n13125_), .ZN(new_n13127_));
  NOR3_X1    g12125(.A1(new_n12924_), .A2(new_n12923_), .A3(new_n12922_), .ZN(new_n13128_));
  AOI21_X1   g12126(.A1(new_n12908_), .A2(new_n12903_), .B(new_n12824_), .ZN(new_n13129_));
  NOR2_X1    g12127(.A1(new_n13128_), .A2(new_n13129_), .ZN(new_n13130_));
  NAND2_X1   g12128(.A1(new_n12927_), .A2(new_n12928_), .ZN(new_n13131_));
  INV_X1     g12129(.I(new_n12934_), .ZN(new_n13132_));
  INV_X1     g12130(.I(new_n12935_), .ZN(new_n13133_));
  NOR3_X1    g12131(.A1(new_n11752_), .A2(new_n11727_), .A3(new_n11712_), .ZN(new_n13134_));
  OAI21_X1   g12132(.A1(new_n13133_), .A2(new_n13134_), .B(new_n13132_), .ZN(new_n13135_));
  NOR3_X1    g12133(.A1(new_n13133_), .A2(new_n13132_), .A3(new_n13134_), .ZN(new_n13136_));
  AOI21_X1   g12134(.A1(new_n13131_), .A2(new_n13135_), .B(new_n13136_), .ZN(new_n13137_));
  NAND3_X1   g12135(.A1(new_n12915_), .A2(new_n12808_), .A3(new_n12921_), .ZN(new_n13138_));
  OAI21_X1   g12136(.A1(new_n12914_), .A2(new_n12809_), .B(new_n12823_), .ZN(new_n13139_));
  NAND3_X1   g12137(.A1(new_n11742_), .A2(new_n11758_), .A3(new_n11729_), .ZN(new_n13140_));
  OAI21_X1   g12138(.A1(new_n11741_), .A2(new_n11759_), .B(new_n11753_), .ZN(new_n13141_));
  NAND4_X1   g12139(.A1(new_n13139_), .A2(new_n13138_), .A3(new_n13141_), .A4(new_n13140_), .ZN(new_n13142_));
  AOI22_X1   g12140(.A1(new_n13139_), .A2(new_n13138_), .B1(new_n13141_), .B2(new_n13140_), .ZN(new_n13143_));
  OAI21_X1   g12141(.A1(new_n13143_), .A2(new_n13137_), .B(new_n13142_), .ZN(new_n13144_));
  NAND2_X1   g12142(.A1(new_n13130_), .A2(new_n13144_), .ZN(new_n13145_));
  NOR2_X1    g12143(.A1(new_n13130_), .A2(new_n13144_), .ZN(new_n13146_));
  OAI21_X1   g12144(.A1(new_n13127_), .A2(new_n13146_), .B(new_n13145_), .ZN(new_n13147_));
  AOI21_X1   g12145(.A1(new_n12998_), .A2(new_n13005_), .B(new_n13009_), .ZN(new_n13148_));
  NOR2_X1    g12146(.A1(new_n13006_), .A2(new_n12951_), .ZN(new_n13149_));
  NOR3_X1    g12147(.A1(new_n13077_), .A2(new_n13076_), .A3(new_n13075_), .ZN(new_n13150_));
  AOI22_X1   g12148(.A1(new_n13064_), .A2(new_n13073_), .B1(new_n12903_), .B2(new_n13011_), .ZN(new_n13151_));
  NOR2_X1    g12149(.A1(new_n13151_), .A2(new_n13150_), .ZN(new_n13152_));
  NOR3_X1    g12150(.A1(new_n13148_), .A2(new_n13152_), .A3(new_n13149_), .ZN(new_n13153_));
  OAI21_X1   g12151(.A1(new_n13148_), .A2(new_n13149_), .B(new_n13152_), .ZN(new_n13154_));
  AOI21_X1   g12152(.A1(new_n13154_), .A2(new_n13147_), .B(new_n13153_), .ZN(new_n13155_));
  NAND4_X1   g12153(.A1(new_n13120_), .A2(new_n13121_), .A3(new_n13118_), .A4(new_n13119_), .ZN(new_n13156_));
  OAI22_X1   g12154(.A1(new_n13116_), .A2(new_n13112_), .B1(new_n13096_), .B2(new_n13099_), .ZN(new_n13157_));
  NAND2_X1   g12155(.A1(new_n13157_), .A2(new_n13156_), .ZN(new_n13158_));
  NAND2_X1   g12156(.A1(new_n13155_), .A2(new_n13158_), .ZN(new_n13159_));
  INV_X1     g12157(.I(\A[583] ), .ZN(new_n13160_));
  INV_X1     g12158(.I(\A[584] ), .ZN(new_n13161_));
  NAND2_X1   g12159(.A1(new_n13161_), .A2(\A[585] ), .ZN(new_n13162_));
  INV_X1     g12160(.I(\A[585] ), .ZN(new_n13163_));
  NAND2_X1   g12161(.A1(new_n13163_), .A2(\A[584] ), .ZN(new_n13164_));
  AOI21_X1   g12162(.A1(new_n13162_), .A2(new_n13164_), .B(new_n13160_), .ZN(new_n13165_));
  NAND2_X1   g12163(.A1(\A[584] ), .A2(\A[585] ), .ZN(new_n13166_));
  NOR2_X1    g12164(.A1(\A[584] ), .A2(\A[585] ), .ZN(new_n13167_));
  INV_X1     g12165(.I(new_n13167_), .ZN(new_n13168_));
  AOI21_X1   g12166(.A1(new_n13168_), .A2(new_n13166_), .B(\A[583] ), .ZN(new_n13169_));
  INV_X1     g12167(.I(\A[586] ), .ZN(new_n13170_));
  INV_X1     g12168(.I(\A[587] ), .ZN(new_n13171_));
  NAND2_X1   g12169(.A1(new_n13171_), .A2(\A[588] ), .ZN(new_n13172_));
  INV_X1     g12170(.I(\A[588] ), .ZN(new_n13173_));
  NAND2_X1   g12171(.A1(new_n13173_), .A2(\A[587] ), .ZN(new_n13174_));
  AOI21_X1   g12172(.A1(new_n13172_), .A2(new_n13174_), .B(new_n13170_), .ZN(new_n13175_));
  NAND2_X1   g12173(.A1(\A[587] ), .A2(\A[588] ), .ZN(new_n13176_));
  NOR2_X1    g12174(.A1(\A[587] ), .A2(\A[588] ), .ZN(new_n13177_));
  INV_X1     g12175(.I(new_n13177_), .ZN(new_n13178_));
  AOI21_X1   g12176(.A1(new_n13178_), .A2(new_n13176_), .B(\A[586] ), .ZN(new_n13179_));
  NOR4_X1    g12177(.A1(new_n13165_), .A2(new_n13169_), .A3(new_n13179_), .A4(new_n13175_), .ZN(new_n13180_));
  AOI21_X1   g12178(.A1(new_n13170_), .A2(new_n13176_), .B(new_n13177_), .ZN(new_n13181_));
  AOI21_X1   g12179(.A1(\A[584] ), .A2(\A[585] ), .B(\A[583] ), .ZN(new_n13182_));
  NOR2_X1    g12180(.A1(new_n13182_), .A2(new_n13167_), .ZN(new_n13183_));
  NOR2_X1    g12181(.A1(new_n13181_), .A2(new_n13183_), .ZN(new_n13184_));
  INV_X1     g12182(.I(new_n13184_), .ZN(new_n13185_));
  NAND2_X1   g12183(.A1(new_n13181_), .A2(new_n13183_), .ZN(new_n13186_));
  NAND2_X1   g12184(.A1(new_n13185_), .A2(new_n13186_), .ZN(new_n13187_));
  XOR2_X1    g12185(.A1(new_n13187_), .A2(new_n13180_), .Z(new_n13188_));
  INV_X1     g12186(.I(\A[591] ), .ZN(new_n13189_));
  NOR2_X1    g12187(.A1(new_n13189_), .A2(\A[590] ), .ZN(new_n13190_));
  INV_X1     g12188(.I(\A[590] ), .ZN(new_n13191_));
  NOR2_X1    g12189(.A1(new_n13191_), .A2(\A[591] ), .ZN(new_n13192_));
  OAI21_X1   g12190(.A1(new_n13190_), .A2(new_n13192_), .B(\A[589] ), .ZN(new_n13193_));
  INV_X1     g12191(.I(\A[589] ), .ZN(new_n13194_));
  NOR2_X1    g12192(.A1(\A[590] ), .A2(\A[591] ), .ZN(new_n13195_));
  NOR2_X1    g12193(.A1(new_n13191_), .A2(new_n13189_), .ZN(new_n13196_));
  OAI21_X1   g12194(.A1(new_n13196_), .A2(new_n13195_), .B(new_n13194_), .ZN(new_n13197_));
  INV_X1     g12195(.I(\A[594] ), .ZN(new_n13198_));
  NOR2_X1    g12196(.A1(new_n13198_), .A2(\A[593] ), .ZN(new_n13199_));
  INV_X1     g12197(.I(\A[593] ), .ZN(new_n13200_));
  NOR2_X1    g12198(.A1(new_n13200_), .A2(\A[594] ), .ZN(new_n13201_));
  OAI21_X1   g12199(.A1(new_n13199_), .A2(new_n13201_), .B(\A[592] ), .ZN(new_n13202_));
  INV_X1     g12200(.I(\A[592] ), .ZN(new_n13203_));
  NOR2_X1    g12201(.A1(\A[593] ), .A2(\A[594] ), .ZN(new_n13204_));
  NOR2_X1    g12202(.A1(new_n13200_), .A2(new_n13198_), .ZN(new_n13205_));
  OAI21_X1   g12203(.A1(new_n13205_), .A2(new_n13204_), .B(new_n13203_), .ZN(new_n13206_));
  NAND4_X1   g12204(.A1(new_n13193_), .A2(new_n13197_), .A3(new_n13206_), .A4(new_n13202_), .ZN(new_n13207_));
  AOI21_X1   g12205(.A1(\A[593] ), .A2(\A[594] ), .B(\A[592] ), .ZN(new_n13208_));
  NOR2_X1    g12206(.A1(new_n13208_), .A2(new_n13204_), .ZN(new_n13209_));
  AOI21_X1   g12207(.A1(\A[590] ), .A2(\A[591] ), .B(\A[589] ), .ZN(new_n13210_));
  NOR2_X1    g12208(.A1(new_n13210_), .A2(new_n13195_), .ZN(new_n13211_));
  XNOR2_X1   g12209(.A1(new_n13209_), .A2(new_n13211_), .ZN(new_n13212_));
  XNOR2_X1   g12210(.A1(new_n13212_), .A2(new_n13207_), .ZN(new_n13213_));
  NAND2_X1   g12211(.A1(new_n13197_), .A2(new_n13193_), .ZN(new_n13214_));
  NAND2_X1   g12212(.A1(new_n13206_), .A2(new_n13202_), .ZN(new_n13215_));
  NAND2_X1   g12213(.A1(new_n13214_), .A2(new_n13215_), .ZN(new_n13216_));
  OAI22_X1   g12214(.A1(new_n13165_), .A2(new_n13169_), .B1(new_n13179_), .B2(new_n13175_), .ZN(new_n13217_));
  INV_X1     g12215(.I(new_n13217_), .ZN(new_n13218_));
  NOR2_X1    g12216(.A1(new_n13218_), .A2(new_n13180_), .ZN(new_n13219_));
  NAND3_X1   g12217(.A1(new_n13219_), .A2(new_n13207_), .A3(new_n13216_), .ZN(new_n13220_));
  AOI21_X1   g12218(.A1(new_n13213_), .A2(new_n13220_), .B(new_n13188_), .ZN(new_n13221_));
  XOR2_X1    g12219(.A1(new_n13212_), .A2(new_n13207_), .Z(new_n13222_));
  NAND2_X1   g12220(.A1(new_n13216_), .A2(new_n13207_), .ZN(new_n13223_));
  INV_X1     g12221(.I(new_n13180_), .ZN(new_n13224_));
  NAND2_X1   g12222(.A1(new_n13224_), .A2(new_n13217_), .ZN(new_n13225_));
  NOR2_X1    g12223(.A1(new_n13225_), .A2(new_n13223_), .ZN(new_n13226_));
  NAND2_X1   g12224(.A1(new_n13222_), .A2(new_n13226_), .ZN(new_n13227_));
  NAND2_X1   g12225(.A1(new_n13213_), .A2(new_n13220_), .ZN(new_n13228_));
  NAND2_X1   g12226(.A1(new_n13228_), .A2(new_n13227_), .ZN(new_n13229_));
  AOI22_X1   g12227(.A1(new_n13229_), .A2(new_n13188_), .B1(new_n13221_), .B2(new_n13227_), .ZN(new_n13230_));
  INV_X1     g12228(.I(\A[603] ), .ZN(new_n13231_));
  NOR2_X1    g12229(.A1(new_n13231_), .A2(\A[602] ), .ZN(new_n13232_));
  INV_X1     g12230(.I(\A[602] ), .ZN(new_n13233_));
  NOR2_X1    g12231(.A1(new_n13233_), .A2(\A[603] ), .ZN(new_n13234_));
  OAI21_X1   g12232(.A1(new_n13232_), .A2(new_n13234_), .B(\A[601] ), .ZN(new_n13235_));
  INV_X1     g12233(.I(\A[601] ), .ZN(new_n13236_));
  NOR2_X1    g12234(.A1(\A[602] ), .A2(\A[603] ), .ZN(new_n13237_));
  NAND2_X1   g12235(.A1(\A[602] ), .A2(\A[603] ), .ZN(new_n13238_));
  INV_X1     g12236(.I(new_n13238_), .ZN(new_n13239_));
  OAI21_X1   g12237(.A1(new_n13239_), .A2(new_n13237_), .B(new_n13236_), .ZN(new_n13240_));
  NAND2_X1   g12238(.A1(new_n13235_), .A2(new_n13240_), .ZN(new_n13241_));
  INV_X1     g12239(.I(\A[606] ), .ZN(new_n13242_));
  NOR2_X1    g12240(.A1(new_n13242_), .A2(\A[605] ), .ZN(new_n13243_));
  INV_X1     g12241(.I(\A[605] ), .ZN(new_n13244_));
  NOR2_X1    g12242(.A1(new_n13244_), .A2(\A[606] ), .ZN(new_n13245_));
  OAI21_X1   g12243(.A1(new_n13243_), .A2(new_n13245_), .B(\A[604] ), .ZN(new_n13246_));
  INV_X1     g12244(.I(\A[604] ), .ZN(new_n13247_));
  NOR2_X1    g12245(.A1(\A[605] ), .A2(\A[606] ), .ZN(new_n13248_));
  NAND2_X1   g12246(.A1(\A[605] ), .A2(\A[606] ), .ZN(new_n13249_));
  INV_X1     g12247(.I(new_n13249_), .ZN(new_n13250_));
  OAI21_X1   g12248(.A1(new_n13250_), .A2(new_n13248_), .B(new_n13247_), .ZN(new_n13251_));
  NAND2_X1   g12249(.A1(new_n13246_), .A2(new_n13251_), .ZN(new_n13252_));
  NOR2_X1    g12250(.A1(new_n13241_), .A2(new_n13252_), .ZN(new_n13253_));
  NAND2_X1   g12251(.A1(new_n13233_), .A2(\A[603] ), .ZN(new_n13254_));
  NAND2_X1   g12252(.A1(new_n13231_), .A2(\A[602] ), .ZN(new_n13255_));
  AOI21_X1   g12253(.A1(new_n13254_), .A2(new_n13255_), .B(new_n13236_), .ZN(new_n13256_));
  INV_X1     g12254(.I(new_n13237_), .ZN(new_n13257_));
  AOI21_X1   g12255(.A1(new_n13257_), .A2(new_n13238_), .B(\A[601] ), .ZN(new_n13258_));
  NOR2_X1    g12256(.A1(new_n13258_), .A2(new_n13256_), .ZN(new_n13259_));
  NAND2_X1   g12257(.A1(new_n13244_), .A2(\A[606] ), .ZN(new_n13260_));
  NAND2_X1   g12258(.A1(new_n13242_), .A2(\A[605] ), .ZN(new_n13261_));
  AOI21_X1   g12259(.A1(new_n13260_), .A2(new_n13261_), .B(new_n13247_), .ZN(new_n13262_));
  INV_X1     g12260(.I(new_n13248_), .ZN(new_n13263_));
  AOI21_X1   g12261(.A1(new_n13263_), .A2(new_n13249_), .B(\A[604] ), .ZN(new_n13264_));
  NOR2_X1    g12262(.A1(new_n13264_), .A2(new_n13262_), .ZN(new_n13265_));
  NOR2_X1    g12263(.A1(new_n13259_), .A2(new_n13265_), .ZN(new_n13266_));
  NOR2_X1    g12264(.A1(new_n13266_), .A2(new_n13253_), .ZN(new_n13267_));
  INV_X1     g12265(.I(\A[595] ), .ZN(new_n13268_));
  INV_X1     g12266(.I(\A[596] ), .ZN(new_n13269_));
  NAND2_X1   g12267(.A1(new_n13269_), .A2(\A[597] ), .ZN(new_n13270_));
  INV_X1     g12268(.I(\A[597] ), .ZN(new_n13271_));
  NAND2_X1   g12269(.A1(new_n13271_), .A2(\A[596] ), .ZN(new_n13272_));
  AOI21_X1   g12270(.A1(new_n13270_), .A2(new_n13272_), .B(new_n13268_), .ZN(new_n13273_));
  NAND2_X1   g12271(.A1(\A[596] ), .A2(\A[597] ), .ZN(new_n13274_));
  NOR2_X1    g12272(.A1(\A[596] ), .A2(\A[597] ), .ZN(new_n13275_));
  INV_X1     g12273(.I(new_n13275_), .ZN(new_n13276_));
  AOI21_X1   g12274(.A1(new_n13276_), .A2(new_n13274_), .B(\A[595] ), .ZN(new_n13277_));
  NOR2_X1    g12275(.A1(new_n13277_), .A2(new_n13273_), .ZN(new_n13278_));
  INV_X1     g12276(.I(\A[598] ), .ZN(new_n13279_));
  INV_X1     g12277(.I(\A[599] ), .ZN(new_n13280_));
  NAND2_X1   g12278(.A1(new_n13280_), .A2(\A[600] ), .ZN(new_n13281_));
  INV_X1     g12279(.I(\A[600] ), .ZN(new_n13282_));
  NAND2_X1   g12280(.A1(new_n13282_), .A2(\A[599] ), .ZN(new_n13283_));
  AOI21_X1   g12281(.A1(new_n13281_), .A2(new_n13283_), .B(new_n13279_), .ZN(new_n13284_));
  NAND2_X1   g12282(.A1(\A[599] ), .A2(\A[600] ), .ZN(new_n13285_));
  NOR2_X1    g12283(.A1(\A[599] ), .A2(\A[600] ), .ZN(new_n13286_));
  INV_X1     g12284(.I(new_n13286_), .ZN(new_n13287_));
  AOI21_X1   g12285(.A1(new_n13287_), .A2(new_n13285_), .B(\A[598] ), .ZN(new_n13288_));
  NOR2_X1    g12286(.A1(new_n13288_), .A2(new_n13284_), .ZN(new_n13289_));
  NAND2_X1   g12287(.A1(new_n13278_), .A2(new_n13289_), .ZN(new_n13290_));
  NOR2_X1    g12288(.A1(new_n13271_), .A2(\A[596] ), .ZN(new_n13291_));
  NOR2_X1    g12289(.A1(new_n13269_), .A2(\A[597] ), .ZN(new_n13292_));
  OAI21_X1   g12290(.A1(new_n13291_), .A2(new_n13292_), .B(\A[595] ), .ZN(new_n13293_));
  INV_X1     g12291(.I(new_n13274_), .ZN(new_n13294_));
  OAI21_X1   g12292(.A1(new_n13294_), .A2(new_n13275_), .B(new_n13268_), .ZN(new_n13295_));
  NAND2_X1   g12293(.A1(new_n13293_), .A2(new_n13295_), .ZN(new_n13296_));
  NOR2_X1    g12294(.A1(new_n13282_), .A2(\A[599] ), .ZN(new_n13297_));
  NOR2_X1    g12295(.A1(new_n13280_), .A2(\A[600] ), .ZN(new_n13298_));
  OAI21_X1   g12296(.A1(new_n13297_), .A2(new_n13298_), .B(\A[598] ), .ZN(new_n13299_));
  INV_X1     g12297(.I(new_n13285_), .ZN(new_n13300_));
  OAI21_X1   g12298(.A1(new_n13300_), .A2(new_n13286_), .B(new_n13279_), .ZN(new_n13301_));
  NAND2_X1   g12299(.A1(new_n13299_), .A2(new_n13301_), .ZN(new_n13302_));
  NAND2_X1   g12300(.A1(new_n13296_), .A2(new_n13302_), .ZN(new_n13303_));
  NAND2_X1   g12301(.A1(new_n13290_), .A2(new_n13303_), .ZN(new_n13304_));
  NAND2_X1   g12302(.A1(new_n13267_), .A2(new_n13304_), .ZN(new_n13305_));
  NAND2_X1   g12303(.A1(new_n13259_), .A2(new_n13265_), .ZN(new_n13306_));
  NAND2_X1   g12304(.A1(new_n13241_), .A2(new_n13252_), .ZN(new_n13307_));
  NAND2_X1   g12305(.A1(new_n13306_), .A2(new_n13307_), .ZN(new_n13308_));
  NOR2_X1    g12306(.A1(new_n13296_), .A2(new_n13302_), .ZN(new_n13309_));
  NOR2_X1    g12307(.A1(new_n13278_), .A2(new_n13289_), .ZN(new_n13310_));
  NOR2_X1    g12308(.A1(new_n13310_), .A2(new_n13309_), .ZN(new_n13311_));
  NAND2_X1   g12309(.A1(new_n13311_), .A2(new_n13308_), .ZN(new_n13312_));
  NAND3_X1   g12310(.A1(new_n13225_), .A2(new_n13207_), .A3(new_n13216_), .ZN(new_n13313_));
  NAND2_X1   g12311(.A1(new_n13219_), .A2(new_n13223_), .ZN(new_n13314_));
  AOI22_X1   g12312(.A1(new_n13305_), .A2(new_n13312_), .B1(new_n13313_), .B2(new_n13314_), .ZN(new_n13315_));
  INV_X1     g12313(.I(new_n13315_), .ZN(new_n13316_));
  AOI21_X1   g12314(.A1(\A[599] ), .A2(\A[600] ), .B(\A[598] ), .ZN(new_n13317_));
  AOI21_X1   g12315(.A1(\A[596] ), .A2(\A[597] ), .B(\A[595] ), .ZN(new_n13318_));
  OAI22_X1   g12316(.A1(new_n13275_), .A2(new_n13318_), .B1(new_n13317_), .B2(new_n13286_), .ZN(new_n13319_));
  NOR4_X1    g12317(.A1(new_n13317_), .A2(new_n13318_), .A3(new_n13275_), .A4(new_n13286_), .ZN(new_n13320_));
  INV_X1     g12318(.I(new_n13320_), .ZN(new_n13321_));
  NAND2_X1   g12319(.A1(new_n13321_), .A2(new_n13319_), .ZN(new_n13322_));
  XOR2_X1    g12320(.A1(new_n13309_), .A2(new_n13322_), .Z(new_n13323_));
  AOI21_X1   g12321(.A1(new_n13247_), .A2(new_n13249_), .B(new_n13248_), .ZN(new_n13324_));
  AOI21_X1   g12322(.A1(new_n13236_), .A2(new_n13238_), .B(new_n13237_), .ZN(new_n13325_));
  XOR2_X1    g12323(.A1(new_n13324_), .A2(new_n13325_), .Z(new_n13326_));
  NOR2_X1    g12324(.A1(new_n13253_), .A2(new_n13326_), .ZN(new_n13327_));
  XNOR2_X1   g12325(.A1(new_n13324_), .A2(new_n13325_), .ZN(new_n13328_));
  NOR2_X1    g12326(.A1(new_n13306_), .A2(new_n13328_), .ZN(new_n13329_));
  OAI22_X1   g12327(.A1(new_n13308_), .A2(new_n13304_), .B1(new_n13329_), .B2(new_n13327_), .ZN(new_n13330_));
  NAND4_X1   g12328(.A1(new_n13311_), .A2(new_n13306_), .A3(new_n13307_), .A4(new_n13326_), .ZN(new_n13331_));
  NAND3_X1   g12329(.A1(new_n13330_), .A2(new_n13323_), .A3(new_n13331_), .ZN(new_n13332_));
  AOI21_X1   g12330(.A1(new_n13330_), .A2(new_n13331_), .B(new_n13323_), .ZN(new_n13333_));
  INV_X1     g12331(.I(new_n13333_), .ZN(new_n13334_));
  AOI21_X1   g12332(.A1(new_n13334_), .A2(new_n13332_), .B(new_n13316_), .ZN(new_n13335_));
  INV_X1     g12333(.I(new_n13332_), .ZN(new_n13336_));
  NOR3_X1    g12334(.A1(new_n13336_), .A2(new_n13315_), .A3(new_n13333_), .ZN(new_n13337_));
  NOR3_X1    g12335(.A1(new_n13335_), .A2(new_n13337_), .A3(new_n13230_), .ZN(new_n13338_));
  XNOR2_X1   g12336(.A1(new_n13187_), .A2(new_n13180_), .ZN(new_n13339_));
  OAI21_X1   g12337(.A1(new_n13222_), .A2(new_n13226_), .B(new_n13339_), .ZN(new_n13340_));
  NOR2_X1    g12338(.A1(new_n13213_), .A2(new_n13220_), .ZN(new_n13341_));
  NOR2_X1    g12339(.A1(new_n13222_), .A2(new_n13226_), .ZN(new_n13342_));
  NOR2_X1    g12340(.A1(new_n13341_), .A2(new_n13342_), .ZN(new_n13343_));
  OAI22_X1   g12341(.A1(new_n13343_), .A2(new_n13339_), .B1(new_n13340_), .B2(new_n13341_), .ZN(new_n13344_));
  OAI21_X1   g12342(.A1(new_n13336_), .A2(new_n13333_), .B(new_n13315_), .ZN(new_n13345_));
  NAND3_X1   g12343(.A1(new_n13316_), .A2(new_n13334_), .A3(new_n13332_), .ZN(new_n13346_));
  AOI21_X1   g12344(.A1(new_n13346_), .A2(new_n13345_), .B(new_n13344_), .ZN(new_n13347_));
  NOR2_X1    g12345(.A1(new_n13338_), .A2(new_n13347_), .ZN(new_n13348_));
  INV_X1     g12346(.I(new_n13348_), .ZN(new_n13349_));
  INV_X1     g12347(.I(\A[571] ), .ZN(new_n13350_));
  INV_X1     g12348(.I(\A[572] ), .ZN(new_n13351_));
  NAND2_X1   g12349(.A1(new_n13351_), .A2(\A[573] ), .ZN(new_n13352_));
  INV_X1     g12350(.I(\A[573] ), .ZN(new_n13353_));
  NAND2_X1   g12351(.A1(new_n13353_), .A2(\A[572] ), .ZN(new_n13354_));
  AOI21_X1   g12352(.A1(new_n13352_), .A2(new_n13354_), .B(new_n13350_), .ZN(new_n13355_));
  NAND2_X1   g12353(.A1(\A[572] ), .A2(\A[573] ), .ZN(new_n13356_));
  NOR2_X1    g12354(.A1(\A[572] ), .A2(\A[573] ), .ZN(new_n13357_));
  INV_X1     g12355(.I(new_n13357_), .ZN(new_n13358_));
  AOI21_X1   g12356(.A1(new_n13358_), .A2(new_n13356_), .B(\A[571] ), .ZN(new_n13359_));
  NOR2_X1    g12357(.A1(new_n13359_), .A2(new_n13355_), .ZN(new_n13360_));
  INV_X1     g12358(.I(\A[574] ), .ZN(new_n13361_));
  INV_X1     g12359(.I(\A[575] ), .ZN(new_n13362_));
  NAND2_X1   g12360(.A1(new_n13362_), .A2(\A[576] ), .ZN(new_n13363_));
  INV_X1     g12361(.I(\A[576] ), .ZN(new_n13364_));
  NAND2_X1   g12362(.A1(new_n13364_), .A2(\A[575] ), .ZN(new_n13365_));
  AOI21_X1   g12363(.A1(new_n13363_), .A2(new_n13365_), .B(new_n13361_), .ZN(new_n13366_));
  NAND2_X1   g12364(.A1(\A[575] ), .A2(\A[576] ), .ZN(new_n13367_));
  NOR2_X1    g12365(.A1(\A[575] ), .A2(\A[576] ), .ZN(new_n13368_));
  INV_X1     g12366(.I(new_n13368_), .ZN(new_n13369_));
  AOI21_X1   g12367(.A1(new_n13369_), .A2(new_n13367_), .B(\A[574] ), .ZN(new_n13370_));
  NOR2_X1    g12368(.A1(new_n13370_), .A2(new_n13366_), .ZN(new_n13371_));
  NAND2_X1   g12369(.A1(new_n13360_), .A2(new_n13371_), .ZN(new_n13372_));
  AOI21_X1   g12370(.A1(new_n13361_), .A2(new_n13367_), .B(new_n13368_), .ZN(new_n13373_));
  AOI21_X1   g12371(.A1(new_n13350_), .A2(new_n13356_), .B(new_n13357_), .ZN(new_n13374_));
  NOR2_X1    g12372(.A1(new_n13373_), .A2(new_n13374_), .ZN(new_n13375_));
  NAND2_X1   g12373(.A1(new_n13373_), .A2(new_n13374_), .ZN(new_n13376_));
  INV_X1     g12374(.I(new_n13376_), .ZN(new_n13377_));
  NOR2_X1    g12375(.A1(new_n13377_), .A2(new_n13375_), .ZN(new_n13378_));
  XOR2_X1    g12376(.A1(new_n13378_), .A2(new_n13372_), .Z(new_n13379_));
  INV_X1     g12377(.I(\A[579] ), .ZN(new_n13380_));
  NOR2_X1    g12378(.A1(new_n13380_), .A2(\A[578] ), .ZN(new_n13381_));
  INV_X1     g12379(.I(\A[578] ), .ZN(new_n13382_));
  NOR2_X1    g12380(.A1(new_n13382_), .A2(\A[579] ), .ZN(new_n13383_));
  OAI21_X1   g12381(.A1(new_n13381_), .A2(new_n13383_), .B(\A[577] ), .ZN(new_n13384_));
  INV_X1     g12382(.I(\A[577] ), .ZN(new_n13385_));
  NOR2_X1    g12383(.A1(\A[578] ), .A2(\A[579] ), .ZN(new_n13386_));
  NAND2_X1   g12384(.A1(\A[578] ), .A2(\A[579] ), .ZN(new_n13387_));
  INV_X1     g12385(.I(new_n13387_), .ZN(new_n13388_));
  OAI21_X1   g12386(.A1(new_n13388_), .A2(new_n13386_), .B(new_n13385_), .ZN(new_n13389_));
  NAND2_X1   g12387(.A1(new_n13384_), .A2(new_n13389_), .ZN(new_n13390_));
  INV_X1     g12388(.I(\A[582] ), .ZN(new_n13391_));
  NOR2_X1    g12389(.A1(new_n13391_), .A2(\A[581] ), .ZN(new_n13392_));
  INV_X1     g12390(.I(\A[581] ), .ZN(new_n13393_));
  NOR2_X1    g12391(.A1(new_n13393_), .A2(\A[582] ), .ZN(new_n13394_));
  OAI21_X1   g12392(.A1(new_n13392_), .A2(new_n13394_), .B(\A[580] ), .ZN(new_n13395_));
  INV_X1     g12393(.I(\A[580] ), .ZN(new_n13396_));
  NOR2_X1    g12394(.A1(\A[581] ), .A2(\A[582] ), .ZN(new_n13397_));
  NAND2_X1   g12395(.A1(\A[581] ), .A2(\A[582] ), .ZN(new_n13398_));
  INV_X1     g12396(.I(new_n13398_), .ZN(new_n13399_));
  OAI21_X1   g12397(.A1(new_n13399_), .A2(new_n13397_), .B(new_n13396_), .ZN(new_n13400_));
  NAND2_X1   g12398(.A1(new_n13395_), .A2(new_n13400_), .ZN(new_n13401_));
  NOR2_X1    g12399(.A1(new_n13390_), .A2(new_n13401_), .ZN(new_n13402_));
  AOI21_X1   g12400(.A1(new_n13396_), .A2(new_n13398_), .B(new_n13397_), .ZN(new_n13403_));
  AOI21_X1   g12401(.A1(new_n13385_), .A2(new_n13387_), .B(new_n13386_), .ZN(new_n13404_));
  XNOR2_X1   g12402(.A1(new_n13403_), .A2(new_n13404_), .ZN(new_n13405_));
  XOR2_X1    g12403(.A1(new_n13402_), .A2(new_n13405_), .Z(new_n13406_));
  NAND2_X1   g12404(.A1(new_n13382_), .A2(\A[579] ), .ZN(new_n13407_));
  NAND2_X1   g12405(.A1(new_n13380_), .A2(\A[578] ), .ZN(new_n13408_));
  AOI21_X1   g12406(.A1(new_n13407_), .A2(new_n13408_), .B(new_n13385_), .ZN(new_n13409_));
  INV_X1     g12407(.I(new_n13386_), .ZN(new_n13410_));
  AOI21_X1   g12408(.A1(new_n13410_), .A2(new_n13387_), .B(\A[577] ), .ZN(new_n13411_));
  NOR2_X1    g12409(.A1(new_n13411_), .A2(new_n13409_), .ZN(new_n13412_));
  NAND2_X1   g12410(.A1(new_n13393_), .A2(\A[582] ), .ZN(new_n13413_));
  NAND2_X1   g12411(.A1(new_n13391_), .A2(\A[581] ), .ZN(new_n13414_));
  AOI21_X1   g12412(.A1(new_n13413_), .A2(new_n13414_), .B(new_n13396_), .ZN(new_n13415_));
  INV_X1     g12413(.I(new_n13397_), .ZN(new_n13416_));
  AOI21_X1   g12414(.A1(new_n13416_), .A2(new_n13398_), .B(\A[580] ), .ZN(new_n13417_));
  NOR2_X1    g12415(.A1(new_n13417_), .A2(new_n13415_), .ZN(new_n13418_));
  NOR2_X1    g12416(.A1(new_n13412_), .A2(new_n13418_), .ZN(new_n13419_));
  NOR2_X1    g12417(.A1(new_n13419_), .A2(new_n13402_), .ZN(new_n13420_));
  NOR2_X1    g12418(.A1(new_n13353_), .A2(\A[572] ), .ZN(new_n13421_));
  NOR2_X1    g12419(.A1(new_n13351_), .A2(\A[573] ), .ZN(new_n13422_));
  OAI21_X1   g12420(.A1(new_n13421_), .A2(new_n13422_), .B(\A[571] ), .ZN(new_n13423_));
  INV_X1     g12421(.I(new_n13356_), .ZN(new_n13424_));
  OAI21_X1   g12422(.A1(new_n13424_), .A2(new_n13357_), .B(new_n13350_), .ZN(new_n13425_));
  NAND2_X1   g12423(.A1(new_n13423_), .A2(new_n13425_), .ZN(new_n13426_));
  NOR2_X1    g12424(.A1(new_n13364_), .A2(\A[575] ), .ZN(new_n13427_));
  NOR2_X1    g12425(.A1(new_n13362_), .A2(\A[576] ), .ZN(new_n13428_));
  OAI21_X1   g12426(.A1(new_n13427_), .A2(new_n13428_), .B(\A[574] ), .ZN(new_n13429_));
  INV_X1     g12427(.I(new_n13367_), .ZN(new_n13430_));
  OAI21_X1   g12428(.A1(new_n13430_), .A2(new_n13368_), .B(new_n13361_), .ZN(new_n13431_));
  NAND2_X1   g12429(.A1(new_n13429_), .A2(new_n13431_), .ZN(new_n13432_));
  NOR2_X1    g12430(.A1(new_n13426_), .A2(new_n13432_), .ZN(new_n13433_));
  NOR2_X1    g12431(.A1(new_n13360_), .A2(new_n13371_), .ZN(new_n13434_));
  NOR2_X1    g12432(.A1(new_n13434_), .A2(new_n13433_), .ZN(new_n13435_));
  NAND2_X1   g12433(.A1(new_n13435_), .A2(new_n13420_), .ZN(new_n13436_));
  NAND2_X1   g12434(.A1(new_n13406_), .A2(new_n13436_), .ZN(new_n13437_));
  NAND2_X1   g12435(.A1(new_n13426_), .A2(new_n13432_), .ZN(new_n13438_));
  NAND2_X1   g12436(.A1(new_n13372_), .A2(new_n13438_), .ZN(new_n13439_));
  NOR4_X1    g12437(.A1(new_n13439_), .A2(new_n13402_), .A3(new_n13405_), .A4(new_n13419_), .ZN(new_n13440_));
  INV_X1     g12438(.I(new_n13440_), .ZN(new_n13441_));
  NAND3_X1   g12439(.A1(new_n13437_), .A2(new_n13441_), .A3(new_n13379_), .ZN(new_n13442_));
  NAND2_X1   g12440(.A1(new_n13378_), .A2(new_n13372_), .ZN(new_n13443_));
  OAI21_X1   g12441(.A1(new_n13375_), .A2(new_n13377_), .B(new_n13433_), .ZN(new_n13444_));
  NAND2_X1   g12442(.A1(new_n13444_), .A2(new_n13443_), .ZN(new_n13445_));
  NAND2_X1   g12443(.A1(new_n13412_), .A2(new_n13418_), .ZN(new_n13446_));
  XOR2_X1    g12444(.A1(new_n13446_), .A2(new_n13405_), .Z(new_n13447_));
  NAND2_X1   g12445(.A1(new_n13390_), .A2(new_n13401_), .ZN(new_n13448_));
  NAND2_X1   g12446(.A1(new_n13446_), .A2(new_n13448_), .ZN(new_n13449_));
  NOR2_X1    g12447(.A1(new_n13449_), .A2(new_n13439_), .ZN(new_n13450_));
  NOR2_X1    g12448(.A1(new_n13447_), .A2(new_n13450_), .ZN(new_n13451_));
  OAI21_X1   g12449(.A1(new_n13451_), .A2(new_n13440_), .B(new_n13445_), .ZN(new_n13452_));
  NAND2_X1   g12450(.A1(new_n13452_), .A2(new_n13442_), .ZN(new_n13453_));
  INV_X1     g12451(.I(\A[559] ), .ZN(new_n13454_));
  INV_X1     g12452(.I(\A[560] ), .ZN(new_n13455_));
  NAND2_X1   g12453(.A1(new_n13455_), .A2(\A[561] ), .ZN(new_n13456_));
  INV_X1     g12454(.I(\A[561] ), .ZN(new_n13457_));
  NAND2_X1   g12455(.A1(new_n13457_), .A2(\A[560] ), .ZN(new_n13458_));
  AOI21_X1   g12456(.A1(new_n13456_), .A2(new_n13458_), .B(new_n13454_), .ZN(new_n13459_));
  NAND2_X1   g12457(.A1(\A[560] ), .A2(\A[561] ), .ZN(new_n13460_));
  NOR2_X1    g12458(.A1(\A[560] ), .A2(\A[561] ), .ZN(new_n13461_));
  INV_X1     g12459(.I(new_n13461_), .ZN(new_n13462_));
  AOI21_X1   g12460(.A1(new_n13462_), .A2(new_n13460_), .B(\A[559] ), .ZN(new_n13463_));
  INV_X1     g12461(.I(\A[562] ), .ZN(new_n13464_));
  INV_X1     g12462(.I(\A[563] ), .ZN(new_n13465_));
  NAND2_X1   g12463(.A1(new_n13465_), .A2(\A[564] ), .ZN(new_n13466_));
  INV_X1     g12464(.I(\A[564] ), .ZN(new_n13467_));
  NAND2_X1   g12465(.A1(new_n13467_), .A2(\A[563] ), .ZN(new_n13468_));
  AOI21_X1   g12466(.A1(new_n13466_), .A2(new_n13468_), .B(new_n13464_), .ZN(new_n13469_));
  NAND2_X1   g12467(.A1(\A[563] ), .A2(\A[564] ), .ZN(new_n13470_));
  NOR2_X1    g12468(.A1(\A[563] ), .A2(\A[564] ), .ZN(new_n13471_));
  INV_X1     g12469(.I(new_n13471_), .ZN(new_n13472_));
  AOI21_X1   g12470(.A1(new_n13472_), .A2(new_n13470_), .B(\A[562] ), .ZN(new_n13473_));
  NOR4_X1    g12471(.A1(new_n13459_), .A2(new_n13463_), .A3(new_n13473_), .A4(new_n13469_), .ZN(new_n13474_));
  AOI21_X1   g12472(.A1(new_n13464_), .A2(new_n13470_), .B(new_n13471_), .ZN(new_n13475_));
  AOI21_X1   g12473(.A1(new_n13454_), .A2(new_n13460_), .B(new_n13461_), .ZN(new_n13476_));
  NOR2_X1    g12474(.A1(new_n13475_), .A2(new_n13476_), .ZN(new_n13477_));
  NAND2_X1   g12475(.A1(new_n13475_), .A2(new_n13476_), .ZN(new_n13478_));
  INV_X1     g12476(.I(new_n13478_), .ZN(new_n13479_));
  NOR2_X1    g12477(.A1(new_n13479_), .A2(new_n13477_), .ZN(new_n13480_));
  XOR2_X1    g12478(.A1(new_n13480_), .A2(new_n13474_), .Z(new_n13481_));
  INV_X1     g12479(.I(\A[567] ), .ZN(new_n13482_));
  NOR2_X1    g12480(.A1(new_n13482_), .A2(\A[566] ), .ZN(new_n13483_));
  INV_X1     g12481(.I(\A[566] ), .ZN(new_n13484_));
  NOR2_X1    g12482(.A1(new_n13484_), .A2(\A[567] ), .ZN(new_n13485_));
  OAI21_X1   g12483(.A1(new_n13483_), .A2(new_n13485_), .B(\A[565] ), .ZN(new_n13486_));
  INV_X1     g12484(.I(\A[565] ), .ZN(new_n13487_));
  NOR2_X1    g12485(.A1(\A[566] ), .A2(\A[567] ), .ZN(new_n13488_));
  NAND2_X1   g12486(.A1(\A[566] ), .A2(\A[567] ), .ZN(new_n13489_));
  INV_X1     g12487(.I(new_n13489_), .ZN(new_n13490_));
  OAI21_X1   g12488(.A1(new_n13490_), .A2(new_n13488_), .B(new_n13487_), .ZN(new_n13491_));
  NAND2_X1   g12489(.A1(new_n13486_), .A2(new_n13491_), .ZN(new_n13492_));
  INV_X1     g12490(.I(\A[570] ), .ZN(new_n13493_));
  NOR2_X1    g12491(.A1(new_n13493_), .A2(\A[569] ), .ZN(new_n13494_));
  INV_X1     g12492(.I(\A[569] ), .ZN(new_n13495_));
  NOR2_X1    g12493(.A1(new_n13495_), .A2(\A[570] ), .ZN(new_n13496_));
  OAI21_X1   g12494(.A1(new_n13494_), .A2(new_n13496_), .B(\A[568] ), .ZN(new_n13497_));
  INV_X1     g12495(.I(\A[568] ), .ZN(new_n13498_));
  NOR2_X1    g12496(.A1(\A[569] ), .A2(\A[570] ), .ZN(new_n13499_));
  NAND2_X1   g12497(.A1(\A[569] ), .A2(\A[570] ), .ZN(new_n13500_));
  INV_X1     g12498(.I(new_n13500_), .ZN(new_n13501_));
  OAI21_X1   g12499(.A1(new_n13501_), .A2(new_n13499_), .B(new_n13498_), .ZN(new_n13502_));
  NAND2_X1   g12500(.A1(new_n13497_), .A2(new_n13502_), .ZN(new_n13503_));
  NOR2_X1    g12501(.A1(new_n13492_), .A2(new_n13503_), .ZN(new_n13504_));
  AOI21_X1   g12502(.A1(new_n13498_), .A2(new_n13500_), .B(new_n13499_), .ZN(new_n13505_));
  AOI21_X1   g12503(.A1(new_n13487_), .A2(new_n13489_), .B(new_n13488_), .ZN(new_n13506_));
  XOR2_X1    g12504(.A1(new_n13505_), .A2(new_n13506_), .Z(new_n13507_));
  NOR2_X1    g12505(.A1(new_n13504_), .A2(new_n13507_), .ZN(new_n13508_));
  NAND2_X1   g12506(.A1(new_n13484_), .A2(\A[567] ), .ZN(new_n13509_));
  NAND2_X1   g12507(.A1(new_n13482_), .A2(\A[566] ), .ZN(new_n13510_));
  AOI21_X1   g12508(.A1(new_n13509_), .A2(new_n13510_), .B(new_n13487_), .ZN(new_n13511_));
  INV_X1     g12509(.I(new_n13488_), .ZN(new_n13512_));
  AOI21_X1   g12510(.A1(new_n13512_), .A2(new_n13489_), .B(\A[565] ), .ZN(new_n13513_));
  NOR2_X1    g12511(.A1(new_n13513_), .A2(new_n13511_), .ZN(new_n13514_));
  NAND2_X1   g12512(.A1(new_n13495_), .A2(\A[570] ), .ZN(new_n13515_));
  NAND2_X1   g12513(.A1(new_n13493_), .A2(\A[569] ), .ZN(new_n13516_));
  AOI21_X1   g12514(.A1(new_n13515_), .A2(new_n13516_), .B(new_n13498_), .ZN(new_n13517_));
  INV_X1     g12515(.I(new_n13499_), .ZN(new_n13518_));
  AOI21_X1   g12516(.A1(new_n13518_), .A2(new_n13500_), .B(\A[568] ), .ZN(new_n13519_));
  NOR2_X1    g12517(.A1(new_n13519_), .A2(new_n13517_), .ZN(new_n13520_));
  NAND2_X1   g12518(.A1(new_n13514_), .A2(new_n13520_), .ZN(new_n13521_));
  XNOR2_X1   g12519(.A1(new_n13505_), .A2(new_n13506_), .ZN(new_n13522_));
  NOR2_X1    g12520(.A1(new_n13521_), .A2(new_n13522_), .ZN(new_n13523_));
  NAND2_X1   g12521(.A1(new_n13492_), .A2(new_n13503_), .ZN(new_n13524_));
  NAND2_X1   g12522(.A1(new_n13521_), .A2(new_n13524_), .ZN(new_n13525_));
  INV_X1     g12523(.I(new_n13474_), .ZN(new_n13526_));
  OAI22_X1   g12524(.A1(new_n13459_), .A2(new_n13463_), .B1(new_n13473_), .B2(new_n13469_), .ZN(new_n13527_));
  NAND2_X1   g12525(.A1(new_n13526_), .A2(new_n13527_), .ZN(new_n13528_));
  OAI22_X1   g12526(.A1(new_n13525_), .A2(new_n13528_), .B1(new_n13523_), .B2(new_n13508_), .ZN(new_n13529_));
  NOR2_X1    g12527(.A1(new_n13514_), .A2(new_n13520_), .ZN(new_n13530_));
  NOR4_X1    g12528(.A1(new_n13528_), .A2(new_n13504_), .A3(new_n13522_), .A4(new_n13530_), .ZN(new_n13531_));
  INV_X1     g12529(.I(new_n13531_), .ZN(new_n13532_));
  NAND3_X1   g12530(.A1(new_n13532_), .A2(new_n13529_), .A3(new_n13481_), .ZN(new_n13533_));
  XNOR2_X1   g12531(.A1(new_n13480_), .A2(new_n13474_), .ZN(new_n13534_));
  INV_X1     g12532(.I(new_n13529_), .ZN(new_n13535_));
  OAI21_X1   g12533(.A1(new_n13535_), .A2(new_n13531_), .B(new_n13534_), .ZN(new_n13536_));
  NOR2_X1    g12534(.A1(new_n13435_), .A2(new_n13449_), .ZN(new_n13537_));
  NOR2_X1    g12535(.A1(new_n13420_), .A2(new_n13439_), .ZN(new_n13538_));
  INV_X1     g12536(.I(new_n13527_), .ZN(new_n13539_));
  NOR2_X1    g12537(.A1(new_n13539_), .A2(new_n13474_), .ZN(new_n13540_));
  NOR2_X1    g12538(.A1(new_n13540_), .A2(new_n13525_), .ZN(new_n13541_));
  NOR2_X1    g12539(.A1(new_n13530_), .A2(new_n13504_), .ZN(new_n13542_));
  NOR2_X1    g12540(.A1(new_n13528_), .A2(new_n13542_), .ZN(new_n13543_));
  OAI22_X1   g12541(.A1(new_n13537_), .A2(new_n13538_), .B1(new_n13543_), .B2(new_n13541_), .ZN(new_n13544_));
  INV_X1     g12542(.I(new_n13544_), .ZN(new_n13545_));
  NAND3_X1   g12543(.A1(new_n13545_), .A2(new_n13536_), .A3(new_n13533_), .ZN(new_n13546_));
  NOR3_X1    g12544(.A1(new_n13535_), .A2(new_n13534_), .A3(new_n13531_), .ZN(new_n13547_));
  AOI21_X1   g12545(.A1(new_n13532_), .A2(new_n13529_), .B(new_n13481_), .ZN(new_n13548_));
  OAI21_X1   g12546(.A1(new_n13547_), .A2(new_n13548_), .B(new_n13544_), .ZN(new_n13549_));
  NAND3_X1   g12547(.A1(new_n13546_), .A2(new_n13549_), .A3(new_n13453_), .ZN(new_n13550_));
  AND2_X2    g12548(.A1(new_n13452_), .A2(new_n13442_), .Z(new_n13551_));
  NOR3_X1    g12549(.A1(new_n13547_), .A2(new_n13548_), .A3(new_n13544_), .ZN(new_n13552_));
  AOI21_X1   g12550(.A1(new_n13536_), .A2(new_n13533_), .B(new_n13545_), .ZN(new_n13553_));
  OAI21_X1   g12551(.A1(new_n13552_), .A2(new_n13553_), .B(new_n13551_), .ZN(new_n13554_));
  NAND2_X1   g12552(.A1(new_n13305_), .A2(new_n13312_), .ZN(new_n13555_));
  NAND2_X1   g12553(.A1(new_n13313_), .A2(new_n13314_), .ZN(new_n13556_));
  NOR2_X1    g12554(.A1(new_n13555_), .A2(new_n13556_), .ZN(new_n13557_));
  NOR2_X1    g12555(.A1(new_n13557_), .A2(new_n13315_), .ZN(new_n13558_));
  OR4_X2     g12556(.A1(new_n13537_), .A2(new_n13538_), .A3(new_n13541_), .A4(new_n13543_), .Z(new_n13559_));
  NAND3_X1   g12557(.A1(new_n13558_), .A2(new_n13544_), .A3(new_n13559_), .ZN(new_n13560_));
  INV_X1     g12558(.I(new_n13560_), .ZN(new_n13561_));
  NAND3_X1   g12559(.A1(new_n13554_), .A2(new_n13550_), .A3(new_n13561_), .ZN(new_n13562_));
  NOR3_X1    g12560(.A1(new_n13551_), .A2(new_n13553_), .A3(new_n13552_), .ZN(new_n13563_));
  AOI21_X1   g12561(.A1(new_n13546_), .A2(new_n13549_), .B(new_n13453_), .ZN(new_n13564_));
  OAI21_X1   g12562(.A1(new_n13563_), .A2(new_n13564_), .B(new_n13560_), .ZN(new_n13565_));
  NAND3_X1   g12563(.A1(new_n13349_), .A2(new_n13562_), .A3(new_n13565_), .ZN(new_n13566_));
  NOR3_X1    g12564(.A1(new_n13563_), .A2(new_n13564_), .A3(new_n13560_), .ZN(new_n13567_));
  AOI21_X1   g12565(.A1(new_n13554_), .A2(new_n13550_), .B(new_n13561_), .ZN(new_n13568_));
  OAI21_X1   g12566(.A1(new_n13568_), .A2(new_n13567_), .B(new_n13348_), .ZN(new_n13569_));
  NAND2_X1   g12567(.A1(new_n13566_), .A2(new_n13569_), .ZN(new_n13570_));
  INV_X1     g12568(.I(\A[649] ), .ZN(new_n13571_));
  INV_X1     g12569(.I(\A[650] ), .ZN(new_n13572_));
  NAND2_X1   g12570(.A1(new_n13572_), .A2(\A[651] ), .ZN(new_n13573_));
  INV_X1     g12571(.I(\A[651] ), .ZN(new_n13574_));
  NAND2_X1   g12572(.A1(new_n13574_), .A2(\A[650] ), .ZN(new_n13575_));
  AOI21_X1   g12573(.A1(new_n13573_), .A2(new_n13575_), .B(new_n13571_), .ZN(new_n13576_));
  NOR2_X1    g12574(.A1(\A[650] ), .A2(\A[651] ), .ZN(new_n13577_));
  INV_X1     g12575(.I(new_n13577_), .ZN(new_n13578_));
  NAND2_X1   g12576(.A1(\A[650] ), .A2(\A[651] ), .ZN(new_n13579_));
  AOI21_X1   g12577(.A1(new_n13578_), .A2(new_n13579_), .B(\A[649] ), .ZN(new_n13580_));
  NOR2_X1    g12578(.A1(new_n13580_), .A2(new_n13576_), .ZN(new_n13581_));
  INV_X1     g12579(.I(\A[652] ), .ZN(new_n13582_));
  INV_X1     g12580(.I(\A[653] ), .ZN(new_n13583_));
  NAND2_X1   g12581(.A1(new_n13583_), .A2(\A[654] ), .ZN(new_n13584_));
  INV_X1     g12582(.I(\A[654] ), .ZN(new_n13585_));
  NAND2_X1   g12583(.A1(new_n13585_), .A2(\A[653] ), .ZN(new_n13586_));
  AOI21_X1   g12584(.A1(new_n13584_), .A2(new_n13586_), .B(new_n13582_), .ZN(new_n13587_));
  NOR2_X1    g12585(.A1(\A[653] ), .A2(\A[654] ), .ZN(new_n13588_));
  INV_X1     g12586(.I(new_n13588_), .ZN(new_n13589_));
  NAND2_X1   g12587(.A1(\A[653] ), .A2(\A[654] ), .ZN(new_n13590_));
  AOI21_X1   g12588(.A1(new_n13589_), .A2(new_n13590_), .B(\A[652] ), .ZN(new_n13591_));
  NOR2_X1    g12589(.A1(new_n13591_), .A2(new_n13587_), .ZN(new_n13592_));
  NAND2_X1   g12590(.A1(new_n13581_), .A2(new_n13592_), .ZN(new_n13593_));
  NOR2_X1    g12591(.A1(new_n13574_), .A2(\A[650] ), .ZN(new_n13594_));
  NOR2_X1    g12592(.A1(new_n13572_), .A2(\A[651] ), .ZN(new_n13595_));
  OAI21_X1   g12593(.A1(new_n13594_), .A2(new_n13595_), .B(\A[649] ), .ZN(new_n13596_));
  INV_X1     g12594(.I(new_n13579_), .ZN(new_n13597_));
  OAI21_X1   g12595(.A1(new_n13597_), .A2(new_n13577_), .B(new_n13571_), .ZN(new_n13598_));
  NAND2_X1   g12596(.A1(new_n13596_), .A2(new_n13598_), .ZN(new_n13599_));
  NOR2_X1    g12597(.A1(new_n13585_), .A2(\A[653] ), .ZN(new_n13600_));
  NOR2_X1    g12598(.A1(new_n13583_), .A2(\A[654] ), .ZN(new_n13601_));
  OAI21_X1   g12599(.A1(new_n13600_), .A2(new_n13601_), .B(\A[652] ), .ZN(new_n13602_));
  INV_X1     g12600(.I(new_n13590_), .ZN(new_n13603_));
  OAI21_X1   g12601(.A1(new_n13603_), .A2(new_n13588_), .B(new_n13582_), .ZN(new_n13604_));
  NAND2_X1   g12602(.A1(new_n13602_), .A2(new_n13604_), .ZN(new_n13605_));
  NAND2_X1   g12603(.A1(new_n13599_), .A2(new_n13605_), .ZN(new_n13606_));
  NAND2_X1   g12604(.A1(new_n13593_), .A2(new_n13606_), .ZN(new_n13607_));
  INV_X1     g12605(.I(\A[645] ), .ZN(new_n13608_));
  NOR2_X1    g12606(.A1(new_n13608_), .A2(\A[644] ), .ZN(new_n13609_));
  INV_X1     g12607(.I(\A[644] ), .ZN(new_n13610_));
  NOR2_X1    g12608(.A1(new_n13610_), .A2(\A[645] ), .ZN(new_n13611_));
  OAI21_X1   g12609(.A1(new_n13609_), .A2(new_n13611_), .B(\A[643] ), .ZN(new_n13612_));
  INV_X1     g12610(.I(\A[643] ), .ZN(new_n13613_));
  NAND2_X1   g12611(.A1(\A[644] ), .A2(\A[645] ), .ZN(new_n13614_));
  INV_X1     g12612(.I(new_n13614_), .ZN(new_n13615_));
  NOR2_X1    g12613(.A1(\A[644] ), .A2(\A[645] ), .ZN(new_n13616_));
  OAI21_X1   g12614(.A1(new_n13615_), .A2(new_n13616_), .B(new_n13613_), .ZN(new_n13617_));
  NAND2_X1   g12615(.A1(new_n13612_), .A2(new_n13617_), .ZN(new_n13618_));
  INV_X1     g12616(.I(\A[648] ), .ZN(new_n13619_));
  NOR2_X1    g12617(.A1(new_n13619_), .A2(\A[647] ), .ZN(new_n13620_));
  INV_X1     g12618(.I(\A[647] ), .ZN(new_n13621_));
  NOR2_X1    g12619(.A1(new_n13621_), .A2(\A[648] ), .ZN(new_n13622_));
  OAI21_X1   g12620(.A1(new_n13620_), .A2(new_n13622_), .B(\A[646] ), .ZN(new_n13623_));
  INV_X1     g12621(.I(\A[646] ), .ZN(new_n13624_));
  NAND2_X1   g12622(.A1(\A[647] ), .A2(\A[648] ), .ZN(new_n13625_));
  INV_X1     g12623(.I(new_n13625_), .ZN(new_n13626_));
  NOR2_X1    g12624(.A1(\A[647] ), .A2(\A[648] ), .ZN(new_n13627_));
  OAI21_X1   g12625(.A1(new_n13626_), .A2(new_n13627_), .B(new_n13624_), .ZN(new_n13628_));
  NAND2_X1   g12626(.A1(new_n13623_), .A2(new_n13628_), .ZN(new_n13629_));
  NOR2_X1    g12627(.A1(new_n13618_), .A2(new_n13629_), .ZN(new_n13630_));
  NAND2_X1   g12628(.A1(new_n13610_), .A2(\A[645] ), .ZN(new_n13631_));
  NAND2_X1   g12629(.A1(new_n13608_), .A2(\A[644] ), .ZN(new_n13632_));
  AOI21_X1   g12630(.A1(new_n13631_), .A2(new_n13632_), .B(new_n13613_), .ZN(new_n13633_));
  INV_X1     g12631(.I(new_n13616_), .ZN(new_n13634_));
  AOI21_X1   g12632(.A1(new_n13634_), .A2(new_n13614_), .B(\A[643] ), .ZN(new_n13635_));
  NOR2_X1    g12633(.A1(new_n13635_), .A2(new_n13633_), .ZN(new_n13636_));
  NAND2_X1   g12634(.A1(new_n13621_), .A2(\A[648] ), .ZN(new_n13637_));
  NAND2_X1   g12635(.A1(new_n13619_), .A2(\A[647] ), .ZN(new_n13638_));
  AOI21_X1   g12636(.A1(new_n13637_), .A2(new_n13638_), .B(new_n13624_), .ZN(new_n13639_));
  INV_X1     g12637(.I(new_n13627_), .ZN(new_n13640_));
  AOI21_X1   g12638(.A1(new_n13640_), .A2(new_n13625_), .B(\A[646] ), .ZN(new_n13641_));
  NOR2_X1    g12639(.A1(new_n13641_), .A2(new_n13639_), .ZN(new_n13642_));
  NOR2_X1    g12640(.A1(new_n13636_), .A2(new_n13642_), .ZN(new_n13643_));
  NOR2_X1    g12641(.A1(new_n13643_), .A2(new_n13630_), .ZN(new_n13644_));
  NOR2_X1    g12642(.A1(new_n13644_), .A2(new_n13607_), .ZN(new_n13645_));
  NOR2_X1    g12643(.A1(new_n13599_), .A2(new_n13605_), .ZN(new_n13646_));
  NOR2_X1    g12644(.A1(new_n13581_), .A2(new_n13592_), .ZN(new_n13647_));
  NOR2_X1    g12645(.A1(new_n13647_), .A2(new_n13646_), .ZN(new_n13648_));
  NAND2_X1   g12646(.A1(new_n13636_), .A2(new_n13642_), .ZN(new_n13649_));
  NAND2_X1   g12647(.A1(new_n13618_), .A2(new_n13629_), .ZN(new_n13650_));
  NAND2_X1   g12648(.A1(new_n13649_), .A2(new_n13650_), .ZN(new_n13651_));
  NOR2_X1    g12649(.A1(new_n13648_), .A2(new_n13651_), .ZN(new_n13652_));
  NOR2_X1    g12650(.A1(new_n13645_), .A2(new_n13652_), .ZN(new_n13653_));
  INV_X1     g12651(.I(\A[637] ), .ZN(new_n13654_));
  INV_X1     g12652(.I(\A[638] ), .ZN(new_n13655_));
  NAND2_X1   g12653(.A1(new_n13655_), .A2(\A[639] ), .ZN(new_n13656_));
  INV_X1     g12654(.I(\A[639] ), .ZN(new_n13657_));
  NAND2_X1   g12655(.A1(new_n13657_), .A2(\A[638] ), .ZN(new_n13658_));
  AOI21_X1   g12656(.A1(new_n13656_), .A2(new_n13658_), .B(new_n13654_), .ZN(new_n13659_));
  NOR2_X1    g12657(.A1(\A[638] ), .A2(\A[639] ), .ZN(new_n13660_));
  INV_X1     g12658(.I(new_n13660_), .ZN(new_n13661_));
  NAND2_X1   g12659(.A1(\A[638] ), .A2(\A[639] ), .ZN(new_n13662_));
  AOI21_X1   g12660(.A1(new_n13661_), .A2(new_n13662_), .B(\A[637] ), .ZN(new_n13663_));
  NOR2_X1    g12661(.A1(new_n13663_), .A2(new_n13659_), .ZN(new_n13664_));
  INV_X1     g12662(.I(\A[640] ), .ZN(new_n13665_));
  INV_X1     g12663(.I(\A[641] ), .ZN(new_n13666_));
  NAND2_X1   g12664(.A1(new_n13666_), .A2(\A[642] ), .ZN(new_n13667_));
  INV_X1     g12665(.I(\A[642] ), .ZN(new_n13668_));
  NAND2_X1   g12666(.A1(new_n13668_), .A2(\A[641] ), .ZN(new_n13669_));
  AOI21_X1   g12667(.A1(new_n13667_), .A2(new_n13669_), .B(new_n13665_), .ZN(new_n13670_));
  NOR2_X1    g12668(.A1(\A[641] ), .A2(\A[642] ), .ZN(new_n13671_));
  INV_X1     g12669(.I(new_n13671_), .ZN(new_n13672_));
  NAND2_X1   g12670(.A1(\A[641] ), .A2(\A[642] ), .ZN(new_n13673_));
  AOI21_X1   g12671(.A1(new_n13672_), .A2(new_n13673_), .B(\A[640] ), .ZN(new_n13674_));
  NOR2_X1    g12672(.A1(new_n13674_), .A2(new_n13670_), .ZN(new_n13675_));
  NAND2_X1   g12673(.A1(new_n13664_), .A2(new_n13675_), .ZN(new_n13676_));
  NOR2_X1    g12674(.A1(new_n13657_), .A2(\A[638] ), .ZN(new_n13677_));
  NOR2_X1    g12675(.A1(new_n13655_), .A2(\A[639] ), .ZN(new_n13678_));
  OAI21_X1   g12676(.A1(new_n13677_), .A2(new_n13678_), .B(\A[637] ), .ZN(new_n13679_));
  INV_X1     g12677(.I(new_n13662_), .ZN(new_n13680_));
  OAI21_X1   g12678(.A1(new_n13680_), .A2(new_n13660_), .B(new_n13654_), .ZN(new_n13681_));
  NAND2_X1   g12679(.A1(new_n13679_), .A2(new_n13681_), .ZN(new_n13682_));
  NOR2_X1    g12680(.A1(new_n13668_), .A2(\A[641] ), .ZN(new_n13683_));
  NOR2_X1    g12681(.A1(new_n13666_), .A2(\A[642] ), .ZN(new_n13684_));
  OAI21_X1   g12682(.A1(new_n13683_), .A2(new_n13684_), .B(\A[640] ), .ZN(new_n13685_));
  INV_X1     g12683(.I(new_n13673_), .ZN(new_n13686_));
  OAI21_X1   g12684(.A1(new_n13686_), .A2(new_n13671_), .B(new_n13665_), .ZN(new_n13687_));
  NAND2_X1   g12685(.A1(new_n13685_), .A2(new_n13687_), .ZN(new_n13688_));
  NAND2_X1   g12686(.A1(new_n13682_), .A2(new_n13688_), .ZN(new_n13689_));
  NAND2_X1   g12687(.A1(new_n13676_), .A2(new_n13689_), .ZN(new_n13690_));
  INV_X1     g12688(.I(\A[631] ), .ZN(new_n13691_));
  INV_X1     g12689(.I(\A[632] ), .ZN(new_n13692_));
  NAND2_X1   g12690(.A1(new_n13692_), .A2(\A[633] ), .ZN(new_n13693_));
  INV_X1     g12691(.I(\A[633] ), .ZN(new_n13694_));
  NAND2_X1   g12692(.A1(new_n13694_), .A2(\A[632] ), .ZN(new_n13695_));
  AOI21_X1   g12693(.A1(new_n13693_), .A2(new_n13695_), .B(new_n13691_), .ZN(new_n13696_));
  NAND2_X1   g12694(.A1(\A[632] ), .A2(\A[633] ), .ZN(new_n13697_));
  NOR2_X1    g12695(.A1(\A[632] ), .A2(\A[633] ), .ZN(new_n13698_));
  INV_X1     g12696(.I(new_n13698_), .ZN(new_n13699_));
  AOI21_X1   g12697(.A1(new_n13699_), .A2(new_n13697_), .B(\A[631] ), .ZN(new_n13700_));
  INV_X1     g12698(.I(\A[634] ), .ZN(new_n13701_));
  INV_X1     g12699(.I(\A[635] ), .ZN(new_n13702_));
  NAND2_X1   g12700(.A1(new_n13702_), .A2(\A[636] ), .ZN(new_n13703_));
  INV_X1     g12701(.I(\A[636] ), .ZN(new_n13704_));
  NAND2_X1   g12702(.A1(new_n13704_), .A2(\A[635] ), .ZN(new_n13705_));
  AOI21_X1   g12703(.A1(new_n13703_), .A2(new_n13705_), .B(new_n13701_), .ZN(new_n13706_));
  NAND2_X1   g12704(.A1(\A[635] ), .A2(\A[636] ), .ZN(new_n13707_));
  NOR2_X1    g12705(.A1(\A[635] ), .A2(\A[636] ), .ZN(new_n13708_));
  INV_X1     g12706(.I(new_n13708_), .ZN(new_n13709_));
  AOI21_X1   g12707(.A1(new_n13709_), .A2(new_n13707_), .B(\A[634] ), .ZN(new_n13710_));
  NOR4_X1    g12708(.A1(new_n13696_), .A2(new_n13700_), .A3(new_n13710_), .A4(new_n13706_), .ZN(new_n13711_));
  OAI22_X1   g12709(.A1(new_n13696_), .A2(new_n13700_), .B1(new_n13710_), .B2(new_n13706_), .ZN(new_n13712_));
  INV_X1     g12710(.I(new_n13712_), .ZN(new_n13713_));
  NOR2_X1    g12711(.A1(new_n13713_), .A2(new_n13711_), .ZN(new_n13714_));
  NOR2_X1    g12712(.A1(new_n13714_), .A2(new_n13690_), .ZN(new_n13715_));
  NOR2_X1    g12713(.A1(new_n13682_), .A2(new_n13688_), .ZN(new_n13716_));
  NOR2_X1    g12714(.A1(new_n13664_), .A2(new_n13675_), .ZN(new_n13717_));
  NOR2_X1    g12715(.A1(new_n13717_), .A2(new_n13716_), .ZN(new_n13718_));
  NOR2_X1    g12716(.A1(new_n13700_), .A2(new_n13696_), .ZN(new_n13719_));
  NOR2_X1    g12717(.A1(new_n13710_), .A2(new_n13706_), .ZN(new_n13720_));
  NAND2_X1   g12718(.A1(new_n13719_), .A2(new_n13720_), .ZN(new_n13721_));
  NAND2_X1   g12719(.A1(new_n13721_), .A2(new_n13712_), .ZN(new_n13722_));
  NOR2_X1    g12720(.A1(new_n13718_), .A2(new_n13722_), .ZN(new_n13723_));
  NOR2_X1    g12721(.A1(new_n13715_), .A2(new_n13723_), .ZN(new_n13724_));
  NOR2_X1    g12722(.A1(new_n13653_), .A2(new_n13724_), .ZN(new_n13725_));
  NAND2_X1   g12723(.A1(new_n13653_), .A2(new_n13724_), .ZN(new_n13726_));
  INV_X1     g12724(.I(new_n13726_), .ZN(new_n13727_));
  INV_X1     g12725(.I(\A[627] ), .ZN(new_n13728_));
  NOR2_X1    g12726(.A1(new_n13728_), .A2(\A[626] ), .ZN(new_n13729_));
  INV_X1     g12727(.I(\A[626] ), .ZN(new_n13730_));
  NOR2_X1    g12728(.A1(new_n13730_), .A2(\A[627] ), .ZN(new_n13731_));
  OAI21_X1   g12729(.A1(new_n13729_), .A2(new_n13731_), .B(\A[625] ), .ZN(new_n13732_));
  INV_X1     g12730(.I(\A[625] ), .ZN(new_n13733_));
  NOR2_X1    g12731(.A1(\A[626] ), .A2(\A[627] ), .ZN(new_n13734_));
  NAND2_X1   g12732(.A1(\A[626] ), .A2(\A[627] ), .ZN(new_n13735_));
  INV_X1     g12733(.I(new_n13735_), .ZN(new_n13736_));
  OAI21_X1   g12734(.A1(new_n13736_), .A2(new_n13734_), .B(new_n13733_), .ZN(new_n13737_));
  NAND2_X1   g12735(.A1(new_n13732_), .A2(new_n13737_), .ZN(new_n13738_));
  INV_X1     g12736(.I(\A[630] ), .ZN(new_n13739_));
  NOR2_X1    g12737(.A1(new_n13739_), .A2(\A[629] ), .ZN(new_n13740_));
  INV_X1     g12738(.I(\A[629] ), .ZN(new_n13741_));
  NOR2_X1    g12739(.A1(new_n13741_), .A2(\A[630] ), .ZN(new_n13742_));
  OAI21_X1   g12740(.A1(new_n13740_), .A2(new_n13742_), .B(\A[628] ), .ZN(new_n13743_));
  INV_X1     g12741(.I(\A[628] ), .ZN(new_n13744_));
  NOR2_X1    g12742(.A1(\A[629] ), .A2(\A[630] ), .ZN(new_n13745_));
  NAND2_X1   g12743(.A1(\A[629] ), .A2(\A[630] ), .ZN(new_n13746_));
  INV_X1     g12744(.I(new_n13746_), .ZN(new_n13747_));
  OAI21_X1   g12745(.A1(new_n13747_), .A2(new_n13745_), .B(new_n13744_), .ZN(new_n13748_));
  NAND2_X1   g12746(.A1(new_n13743_), .A2(new_n13748_), .ZN(new_n13749_));
  NOR2_X1    g12747(.A1(new_n13738_), .A2(new_n13749_), .ZN(new_n13750_));
  NAND2_X1   g12748(.A1(new_n13730_), .A2(\A[627] ), .ZN(new_n13751_));
  NAND2_X1   g12749(.A1(new_n13728_), .A2(\A[626] ), .ZN(new_n13752_));
  AOI21_X1   g12750(.A1(new_n13751_), .A2(new_n13752_), .B(new_n13733_), .ZN(new_n13753_));
  INV_X1     g12751(.I(new_n13734_), .ZN(new_n13754_));
  AOI21_X1   g12752(.A1(new_n13754_), .A2(new_n13735_), .B(\A[625] ), .ZN(new_n13755_));
  NOR2_X1    g12753(.A1(new_n13755_), .A2(new_n13753_), .ZN(new_n13756_));
  NAND2_X1   g12754(.A1(new_n13741_), .A2(\A[630] ), .ZN(new_n13757_));
  NAND2_X1   g12755(.A1(new_n13739_), .A2(\A[629] ), .ZN(new_n13758_));
  AOI21_X1   g12756(.A1(new_n13757_), .A2(new_n13758_), .B(new_n13744_), .ZN(new_n13759_));
  INV_X1     g12757(.I(new_n13745_), .ZN(new_n13760_));
  AOI21_X1   g12758(.A1(new_n13760_), .A2(new_n13746_), .B(\A[628] ), .ZN(new_n13761_));
  NOR2_X1    g12759(.A1(new_n13761_), .A2(new_n13759_), .ZN(new_n13762_));
  NOR2_X1    g12760(.A1(new_n13756_), .A2(new_n13762_), .ZN(new_n13763_));
  NOR2_X1    g12761(.A1(new_n13763_), .A2(new_n13750_), .ZN(new_n13764_));
  INV_X1     g12762(.I(\A[621] ), .ZN(new_n13765_));
  NOR2_X1    g12763(.A1(new_n13765_), .A2(\A[620] ), .ZN(new_n13766_));
  INV_X1     g12764(.I(\A[620] ), .ZN(new_n13767_));
  NOR2_X1    g12765(.A1(new_n13767_), .A2(\A[621] ), .ZN(new_n13768_));
  OAI21_X1   g12766(.A1(new_n13766_), .A2(new_n13768_), .B(\A[619] ), .ZN(new_n13769_));
  INV_X1     g12767(.I(\A[619] ), .ZN(new_n13770_));
  NAND2_X1   g12768(.A1(\A[620] ), .A2(\A[621] ), .ZN(new_n13771_));
  INV_X1     g12769(.I(new_n13771_), .ZN(new_n13772_));
  NOR2_X1    g12770(.A1(\A[620] ), .A2(\A[621] ), .ZN(new_n13773_));
  OAI21_X1   g12771(.A1(new_n13772_), .A2(new_n13773_), .B(new_n13770_), .ZN(new_n13774_));
  INV_X1     g12772(.I(\A[624] ), .ZN(new_n13775_));
  NOR2_X1    g12773(.A1(new_n13775_), .A2(\A[623] ), .ZN(new_n13776_));
  INV_X1     g12774(.I(\A[623] ), .ZN(new_n13777_));
  NOR2_X1    g12775(.A1(new_n13777_), .A2(\A[624] ), .ZN(new_n13778_));
  OAI21_X1   g12776(.A1(new_n13776_), .A2(new_n13778_), .B(\A[622] ), .ZN(new_n13779_));
  INV_X1     g12777(.I(\A[622] ), .ZN(new_n13780_));
  NAND2_X1   g12778(.A1(\A[623] ), .A2(\A[624] ), .ZN(new_n13781_));
  INV_X1     g12779(.I(new_n13781_), .ZN(new_n13782_));
  NOR2_X1    g12780(.A1(\A[623] ), .A2(\A[624] ), .ZN(new_n13783_));
  OAI21_X1   g12781(.A1(new_n13782_), .A2(new_n13783_), .B(new_n13780_), .ZN(new_n13784_));
  NAND4_X1   g12782(.A1(new_n13769_), .A2(new_n13774_), .A3(new_n13779_), .A4(new_n13784_), .ZN(new_n13785_));
  NAND2_X1   g12783(.A1(new_n13769_), .A2(new_n13774_), .ZN(new_n13786_));
  NAND2_X1   g12784(.A1(new_n13779_), .A2(new_n13784_), .ZN(new_n13787_));
  NAND2_X1   g12785(.A1(new_n13786_), .A2(new_n13787_), .ZN(new_n13788_));
  NAND2_X1   g12786(.A1(new_n13788_), .A2(new_n13785_), .ZN(new_n13789_));
  NAND2_X1   g12787(.A1(new_n13764_), .A2(new_n13789_), .ZN(new_n13790_));
  NAND2_X1   g12788(.A1(new_n13756_), .A2(new_n13762_), .ZN(new_n13791_));
  NAND2_X1   g12789(.A1(new_n13738_), .A2(new_n13749_), .ZN(new_n13792_));
  NAND2_X1   g12790(.A1(new_n13791_), .A2(new_n13792_), .ZN(new_n13793_));
  INV_X1     g12791(.I(new_n13789_), .ZN(new_n13794_));
  NAND2_X1   g12792(.A1(new_n13794_), .A2(new_n13793_), .ZN(new_n13795_));
  INV_X1     g12793(.I(\A[615] ), .ZN(new_n13796_));
  NOR2_X1    g12794(.A1(new_n13796_), .A2(\A[614] ), .ZN(new_n13797_));
  INV_X1     g12795(.I(\A[614] ), .ZN(new_n13798_));
  NOR2_X1    g12796(.A1(new_n13798_), .A2(\A[615] ), .ZN(new_n13799_));
  OAI21_X1   g12797(.A1(new_n13797_), .A2(new_n13799_), .B(\A[613] ), .ZN(new_n13800_));
  INV_X1     g12798(.I(\A[613] ), .ZN(new_n13801_));
  NOR2_X1    g12799(.A1(\A[614] ), .A2(\A[615] ), .ZN(new_n13802_));
  NAND2_X1   g12800(.A1(\A[614] ), .A2(\A[615] ), .ZN(new_n13803_));
  INV_X1     g12801(.I(new_n13803_), .ZN(new_n13804_));
  OAI21_X1   g12802(.A1(new_n13804_), .A2(new_n13802_), .B(new_n13801_), .ZN(new_n13805_));
  NAND2_X1   g12803(.A1(new_n13800_), .A2(new_n13805_), .ZN(new_n13806_));
  INV_X1     g12804(.I(\A[618] ), .ZN(new_n13807_));
  NOR2_X1    g12805(.A1(new_n13807_), .A2(\A[617] ), .ZN(new_n13808_));
  INV_X1     g12806(.I(\A[617] ), .ZN(new_n13809_));
  NOR2_X1    g12807(.A1(new_n13809_), .A2(\A[618] ), .ZN(new_n13810_));
  OAI21_X1   g12808(.A1(new_n13808_), .A2(new_n13810_), .B(\A[616] ), .ZN(new_n13811_));
  INV_X1     g12809(.I(\A[616] ), .ZN(new_n13812_));
  NOR2_X1    g12810(.A1(\A[617] ), .A2(\A[618] ), .ZN(new_n13813_));
  NAND2_X1   g12811(.A1(\A[617] ), .A2(\A[618] ), .ZN(new_n13814_));
  INV_X1     g12812(.I(new_n13814_), .ZN(new_n13815_));
  OAI21_X1   g12813(.A1(new_n13815_), .A2(new_n13813_), .B(new_n13812_), .ZN(new_n13816_));
  NAND2_X1   g12814(.A1(new_n13811_), .A2(new_n13816_), .ZN(new_n13817_));
  NOR2_X1    g12815(.A1(new_n13806_), .A2(new_n13817_), .ZN(new_n13818_));
  NAND2_X1   g12816(.A1(new_n13798_), .A2(\A[615] ), .ZN(new_n13819_));
  NAND2_X1   g12817(.A1(new_n13796_), .A2(\A[614] ), .ZN(new_n13820_));
  AOI21_X1   g12818(.A1(new_n13819_), .A2(new_n13820_), .B(new_n13801_), .ZN(new_n13821_));
  INV_X1     g12819(.I(new_n13802_), .ZN(new_n13822_));
  AOI21_X1   g12820(.A1(new_n13822_), .A2(new_n13803_), .B(\A[613] ), .ZN(new_n13823_));
  NOR2_X1    g12821(.A1(new_n13823_), .A2(new_n13821_), .ZN(new_n13824_));
  NAND2_X1   g12822(.A1(new_n13809_), .A2(\A[618] ), .ZN(new_n13825_));
  NAND2_X1   g12823(.A1(new_n13807_), .A2(\A[617] ), .ZN(new_n13826_));
  AOI21_X1   g12824(.A1(new_n13825_), .A2(new_n13826_), .B(new_n13812_), .ZN(new_n13827_));
  INV_X1     g12825(.I(new_n13813_), .ZN(new_n13828_));
  AOI21_X1   g12826(.A1(new_n13828_), .A2(new_n13814_), .B(\A[616] ), .ZN(new_n13829_));
  NOR2_X1    g12827(.A1(new_n13829_), .A2(new_n13827_), .ZN(new_n13830_));
  NOR2_X1    g12828(.A1(new_n13824_), .A2(new_n13830_), .ZN(new_n13831_));
  NOR2_X1    g12829(.A1(new_n13831_), .A2(new_n13818_), .ZN(new_n13832_));
  INV_X1     g12830(.I(\A[607] ), .ZN(new_n13833_));
  INV_X1     g12831(.I(\A[608] ), .ZN(new_n13834_));
  NAND2_X1   g12832(.A1(new_n13834_), .A2(\A[609] ), .ZN(new_n13835_));
  INV_X1     g12833(.I(\A[609] ), .ZN(new_n13836_));
  NAND2_X1   g12834(.A1(new_n13836_), .A2(\A[608] ), .ZN(new_n13837_));
  AOI21_X1   g12835(.A1(new_n13835_), .A2(new_n13837_), .B(new_n13833_), .ZN(new_n13838_));
  NAND2_X1   g12836(.A1(\A[608] ), .A2(\A[609] ), .ZN(new_n13839_));
  NOR2_X1    g12837(.A1(\A[608] ), .A2(\A[609] ), .ZN(new_n13840_));
  INV_X1     g12838(.I(new_n13840_), .ZN(new_n13841_));
  AOI21_X1   g12839(.A1(new_n13841_), .A2(new_n13839_), .B(\A[607] ), .ZN(new_n13842_));
  INV_X1     g12840(.I(\A[610] ), .ZN(new_n13843_));
  INV_X1     g12841(.I(\A[611] ), .ZN(new_n13844_));
  NAND2_X1   g12842(.A1(new_n13844_), .A2(\A[612] ), .ZN(new_n13845_));
  INV_X1     g12843(.I(\A[612] ), .ZN(new_n13846_));
  NAND2_X1   g12844(.A1(new_n13846_), .A2(\A[611] ), .ZN(new_n13847_));
  AOI21_X1   g12845(.A1(new_n13845_), .A2(new_n13847_), .B(new_n13843_), .ZN(new_n13848_));
  NAND2_X1   g12846(.A1(\A[611] ), .A2(\A[612] ), .ZN(new_n13849_));
  NOR2_X1    g12847(.A1(\A[611] ), .A2(\A[612] ), .ZN(new_n13850_));
  INV_X1     g12848(.I(new_n13850_), .ZN(new_n13851_));
  AOI21_X1   g12849(.A1(new_n13851_), .A2(new_n13849_), .B(\A[610] ), .ZN(new_n13852_));
  NOR4_X1    g12850(.A1(new_n13838_), .A2(new_n13842_), .A3(new_n13852_), .A4(new_n13848_), .ZN(new_n13853_));
  INV_X1     g12851(.I(new_n13853_), .ZN(new_n13854_));
  OAI22_X1   g12852(.A1(new_n13838_), .A2(new_n13842_), .B1(new_n13852_), .B2(new_n13848_), .ZN(new_n13855_));
  NAND2_X1   g12853(.A1(new_n13854_), .A2(new_n13855_), .ZN(new_n13856_));
  NAND2_X1   g12854(.A1(new_n13856_), .A2(new_n13832_), .ZN(new_n13857_));
  NAND2_X1   g12855(.A1(new_n13824_), .A2(new_n13830_), .ZN(new_n13858_));
  NAND2_X1   g12856(.A1(new_n13806_), .A2(new_n13817_), .ZN(new_n13859_));
  NAND2_X1   g12857(.A1(new_n13858_), .A2(new_n13859_), .ZN(new_n13860_));
  INV_X1     g12858(.I(new_n13855_), .ZN(new_n13861_));
  NOR2_X1    g12859(.A1(new_n13861_), .A2(new_n13853_), .ZN(new_n13862_));
  NAND2_X1   g12860(.A1(new_n13862_), .A2(new_n13860_), .ZN(new_n13863_));
  AOI22_X1   g12861(.A1(new_n13795_), .A2(new_n13790_), .B1(new_n13857_), .B2(new_n13863_), .ZN(new_n13864_));
  NAND2_X1   g12862(.A1(new_n13795_), .A2(new_n13790_), .ZN(new_n13865_));
  NAND2_X1   g12863(.A1(new_n13857_), .A2(new_n13863_), .ZN(new_n13866_));
  NOR2_X1    g12864(.A1(new_n13865_), .A2(new_n13866_), .ZN(new_n13867_));
  NOR4_X1    g12865(.A1(new_n13867_), .A2(new_n13725_), .A3(new_n13727_), .A4(new_n13864_), .ZN(new_n13868_));
  NOR2_X1    g12866(.A1(new_n13727_), .A2(new_n13725_), .ZN(new_n13869_));
  NOR2_X1    g12867(.A1(new_n13867_), .A2(new_n13864_), .ZN(new_n13870_));
  NOR2_X1    g12868(.A1(new_n13869_), .A2(new_n13870_), .ZN(new_n13871_));
  NOR2_X1    g12869(.A1(new_n13871_), .A2(new_n13868_), .ZN(new_n13872_));
  AOI21_X1   g12870(.A1(new_n13544_), .A2(new_n13559_), .B(new_n13558_), .ZN(new_n13873_));
  NOR2_X1    g12871(.A1(new_n13561_), .A2(new_n13873_), .ZN(new_n13874_));
  NAND2_X1   g12872(.A1(new_n13874_), .A2(new_n13872_), .ZN(new_n13875_));
  INV_X1     g12873(.I(new_n13875_), .ZN(new_n13876_));
  AOI21_X1   g12874(.A1(\A[623] ), .A2(\A[624] ), .B(\A[622] ), .ZN(new_n13877_));
  AOI21_X1   g12875(.A1(\A[620] ), .A2(\A[621] ), .B(\A[619] ), .ZN(new_n13878_));
  OAI22_X1   g12876(.A1(new_n13773_), .A2(new_n13878_), .B1(new_n13877_), .B2(new_n13783_), .ZN(new_n13879_));
  NOR4_X1    g12877(.A1(new_n13877_), .A2(new_n13878_), .A3(new_n13773_), .A4(new_n13783_), .ZN(new_n13880_));
  INV_X1     g12878(.I(new_n13880_), .ZN(new_n13881_));
  NAND2_X1   g12879(.A1(new_n13881_), .A2(new_n13879_), .ZN(new_n13882_));
  XOR2_X1    g12880(.A1(new_n13785_), .A2(new_n13882_), .Z(new_n13883_));
  INV_X1     g12881(.I(new_n13883_), .ZN(new_n13884_));
  AOI21_X1   g12882(.A1(new_n13744_), .A2(new_n13746_), .B(new_n13745_), .ZN(new_n13885_));
  AOI21_X1   g12883(.A1(new_n13733_), .A2(new_n13735_), .B(new_n13734_), .ZN(new_n13886_));
  XNOR2_X1   g12884(.A1(new_n13885_), .A2(new_n13886_), .ZN(new_n13887_));
  XOR2_X1    g12885(.A1(new_n13750_), .A2(new_n13887_), .Z(new_n13888_));
  NOR2_X1    g12886(.A1(new_n13793_), .A2(new_n13789_), .ZN(new_n13889_));
  INV_X1     g12887(.I(new_n13889_), .ZN(new_n13890_));
  NAND2_X1   g12888(.A1(new_n13890_), .A2(new_n13888_), .ZN(new_n13891_));
  NOR4_X1    g12889(.A1(new_n13789_), .A2(new_n13750_), .A3(new_n13763_), .A4(new_n13887_), .ZN(new_n13892_));
  INV_X1     g12890(.I(new_n13892_), .ZN(new_n13893_));
  NAND3_X1   g12891(.A1(new_n13891_), .A2(new_n13893_), .A3(new_n13884_), .ZN(new_n13894_));
  XOR2_X1    g12892(.A1(new_n13791_), .A2(new_n13887_), .Z(new_n13895_));
  NOR2_X1    g12893(.A1(new_n13895_), .A2(new_n13889_), .ZN(new_n13896_));
  OAI21_X1   g12894(.A1(new_n13896_), .A2(new_n13892_), .B(new_n13883_), .ZN(new_n13897_));
  NAND2_X1   g12895(.A1(new_n13894_), .A2(new_n13897_), .ZN(new_n13898_));
  AOI21_X1   g12896(.A1(new_n13843_), .A2(new_n13849_), .B(new_n13850_), .ZN(new_n13899_));
  AOI21_X1   g12897(.A1(new_n13833_), .A2(new_n13839_), .B(new_n13840_), .ZN(new_n13900_));
  XOR2_X1    g12898(.A1(new_n13899_), .A2(new_n13900_), .Z(new_n13901_));
  XNOR2_X1   g12899(.A1(new_n13901_), .A2(new_n13853_), .ZN(new_n13902_));
  AOI21_X1   g12900(.A1(new_n13812_), .A2(new_n13814_), .B(new_n13813_), .ZN(new_n13903_));
  AOI21_X1   g12901(.A1(new_n13801_), .A2(new_n13803_), .B(new_n13802_), .ZN(new_n13904_));
  XOR2_X1    g12902(.A1(new_n13903_), .A2(new_n13904_), .Z(new_n13905_));
  XOR2_X1    g12903(.A1(new_n13858_), .A2(new_n13905_), .Z(new_n13906_));
  NAND2_X1   g12904(.A1(new_n13862_), .A2(new_n13832_), .ZN(new_n13907_));
  AOI21_X1   g12905(.A1(new_n13906_), .A2(new_n13907_), .B(new_n13902_), .ZN(new_n13908_));
  XOR2_X1    g12906(.A1(new_n13818_), .A2(new_n13905_), .Z(new_n13909_));
  NOR2_X1    g12907(.A1(new_n13856_), .A2(new_n13860_), .ZN(new_n13910_));
  NAND2_X1   g12908(.A1(new_n13909_), .A2(new_n13910_), .ZN(new_n13911_));
  NAND2_X1   g12909(.A1(new_n13908_), .A2(new_n13911_), .ZN(new_n13912_));
  NOR2_X1    g12910(.A1(new_n13909_), .A2(new_n13910_), .ZN(new_n13913_));
  NOR2_X1    g12911(.A1(new_n13906_), .A2(new_n13907_), .ZN(new_n13914_));
  OAI21_X1   g12912(.A1(new_n13914_), .A2(new_n13913_), .B(new_n13902_), .ZN(new_n13915_));
  NAND3_X1   g12913(.A1(new_n13912_), .A2(new_n13915_), .A3(new_n13864_), .ZN(new_n13916_));
  NAND2_X1   g12914(.A1(new_n13865_), .A2(new_n13866_), .ZN(new_n13917_));
  XOR2_X1    g12915(.A1(new_n13901_), .A2(new_n13853_), .Z(new_n13918_));
  OAI21_X1   g12916(.A1(new_n13909_), .A2(new_n13910_), .B(new_n13918_), .ZN(new_n13919_));
  NOR2_X1    g12917(.A1(new_n13919_), .A2(new_n13914_), .ZN(new_n13920_));
  NAND2_X1   g12918(.A1(new_n13906_), .A2(new_n13907_), .ZN(new_n13921_));
  AOI21_X1   g12919(.A1(new_n13921_), .A2(new_n13911_), .B(new_n13918_), .ZN(new_n13922_));
  OAI21_X1   g12920(.A1(new_n13922_), .A2(new_n13920_), .B(new_n13917_), .ZN(new_n13923_));
  NAND3_X1   g12921(.A1(new_n13923_), .A2(new_n13916_), .A3(new_n13898_), .ZN(new_n13924_));
  NOR3_X1    g12922(.A1(new_n13896_), .A2(new_n13883_), .A3(new_n13892_), .ZN(new_n13925_));
  AOI21_X1   g12923(.A1(new_n13891_), .A2(new_n13893_), .B(new_n13884_), .ZN(new_n13926_));
  NOR2_X1    g12924(.A1(new_n13926_), .A2(new_n13925_), .ZN(new_n13927_));
  NOR3_X1    g12925(.A1(new_n13922_), .A2(new_n13920_), .A3(new_n13917_), .ZN(new_n13928_));
  AOI21_X1   g12926(.A1(new_n13912_), .A2(new_n13915_), .B(new_n13864_), .ZN(new_n13929_));
  OAI21_X1   g12927(.A1(new_n13929_), .A2(new_n13928_), .B(new_n13927_), .ZN(new_n13930_));
  NAND2_X1   g12928(.A1(new_n13930_), .A2(new_n13924_), .ZN(new_n13931_));
  AOI21_X1   g12929(.A1(\A[635] ), .A2(\A[636] ), .B(\A[634] ), .ZN(new_n13932_));
  AOI21_X1   g12930(.A1(\A[632] ), .A2(\A[633] ), .B(\A[631] ), .ZN(new_n13933_));
  OAI22_X1   g12931(.A1(new_n13698_), .A2(new_n13933_), .B1(new_n13932_), .B2(new_n13708_), .ZN(new_n13934_));
  OR4_X2     g12932(.A1(new_n13698_), .A2(new_n13932_), .A3(new_n13933_), .A4(new_n13708_), .Z(new_n13935_));
  NAND2_X1   g12933(.A1(new_n13935_), .A2(new_n13934_), .ZN(new_n13936_));
  XNOR2_X1   g12934(.A1(new_n13711_), .A2(new_n13936_), .ZN(new_n13937_));
  AOI21_X1   g12935(.A1(new_n13665_), .A2(new_n13673_), .B(new_n13671_), .ZN(new_n13938_));
  AOI21_X1   g12936(.A1(\A[638] ), .A2(\A[639] ), .B(\A[637] ), .ZN(new_n13939_));
  NOR2_X1    g12937(.A1(new_n13939_), .A2(new_n13660_), .ZN(new_n13940_));
  XOR2_X1    g12938(.A1(new_n13938_), .A2(new_n13940_), .Z(new_n13941_));
  XOR2_X1    g12939(.A1(new_n13716_), .A2(new_n13941_), .Z(new_n13942_));
  NOR2_X1    g12940(.A1(new_n13690_), .A2(new_n13722_), .ZN(new_n13943_));
  OAI21_X1   g12941(.A1(new_n13942_), .A2(new_n13943_), .B(new_n13937_), .ZN(new_n13944_));
  XOR2_X1    g12942(.A1(new_n13676_), .A2(new_n13941_), .Z(new_n13945_));
  NAND2_X1   g12943(.A1(new_n13714_), .A2(new_n13718_), .ZN(new_n13946_));
  NOR2_X1    g12944(.A1(new_n13945_), .A2(new_n13946_), .ZN(new_n13947_));
  NOR2_X1    g12945(.A1(new_n13942_), .A2(new_n13943_), .ZN(new_n13948_));
  NOR2_X1    g12946(.A1(new_n13947_), .A2(new_n13948_), .ZN(new_n13949_));
  OAI22_X1   g12947(.A1(new_n13949_), .A2(new_n13937_), .B1(new_n13944_), .B2(new_n13947_), .ZN(new_n13950_));
  AOI21_X1   g12948(.A1(new_n13624_), .A2(new_n13625_), .B(new_n13627_), .ZN(new_n13951_));
  AOI21_X1   g12949(.A1(new_n13613_), .A2(new_n13614_), .B(new_n13616_), .ZN(new_n13952_));
  OR2_X2     g12950(.A1(new_n13951_), .A2(new_n13952_), .Z(new_n13953_));
  NAND2_X1   g12951(.A1(new_n13951_), .A2(new_n13952_), .ZN(new_n13954_));
  NAND2_X1   g12952(.A1(new_n13953_), .A2(new_n13954_), .ZN(new_n13955_));
  XOR2_X1    g12953(.A1(new_n13649_), .A2(new_n13955_), .Z(new_n13956_));
  AOI21_X1   g12954(.A1(new_n13582_), .A2(new_n13590_), .B(new_n13588_), .ZN(new_n13957_));
  AOI21_X1   g12955(.A1(new_n13571_), .A2(new_n13579_), .B(new_n13577_), .ZN(new_n13958_));
  XNOR2_X1   g12956(.A1(new_n13957_), .A2(new_n13958_), .ZN(new_n13959_));
  NAND2_X1   g12957(.A1(new_n13593_), .A2(new_n13959_), .ZN(new_n13960_));
  XOR2_X1    g12958(.A1(new_n13957_), .A2(new_n13958_), .Z(new_n13961_));
  NAND2_X1   g12959(.A1(new_n13646_), .A2(new_n13961_), .ZN(new_n13962_));
  AOI22_X1   g12960(.A1(new_n13644_), .A2(new_n13648_), .B1(new_n13960_), .B2(new_n13962_), .ZN(new_n13963_));
  NOR4_X1    g12961(.A1(new_n13651_), .A2(new_n13646_), .A3(new_n13647_), .A4(new_n13959_), .ZN(new_n13964_));
  NOR3_X1    g12962(.A1(new_n13963_), .A2(new_n13956_), .A3(new_n13964_), .ZN(new_n13965_));
  XOR2_X1    g12963(.A1(new_n13630_), .A2(new_n13955_), .Z(new_n13966_));
  NOR2_X1    g12964(.A1(new_n13646_), .A2(new_n13961_), .ZN(new_n13967_));
  NOR2_X1    g12965(.A1(new_n13593_), .A2(new_n13959_), .ZN(new_n13968_));
  OAI22_X1   g12966(.A1(new_n13607_), .A2(new_n13651_), .B1(new_n13968_), .B2(new_n13967_), .ZN(new_n13969_));
  NAND4_X1   g12967(.A1(new_n13644_), .A2(new_n13593_), .A3(new_n13606_), .A4(new_n13961_), .ZN(new_n13970_));
  AOI21_X1   g12968(.A1(new_n13969_), .A2(new_n13970_), .B(new_n13966_), .ZN(new_n13971_));
  OAI21_X1   g12969(.A1(new_n13965_), .A2(new_n13971_), .B(new_n13725_), .ZN(new_n13972_));
  XOR2_X1    g12970(.A1(new_n13607_), .A2(new_n13651_), .Z(new_n13973_));
  XOR2_X1    g12971(.A1(new_n13690_), .A2(new_n13722_), .Z(new_n13974_));
  NAND2_X1   g12972(.A1(new_n13973_), .A2(new_n13974_), .ZN(new_n13975_));
  NAND3_X1   g12973(.A1(new_n13969_), .A2(new_n13966_), .A3(new_n13970_), .ZN(new_n13976_));
  OAI21_X1   g12974(.A1(new_n13963_), .A2(new_n13964_), .B(new_n13956_), .ZN(new_n13977_));
  NAND3_X1   g12975(.A1(new_n13975_), .A2(new_n13977_), .A3(new_n13976_), .ZN(new_n13978_));
  AOI21_X1   g12976(.A1(new_n13972_), .A2(new_n13978_), .B(new_n13950_), .ZN(new_n13979_));
  XOR2_X1    g12977(.A1(new_n13711_), .A2(new_n13936_), .Z(new_n13980_));
  AOI21_X1   g12978(.A1(new_n13945_), .A2(new_n13946_), .B(new_n13980_), .ZN(new_n13981_));
  NAND2_X1   g12979(.A1(new_n13942_), .A2(new_n13943_), .ZN(new_n13982_));
  NAND2_X1   g12980(.A1(new_n13945_), .A2(new_n13946_), .ZN(new_n13983_));
  NAND2_X1   g12981(.A1(new_n13983_), .A2(new_n13982_), .ZN(new_n13984_));
  AOI22_X1   g12982(.A1(new_n13984_), .A2(new_n13980_), .B1(new_n13981_), .B2(new_n13982_), .ZN(new_n13985_));
  AOI21_X1   g12983(.A1(new_n13976_), .A2(new_n13977_), .B(new_n13975_), .ZN(new_n13986_));
  NOR3_X1    g12984(.A1(new_n13725_), .A2(new_n13971_), .A3(new_n13965_), .ZN(new_n13987_));
  NOR3_X1    g12985(.A1(new_n13986_), .A2(new_n13985_), .A3(new_n13987_), .ZN(new_n13988_));
  OAI21_X1   g12986(.A1(new_n13979_), .A2(new_n13988_), .B(new_n13868_), .ZN(new_n13989_));
  NAND2_X1   g12987(.A1(new_n13869_), .A2(new_n13870_), .ZN(new_n13990_));
  OAI21_X1   g12988(.A1(new_n13986_), .A2(new_n13987_), .B(new_n13985_), .ZN(new_n13991_));
  NAND3_X1   g12989(.A1(new_n13950_), .A2(new_n13972_), .A3(new_n13978_), .ZN(new_n13992_));
  NAND3_X1   g12990(.A1(new_n13991_), .A2(new_n13992_), .A3(new_n13990_), .ZN(new_n13993_));
  AOI21_X1   g12991(.A1(new_n13989_), .A2(new_n13993_), .B(new_n13931_), .ZN(new_n13994_));
  NAND3_X1   g12992(.A1(new_n13989_), .A2(new_n13993_), .A3(new_n13931_), .ZN(new_n13995_));
  INV_X1     g12993(.I(new_n13995_), .ZN(new_n13996_));
  OAI21_X1   g12994(.A1(new_n13996_), .A2(new_n13994_), .B(new_n13876_), .ZN(new_n13997_));
  NOR3_X1    g12995(.A1(new_n13996_), .A2(new_n13876_), .A3(new_n13994_), .ZN(new_n13998_));
  AOI21_X1   g12996(.A1(new_n13997_), .A2(new_n13570_), .B(new_n13998_), .ZN(new_n13999_));
  AOI21_X1   g12997(.A1(new_n13406_), .A2(new_n13436_), .B(new_n13379_), .ZN(new_n14000_));
  NAND2_X1   g12998(.A1(new_n13403_), .A2(new_n13404_), .ZN(new_n14001_));
  NOR2_X1    g12999(.A1(new_n13403_), .A2(new_n13404_), .ZN(new_n14002_));
  AOI21_X1   g13000(.A1(new_n13446_), .A2(new_n14001_), .B(new_n14002_), .ZN(new_n14003_));
  AOI21_X1   g13001(.A1(new_n13372_), .A2(new_n13376_), .B(new_n13375_), .ZN(new_n14004_));
  NOR2_X1    g13002(.A1(new_n14003_), .A2(new_n14004_), .ZN(new_n14005_));
  AND2_X2    g13003(.A1(new_n14003_), .A2(new_n14004_), .Z(new_n14006_));
  NOR2_X1    g13004(.A1(new_n14006_), .A2(new_n14005_), .ZN(new_n14007_));
  OAI21_X1   g13005(.A1(new_n14000_), .A2(new_n13440_), .B(new_n14007_), .ZN(new_n14008_));
  OAI21_X1   g13006(.A1(new_n13447_), .A2(new_n13450_), .B(new_n13445_), .ZN(new_n14009_));
  INV_X1     g13007(.I(new_n14005_), .ZN(new_n14010_));
  NAND2_X1   g13008(.A1(new_n14003_), .A2(new_n14004_), .ZN(new_n14011_));
  NAND2_X1   g13009(.A1(new_n14010_), .A2(new_n14011_), .ZN(new_n14012_));
  NAND3_X1   g13010(.A1(new_n14012_), .A2(new_n14009_), .A3(new_n13441_), .ZN(new_n14013_));
  NAND2_X1   g13011(.A1(new_n14008_), .A2(new_n14013_), .ZN(new_n14014_));
  AND2_X2    g13012(.A1(new_n13505_), .A2(new_n13506_), .Z(new_n14015_));
  NOR2_X1    g13013(.A1(new_n13505_), .A2(new_n13506_), .ZN(new_n14016_));
  INV_X1     g13014(.I(new_n14016_), .ZN(new_n14017_));
  OAI21_X1   g13015(.A1(new_n13504_), .A2(new_n14015_), .B(new_n14017_), .ZN(new_n14018_));
  NOR2_X1    g13016(.A1(new_n13523_), .A2(new_n13508_), .ZN(new_n14019_));
  INV_X1     g13017(.I(new_n14019_), .ZN(new_n14020_));
  NAND2_X1   g13018(.A1(new_n13540_), .A2(new_n13542_), .ZN(new_n14021_));
  AOI21_X1   g13019(.A1(new_n14020_), .A2(new_n14021_), .B(new_n13534_), .ZN(new_n14022_));
  AOI21_X1   g13020(.A1(new_n13526_), .A2(new_n13478_), .B(new_n13477_), .ZN(new_n14023_));
  NOR3_X1    g13021(.A1(new_n14022_), .A2(new_n13531_), .A3(new_n14023_), .ZN(new_n14024_));
  AOI21_X1   g13022(.A1(new_n13529_), .A2(new_n13481_), .B(new_n13531_), .ZN(new_n14025_));
  INV_X1     g13023(.I(new_n14023_), .ZN(new_n14026_));
  NOR2_X1    g13024(.A1(new_n14025_), .A2(new_n14026_), .ZN(new_n14027_));
  NOR3_X1    g13025(.A1(new_n14024_), .A2(new_n14027_), .A3(new_n14018_), .ZN(new_n14028_));
  INV_X1     g13026(.I(new_n14018_), .ZN(new_n14029_));
  NAND2_X1   g13027(.A1(new_n14025_), .A2(new_n14026_), .ZN(new_n14030_));
  OAI21_X1   g13028(.A1(new_n14022_), .A2(new_n13531_), .B(new_n14023_), .ZN(new_n14031_));
  AOI21_X1   g13029(.A1(new_n14031_), .A2(new_n14030_), .B(new_n14029_), .ZN(new_n14032_));
  OAI21_X1   g13030(.A1(new_n14028_), .A2(new_n14032_), .B(new_n14014_), .ZN(new_n14033_));
  AOI21_X1   g13031(.A1(new_n14009_), .A2(new_n13441_), .B(new_n14012_), .ZN(new_n14034_));
  NOR3_X1    g13032(.A1(new_n14000_), .A2(new_n14007_), .A3(new_n13440_), .ZN(new_n14035_));
  NOR2_X1    g13033(.A1(new_n14034_), .A2(new_n14035_), .ZN(new_n14036_));
  NAND3_X1   g13034(.A1(new_n14031_), .A2(new_n14030_), .A3(new_n14029_), .ZN(new_n14037_));
  OAI21_X1   g13035(.A1(new_n14024_), .A2(new_n14027_), .B(new_n14018_), .ZN(new_n14038_));
  NAND3_X1   g13036(.A1(new_n14036_), .A2(new_n14038_), .A3(new_n14037_), .ZN(new_n14039_));
  OAI21_X1   g13037(.A1(new_n13453_), .A2(new_n13552_), .B(new_n13549_), .ZN(new_n14040_));
  NAND3_X1   g13038(.A1(new_n14039_), .A2(new_n14033_), .A3(new_n14040_), .ZN(new_n14041_));
  AOI21_X1   g13039(.A1(new_n14037_), .A2(new_n14038_), .B(new_n14036_), .ZN(new_n14042_));
  NOR3_X1    g13040(.A1(new_n14028_), .A2(new_n14032_), .A3(new_n14014_), .ZN(new_n14043_));
  AOI21_X1   g13041(.A1(new_n13551_), .A2(new_n13546_), .B(new_n13553_), .ZN(new_n14044_));
  OAI21_X1   g13042(.A1(new_n14042_), .A2(new_n14043_), .B(new_n14044_), .ZN(new_n14045_));
  OAI21_X1   g13043(.A1(new_n13335_), .A2(new_n13230_), .B(new_n13346_), .ZN(new_n14046_));
  INV_X1     g13044(.I(new_n13331_), .ZN(new_n14047_));
  OR2_X2     g13045(.A1(new_n13329_), .A2(new_n13327_), .Z(new_n14048_));
  NAND2_X1   g13046(.A1(new_n13311_), .A2(new_n13267_), .ZN(new_n14049_));
  AOI21_X1   g13047(.A1(new_n14048_), .A2(new_n14049_), .B(new_n13323_), .ZN(new_n14050_));
  INV_X1     g13048(.I(new_n13324_), .ZN(new_n14051_));
  INV_X1     g13049(.I(new_n13325_), .ZN(new_n14052_));
  NOR2_X1    g13050(.A1(new_n14051_), .A2(new_n14052_), .ZN(new_n14053_));
  INV_X1     g13051(.I(new_n14053_), .ZN(new_n14054_));
  NOR2_X1    g13052(.A1(new_n13324_), .A2(new_n13325_), .ZN(new_n14055_));
  AOI21_X1   g13053(.A1(new_n13306_), .A2(new_n14054_), .B(new_n14055_), .ZN(new_n14056_));
  INV_X1     g13054(.I(new_n13319_), .ZN(new_n14057_));
  AOI21_X1   g13055(.A1(new_n13290_), .A2(new_n13321_), .B(new_n14057_), .ZN(new_n14058_));
  NOR2_X1    g13056(.A1(new_n14056_), .A2(new_n14058_), .ZN(new_n14059_));
  INV_X1     g13057(.I(new_n14055_), .ZN(new_n14060_));
  OAI21_X1   g13058(.A1(new_n13253_), .A2(new_n14053_), .B(new_n14060_), .ZN(new_n14061_));
  OAI21_X1   g13059(.A1(new_n13309_), .A2(new_n13320_), .B(new_n13319_), .ZN(new_n14062_));
  NOR2_X1    g13060(.A1(new_n14061_), .A2(new_n14062_), .ZN(new_n14063_));
  NOR2_X1    g13061(.A1(new_n14059_), .A2(new_n14063_), .ZN(new_n14064_));
  OAI21_X1   g13062(.A1(new_n14050_), .A2(new_n14047_), .B(new_n14064_), .ZN(new_n14065_));
  XOR2_X1    g13063(.A1(new_n13290_), .A2(new_n13322_), .Z(new_n14066_));
  NAND2_X1   g13064(.A1(new_n13330_), .A2(new_n14066_), .ZN(new_n14067_));
  NAND2_X1   g13065(.A1(new_n14061_), .A2(new_n14062_), .ZN(new_n14068_));
  NAND2_X1   g13066(.A1(new_n14056_), .A2(new_n14058_), .ZN(new_n14069_));
  NAND2_X1   g13067(.A1(new_n14069_), .A2(new_n14068_), .ZN(new_n14070_));
  NAND3_X1   g13068(.A1(new_n14067_), .A2(new_n14070_), .A3(new_n13331_), .ZN(new_n14071_));
  NAND2_X1   g13069(.A1(new_n14065_), .A2(new_n14071_), .ZN(new_n14072_));
  NOR4_X1    g13070(.A1(new_n13208_), .A2(new_n13210_), .A3(new_n13195_), .A4(new_n13204_), .ZN(new_n14073_));
  INV_X1     g13071(.I(new_n14073_), .ZN(new_n14074_));
  NOR2_X1    g13072(.A1(new_n13209_), .A2(new_n13211_), .ZN(new_n14075_));
  AOI21_X1   g13073(.A1(new_n13207_), .A2(new_n14074_), .B(new_n14075_), .ZN(new_n14076_));
  INV_X1     g13074(.I(new_n14076_), .ZN(new_n14077_));
  AOI21_X1   g13075(.A1(new_n13224_), .A2(new_n13186_), .B(new_n13184_), .ZN(new_n14078_));
  NOR3_X1    g13076(.A1(new_n13221_), .A2(new_n13341_), .A3(new_n14078_), .ZN(new_n14079_));
  INV_X1     g13077(.I(new_n14078_), .ZN(new_n14080_));
  AOI21_X1   g13078(.A1(new_n13340_), .A2(new_n13227_), .B(new_n14080_), .ZN(new_n14081_));
  NOR3_X1    g13079(.A1(new_n14081_), .A2(new_n14079_), .A3(new_n14077_), .ZN(new_n14082_));
  NAND3_X1   g13080(.A1(new_n13340_), .A2(new_n13227_), .A3(new_n14080_), .ZN(new_n14083_));
  OAI21_X1   g13081(.A1(new_n13221_), .A2(new_n13341_), .B(new_n14078_), .ZN(new_n14084_));
  AOI21_X1   g13082(.A1(new_n14083_), .A2(new_n14084_), .B(new_n14076_), .ZN(new_n14085_));
  OAI21_X1   g13083(.A1(new_n14085_), .A2(new_n14082_), .B(new_n14072_), .ZN(new_n14086_));
  AOI21_X1   g13084(.A1(new_n14067_), .A2(new_n13331_), .B(new_n14070_), .ZN(new_n14087_));
  NOR3_X1    g13085(.A1(new_n14050_), .A2(new_n14047_), .A3(new_n14064_), .ZN(new_n14088_));
  NOR2_X1    g13086(.A1(new_n14088_), .A2(new_n14087_), .ZN(new_n14089_));
  NAND3_X1   g13087(.A1(new_n14083_), .A2(new_n14084_), .A3(new_n14076_), .ZN(new_n14090_));
  OAI21_X1   g13088(.A1(new_n14081_), .A2(new_n14079_), .B(new_n14077_), .ZN(new_n14091_));
  NAND3_X1   g13089(.A1(new_n14091_), .A2(new_n14090_), .A3(new_n14089_), .ZN(new_n14092_));
  NAND3_X1   g13090(.A1(new_n14086_), .A2(new_n14092_), .A3(new_n14046_), .ZN(new_n14093_));
  AOI21_X1   g13091(.A1(new_n13344_), .A2(new_n13345_), .B(new_n13337_), .ZN(new_n14094_));
  AOI21_X1   g13092(.A1(new_n14091_), .A2(new_n14090_), .B(new_n14089_), .ZN(new_n14095_));
  NOR3_X1    g13093(.A1(new_n14085_), .A2(new_n14082_), .A3(new_n14072_), .ZN(new_n14096_));
  OAI21_X1   g13094(.A1(new_n14096_), .A2(new_n14095_), .B(new_n14094_), .ZN(new_n14097_));
  NAND4_X1   g13095(.A1(new_n14045_), .A2(new_n14041_), .A3(new_n14097_), .A4(new_n14093_), .ZN(new_n14098_));
  NOR3_X1    g13096(.A1(new_n14042_), .A2(new_n14043_), .A3(new_n14044_), .ZN(new_n14099_));
  AOI21_X1   g13097(.A1(new_n14039_), .A2(new_n14033_), .B(new_n14040_), .ZN(new_n14100_));
  NOR3_X1    g13098(.A1(new_n14096_), .A2(new_n14095_), .A3(new_n14094_), .ZN(new_n14101_));
  AOI21_X1   g13099(.A1(new_n14086_), .A2(new_n14092_), .B(new_n14046_), .ZN(new_n14102_));
  OAI22_X1   g13100(.A1(new_n14100_), .A2(new_n14099_), .B1(new_n14101_), .B2(new_n14102_), .ZN(new_n14103_));
  OAI21_X1   g13101(.A1(new_n13349_), .A2(new_n13567_), .B(new_n13565_), .ZN(new_n14104_));
  NAND3_X1   g13102(.A1(new_n14103_), .A2(new_n14098_), .A3(new_n14104_), .ZN(new_n14105_));
  NOR4_X1    g13103(.A1(new_n14100_), .A2(new_n14099_), .A3(new_n14101_), .A4(new_n14102_), .ZN(new_n14106_));
  AOI22_X1   g13104(.A1(new_n14045_), .A2(new_n14041_), .B1(new_n14097_), .B2(new_n14093_), .ZN(new_n14107_));
  AOI21_X1   g13105(.A1(new_n13348_), .A2(new_n13562_), .B(new_n13568_), .ZN(new_n14108_));
  OAI21_X1   g13106(.A1(new_n14106_), .A2(new_n14107_), .B(new_n14108_), .ZN(new_n14109_));
  AND2_X2    g13107(.A1(new_n13930_), .A2(new_n13924_), .Z(new_n14110_));
  AOI21_X1   g13108(.A1(new_n13991_), .A2(new_n13992_), .B(new_n13990_), .ZN(new_n14111_));
  OAI21_X1   g13109(.A1(new_n14110_), .A2(new_n14111_), .B(new_n13993_), .ZN(new_n14112_));
  AOI21_X1   g13110(.A1(new_n13890_), .A2(new_n13888_), .B(new_n13884_), .ZN(new_n14113_));
  INV_X1     g13111(.I(new_n13885_), .ZN(new_n14114_));
  INV_X1     g13112(.I(new_n13886_), .ZN(new_n14115_));
  NOR2_X1    g13113(.A1(new_n14114_), .A2(new_n14115_), .ZN(new_n14116_));
  INV_X1     g13114(.I(new_n14116_), .ZN(new_n14117_));
  NOR2_X1    g13115(.A1(new_n13885_), .A2(new_n13886_), .ZN(new_n14118_));
  AOI21_X1   g13116(.A1(new_n13791_), .A2(new_n14117_), .B(new_n14118_), .ZN(new_n14119_));
  INV_X1     g13117(.I(new_n13879_), .ZN(new_n14120_));
  AOI21_X1   g13118(.A1(new_n13785_), .A2(new_n13881_), .B(new_n14120_), .ZN(new_n14121_));
  NOR2_X1    g13119(.A1(new_n14119_), .A2(new_n14121_), .ZN(new_n14122_));
  INV_X1     g13120(.I(new_n14118_), .ZN(new_n14123_));
  OAI21_X1   g13121(.A1(new_n13750_), .A2(new_n14116_), .B(new_n14123_), .ZN(new_n14124_));
  INV_X1     g13122(.I(new_n14121_), .ZN(new_n14125_));
  NOR2_X1    g13123(.A1(new_n14125_), .A2(new_n14124_), .ZN(new_n14126_));
  NOR2_X1    g13124(.A1(new_n14126_), .A2(new_n14122_), .ZN(new_n14127_));
  OAI21_X1   g13125(.A1(new_n14113_), .A2(new_n13892_), .B(new_n14127_), .ZN(new_n14128_));
  OAI21_X1   g13126(.A1(new_n13895_), .A2(new_n13889_), .B(new_n13883_), .ZN(new_n14129_));
  NAND2_X1   g13127(.A1(new_n14125_), .A2(new_n14124_), .ZN(new_n14130_));
  NAND2_X1   g13128(.A1(new_n14119_), .A2(new_n14121_), .ZN(new_n14131_));
  NAND2_X1   g13129(.A1(new_n14130_), .A2(new_n14131_), .ZN(new_n14132_));
  NAND3_X1   g13130(.A1(new_n14129_), .A2(new_n13893_), .A3(new_n14132_), .ZN(new_n14133_));
  NAND2_X1   g13131(.A1(new_n14128_), .A2(new_n14133_), .ZN(new_n14134_));
  AND2_X2    g13132(.A1(new_n13903_), .A2(new_n13904_), .Z(new_n14135_));
  NOR2_X1    g13133(.A1(new_n13903_), .A2(new_n13904_), .ZN(new_n14136_));
  INV_X1     g13134(.I(new_n14136_), .ZN(new_n14137_));
  OAI21_X1   g13135(.A1(new_n13818_), .A2(new_n14135_), .B(new_n14137_), .ZN(new_n14138_));
  NOR2_X1    g13136(.A1(new_n13899_), .A2(new_n13900_), .ZN(new_n14139_));
  NAND2_X1   g13137(.A1(new_n13899_), .A2(new_n13900_), .ZN(new_n14140_));
  AOI21_X1   g13138(.A1(new_n13854_), .A2(new_n14140_), .B(new_n14139_), .ZN(new_n14141_));
  NOR3_X1    g13139(.A1(new_n13908_), .A2(new_n13914_), .A3(new_n14141_), .ZN(new_n14142_));
  INV_X1     g13140(.I(new_n14141_), .ZN(new_n14143_));
  AOI21_X1   g13141(.A1(new_n13919_), .A2(new_n13911_), .B(new_n14143_), .ZN(new_n14144_));
  NOR3_X1    g13142(.A1(new_n14142_), .A2(new_n14144_), .A3(new_n14138_), .ZN(new_n14145_));
  INV_X1     g13143(.I(new_n14138_), .ZN(new_n14146_));
  NAND3_X1   g13144(.A1(new_n13919_), .A2(new_n13911_), .A3(new_n14143_), .ZN(new_n14147_));
  OAI21_X1   g13145(.A1(new_n13908_), .A2(new_n13914_), .B(new_n14141_), .ZN(new_n14148_));
  AOI21_X1   g13146(.A1(new_n14148_), .A2(new_n14147_), .B(new_n14146_), .ZN(new_n14149_));
  OAI21_X1   g13147(.A1(new_n14145_), .A2(new_n14149_), .B(new_n14134_), .ZN(new_n14150_));
  AOI21_X1   g13148(.A1(new_n14129_), .A2(new_n13893_), .B(new_n14132_), .ZN(new_n14151_));
  NOR3_X1    g13149(.A1(new_n14113_), .A2(new_n13892_), .A3(new_n14127_), .ZN(new_n14152_));
  NOR2_X1    g13150(.A1(new_n14152_), .A2(new_n14151_), .ZN(new_n14153_));
  NAND3_X1   g13151(.A1(new_n14148_), .A2(new_n14147_), .A3(new_n14146_), .ZN(new_n14154_));
  OAI21_X1   g13152(.A1(new_n14142_), .A2(new_n14144_), .B(new_n14138_), .ZN(new_n14155_));
  NAND3_X1   g13153(.A1(new_n14153_), .A2(new_n14155_), .A3(new_n14154_), .ZN(new_n14156_));
  OAI21_X1   g13154(.A1(new_n13898_), .A2(new_n13928_), .B(new_n13923_), .ZN(new_n14157_));
  NAND3_X1   g13155(.A1(new_n14150_), .A2(new_n14156_), .A3(new_n14157_), .ZN(new_n14158_));
  AOI21_X1   g13156(.A1(new_n14154_), .A2(new_n14155_), .B(new_n14153_), .ZN(new_n14159_));
  NOR3_X1    g13157(.A1(new_n14134_), .A2(new_n14145_), .A3(new_n14149_), .ZN(new_n14160_));
  AOI21_X1   g13158(.A1(new_n13927_), .A2(new_n13916_), .B(new_n13929_), .ZN(new_n14161_));
  OAI21_X1   g13159(.A1(new_n14159_), .A2(new_n14160_), .B(new_n14161_), .ZN(new_n14162_));
  OAI21_X1   g13160(.A1(new_n13986_), .A2(new_n13985_), .B(new_n13978_), .ZN(new_n14163_));
  NOR2_X1    g13161(.A1(new_n13963_), .A2(new_n13966_), .ZN(new_n14164_));
  INV_X1     g13162(.I(new_n13957_), .ZN(new_n14165_));
  INV_X1     g13163(.I(new_n13958_), .ZN(new_n14166_));
  NOR2_X1    g13164(.A1(new_n14165_), .A2(new_n14166_), .ZN(new_n14167_));
  INV_X1     g13165(.I(new_n14167_), .ZN(new_n14168_));
  NOR2_X1    g13166(.A1(new_n13957_), .A2(new_n13958_), .ZN(new_n14169_));
  AOI21_X1   g13167(.A1(new_n13593_), .A2(new_n14168_), .B(new_n14169_), .ZN(new_n14170_));
  INV_X1     g13168(.I(new_n13953_), .ZN(new_n14171_));
  AOI21_X1   g13169(.A1(new_n13649_), .A2(new_n13954_), .B(new_n14171_), .ZN(new_n14172_));
  NOR2_X1    g13170(.A1(new_n14170_), .A2(new_n14172_), .ZN(new_n14173_));
  INV_X1     g13171(.I(new_n14169_), .ZN(new_n14174_));
  OAI21_X1   g13172(.A1(new_n13646_), .A2(new_n14167_), .B(new_n14174_), .ZN(new_n14175_));
  INV_X1     g13173(.I(new_n13954_), .ZN(new_n14176_));
  OAI21_X1   g13174(.A1(new_n13630_), .A2(new_n14176_), .B(new_n13953_), .ZN(new_n14177_));
  NOR2_X1    g13175(.A1(new_n14175_), .A2(new_n14177_), .ZN(new_n14178_));
  NOR2_X1    g13176(.A1(new_n14173_), .A2(new_n14178_), .ZN(new_n14179_));
  OAI21_X1   g13177(.A1(new_n14164_), .A2(new_n13964_), .B(new_n14179_), .ZN(new_n14180_));
  NAND2_X1   g13178(.A1(new_n13969_), .A2(new_n13956_), .ZN(new_n14181_));
  NAND2_X1   g13179(.A1(new_n14175_), .A2(new_n14177_), .ZN(new_n14182_));
  NAND2_X1   g13180(.A1(new_n14170_), .A2(new_n14172_), .ZN(new_n14183_));
  NAND2_X1   g13181(.A1(new_n14183_), .A2(new_n14182_), .ZN(new_n14184_));
  NAND3_X1   g13182(.A1(new_n14181_), .A2(new_n14184_), .A3(new_n13970_), .ZN(new_n14185_));
  NAND2_X1   g13183(.A1(new_n14180_), .A2(new_n14185_), .ZN(new_n14186_));
  AND2_X2    g13184(.A1(new_n13938_), .A2(new_n13940_), .Z(new_n14187_));
  NOR2_X1    g13185(.A1(new_n13938_), .A2(new_n13940_), .ZN(new_n14188_));
  INV_X1     g13186(.I(new_n14188_), .ZN(new_n14189_));
  OAI21_X1   g13187(.A1(new_n13716_), .A2(new_n14187_), .B(new_n14189_), .ZN(new_n14190_));
  NAND2_X1   g13188(.A1(new_n13721_), .A2(new_n13935_), .ZN(new_n14191_));
  NAND2_X1   g13189(.A1(new_n14191_), .A2(new_n13934_), .ZN(new_n14192_));
  INV_X1     g13190(.I(new_n14192_), .ZN(new_n14193_));
  NOR3_X1    g13191(.A1(new_n13981_), .A2(new_n13947_), .A3(new_n14193_), .ZN(new_n14194_));
  AOI21_X1   g13192(.A1(new_n13944_), .A2(new_n13982_), .B(new_n14192_), .ZN(new_n14195_));
  NOR3_X1    g13193(.A1(new_n14194_), .A2(new_n14195_), .A3(new_n14190_), .ZN(new_n14196_));
  INV_X1     g13194(.I(new_n14190_), .ZN(new_n14197_));
  NAND3_X1   g13195(.A1(new_n13944_), .A2(new_n13982_), .A3(new_n14192_), .ZN(new_n14198_));
  OAI21_X1   g13196(.A1(new_n13981_), .A2(new_n13947_), .B(new_n14193_), .ZN(new_n14199_));
  AOI21_X1   g13197(.A1(new_n14199_), .A2(new_n14198_), .B(new_n14197_), .ZN(new_n14200_));
  OAI21_X1   g13198(.A1(new_n14196_), .A2(new_n14200_), .B(new_n14186_), .ZN(new_n14201_));
  AOI21_X1   g13199(.A1(new_n14181_), .A2(new_n13970_), .B(new_n14184_), .ZN(new_n14202_));
  NOR3_X1    g13200(.A1(new_n14164_), .A2(new_n14179_), .A3(new_n13964_), .ZN(new_n14203_));
  NOR2_X1    g13201(.A1(new_n14203_), .A2(new_n14202_), .ZN(new_n14204_));
  NAND3_X1   g13202(.A1(new_n14199_), .A2(new_n14198_), .A3(new_n14197_), .ZN(new_n14205_));
  OAI21_X1   g13203(.A1(new_n14194_), .A2(new_n14195_), .B(new_n14190_), .ZN(new_n14206_));
  NAND3_X1   g13204(.A1(new_n14204_), .A2(new_n14206_), .A3(new_n14205_), .ZN(new_n14207_));
  NAND3_X1   g13205(.A1(new_n14207_), .A2(new_n14201_), .A3(new_n14163_), .ZN(new_n14208_));
  AOI21_X1   g13206(.A1(new_n13950_), .A2(new_n13972_), .B(new_n13987_), .ZN(new_n14209_));
  AOI21_X1   g13207(.A1(new_n14205_), .A2(new_n14206_), .B(new_n14204_), .ZN(new_n14210_));
  NOR3_X1    g13208(.A1(new_n14196_), .A2(new_n14200_), .A3(new_n14186_), .ZN(new_n14211_));
  OAI21_X1   g13209(.A1(new_n14210_), .A2(new_n14211_), .B(new_n14209_), .ZN(new_n14212_));
  NAND4_X1   g13210(.A1(new_n14158_), .A2(new_n14162_), .A3(new_n14212_), .A4(new_n14208_), .ZN(new_n14213_));
  NOR3_X1    g13211(.A1(new_n14159_), .A2(new_n14160_), .A3(new_n14161_), .ZN(new_n14214_));
  AOI21_X1   g13212(.A1(new_n14150_), .A2(new_n14156_), .B(new_n14157_), .ZN(new_n14215_));
  NOR3_X1    g13213(.A1(new_n14210_), .A2(new_n14211_), .A3(new_n14209_), .ZN(new_n14216_));
  AOI21_X1   g13214(.A1(new_n14207_), .A2(new_n14201_), .B(new_n14163_), .ZN(new_n14217_));
  OAI22_X1   g13215(.A1(new_n14214_), .A2(new_n14215_), .B1(new_n14217_), .B2(new_n14216_), .ZN(new_n14218_));
  NAND3_X1   g13216(.A1(new_n14218_), .A2(new_n14213_), .A3(new_n14112_), .ZN(new_n14219_));
  NOR3_X1    g13217(.A1(new_n13979_), .A2(new_n13988_), .A3(new_n13868_), .ZN(new_n14220_));
  AOI21_X1   g13218(.A1(new_n13931_), .A2(new_n13989_), .B(new_n14220_), .ZN(new_n14221_));
  NOR4_X1    g13219(.A1(new_n14214_), .A2(new_n14215_), .A3(new_n14217_), .A4(new_n14216_), .ZN(new_n14222_));
  AOI22_X1   g13220(.A1(new_n14162_), .A2(new_n14158_), .B1(new_n14212_), .B2(new_n14208_), .ZN(new_n14223_));
  OAI21_X1   g13221(.A1(new_n14222_), .A2(new_n14223_), .B(new_n14221_), .ZN(new_n14224_));
  NAND4_X1   g13222(.A1(new_n14105_), .A2(new_n14109_), .A3(new_n14224_), .A4(new_n14219_), .ZN(new_n14225_));
  AOI22_X1   g13223(.A1(new_n14109_), .A2(new_n14105_), .B1(new_n14224_), .B2(new_n14219_), .ZN(new_n14226_));
  OAI21_X1   g13224(.A1(new_n13999_), .A2(new_n14226_), .B(new_n14225_), .ZN(new_n14227_));
  OAI21_X1   g13225(.A1(new_n14221_), .A2(new_n14223_), .B(new_n14213_), .ZN(new_n14228_));
  NOR2_X1    g13226(.A1(new_n14210_), .A2(new_n14163_), .ZN(new_n14229_));
  OAI21_X1   g13227(.A1(new_n14197_), .A2(new_n14195_), .B(new_n14198_), .ZN(new_n14230_));
  NOR2_X1    g13228(.A1(new_n14164_), .A2(new_n13964_), .ZN(new_n14231_));
  AOI21_X1   g13229(.A1(new_n14231_), .A2(new_n14183_), .B(new_n14173_), .ZN(new_n14232_));
  NAND2_X1   g13230(.A1(new_n14230_), .A2(new_n14232_), .ZN(new_n14233_));
  INV_X1     g13231(.I(new_n14233_), .ZN(new_n14234_));
  NOR2_X1    g13232(.A1(new_n14230_), .A2(new_n14232_), .ZN(new_n14235_));
  NOR2_X1    g13233(.A1(new_n14234_), .A2(new_n14235_), .ZN(new_n14236_));
  OAI21_X1   g13234(.A1(new_n14211_), .A2(new_n14229_), .B(new_n14236_), .ZN(new_n14237_));
  NAND2_X1   g13235(.A1(new_n14201_), .A2(new_n14209_), .ZN(new_n14238_));
  INV_X1     g13236(.I(new_n14235_), .ZN(new_n14239_));
  NAND2_X1   g13237(.A1(new_n14239_), .A2(new_n14233_), .ZN(new_n14240_));
  NAND3_X1   g13238(.A1(new_n14240_), .A2(new_n14238_), .A3(new_n14207_), .ZN(new_n14241_));
  NOR2_X1    g13239(.A1(new_n14159_), .A2(new_n14157_), .ZN(new_n14242_));
  NAND2_X1   g13240(.A1(new_n14148_), .A2(new_n14138_), .ZN(new_n14243_));
  NAND2_X1   g13241(.A1(new_n14129_), .A2(new_n13893_), .ZN(new_n14244_));
  OAI21_X1   g13242(.A1(new_n14244_), .A2(new_n14126_), .B(new_n14130_), .ZN(new_n14245_));
  AOI21_X1   g13243(.A1(new_n14243_), .A2(new_n14147_), .B(new_n14245_), .ZN(new_n14246_));
  NOR2_X1    g13244(.A1(new_n14144_), .A2(new_n14146_), .ZN(new_n14247_));
  NOR2_X1    g13245(.A1(new_n14113_), .A2(new_n13892_), .ZN(new_n14248_));
  AOI21_X1   g13246(.A1(new_n14248_), .A2(new_n14131_), .B(new_n14122_), .ZN(new_n14249_));
  NOR3_X1    g13247(.A1(new_n14249_), .A2(new_n14247_), .A3(new_n14142_), .ZN(new_n14250_));
  NOR2_X1    g13248(.A1(new_n14250_), .A2(new_n14246_), .ZN(new_n14251_));
  OAI21_X1   g13249(.A1(new_n14242_), .A2(new_n14160_), .B(new_n14251_), .ZN(new_n14252_));
  NAND2_X1   g13250(.A1(new_n14150_), .A2(new_n14161_), .ZN(new_n14253_));
  OAI21_X1   g13251(.A1(new_n14142_), .A2(new_n14247_), .B(new_n14249_), .ZN(new_n14254_));
  NAND3_X1   g13252(.A1(new_n14243_), .A2(new_n14245_), .A3(new_n14147_), .ZN(new_n14255_));
  NAND2_X1   g13253(.A1(new_n14254_), .A2(new_n14255_), .ZN(new_n14256_));
  NAND3_X1   g13254(.A1(new_n14253_), .A2(new_n14256_), .A3(new_n14156_), .ZN(new_n14257_));
  NAND4_X1   g13255(.A1(new_n14237_), .A2(new_n14241_), .A3(new_n14257_), .A4(new_n14252_), .ZN(new_n14258_));
  AOI21_X1   g13256(.A1(new_n14207_), .A2(new_n14238_), .B(new_n14240_), .ZN(new_n14259_));
  NOR3_X1    g13257(.A1(new_n14236_), .A2(new_n14229_), .A3(new_n14211_), .ZN(new_n14260_));
  AOI21_X1   g13258(.A1(new_n14253_), .A2(new_n14156_), .B(new_n14256_), .ZN(new_n14261_));
  NOR3_X1    g13259(.A1(new_n14242_), .A2(new_n14251_), .A3(new_n14160_), .ZN(new_n14262_));
  OAI22_X1   g13260(.A1(new_n14259_), .A2(new_n14260_), .B1(new_n14261_), .B2(new_n14262_), .ZN(new_n14263_));
  NAND3_X1   g13261(.A1(new_n14228_), .A2(new_n14263_), .A3(new_n14258_), .ZN(new_n14264_));
  AOI21_X1   g13262(.A1(new_n14112_), .A2(new_n14218_), .B(new_n14222_), .ZN(new_n14265_));
  NAND2_X1   g13263(.A1(new_n14263_), .A2(new_n14258_), .ZN(new_n14266_));
  NAND2_X1   g13264(.A1(new_n14266_), .A2(new_n14265_), .ZN(new_n14267_));
  OAI21_X1   g13265(.A1(new_n14107_), .A2(new_n14108_), .B(new_n14098_), .ZN(new_n14268_));
  NOR2_X1    g13266(.A1(new_n14095_), .A2(new_n14046_), .ZN(new_n14269_));
  NAND2_X1   g13267(.A1(new_n14084_), .A2(new_n14077_), .ZN(new_n14270_));
  NAND2_X1   g13268(.A1(new_n14067_), .A2(new_n13331_), .ZN(new_n14271_));
  OAI21_X1   g13269(.A1(new_n14271_), .A2(new_n14063_), .B(new_n14068_), .ZN(new_n14272_));
  AOI21_X1   g13270(.A1(new_n14270_), .A2(new_n14083_), .B(new_n14272_), .ZN(new_n14273_));
  NOR2_X1    g13271(.A1(new_n14081_), .A2(new_n14076_), .ZN(new_n14274_));
  NOR2_X1    g13272(.A1(new_n14050_), .A2(new_n14047_), .ZN(new_n14275_));
  AOI21_X1   g13273(.A1(new_n14275_), .A2(new_n14069_), .B(new_n14059_), .ZN(new_n14276_));
  NOR3_X1    g13274(.A1(new_n14276_), .A2(new_n14274_), .A3(new_n14079_), .ZN(new_n14277_));
  NOR2_X1    g13275(.A1(new_n14277_), .A2(new_n14273_), .ZN(new_n14278_));
  OAI21_X1   g13276(.A1(new_n14269_), .A2(new_n14096_), .B(new_n14278_), .ZN(new_n14279_));
  NAND2_X1   g13277(.A1(new_n14086_), .A2(new_n14094_), .ZN(new_n14280_));
  OAI21_X1   g13278(.A1(new_n14079_), .A2(new_n14274_), .B(new_n14276_), .ZN(new_n14281_));
  NAND3_X1   g13279(.A1(new_n14270_), .A2(new_n14272_), .A3(new_n14083_), .ZN(new_n14282_));
  NAND2_X1   g13280(.A1(new_n14281_), .A2(new_n14282_), .ZN(new_n14283_));
  NAND3_X1   g13281(.A1(new_n14280_), .A2(new_n14283_), .A3(new_n14092_), .ZN(new_n14284_));
  NOR2_X1    g13282(.A1(new_n14042_), .A2(new_n14040_), .ZN(new_n14285_));
  OAI21_X1   g13283(.A1(new_n14025_), .A2(new_n14026_), .B(new_n14018_), .ZN(new_n14286_));
  NAND2_X1   g13284(.A1(new_n14286_), .A2(new_n14030_), .ZN(new_n14287_));
  AOI21_X1   g13285(.A1(new_n13437_), .A2(new_n13445_), .B(new_n13440_), .ZN(new_n14288_));
  AOI21_X1   g13286(.A1(new_n14288_), .A2(new_n14011_), .B(new_n14005_), .ZN(new_n14289_));
  XOR2_X1    g13287(.A1(new_n14287_), .A2(new_n14289_), .Z(new_n14290_));
  OAI21_X1   g13288(.A1(new_n14285_), .A2(new_n14043_), .B(new_n14290_), .ZN(new_n14291_));
  NAND2_X1   g13289(.A1(new_n14033_), .A2(new_n14044_), .ZN(new_n14292_));
  NAND2_X1   g13290(.A1(new_n14287_), .A2(new_n14289_), .ZN(new_n14293_));
  INV_X1     g13291(.I(new_n14289_), .ZN(new_n14294_));
  NAND3_X1   g13292(.A1(new_n14294_), .A2(new_n14030_), .A3(new_n14286_), .ZN(new_n14295_));
  NAND2_X1   g13293(.A1(new_n14295_), .A2(new_n14293_), .ZN(new_n14296_));
  NAND3_X1   g13294(.A1(new_n14292_), .A2(new_n14296_), .A3(new_n14039_), .ZN(new_n14297_));
  NAND4_X1   g13295(.A1(new_n14291_), .A2(new_n14297_), .A3(new_n14279_), .A4(new_n14284_), .ZN(new_n14298_));
  AOI21_X1   g13296(.A1(new_n14280_), .A2(new_n14092_), .B(new_n14283_), .ZN(new_n14299_));
  NOR3_X1    g13297(.A1(new_n14269_), .A2(new_n14278_), .A3(new_n14096_), .ZN(new_n14300_));
  AOI21_X1   g13298(.A1(new_n14292_), .A2(new_n14039_), .B(new_n14296_), .ZN(new_n14301_));
  NOR3_X1    g13299(.A1(new_n14285_), .A2(new_n14290_), .A3(new_n14043_), .ZN(new_n14302_));
  OAI22_X1   g13300(.A1(new_n14301_), .A2(new_n14302_), .B1(new_n14299_), .B2(new_n14300_), .ZN(new_n14303_));
  NAND3_X1   g13301(.A1(new_n14268_), .A2(new_n14298_), .A3(new_n14303_), .ZN(new_n14304_));
  AOI21_X1   g13302(.A1(new_n14103_), .A2(new_n14104_), .B(new_n14106_), .ZN(new_n14305_));
  NOR4_X1    g13303(.A1(new_n14301_), .A2(new_n14302_), .A3(new_n14299_), .A4(new_n14300_), .ZN(new_n14306_));
  AOI22_X1   g13304(.A1(new_n14291_), .A2(new_n14297_), .B1(new_n14279_), .B2(new_n14284_), .ZN(new_n14307_));
  OAI21_X1   g13305(.A1(new_n14306_), .A2(new_n14307_), .B(new_n14305_), .ZN(new_n14308_));
  NAND4_X1   g13306(.A1(new_n14267_), .A2(new_n14308_), .A3(new_n14264_), .A4(new_n14304_), .ZN(new_n14309_));
  NOR2_X1    g13307(.A1(new_n14266_), .A2(new_n14265_), .ZN(new_n14310_));
  AOI21_X1   g13308(.A1(new_n14258_), .A2(new_n14263_), .B(new_n14228_), .ZN(new_n14311_));
  NOR3_X1    g13309(.A1(new_n14305_), .A2(new_n14306_), .A3(new_n14307_), .ZN(new_n14312_));
  AOI21_X1   g13310(.A1(new_n14298_), .A2(new_n14303_), .B(new_n14268_), .ZN(new_n14313_));
  OAI22_X1   g13311(.A1(new_n14310_), .A2(new_n14311_), .B1(new_n14313_), .B2(new_n14312_), .ZN(new_n14314_));
  NAND3_X1   g13312(.A1(new_n14314_), .A2(new_n14309_), .A3(new_n14227_), .ZN(new_n14315_));
  INV_X1     g13313(.I(new_n13570_), .ZN(new_n14316_));
  INV_X1     g13314(.I(new_n13994_), .ZN(new_n14317_));
  AOI21_X1   g13315(.A1(new_n14317_), .A2(new_n13995_), .B(new_n13875_), .ZN(new_n14318_));
  NAND3_X1   g13316(.A1(new_n14317_), .A2(new_n13875_), .A3(new_n13995_), .ZN(new_n14319_));
  OAI21_X1   g13317(.A1(new_n14316_), .A2(new_n14318_), .B(new_n14319_), .ZN(new_n14320_));
  NOR3_X1    g13318(.A1(new_n14106_), .A2(new_n14107_), .A3(new_n14108_), .ZN(new_n14321_));
  AOI21_X1   g13319(.A1(new_n14103_), .A2(new_n14098_), .B(new_n14104_), .ZN(new_n14322_));
  NOR3_X1    g13320(.A1(new_n14222_), .A2(new_n14223_), .A3(new_n14221_), .ZN(new_n14323_));
  AOI21_X1   g13321(.A1(new_n14218_), .A2(new_n14213_), .B(new_n14112_), .ZN(new_n14324_));
  NOR4_X1    g13322(.A1(new_n14321_), .A2(new_n14322_), .A3(new_n14323_), .A4(new_n14324_), .ZN(new_n14325_));
  OAI22_X1   g13323(.A1(new_n14321_), .A2(new_n14322_), .B1(new_n14323_), .B2(new_n14324_), .ZN(new_n14326_));
  AOI21_X1   g13324(.A1(new_n14320_), .A2(new_n14326_), .B(new_n14325_), .ZN(new_n14327_));
  NOR4_X1    g13325(.A1(new_n14310_), .A2(new_n14313_), .A3(new_n14311_), .A4(new_n14312_), .ZN(new_n14328_));
  AOI22_X1   g13326(.A1(new_n14267_), .A2(new_n14264_), .B1(new_n14308_), .B2(new_n14304_), .ZN(new_n14329_));
  OAI21_X1   g13327(.A1(new_n14329_), .A2(new_n14328_), .B(new_n14327_), .ZN(new_n14330_));
  INV_X1     g13328(.I(\A[477] ), .ZN(new_n14331_));
  NOR2_X1    g13329(.A1(new_n14331_), .A2(\A[476] ), .ZN(new_n14332_));
  INV_X1     g13330(.I(\A[476] ), .ZN(new_n14333_));
  NOR2_X1    g13331(.A1(new_n14333_), .A2(\A[477] ), .ZN(new_n14334_));
  OAI21_X1   g13332(.A1(new_n14332_), .A2(new_n14334_), .B(\A[475] ), .ZN(new_n14335_));
  INV_X1     g13333(.I(\A[475] ), .ZN(new_n14336_));
  NAND2_X1   g13334(.A1(\A[476] ), .A2(\A[477] ), .ZN(new_n14337_));
  INV_X1     g13335(.I(new_n14337_), .ZN(new_n14338_));
  NOR2_X1    g13336(.A1(\A[476] ), .A2(\A[477] ), .ZN(new_n14339_));
  OAI21_X1   g13337(.A1(new_n14338_), .A2(new_n14339_), .B(new_n14336_), .ZN(new_n14340_));
  NAND2_X1   g13338(.A1(new_n14335_), .A2(new_n14340_), .ZN(new_n14341_));
  INV_X1     g13339(.I(\A[480] ), .ZN(new_n14342_));
  NOR2_X1    g13340(.A1(new_n14342_), .A2(\A[479] ), .ZN(new_n14343_));
  INV_X1     g13341(.I(\A[479] ), .ZN(new_n14344_));
  NOR2_X1    g13342(.A1(new_n14344_), .A2(\A[480] ), .ZN(new_n14345_));
  OAI21_X1   g13343(.A1(new_n14343_), .A2(new_n14345_), .B(\A[478] ), .ZN(new_n14346_));
  INV_X1     g13344(.I(\A[478] ), .ZN(new_n14347_));
  NAND2_X1   g13345(.A1(\A[479] ), .A2(\A[480] ), .ZN(new_n14348_));
  INV_X1     g13346(.I(new_n14348_), .ZN(new_n14349_));
  NOR2_X1    g13347(.A1(\A[479] ), .A2(\A[480] ), .ZN(new_n14350_));
  OAI21_X1   g13348(.A1(new_n14349_), .A2(new_n14350_), .B(new_n14347_), .ZN(new_n14351_));
  NAND2_X1   g13349(.A1(new_n14346_), .A2(new_n14351_), .ZN(new_n14352_));
  NOR2_X1    g13350(.A1(new_n14341_), .A2(new_n14352_), .ZN(new_n14353_));
  AOI21_X1   g13351(.A1(\A[479] ), .A2(\A[480] ), .B(\A[478] ), .ZN(new_n14354_));
  AOI21_X1   g13352(.A1(\A[476] ), .A2(\A[477] ), .B(\A[475] ), .ZN(new_n14355_));
  OAI22_X1   g13353(.A1(new_n14339_), .A2(new_n14355_), .B1(new_n14354_), .B2(new_n14350_), .ZN(new_n14356_));
  NOR4_X1    g13354(.A1(new_n14354_), .A2(new_n14355_), .A3(new_n14339_), .A4(new_n14350_), .ZN(new_n14357_));
  INV_X1     g13355(.I(new_n14357_), .ZN(new_n14358_));
  NAND2_X1   g13356(.A1(new_n14358_), .A2(new_n14356_), .ZN(new_n14359_));
  XOR2_X1    g13357(.A1(new_n14353_), .A2(new_n14359_), .Z(new_n14360_));
  INV_X1     g13358(.I(\A[483] ), .ZN(new_n14361_));
  NOR2_X1    g13359(.A1(new_n14361_), .A2(\A[482] ), .ZN(new_n14362_));
  INV_X1     g13360(.I(\A[482] ), .ZN(new_n14363_));
  NOR2_X1    g13361(.A1(new_n14363_), .A2(\A[483] ), .ZN(new_n14364_));
  OAI21_X1   g13362(.A1(new_n14362_), .A2(new_n14364_), .B(\A[481] ), .ZN(new_n14365_));
  INV_X1     g13363(.I(\A[481] ), .ZN(new_n14366_));
  NOR2_X1    g13364(.A1(\A[482] ), .A2(\A[483] ), .ZN(new_n14367_));
  NAND2_X1   g13365(.A1(\A[482] ), .A2(\A[483] ), .ZN(new_n14368_));
  INV_X1     g13366(.I(new_n14368_), .ZN(new_n14369_));
  OAI21_X1   g13367(.A1(new_n14369_), .A2(new_n14367_), .B(new_n14366_), .ZN(new_n14370_));
  NAND2_X1   g13368(.A1(new_n14365_), .A2(new_n14370_), .ZN(new_n14371_));
  INV_X1     g13369(.I(\A[486] ), .ZN(new_n14372_));
  NOR2_X1    g13370(.A1(new_n14372_), .A2(\A[485] ), .ZN(new_n14373_));
  INV_X1     g13371(.I(\A[485] ), .ZN(new_n14374_));
  NOR2_X1    g13372(.A1(new_n14374_), .A2(\A[486] ), .ZN(new_n14375_));
  OAI21_X1   g13373(.A1(new_n14373_), .A2(new_n14375_), .B(\A[484] ), .ZN(new_n14376_));
  INV_X1     g13374(.I(\A[484] ), .ZN(new_n14377_));
  NOR2_X1    g13375(.A1(\A[485] ), .A2(\A[486] ), .ZN(new_n14378_));
  NAND2_X1   g13376(.A1(\A[485] ), .A2(\A[486] ), .ZN(new_n14379_));
  INV_X1     g13377(.I(new_n14379_), .ZN(new_n14380_));
  OAI21_X1   g13378(.A1(new_n14380_), .A2(new_n14378_), .B(new_n14377_), .ZN(new_n14381_));
  NAND2_X1   g13379(.A1(new_n14376_), .A2(new_n14381_), .ZN(new_n14382_));
  NOR2_X1    g13380(.A1(new_n14371_), .A2(new_n14382_), .ZN(new_n14383_));
  AOI21_X1   g13381(.A1(new_n14377_), .A2(new_n14379_), .B(new_n14378_), .ZN(new_n14384_));
  AOI21_X1   g13382(.A1(\A[482] ), .A2(\A[483] ), .B(\A[481] ), .ZN(new_n14385_));
  NOR2_X1    g13383(.A1(new_n14385_), .A2(new_n14367_), .ZN(new_n14386_));
  XOR2_X1    g13384(.A1(new_n14384_), .A2(new_n14386_), .Z(new_n14387_));
  NOR2_X1    g13385(.A1(new_n14383_), .A2(new_n14387_), .ZN(new_n14388_));
  NAND2_X1   g13386(.A1(new_n14363_), .A2(\A[483] ), .ZN(new_n14389_));
  NAND2_X1   g13387(.A1(new_n14361_), .A2(\A[482] ), .ZN(new_n14390_));
  AOI21_X1   g13388(.A1(new_n14389_), .A2(new_n14390_), .B(new_n14366_), .ZN(new_n14391_));
  INV_X1     g13389(.I(new_n14367_), .ZN(new_n14392_));
  AOI21_X1   g13390(.A1(new_n14392_), .A2(new_n14368_), .B(\A[481] ), .ZN(new_n14393_));
  NOR2_X1    g13391(.A1(new_n14393_), .A2(new_n14391_), .ZN(new_n14394_));
  NAND2_X1   g13392(.A1(new_n14374_), .A2(\A[486] ), .ZN(new_n14395_));
  NAND2_X1   g13393(.A1(new_n14372_), .A2(\A[485] ), .ZN(new_n14396_));
  AOI21_X1   g13394(.A1(new_n14395_), .A2(new_n14396_), .B(new_n14377_), .ZN(new_n14397_));
  INV_X1     g13395(.I(new_n14378_), .ZN(new_n14398_));
  AOI21_X1   g13396(.A1(new_n14398_), .A2(new_n14379_), .B(\A[484] ), .ZN(new_n14399_));
  NOR2_X1    g13397(.A1(new_n14399_), .A2(new_n14397_), .ZN(new_n14400_));
  NAND2_X1   g13398(.A1(new_n14394_), .A2(new_n14400_), .ZN(new_n14401_));
  XNOR2_X1   g13399(.A1(new_n14384_), .A2(new_n14386_), .ZN(new_n14402_));
  NOR2_X1    g13400(.A1(new_n14401_), .A2(new_n14402_), .ZN(new_n14403_));
  OR2_X2     g13401(.A1(new_n14403_), .A2(new_n14388_), .Z(new_n14404_));
  NOR2_X1    g13402(.A1(new_n14394_), .A2(new_n14400_), .ZN(new_n14405_));
  NOR2_X1    g13403(.A1(new_n14405_), .A2(new_n14383_), .ZN(new_n14406_));
  NAND2_X1   g13404(.A1(new_n14333_), .A2(\A[477] ), .ZN(new_n14407_));
  NAND2_X1   g13405(.A1(new_n14331_), .A2(\A[476] ), .ZN(new_n14408_));
  AOI21_X1   g13406(.A1(new_n14407_), .A2(new_n14408_), .B(new_n14336_), .ZN(new_n14409_));
  INV_X1     g13407(.I(new_n14339_), .ZN(new_n14410_));
  AOI21_X1   g13408(.A1(new_n14410_), .A2(new_n14337_), .B(\A[475] ), .ZN(new_n14411_));
  NOR2_X1    g13409(.A1(new_n14411_), .A2(new_n14409_), .ZN(new_n14412_));
  NAND2_X1   g13410(.A1(new_n14344_), .A2(\A[480] ), .ZN(new_n14413_));
  NAND2_X1   g13411(.A1(new_n14342_), .A2(\A[479] ), .ZN(new_n14414_));
  AOI21_X1   g13412(.A1(new_n14413_), .A2(new_n14414_), .B(new_n14347_), .ZN(new_n14415_));
  INV_X1     g13413(.I(new_n14350_), .ZN(new_n14416_));
  AOI21_X1   g13414(.A1(new_n14416_), .A2(new_n14348_), .B(\A[478] ), .ZN(new_n14417_));
  NOR2_X1    g13415(.A1(new_n14417_), .A2(new_n14415_), .ZN(new_n14418_));
  NOR2_X1    g13416(.A1(new_n14412_), .A2(new_n14418_), .ZN(new_n14419_));
  NOR2_X1    g13417(.A1(new_n14419_), .A2(new_n14353_), .ZN(new_n14420_));
  NAND2_X1   g13418(.A1(new_n14420_), .A2(new_n14406_), .ZN(new_n14421_));
  AOI21_X1   g13419(.A1(new_n14404_), .A2(new_n14421_), .B(new_n14360_), .ZN(new_n14422_));
  NAND2_X1   g13420(.A1(new_n14412_), .A2(new_n14418_), .ZN(new_n14423_));
  NAND2_X1   g13421(.A1(new_n14341_), .A2(new_n14352_), .ZN(new_n14424_));
  NAND2_X1   g13422(.A1(new_n14423_), .A2(new_n14424_), .ZN(new_n14425_));
  NOR4_X1    g13423(.A1(new_n14425_), .A2(new_n14383_), .A3(new_n14402_), .A4(new_n14405_), .ZN(new_n14426_));
  INV_X1     g13424(.I(new_n14384_), .ZN(new_n14427_));
  INV_X1     g13425(.I(new_n14386_), .ZN(new_n14428_));
  NOR2_X1    g13426(.A1(new_n14427_), .A2(new_n14428_), .ZN(new_n14429_));
  INV_X1     g13427(.I(new_n14429_), .ZN(new_n14430_));
  NOR2_X1    g13428(.A1(new_n14384_), .A2(new_n14386_), .ZN(new_n14431_));
  AOI21_X1   g13429(.A1(new_n14401_), .A2(new_n14430_), .B(new_n14431_), .ZN(new_n14432_));
  INV_X1     g13430(.I(new_n14356_), .ZN(new_n14433_));
  AOI21_X1   g13431(.A1(new_n14423_), .A2(new_n14358_), .B(new_n14433_), .ZN(new_n14434_));
  NOR2_X1    g13432(.A1(new_n14432_), .A2(new_n14434_), .ZN(new_n14435_));
  INV_X1     g13433(.I(new_n14431_), .ZN(new_n14436_));
  OAI21_X1   g13434(.A1(new_n14383_), .A2(new_n14429_), .B(new_n14436_), .ZN(new_n14437_));
  OAI21_X1   g13435(.A1(new_n14353_), .A2(new_n14357_), .B(new_n14356_), .ZN(new_n14438_));
  NOR2_X1    g13436(.A1(new_n14437_), .A2(new_n14438_), .ZN(new_n14439_));
  NOR2_X1    g13437(.A1(new_n14435_), .A2(new_n14439_), .ZN(new_n14440_));
  OAI21_X1   g13438(.A1(new_n14422_), .A2(new_n14426_), .B(new_n14440_), .ZN(new_n14441_));
  XOR2_X1    g13439(.A1(new_n14423_), .A2(new_n14359_), .Z(new_n14442_));
  NAND2_X1   g13440(.A1(new_n14371_), .A2(new_n14382_), .ZN(new_n14443_));
  NAND2_X1   g13441(.A1(new_n14401_), .A2(new_n14443_), .ZN(new_n14444_));
  OAI22_X1   g13442(.A1(new_n14444_), .A2(new_n14425_), .B1(new_n14403_), .B2(new_n14388_), .ZN(new_n14445_));
  AOI21_X1   g13443(.A1(new_n14445_), .A2(new_n14442_), .B(new_n14426_), .ZN(new_n14446_));
  NAND2_X1   g13444(.A1(new_n14437_), .A2(new_n14438_), .ZN(new_n14447_));
  NAND2_X1   g13445(.A1(new_n14432_), .A2(new_n14434_), .ZN(new_n14448_));
  NAND2_X1   g13446(.A1(new_n14448_), .A2(new_n14447_), .ZN(new_n14449_));
  NAND2_X1   g13447(.A1(new_n14446_), .A2(new_n14449_), .ZN(new_n14450_));
  NAND2_X1   g13448(.A1(new_n14441_), .A2(new_n14450_), .ZN(new_n14451_));
  INV_X1     g13449(.I(\A[471] ), .ZN(new_n14452_));
  NOR2_X1    g13450(.A1(new_n14452_), .A2(\A[470] ), .ZN(new_n14453_));
  INV_X1     g13451(.I(\A[470] ), .ZN(new_n14454_));
  NOR2_X1    g13452(.A1(new_n14454_), .A2(\A[471] ), .ZN(new_n14455_));
  OAI21_X1   g13453(.A1(new_n14453_), .A2(new_n14455_), .B(\A[469] ), .ZN(new_n14456_));
  INV_X1     g13454(.I(\A[469] ), .ZN(new_n14457_));
  NOR2_X1    g13455(.A1(\A[470] ), .A2(\A[471] ), .ZN(new_n14458_));
  NAND2_X1   g13456(.A1(\A[470] ), .A2(\A[471] ), .ZN(new_n14459_));
  INV_X1     g13457(.I(new_n14459_), .ZN(new_n14460_));
  OAI21_X1   g13458(.A1(new_n14460_), .A2(new_n14458_), .B(new_n14457_), .ZN(new_n14461_));
  NAND2_X1   g13459(.A1(new_n14456_), .A2(new_n14461_), .ZN(new_n14462_));
  INV_X1     g13460(.I(\A[474] ), .ZN(new_n14463_));
  NOR2_X1    g13461(.A1(new_n14463_), .A2(\A[473] ), .ZN(new_n14464_));
  INV_X1     g13462(.I(\A[473] ), .ZN(new_n14465_));
  NOR2_X1    g13463(.A1(new_n14465_), .A2(\A[474] ), .ZN(new_n14466_));
  OAI21_X1   g13464(.A1(new_n14464_), .A2(new_n14466_), .B(\A[472] ), .ZN(new_n14467_));
  INV_X1     g13465(.I(\A[472] ), .ZN(new_n14468_));
  NOR2_X1    g13466(.A1(\A[473] ), .A2(\A[474] ), .ZN(new_n14469_));
  NAND2_X1   g13467(.A1(\A[473] ), .A2(\A[474] ), .ZN(new_n14470_));
  INV_X1     g13468(.I(new_n14470_), .ZN(new_n14471_));
  OAI21_X1   g13469(.A1(new_n14471_), .A2(new_n14469_), .B(new_n14468_), .ZN(new_n14472_));
  NAND2_X1   g13470(.A1(new_n14467_), .A2(new_n14472_), .ZN(new_n14473_));
  NOR2_X1    g13471(.A1(new_n14462_), .A2(new_n14473_), .ZN(new_n14474_));
  AOI21_X1   g13472(.A1(new_n14468_), .A2(new_n14470_), .B(new_n14469_), .ZN(new_n14475_));
  AOI21_X1   g13473(.A1(\A[470] ), .A2(\A[471] ), .B(\A[469] ), .ZN(new_n14476_));
  NOR2_X1    g13474(.A1(new_n14476_), .A2(new_n14458_), .ZN(new_n14477_));
  AND2_X2    g13475(.A1(new_n14475_), .A2(new_n14477_), .Z(new_n14478_));
  NOR2_X1    g13476(.A1(new_n14475_), .A2(new_n14477_), .ZN(new_n14479_));
  INV_X1     g13477(.I(new_n14479_), .ZN(new_n14480_));
  OAI21_X1   g13478(.A1(new_n14474_), .A2(new_n14478_), .B(new_n14480_), .ZN(new_n14481_));
  INV_X1     g13479(.I(\A[466] ), .ZN(new_n14482_));
  INV_X1     g13480(.I(\A[467] ), .ZN(new_n14483_));
  NAND2_X1   g13481(.A1(new_n14483_), .A2(\A[468] ), .ZN(new_n14484_));
  INV_X1     g13482(.I(\A[468] ), .ZN(new_n14485_));
  NAND2_X1   g13483(.A1(new_n14485_), .A2(\A[467] ), .ZN(new_n14486_));
  AOI21_X1   g13484(.A1(new_n14484_), .A2(new_n14486_), .B(new_n14482_), .ZN(new_n14487_));
  NAND2_X1   g13485(.A1(\A[467] ), .A2(\A[468] ), .ZN(new_n14488_));
  NOR2_X1    g13486(.A1(\A[467] ), .A2(\A[468] ), .ZN(new_n14489_));
  INV_X1     g13487(.I(new_n14489_), .ZN(new_n14490_));
  AOI21_X1   g13488(.A1(new_n14490_), .A2(new_n14488_), .B(\A[466] ), .ZN(new_n14491_));
  INV_X1     g13489(.I(\A[463] ), .ZN(new_n14492_));
  INV_X1     g13490(.I(\A[464] ), .ZN(new_n14493_));
  NAND2_X1   g13491(.A1(new_n14493_), .A2(\A[465] ), .ZN(new_n14494_));
  INV_X1     g13492(.I(\A[465] ), .ZN(new_n14495_));
  NAND2_X1   g13493(.A1(new_n14495_), .A2(\A[464] ), .ZN(new_n14496_));
  AOI21_X1   g13494(.A1(new_n14494_), .A2(new_n14496_), .B(new_n14492_), .ZN(new_n14497_));
  NAND2_X1   g13495(.A1(\A[464] ), .A2(\A[465] ), .ZN(new_n14498_));
  NOR2_X1    g13496(.A1(\A[464] ), .A2(\A[465] ), .ZN(new_n14499_));
  INV_X1     g13497(.I(new_n14499_), .ZN(new_n14500_));
  AOI21_X1   g13498(.A1(new_n14500_), .A2(new_n14498_), .B(\A[463] ), .ZN(new_n14501_));
  NOR4_X1    g13499(.A1(new_n14487_), .A2(new_n14491_), .A3(new_n14501_), .A4(new_n14497_), .ZN(new_n14502_));
  AOI21_X1   g13500(.A1(new_n14482_), .A2(new_n14488_), .B(new_n14489_), .ZN(new_n14503_));
  AOI21_X1   g13501(.A1(\A[464] ), .A2(\A[465] ), .B(\A[463] ), .ZN(new_n14504_));
  NOR2_X1    g13502(.A1(new_n14504_), .A2(new_n14499_), .ZN(new_n14505_));
  NOR2_X1    g13503(.A1(new_n14503_), .A2(new_n14505_), .ZN(new_n14506_));
  INV_X1     g13504(.I(new_n14506_), .ZN(new_n14507_));
  NAND2_X1   g13505(.A1(new_n14503_), .A2(new_n14505_), .ZN(new_n14508_));
  NAND2_X1   g13506(.A1(new_n14507_), .A2(new_n14508_), .ZN(new_n14509_));
  NOR2_X1    g13507(.A1(new_n14509_), .A2(new_n14502_), .ZN(new_n14510_));
  NOR2_X1    g13508(.A1(new_n14491_), .A2(new_n14487_), .ZN(new_n14511_));
  NOR2_X1    g13509(.A1(new_n14501_), .A2(new_n14497_), .ZN(new_n14512_));
  NAND2_X1   g13510(.A1(new_n14511_), .A2(new_n14512_), .ZN(new_n14513_));
  INV_X1     g13511(.I(new_n14508_), .ZN(new_n14514_));
  NOR2_X1    g13512(.A1(new_n14514_), .A2(new_n14506_), .ZN(new_n14515_));
  NOR2_X1    g13513(.A1(new_n14513_), .A2(new_n14515_), .ZN(new_n14516_));
  NOR2_X1    g13514(.A1(new_n14516_), .A2(new_n14510_), .ZN(new_n14517_));
  NAND2_X1   g13515(.A1(new_n14454_), .A2(\A[471] ), .ZN(new_n14518_));
  NAND2_X1   g13516(.A1(new_n14452_), .A2(\A[470] ), .ZN(new_n14519_));
  AOI21_X1   g13517(.A1(new_n14518_), .A2(new_n14519_), .B(new_n14457_), .ZN(new_n14520_));
  INV_X1     g13518(.I(new_n14458_), .ZN(new_n14521_));
  AOI21_X1   g13519(.A1(new_n14521_), .A2(new_n14459_), .B(\A[469] ), .ZN(new_n14522_));
  NOR2_X1    g13520(.A1(new_n14522_), .A2(new_n14520_), .ZN(new_n14523_));
  NAND2_X1   g13521(.A1(new_n14465_), .A2(\A[474] ), .ZN(new_n14524_));
  NAND2_X1   g13522(.A1(new_n14463_), .A2(\A[473] ), .ZN(new_n14525_));
  AOI21_X1   g13523(.A1(new_n14524_), .A2(new_n14525_), .B(new_n14468_), .ZN(new_n14526_));
  INV_X1     g13524(.I(new_n14469_), .ZN(new_n14527_));
  AOI21_X1   g13525(.A1(new_n14527_), .A2(new_n14470_), .B(\A[472] ), .ZN(new_n14528_));
  NOR2_X1    g13526(.A1(new_n14528_), .A2(new_n14526_), .ZN(new_n14529_));
  NAND2_X1   g13527(.A1(new_n14523_), .A2(new_n14529_), .ZN(new_n14530_));
  XOR2_X1    g13528(.A1(new_n14475_), .A2(new_n14477_), .Z(new_n14531_));
  XOR2_X1    g13529(.A1(new_n14530_), .A2(new_n14531_), .Z(new_n14532_));
  NOR2_X1    g13530(.A1(new_n14523_), .A2(new_n14529_), .ZN(new_n14533_));
  NOR2_X1    g13531(.A1(new_n14533_), .A2(new_n14474_), .ZN(new_n14534_));
  NOR2_X1    g13532(.A1(new_n14511_), .A2(new_n14512_), .ZN(new_n14535_));
  NOR2_X1    g13533(.A1(new_n14535_), .A2(new_n14502_), .ZN(new_n14536_));
  NAND2_X1   g13534(.A1(new_n14534_), .A2(new_n14536_), .ZN(new_n14537_));
  AOI21_X1   g13535(.A1(new_n14532_), .A2(new_n14537_), .B(new_n14517_), .ZN(new_n14538_));
  NAND2_X1   g13536(.A1(new_n14462_), .A2(new_n14473_), .ZN(new_n14539_));
  NAND4_X1   g13537(.A1(new_n14536_), .A2(new_n14530_), .A3(new_n14531_), .A4(new_n14539_), .ZN(new_n14540_));
  INV_X1     g13538(.I(new_n14540_), .ZN(new_n14541_));
  AOI21_X1   g13539(.A1(new_n14513_), .A2(new_n14508_), .B(new_n14506_), .ZN(new_n14542_));
  NOR3_X1    g13540(.A1(new_n14538_), .A2(new_n14541_), .A3(new_n14542_), .ZN(new_n14543_));
  NAND2_X1   g13541(.A1(new_n14513_), .A2(new_n14515_), .ZN(new_n14544_));
  NAND2_X1   g13542(.A1(new_n14509_), .A2(new_n14502_), .ZN(new_n14545_));
  NAND2_X1   g13543(.A1(new_n14544_), .A2(new_n14545_), .ZN(new_n14546_));
  NOR2_X1    g13544(.A1(new_n14474_), .A2(new_n14531_), .ZN(new_n14547_));
  XNOR2_X1   g13545(.A1(new_n14475_), .A2(new_n14477_), .ZN(new_n14548_));
  NOR2_X1    g13546(.A1(new_n14530_), .A2(new_n14548_), .ZN(new_n14549_));
  NOR2_X1    g13547(.A1(new_n14549_), .A2(new_n14547_), .ZN(new_n14550_));
  NAND2_X1   g13548(.A1(new_n14530_), .A2(new_n14539_), .ZN(new_n14551_));
  OAI22_X1   g13549(.A1(new_n14487_), .A2(new_n14491_), .B1(new_n14501_), .B2(new_n14497_), .ZN(new_n14552_));
  NAND2_X1   g13550(.A1(new_n14513_), .A2(new_n14552_), .ZN(new_n14553_));
  NOR2_X1    g13551(.A1(new_n14551_), .A2(new_n14553_), .ZN(new_n14554_));
  OAI21_X1   g13552(.A1(new_n14550_), .A2(new_n14554_), .B(new_n14546_), .ZN(new_n14555_));
  INV_X1     g13553(.I(new_n14542_), .ZN(new_n14556_));
  AOI21_X1   g13554(.A1(new_n14555_), .A2(new_n14540_), .B(new_n14556_), .ZN(new_n14557_));
  NOR3_X1    g13555(.A1(new_n14543_), .A2(new_n14557_), .A3(new_n14481_), .ZN(new_n14558_));
  INV_X1     g13556(.I(new_n14481_), .ZN(new_n14559_));
  NAND3_X1   g13557(.A1(new_n14555_), .A2(new_n14540_), .A3(new_n14556_), .ZN(new_n14560_));
  OAI21_X1   g13558(.A1(new_n14538_), .A2(new_n14541_), .B(new_n14542_), .ZN(new_n14561_));
  AOI21_X1   g13559(.A1(new_n14561_), .A2(new_n14560_), .B(new_n14559_), .ZN(new_n14562_));
  OAI21_X1   g13560(.A1(new_n14558_), .A2(new_n14562_), .B(new_n14451_), .ZN(new_n14563_));
  XOR2_X1    g13561(.A1(new_n14446_), .A2(new_n14449_), .Z(new_n14564_));
  NAND3_X1   g13562(.A1(new_n14561_), .A2(new_n14560_), .A3(new_n14559_), .ZN(new_n14565_));
  OAI21_X1   g13563(.A1(new_n14543_), .A2(new_n14557_), .B(new_n14481_), .ZN(new_n14566_));
  NAND3_X1   g13564(.A1(new_n14564_), .A2(new_n14566_), .A3(new_n14565_), .ZN(new_n14567_));
  NOR2_X1    g13565(.A1(new_n14555_), .A2(new_n14541_), .ZN(new_n14568_));
  OAI22_X1   g13566(.A1(new_n14551_), .A2(new_n14553_), .B1(new_n14549_), .B2(new_n14547_), .ZN(new_n14569_));
  AOI21_X1   g13567(.A1(new_n14569_), .A2(new_n14540_), .B(new_n14546_), .ZN(new_n14570_));
  NOR2_X1    g13568(.A1(new_n14551_), .A2(new_n14536_), .ZN(new_n14571_));
  NOR2_X1    g13569(.A1(new_n14534_), .A2(new_n14553_), .ZN(new_n14572_));
  NOR2_X1    g13570(.A1(new_n14420_), .A2(new_n14444_), .ZN(new_n14573_));
  NOR2_X1    g13571(.A1(new_n14406_), .A2(new_n14425_), .ZN(new_n14574_));
  OAI22_X1   g13572(.A1(new_n14573_), .A2(new_n14574_), .B1(new_n14571_), .B2(new_n14572_), .ZN(new_n14575_));
  OAI21_X1   g13573(.A1(new_n14568_), .A2(new_n14570_), .B(new_n14575_), .ZN(new_n14576_));
  INV_X1     g13574(.I(new_n14426_), .ZN(new_n14577_));
  NAND3_X1   g13575(.A1(new_n14577_), .A2(new_n14445_), .A3(new_n14360_), .ZN(new_n14578_));
  INV_X1     g13576(.I(new_n14445_), .ZN(new_n14579_));
  OAI21_X1   g13577(.A1(new_n14579_), .A2(new_n14426_), .B(new_n14442_), .ZN(new_n14580_));
  NAND2_X1   g13578(.A1(new_n14580_), .A2(new_n14578_), .ZN(new_n14581_));
  NOR3_X1    g13579(.A1(new_n14568_), .A2(new_n14575_), .A3(new_n14570_), .ZN(new_n14582_));
  OAI21_X1   g13580(.A1(new_n14581_), .A2(new_n14582_), .B(new_n14576_), .ZN(new_n14583_));
  NAND3_X1   g13581(.A1(new_n14567_), .A2(new_n14563_), .A3(new_n14583_), .ZN(new_n14584_));
  AOI21_X1   g13582(.A1(new_n14565_), .A2(new_n14566_), .B(new_n14564_), .ZN(new_n14585_));
  NOR3_X1    g13583(.A1(new_n14451_), .A2(new_n14558_), .A3(new_n14562_), .ZN(new_n14586_));
  NAND2_X1   g13584(.A1(new_n14538_), .A2(new_n14540_), .ZN(new_n14587_));
  INV_X1     g13585(.I(new_n14570_), .ZN(new_n14588_));
  NOR2_X1    g13586(.A1(new_n14571_), .A2(new_n14572_), .ZN(new_n14589_));
  NOR2_X1    g13587(.A1(new_n14573_), .A2(new_n14574_), .ZN(new_n14590_));
  NOR2_X1    g13588(.A1(new_n14590_), .A2(new_n14589_), .ZN(new_n14591_));
  AOI21_X1   g13589(.A1(new_n14588_), .A2(new_n14587_), .B(new_n14591_), .ZN(new_n14592_));
  INV_X1     g13590(.I(new_n14578_), .ZN(new_n14593_));
  AOI21_X1   g13591(.A1(new_n14577_), .A2(new_n14445_), .B(new_n14360_), .ZN(new_n14594_));
  NOR2_X1    g13592(.A1(new_n14593_), .A2(new_n14594_), .ZN(new_n14595_));
  NAND3_X1   g13593(.A1(new_n14588_), .A2(new_n14587_), .A3(new_n14591_), .ZN(new_n14596_));
  AOI21_X1   g13594(.A1(new_n14595_), .A2(new_n14596_), .B(new_n14592_), .ZN(new_n14597_));
  OAI21_X1   g13595(.A1(new_n14585_), .A2(new_n14586_), .B(new_n14597_), .ZN(new_n14598_));
  INV_X1     g13596(.I(\A[487] ), .ZN(new_n14599_));
  INV_X1     g13597(.I(\A[488] ), .ZN(new_n14600_));
  NAND2_X1   g13598(.A1(new_n14600_), .A2(\A[489] ), .ZN(new_n14601_));
  INV_X1     g13599(.I(\A[489] ), .ZN(new_n14602_));
  NAND2_X1   g13600(.A1(new_n14602_), .A2(\A[488] ), .ZN(new_n14603_));
  AOI21_X1   g13601(.A1(new_n14601_), .A2(new_n14603_), .B(new_n14599_), .ZN(new_n14604_));
  NAND2_X1   g13602(.A1(\A[488] ), .A2(\A[489] ), .ZN(new_n14605_));
  NOR2_X1    g13603(.A1(\A[488] ), .A2(\A[489] ), .ZN(new_n14606_));
  INV_X1     g13604(.I(new_n14606_), .ZN(new_n14607_));
  AOI21_X1   g13605(.A1(new_n14607_), .A2(new_n14605_), .B(\A[487] ), .ZN(new_n14608_));
  INV_X1     g13606(.I(\A[490] ), .ZN(new_n14609_));
  INV_X1     g13607(.I(\A[491] ), .ZN(new_n14610_));
  NAND2_X1   g13608(.A1(new_n14610_), .A2(\A[492] ), .ZN(new_n14611_));
  INV_X1     g13609(.I(\A[492] ), .ZN(new_n14612_));
  NAND2_X1   g13610(.A1(new_n14612_), .A2(\A[491] ), .ZN(new_n14613_));
  AOI21_X1   g13611(.A1(new_n14611_), .A2(new_n14613_), .B(new_n14609_), .ZN(new_n14614_));
  NAND2_X1   g13612(.A1(\A[491] ), .A2(\A[492] ), .ZN(new_n14615_));
  NOR2_X1    g13613(.A1(\A[491] ), .A2(\A[492] ), .ZN(new_n14616_));
  INV_X1     g13614(.I(new_n14616_), .ZN(new_n14617_));
  AOI21_X1   g13615(.A1(new_n14617_), .A2(new_n14615_), .B(\A[490] ), .ZN(new_n14618_));
  NOR4_X1    g13616(.A1(new_n14604_), .A2(new_n14608_), .A3(new_n14618_), .A4(new_n14614_), .ZN(new_n14619_));
  AOI21_X1   g13617(.A1(new_n14609_), .A2(new_n14615_), .B(new_n14616_), .ZN(new_n14620_));
  AOI21_X1   g13618(.A1(\A[488] ), .A2(\A[489] ), .B(\A[487] ), .ZN(new_n14621_));
  NOR2_X1    g13619(.A1(new_n14621_), .A2(new_n14606_), .ZN(new_n14622_));
  NOR2_X1    g13620(.A1(new_n14620_), .A2(new_n14622_), .ZN(new_n14623_));
  NAND2_X1   g13621(.A1(new_n14620_), .A2(new_n14622_), .ZN(new_n14624_));
  INV_X1     g13622(.I(new_n14624_), .ZN(new_n14625_));
  NOR2_X1    g13623(.A1(new_n14625_), .A2(new_n14623_), .ZN(new_n14626_));
  XNOR2_X1   g13624(.A1(new_n14626_), .A2(new_n14619_), .ZN(new_n14627_));
  INV_X1     g13625(.I(\A[495] ), .ZN(new_n14628_));
  NOR2_X1    g13626(.A1(new_n14628_), .A2(\A[494] ), .ZN(new_n14629_));
  INV_X1     g13627(.I(\A[494] ), .ZN(new_n14630_));
  NOR2_X1    g13628(.A1(new_n14630_), .A2(\A[495] ), .ZN(new_n14631_));
  OAI21_X1   g13629(.A1(new_n14629_), .A2(new_n14631_), .B(\A[493] ), .ZN(new_n14632_));
  INV_X1     g13630(.I(\A[493] ), .ZN(new_n14633_));
  NOR2_X1    g13631(.A1(\A[494] ), .A2(\A[495] ), .ZN(new_n14634_));
  NAND2_X1   g13632(.A1(\A[494] ), .A2(\A[495] ), .ZN(new_n14635_));
  INV_X1     g13633(.I(new_n14635_), .ZN(new_n14636_));
  OAI21_X1   g13634(.A1(new_n14636_), .A2(new_n14634_), .B(new_n14633_), .ZN(new_n14637_));
  NAND2_X1   g13635(.A1(new_n14632_), .A2(new_n14637_), .ZN(new_n14638_));
  INV_X1     g13636(.I(\A[498] ), .ZN(new_n14639_));
  NOR2_X1    g13637(.A1(new_n14639_), .A2(\A[497] ), .ZN(new_n14640_));
  INV_X1     g13638(.I(\A[497] ), .ZN(new_n14641_));
  NOR2_X1    g13639(.A1(new_n14641_), .A2(\A[498] ), .ZN(new_n14642_));
  OAI21_X1   g13640(.A1(new_n14640_), .A2(new_n14642_), .B(\A[496] ), .ZN(new_n14643_));
  INV_X1     g13641(.I(\A[496] ), .ZN(new_n14644_));
  NOR2_X1    g13642(.A1(\A[497] ), .A2(\A[498] ), .ZN(new_n14645_));
  NAND2_X1   g13643(.A1(\A[497] ), .A2(\A[498] ), .ZN(new_n14646_));
  INV_X1     g13644(.I(new_n14646_), .ZN(new_n14647_));
  OAI21_X1   g13645(.A1(new_n14647_), .A2(new_n14645_), .B(new_n14644_), .ZN(new_n14648_));
  NAND2_X1   g13646(.A1(new_n14643_), .A2(new_n14648_), .ZN(new_n14649_));
  NOR2_X1    g13647(.A1(new_n14638_), .A2(new_n14649_), .ZN(new_n14650_));
  AOI21_X1   g13648(.A1(new_n14644_), .A2(new_n14646_), .B(new_n14645_), .ZN(new_n14651_));
  AOI21_X1   g13649(.A1(new_n14633_), .A2(new_n14635_), .B(new_n14634_), .ZN(new_n14652_));
  XNOR2_X1   g13650(.A1(new_n14651_), .A2(new_n14652_), .ZN(new_n14653_));
  XOR2_X1    g13651(.A1(new_n14650_), .A2(new_n14653_), .Z(new_n14654_));
  NAND2_X1   g13652(.A1(new_n14630_), .A2(\A[495] ), .ZN(new_n14655_));
  NAND2_X1   g13653(.A1(new_n14628_), .A2(\A[494] ), .ZN(new_n14656_));
  AOI21_X1   g13654(.A1(new_n14655_), .A2(new_n14656_), .B(new_n14633_), .ZN(new_n14657_));
  INV_X1     g13655(.I(new_n14634_), .ZN(new_n14658_));
  AOI21_X1   g13656(.A1(new_n14658_), .A2(new_n14635_), .B(\A[493] ), .ZN(new_n14659_));
  NOR2_X1    g13657(.A1(new_n14659_), .A2(new_n14657_), .ZN(new_n14660_));
  NAND2_X1   g13658(.A1(new_n14641_), .A2(\A[498] ), .ZN(new_n14661_));
  NAND2_X1   g13659(.A1(new_n14639_), .A2(\A[497] ), .ZN(new_n14662_));
  AOI21_X1   g13660(.A1(new_n14661_), .A2(new_n14662_), .B(new_n14644_), .ZN(new_n14663_));
  INV_X1     g13661(.I(new_n14645_), .ZN(new_n14664_));
  AOI21_X1   g13662(.A1(new_n14664_), .A2(new_n14646_), .B(\A[496] ), .ZN(new_n14665_));
  NOR2_X1    g13663(.A1(new_n14665_), .A2(new_n14663_), .ZN(new_n14666_));
  NOR2_X1    g13664(.A1(new_n14660_), .A2(new_n14666_), .ZN(new_n14667_));
  NOR2_X1    g13665(.A1(new_n14667_), .A2(new_n14650_), .ZN(new_n14668_));
  OAI22_X1   g13666(.A1(new_n14604_), .A2(new_n14608_), .B1(new_n14618_), .B2(new_n14614_), .ZN(new_n14669_));
  INV_X1     g13667(.I(new_n14669_), .ZN(new_n14670_));
  NOR2_X1    g13668(.A1(new_n14670_), .A2(new_n14619_), .ZN(new_n14671_));
  NAND2_X1   g13669(.A1(new_n14671_), .A2(new_n14668_), .ZN(new_n14672_));
  AOI21_X1   g13670(.A1(new_n14654_), .A2(new_n14672_), .B(new_n14627_), .ZN(new_n14673_));
  NAND2_X1   g13671(.A1(new_n14660_), .A2(new_n14666_), .ZN(new_n14674_));
  XOR2_X1    g13672(.A1(new_n14674_), .A2(new_n14653_), .Z(new_n14675_));
  NAND2_X1   g13673(.A1(new_n14638_), .A2(new_n14649_), .ZN(new_n14676_));
  NAND2_X1   g13674(.A1(new_n14674_), .A2(new_n14676_), .ZN(new_n14677_));
  INV_X1     g13675(.I(new_n14619_), .ZN(new_n14678_));
  NAND2_X1   g13676(.A1(new_n14678_), .A2(new_n14669_), .ZN(new_n14679_));
  NOR2_X1    g13677(.A1(new_n14679_), .A2(new_n14677_), .ZN(new_n14680_));
  NAND2_X1   g13678(.A1(new_n14675_), .A2(new_n14680_), .ZN(new_n14681_));
  NAND2_X1   g13679(.A1(new_n14654_), .A2(new_n14672_), .ZN(new_n14682_));
  NAND2_X1   g13680(.A1(new_n14681_), .A2(new_n14682_), .ZN(new_n14683_));
  AOI22_X1   g13681(.A1(new_n14683_), .A2(new_n14627_), .B1(new_n14673_), .B2(new_n14681_), .ZN(new_n14684_));
  INV_X1     g13682(.I(\A[507] ), .ZN(new_n14685_));
  NOR2_X1    g13683(.A1(new_n14685_), .A2(\A[506] ), .ZN(new_n14686_));
  INV_X1     g13684(.I(\A[506] ), .ZN(new_n14687_));
  NOR2_X1    g13685(.A1(new_n14687_), .A2(\A[507] ), .ZN(new_n14688_));
  OAI21_X1   g13686(.A1(new_n14686_), .A2(new_n14688_), .B(\A[505] ), .ZN(new_n14689_));
  INV_X1     g13687(.I(\A[505] ), .ZN(new_n14690_));
  NOR2_X1    g13688(.A1(\A[506] ), .A2(\A[507] ), .ZN(new_n14691_));
  NAND2_X1   g13689(.A1(\A[506] ), .A2(\A[507] ), .ZN(new_n14692_));
  INV_X1     g13690(.I(new_n14692_), .ZN(new_n14693_));
  OAI21_X1   g13691(.A1(new_n14693_), .A2(new_n14691_), .B(new_n14690_), .ZN(new_n14694_));
  NAND2_X1   g13692(.A1(new_n14689_), .A2(new_n14694_), .ZN(new_n14695_));
  INV_X1     g13693(.I(\A[510] ), .ZN(new_n14696_));
  NOR2_X1    g13694(.A1(new_n14696_), .A2(\A[509] ), .ZN(new_n14697_));
  INV_X1     g13695(.I(\A[509] ), .ZN(new_n14698_));
  NOR2_X1    g13696(.A1(new_n14698_), .A2(\A[510] ), .ZN(new_n14699_));
  OAI21_X1   g13697(.A1(new_n14697_), .A2(new_n14699_), .B(\A[508] ), .ZN(new_n14700_));
  INV_X1     g13698(.I(\A[508] ), .ZN(new_n14701_));
  NOR2_X1    g13699(.A1(\A[509] ), .A2(\A[510] ), .ZN(new_n14702_));
  NAND2_X1   g13700(.A1(\A[509] ), .A2(\A[510] ), .ZN(new_n14703_));
  INV_X1     g13701(.I(new_n14703_), .ZN(new_n14704_));
  OAI21_X1   g13702(.A1(new_n14704_), .A2(new_n14702_), .B(new_n14701_), .ZN(new_n14705_));
  NAND2_X1   g13703(.A1(new_n14700_), .A2(new_n14705_), .ZN(new_n14706_));
  NOR2_X1    g13704(.A1(new_n14695_), .A2(new_n14706_), .ZN(new_n14707_));
  NAND2_X1   g13705(.A1(new_n14687_), .A2(\A[507] ), .ZN(new_n14708_));
  NAND2_X1   g13706(.A1(new_n14685_), .A2(\A[506] ), .ZN(new_n14709_));
  AOI21_X1   g13707(.A1(new_n14708_), .A2(new_n14709_), .B(new_n14690_), .ZN(new_n14710_));
  INV_X1     g13708(.I(new_n14691_), .ZN(new_n14711_));
  AOI21_X1   g13709(.A1(new_n14711_), .A2(new_n14692_), .B(\A[505] ), .ZN(new_n14712_));
  NOR2_X1    g13710(.A1(new_n14712_), .A2(new_n14710_), .ZN(new_n14713_));
  NAND2_X1   g13711(.A1(new_n14698_), .A2(\A[510] ), .ZN(new_n14714_));
  NAND2_X1   g13712(.A1(new_n14696_), .A2(\A[509] ), .ZN(new_n14715_));
  AOI21_X1   g13713(.A1(new_n14714_), .A2(new_n14715_), .B(new_n14701_), .ZN(new_n14716_));
  INV_X1     g13714(.I(new_n14702_), .ZN(new_n14717_));
  AOI21_X1   g13715(.A1(new_n14717_), .A2(new_n14703_), .B(\A[508] ), .ZN(new_n14718_));
  NOR2_X1    g13716(.A1(new_n14718_), .A2(new_n14716_), .ZN(new_n14719_));
  NOR2_X1    g13717(.A1(new_n14713_), .A2(new_n14719_), .ZN(new_n14720_));
  NOR2_X1    g13718(.A1(new_n14720_), .A2(new_n14707_), .ZN(new_n14721_));
  INV_X1     g13719(.I(\A[501] ), .ZN(new_n14722_));
  NOR2_X1    g13720(.A1(new_n14722_), .A2(\A[500] ), .ZN(new_n14723_));
  INV_X1     g13721(.I(\A[500] ), .ZN(new_n14724_));
  NOR2_X1    g13722(.A1(new_n14724_), .A2(\A[501] ), .ZN(new_n14725_));
  OAI21_X1   g13723(.A1(new_n14723_), .A2(new_n14725_), .B(\A[499] ), .ZN(new_n14726_));
  INV_X1     g13724(.I(\A[499] ), .ZN(new_n14727_));
  NAND2_X1   g13725(.A1(\A[500] ), .A2(\A[501] ), .ZN(new_n14728_));
  INV_X1     g13726(.I(new_n14728_), .ZN(new_n14729_));
  NOR2_X1    g13727(.A1(\A[500] ), .A2(\A[501] ), .ZN(new_n14730_));
  OAI21_X1   g13728(.A1(new_n14729_), .A2(new_n14730_), .B(new_n14727_), .ZN(new_n14731_));
  INV_X1     g13729(.I(\A[504] ), .ZN(new_n14732_));
  NOR2_X1    g13730(.A1(new_n14732_), .A2(\A[503] ), .ZN(new_n14733_));
  INV_X1     g13731(.I(\A[503] ), .ZN(new_n14734_));
  NOR2_X1    g13732(.A1(new_n14734_), .A2(\A[504] ), .ZN(new_n14735_));
  OAI21_X1   g13733(.A1(new_n14733_), .A2(new_n14735_), .B(\A[502] ), .ZN(new_n14736_));
  INV_X1     g13734(.I(\A[502] ), .ZN(new_n14737_));
  NAND2_X1   g13735(.A1(\A[503] ), .A2(\A[504] ), .ZN(new_n14738_));
  INV_X1     g13736(.I(new_n14738_), .ZN(new_n14739_));
  NOR2_X1    g13737(.A1(\A[503] ), .A2(\A[504] ), .ZN(new_n14740_));
  OAI21_X1   g13738(.A1(new_n14739_), .A2(new_n14740_), .B(new_n14737_), .ZN(new_n14741_));
  NAND4_X1   g13739(.A1(new_n14726_), .A2(new_n14731_), .A3(new_n14736_), .A4(new_n14741_), .ZN(new_n14742_));
  NAND2_X1   g13740(.A1(new_n14726_), .A2(new_n14731_), .ZN(new_n14743_));
  NAND2_X1   g13741(.A1(new_n14736_), .A2(new_n14741_), .ZN(new_n14744_));
  NAND2_X1   g13742(.A1(new_n14743_), .A2(new_n14744_), .ZN(new_n14745_));
  NAND2_X1   g13743(.A1(new_n14745_), .A2(new_n14742_), .ZN(new_n14746_));
  NAND2_X1   g13744(.A1(new_n14721_), .A2(new_n14746_), .ZN(new_n14747_));
  NAND2_X1   g13745(.A1(new_n14713_), .A2(new_n14719_), .ZN(new_n14748_));
  NAND2_X1   g13746(.A1(new_n14695_), .A2(new_n14706_), .ZN(new_n14749_));
  NAND2_X1   g13747(.A1(new_n14748_), .A2(new_n14749_), .ZN(new_n14750_));
  INV_X1     g13748(.I(new_n14746_), .ZN(new_n14751_));
  NAND2_X1   g13749(.A1(new_n14751_), .A2(new_n14750_), .ZN(new_n14752_));
  NAND2_X1   g13750(.A1(new_n14679_), .A2(new_n14668_), .ZN(new_n14753_));
  NAND2_X1   g13751(.A1(new_n14671_), .A2(new_n14677_), .ZN(new_n14754_));
  AOI22_X1   g13752(.A1(new_n14752_), .A2(new_n14747_), .B1(new_n14753_), .B2(new_n14754_), .ZN(new_n14755_));
  INV_X1     g13753(.I(new_n14755_), .ZN(new_n14756_));
  AOI21_X1   g13754(.A1(\A[503] ), .A2(\A[504] ), .B(\A[502] ), .ZN(new_n14757_));
  AOI21_X1   g13755(.A1(\A[500] ), .A2(\A[501] ), .B(\A[499] ), .ZN(new_n14758_));
  OAI22_X1   g13756(.A1(new_n14730_), .A2(new_n14758_), .B1(new_n14757_), .B2(new_n14740_), .ZN(new_n14759_));
  NOR4_X1    g13757(.A1(new_n14757_), .A2(new_n14758_), .A3(new_n14730_), .A4(new_n14740_), .ZN(new_n14760_));
  INV_X1     g13758(.I(new_n14760_), .ZN(new_n14761_));
  NAND2_X1   g13759(.A1(new_n14761_), .A2(new_n14759_), .ZN(new_n14762_));
  XNOR2_X1   g13760(.A1(new_n14742_), .A2(new_n14762_), .ZN(new_n14763_));
  AOI21_X1   g13761(.A1(new_n14701_), .A2(new_n14703_), .B(new_n14702_), .ZN(new_n14764_));
  AOI21_X1   g13762(.A1(new_n14690_), .A2(new_n14692_), .B(new_n14691_), .ZN(new_n14765_));
  XOR2_X1    g13763(.A1(new_n14764_), .A2(new_n14765_), .Z(new_n14766_));
  NOR2_X1    g13764(.A1(new_n14707_), .A2(new_n14766_), .ZN(new_n14767_));
  XNOR2_X1   g13765(.A1(new_n14764_), .A2(new_n14765_), .ZN(new_n14768_));
  NOR2_X1    g13766(.A1(new_n14748_), .A2(new_n14768_), .ZN(new_n14769_));
  OAI22_X1   g13767(.A1(new_n14750_), .A2(new_n14746_), .B1(new_n14769_), .B2(new_n14767_), .ZN(new_n14770_));
  NOR4_X1    g13768(.A1(new_n14746_), .A2(new_n14707_), .A3(new_n14720_), .A4(new_n14768_), .ZN(new_n14771_));
  INV_X1     g13769(.I(new_n14771_), .ZN(new_n14772_));
  NAND3_X1   g13770(.A1(new_n14772_), .A2(new_n14770_), .A3(new_n14763_), .ZN(new_n14773_));
  XOR2_X1    g13771(.A1(new_n14742_), .A2(new_n14762_), .Z(new_n14774_));
  INV_X1     g13772(.I(new_n14770_), .ZN(new_n14775_));
  OAI21_X1   g13773(.A1(new_n14775_), .A2(new_n14771_), .B(new_n14774_), .ZN(new_n14776_));
  AOI21_X1   g13774(.A1(new_n14776_), .A2(new_n14773_), .B(new_n14756_), .ZN(new_n14777_));
  NAND3_X1   g13775(.A1(new_n14756_), .A2(new_n14776_), .A3(new_n14773_), .ZN(new_n14778_));
  OAI21_X1   g13776(.A1(new_n14777_), .A2(new_n14684_), .B(new_n14778_), .ZN(new_n14779_));
  NOR2_X1    g13777(.A1(new_n14769_), .A2(new_n14767_), .ZN(new_n14780_));
  INV_X1     g13778(.I(new_n14780_), .ZN(new_n14781_));
  NAND2_X1   g13779(.A1(new_n14751_), .A2(new_n14721_), .ZN(new_n14782_));
  AOI21_X1   g13780(.A1(new_n14781_), .A2(new_n14782_), .B(new_n14763_), .ZN(new_n14783_));
  INV_X1     g13781(.I(new_n14764_), .ZN(new_n14784_));
  INV_X1     g13782(.I(new_n14765_), .ZN(new_n14785_));
  NOR2_X1    g13783(.A1(new_n14784_), .A2(new_n14785_), .ZN(new_n14786_));
  INV_X1     g13784(.I(new_n14786_), .ZN(new_n14787_));
  NOR2_X1    g13785(.A1(new_n14764_), .A2(new_n14765_), .ZN(new_n14788_));
  AOI21_X1   g13786(.A1(new_n14748_), .A2(new_n14787_), .B(new_n14788_), .ZN(new_n14789_));
  INV_X1     g13787(.I(new_n14759_), .ZN(new_n14790_));
  AOI21_X1   g13788(.A1(new_n14742_), .A2(new_n14761_), .B(new_n14790_), .ZN(new_n14791_));
  NOR2_X1    g13789(.A1(new_n14789_), .A2(new_n14791_), .ZN(new_n14792_));
  INV_X1     g13790(.I(new_n14788_), .ZN(new_n14793_));
  OAI21_X1   g13791(.A1(new_n14707_), .A2(new_n14786_), .B(new_n14793_), .ZN(new_n14794_));
  INV_X1     g13792(.I(new_n14791_), .ZN(new_n14795_));
  NOR2_X1    g13793(.A1(new_n14795_), .A2(new_n14794_), .ZN(new_n14796_));
  NOR2_X1    g13794(.A1(new_n14796_), .A2(new_n14792_), .ZN(new_n14797_));
  OAI21_X1   g13795(.A1(new_n14783_), .A2(new_n14771_), .B(new_n14797_), .ZN(new_n14798_));
  AOI21_X1   g13796(.A1(new_n14770_), .A2(new_n14774_), .B(new_n14771_), .ZN(new_n14799_));
  NAND2_X1   g13797(.A1(new_n14795_), .A2(new_n14794_), .ZN(new_n14800_));
  NAND2_X1   g13798(.A1(new_n14789_), .A2(new_n14791_), .ZN(new_n14801_));
  NAND2_X1   g13799(.A1(new_n14800_), .A2(new_n14801_), .ZN(new_n14802_));
  NAND2_X1   g13800(.A1(new_n14799_), .A2(new_n14802_), .ZN(new_n14803_));
  NAND2_X1   g13801(.A1(new_n14798_), .A2(new_n14803_), .ZN(new_n14804_));
  AND2_X2    g13802(.A1(new_n14651_), .A2(new_n14652_), .Z(new_n14805_));
  NOR2_X1    g13803(.A1(new_n14651_), .A2(new_n14652_), .ZN(new_n14806_));
  INV_X1     g13804(.I(new_n14806_), .ZN(new_n14807_));
  OAI21_X1   g13805(.A1(new_n14650_), .A2(new_n14805_), .B(new_n14807_), .ZN(new_n14808_));
  NOR2_X1    g13806(.A1(new_n14654_), .A2(new_n14672_), .ZN(new_n14809_));
  INV_X1     g13807(.I(new_n14623_), .ZN(new_n14810_));
  OAI21_X1   g13808(.A1(new_n14619_), .A2(new_n14625_), .B(new_n14810_), .ZN(new_n14811_));
  INV_X1     g13809(.I(new_n14811_), .ZN(new_n14812_));
  NOR3_X1    g13810(.A1(new_n14673_), .A2(new_n14809_), .A3(new_n14812_), .ZN(new_n14813_));
  XOR2_X1    g13811(.A1(new_n14626_), .A2(new_n14619_), .Z(new_n14814_));
  OAI21_X1   g13812(.A1(new_n14675_), .A2(new_n14680_), .B(new_n14814_), .ZN(new_n14815_));
  AOI21_X1   g13813(.A1(new_n14815_), .A2(new_n14681_), .B(new_n14811_), .ZN(new_n14816_));
  NOR3_X1    g13814(.A1(new_n14813_), .A2(new_n14816_), .A3(new_n14808_), .ZN(new_n14817_));
  INV_X1     g13815(.I(new_n14808_), .ZN(new_n14818_));
  NAND3_X1   g13816(.A1(new_n14815_), .A2(new_n14681_), .A3(new_n14811_), .ZN(new_n14819_));
  OAI21_X1   g13817(.A1(new_n14673_), .A2(new_n14809_), .B(new_n14812_), .ZN(new_n14820_));
  AOI21_X1   g13818(.A1(new_n14820_), .A2(new_n14819_), .B(new_n14818_), .ZN(new_n14821_));
  OAI21_X1   g13819(.A1(new_n14817_), .A2(new_n14821_), .B(new_n14804_), .ZN(new_n14822_));
  NOR2_X1    g13820(.A1(new_n14799_), .A2(new_n14802_), .ZN(new_n14823_));
  NOR3_X1    g13821(.A1(new_n14783_), .A2(new_n14771_), .A3(new_n14797_), .ZN(new_n14824_));
  NOR2_X1    g13822(.A1(new_n14824_), .A2(new_n14823_), .ZN(new_n14825_));
  NAND3_X1   g13823(.A1(new_n14820_), .A2(new_n14819_), .A3(new_n14818_), .ZN(new_n14826_));
  OAI21_X1   g13824(.A1(new_n14813_), .A2(new_n14816_), .B(new_n14808_), .ZN(new_n14827_));
  NAND3_X1   g13825(.A1(new_n14826_), .A2(new_n14827_), .A3(new_n14825_), .ZN(new_n14828_));
  NAND3_X1   g13826(.A1(new_n14828_), .A2(new_n14822_), .A3(new_n14779_), .ZN(new_n14829_));
  NOR2_X1    g13827(.A1(new_n14675_), .A2(new_n14680_), .ZN(new_n14830_));
  NOR2_X1    g13828(.A1(new_n14830_), .A2(new_n14809_), .ZN(new_n14831_));
  OAI22_X1   g13829(.A1(new_n14831_), .A2(new_n14814_), .B1(new_n14815_), .B2(new_n14809_), .ZN(new_n14832_));
  NOR3_X1    g13830(.A1(new_n14775_), .A2(new_n14774_), .A3(new_n14771_), .ZN(new_n14833_));
  AOI21_X1   g13831(.A1(new_n14772_), .A2(new_n14770_), .B(new_n14763_), .ZN(new_n14834_));
  OAI21_X1   g13832(.A1(new_n14833_), .A2(new_n14834_), .B(new_n14755_), .ZN(new_n14835_));
  NOR3_X1    g13833(.A1(new_n14833_), .A2(new_n14755_), .A3(new_n14834_), .ZN(new_n14836_));
  AOI21_X1   g13834(.A1(new_n14832_), .A2(new_n14835_), .B(new_n14836_), .ZN(new_n14837_));
  AOI21_X1   g13835(.A1(new_n14827_), .A2(new_n14826_), .B(new_n14825_), .ZN(new_n14838_));
  NOR3_X1    g13836(.A1(new_n14817_), .A2(new_n14821_), .A3(new_n14804_), .ZN(new_n14839_));
  OAI21_X1   g13837(.A1(new_n14838_), .A2(new_n14839_), .B(new_n14837_), .ZN(new_n14840_));
  NAND4_X1   g13838(.A1(new_n14598_), .A2(new_n14840_), .A3(new_n14829_), .A4(new_n14584_), .ZN(new_n14841_));
  NOR3_X1    g13839(.A1(new_n14585_), .A2(new_n14586_), .A3(new_n14597_), .ZN(new_n14842_));
  AOI21_X1   g13840(.A1(new_n14567_), .A2(new_n14563_), .B(new_n14583_), .ZN(new_n14843_));
  NOR3_X1    g13841(.A1(new_n14838_), .A2(new_n14839_), .A3(new_n14837_), .ZN(new_n14844_));
  AOI21_X1   g13842(.A1(new_n14828_), .A2(new_n14822_), .B(new_n14779_), .ZN(new_n14845_));
  OAI22_X1   g13843(.A1(new_n14844_), .A2(new_n14845_), .B1(new_n14842_), .B2(new_n14843_), .ZN(new_n14846_));
  NAND3_X1   g13844(.A1(new_n14596_), .A2(new_n14581_), .A3(new_n14576_), .ZN(new_n14847_));
  INV_X1     g13845(.I(new_n14847_), .ZN(new_n14848_));
  AOI21_X1   g13846(.A1(new_n14596_), .A2(new_n14576_), .B(new_n14581_), .ZN(new_n14849_));
  NAND2_X1   g13847(.A1(new_n14590_), .A2(new_n14589_), .ZN(new_n14850_));
  NAND2_X1   g13848(.A1(new_n14752_), .A2(new_n14747_), .ZN(new_n14851_));
  NAND2_X1   g13849(.A1(new_n14753_), .A2(new_n14754_), .ZN(new_n14852_));
  NOR2_X1    g13850(.A1(new_n14851_), .A2(new_n14852_), .ZN(new_n14853_));
  NOR2_X1    g13851(.A1(new_n14853_), .A2(new_n14755_), .ZN(new_n14854_));
  NAND3_X1   g13852(.A1(new_n14854_), .A2(new_n14575_), .A3(new_n14850_), .ZN(new_n14855_));
  OAI21_X1   g13853(.A1(new_n14848_), .A2(new_n14849_), .B(new_n14855_), .ZN(new_n14856_));
  NAND3_X1   g13854(.A1(new_n14832_), .A2(new_n14778_), .A3(new_n14835_), .ZN(new_n14857_));
  OAI21_X1   g13855(.A1(new_n14777_), .A2(new_n14836_), .B(new_n14684_), .ZN(new_n14858_));
  NAND2_X1   g13856(.A1(new_n14858_), .A2(new_n14857_), .ZN(new_n14859_));
  NOR3_X1    g13857(.A1(new_n14848_), .A2(new_n14849_), .A3(new_n14855_), .ZN(new_n14860_));
  OAI21_X1   g13858(.A1(new_n14859_), .A2(new_n14860_), .B(new_n14856_), .ZN(new_n14861_));
  NAND3_X1   g13859(.A1(new_n14846_), .A2(new_n14841_), .A3(new_n14861_), .ZN(new_n14862_));
  NOR4_X1    g13860(.A1(new_n14842_), .A2(new_n14845_), .A3(new_n14844_), .A4(new_n14843_), .ZN(new_n14863_));
  AOI22_X1   g13861(.A1(new_n14829_), .A2(new_n14840_), .B1(new_n14598_), .B2(new_n14584_), .ZN(new_n14864_));
  OAI21_X1   g13862(.A1(new_n14592_), .A2(new_n14582_), .B(new_n14595_), .ZN(new_n14865_));
  INV_X1     g13863(.I(new_n14855_), .ZN(new_n14866_));
  AOI21_X1   g13864(.A1(new_n14847_), .A2(new_n14865_), .B(new_n14866_), .ZN(new_n14867_));
  INV_X1     g13865(.I(new_n14859_), .ZN(new_n14868_));
  NAND3_X1   g13866(.A1(new_n14865_), .A2(new_n14866_), .A3(new_n14847_), .ZN(new_n14869_));
  AOI21_X1   g13867(.A1(new_n14868_), .A2(new_n14869_), .B(new_n14867_), .ZN(new_n14870_));
  OAI21_X1   g13868(.A1(new_n14864_), .A2(new_n14863_), .B(new_n14870_), .ZN(new_n14871_));
  INV_X1     g13869(.I(\A[525] ), .ZN(new_n14872_));
  NOR2_X1    g13870(.A1(new_n14872_), .A2(\A[524] ), .ZN(new_n14873_));
  INV_X1     g13871(.I(\A[524] ), .ZN(new_n14874_));
  NOR2_X1    g13872(.A1(new_n14874_), .A2(\A[525] ), .ZN(new_n14875_));
  OAI21_X1   g13873(.A1(new_n14873_), .A2(new_n14875_), .B(\A[523] ), .ZN(new_n14876_));
  INV_X1     g13874(.I(\A[523] ), .ZN(new_n14877_));
  NAND2_X1   g13875(.A1(\A[524] ), .A2(\A[525] ), .ZN(new_n14878_));
  INV_X1     g13876(.I(new_n14878_), .ZN(new_n14879_));
  NOR2_X1    g13877(.A1(\A[524] ), .A2(\A[525] ), .ZN(new_n14880_));
  OAI21_X1   g13878(.A1(new_n14879_), .A2(new_n14880_), .B(new_n14877_), .ZN(new_n14881_));
  INV_X1     g13879(.I(\A[528] ), .ZN(new_n14882_));
  NOR2_X1    g13880(.A1(new_n14882_), .A2(\A[527] ), .ZN(new_n14883_));
  INV_X1     g13881(.I(\A[527] ), .ZN(new_n14884_));
  NOR2_X1    g13882(.A1(new_n14884_), .A2(\A[528] ), .ZN(new_n14885_));
  OAI21_X1   g13883(.A1(new_n14883_), .A2(new_n14885_), .B(\A[526] ), .ZN(new_n14886_));
  INV_X1     g13884(.I(\A[526] ), .ZN(new_n14887_));
  NAND2_X1   g13885(.A1(\A[527] ), .A2(\A[528] ), .ZN(new_n14888_));
  INV_X1     g13886(.I(new_n14888_), .ZN(new_n14889_));
  NOR2_X1    g13887(.A1(\A[527] ), .A2(\A[528] ), .ZN(new_n14890_));
  OAI21_X1   g13888(.A1(new_n14889_), .A2(new_n14890_), .B(new_n14887_), .ZN(new_n14891_));
  NAND4_X1   g13889(.A1(new_n14876_), .A2(new_n14881_), .A3(new_n14886_), .A4(new_n14891_), .ZN(new_n14892_));
  AOI21_X1   g13890(.A1(\A[527] ), .A2(\A[528] ), .B(\A[526] ), .ZN(new_n14893_));
  NOR2_X1    g13891(.A1(new_n14893_), .A2(new_n14890_), .ZN(new_n14894_));
  AOI21_X1   g13892(.A1(\A[524] ), .A2(\A[525] ), .B(\A[523] ), .ZN(new_n14895_));
  NOR2_X1    g13893(.A1(new_n14895_), .A2(new_n14880_), .ZN(new_n14896_));
  NOR2_X1    g13894(.A1(new_n14894_), .A2(new_n14896_), .ZN(new_n14897_));
  NOR4_X1    g13895(.A1(new_n14893_), .A2(new_n14895_), .A3(new_n14880_), .A4(new_n14890_), .ZN(new_n14898_));
  NOR2_X1    g13896(.A1(new_n14897_), .A2(new_n14898_), .ZN(new_n14899_));
  XOR2_X1    g13897(.A1(new_n14892_), .A2(new_n14899_), .Z(new_n14900_));
  INV_X1     g13898(.I(\A[531] ), .ZN(new_n14901_));
  NOR2_X1    g13899(.A1(new_n14901_), .A2(\A[530] ), .ZN(new_n14902_));
  INV_X1     g13900(.I(\A[530] ), .ZN(new_n14903_));
  NOR2_X1    g13901(.A1(new_n14903_), .A2(\A[531] ), .ZN(new_n14904_));
  OAI21_X1   g13902(.A1(new_n14902_), .A2(new_n14904_), .B(\A[529] ), .ZN(new_n14905_));
  INV_X1     g13903(.I(\A[529] ), .ZN(new_n14906_));
  NOR2_X1    g13904(.A1(\A[530] ), .A2(\A[531] ), .ZN(new_n14907_));
  NAND2_X1   g13905(.A1(\A[530] ), .A2(\A[531] ), .ZN(new_n14908_));
  INV_X1     g13906(.I(new_n14908_), .ZN(new_n14909_));
  OAI21_X1   g13907(.A1(new_n14909_), .A2(new_n14907_), .B(new_n14906_), .ZN(new_n14910_));
  NAND2_X1   g13908(.A1(new_n14905_), .A2(new_n14910_), .ZN(new_n14911_));
  INV_X1     g13909(.I(\A[534] ), .ZN(new_n14912_));
  NOR2_X1    g13910(.A1(new_n14912_), .A2(\A[533] ), .ZN(new_n14913_));
  INV_X1     g13911(.I(\A[533] ), .ZN(new_n14914_));
  NOR2_X1    g13912(.A1(new_n14914_), .A2(\A[534] ), .ZN(new_n14915_));
  OAI21_X1   g13913(.A1(new_n14913_), .A2(new_n14915_), .B(\A[532] ), .ZN(new_n14916_));
  INV_X1     g13914(.I(\A[532] ), .ZN(new_n14917_));
  NOR2_X1    g13915(.A1(\A[533] ), .A2(\A[534] ), .ZN(new_n14918_));
  NAND2_X1   g13916(.A1(\A[533] ), .A2(\A[534] ), .ZN(new_n14919_));
  INV_X1     g13917(.I(new_n14919_), .ZN(new_n14920_));
  OAI21_X1   g13918(.A1(new_n14920_), .A2(new_n14918_), .B(new_n14917_), .ZN(new_n14921_));
  NAND2_X1   g13919(.A1(new_n14916_), .A2(new_n14921_), .ZN(new_n14922_));
  NOR2_X1    g13920(.A1(new_n14911_), .A2(new_n14922_), .ZN(new_n14923_));
  AOI21_X1   g13921(.A1(new_n14917_), .A2(new_n14919_), .B(new_n14918_), .ZN(new_n14924_));
  AOI21_X1   g13922(.A1(new_n14906_), .A2(new_n14908_), .B(new_n14907_), .ZN(new_n14925_));
  XOR2_X1    g13923(.A1(new_n14924_), .A2(new_n14925_), .Z(new_n14926_));
  NOR2_X1    g13924(.A1(new_n14923_), .A2(new_n14926_), .ZN(new_n14927_));
  NAND2_X1   g13925(.A1(new_n14903_), .A2(\A[531] ), .ZN(new_n14928_));
  NAND2_X1   g13926(.A1(new_n14901_), .A2(\A[530] ), .ZN(new_n14929_));
  AOI21_X1   g13927(.A1(new_n14928_), .A2(new_n14929_), .B(new_n14906_), .ZN(new_n14930_));
  INV_X1     g13928(.I(new_n14907_), .ZN(new_n14931_));
  AOI21_X1   g13929(.A1(new_n14931_), .A2(new_n14908_), .B(\A[529] ), .ZN(new_n14932_));
  NOR2_X1    g13930(.A1(new_n14932_), .A2(new_n14930_), .ZN(new_n14933_));
  NAND2_X1   g13931(.A1(new_n14914_), .A2(\A[534] ), .ZN(new_n14934_));
  NAND2_X1   g13932(.A1(new_n14912_), .A2(\A[533] ), .ZN(new_n14935_));
  AOI21_X1   g13933(.A1(new_n14934_), .A2(new_n14935_), .B(new_n14917_), .ZN(new_n14936_));
  INV_X1     g13934(.I(new_n14918_), .ZN(new_n14937_));
  AOI21_X1   g13935(.A1(new_n14937_), .A2(new_n14919_), .B(\A[532] ), .ZN(new_n14938_));
  NOR2_X1    g13936(.A1(new_n14938_), .A2(new_n14936_), .ZN(new_n14939_));
  NAND2_X1   g13937(.A1(new_n14933_), .A2(new_n14939_), .ZN(new_n14940_));
  XNOR2_X1   g13938(.A1(new_n14924_), .A2(new_n14925_), .ZN(new_n14941_));
  NOR2_X1    g13939(.A1(new_n14940_), .A2(new_n14941_), .ZN(new_n14942_));
  NAND2_X1   g13940(.A1(new_n14911_), .A2(new_n14922_), .ZN(new_n14943_));
  NAND2_X1   g13941(.A1(new_n14940_), .A2(new_n14943_), .ZN(new_n14944_));
  NAND2_X1   g13942(.A1(new_n14876_), .A2(new_n14881_), .ZN(new_n14945_));
  NAND2_X1   g13943(.A1(new_n14886_), .A2(new_n14891_), .ZN(new_n14946_));
  NAND2_X1   g13944(.A1(new_n14945_), .A2(new_n14946_), .ZN(new_n14947_));
  NAND2_X1   g13945(.A1(new_n14947_), .A2(new_n14892_), .ZN(new_n14948_));
  OAI22_X1   g13946(.A1(new_n14944_), .A2(new_n14948_), .B1(new_n14942_), .B2(new_n14927_), .ZN(new_n14949_));
  NOR2_X1    g13947(.A1(new_n14933_), .A2(new_n14939_), .ZN(new_n14950_));
  NOR4_X1    g13948(.A1(new_n14948_), .A2(new_n14923_), .A3(new_n14941_), .A4(new_n14950_), .ZN(new_n14951_));
  INV_X1     g13949(.I(new_n14951_), .ZN(new_n14952_));
  NAND3_X1   g13950(.A1(new_n14952_), .A2(new_n14949_), .A3(new_n14900_), .ZN(new_n14953_));
  INV_X1     g13951(.I(new_n14953_), .ZN(new_n14954_));
  AOI21_X1   g13952(.A1(new_n14952_), .A2(new_n14949_), .B(new_n14900_), .ZN(new_n14955_));
  NOR2_X1    g13953(.A1(new_n14954_), .A2(new_n14955_), .ZN(new_n14956_));
  INV_X1     g13954(.I(\A[511] ), .ZN(new_n14957_));
  INV_X1     g13955(.I(\A[512] ), .ZN(new_n14958_));
  NAND2_X1   g13956(.A1(new_n14958_), .A2(\A[513] ), .ZN(new_n14959_));
  INV_X1     g13957(.I(\A[513] ), .ZN(new_n14960_));
  NAND2_X1   g13958(.A1(new_n14960_), .A2(\A[512] ), .ZN(new_n14961_));
  AOI21_X1   g13959(.A1(new_n14959_), .A2(new_n14961_), .B(new_n14957_), .ZN(new_n14962_));
  NAND2_X1   g13960(.A1(\A[512] ), .A2(\A[513] ), .ZN(new_n14963_));
  NOR2_X1    g13961(.A1(\A[512] ), .A2(\A[513] ), .ZN(new_n14964_));
  INV_X1     g13962(.I(new_n14964_), .ZN(new_n14965_));
  AOI21_X1   g13963(.A1(new_n14965_), .A2(new_n14963_), .B(\A[511] ), .ZN(new_n14966_));
  INV_X1     g13964(.I(\A[514] ), .ZN(new_n14967_));
  INV_X1     g13965(.I(\A[515] ), .ZN(new_n14968_));
  NAND2_X1   g13966(.A1(new_n14968_), .A2(\A[516] ), .ZN(new_n14969_));
  INV_X1     g13967(.I(\A[516] ), .ZN(new_n14970_));
  NAND2_X1   g13968(.A1(new_n14970_), .A2(\A[515] ), .ZN(new_n14971_));
  AOI21_X1   g13969(.A1(new_n14969_), .A2(new_n14971_), .B(new_n14967_), .ZN(new_n14972_));
  NAND2_X1   g13970(.A1(\A[515] ), .A2(\A[516] ), .ZN(new_n14973_));
  NOR2_X1    g13971(.A1(\A[515] ), .A2(\A[516] ), .ZN(new_n14974_));
  INV_X1     g13972(.I(new_n14974_), .ZN(new_n14975_));
  AOI21_X1   g13973(.A1(new_n14975_), .A2(new_n14973_), .B(\A[514] ), .ZN(new_n14976_));
  NOR4_X1    g13974(.A1(new_n14962_), .A2(new_n14966_), .A3(new_n14976_), .A4(new_n14972_), .ZN(new_n14977_));
  AOI21_X1   g13975(.A1(new_n14967_), .A2(new_n14973_), .B(new_n14974_), .ZN(new_n14978_));
  AOI21_X1   g13976(.A1(new_n14957_), .A2(new_n14963_), .B(new_n14964_), .ZN(new_n14979_));
  XOR2_X1    g13977(.A1(new_n14978_), .A2(new_n14979_), .Z(new_n14980_));
  XNOR2_X1   g13978(.A1(new_n14980_), .A2(new_n14977_), .ZN(new_n14981_));
  INV_X1     g13979(.I(\A[519] ), .ZN(new_n14982_));
  NOR2_X1    g13980(.A1(new_n14982_), .A2(\A[518] ), .ZN(new_n14983_));
  INV_X1     g13981(.I(\A[518] ), .ZN(new_n14984_));
  NOR2_X1    g13982(.A1(new_n14984_), .A2(\A[519] ), .ZN(new_n14985_));
  OAI21_X1   g13983(.A1(new_n14983_), .A2(new_n14985_), .B(\A[517] ), .ZN(new_n14986_));
  INV_X1     g13984(.I(\A[517] ), .ZN(new_n14987_));
  NOR2_X1    g13985(.A1(\A[518] ), .A2(\A[519] ), .ZN(new_n14988_));
  NAND2_X1   g13986(.A1(\A[518] ), .A2(\A[519] ), .ZN(new_n14989_));
  INV_X1     g13987(.I(new_n14989_), .ZN(new_n14990_));
  OAI21_X1   g13988(.A1(new_n14990_), .A2(new_n14988_), .B(new_n14987_), .ZN(new_n14991_));
  NAND2_X1   g13989(.A1(new_n14986_), .A2(new_n14991_), .ZN(new_n14992_));
  INV_X1     g13990(.I(\A[522] ), .ZN(new_n14993_));
  NOR2_X1    g13991(.A1(new_n14993_), .A2(\A[521] ), .ZN(new_n14994_));
  INV_X1     g13992(.I(\A[521] ), .ZN(new_n14995_));
  NOR2_X1    g13993(.A1(new_n14995_), .A2(\A[522] ), .ZN(new_n14996_));
  OAI21_X1   g13994(.A1(new_n14994_), .A2(new_n14996_), .B(\A[520] ), .ZN(new_n14997_));
  INV_X1     g13995(.I(\A[520] ), .ZN(new_n14998_));
  NOR2_X1    g13996(.A1(\A[521] ), .A2(\A[522] ), .ZN(new_n14999_));
  NAND2_X1   g13997(.A1(\A[521] ), .A2(\A[522] ), .ZN(new_n15000_));
  INV_X1     g13998(.I(new_n15000_), .ZN(new_n15001_));
  OAI21_X1   g13999(.A1(new_n15001_), .A2(new_n14999_), .B(new_n14998_), .ZN(new_n15002_));
  NAND2_X1   g14000(.A1(new_n14997_), .A2(new_n15002_), .ZN(new_n15003_));
  NOR2_X1    g14001(.A1(new_n14992_), .A2(new_n15003_), .ZN(new_n15004_));
  AOI21_X1   g14002(.A1(new_n14998_), .A2(new_n15000_), .B(new_n14999_), .ZN(new_n15005_));
  AOI21_X1   g14003(.A1(new_n14987_), .A2(new_n14989_), .B(new_n14988_), .ZN(new_n15006_));
  XOR2_X1    g14004(.A1(new_n15005_), .A2(new_n15006_), .Z(new_n15007_));
  NOR2_X1    g14005(.A1(new_n15004_), .A2(new_n15007_), .ZN(new_n15008_));
  NAND2_X1   g14006(.A1(new_n14984_), .A2(\A[519] ), .ZN(new_n15009_));
  NAND2_X1   g14007(.A1(new_n14982_), .A2(\A[518] ), .ZN(new_n15010_));
  AOI21_X1   g14008(.A1(new_n15009_), .A2(new_n15010_), .B(new_n14987_), .ZN(new_n15011_));
  INV_X1     g14009(.I(new_n14988_), .ZN(new_n15012_));
  AOI21_X1   g14010(.A1(new_n15012_), .A2(new_n14989_), .B(\A[517] ), .ZN(new_n15013_));
  NOR2_X1    g14011(.A1(new_n15013_), .A2(new_n15011_), .ZN(new_n15014_));
  NAND2_X1   g14012(.A1(new_n14995_), .A2(\A[522] ), .ZN(new_n15015_));
  NAND2_X1   g14013(.A1(new_n14993_), .A2(\A[521] ), .ZN(new_n15016_));
  AOI21_X1   g14014(.A1(new_n15015_), .A2(new_n15016_), .B(new_n14998_), .ZN(new_n15017_));
  INV_X1     g14015(.I(new_n14999_), .ZN(new_n15018_));
  AOI21_X1   g14016(.A1(new_n15018_), .A2(new_n15000_), .B(\A[520] ), .ZN(new_n15019_));
  NOR2_X1    g14017(.A1(new_n15019_), .A2(new_n15017_), .ZN(new_n15020_));
  NAND2_X1   g14018(.A1(new_n15014_), .A2(new_n15020_), .ZN(new_n15021_));
  XNOR2_X1   g14019(.A1(new_n15005_), .A2(new_n15006_), .ZN(new_n15022_));
  NOR2_X1    g14020(.A1(new_n15021_), .A2(new_n15022_), .ZN(new_n15023_));
  NAND2_X1   g14021(.A1(new_n14992_), .A2(new_n15003_), .ZN(new_n15024_));
  NAND2_X1   g14022(.A1(new_n15021_), .A2(new_n15024_), .ZN(new_n15025_));
  OR4_X2     g14023(.A1(new_n14962_), .A2(new_n14966_), .A3(new_n14976_), .A4(new_n14972_), .Z(new_n15026_));
  OAI22_X1   g14024(.A1(new_n14962_), .A2(new_n14966_), .B1(new_n14976_), .B2(new_n14972_), .ZN(new_n15027_));
  NAND2_X1   g14025(.A1(new_n15026_), .A2(new_n15027_), .ZN(new_n15028_));
  OAI22_X1   g14026(.A1(new_n15025_), .A2(new_n15028_), .B1(new_n15023_), .B2(new_n15008_), .ZN(new_n15029_));
  INV_X1     g14027(.I(new_n15029_), .ZN(new_n15030_));
  NOR2_X1    g14028(.A1(new_n15014_), .A2(new_n15020_), .ZN(new_n15031_));
  NOR4_X1    g14029(.A1(new_n15028_), .A2(new_n15004_), .A3(new_n15022_), .A4(new_n15031_), .ZN(new_n15032_));
  NOR3_X1    g14030(.A1(new_n15030_), .A2(new_n14981_), .A3(new_n15032_), .ZN(new_n15033_));
  XOR2_X1    g14031(.A1(new_n14980_), .A2(new_n14977_), .Z(new_n15034_));
  INV_X1     g14032(.I(new_n15032_), .ZN(new_n15035_));
  AOI21_X1   g14033(.A1(new_n15035_), .A2(new_n15029_), .B(new_n15034_), .ZN(new_n15036_));
  NOR2_X1    g14034(.A1(new_n14950_), .A2(new_n14923_), .ZN(new_n15037_));
  NAND2_X1   g14035(.A1(new_n15037_), .A2(new_n14948_), .ZN(new_n15038_));
  INV_X1     g14036(.I(new_n15038_), .ZN(new_n15039_));
  NOR2_X1    g14037(.A1(new_n15037_), .A2(new_n14948_), .ZN(new_n15040_));
  NOR2_X1    g14038(.A1(new_n15031_), .A2(new_n15004_), .ZN(new_n15041_));
  NAND2_X1   g14039(.A1(new_n15041_), .A2(new_n15028_), .ZN(new_n15042_));
  INV_X1     g14040(.I(new_n15042_), .ZN(new_n15043_));
  NOR2_X1    g14041(.A1(new_n15041_), .A2(new_n15028_), .ZN(new_n15044_));
  OAI22_X1   g14042(.A1(new_n15039_), .A2(new_n15040_), .B1(new_n15043_), .B2(new_n15044_), .ZN(new_n15045_));
  NOR3_X1    g14043(.A1(new_n15033_), .A2(new_n15045_), .A3(new_n15036_), .ZN(new_n15046_));
  NAND3_X1   g14044(.A1(new_n15035_), .A2(new_n15029_), .A3(new_n15034_), .ZN(new_n15047_));
  OAI21_X1   g14045(.A1(new_n15030_), .A2(new_n15032_), .B(new_n14981_), .ZN(new_n15048_));
  INV_X1     g14046(.I(new_n15040_), .ZN(new_n15049_));
  INV_X1     g14047(.I(new_n15044_), .ZN(new_n15050_));
  AOI22_X1   g14048(.A1(new_n15038_), .A2(new_n15049_), .B1(new_n15050_), .B2(new_n15042_), .ZN(new_n15051_));
  AOI21_X1   g14049(.A1(new_n15048_), .A2(new_n15047_), .B(new_n15051_), .ZN(new_n15052_));
  NOR3_X1    g14050(.A1(new_n14956_), .A2(new_n15052_), .A3(new_n15046_), .ZN(new_n15053_));
  INV_X1     g14051(.I(new_n14955_), .ZN(new_n15054_));
  NAND2_X1   g14052(.A1(new_n15054_), .A2(new_n14953_), .ZN(new_n15055_));
  NAND3_X1   g14053(.A1(new_n15048_), .A2(new_n15051_), .A3(new_n15047_), .ZN(new_n15056_));
  OAI21_X1   g14054(.A1(new_n15033_), .A2(new_n15036_), .B(new_n15045_), .ZN(new_n15057_));
  AOI21_X1   g14055(.A1(new_n15057_), .A2(new_n15056_), .B(new_n15055_), .ZN(new_n15058_));
  NOR2_X1    g14056(.A1(new_n15058_), .A2(new_n15053_), .ZN(new_n15059_));
  INV_X1     g14057(.I(\A[555] ), .ZN(new_n15060_));
  NOR2_X1    g14058(.A1(new_n15060_), .A2(\A[554] ), .ZN(new_n15061_));
  INV_X1     g14059(.I(\A[554] ), .ZN(new_n15062_));
  NOR2_X1    g14060(.A1(new_n15062_), .A2(\A[555] ), .ZN(new_n15063_));
  OAI21_X1   g14061(.A1(new_n15061_), .A2(new_n15063_), .B(\A[553] ), .ZN(new_n15064_));
  INV_X1     g14062(.I(\A[553] ), .ZN(new_n15065_));
  NOR2_X1    g14063(.A1(\A[554] ), .A2(\A[555] ), .ZN(new_n15066_));
  NAND2_X1   g14064(.A1(\A[554] ), .A2(\A[555] ), .ZN(new_n15067_));
  INV_X1     g14065(.I(new_n15067_), .ZN(new_n15068_));
  OAI21_X1   g14066(.A1(new_n15068_), .A2(new_n15066_), .B(new_n15065_), .ZN(new_n15069_));
  NAND2_X1   g14067(.A1(new_n15064_), .A2(new_n15069_), .ZN(new_n15070_));
  INV_X1     g14068(.I(\A[558] ), .ZN(new_n15071_));
  NOR2_X1    g14069(.A1(new_n15071_), .A2(\A[557] ), .ZN(new_n15072_));
  INV_X1     g14070(.I(\A[557] ), .ZN(new_n15073_));
  NOR2_X1    g14071(.A1(new_n15073_), .A2(\A[558] ), .ZN(new_n15074_));
  OAI21_X1   g14072(.A1(new_n15072_), .A2(new_n15074_), .B(\A[556] ), .ZN(new_n15075_));
  INV_X1     g14073(.I(\A[556] ), .ZN(new_n15076_));
  NOR2_X1    g14074(.A1(\A[557] ), .A2(\A[558] ), .ZN(new_n15077_));
  NAND2_X1   g14075(.A1(\A[557] ), .A2(\A[558] ), .ZN(new_n15078_));
  INV_X1     g14076(.I(new_n15078_), .ZN(new_n15079_));
  OAI21_X1   g14077(.A1(new_n15079_), .A2(new_n15077_), .B(new_n15076_), .ZN(new_n15080_));
  NAND2_X1   g14078(.A1(new_n15075_), .A2(new_n15080_), .ZN(new_n15081_));
  NOR2_X1    g14079(.A1(new_n15070_), .A2(new_n15081_), .ZN(new_n15082_));
  NAND2_X1   g14080(.A1(new_n15062_), .A2(\A[555] ), .ZN(new_n15083_));
  NAND2_X1   g14081(.A1(new_n15060_), .A2(\A[554] ), .ZN(new_n15084_));
  AOI21_X1   g14082(.A1(new_n15083_), .A2(new_n15084_), .B(new_n15065_), .ZN(new_n15085_));
  INV_X1     g14083(.I(new_n15066_), .ZN(new_n15086_));
  AOI21_X1   g14084(.A1(new_n15086_), .A2(new_n15067_), .B(\A[553] ), .ZN(new_n15087_));
  NOR2_X1    g14085(.A1(new_n15087_), .A2(new_n15085_), .ZN(new_n15088_));
  NAND2_X1   g14086(.A1(new_n15073_), .A2(\A[558] ), .ZN(new_n15089_));
  NAND2_X1   g14087(.A1(new_n15071_), .A2(\A[557] ), .ZN(new_n15090_));
  AOI21_X1   g14088(.A1(new_n15089_), .A2(new_n15090_), .B(new_n15076_), .ZN(new_n15091_));
  INV_X1     g14089(.I(new_n15077_), .ZN(new_n15092_));
  AOI21_X1   g14090(.A1(new_n15092_), .A2(new_n15078_), .B(\A[556] ), .ZN(new_n15093_));
  NOR2_X1    g14091(.A1(new_n15093_), .A2(new_n15091_), .ZN(new_n15094_));
  NOR2_X1    g14092(.A1(new_n15088_), .A2(new_n15094_), .ZN(new_n15095_));
  NOR2_X1    g14093(.A1(new_n15095_), .A2(new_n15082_), .ZN(new_n15096_));
  INV_X1     g14094(.I(\A[547] ), .ZN(new_n15097_));
  INV_X1     g14095(.I(\A[548] ), .ZN(new_n15098_));
  NAND2_X1   g14096(.A1(new_n15098_), .A2(\A[549] ), .ZN(new_n15099_));
  INV_X1     g14097(.I(\A[549] ), .ZN(new_n15100_));
  NAND2_X1   g14098(.A1(new_n15100_), .A2(\A[548] ), .ZN(new_n15101_));
  AOI21_X1   g14099(.A1(new_n15099_), .A2(new_n15101_), .B(new_n15097_), .ZN(new_n15102_));
  NAND2_X1   g14100(.A1(\A[548] ), .A2(\A[549] ), .ZN(new_n15103_));
  NOR2_X1    g14101(.A1(\A[548] ), .A2(\A[549] ), .ZN(new_n15104_));
  INV_X1     g14102(.I(new_n15104_), .ZN(new_n15105_));
  AOI21_X1   g14103(.A1(new_n15105_), .A2(new_n15103_), .B(\A[547] ), .ZN(new_n15106_));
  NOR2_X1    g14104(.A1(new_n15106_), .A2(new_n15102_), .ZN(new_n15107_));
  INV_X1     g14105(.I(\A[550] ), .ZN(new_n15108_));
  INV_X1     g14106(.I(\A[551] ), .ZN(new_n15109_));
  NAND2_X1   g14107(.A1(new_n15109_), .A2(\A[552] ), .ZN(new_n15110_));
  INV_X1     g14108(.I(\A[552] ), .ZN(new_n15111_));
  NAND2_X1   g14109(.A1(new_n15111_), .A2(\A[551] ), .ZN(new_n15112_));
  AOI21_X1   g14110(.A1(new_n15110_), .A2(new_n15112_), .B(new_n15108_), .ZN(new_n15113_));
  NAND2_X1   g14111(.A1(\A[551] ), .A2(\A[552] ), .ZN(new_n15114_));
  NOR2_X1    g14112(.A1(\A[551] ), .A2(\A[552] ), .ZN(new_n15115_));
  INV_X1     g14113(.I(new_n15115_), .ZN(new_n15116_));
  AOI21_X1   g14114(.A1(new_n15116_), .A2(new_n15114_), .B(\A[550] ), .ZN(new_n15117_));
  NOR2_X1    g14115(.A1(new_n15117_), .A2(new_n15113_), .ZN(new_n15118_));
  NAND2_X1   g14116(.A1(new_n15107_), .A2(new_n15118_), .ZN(new_n15119_));
  NOR2_X1    g14117(.A1(new_n15100_), .A2(\A[548] ), .ZN(new_n15120_));
  NOR2_X1    g14118(.A1(new_n15098_), .A2(\A[549] ), .ZN(new_n15121_));
  OAI21_X1   g14119(.A1(new_n15120_), .A2(new_n15121_), .B(\A[547] ), .ZN(new_n15122_));
  INV_X1     g14120(.I(new_n15103_), .ZN(new_n15123_));
  OAI21_X1   g14121(.A1(new_n15123_), .A2(new_n15104_), .B(new_n15097_), .ZN(new_n15124_));
  NAND2_X1   g14122(.A1(new_n15122_), .A2(new_n15124_), .ZN(new_n15125_));
  NOR2_X1    g14123(.A1(new_n15111_), .A2(\A[551] ), .ZN(new_n15126_));
  NOR2_X1    g14124(.A1(new_n15109_), .A2(\A[552] ), .ZN(new_n15127_));
  OAI21_X1   g14125(.A1(new_n15126_), .A2(new_n15127_), .B(\A[550] ), .ZN(new_n15128_));
  INV_X1     g14126(.I(new_n15114_), .ZN(new_n15129_));
  OAI21_X1   g14127(.A1(new_n15129_), .A2(new_n15115_), .B(new_n15108_), .ZN(new_n15130_));
  NAND2_X1   g14128(.A1(new_n15128_), .A2(new_n15130_), .ZN(new_n15131_));
  NAND2_X1   g14129(.A1(new_n15125_), .A2(new_n15131_), .ZN(new_n15132_));
  NAND2_X1   g14130(.A1(new_n15119_), .A2(new_n15132_), .ZN(new_n15133_));
  NAND2_X1   g14131(.A1(new_n15096_), .A2(new_n15133_), .ZN(new_n15134_));
  NAND2_X1   g14132(.A1(new_n15088_), .A2(new_n15094_), .ZN(new_n15135_));
  NAND2_X1   g14133(.A1(new_n15070_), .A2(new_n15081_), .ZN(new_n15136_));
  NAND2_X1   g14134(.A1(new_n15135_), .A2(new_n15136_), .ZN(new_n15137_));
  NOR2_X1    g14135(.A1(new_n15125_), .A2(new_n15131_), .ZN(new_n15138_));
  NOR2_X1    g14136(.A1(new_n15107_), .A2(new_n15118_), .ZN(new_n15139_));
  NOR2_X1    g14137(.A1(new_n15139_), .A2(new_n15138_), .ZN(new_n15140_));
  NAND2_X1   g14138(.A1(new_n15140_), .A2(new_n15137_), .ZN(new_n15141_));
  NAND2_X1   g14139(.A1(new_n15134_), .A2(new_n15141_), .ZN(new_n15142_));
  INV_X1     g14140(.I(\A[543] ), .ZN(new_n15143_));
  NOR2_X1    g14141(.A1(new_n15143_), .A2(\A[542] ), .ZN(new_n15144_));
  INV_X1     g14142(.I(\A[542] ), .ZN(new_n15145_));
  NOR2_X1    g14143(.A1(new_n15145_), .A2(\A[543] ), .ZN(new_n15146_));
  OAI21_X1   g14144(.A1(new_n15144_), .A2(new_n15146_), .B(\A[541] ), .ZN(new_n15147_));
  INV_X1     g14145(.I(\A[541] ), .ZN(new_n15148_));
  NOR2_X1    g14146(.A1(\A[542] ), .A2(\A[543] ), .ZN(new_n15149_));
  NOR2_X1    g14147(.A1(new_n15145_), .A2(new_n15143_), .ZN(new_n15150_));
  OAI21_X1   g14148(.A1(new_n15150_), .A2(new_n15149_), .B(new_n15148_), .ZN(new_n15151_));
  INV_X1     g14149(.I(\A[546] ), .ZN(new_n15152_));
  NOR2_X1    g14150(.A1(new_n15152_), .A2(\A[545] ), .ZN(new_n15153_));
  INV_X1     g14151(.I(\A[545] ), .ZN(new_n15154_));
  NOR2_X1    g14152(.A1(new_n15154_), .A2(\A[546] ), .ZN(new_n15155_));
  OAI21_X1   g14153(.A1(new_n15153_), .A2(new_n15155_), .B(\A[544] ), .ZN(new_n15156_));
  INV_X1     g14154(.I(\A[544] ), .ZN(new_n15157_));
  NOR2_X1    g14155(.A1(\A[545] ), .A2(\A[546] ), .ZN(new_n15158_));
  NOR2_X1    g14156(.A1(new_n15154_), .A2(new_n15152_), .ZN(new_n15159_));
  OAI21_X1   g14157(.A1(new_n15159_), .A2(new_n15158_), .B(new_n15157_), .ZN(new_n15160_));
  NAND4_X1   g14158(.A1(new_n15147_), .A2(new_n15151_), .A3(new_n15160_), .A4(new_n15156_), .ZN(new_n15161_));
  NAND2_X1   g14159(.A1(new_n15151_), .A2(new_n15147_), .ZN(new_n15162_));
  NAND2_X1   g14160(.A1(new_n15160_), .A2(new_n15156_), .ZN(new_n15163_));
  NAND2_X1   g14161(.A1(new_n15162_), .A2(new_n15163_), .ZN(new_n15164_));
  INV_X1     g14162(.I(\A[535] ), .ZN(new_n15165_));
  INV_X1     g14163(.I(\A[536] ), .ZN(new_n15166_));
  NAND2_X1   g14164(.A1(new_n15166_), .A2(\A[537] ), .ZN(new_n15167_));
  INV_X1     g14165(.I(\A[537] ), .ZN(new_n15168_));
  NAND2_X1   g14166(.A1(new_n15168_), .A2(\A[536] ), .ZN(new_n15169_));
  AOI21_X1   g14167(.A1(new_n15167_), .A2(new_n15169_), .B(new_n15165_), .ZN(new_n15170_));
  NAND2_X1   g14168(.A1(\A[536] ), .A2(\A[537] ), .ZN(new_n15171_));
  NOR2_X1    g14169(.A1(\A[536] ), .A2(\A[537] ), .ZN(new_n15172_));
  INV_X1     g14170(.I(new_n15172_), .ZN(new_n15173_));
  AOI21_X1   g14171(.A1(new_n15173_), .A2(new_n15171_), .B(\A[535] ), .ZN(new_n15174_));
  INV_X1     g14172(.I(\A[538] ), .ZN(new_n15175_));
  INV_X1     g14173(.I(\A[539] ), .ZN(new_n15176_));
  NAND2_X1   g14174(.A1(new_n15176_), .A2(\A[540] ), .ZN(new_n15177_));
  INV_X1     g14175(.I(\A[540] ), .ZN(new_n15178_));
  NAND2_X1   g14176(.A1(new_n15178_), .A2(\A[539] ), .ZN(new_n15179_));
  AOI21_X1   g14177(.A1(new_n15177_), .A2(new_n15179_), .B(new_n15175_), .ZN(new_n15180_));
  NAND2_X1   g14178(.A1(\A[539] ), .A2(\A[540] ), .ZN(new_n15181_));
  NOR2_X1    g14179(.A1(\A[539] ), .A2(\A[540] ), .ZN(new_n15182_));
  INV_X1     g14180(.I(new_n15182_), .ZN(new_n15183_));
  AOI21_X1   g14181(.A1(new_n15183_), .A2(new_n15181_), .B(\A[538] ), .ZN(new_n15184_));
  NOR4_X1    g14182(.A1(new_n15170_), .A2(new_n15174_), .A3(new_n15184_), .A4(new_n15180_), .ZN(new_n15185_));
  INV_X1     g14183(.I(new_n15185_), .ZN(new_n15186_));
  OAI22_X1   g14184(.A1(new_n15170_), .A2(new_n15174_), .B1(new_n15184_), .B2(new_n15180_), .ZN(new_n15187_));
  NAND2_X1   g14185(.A1(new_n15186_), .A2(new_n15187_), .ZN(new_n15188_));
  NAND3_X1   g14186(.A1(new_n15188_), .A2(new_n15161_), .A3(new_n15164_), .ZN(new_n15189_));
  NAND2_X1   g14187(.A1(new_n15164_), .A2(new_n15161_), .ZN(new_n15190_));
  NOR2_X1    g14188(.A1(new_n15174_), .A2(new_n15170_), .ZN(new_n15191_));
  NOR2_X1    g14189(.A1(new_n15184_), .A2(new_n15180_), .ZN(new_n15192_));
  NOR2_X1    g14190(.A1(new_n15191_), .A2(new_n15192_), .ZN(new_n15193_));
  NOR2_X1    g14191(.A1(new_n15193_), .A2(new_n15185_), .ZN(new_n15194_));
  NAND2_X1   g14192(.A1(new_n15194_), .A2(new_n15190_), .ZN(new_n15195_));
  NAND2_X1   g14193(.A1(new_n15189_), .A2(new_n15195_), .ZN(new_n15196_));
  NAND2_X1   g14194(.A1(new_n15142_), .A2(new_n15196_), .ZN(new_n15197_));
  NAND4_X1   g14195(.A1(new_n15134_), .A2(new_n15189_), .A3(new_n15141_), .A4(new_n15195_), .ZN(new_n15198_));
  NAND2_X1   g14196(.A1(new_n15197_), .A2(new_n15198_), .ZN(new_n15199_));
  NAND4_X1   g14197(.A1(new_n15049_), .A2(new_n15050_), .A3(new_n15038_), .A4(new_n15042_), .ZN(new_n15200_));
  NAND2_X1   g14198(.A1(new_n15045_), .A2(new_n15200_), .ZN(new_n15201_));
  NOR2_X1    g14199(.A1(new_n15201_), .A2(new_n15199_), .ZN(new_n15202_));
  INV_X1     g14200(.I(new_n15202_), .ZN(new_n15203_));
  AOI21_X1   g14201(.A1(new_n15175_), .A2(new_n15181_), .B(new_n15182_), .ZN(new_n15204_));
  AOI21_X1   g14202(.A1(\A[536] ), .A2(\A[537] ), .B(\A[535] ), .ZN(new_n15205_));
  NOR2_X1    g14203(.A1(new_n15205_), .A2(new_n15172_), .ZN(new_n15206_));
  NOR2_X1    g14204(.A1(new_n15204_), .A2(new_n15206_), .ZN(new_n15207_));
  INV_X1     g14205(.I(new_n15207_), .ZN(new_n15208_));
  NAND2_X1   g14206(.A1(new_n15204_), .A2(new_n15206_), .ZN(new_n15209_));
  NAND2_X1   g14207(.A1(new_n15208_), .A2(new_n15209_), .ZN(new_n15210_));
  NOR2_X1    g14208(.A1(new_n15210_), .A2(new_n15185_), .ZN(new_n15211_));
  INV_X1     g14209(.I(new_n15209_), .ZN(new_n15212_));
  NOR2_X1    g14210(.A1(new_n15212_), .A2(new_n15207_), .ZN(new_n15213_));
  NOR2_X1    g14211(.A1(new_n15186_), .A2(new_n15213_), .ZN(new_n15214_));
  NOR2_X1    g14212(.A1(new_n15214_), .A2(new_n15211_), .ZN(new_n15215_));
  AOI21_X1   g14213(.A1(\A[545] ), .A2(\A[546] ), .B(\A[544] ), .ZN(new_n15216_));
  NOR2_X1    g14214(.A1(new_n15216_), .A2(new_n15158_), .ZN(new_n15217_));
  AOI21_X1   g14215(.A1(\A[542] ), .A2(\A[543] ), .B(\A[541] ), .ZN(new_n15218_));
  NOR2_X1    g14216(.A1(new_n15218_), .A2(new_n15149_), .ZN(new_n15219_));
  XNOR2_X1   g14217(.A1(new_n15217_), .A2(new_n15219_), .ZN(new_n15220_));
  XNOR2_X1   g14218(.A1(new_n15220_), .A2(new_n15161_), .ZN(new_n15221_));
  NAND3_X1   g14219(.A1(new_n15194_), .A2(new_n15161_), .A3(new_n15164_), .ZN(new_n15222_));
  AOI21_X1   g14220(.A1(new_n15221_), .A2(new_n15222_), .B(new_n15215_), .ZN(new_n15223_));
  XOR2_X1    g14221(.A1(new_n15220_), .A2(new_n15161_), .Z(new_n15224_));
  NOR2_X1    g14222(.A1(new_n15188_), .A2(new_n15190_), .ZN(new_n15225_));
  NAND2_X1   g14223(.A1(new_n15224_), .A2(new_n15225_), .ZN(new_n15226_));
  NAND2_X1   g14224(.A1(new_n15221_), .A2(new_n15222_), .ZN(new_n15227_));
  NAND2_X1   g14225(.A1(new_n15227_), .A2(new_n15226_), .ZN(new_n15228_));
  AOI22_X1   g14226(.A1(new_n15228_), .A2(new_n15215_), .B1(new_n15223_), .B2(new_n15226_), .ZN(new_n15229_));
  AOI21_X1   g14227(.A1(\A[551] ), .A2(\A[552] ), .B(\A[550] ), .ZN(new_n15230_));
  AOI21_X1   g14228(.A1(\A[548] ), .A2(\A[549] ), .B(\A[547] ), .ZN(new_n15231_));
  OAI22_X1   g14229(.A1(new_n15104_), .A2(new_n15231_), .B1(new_n15230_), .B2(new_n15115_), .ZN(new_n15232_));
  NOR4_X1    g14230(.A1(new_n15230_), .A2(new_n15231_), .A3(new_n15104_), .A4(new_n15115_), .ZN(new_n15233_));
  INV_X1     g14231(.I(new_n15233_), .ZN(new_n15234_));
  NAND2_X1   g14232(.A1(new_n15234_), .A2(new_n15232_), .ZN(new_n15235_));
  XOR2_X1    g14233(.A1(new_n15138_), .A2(new_n15235_), .Z(new_n15236_));
  AOI21_X1   g14234(.A1(new_n15076_), .A2(new_n15078_), .B(new_n15077_), .ZN(new_n15237_));
  AOI21_X1   g14235(.A1(\A[554] ), .A2(\A[555] ), .B(\A[553] ), .ZN(new_n15238_));
  NOR2_X1    g14236(.A1(new_n15238_), .A2(new_n15066_), .ZN(new_n15239_));
  XOR2_X1    g14237(.A1(new_n15237_), .A2(new_n15239_), .Z(new_n15240_));
  NOR2_X1    g14238(.A1(new_n15082_), .A2(new_n15240_), .ZN(new_n15241_));
  XNOR2_X1   g14239(.A1(new_n15237_), .A2(new_n15239_), .ZN(new_n15242_));
  NOR2_X1    g14240(.A1(new_n15135_), .A2(new_n15242_), .ZN(new_n15243_));
  OAI22_X1   g14241(.A1(new_n15137_), .A2(new_n15133_), .B1(new_n15243_), .B2(new_n15241_), .ZN(new_n15244_));
  NAND4_X1   g14242(.A1(new_n15140_), .A2(new_n15135_), .A3(new_n15136_), .A4(new_n15240_), .ZN(new_n15245_));
  NAND3_X1   g14243(.A1(new_n15244_), .A2(new_n15245_), .A3(new_n15236_), .ZN(new_n15246_));
  XOR2_X1    g14244(.A1(new_n15119_), .A2(new_n15235_), .Z(new_n15247_));
  NOR2_X1    g14245(.A1(new_n15243_), .A2(new_n15241_), .ZN(new_n15248_));
  NOR2_X1    g14246(.A1(new_n15137_), .A2(new_n15133_), .ZN(new_n15249_));
  NOR2_X1    g14247(.A1(new_n15249_), .A2(new_n15248_), .ZN(new_n15250_));
  INV_X1     g14248(.I(new_n15245_), .ZN(new_n15251_));
  OAI21_X1   g14249(.A1(new_n15250_), .A2(new_n15251_), .B(new_n15247_), .ZN(new_n15252_));
  AOI21_X1   g14250(.A1(new_n15252_), .A2(new_n15246_), .B(new_n15197_), .ZN(new_n15253_));
  AOI22_X1   g14251(.A1(new_n15134_), .A2(new_n15141_), .B1(new_n15189_), .B2(new_n15195_), .ZN(new_n15254_));
  INV_X1     g14252(.I(new_n15246_), .ZN(new_n15255_));
  AOI21_X1   g14253(.A1(new_n15244_), .A2(new_n15245_), .B(new_n15236_), .ZN(new_n15256_));
  NOR3_X1    g14254(.A1(new_n15255_), .A2(new_n15254_), .A3(new_n15256_), .ZN(new_n15257_));
  OAI21_X1   g14255(.A1(new_n15253_), .A2(new_n15257_), .B(new_n15229_), .ZN(new_n15258_));
  NAND2_X1   g14256(.A1(new_n15186_), .A2(new_n15213_), .ZN(new_n15259_));
  NAND2_X1   g14257(.A1(new_n15210_), .A2(new_n15185_), .ZN(new_n15260_));
  NAND2_X1   g14258(.A1(new_n15259_), .A2(new_n15260_), .ZN(new_n15261_));
  OAI21_X1   g14259(.A1(new_n15224_), .A2(new_n15225_), .B(new_n15261_), .ZN(new_n15262_));
  NOR2_X1    g14260(.A1(new_n15221_), .A2(new_n15222_), .ZN(new_n15263_));
  NOR2_X1    g14261(.A1(new_n15224_), .A2(new_n15225_), .ZN(new_n15264_));
  NOR2_X1    g14262(.A1(new_n15263_), .A2(new_n15264_), .ZN(new_n15265_));
  OAI22_X1   g14263(.A1(new_n15265_), .A2(new_n15261_), .B1(new_n15262_), .B2(new_n15263_), .ZN(new_n15266_));
  OAI21_X1   g14264(.A1(new_n15255_), .A2(new_n15256_), .B(new_n15254_), .ZN(new_n15267_));
  NAND3_X1   g14265(.A1(new_n15252_), .A2(new_n15197_), .A3(new_n15246_), .ZN(new_n15268_));
  NAND3_X1   g14266(.A1(new_n15266_), .A2(new_n15267_), .A3(new_n15268_), .ZN(new_n15269_));
  AOI21_X1   g14267(.A1(new_n15258_), .A2(new_n15269_), .B(new_n15203_), .ZN(new_n15270_));
  NAND3_X1   g14268(.A1(new_n15203_), .A2(new_n15258_), .A3(new_n15269_), .ZN(new_n15271_));
  OAI21_X1   g14269(.A1(new_n15270_), .A2(new_n15059_), .B(new_n15271_), .ZN(new_n15272_));
  OR2_X2     g14270(.A1(new_n14942_), .A2(new_n14927_), .Z(new_n15273_));
  INV_X1     g14271(.I(new_n14948_), .ZN(new_n15274_));
  NAND2_X1   g14272(.A1(new_n15274_), .A2(new_n15037_), .ZN(new_n15275_));
  AOI21_X1   g14273(.A1(new_n15273_), .A2(new_n15275_), .B(new_n14900_), .ZN(new_n15276_));
  NAND2_X1   g14274(.A1(new_n14924_), .A2(new_n14925_), .ZN(new_n15277_));
  NOR2_X1    g14275(.A1(new_n14924_), .A2(new_n14925_), .ZN(new_n15278_));
  AOI21_X1   g14276(.A1(new_n14940_), .A2(new_n15277_), .B(new_n15278_), .ZN(new_n15279_));
  INV_X1     g14277(.I(new_n14898_), .ZN(new_n15280_));
  AOI21_X1   g14278(.A1(new_n14892_), .A2(new_n15280_), .B(new_n14897_), .ZN(new_n15281_));
  NOR2_X1    g14279(.A1(new_n15279_), .A2(new_n15281_), .ZN(new_n15282_));
  NAND2_X1   g14280(.A1(new_n15279_), .A2(new_n15281_), .ZN(new_n15283_));
  INV_X1     g14281(.I(new_n15283_), .ZN(new_n15284_));
  NOR2_X1    g14282(.A1(new_n15284_), .A2(new_n15282_), .ZN(new_n15285_));
  OAI21_X1   g14283(.A1(new_n15276_), .A2(new_n14951_), .B(new_n15285_), .ZN(new_n15286_));
  INV_X1     g14284(.I(new_n14900_), .ZN(new_n15287_));
  AOI21_X1   g14285(.A1(new_n14949_), .A2(new_n15287_), .B(new_n14951_), .ZN(new_n15288_));
  INV_X1     g14286(.I(new_n15282_), .ZN(new_n15289_));
  NAND2_X1   g14287(.A1(new_n15289_), .A2(new_n15283_), .ZN(new_n15290_));
  NAND2_X1   g14288(.A1(new_n15288_), .A2(new_n15290_), .ZN(new_n15291_));
  NAND2_X1   g14289(.A1(new_n15286_), .A2(new_n15291_), .ZN(new_n15292_));
  AND2_X2    g14290(.A1(new_n15005_), .A2(new_n15006_), .Z(new_n15293_));
  NOR2_X1    g14291(.A1(new_n15005_), .A2(new_n15006_), .ZN(new_n15294_));
  INV_X1     g14292(.I(new_n15294_), .ZN(new_n15295_));
  OAI21_X1   g14293(.A1(new_n15004_), .A2(new_n15293_), .B(new_n15295_), .ZN(new_n15296_));
  OR2_X2     g14294(.A1(new_n15023_), .A2(new_n15008_), .Z(new_n15297_));
  INV_X1     g14295(.I(new_n15028_), .ZN(new_n15298_));
  NAND2_X1   g14296(.A1(new_n15298_), .A2(new_n15041_), .ZN(new_n15299_));
  AOI21_X1   g14297(.A1(new_n15297_), .A2(new_n15299_), .B(new_n14981_), .ZN(new_n15300_));
  NOR2_X1    g14298(.A1(new_n14978_), .A2(new_n14979_), .ZN(new_n15301_));
  NAND2_X1   g14299(.A1(new_n14978_), .A2(new_n14979_), .ZN(new_n15302_));
  AOI21_X1   g14300(.A1(new_n15026_), .A2(new_n15302_), .B(new_n15301_), .ZN(new_n15303_));
  NOR3_X1    g14301(.A1(new_n15300_), .A2(new_n15032_), .A3(new_n15303_), .ZN(new_n15304_));
  AOI21_X1   g14302(.A1(new_n15029_), .A2(new_n15034_), .B(new_n15032_), .ZN(new_n15305_));
  INV_X1     g14303(.I(new_n15303_), .ZN(new_n15306_));
  NOR2_X1    g14304(.A1(new_n15305_), .A2(new_n15306_), .ZN(new_n15307_));
  NOR3_X1    g14305(.A1(new_n15304_), .A2(new_n15307_), .A3(new_n15296_), .ZN(new_n15308_));
  INV_X1     g14306(.I(new_n15296_), .ZN(new_n15309_));
  NAND2_X1   g14307(.A1(new_n15305_), .A2(new_n15306_), .ZN(new_n15310_));
  OAI21_X1   g14308(.A1(new_n15300_), .A2(new_n15032_), .B(new_n15303_), .ZN(new_n15311_));
  AOI21_X1   g14309(.A1(new_n15311_), .A2(new_n15310_), .B(new_n15309_), .ZN(new_n15312_));
  OAI21_X1   g14310(.A1(new_n15308_), .A2(new_n15312_), .B(new_n15292_), .ZN(new_n15313_));
  NOR2_X1    g14311(.A1(new_n15288_), .A2(new_n15290_), .ZN(new_n15314_));
  NOR3_X1    g14312(.A1(new_n15276_), .A2(new_n15285_), .A3(new_n14951_), .ZN(new_n15315_));
  NOR2_X1    g14313(.A1(new_n15315_), .A2(new_n15314_), .ZN(new_n15316_));
  NAND3_X1   g14314(.A1(new_n15311_), .A2(new_n15310_), .A3(new_n15309_), .ZN(new_n15317_));
  OAI21_X1   g14315(.A1(new_n15304_), .A2(new_n15307_), .B(new_n15296_), .ZN(new_n15318_));
  NAND3_X1   g14316(.A1(new_n15317_), .A2(new_n15318_), .A3(new_n15316_), .ZN(new_n15319_));
  OAI21_X1   g14317(.A1(new_n15055_), .A2(new_n15046_), .B(new_n15057_), .ZN(new_n15320_));
  NAND3_X1   g14318(.A1(new_n15313_), .A2(new_n15319_), .A3(new_n15320_), .ZN(new_n15321_));
  AOI21_X1   g14319(.A1(new_n15318_), .A2(new_n15317_), .B(new_n15316_), .ZN(new_n15322_));
  NOR3_X1    g14320(.A1(new_n15308_), .A2(new_n15312_), .A3(new_n15292_), .ZN(new_n15323_));
  AOI21_X1   g14321(.A1(new_n14956_), .A2(new_n15056_), .B(new_n15052_), .ZN(new_n15324_));
  OAI21_X1   g14322(.A1(new_n15323_), .A2(new_n15322_), .B(new_n15324_), .ZN(new_n15325_));
  OAI21_X1   g14323(.A1(new_n15253_), .A2(new_n15229_), .B(new_n15268_), .ZN(new_n15326_));
  OR2_X2     g14324(.A1(new_n15243_), .A2(new_n15241_), .Z(new_n15327_));
  NAND2_X1   g14325(.A1(new_n15140_), .A2(new_n15096_), .ZN(new_n15328_));
  AOI21_X1   g14326(.A1(new_n15327_), .A2(new_n15328_), .B(new_n15236_), .ZN(new_n15329_));
  INV_X1     g14327(.I(new_n15237_), .ZN(new_n15330_));
  INV_X1     g14328(.I(new_n15239_), .ZN(new_n15331_));
  NOR2_X1    g14329(.A1(new_n15330_), .A2(new_n15331_), .ZN(new_n15332_));
  INV_X1     g14330(.I(new_n15332_), .ZN(new_n15333_));
  NOR2_X1    g14331(.A1(new_n15237_), .A2(new_n15239_), .ZN(new_n15334_));
  AOI21_X1   g14332(.A1(new_n15135_), .A2(new_n15333_), .B(new_n15334_), .ZN(new_n15335_));
  INV_X1     g14333(.I(new_n15232_), .ZN(new_n15336_));
  AOI21_X1   g14334(.A1(new_n15119_), .A2(new_n15234_), .B(new_n15336_), .ZN(new_n15337_));
  NOR2_X1    g14335(.A1(new_n15335_), .A2(new_n15337_), .ZN(new_n15338_));
  INV_X1     g14336(.I(new_n15334_), .ZN(new_n15339_));
  OAI21_X1   g14337(.A1(new_n15082_), .A2(new_n15332_), .B(new_n15339_), .ZN(new_n15340_));
  OAI21_X1   g14338(.A1(new_n15138_), .A2(new_n15233_), .B(new_n15232_), .ZN(new_n15341_));
  NOR2_X1    g14339(.A1(new_n15340_), .A2(new_n15341_), .ZN(new_n15342_));
  NOR2_X1    g14340(.A1(new_n15338_), .A2(new_n15342_), .ZN(new_n15343_));
  OAI21_X1   g14341(.A1(new_n15329_), .A2(new_n15251_), .B(new_n15343_), .ZN(new_n15344_));
  NAND2_X1   g14342(.A1(new_n15244_), .A2(new_n15247_), .ZN(new_n15345_));
  NAND2_X1   g14343(.A1(new_n15340_), .A2(new_n15341_), .ZN(new_n15346_));
  NAND2_X1   g14344(.A1(new_n15335_), .A2(new_n15337_), .ZN(new_n15347_));
  NAND2_X1   g14345(.A1(new_n15347_), .A2(new_n15346_), .ZN(new_n15348_));
  NAND3_X1   g14346(.A1(new_n15345_), .A2(new_n15348_), .A3(new_n15245_), .ZN(new_n15349_));
  NAND2_X1   g14347(.A1(new_n15344_), .A2(new_n15349_), .ZN(new_n15350_));
  NOR4_X1    g14348(.A1(new_n15216_), .A2(new_n15218_), .A3(new_n15149_), .A4(new_n15158_), .ZN(new_n15351_));
  INV_X1     g14349(.I(new_n15351_), .ZN(new_n15352_));
  NOR2_X1    g14350(.A1(new_n15217_), .A2(new_n15219_), .ZN(new_n15353_));
  AOI21_X1   g14351(.A1(new_n15161_), .A2(new_n15352_), .B(new_n15353_), .ZN(new_n15354_));
  INV_X1     g14352(.I(new_n15354_), .ZN(new_n15355_));
  AOI21_X1   g14353(.A1(new_n15186_), .A2(new_n15209_), .B(new_n15207_), .ZN(new_n15356_));
  NOR3_X1    g14354(.A1(new_n15223_), .A2(new_n15263_), .A3(new_n15356_), .ZN(new_n15357_));
  INV_X1     g14355(.I(new_n15356_), .ZN(new_n15358_));
  AOI21_X1   g14356(.A1(new_n15262_), .A2(new_n15226_), .B(new_n15358_), .ZN(new_n15359_));
  NOR3_X1    g14357(.A1(new_n15357_), .A2(new_n15359_), .A3(new_n15355_), .ZN(new_n15360_));
  NAND3_X1   g14358(.A1(new_n15262_), .A2(new_n15226_), .A3(new_n15358_), .ZN(new_n15361_));
  OAI21_X1   g14359(.A1(new_n15223_), .A2(new_n15263_), .B(new_n15356_), .ZN(new_n15362_));
  AOI21_X1   g14360(.A1(new_n15362_), .A2(new_n15361_), .B(new_n15354_), .ZN(new_n15363_));
  OAI21_X1   g14361(.A1(new_n15363_), .A2(new_n15360_), .B(new_n15350_), .ZN(new_n15364_));
  AOI21_X1   g14362(.A1(new_n15345_), .A2(new_n15245_), .B(new_n15348_), .ZN(new_n15365_));
  NOR3_X1    g14363(.A1(new_n15329_), .A2(new_n15251_), .A3(new_n15343_), .ZN(new_n15366_));
  NOR2_X1    g14364(.A1(new_n15366_), .A2(new_n15365_), .ZN(new_n15367_));
  NAND3_X1   g14365(.A1(new_n15362_), .A2(new_n15361_), .A3(new_n15354_), .ZN(new_n15368_));
  OAI21_X1   g14366(.A1(new_n15357_), .A2(new_n15359_), .B(new_n15355_), .ZN(new_n15369_));
  NAND3_X1   g14367(.A1(new_n15367_), .A2(new_n15369_), .A3(new_n15368_), .ZN(new_n15370_));
  NAND3_X1   g14368(.A1(new_n15364_), .A2(new_n15370_), .A3(new_n15326_), .ZN(new_n15371_));
  AOI21_X1   g14369(.A1(new_n15266_), .A2(new_n15267_), .B(new_n15257_), .ZN(new_n15372_));
  AOI21_X1   g14370(.A1(new_n15368_), .A2(new_n15369_), .B(new_n15367_), .ZN(new_n15373_));
  NOR3_X1    g14371(.A1(new_n15360_), .A2(new_n15363_), .A3(new_n15350_), .ZN(new_n15374_));
  OAI21_X1   g14372(.A1(new_n15373_), .A2(new_n15374_), .B(new_n15372_), .ZN(new_n15375_));
  NAND4_X1   g14373(.A1(new_n15325_), .A2(new_n15321_), .A3(new_n15375_), .A4(new_n15371_), .ZN(new_n15376_));
  NOR3_X1    g14374(.A1(new_n15323_), .A2(new_n15322_), .A3(new_n15324_), .ZN(new_n15377_));
  AOI21_X1   g14375(.A1(new_n15313_), .A2(new_n15319_), .B(new_n15320_), .ZN(new_n15378_));
  NOR3_X1    g14376(.A1(new_n15373_), .A2(new_n15374_), .A3(new_n15372_), .ZN(new_n15379_));
  AOI21_X1   g14377(.A1(new_n15364_), .A2(new_n15370_), .B(new_n15326_), .ZN(new_n15380_));
  OAI22_X1   g14378(.A1(new_n15378_), .A2(new_n15377_), .B1(new_n15379_), .B2(new_n15380_), .ZN(new_n15381_));
  NAND3_X1   g14379(.A1(new_n15381_), .A2(new_n15376_), .A3(new_n15272_), .ZN(new_n15382_));
  OR2_X2     g14380(.A1(new_n15058_), .A2(new_n15053_), .Z(new_n15383_));
  AOI21_X1   g14381(.A1(new_n15267_), .A2(new_n15268_), .B(new_n15266_), .ZN(new_n15384_));
  NOR3_X1    g14382(.A1(new_n15253_), .A2(new_n15229_), .A3(new_n15257_), .ZN(new_n15385_));
  OAI21_X1   g14383(.A1(new_n15384_), .A2(new_n15385_), .B(new_n15202_), .ZN(new_n15386_));
  NOR3_X1    g14384(.A1(new_n15384_), .A2(new_n15385_), .A3(new_n15202_), .ZN(new_n15387_));
  AOI21_X1   g14385(.A1(new_n15383_), .A2(new_n15386_), .B(new_n15387_), .ZN(new_n15388_));
  NOR4_X1    g14386(.A1(new_n15378_), .A2(new_n15377_), .A3(new_n15379_), .A4(new_n15380_), .ZN(new_n15389_));
  AOI22_X1   g14387(.A1(new_n15325_), .A2(new_n15321_), .B1(new_n15375_), .B2(new_n15371_), .ZN(new_n15390_));
  OAI21_X1   g14388(.A1(new_n15389_), .A2(new_n15390_), .B(new_n15388_), .ZN(new_n15391_));
  NAND4_X1   g14389(.A1(new_n14871_), .A2(new_n14862_), .A3(new_n15391_), .A4(new_n15382_), .ZN(new_n15392_));
  AOI22_X1   g14390(.A1(new_n14871_), .A2(new_n14862_), .B1(new_n15391_), .B2(new_n15382_), .ZN(new_n15393_));
  NAND3_X1   g14391(.A1(new_n14856_), .A2(new_n14869_), .A3(new_n14859_), .ZN(new_n15394_));
  OAI21_X1   g14392(.A1(new_n14867_), .A2(new_n14860_), .B(new_n14868_), .ZN(new_n15395_));
  NAND2_X1   g14393(.A1(new_n14850_), .A2(new_n14575_), .ZN(new_n15396_));
  OAI21_X1   g14394(.A1(new_n14755_), .A2(new_n14853_), .B(new_n15396_), .ZN(new_n15397_));
  NAND2_X1   g14395(.A1(new_n15397_), .A2(new_n14855_), .ZN(new_n15398_));
  NAND2_X1   g14396(.A1(new_n15201_), .A2(new_n15199_), .ZN(new_n15399_));
  NAND2_X1   g14397(.A1(new_n15203_), .A2(new_n15399_), .ZN(new_n15400_));
  NOR2_X1    g14398(.A1(new_n15400_), .A2(new_n15398_), .ZN(new_n15401_));
  AOI21_X1   g14399(.A1(new_n15395_), .A2(new_n15394_), .B(new_n15401_), .ZN(new_n15402_));
  NOR2_X1    g14400(.A1(new_n15270_), .A2(new_n15059_), .ZN(new_n15403_));
  NAND2_X1   g14401(.A1(new_n15386_), .A2(new_n15271_), .ZN(new_n15404_));
  AOI22_X1   g14402(.A1(new_n15403_), .A2(new_n15271_), .B1(new_n15404_), .B2(new_n15059_), .ZN(new_n15405_));
  NAND3_X1   g14403(.A1(new_n15395_), .A2(new_n15394_), .A3(new_n15401_), .ZN(new_n15406_));
  AOI21_X1   g14404(.A1(new_n15405_), .A2(new_n15406_), .B(new_n15402_), .ZN(new_n15407_));
  OAI21_X1   g14405(.A1(new_n15393_), .A2(new_n15407_), .B(new_n15392_), .ZN(new_n15408_));
  OAI21_X1   g14406(.A1(new_n15390_), .A2(new_n15388_), .B(new_n15376_), .ZN(new_n15409_));
  NOR2_X1    g14407(.A1(new_n15373_), .A2(new_n15326_), .ZN(new_n15410_));
  NAND2_X1   g14408(.A1(new_n15362_), .A2(new_n15355_), .ZN(new_n15411_));
  NAND2_X1   g14409(.A1(new_n15345_), .A2(new_n15245_), .ZN(new_n15412_));
  OAI21_X1   g14410(.A1(new_n15412_), .A2(new_n15342_), .B(new_n15346_), .ZN(new_n15413_));
  AOI21_X1   g14411(.A1(new_n15361_), .A2(new_n15411_), .B(new_n15413_), .ZN(new_n15414_));
  NAND2_X1   g14412(.A1(new_n15411_), .A2(new_n15361_), .ZN(new_n15415_));
  NOR2_X1    g14413(.A1(new_n15329_), .A2(new_n15251_), .ZN(new_n15416_));
  AOI21_X1   g14414(.A1(new_n15416_), .A2(new_n15347_), .B(new_n15338_), .ZN(new_n15417_));
  NOR2_X1    g14415(.A1(new_n15415_), .A2(new_n15417_), .ZN(new_n15418_));
  NOR2_X1    g14416(.A1(new_n15418_), .A2(new_n15414_), .ZN(new_n15419_));
  OAI21_X1   g14417(.A1(new_n15410_), .A2(new_n15374_), .B(new_n15419_), .ZN(new_n15420_));
  NAND2_X1   g14418(.A1(new_n15364_), .A2(new_n15372_), .ZN(new_n15421_));
  NAND2_X1   g14419(.A1(new_n15415_), .A2(new_n15417_), .ZN(new_n15422_));
  NAND3_X1   g14420(.A1(new_n15413_), .A2(new_n15411_), .A3(new_n15361_), .ZN(new_n15423_));
  NAND2_X1   g14421(.A1(new_n15422_), .A2(new_n15423_), .ZN(new_n15424_));
  NAND3_X1   g14422(.A1(new_n15424_), .A2(new_n15421_), .A3(new_n15370_), .ZN(new_n15425_));
  NOR2_X1    g14423(.A1(new_n15322_), .A2(new_n15320_), .ZN(new_n15426_));
  OAI21_X1   g14424(.A1(new_n15305_), .A2(new_n15306_), .B(new_n15296_), .ZN(new_n15427_));
  NAND2_X1   g14425(.A1(new_n15427_), .A2(new_n15310_), .ZN(new_n15428_));
  AOI21_X1   g14426(.A1(new_n15288_), .A2(new_n15283_), .B(new_n15282_), .ZN(new_n15429_));
  XOR2_X1    g14427(.A1(new_n15428_), .A2(new_n15429_), .Z(new_n15430_));
  OAI21_X1   g14428(.A1(new_n15426_), .A2(new_n15323_), .B(new_n15430_), .ZN(new_n15431_));
  NAND2_X1   g14429(.A1(new_n15313_), .A2(new_n15324_), .ZN(new_n15432_));
  NAND2_X1   g14430(.A1(new_n15428_), .A2(new_n15429_), .ZN(new_n15433_));
  INV_X1     g14431(.I(new_n15429_), .ZN(new_n15434_));
  NAND3_X1   g14432(.A1(new_n15434_), .A2(new_n15310_), .A3(new_n15427_), .ZN(new_n15435_));
  NAND2_X1   g14433(.A1(new_n15435_), .A2(new_n15433_), .ZN(new_n15436_));
  NAND3_X1   g14434(.A1(new_n15432_), .A2(new_n15319_), .A3(new_n15436_), .ZN(new_n15437_));
  NAND4_X1   g14435(.A1(new_n15420_), .A2(new_n15431_), .A3(new_n15437_), .A4(new_n15425_), .ZN(new_n15438_));
  AOI21_X1   g14436(.A1(new_n15370_), .A2(new_n15421_), .B(new_n15424_), .ZN(new_n15439_));
  NOR3_X1    g14437(.A1(new_n15419_), .A2(new_n15410_), .A3(new_n15374_), .ZN(new_n15440_));
  AOI21_X1   g14438(.A1(new_n15432_), .A2(new_n15319_), .B(new_n15436_), .ZN(new_n15441_));
  NOR3_X1    g14439(.A1(new_n15426_), .A2(new_n15430_), .A3(new_n15323_), .ZN(new_n15442_));
  OAI22_X1   g14440(.A1(new_n15439_), .A2(new_n15440_), .B1(new_n15442_), .B2(new_n15441_), .ZN(new_n15443_));
  NAND3_X1   g14441(.A1(new_n15409_), .A2(new_n15443_), .A3(new_n15438_), .ZN(new_n15444_));
  AOI21_X1   g14442(.A1(new_n15272_), .A2(new_n15381_), .B(new_n15389_), .ZN(new_n15445_));
  NOR4_X1    g14443(.A1(new_n15439_), .A2(new_n15440_), .A3(new_n15442_), .A4(new_n15441_), .ZN(new_n15446_));
  AOI22_X1   g14444(.A1(new_n15420_), .A2(new_n15425_), .B1(new_n15431_), .B2(new_n15437_), .ZN(new_n15447_));
  OAI21_X1   g14445(.A1(new_n15446_), .A2(new_n15447_), .B(new_n15445_), .ZN(new_n15448_));
  OAI21_X1   g14446(.A1(new_n14864_), .A2(new_n14870_), .B(new_n14841_), .ZN(new_n15449_));
  NOR2_X1    g14447(.A1(new_n14838_), .A2(new_n14779_), .ZN(new_n15450_));
  NAND2_X1   g14448(.A1(new_n14820_), .A2(new_n14808_), .ZN(new_n15451_));
  AOI21_X1   g14449(.A1(new_n14799_), .A2(new_n14801_), .B(new_n14792_), .ZN(new_n15452_));
  INV_X1     g14450(.I(new_n15452_), .ZN(new_n15453_));
  AOI21_X1   g14451(.A1(new_n15451_), .A2(new_n14819_), .B(new_n15453_), .ZN(new_n15454_));
  NOR2_X1    g14452(.A1(new_n14816_), .A2(new_n14818_), .ZN(new_n15455_));
  NOR3_X1    g14453(.A1(new_n15455_), .A2(new_n14813_), .A3(new_n15452_), .ZN(new_n15456_));
  NOR2_X1    g14454(.A1(new_n15454_), .A2(new_n15456_), .ZN(new_n15457_));
  OAI21_X1   g14455(.A1(new_n15450_), .A2(new_n14839_), .B(new_n15457_), .ZN(new_n15458_));
  NAND2_X1   g14456(.A1(new_n14822_), .A2(new_n14837_), .ZN(new_n15459_));
  OAI21_X1   g14457(.A1(new_n15455_), .A2(new_n14813_), .B(new_n15452_), .ZN(new_n15460_));
  NAND3_X1   g14458(.A1(new_n15451_), .A2(new_n15453_), .A3(new_n14819_), .ZN(new_n15461_));
  NAND2_X1   g14459(.A1(new_n15461_), .A2(new_n15460_), .ZN(new_n15462_));
  NAND3_X1   g14460(.A1(new_n15459_), .A2(new_n14828_), .A3(new_n15462_), .ZN(new_n15463_));
  NAND2_X1   g14461(.A1(new_n14566_), .A2(new_n14565_), .ZN(new_n15464_));
  AOI21_X1   g14462(.A1(new_n15464_), .A2(new_n14451_), .B(new_n14583_), .ZN(new_n15465_));
  NAND2_X1   g14463(.A1(new_n14561_), .A2(new_n14481_), .ZN(new_n15466_));
  AOI21_X1   g14464(.A1(new_n14446_), .A2(new_n14448_), .B(new_n14435_), .ZN(new_n15467_));
  INV_X1     g14465(.I(new_n15467_), .ZN(new_n15468_));
  AOI21_X1   g14466(.A1(new_n14560_), .A2(new_n15466_), .B(new_n15468_), .ZN(new_n15469_));
  NOR2_X1    g14467(.A1(new_n14557_), .A2(new_n14559_), .ZN(new_n15470_));
  NOR3_X1    g14468(.A1(new_n15470_), .A2(new_n14543_), .A3(new_n15467_), .ZN(new_n15471_));
  NOR2_X1    g14469(.A1(new_n15469_), .A2(new_n15471_), .ZN(new_n15472_));
  OAI21_X1   g14470(.A1(new_n15465_), .A2(new_n14586_), .B(new_n15472_), .ZN(new_n15473_));
  NAND2_X1   g14471(.A1(new_n14563_), .A2(new_n14597_), .ZN(new_n15474_));
  OAI21_X1   g14472(.A1(new_n15470_), .A2(new_n14543_), .B(new_n15467_), .ZN(new_n15475_));
  NAND3_X1   g14473(.A1(new_n15468_), .A2(new_n15466_), .A3(new_n14560_), .ZN(new_n15476_));
  NAND2_X1   g14474(.A1(new_n15476_), .A2(new_n15475_), .ZN(new_n15477_));
  NAND3_X1   g14475(.A1(new_n15474_), .A2(new_n14567_), .A3(new_n15477_), .ZN(new_n15478_));
  NAND4_X1   g14476(.A1(new_n15458_), .A2(new_n15463_), .A3(new_n15473_), .A4(new_n15478_), .ZN(new_n15479_));
  AOI21_X1   g14477(.A1(new_n15459_), .A2(new_n14828_), .B(new_n15462_), .ZN(new_n15480_));
  NOR3_X1    g14478(.A1(new_n15450_), .A2(new_n14839_), .A3(new_n15457_), .ZN(new_n15481_));
  AOI21_X1   g14479(.A1(new_n15474_), .A2(new_n14567_), .B(new_n15477_), .ZN(new_n15482_));
  NOR3_X1    g14480(.A1(new_n15465_), .A2(new_n15472_), .A3(new_n14586_), .ZN(new_n15483_));
  OAI22_X1   g14481(.A1(new_n15480_), .A2(new_n15481_), .B1(new_n15482_), .B2(new_n15483_), .ZN(new_n15484_));
  NAND3_X1   g14482(.A1(new_n15449_), .A2(new_n15479_), .A3(new_n15484_), .ZN(new_n15485_));
  AOI21_X1   g14483(.A1(new_n14846_), .A2(new_n14861_), .B(new_n14863_), .ZN(new_n15486_));
  NAND2_X1   g14484(.A1(new_n15484_), .A2(new_n15479_), .ZN(new_n15487_));
  NAND2_X1   g14485(.A1(new_n15487_), .A2(new_n15486_), .ZN(new_n15488_));
  NAND4_X1   g14486(.A1(new_n15488_), .A2(new_n15448_), .A3(new_n15444_), .A4(new_n15485_), .ZN(new_n15489_));
  NOR3_X1    g14487(.A1(new_n15445_), .A2(new_n15446_), .A3(new_n15447_), .ZN(new_n15490_));
  AOI21_X1   g14488(.A1(new_n15438_), .A2(new_n15443_), .B(new_n15409_), .ZN(new_n15491_));
  NOR4_X1    g14489(.A1(new_n15480_), .A2(new_n15481_), .A3(new_n15483_), .A4(new_n15482_), .ZN(new_n15492_));
  AOI22_X1   g14490(.A1(new_n15458_), .A2(new_n15463_), .B1(new_n15473_), .B2(new_n15478_), .ZN(new_n15493_));
  NOR3_X1    g14491(.A1(new_n15486_), .A2(new_n15492_), .A3(new_n15493_), .ZN(new_n15494_));
  AOI21_X1   g14492(.A1(new_n15479_), .A2(new_n15484_), .B(new_n15449_), .ZN(new_n15495_));
  OAI22_X1   g14493(.A1(new_n15494_), .A2(new_n15495_), .B1(new_n15491_), .B2(new_n15490_), .ZN(new_n15496_));
  NAND3_X1   g14494(.A1(new_n15408_), .A2(new_n15496_), .A3(new_n15489_), .ZN(new_n15497_));
  NOR3_X1    g14495(.A1(new_n14864_), .A2(new_n14863_), .A3(new_n14870_), .ZN(new_n15498_));
  AOI21_X1   g14496(.A1(new_n14846_), .A2(new_n14841_), .B(new_n14861_), .ZN(new_n15499_));
  NOR3_X1    g14497(.A1(new_n15389_), .A2(new_n15390_), .A3(new_n15388_), .ZN(new_n15500_));
  AOI21_X1   g14498(.A1(new_n15381_), .A2(new_n15376_), .B(new_n15272_), .ZN(new_n15501_));
  NOR4_X1    g14499(.A1(new_n15498_), .A2(new_n15499_), .A3(new_n15500_), .A4(new_n15501_), .ZN(new_n15502_));
  OAI22_X1   g14500(.A1(new_n15498_), .A2(new_n15499_), .B1(new_n15500_), .B2(new_n15501_), .ZN(new_n15503_));
  NOR3_X1    g14501(.A1(new_n14868_), .A2(new_n14860_), .A3(new_n14867_), .ZN(new_n15504_));
  AOI21_X1   g14502(.A1(new_n14856_), .A2(new_n14869_), .B(new_n14859_), .ZN(new_n15505_));
  INV_X1     g14503(.I(new_n15401_), .ZN(new_n15506_));
  OAI21_X1   g14504(.A1(new_n15504_), .A2(new_n15505_), .B(new_n15506_), .ZN(new_n15507_));
  NAND2_X1   g14505(.A1(new_n15404_), .A2(new_n15059_), .ZN(new_n15508_));
  NAND2_X1   g14506(.A1(new_n15403_), .A2(new_n15271_), .ZN(new_n15509_));
  NAND2_X1   g14507(.A1(new_n15509_), .A2(new_n15508_), .ZN(new_n15510_));
  NOR3_X1    g14508(.A1(new_n15504_), .A2(new_n15505_), .A3(new_n15506_), .ZN(new_n15511_));
  OAI21_X1   g14509(.A1(new_n15510_), .A2(new_n15511_), .B(new_n15507_), .ZN(new_n15512_));
  AOI21_X1   g14510(.A1(new_n15503_), .A2(new_n15512_), .B(new_n15502_), .ZN(new_n15513_));
  NOR4_X1    g14511(.A1(new_n15494_), .A2(new_n15495_), .A3(new_n15491_), .A4(new_n15490_), .ZN(new_n15514_));
  AOI22_X1   g14512(.A1(new_n15485_), .A2(new_n15488_), .B1(new_n15448_), .B2(new_n15444_), .ZN(new_n15515_));
  OAI21_X1   g14513(.A1(new_n15515_), .A2(new_n15514_), .B(new_n15513_), .ZN(new_n15516_));
  NAND4_X1   g14514(.A1(new_n14330_), .A2(new_n15516_), .A3(new_n14315_), .A4(new_n15497_), .ZN(new_n15517_));
  NAND3_X1   g14515(.A1(new_n15503_), .A2(new_n15392_), .A3(new_n15512_), .ZN(new_n15518_));
  OAI21_X1   g14516(.A1(new_n15502_), .A2(new_n15393_), .B(new_n15407_), .ZN(new_n15519_));
  NAND3_X1   g14517(.A1(new_n14326_), .A2(new_n14225_), .A3(new_n14320_), .ZN(new_n15520_));
  OAI21_X1   g14518(.A1(new_n14325_), .A2(new_n14226_), .B(new_n13999_), .ZN(new_n15521_));
  NAND4_X1   g14519(.A1(new_n15519_), .A2(new_n15521_), .A3(new_n15520_), .A4(new_n15518_), .ZN(new_n15522_));
  AOI22_X1   g14520(.A1(new_n15520_), .A2(new_n15521_), .B1(new_n15519_), .B2(new_n15518_), .ZN(new_n15523_));
  NAND3_X1   g14521(.A1(new_n15510_), .A2(new_n15406_), .A3(new_n15507_), .ZN(new_n15524_));
  OAI21_X1   g14522(.A1(new_n15402_), .A2(new_n15511_), .B(new_n15405_), .ZN(new_n15525_));
  NAND2_X1   g14523(.A1(new_n15400_), .A2(new_n15398_), .ZN(new_n15526_));
  NAND2_X1   g14524(.A1(new_n15506_), .A2(new_n15526_), .ZN(new_n15527_));
  NOR2_X1    g14525(.A1(new_n13874_), .A2(new_n13872_), .ZN(new_n15528_));
  NOR3_X1    g14526(.A1(new_n15527_), .A2(new_n13876_), .A3(new_n15528_), .ZN(new_n15529_));
  AOI21_X1   g14527(.A1(new_n15524_), .A2(new_n15525_), .B(new_n15529_), .ZN(new_n15530_));
  AOI21_X1   g14528(.A1(new_n13997_), .A2(new_n14319_), .B(new_n13570_), .ZN(new_n15531_));
  NOR3_X1    g14529(.A1(new_n14316_), .A2(new_n14318_), .A3(new_n13998_), .ZN(new_n15532_));
  NOR2_X1    g14530(.A1(new_n15532_), .A2(new_n15531_), .ZN(new_n15533_));
  NAND3_X1   g14531(.A1(new_n15524_), .A2(new_n15525_), .A3(new_n15529_), .ZN(new_n15534_));
  AOI21_X1   g14532(.A1(new_n15533_), .A2(new_n15534_), .B(new_n15530_), .ZN(new_n15535_));
  OAI21_X1   g14533(.A1(new_n15523_), .A2(new_n15535_), .B(new_n15522_), .ZN(new_n15536_));
  NOR3_X1    g14534(.A1(new_n14329_), .A2(new_n14328_), .A3(new_n14327_), .ZN(new_n15537_));
  AOI21_X1   g14535(.A1(new_n14314_), .A2(new_n14309_), .B(new_n14227_), .ZN(new_n15538_));
  NOR3_X1    g14536(.A1(new_n15515_), .A2(new_n15513_), .A3(new_n15514_), .ZN(new_n15539_));
  AOI21_X1   g14537(.A1(new_n15496_), .A2(new_n15489_), .B(new_n15408_), .ZN(new_n15540_));
  OAI22_X1   g14538(.A1(new_n15537_), .A2(new_n15538_), .B1(new_n15539_), .B2(new_n15540_), .ZN(new_n15541_));
  NAND2_X1   g14539(.A1(new_n15541_), .A2(new_n15536_), .ZN(new_n15542_));
  NAND2_X1   g14540(.A1(new_n15542_), .A2(new_n15517_), .ZN(new_n15543_));
  NAND2_X1   g14541(.A1(new_n14314_), .A2(new_n14227_), .ZN(new_n15544_));
  NAND2_X1   g14542(.A1(new_n14265_), .A2(new_n14258_), .ZN(new_n15545_));
  NAND2_X1   g14543(.A1(new_n15545_), .A2(new_n14263_), .ZN(new_n15546_));
  INV_X1     g14544(.I(new_n14230_), .ZN(new_n15547_));
  NAND2_X1   g14545(.A1(new_n15547_), .A2(new_n14232_), .ZN(new_n15548_));
  OAI22_X1   g14546(.A1(new_n14229_), .A2(new_n14211_), .B1(new_n15547_), .B2(new_n14232_), .ZN(new_n15549_));
  NAND2_X1   g14547(.A1(new_n15549_), .A2(new_n15548_), .ZN(new_n15550_));
  NAND2_X1   g14548(.A1(new_n14243_), .A2(new_n14147_), .ZN(new_n15551_));
  NOR2_X1    g14549(.A1(new_n15551_), .A2(new_n14245_), .ZN(new_n15552_));
  AOI22_X1   g14550(.A1(new_n14253_), .A2(new_n14156_), .B1(new_n15551_), .B2(new_n14245_), .ZN(new_n15553_));
  NOR2_X1    g14551(.A1(new_n15553_), .A2(new_n15552_), .ZN(new_n15554_));
  XOR2_X1    g14552(.A1(new_n15554_), .A2(new_n15550_), .Z(new_n15555_));
  NAND2_X1   g14553(.A1(new_n15546_), .A2(new_n15555_), .ZN(new_n15556_));
  XNOR2_X1   g14554(.A1(new_n15554_), .A2(new_n15550_), .ZN(new_n15557_));
  NAND3_X1   g14555(.A1(new_n15557_), .A2(new_n14263_), .A3(new_n15545_), .ZN(new_n15558_));
  AOI21_X1   g14556(.A1(new_n14305_), .A2(new_n14298_), .B(new_n14307_), .ZN(new_n15559_));
  INV_X1     g14557(.I(new_n15559_), .ZN(new_n15560_));
  NAND2_X1   g14558(.A1(new_n14280_), .A2(new_n14092_), .ZN(new_n15561_));
  NAND2_X1   g14559(.A1(new_n14270_), .A2(new_n14083_), .ZN(new_n15562_));
  NOR2_X1    g14560(.A1(new_n15562_), .A2(new_n14272_), .ZN(new_n15563_));
  NAND2_X1   g14561(.A1(new_n15562_), .A2(new_n14272_), .ZN(new_n15564_));
  AOI21_X1   g14562(.A1(new_n15561_), .A2(new_n15564_), .B(new_n15563_), .ZN(new_n15565_));
  NAND2_X1   g14563(.A1(new_n14292_), .A2(new_n14039_), .ZN(new_n15566_));
  NOR2_X1    g14564(.A1(new_n14294_), .A2(new_n14287_), .ZN(new_n15567_));
  NAND2_X1   g14565(.A1(new_n14294_), .A2(new_n14287_), .ZN(new_n15568_));
  AOI21_X1   g14566(.A1(new_n15566_), .A2(new_n15568_), .B(new_n15567_), .ZN(new_n15569_));
  XNOR2_X1   g14567(.A1(new_n15569_), .A2(new_n15565_), .ZN(new_n15570_));
  NAND2_X1   g14568(.A1(new_n15560_), .A2(new_n15570_), .ZN(new_n15571_));
  XOR2_X1    g14569(.A1(new_n15569_), .A2(new_n15565_), .Z(new_n15572_));
  NAND2_X1   g14570(.A1(new_n15572_), .A2(new_n15559_), .ZN(new_n15573_));
  NAND4_X1   g14571(.A1(new_n15571_), .A2(new_n15556_), .A3(new_n15558_), .A4(new_n15573_), .ZN(new_n15574_));
  INV_X1     g14572(.I(new_n15556_), .ZN(new_n15575_));
  NOR2_X1    g14573(.A1(new_n15546_), .A2(new_n15555_), .ZN(new_n15576_));
  NOR2_X1    g14574(.A1(new_n15572_), .A2(new_n15559_), .ZN(new_n15577_));
  INV_X1     g14575(.I(new_n15573_), .ZN(new_n15578_));
  OAI22_X1   g14576(.A1(new_n15575_), .A2(new_n15576_), .B1(new_n15577_), .B2(new_n15578_), .ZN(new_n15579_));
  NAND4_X1   g14577(.A1(new_n15579_), .A2(new_n14309_), .A3(new_n15574_), .A4(new_n15544_), .ZN(new_n15580_));
  NAND2_X1   g14578(.A1(new_n15544_), .A2(new_n14309_), .ZN(new_n15581_));
  NOR4_X1    g14579(.A1(new_n15575_), .A2(new_n15576_), .A3(new_n15577_), .A4(new_n15578_), .ZN(new_n15582_));
  AOI22_X1   g14580(.A1(new_n15571_), .A2(new_n15573_), .B1(new_n15556_), .B2(new_n15558_), .ZN(new_n15583_));
  OAI21_X1   g14581(.A1(new_n15582_), .A2(new_n15583_), .B(new_n15581_), .ZN(new_n15584_));
  NAND2_X1   g14582(.A1(new_n15584_), .A2(new_n15580_), .ZN(new_n15585_));
  NAND2_X1   g14583(.A1(new_n15543_), .A2(new_n15585_), .ZN(new_n15586_));
  OAI21_X1   g14584(.A1(new_n15515_), .A2(new_n15513_), .B(new_n15489_), .ZN(new_n15587_));
  AOI21_X1   g14585(.A1(new_n15445_), .A2(new_n15438_), .B(new_n15447_), .ZN(new_n15588_));
  NAND2_X1   g14586(.A1(new_n15415_), .A2(new_n15413_), .ZN(new_n15589_));
  OAI21_X1   g14587(.A1(new_n15410_), .A2(new_n15374_), .B(new_n15589_), .ZN(new_n15590_));
  OAI21_X1   g14588(.A1(new_n15415_), .A2(new_n15413_), .B(new_n15590_), .ZN(new_n15591_));
  INV_X1     g14589(.I(new_n15428_), .ZN(new_n15592_));
  OAI22_X1   g14590(.A1(new_n15426_), .A2(new_n15323_), .B1(new_n15592_), .B2(new_n15429_), .ZN(new_n15593_));
  OAI21_X1   g14591(.A1(new_n15428_), .A2(new_n15434_), .B(new_n15593_), .ZN(new_n15594_));
  XOR2_X1    g14592(.A1(new_n15594_), .A2(new_n15591_), .Z(new_n15595_));
  NOR2_X1    g14593(.A1(new_n15595_), .A2(new_n15588_), .ZN(new_n15596_));
  INV_X1     g14594(.I(new_n15588_), .ZN(new_n15597_));
  XNOR2_X1   g14595(.A1(new_n15594_), .A2(new_n15591_), .ZN(new_n15598_));
  NOR2_X1    g14596(.A1(new_n15598_), .A2(new_n15597_), .ZN(new_n15599_));
  AOI21_X1   g14597(.A1(new_n15486_), .A2(new_n15479_), .B(new_n15493_), .ZN(new_n15600_));
  NAND2_X1   g14598(.A1(new_n15451_), .A2(new_n14819_), .ZN(new_n15601_));
  NOR2_X1    g14599(.A1(new_n15601_), .A2(new_n15453_), .ZN(new_n15602_));
  AOI22_X1   g14600(.A1(new_n15459_), .A2(new_n14828_), .B1(new_n15601_), .B2(new_n15453_), .ZN(new_n15603_));
  NOR2_X1    g14601(.A1(new_n15603_), .A2(new_n15602_), .ZN(new_n15604_));
  NAND2_X1   g14602(.A1(new_n15474_), .A2(new_n14567_), .ZN(new_n15605_));
  NAND2_X1   g14603(.A1(new_n15466_), .A2(new_n14560_), .ZN(new_n15606_));
  NOR2_X1    g14604(.A1(new_n15606_), .A2(new_n15468_), .ZN(new_n15607_));
  NAND2_X1   g14605(.A1(new_n15606_), .A2(new_n15468_), .ZN(new_n15608_));
  AOI21_X1   g14606(.A1(new_n15605_), .A2(new_n15608_), .B(new_n15607_), .ZN(new_n15609_));
  XOR2_X1    g14607(.A1(new_n15604_), .A2(new_n15609_), .Z(new_n15610_));
  NOR2_X1    g14608(.A1(new_n15610_), .A2(new_n15600_), .ZN(new_n15611_));
  INV_X1     g14609(.I(new_n15600_), .ZN(new_n15612_));
  XNOR2_X1   g14610(.A1(new_n15604_), .A2(new_n15609_), .ZN(new_n15613_));
  NOR2_X1    g14611(.A1(new_n15612_), .A2(new_n15613_), .ZN(new_n15614_));
  NOR4_X1    g14612(.A1(new_n15599_), .A2(new_n15614_), .A3(new_n15596_), .A4(new_n15611_), .ZN(new_n15615_));
  NAND2_X1   g14613(.A1(new_n15598_), .A2(new_n15597_), .ZN(new_n15616_));
  NAND2_X1   g14614(.A1(new_n15595_), .A2(new_n15588_), .ZN(new_n15617_));
  INV_X1     g14615(.I(new_n15611_), .ZN(new_n15618_));
  NAND2_X1   g14616(.A1(new_n15610_), .A2(new_n15600_), .ZN(new_n15619_));
  AOI22_X1   g14617(.A1(new_n15618_), .A2(new_n15619_), .B1(new_n15616_), .B2(new_n15617_), .ZN(new_n15620_));
  NOR3_X1    g14618(.A1(new_n15620_), .A2(new_n15615_), .A3(new_n15587_), .ZN(new_n15621_));
  AOI21_X1   g14619(.A1(new_n15408_), .A2(new_n15496_), .B(new_n15514_), .ZN(new_n15622_));
  NAND4_X1   g14620(.A1(new_n15618_), .A2(new_n15616_), .A3(new_n15617_), .A4(new_n15619_), .ZN(new_n15623_));
  OAI22_X1   g14621(.A1(new_n15596_), .A2(new_n15599_), .B1(new_n15614_), .B2(new_n15611_), .ZN(new_n15624_));
  AOI21_X1   g14622(.A1(new_n15624_), .A2(new_n15623_), .B(new_n15622_), .ZN(new_n15625_));
  NOR2_X1    g14623(.A1(new_n15625_), .A2(new_n15621_), .ZN(new_n15626_));
  INV_X1     g14624(.I(new_n15626_), .ZN(new_n15627_));
  OAI21_X1   g14625(.A1(new_n15543_), .A2(new_n15585_), .B(new_n15627_), .ZN(new_n15628_));
  NAND2_X1   g14626(.A1(new_n15628_), .A2(new_n15586_), .ZN(new_n15629_));
  NAND2_X1   g14627(.A1(new_n15623_), .A2(new_n15622_), .ZN(new_n15630_));
  NAND2_X1   g14628(.A1(new_n15594_), .A2(new_n15591_), .ZN(new_n15631_));
  INV_X1     g14629(.I(new_n15631_), .ZN(new_n15632_));
  NOR2_X1    g14630(.A1(new_n15594_), .A2(new_n15591_), .ZN(new_n15633_));
  NOR3_X1    g14631(.A1(new_n15632_), .A2(new_n15588_), .A3(new_n15633_), .ZN(new_n15634_));
  NOR2_X1    g14632(.A1(new_n15604_), .A2(new_n15609_), .ZN(new_n15635_));
  NAND2_X1   g14633(.A1(new_n15604_), .A2(new_n15609_), .ZN(new_n15636_));
  INV_X1     g14634(.I(new_n15636_), .ZN(new_n15637_));
  NOR3_X1    g14635(.A1(new_n15600_), .A2(new_n15635_), .A3(new_n15637_), .ZN(new_n15638_));
  NOR2_X1    g14636(.A1(new_n15612_), .A2(new_n15610_), .ZN(new_n15639_));
  NOR2_X1    g14637(.A1(new_n15595_), .A2(new_n15597_), .ZN(new_n15640_));
  NOR4_X1    g14638(.A1(new_n15640_), .A2(new_n15639_), .A3(new_n15634_), .A4(new_n15638_), .ZN(new_n15641_));
  INV_X1     g14639(.I(new_n15641_), .ZN(new_n15642_));
  OAI21_X1   g14640(.A1(new_n15588_), .A2(new_n15633_), .B(new_n15631_), .ZN(new_n15643_));
  INV_X1     g14641(.I(new_n15635_), .ZN(new_n15644_));
  OAI21_X1   g14642(.A1(new_n15600_), .A2(new_n15637_), .B(new_n15644_), .ZN(new_n15645_));
  XNOR2_X1   g14643(.A1(new_n15645_), .A2(new_n15643_), .ZN(new_n15646_));
  INV_X1     g14644(.I(new_n15646_), .ZN(new_n15647_));
  AOI21_X1   g14645(.A1(new_n15642_), .A2(new_n15630_), .B(new_n15647_), .ZN(new_n15648_));
  NOR2_X1    g14646(.A1(new_n15615_), .A2(new_n15587_), .ZN(new_n15649_));
  NOR3_X1    g14647(.A1(new_n15649_), .A2(new_n15646_), .A3(new_n15641_), .ZN(new_n15650_));
  NAND3_X1   g14648(.A1(new_n15574_), .A2(new_n15544_), .A3(new_n14309_), .ZN(new_n15651_));
  INV_X1     g14649(.I(new_n15546_), .ZN(new_n15652_));
  INV_X1     g14650(.I(new_n15554_), .ZN(new_n15653_));
  NAND2_X1   g14651(.A1(new_n15653_), .A2(new_n15550_), .ZN(new_n15654_));
  INV_X1     g14652(.I(new_n15654_), .ZN(new_n15655_));
  NOR2_X1    g14653(.A1(new_n15653_), .A2(new_n15550_), .ZN(new_n15656_));
  NOR3_X1    g14654(.A1(new_n15652_), .A2(new_n15655_), .A3(new_n15656_), .ZN(new_n15657_));
  NOR2_X1    g14655(.A1(new_n15569_), .A2(new_n15565_), .ZN(new_n15658_));
  AND2_X2    g14656(.A1(new_n15569_), .A2(new_n15565_), .Z(new_n15659_));
  NOR3_X1    g14657(.A1(new_n15559_), .A2(new_n15658_), .A3(new_n15659_), .ZN(new_n15660_));
  NOR2_X1    g14658(.A1(new_n15560_), .A2(new_n15572_), .ZN(new_n15661_));
  NOR2_X1    g14659(.A1(new_n15546_), .A2(new_n15557_), .ZN(new_n15662_));
  NOR4_X1    g14660(.A1(new_n15657_), .A2(new_n15660_), .A3(new_n15661_), .A4(new_n15662_), .ZN(new_n15663_));
  INV_X1     g14661(.I(new_n15663_), .ZN(new_n15664_));
  INV_X1     g14662(.I(new_n15656_), .ZN(new_n15665_));
  AOI21_X1   g14663(.A1(new_n15546_), .A2(new_n15665_), .B(new_n15655_), .ZN(new_n15666_));
  INV_X1     g14664(.I(new_n15658_), .ZN(new_n15667_));
  OAI21_X1   g14665(.A1(new_n15559_), .A2(new_n15659_), .B(new_n15667_), .ZN(new_n15668_));
  XNOR2_X1   g14666(.A1(new_n15666_), .A2(new_n15668_), .ZN(new_n15669_));
  AOI21_X1   g14667(.A1(new_n15664_), .A2(new_n15651_), .B(new_n15669_), .ZN(new_n15670_));
  NOR2_X1    g14668(.A1(new_n15581_), .A2(new_n15582_), .ZN(new_n15671_));
  XOR2_X1    g14669(.A1(new_n15666_), .A2(new_n15668_), .Z(new_n15672_));
  NOR3_X1    g14670(.A1(new_n15671_), .A2(new_n15663_), .A3(new_n15672_), .ZN(new_n15673_));
  NOR4_X1    g14671(.A1(new_n15673_), .A2(new_n15648_), .A3(new_n15670_), .A4(new_n15650_), .ZN(new_n15674_));
  OAI21_X1   g14672(.A1(new_n15649_), .A2(new_n15641_), .B(new_n15646_), .ZN(new_n15675_));
  NAND3_X1   g14673(.A1(new_n15647_), .A2(new_n15630_), .A3(new_n15642_), .ZN(new_n15676_));
  OAI21_X1   g14674(.A1(new_n15671_), .A2(new_n15663_), .B(new_n15672_), .ZN(new_n15677_));
  NAND3_X1   g14675(.A1(new_n15664_), .A2(new_n15669_), .A3(new_n15651_), .ZN(new_n15678_));
  AOI22_X1   g14676(.A1(new_n15677_), .A2(new_n15678_), .B1(new_n15675_), .B2(new_n15676_), .ZN(new_n15679_));
  NOR2_X1    g14677(.A1(new_n15674_), .A2(new_n15679_), .ZN(new_n15680_));
  NAND2_X1   g14678(.A1(new_n15629_), .A2(new_n15680_), .ZN(new_n15681_));
  NAND4_X1   g14679(.A1(new_n15677_), .A2(new_n15678_), .A3(new_n15676_), .A4(new_n15675_), .ZN(new_n15682_));
  OAI22_X1   g14680(.A1(new_n15673_), .A2(new_n15670_), .B1(new_n15648_), .B2(new_n15650_), .ZN(new_n15683_));
  NAND2_X1   g14681(.A1(new_n15683_), .A2(new_n15682_), .ZN(new_n15684_));
  NAND3_X1   g14682(.A1(new_n15684_), .A2(new_n15586_), .A3(new_n15628_), .ZN(new_n15685_));
  NAND4_X1   g14683(.A1(new_n13159_), .A2(new_n13124_), .A3(new_n15681_), .A4(new_n15685_), .ZN(new_n15686_));
  NOR3_X1    g14684(.A1(new_n12947_), .A2(new_n13146_), .A3(new_n13127_), .ZN(new_n15687_));
  AOI21_X1   g14685(.A1(new_n12948_), .A2(new_n13145_), .B(new_n11766_), .ZN(new_n15688_));
  NOR2_X1    g14686(.A1(new_n15688_), .A2(new_n15687_), .ZN(new_n15689_));
  NOR3_X1    g14687(.A1(new_n15502_), .A2(new_n15393_), .A3(new_n15407_), .ZN(new_n15690_));
  AOI21_X1   g14688(.A1(new_n15503_), .A2(new_n15392_), .B(new_n15512_), .ZN(new_n15691_));
  NOR3_X1    g14689(.A1(new_n14325_), .A2(new_n14226_), .A3(new_n13999_), .ZN(new_n15692_));
  AOI21_X1   g14690(.A1(new_n14326_), .A2(new_n14225_), .B(new_n14320_), .ZN(new_n15693_));
  OAI22_X1   g14691(.A1(new_n15692_), .A2(new_n15693_), .B1(new_n15690_), .B2(new_n15691_), .ZN(new_n15694_));
  NOR3_X1    g14692(.A1(new_n15402_), .A2(new_n15511_), .A3(new_n15405_), .ZN(new_n15695_));
  AOI21_X1   g14693(.A1(new_n15406_), .A2(new_n15507_), .B(new_n15510_), .ZN(new_n15696_));
  INV_X1     g14694(.I(new_n15529_), .ZN(new_n15697_));
  OAI21_X1   g14695(.A1(new_n15696_), .A2(new_n15695_), .B(new_n15697_), .ZN(new_n15698_));
  NAND2_X1   g14696(.A1(new_n13997_), .A2(new_n13570_), .ZN(new_n15699_));
  NOR2_X1    g14697(.A1(new_n14318_), .A2(new_n13998_), .ZN(new_n15700_));
  OAI22_X1   g14698(.A1(new_n15700_), .A2(new_n13570_), .B1(new_n15699_), .B2(new_n13998_), .ZN(new_n15701_));
  NOR3_X1    g14699(.A1(new_n15696_), .A2(new_n15695_), .A3(new_n15697_), .ZN(new_n15702_));
  OAI21_X1   g14700(.A1(new_n15701_), .A2(new_n15702_), .B(new_n15698_), .ZN(new_n15703_));
  NAND3_X1   g14701(.A1(new_n15694_), .A2(new_n15522_), .A3(new_n15703_), .ZN(new_n15704_));
  NOR4_X1    g14702(.A1(new_n15690_), .A2(new_n15692_), .A3(new_n15693_), .A4(new_n15691_), .ZN(new_n15705_));
  OAI21_X1   g14703(.A1(new_n15705_), .A2(new_n15523_), .B(new_n15535_), .ZN(new_n15706_));
  NAND3_X1   g14704(.A1(new_n12945_), .A2(new_n13142_), .A3(new_n12939_), .ZN(new_n15707_));
  OAI21_X1   g14705(.A1(new_n12944_), .A2(new_n13143_), .B(new_n13137_), .ZN(new_n15708_));
  NAND4_X1   g14706(.A1(new_n15706_), .A2(new_n15708_), .A3(new_n15704_), .A4(new_n15707_), .ZN(new_n15709_));
  NAND3_X1   g14707(.A1(new_n15541_), .A2(new_n15517_), .A3(new_n15536_), .ZN(new_n15710_));
  AOI21_X1   g14708(.A1(new_n15694_), .A2(new_n15703_), .B(new_n15705_), .ZN(new_n15711_));
  NOR4_X1    g14709(.A1(new_n15537_), .A2(new_n15538_), .A3(new_n15539_), .A4(new_n15540_), .ZN(new_n15712_));
  AOI22_X1   g14710(.A1(new_n14315_), .A2(new_n14330_), .B1(new_n15516_), .B2(new_n15497_), .ZN(new_n15713_));
  OAI21_X1   g14711(.A1(new_n15712_), .A2(new_n15713_), .B(new_n15711_), .ZN(new_n15714_));
  NAND2_X1   g14712(.A1(new_n15714_), .A2(new_n15710_), .ZN(new_n15715_));
  NOR3_X1    g14713(.A1(new_n15705_), .A2(new_n15523_), .A3(new_n15535_), .ZN(new_n15716_));
  AOI21_X1   g14714(.A1(new_n15694_), .A2(new_n15522_), .B(new_n15703_), .ZN(new_n15717_));
  NOR2_X1    g14715(.A1(new_n15716_), .A2(new_n15717_), .ZN(new_n15718_));
  NOR3_X1    g14716(.A1(new_n12944_), .A2(new_n13143_), .A3(new_n13137_), .ZN(new_n15719_));
  AOI21_X1   g14717(.A1(new_n12945_), .A2(new_n13142_), .B(new_n12939_), .ZN(new_n15720_));
  NOR2_X1    g14718(.A1(new_n15719_), .A2(new_n15720_), .ZN(new_n15721_));
  NOR2_X1    g14719(.A1(new_n12933_), .A2(new_n12931_), .ZN(new_n15722_));
  NOR2_X1    g14720(.A1(new_n13132_), .A2(new_n15722_), .ZN(new_n15723_));
  NOR2_X1    g14721(.A1(new_n13876_), .A2(new_n15528_), .ZN(new_n15724_));
  AOI21_X1   g14722(.A1(new_n15506_), .A2(new_n15526_), .B(new_n15724_), .ZN(new_n15725_));
  NOR2_X1    g14723(.A1(new_n15725_), .A2(new_n15529_), .ZN(new_n15726_));
  NAND2_X1   g14724(.A1(new_n15723_), .A2(new_n15726_), .ZN(new_n15727_));
  NOR3_X1    g14725(.A1(new_n15533_), .A2(new_n15702_), .A3(new_n15530_), .ZN(new_n15728_));
  AOI21_X1   g14726(.A1(new_n15534_), .A2(new_n15698_), .B(new_n15701_), .ZN(new_n15729_));
  OAI21_X1   g14727(.A1(new_n15729_), .A2(new_n15728_), .B(new_n15727_), .ZN(new_n15730_));
  OAI21_X1   g14728(.A1(new_n13136_), .A2(new_n12937_), .B(new_n12929_), .ZN(new_n15731_));
  NAND3_X1   g14729(.A1(new_n13135_), .A2(new_n12938_), .A3(new_n13131_), .ZN(new_n15732_));
  NAND2_X1   g14730(.A1(new_n15731_), .A2(new_n15732_), .ZN(new_n15733_));
  NOR3_X1    g14731(.A1(new_n15729_), .A2(new_n15728_), .A3(new_n15727_), .ZN(new_n15734_));
  OAI21_X1   g14732(.A1(new_n15733_), .A2(new_n15734_), .B(new_n15730_), .ZN(new_n15735_));
  OAI21_X1   g14733(.A1(new_n15718_), .A2(new_n15721_), .B(new_n15735_), .ZN(new_n15736_));
  AOI21_X1   g14734(.A1(new_n15709_), .A2(new_n15736_), .B(new_n15715_), .ZN(new_n15737_));
  NAND3_X1   g14735(.A1(new_n15715_), .A2(new_n15736_), .A3(new_n15709_), .ZN(new_n15738_));
  AOI21_X1   g14736(.A1(new_n15689_), .A2(new_n15738_), .B(new_n15737_), .ZN(new_n15739_));
  AOI21_X1   g14737(.A1(new_n15517_), .A2(new_n15542_), .B(new_n15585_), .ZN(new_n15740_));
  NOR3_X1    g14738(.A1(new_n15581_), .A2(new_n15582_), .A3(new_n15583_), .ZN(new_n15741_));
  AOI22_X1   g14739(.A1(new_n15579_), .A2(new_n15574_), .B1(new_n14309_), .B2(new_n15544_), .ZN(new_n15742_));
  NOR2_X1    g14740(.A1(new_n15742_), .A2(new_n15741_), .ZN(new_n15743_));
  NOR2_X1    g14741(.A1(new_n15543_), .A2(new_n15743_), .ZN(new_n15744_));
  OAI21_X1   g14742(.A1(new_n15744_), .A2(new_n15740_), .B(new_n15627_), .ZN(new_n15745_));
  NAND2_X1   g14743(.A1(new_n15543_), .A2(new_n15743_), .ZN(new_n15746_));
  NAND3_X1   g14744(.A1(new_n15585_), .A2(new_n15517_), .A3(new_n15542_), .ZN(new_n15747_));
  NAND3_X1   g14745(.A1(new_n15746_), .A2(new_n15747_), .A3(new_n15626_), .ZN(new_n15748_));
  OAI21_X1   g14746(.A1(new_n13081_), .A2(new_n13153_), .B(new_n12949_), .ZN(new_n15749_));
  NAND3_X1   g14747(.A1(new_n13154_), .A2(new_n13080_), .A3(new_n13147_), .ZN(new_n15750_));
  NAND4_X1   g14748(.A1(new_n15745_), .A2(new_n15748_), .A3(new_n15749_), .A4(new_n15750_), .ZN(new_n15751_));
  AOI22_X1   g14749(.A1(new_n15745_), .A2(new_n15748_), .B1(new_n15749_), .B2(new_n15750_), .ZN(new_n15752_));
  OAI21_X1   g14750(.A1(new_n15739_), .A2(new_n15752_), .B(new_n15751_), .ZN(new_n15753_));
  NOR2_X1    g14751(.A1(new_n13155_), .A2(new_n13158_), .ZN(new_n15754_));
  NOR2_X1    g14752(.A1(new_n13123_), .A2(new_n13082_), .ZN(new_n15755_));
  AOI21_X1   g14753(.A1(new_n15586_), .A2(new_n15628_), .B(new_n15684_), .ZN(new_n15756_));
  NOR2_X1    g14754(.A1(new_n15629_), .A2(new_n15680_), .ZN(new_n15757_));
  OAI22_X1   g14755(.A1(new_n15754_), .A2(new_n15755_), .B1(new_n15756_), .B2(new_n15757_), .ZN(new_n15758_));
  NAND2_X1   g14756(.A1(new_n15753_), .A2(new_n15758_), .ZN(new_n15759_));
  NOR2_X1    g14757(.A1(new_n13097_), .A2(new_n13091_), .ZN(new_n15760_));
  NOR2_X1    g14758(.A1(new_n13094_), .A2(new_n13093_), .ZN(new_n15761_));
  AND2_X2    g14759(.A1(new_n13094_), .A2(new_n13093_), .Z(new_n15762_));
  NOR3_X1    g14760(.A1(new_n15760_), .A2(new_n15761_), .A3(new_n15762_), .ZN(new_n15763_));
  NOR2_X1    g14761(.A1(new_n13114_), .A2(new_n13107_), .ZN(new_n15764_));
  NOR2_X1    g14762(.A1(new_n13110_), .A2(new_n13109_), .ZN(new_n15765_));
  AND2_X2    g14763(.A1(new_n13110_), .A2(new_n13109_), .Z(new_n15766_));
  NOR3_X1    g14764(.A1(new_n15764_), .A2(new_n15765_), .A3(new_n15766_), .ZN(new_n15767_));
  NOR3_X1    g14765(.A1(new_n13114_), .A2(new_n13107_), .A3(new_n13111_), .ZN(new_n15768_));
  NOR3_X1    g14766(.A1(new_n13097_), .A2(new_n13095_), .A3(new_n13091_), .ZN(new_n15769_));
  NOR4_X1    g14767(.A1(new_n15767_), .A2(new_n15763_), .A3(new_n15768_), .A4(new_n15769_), .ZN(new_n15770_));
  AOI21_X1   g14768(.A1(new_n13155_), .A2(new_n13156_), .B(new_n15770_), .ZN(new_n15771_));
  INV_X1     g14769(.I(new_n15771_), .ZN(new_n15772_));
  INV_X1     g14770(.I(new_n15765_), .ZN(new_n15773_));
  OAI21_X1   g14771(.A1(new_n15764_), .A2(new_n15766_), .B(new_n15773_), .ZN(new_n15774_));
  NOR2_X1    g14772(.A1(new_n15760_), .A2(new_n15762_), .ZN(new_n15775_));
  NOR2_X1    g14773(.A1(new_n15775_), .A2(new_n15761_), .ZN(new_n15776_));
  XOR2_X1    g14774(.A1(new_n15776_), .A2(new_n15774_), .Z(new_n15777_));
  NAND2_X1   g14775(.A1(new_n15772_), .A2(new_n15777_), .ZN(new_n15778_));
  INV_X1     g14776(.I(new_n15777_), .ZN(new_n15779_));
  NAND2_X1   g14777(.A1(new_n15779_), .A2(new_n15771_), .ZN(new_n15780_));
  NAND3_X1   g14778(.A1(new_n15628_), .A2(new_n15586_), .A3(new_n15682_), .ZN(new_n15781_));
  NOR2_X1    g14779(.A1(new_n15649_), .A2(new_n15641_), .ZN(new_n15782_));
  NAND2_X1   g14780(.A1(new_n15645_), .A2(new_n15643_), .ZN(new_n15783_));
  INV_X1     g14781(.I(new_n15783_), .ZN(new_n15784_));
  NOR2_X1    g14782(.A1(new_n15645_), .A2(new_n15643_), .ZN(new_n15785_));
  OR3_X2     g14783(.A1(new_n15782_), .A2(new_n15784_), .A3(new_n15785_), .Z(new_n15786_));
  NOR2_X1    g14784(.A1(new_n15671_), .A2(new_n15663_), .ZN(new_n15787_));
  INV_X1     g14785(.I(new_n15666_), .ZN(new_n15788_));
  NAND2_X1   g14786(.A1(new_n15788_), .A2(new_n15668_), .ZN(new_n15789_));
  INV_X1     g14787(.I(new_n15789_), .ZN(new_n15790_));
  NOR2_X1    g14788(.A1(new_n15788_), .A2(new_n15668_), .ZN(new_n15791_));
  OR3_X2     g14789(.A1(new_n15787_), .A2(new_n15790_), .A3(new_n15791_), .Z(new_n15792_));
  NAND2_X1   g14790(.A1(new_n15787_), .A2(new_n15672_), .ZN(new_n15793_));
  NAND2_X1   g14791(.A1(new_n15782_), .A2(new_n15646_), .ZN(new_n15794_));
  NAND4_X1   g14792(.A1(new_n15792_), .A2(new_n15786_), .A3(new_n15793_), .A4(new_n15794_), .ZN(new_n15795_));
  OAI21_X1   g14793(.A1(new_n15787_), .A2(new_n15791_), .B(new_n15789_), .ZN(new_n15796_));
  OAI21_X1   g14794(.A1(new_n15782_), .A2(new_n15785_), .B(new_n15783_), .ZN(new_n15797_));
  XOR2_X1    g14795(.A1(new_n15796_), .A2(new_n15797_), .Z(new_n15798_));
  AOI21_X1   g14796(.A1(new_n15781_), .A2(new_n15795_), .B(new_n15798_), .ZN(new_n15799_));
  INV_X1     g14797(.I(new_n15799_), .ZN(new_n15800_));
  NAND3_X1   g14798(.A1(new_n15798_), .A2(new_n15795_), .A3(new_n15781_), .ZN(new_n15801_));
  NAND4_X1   g14799(.A1(new_n15778_), .A2(new_n15780_), .A3(new_n15800_), .A4(new_n15801_), .ZN(new_n15802_));
  NAND3_X1   g14800(.A1(new_n15802_), .A2(new_n15759_), .A3(new_n15686_), .ZN(new_n15803_));
  OAI21_X1   g14801(.A1(new_n15761_), .A2(new_n15775_), .B(new_n15774_), .ZN(new_n15804_));
  NOR3_X1    g14802(.A1(new_n15774_), .A2(new_n15761_), .A3(new_n15775_), .ZN(new_n15805_));
  INV_X1     g14803(.I(new_n15805_), .ZN(new_n15806_));
  NAND3_X1   g14804(.A1(new_n15772_), .A2(new_n15804_), .A3(new_n15806_), .ZN(new_n15807_));
  AND2_X2    g14805(.A1(new_n15796_), .A2(new_n15797_), .Z(new_n15808_));
  NAND2_X1   g14806(.A1(new_n15781_), .A2(new_n15795_), .ZN(new_n15809_));
  OR2_X2     g14807(.A1(new_n15796_), .A2(new_n15797_), .Z(new_n15810_));
  NAND2_X1   g14808(.A1(new_n15809_), .A2(new_n15810_), .ZN(new_n15811_));
  NOR2_X1    g14809(.A1(new_n15811_), .A2(new_n15808_), .ZN(new_n15812_));
  NOR2_X1    g14810(.A1(new_n15809_), .A2(new_n15798_), .ZN(new_n15813_));
  NOR2_X1    g14811(.A1(new_n15812_), .A2(new_n15813_), .ZN(new_n15814_));
  NOR2_X1    g14812(.A1(new_n15772_), .A2(new_n15779_), .ZN(new_n15815_));
  INV_X1     g14813(.I(new_n15815_), .ZN(new_n15816_));
  NAND3_X1   g14814(.A1(new_n15814_), .A2(new_n15807_), .A3(new_n15816_), .ZN(new_n15817_));
  NAND2_X1   g14815(.A1(new_n15803_), .A2(new_n15817_), .ZN(new_n15818_));
  OAI21_X1   g14816(.A1(new_n15771_), .A2(new_n15805_), .B(new_n15804_), .ZN(new_n15819_));
  AOI21_X1   g14817(.A1(new_n15809_), .A2(new_n15810_), .B(new_n15808_), .ZN(new_n15820_));
  INV_X1     g14818(.I(new_n15820_), .ZN(new_n15821_));
  NAND2_X1   g14819(.A1(new_n15821_), .A2(new_n15819_), .ZN(new_n15822_));
  INV_X1     g14820(.I(new_n15822_), .ZN(new_n15823_));
  NOR2_X1    g14821(.A1(new_n15821_), .A2(new_n15819_), .ZN(new_n15824_));
  INV_X1     g14822(.I(new_n15824_), .ZN(new_n15825_));
  AOI21_X1   g14823(.A1(new_n15818_), .A2(new_n15825_), .B(new_n15823_), .ZN(new_n15826_));
  NAND2_X1   g14824(.A1(new_n10543_), .A2(new_n10544_), .ZN(new_n15827_));
  OAI21_X1   g14825(.A1(new_n10530_), .A2(new_n10539_), .B(new_n15827_), .ZN(new_n15828_));
  NAND3_X1   g14826(.A1(new_n6842_), .A2(new_n6841_), .A3(new_n6840_), .ZN(new_n15829_));
  OAI21_X1   g14827(.A1(new_n6820_), .A2(new_n6825_), .B(new_n6525_), .ZN(new_n15830_));
  NAND2_X1   g14828(.A1(new_n15830_), .A2(new_n15829_), .ZN(new_n15831_));
  AOI21_X1   g14829(.A1(new_n10165_), .A2(new_n10160_), .B(new_n10159_), .ZN(new_n15832_));
  NOR3_X1    g14830(.A1(new_n10139_), .A2(new_n8760_), .A3(new_n10155_), .ZN(new_n15833_));
  NOR2_X1    g14831(.A1(new_n15833_), .A2(new_n15832_), .ZN(new_n15834_));
  NOR2_X1    g14832(.A1(new_n15834_), .A2(new_n15831_), .ZN(new_n15835_));
  NOR3_X1    g14833(.A1(new_n6831_), .A2(new_n6125_), .A3(new_n5194_), .ZN(new_n15836_));
  AOI21_X1   g14834(.A1(new_n6832_), .A2(new_n6124_), .B(new_n5193_), .ZN(new_n15837_));
  NOR2_X1    g14835(.A1(new_n15836_), .A2(new_n15837_), .ZN(new_n15838_));
  NAND2_X1   g14836(.A1(new_n10177_), .A2(new_n10180_), .ZN(new_n15839_));
  NAND2_X1   g14837(.A1(new_n10172_), .A2(new_n10175_), .ZN(new_n15840_));
  NAND2_X1   g14838(.A1(new_n15840_), .A2(new_n15839_), .ZN(new_n15841_));
  NAND2_X1   g14839(.A1(new_n15838_), .A2(new_n15841_), .ZN(new_n15842_));
  INV_X1     g14840(.I(new_n10192_), .ZN(new_n15843_));
  OAI21_X1   g14841(.A1(new_n10201_), .A2(new_n5191_), .B(new_n3089_), .ZN(new_n15844_));
  NAND3_X1   g14842(.A1(new_n10199_), .A2(new_n5192_), .A3(new_n10195_), .ZN(new_n15845_));
  AOI21_X1   g14843(.A1(new_n15844_), .A2(new_n15845_), .B(new_n15843_), .ZN(new_n15846_));
  NAND3_X1   g14844(.A1(new_n15844_), .A2(new_n15845_), .A3(new_n15843_), .ZN(new_n15847_));
  OAI21_X1   g14845(.A1(new_n10186_), .A2(new_n15846_), .B(new_n15847_), .ZN(new_n15848_));
  OAI21_X1   g14846(.A1(new_n15838_), .A2(new_n15841_), .B(new_n15848_), .ZN(new_n15849_));
  NAND2_X1   g14847(.A1(new_n15849_), .A2(new_n15842_), .ZN(new_n15850_));
  NOR3_X1    g14848(.A1(new_n6523_), .A2(new_n6839_), .A3(new_n6833_), .ZN(new_n15851_));
  AOI21_X1   g14849(.A1(new_n6524_), .A2(new_n6838_), .B(new_n6126_), .ZN(new_n15852_));
  AOI21_X1   g14850(.A1(new_n10223_), .A2(new_n10222_), .B(new_n10221_), .ZN(new_n15853_));
  NOR3_X1    g14851(.A1(new_n10214_), .A2(new_n10216_), .A3(new_n10212_), .ZN(new_n15854_));
  NOR4_X1    g14852(.A1(new_n15851_), .A2(new_n15852_), .A3(new_n15854_), .A4(new_n15853_), .ZN(new_n15855_));
  OAI22_X1   g14853(.A1(new_n15851_), .A2(new_n15852_), .B1(new_n15854_), .B2(new_n15853_), .ZN(new_n15856_));
  AOI21_X1   g14854(.A1(new_n15850_), .A2(new_n15856_), .B(new_n15855_), .ZN(new_n15857_));
  AOI21_X1   g14855(.A1(new_n15834_), .A2(new_n15831_), .B(new_n15857_), .ZN(new_n15858_));
  NOR2_X1    g14856(.A1(new_n15858_), .A2(new_n15835_), .ZN(new_n15859_));
  NAND3_X1   g14857(.A1(new_n10324_), .A2(new_n10326_), .A3(new_n10325_), .ZN(new_n15860_));
  OAI21_X1   g14858(.A1(new_n10322_), .A2(new_n10317_), .B(new_n10230_), .ZN(new_n15861_));
  NAND2_X1   g14859(.A1(new_n10410_), .A2(new_n10407_), .ZN(new_n15862_));
  NAND2_X1   g14860(.A1(new_n10402_), .A2(new_n10332_), .ZN(new_n15863_));
  AOI22_X1   g14861(.A1(new_n15862_), .A2(new_n15863_), .B1(new_n15861_), .B2(new_n15860_), .ZN(new_n15864_));
  NAND4_X1   g14862(.A1(new_n15862_), .A2(new_n15863_), .A3(new_n15861_), .A4(new_n15860_), .ZN(new_n15865_));
  AOI21_X1   g14863(.A1(new_n15859_), .A2(new_n15865_), .B(new_n15864_), .ZN(new_n15866_));
  INV_X1     g14864(.I(new_n10465_), .ZN(new_n15867_));
  NOR2_X1    g14865(.A1(new_n15867_), .A2(new_n10466_), .ZN(new_n15868_));
  NAND2_X1   g14866(.A1(new_n15866_), .A2(new_n15868_), .ZN(new_n15869_));
  NAND2_X1   g14867(.A1(new_n10486_), .A2(new_n10487_), .ZN(new_n15870_));
  NAND2_X1   g14868(.A1(new_n10471_), .A2(new_n10483_), .ZN(new_n15871_));
  NAND2_X1   g14869(.A1(new_n15871_), .A2(new_n15870_), .ZN(new_n15872_));
  OAI21_X1   g14870(.A1(new_n15866_), .A2(new_n15868_), .B(new_n15872_), .ZN(new_n15873_));
  NAND2_X1   g14871(.A1(new_n10528_), .A2(new_n10508_), .ZN(new_n15874_));
  NAND2_X1   g14872(.A1(new_n15874_), .A2(new_n10538_), .ZN(new_n15875_));
  NAND3_X1   g14873(.A1(new_n15873_), .A2(new_n15869_), .A3(new_n15875_), .ZN(new_n15876_));
  INV_X1     g14874(.I(new_n10539_), .ZN(new_n15877_));
  NOR2_X1    g14875(.A1(new_n10545_), .A2(new_n10542_), .ZN(new_n15878_));
  NAND3_X1   g14876(.A1(new_n15876_), .A2(new_n15877_), .A3(new_n15878_), .ZN(new_n15879_));
  AOI21_X1   g14877(.A1(new_n15828_), .A2(new_n15879_), .B(new_n15826_), .ZN(new_n15880_));
  INV_X1     g14878(.I(new_n15880_), .ZN(new_n15881_));
  INV_X1     g14879(.I(new_n15709_), .ZN(new_n15882_));
  AOI22_X1   g14880(.A1(new_n15706_), .A2(new_n15704_), .B1(new_n15708_), .B2(new_n15707_), .ZN(new_n15883_));
  INV_X1     g14881(.I(new_n15727_), .ZN(new_n15884_));
  NAND3_X1   g14882(.A1(new_n15701_), .A2(new_n15698_), .A3(new_n15534_), .ZN(new_n15885_));
  INV_X1     g14883(.I(new_n15729_), .ZN(new_n15886_));
  AOI21_X1   g14884(.A1(new_n15886_), .A2(new_n15885_), .B(new_n15884_), .ZN(new_n15887_));
  NOR2_X1    g14885(.A1(new_n15733_), .A2(new_n15734_), .ZN(new_n15888_));
  NOR2_X1    g14886(.A1(new_n15888_), .A2(new_n15887_), .ZN(new_n15889_));
  NOR3_X1    g14887(.A1(new_n15882_), .A2(new_n15883_), .A3(new_n15889_), .ZN(new_n15890_));
  OAI22_X1   g14888(.A1(new_n15716_), .A2(new_n15717_), .B1(new_n15719_), .B2(new_n15720_), .ZN(new_n15891_));
  AOI21_X1   g14889(.A1(new_n15891_), .A2(new_n15709_), .B(new_n15735_), .ZN(new_n15892_));
  NOR2_X1    g14890(.A1(new_n15890_), .A2(new_n15892_), .ZN(new_n15893_));
  NAND2_X1   g14891(.A1(new_n10182_), .A2(new_n10205_), .ZN(new_n15894_));
  NAND2_X1   g14892(.A1(new_n15841_), .A2(new_n15848_), .ZN(new_n15895_));
  AOI21_X1   g14893(.A1(new_n15894_), .A2(new_n15895_), .B(new_n10171_), .ZN(new_n15896_));
  NOR3_X1    g14894(.A1(new_n15848_), .A2(new_n10176_), .A3(new_n10181_), .ZN(new_n15897_));
  NOR2_X1    g14895(.A1(new_n10182_), .A2(new_n10205_), .ZN(new_n15898_));
  NOR3_X1    g14896(.A1(new_n15898_), .A2(new_n15897_), .A3(new_n15838_), .ZN(new_n15899_));
  NOR3_X1    g14897(.A1(new_n15896_), .A2(new_n15899_), .A3(new_n15893_), .ZN(new_n15900_));
  NOR2_X1    g14898(.A1(new_n15887_), .A2(new_n15734_), .ZN(new_n15901_));
  XNOR2_X1   g14899(.A1(new_n15901_), .A2(new_n15733_), .ZN(new_n15902_));
  NOR2_X1    g14900(.A1(new_n15723_), .A2(new_n15726_), .ZN(new_n15903_));
  NOR2_X1    g14901(.A1(new_n15884_), .A2(new_n15903_), .ZN(new_n15904_));
  NOR2_X1    g14902(.A1(new_n10191_), .A2(new_n9973_), .ZN(new_n15905_));
  XNOR2_X1   g14903(.A1(new_n10190_), .A2(new_n15905_), .ZN(new_n15906_));
  AND2_X2    g14904(.A1(new_n15906_), .A2(new_n15904_), .Z(new_n15907_));
  AOI21_X1   g14905(.A1(new_n10203_), .A2(new_n15847_), .B(new_n10187_), .ZN(new_n15908_));
  NOR3_X1    g14906(.A1(new_n15846_), .A2(new_n10204_), .A3(new_n10186_), .ZN(new_n15909_));
  OAI21_X1   g14907(.A1(new_n15908_), .A2(new_n15909_), .B(new_n15907_), .ZN(new_n15910_));
  NAND2_X1   g14908(.A1(new_n15910_), .A2(new_n15902_), .ZN(new_n15911_));
  NOR3_X1    g14909(.A1(new_n15908_), .A2(new_n15909_), .A3(new_n15907_), .ZN(new_n15912_));
  INV_X1     g14910(.I(new_n15912_), .ZN(new_n15913_));
  NAND2_X1   g14911(.A1(new_n15911_), .A2(new_n15913_), .ZN(new_n15914_));
  INV_X1     g14912(.I(new_n15914_), .ZN(new_n15915_));
  OAI21_X1   g14913(.A1(new_n15896_), .A2(new_n15899_), .B(new_n15893_), .ZN(new_n15916_));
  AOI21_X1   g14914(.A1(new_n15915_), .A2(new_n15916_), .B(new_n15900_), .ZN(new_n15917_));
  NAND3_X1   g14915(.A1(new_n10207_), .A2(new_n15856_), .A3(new_n10225_), .ZN(new_n15918_));
  OAI22_X1   g14916(.A1(new_n15855_), .A2(new_n10226_), .B1(new_n10183_), .B2(new_n10206_), .ZN(new_n15919_));
  NOR3_X1    g14917(.A1(new_n15712_), .A2(new_n15713_), .A3(new_n15711_), .ZN(new_n15920_));
  AOI21_X1   g14918(.A1(new_n15541_), .A2(new_n15517_), .B(new_n15536_), .ZN(new_n15921_));
  NOR2_X1    g14919(.A1(new_n15920_), .A2(new_n15921_), .ZN(new_n15922_));
  OAI21_X1   g14920(.A1(new_n15883_), .A2(new_n15889_), .B(new_n15709_), .ZN(new_n15923_));
  NAND2_X1   g14921(.A1(new_n15923_), .A2(new_n15922_), .ZN(new_n15924_));
  NAND3_X1   g14922(.A1(new_n15924_), .A2(new_n15738_), .A3(new_n15689_), .ZN(new_n15925_));
  NAND3_X1   g14923(.A1(new_n12948_), .A2(new_n13145_), .A3(new_n11766_), .ZN(new_n15926_));
  OAI21_X1   g14924(.A1(new_n12947_), .A2(new_n13146_), .B(new_n13127_), .ZN(new_n15927_));
  NAND2_X1   g14925(.A1(new_n15927_), .A2(new_n15926_), .ZN(new_n15928_));
  NOR2_X1    g14926(.A1(new_n15923_), .A2(new_n15922_), .ZN(new_n15929_));
  OAI21_X1   g14927(.A1(new_n15737_), .A2(new_n15929_), .B(new_n15928_), .ZN(new_n15930_));
  NAND2_X1   g14928(.A1(new_n15930_), .A2(new_n15925_), .ZN(new_n15931_));
  AOI21_X1   g14929(.A1(new_n15919_), .A2(new_n15918_), .B(new_n15931_), .ZN(new_n15932_));
  NAND3_X1   g14930(.A1(new_n15919_), .A2(new_n15918_), .A3(new_n15931_), .ZN(new_n15933_));
  OAI21_X1   g14931(.A1(new_n15917_), .A2(new_n15932_), .B(new_n15933_), .ZN(new_n15934_));
  INV_X1     g14932(.I(new_n15739_), .ZN(new_n15935_));
  AOI21_X1   g14933(.A1(new_n15746_), .A2(new_n15747_), .B(new_n15626_), .ZN(new_n15936_));
  NOR3_X1    g14934(.A1(new_n15744_), .A2(new_n15740_), .A3(new_n15627_), .ZN(new_n15937_));
  AOI21_X1   g14935(.A1(new_n13154_), .A2(new_n13080_), .B(new_n13147_), .ZN(new_n15938_));
  NOR3_X1    g14936(.A1(new_n13081_), .A2(new_n13153_), .A3(new_n12949_), .ZN(new_n15939_));
  OAI22_X1   g14937(.A1(new_n15936_), .A2(new_n15937_), .B1(new_n15939_), .B2(new_n15938_), .ZN(new_n15940_));
  NAND3_X1   g14938(.A1(new_n15935_), .A2(new_n15940_), .A3(new_n15751_), .ZN(new_n15941_));
  NOR4_X1    g14939(.A1(new_n15936_), .A2(new_n15937_), .A3(new_n15939_), .A4(new_n15938_), .ZN(new_n15942_));
  OAI21_X1   g14940(.A1(new_n15942_), .A2(new_n15752_), .B(new_n15739_), .ZN(new_n15943_));
  NAND2_X1   g14941(.A1(new_n15941_), .A2(new_n15943_), .ZN(new_n15944_));
  NOR3_X1    g14942(.A1(new_n6844_), .A2(new_n15832_), .A3(new_n15833_), .ZN(new_n15945_));
  OAI21_X1   g14943(.A1(new_n15835_), .A2(new_n15945_), .B(new_n10227_), .ZN(new_n15946_));
  NAND3_X1   g14944(.A1(new_n15831_), .A2(new_n10156_), .A3(new_n10166_), .ZN(new_n15947_));
  NAND3_X1   g14945(.A1(new_n10168_), .A2(new_n15947_), .A3(new_n15857_), .ZN(new_n15948_));
  AOI22_X1   g14946(.A1(new_n15934_), .A2(new_n15944_), .B1(new_n15946_), .B2(new_n15948_), .ZN(new_n15949_));
  NOR2_X1    g14947(.A1(new_n15934_), .A2(new_n15944_), .ZN(new_n15950_));
  AOI21_X1   g14948(.A1(new_n15935_), .A2(new_n15940_), .B(new_n15942_), .ZN(new_n15951_));
  INV_X1     g14949(.I(new_n15686_), .ZN(new_n15952_));
  AOI22_X1   g14950(.A1(new_n13159_), .A2(new_n13124_), .B1(new_n15681_), .B2(new_n15685_), .ZN(new_n15953_));
  NOR3_X1    g14951(.A1(new_n15952_), .A2(new_n15951_), .A3(new_n15953_), .ZN(new_n15954_));
  AOI21_X1   g14952(.A1(new_n15686_), .A2(new_n15758_), .B(new_n15753_), .ZN(new_n15955_));
  NOR2_X1    g14953(.A1(new_n15954_), .A2(new_n15955_), .ZN(new_n15956_));
  OAI21_X1   g14954(.A1(new_n15949_), .A2(new_n15950_), .B(new_n15956_), .ZN(new_n15957_));
  OR2_X2     g14955(.A1(new_n15890_), .A2(new_n15892_), .Z(new_n15958_));
  OAI21_X1   g14956(.A1(new_n15898_), .A2(new_n15897_), .B(new_n15838_), .ZN(new_n15959_));
  NAND3_X1   g14957(.A1(new_n15894_), .A2(new_n15895_), .A3(new_n10171_), .ZN(new_n15960_));
  NAND3_X1   g14958(.A1(new_n15958_), .A2(new_n15959_), .A3(new_n15960_), .ZN(new_n15961_));
  AOI21_X1   g14959(.A1(new_n15960_), .A2(new_n15959_), .B(new_n15958_), .ZN(new_n15962_));
  OAI21_X1   g14960(.A1(new_n15962_), .A2(new_n15914_), .B(new_n15961_), .ZN(new_n15963_));
  NOR3_X1    g14961(.A1(new_n15850_), .A2(new_n15855_), .A3(new_n10226_), .ZN(new_n15964_));
  AOI21_X1   g14962(.A1(new_n10225_), .A2(new_n15856_), .B(new_n10207_), .ZN(new_n15965_));
  NOR3_X1    g14963(.A1(new_n15737_), .A2(new_n15929_), .A3(new_n15928_), .ZN(new_n15966_));
  AOI21_X1   g14964(.A1(new_n15924_), .A2(new_n15738_), .B(new_n15689_), .ZN(new_n15967_));
  NOR2_X1    g14965(.A1(new_n15966_), .A2(new_n15967_), .ZN(new_n15968_));
  OAI21_X1   g14966(.A1(new_n15965_), .A2(new_n15964_), .B(new_n15968_), .ZN(new_n15969_));
  NOR3_X1    g14967(.A1(new_n15965_), .A2(new_n15964_), .A3(new_n15968_), .ZN(new_n15970_));
  AOI21_X1   g14968(.A1(new_n15963_), .A2(new_n15969_), .B(new_n15970_), .ZN(new_n15971_));
  NOR3_X1    g14969(.A1(new_n15942_), .A2(new_n15752_), .A3(new_n15739_), .ZN(new_n15972_));
  AOI21_X1   g14970(.A1(new_n15940_), .A2(new_n15751_), .B(new_n15935_), .ZN(new_n15973_));
  NOR2_X1    g14971(.A1(new_n15973_), .A2(new_n15972_), .ZN(new_n15974_));
  AOI21_X1   g14972(.A1(new_n10168_), .A2(new_n15947_), .B(new_n15857_), .ZN(new_n15975_));
  NOR3_X1    g14973(.A1(new_n15835_), .A2(new_n15945_), .A3(new_n10227_), .ZN(new_n15976_));
  OAI22_X1   g14974(.A1(new_n15971_), .A2(new_n15974_), .B1(new_n15975_), .B2(new_n15976_), .ZN(new_n15977_));
  NAND2_X1   g14975(.A1(new_n15971_), .A2(new_n15974_), .ZN(new_n15978_));
  NAND3_X1   g14976(.A1(new_n15753_), .A2(new_n15758_), .A3(new_n15686_), .ZN(new_n15979_));
  OAI21_X1   g14977(.A1(new_n15952_), .A2(new_n15953_), .B(new_n15951_), .ZN(new_n15980_));
  NAND2_X1   g14978(.A1(new_n15980_), .A2(new_n15979_), .ZN(new_n15981_));
  NAND3_X1   g14979(.A1(new_n15977_), .A2(new_n15978_), .A3(new_n15981_), .ZN(new_n15982_));
  NAND2_X1   g14980(.A1(new_n10412_), .A2(new_n15865_), .ZN(new_n15983_));
  NAND2_X1   g14981(.A1(new_n15983_), .A2(new_n10229_), .ZN(new_n15984_));
  NAND3_X1   g14982(.A1(new_n15859_), .A2(new_n10412_), .A3(new_n15865_), .ZN(new_n15985_));
  NAND2_X1   g14983(.A1(new_n15984_), .A2(new_n15985_), .ZN(new_n15986_));
  NAND2_X1   g14984(.A1(new_n15982_), .A2(new_n15986_), .ZN(new_n15987_));
  NAND2_X1   g14985(.A1(new_n15759_), .A2(new_n15686_), .ZN(new_n15988_));
  NOR2_X1    g14986(.A1(new_n15779_), .A2(new_n15771_), .ZN(new_n15989_));
  NOR2_X1    g14987(.A1(new_n15772_), .A2(new_n15777_), .ZN(new_n15990_));
  INV_X1     g14988(.I(new_n15801_), .ZN(new_n15991_));
  OAI22_X1   g14989(.A1(new_n15990_), .A2(new_n15989_), .B1(new_n15991_), .B2(new_n15799_), .ZN(new_n15992_));
  NAND2_X1   g14990(.A1(new_n15992_), .A2(new_n15802_), .ZN(new_n15993_));
  XOR2_X1    g14991(.A1(new_n15993_), .A2(new_n15988_), .Z(new_n15994_));
  AOI21_X1   g14992(.A1(new_n15987_), .A2(new_n15957_), .B(new_n15994_), .ZN(new_n15995_));
  AOI21_X1   g14993(.A1(new_n15977_), .A2(new_n15978_), .B(new_n15981_), .ZN(new_n15996_));
  AOI21_X1   g14994(.A1(new_n15982_), .A2(new_n15986_), .B(new_n15996_), .ZN(new_n15997_));
  NOR3_X1    g14995(.A1(new_n15872_), .A2(new_n15867_), .A3(new_n10466_), .ZN(new_n15998_));
  AOI22_X1   g14996(.A1(new_n10467_), .A2(new_n10465_), .B1(new_n15870_), .B2(new_n15871_), .ZN(new_n15999_));
  NOR3_X1    g14997(.A1(new_n15998_), .A2(new_n15999_), .A3(new_n10414_), .ZN(new_n16000_));
  NAND4_X1   g14998(.A1(new_n10467_), .A2(new_n10465_), .A3(new_n15871_), .A4(new_n15870_), .ZN(new_n16001_));
  OAI22_X1   g14999(.A1(new_n15867_), .A2(new_n10466_), .B1(new_n10484_), .B2(new_n10488_), .ZN(new_n16002_));
  AOI21_X1   g15000(.A1(new_n16001_), .A2(new_n16002_), .B(new_n15866_), .ZN(new_n16003_));
  NOR2_X1    g15001(.A1(new_n16000_), .A2(new_n16003_), .ZN(new_n16004_));
  AOI21_X1   g15002(.A1(new_n15997_), .A2(new_n15994_), .B(new_n16004_), .ZN(new_n16005_));
  NOR4_X1    g15003(.A1(new_n15990_), .A2(new_n15989_), .A3(new_n15991_), .A4(new_n15799_), .ZN(new_n16006_));
  NOR2_X1    g15004(.A1(new_n15988_), .A2(new_n16006_), .ZN(new_n16007_));
  INV_X1     g15005(.I(new_n15807_), .ZN(new_n16008_));
  NOR4_X1    g15006(.A1(new_n16008_), .A2(new_n15812_), .A3(new_n15813_), .A4(new_n15815_), .ZN(new_n16009_));
  XOR2_X1    g15007(.A1(new_n15819_), .A2(new_n15820_), .Z(new_n16010_));
  OAI21_X1   g15008(.A1(new_n16007_), .A2(new_n16009_), .B(new_n16010_), .ZN(new_n16011_));
  XNOR2_X1   g15009(.A1(new_n15819_), .A2(new_n15820_), .ZN(new_n16012_));
  NAND3_X1   g15010(.A1(new_n15803_), .A2(new_n15817_), .A3(new_n16012_), .ZN(new_n16013_));
  NAND2_X1   g15011(.A1(new_n16011_), .A2(new_n16013_), .ZN(new_n16014_));
  NAND2_X1   g15012(.A1(new_n10535_), .A2(new_n10524_), .ZN(new_n16015_));
  NAND3_X1   g15013(.A1(new_n10538_), .A2(new_n10534_), .A3(new_n10508_), .ZN(new_n16016_));
  AOI22_X1   g15014(.A1(new_n15873_), .A2(new_n15869_), .B1(new_n16015_), .B2(new_n16016_), .ZN(new_n16017_));
  AOI21_X1   g15015(.A1(new_n10534_), .A2(new_n10508_), .B(new_n10538_), .ZN(new_n16018_));
  AND3_X2    g15016(.A1(new_n10500_), .A2(new_n10496_), .A3(new_n10499_), .Z(new_n16019_));
  AOI22_X1   g15017(.A1(new_n16019_), .A2(new_n10501_), .B1(new_n10491_), .B2(new_n10459_), .ZN(new_n16020_));
  INV_X1     g15018(.I(new_n10533_), .ZN(new_n16021_));
  NOR3_X1    g15019(.A1(new_n16020_), .A2(new_n10531_), .A3(new_n16021_), .ZN(new_n16022_));
  NOR2_X1    g15020(.A1(new_n10526_), .A2(new_n10527_), .ZN(new_n16023_));
  NOR3_X1    g15021(.A1(new_n10524_), .A2(new_n16022_), .A3(new_n16023_), .ZN(new_n16024_));
  NOR4_X1    g15022(.A1(new_n10490_), .A2(new_n10469_), .A3(new_n16018_), .A4(new_n16024_), .ZN(new_n16025_));
  NOR3_X1    g15023(.A1(new_n16017_), .A2(new_n16025_), .A3(new_n16014_), .ZN(new_n16026_));
  NOR3_X1    g15024(.A1(new_n16005_), .A2(new_n15995_), .A3(new_n16026_), .ZN(new_n16027_));
  AOI21_X1   g15025(.A1(new_n15803_), .A2(new_n15817_), .B(new_n16012_), .ZN(new_n16028_));
  NOR3_X1    g15026(.A1(new_n16007_), .A2(new_n16009_), .A3(new_n16010_), .ZN(new_n16029_));
  NOR2_X1    g15027(.A1(new_n16029_), .A2(new_n16028_), .ZN(new_n16030_));
  OAI22_X1   g15028(.A1(new_n10490_), .A2(new_n10469_), .B1(new_n16018_), .B2(new_n16024_), .ZN(new_n16031_));
  NAND4_X1   g15029(.A1(new_n15873_), .A2(new_n15869_), .A3(new_n16015_), .A4(new_n16016_), .ZN(new_n16032_));
  AOI21_X1   g15030(.A1(new_n16031_), .A2(new_n16032_), .B(new_n16030_), .ZN(new_n16033_));
  NAND3_X1   g15031(.A1(new_n15828_), .A2(new_n15879_), .A3(new_n15826_), .ZN(new_n16034_));
  OAI21_X1   g15032(.A1(new_n16027_), .A2(new_n16033_), .B(new_n16034_), .ZN(new_n16035_));
  AOI21_X1   g15033(.A1(new_n16035_), .A2(new_n15881_), .B(new_n10547_), .ZN(new_n16036_));
  AOI21_X1   g15034(.A1(new_n15969_), .A2(new_n15933_), .B(new_n15963_), .ZN(new_n16037_));
  NOR3_X1    g15035(.A1(new_n15917_), .A2(new_n15970_), .A3(new_n15932_), .ZN(new_n16038_));
  AOI21_X1   g15036(.A1(new_n15913_), .A2(new_n15910_), .B(new_n15902_), .ZN(new_n16039_));
  NOR2_X1    g15037(.A1(new_n15911_), .A2(new_n15912_), .ZN(new_n16040_));
  NOR2_X1    g15038(.A1(new_n16040_), .A2(new_n16039_), .ZN(new_n16041_));
  INV_X1     g15039(.I(\A[1000] ), .ZN(new_n16042_));
  NOR2_X1    g15040(.A1(new_n15906_), .A2(new_n15904_), .ZN(new_n16043_));
  NOR3_X1    g15041(.A1(new_n15907_), .A2(new_n16042_), .A3(new_n16043_), .ZN(new_n16044_));
  INV_X1     g15042(.I(new_n16044_), .ZN(new_n16045_));
  NOR2_X1    g15043(.A1(new_n16041_), .A2(new_n16045_), .ZN(new_n16046_));
  NAND3_X1   g15044(.A1(new_n15915_), .A2(new_n15961_), .A3(new_n15916_), .ZN(new_n16047_));
  OAI21_X1   g15045(.A1(new_n15962_), .A2(new_n15900_), .B(new_n15914_), .ZN(new_n16048_));
  NAND3_X1   g15046(.A1(new_n16046_), .A2(new_n16048_), .A3(new_n16047_), .ZN(new_n16049_));
  OR3_X2     g15047(.A1(new_n16037_), .A2(new_n16038_), .A3(new_n16049_), .Z(new_n16050_));
  NAND2_X1   g15048(.A1(new_n15946_), .A2(new_n15948_), .ZN(new_n16051_));
  NOR2_X1    g15049(.A1(new_n16051_), .A2(new_n15944_), .ZN(new_n16052_));
  NOR2_X1    g15050(.A1(new_n15976_), .A2(new_n15975_), .ZN(new_n16053_));
  NOR2_X1    g15051(.A1(new_n16053_), .A2(new_n15974_), .ZN(new_n16054_));
  NOR3_X1    g15052(.A1(new_n16054_), .A2(new_n16052_), .A3(new_n15934_), .ZN(new_n16055_));
  NAND2_X1   g15053(.A1(new_n16053_), .A2(new_n15974_), .ZN(new_n16056_));
  NAND2_X1   g15054(.A1(new_n16051_), .A2(new_n15944_), .ZN(new_n16057_));
  AOI21_X1   g15055(.A1(new_n16056_), .A2(new_n16057_), .B(new_n15971_), .ZN(new_n16058_));
  NOR3_X1    g15056(.A1(new_n16058_), .A2(new_n16055_), .A3(new_n16050_), .ZN(new_n16059_));
  XOR2_X1    g15057(.A1(new_n15983_), .A2(new_n15859_), .Z(new_n16060_));
  NOR3_X1    g15058(.A1(new_n15949_), .A2(new_n15950_), .A3(new_n15956_), .ZN(new_n16061_));
  OAI21_X1   g15059(.A1(new_n16061_), .A2(new_n15996_), .B(new_n16060_), .ZN(new_n16062_));
  XOR2_X1    g15060(.A1(new_n15983_), .A2(new_n10229_), .Z(new_n16063_));
  NAND3_X1   g15061(.A1(new_n16063_), .A2(new_n15982_), .A3(new_n15957_), .ZN(new_n16064_));
  NAND3_X1   g15062(.A1(new_n16062_), .A2(new_n16059_), .A3(new_n16064_), .ZN(new_n16065_));
  NAND2_X1   g15063(.A1(new_n16002_), .A2(new_n16001_), .ZN(new_n16066_));
  XOR2_X1    g15064(.A1(new_n16066_), .A2(new_n10414_), .Z(new_n16067_));
  NAND3_X1   g15065(.A1(new_n15987_), .A2(new_n15994_), .A3(new_n15957_), .ZN(new_n16068_));
  AOI21_X1   g15066(.A1(new_n10412_), .A2(new_n15865_), .B(new_n15859_), .ZN(new_n16069_));
  NOR2_X1    g15067(.A1(new_n15983_), .A2(new_n10229_), .ZN(new_n16070_));
  NOR2_X1    g15068(.A1(new_n16070_), .A2(new_n16069_), .ZN(new_n16071_));
  OAI21_X1   g15069(.A1(new_n16061_), .A2(new_n16071_), .B(new_n15957_), .ZN(new_n16072_));
  XNOR2_X1   g15070(.A1(new_n15993_), .A2(new_n15988_), .ZN(new_n16073_));
  NAND2_X1   g15071(.A1(new_n16072_), .A2(new_n16073_), .ZN(new_n16074_));
  AOI21_X1   g15072(.A1(new_n16074_), .A2(new_n16068_), .B(new_n16067_), .ZN(new_n16075_));
  XOR2_X1    g15073(.A1(new_n16066_), .A2(new_n15866_), .Z(new_n16076_));
  NOR2_X1    g15074(.A1(new_n16072_), .A2(new_n16073_), .ZN(new_n16077_));
  NOR3_X1    g15075(.A1(new_n16077_), .A2(new_n15995_), .A3(new_n16076_), .ZN(new_n16078_));
  NOR3_X1    g15076(.A1(new_n16078_), .A2(new_n16075_), .A3(new_n16065_), .ZN(new_n16079_));
  NAND2_X1   g15077(.A1(new_n15873_), .A2(new_n15869_), .ZN(new_n16080_));
  XOR2_X1    g15078(.A1(new_n16014_), .A2(new_n16080_), .Z(new_n16081_));
  NOR2_X1    g15079(.A1(new_n16018_), .A2(new_n16024_), .ZN(new_n16082_));
  INV_X1     g15080(.I(new_n16082_), .ZN(new_n16083_));
  NAND3_X1   g15081(.A1(new_n16001_), .A2(new_n16002_), .A3(new_n15866_), .ZN(new_n16084_));
  OAI21_X1   g15082(.A1(new_n15998_), .A2(new_n15999_), .B(new_n10414_), .ZN(new_n16085_));
  NAND2_X1   g15083(.A1(new_n16085_), .A2(new_n16084_), .ZN(new_n16086_));
  OAI21_X1   g15084(.A1(new_n16072_), .A2(new_n16073_), .B(new_n16086_), .ZN(new_n16087_));
  NAND3_X1   g15085(.A1(new_n16087_), .A2(new_n16074_), .A3(new_n16083_), .ZN(new_n16088_));
  OAI21_X1   g15086(.A1(new_n16005_), .A2(new_n15995_), .B(new_n16082_), .ZN(new_n16089_));
  AOI21_X1   g15087(.A1(new_n16089_), .A2(new_n16088_), .B(new_n16081_), .ZN(new_n16090_));
  XOR2_X1    g15088(.A1(new_n16030_), .A2(new_n16080_), .Z(new_n16091_));
  NOR3_X1    g15089(.A1(new_n16005_), .A2(new_n15995_), .A3(new_n16082_), .ZN(new_n16092_));
  AOI21_X1   g15090(.A1(new_n16087_), .A2(new_n16074_), .B(new_n16083_), .ZN(new_n16093_));
  NOR3_X1    g15091(.A1(new_n16092_), .A2(new_n16093_), .A3(new_n16091_), .ZN(new_n16094_));
  OAI21_X1   g15092(.A1(new_n16094_), .A2(new_n16090_), .B(new_n16079_), .ZN(new_n16095_));
  AOI21_X1   g15093(.A1(new_n15876_), .A2(new_n15877_), .B(new_n15878_), .ZN(new_n16096_));
  NOR3_X1    g15094(.A1(new_n10530_), .A2(new_n10539_), .A3(new_n15827_), .ZN(new_n16097_));
  NOR3_X1    g15095(.A1(new_n16097_), .A2(new_n16096_), .A3(new_n15826_), .ZN(new_n16098_));
  INV_X1     g15096(.I(new_n15826_), .ZN(new_n16099_));
  AOI21_X1   g15097(.A1(new_n15828_), .A2(new_n15879_), .B(new_n16099_), .ZN(new_n16100_));
  NOR4_X1    g15098(.A1(new_n16027_), .A2(new_n16033_), .A3(new_n16098_), .A4(new_n16100_), .ZN(new_n16101_));
  NAND3_X1   g15099(.A1(new_n16032_), .A2(new_n16031_), .A3(new_n16030_), .ZN(new_n16102_));
  NAND3_X1   g15100(.A1(new_n16087_), .A2(new_n16074_), .A3(new_n16102_), .ZN(new_n16103_));
  INV_X1     g15101(.I(new_n16033_), .ZN(new_n16104_));
  NOR3_X1    g15102(.A1(new_n16097_), .A2(new_n16096_), .A3(new_n16099_), .ZN(new_n16105_));
  AOI21_X1   g15103(.A1(new_n16103_), .A2(new_n16104_), .B(new_n16105_), .ZN(new_n16106_));
  NAND2_X1   g15104(.A1(new_n10547_), .A2(new_n15880_), .ZN(new_n16107_));
  NOR4_X1    g15105(.A1(new_n16095_), .A2(new_n10547_), .A3(new_n16101_), .A4(new_n16107_), .ZN(new_n16108_));
  NOR3_X1    g15106(.A1(new_n16106_), .A2(new_n10546_), .A3(new_n15880_), .ZN(new_n16109_));
  NAND3_X1   g15107(.A1(new_n15828_), .A2(new_n15879_), .A3(new_n16099_), .ZN(new_n16110_));
  OAI21_X1   g15108(.A1(new_n16097_), .A2(new_n16096_), .B(new_n15826_), .ZN(new_n16111_));
  NAND4_X1   g15109(.A1(new_n16103_), .A2(new_n16104_), .A3(new_n16110_), .A4(new_n16111_), .ZN(new_n16112_));
  OAI22_X1   g15110(.A1(new_n16027_), .A2(new_n16033_), .B1(new_n16098_), .B2(new_n16100_), .ZN(new_n16113_));
  NAND2_X1   g15111(.A1(new_n16113_), .A2(new_n16112_), .ZN(new_n16114_));
  NOR4_X1    g15112(.A1(new_n16095_), .A2(new_n16036_), .A3(new_n16114_), .A4(new_n16109_), .ZN(new_n16115_));
  OAI21_X1   g15113(.A1(new_n16106_), .A2(new_n15880_), .B(new_n10546_), .ZN(new_n16116_));
  NAND3_X1   g15114(.A1(new_n16035_), .A2(new_n10547_), .A3(new_n15881_), .ZN(new_n16117_));
  NAND2_X1   g15115(.A1(new_n16117_), .A2(new_n16116_), .ZN(new_n16118_));
  NOR2_X1    g15116(.A1(new_n16095_), .A2(new_n16114_), .ZN(new_n16119_));
  NAND3_X1   g15117(.A1(new_n16056_), .A2(new_n16057_), .A3(new_n15971_), .ZN(new_n16120_));
  OAI21_X1   g15118(.A1(new_n16054_), .A2(new_n16052_), .B(new_n15934_), .ZN(new_n16121_));
  NAND2_X1   g15119(.A1(new_n16121_), .A2(new_n16120_), .ZN(new_n16122_));
  AOI21_X1   g15120(.A1(new_n15982_), .A2(new_n15957_), .B(new_n16063_), .ZN(new_n16123_));
  NOR3_X1    g15121(.A1(new_n16060_), .A2(new_n16061_), .A3(new_n15996_), .ZN(new_n16124_));
  NOR4_X1    g15122(.A1(new_n16123_), .A2(new_n16122_), .A3(new_n16124_), .A4(new_n16050_), .ZN(new_n16125_));
  OAI21_X1   g15123(.A1(new_n16077_), .A2(new_n15995_), .B(new_n16076_), .ZN(new_n16126_));
  NAND3_X1   g15124(.A1(new_n16074_), .A2(new_n16068_), .A3(new_n16067_), .ZN(new_n16127_));
  NAND2_X1   g15125(.A1(new_n16126_), .A2(new_n16127_), .ZN(new_n16128_));
  AND3_X2    g15126(.A1(new_n16121_), .A2(new_n16120_), .A3(new_n16050_), .Z(new_n16129_));
  AOI21_X1   g15127(.A1(new_n16121_), .A2(new_n16120_), .B(new_n16050_), .ZN(new_n16130_));
  INV_X1     g15128(.I(new_n16049_), .ZN(new_n16131_));
  XOR2_X1    g15129(.A1(new_n16041_), .A2(new_n16044_), .Z(new_n16132_));
  AOI21_X1   g15130(.A1(new_n16048_), .A2(new_n16047_), .B(new_n16046_), .ZN(new_n16133_));
  OAI21_X1   g15131(.A1(new_n16131_), .A2(new_n16133_), .B(new_n16132_), .ZN(new_n16134_));
  OAI21_X1   g15132(.A1(new_n16037_), .A2(new_n16038_), .B(new_n16049_), .ZN(new_n16135_));
  AND3_X2    g15133(.A1(new_n16050_), .A2(new_n16134_), .A3(new_n16135_), .Z(new_n16136_));
  NOR3_X1    g15134(.A1(new_n16129_), .A2(new_n16130_), .A3(new_n16136_), .ZN(new_n16137_));
  AOI21_X1   g15135(.A1(new_n16062_), .A2(new_n16064_), .B(new_n16059_), .ZN(new_n16138_));
  NOR4_X1    g15136(.A1(new_n16128_), .A2(new_n16125_), .A3(new_n16137_), .A4(new_n16138_), .ZN(new_n16139_));
  NAND3_X1   g15137(.A1(new_n16126_), .A2(new_n16127_), .A3(new_n16125_), .ZN(new_n16140_));
  OAI21_X1   g15138(.A1(new_n16092_), .A2(new_n16093_), .B(new_n16091_), .ZN(new_n16141_));
  NAND3_X1   g15139(.A1(new_n16089_), .A2(new_n16088_), .A3(new_n16081_), .ZN(new_n16142_));
  NAND3_X1   g15140(.A1(new_n16141_), .A2(new_n16142_), .A3(new_n16140_), .ZN(new_n16143_));
  NAND3_X1   g15141(.A1(new_n16095_), .A2(new_n16143_), .A3(new_n16139_), .ZN(new_n16144_));
  AOI21_X1   g15142(.A1(new_n16141_), .A2(new_n16142_), .B(new_n16140_), .ZN(new_n16145_));
  AOI22_X1   g15143(.A1(new_n16103_), .A2(new_n16104_), .B1(new_n16110_), .B2(new_n16111_), .ZN(new_n16146_));
  NOR2_X1    g15144(.A1(new_n16101_), .A2(new_n16146_), .ZN(new_n16147_));
  NOR2_X1    g15145(.A1(new_n16145_), .A2(new_n16147_), .ZN(new_n16148_));
  NOR4_X1    g15146(.A1(new_n16144_), .A2(new_n16148_), .A3(new_n16119_), .A4(new_n16118_), .ZN(new_n16149_));
  NOR4_X1    g15147(.A1(new_n16149_), .A2(new_n16036_), .A3(new_n16108_), .A4(new_n16115_), .ZN(new_n16150_));
  AOI22_X1   g15148(.A1(new_n16145_), .A2(new_n16147_), .B1(new_n16117_), .B2(new_n16116_), .ZN(new_n16151_));
  NOR2_X1    g15149(.A1(new_n16115_), .A2(new_n16151_), .ZN(new_n16152_));
  NOR2_X1    g15150(.A1(new_n16036_), .A2(new_n16109_), .ZN(new_n16153_));
  NAND2_X1   g15151(.A1(new_n16145_), .A2(new_n16147_), .ZN(new_n16154_));
  NOR2_X1    g15152(.A1(new_n16094_), .A2(new_n16090_), .ZN(new_n16155_));
  NOR3_X1    g15153(.A1(new_n16137_), .A2(new_n16125_), .A3(new_n16138_), .ZN(new_n16156_));
  INV_X1     g15154(.I(new_n16156_), .ZN(new_n16157_));
  OAI21_X1   g15155(.A1(new_n16078_), .A2(new_n16075_), .B(new_n16065_), .ZN(new_n16158_));
  INV_X1     g15156(.I(new_n16158_), .ZN(new_n16159_));
  NOR4_X1    g15157(.A1(new_n16155_), .A2(new_n16079_), .A3(new_n16157_), .A4(new_n16159_), .ZN(new_n16160_));
  NAND2_X1   g15158(.A1(new_n16095_), .A2(new_n16114_), .ZN(new_n16161_));
  NAND4_X1   g15159(.A1(new_n16160_), .A2(new_n16154_), .A3(new_n16161_), .A4(new_n16153_), .ZN(new_n16162_));
  NAND4_X1   g15160(.A1(new_n16095_), .A2(new_n16143_), .A3(new_n16147_), .A4(new_n16139_), .ZN(new_n16163_));
  NAND3_X1   g15161(.A1(new_n16158_), .A2(new_n16140_), .A3(new_n16156_), .ZN(new_n16164_));
  NAND3_X1   g15162(.A1(new_n16095_), .A2(new_n16143_), .A3(new_n16164_), .ZN(new_n16165_));
  NOR2_X1    g15163(.A1(new_n16129_), .A2(new_n16130_), .ZN(new_n16166_));
  NOR2_X1    g15164(.A1(new_n16131_), .A2(new_n16133_), .ZN(new_n16167_));
  XOR2_X1    g15165(.A1(new_n15905_), .A2(\A[1000] ), .Z(new_n16168_));
  XOR2_X1    g15166(.A1(new_n15904_), .A2(new_n10190_), .Z(new_n16169_));
  XOR2_X1    g15167(.A1(new_n16169_), .A2(new_n16168_), .Z(new_n16170_));
  NAND2_X1   g15168(.A1(new_n16132_), .A2(new_n16170_), .ZN(new_n16171_));
  AOI22_X1   g15169(.A1(new_n16050_), .A2(new_n16135_), .B1(new_n16167_), .B2(new_n16171_), .ZN(new_n16172_));
  NOR4_X1    g15170(.A1(new_n16125_), .A2(new_n16166_), .A3(new_n16138_), .A4(new_n16172_), .ZN(new_n16173_));
  NAND2_X1   g15171(.A1(new_n16139_), .A2(new_n16173_), .ZN(new_n16174_));
  AOI21_X1   g15172(.A1(new_n16165_), .A2(new_n16174_), .B(new_n16163_), .ZN(new_n16175_));
  OAI22_X1   g15173(.A1(new_n16175_), .A2(new_n16152_), .B1(new_n16162_), .B2(new_n16036_), .ZN(new_n16176_));
  NAND2_X1   g15174(.A1(new_n16176_), .A2(new_n16150_), .ZN(maj));
endmodule


