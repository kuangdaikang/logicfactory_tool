// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:27 2022

module jbp  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35,
    \v36.0 , \v36.1 , \v36.2 , \v36.3 , \v36.4 , \v36.5 , \v36.6 , \v36.7 ,
    \v36.8 , \v36.9 , \v36.10 , \v36.11 , \v36.12 , \v36.13 , \v36.14 ,
    \v36.15 , \v36.16 , \v36.17 , \v36.18 , \v36.19 , \v36.20 , \v36.21 ,
    \v36.22 , \v36.23 , \v36.24 , \v36.25 , \v36.26 , \v36.27 , \v36.28 ,
    \v36.29 , \v36.30 , \v36.31 , \v36.32 , \v36.33 , \v36.34 , \v36.35 ,
    \v36.36 , \v36.37 , \v36.38 , \v36.39 , \v36.40 , \v36.41 , \v36.42 ,
    \v36.43 , \v36.44 , \v36.45 , \v36.46 , \v36.47 , \v36.48 , \v36.49 ,
    \v36.50 , \v36.51 , \v36.52 , \v36.53 , \v36.54 , \v36.55 , \v36.56   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35;
  output \v36.0 , \v36.1 , \v36.2 , \v36.3 , \v36.4 , \v36.5 , \v36.6 ,
    \v36.7 , \v36.8 , \v36.9 , \v36.10 , \v36.11 , \v36.12 , \v36.13 ,
    \v36.14 , \v36.15 , \v36.16 , \v36.17 , \v36.18 , \v36.19 , \v36.20 ,
    \v36.21 , \v36.22 , \v36.23 , \v36.24 , \v36.25 , \v36.26 , \v36.27 ,
    \v36.28 , \v36.29 , \v36.30 , \v36.31 , \v36.32 , \v36.33 , \v36.34 ,
    \v36.35 , \v36.36 , \v36.37 , \v36.38 , \v36.39 , \v36.40 , \v36.41 ,
    \v36.42 , \v36.43 , \v36.44 , \v36.45 , \v36.46 , \v36.47 , \v36.48 ,
    \v36.49 , \v36.50 , \v36.51 , \v36.52 , \v36.53 , \v36.54 , \v36.55 ,
    \v36.56 ;
  wire new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n115_,
    new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n267_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n306_, new_n308_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n443_, new_n444_, new_n445_,
    new_n447_, new_n448_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n456_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n472_, new_n473_, new_n474_, new_n475_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_;
  assign new_n94_ = v1 & ~v9;
  assign new_n95_ = v8 & ~new_n94_;
  assign new_n96_ = ~v0 & ~new_n95_;
  assign new_n97_ = ~v34 & ~new_n96_;
  assign new_n98_ = ~v30 & new_n97_;
  assign new_n99_ = ~v29 & new_n98_;
  assign \v36.0  = v20 & new_n99_;
  assign new_n101_ = v3 & v10;
  assign new_n102_ = ~v12 & ~v13;
  assign new_n103_ = v11 & new_n102_;
  assign new_n104_ = new_n101_ & new_n103_;
  assign new_n105_ = ~v8 & ~new_n104_;
  assign new_n106_ = ~v34 & ~new_n105_;
  assign new_n107_ = ~v30 & new_n106_;
  assign new_n108_ = ~v29 & new_n107_;
  assign new_n109_ = v20 & new_n108_;
  assign new_n110_ = ~v9 & new_n109_;
  assign new_n111_ = v1 & new_n110_;
  assign new_n112_ = ~v0 & new_n111_;
  assign \v36.48  = v28 & v29;
  assign \v36.1  = new_n112_ | \v36.48 ;
  assign new_n115_ = ~v1 & v8;
  assign new_n116_ = v9 & ~new_n115_;
  assign new_n117_ = v11 & ~v12;
  assign new_n118_ = v3 & ~new_n117_;
  assign new_n119_ = v10 & ~new_n118_;
  assign new_n120_ = ~v11 & ~v12;
  assign new_n121_ = ~v10 & new_n120_;
  assign new_n122_ = ~new_n119_ & ~new_n121_;
  assign new_n123_ = ~v13 & ~new_n122_;
  assign new_n124_ = ~v8 & new_n123_;
  assign new_n125_ = v1 & new_n124_;
  assign new_n126_ = ~new_n116_ & ~new_n125_;
  assign new_n127_ = ~v34 & ~new_n126_;
  assign new_n128_ = ~v30 & new_n127_;
  assign new_n129_ = ~v29 & new_n128_;
  assign new_n130_ = v20 & new_n129_;
  assign new_n131_ = ~v0 & new_n130_;
  assign \v36.53  = ~v28 & v29;
  assign \v36.2  = new_n131_ | \v36.53 ;
  assign new_n134_ = ~v24 & v33;
  assign new_n135_ = v24 & ~v33;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = v29 & ~new_n136_;
  assign new_n138_ = ~v23 & new_n137_;
  assign new_n139_ = ~v29 & v33;
  assign new_n140_ = v23 & new_n139_;
  assign new_n141_ = ~new_n138_ & ~new_n140_;
  assign new_n142_ = ~v22 & ~new_n141_;
  assign new_n143_ = ~v29 & ~v33;
  assign new_n144_ = v22 & new_n143_;
  assign new_n145_ = ~new_n142_ & ~new_n144_;
  assign new_n146_ = v28 & ~new_n145_;
  assign new_n147_ = ~v21 & new_n146_;
  assign new_n148_ = v21 & ~v28;
  assign new_n149_ = v29 & v33;
  assign new_n150_ = new_n148_ & new_n149_;
  assign new_n151_ = ~new_n147_ & ~new_n150_;
  assign new_n152_ = ~v27 & ~new_n151_;
  assign new_n153_ = v27 & ~v28;
  assign new_n154_ = v29 & ~v33;
  assign new_n155_ = new_n153_ & new_n154_;
  assign new_n156_ = ~new_n152_ & ~new_n155_;
  assign new_n157_ = ~v26 & ~new_n156_;
  assign new_n158_ = v26 & ~v28;
  assign new_n159_ = new_n139_ & new_n158_;
  assign new_n160_ = ~new_n157_ & ~new_n159_;
  assign new_n161_ = ~v32 & ~new_n160_;
  assign new_n162_ = ~v28 & ~v29;
  assign new_n163_ = v32 & ~v33;
  assign new_n164_ = new_n162_ & new_n163_;
  assign new_n165_ = v31 & ~new_n164_;
  assign \v36.3  = new_n161_ | ~new_n165_;
  assign \v36.4  = v16 & v25;
  assign new_n168_ = ~v0 & v1;
  assign new_n169_ = ~v3 & new_n168_;
  assign new_n170_ = ~v8 & new_n169_;
  assign new_n171_ = ~v9 & new_n170_;
  assign new_n172_ = v10 & new_n171_;
  assign new_n173_ = v12 & new_n172_;
  assign new_n174_ = ~v13 & new_n173_;
  assign new_n175_ = v20 & new_n174_;
  assign new_n176_ = ~v29 & new_n175_;
  assign new_n177_ = ~v30 & new_n176_;
  assign \v36.5  = ~v34 & new_n177_;
  assign new_n179_ = v8 & ~v10;
  assign new_n180_ = v11 & v12;
  assign new_n181_ = new_n179_ & new_n180_;
  assign new_n182_ = ~v11 & v13;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = ~v1 & ~new_n183_;
  assign new_n185_ = v12 & v13;
  assign new_n186_ = ~new_n184_ & ~new_n185_;
  assign new_n187_ = v9 & ~new_n186_;
  assign new_n188_ = v10 & v13;
  assign new_n189_ = ~new_n187_ & ~new_n188_;
  assign new_n190_ = ~v30 & ~new_n189_;
  assign new_n191_ = ~v29 & new_n190_;
  assign \v36.6  = v0 & new_n191_;
  assign new_n193_ = v9 & ~new_n117_;
  assign new_n194_ = ~v10 & ~new_n193_;
  assign new_n195_ = ~v13 & ~new_n194_;
  assign new_n196_ = v1 & new_n195_;
  assign new_n197_ = v0 & new_n196_;
  assign new_n198_ = ~v8 & v11;
  assign new_n199_ = v12 & ~new_n198_;
  assign new_n200_ = ~v10 & new_n199_;
  assign new_n201_ = ~v9 & new_n200_;
  assign new_n202_ = ~new_n197_ & ~new_n201_;
  assign new_n203_ = ~v30 & ~new_n202_;
  assign \v36.7  = ~v29 & new_n203_;
  assign new_n205_ = ~v0 & ~new_n117_;
  assign new_n206_ = ~new_n181_ & ~new_n205_;
  assign new_n207_ = ~v13 & ~new_n206_;
  assign new_n208_ = ~v1 & new_n207_;
  assign new_n209_ = ~v0 & v12;
  assign new_n210_ = v13 & ~new_n209_;
  assign new_n211_ = ~v11 & new_n210_;
  assign new_n212_ = ~v10 & new_n211_;
  assign new_n213_ = v1 & new_n212_;
  assign new_n214_ = ~new_n208_ & ~new_n213_;
  assign new_n215_ = v9 & ~new_n214_;
  assign new_n216_ = ~v8 & ~v9;
  assign new_n217_ = ~v10 & new_n180_;
  assign new_n218_ = new_n216_ & new_n217_;
  assign new_n219_ = ~v0 & ~v1;
  assign new_n220_ = v10 & ~v13;
  assign new_n221_ = new_n219_ & new_n220_;
  assign new_n222_ = ~new_n218_ & ~new_n221_;
  assign new_n223_ = ~new_n215_ & new_n222_;
  assign new_n224_ = ~v30 & ~new_n223_;
  assign \v36.8  = v29 | new_n224_;
  assign new_n226_ = v1 & ~new_n185_;
  assign new_n227_ = ~v0 & ~new_n226_;
  assign new_n228_ = ~v10 & ~v11;
  assign new_n229_ = v1 & new_n228_;
  assign new_n230_ = v13 & ~new_n229_;
  assign new_n231_ = ~v30 & ~new_n230_;
  assign new_n232_ = ~new_n194_ & new_n231_;
  assign new_n233_ = ~new_n227_ & new_n232_;
  assign \v36.9  = ~v29 & ~new_n233_;
  assign new_n235_ = v1 & ~v13;
  assign new_n236_ = ~new_n198_ & ~new_n235_;
  assign new_n237_ = v0 & ~new_n236_;
  assign new_n238_ = ~v1 & v13;
  assign new_n239_ = ~v0 & new_n238_;
  assign new_n240_ = ~new_n237_ & ~new_n239_;
  assign new_n241_ = v9 & ~new_n240_;
  assign new_n242_ = ~v1 & v11;
  assign new_n243_ = ~v0 & new_n242_;
  assign new_n244_ = v9 & ~new_n243_;
  assign new_n245_ = v8 & ~new_n244_;
  assign new_n246_ = ~v9 & ~v11;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = ~v10 & ~new_n247_;
  assign new_n249_ = ~new_n241_ & ~new_n248_;
  assign new_n250_ = v12 & ~new_n249_;
  assign new_n251_ = v9 & ~v11;
  assign new_n252_ = v0 & new_n251_;
  assign new_n253_ = ~new_n188_ & ~new_n252_;
  assign new_n254_ = ~v1 & ~new_n253_;
  assign new_n255_ = v9 & new_n120_;
  assign new_n256_ = ~v10 & ~new_n255_;
  assign new_n257_ = v0 & ~new_n256_;
  assign new_n258_ = v9 & ~v10;
  assign new_n259_ = ~v12 & v13;
  assign new_n260_ = ~v11 & new_n259_;
  assign new_n261_ = new_n258_ & new_n260_;
  assign new_n262_ = ~new_n257_ & ~new_n261_;
  assign new_n263_ = ~new_n254_ & new_n262_;
  assign new_n264_ = ~new_n250_ & new_n263_;
  assign new_n265_ = ~v30 & ~new_n264_;
  assign \v36.10  = v29 | new_n265_;
  assign new_n267_ = ~v30 & ~new_n194_;
  assign \v36.11  = ~v29 & new_n267_;
  assign new_n269_ = ~v11 & v30;
  assign new_n270_ = v7 & new_n269_;
  assign new_n271_ = v1 & v3;
  assign new_n272_ = ~v0 & new_n271_;
  assign new_n273_ = ~v9 & ~v10;
  assign new_n274_ = ~v8 & new_n273_;
  assign new_n275_ = new_n272_ & new_n274_;
  assign new_n276_ = v12 & ~v13;
  assign new_n277_ = v11 & new_n276_;
  assign new_n278_ = v20 & ~v29;
  assign new_n279_ = ~v30 & ~v34;
  assign new_n280_ = new_n278_ & new_n279_;
  assign new_n281_ = new_n277_ & new_n280_;
  assign new_n282_ = new_n275_ & new_n281_;
  assign \v36.12  = new_n270_ | new_n282_;
  assign new_n284_ = ~v8 & new_n168_;
  assign new_n285_ = v9 & new_n284_;
  assign new_n286_ = v20 & new_n285_;
  assign new_n287_ = ~v29 & new_n286_;
  assign new_n288_ = ~v30 & new_n287_;
  assign \v36.13  = ~v34 & new_n288_;
  assign new_n290_ = ~v11 & v12;
  assign new_n291_ = ~v10 & new_n290_;
  assign new_n292_ = v3 & v11;
  assign new_n293_ = ~v3 & v12;
  assign new_n294_ = ~new_n292_ & ~new_n293_;
  assign new_n295_ = v10 & ~new_n294_;
  assign new_n296_ = ~new_n291_ & ~new_n295_;
  assign new_n297_ = ~v34 & ~new_n296_;
  assign new_n298_ = ~v30 & new_n297_;
  assign new_n299_ = ~v29 & new_n298_;
  assign new_n300_ = v20 & new_n299_;
  assign new_n301_ = ~v13 & new_n300_;
  assign new_n302_ = ~v9 & new_n301_;
  assign new_n303_ = ~v8 & new_n302_;
  assign new_n304_ = v1 & new_n303_;
  assign \v36.14  = ~v0 & new_n304_;
  assign new_n306_ = v19 & v28;
  assign \v36.15  = v29 & new_n306_;
  assign new_n308_ = ~v30 & new_n162_;
  assign \v36.16  = v34 & new_n308_;
  assign new_n310_ = v8 & new_n168_;
  assign new_n311_ = ~v9 & new_n310_;
  assign new_n312_ = v20 & new_n311_;
  assign new_n313_ = ~v29 & new_n312_;
  assign new_n314_ = ~v30 & new_n313_;
  assign \v36.17  = ~v34 & new_n314_;
  assign new_n316_ = ~v7 & v30;
  assign new_n317_ = v3 & new_n216_;
  assign new_n318_ = new_n168_ & new_n317_;
  assign new_n319_ = ~v13 & v20;
  assign new_n320_ = ~v10 & new_n319_;
  assign new_n321_ = ~v29 & new_n279_;
  assign new_n322_ = new_n320_ & new_n321_;
  assign new_n323_ = new_n318_ & new_n322_;
  assign new_n324_ = ~new_n316_ & ~new_n323_;
  assign new_n325_ = v11 & ~new_n324_;
  assign \v36.18  = new_n270_ | new_n325_;
  assign new_n327_ = v20 & new_n279_;
  assign new_n328_ = ~v29 & ~new_n327_;
  assign new_n329_ = v2 & ~v3;
  assign new_n330_ = ~v2 & v3;
  assign new_n331_ = ~new_n329_ & ~new_n330_;
  assign new_n332_ = ~new_n328_ & ~new_n331_;
  assign new_n333_ = v15 & new_n332_;
  assign new_n334_ = v14 & new_n333_;
  assign new_n335_ = v13 & new_n334_;
  assign new_n336_ = v8 & new_n335_;
  assign new_n337_ = ~v1 & new_n336_;
  assign new_n338_ = ~v0 & new_n337_;
  assign \v36.19  = \v36.53  | new_n338_;
  assign \v36.21  = ~v16 & v25;
  assign new_n341_ = v7 & ~v9;
  assign new_n342_ = v3 & new_n341_;
  assign new_n343_ = new_n120_ & new_n258_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign new_n345_ = ~v8 & ~new_n344_;
  assign new_n346_ = ~v7 & v9;
  assign new_n347_ = new_n121_ & new_n346_;
  assign new_n348_ = ~new_n345_ & ~new_n347_;
  assign new_n349_ = ~v1 & ~new_n348_;
  assign new_n350_ = v1 & v8;
  assign \v36.22  = new_n349_ | new_n350_;
  assign new_n352_ = v4 & ~v9;
  assign new_n353_ = ~new_n343_ & ~new_n352_;
  assign new_n354_ = ~v8 & ~new_n353_;
  assign new_n355_ = ~v1 & ~new_n354_;
  assign new_n356_ = v7 & ~new_n355_;
  assign new_n357_ = ~v1 & new_n346_;
  assign new_n358_ = new_n291_ & new_n357_;
  assign \v36.23  = new_n356_ | new_n358_;
  assign new_n360_ = v5 & ~v9;
  assign new_n361_ = ~v1 & new_n360_;
  assign new_n362_ = ~new_n343_ & ~new_n361_;
  assign new_n363_ = ~v8 & ~new_n362_;
  assign new_n364_ = v7 & new_n363_;
  assign new_n365_ = ~v7 & ~v10;
  assign new_n366_ = new_n117_ & new_n365_;
  assign new_n367_ = ~v1 & ~new_n366_;
  assign new_n368_ = v9 & ~new_n367_;
  assign \v36.24  = new_n364_ | new_n368_;
  assign new_n370_ = v6 & ~v9;
  assign new_n371_ = ~new_n343_ & ~new_n370_;
  assign new_n372_ = ~v8 & ~new_n371_;
  assign new_n373_ = v7 & new_n372_;
  assign new_n374_ = new_n217_ & new_n346_;
  assign new_n375_ = ~new_n373_ & ~new_n374_;
  assign new_n376_ = ~v1 & ~new_n375_;
  assign new_n377_ = v1 & v13;
  assign \v36.25  = new_n376_ | new_n377_;
  assign new_n379_ = v1 & v14;
  assign new_n380_ = v3 & v9;
  assign new_n381_ = new_n120_ & new_n273_;
  assign new_n382_ = ~new_n380_ & ~new_n381_;
  assign new_n383_ = ~v8 & ~new_n382_;
  assign new_n384_ = v7 & new_n383_;
  assign new_n385_ = v10 & new_n120_;
  assign new_n386_ = new_n346_ & new_n385_;
  assign new_n387_ = ~new_n384_ & ~new_n386_;
  assign new_n388_ = ~v1 & ~new_n387_;
  assign \v36.26  = new_n379_ | new_n388_;
  assign new_n390_ = v1 & v15;
  assign new_n391_ = v4 & v9;
  assign new_n392_ = ~new_n381_ & ~new_n391_;
  assign new_n393_ = ~v8 & ~new_n392_;
  assign new_n394_ = v7 & new_n393_;
  assign new_n395_ = v10 & new_n290_;
  assign new_n396_ = new_n346_ & new_n395_;
  assign new_n397_ = ~new_n394_ & ~new_n396_;
  assign new_n398_ = ~v1 & ~new_n397_;
  assign \v36.27  = new_n390_ | new_n398_;
  assign new_n400_ = v0 & v1;
  assign new_n401_ = v5 & v9;
  assign new_n402_ = ~new_n381_ & ~new_n401_;
  assign new_n403_ = ~v8 & ~new_n402_;
  assign new_n404_ = v7 & new_n403_;
  assign new_n405_ = v10 & new_n117_;
  assign new_n406_ = new_n346_ & new_n405_;
  assign new_n407_ = ~new_n404_ & ~new_n406_;
  assign new_n408_ = ~v1 & ~new_n407_;
  assign \v36.28  = new_n400_ | new_n408_;
  assign new_n410_ = v1 & v2;
  assign new_n411_ = v6 & v9;
  assign new_n412_ = ~new_n381_ & ~new_n411_;
  assign new_n413_ = ~v8 & ~new_n412_;
  assign new_n414_ = v7 & new_n413_;
  assign new_n415_ = v10 & new_n180_;
  assign new_n416_ = new_n346_ & new_n415_;
  assign new_n417_ = ~new_n414_ & ~new_n416_;
  assign new_n418_ = ~v1 & ~new_n417_;
  assign \v36.29  = new_n410_ | new_n418_;
  assign new_n420_ = v10 & ~v12;
  assign new_n421_ = ~v34 & ~new_n420_;
  assign new_n422_ = ~v29 & new_n421_;
  assign new_n423_ = v20 & new_n422_;
  assign new_n424_ = ~v13 & new_n423_;
  assign new_n425_ = v11 & new_n424_;
  assign new_n426_ = ~v9 & new_n425_;
  assign new_n427_ = ~v8 & new_n426_;
  assign new_n428_ = v3 & new_n427_;
  assign new_n429_ = v1 & new_n428_;
  assign new_n430_ = ~v0 & new_n429_;
  assign \v36.30  = v30 | new_n430_;
  assign new_n432_ = ~v34 & ~new_n118_;
  assign new_n433_ = ~v30 & new_n432_;
  assign new_n434_ = ~v29 & new_n433_;
  assign new_n435_ = v20 & new_n434_;
  assign new_n436_ = ~v13 & new_n435_;
  assign new_n437_ = v10 & new_n436_;
  assign new_n438_ = ~v9 & new_n437_;
  assign new_n439_ = ~v8 & new_n438_;
  assign new_n440_ = v1 & new_n439_;
  assign new_n441_ = ~v0 & new_n440_;
  assign \v36.31  = \v36.53  | new_n441_;
  assign new_n443_ = ~v21 & ~v26;
  assign new_n444_ = ~v27 & ~v32;
  assign new_n445_ = new_n443_ & new_n444_;
  assign \v36.32  = ~v31 | new_n445_;
  assign new_n447_ = ~v27 & new_n443_;
  assign new_n448_ = v31 & new_n447_;
  assign \v36.33  = ~v32 & new_n448_;
  assign new_n450_ = ~v22 & ~v23;
  assign new_n451_ = ~v27 & ~new_n450_;
  assign new_n452_ = ~v21 & new_n451_;
  assign new_n453_ = ~v32 & ~new_n452_;
  assign new_n454_ = ~v26 & new_n453_;
  assign \v36.34  = ~v31 | new_n454_;
  assign new_n456_ = v31 & new_n453_;
  assign \v36.35  = ~v26 & new_n456_;
  assign new_n458_ = ~v23 & v24;
  assign new_n459_ = ~v22 & ~new_n458_;
  assign new_n460_ = ~v21 & ~new_n459_;
  assign new_n461_ = ~v27 & ~new_n460_;
  assign new_n462_ = ~v26 & ~new_n461_;
  assign new_n463_ = ~v32 & ~new_n462_;
  assign \v36.36  = v31 & ~new_n463_;
  assign \v36.37  = v31 & new_n463_;
  assign new_n466_ = ~v0 & ~v8;
  assign new_n467_ = v9 & new_n466_;
  assign new_n468_ = v20 & new_n467_;
  assign new_n469_ = ~v29 & new_n468_;
  assign new_n470_ = ~v30 & new_n469_;
  assign \v36.38  = ~v34 & new_n470_;
  assign new_n472_ = ~v13 & new_n172_;
  assign new_n473_ = v20 & new_n472_;
  assign new_n474_ = ~v29 & new_n473_;
  assign new_n475_ = ~v30 & new_n474_;
  assign \v36.39  = ~v34 & new_n475_;
  assign new_n477_ = v3 & new_n168_;
  assign new_n478_ = ~v8 & new_n477_;
  assign new_n479_ = ~v9 & new_n478_;
  assign new_n480_ = ~v10 & new_n479_;
  assign new_n481_ = ~v11 & new_n480_;
  assign new_n482_ = ~v13 & new_n481_;
  assign new_n483_ = v20 & new_n482_;
  assign new_n484_ = ~v29 & new_n483_;
  assign new_n485_ = ~v30 & new_n484_;
  assign \v36.40  = ~v34 & new_n485_;
  assign new_n487_ = v9 & v12;
  assign new_n488_ = ~v10 & ~new_n487_;
  assign new_n489_ = v17 & ~new_n488_;
  assign new_n490_ = v1 & new_n489_;
  assign new_n491_ = v8 & v9;
  assign new_n492_ = ~v1 & new_n491_;
  assign new_n493_ = new_n217_ & new_n492_;
  assign new_n494_ = ~new_n490_ & ~new_n493_;
  assign new_n495_ = v13 & ~new_n494_;
  assign new_n496_ = ~v10 & v11;
  assign new_n497_ = v12 & v17;
  assign new_n498_ = new_n496_ & new_n497_;
  assign new_n499_ = new_n492_ & new_n498_;
  assign new_n500_ = ~new_n495_ & ~new_n499_;
  assign new_n501_ = ~v30 & ~new_n500_;
  assign new_n502_ = ~v29 & new_n501_;
  assign \v36.41  = v0 & new_n502_;
  assign new_n504_ = ~v9 & new_n284_;
  assign new_n505_ = ~v10 & new_n504_;
  assign new_n506_ = ~v11 & new_n505_;
  assign new_n507_ = v12 & new_n506_;
  assign new_n508_ = ~v13 & new_n507_;
  assign new_n509_ = v20 & new_n508_;
  assign new_n510_ = ~v29 & new_n509_;
  assign new_n511_ = ~v30 & new_n510_;
  assign \v36.42  = ~v34 & new_n511_;
  assign new_n513_ = ~v13 & new_n506_;
  assign new_n514_ = v20 & new_n513_;
  assign new_n515_ = ~v29 & new_n514_;
  assign new_n516_ = ~v30 & new_n515_;
  assign \v36.43  = ~v34 & new_n516_;
  assign new_n518_ = ~v1 & ~new_n405_;
  assign new_n519_ = ~v34 & ~new_n518_;
  assign new_n520_ = ~v30 & new_n519_;
  assign new_n521_ = ~v29 & new_n520_;
  assign new_n522_ = v20 & new_n521_;
  assign new_n523_ = v9 & new_n522_;
  assign new_n524_ = v8 & new_n523_;
  assign \v36.44  = ~v0 & new_n524_;
  assign new_n526_ = v1 & v9;
  assign new_n527_ = new_n115_ & new_n415_;
  assign new_n528_ = ~new_n526_ & ~new_n527_;
  assign new_n529_ = ~v0 & new_n528_;
  assign new_n530_ = ~v34 & ~new_n529_;
  assign new_n531_ = ~v30 & new_n530_;
  assign new_n532_ = ~v29 & new_n531_;
  assign \v36.45  = v20 & new_n532_;
  assign new_n534_ = ~v12 & v18;
  assign new_n535_ = v12 & ~v18;
  assign new_n536_ = ~new_n534_ & ~new_n535_;
  assign new_n537_ = v10 & ~new_n536_;
  assign new_n538_ = ~v12 & v35;
  assign new_n539_ = v12 & ~v35;
  assign new_n540_ = ~new_n538_ & ~new_n539_;
  assign new_n541_ = ~v10 & ~new_n540_;
  assign new_n542_ = ~new_n537_ & ~new_n541_;
  assign new_n543_ = ~v11 & ~new_n542_;
  assign new_n544_ = ~v12 & v17;
  assign new_n545_ = v12 & ~v17;
  assign new_n546_ = ~new_n544_ & ~new_n545_;
  assign new_n547_ = v11 & ~new_n546_;
  assign new_n548_ = ~v10 & new_n547_;
  assign new_n549_ = ~new_n543_ & ~new_n548_;
  assign new_n550_ = ~v34 & ~new_n549_;
  assign new_n551_ = ~v30 & new_n550_;
  assign new_n552_ = ~v29 & new_n551_;
  assign new_n553_ = v20 & new_n552_;
  assign new_n554_ = v13 & new_n553_;
  assign new_n555_ = ~v9 & new_n554_;
  assign new_n556_ = ~v8 & new_n555_;
  assign new_n557_ = v1 & new_n556_;
  assign \v36.46  = ~v0 & new_n557_;
  assign new_n559_ = v1 & new_n491_;
  assign new_n560_ = ~v0 & ~new_n559_;
  assign new_n561_ = ~new_n420_ & ~new_n560_;
  assign new_n562_ = ~v9 & ~v12;
  assign new_n563_ = new_n219_ & new_n562_;
  assign new_n564_ = ~new_n487_ & ~new_n563_;
  assign new_n565_ = v11 & ~new_n564_;
  assign new_n566_ = v10 & new_n565_;
  assign new_n567_ = v8 & new_n566_;
  assign new_n568_ = v1 & new_n216_;
  assign new_n569_ = new_n228_ & new_n276_;
  assign new_n570_ = new_n568_ & new_n569_;
  assign new_n571_ = ~new_n567_ & ~new_n570_;
  assign new_n572_ = ~new_n561_ & new_n571_;
  assign new_n573_ = ~v34 & ~new_n572_;
  assign new_n574_ = ~v30 & new_n573_;
  assign new_n575_ = ~v29 & new_n574_;
  assign \v36.47  = v20 & new_n575_;
  assign new_n577_ = ~v12 & new_n172_;
  assign new_n578_ = ~v13 & new_n577_;
  assign new_n579_ = v20 & new_n578_;
  assign new_n580_ = ~v29 & new_n579_;
  assign new_n581_ = ~v30 & new_n580_;
  assign \v36.49  = ~v34 & new_n581_;
  assign new_n583_ = ~v12 & new_n506_;
  assign new_n584_ = ~v13 & new_n583_;
  assign new_n585_ = v20 & new_n584_;
  assign new_n586_ = ~v29 & new_n585_;
  assign new_n587_ = ~v30 & new_n586_;
  assign \v36.50  = ~v34 & new_n587_;
  assign new_n589_ = ~v0 & ~new_n350_;
  assign new_n590_ = ~new_n420_ & ~new_n589_;
  assign new_n591_ = v11 & ~v13;
  assign new_n592_ = v3 & new_n591_;
  assign new_n593_ = ~v8 & ~new_n592_;
  assign new_n594_ = v1 & ~new_n593_;
  assign new_n595_ = v8 & v10;
  assign new_n596_ = new_n117_ & new_n595_;
  assign new_n597_ = ~new_n594_ & ~new_n596_;
  assign new_n598_ = ~v0 & ~new_n597_;
  assign new_n599_ = ~v3 & v10;
  assign new_n600_ = ~new_n228_ & ~new_n599_;
  assign new_n601_ = ~v13 & ~new_n600_;
  assign new_n602_ = v12 & new_n601_;
  assign new_n603_ = v1 & new_n602_;
  assign new_n604_ = ~new_n598_ & ~new_n603_;
  assign new_n605_ = ~v9 & ~new_n604_;
  assign new_n606_ = new_n415_ & new_n491_;
  assign new_n607_ = ~new_n605_ & ~new_n606_;
  assign new_n608_ = ~new_n590_ & new_n607_;
  assign new_n609_ = ~v34 & ~new_n608_;
  assign new_n610_ = v20 & new_n609_;
  assign new_n611_ = ~v29 & ~v30;
  assign \v36.51  = new_n610_ | ~new_n611_;
  assign new_n613_ = ~v34 & ~new_n216_;
  assign new_n614_ = ~v30 & new_n613_;
  assign new_n615_ = ~v29 & new_n614_;
  assign new_n616_ = v20 & new_n615_;
  assign new_n617_ = ~v1 & new_n616_;
  assign \v36.52  = ~v0 & new_n617_;
  assign new_n619_ = ~v1 & ~v8;
  assign new_n620_ = ~new_n350_ & ~new_n619_;
  assign new_n621_ = ~v34 & ~new_n620_;
  assign new_n622_ = ~v30 & new_n621_;
  assign new_n623_ = ~v29 & new_n622_;
  assign new_n624_ = v20 & new_n623_;
  assign new_n625_ = ~v9 & new_n624_;
  assign \v36.54  = ~v0 & new_n625_;
  assign new_n627_ = ~v30 & new_n421_;
  assign new_n628_ = ~v29 & new_n627_;
  assign new_n629_ = v20 & new_n628_;
  assign new_n630_ = v8 & new_n629_;
  assign new_n631_ = ~v1 & new_n630_;
  assign \v36.55  = ~v0 & new_n631_;
  assign new_n633_ = ~v10 & new_n591_;
  assign new_n634_ = ~v29 & ~v34;
  assign new_n635_ = v20 & new_n634_;
  assign new_n636_ = new_n633_ & new_n635_;
  assign new_n637_ = new_n318_ & new_n636_;
  assign \v36.56  = v30 | new_n637_;
  assign \v36.20  = v31;
endmodule


