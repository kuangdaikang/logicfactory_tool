// Benchmark "square" written by ABC on Mon Sep  4 17:36:38 2023

module square ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ;
  output \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127] ;
  wire new_n194_, new_n196_, new_n197_, new_n198_, new_n199_, new_n201_,
    new_n202_, new_n203_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_,
    new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_,
    new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_,
    new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_,
    new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_,
    new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_,
    new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_,
    new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_,
    new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_,
    new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_,
    new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_,
    new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_,
    new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_,
    new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2886_, new_n2887_, new_n2888_,
    new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_,
    new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3019_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_,
    new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_,
    new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_,
    new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_,
    new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_,
    new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_,
    new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_,
    new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_,
    new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_,
    new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_,
    new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_,
    new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_,
    new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_,
    new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_,
    new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_,
    new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_,
    new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_,
    new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_,
    new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_,
    new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_,
    new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_,
    new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_,
    new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_,
    new_n3311_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_,
    new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_,
    new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_,
    new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_,
    new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_,
    new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_,
    new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_,
    new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_,
    new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_,
    new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_,
    new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_,
    new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_,
    new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_,
    new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_,
    new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_,
    new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_,
    new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_,
    new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_,
    new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_,
    new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_,
    new_n3770_, new_n3771_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_,
    new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_,
    new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_,
    new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_,
    new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_,
    new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_,
    new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_,
    new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_,
    new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_,
    new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_,
    new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_,
    new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4075_, new_n4076_, new_n4077_, new_n4078_,
    new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_,
    new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_,
    new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_,
    new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_,
    new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_,
    new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_,
    new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_,
    new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_,
    new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_,
    new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_,
    new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_,
    new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_,
    new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_,
    new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_,
    new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_,
    new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_,
    new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_,
    new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_,
    new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_,
    new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_,
    new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_,
    new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_,
    new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_,
    new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_,
    new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_,
    new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_,
    new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_,
    new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_,
    new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_,
    new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_,
    new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_,
    new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_,
    new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_,
    new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_,
    new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_,
    new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_,
    new_n4585_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_,
    new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_,
    new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_,
    new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_,
    new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_,
    new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_,
    new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_,
    new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_,
    new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_,
    new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_,
    new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_,
    new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_,
    new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_,
    new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_,
    new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_,
    new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_,
    new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_,
    new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_,
    new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_,
    new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_,
    new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_,
    new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_,
    new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_,
    new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_,
    new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_,
    new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_,
    new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_,
    new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_,
    new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_,
    new_n5122_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_,
    new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_,
    new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_,
    new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_,
    new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_,
    new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_,
    new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_,
    new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_,
    new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_,
    new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_,
    new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_,
    new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_,
    new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_,
    new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_,
    new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_,
    new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_,
    new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_,
    new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_,
    new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_,
    new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_,
    new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_,
    new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_,
    new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_,
    new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_,
    new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_,
    new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_,
    new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_,
    new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_,
    new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_,
    new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_,
    new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_,
    new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_,
    new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_,
    new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_,
    new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_,
    new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_,
    new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_,
    new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_,
    new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_,
    new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_,
    new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_,
    new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5851_, new_n5852_,
    new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_,
    new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_,
    new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_,
    new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_,
    new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_,
    new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_,
    new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_,
    new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_,
    new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_,
    new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_,
    new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_,
    new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_,
    new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_,
    new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_,
    new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_,
    new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_,
    new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_,
    new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_,
    new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_,
    new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_,
    new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_,
    new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_,
    new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_,
    new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_,
    new_n6045_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_,
    new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_,
    new_n6256_, new_n6257_, new_n6258_, new_n6260_, new_n6261_, new_n6262_,
    new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_,
    new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_,
    new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_,
    new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_,
    new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_,
    new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_,
    new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_,
    new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_,
    new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_,
    new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_,
    new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_,
    new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_,
    new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_,
    new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_,
    new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_,
    new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_,
    new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_,
    new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_,
    new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_,
    new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_,
    new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_,
    new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_,
    new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_,
    new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_,
    new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7104_, new_n7105_, new_n7106_,
    new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_,
    new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_,
    new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_,
    new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_,
    new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_,
    new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_,
    new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_,
    new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_,
    new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_,
    new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_,
    new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_,
    new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_,
    new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_,
    new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_,
    new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_,
    new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_,
    new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_,
    new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_,
    new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_,
    new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_,
    new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_,
    new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_,
    new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_,
    new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_,
    new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_,
    new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_,
    new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_,
    new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7538_, new_n7539_, new_n7540_,
    new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_,
    new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_,
    new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_,
    new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_,
    new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_,
    new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_,
    new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_,
    new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_,
    new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_,
    new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_,
    new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_,
    new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_,
    new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_,
    new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_,
    new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_,
    new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_,
    new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_,
    new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_,
    new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_,
    new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_,
    new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_,
    new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_,
    new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_,
    new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_,
    new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_,
    new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_,
    new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_,
    new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_,
    new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_,
    new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_,
    new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_,
    new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_,
    new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_,
    new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_,
    new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_,
    new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_,
    new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_,
    new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_,
    new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_,
    new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7949_, new_n7950_,
    new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_,
    new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_,
    new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_,
    new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_,
    new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_,
    new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_,
    new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_,
    new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_,
    new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_,
    new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_,
    new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_,
    new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_,
    new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_,
    new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_,
    new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_,
    new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_,
    new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_,
    new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_,
    new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_,
    new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_,
    new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_,
    new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_,
    new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_,
    new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_,
    new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_,
    new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_,
    new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_,
    new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_,
    new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_,
    new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_,
    new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_,
    new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_,
    new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_,
    new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_,
    new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_,
    new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_,
    new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_,
    new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_,
    new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_,
    new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_,
    new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_,
    new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_,
    new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_,
    new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_,
    new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_,
    new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_,
    new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_,
    new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_,
    new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_,
    new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_,
    new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_,
    new_n8342_, new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_,
    new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_,
    new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_,
    new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_,
    new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_,
    new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_,
    new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_,
    new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_,
    new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_,
    new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_, new_n8402_,
    new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_,
    new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_,
    new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_,
    new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_,
    new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_, new_n8432_,
    new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_, new_n8438_,
    new_n8439_, new_n8440_, new_n8441_, new_n8442_, new_n8443_, new_n8444_,
    new_n8445_, new_n8446_, new_n8447_, new_n8448_, new_n8449_, new_n8450_,
    new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_,
    new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8461_, new_n8462_,
    new_n8463_, new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_,
    new_n8469_, new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_,
    new_n8475_, new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_,
    new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_,
    new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_,
    new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_,
    new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_,
    new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_,
    new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_,
    new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_,
    new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_,
    new_n8529_, new_n8530_, new_n8531_, new_n8533_, new_n8534_, new_n8535_,
    new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_,
    new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_,
    new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_,
    new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_,
    new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_,
    new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_,
    new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_,
    new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_,
    new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_,
    new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_,
    new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_,
    new_n8632_, new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_,
    new_n8638_, new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_,
    new_n8644_, new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_,
    new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_,
    new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_,
    new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_,
    new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_,
    new_n8674_, new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_,
    new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_,
    new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_,
    new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_,
    new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_,
    new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_,
    new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_,
    new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_,
    new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_,
    new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_,
    new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_,
    new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_,
    new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_,
    new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_,
    new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_,
    new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_,
    new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_,
    new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_,
    new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_,
    new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_,
    new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_,
    new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_,
    new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_,
    new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_,
    new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_,
    new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_,
    new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_,
    new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_,
    new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_,
    new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_,
    new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_,
    new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_,
    new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_,
    new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_,
    new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_,
    new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_,
    new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_,
    new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_,
    new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_,
    new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_,
    new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_,
    new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_,
    new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_,
    new_n8933_, new_n8934_, new_n8935_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_,
    new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_,
    new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_,
    new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_,
    new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_,
    new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_,
    new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_,
    new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_,
    new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_,
    new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_,
    new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9120_,
    new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_,
    new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_,
    new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_,
    new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_,
    new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_,
    new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_,
    new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_,
    new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_,
    new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_,
    new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_,
    new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_,
    new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_,
    new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_,
    new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_,
    new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_,
    new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_,
    new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_,
    new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9300_, new_n9301_,
    new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_,
    new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_,
    new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_,
    new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_,
    new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_,
    new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_,
    new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_,
    new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_,
    new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_,
    new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_,
    new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_,
    new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_,
    new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_,
    new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_,
    new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_,
    new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_,
    new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_,
    new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_,
    new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_,
    new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_,
    new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_,
    new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_,
    new_n9464_, new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_,
    new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_,
    new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_,
    new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_,
    new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_,
    new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_,
    new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_,
    new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_,
    new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_,
    new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_,
    new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_,
    new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_,
    new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_,
    new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_,
    new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_,
    new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_,
    new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_,
    new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_,
    new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_,
    new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_,
    new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_,
    new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_,
    new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_,
    new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_,
    new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_,
    new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_,
    new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_,
    new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_,
    new_n9633_, new_n9634_, new_n9635_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_,
    new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_,
    new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_,
    new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_,
    new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_,
    new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_,
    new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_,
    new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9814_,
    new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_,
    new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_,
    new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_,
    new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_,
    new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_,
    new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_,
    new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_,
    new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_,
    new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_,
    new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_,
    new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_,
    new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_,
    new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_,
    new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_,
    new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_,
    new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_,
    new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_,
    new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_,
    new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_,
    new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_,
    new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_,
    new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_,
    new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_,
    new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_,
    new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_,
    new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_,
    new_n9977_, new_n9978_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10147_, new_n10148_, new_n10149_, new_n10150_, new_n10151_,
    new_n10152_, new_n10153_, new_n10154_, new_n10155_, new_n10156_,
    new_n10157_, new_n10158_, new_n10159_, new_n10160_, new_n10161_,
    new_n10162_, new_n10163_, new_n10164_, new_n10165_, new_n10166_,
    new_n10167_, new_n10168_, new_n10169_, new_n10170_, new_n10171_,
    new_n10172_, new_n10173_, new_n10174_, new_n10175_, new_n10176_,
    new_n10177_, new_n10178_, new_n10179_, new_n10180_, new_n10181_,
    new_n10182_, new_n10183_, new_n10184_, new_n10185_, new_n10186_,
    new_n10187_, new_n10188_, new_n10189_, new_n10190_, new_n10191_,
    new_n10192_, new_n10193_, new_n10194_, new_n10195_, new_n10196_,
    new_n10197_, new_n10198_, new_n10199_, new_n10200_, new_n10201_,
    new_n10202_, new_n10203_, new_n10204_, new_n10205_, new_n10206_,
    new_n10207_, new_n10208_, new_n10209_, new_n10210_, new_n10211_,
    new_n10212_, new_n10213_, new_n10214_, new_n10215_, new_n10216_,
    new_n10217_, new_n10218_, new_n10219_, new_n10220_, new_n10221_,
    new_n10222_, new_n10223_, new_n10224_, new_n10225_, new_n10226_,
    new_n10227_, new_n10228_, new_n10229_, new_n10230_, new_n10231_,
    new_n10232_, new_n10233_, new_n10234_, new_n10235_, new_n10236_,
    new_n10237_, new_n10238_, new_n10239_, new_n10240_, new_n10241_,
    new_n10242_, new_n10243_, new_n10244_, new_n10245_, new_n10246_,
    new_n10247_, new_n10248_, new_n10249_, new_n10250_, new_n10251_,
    new_n10252_, new_n10253_, new_n10254_, new_n10255_, new_n10256_,
    new_n10257_, new_n10258_, new_n10259_, new_n10260_, new_n10261_,
    new_n10262_, new_n10263_, new_n10264_, new_n10265_, new_n10266_,
    new_n10267_, new_n10268_, new_n10269_, new_n10270_, new_n10271_,
    new_n10272_, new_n10273_, new_n10274_, new_n10275_, new_n10276_,
    new_n10277_, new_n10278_, new_n10279_, new_n10280_, new_n10281_,
    new_n10282_, new_n10283_, new_n10284_, new_n10285_, new_n10286_,
    new_n10287_, new_n10288_, new_n10289_, new_n10290_, new_n10291_,
    new_n10292_, new_n10293_, new_n10294_, new_n10295_, new_n10296_,
    new_n10297_, new_n10298_, new_n10299_, new_n10300_, new_n10301_,
    new_n10302_, new_n10303_, new_n10304_, new_n10305_, new_n10306_,
    new_n10307_, new_n10308_, new_n10309_, new_n10310_, new_n10312_,
    new_n10313_, new_n10314_, new_n10315_, new_n10316_, new_n10317_,
    new_n10318_, new_n10319_, new_n10320_, new_n10321_, new_n10322_,
    new_n10323_, new_n10324_, new_n10325_, new_n10326_, new_n10327_,
    new_n10328_, new_n10329_, new_n10330_, new_n10331_, new_n10332_,
    new_n10333_, new_n10334_, new_n10335_, new_n10336_, new_n10337_,
    new_n10338_, new_n10339_, new_n10340_, new_n10341_, new_n10342_,
    new_n10343_, new_n10344_, new_n10345_, new_n10346_, new_n10347_,
    new_n10348_, new_n10349_, new_n10350_, new_n10351_, new_n10352_,
    new_n10353_, new_n10354_, new_n10355_, new_n10356_, new_n10357_,
    new_n10358_, new_n10359_, new_n10360_, new_n10361_, new_n10362_,
    new_n10363_, new_n10364_, new_n10365_, new_n10366_, new_n10367_,
    new_n10368_, new_n10369_, new_n10370_, new_n10371_, new_n10372_,
    new_n10373_, new_n10374_, new_n10375_, new_n10376_, new_n10377_,
    new_n10378_, new_n10379_, new_n10380_, new_n10381_, new_n10382_,
    new_n10383_, new_n10384_, new_n10385_, new_n10386_, new_n10387_,
    new_n10388_, new_n10389_, new_n10390_, new_n10391_, new_n10392_,
    new_n10393_, new_n10394_, new_n10395_, new_n10396_, new_n10397_,
    new_n10398_, new_n10399_, new_n10400_, new_n10401_, new_n10402_,
    new_n10403_, new_n10404_, new_n10405_, new_n10406_, new_n10407_,
    new_n10408_, new_n10409_, new_n10410_, new_n10411_, new_n10412_,
    new_n10413_, new_n10414_, new_n10415_, new_n10416_, new_n10417_,
    new_n10418_, new_n10419_, new_n10420_, new_n10421_, new_n10422_,
    new_n10423_, new_n10424_, new_n10425_, new_n10426_, new_n10427_,
    new_n10428_, new_n10429_, new_n10430_, new_n10431_, new_n10432_,
    new_n10433_, new_n10434_, new_n10435_, new_n10436_, new_n10437_,
    new_n10438_, new_n10439_, new_n10440_, new_n10441_, new_n10442_,
    new_n10443_, new_n10444_, new_n10445_, new_n10446_, new_n10447_,
    new_n10448_, new_n10449_, new_n10450_, new_n10451_, new_n10452_,
    new_n10453_, new_n10454_, new_n10455_, new_n10456_, new_n10457_,
    new_n10458_, new_n10459_, new_n10460_, new_n10461_, new_n10462_,
    new_n10463_, new_n10464_, new_n10465_, new_n10466_, new_n10467_,
    new_n10468_, new_n10469_, new_n10470_, new_n10471_, new_n10472_,
    new_n10473_, new_n10474_, new_n10475_, new_n10476_, new_n10477_,
    new_n10478_, new_n10479_, new_n10480_, new_n10481_, new_n10482_,
    new_n10483_, new_n10484_, new_n10485_, new_n10486_, new_n10487_,
    new_n10488_, new_n10489_, new_n10491_, new_n10492_, new_n10493_,
    new_n10494_, new_n10495_, new_n10496_, new_n10497_, new_n10498_,
    new_n10499_, new_n10500_, new_n10501_, new_n10502_, new_n10503_,
    new_n10504_, new_n10505_, new_n10506_, new_n10507_, new_n10508_,
    new_n10509_, new_n10510_, new_n10511_, new_n10512_, new_n10513_,
    new_n10514_, new_n10515_, new_n10516_, new_n10517_, new_n10518_,
    new_n10519_, new_n10520_, new_n10521_, new_n10522_, new_n10523_,
    new_n10524_, new_n10525_, new_n10526_, new_n10527_, new_n10528_,
    new_n10529_, new_n10530_, new_n10531_, new_n10532_, new_n10533_,
    new_n10534_, new_n10535_, new_n10536_, new_n10537_, new_n10538_,
    new_n10539_, new_n10540_, new_n10541_, new_n10542_, new_n10543_,
    new_n10544_, new_n10545_, new_n10546_, new_n10547_, new_n10548_,
    new_n10549_, new_n10550_, new_n10551_, new_n10552_, new_n10553_,
    new_n10554_, new_n10555_, new_n10556_, new_n10557_, new_n10558_,
    new_n10559_, new_n10560_, new_n10561_, new_n10562_, new_n10563_,
    new_n10564_, new_n10565_, new_n10566_, new_n10567_, new_n10568_,
    new_n10569_, new_n10570_, new_n10571_, new_n10572_, new_n10573_,
    new_n10574_, new_n10575_, new_n10576_, new_n10577_, new_n10578_,
    new_n10579_, new_n10580_, new_n10581_, new_n10582_, new_n10583_,
    new_n10584_, new_n10585_, new_n10586_, new_n10587_, new_n10588_,
    new_n10589_, new_n10590_, new_n10591_, new_n10592_, new_n10593_,
    new_n10594_, new_n10595_, new_n10596_, new_n10597_, new_n10598_,
    new_n10599_, new_n10600_, new_n10601_, new_n10602_, new_n10603_,
    new_n10604_, new_n10605_, new_n10606_, new_n10607_, new_n10608_,
    new_n10609_, new_n10610_, new_n10611_, new_n10612_, new_n10613_,
    new_n10614_, new_n10615_, new_n10616_, new_n10617_, new_n10618_,
    new_n10619_, new_n10620_, new_n10621_, new_n10622_, new_n10623_,
    new_n10624_, new_n10625_, new_n10626_, new_n10627_, new_n10628_,
    new_n10629_, new_n10630_, new_n10631_, new_n10632_, new_n10633_,
    new_n10634_, new_n10635_, new_n10636_, new_n10637_, new_n10638_,
    new_n10639_, new_n10640_, new_n10641_, new_n10642_, new_n10643_,
    new_n10644_, new_n10645_, new_n10646_, new_n10647_, new_n10648_,
    new_n10649_, new_n10650_, new_n10651_, new_n10652_, new_n10653_,
    new_n10654_, new_n10655_, new_n10656_, new_n10657_, new_n10658_,
    new_n10659_, new_n10660_, new_n10661_, new_n10662_, new_n10663_,
    new_n10664_, new_n10665_, new_n10666_, new_n10667_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11025_, new_n11026_,
    new_n11027_, new_n11028_, new_n11029_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11094_, new_n11095_, new_n11096_, new_n11097_,
    new_n11098_, new_n11099_, new_n11100_, new_n11101_, new_n11102_,
    new_n11103_, new_n11104_, new_n11105_, new_n11106_, new_n11107_,
    new_n11108_, new_n11109_, new_n11110_, new_n11111_, new_n11112_,
    new_n11113_, new_n11114_, new_n11115_, new_n11116_, new_n11117_,
    new_n11118_, new_n11119_, new_n11120_, new_n11121_, new_n11122_,
    new_n11123_, new_n11124_, new_n11125_, new_n11126_, new_n11127_,
    new_n11128_, new_n11129_, new_n11130_, new_n11131_, new_n11132_,
    new_n11133_, new_n11134_, new_n11135_, new_n11136_, new_n11137_,
    new_n11138_, new_n11139_, new_n11140_, new_n11141_, new_n11142_,
    new_n11143_, new_n11144_, new_n11145_, new_n11146_, new_n11147_,
    new_n11148_, new_n11149_, new_n11150_, new_n11151_, new_n11152_,
    new_n11153_, new_n11154_, new_n11155_, new_n11156_, new_n11157_,
    new_n11158_, new_n11159_, new_n11160_, new_n11161_, new_n11162_,
    new_n11163_, new_n11164_, new_n11165_, new_n11166_, new_n11167_,
    new_n11168_, new_n11169_, new_n11170_, new_n11171_, new_n11172_,
    new_n11173_, new_n11174_, new_n11175_, new_n11176_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11188_, new_n11189_, new_n11190_, new_n11191_, new_n11192_,
    new_n11193_, new_n11194_, new_n11195_, new_n11196_, new_n11197_,
    new_n11198_, new_n11199_, new_n11200_, new_n11201_, new_n11202_,
    new_n11203_, new_n11204_, new_n11205_, new_n11206_, new_n11207_,
    new_n11208_, new_n11209_, new_n11210_, new_n11211_, new_n11212_,
    new_n11213_, new_n11214_, new_n11215_, new_n11216_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11227_,
    new_n11228_, new_n11229_, new_n11230_, new_n11231_, new_n11232_,
    new_n11233_, new_n11234_, new_n11235_, new_n11237_, new_n11238_,
    new_n11239_, new_n11240_, new_n11241_, new_n11242_, new_n11243_,
    new_n11244_, new_n11245_, new_n11246_, new_n11247_, new_n11248_,
    new_n11249_, new_n11250_, new_n11251_, new_n11252_, new_n11253_,
    new_n11254_, new_n11255_, new_n11256_, new_n11257_, new_n11258_,
    new_n11259_, new_n11260_, new_n11261_, new_n11262_, new_n11263_,
    new_n11264_, new_n11265_, new_n11266_, new_n11267_, new_n11268_,
    new_n11269_, new_n11270_, new_n11271_, new_n11272_, new_n11273_,
    new_n11274_, new_n11275_, new_n11276_, new_n11277_, new_n11278_,
    new_n11279_, new_n11280_, new_n11281_, new_n11282_, new_n11283_,
    new_n11284_, new_n11285_, new_n11286_, new_n11287_, new_n11288_,
    new_n11289_, new_n11290_, new_n11291_, new_n11292_, new_n11293_,
    new_n11294_, new_n11295_, new_n11296_, new_n11297_, new_n11298_,
    new_n11299_, new_n11300_, new_n11301_, new_n11302_, new_n11303_,
    new_n11304_, new_n11305_, new_n11306_, new_n11307_, new_n11308_,
    new_n11309_, new_n11310_, new_n11311_, new_n11312_, new_n11313_,
    new_n11314_, new_n11315_, new_n11316_, new_n11317_, new_n11318_,
    new_n11319_, new_n11320_, new_n11321_, new_n11322_, new_n11323_,
    new_n11324_, new_n11325_, new_n11326_, new_n11327_, new_n11328_,
    new_n11329_, new_n11330_, new_n11331_, new_n11332_, new_n11333_,
    new_n11334_, new_n11335_, new_n11336_, new_n11337_, new_n11338_,
    new_n11339_, new_n11340_, new_n11341_, new_n11342_, new_n11343_,
    new_n11344_, new_n11345_, new_n11346_, new_n11347_, new_n11348_,
    new_n11349_, new_n11350_, new_n11351_, new_n11352_, new_n11353_,
    new_n11354_, new_n11355_, new_n11356_, new_n11357_, new_n11358_,
    new_n11359_, new_n11360_, new_n11361_, new_n11362_, new_n11363_,
    new_n11364_, new_n11365_, new_n11366_, new_n11367_, new_n11368_,
    new_n11369_, new_n11370_, new_n11371_, new_n11372_, new_n11373_,
    new_n11374_, new_n11375_, new_n11376_, new_n11377_, new_n11378_,
    new_n11379_, new_n11380_, new_n11381_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11528_, new_n11529_,
    new_n11530_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11790_, new_n11791_,
    new_n11792_, new_n11793_, new_n11794_, new_n11795_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11813_, new_n11814_, new_n11815_, new_n11816_, new_n11817_,
    new_n11818_, new_n11819_, new_n11820_, new_n11821_, new_n11822_,
    new_n11823_, new_n11824_, new_n11825_, new_n11826_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11844_, new_n11845_, new_n11846_, new_n11847_,
    new_n11848_, new_n11849_, new_n11850_, new_n11851_, new_n11852_,
    new_n11853_, new_n11854_, new_n11855_, new_n11856_, new_n11857_,
    new_n11858_, new_n11859_, new_n11860_, new_n11861_, new_n11862_,
    new_n11863_, new_n11864_, new_n11865_, new_n11866_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11873_, new_n11874_, new_n11875_, new_n11876_, new_n11877_,
    new_n11878_, new_n11879_, new_n11880_, new_n11881_, new_n11882_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11926_, new_n11927_, new_n11928_,
    new_n11929_, new_n11930_, new_n11931_, new_n11932_, new_n11933_,
    new_n11934_, new_n11935_, new_n11936_, new_n11937_, new_n11938_,
    new_n11939_, new_n11940_, new_n11941_, new_n11942_, new_n11943_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11950_, new_n11951_, new_n11952_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11958_,
    new_n11959_, new_n11960_, new_n11961_, new_n11962_, new_n11963_,
    new_n11964_, new_n11965_, new_n11966_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12061_, new_n12062_, new_n12063_, new_n12064_,
    new_n12065_, new_n12066_, new_n12067_, new_n12068_, new_n12069_,
    new_n12070_, new_n12071_, new_n12072_, new_n12073_, new_n12074_,
    new_n12075_, new_n12076_, new_n12077_, new_n12078_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12084_,
    new_n12085_, new_n12086_, new_n12087_, new_n12088_, new_n12089_,
    new_n12090_, new_n12091_, new_n12092_, new_n12093_, new_n12094_,
    new_n12095_, new_n12096_, new_n12097_, new_n12098_, new_n12099_,
    new_n12100_, new_n12101_, new_n12102_, new_n12103_, new_n12104_,
    new_n12105_, new_n12106_, new_n12107_, new_n12108_, new_n12109_,
    new_n12110_, new_n12111_, new_n12112_, new_n12113_, new_n12114_,
    new_n12115_, new_n12116_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12302_, new_n12303_, new_n12304_, new_n12305_, new_n12306_,
    new_n12307_, new_n12308_, new_n12309_, new_n12310_, new_n12311_,
    new_n12312_, new_n12313_, new_n12314_, new_n12315_, new_n12316_,
    new_n12317_, new_n12318_, new_n12319_, new_n12320_, new_n12321_,
    new_n12322_, new_n12323_, new_n12324_, new_n12325_, new_n12326_,
    new_n12327_, new_n12328_, new_n12329_, new_n12330_, new_n12331_,
    new_n12332_, new_n12333_, new_n12334_, new_n12335_, new_n12336_,
    new_n12337_, new_n12338_, new_n12339_, new_n12340_, new_n12341_,
    new_n12342_, new_n12343_, new_n12344_, new_n12345_, new_n12346_,
    new_n12347_, new_n12348_, new_n12349_, new_n12350_, new_n12351_,
    new_n12352_, new_n12353_, new_n12354_, new_n12355_, new_n12356_,
    new_n12357_, new_n12358_, new_n12359_, new_n12360_, new_n12361_,
    new_n12362_, new_n12363_, new_n12364_, new_n12365_, new_n12366_,
    new_n12367_, new_n12368_, new_n12369_, new_n12370_, new_n12371_,
    new_n12372_, new_n12373_, new_n12374_, new_n12375_, new_n12376_,
    new_n12377_, new_n12378_, new_n12379_, new_n12380_, new_n12381_,
    new_n12382_, new_n12383_, new_n12384_, new_n12385_, new_n12386_,
    new_n12387_, new_n12388_, new_n12389_, new_n12390_, new_n12391_,
    new_n12392_, new_n12393_, new_n12394_, new_n12395_, new_n12396_,
    new_n12397_, new_n12398_, new_n12399_, new_n12400_, new_n12401_,
    new_n12402_, new_n12403_, new_n12404_, new_n12405_, new_n12406_,
    new_n12407_, new_n12408_, new_n12409_, new_n12410_, new_n12411_,
    new_n12412_, new_n12413_, new_n12414_, new_n12415_, new_n12416_,
    new_n12418_, new_n12419_, new_n12420_, new_n12421_, new_n12422_,
    new_n12423_, new_n12424_, new_n12425_, new_n12426_, new_n12427_,
    new_n12428_, new_n12429_, new_n12430_, new_n12431_, new_n12432_,
    new_n12433_, new_n12434_, new_n12435_, new_n12436_, new_n12437_,
    new_n12438_, new_n12439_, new_n12440_, new_n12441_, new_n12442_,
    new_n12443_, new_n12444_, new_n12445_, new_n12446_, new_n12447_,
    new_n12448_, new_n12449_, new_n12450_, new_n12451_, new_n12452_,
    new_n12453_, new_n12454_, new_n12455_, new_n12456_, new_n12457_,
    new_n12458_, new_n12459_, new_n12460_, new_n12461_, new_n12462_,
    new_n12463_, new_n12464_, new_n12465_, new_n12466_, new_n12467_,
    new_n12468_, new_n12469_, new_n12470_, new_n12471_, new_n12472_,
    new_n12473_, new_n12474_, new_n12475_, new_n12476_, new_n12477_,
    new_n12478_, new_n12479_, new_n12480_, new_n12481_, new_n12482_,
    new_n12483_, new_n12484_, new_n12485_, new_n12486_, new_n12487_,
    new_n12488_, new_n12489_, new_n12490_, new_n12491_, new_n12492_,
    new_n12493_, new_n12494_, new_n12495_, new_n12496_, new_n12497_,
    new_n12498_, new_n12499_, new_n12500_, new_n12501_, new_n12502_,
    new_n12503_, new_n12504_, new_n12505_, new_n12506_, new_n12507_,
    new_n12508_, new_n12509_, new_n12510_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12522_,
    new_n12523_, new_n12524_, new_n12525_, new_n12526_, new_n12527_,
    new_n12528_, new_n12529_, new_n12530_, new_n12531_, new_n12532_,
    new_n12533_, new_n12534_, new_n12535_, new_n12537_, new_n12538_,
    new_n12539_, new_n12540_, new_n12541_, new_n12542_, new_n12543_,
    new_n12544_, new_n12545_, new_n12546_, new_n12547_, new_n12548_,
    new_n12549_, new_n12550_, new_n12551_, new_n12552_, new_n12553_,
    new_n12554_, new_n12555_, new_n12556_, new_n12557_, new_n12558_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12566_, new_n12567_, new_n12568_,
    new_n12569_, new_n12570_, new_n12571_, new_n12572_, new_n12573_,
    new_n12574_, new_n12575_, new_n12576_, new_n12577_, new_n12578_,
    new_n12579_, new_n12580_, new_n12581_, new_n12582_, new_n12583_,
    new_n12584_, new_n12585_, new_n12586_, new_n12587_, new_n12588_,
    new_n12589_, new_n12590_, new_n12591_, new_n12592_, new_n12593_,
    new_n12594_, new_n12595_, new_n12596_, new_n12597_, new_n12598_,
    new_n12599_, new_n12600_, new_n12601_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12608_,
    new_n12609_, new_n12610_, new_n12611_, new_n12612_, new_n12613_,
    new_n12614_, new_n12615_, new_n12616_, new_n12617_, new_n12618_,
    new_n12619_, new_n12620_, new_n12621_, new_n12622_, new_n12623_,
    new_n12624_, new_n12625_, new_n12626_, new_n12627_, new_n12628_,
    new_n12629_, new_n12630_, new_n12631_, new_n12632_, new_n12633_,
    new_n12634_, new_n12635_, new_n12636_, new_n12637_, new_n12638_,
    new_n12640_, new_n12641_, new_n12642_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12649_,
    new_n12650_, new_n12651_, new_n12652_, new_n12653_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12663_, new_n12664_,
    new_n12665_, new_n12666_, new_n12667_, new_n12668_, new_n12669_,
    new_n12670_, new_n12671_, new_n12672_, new_n12673_, new_n12674_,
    new_n12675_, new_n12676_, new_n12677_, new_n12678_, new_n12679_,
    new_n12680_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12687_, new_n12688_, new_n12689_,
    new_n12690_, new_n12691_, new_n12692_, new_n12693_, new_n12694_,
    new_n12695_, new_n12696_, new_n12697_, new_n12698_, new_n12699_,
    new_n12700_, new_n12701_, new_n12702_, new_n12703_, new_n12704_,
    new_n12705_, new_n12706_, new_n12707_, new_n12708_, new_n12709_,
    new_n12710_, new_n12711_, new_n12712_, new_n12713_, new_n12714_,
    new_n12715_, new_n12716_, new_n12717_, new_n12718_, new_n12719_,
    new_n12720_, new_n12721_, new_n12722_, new_n12723_, new_n12724_,
    new_n12725_, new_n12726_, new_n12727_, new_n12728_, new_n12729_,
    new_n12730_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12852_, new_n12853_, new_n12854_, new_n12855_, new_n12856_,
    new_n12857_, new_n12858_, new_n12859_, new_n12860_, new_n12861_,
    new_n12862_, new_n12863_, new_n12864_, new_n12865_, new_n12866_,
    new_n12867_, new_n12868_, new_n12869_, new_n12870_, new_n12871_,
    new_n12872_, new_n12873_, new_n12874_, new_n12875_, new_n12876_,
    new_n12877_, new_n12878_, new_n12879_, new_n12880_, new_n12881_,
    new_n12882_, new_n12883_, new_n12884_, new_n12885_, new_n12886_,
    new_n12887_, new_n12888_, new_n12889_, new_n12890_, new_n12891_,
    new_n12892_, new_n12893_, new_n12894_, new_n12895_, new_n12896_,
    new_n12897_, new_n12898_, new_n12899_, new_n12900_, new_n12901_,
    new_n12902_, new_n12903_, new_n12904_, new_n12905_, new_n12906_,
    new_n12907_, new_n12908_, new_n12909_, new_n12910_, new_n12911_,
    new_n12912_, new_n12913_, new_n12914_, new_n12915_, new_n12916_,
    new_n12917_, new_n12918_, new_n12919_, new_n12920_, new_n12921_,
    new_n12922_, new_n12923_, new_n12924_, new_n12925_, new_n12926_,
    new_n12927_, new_n12928_, new_n12929_, new_n12930_, new_n12931_,
    new_n12932_, new_n12933_, new_n12934_, new_n12935_, new_n12936_,
    new_n12937_, new_n12938_, new_n12939_, new_n12940_, new_n12941_,
    new_n12942_, new_n12943_, new_n12944_, new_n12945_, new_n12946_,
    new_n12947_, new_n12948_, new_n12949_, new_n12950_, new_n12951_,
    new_n12952_, new_n12953_, new_n12954_, new_n12955_, new_n12956_,
    new_n12957_, new_n12958_, new_n12959_, new_n12960_, new_n12961_,
    new_n12962_, new_n12964_, new_n12965_, new_n12966_, new_n12967_,
    new_n12968_, new_n12969_, new_n12970_, new_n12971_, new_n12972_,
    new_n12973_, new_n12974_, new_n12975_, new_n12976_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12983_, new_n12984_, new_n12985_, new_n12986_, new_n12987_,
    new_n12988_, new_n12989_, new_n12990_, new_n12991_, new_n12992_,
    new_n12993_, new_n12994_, new_n12995_, new_n12996_, new_n12997_,
    new_n12998_, new_n12999_, new_n13000_, new_n13001_, new_n13002_,
    new_n13003_, new_n13004_, new_n13005_, new_n13006_, new_n13007_,
    new_n13008_, new_n13009_, new_n13010_, new_n13011_, new_n13012_,
    new_n13013_, new_n13014_, new_n13015_, new_n13016_, new_n13017_,
    new_n13018_, new_n13019_, new_n13020_, new_n13021_, new_n13022_,
    new_n13023_, new_n13024_, new_n13025_, new_n13026_, new_n13027_,
    new_n13028_, new_n13029_, new_n13030_, new_n13031_, new_n13032_,
    new_n13033_, new_n13034_, new_n13035_, new_n13036_, new_n13037_,
    new_n13038_, new_n13039_, new_n13040_, new_n13041_, new_n13042_,
    new_n13043_, new_n13044_, new_n13045_, new_n13046_, new_n13047_,
    new_n13048_, new_n13049_, new_n13050_, new_n13051_, new_n13052_,
    new_n13053_, new_n13054_, new_n13055_, new_n13056_, new_n13057_,
    new_n13058_, new_n13059_, new_n13060_, new_n13061_, new_n13062_,
    new_n13063_, new_n13065_, new_n13066_, new_n13067_, new_n13068_,
    new_n13069_, new_n13070_, new_n13071_, new_n13072_, new_n13073_,
    new_n13074_, new_n13075_, new_n13076_, new_n13077_, new_n13078_,
    new_n13079_, new_n13080_, new_n13081_, new_n13082_, new_n13083_,
    new_n13084_, new_n13085_, new_n13086_, new_n13087_, new_n13088_,
    new_n13089_, new_n13090_, new_n13091_, new_n13092_, new_n13093_,
    new_n13094_, new_n13095_, new_n13096_, new_n13097_, new_n13098_,
    new_n13099_, new_n13100_, new_n13101_, new_n13102_, new_n13103_,
    new_n13104_, new_n13105_, new_n13106_, new_n13107_, new_n13108_,
    new_n13109_, new_n13110_, new_n13111_, new_n13112_, new_n13113_,
    new_n13114_, new_n13115_, new_n13116_, new_n13117_, new_n13118_,
    new_n13119_, new_n13120_, new_n13121_, new_n13122_, new_n13123_,
    new_n13124_, new_n13125_, new_n13126_, new_n13127_, new_n13128_,
    new_n13129_, new_n13130_, new_n13131_, new_n13132_, new_n13133_,
    new_n13134_, new_n13135_, new_n13136_, new_n13137_, new_n13138_,
    new_n13139_, new_n13140_, new_n13141_, new_n13142_, new_n13143_,
    new_n13144_, new_n13145_, new_n13146_, new_n13147_, new_n13148_,
    new_n13149_, new_n13150_, new_n13151_, new_n13152_, new_n13153_,
    new_n13154_, new_n13155_, new_n13156_, new_n13157_, new_n13158_,
    new_n13159_, new_n13160_, new_n13161_, new_n13162_, new_n13163_,
    new_n13164_, new_n13165_, new_n13166_, new_n13167_, new_n13169_,
    new_n13170_, new_n13171_, new_n13172_, new_n13173_, new_n13174_,
    new_n13175_, new_n13176_, new_n13177_, new_n13178_, new_n13179_,
    new_n13180_, new_n13181_, new_n13182_, new_n13183_, new_n13184_,
    new_n13185_, new_n13186_, new_n13187_, new_n13188_, new_n13189_,
    new_n13190_, new_n13191_, new_n13192_, new_n13193_, new_n13194_,
    new_n13195_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13200_, new_n13201_, new_n13202_, new_n13203_, new_n13204_,
    new_n13205_, new_n13206_, new_n13207_, new_n13208_, new_n13209_,
    new_n13210_, new_n13211_, new_n13212_, new_n13213_, new_n13214_,
    new_n13215_, new_n13216_, new_n13217_, new_n13218_, new_n13219_,
    new_n13220_, new_n13221_, new_n13222_, new_n13223_, new_n13224_,
    new_n13225_, new_n13226_, new_n13227_, new_n13228_, new_n13229_,
    new_n13230_, new_n13231_, new_n13232_, new_n13233_, new_n13234_,
    new_n13235_, new_n13236_, new_n13237_, new_n13238_, new_n13239_,
    new_n13240_, new_n13241_, new_n13242_, new_n13243_, new_n13244_,
    new_n13245_, new_n13246_, new_n13247_, new_n13248_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13344_, new_n13345_, new_n13346_,
    new_n13347_, new_n13348_, new_n13349_, new_n13350_, new_n13351_,
    new_n13352_, new_n13353_, new_n13354_, new_n13355_, new_n13356_,
    new_n13357_, new_n13358_, new_n13359_, new_n13360_, new_n13361_,
    new_n13362_, new_n13363_, new_n13364_, new_n13365_, new_n13366_,
    new_n13367_, new_n13368_, new_n13369_, new_n13370_, new_n13371_,
    new_n13372_, new_n13373_, new_n13374_, new_n13375_, new_n13376_,
    new_n13377_, new_n13378_, new_n13379_, new_n13380_, new_n13381_,
    new_n13382_, new_n13383_, new_n13384_, new_n13385_, new_n13386_,
    new_n13387_, new_n13388_, new_n13389_, new_n13390_, new_n13391_,
    new_n13392_, new_n13393_, new_n13394_, new_n13395_, new_n13396_,
    new_n13397_, new_n13398_, new_n13399_, new_n13400_, new_n13401_,
    new_n13402_, new_n13403_, new_n13404_, new_n13405_, new_n13406_,
    new_n13407_, new_n13408_, new_n13409_, new_n13410_, new_n13411_,
    new_n13412_, new_n13413_, new_n13414_, new_n13415_, new_n13416_,
    new_n13417_, new_n13418_, new_n13419_, new_n13421_, new_n13422_,
    new_n13423_, new_n13424_, new_n13425_, new_n13426_, new_n13427_,
    new_n13428_, new_n13429_, new_n13430_, new_n13431_, new_n13432_,
    new_n13433_, new_n13434_, new_n13435_, new_n13436_, new_n13437_,
    new_n13438_, new_n13439_, new_n13440_, new_n13441_, new_n13442_,
    new_n13443_, new_n13444_, new_n13445_, new_n13446_, new_n13447_,
    new_n13448_, new_n13449_, new_n13450_, new_n13451_, new_n13452_,
    new_n13453_, new_n13454_, new_n13455_, new_n13456_, new_n13457_,
    new_n13458_, new_n13459_, new_n13460_, new_n13461_, new_n13462_,
    new_n13463_, new_n13464_, new_n13465_, new_n13466_, new_n13467_,
    new_n13468_, new_n13469_, new_n13470_, new_n13471_, new_n13472_,
    new_n13473_, new_n13474_, new_n13475_, new_n13476_, new_n13477_,
    new_n13478_, new_n13479_, new_n13480_, new_n13481_, new_n13482_,
    new_n13483_, new_n13484_, new_n13485_, new_n13486_, new_n13487_,
    new_n13488_, new_n13489_, new_n13490_, new_n13491_, new_n13492_,
    new_n13493_, new_n13494_, new_n13495_, new_n13496_, new_n13497_,
    new_n13498_, new_n13500_, new_n13501_, new_n13502_, new_n13503_,
    new_n13504_, new_n13505_, new_n13506_, new_n13507_, new_n13508_,
    new_n13509_, new_n13510_, new_n13511_, new_n13512_, new_n13513_,
    new_n13514_, new_n13515_, new_n13516_, new_n13517_, new_n13518_,
    new_n13519_, new_n13520_, new_n13521_, new_n13522_, new_n13523_,
    new_n13524_, new_n13525_, new_n13526_, new_n13527_, new_n13528_,
    new_n13529_, new_n13530_, new_n13531_, new_n13532_, new_n13533_,
    new_n13534_, new_n13535_, new_n13536_, new_n13537_, new_n13538_,
    new_n13539_, new_n13540_, new_n13541_, new_n13542_, new_n13543_,
    new_n13544_, new_n13545_, new_n13546_, new_n13547_, new_n13548_,
    new_n13549_, new_n13550_, new_n13551_, new_n13552_, new_n13553_,
    new_n13554_, new_n13555_, new_n13556_, new_n13557_, new_n13558_,
    new_n13559_, new_n13560_, new_n13561_, new_n13562_, new_n13563_,
    new_n13564_, new_n13565_, new_n13567_, new_n13568_, new_n13569_,
    new_n13570_, new_n13571_, new_n13572_, new_n13573_, new_n13574_,
    new_n13575_, new_n13576_, new_n13577_, new_n13578_, new_n13579_,
    new_n13580_, new_n13581_, new_n13582_, new_n13583_, new_n13584_,
    new_n13585_, new_n13586_, new_n13587_, new_n13588_, new_n13589_,
    new_n13590_, new_n13591_, new_n13592_, new_n13593_, new_n13594_,
    new_n13595_, new_n13596_, new_n13597_, new_n13598_, new_n13599_,
    new_n13600_, new_n13601_, new_n13602_, new_n13603_, new_n13604_,
    new_n13605_, new_n13606_, new_n13607_, new_n13608_, new_n13609_,
    new_n13610_, new_n13611_, new_n13612_, new_n13613_, new_n13614_,
    new_n13615_, new_n13616_, new_n13617_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13627_, new_n13628_, new_n13629_,
    new_n13630_, new_n13631_, new_n13632_, new_n13633_, new_n13634_,
    new_n13635_, new_n13636_, new_n13637_, new_n13638_, new_n13639_,
    new_n13640_, new_n13641_, new_n13642_, new_n13643_, new_n13644_,
    new_n13645_, new_n13646_, new_n13647_, new_n13648_, new_n13649_,
    new_n13650_, new_n13651_, new_n13652_, new_n13653_, new_n13654_,
    new_n13655_, new_n13656_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13786_, new_n13787_,
    new_n13788_, new_n13789_, new_n13790_, new_n13791_, new_n13792_,
    new_n13793_, new_n13794_, new_n13795_, new_n13796_, new_n13797_,
    new_n13798_, new_n13799_, new_n13800_, new_n13801_, new_n13802_,
    new_n13803_, new_n13804_, new_n13805_, new_n13806_, new_n13807_,
    new_n13808_, new_n13809_, new_n13810_, new_n13811_, new_n13812_,
    new_n13813_, new_n13814_, new_n13815_, new_n13816_, new_n13817_,
    new_n13818_, new_n13819_, new_n13820_, new_n13821_, new_n13822_,
    new_n13823_, new_n13824_, new_n13825_, new_n13826_, new_n13827_,
    new_n13828_, new_n13829_, new_n13830_, new_n13831_, new_n13832_,
    new_n13833_, new_n13834_, new_n13835_, new_n13836_, new_n13837_,
    new_n13838_, new_n13839_, new_n13840_, new_n13841_, new_n13843_,
    new_n13844_, new_n13845_, new_n13846_, new_n13847_, new_n13848_,
    new_n13849_, new_n13850_, new_n13851_, new_n13852_, new_n13853_,
    new_n13854_, new_n13855_, new_n13856_, new_n13857_, new_n13858_,
    new_n13859_, new_n13860_, new_n13861_, new_n13862_, new_n13863_,
    new_n13864_, new_n13865_, new_n13866_, new_n13867_, new_n13868_,
    new_n13869_, new_n13870_, new_n13871_, new_n13872_, new_n13873_,
    new_n13874_, new_n13875_, new_n13876_, new_n13877_, new_n13878_,
    new_n13879_, new_n13880_, new_n13881_, new_n13882_, new_n13883_,
    new_n13884_, new_n13885_, new_n13886_, new_n13887_, new_n13888_,
    new_n13889_, new_n13890_, new_n13891_, new_n13892_, new_n13893_,
    new_n13894_, new_n13895_, new_n13896_, new_n13897_, new_n13898_,
    new_n13899_, new_n13900_, new_n13901_, new_n13902_, new_n13903_,
    new_n13904_, new_n13905_, new_n13906_, new_n13907_, new_n13908_,
    new_n13909_, new_n13910_, new_n13912_, new_n13913_, new_n13914_,
    new_n13915_, new_n13916_, new_n13917_, new_n13918_, new_n13919_,
    new_n13920_, new_n13921_, new_n13922_, new_n13923_, new_n13924_,
    new_n13925_, new_n13926_, new_n13927_, new_n13928_, new_n13929_,
    new_n13930_, new_n13931_, new_n13932_, new_n13933_, new_n13934_,
    new_n13935_, new_n13936_, new_n13937_, new_n13938_, new_n13939_,
    new_n13940_, new_n13941_, new_n13942_, new_n13943_, new_n13944_,
    new_n13945_, new_n13946_, new_n13947_, new_n13948_, new_n13949_,
    new_n13950_, new_n13951_, new_n13952_, new_n13953_, new_n13954_,
    new_n13955_, new_n13956_, new_n13957_, new_n13958_, new_n13959_,
    new_n13960_, new_n13961_, new_n13962_, new_n13963_, new_n13964_,
    new_n13965_, new_n13966_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14123_,
    new_n14124_, new_n14125_, new_n14126_, new_n14127_, new_n14128_,
    new_n14129_, new_n14130_, new_n14131_, new_n14132_, new_n14133_,
    new_n14134_, new_n14135_, new_n14136_, new_n14137_, new_n14138_,
    new_n14139_, new_n14140_, new_n14141_, new_n14142_, new_n14143_,
    new_n14144_, new_n14145_, new_n14146_, new_n14147_, new_n14148_,
    new_n14149_, new_n14150_, new_n14151_, new_n14152_, new_n14153_,
    new_n14154_, new_n14155_, new_n14156_, new_n14157_, new_n14158_,
    new_n14159_, new_n14160_, new_n14161_, new_n14162_, new_n14163_,
    new_n14164_, new_n14165_, new_n14166_, new_n14168_, new_n14169_,
    new_n14170_, new_n14171_, new_n14172_, new_n14173_, new_n14174_,
    new_n14175_, new_n14176_, new_n14177_, new_n14178_, new_n14179_,
    new_n14180_, new_n14181_, new_n14182_, new_n14183_, new_n14184_,
    new_n14185_, new_n14186_, new_n14187_, new_n14188_, new_n14189_,
    new_n14190_, new_n14191_, new_n14192_, new_n14193_, new_n14194_,
    new_n14195_, new_n14196_, new_n14197_, new_n14198_, new_n14199_,
    new_n14200_, new_n14201_, new_n14202_, new_n14203_, new_n14204_,
    new_n14205_, new_n14206_, new_n14207_, new_n14208_, new_n14209_,
    new_n14210_, new_n14212_, new_n14213_, new_n14214_, new_n14215_,
    new_n14216_, new_n14217_, new_n14218_, new_n14219_, new_n14220_,
    new_n14221_, new_n14222_, new_n14223_, new_n14224_, new_n14225_,
    new_n14226_, new_n14227_, new_n14228_, new_n14229_, new_n14230_,
    new_n14231_, new_n14232_, new_n14233_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14240_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14297_, new_n14298_,
    new_n14299_, new_n14300_, new_n14301_, new_n14302_, new_n14303_,
    new_n14304_, new_n14305_, new_n14306_, new_n14307_, new_n14308_,
    new_n14309_, new_n14310_, new_n14311_, new_n14312_, new_n14313_,
    new_n14314_, new_n14315_, new_n14316_, new_n14317_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14324_, new_n14325_, new_n14326_, new_n14327_, new_n14328_,
    new_n14329_, new_n14330_, new_n14331_, new_n14333_, new_n14334_,
    new_n14335_, new_n14336_, new_n14337_, new_n14338_, new_n14339_,
    new_n14340_, new_n14341_, new_n14342_, new_n14343_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14350_,
    new_n14351_, new_n14352_, new_n14353_, new_n14354_, new_n14355_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14367_, new_n14368_, new_n14369_, new_n14370_, new_n14371_,
    new_n14372_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14386_, new_n14387_, new_n14388_,
    new_n14389_, new_n14390_, new_n14391_, new_n14392_, new_n14393_,
    new_n14394_, new_n14395_, new_n14396_, new_n14398_;
  INV_X1     g00000(.I(\a[1] ), .ZN(new_n194_));
  NOR2_X1    g00001(.A1(new_n194_), .A2(\a[0] ), .ZN(\asquared[2] ));
  INV_X1     g00002(.I(\a[0] ), .ZN(new_n196_));
  INV_X1     g00003(.I(\a[2] ), .ZN(new_n197_));
  NOR3_X1    g00004(.A1(new_n196_), .A2(new_n194_), .A3(new_n197_), .ZN(new_n198_));
  OAI21_X1   g00005(.A1(\a[1] ), .A2(\a[2] ), .B(\a[0] ), .ZN(new_n199_));
  NOR2_X1    g00006(.A1(new_n198_), .A2(new_n199_), .ZN(\asquared[3] ));
  NAND2_X1   g00007(.A1(new_n194_), .A2(\a[2] ), .ZN(new_n201_));
  NAND2_X1   g00008(.A1(\a[0] ), .A2(\a[3] ), .ZN(new_n202_));
  XOR2_X1    g00009(.A1(new_n201_), .A2(new_n202_), .Z(new_n203_));
  XOR2_X1    g00010(.A1(new_n203_), .A2(new_n198_), .Z(\asquared[4] ));
  AND3_X2    g00011(.A1(\a[0] ), .A2(\a[2] ), .A3(\a[3] ), .Z(new_n205_));
  INV_X1     g00012(.I(new_n205_), .ZN(new_n206_));
  NAND2_X1   g00013(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n207_));
  AND4_X2    g00014(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[3] ), .A4(\a[4] ), .Z(new_n208_));
  AOI22_X1   g00015(.A1(\a[0] ), .A2(\a[4] ), .B1(\a[1] ), .B2(\a[3] ), .ZN(new_n209_));
  OAI21_X1   g00016(.A1(new_n208_), .A2(new_n209_), .B(new_n207_), .ZN(new_n210_));
  INV_X1     g00017(.I(new_n207_), .ZN(new_n211_));
  NAND4_X1   g00018(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[3] ), .A4(\a[4] ), .ZN(new_n212_));
  INV_X1     g00019(.I(new_n209_), .ZN(new_n213_));
  NAND3_X1   g00020(.A1(new_n213_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n214_));
  NAND2_X1   g00021(.A1(new_n214_), .A2(new_n210_), .ZN(new_n215_));
  XOR2_X1    g00022(.A1(new_n215_), .A2(new_n206_), .Z(\asquared[5] ));
  AOI21_X1   g00023(.A1(new_n213_), .A2(new_n212_), .B(new_n211_), .ZN(new_n217_));
  OAI21_X1   g00024(.A1(new_n206_), .A2(new_n217_), .B(new_n214_), .ZN(new_n218_));
  AOI22_X1   g00025(.A1(\a[0] ), .A2(\a[5] ), .B1(\a[1] ), .B2(\a[4] ), .ZN(new_n219_));
  AND4_X2    g00026(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[4] ), .A4(\a[5] ), .Z(new_n220_));
  NOR3_X1    g00027(.A1(new_n208_), .A2(new_n220_), .A3(new_n219_), .ZN(new_n221_));
  NAND4_X1   g00028(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[4] ), .A4(\a[5] ), .ZN(new_n222_));
  AND4_X2    g00029(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[3] ), .A4(\a[4] ), .Z(new_n223_));
  AOI21_X1   g00030(.A1(new_n223_), .A2(new_n222_), .B(new_n212_), .ZN(new_n224_));
  INV_X1     g00031(.I(\a[3] ), .ZN(new_n225_));
  NOR2_X1    g00032(.A1(new_n225_), .A2(\a[2] ), .ZN(new_n226_));
  NOR3_X1    g00033(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1   g00034(.A1(\a[1] ), .A2(\a[4] ), .ZN(new_n228_));
  NAND2_X1   g00035(.A1(\a[0] ), .A2(\a[5] ), .ZN(new_n229_));
  NAND2_X1   g00036(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1   g00037(.A1(new_n230_), .A2(new_n212_), .A3(new_n222_), .ZN(new_n231_));
  OAI21_X1   g00038(.A1(new_n219_), .A2(new_n220_), .B(new_n208_), .ZN(new_n232_));
  INV_X1     g00039(.I(new_n226_), .ZN(new_n233_));
  AOI21_X1   g00040(.A1(new_n232_), .A2(new_n231_), .B(new_n233_), .ZN(new_n234_));
  NOR2_X1    g00041(.A1(new_n234_), .A2(new_n227_), .ZN(new_n235_));
  XOR2_X1    g00042(.A1(new_n235_), .A2(new_n218_), .Z(\asquared[6] ));
  NOR3_X1    g00043(.A1(new_n208_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n237_));
  AOI21_X1   g00044(.A1(new_n205_), .A2(new_n210_), .B(new_n237_), .ZN(new_n238_));
  NOR2_X1    g00045(.A1(new_n238_), .A2(new_n227_), .ZN(new_n239_));
  NOR2_X1    g00046(.A1(new_n239_), .A2(new_n234_), .ZN(new_n240_));
  NOR2_X1    g00047(.A1(new_n220_), .A2(new_n223_), .ZN(new_n241_));
  NAND2_X1   g00048(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n242_));
  INV_X1     g00049(.I(new_n242_), .ZN(new_n243_));
  AOI22_X1   g00050(.A1(\a[1] ), .A2(\a[5] ), .B1(\a[2] ), .B2(\a[4] ), .ZN(new_n244_));
  AOI21_X1   g00051(.A1(new_n211_), .A2(new_n243_), .B(new_n244_), .ZN(new_n245_));
  NAND2_X1   g00052(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n246_));
  NAND2_X1   g00053(.A1(\a[0] ), .A2(\a[6] ), .ZN(new_n247_));
  AOI22_X1   g00054(.A1(new_n205_), .A2(\a[6] ), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NOR2_X1    g00055(.A1(new_n248_), .A2(new_n245_), .ZN(new_n249_));
  NAND4_X1   g00056(.A1(\a[1] ), .A2(\a[2] ), .A3(\a[4] ), .A4(\a[5] ), .ZN(new_n250_));
  NAND2_X1   g00057(.A1(\a[2] ), .A2(\a[4] ), .ZN(new_n251_));
  INV_X1     g00058(.I(new_n251_), .ZN(new_n252_));
  INV_X1     g00059(.I(\a[5] ), .ZN(new_n253_));
  NOR2_X1    g00060(.A1(new_n194_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1   g00061(.A1(new_n254_), .A2(new_n252_), .B(new_n250_), .ZN(new_n255_));
  INV_X1     g00062(.I(new_n246_), .ZN(new_n256_));
  NAND4_X1   g00063(.A1(\a[0] ), .A2(\a[2] ), .A3(\a[3] ), .A4(\a[6] ), .ZN(new_n257_));
  AND2_X2    g00064(.A1(\a[0] ), .A2(\a[6] ), .Z(new_n258_));
  OAI21_X1   g00065(.A1(new_n256_), .A2(new_n258_), .B(new_n257_), .ZN(new_n259_));
  NOR2_X1    g00066(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  NOR3_X1    g00067(.A1(new_n249_), .A2(new_n260_), .A3(new_n241_), .ZN(new_n261_));
  INV_X1     g00068(.I(new_n261_), .ZN(new_n262_));
  OAI21_X1   g00069(.A1(new_n249_), .A2(new_n260_), .B(new_n241_), .ZN(new_n263_));
  NAND2_X1   g00070(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1     g00071(.I(new_n234_), .ZN(new_n265_));
  NAND3_X1   g00072(.A1(new_n232_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n266_));
  NAND2_X1   g00073(.A1(new_n218_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1     g00074(.I(new_n241_), .ZN(new_n268_));
  NAND2_X1   g00075(.A1(new_n255_), .A2(new_n259_), .ZN(new_n269_));
  NAND2_X1   g00076(.A1(new_n248_), .A2(new_n245_), .ZN(new_n270_));
  AOI21_X1   g00077(.A1(new_n270_), .A2(new_n269_), .B(new_n268_), .ZN(new_n271_));
  AOI21_X1   g00078(.A1(new_n267_), .A2(new_n265_), .B(new_n271_), .ZN(new_n272_));
  AOI22_X1   g00079(.A1(new_n264_), .A2(new_n240_), .B1(new_n272_), .B2(new_n262_), .ZN(\asquared[7] ));
  OAI21_X1   g00080(.A1(new_n239_), .A2(new_n234_), .B(new_n263_), .ZN(new_n274_));
  NAND2_X1   g00081(.A1(new_n274_), .A2(new_n262_), .ZN(new_n275_));
  AOI22_X1   g00082(.A1(\a[2] ), .A2(\a[5] ), .B1(\a[3] ), .B2(\a[4] ), .ZN(new_n276_));
  NAND2_X1   g00083(.A1(\a[0] ), .A2(\a[7] ), .ZN(new_n277_));
  NAND4_X1   g00084(.A1(\a[0] ), .A2(\a[3] ), .A3(\a[4] ), .A4(\a[7] ), .ZN(new_n278_));
  NAND4_X1   g00085(.A1(\a[0] ), .A2(\a[2] ), .A3(\a[5] ), .A4(\a[7] ), .ZN(new_n279_));
  AOI22_X1   g00086(.A1(new_n256_), .A2(new_n243_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND4_X1   g00087(.A1(\a[2] ), .A2(\a[3] ), .A3(\a[4] ), .A4(\a[5] ), .ZN(new_n281_));
  NAND3_X1   g00088(.A1(new_n281_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n282_));
  OAI22_X1   g00089(.A1(new_n280_), .A2(new_n277_), .B1(new_n282_), .B2(new_n276_), .ZN(new_n283_));
  INV_X1     g00090(.I(new_n257_), .ZN(new_n284_));
  AOI21_X1   g00091(.A1(new_n248_), .A2(new_n245_), .B(new_n284_), .ZN(new_n285_));
  NOR4_X1    g00092(.A1(new_n242_), .A2(new_n194_), .A3(new_n197_), .A4(\a[6] ), .ZN(new_n286_));
  INV_X1     g00093(.I(new_n286_), .ZN(new_n287_));
  NAND2_X1   g00094(.A1(\a[1] ), .A2(\a[6] ), .ZN(new_n288_));
  NOR2_X1    g00095(.A1(new_n250_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1     g00096(.I(\a[4] ), .ZN(new_n290_));
  NOR2_X1    g00097(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1   g00098(.A1(\a[1] ), .A2(\a[6] ), .B(\a[4] ), .ZN(new_n292_));
  NOR2_X1    g00099(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1   g00100(.A1(new_n287_), .A2(new_n293_), .B(new_n289_), .ZN(new_n294_));
  NAND2_X1   g00101(.A1(new_n285_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1   g00102(.A1(new_n255_), .A2(new_n259_), .B(new_n257_), .ZN(new_n296_));
  NAND3_X1   g00103(.A1(\a[1] ), .A2(\a[4] ), .A3(\a[6] ), .ZN(new_n297_));
  NAND2_X1   g00104(.A1(new_n288_), .A2(new_n290_), .ZN(new_n298_));
  NAND2_X1   g00105(.A1(new_n298_), .A2(new_n297_), .ZN(new_n299_));
  AOI21_X1   g00106(.A1(new_n299_), .A2(new_n250_), .B(new_n286_), .ZN(new_n300_));
  NAND2_X1   g00107(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1   g00108(.A1(new_n295_), .A2(new_n301_), .B(new_n283_), .ZN(new_n302_));
  NOR2_X1    g00109(.A1(new_n282_), .A2(new_n276_), .ZN(new_n303_));
  NOR2_X1    g00110(.A1(new_n280_), .A2(new_n277_), .ZN(new_n304_));
  NOR2_X1    g00111(.A1(new_n304_), .A2(new_n303_), .ZN(new_n305_));
  NOR2_X1    g00112(.A1(new_n296_), .A2(new_n300_), .ZN(new_n306_));
  NOR2_X1    g00113(.A1(new_n285_), .A2(new_n294_), .ZN(new_n307_));
  NOR3_X1    g00114(.A1(new_n307_), .A2(new_n306_), .A3(new_n305_), .ZN(new_n308_));
  NOR2_X1    g00115(.A1(new_n308_), .A2(new_n302_), .ZN(new_n309_));
  XOR2_X1    g00116(.A1(new_n275_), .A2(new_n309_), .Z(\asquared[8] ));
  AOI22_X1   g00117(.A1(\a[0] ), .A2(\a[8] ), .B1(\a[2] ), .B2(\a[6] ), .ZN(new_n311_));
  NAND4_X1   g00118(.A1(\a[0] ), .A2(\a[2] ), .A3(\a[6] ), .A4(\a[8] ), .ZN(new_n312_));
  INV_X1     g00119(.I(new_n312_), .ZN(new_n313_));
  NOR3_X1    g00120(.A1(new_n313_), .A2(new_n297_), .A3(new_n311_), .ZN(new_n314_));
  OAI21_X1   g00121(.A1(new_n297_), .A2(new_n311_), .B(new_n312_), .ZN(new_n315_));
  OAI22_X1   g00122(.A1(new_n314_), .A2(new_n297_), .B1(new_n315_), .B2(new_n311_), .ZN(new_n316_));
  INV_X1     g00123(.I(new_n282_), .ZN(new_n317_));
  NAND2_X1   g00124(.A1(\a[3] ), .A2(\a[5] ), .ZN(new_n318_));
  NAND2_X1   g00125(.A1(\a[1] ), .A2(\a[7] ), .ZN(new_n319_));
  XOR2_X1    g00126(.A1(new_n318_), .A2(new_n319_), .Z(new_n320_));
  NOR2_X1    g00127(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1   g00128(.A1(new_n318_), .A2(new_n319_), .ZN(new_n322_));
  NOR2_X1    g00129(.A1(new_n322_), .A2(new_n282_), .ZN(new_n323_));
  OAI21_X1   g00130(.A1(new_n321_), .A2(new_n323_), .B(new_n316_), .ZN(new_n324_));
  INV_X1     g00131(.I(new_n311_), .ZN(new_n325_));
  NAND3_X1   g00132(.A1(new_n325_), .A2(new_n291_), .A3(new_n312_), .ZN(new_n326_));
  INV_X1     g00133(.I(new_n315_), .ZN(new_n327_));
  AOI22_X1   g00134(.A1(new_n327_), .A2(new_n325_), .B1(new_n326_), .B2(new_n291_), .ZN(new_n328_));
  NAND2_X1   g00135(.A1(new_n322_), .A2(new_n282_), .ZN(new_n329_));
  NAND2_X1   g00136(.A1(new_n317_), .A2(new_n320_), .ZN(new_n330_));
  NAND3_X1   g00137(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1   g00138(.A1(new_n296_), .A2(new_n300_), .B(new_n286_), .ZN(new_n332_));
  INV_X1     g00139(.I(new_n332_), .ZN(new_n333_));
  AOI21_X1   g00140(.A1(new_n324_), .A2(new_n331_), .B(new_n333_), .ZN(new_n334_));
  AOI21_X1   g00141(.A1(new_n329_), .A2(new_n330_), .B(new_n328_), .ZN(new_n335_));
  NOR3_X1    g00142(.A1(new_n316_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n336_));
  NOR3_X1    g00143(.A1(new_n335_), .A2(new_n336_), .A3(new_n332_), .ZN(new_n337_));
  NOR2_X1    g00144(.A1(new_n337_), .A2(new_n334_), .ZN(new_n338_));
  INV_X1     g00145(.I(new_n308_), .ZN(new_n339_));
  OAI21_X1   g00146(.A1(new_n307_), .A2(new_n306_), .B(new_n305_), .ZN(new_n340_));
  OAI21_X1   g00147(.A1(new_n272_), .A2(new_n261_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1   g00148(.A1(new_n341_), .A2(new_n339_), .ZN(new_n342_));
  XOR2_X1    g00149(.A1(new_n342_), .A2(new_n338_), .Z(\asquared[9] ));
  INV_X1     g00150(.I(new_n337_), .ZN(new_n344_));
  OAI21_X1   g00151(.A1(new_n335_), .A2(new_n336_), .B(new_n332_), .ZN(new_n345_));
  AOI21_X1   g00152(.A1(new_n274_), .A2(new_n262_), .B(new_n302_), .ZN(new_n346_));
  OAI21_X1   g00153(.A1(new_n346_), .A2(new_n308_), .B(new_n345_), .ZN(new_n347_));
  NAND2_X1   g00154(.A1(new_n347_), .A2(new_n344_), .ZN(new_n348_));
  NOR2_X1    g00155(.A1(new_n317_), .A2(new_n322_), .ZN(new_n349_));
  INV_X1     g00156(.I(new_n349_), .ZN(new_n350_));
  NAND2_X1   g00157(.A1(new_n324_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1   g00158(.A1(\a[5] ), .A2(\a[8] ), .ZN(new_n352_));
  NOR2_X1    g00159(.A1(new_n352_), .A2(new_n194_), .ZN(new_n353_));
  INV_X1     g00160(.I(new_n353_), .ZN(new_n354_));
  INV_X1     g00161(.I(\a[8] ), .ZN(new_n355_));
  NOR2_X1    g00162(.A1(new_n194_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1   g00163(.A1(new_n356_), .A2(\a[5] ), .B(new_n354_), .ZN(new_n357_));
  NAND4_X1   g00164(.A1(\a[1] ), .A2(\a[3] ), .A3(\a[5] ), .A4(\a[7] ), .ZN(new_n358_));
  NAND2_X1   g00165(.A1(\a[0] ), .A2(\a[9] ), .ZN(new_n359_));
  XNOR2_X1   g00166(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1    g00167(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1     g00168(.I(new_n356_), .ZN(new_n362_));
  AOI21_X1   g00169(.A1(new_n362_), .A2(new_n253_), .B(new_n353_), .ZN(new_n363_));
  XOR2_X1    g00170(.A1(new_n358_), .A2(new_n359_), .Z(new_n364_));
  NOR2_X1    g00171(.A1(new_n364_), .A2(new_n363_), .ZN(new_n365_));
  NOR2_X1    g00172(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1     g00173(.I(\a[6] ), .ZN(new_n367_));
  NOR2_X1    g00174(.A1(new_n225_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1    g00175(.A1(new_n368_), .A2(new_n243_), .ZN(new_n369_));
  NAND2_X1   g00176(.A1(\a[3] ), .A2(\a[4] ), .ZN(new_n370_));
  NAND2_X1   g00177(.A1(\a[5] ), .A2(\a[6] ), .ZN(new_n371_));
  NOR2_X1    g00178(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1   g00179(.A1(\a[5] ), .A2(\a[7] ), .ZN(new_n373_));
  NAND2_X1   g00180(.A1(\a[6] ), .A2(\a[7] ), .ZN(new_n374_));
  OAI22_X1   g00181(.A1(new_n246_), .A2(new_n374_), .B1(new_n251_), .B2(new_n373_), .ZN(new_n375_));
  NOR3_X1    g00182(.A1(new_n369_), .A2(new_n375_), .A3(new_n372_), .ZN(new_n376_));
  INV_X1     g00183(.I(new_n372_), .ZN(new_n377_));
  NAND2_X1   g00184(.A1(\a[2] ), .A2(\a[7] ), .ZN(new_n378_));
  AOI21_X1   g00185(.A1(new_n377_), .A2(new_n375_), .B(new_n378_), .ZN(new_n379_));
  NOR3_X1    g00186(.A1(new_n379_), .A2(new_n376_), .A3(new_n327_), .ZN(new_n380_));
  OAI21_X1   g00187(.A1(new_n379_), .A2(new_n376_), .B(new_n327_), .ZN(new_n381_));
  INV_X1     g00188(.I(new_n381_), .ZN(new_n382_));
  OAI21_X1   g00189(.A1(new_n380_), .A2(new_n382_), .B(new_n366_), .ZN(new_n383_));
  NAND2_X1   g00190(.A1(new_n364_), .A2(new_n363_), .ZN(new_n384_));
  NAND2_X1   g00191(.A1(new_n357_), .A2(new_n360_), .ZN(new_n385_));
  NAND2_X1   g00192(.A1(new_n385_), .A2(new_n384_), .ZN(new_n386_));
  INV_X1     g00193(.I(new_n380_), .ZN(new_n387_));
  NAND3_X1   g00194(.A1(new_n386_), .A2(new_n387_), .A3(new_n381_), .ZN(new_n388_));
  AOI21_X1   g00195(.A1(new_n383_), .A2(new_n388_), .B(new_n351_), .ZN(new_n389_));
  NOR2_X1    g00196(.A1(new_n335_), .A2(new_n349_), .ZN(new_n390_));
  AOI21_X1   g00197(.A1(new_n387_), .A2(new_n381_), .B(new_n386_), .ZN(new_n391_));
  NOR3_X1    g00198(.A1(new_n366_), .A2(new_n382_), .A3(new_n380_), .ZN(new_n392_));
  NOR3_X1    g00199(.A1(new_n391_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  NOR2_X1    g00200(.A1(new_n393_), .A2(new_n389_), .ZN(new_n394_));
  XOR2_X1    g00201(.A1(new_n348_), .A2(new_n394_), .Z(\asquared[10] ));
  AOI21_X1   g00202(.A1(new_n347_), .A2(new_n344_), .B(new_n389_), .ZN(new_n396_));
  NOR2_X1    g00203(.A1(new_n396_), .A2(new_n393_), .ZN(new_n397_));
  OAI21_X1   g00204(.A1(new_n379_), .A2(new_n376_), .B(new_n315_), .ZN(new_n398_));
  INV_X1     g00205(.I(new_n398_), .ZN(new_n399_));
  NOR2_X1    g00206(.A1(new_n391_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1    g00207(.A1(new_n375_), .A2(new_n372_), .ZN(new_n401_));
  AOI22_X1   g00208(.A1(\a[1] ), .A2(\a[9] ), .B1(\a[4] ), .B2(\a[6] ), .ZN(new_n402_));
  INV_X1     g00209(.I(\a[9] ), .ZN(new_n403_));
  NOR2_X1    g00210(.A1(new_n297_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1    g00211(.A1(new_n404_), .A2(new_n402_), .ZN(new_n405_));
  NAND2_X1   g00212(.A1(new_n405_), .A2(new_n354_), .ZN(new_n406_));
  OAI21_X1   g00213(.A1(new_n404_), .A2(new_n402_), .B(new_n353_), .ZN(new_n407_));
  AOI21_X1   g00214(.A1(new_n406_), .A2(new_n407_), .B(new_n401_), .ZN(new_n408_));
  INV_X1     g00215(.I(new_n408_), .ZN(new_n409_));
  NAND3_X1   g00216(.A1(new_n406_), .A2(new_n401_), .A3(new_n407_), .ZN(new_n410_));
  NAND2_X1   g00217(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1   g00218(.A1(\a[0] ), .A2(\a[2] ), .ZN(new_n412_));
  NAND2_X1   g00219(.A1(\a[8] ), .A2(\a[10] ), .ZN(new_n413_));
  NOR2_X1    g00220(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1   g00221(.A1(\a[7] ), .A2(\a[8] ), .ZN(new_n415_));
  NOR2_X1    g00222(.A1(new_n246_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1     g00223(.I(\a[10] ), .ZN(new_n417_));
  NOR2_X1    g00224(.A1(new_n196_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1   g00225(.A1(new_n418_), .A2(\a[3] ), .A3(\a[7] ), .ZN(new_n419_));
  OAI21_X1   g00226(.A1(new_n414_), .A2(new_n416_), .B(new_n419_), .ZN(new_n420_));
  NOR2_X1    g00227(.A1(new_n197_), .A2(new_n355_), .ZN(new_n421_));
  INV_X1     g00228(.I(\a[7] ), .ZN(new_n422_));
  OAI22_X1   g00229(.A1(new_n196_), .A2(new_n417_), .B1(new_n225_), .B2(new_n422_), .ZN(new_n423_));
  NOR4_X1    g00230(.A1(new_n196_), .A2(new_n225_), .A3(new_n422_), .A4(new_n417_), .ZN(new_n424_));
  NOR3_X1    g00231(.A1(new_n424_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n425_));
  AOI22_X1   g00232(.A1(new_n420_), .A2(new_n421_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1    g00233(.A1(new_n358_), .A2(new_n359_), .ZN(new_n427_));
  INV_X1     g00234(.I(new_n427_), .ZN(new_n428_));
  NAND2_X1   g00235(.A1(new_n384_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1   g00236(.A1(new_n429_), .A2(new_n426_), .ZN(new_n430_));
  NOR2_X1    g00237(.A1(new_n429_), .A2(new_n426_), .ZN(new_n431_));
  INV_X1     g00238(.I(new_n431_), .ZN(new_n432_));
  AOI21_X1   g00239(.A1(new_n432_), .A2(new_n430_), .B(new_n411_), .ZN(new_n433_));
  INV_X1     g00240(.I(new_n410_), .ZN(new_n434_));
  NOR2_X1    g00241(.A1(new_n434_), .A2(new_n408_), .ZN(new_n435_));
  NAND2_X1   g00242(.A1(new_n420_), .A2(new_n421_), .ZN(new_n436_));
  NAND2_X1   g00243(.A1(new_n425_), .A2(new_n423_), .ZN(new_n437_));
  NAND2_X1   g00244(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1    g00245(.A1(new_n361_), .A2(new_n427_), .ZN(new_n439_));
  NOR2_X1    g00246(.A1(new_n439_), .A2(new_n438_), .ZN(new_n440_));
  NOR3_X1    g00247(.A1(new_n440_), .A2(new_n435_), .A3(new_n431_), .ZN(new_n441_));
  NOR3_X1    g00248(.A1(new_n400_), .A2(new_n433_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1     g00249(.I(new_n442_), .ZN(new_n443_));
  OAI21_X1   g00250(.A1(new_n433_), .A2(new_n441_), .B(new_n400_), .ZN(new_n444_));
  NAND2_X1   g00251(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1     g00252(.I(new_n393_), .ZN(new_n446_));
  AOI21_X1   g00253(.A1(new_n341_), .A2(new_n339_), .B(new_n334_), .ZN(new_n447_));
  OAI21_X1   g00254(.A1(new_n391_), .A2(new_n392_), .B(new_n390_), .ZN(new_n448_));
  OAI21_X1   g00255(.A1(new_n447_), .A2(new_n337_), .B(new_n448_), .ZN(new_n449_));
  NAND2_X1   g00256(.A1(new_n383_), .A2(new_n398_), .ZN(new_n450_));
  OAI21_X1   g00257(.A1(new_n440_), .A2(new_n431_), .B(new_n435_), .ZN(new_n451_));
  NAND3_X1   g00258(.A1(new_n432_), .A2(new_n411_), .A3(new_n430_), .ZN(new_n452_));
  AOI21_X1   g00259(.A1(new_n452_), .A2(new_n451_), .B(new_n450_), .ZN(new_n453_));
  AOI21_X1   g00260(.A1(new_n449_), .A2(new_n446_), .B(new_n453_), .ZN(new_n454_));
  AOI22_X1   g00261(.A1(new_n445_), .A2(new_n397_), .B1(new_n454_), .B2(new_n443_), .ZN(\asquared[11] ));
  OAI21_X1   g00262(.A1(new_n396_), .A2(new_n393_), .B(new_n444_), .ZN(new_n456_));
  NAND2_X1   g00263(.A1(new_n456_), .A2(new_n443_), .ZN(new_n457_));
  NOR2_X1    g00264(.A1(new_n288_), .A2(new_n417_), .ZN(new_n458_));
  NOR2_X1    g00265(.A1(new_n194_), .A2(new_n417_), .ZN(new_n459_));
  INV_X1     g00266(.I(new_n459_), .ZN(new_n460_));
  AOI21_X1   g00267(.A1(new_n460_), .A2(new_n367_), .B(new_n458_), .ZN(new_n461_));
  NAND2_X1   g00268(.A1(new_n461_), .A2(new_n425_), .ZN(new_n462_));
  INV_X1     g00269(.I(new_n462_), .ZN(new_n463_));
  NOR2_X1    g00270(.A1(new_n461_), .A2(new_n425_), .ZN(new_n464_));
  AOI22_X1   g00271(.A1(\a[2] ), .A2(\a[9] ), .B1(\a[3] ), .B2(\a[8] ), .ZN(new_n465_));
  INV_X1     g00272(.I(new_n465_), .ZN(new_n466_));
  NOR2_X1    g00273(.A1(new_n355_), .A2(new_n403_), .ZN(new_n467_));
  NAND2_X1   g00274(.A1(new_n467_), .A2(new_n256_), .ZN(new_n468_));
  NAND2_X1   g00275(.A1(new_n468_), .A2(new_n466_), .ZN(new_n469_));
  AOI22_X1   g00276(.A1(new_n466_), .A2(new_n404_), .B1(new_n256_), .B2(new_n467_), .ZN(new_n470_));
  AOI22_X1   g00277(.A1(new_n404_), .A2(new_n469_), .B1(new_n470_), .B2(new_n466_), .ZN(new_n471_));
  OAI21_X1   g00278(.A1(new_n463_), .A2(new_n464_), .B(new_n471_), .ZN(new_n472_));
  OR3_X2     g00279(.A1(new_n463_), .A2(new_n471_), .A3(new_n464_), .Z(new_n473_));
  INV_X1     g00280(.I(new_n405_), .ZN(new_n474_));
  NOR2_X1    g00281(.A1(new_n474_), .A2(new_n354_), .ZN(new_n475_));
  OAI21_X1   g00282(.A1(new_n290_), .A2(new_n422_), .B(new_n371_), .ZN(new_n476_));
  NAND2_X1   g00283(.A1(\a[0] ), .A2(\a[11] ), .ZN(new_n477_));
  INV_X1     g00284(.I(new_n477_), .ZN(new_n478_));
  INV_X1     g00285(.I(new_n374_), .ZN(new_n479_));
  NAND2_X1   g00286(.A1(new_n243_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1   g00287(.A1(new_n480_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n481_));
  AOI22_X1   g00288(.A1(new_n476_), .A2(new_n478_), .B1(new_n243_), .B2(new_n479_), .ZN(new_n482_));
  AOI22_X1   g00289(.A1(new_n481_), .A2(new_n478_), .B1(new_n482_), .B2(new_n476_), .ZN(new_n483_));
  OAI21_X1   g00290(.A1(new_n475_), .A2(new_n408_), .B(new_n483_), .ZN(new_n484_));
  NOR3_X1    g00291(.A1(new_n483_), .A2(new_n408_), .A3(new_n475_), .ZN(new_n485_));
  INV_X1     g00292(.I(new_n485_), .ZN(new_n486_));
  AOI22_X1   g00293(.A1(new_n486_), .A2(new_n484_), .B1(new_n473_), .B2(new_n472_), .ZN(new_n487_));
  INV_X1     g00294(.I(new_n472_), .ZN(new_n488_));
  NOR3_X1    g00295(.A1(new_n463_), .A2(new_n471_), .A3(new_n464_), .ZN(new_n489_));
  INV_X1     g00296(.I(new_n484_), .ZN(new_n490_));
  NOR4_X1    g00297(.A1(new_n488_), .A2(new_n490_), .A3(new_n489_), .A4(new_n485_), .ZN(new_n491_));
  NOR2_X1    g00298(.A1(new_n491_), .A2(new_n487_), .ZN(new_n492_));
  OAI21_X1   g00299(.A1(new_n426_), .A2(new_n439_), .B(new_n451_), .ZN(new_n493_));
  NOR2_X1    g00300(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI22_X1   g00301(.A1(new_n488_), .A2(new_n489_), .B1(new_n490_), .B2(new_n485_), .ZN(new_n495_));
  NAND4_X1   g00302(.A1(new_n486_), .A2(new_n473_), .A3(new_n472_), .A4(new_n484_), .ZN(new_n496_));
  NAND2_X1   g00303(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1   g00304(.A1(new_n438_), .A2(new_n429_), .B(new_n433_), .ZN(new_n498_));
  NOR2_X1    g00305(.A1(new_n498_), .A2(new_n497_), .ZN(new_n499_));
  NOR2_X1    g00306(.A1(new_n499_), .A2(new_n494_), .ZN(new_n500_));
  XOR2_X1    g00307(.A1(new_n457_), .A2(new_n500_), .Z(\asquared[12] ));
  AOI21_X1   g00308(.A1(new_n456_), .A2(new_n443_), .B(new_n494_), .ZN(new_n502_));
  NOR2_X1    g00309(.A1(new_n502_), .A2(new_n499_), .ZN(new_n503_));
  NOR2_X1    g00310(.A1(new_n408_), .A2(new_n475_), .ZN(new_n504_));
  NOR2_X1    g00311(.A1(new_n504_), .A2(new_n483_), .ZN(new_n505_));
  NOR2_X1    g00312(.A1(new_n487_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1     g00313(.I(new_n461_), .ZN(new_n507_));
  NOR2_X1    g00314(.A1(new_n507_), .A2(new_n425_), .ZN(new_n508_));
  INV_X1     g00315(.I(new_n464_), .ZN(new_n509_));
  AOI21_X1   g00316(.A1(new_n462_), .A2(new_n509_), .B(new_n471_), .ZN(new_n510_));
  NOR2_X1    g00317(.A1(new_n510_), .A2(new_n508_), .ZN(new_n511_));
  AOI21_X1   g00318(.A1(\a[4] ), .A2(\a[8] ), .B(new_n458_), .ZN(new_n512_));
  INV_X1     g00319(.I(\a[11] ), .ZN(new_n513_));
  OAI21_X1   g00320(.A1(new_n194_), .A2(new_n513_), .B(new_n373_), .ZN(new_n514_));
  NAND2_X1   g00321(.A1(\a[5] ), .A2(\a[11] ), .ZN(new_n515_));
  NOR2_X1    g00322(.A1(new_n319_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1     g00323(.I(new_n516_), .ZN(new_n517_));
  NAND2_X1   g00324(.A1(new_n517_), .A2(new_n514_), .ZN(new_n518_));
  NAND3_X1   g00325(.A1(new_n458_), .A2(\a[4] ), .A3(\a[8] ), .ZN(new_n519_));
  INV_X1     g00326(.I(new_n519_), .ZN(new_n520_));
  NOR3_X1    g00327(.A1(new_n518_), .A2(new_n520_), .A3(new_n512_), .ZN(new_n521_));
  OAI21_X1   g00328(.A1(new_n518_), .A2(new_n512_), .B(new_n519_), .ZN(new_n522_));
  OAI22_X1   g00329(.A1(new_n521_), .A2(new_n518_), .B1(new_n522_), .B2(new_n512_), .ZN(new_n523_));
  INV_X1     g00330(.I(new_n523_), .ZN(new_n524_));
  NAND2_X1   g00331(.A1(new_n511_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1     g00332(.I(new_n525_), .ZN(new_n526_));
  NOR2_X1    g00333(.A1(new_n511_), .A2(new_n524_), .ZN(new_n527_));
  NAND2_X1   g00334(.A1(new_n470_), .A2(new_n482_), .ZN(new_n528_));
  NOR2_X1    g00335(.A1(new_n470_), .A2(new_n482_), .ZN(new_n529_));
  INV_X1     g00336(.I(new_n529_), .ZN(new_n530_));
  NAND2_X1   g00337(.A1(new_n530_), .A2(new_n528_), .ZN(new_n531_));
  NAND2_X1   g00338(.A1(\a[3] ), .A2(\a[9] ), .ZN(new_n532_));
  INV_X1     g00339(.I(new_n412_), .ZN(new_n533_));
  NAND2_X1   g00340(.A1(\a[10] ), .A2(\a[12] ), .ZN(new_n534_));
  INV_X1     g00341(.I(new_n534_), .ZN(new_n535_));
  INV_X1     g00342(.I(\a[12] ), .ZN(new_n536_));
  NOR2_X1    g00343(.A1(new_n196_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1   g00344(.A1(new_n537_), .A2(\a[3] ), .A3(\a[9] ), .ZN(new_n538_));
  NAND2_X1   g00345(.A1(\a[9] ), .A2(\a[10] ), .ZN(new_n539_));
  INV_X1     g00346(.I(new_n539_), .ZN(new_n540_));
  NAND2_X1   g00347(.A1(new_n256_), .A2(new_n540_), .ZN(new_n541_));
  AOI22_X1   g00348(.A1(new_n538_), .A2(new_n541_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n542_));
  AOI21_X1   g00349(.A1(\a[2] ), .A2(\a[10] ), .B(new_n537_), .ZN(new_n543_));
  NAND2_X1   g00350(.A1(new_n533_), .A2(new_n535_), .ZN(new_n544_));
  NAND3_X1   g00351(.A1(new_n544_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n545_));
  OAI22_X1   g00352(.A1(new_n542_), .A2(new_n532_), .B1(new_n545_), .B2(new_n543_), .ZN(new_n546_));
  XOR2_X1    g00353(.A1(new_n531_), .A2(new_n546_), .Z(new_n547_));
  NOR3_X1    g00354(.A1(new_n526_), .A2(new_n527_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1     g00355(.I(new_n527_), .ZN(new_n549_));
  XNOR2_X1   g00356(.A1(new_n531_), .A2(new_n546_), .ZN(new_n550_));
  AOI21_X1   g00357(.A1(new_n549_), .A2(new_n525_), .B(new_n550_), .ZN(new_n551_));
  NOR3_X1    g00358(.A1(new_n551_), .A2(new_n548_), .A3(new_n506_), .ZN(new_n552_));
  INV_X1     g00359(.I(new_n552_), .ZN(new_n553_));
  OAI21_X1   g00360(.A1(new_n551_), .A2(new_n548_), .B(new_n506_), .ZN(new_n554_));
  NAND2_X1   g00361(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1     g00362(.I(new_n499_), .ZN(new_n556_));
  NAND2_X1   g00363(.A1(new_n498_), .A2(new_n497_), .ZN(new_n557_));
  OAI21_X1   g00364(.A1(new_n454_), .A2(new_n442_), .B(new_n557_), .ZN(new_n558_));
  INV_X1     g00365(.I(new_n506_), .ZN(new_n559_));
  NAND3_X1   g00366(.A1(new_n549_), .A2(new_n525_), .A3(new_n550_), .ZN(new_n560_));
  OAI21_X1   g00367(.A1(new_n526_), .A2(new_n527_), .B(new_n547_), .ZN(new_n561_));
  AOI21_X1   g00368(.A1(new_n561_), .A2(new_n560_), .B(new_n559_), .ZN(new_n562_));
  AOI21_X1   g00369(.A1(new_n558_), .A2(new_n556_), .B(new_n562_), .ZN(new_n563_));
  AOI22_X1   g00370(.A1(new_n563_), .A2(new_n553_), .B1(new_n555_), .B2(new_n503_), .ZN(\asquared[13] ));
  OAI21_X1   g00371(.A1(new_n502_), .A2(new_n499_), .B(new_n554_), .ZN(new_n565_));
  NAND2_X1   g00372(.A1(new_n565_), .A2(new_n553_), .ZN(new_n566_));
  OAI21_X1   g00373(.A1(new_n547_), .A2(new_n526_), .B(new_n549_), .ZN(new_n567_));
  INV_X1     g00374(.I(new_n545_), .ZN(new_n568_));
  NOR2_X1    g00375(.A1(new_n517_), .A2(\a[12] ), .ZN(new_n569_));
  NOR2_X1    g00376(.A1(new_n319_), .A2(new_n536_), .ZN(new_n570_));
  INV_X1     g00377(.I(new_n570_), .ZN(new_n571_));
  OAI21_X1   g00378(.A1(new_n194_), .A2(new_n536_), .B(new_n422_), .ZN(new_n572_));
  AOI21_X1   g00379(.A1(new_n571_), .A2(new_n572_), .B(new_n516_), .ZN(new_n573_));
  OR2_X2     g00380(.A1(new_n573_), .A2(new_n569_), .Z(new_n574_));
  XOR2_X1    g00381(.A1(new_n574_), .A2(new_n568_), .Z(new_n575_));
  AOI21_X1   g00382(.A1(new_n546_), .A2(new_n528_), .B(new_n529_), .ZN(new_n576_));
  INV_X1     g00383(.I(new_n576_), .ZN(new_n577_));
  NOR2_X1    g00384(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1    g00385(.A1(new_n574_), .A2(new_n545_), .Z(new_n579_));
  NOR2_X1    g00386(.A1(new_n579_), .A2(new_n576_), .ZN(new_n580_));
  NOR2_X1    g00387(.A1(new_n580_), .A2(new_n578_), .ZN(new_n581_));
  NOR2_X1    g00388(.A1(new_n567_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1   g00389(.A1(new_n550_), .A2(new_n525_), .B(new_n527_), .ZN(new_n583_));
  INV_X1     g00390(.I(new_n581_), .ZN(new_n584_));
  NOR2_X1    g00391(.A1(new_n584_), .A2(new_n583_), .ZN(new_n585_));
  INV_X1     g00392(.I(new_n352_), .ZN(new_n586_));
  NOR2_X1    g00393(.A1(new_n586_), .A2(new_n479_), .ZN(new_n587_));
  NAND2_X1   g00394(.A1(\a[2] ), .A2(\a[11] ), .ZN(new_n588_));
  NOR2_X1    g00395(.A1(new_n371_), .A2(new_n415_), .ZN(new_n589_));
  NOR3_X1    g00396(.A1(new_n587_), .A2(new_n589_), .A3(new_n588_), .ZN(new_n590_));
  NOR2_X1    g00397(.A1(new_n590_), .A2(new_n589_), .ZN(new_n591_));
  INV_X1     g00398(.I(new_n591_), .ZN(new_n592_));
  OAI22_X1   g00399(.A1(new_n592_), .A2(new_n587_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n593_));
  INV_X1     g00400(.I(new_n593_), .ZN(new_n594_));
  NAND2_X1   g00401(.A1(\a[0] ), .A2(\a[4] ), .ZN(new_n595_));
  NAND2_X1   g00402(.A1(\a[9] ), .A2(\a[13] ), .ZN(new_n596_));
  INV_X1     g00403(.I(\a[13] ), .ZN(new_n597_));
  NOR4_X1    g00404(.A1(new_n196_), .A2(new_n225_), .A3(new_n417_), .A4(new_n597_), .ZN(new_n598_));
  NOR2_X1    g00405(.A1(new_n370_), .A2(new_n539_), .ZN(new_n599_));
  OAI22_X1   g00406(.A1(new_n598_), .A2(new_n599_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n600_));
  NAND3_X1   g00407(.A1(new_n600_), .A2(\a[3] ), .A3(\a[10] ), .ZN(new_n601_));
  OAI22_X1   g00408(.A1(new_n196_), .A2(new_n597_), .B1(new_n290_), .B2(new_n403_), .ZN(new_n602_));
  NOR2_X1    g00409(.A1(new_n595_), .A2(new_n596_), .ZN(new_n603_));
  NOR3_X1    g00410(.A1(new_n598_), .A2(new_n603_), .A3(new_n599_), .ZN(new_n604_));
  NAND2_X1   g00411(.A1(new_n604_), .A2(new_n602_), .ZN(new_n605_));
  NAND2_X1   g00412(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1   g00413(.A1(new_n606_), .A2(new_n522_), .ZN(new_n607_));
  NOR2_X1    g00414(.A1(new_n607_), .A2(new_n594_), .ZN(new_n608_));
  INV_X1     g00415(.I(new_n608_), .ZN(new_n609_));
  NAND2_X1   g00416(.A1(new_n607_), .A2(new_n594_), .ZN(new_n610_));
  NAND2_X1   g00417(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR3_X1    g00418(.A1(new_n582_), .A2(new_n585_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1   g00419(.A1(new_n584_), .A2(new_n583_), .ZN(new_n613_));
  NAND2_X1   g00420(.A1(new_n567_), .A2(new_n581_), .ZN(new_n614_));
  AOI22_X1   g00421(.A1(new_n613_), .A2(new_n614_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n615_));
  NOR2_X1    g00422(.A1(new_n615_), .A2(new_n612_), .ZN(new_n616_));
  XOR2_X1    g00423(.A1(new_n566_), .A2(new_n616_), .Z(\asquared[14] ));
  OAI22_X1   g00424(.A1(new_n568_), .A2(new_n573_), .B1(\a[12] ), .B2(new_n517_), .ZN(new_n618_));
  NAND2_X1   g00425(.A1(\a[11] ), .A2(\a[12] ), .ZN(new_n619_));
  NOR2_X1    g00426(.A1(new_n246_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1     g00427(.I(new_n620_), .ZN(new_n621_));
  NAND2_X1   g00428(.A1(\a[3] ), .A2(\a[14] ), .ZN(new_n622_));
  NAND2_X1   g00429(.A1(\a[12] ), .A2(\a[14] ), .ZN(new_n623_));
  OAI22_X1   g00430(.A1(new_n412_), .A2(new_n623_), .B1(new_n477_), .B2(new_n622_), .ZN(new_n624_));
  NAND2_X1   g00431(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1   g00432(.A1(new_n625_), .A2(\a[0] ), .A3(\a[14] ), .ZN(new_n626_));
  OAI22_X1   g00433(.A1(new_n197_), .A2(new_n536_), .B1(new_n225_), .B2(new_n513_), .ZN(new_n627_));
  NOR2_X1    g00434(.A1(new_n624_), .A2(new_n620_), .ZN(new_n628_));
  NAND2_X1   g00435(.A1(new_n628_), .A2(new_n627_), .ZN(new_n629_));
  NAND2_X1   g00436(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1    g00437(.A1(new_n242_), .A2(new_n539_), .ZN(new_n631_));
  AOI22_X1   g00438(.A1(\a[4] ), .A2(\a[10] ), .B1(\a[5] ), .B2(\a[9] ), .ZN(new_n632_));
  OAI21_X1   g00439(.A1(new_n631_), .A2(new_n632_), .B(new_n570_), .ZN(new_n633_));
  INV_X1     g00440(.I(new_n632_), .ZN(new_n634_));
  AOI21_X1   g00441(.A1(new_n634_), .A2(new_n570_), .B(new_n631_), .ZN(new_n635_));
  NAND2_X1   g00442(.A1(new_n635_), .A2(new_n634_), .ZN(new_n636_));
  NAND2_X1   g00443(.A1(new_n636_), .A2(new_n633_), .ZN(new_n637_));
  XOR2_X1    g00444(.A1(new_n630_), .A2(new_n637_), .Z(new_n638_));
  NAND2_X1   g00445(.A1(new_n638_), .A2(new_n618_), .ZN(new_n639_));
  OR2_X2     g00446(.A1(new_n638_), .A2(new_n618_), .Z(new_n640_));
  NAND2_X1   g00447(.A1(new_n640_), .A2(new_n639_), .ZN(new_n641_));
  INV_X1     g00448(.I(new_n641_), .ZN(new_n642_));
  NAND2_X1   g00449(.A1(\a[6] ), .A2(\a[8] ), .ZN(new_n643_));
  NOR3_X1    g00450(.A1(new_n643_), .A2(new_n194_), .A3(new_n597_), .ZN(new_n644_));
  INV_X1     g00451(.I(new_n643_), .ZN(new_n645_));
  AOI21_X1   g00452(.A1(\a[1] ), .A2(\a[13] ), .B(new_n645_), .ZN(new_n646_));
  NOR2_X1    g00453(.A1(new_n646_), .A2(new_n644_), .ZN(new_n647_));
  XNOR2_X1   g00454(.A1(new_n591_), .A2(new_n647_), .ZN(new_n648_));
  XOR2_X1    g00455(.A1(new_n648_), .A2(new_n604_), .Z(new_n649_));
  INV_X1     g00456(.I(new_n649_), .ZN(new_n650_));
  NAND2_X1   g00457(.A1(new_n606_), .A2(new_n522_), .ZN(new_n651_));
  NAND2_X1   g00458(.A1(new_n609_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1    g00459(.A1(new_n652_), .A2(new_n650_), .ZN(new_n653_));
  AOI21_X1   g00460(.A1(new_n522_), .A2(new_n606_), .B(new_n608_), .ZN(new_n654_));
  NOR2_X1    g00461(.A1(new_n654_), .A2(new_n649_), .ZN(new_n655_));
  OAI21_X1   g00462(.A1(new_n653_), .A2(new_n655_), .B(new_n642_), .ZN(new_n656_));
  NAND2_X1   g00463(.A1(new_n654_), .A2(new_n649_), .ZN(new_n657_));
  NAND2_X1   g00464(.A1(new_n652_), .A2(new_n650_), .ZN(new_n658_));
  NAND3_X1   g00465(.A1(new_n658_), .A2(new_n657_), .A3(new_n641_), .ZN(new_n659_));
  NOR2_X1    g00466(.A1(new_n585_), .A2(new_n580_), .ZN(new_n660_));
  AOI21_X1   g00467(.A1(new_n656_), .A2(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1     g00468(.I(new_n661_), .ZN(new_n662_));
  NAND3_X1   g00469(.A1(new_n656_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n663_));
  NAND2_X1   g00470(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1   g00471(.A1(new_n565_), .A2(new_n553_), .B(new_n615_), .ZN(new_n665_));
  NOR2_X1    g00472(.A1(new_n665_), .A2(new_n612_), .ZN(new_n666_));
  INV_X1     g00473(.I(new_n612_), .ZN(new_n667_));
  AOI21_X1   g00474(.A1(new_n658_), .A2(new_n657_), .B(new_n641_), .ZN(new_n668_));
  NOR3_X1    g00475(.A1(new_n653_), .A2(new_n642_), .A3(new_n655_), .ZN(new_n669_));
  NOR4_X1    g00476(.A1(new_n669_), .A2(new_n668_), .A3(new_n580_), .A4(new_n585_), .ZN(new_n670_));
  OAI21_X1   g00477(.A1(new_n582_), .A2(new_n585_), .B(new_n611_), .ZN(new_n671_));
  OAI21_X1   g00478(.A1(new_n563_), .A2(new_n552_), .B(new_n671_), .ZN(new_n672_));
  AOI21_X1   g00479(.A1(new_n672_), .A2(new_n667_), .B(new_n670_), .ZN(new_n673_));
  AOI22_X1   g00480(.A1(new_n673_), .A2(new_n662_), .B1(new_n664_), .B2(new_n666_), .ZN(\asquared[15] ));
  OAI21_X1   g00481(.A1(new_n665_), .A2(new_n612_), .B(new_n663_), .ZN(new_n675_));
  NAND2_X1   g00482(.A1(new_n675_), .A2(new_n662_), .ZN(new_n676_));
  AOI21_X1   g00483(.A1(new_n642_), .A2(new_n657_), .B(new_n655_), .ZN(new_n677_));
  INV_X1     g00484(.I(new_n677_), .ZN(new_n678_));
  NAND2_X1   g00485(.A1(new_n592_), .A2(new_n647_), .ZN(new_n679_));
  INV_X1     g00486(.I(new_n648_), .ZN(new_n680_));
  OAI21_X1   g00487(.A1(new_n680_), .A2(new_n604_), .B(new_n679_), .ZN(new_n681_));
  NOR2_X1    g00488(.A1(new_n290_), .A2(new_n513_), .ZN(new_n682_));
  NOR2_X1    g00489(.A1(new_n644_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1     g00490(.I(new_n683_), .ZN(new_n684_));
  AND2_X2    g00491(.A1(new_n644_), .A2(new_n682_), .Z(new_n685_));
  NAND2_X1   g00492(.A1(\a[1] ), .A2(\a[14] ), .ZN(new_n686_));
  XOR2_X1    g00493(.A1(new_n686_), .A2(new_n355_), .Z(new_n687_));
  AOI21_X1   g00494(.A1(new_n684_), .A2(new_n687_), .B(new_n685_), .ZN(new_n688_));
  NAND2_X1   g00495(.A1(new_n688_), .A2(new_n684_), .ZN(new_n689_));
  OAI21_X1   g00496(.A1(new_n685_), .A2(new_n683_), .B(new_n687_), .ZN(new_n690_));
  NAND2_X1   g00497(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1   g00498(.A1(\a[2] ), .A2(\a[13] ), .ZN(new_n692_));
  INV_X1     g00499(.I(new_n415_), .ZN(new_n693_));
  AOI21_X1   g00500(.A1(\a[6] ), .A2(\a[9] ), .B(new_n693_), .ZN(new_n694_));
  INV_X1     g00501(.I(new_n694_), .ZN(new_n695_));
  NAND3_X1   g00502(.A1(new_n693_), .A2(\a[6] ), .A3(\a[9] ), .ZN(new_n696_));
  AOI21_X1   g00503(.A1(new_n695_), .A2(new_n696_), .B(new_n692_), .ZN(new_n697_));
  OAI21_X1   g00504(.A1(new_n694_), .A2(new_n692_), .B(new_n696_), .ZN(new_n698_));
  NOR2_X1    g00505(.A1(new_n698_), .A2(new_n694_), .ZN(new_n699_));
  NOR2_X1    g00506(.A1(new_n699_), .A2(new_n697_), .ZN(new_n700_));
  XNOR2_X1   g00507(.A1(new_n691_), .A2(new_n700_), .ZN(new_n701_));
  XOR2_X1    g00508(.A1(new_n701_), .A2(new_n681_), .Z(new_n702_));
  INV_X1     g00509(.I(new_n702_), .ZN(new_n703_));
  NAND2_X1   g00510(.A1(new_n630_), .A2(new_n637_), .ZN(new_n704_));
  NAND2_X1   g00511(.A1(new_n639_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1   g00512(.A1(new_n628_), .A2(new_n635_), .ZN(new_n706_));
  NOR2_X1    g00513(.A1(new_n628_), .A2(new_n635_), .ZN(new_n707_));
  INV_X1     g00514(.I(new_n707_), .ZN(new_n708_));
  NAND2_X1   g00515(.A1(new_n708_), .A2(new_n706_), .ZN(new_n709_));
  NAND2_X1   g00516(.A1(\a[10] ), .A2(\a[15] ), .ZN(new_n710_));
  OAI22_X1   g00517(.A1(new_n196_), .A2(new_n710_), .B1(new_n534_), .B2(new_n225_), .ZN(new_n711_));
  NAND4_X1   g00518(.A1(\a[0] ), .A2(\a[3] ), .A3(\a[12] ), .A4(\a[15] ), .ZN(new_n712_));
  NAND3_X1   g00519(.A1(new_n711_), .A2(\a[5] ), .A3(new_n712_), .ZN(new_n713_));
  NAND3_X1   g00520(.A1(new_n713_), .A2(\a[5] ), .A3(\a[10] ), .ZN(new_n714_));
  INV_X1     g00521(.I(new_n712_), .ZN(new_n715_));
  AOI21_X1   g00522(.A1(new_n711_), .A2(\a[5] ), .B(new_n715_), .ZN(new_n716_));
  INV_X1     g00523(.I(\a[15] ), .ZN(new_n717_));
  OAI22_X1   g00524(.A1(new_n196_), .A2(new_n717_), .B1(new_n225_), .B2(new_n536_), .ZN(new_n718_));
  NAND2_X1   g00525(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1   g00526(.A1(new_n714_), .A2(new_n719_), .ZN(new_n720_));
  XOR2_X1    g00527(.A1(new_n709_), .A2(new_n720_), .Z(new_n721_));
  XNOR2_X1   g00528(.A1(new_n705_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1    g00529(.A1(new_n703_), .A2(new_n722_), .ZN(new_n723_));
  XOR2_X1    g00530(.A1(new_n705_), .A2(new_n721_), .Z(new_n724_));
  NOR2_X1    g00531(.A1(new_n724_), .A2(new_n702_), .ZN(new_n725_));
  NOR3_X1    g00532(.A1(new_n723_), .A2(new_n678_), .A3(new_n725_), .ZN(new_n726_));
  NOR2_X1    g00533(.A1(new_n723_), .A2(new_n725_), .ZN(new_n727_));
  NOR2_X1    g00534(.A1(new_n727_), .A2(new_n677_), .ZN(new_n728_));
  NOR2_X1    g00535(.A1(new_n728_), .A2(new_n726_), .ZN(new_n729_));
  XOR2_X1    g00536(.A1(new_n676_), .A2(new_n729_), .Z(\asquared[16] ));
  INV_X1     g00537(.I(new_n728_), .ZN(new_n731_));
  NAND2_X1   g00538(.A1(new_n727_), .A2(new_n677_), .ZN(new_n732_));
  OAI21_X1   g00539(.A1(new_n673_), .A2(new_n661_), .B(new_n732_), .ZN(new_n733_));
  NAND2_X1   g00540(.A1(new_n733_), .A2(new_n731_), .ZN(new_n734_));
  AOI21_X1   g00541(.A1(new_n639_), .A2(new_n704_), .B(new_n721_), .ZN(new_n735_));
  AOI21_X1   g00542(.A1(new_n722_), .A2(new_n702_), .B(new_n735_), .ZN(new_n736_));
  INV_X1     g00543(.I(new_n736_), .ZN(new_n737_));
  INV_X1     g00544(.I(new_n691_), .ZN(new_n738_));
  NAND2_X1   g00545(.A1(new_n701_), .A2(new_n681_), .ZN(new_n739_));
  OAI21_X1   g00546(.A1(new_n738_), .A2(new_n700_), .B(new_n739_), .ZN(new_n740_));
  XOR2_X1    g00547(.A1(new_n688_), .A2(new_n716_), .Z(new_n741_));
  INV_X1     g00548(.I(\a[16] ), .ZN(new_n742_));
  NOR2_X1    g00549(.A1(new_n367_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1     g00550(.I(new_n515_), .ZN(new_n744_));
  NAND3_X1   g00551(.A1(new_n744_), .A2(\a[0] ), .A3(\a[16] ), .ZN(new_n745_));
  INV_X1     g00552(.I(new_n371_), .ZN(new_n746_));
  NOR2_X1    g00553(.A1(new_n417_), .A2(new_n513_), .ZN(new_n747_));
  NAND2_X1   g00554(.A1(new_n747_), .A2(new_n746_), .ZN(new_n748_));
  AOI22_X1   g00555(.A1(new_n748_), .A2(new_n745_), .B1(new_n418_), .B2(new_n743_), .ZN(new_n749_));
  AOI22_X1   g00556(.A1(\a[0] ), .A2(\a[16] ), .B1(\a[6] ), .B2(\a[10] ), .ZN(new_n750_));
  NAND2_X1   g00557(.A1(new_n418_), .A2(new_n743_), .ZN(new_n751_));
  NAND3_X1   g00558(.A1(new_n751_), .A2(new_n748_), .A3(new_n745_), .ZN(new_n752_));
  OAI22_X1   g00559(.A1(new_n749_), .A2(new_n515_), .B1(new_n752_), .B2(new_n750_), .ZN(new_n753_));
  XOR2_X1    g00560(.A1(new_n741_), .A2(new_n753_), .Z(new_n754_));
  XNOR2_X1   g00561(.A1(new_n740_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1     g00562(.I(new_n720_), .ZN(new_n756_));
  OAI21_X1   g00563(.A1(new_n756_), .A2(new_n709_), .B(new_n708_), .ZN(new_n757_));
  NAND2_X1   g00564(.A1(\a[4] ), .A2(\a[12] ), .ZN(new_n758_));
  INV_X1     g00565(.I(\a[14] ), .ZN(new_n759_));
  NOR2_X1    g00566(.A1(new_n597_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1     g00567(.I(new_n370_), .ZN(new_n761_));
  INV_X1     g00568(.I(new_n623_), .ZN(new_n762_));
  NOR2_X1    g00569(.A1(new_n536_), .A2(new_n597_), .ZN(new_n763_));
  AOI22_X1   g00570(.A1(new_n761_), .A2(new_n763_), .B1(new_n252_), .B2(new_n762_), .ZN(new_n764_));
  AOI21_X1   g00571(.A1(new_n256_), .A2(new_n760_), .B(new_n764_), .ZN(new_n765_));
  AOI22_X1   g00572(.A1(\a[2] ), .A2(\a[14] ), .B1(\a[3] ), .B2(\a[13] ), .ZN(new_n766_));
  INV_X1     g00573(.I(new_n760_), .ZN(new_n767_));
  OAI21_X1   g00574(.A1(new_n246_), .A2(new_n767_), .B(new_n764_), .ZN(new_n768_));
  OAI22_X1   g00575(.A1(new_n758_), .A2(new_n765_), .B1(new_n768_), .B2(new_n766_), .ZN(new_n769_));
  XOR2_X1    g00576(.A1(new_n757_), .A2(new_n769_), .Z(new_n770_));
  NOR2_X1    g00577(.A1(new_n686_), .A2(new_n355_), .ZN(new_n771_));
  INV_X1     g00578(.I(new_n771_), .ZN(new_n772_));
  NAND2_X1   g00579(.A1(\a[7] ), .A2(\a[9] ), .ZN(new_n773_));
  NAND2_X1   g00580(.A1(\a[1] ), .A2(\a[15] ), .ZN(new_n774_));
  XNOR2_X1   g00581(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  XOR2_X1    g00582(.A1(new_n775_), .A2(new_n772_), .Z(new_n776_));
  XOR2_X1    g00583(.A1(new_n776_), .A2(new_n698_), .Z(new_n777_));
  XNOR2_X1   g00584(.A1(new_n770_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1   g00585(.A1(new_n755_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1    g00586(.A1(new_n740_), .A2(new_n754_), .ZN(new_n780_));
  NAND2_X1   g00587(.A1(new_n740_), .A2(new_n754_), .ZN(new_n781_));
  INV_X1     g00588(.I(new_n781_), .ZN(new_n782_));
  NOR2_X1    g00589(.A1(new_n782_), .A2(new_n780_), .ZN(new_n783_));
  INV_X1     g00590(.I(new_n778_), .ZN(new_n784_));
  NAND2_X1   g00591(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1   g00592(.A1(new_n785_), .A2(new_n779_), .B(new_n737_), .ZN(new_n786_));
  NOR2_X1    g00593(.A1(new_n783_), .A2(new_n784_), .ZN(new_n787_));
  NOR2_X1    g00594(.A1(new_n755_), .A2(new_n778_), .ZN(new_n788_));
  NOR3_X1    g00595(.A1(new_n787_), .A2(new_n788_), .A3(new_n736_), .ZN(new_n789_));
  NOR2_X1    g00596(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  XOR2_X1    g00597(.A1(new_n734_), .A2(new_n790_), .Z(\asquared[17] ));
  INV_X1     g00598(.I(new_n789_), .ZN(new_n792_));
  AOI21_X1   g00599(.A1(new_n675_), .A2(new_n662_), .B(new_n726_), .ZN(new_n793_));
  OAI21_X1   g00600(.A1(new_n787_), .A2(new_n788_), .B(new_n736_), .ZN(new_n794_));
  OAI21_X1   g00601(.A1(new_n793_), .A2(new_n728_), .B(new_n794_), .ZN(new_n795_));
  NAND2_X1   g00602(.A1(new_n795_), .A2(new_n792_), .ZN(new_n796_));
  NOR2_X1    g00603(.A1(new_n788_), .A2(new_n782_), .ZN(new_n797_));
  NAND2_X1   g00604(.A1(\a[9] ), .A2(\a[16] ), .ZN(new_n798_));
  NOR2_X1    g00605(.A1(new_n798_), .A2(new_n194_), .ZN(new_n799_));
  INV_X1     g00606(.I(new_n799_), .ZN(new_n800_));
  NOR2_X1    g00607(.A1(new_n194_), .A2(new_n742_), .ZN(new_n801_));
  OAI21_X1   g00608(.A1(\a[9] ), .A2(new_n801_), .B(new_n800_), .ZN(new_n802_));
  XNOR2_X1   g00609(.A1(new_n768_), .A2(new_n802_), .ZN(new_n803_));
  XNOR2_X1   g00610(.A1(new_n803_), .A2(new_n752_), .ZN(new_n804_));
  NOR2_X1    g00611(.A1(new_n688_), .A2(new_n716_), .ZN(new_n805_));
  AOI21_X1   g00612(.A1(new_n741_), .A2(new_n753_), .B(new_n805_), .ZN(new_n806_));
  NOR2_X1    g00613(.A1(new_n775_), .A2(new_n772_), .ZN(new_n807_));
  INV_X1     g00614(.I(new_n807_), .ZN(new_n808_));
  NAND2_X1   g00615(.A1(new_n776_), .A2(new_n698_), .ZN(new_n809_));
  NAND2_X1   g00616(.A1(new_n809_), .A2(new_n808_), .ZN(new_n810_));
  XOR2_X1    g00617(.A1(new_n806_), .A2(new_n810_), .Z(new_n811_));
  XOR2_X1    g00618(.A1(new_n811_), .A2(new_n804_), .Z(new_n812_));
  INV_X1     g00619(.I(new_n812_), .ZN(new_n813_));
  NAND2_X1   g00620(.A1(\a[0] ), .A2(\a[17] ), .ZN(new_n814_));
  NAND2_X1   g00621(.A1(\a[5] ), .A2(\a[12] ), .ZN(new_n815_));
  NAND2_X1   g00622(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1    g00623(.A1(new_n773_), .A2(new_n774_), .ZN(new_n817_));
  NOR2_X1    g00624(.A1(new_n814_), .A2(new_n815_), .ZN(new_n818_));
  AOI21_X1   g00625(.A1(new_n817_), .A2(new_n816_), .B(new_n818_), .ZN(new_n819_));
  NAND2_X1   g00626(.A1(new_n819_), .A2(new_n816_), .ZN(new_n820_));
  NAND2_X1   g00627(.A1(new_n817_), .A2(new_n816_), .ZN(new_n821_));
  OAI21_X1   g00628(.A1(new_n821_), .A2(new_n818_), .B(new_n817_), .ZN(new_n822_));
  NAND2_X1   g00629(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1   g00630(.A1(\a[7] ), .A2(\a[10] ), .B(new_n467_), .ZN(new_n824_));
  NAND2_X1   g00631(.A1(new_n693_), .A2(new_n540_), .ZN(new_n825_));
  OAI21_X1   g00632(.A1(new_n824_), .A2(new_n622_), .B(new_n825_), .ZN(new_n826_));
  NOR2_X1    g00633(.A1(new_n826_), .A2(new_n824_), .ZN(new_n827_));
  NOR2_X1    g00634(.A1(new_n824_), .A2(new_n622_), .ZN(new_n828_));
  AOI21_X1   g00635(.A1(new_n828_), .A2(new_n825_), .B(new_n622_), .ZN(new_n829_));
  NOR2_X1    g00636(.A1(new_n829_), .A2(new_n827_), .ZN(new_n830_));
  XNOR2_X1   g00637(.A1(new_n830_), .A2(new_n823_), .ZN(new_n831_));
  NOR2_X1    g00638(.A1(new_n513_), .A2(new_n717_), .ZN(new_n832_));
  NAND2_X1   g00639(.A1(\a[11] ), .A2(\a[13] ), .ZN(new_n833_));
  INV_X1     g00640(.I(new_n833_), .ZN(new_n834_));
  AOI22_X1   g00641(.A1(\a[2] ), .A2(new_n832_), .B1(new_n834_), .B2(\a[4] ), .ZN(new_n835_));
  NAND2_X1   g00642(.A1(\a[13] ), .A2(\a[15] ), .ZN(new_n836_));
  NOR2_X1    g00643(.A1(new_n251_), .A2(new_n836_), .ZN(new_n837_));
  NOR3_X1    g00644(.A1(new_n835_), .A2(new_n367_), .A3(new_n837_), .ZN(new_n838_));
  NOR2_X1    g00645(.A1(new_n367_), .A2(new_n513_), .ZN(new_n839_));
  INV_X1     g00646(.I(new_n839_), .ZN(new_n840_));
  NOR2_X1    g00647(.A1(new_n838_), .A2(new_n837_), .ZN(new_n841_));
  OAI22_X1   g00648(.A1(new_n197_), .A2(new_n717_), .B1(new_n290_), .B2(new_n597_), .ZN(new_n842_));
  NAND2_X1   g00649(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1   g00650(.A1(new_n838_), .A2(new_n840_), .B(new_n843_), .ZN(new_n844_));
  XNOR2_X1   g00651(.A1(new_n831_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1   g00652(.A1(new_n757_), .A2(new_n769_), .ZN(new_n846_));
  INV_X1     g00653(.I(new_n846_), .ZN(new_n847_));
  AND2_X2    g00654(.A1(new_n770_), .A2(new_n777_), .Z(new_n848_));
  NOR2_X1    g00655(.A1(new_n848_), .A2(new_n847_), .ZN(new_n849_));
  NAND2_X1   g00656(.A1(new_n849_), .A2(new_n845_), .ZN(new_n850_));
  NOR2_X1    g00657(.A1(new_n849_), .A2(new_n845_), .ZN(new_n851_));
  INV_X1     g00658(.I(new_n851_), .ZN(new_n852_));
  NAND2_X1   g00659(.A1(new_n852_), .A2(new_n850_), .ZN(new_n853_));
  NOR2_X1    g00660(.A1(new_n853_), .A2(new_n813_), .ZN(new_n854_));
  INV_X1     g00661(.I(new_n850_), .ZN(new_n855_));
  NOR2_X1    g00662(.A1(new_n855_), .A2(new_n851_), .ZN(new_n856_));
  NOR2_X1    g00663(.A1(new_n856_), .A2(new_n812_), .ZN(new_n857_));
  NOR3_X1    g00664(.A1(new_n857_), .A2(new_n854_), .A3(new_n797_), .ZN(new_n858_));
  NAND2_X1   g00665(.A1(new_n785_), .A2(new_n781_), .ZN(new_n859_));
  NAND2_X1   g00666(.A1(new_n856_), .A2(new_n812_), .ZN(new_n860_));
  NAND2_X1   g00667(.A1(new_n853_), .A2(new_n813_), .ZN(new_n861_));
  AOI21_X1   g00668(.A1(new_n860_), .A2(new_n861_), .B(new_n859_), .ZN(new_n862_));
  NOR2_X1    g00669(.A1(new_n862_), .A2(new_n858_), .ZN(new_n863_));
  XOR2_X1    g00670(.A1(new_n796_), .A2(new_n863_), .Z(\asquared[18] ));
  AOI21_X1   g00671(.A1(new_n795_), .A2(new_n792_), .B(new_n862_), .ZN(new_n865_));
  NOR2_X1    g00672(.A1(new_n865_), .A2(new_n858_), .ZN(new_n866_));
  XOR2_X1    g00673(.A1(new_n841_), .A2(new_n826_), .Z(new_n867_));
  XOR2_X1    g00674(.A1(new_n867_), .A2(new_n819_), .Z(new_n868_));
  INV_X1     g00675(.I(new_n802_), .ZN(new_n869_));
  NAND2_X1   g00676(.A1(new_n768_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1   g00677(.A1(new_n803_), .A2(new_n752_), .ZN(new_n871_));
  OAI21_X1   g00678(.A1(new_n827_), .A2(new_n829_), .B(new_n823_), .ZN(new_n872_));
  NAND2_X1   g00679(.A1(new_n831_), .A2(new_n844_), .ZN(new_n873_));
  NAND4_X1   g00680(.A1(new_n873_), .A2(new_n870_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n874_));
  NAND2_X1   g00681(.A1(new_n873_), .A2(new_n872_), .ZN(new_n875_));
  NAND2_X1   g00682(.A1(new_n871_), .A2(new_n870_), .ZN(new_n876_));
  NAND2_X1   g00683(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1   g00684(.A1(new_n877_), .A2(new_n868_), .A3(new_n874_), .ZN(new_n878_));
  INV_X1     g00685(.I(new_n868_), .ZN(new_n879_));
  XNOR2_X1   g00686(.A1(new_n875_), .A2(new_n876_), .ZN(new_n880_));
  NAND2_X1   g00687(.A1(new_n880_), .A2(new_n879_), .ZN(new_n881_));
  NAND2_X1   g00688(.A1(new_n881_), .A2(new_n878_), .ZN(new_n882_));
  NAND4_X1   g00689(.A1(\a[0] ), .A2(\a[5] ), .A3(\a[13] ), .A4(\a[18] ), .ZN(new_n883_));
  INV_X1     g00690(.I(\a[18] ), .ZN(new_n884_));
  NOR3_X1    g00691(.A1(new_n477_), .A2(new_n422_), .A3(new_n884_), .ZN(new_n885_));
  NOR2_X1    g00692(.A1(new_n373_), .A2(new_n833_), .ZN(new_n886_));
  OAI21_X1   g00693(.A1(new_n885_), .A2(new_n886_), .B(new_n883_), .ZN(new_n887_));
  NAND3_X1   g00694(.A1(new_n887_), .A2(\a[7] ), .A3(\a[11] ), .ZN(new_n888_));
  NAND2_X1   g00695(.A1(new_n887_), .A2(new_n883_), .ZN(new_n889_));
  AOI22_X1   g00696(.A1(\a[0] ), .A2(\a[18] ), .B1(\a[5] ), .B2(\a[13] ), .ZN(new_n890_));
  OAI21_X1   g00697(.A1(new_n889_), .A2(new_n890_), .B(new_n888_), .ZN(new_n891_));
  NAND2_X1   g00698(.A1(\a[4] ), .A2(\a[14] ), .ZN(new_n892_));
  NAND2_X1   g00699(.A1(\a[15] ), .A2(\a[16] ), .ZN(new_n893_));
  NOR2_X1    g00700(.A1(new_n246_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1    g00701(.A1(new_n759_), .A2(new_n742_), .ZN(new_n895_));
  NAND2_X1   g00702(.A1(new_n895_), .A2(new_n252_), .ZN(new_n896_));
  NOR2_X1    g00703(.A1(new_n759_), .A2(new_n717_), .ZN(new_n897_));
  NAND2_X1   g00704(.A1(new_n897_), .A2(new_n761_), .ZN(new_n898_));
  AOI21_X1   g00705(.A1(new_n896_), .A2(new_n898_), .B(new_n894_), .ZN(new_n899_));
  NOR2_X1    g00706(.A1(new_n197_), .A2(new_n742_), .ZN(new_n900_));
  AOI21_X1   g00707(.A1(\a[3] ), .A2(\a[15] ), .B(new_n900_), .ZN(new_n901_));
  INV_X1     g00708(.I(new_n894_), .ZN(new_n902_));
  NAND3_X1   g00709(.A1(new_n902_), .A2(new_n896_), .A3(new_n898_), .ZN(new_n903_));
  OAI22_X1   g00710(.A1(new_n901_), .A2(new_n903_), .B1(new_n899_), .B2(new_n892_), .ZN(new_n904_));
  XOR2_X1    g00711(.A1(new_n891_), .A2(new_n904_), .Z(new_n905_));
  AOI21_X1   g00712(.A1(\a[6] ), .A2(\a[12] ), .B(new_n799_), .ZN(new_n906_));
  NAND2_X1   g00713(.A1(\a[1] ), .A2(\a[17] ), .ZN(new_n907_));
  XNOR2_X1   g00714(.A1(new_n413_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1   g00715(.A1(new_n799_), .A2(\a[6] ), .A3(\a[12] ), .ZN(new_n909_));
  INV_X1     g00716(.I(new_n909_), .ZN(new_n910_));
  NOR2_X1    g00717(.A1(new_n910_), .A2(new_n906_), .ZN(new_n911_));
  OAI21_X1   g00718(.A1(new_n908_), .A2(new_n906_), .B(new_n909_), .ZN(new_n912_));
  OAI22_X1   g00719(.A1(new_n908_), .A2(new_n911_), .B1(new_n912_), .B2(new_n906_), .ZN(new_n913_));
  XNOR2_X1   g00720(.A1(new_n905_), .A2(new_n913_), .ZN(new_n914_));
  AOI21_X1   g00721(.A1(new_n808_), .A2(new_n809_), .B(new_n806_), .ZN(new_n915_));
  NOR2_X1    g00722(.A1(new_n811_), .A2(new_n804_), .ZN(new_n916_));
  NOR2_X1    g00723(.A1(new_n916_), .A2(new_n915_), .ZN(new_n917_));
  XNOR2_X1   g00724(.A1(new_n917_), .A2(new_n914_), .ZN(new_n918_));
  NOR2_X1    g00725(.A1(new_n918_), .A2(new_n882_), .ZN(new_n919_));
  NAND2_X1   g00726(.A1(new_n918_), .A2(new_n882_), .ZN(new_n920_));
  INV_X1     g00727(.I(new_n920_), .ZN(new_n921_));
  NOR2_X1    g00728(.A1(new_n854_), .A2(new_n851_), .ZN(new_n922_));
  NOR3_X1    g00729(.A1(new_n921_), .A2(new_n922_), .A3(new_n919_), .ZN(new_n923_));
  INV_X1     g00730(.I(new_n923_), .ZN(new_n924_));
  OAI21_X1   g00731(.A1(new_n919_), .A2(new_n921_), .B(new_n922_), .ZN(new_n925_));
  NAND2_X1   g00732(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  INV_X1     g00733(.I(new_n858_), .ZN(new_n927_));
  AOI21_X1   g00734(.A1(new_n733_), .A2(new_n731_), .B(new_n786_), .ZN(new_n928_));
  OAI21_X1   g00735(.A1(new_n857_), .A2(new_n854_), .B(new_n797_), .ZN(new_n929_));
  OAI21_X1   g00736(.A1(new_n928_), .A2(new_n789_), .B(new_n929_), .ZN(new_n930_));
  INV_X1     g00737(.I(new_n919_), .ZN(new_n931_));
  NAND2_X1   g00738(.A1(new_n860_), .A2(new_n852_), .ZN(new_n932_));
  AOI21_X1   g00739(.A1(new_n931_), .A2(new_n920_), .B(new_n932_), .ZN(new_n933_));
  AOI21_X1   g00740(.A1(new_n930_), .A2(new_n927_), .B(new_n933_), .ZN(new_n934_));
  AOI22_X1   g00741(.A1(new_n934_), .A2(new_n924_), .B1(new_n866_), .B2(new_n926_), .ZN(\asquared[19] ));
  OAI21_X1   g00742(.A1(new_n865_), .A2(new_n858_), .B(new_n925_), .ZN(new_n936_));
  NAND2_X1   g00743(.A1(new_n936_), .A2(new_n924_), .ZN(new_n937_));
  NOR2_X1    g00744(.A1(new_n912_), .A2(new_n889_), .ZN(new_n938_));
  AND2_X2    g00745(.A1(new_n912_), .A2(new_n889_), .Z(new_n939_));
  NOR2_X1    g00746(.A1(new_n939_), .A2(new_n938_), .ZN(new_n940_));
  NAND2_X1   g00747(.A1(\a[3] ), .A2(\a[16] ), .ZN(new_n941_));
  NOR2_X1    g00748(.A1(new_n355_), .A2(new_n513_), .ZN(new_n942_));
  NOR2_X1    g00749(.A1(new_n942_), .A2(new_n540_), .ZN(new_n943_));
  NAND2_X1   g00750(.A1(new_n942_), .A2(new_n540_), .ZN(new_n944_));
  INV_X1     g00751(.I(new_n944_), .ZN(new_n945_));
  NOR3_X1    g00752(.A1(new_n945_), .A2(new_n941_), .A3(new_n943_), .ZN(new_n946_));
  OAI21_X1   g00753(.A1(new_n941_), .A2(new_n943_), .B(new_n944_), .ZN(new_n947_));
  OAI22_X1   g00754(.A1(new_n946_), .A2(new_n941_), .B1(new_n943_), .B2(new_n947_), .ZN(new_n948_));
  XNOR2_X1   g00755(.A1(new_n940_), .A2(new_n948_), .ZN(new_n949_));
  INV_X1     g00756(.I(new_n949_), .ZN(new_n950_));
  NAND2_X1   g00757(.A1(new_n891_), .A2(new_n904_), .ZN(new_n951_));
  NAND2_X1   g00758(.A1(new_n905_), .A2(new_n913_), .ZN(new_n952_));
  NAND2_X1   g00759(.A1(new_n952_), .A2(new_n951_), .ZN(new_n953_));
  NOR2_X1    g00760(.A1(new_n413_), .A2(new_n907_), .ZN(new_n954_));
  NAND2_X1   g00761(.A1(\a[1] ), .A2(\a[18] ), .ZN(new_n955_));
  NAND2_X1   g00762(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  XOR2_X1    g00763(.A1(new_n955_), .A2(new_n417_), .Z(new_n957_));
  OAI21_X1   g00764(.A1(new_n957_), .A2(new_n954_), .B(new_n956_), .ZN(new_n958_));
  XNOR2_X1   g00765(.A1(new_n958_), .A2(new_n903_), .ZN(new_n959_));
  XOR2_X1    g00766(.A1(new_n953_), .A2(new_n959_), .Z(new_n960_));
  NAND2_X1   g00767(.A1(new_n960_), .A2(new_n950_), .ZN(new_n961_));
  OR2_X2     g00768(.A1(new_n960_), .A2(new_n950_), .Z(new_n962_));
  NAND2_X1   g00769(.A1(new_n962_), .A2(new_n961_), .ZN(new_n963_));
  NAND2_X1   g00770(.A1(new_n878_), .A2(new_n877_), .ZN(new_n964_));
  INV_X1     g00771(.I(new_n826_), .ZN(new_n965_));
  NOR2_X1    g00772(.A1(new_n841_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1    g00773(.A1(new_n867_), .A2(new_n819_), .ZN(new_n967_));
  NOR2_X1    g00774(.A1(new_n967_), .A2(new_n966_), .ZN(new_n968_));
  INV_X1     g00775(.I(new_n373_), .ZN(new_n969_));
  NAND2_X1   g00776(.A1(new_n969_), .A2(new_n762_), .ZN(new_n970_));
  NAND2_X1   g00777(.A1(new_n760_), .A2(new_n746_), .ZN(new_n971_));
  AOI22_X1   g00778(.A1(new_n970_), .A2(new_n971_), .B1(new_n479_), .B2(new_n763_), .ZN(new_n972_));
  NOR2_X1    g00779(.A1(new_n253_), .A2(new_n759_), .ZN(new_n973_));
  INV_X1     g00780(.I(new_n973_), .ZN(new_n974_));
  AOI22_X1   g00781(.A1(\a[6] ), .A2(\a[13] ), .B1(\a[7] ), .B2(\a[12] ), .ZN(new_n975_));
  NAND2_X1   g00782(.A1(new_n763_), .A2(new_n479_), .ZN(new_n976_));
  NAND3_X1   g00783(.A1(new_n976_), .A2(new_n970_), .A3(new_n971_), .ZN(new_n977_));
  OAI22_X1   g00784(.A1(new_n972_), .A2(new_n974_), .B1(new_n977_), .B2(new_n975_), .ZN(new_n978_));
  INV_X1     g00785(.I(\a[19] ), .ZN(new_n979_));
  INV_X1     g00786(.I(new_n595_), .ZN(new_n980_));
  AOI22_X1   g00787(.A1(\a[15] ), .A2(new_n980_), .B1(new_n533_), .B2(\a[17] ), .ZN(new_n981_));
  NAND2_X1   g00788(.A1(\a[15] ), .A2(\a[17] ), .ZN(new_n982_));
  NOR2_X1    g00789(.A1(new_n251_), .A2(new_n982_), .ZN(new_n983_));
  NOR3_X1    g00790(.A1(new_n981_), .A2(new_n979_), .A3(new_n983_), .ZN(new_n984_));
  NOR3_X1    g00791(.A1(new_n984_), .A2(new_n196_), .A3(new_n979_), .ZN(new_n985_));
  OAI22_X1   g00792(.A1(new_n981_), .A2(new_n979_), .B1(new_n251_), .B2(new_n982_), .ZN(new_n986_));
  AOI22_X1   g00793(.A1(\a[2] ), .A2(\a[17] ), .B1(\a[4] ), .B2(\a[15] ), .ZN(new_n987_));
  NOR2_X1    g00794(.A1(new_n986_), .A2(new_n987_), .ZN(new_n988_));
  NOR2_X1    g00795(.A1(new_n988_), .A2(new_n985_), .ZN(new_n989_));
  XOR2_X1    g00796(.A1(new_n989_), .A2(new_n978_), .Z(new_n990_));
  NOR2_X1    g00797(.A1(new_n968_), .A2(new_n990_), .ZN(new_n991_));
  INV_X1     g00798(.I(new_n991_), .ZN(new_n992_));
  NAND2_X1   g00799(.A1(new_n968_), .A2(new_n990_), .ZN(new_n993_));
  NAND2_X1   g00800(.A1(new_n992_), .A2(new_n993_), .ZN(new_n994_));
  INV_X1     g00801(.I(new_n994_), .ZN(new_n995_));
  NOR2_X1    g00802(.A1(new_n964_), .A2(new_n995_), .ZN(new_n996_));
  NAND2_X1   g00803(.A1(new_n964_), .A2(new_n995_), .ZN(new_n997_));
  INV_X1     g00804(.I(new_n997_), .ZN(new_n998_));
  NOR2_X1    g00805(.A1(new_n998_), .A2(new_n996_), .ZN(new_n999_));
  INV_X1     g00806(.I(new_n999_), .ZN(new_n1000_));
  NOR2_X1    g00807(.A1(new_n1000_), .A2(new_n963_), .ZN(new_n1001_));
  NAND2_X1   g00808(.A1(new_n1000_), .A2(new_n963_), .ZN(new_n1002_));
  INV_X1     g00809(.I(new_n1002_), .ZN(new_n1003_));
  NOR2_X1    g00810(.A1(new_n917_), .A2(new_n914_), .ZN(new_n1004_));
  NOR2_X1    g00811(.A1(new_n919_), .A2(new_n1004_), .ZN(new_n1005_));
  NOR3_X1    g00812(.A1(new_n1003_), .A2(new_n1001_), .A3(new_n1005_), .ZN(new_n1006_));
  INV_X1     g00813(.I(new_n1001_), .ZN(new_n1007_));
  INV_X1     g00814(.I(new_n1005_), .ZN(new_n1008_));
  AOI21_X1   g00815(.A1(new_n1007_), .A2(new_n1002_), .B(new_n1008_), .ZN(new_n1009_));
  NOR2_X1    g00816(.A1(new_n1009_), .A2(new_n1006_), .ZN(new_n1010_));
  XOR2_X1    g00817(.A1(new_n937_), .A2(new_n1010_), .Z(\asquared[20] ));
  INV_X1     g00818(.I(new_n1006_), .ZN(new_n1012_));
  OAI21_X1   g00819(.A1(new_n1003_), .A2(new_n1001_), .B(new_n1005_), .ZN(new_n1013_));
  OAI21_X1   g00820(.A1(new_n934_), .A2(new_n923_), .B(new_n1013_), .ZN(new_n1014_));
  NAND2_X1   g00821(.A1(new_n1014_), .A2(new_n1012_), .ZN(new_n1015_));
  NAND2_X1   g00822(.A1(new_n953_), .A2(new_n959_), .ZN(new_n1016_));
  NAND2_X1   g00823(.A1(new_n961_), .A2(new_n1016_), .ZN(new_n1017_));
  INV_X1     g00824(.I(new_n939_), .ZN(new_n1018_));
  NAND2_X1   g00825(.A1(new_n940_), .A2(new_n948_), .ZN(new_n1019_));
  NAND2_X1   g00826(.A1(new_n1019_), .A2(new_n1018_), .ZN(new_n1020_));
  INV_X1     g00827(.I(new_n903_), .ZN(new_n1021_));
  OAI21_X1   g00828(.A1(new_n1021_), .A2(new_n958_), .B(new_n956_), .ZN(new_n1022_));
  INV_X1     g00829(.I(\a[17] ), .ZN(new_n1023_));
  NOR2_X1    g00830(.A1(new_n742_), .A2(new_n1023_), .ZN(new_n1024_));
  NOR2_X1    g00831(.A1(new_n742_), .A2(new_n884_), .ZN(new_n1025_));
  NAND2_X1   g00832(.A1(new_n1025_), .A2(new_n252_), .ZN(new_n1026_));
  NOR2_X1    g00833(.A1(new_n1023_), .A2(new_n884_), .ZN(new_n1027_));
  NAND2_X1   g00834(.A1(new_n1027_), .A2(new_n256_), .ZN(new_n1028_));
  AOI22_X1   g00835(.A1(new_n1026_), .A2(new_n1028_), .B1(new_n761_), .B2(new_n1024_), .ZN(new_n1029_));
  NAND2_X1   g00836(.A1(\a[2] ), .A2(\a[18] ), .ZN(new_n1030_));
  AOI22_X1   g00837(.A1(\a[3] ), .A2(\a[17] ), .B1(\a[4] ), .B2(\a[16] ), .ZN(new_n1031_));
  NAND2_X1   g00838(.A1(new_n1024_), .A2(new_n761_), .ZN(new_n1032_));
  NAND3_X1   g00839(.A1(new_n1032_), .A2(new_n1026_), .A3(new_n1028_), .ZN(new_n1033_));
  OAI22_X1   g00840(.A1(new_n1029_), .A2(new_n1030_), .B1(new_n1033_), .B2(new_n1031_), .ZN(new_n1034_));
  XOR2_X1    g00841(.A1(new_n1022_), .A2(new_n1034_), .Z(new_n1035_));
  XOR2_X1    g00842(.A1(new_n1020_), .A2(new_n1035_), .Z(new_n1036_));
  NOR2_X1    g00843(.A1(new_n1017_), .A2(new_n1036_), .ZN(new_n1037_));
  NAND2_X1   g00844(.A1(new_n1017_), .A2(new_n1036_), .ZN(new_n1038_));
  INV_X1     g00845(.I(new_n1038_), .ZN(new_n1039_));
  NOR2_X1    g00846(.A1(new_n1039_), .A2(new_n1037_), .ZN(new_n1040_));
  NOR2_X1    g00847(.A1(new_n955_), .A2(new_n417_), .ZN(new_n1041_));
  AOI22_X1   g00848(.A1(\a[0] ), .A2(\a[20] ), .B1(\a[7] ), .B2(\a[13] ), .ZN(new_n1042_));
  INV_X1     g00849(.I(\a[20] ), .ZN(new_n1043_));
  NOR4_X1    g00850(.A1(new_n196_), .A2(new_n422_), .A3(new_n597_), .A4(new_n1043_), .ZN(new_n1044_));
  NOR2_X1    g00851(.A1(new_n1044_), .A2(new_n1042_), .ZN(new_n1045_));
  XOR2_X1    g00852(.A1(new_n1045_), .A2(new_n1041_), .Z(new_n1046_));
  XOR2_X1    g00853(.A1(new_n1046_), .A2(new_n977_), .Z(new_n1047_));
  NAND2_X1   g00854(.A1(new_n645_), .A2(new_n762_), .ZN(new_n1048_));
  NAND4_X1   g00855(.A1(\a[5] ), .A2(\a[8] ), .A3(\a[12] ), .A4(\a[15] ), .ZN(new_n1049_));
  AOI22_X1   g00856(.A1(new_n1048_), .A2(new_n1049_), .B1(new_n746_), .B2(new_n897_), .ZN(new_n1050_));
  NAND2_X1   g00857(.A1(new_n897_), .A2(new_n746_), .ZN(new_n1051_));
  NAND3_X1   g00858(.A1(new_n1051_), .A2(new_n1048_), .A3(new_n1049_), .ZN(new_n1052_));
  NOR2_X1    g00859(.A1(new_n367_), .A2(new_n759_), .ZN(new_n1053_));
  NOR2_X1    g00860(.A1(new_n253_), .A2(new_n717_), .ZN(new_n1054_));
  NOR2_X1    g00861(.A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_));
  NAND2_X1   g00862(.A1(\a[8] ), .A2(\a[12] ), .ZN(new_n1056_));
  OAI22_X1   g00863(.A1(new_n1050_), .A2(new_n1056_), .B1(new_n1052_), .B2(new_n1055_), .ZN(new_n1057_));
  XNOR2_X1   g00864(.A1(new_n1047_), .A2(new_n1057_), .ZN(new_n1058_));
  OAI21_X1   g00865(.A1(new_n985_), .A2(new_n988_), .B(new_n978_), .ZN(new_n1059_));
  NOR2_X1    g00866(.A1(new_n403_), .A2(new_n513_), .ZN(new_n1060_));
  NOR2_X1    g00867(.A1(new_n194_), .A2(new_n979_), .ZN(new_n1061_));
  NAND2_X1   g00868(.A1(new_n1060_), .A2(new_n1061_), .ZN(new_n1062_));
  INV_X1     g00869(.I(new_n1060_), .ZN(new_n1063_));
  INV_X1     g00870(.I(new_n1061_), .ZN(new_n1064_));
  NAND2_X1   g00871(.A1(new_n1063_), .A2(new_n1064_), .ZN(new_n1065_));
  NAND2_X1   g00872(.A1(new_n1065_), .A2(new_n1062_), .ZN(new_n1066_));
  XOR2_X1    g00873(.A1(new_n1066_), .A2(new_n947_), .Z(new_n1067_));
  XOR2_X1    g00874(.A1(new_n1067_), .A2(new_n986_), .Z(new_n1068_));
  NAND3_X1   g00875(.A1(new_n992_), .A2(new_n1059_), .A3(new_n1068_), .ZN(new_n1069_));
  INV_X1     g00876(.I(new_n1059_), .ZN(new_n1070_));
  INV_X1     g00877(.I(new_n1068_), .ZN(new_n1071_));
  OAI21_X1   g00878(.A1(new_n991_), .A2(new_n1070_), .B(new_n1071_), .ZN(new_n1072_));
  NAND2_X1   g00879(.A1(new_n1069_), .A2(new_n1072_), .ZN(new_n1073_));
  XOR2_X1    g00880(.A1(new_n1073_), .A2(new_n1058_), .Z(new_n1074_));
  XOR2_X1    g00881(.A1(new_n1040_), .A2(new_n1074_), .Z(new_n1075_));
  NOR2_X1    g00882(.A1(new_n1001_), .A2(new_n998_), .ZN(new_n1076_));
  INV_X1     g00883(.I(new_n1076_), .ZN(new_n1077_));
  NOR2_X1    g00884(.A1(new_n1077_), .A2(new_n1075_), .ZN(new_n1078_));
  INV_X1     g00885(.I(new_n1075_), .ZN(new_n1079_));
  NOR2_X1    g00886(.A1(new_n1079_), .A2(new_n1076_), .ZN(new_n1080_));
  NOR2_X1    g00887(.A1(new_n1080_), .A2(new_n1078_), .ZN(new_n1081_));
  XOR2_X1    g00888(.A1(new_n1015_), .A2(new_n1081_), .Z(\asquared[21] ));
  INV_X1     g00889(.I(new_n1080_), .ZN(new_n1083_));
  AOI21_X1   g00890(.A1(new_n936_), .A2(new_n924_), .B(new_n1009_), .ZN(new_n1084_));
  NAND2_X1   g00891(.A1(new_n1079_), .A2(new_n1076_), .ZN(new_n1085_));
  OAI21_X1   g00892(.A1(new_n1084_), .A2(new_n1006_), .B(new_n1085_), .ZN(new_n1086_));
  NAND2_X1   g00893(.A1(new_n1086_), .A2(new_n1083_), .ZN(new_n1087_));
  AND2_X2    g00894(.A1(new_n1040_), .A2(new_n1074_), .Z(new_n1088_));
  NOR2_X1    g00895(.A1(new_n1088_), .A2(new_n1039_), .ZN(new_n1089_));
  INV_X1     g00896(.I(new_n1089_), .ZN(new_n1090_));
  AOI22_X1   g00897(.A1(\a[3] ), .A2(new_n1025_), .B1(new_n900_), .B2(\a[19] ), .ZN(new_n1091_));
  NAND2_X1   g00898(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n1092_));
  NOR2_X1    g00899(.A1(new_n246_), .A2(new_n1092_), .ZN(new_n1093_));
  NOR3_X1    g00900(.A1(new_n1091_), .A2(new_n253_), .A3(new_n1093_), .ZN(new_n1094_));
  NAND2_X1   g00901(.A1(\a[5] ), .A2(\a[16] ), .ZN(new_n1095_));
  NOR2_X1    g00902(.A1(new_n1094_), .A2(new_n1093_), .ZN(new_n1096_));
  INV_X1     g00903(.I(new_n1096_), .ZN(new_n1097_));
  AOI22_X1   g00904(.A1(\a[2] ), .A2(\a[19] ), .B1(\a[3] ), .B2(\a[18] ), .ZN(new_n1098_));
  OAI22_X1   g00905(.A1(new_n1097_), .A2(new_n1098_), .B1(new_n1094_), .B2(new_n1095_), .ZN(new_n1099_));
  NOR2_X1    g00906(.A1(new_n767_), .A2(new_n415_), .ZN(new_n1100_));
  INV_X1     g00907(.I(new_n836_), .ZN(new_n1101_));
  AOI22_X1   g00908(.A1(new_n479_), .A2(new_n897_), .B1(new_n645_), .B2(new_n1101_), .ZN(new_n1102_));
  NOR2_X1    g00909(.A1(new_n1100_), .A2(new_n1102_), .ZN(new_n1103_));
  NAND2_X1   g00910(.A1(\a[6] ), .A2(\a[15] ), .ZN(new_n1104_));
  AOI22_X1   g00911(.A1(\a[7] ), .A2(\a[14] ), .B1(\a[8] ), .B2(\a[13] ), .ZN(new_n1105_));
  OAI21_X1   g00912(.A1(new_n415_), .A2(new_n767_), .B(new_n1102_), .ZN(new_n1106_));
  OAI22_X1   g00913(.A1(new_n1106_), .A2(new_n1105_), .B1(new_n1103_), .B2(new_n1104_), .ZN(new_n1107_));
  XOR2_X1    g00914(.A1(new_n1099_), .A2(new_n1107_), .Z(new_n1108_));
  AOI21_X1   g00915(.A1(\a[9] ), .A2(\a[12] ), .B(new_n747_), .ZN(new_n1109_));
  NOR2_X1    g00916(.A1(new_n290_), .A2(new_n1023_), .ZN(new_n1110_));
  INV_X1     g00917(.I(new_n1110_), .ZN(new_n1111_));
  OAI22_X1   g00918(.A1(new_n1109_), .A2(new_n1111_), .B1(new_n539_), .B2(new_n619_), .ZN(new_n1112_));
  NOR2_X1    g00919(.A1(new_n539_), .A2(new_n619_), .ZN(new_n1113_));
  OAI21_X1   g00920(.A1(new_n1109_), .A2(new_n1113_), .B(new_n1110_), .ZN(new_n1114_));
  OAI21_X1   g00921(.A1(new_n1112_), .A2(new_n1109_), .B(new_n1114_), .ZN(new_n1115_));
  XOR2_X1    g00922(.A1(new_n1108_), .A2(new_n1115_), .Z(new_n1116_));
  INV_X1     g00923(.I(new_n1116_), .ZN(new_n1117_));
  NAND2_X1   g00924(.A1(new_n1022_), .A2(new_n1034_), .ZN(new_n1118_));
  NAND2_X1   g00925(.A1(new_n1020_), .A2(new_n1035_), .ZN(new_n1119_));
  NAND2_X1   g00926(.A1(new_n1119_), .A2(new_n1118_), .ZN(new_n1120_));
  INV_X1     g00927(.I(new_n1044_), .ZN(new_n1121_));
  NAND2_X1   g00928(.A1(new_n1045_), .A2(new_n1041_), .ZN(new_n1122_));
  NAND2_X1   g00929(.A1(new_n1122_), .A2(new_n1121_), .ZN(new_n1123_));
  XOR2_X1    g00930(.A1(new_n1033_), .A2(new_n1052_), .Z(new_n1124_));
  XOR2_X1    g00931(.A1(new_n1124_), .A2(new_n1123_), .Z(new_n1125_));
  XNOR2_X1   g00932(.A1(new_n1120_), .A2(new_n1125_), .ZN(new_n1126_));
  OR2_X2     g00933(.A1(new_n1126_), .A2(new_n1117_), .Z(new_n1127_));
  NAND2_X1   g00934(.A1(new_n1126_), .A2(new_n1117_), .ZN(new_n1128_));
  NAND2_X1   g00935(.A1(new_n1127_), .A2(new_n1128_), .ZN(new_n1129_));
  NAND2_X1   g00936(.A1(new_n1046_), .A2(new_n977_), .ZN(new_n1130_));
  NAND2_X1   g00937(.A1(new_n1047_), .A2(new_n1057_), .ZN(new_n1131_));
  NAND3_X1   g00938(.A1(new_n947_), .A2(new_n1062_), .A3(new_n1065_), .ZN(new_n1132_));
  INV_X1     g00939(.I(new_n1132_), .ZN(new_n1133_));
  INV_X1     g00940(.I(new_n986_), .ZN(new_n1134_));
  NOR2_X1    g00941(.A1(new_n1067_), .A2(new_n1134_), .ZN(new_n1135_));
  NOR2_X1    g00942(.A1(new_n1135_), .A2(new_n1133_), .ZN(new_n1136_));
  NAND2_X1   g00943(.A1(\a[1] ), .A2(\a[20] ), .ZN(new_n1137_));
  XOR2_X1    g00944(.A1(new_n1137_), .A2(\a[11] ), .Z(new_n1138_));
  NAND2_X1   g00945(.A1(\a[0] ), .A2(\a[21] ), .ZN(new_n1139_));
  INV_X1     g00946(.I(new_n1139_), .ZN(new_n1140_));
  XOR2_X1    g00947(.A1(new_n1062_), .A2(new_n1140_), .Z(new_n1141_));
  NOR2_X1    g00948(.A1(new_n1141_), .A2(new_n1138_), .ZN(new_n1142_));
  INV_X1     g00949(.I(new_n1142_), .ZN(new_n1143_));
  NAND2_X1   g00950(.A1(new_n1141_), .A2(new_n1138_), .ZN(new_n1144_));
  NAND2_X1   g00951(.A1(new_n1143_), .A2(new_n1144_), .ZN(new_n1145_));
  NAND2_X1   g00952(.A1(new_n1136_), .A2(new_n1145_), .ZN(new_n1146_));
  INV_X1     g00953(.I(new_n1145_), .ZN(new_n1147_));
  OAI21_X1   g00954(.A1(new_n1133_), .A2(new_n1135_), .B(new_n1147_), .ZN(new_n1148_));
  NAND2_X1   g00955(.A1(new_n1148_), .A2(new_n1146_), .ZN(new_n1149_));
  NAND3_X1   g00956(.A1(new_n1149_), .A2(new_n1130_), .A3(new_n1131_), .ZN(new_n1150_));
  NAND2_X1   g00957(.A1(new_n1131_), .A2(new_n1130_), .ZN(new_n1151_));
  NAND3_X1   g00958(.A1(new_n1151_), .A2(new_n1148_), .A3(new_n1146_), .ZN(new_n1152_));
  NAND2_X1   g00959(.A1(new_n1150_), .A2(new_n1152_), .ZN(new_n1153_));
  INV_X1     g00960(.I(new_n1153_), .ZN(new_n1154_));
  OAI21_X1   g00961(.A1(new_n1073_), .A2(new_n1058_), .B(new_n1072_), .ZN(new_n1155_));
  NAND2_X1   g00962(.A1(new_n1155_), .A2(new_n1154_), .ZN(new_n1156_));
  INV_X1     g00963(.I(new_n1156_), .ZN(new_n1157_));
  NOR2_X1    g00964(.A1(new_n1155_), .A2(new_n1154_), .ZN(new_n1158_));
  NOR2_X1    g00965(.A1(new_n1157_), .A2(new_n1158_), .ZN(new_n1159_));
  INV_X1     g00966(.I(new_n1159_), .ZN(new_n1160_));
  NAND2_X1   g00967(.A1(new_n1160_), .A2(new_n1129_), .ZN(new_n1161_));
  NAND3_X1   g00968(.A1(new_n1159_), .A2(new_n1127_), .A3(new_n1128_), .ZN(new_n1162_));
  AND2_X2    g00969(.A1(new_n1161_), .A2(new_n1162_), .Z(new_n1163_));
  NOR2_X1    g00970(.A1(new_n1163_), .A2(new_n1090_), .ZN(new_n1164_));
  NAND2_X1   g00971(.A1(new_n1163_), .A2(new_n1090_), .ZN(new_n1165_));
  INV_X1     g00972(.I(new_n1165_), .ZN(new_n1166_));
  NOR2_X1    g00973(.A1(new_n1166_), .A2(new_n1164_), .ZN(new_n1167_));
  XOR2_X1    g00974(.A1(new_n1087_), .A2(new_n1167_), .Z(\asquared[22] ));
  AOI21_X1   g00975(.A1(new_n1086_), .A2(new_n1083_), .B(new_n1164_), .ZN(new_n1169_));
  NOR2_X1    g00976(.A1(new_n1169_), .A2(new_n1166_), .ZN(new_n1170_));
  AOI22_X1   g00977(.A1(\a[7] ), .A2(\a[15] ), .B1(\a[8] ), .B2(\a[14] ), .ZN(new_n1171_));
  INV_X1     g00978(.I(new_n1171_), .ZN(new_n1172_));
  INV_X1     g00979(.I(new_n897_), .ZN(new_n1173_));
  NOR2_X1    g00980(.A1(new_n1173_), .A2(new_n415_), .ZN(new_n1174_));
  INV_X1     g00981(.I(\a[22] ), .ZN(new_n1175_));
  NOR2_X1    g00982(.A1(new_n196_), .A2(new_n1175_), .ZN(new_n1176_));
  AOI21_X1   g00983(.A1(new_n1172_), .A2(new_n1176_), .B(new_n1174_), .ZN(new_n1177_));
  NAND2_X1   g00984(.A1(new_n1177_), .A2(new_n1172_), .ZN(new_n1178_));
  OAI21_X1   g00985(.A1(new_n1174_), .A2(new_n1171_), .B(new_n1176_), .ZN(new_n1179_));
  NAND2_X1   g00986(.A1(new_n1178_), .A2(new_n1179_), .ZN(new_n1180_));
  INV_X1     g00987(.I(new_n743_), .ZN(new_n1181_));
  OAI21_X1   g00988(.A1(new_n197_), .A2(new_n1043_), .B(new_n1181_), .ZN(new_n1182_));
  INV_X1     g00989(.I(new_n1182_), .ZN(new_n1183_));
  INV_X1     g00990(.I(new_n596_), .ZN(new_n1184_));
  NOR3_X1    g00991(.A1(new_n1181_), .A2(new_n197_), .A3(new_n1043_), .ZN(new_n1185_));
  AOI21_X1   g00992(.A1(new_n1182_), .A2(new_n1184_), .B(new_n1185_), .ZN(new_n1186_));
  INV_X1     g00993(.I(new_n1186_), .ZN(new_n1187_));
  OAI21_X1   g00994(.A1(new_n1183_), .A2(new_n1185_), .B(new_n1184_), .ZN(new_n1188_));
  OAI21_X1   g00995(.A1(new_n1183_), .A2(new_n1187_), .B(new_n1188_), .ZN(new_n1189_));
  XOR2_X1    g00996(.A1(new_n1189_), .A2(new_n1180_), .Z(new_n1190_));
  NOR2_X1    g00997(.A1(new_n225_), .A2(new_n979_), .ZN(new_n1191_));
  INV_X1     g00998(.I(new_n1191_), .ZN(new_n1192_));
  NAND3_X1   g00999(.A1(new_n1191_), .A2(\a[5] ), .A3(\a[17] ), .ZN(new_n1193_));
  INV_X1     g01000(.I(new_n1092_), .ZN(new_n1194_));
  NAND2_X1   g01001(.A1(new_n761_), .A2(new_n1194_), .ZN(new_n1195_));
  AOI22_X1   g01002(.A1(new_n1193_), .A2(new_n1195_), .B1(new_n243_), .B2(new_n1027_), .ZN(new_n1196_));
  AOI22_X1   g01003(.A1(\a[4] ), .A2(\a[18] ), .B1(\a[5] ), .B2(\a[17] ), .ZN(new_n1197_));
  NAND2_X1   g01004(.A1(new_n1027_), .A2(new_n243_), .ZN(new_n1198_));
  NAND3_X1   g01005(.A1(new_n1198_), .A2(new_n1193_), .A3(new_n1195_), .ZN(new_n1199_));
  OAI22_X1   g01006(.A1(new_n1196_), .A2(new_n1192_), .B1(new_n1199_), .B2(new_n1197_), .ZN(new_n1200_));
  XNOR2_X1   g01007(.A1(new_n1190_), .A2(new_n1200_), .ZN(new_n1201_));
  INV_X1     g01008(.I(new_n1201_), .ZN(new_n1202_));
  NAND2_X1   g01009(.A1(new_n1152_), .A2(new_n1148_), .ZN(new_n1203_));
  NOR2_X1    g01010(.A1(new_n1062_), .A2(new_n1139_), .ZN(new_n1204_));
  NOR2_X1    g01011(.A1(new_n1142_), .A2(new_n1204_), .ZN(new_n1205_));
  NOR2_X1    g01012(.A1(new_n1097_), .A2(new_n1106_), .ZN(new_n1206_));
  NAND2_X1   g01013(.A1(new_n1097_), .A2(new_n1106_), .ZN(new_n1207_));
  INV_X1     g01014(.I(new_n1207_), .ZN(new_n1208_));
  NOR2_X1    g01015(.A1(new_n1208_), .A2(new_n1206_), .ZN(new_n1209_));
  XNOR2_X1   g01016(.A1(new_n1209_), .A2(new_n1205_), .ZN(new_n1210_));
  XOR2_X1    g01017(.A1(new_n1203_), .A2(new_n1210_), .Z(new_n1211_));
  XOR2_X1    g01018(.A1(new_n1211_), .A2(new_n1202_), .Z(new_n1212_));
  NAND2_X1   g01019(.A1(new_n1099_), .A2(new_n1107_), .ZN(new_n1213_));
  NAND2_X1   g01020(.A1(new_n1108_), .A2(new_n1115_), .ZN(new_n1214_));
  NAND2_X1   g01021(.A1(new_n1214_), .A2(new_n1213_), .ZN(new_n1215_));
  NAND2_X1   g01022(.A1(new_n1033_), .A2(new_n1052_), .ZN(new_n1216_));
  NAND2_X1   g01023(.A1(new_n1124_), .A2(new_n1123_), .ZN(new_n1217_));
  NAND2_X1   g01024(.A1(new_n1217_), .A2(new_n1216_), .ZN(new_n1218_));
  NOR2_X1    g01025(.A1(new_n1137_), .A2(new_n513_), .ZN(new_n1219_));
  INV_X1     g01026(.I(\a[21] ), .ZN(new_n1220_));
  NOR2_X1    g01027(.A1(new_n194_), .A2(new_n1220_), .ZN(new_n1221_));
  NAND2_X1   g01028(.A1(new_n1221_), .A2(new_n535_), .ZN(new_n1222_));
  NOR2_X1    g01029(.A1(new_n1221_), .A2(new_n535_), .ZN(new_n1223_));
  INV_X1     g01030(.I(new_n1223_), .ZN(new_n1224_));
  NAND2_X1   g01031(.A1(new_n1224_), .A2(new_n1222_), .ZN(new_n1225_));
  XNOR2_X1   g01032(.A1(new_n1225_), .A2(new_n1219_), .ZN(new_n1226_));
  XOR2_X1    g01033(.A1(new_n1226_), .A2(new_n1112_), .Z(new_n1227_));
  XOR2_X1    g01034(.A1(new_n1227_), .A2(new_n1218_), .Z(new_n1228_));
  XOR2_X1    g01035(.A1(new_n1228_), .A2(new_n1215_), .Z(new_n1229_));
  NAND2_X1   g01036(.A1(new_n1120_), .A2(new_n1125_), .ZN(new_n1230_));
  NAND2_X1   g01037(.A1(new_n1127_), .A2(new_n1230_), .ZN(new_n1231_));
  NAND2_X1   g01038(.A1(new_n1231_), .A2(new_n1229_), .ZN(new_n1232_));
  NAND2_X1   g01039(.A1(new_n1232_), .A2(new_n1229_), .ZN(new_n1233_));
  NAND2_X1   g01040(.A1(new_n1232_), .A2(new_n1231_), .ZN(new_n1234_));
  NAND2_X1   g01041(.A1(new_n1234_), .A2(new_n1233_), .ZN(new_n1235_));
  AOI21_X1   g01042(.A1(new_n1232_), .A2(new_n1231_), .B(new_n1212_), .ZN(new_n1236_));
  AOI22_X1   g01043(.A1(new_n1235_), .A2(new_n1212_), .B1(new_n1236_), .B2(new_n1233_), .ZN(new_n1237_));
  INV_X1     g01044(.I(new_n1237_), .ZN(new_n1238_));
  NAND2_X1   g01045(.A1(new_n1162_), .A2(new_n1156_), .ZN(new_n1239_));
  INV_X1     g01046(.I(new_n1239_), .ZN(new_n1240_));
  NOR2_X1    g01047(.A1(new_n1238_), .A2(new_n1240_), .ZN(new_n1241_));
  INV_X1     g01048(.I(new_n1241_), .ZN(new_n1242_));
  NOR2_X1    g01049(.A1(new_n1237_), .A2(new_n1239_), .ZN(new_n1243_));
  INV_X1     g01050(.I(new_n1243_), .ZN(new_n1244_));
  NAND2_X1   g01051(.A1(new_n1242_), .A2(new_n1244_), .ZN(new_n1245_));
  AOI21_X1   g01052(.A1(new_n1014_), .A2(new_n1012_), .B(new_n1078_), .ZN(new_n1246_));
  INV_X1     g01053(.I(new_n1164_), .ZN(new_n1247_));
  OAI21_X1   g01054(.A1(new_n1246_), .A2(new_n1080_), .B(new_n1247_), .ZN(new_n1248_));
  AOI21_X1   g01055(.A1(new_n1248_), .A2(new_n1165_), .B(new_n1243_), .ZN(new_n1249_));
  AOI22_X1   g01056(.A1(new_n1249_), .A2(new_n1242_), .B1(new_n1170_), .B2(new_n1245_), .ZN(\asquared[23] ));
  OAI21_X1   g01057(.A1(new_n1169_), .A2(new_n1166_), .B(new_n1244_), .ZN(new_n1251_));
  NAND2_X1   g01058(.A1(new_n1251_), .A2(new_n1242_), .ZN(new_n1252_));
  NAND2_X1   g01059(.A1(new_n1235_), .A2(new_n1212_), .ZN(new_n1253_));
  AND2_X2    g01060(.A1(new_n1253_), .A2(new_n1232_), .Z(new_n1254_));
  NAND2_X1   g01061(.A1(new_n1227_), .A2(new_n1218_), .ZN(new_n1255_));
  NAND2_X1   g01062(.A1(new_n1228_), .A2(new_n1215_), .ZN(new_n1256_));
  NAND2_X1   g01063(.A1(new_n1256_), .A2(new_n1255_), .ZN(new_n1257_));
  NAND3_X1   g01064(.A1(new_n1224_), .A2(new_n1219_), .A3(new_n1222_), .ZN(new_n1258_));
  NAND2_X1   g01065(.A1(new_n1226_), .A2(new_n1112_), .ZN(new_n1259_));
  NAND2_X1   g01066(.A1(new_n1259_), .A2(new_n1258_), .ZN(new_n1260_));
  INV_X1     g01067(.I(new_n619_), .ZN(new_n1261_));
  AOI21_X1   g01068(.A1(\a[10] ), .A2(\a[13] ), .B(new_n1261_), .ZN(new_n1262_));
  INV_X1     g01069(.I(new_n1262_), .ZN(new_n1263_));
  INV_X1     g01070(.I(new_n747_), .ZN(new_n1264_));
  INV_X1     g01071(.I(new_n763_), .ZN(new_n1265_));
  NOR2_X1    g01072(.A1(new_n1264_), .A2(new_n1265_), .ZN(new_n1266_));
  NOR2_X1    g01073(.A1(new_n290_), .A2(new_n979_), .ZN(new_n1267_));
  AOI21_X1   g01074(.A1(new_n1263_), .A2(new_n1267_), .B(new_n1266_), .ZN(new_n1268_));
  INV_X1     g01075(.I(new_n1268_), .ZN(new_n1269_));
  OAI21_X1   g01076(.A1(new_n1266_), .A2(new_n1262_), .B(new_n1267_), .ZN(new_n1270_));
  OAI21_X1   g01077(.A1(new_n1269_), .A2(new_n1262_), .B(new_n1270_), .ZN(new_n1271_));
  INV_X1     g01078(.I(new_n318_), .ZN(new_n1272_));
  NOR2_X1    g01079(.A1(new_n884_), .A2(new_n1043_), .ZN(new_n1273_));
  INV_X1     g01080(.I(new_n368_), .ZN(new_n1274_));
  INV_X1     g01081(.I(new_n1027_), .ZN(new_n1275_));
  NAND2_X1   g01082(.A1(\a[17] ), .A2(\a[20] ), .ZN(new_n1276_));
  OAI22_X1   g01083(.A1(new_n1275_), .A2(new_n371_), .B1(new_n1274_), .B2(new_n1276_), .ZN(new_n1277_));
  AOI21_X1   g01084(.A1(new_n1272_), .A2(new_n1273_), .B(new_n1277_), .ZN(new_n1278_));
  INV_X1     g01085(.I(new_n1278_), .ZN(new_n1279_));
  AOI22_X1   g01086(.A1(\a[3] ), .A2(\a[20] ), .B1(\a[5] ), .B2(\a[18] ), .ZN(new_n1280_));
  INV_X1     g01087(.I(new_n1273_), .ZN(new_n1281_));
  OAI21_X1   g01088(.A1(new_n318_), .A2(new_n1281_), .B(new_n1277_), .ZN(new_n1282_));
  NAND3_X1   g01089(.A1(new_n1282_), .A2(\a[6] ), .A3(\a[17] ), .ZN(new_n1283_));
  OAI21_X1   g01090(.A1(new_n1279_), .A2(new_n1280_), .B(new_n1283_), .ZN(new_n1284_));
  XOR2_X1    g01091(.A1(new_n1284_), .A2(new_n1271_), .Z(new_n1285_));
  XOR2_X1    g01092(.A1(new_n1285_), .A2(new_n1260_), .Z(new_n1286_));
  INV_X1     g01093(.I(new_n1286_), .ZN(new_n1287_));
  INV_X1     g01094(.I(new_n893_), .ZN(new_n1288_));
  NAND2_X1   g01095(.A1(new_n693_), .A2(new_n1288_), .ZN(new_n1289_));
  INV_X1     g01096(.I(new_n773_), .ZN(new_n1290_));
  NAND2_X1   g01097(.A1(new_n895_), .A2(new_n1290_), .ZN(new_n1291_));
  AOI22_X1   g01098(.A1(new_n1289_), .A2(new_n1291_), .B1(new_n467_), .B2(new_n897_), .ZN(new_n1292_));
  NAND2_X1   g01099(.A1(\a[7] ), .A2(\a[16] ), .ZN(new_n1293_));
  AOI22_X1   g01100(.A1(\a[8] ), .A2(\a[15] ), .B1(\a[9] ), .B2(\a[14] ), .ZN(new_n1294_));
  NAND2_X1   g01101(.A1(new_n467_), .A2(new_n897_), .ZN(new_n1295_));
  NAND3_X1   g01102(.A1(new_n1295_), .A2(new_n1289_), .A3(new_n1291_), .ZN(new_n1296_));
  OAI22_X1   g01103(.A1(new_n1292_), .A2(new_n1293_), .B1(new_n1296_), .B2(new_n1294_), .ZN(new_n1297_));
  AOI22_X1   g01104(.A1(\a[0] ), .A2(\a[23] ), .B1(\a[2] ), .B2(\a[21] ), .ZN(new_n1298_));
  INV_X1     g01105(.I(\a[23] ), .ZN(new_n1299_));
  NOR2_X1    g01106(.A1(new_n1220_), .A2(new_n1299_), .ZN(new_n1300_));
  INV_X1     g01107(.I(new_n1300_), .ZN(new_n1301_));
  NOR2_X1    g01108(.A1(new_n1301_), .A2(new_n412_), .ZN(new_n1302_));
  INV_X1     g01109(.I(new_n1302_), .ZN(new_n1303_));
  OAI21_X1   g01110(.A1(new_n1222_), .A2(new_n1298_), .B(new_n1303_), .ZN(new_n1304_));
  NOR2_X1    g01111(.A1(new_n1304_), .A2(new_n1298_), .ZN(new_n1305_));
  INV_X1     g01112(.I(new_n1298_), .ZN(new_n1306_));
  AOI21_X1   g01113(.A1(new_n1303_), .A2(new_n1306_), .B(new_n1222_), .ZN(new_n1307_));
  NOR2_X1    g01114(.A1(new_n1305_), .A2(new_n1307_), .ZN(new_n1308_));
  XOR2_X1    g01115(.A1(new_n1308_), .A2(new_n1177_), .Z(new_n1309_));
  XNOR2_X1   g01116(.A1(new_n1309_), .A2(new_n1297_), .ZN(new_n1310_));
  OR2_X2     g01117(.A1(new_n1287_), .A2(new_n1310_), .Z(new_n1311_));
  NAND2_X1   g01118(.A1(new_n1287_), .A2(new_n1310_), .ZN(new_n1312_));
  NAND2_X1   g01119(.A1(new_n1311_), .A2(new_n1312_), .ZN(new_n1313_));
  XOR2_X1    g01120(.A1(new_n1313_), .A2(new_n1257_), .Z(new_n1314_));
  NAND2_X1   g01121(.A1(new_n1203_), .A2(new_n1210_), .ZN(new_n1315_));
  NAND2_X1   g01122(.A1(new_n1211_), .A2(new_n1202_), .ZN(new_n1316_));
  NAND2_X1   g01123(.A1(new_n1316_), .A2(new_n1315_), .ZN(new_n1317_));
  NOR2_X1    g01124(.A1(new_n194_), .A2(new_n1175_), .ZN(new_n1318_));
  INV_X1     g01125(.I(new_n1318_), .ZN(new_n1319_));
  NOR2_X1    g01126(.A1(new_n1319_), .A2(new_n536_), .ZN(new_n1320_));
  NOR2_X1    g01127(.A1(new_n1318_), .A2(\a[12] ), .ZN(new_n1321_));
  NOR2_X1    g01128(.A1(new_n1320_), .A2(new_n1321_), .ZN(new_n1322_));
  XOR2_X1    g01129(.A1(new_n1322_), .A2(new_n1199_), .Z(new_n1323_));
  XOR2_X1    g01130(.A1(new_n1323_), .A2(new_n1187_), .Z(new_n1324_));
  INV_X1     g01131(.I(new_n1324_), .ZN(new_n1325_));
  OAI21_X1   g01132(.A1(new_n1205_), .A2(new_n1206_), .B(new_n1207_), .ZN(new_n1326_));
  NAND2_X1   g01133(.A1(new_n1189_), .A2(new_n1180_), .ZN(new_n1327_));
  NAND2_X1   g01134(.A1(new_n1190_), .A2(new_n1200_), .ZN(new_n1328_));
  NAND2_X1   g01135(.A1(new_n1328_), .A2(new_n1327_), .ZN(new_n1329_));
  XNOR2_X1   g01136(.A1(new_n1329_), .A2(new_n1326_), .ZN(new_n1330_));
  XOR2_X1    g01137(.A1(new_n1330_), .A2(new_n1325_), .Z(new_n1331_));
  XOR2_X1    g01138(.A1(new_n1317_), .A2(new_n1331_), .Z(new_n1332_));
  XOR2_X1    g01139(.A1(new_n1332_), .A2(new_n1314_), .Z(new_n1333_));
  NOR2_X1    g01140(.A1(new_n1254_), .A2(new_n1333_), .ZN(new_n1334_));
  NAND2_X1   g01141(.A1(new_n1254_), .A2(new_n1333_), .ZN(new_n1335_));
  INV_X1     g01142(.I(new_n1335_), .ZN(new_n1336_));
  NOR2_X1    g01143(.A1(new_n1336_), .A2(new_n1334_), .ZN(new_n1337_));
  XOR2_X1    g01144(.A1(new_n1252_), .A2(new_n1337_), .Z(\asquared[24] ));
  AOI21_X1   g01145(.A1(new_n1251_), .A2(new_n1242_), .B(new_n1336_), .ZN(new_n1339_));
  NOR2_X1    g01146(.A1(new_n1339_), .A2(new_n1334_), .ZN(new_n1340_));
  INV_X1     g01147(.I(new_n1314_), .ZN(new_n1341_));
  AND2_X2    g01148(.A1(new_n1317_), .A2(new_n1331_), .Z(new_n1342_));
  AOI21_X1   g01149(.A1(new_n1332_), .A2(new_n1341_), .B(new_n1342_), .ZN(new_n1343_));
  NAND2_X1   g01150(.A1(new_n1329_), .A2(new_n1326_), .ZN(new_n1344_));
  OAI21_X1   g01151(.A1(new_n1330_), .A2(new_n1325_), .B(new_n1344_), .ZN(new_n1345_));
  NAND2_X1   g01152(.A1(new_n1322_), .A2(new_n1199_), .ZN(new_n1346_));
  NAND2_X1   g01153(.A1(new_n1323_), .A2(new_n1187_), .ZN(new_n1347_));
  NAND2_X1   g01154(.A1(new_n1347_), .A2(new_n1346_), .ZN(new_n1348_));
  NAND2_X1   g01155(.A1(\a[7] ), .A2(\a[17] ), .ZN(new_n1349_));
  NOR4_X1    g01156(.A1(new_n197_), .A2(new_n367_), .A3(new_n884_), .A4(new_n1175_), .ZN(new_n1350_));
  NAND4_X1   g01157(.A1(\a[2] ), .A2(\a[7] ), .A3(\a[17] ), .A4(\a[22] ), .ZN(new_n1351_));
  NAND2_X1   g01158(.A1(new_n1027_), .A2(new_n479_), .ZN(new_n1352_));
  AOI21_X1   g01159(.A1(new_n1352_), .A2(new_n1351_), .B(new_n1350_), .ZN(new_n1353_));
  AOI22_X1   g01160(.A1(\a[2] ), .A2(\a[22] ), .B1(\a[6] ), .B2(\a[18] ), .ZN(new_n1354_));
  OR2_X2     g01161(.A1(new_n1353_), .A2(new_n1350_), .Z(new_n1355_));
  OAI22_X1   g01162(.A1(new_n1355_), .A2(new_n1354_), .B1(new_n1349_), .B2(new_n1353_), .ZN(new_n1356_));
  INV_X1     g01163(.I(\a[24] ), .ZN(new_n1357_));
  NOR2_X1    g01164(.A1(new_n196_), .A2(new_n1357_), .ZN(new_n1358_));
  XOR2_X1    g01165(.A1(new_n1320_), .A2(new_n1358_), .Z(new_n1359_));
  NOR2_X1    g01166(.A1(new_n194_), .A2(new_n1299_), .ZN(new_n1360_));
  XNOR2_X1   g01167(.A1(new_n1360_), .A2(new_n833_), .ZN(new_n1361_));
  XOR2_X1    g01168(.A1(new_n1359_), .A2(new_n1361_), .Z(new_n1362_));
  XOR2_X1    g01169(.A1(new_n1362_), .A2(new_n1356_), .Z(new_n1363_));
  XOR2_X1    g01170(.A1(new_n1363_), .A2(new_n1348_), .Z(new_n1364_));
  NAND2_X1   g01171(.A1(\a[8] ), .A2(\a[16] ), .ZN(new_n1365_));
  NAND2_X1   g01172(.A1(new_n467_), .A2(new_n1288_), .ZN(new_n1366_));
  INV_X1     g01173(.I(new_n413_), .ZN(new_n1367_));
  NAND2_X1   g01174(.A1(new_n895_), .A2(new_n1367_), .ZN(new_n1368_));
  AOI22_X1   g01175(.A1(new_n1366_), .A2(new_n1368_), .B1(new_n540_), .B2(new_n897_), .ZN(new_n1369_));
  NOR2_X1    g01176(.A1(new_n403_), .A2(new_n717_), .ZN(new_n1370_));
  AOI21_X1   g01177(.A1(\a[10] ), .A2(\a[14] ), .B(new_n1370_), .ZN(new_n1371_));
  NAND2_X1   g01178(.A1(new_n897_), .A2(new_n540_), .ZN(new_n1372_));
  NAND3_X1   g01179(.A1(new_n1372_), .A2(new_n1366_), .A3(new_n1368_), .ZN(new_n1373_));
  OAI22_X1   g01180(.A1(new_n1369_), .A2(new_n1365_), .B1(new_n1373_), .B2(new_n1371_), .ZN(new_n1374_));
  NOR2_X1    g01181(.A1(new_n979_), .A2(new_n1043_), .ZN(new_n1375_));
  INV_X1     g01182(.I(new_n1375_), .ZN(new_n1376_));
  NOR2_X1    g01183(.A1(new_n1376_), .A2(new_n242_), .ZN(new_n1377_));
  NOR2_X1    g01184(.A1(new_n979_), .A2(new_n1220_), .ZN(new_n1378_));
  INV_X1     g01185(.I(new_n1378_), .ZN(new_n1379_));
  NOR2_X1    g01186(.A1(new_n1379_), .A2(new_n318_), .ZN(new_n1380_));
  NOR2_X1    g01187(.A1(new_n1043_), .A2(new_n1220_), .ZN(new_n1381_));
  INV_X1     g01188(.I(new_n1381_), .ZN(new_n1382_));
  NOR2_X1    g01189(.A1(new_n1382_), .A2(new_n370_), .ZN(new_n1383_));
  NOR2_X1    g01190(.A1(new_n1380_), .A2(new_n1383_), .ZN(new_n1384_));
  NOR2_X1    g01191(.A1(new_n1384_), .A2(new_n1377_), .ZN(new_n1385_));
  NAND2_X1   g01192(.A1(\a[3] ), .A2(\a[21] ), .ZN(new_n1386_));
  AOI22_X1   g01193(.A1(\a[4] ), .A2(\a[20] ), .B1(\a[5] ), .B2(\a[19] ), .ZN(new_n1387_));
  NOR2_X1    g01194(.A1(new_n1385_), .A2(new_n1377_), .ZN(new_n1388_));
  INV_X1     g01195(.I(new_n1388_), .ZN(new_n1389_));
  OAI22_X1   g01196(.A1(new_n1389_), .A2(new_n1387_), .B1(new_n1385_), .B2(new_n1386_), .ZN(new_n1390_));
  XOR2_X1    g01197(.A1(new_n1390_), .A2(new_n1304_), .Z(new_n1391_));
  XOR2_X1    g01198(.A1(new_n1391_), .A2(new_n1374_), .Z(new_n1392_));
  XOR2_X1    g01199(.A1(new_n1364_), .A2(new_n1392_), .Z(new_n1393_));
  XOR2_X1    g01200(.A1(new_n1393_), .A2(new_n1345_), .Z(new_n1394_));
  NAND3_X1   g01201(.A1(new_n1311_), .A2(new_n1257_), .A3(new_n1312_), .ZN(new_n1395_));
  NAND2_X1   g01202(.A1(new_n1395_), .A2(new_n1311_), .ZN(new_n1396_));
  XOR2_X1    g01203(.A1(new_n1278_), .A2(new_n1268_), .Z(new_n1397_));
  XOR2_X1    g01204(.A1(new_n1397_), .A2(new_n1296_), .Z(new_n1398_));
  NAND2_X1   g01205(.A1(new_n1284_), .A2(new_n1271_), .ZN(new_n1399_));
  NAND2_X1   g01206(.A1(new_n1285_), .A2(new_n1260_), .ZN(new_n1400_));
  NAND2_X1   g01207(.A1(new_n1400_), .A2(new_n1399_), .ZN(new_n1401_));
  NAND2_X1   g01208(.A1(new_n1309_), .A2(new_n1297_), .ZN(new_n1402_));
  OAI21_X1   g01209(.A1(new_n1177_), .A2(new_n1308_), .B(new_n1402_), .ZN(new_n1403_));
  XOR2_X1    g01210(.A1(new_n1401_), .A2(new_n1403_), .Z(new_n1404_));
  NAND2_X1   g01211(.A1(new_n1404_), .A2(new_n1398_), .ZN(new_n1405_));
  OR2_X2     g01212(.A1(new_n1404_), .A2(new_n1398_), .Z(new_n1406_));
  NAND2_X1   g01213(.A1(new_n1406_), .A2(new_n1405_), .ZN(new_n1407_));
  XOR2_X1    g01214(.A1(new_n1407_), .A2(new_n1396_), .Z(new_n1408_));
  XOR2_X1    g01215(.A1(new_n1408_), .A2(new_n1394_), .Z(new_n1409_));
  NOR2_X1    g01216(.A1(new_n1409_), .A2(new_n1343_), .ZN(new_n1410_));
  INV_X1     g01217(.I(new_n1410_), .ZN(new_n1411_));
  NAND2_X1   g01218(.A1(new_n1409_), .A2(new_n1343_), .ZN(new_n1412_));
  NAND2_X1   g01219(.A1(new_n1411_), .A2(new_n1412_), .ZN(new_n1413_));
  INV_X1     g01220(.I(new_n1334_), .ZN(new_n1414_));
  OAI21_X1   g01221(.A1(new_n1249_), .A2(new_n1241_), .B(new_n1335_), .ZN(new_n1415_));
  INV_X1     g01222(.I(new_n1412_), .ZN(new_n1416_));
  AOI21_X1   g01223(.A1(new_n1415_), .A2(new_n1414_), .B(new_n1416_), .ZN(new_n1417_));
  AOI22_X1   g01224(.A1(new_n1417_), .A2(new_n1411_), .B1(new_n1340_), .B2(new_n1413_), .ZN(\asquared[25] ));
  OAI21_X1   g01225(.A1(new_n1339_), .A2(new_n1334_), .B(new_n1412_), .ZN(new_n1419_));
  NAND2_X1   g01226(.A1(new_n1419_), .A2(new_n1411_), .ZN(new_n1420_));
  AOI21_X1   g01227(.A1(new_n1311_), .A2(new_n1395_), .B(new_n1407_), .ZN(new_n1421_));
  INV_X1     g01228(.I(new_n1394_), .ZN(new_n1422_));
  NOR2_X1    g01229(.A1(new_n1408_), .A2(new_n1422_), .ZN(new_n1423_));
  NOR2_X1    g01230(.A1(new_n1423_), .A2(new_n1421_), .ZN(new_n1424_));
  NAND2_X1   g01231(.A1(new_n1401_), .A2(new_n1403_), .ZN(new_n1425_));
  NAND2_X1   g01232(.A1(new_n1405_), .A2(new_n1425_), .ZN(new_n1426_));
  INV_X1     g01233(.I(new_n467_), .ZN(new_n1427_));
  INV_X1     g01234(.I(new_n1024_), .ZN(new_n1428_));
  INV_X1     g01235(.I(new_n1025_), .ZN(new_n1429_));
  OAI22_X1   g01236(.A1(new_n415_), .A2(new_n1275_), .B1(new_n1429_), .B2(new_n773_), .ZN(new_n1430_));
  OAI21_X1   g01237(.A1(new_n1427_), .A2(new_n1428_), .B(new_n1430_), .ZN(new_n1431_));
  NAND3_X1   g01238(.A1(new_n1431_), .A2(\a[7] ), .A3(\a[18] ), .ZN(new_n1432_));
  AOI22_X1   g01239(.A1(\a[8] ), .A2(\a[17] ), .B1(\a[9] ), .B2(\a[16] ), .ZN(new_n1433_));
  NOR2_X1    g01240(.A1(new_n1428_), .A2(new_n1427_), .ZN(new_n1434_));
  NOR2_X1    g01241(.A1(new_n1430_), .A2(new_n1434_), .ZN(new_n1435_));
  INV_X1     g01242(.I(new_n1435_), .ZN(new_n1436_));
  OAI21_X1   g01243(.A1(new_n1433_), .A2(new_n1436_), .B(new_n1432_), .ZN(new_n1437_));
  AOI22_X1   g01244(.A1(\a[0] ), .A2(\a[25] ), .B1(\a[2] ), .B2(\a[23] ), .ZN(new_n1438_));
  INV_X1     g01245(.I(new_n710_), .ZN(new_n1439_));
  INV_X1     g01246(.I(new_n1438_), .ZN(new_n1440_));
  INV_X1     g01247(.I(\a[25] ), .ZN(new_n1441_));
  NOR2_X1    g01248(.A1(new_n1299_), .A2(new_n1441_), .ZN(new_n1442_));
  INV_X1     g01249(.I(new_n1442_), .ZN(new_n1443_));
  NOR2_X1    g01250(.A1(new_n1443_), .A2(new_n412_), .ZN(new_n1444_));
  AOI21_X1   g01251(.A1(new_n1439_), .A2(new_n1440_), .B(new_n1444_), .ZN(new_n1445_));
  INV_X1     g01252(.I(new_n1445_), .ZN(new_n1446_));
  OAI21_X1   g01253(.A1(new_n1444_), .A2(new_n1438_), .B(new_n1439_), .ZN(new_n1447_));
  OAI21_X1   g01254(.A1(new_n1446_), .A2(new_n1438_), .B(new_n1447_), .ZN(new_n1448_));
  XNOR2_X1   g01255(.A1(new_n1437_), .A2(new_n1448_), .ZN(new_n1449_));
  AOI22_X1   g01256(.A1(\a[4] ), .A2(new_n1378_), .B1(new_n1191_), .B2(\a[22] ), .ZN(new_n1450_));
  INV_X1     g01257(.I(new_n1450_), .ZN(new_n1451_));
  NOR2_X1    g01258(.A1(new_n1220_), .A2(new_n1175_), .ZN(new_n1452_));
  AOI21_X1   g01259(.A1(new_n1452_), .A2(new_n761_), .B(new_n367_), .ZN(new_n1453_));
  NAND2_X1   g01260(.A1(new_n1451_), .A2(new_n1453_), .ZN(new_n1454_));
  NOR2_X1    g01261(.A1(new_n367_), .A2(new_n979_), .ZN(new_n1455_));
  INV_X1     g01262(.I(new_n1452_), .ZN(new_n1456_));
  OAI21_X1   g01263(.A1(new_n370_), .A2(new_n1456_), .B(new_n1454_), .ZN(new_n1457_));
  INV_X1     g01264(.I(new_n1457_), .ZN(new_n1458_));
  OAI22_X1   g01265(.A1(new_n225_), .A2(new_n1175_), .B1(new_n290_), .B2(new_n1220_), .ZN(new_n1459_));
  AOI22_X1   g01266(.A1(new_n1458_), .A2(new_n1459_), .B1(new_n1454_), .B2(new_n1455_), .ZN(new_n1460_));
  XNOR2_X1   g01267(.A1(new_n1449_), .A2(new_n1460_), .ZN(new_n1461_));
  INV_X1     g01268(.I(new_n1461_), .ZN(new_n1462_));
  XOR2_X1    g01269(.A1(new_n1426_), .A2(new_n1462_), .Z(new_n1463_));
  INV_X1     g01270(.I(new_n1360_), .ZN(new_n1464_));
  NOR2_X1    g01271(.A1(new_n1464_), .A2(new_n833_), .ZN(new_n1465_));
  INV_X1     g01272(.I(new_n1465_), .ZN(new_n1466_));
  NOR2_X1    g01273(.A1(new_n194_), .A2(new_n1357_), .ZN(new_n1467_));
  INV_X1     g01274(.I(new_n1467_), .ZN(new_n1468_));
  NAND2_X1   g01275(.A1(new_n1468_), .A2(new_n597_), .ZN(new_n1469_));
  NOR2_X1    g01276(.A1(new_n1468_), .A2(new_n597_), .ZN(new_n1470_));
  INV_X1     g01277(.I(new_n1470_), .ZN(new_n1471_));
  AND2_X2    g01278(.A1(new_n1471_), .A2(new_n1469_), .Z(new_n1472_));
  INV_X1     g01279(.I(new_n1472_), .ZN(new_n1473_));
  NOR2_X1    g01280(.A1(new_n1473_), .A2(new_n1466_), .ZN(new_n1474_));
  NOR2_X1    g01281(.A1(new_n1472_), .A2(new_n1465_), .ZN(new_n1475_));
  NOR2_X1    g01282(.A1(new_n1474_), .A2(new_n1475_), .ZN(new_n1476_));
  XOR2_X1    g01283(.A1(new_n1476_), .A2(new_n1389_), .Z(new_n1477_));
  NAND2_X1   g01284(.A1(new_n1397_), .A2(new_n1296_), .ZN(new_n1478_));
  OAI21_X1   g01285(.A1(new_n1268_), .A2(new_n1278_), .B(new_n1478_), .ZN(new_n1479_));
  NOR2_X1    g01286(.A1(new_n253_), .A2(new_n1043_), .ZN(new_n1480_));
  INV_X1     g01287(.I(new_n1480_), .ZN(new_n1481_));
  NOR2_X1    g01288(.A1(new_n513_), .A2(new_n759_), .ZN(new_n1482_));
  NOR2_X1    g01289(.A1(new_n763_), .A2(new_n1482_), .ZN(new_n1483_));
  NAND2_X1   g01290(.A1(new_n763_), .A2(new_n1482_), .ZN(new_n1484_));
  INV_X1     g01291(.I(new_n1484_), .ZN(new_n1485_));
  NOR3_X1    g01292(.A1(new_n1485_), .A2(new_n1481_), .A3(new_n1483_), .ZN(new_n1486_));
  NOR2_X1    g01293(.A1(new_n1486_), .A2(new_n1485_), .ZN(new_n1487_));
  INV_X1     g01294(.I(new_n1487_), .ZN(new_n1488_));
  OAI22_X1   g01295(.A1(new_n1488_), .A2(new_n1483_), .B1(new_n1481_), .B2(new_n1486_), .ZN(new_n1489_));
  XOR2_X1    g01296(.A1(new_n1479_), .A2(new_n1489_), .Z(new_n1490_));
  XNOR2_X1   g01297(.A1(new_n1490_), .A2(new_n1477_), .ZN(new_n1491_));
  XOR2_X1    g01298(.A1(new_n1463_), .A2(new_n1491_), .Z(new_n1492_));
  NAND2_X1   g01299(.A1(new_n1362_), .A2(new_n1356_), .ZN(new_n1493_));
  NAND2_X1   g01300(.A1(new_n1363_), .A2(new_n1348_), .ZN(new_n1494_));
  NAND2_X1   g01301(.A1(new_n1494_), .A2(new_n1493_), .ZN(new_n1495_));
  NAND2_X1   g01302(.A1(new_n1320_), .A2(new_n1358_), .ZN(new_n1496_));
  NAND2_X1   g01303(.A1(new_n1359_), .A2(new_n1361_), .ZN(new_n1497_));
  NAND2_X1   g01304(.A1(new_n1497_), .A2(new_n1496_), .ZN(new_n1498_));
  XOR2_X1    g01305(.A1(new_n1355_), .A2(new_n1373_), .Z(new_n1499_));
  XOR2_X1    g01306(.A1(new_n1499_), .A2(new_n1498_), .Z(new_n1500_));
  NAND2_X1   g01307(.A1(new_n1391_), .A2(new_n1374_), .ZN(new_n1501_));
  NAND2_X1   g01308(.A1(new_n1390_), .A2(new_n1304_), .ZN(new_n1502_));
  NAND2_X1   g01309(.A1(new_n1501_), .A2(new_n1502_), .ZN(new_n1503_));
  XOR2_X1    g01310(.A1(new_n1503_), .A2(new_n1500_), .Z(new_n1504_));
  XOR2_X1    g01311(.A1(new_n1504_), .A2(new_n1495_), .Z(new_n1505_));
  NAND2_X1   g01312(.A1(new_n1392_), .A2(new_n1364_), .ZN(new_n1506_));
  NAND2_X1   g01313(.A1(new_n1393_), .A2(new_n1345_), .ZN(new_n1507_));
  NAND2_X1   g01314(.A1(new_n1507_), .A2(new_n1506_), .ZN(new_n1508_));
  XNOR2_X1   g01315(.A1(new_n1508_), .A2(new_n1505_), .ZN(new_n1509_));
  NOR2_X1    g01316(.A1(new_n1492_), .A2(new_n1509_), .ZN(new_n1510_));
  INV_X1     g01317(.I(new_n1510_), .ZN(new_n1511_));
  NAND2_X1   g01318(.A1(new_n1492_), .A2(new_n1509_), .ZN(new_n1512_));
  NAND2_X1   g01319(.A1(new_n1511_), .A2(new_n1512_), .ZN(new_n1513_));
  NAND2_X1   g01320(.A1(new_n1513_), .A2(new_n1424_), .ZN(new_n1514_));
  INV_X1     g01321(.I(new_n1514_), .ZN(new_n1515_));
  NOR2_X1    g01322(.A1(new_n1513_), .A2(new_n1424_), .ZN(new_n1516_));
  NOR2_X1    g01323(.A1(new_n1515_), .A2(new_n1516_), .ZN(new_n1517_));
  XOR2_X1    g01324(.A1(new_n1420_), .A2(new_n1517_), .Z(\asquared[26] ));
  AOI21_X1   g01325(.A1(new_n1419_), .A2(new_n1411_), .B(new_n1515_), .ZN(new_n1519_));
  NOR2_X1    g01326(.A1(new_n1519_), .A2(new_n1516_), .ZN(new_n1520_));
  NAND2_X1   g01327(.A1(new_n1508_), .A2(new_n1505_), .ZN(new_n1521_));
  NAND2_X1   g01328(.A1(new_n1511_), .A2(new_n1521_), .ZN(new_n1522_));
  INV_X1     g01329(.I(new_n1522_), .ZN(new_n1523_));
  NAND2_X1   g01330(.A1(new_n1503_), .A2(new_n1500_), .ZN(new_n1524_));
  NAND2_X1   g01331(.A1(new_n1504_), .A2(new_n1495_), .ZN(new_n1525_));
  NAND2_X1   g01332(.A1(new_n1525_), .A2(new_n1524_), .ZN(new_n1526_));
  NOR3_X1    g01333(.A1(new_n378_), .A2(new_n979_), .A3(new_n1357_), .ZN(new_n1527_));
  NOR2_X1    g01334(.A1(new_n1299_), .A2(new_n1357_), .ZN(new_n1528_));
  INV_X1     g01335(.I(new_n1528_), .ZN(new_n1529_));
  NOR2_X1    g01336(.A1(new_n1529_), .A2(new_n246_), .ZN(new_n1530_));
  NOR2_X1    g01337(.A1(new_n1530_), .A2(new_n1527_), .ZN(new_n1531_));
  NOR2_X1    g01338(.A1(new_n225_), .A2(new_n1299_), .ZN(new_n1532_));
  NOR2_X1    g01339(.A1(new_n422_), .A2(new_n979_), .ZN(new_n1533_));
  NAND2_X1   g01340(.A1(new_n1532_), .A2(new_n1533_), .ZN(new_n1534_));
  INV_X1     g01341(.I(new_n1534_), .ZN(new_n1535_));
  NOR2_X1    g01342(.A1(new_n1531_), .A2(new_n1535_), .ZN(new_n1536_));
  NAND2_X1   g01343(.A1(\a[2] ), .A2(\a[24] ), .ZN(new_n1537_));
  NOR2_X1    g01344(.A1(new_n1532_), .A2(new_n1533_), .ZN(new_n1538_));
  NOR2_X1    g01345(.A1(new_n1536_), .A2(new_n1535_), .ZN(new_n1539_));
  INV_X1     g01346(.I(new_n1539_), .ZN(new_n1540_));
  OAI22_X1   g01347(.A1(new_n1540_), .A2(new_n1538_), .B1(new_n1536_), .B2(new_n1537_), .ZN(new_n1541_));
  NOR2_X1    g01348(.A1(new_n403_), .A2(new_n1023_), .ZN(new_n1542_));
  INV_X1     g01349(.I(new_n1542_), .ZN(new_n1543_));
  NAND2_X1   g01350(.A1(new_n1024_), .A2(new_n540_), .ZN(new_n1544_));
  NAND2_X1   g01351(.A1(new_n832_), .A2(new_n1542_), .ZN(new_n1545_));
  AOI22_X1   g01352(.A1(new_n1545_), .A2(new_n1544_), .B1(new_n747_), .B2(new_n1288_), .ZN(new_n1546_));
  AOI21_X1   g01353(.A1(\a[10] ), .A2(\a[16] ), .B(new_n832_), .ZN(new_n1547_));
  NAND2_X1   g01354(.A1(new_n747_), .A2(new_n1288_), .ZN(new_n1548_));
  NAND3_X1   g01355(.A1(new_n1548_), .A2(new_n1545_), .A3(new_n1544_), .ZN(new_n1549_));
  OAI22_X1   g01356(.A1(new_n1546_), .A2(new_n1543_), .B1(new_n1549_), .B2(new_n1547_), .ZN(new_n1550_));
  XOR2_X1    g01357(.A1(new_n1541_), .A2(new_n1550_), .Z(new_n1551_));
  NOR2_X1    g01358(.A1(new_n1043_), .A2(new_n1175_), .ZN(new_n1552_));
  NAND3_X1   g01359(.A1(new_n1552_), .A2(\a[4] ), .A3(\a[6] ), .ZN(new_n1553_));
  NAND2_X1   g01360(.A1(new_n1452_), .A2(new_n243_), .ZN(new_n1554_));
  AOI22_X1   g01361(.A1(new_n1553_), .A2(new_n1554_), .B1(new_n746_), .B2(new_n1381_), .ZN(new_n1555_));
  NAND2_X1   g01362(.A1(\a[4] ), .A2(\a[22] ), .ZN(new_n1556_));
  AOI22_X1   g01363(.A1(\a[5] ), .A2(\a[21] ), .B1(\a[6] ), .B2(\a[20] ), .ZN(new_n1557_));
  NAND2_X1   g01364(.A1(new_n1381_), .A2(new_n746_), .ZN(new_n1558_));
  NAND3_X1   g01365(.A1(new_n1558_), .A2(new_n1553_), .A3(new_n1554_), .ZN(new_n1559_));
  OAI22_X1   g01366(.A1(new_n1555_), .A2(new_n1556_), .B1(new_n1559_), .B2(new_n1557_), .ZN(new_n1560_));
  XNOR2_X1   g01367(.A1(new_n1551_), .A2(new_n1560_), .ZN(new_n1561_));
  INV_X1     g01368(.I(new_n1561_), .ZN(new_n1562_));
  XOR2_X1    g01369(.A1(new_n1526_), .A2(new_n1562_), .Z(new_n1563_));
  XOR2_X1    g01370(.A1(new_n1435_), .A2(new_n1445_), .Z(new_n1564_));
  AOI22_X1   g01371(.A1(\a[0] ), .A2(\a[26] ), .B1(\a[8] ), .B2(\a[18] ), .ZN(new_n1565_));
  INV_X1     g01372(.I(\a[26] ), .ZN(new_n1566_));
  NOR4_X1    g01373(.A1(new_n196_), .A2(new_n355_), .A3(new_n884_), .A4(new_n1566_), .ZN(new_n1567_));
  NOR3_X1    g01374(.A1(new_n1471_), .A2(new_n1565_), .A3(new_n1567_), .ZN(new_n1568_));
  NOR2_X1    g01375(.A1(new_n1568_), .A2(new_n1567_), .ZN(new_n1569_));
  INV_X1     g01376(.I(new_n1569_), .ZN(new_n1570_));
  OAI22_X1   g01377(.A1(new_n1570_), .A2(new_n1565_), .B1(new_n1471_), .B2(new_n1568_), .ZN(new_n1571_));
  XNOR2_X1   g01378(.A1(new_n1571_), .A2(new_n1564_), .ZN(new_n1572_));
  INV_X1     g01379(.I(new_n1572_), .ZN(new_n1573_));
  NAND2_X1   g01380(.A1(new_n1355_), .A2(new_n1373_), .ZN(new_n1574_));
  NAND2_X1   g01381(.A1(new_n1499_), .A2(new_n1498_), .ZN(new_n1575_));
  NAND2_X1   g01382(.A1(new_n1575_), .A2(new_n1574_), .ZN(new_n1576_));
  INV_X1     g01383(.I(new_n1474_), .ZN(new_n1577_));
  OAI21_X1   g01384(.A1(new_n1388_), .A2(new_n1475_), .B(new_n1577_), .ZN(new_n1578_));
  XOR2_X1    g01385(.A1(new_n1576_), .A2(new_n1578_), .Z(new_n1579_));
  XOR2_X1    g01386(.A1(new_n1579_), .A2(new_n1573_), .Z(new_n1580_));
  XNOR2_X1   g01387(.A1(new_n1563_), .A2(new_n1580_), .ZN(new_n1581_));
  NAND2_X1   g01388(.A1(new_n1426_), .A2(new_n1462_), .ZN(new_n1582_));
  INV_X1     g01389(.I(new_n1491_), .ZN(new_n1583_));
  NAND2_X1   g01390(.A1(new_n1463_), .A2(new_n1583_), .ZN(new_n1584_));
  NAND2_X1   g01391(.A1(new_n1584_), .A2(new_n1582_), .ZN(new_n1585_));
  NAND2_X1   g01392(.A1(new_n1479_), .A2(new_n1489_), .ZN(new_n1586_));
  NAND2_X1   g01393(.A1(new_n1490_), .A2(new_n1477_), .ZN(new_n1587_));
  NAND2_X1   g01394(.A1(new_n1587_), .A2(new_n1586_), .ZN(new_n1588_));
  NAND2_X1   g01395(.A1(new_n1437_), .A2(new_n1448_), .ZN(new_n1589_));
  OAI21_X1   g01396(.A1(new_n1449_), .A2(new_n1460_), .B(new_n1589_), .ZN(new_n1590_));
  NOR2_X1    g01397(.A1(new_n194_), .A2(new_n1441_), .ZN(new_n1591_));
  NAND2_X1   g01398(.A1(new_n1591_), .A2(new_n762_), .ZN(new_n1592_));
  INV_X1     g01399(.I(new_n1591_), .ZN(new_n1593_));
  NAND2_X1   g01400(.A1(new_n1593_), .A2(new_n623_), .ZN(new_n1594_));
  AND2_X2    g01401(.A1(new_n1594_), .A2(new_n1592_), .Z(new_n1595_));
  NOR2_X1    g01402(.A1(new_n1487_), .A2(new_n1595_), .ZN(new_n1596_));
  INV_X1     g01403(.I(new_n1595_), .ZN(new_n1597_));
  NOR2_X1    g01404(.A1(new_n1488_), .A2(new_n1597_), .ZN(new_n1598_));
  NOR2_X1    g01405(.A1(new_n1598_), .A2(new_n1596_), .ZN(new_n1599_));
  NOR2_X1    g01406(.A1(new_n1599_), .A2(new_n1458_), .ZN(new_n1600_));
  NOR3_X1    g01407(.A1(new_n1598_), .A2(new_n1457_), .A3(new_n1596_), .ZN(new_n1601_));
  NOR2_X1    g01408(.A1(new_n1600_), .A2(new_n1601_), .ZN(new_n1602_));
  XOR2_X1    g01409(.A1(new_n1590_), .A2(new_n1602_), .Z(new_n1603_));
  XOR2_X1    g01410(.A1(new_n1588_), .A2(new_n1603_), .Z(new_n1604_));
  XNOR2_X1   g01411(.A1(new_n1585_), .A2(new_n1604_), .ZN(new_n1605_));
  XNOR2_X1   g01412(.A1(new_n1605_), .A2(new_n1581_), .ZN(new_n1606_));
  NAND2_X1   g01413(.A1(new_n1606_), .A2(new_n1523_), .ZN(new_n1607_));
  NOR2_X1    g01414(.A1(new_n1606_), .A2(new_n1523_), .ZN(new_n1608_));
  INV_X1     g01415(.I(new_n1608_), .ZN(new_n1609_));
  NAND2_X1   g01416(.A1(new_n1609_), .A2(new_n1607_), .ZN(new_n1610_));
  XOR2_X1    g01417(.A1(new_n1520_), .A2(new_n1610_), .Z(\asquared[27] ));
  OAI21_X1   g01418(.A1(new_n1519_), .A2(new_n1516_), .B(new_n1607_), .ZN(new_n1612_));
  NAND2_X1   g01419(.A1(new_n1612_), .A2(new_n1609_), .ZN(new_n1613_));
  NAND2_X1   g01420(.A1(new_n1585_), .A2(new_n1604_), .ZN(new_n1614_));
  OAI21_X1   g01421(.A1(new_n1605_), .A2(new_n1581_), .B(new_n1614_), .ZN(new_n1615_));
  NAND2_X1   g01422(.A1(new_n1541_), .A2(new_n1550_), .ZN(new_n1616_));
  NAND2_X1   g01423(.A1(new_n1551_), .A2(new_n1560_), .ZN(new_n1617_));
  NAND2_X1   g01424(.A1(new_n1617_), .A2(new_n1616_), .ZN(new_n1618_));
  NOR2_X1    g01425(.A1(new_n1597_), .A2(new_n1487_), .ZN(new_n1619_));
  NOR2_X1    g01426(.A1(new_n1600_), .A2(new_n1619_), .ZN(new_n1620_));
  NAND2_X1   g01427(.A1(new_n1571_), .A2(new_n1564_), .ZN(new_n1621_));
  OAI21_X1   g01428(.A1(new_n1435_), .A2(new_n1445_), .B(new_n1621_), .ZN(new_n1622_));
  XNOR2_X1   g01429(.A1(new_n1622_), .A2(new_n1620_), .ZN(new_n1623_));
  XOR2_X1    g01430(.A1(new_n1623_), .A2(new_n1618_), .Z(new_n1624_));
  NAND2_X1   g01431(.A1(new_n1590_), .A2(new_n1602_), .ZN(new_n1625_));
  NAND2_X1   g01432(.A1(new_n1588_), .A2(new_n1603_), .ZN(new_n1626_));
  NAND2_X1   g01433(.A1(new_n1626_), .A2(new_n1625_), .ZN(new_n1627_));
  NOR2_X1    g01434(.A1(new_n513_), .A2(new_n742_), .ZN(new_n1628_));
  NOR3_X1    g01435(.A1(new_n378_), .A2(new_n1043_), .A3(new_n1441_), .ZN(new_n1629_));
  AOI22_X1   g01436(.A1(\a[2] ), .A2(\a[25] ), .B1(\a[7] ), .B2(\a[20] ), .ZN(new_n1630_));
  NOR2_X1    g01437(.A1(new_n1629_), .A2(new_n1630_), .ZN(new_n1631_));
  XOR2_X1    g01438(.A1(new_n1631_), .A2(new_n1628_), .Z(new_n1632_));
  INV_X1     g01439(.I(new_n1632_), .ZN(new_n1633_));
  NOR2_X1    g01440(.A1(new_n1569_), .A2(new_n1633_), .ZN(new_n1634_));
  NOR2_X1    g01441(.A1(new_n1570_), .A2(new_n1632_), .ZN(new_n1635_));
  NOR2_X1    g01442(.A1(new_n1635_), .A2(new_n1634_), .ZN(new_n1636_));
  NAND2_X1   g01443(.A1(\a[8] ), .A2(\a[19] ), .ZN(new_n1637_));
  NAND4_X1   g01444(.A1(\a[8] ), .A2(\a[10] ), .A3(\a[17] ), .A4(\a[19] ), .ZN(new_n1638_));
  NAND2_X1   g01445(.A1(new_n467_), .A2(new_n1194_), .ZN(new_n1639_));
  AOI22_X1   g01446(.A1(new_n1639_), .A2(new_n1638_), .B1(new_n540_), .B2(new_n1027_), .ZN(new_n1640_));
  AOI22_X1   g01447(.A1(\a[9] ), .A2(\a[18] ), .B1(\a[10] ), .B2(\a[17] ), .ZN(new_n1641_));
  NAND2_X1   g01448(.A1(new_n1027_), .A2(new_n540_), .ZN(new_n1642_));
  NAND3_X1   g01449(.A1(new_n1642_), .A2(new_n1639_), .A3(new_n1638_), .ZN(new_n1643_));
  OAI22_X1   g01450(.A1(new_n1640_), .A2(new_n1637_), .B1(new_n1643_), .B2(new_n1641_), .ZN(new_n1644_));
  XNOR2_X1   g01451(.A1(new_n1636_), .A2(new_n1644_), .ZN(new_n1645_));
  INV_X1     g01452(.I(new_n1645_), .ZN(new_n1646_));
  XOR2_X1    g01453(.A1(new_n1627_), .A2(new_n1646_), .Z(new_n1647_));
  NAND2_X1   g01454(.A1(new_n1647_), .A2(new_n1624_), .ZN(new_n1648_));
  INV_X1     g01455(.I(new_n1648_), .ZN(new_n1649_));
  NOR2_X1    g01456(.A1(new_n1647_), .A2(new_n1624_), .ZN(new_n1650_));
  NOR2_X1    g01457(.A1(new_n1649_), .A2(new_n1650_), .ZN(new_n1651_));
  NAND2_X1   g01458(.A1(new_n1526_), .A2(new_n1562_), .ZN(new_n1652_));
  NAND2_X1   g01459(.A1(new_n1563_), .A2(new_n1580_), .ZN(new_n1653_));
  NAND2_X1   g01460(.A1(new_n1653_), .A2(new_n1652_), .ZN(new_n1654_));
  NOR2_X1    g01461(.A1(new_n686_), .A2(new_n1566_), .ZN(new_n1655_));
  INV_X1     g01462(.I(new_n1655_), .ZN(new_n1656_));
  NOR2_X1    g01463(.A1(new_n194_), .A2(new_n1566_), .ZN(new_n1657_));
  OAI21_X1   g01464(.A1(\a[14] ), .A2(new_n1657_), .B(new_n1656_), .ZN(new_n1658_));
  NAND2_X1   g01465(.A1(\a[0] ), .A2(\a[27] ), .ZN(new_n1659_));
  XNOR2_X1   g01466(.A1(new_n1592_), .A2(new_n1659_), .ZN(new_n1660_));
  XOR2_X1    g01467(.A1(new_n1660_), .A2(new_n1658_), .Z(new_n1661_));
  NOR2_X1    g01468(.A1(new_n367_), .A2(new_n1220_), .ZN(new_n1662_));
  NOR2_X1    g01469(.A1(new_n290_), .A2(new_n1299_), .ZN(new_n1663_));
  NAND2_X1   g01470(.A1(new_n1662_), .A2(new_n1663_), .ZN(new_n1664_));
  NAND2_X1   g01471(.A1(\a[21] ), .A2(\a[24] ), .ZN(new_n1665_));
  OAI22_X1   g01472(.A1(new_n1529_), .A2(new_n370_), .B1(new_n1274_), .B2(new_n1665_), .ZN(new_n1666_));
  NAND2_X1   g01473(.A1(new_n1666_), .A2(new_n1664_), .ZN(new_n1667_));
  NAND3_X1   g01474(.A1(new_n1667_), .A2(\a[3] ), .A3(\a[24] ), .ZN(new_n1668_));
  NAND2_X1   g01475(.A1(new_n1667_), .A2(new_n1664_), .ZN(new_n1669_));
  NOR2_X1    g01476(.A1(new_n1662_), .A2(new_n1663_), .ZN(new_n1670_));
  OAI21_X1   g01477(.A1(new_n1669_), .A2(new_n1670_), .B(new_n1668_), .ZN(new_n1671_));
  AOI21_X1   g01478(.A1(\a[12] ), .A2(\a[15] ), .B(new_n760_), .ZN(new_n1672_));
  NOR2_X1    g01479(.A1(new_n253_), .A2(new_n1175_), .ZN(new_n1673_));
  INV_X1     g01480(.I(new_n1673_), .ZN(new_n1674_));
  OAI22_X1   g01481(.A1(new_n1672_), .A2(new_n1674_), .B1(new_n1265_), .B2(new_n1173_), .ZN(new_n1675_));
  NOR2_X1    g01482(.A1(new_n1265_), .A2(new_n1173_), .ZN(new_n1676_));
  OAI21_X1   g01483(.A1(new_n1676_), .A2(new_n1672_), .B(new_n1673_), .ZN(new_n1677_));
  OAI21_X1   g01484(.A1(new_n1675_), .A2(new_n1672_), .B(new_n1677_), .ZN(new_n1678_));
  XOR2_X1    g01485(.A1(new_n1671_), .A2(new_n1678_), .Z(new_n1679_));
  XNOR2_X1   g01486(.A1(new_n1679_), .A2(new_n1661_), .ZN(new_n1680_));
  INV_X1     g01487(.I(new_n1680_), .ZN(new_n1681_));
  NAND2_X1   g01488(.A1(new_n1576_), .A2(new_n1578_), .ZN(new_n1682_));
  NAND2_X1   g01489(.A1(new_n1579_), .A2(new_n1573_), .ZN(new_n1683_));
  NAND2_X1   g01490(.A1(new_n1683_), .A2(new_n1682_), .ZN(new_n1684_));
  XOR2_X1    g01491(.A1(new_n1549_), .A2(new_n1559_), .Z(new_n1685_));
  XNOR2_X1   g01492(.A1(new_n1685_), .A2(new_n1539_), .ZN(new_n1686_));
  XOR2_X1    g01493(.A1(new_n1684_), .A2(new_n1686_), .Z(new_n1687_));
  XOR2_X1    g01494(.A1(new_n1687_), .A2(new_n1681_), .Z(new_n1688_));
  NOR2_X1    g01495(.A1(new_n1654_), .A2(new_n1688_), .ZN(new_n1689_));
  NAND2_X1   g01496(.A1(new_n1654_), .A2(new_n1688_), .ZN(new_n1690_));
  INV_X1     g01497(.I(new_n1690_), .ZN(new_n1691_));
  NOR2_X1    g01498(.A1(new_n1691_), .A2(new_n1689_), .ZN(new_n1692_));
  XOR2_X1    g01499(.A1(new_n1692_), .A2(new_n1651_), .Z(new_n1693_));
  NOR2_X1    g01500(.A1(new_n1693_), .A2(new_n1615_), .ZN(new_n1694_));
  NAND2_X1   g01501(.A1(new_n1693_), .A2(new_n1615_), .ZN(new_n1695_));
  INV_X1     g01502(.I(new_n1695_), .ZN(new_n1696_));
  NOR2_X1    g01503(.A1(new_n1696_), .A2(new_n1694_), .ZN(new_n1697_));
  XOR2_X1    g01504(.A1(new_n1613_), .A2(new_n1697_), .Z(\asquared[28] ));
  AOI21_X1   g01505(.A1(new_n1612_), .A2(new_n1609_), .B(new_n1694_), .ZN(new_n1699_));
  NOR2_X1    g01506(.A1(new_n1699_), .A2(new_n1696_), .ZN(new_n1700_));
  INV_X1     g01507(.I(new_n1651_), .ZN(new_n1701_));
  OAI21_X1   g01508(.A1(new_n1701_), .A2(new_n1689_), .B(new_n1690_), .ZN(new_n1702_));
  NAND2_X1   g01509(.A1(new_n1627_), .A2(new_n1646_), .ZN(new_n1703_));
  NAND2_X1   g01510(.A1(new_n1648_), .A2(new_n1703_), .ZN(new_n1704_));
  INV_X1     g01511(.I(new_n1704_), .ZN(new_n1705_));
  NAND2_X1   g01512(.A1(new_n1549_), .A2(new_n1559_), .ZN(new_n1706_));
  NAND2_X1   g01513(.A1(new_n1540_), .A2(new_n1685_), .ZN(new_n1707_));
  NAND2_X1   g01514(.A1(new_n1707_), .A2(new_n1706_), .ZN(new_n1708_));
  AOI22_X1   g01515(.A1(\a[9] ), .A2(\a[19] ), .B1(\a[10] ), .B2(\a[18] ), .ZN(new_n1709_));
  NOR2_X1    g01516(.A1(new_n197_), .A2(new_n1566_), .ZN(new_n1710_));
  NOR2_X1    g01517(.A1(new_n539_), .A2(new_n1092_), .ZN(new_n1711_));
  OAI21_X1   g01518(.A1(new_n1711_), .A2(new_n1709_), .B(new_n1710_), .ZN(new_n1712_));
  INV_X1     g01519(.I(new_n1709_), .ZN(new_n1713_));
  AOI21_X1   g01520(.A1(new_n1713_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n1714_));
  INV_X1     g01521(.I(new_n1714_), .ZN(new_n1715_));
  OAI21_X1   g01522(.A1(new_n1715_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n1716_));
  NOR2_X1    g01523(.A1(new_n536_), .A2(new_n742_), .ZN(new_n1717_));
  INV_X1     g01524(.I(\a[28] ), .ZN(new_n1718_));
  NOR2_X1    g01525(.A1(new_n196_), .A2(new_n1718_), .ZN(new_n1719_));
  NAND2_X1   g01526(.A1(new_n1717_), .A2(new_n1719_), .ZN(new_n1720_));
  NOR2_X1    g01527(.A1(new_n513_), .A2(new_n1718_), .ZN(new_n1721_));
  INV_X1     g01528(.I(new_n1721_), .ZN(new_n1722_));
  OAI22_X1   g01529(.A1(new_n619_), .A2(new_n1428_), .B1(new_n1722_), .B2(new_n814_), .ZN(new_n1723_));
  NAND2_X1   g01530(.A1(new_n1723_), .A2(new_n1720_), .ZN(new_n1724_));
  NAND3_X1   g01531(.A1(new_n1724_), .A2(\a[11] ), .A3(\a[17] ), .ZN(new_n1725_));
  NAND2_X1   g01532(.A1(new_n1724_), .A2(new_n1720_), .ZN(new_n1726_));
  NOR2_X1    g01533(.A1(new_n1717_), .A2(new_n1719_), .ZN(new_n1727_));
  OAI21_X1   g01534(.A1(new_n1726_), .A2(new_n1727_), .B(new_n1725_), .ZN(new_n1728_));
  XNOR2_X1   g01535(.A1(new_n1728_), .A2(new_n1716_), .ZN(new_n1729_));
  XNOR2_X1   g01536(.A1(new_n1729_), .A2(new_n1708_), .ZN(new_n1730_));
  OAI21_X1   g01537(.A1(new_n1619_), .A2(new_n1600_), .B(new_n1622_), .ZN(new_n1731_));
  NAND2_X1   g01538(.A1(new_n1623_), .A2(new_n1618_), .ZN(new_n1732_));
  NAND2_X1   g01539(.A1(new_n1732_), .A2(new_n1731_), .ZN(new_n1733_));
  INV_X1     g01540(.I(new_n1628_), .ZN(new_n1734_));
  INV_X1     g01541(.I(new_n1629_), .ZN(new_n1735_));
  OAI21_X1   g01542(.A1(new_n1734_), .A2(new_n1630_), .B(new_n1735_), .ZN(new_n1736_));
  XOR2_X1    g01543(.A1(new_n1669_), .A2(new_n1643_), .Z(new_n1737_));
  XOR2_X1    g01544(.A1(new_n1737_), .A2(new_n1736_), .Z(new_n1738_));
  XOR2_X1    g01545(.A1(new_n1733_), .A2(new_n1738_), .Z(new_n1739_));
  XNOR2_X1   g01546(.A1(new_n1739_), .A2(new_n1730_), .ZN(new_n1740_));
  NAND2_X1   g01547(.A1(new_n1705_), .A2(new_n1740_), .ZN(new_n1741_));
  NOR2_X1    g01548(.A1(new_n1705_), .A2(new_n1740_), .ZN(new_n1742_));
  INV_X1     g01549(.I(new_n1742_), .ZN(new_n1743_));
  NAND2_X1   g01550(.A1(new_n1743_), .A2(new_n1741_), .ZN(new_n1744_));
  XOR2_X1    g01551(.A1(new_n1744_), .A2(new_n1702_), .Z(new_n1745_));
  NAND2_X1   g01552(.A1(new_n1671_), .A2(new_n1678_), .ZN(new_n1746_));
  INV_X1     g01553(.I(new_n1746_), .ZN(new_n1747_));
  AOI21_X1   g01554(.A1(new_n1679_), .A2(new_n1661_), .B(new_n1747_), .ZN(new_n1748_));
  AOI21_X1   g01555(.A1(new_n1636_), .A2(new_n1644_), .B(new_n1634_), .ZN(new_n1749_));
  INV_X1     g01556(.I(\a[27] ), .ZN(new_n1750_));
  NOR2_X1    g01557(.A1(new_n194_), .A2(new_n1750_), .ZN(new_n1751_));
  INV_X1     g01558(.I(new_n1751_), .ZN(new_n1752_));
  NOR2_X1    g01559(.A1(new_n1752_), .A2(new_n836_), .ZN(new_n1753_));
  NOR2_X1    g01560(.A1(new_n1751_), .A2(new_n1101_), .ZN(new_n1754_));
  NOR2_X1    g01561(.A1(new_n1753_), .A2(new_n1754_), .ZN(new_n1755_));
  XOR2_X1    g01562(.A1(new_n1755_), .A2(new_n1656_), .Z(new_n1756_));
  XNOR2_X1   g01563(.A1(new_n1756_), .A2(new_n1675_), .ZN(new_n1757_));
  XNOR2_X1   g01564(.A1(new_n1757_), .A2(new_n1749_), .ZN(new_n1758_));
  INV_X1     g01565(.I(new_n1758_), .ZN(new_n1759_));
  NAND2_X1   g01566(.A1(new_n1759_), .A2(new_n1748_), .ZN(new_n1760_));
  NOR2_X1    g01567(.A1(new_n1759_), .A2(new_n1748_), .ZN(new_n1761_));
  INV_X1     g01568(.I(new_n1761_), .ZN(new_n1762_));
  AND2_X2    g01569(.A1(new_n1762_), .A2(new_n1760_), .Z(new_n1763_));
  NAND2_X1   g01570(.A1(new_n1684_), .A2(new_n1686_), .ZN(new_n1764_));
  NAND2_X1   g01571(.A1(new_n1687_), .A2(new_n1681_), .ZN(new_n1765_));
  NAND2_X1   g01572(.A1(new_n1765_), .A2(new_n1764_), .ZN(new_n1766_));
  NOR2_X1    g01573(.A1(new_n1175_), .A2(new_n1299_), .ZN(new_n1767_));
  NAND2_X1   g01574(.A1(new_n1300_), .A2(new_n969_), .ZN(new_n1768_));
  NAND2_X1   g01575(.A1(new_n1452_), .A2(new_n479_), .ZN(new_n1769_));
  AOI22_X1   g01576(.A1(new_n1768_), .A2(new_n1769_), .B1(new_n746_), .B2(new_n1767_), .ZN(new_n1770_));
  NAND2_X1   g01577(.A1(\a[7] ), .A2(\a[21] ), .ZN(new_n1771_));
  AOI22_X1   g01578(.A1(\a[5] ), .A2(\a[23] ), .B1(\a[6] ), .B2(\a[22] ), .ZN(new_n1772_));
  NAND2_X1   g01579(.A1(new_n1767_), .A2(new_n746_), .ZN(new_n1773_));
  NAND3_X1   g01580(.A1(new_n1773_), .A2(new_n1768_), .A3(new_n1769_), .ZN(new_n1774_));
  OAI22_X1   g01581(.A1(new_n1770_), .A2(new_n1771_), .B1(new_n1774_), .B2(new_n1772_), .ZN(new_n1775_));
  AOI22_X1   g01582(.A1(\a[3] ), .A2(\a[25] ), .B1(\a[4] ), .B2(\a[24] ), .ZN(new_n1776_));
  INV_X1     g01583(.I(new_n1776_), .ZN(new_n1777_));
  NOR2_X1    g01584(.A1(new_n1357_), .A2(new_n1441_), .ZN(new_n1778_));
  INV_X1     g01585(.I(new_n1778_), .ZN(new_n1779_));
  NOR2_X1    g01586(.A1(new_n1779_), .A2(new_n370_), .ZN(new_n1780_));
  NOR2_X1    g01587(.A1(new_n355_), .A2(new_n1043_), .ZN(new_n1781_));
  AOI21_X1   g01588(.A1(new_n1777_), .A2(new_n1781_), .B(new_n1780_), .ZN(new_n1782_));
  INV_X1     g01589(.I(new_n1782_), .ZN(new_n1783_));
  OAI21_X1   g01590(.A1(new_n1780_), .A2(new_n1776_), .B(new_n1781_), .ZN(new_n1784_));
  OAI21_X1   g01591(.A1(new_n1783_), .A2(new_n1776_), .B(new_n1784_), .ZN(new_n1785_));
  NOR2_X1    g01592(.A1(new_n1660_), .A2(new_n1658_), .ZN(new_n1786_));
  NOR2_X1    g01593(.A1(new_n1592_), .A2(new_n1659_), .ZN(new_n1787_));
  NOR2_X1    g01594(.A1(new_n1786_), .A2(new_n1787_), .ZN(new_n1788_));
  XOR2_X1    g01595(.A1(new_n1788_), .A2(new_n1785_), .Z(new_n1789_));
  XNOR2_X1   g01596(.A1(new_n1789_), .A2(new_n1775_), .ZN(new_n1790_));
  XOR2_X1    g01597(.A1(new_n1766_), .A2(new_n1790_), .Z(new_n1791_));
  XOR2_X1    g01598(.A1(new_n1791_), .A2(new_n1763_), .Z(new_n1792_));
  INV_X1     g01599(.I(new_n1792_), .ZN(new_n1793_));
  NOR2_X1    g01600(.A1(new_n1745_), .A2(new_n1793_), .ZN(new_n1794_));
  INV_X1     g01601(.I(new_n1794_), .ZN(new_n1795_));
  NAND2_X1   g01602(.A1(new_n1745_), .A2(new_n1793_), .ZN(new_n1796_));
  NAND2_X1   g01603(.A1(new_n1795_), .A2(new_n1796_), .ZN(new_n1797_));
  XOR2_X1    g01604(.A1(new_n1700_), .A2(new_n1797_), .Z(\asquared[29] ));
  OAI21_X1   g01605(.A1(new_n1699_), .A2(new_n1696_), .B(new_n1796_), .ZN(new_n1799_));
  NAND2_X1   g01606(.A1(new_n1799_), .A2(new_n1795_), .ZN(new_n1800_));
  NAND3_X1   g01607(.A1(new_n1702_), .A2(new_n1743_), .A3(new_n1741_), .ZN(new_n1801_));
  NAND2_X1   g01608(.A1(new_n1801_), .A2(new_n1743_), .ZN(new_n1802_));
  INV_X1     g01609(.I(new_n1802_), .ZN(new_n1803_));
  NAND2_X1   g01610(.A1(new_n1733_), .A2(new_n1738_), .ZN(new_n1804_));
  NAND2_X1   g01611(.A1(new_n1739_), .A2(new_n1730_), .ZN(new_n1805_));
  NAND2_X1   g01612(.A1(new_n1805_), .A2(new_n1804_), .ZN(new_n1806_));
  INV_X1     g01613(.I(new_n1757_), .ZN(new_n1807_));
  NOR2_X1    g01614(.A1(new_n1749_), .A2(new_n1807_), .ZN(new_n1808_));
  NOR2_X1    g01615(.A1(new_n1761_), .A2(new_n1808_), .ZN(new_n1809_));
  XNOR2_X1   g01616(.A1(new_n1806_), .A2(new_n1809_), .ZN(new_n1810_));
  XOR2_X1    g01617(.A1(new_n1726_), .A2(new_n1715_), .Z(new_n1811_));
  INV_X1     g01618(.I(new_n1753_), .ZN(new_n1812_));
  AOI22_X1   g01619(.A1(\a[0] ), .A2(\a[29] ), .B1(\a[2] ), .B2(\a[27] ), .ZN(new_n1813_));
  INV_X1     g01620(.I(\a[29] ), .ZN(new_n1814_));
  NOR2_X1    g01621(.A1(new_n1750_), .A2(new_n1814_), .ZN(new_n1815_));
  INV_X1     g01622(.I(new_n1815_), .ZN(new_n1816_));
  NOR2_X1    g01623(.A1(new_n1816_), .A2(new_n412_), .ZN(new_n1817_));
  NOR3_X1    g01624(.A1(new_n1812_), .A2(new_n1817_), .A3(new_n1813_), .ZN(new_n1818_));
  NOR2_X1    g01625(.A1(new_n1818_), .A2(new_n1817_), .ZN(new_n1819_));
  INV_X1     g01626(.I(new_n1819_), .ZN(new_n1820_));
  OAI22_X1   g01627(.A1(new_n1820_), .A2(new_n1813_), .B1(new_n1818_), .B2(new_n1812_), .ZN(new_n1821_));
  XNOR2_X1   g01628(.A1(new_n1821_), .A2(new_n1811_), .ZN(new_n1822_));
  INV_X1     g01629(.I(new_n1822_), .ZN(new_n1823_));
  NAND2_X1   g01630(.A1(new_n1728_), .A2(new_n1716_), .ZN(new_n1824_));
  INV_X1     g01631(.I(new_n1729_), .ZN(new_n1825_));
  NAND2_X1   g01632(.A1(new_n1825_), .A2(new_n1708_), .ZN(new_n1826_));
  NAND2_X1   g01633(.A1(new_n1826_), .A2(new_n1824_), .ZN(new_n1827_));
  INV_X1     g01634(.I(new_n1785_), .ZN(new_n1828_));
  INV_X1     g01635(.I(new_n1789_), .ZN(new_n1829_));
  NAND2_X1   g01636(.A1(new_n1829_), .A2(new_n1775_), .ZN(new_n1830_));
  OAI21_X1   g01637(.A1(new_n1828_), .A2(new_n1788_), .B(new_n1830_), .ZN(new_n1831_));
  NOR2_X1    g01638(.A1(new_n1831_), .A2(new_n1827_), .ZN(new_n1832_));
  NAND2_X1   g01639(.A1(new_n1831_), .A2(new_n1827_), .ZN(new_n1833_));
  INV_X1     g01640(.I(new_n1833_), .ZN(new_n1834_));
  NOR2_X1    g01641(.A1(new_n1834_), .A2(new_n1832_), .ZN(new_n1835_));
  NAND2_X1   g01642(.A1(new_n1835_), .A2(new_n1823_), .ZN(new_n1836_));
  INV_X1     g01643(.I(new_n1836_), .ZN(new_n1837_));
  NOR2_X1    g01644(.A1(new_n1835_), .A2(new_n1823_), .ZN(new_n1838_));
  NOR2_X1    g01645(.A1(new_n1837_), .A2(new_n1838_), .ZN(new_n1839_));
  XNOR2_X1   g01646(.A1(new_n1810_), .A2(new_n1839_), .ZN(new_n1840_));
  NAND2_X1   g01647(.A1(new_n1766_), .A2(new_n1790_), .ZN(new_n1841_));
  NAND2_X1   g01648(.A1(new_n1791_), .A2(new_n1763_), .ZN(new_n1842_));
  NAND2_X1   g01649(.A1(new_n1842_), .A2(new_n1841_), .ZN(new_n1843_));
  NAND2_X1   g01650(.A1(new_n1669_), .A2(new_n1643_), .ZN(new_n1844_));
  NAND2_X1   g01651(.A1(new_n1737_), .A2(new_n1736_), .ZN(new_n1845_));
  NAND2_X1   g01652(.A1(new_n1845_), .A2(new_n1844_), .ZN(new_n1846_));
  NAND2_X1   g01653(.A1(new_n1755_), .A2(new_n1655_), .ZN(new_n1847_));
  INV_X1     g01654(.I(new_n1756_), .ZN(new_n1848_));
  NAND2_X1   g01655(.A1(new_n1848_), .A2(new_n1675_), .ZN(new_n1849_));
  NAND2_X1   g01656(.A1(new_n1849_), .A2(new_n1847_), .ZN(new_n1850_));
  NOR2_X1    g01657(.A1(new_n367_), .A2(new_n1299_), .ZN(new_n1851_));
  INV_X1     g01658(.I(new_n1851_), .ZN(new_n1852_));
  AOI21_X1   g01659(.A1(\a[13] ), .A2(\a[16] ), .B(new_n897_), .ZN(new_n1853_));
  NOR3_X1    g01660(.A1(new_n1173_), .A2(new_n597_), .A3(new_n742_), .ZN(new_n1854_));
  NOR3_X1    g01661(.A1(new_n1854_), .A2(new_n1852_), .A3(new_n1853_), .ZN(new_n1855_));
  NOR2_X1    g01662(.A1(new_n1855_), .A2(new_n1854_), .ZN(new_n1856_));
  INV_X1     g01663(.I(new_n1856_), .ZN(new_n1857_));
  OAI22_X1   g01664(.A1(new_n1857_), .A2(new_n1853_), .B1(new_n1852_), .B2(new_n1855_), .ZN(new_n1858_));
  XNOR2_X1   g01665(.A1(new_n1850_), .A2(new_n1858_), .ZN(new_n1859_));
  XOR2_X1    g01666(.A1(new_n1859_), .A2(new_n1846_), .Z(new_n1860_));
  OAI22_X1   g01667(.A1(new_n1063_), .A2(new_n1281_), .B1(new_n1376_), .B2(new_n539_), .ZN(new_n1861_));
  OAI21_X1   g01668(.A1(new_n1264_), .A2(new_n1092_), .B(new_n1861_), .ZN(new_n1862_));
  NAND3_X1   g01669(.A1(new_n1862_), .A2(\a[9] ), .A3(\a[20] ), .ZN(new_n1863_));
  AOI22_X1   g01670(.A1(\a[10] ), .A2(\a[19] ), .B1(\a[11] ), .B2(\a[18] ), .ZN(new_n1864_));
  NOR2_X1    g01671(.A1(new_n1264_), .A2(new_n1092_), .ZN(new_n1865_));
  NOR2_X1    g01672(.A1(new_n1861_), .A2(new_n1865_), .ZN(new_n1866_));
  INV_X1     g01673(.I(new_n1866_), .ZN(new_n1867_));
  OAI21_X1   g01674(.A1(new_n1864_), .A2(new_n1867_), .B(new_n1863_), .ZN(new_n1868_));
  AOI22_X1   g01675(.A1(\a[3] ), .A2(\a[26] ), .B1(\a[8] ), .B2(\a[21] ), .ZN(new_n1869_));
  NOR4_X1    g01676(.A1(new_n225_), .A2(new_n355_), .A3(new_n1220_), .A4(new_n1566_), .ZN(new_n1870_));
  NOR3_X1    g01677(.A1(new_n1869_), .A2(new_n536_), .A3(new_n1023_), .ZN(new_n1871_));
  NOR2_X1    g01678(.A1(new_n1871_), .A2(new_n1870_), .ZN(new_n1872_));
  INV_X1     g01679(.I(new_n1872_), .ZN(new_n1873_));
  NOR2_X1    g01680(.A1(new_n536_), .A2(new_n1023_), .ZN(new_n1874_));
  OAI21_X1   g01681(.A1(new_n1870_), .A2(new_n1869_), .B(new_n1874_), .ZN(new_n1875_));
  OAI21_X1   g01682(.A1(new_n1873_), .A2(new_n1869_), .B(new_n1875_), .ZN(new_n1876_));
  XNOR2_X1   g01683(.A1(new_n1868_), .A2(new_n1876_), .ZN(new_n1877_));
  NAND2_X1   g01684(.A1(\a[4] ), .A2(\a[25] ), .ZN(new_n1878_));
  NOR2_X1    g01685(.A1(new_n1175_), .A2(new_n1357_), .ZN(new_n1879_));
  INV_X1     g01686(.I(new_n1879_), .ZN(new_n1880_));
  NOR2_X1    g01687(.A1(new_n1880_), .A2(new_n373_), .ZN(new_n1881_));
  NAND4_X1   g01688(.A1(\a[4] ), .A2(\a[7] ), .A3(\a[22] ), .A4(\a[25] ), .ZN(new_n1882_));
  NAND2_X1   g01689(.A1(new_n1778_), .A2(new_n243_), .ZN(new_n1883_));
  AOI21_X1   g01690(.A1(new_n1882_), .A2(new_n1883_), .B(new_n1881_), .ZN(new_n1884_));
  AOI22_X1   g01691(.A1(\a[5] ), .A2(\a[24] ), .B1(\a[7] ), .B2(\a[22] ), .ZN(new_n1885_));
  NOR2_X1    g01692(.A1(new_n1884_), .A2(new_n1881_), .ZN(new_n1886_));
  INV_X1     g01693(.I(new_n1886_), .ZN(new_n1887_));
  OAI22_X1   g01694(.A1(new_n1887_), .A2(new_n1885_), .B1(new_n1878_), .B2(new_n1884_), .ZN(new_n1888_));
  XOR2_X1    g01695(.A1(new_n1877_), .A2(new_n1888_), .Z(new_n1889_));
  NOR2_X1    g01696(.A1(new_n194_), .A2(new_n1718_), .ZN(new_n1890_));
  NOR2_X1    g01697(.A1(new_n774_), .A2(new_n1718_), .ZN(new_n1891_));
  INV_X1     g01698(.I(new_n1891_), .ZN(new_n1892_));
  OAI21_X1   g01699(.A1(\a[15] ), .A2(new_n1890_), .B(new_n1892_), .ZN(new_n1893_));
  XNOR2_X1   g01700(.A1(new_n1774_), .A2(new_n1893_), .ZN(new_n1894_));
  XOR2_X1    g01701(.A1(new_n1894_), .A2(new_n1783_), .Z(new_n1895_));
  INV_X1     g01702(.I(new_n1895_), .ZN(new_n1896_));
  XOR2_X1    g01703(.A1(new_n1889_), .A2(new_n1896_), .Z(new_n1897_));
  XNOR2_X1   g01704(.A1(new_n1897_), .A2(new_n1860_), .ZN(new_n1898_));
  INV_X1     g01705(.I(new_n1898_), .ZN(new_n1899_));
  NAND2_X1   g01706(.A1(new_n1843_), .A2(new_n1899_), .ZN(new_n1900_));
  NOR2_X1    g01707(.A1(new_n1843_), .A2(new_n1899_), .ZN(new_n1901_));
  INV_X1     g01708(.I(new_n1901_), .ZN(new_n1902_));
  AOI21_X1   g01709(.A1(new_n1902_), .A2(new_n1900_), .B(new_n1840_), .ZN(new_n1903_));
  INV_X1     g01710(.I(new_n1903_), .ZN(new_n1904_));
  NAND3_X1   g01711(.A1(new_n1840_), .A2(new_n1902_), .A3(new_n1900_), .ZN(new_n1905_));
  NAND2_X1   g01712(.A1(new_n1904_), .A2(new_n1905_), .ZN(new_n1906_));
  NOR2_X1    g01713(.A1(new_n1906_), .A2(new_n1803_), .ZN(new_n1907_));
  AOI21_X1   g01714(.A1(new_n1904_), .A2(new_n1905_), .B(new_n1802_), .ZN(new_n1908_));
  NOR2_X1    g01715(.A1(new_n1907_), .A2(new_n1908_), .ZN(new_n1909_));
  XOR2_X1    g01716(.A1(new_n1800_), .A2(new_n1909_), .Z(\asquared[30] ));
  AOI21_X1   g01717(.A1(new_n1799_), .A2(new_n1795_), .B(new_n1908_), .ZN(new_n1911_));
  NOR2_X1    g01718(.A1(new_n1911_), .A2(new_n1907_), .ZN(new_n1912_));
  NAND2_X1   g01719(.A1(new_n1843_), .A2(new_n1898_), .ZN(new_n1913_));
  NAND2_X1   g01720(.A1(new_n1904_), .A2(new_n1913_), .ZN(new_n1914_));
  XOR2_X1    g01721(.A1(new_n1866_), .A2(new_n1872_), .Z(new_n1915_));
  XOR2_X1    g01722(.A1(new_n1915_), .A2(new_n1820_), .Z(new_n1916_));
  XOR2_X1    g01723(.A1(new_n1886_), .A2(new_n1856_), .Z(new_n1917_));
  NOR2_X1    g01724(.A1(new_n597_), .A2(new_n1023_), .ZN(new_n1918_));
  INV_X1     g01725(.I(new_n1918_), .ZN(new_n1919_));
  AOI22_X1   g01726(.A1(\a[2] ), .A2(\a[28] ), .B1(\a[9] ), .B2(\a[21] ), .ZN(new_n1920_));
  NOR4_X1    g01727(.A1(new_n197_), .A2(new_n403_), .A3(new_n1220_), .A4(new_n1718_), .ZN(new_n1921_));
  NOR3_X1    g01728(.A1(new_n1919_), .A2(new_n1921_), .A3(new_n1920_), .ZN(new_n1922_));
  NOR2_X1    g01729(.A1(new_n1922_), .A2(new_n1921_), .ZN(new_n1923_));
  INV_X1     g01730(.I(new_n1923_), .ZN(new_n1924_));
  OAI22_X1   g01731(.A1(new_n1924_), .A2(new_n1920_), .B1(new_n1919_), .B2(new_n1922_), .ZN(new_n1925_));
  XOR2_X1    g01732(.A1(new_n1917_), .A2(new_n1925_), .Z(new_n1926_));
  NAND2_X1   g01733(.A1(new_n1868_), .A2(new_n1876_), .ZN(new_n1927_));
  INV_X1     g01734(.I(new_n1877_), .ZN(new_n1928_));
  NAND2_X1   g01735(.A1(new_n1928_), .A2(new_n1888_), .ZN(new_n1929_));
  NAND2_X1   g01736(.A1(new_n1929_), .A2(new_n1927_), .ZN(new_n1930_));
  XOR2_X1    g01737(.A1(new_n1930_), .A2(new_n1926_), .Z(new_n1931_));
  XOR2_X1    g01738(.A1(new_n1931_), .A2(new_n1916_), .Z(new_n1932_));
  NOR2_X1    g01739(.A1(new_n1889_), .A2(new_n1896_), .ZN(new_n1933_));
  INV_X1     g01740(.I(new_n1897_), .ZN(new_n1934_));
  NOR2_X1    g01741(.A1(new_n1934_), .A2(new_n1860_), .ZN(new_n1935_));
  NOR2_X1    g01742(.A1(new_n1935_), .A2(new_n1933_), .ZN(new_n1936_));
  NAND2_X1   g01743(.A1(new_n1726_), .A2(new_n1715_), .ZN(new_n1937_));
  NAND2_X1   g01744(.A1(new_n1821_), .A2(new_n1811_), .ZN(new_n1938_));
  NAND2_X1   g01745(.A1(new_n1938_), .A2(new_n1937_), .ZN(new_n1939_));
  INV_X1     g01746(.I(new_n1893_), .ZN(new_n1940_));
  NAND2_X1   g01747(.A1(new_n1940_), .A2(new_n1774_), .ZN(new_n1941_));
  NAND2_X1   g01748(.A1(new_n1894_), .A2(new_n1783_), .ZN(new_n1942_));
  NAND2_X1   g01749(.A1(new_n1942_), .A2(new_n1941_), .ZN(new_n1943_));
  NAND2_X1   g01750(.A1(\a[0] ), .A2(\a[30] ), .ZN(new_n1944_));
  XOR2_X1    g01751(.A1(new_n1891_), .A2(new_n1944_), .Z(new_n1945_));
  NOR2_X1    g01752(.A1(new_n194_), .A2(new_n1814_), .ZN(new_n1946_));
  XNOR2_X1   g01753(.A1(new_n895_), .A2(new_n1946_), .ZN(new_n1947_));
  XOR2_X1    g01754(.A1(new_n1947_), .A2(new_n1945_), .Z(new_n1948_));
  NOR2_X1    g01755(.A1(new_n1943_), .A2(new_n1948_), .ZN(new_n1949_));
  NAND2_X1   g01756(.A1(new_n1943_), .A2(new_n1948_), .ZN(new_n1950_));
  INV_X1     g01757(.I(new_n1950_), .ZN(new_n1951_));
  NOR2_X1    g01758(.A1(new_n1951_), .A2(new_n1949_), .ZN(new_n1952_));
  NOR2_X1    g01759(.A1(new_n1952_), .A2(new_n1939_), .ZN(new_n1953_));
  NAND2_X1   g01760(.A1(new_n1952_), .A2(new_n1939_), .ZN(new_n1954_));
  INV_X1     g01761(.I(new_n1954_), .ZN(new_n1955_));
  NOR2_X1    g01762(.A1(new_n1955_), .A2(new_n1953_), .ZN(new_n1956_));
  INV_X1     g01763(.I(new_n1956_), .ZN(new_n1957_));
  XOR2_X1    g01764(.A1(new_n1936_), .A2(new_n1957_), .Z(new_n1958_));
  NOR2_X1    g01765(.A1(new_n1958_), .A2(new_n1932_), .ZN(new_n1959_));
  AND2_X2    g01766(.A1(new_n1958_), .A2(new_n1932_), .Z(new_n1960_));
  NOR2_X1    g01767(.A1(new_n1960_), .A2(new_n1959_), .ZN(new_n1961_));
  OAI21_X1   g01768(.A1(new_n1808_), .A2(new_n1761_), .B(new_n1806_), .ZN(new_n1962_));
  NAND2_X1   g01769(.A1(new_n1810_), .A2(new_n1839_), .ZN(new_n1963_));
  NAND2_X1   g01770(.A1(new_n1963_), .A2(new_n1962_), .ZN(new_n1964_));
  NOR2_X1    g01771(.A1(new_n1837_), .A2(new_n1834_), .ZN(new_n1965_));
  NAND2_X1   g01772(.A1(new_n1850_), .A2(new_n1858_), .ZN(new_n1966_));
  INV_X1     g01773(.I(new_n1859_), .ZN(new_n1967_));
  NAND2_X1   g01774(.A1(new_n1967_), .A2(new_n1846_), .ZN(new_n1968_));
  NAND2_X1   g01775(.A1(new_n1968_), .A2(new_n1966_), .ZN(new_n1969_));
  NOR4_X1    g01776(.A1(new_n225_), .A2(new_n355_), .A3(new_n1175_), .A4(new_n1750_), .ZN(new_n1970_));
  NOR2_X1    g01777(.A1(new_n1566_), .A2(new_n1750_), .ZN(new_n1971_));
  INV_X1     g01778(.I(new_n1971_), .ZN(new_n1972_));
  NOR2_X1    g01779(.A1(new_n1972_), .A2(new_n370_), .ZN(new_n1973_));
  NOR2_X1    g01780(.A1(new_n290_), .A2(new_n1566_), .ZN(new_n1974_));
  NAND3_X1   g01781(.A1(new_n1974_), .A2(\a[8] ), .A3(\a[22] ), .ZN(new_n1975_));
  OAI21_X1   g01782(.A1(new_n1973_), .A2(new_n1970_), .B(new_n1975_), .ZN(new_n1976_));
  NAND3_X1   g01783(.A1(new_n1976_), .A2(\a[3] ), .A3(\a[27] ), .ZN(new_n1977_));
  AOI21_X1   g01784(.A1(\a[8] ), .A2(\a[22] ), .B(new_n1974_), .ZN(new_n1978_));
  NAND2_X1   g01785(.A1(new_n1976_), .A2(new_n1975_), .ZN(new_n1979_));
  OAI21_X1   g01786(.A1(new_n1978_), .A2(new_n1979_), .B(new_n1977_), .ZN(new_n1980_));
  NAND2_X1   g01787(.A1(new_n1528_), .A2(new_n479_), .ZN(new_n1981_));
  OAI22_X1   g01788(.A1(new_n373_), .A2(new_n1443_), .B1(new_n1779_), .B2(new_n371_), .ZN(new_n1982_));
  NAND2_X1   g01789(.A1(new_n1982_), .A2(new_n1981_), .ZN(new_n1983_));
  NAND3_X1   g01790(.A1(new_n1983_), .A2(\a[5] ), .A3(\a[25] ), .ZN(new_n1984_));
  AOI22_X1   g01791(.A1(\a[6] ), .A2(\a[24] ), .B1(\a[7] ), .B2(\a[23] ), .ZN(new_n1985_));
  NAND2_X1   g01792(.A1(new_n1983_), .A2(new_n1981_), .ZN(new_n1986_));
  OAI21_X1   g01793(.A1(new_n1985_), .A2(new_n1986_), .B(new_n1984_), .ZN(new_n1987_));
  XNOR2_X1   g01794(.A1(new_n1987_), .A2(new_n1980_), .ZN(new_n1988_));
  NAND2_X1   g01795(.A1(new_n1273_), .A2(new_n535_), .ZN(new_n1989_));
  NAND2_X1   g01796(.A1(new_n747_), .A2(new_n1375_), .ZN(new_n1990_));
  AOI22_X1   g01797(.A1(new_n1990_), .A2(new_n1989_), .B1(new_n1261_), .B2(new_n1194_), .ZN(new_n1991_));
  NAND2_X1   g01798(.A1(\a[10] ), .A2(\a[20] ), .ZN(new_n1992_));
  AOI22_X1   g01799(.A1(\a[11] ), .A2(\a[19] ), .B1(\a[12] ), .B2(\a[18] ), .ZN(new_n1993_));
  NAND2_X1   g01800(.A1(new_n1261_), .A2(new_n1194_), .ZN(new_n1994_));
  NAND3_X1   g01801(.A1(new_n1989_), .A2(new_n1990_), .A3(new_n1994_), .ZN(new_n1995_));
  OAI22_X1   g01802(.A1(new_n1991_), .A2(new_n1992_), .B1(new_n1995_), .B2(new_n1993_), .ZN(new_n1996_));
  XOR2_X1    g01803(.A1(new_n1988_), .A2(new_n1996_), .Z(new_n1997_));
  INV_X1     g01804(.I(new_n1997_), .ZN(new_n1998_));
  XOR2_X1    g01805(.A1(new_n1969_), .A2(new_n1998_), .Z(new_n1999_));
  INV_X1     g01806(.I(new_n1999_), .ZN(new_n2000_));
  XOR2_X1    g01807(.A1(new_n1965_), .A2(new_n2000_), .Z(new_n2001_));
  XOR2_X1    g01808(.A1(new_n1964_), .A2(new_n2001_), .Z(new_n2002_));
  XOR2_X1    g01809(.A1(new_n2002_), .A2(new_n1961_), .Z(new_n2003_));
  NOR2_X1    g01810(.A1(new_n2003_), .A2(new_n1914_), .ZN(new_n2004_));
  INV_X1     g01811(.I(new_n2004_), .ZN(new_n2005_));
  NAND2_X1   g01812(.A1(new_n2003_), .A2(new_n1914_), .ZN(new_n2006_));
  NAND2_X1   g01813(.A1(new_n2005_), .A2(new_n2006_), .ZN(new_n2007_));
  XOR2_X1    g01814(.A1(new_n1912_), .A2(new_n2007_), .Z(\asquared[31] ));
  OAI21_X1   g01815(.A1(new_n1911_), .A2(new_n1907_), .B(new_n2005_), .ZN(new_n2009_));
  NAND2_X1   g01816(.A1(new_n2009_), .A2(new_n2006_), .ZN(new_n2010_));
  NOR2_X1    g01817(.A1(new_n1955_), .A2(new_n1951_), .ZN(new_n2011_));
  XOR2_X1    g01818(.A1(new_n1979_), .A2(new_n1924_), .Z(new_n2012_));
  XOR2_X1    g01819(.A1(new_n2012_), .A2(new_n1995_), .Z(new_n2013_));
  NAND2_X1   g01820(.A1(new_n1987_), .A2(new_n1980_), .ZN(new_n2014_));
  INV_X1     g01821(.I(new_n1996_), .ZN(new_n2015_));
  OAI21_X1   g01822(.A1(new_n1988_), .A2(new_n2015_), .B(new_n2014_), .ZN(new_n2016_));
  NAND2_X1   g01823(.A1(new_n2016_), .A2(new_n2013_), .ZN(new_n2017_));
  INV_X1     g01824(.I(new_n2017_), .ZN(new_n2018_));
  NOR2_X1    g01825(.A1(new_n2016_), .A2(new_n2013_), .ZN(new_n2019_));
  NOR2_X1    g01826(.A1(new_n2018_), .A2(new_n2019_), .ZN(new_n2020_));
  INV_X1     g01827(.I(new_n2020_), .ZN(new_n2021_));
  NAND2_X1   g01828(.A1(new_n2021_), .A2(new_n2011_), .ZN(new_n2022_));
  NOR2_X1    g01829(.A1(new_n2021_), .A2(new_n2011_), .ZN(new_n2023_));
  INV_X1     g01830(.I(new_n2023_), .ZN(new_n2024_));
  AND2_X2    g01831(.A1(new_n2024_), .A2(new_n2022_), .Z(new_n2025_));
  NAND2_X1   g01832(.A1(new_n1969_), .A2(new_n1998_), .ZN(new_n2026_));
  OAI21_X1   g01833(.A1(new_n1965_), .A2(new_n2000_), .B(new_n2026_), .ZN(new_n2027_));
  INV_X1     g01834(.I(new_n895_), .ZN(new_n2028_));
  NOR3_X1    g01835(.A1(new_n2028_), .A2(new_n194_), .A3(new_n1814_), .ZN(new_n2029_));
  INV_X1     g01836(.I(\a[30] ), .ZN(new_n2030_));
  NOR2_X1    g01837(.A1(new_n194_), .A2(new_n2030_), .ZN(new_n2031_));
  INV_X1     g01838(.I(new_n2031_), .ZN(new_n2032_));
  NOR2_X1    g01839(.A1(new_n2032_), .A2(new_n742_), .ZN(new_n2033_));
  NOR2_X1    g01840(.A1(new_n2031_), .A2(\a[16] ), .ZN(new_n2034_));
  NOR2_X1    g01841(.A1(new_n2033_), .A2(new_n2034_), .ZN(new_n2035_));
  XOR2_X1    g01842(.A1(new_n2035_), .A2(new_n2029_), .Z(new_n2036_));
  XOR2_X1    g01843(.A1(new_n2036_), .A2(new_n1986_), .Z(new_n2037_));
  NAND2_X1   g01844(.A1(new_n1917_), .A2(new_n1925_), .ZN(new_n2038_));
  OAI21_X1   g01845(.A1(new_n1856_), .A2(new_n1886_), .B(new_n2038_), .ZN(new_n2039_));
  NAND2_X1   g01846(.A1(new_n1915_), .A2(new_n1820_), .ZN(new_n2040_));
  OAI21_X1   g01847(.A1(new_n1866_), .A2(new_n1872_), .B(new_n2040_), .ZN(new_n2041_));
  XOR2_X1    g01848(.A1(new_n2039_), .A2(new_n2041_), .Z(new_n2042_));
  XOR2_X1    g01849(.A1(new_n2042_), .A2(new_n2037_), .Z(new_n2043_));
  XOR2_X1    g01850(.A1(new_n2027_), .A2(new_n2043_), .Z(new_n2044_));
  XOR2_X1    g01851(.A1(new_n2044_), .A2(new_n2025_), .Z(new_n2045_));
  NOR2_X1    g01852(.A1(new_n1936_), .A2(new_n1957_), .ZN(new_n2046_));
  NOR2_X1    g01853(.A1(new_n1960_), .A2(new_n2046_), .ZN(new_n2047_));
  NAND2_X1   g01854(.A1(new_n1930_), .A2(new_n1926_), .ZN(new_n2048_));
  NAND2_X1   g01855(.A1(new_n1931_), .A2(new_n1916_), .ZN(new_n2049_));
  NAND2_X1   g01856(.A1(new_n2049_), .A2(new_n2048_), .ZN(new_n2050_));
  INV_X1     g01857(.I(\a[31] ), .ZN(new_n2051_));
  NOR2_X1    g01858(.A1(new_n1175_), .A2(new_n2051_), .ZN(new_n2052_));
  INV_X1     g01859(.I(new_n2052_), .ZN(new_n2053_));
  NOR2_X1    g01860(.A1(new_n2053_), .A2(new_n359_), .ZN(new_n2054_));
  NOR2_X1    g01861(.A1(new_n417_), .A2(new_n2051_), .ZN(new_n2055_));
  AOI22_X1   g01862(.A1(new_n540_), .A2(new_n1452_), .B1(new_n2055_), .B2(new_n1140_), .ZN(new_n2056_));
  NOR2_X1    g01863(.A1(new_n2054_), .A2(new_n2056_), .ZN(new_n2057_));
  NAND2_X1   g01864(.A1(\a[10] ), .A2(\a[21] ), .ZN(new_n2058_));
  OAI21_X1   g01865(.A1(new_n359_), .A2(new_n2053_), .B(new_n2056_), .ZN(new_n2059_));
  AOI22_X1   g01866(.A1(\a[0] ), .A2(\a[31] ), .B1(\a[9] ), .B2(\a[22] ), .ZN(new_n2060_));
  OAI22_X1   g01867(.A1(new_n2059_), .A2(new_n2060_), .B1(new_n2057_), .B2(new_n2058_), .ZN(new_n2061_));
  NOR2_X1    g01868(.A1(new_n1892_), .A2(new_n1944_), .ZN(new_n2062_));
  NOR2_X1    g01869(.A1(new_n1947_), .A2(new_n1945_), .ZN(new_n2063_));
  NOR2_X1    g01870(.A1(new_n2063_), .A2(new_n2062_), .ZN(new_n2064_));
  NAND2_X1   g01871(.A1(new_n1273_), .A2(new_n834_), .ZN(new_n2065_));
  NAND2_X1   g01872(.A1(new_n1375_), .A2(new_n1261_), .ZN(new_n2066_));
  AOI22_X1   g01873(.A1(new_n2065_), .A2(new_n2066_), .B1(new_n763_), .B2(new_n1194_), .ZN(new_n2067_));
  NOR3_X1    g01874(.A1(new_n2067_), .A2(new_n513_), .A3(new_n1043_), .ZN(new_n2068_));
  AOI22_X1   g01875(.A1(\a[12] ), .A2(\a[19] ), .B1(\a[13] ), .B2(\a[18] ), .ZN(new_n2069_));
  NAND2_X1   g01876(.A1(new_n763_), .A2(new_n1194_), .ZN(new_n2070_));
  NAND3_X1   g01877(.A1(new_n2065_), .A2(new_n2066_), .A3(new_n2070_), .ZN(new_n2071_));
  NOR2_X1    g01878(.A1(new_n2071_), .A2(new_n2069_), .ZN(new_n2072_));
  NOR2_X1    g01879(.A1(new_n2068_), .A2(new_n2072_), .ZN(new_n2073_));
  NOR2_X1    g01880(.A1(new_n2073_), .A2(new_n2064_), .ZN(new_n2074_));
  NOR2_X1    g01881(.A1(new_n2074_), .A2(new_n2064_), .ZN(new_n2075_));
  NOR2_X1    g01882(.A1(new_n2074_), .A2(new_n2073_), .ZN(new_n2076_));
  OAI21_X1   g01883(.A1(new_n2075_), .A2(new_n2076_), .B(new_n2061_), .ZN(new_n2077_));
  OR3_X2     g01884(.A1(new_n2075_), .A2(new_n2076_), .A3(new_n2061_), .Z(new_n2078_));
  NAND2_X1   g01885(.A1(new_n2078_), .A2(new_n2077_), .ZN(new_n2079_));
  NOR2_X1    g01886(.A1(new_n1357_), .A2(new_n1566_), .ZN(new_n2080_));
  INV_X1     g01887(.I(new_n2080_), .ZN(new_n2081_));
  NOR2_X1    g01888(.A1(new_n2081_), .A2(new_n373_), .ZN(new_n2082_));
  NOR2_X1    g01889(.A1(new_n1299_), .A2(new_n1566_), .ZN(new_n2083_));
  INV_X1     g01890(.I(new_n2083_), .ZN(new_n2084_));
  NOR2_X1    g01891(.A1(new_n2084_), .A2(new_n352_), .ZN(new_n2085_));
  NOR2_X1    g01892(.A1(new_n1529_), .A2(new_n415_), .ZN(new_n2086_));
  NOR2_X1    g01893(.A1(new_n2085_), .A2(new_n2086_), .ZN(new_n2087_));
  NOR2_X1    g01894(.A1(new_n2087_), .A2(new_n2082_), .ZN(new_n2088_));
  NAND2_X1   g01895(.A1(\a[8] ), .A2(\a[23] ), .ZN(new_n2089_));
  AOI22_X1   g01896(.A1(\a[5] ), .A2(\a[26] ), .B1(\a[7] ), .B2(\a[24] ), .ZN(new_n2090_));
  NOR2_X1    g01897(.A1(new_n2088_), .A2(new_n2082_), .ZN(new_n2091_));
  INV_X1     g01898(.I(new_n2091_), .ZN(new_n2092_));
  OAI22_X1   g01899(.A1(new_n2092_), .A2(new_n2090_), .B1(new_n2088_), .B2(new_n2089_), .ZN(new_n2093_));
  AOI21_X1   g01900(.A1(\a[14] ), .A2(\a[17] ), .B(new_n1288_), .ZN(new_n2094_));
  INV_X1     g01901(.I(new_n2094_), .ZN(new_n2095_));
  NOR2_X1    g01902(.A1(new_n1173_), .A2(new_n1428_), .ZN(new_n2096_));
  NOR2_X1    g01903(.A1(new_n367_), .A2(new_n1441_), .ZN(new_n2097_));
  AOI21_X1   g01904(.A1(new_n2095_), .A2(new_n2097_), .B(new_n2096_), .ZN(new_n2098_));
  INV_X1     g01905(.I(new_n2098_), .ZN(new_n2099_));
  OAI21_X1   g01906(.A1(new_n2096_), .A2(new_n2094_), .B(new_n2097_), .ZN(new_n2100_));
  OAI21_X1   g01907(.A1(new_n2099_), .A2(new_n2094_), .B(new_n2100_), .ZN(new_n2101_));
  XOR2_X1    g01908(.A1(new_n2093_), .A2(new_n2101_), .Z(new_n2102_));
  NOR2_X1    g01909(.A1(new_n1750_), .A2(new_n1718_), .ZN(new_n2103_));
  NAND2_X1   g01910(.A1(new_n1815_), .A2(new_n252_), .ZN(new_n2104_));
  NOR2_X1    g01911(.A1(new_n1718_), .A2(new_n1814_), .ZN(new_n2105_));
  NAND2_X1   g01912(.A1(new_n2105_), .A2(new_n256_), .ZN(new_n2106_));
  AOI22_X1   g01913(.A1(new_n2104_), .A2(new_n2106_), .B1(new_n761_), .B2(new_n2103_), .ZN(new_n2107_));
  NAND2_X1   g01914(.A1(\a[2] ), .A2(\a[29] ), .ZN(new_n2108_));
  AOI22_X1   g01915(.A1(\a[3] ), .A2(\a[28] ), .B1(\a[4] ), .B2(\a[27] ), .ZN(new_n2109_));
  NAND2_X1   g01916(.A1(new_n2103_), .A2(new_n761_), .ZN(new_n2110_));
  NAND3_X1   g01917(.A1(new_n2110_), .A2(new_n2104_), .A3(new_n2106_), .ZN(new_n2111_));
  OAI22_X1   g01918(.A1(new_n2107_), .A2(new_n2108_), .B1(new_n2111_), .B2(new_n2109_), .ZN(new_n2112_));
  XNOR2_X1   g01919(.A1(new_n2102_), .A2(new_n2112_), .ZN(new_n2113_));
  XOR2_X1    g01920(.A1(new_n2113_), .A2(new_n2079_), .Z(new_n2114_));
  XNOR2_X1   g01921(.A1(new_n2050_), .A2(new_n2114_), .ZN(new_n2115_));
  XOR2_X1    g01922(.A1(new_n2047_), .A2(new_n2115_), .Z(new_n2116_));
  NAND2_X1   g01923(.A1(new_n2116_), .A2(new_n2045_), .ZN(new_n2117_));
  INV_X1     g01924(.I(new_n2117_), .ZN(new_n2118_));
  NOR2_X1    g01925(.A1(new_n2116_), .A2(new_n2045_), .ZN(new_n2119_));
  NOR2_X1    g01926(.A1(new_n2118_), .A2(new_n2119_), .ZN(new_n2120_));
  NAND2_X1   g01927(.A1(new_n1964_), .A2(new_n2001_), .ZN(new_n2121_));
  NAND2_X1   g01928(.A1(new_n2002_), .A2(new_n1961_), .ZN(new_n2122_));
  NAND2_X1   g01929(.A1(new_n2122_), .A2(new_n2121_), .ZN(new_n2123_));
  NAND2_X1   g01930(.A1(new_n2123_), .A2(new_n2120_), .ZN(new_n2124_));
  INV_X1     g01931(.I(new_n2124_), .ZN(new_n2125_));
  NOR2_X1    g01932(.A1(new_n2123_), .A2(new_n2120_), .ZN(new_n2126_));
  NOR2_X1    g01933(.A1(new_n2125_), .A2(new_n2126_), .ZN(new_n2127_));
  XOR2_X1    g01934(.A1(new_n2010_), .A2(new_n2127_), .Z(\asquared[32] ));
  AOI21_X1   g01935(.A1(new_n2009_), .A2(new_n2006_), .B(new_n2126_), .ZN(new_n2129_));
  NOR2_X1    g01936(.A1(new_n2129_), .A2(new_n2125_), .ZN(new_n2130_));
  NOR2_X1    g01937(.A1(new_n2047_), .A2(new_n2115_), .ZN(new_n2131_));
  NOR2_X1    g01938(.A1(new_n2118_), .A2(new_n2131_), .ZN(new_n2132_));
  NAND2_X1   g01939(.A1(new_n2039_), .A2(new_n2041_), .ZN(new_n2133_));
  NAND2_X1   g01940(.A1(new_n2042_), .A2(new_n2037_), .ZN(new_n2134_));
  NAND2_X1   g01941(.A1(new_n2134_), .A2(new_n2133_), .ZN(new_n2135_));
  XOR2_X1    g01942(.A1(new_n2059_), .A2(new_n2071_), .Z(new_n2136_));
  XOR2_X1    g01943(.A1(new_n2136_), .A2(new_n2111_), .Z(new_n2137_));
  NAND2_X1   g01944(.A1(\a[1] ), .A2(\a[31] ), .ZN(new_n2138_));
  XOR2_X1    g01945(.A1(new_n982_), .A2(new_n2138_), .Z(new_n2139_));
  NOR2_X1    g01946(.A1(new_n2099_), .A2(new_n2139_), .ZN(new_n2140_));
  INV_X1     g01947(.I(new_n2139_), .ZN(new_n2141_));
  NOR2_X1    g01948(.A1(new_n2098_), .A2(new_n2141_), .ZN(new_n2142_));
  NOR2_X1    g01949(.A1(new_n2140_), .A2(new_n2142_), .ZN(new_n2143_));
  NOR2_X1    g01950(.A1(new_n2143_), .A2(new_n2092_), .ZN(new_n2144_));
  INV_X1     g01951(.I(new_n2143_), .ZN(new_n2145_));
  NOR2_X1    g01952(.A1(new_n2145_), .A2(new_n2091_), .ZN(new_n2146_));
  NOR2_X1    g01953(.A1(new_n2146_), .A2(new_n2144_), .ZN(new_n2147_));
  XOR2_X1    g01954(.A1(new_n2147_), .A2(new_n2137_), .Z(new_n2148_));
  XOR2_X1    g01955(.A1(new_n2135_), .A2(new_n2148_), .Z(new_n2149_));
  NAND2_X1   g01956(.A1(new_n2093_), .A2(new_n2101_), .ZN(new_n2150_));
  NAND2_X1   g01957(.A1(new_n2102_), .A2(new_n2112_), .ZN(new_n2151_));
  NAND2_X1   g01958(.A1(new_n2151_), .A2(new_n2150_), .ZN(new_n2152_));
  OAI21_X1   g01959(.A1(new_n2064_), .A2(new_n2073_), .B(new_n2077_), .ZN(new_n2153_));
  NAND2_X1   g01960(.A1(new_n1979_), .A2(new_n1924_), .ZN(new_n2154_));
  NAND2_X1   g01961(.A1(new_n2012_), .A2(new_n1995_), .ZN(new_n2155_));
  NAND2_X1   g01962(.A1(new_n2155_), .A2(new_n2154_), .ZN(new_n2156_));
  XOR2_X1    g01963(.A1(new_n2153_), .A2(new_n2156_), .Z(new_n2157_));
  XOR2_X1    g01964(.A1(new_n2157_), .A2(new_n2152_), .Z(new_n2158_));
  NAND2_X1   g01965(.A1(new_n2050_), .A2(new_n2114_), .ZN(new_n2159_));
  OAI21_X1   g01966(.A1(new_n2079_), .A2(new_n2113_), .B(new_n2159_), .ZN(new_n2160_));
  NAND2_X1   g01967(.A1(new_n2160_), .A2(new_n2158_), .ZN(new_n2161_));
  INV_X1     g01968(.I(new_n2161_), .ZN(new_n2162_));
  NOR2_X1    g01969(.A1(new_n2160_), .A2(new_n2158_), .ZN(new_n2163_));
  NOR2_X1    g01970(.A1(new_n2162_), .A2(new_n2163_), .ZN(new_n2164_));
  NAND2_X1   g01971(.A1(new_n2164_), .A2(new_n2149_), .ZN(new_n2165_));
  INV_X1     g01972(.I(new_n2165_), .ZN(new_n2166_));
  NOR2_X1    g01973(.A1(new_n2164_), .A2(new_n2149_), .ZN(new_n2167_));
  NOR2_X1    g01974(.A1(new_n2166_), .A2(new_n2167_), .ZN(new_n2168_));
  NAND2_X1   g01975(.A1(new_n2027_), .A2(new_n2043_), .ZN(new_n2169_));
  NAND2_X1   g01976(.A1(new_n2044_), .A2(new_n2025_), .ZN(new_n2170_));
  NAND2_X1   g01977(.A1(new_n2170_), .A2(new_n2169_), .ZN(new_n2171_));
  NOR2_X1    g01978(.A1(new_n2023_), .A2(new_n2018_), .ZN(new_n2172_));
  NAND2_X1   g01979(.A1(new_n2035_), .A2(new_n2029_), .ZN(new_n2173_));
  NAND2_X1   g01980(.A1(new_n2036_), .A2(new_n1986_), .ZN(new_n2174_));
  NAND2_X1   g01981(.A1(new_n2174_), .A2(new_n2173_), .ZN(new_n2175_));
  NOR2_X1    g01982(.A1(new_n1441_), .A2(new_n1566_), .ZN(new_n2176_));
  INV_X1     g01983(.I(new_n2176_), .ZN(new_n2177_));
  OAI22_X1   g01984(.A1(new_n643_), .A2(new_n2081_), .B1(new_n1779_), .B2(new_n415_), .ZN(new_n2178_));
  OAI21_X1   g01985(.A1(new_n374_), .A2(new_n2177_), .B(new_n2178_), .ZN(new_n2179_));
  NAND3_X1   g01986(.A1(new_n2179_), .A2(\a[8] ), .A3(\a[24] ), .ZN(new_n2180_));
  AOI22_X1   g01987(.A1(\a[6] ), .A2(\a[26] ), .B1(\a[7] ), .B2(\a[25] ), .ZN(new_n2181_));
  NOR2_X1    g01988(.A1(new_n2177_), .A2(new_n374_), .ZN(new_n2182_));
  NOR2_X1    g01989(.A1(new_n2178_), .A2(new_n2182_), .ZN(new_n2183_));
  INV_X1     g01990(.I(new_n2183_), .ZN(new_n2184_));
  OAI21_X1   g01991(.A1(new_n2181_), .A2(new_n2184_), .B(new_n2180_), .ZN(new_n2185_));
  NOR2_X1    g01992(.A1(new_n290_), .A2(new_n1718_), .ZN(new_n2186_));
  AOI21_X1   g01993(.A1(\a[5] ), .A2(\a[27] ), .B(new_n2186_), .ZN(new_n2187_));
  INV_X1     g01994(.I(new_n2187_), .ZN(new_n2188_));
  INV_X1     g01995(.I(new_n2103_), .ZN(new_n2189_));
  NOR2_X1    g01996(.A1(new_n2189_), .A2(new_n242_), .ZN(new_n2190_));
  NOR2_X1    g01997(.A1(new_n403_), .A2(new_n1299_), .ZN(new_n2191_));
  AOI21_X1   g01998(.A1(new_n2188_), .A2(new_n2191_), .B(new_n2190_), .ZN(new_n2192_));
  INV_X1     g01999(.I(new_n2192_), .ZN(new_n2193_));
  OAI21_X1   g02000(.A1(new_n2190_), .A2(new_n2187_), .B(new_n2191_), .ZN(new_n2194_));
  OAI21_X1   g02001(.A1(new_n2193_), .A2(new_n2187_), .B(new_n2194_), .ZN(new_n2195_));
  XOR2_X1    g02002(.A1(new_n2185_), .A2(new_n2195_), .Z(new_n2196_));
  XOR2_X1    g02003(.A1(new_n2196_), .A2(new_n2175_), .Z(new_n2197_));
  AOI22_X1   g02004(.A1(\a[0] ), .A2(\a[32] ), .B1(\a[2] ), .B2(\a[30] ), .ZN(new_n2198_));
  INV_X1     g02005(.I(new_n2198_), .ZN(new_n2199_));
  INV_X1     g02006(.I(\a[32] ), .ZN(new_n2200_));
  NOR2_X1    g02007(.A1(new_n2030_), .A2(new_n2200_), .ZN(new_n2201_));
  INV_X1     g02008(.I(new_n2201_), .ZN(new_n2202_));
  NOR2_X1    g02009(.A1(new_n2202_), .A2(new_n412_), .ZN(new_n2203_));
  AOI21_X1   g02010(.A1(new_n2033_), .A2(new_n2199_), .B(new_n2203_), .ZN(new_n2204_));
  INV_X1     g02011(.I(new_n2204_), .ZN(new_n2205_));
  OAI21_X1   g02012(.A1(new_n2203_), .A2(new_n2198_), .B(new_n2033_), .ZN(new_n2206_));
  OAI21_X1   g02013(.A1(new_n2205_), .A2(new_n2198_), .B(new_n2206_), .ZN(new_n2207_));
  OAI22_X1   g02014(.A1(new_n619_), .A2(new_n1382_), .B1(new_n1379_), .B2(new_n833_), .ZN(new_n2208_));
  OAI21_X1   g02015(.A1(new_n1265_), .A2(new_n1376_), .B(new_n2208_), .ZN(new_n2209_));
  NAND3_X1   g02016(.A1(new_n2209_), .A2(\a[11] ), .A3(\a[21] ), .ZN(new_n2210_));
  AOI22_X1   g02017(.A1(\a[12] ), .A2(\a[20] ), .B1(\a[13] ), .B2(\a[19] ), .ZN(new_n2211_));
  NOR2_X1    g02018(.A1(new_n1265_), .A2(new_n1376_), .ZN(new_n2212_));
  NOR2_X1    g02019(.A1(new_n2208_), .A2(new_n2212_), .ZN(new_n2213_));
  INV_X1     g02020(.I(new_n2213_), .ZN(new_n2214_));
  OAI21_X1   g02021(.A1(new_n2211_), .A2(new_n2214_), .B(new_n2210_), .ZN(new_n2215_));
  XNOR2_X1   g02022(.A1(new_n2215_), .A2(new_n2207_), .ZN(new_n2216_));
  NOR2_X1    g02023(.A1(new_n759_), .A2(new_n884_), .ZN(new_n2217_));
  INV_X1     g02024(.I(new_n2217_), .ZN(new_n2218_));
  AOI22_X1   g02025(.A1(\a[3] ), .A2(\a[29] ), .B1(\a[10] ), .B2(\a[22] ), .ZN(new_n2219_));
  NOR4_X1    g02026(.A1(new_n225_), .A2(new_n417_), .A3(new_n1175_), .A4(new_n1814_), .ZN(new_n2220_));
  NOR3_X1    g02027(.A1(new_n2218_), .A2(new_n2220_), .A3(new_n2219_), .ZN(new_n2221_));
  NOR2_X1    g02028(.A1(new_n2221_), .A2(new_n2220_), .ZN(new_n2222_));
  INV_X1     g02029(.I(new_n2222_), .ZN(new_n2223_));
  OAI22_X1   g02030(.A1(new_n2223_), .A2(new_n2219_), .B1(new_n2218_), .B2(new_n2221_), .ZN(new_n2224_));
  INV_X1     g02031(.I(new_n2224_), .ZN(new_n2225_));
  XOR2_X1    g02032(.A1(new_n2216_), .A2(new_n2225_), .Z(new_n2226_));
  XNOR2_X1   g02033(.A1(new_n2226_), .A2(new_n2197_), .ZN(new_n2227_));
  XOR2_X1    g02034(.A1(new_n2172_), .A2(new_n2227_), .Z(new_n2228_));
  NOR2_X1    g02035(.A1(new_n2171_), .A2(new_n2228_), .ZN(new_n2229_));
  NAND2_X1   g02036(.A1(new_n2171_), .A2(new_n2228_), .ZN(new_n2230_));
  INV_X1     g02037(.I(new_n2230_), .ZN(new_n2231_));
  NOR2_X1    g02038(.A1(new_n2231_), .A2(new_n2229_), .ZN(new_n2232_));
  NOR2_X1    g02039(.A1(new_n2232_), .A2(new_n2168_), .ZN(new_n2233_));
  NAND2_X1   g02040(.A1(new_n2232_), .A2(new_n2168_), .ZN(new_n2234_));
  INV_X1     g02041(.I(new_n2234_), .ZN(new_n2235_));
  NOR2_X1    g02042(.A1(new_n2235_), .A2(new_n2233_), .ZN(new_n2236_));
  INV_X1     g02043(.I(new_n2236_), .ZN(new_n2237_));
  NOR2_X1    g02044(.A1(new_n2237_), .A2(new_n2132_), .ZN(new_n2238_));
  INV_X1     g02045(.I(new_n2238_), .ZN(new_n2239_));
  NAND2_X1   g02046(.A1(new_n2237_), .A2(new_n2132_), .ZN(new_n2240_));
  NAND2_X1   g02047(.A1(new_n2239_), .A2(new_n2240_), .ZN(new_n2241_));
  XOR2_X1    g02048(.A1(new_n2130_), .A2(new_n2241_), .Z(\asquared[33] ));
  OAI21_X1   g02049(.A1(new_n2129_), .A2(new_n2125_), .B(new_n2240_), .ZN(new_n2243_));
  NAND2_X1   g02050(.A1(new_n2243_), .A2(new_n2239_), .ZN(new_n2244_));
  NAND2_X1   g02051(.A1(\a[5] ), .A2(\a[28] ), .ZN(new_n2245_));
  NOR2_X1    g02052(.A1(new_n1441_), .A2(new_n1750_), .ZN(new_n2246_));
  NAND4_X1   g02053(.A1(\a[5] ), .A2(\a[8] ), .A3(\a[25] ), .A4(\a[28] ), .ZN(new_n2247_));
  NAND2_X1   g02054(.A1(new_n2103_), .A2(new_n746_), .ZN(new_n2248_));
  AOI22_X1   g02055(.A1(new_n2248_), .A2(new_n2247_), .B1(new_n645_), .B2(new_n2246_), .ZN(new_n2249_));
  AOI22_X1   g02056(.A1(\a[6] ), .A2(\a[27] ), .B1(\a[8] ), .B2(\a[25] ), .ZN(new_n2250_));
  NAND2_X1   g02057(.A1(new_n2246_), .A2(new_n645_), .ZN(new_n2251_));
  NAND3_X1   g02058(.A1(new_n2251_), .A2(new_n2248_), .A3(new_n2247_), .ZN(new_n2252_));
  OAI22_X1   g02059(.A1(new_n2249_), .A2(new_n2245_), .B1(new_n2252_), .B2(new_n2250_), .ZN(new_n2253_));
  NOR2_X1    g02060(.A1(new_n1814_), .A2(new_n2030_), .ZN(new_n2254_));
  INV_X1     g02061(.I(new_n2254_), .ZN(new_n2255_));
  NOR2_X1    g02062(.A1(new_n2255_), .A2(new_n370_), .ZN(new_n2256_));
  NOR3_X1    g02063(.A1(new_n532_), .A2(new_n1357_), .A3(new_n2030_), .ZN(new_n2257_));
  NAND4_X1   g02064(.A1(\a[4] ), .A2(\a[9] ), .A3(\a[24] ), .A4(\a[29] ), .ZN(new_n2258_));
  OAI21_X1   g02065(.A1(new_n2256_), .A2(new_n2257_), .B(new_n2258_), .ZN(new_n2259_));
  NAND3_X1   g02066(.A1(new_n2259_), .A2(\a[3] ), .A3(\a[30] ), .ZN(new_n2260_));
  AOI22_X1   g02067(.A1(\a[4] ), .A2(\a[29] ), .B1(\a[9] ), .B2(\a[24] ), .ZN(new_n2261_));
  NAND2_X1   g02068(.A1(new_n2259_), .A2(new_n2258_), .ZN(new_n2262_));
  OAI21_X1   g02069(.A1(new_n2261_), .A2(new_n2262_), .B(new_n2260_), .ZN(new_n2263_));
  XNOR2_X1   g02070(.A1(new_n2263_), .A2(new_n2253_), .ZN(new_n2264_));
  AOI21_X1   g02071(.A1(\a[15] ), .A2(\a[18] ), .B(new_n1024_), .ZN(new_n2265_));
  NAND2_X1   g02072(.A1(\a[7] ), .A2(\a[26] ), .ZN(new_n2266_));
  NOR2_X1    g02073(.A1(new_n1275_), .A2(new_n893_), .ZN(new_n2267_));
  NOR3_X1    g02074(.A1(new_n2267_), .A2(new_n2265_), .A3(new_n2266_), .ZN(new_n2268_));
  OAI22_X1   g02075(.A1(new_n2265_), .A2(new_n2266_), .B1(new_n893_), .B2(new_n1275_), .ZN(new_n2269_));
  OAI22_X1   g02076(.A1(new_n2266_), .A2(new_n2268_), .B1(new_n2269_), .B2(new_n2265_), .ZN(new_n2270_));
  XOR2_X1    g02077(.A1(new_n2264_), .A2(new_n2270_), .Z(new_n2271_));
  XOR2_X1    g02078(.A1(new_n2183_), .A2(new_n2192_), .Z(new_n2272_));
  NAND3_X1   g02079(.A1(new_n478_), .A2(\a[22] ), .A3(\a[33] ), .ZN(new_n2273_));
  INV_X1     g02080(.I(\a[33] ), .ZN(new_n2274_));
  NOR2_X1    g02081(.A1(new_n2051_), .A2(new_n2274_), .ZN(new_n2275_));
  INV_X1     g02082(.I(new_n2275_), .ZN(new_n2276_));
  OAI22_X1   g02083(.A1(new_n412_), .A2(new_n2276_), .B1(new_n2053_), .B2(new_n588_), .ZN(new_n2277_));
  NAND2_X1   g02084(.A1(new_n2277_), .A2(new_n2273_), .ZN(new_n2278_));
  NAND3_X1   g02085(.A1(new_n2278_), .A2(\a[2] ), .A3(\a[31] ), .ZN(new_n2279_));
  NAND2_X1   g02086(.A1(new_n2278_), .A2(new_n2273_), .ZN(new_n2280_));
  AOI22_X1   g02087(.A1(\a[0] ), .A2(\a[33] ), .B1(\a[11] ), .B2(\a[22] ), .ZN(new_n2281_));
  OAI21_X1   g02088(.A1(new_n2280_), .A2(new_n2281_), .B(new_n2279_), .ZN(new_n2282_));
  XNOR2_X1   g02089(.A1(new_n2272_), .A2(new_n2282_), .ZN(new_n2283_));
  NAND2_X1   g02090(.A1(new_n2213_), .A2(new_n2204_), .ZN(new_n2284_));
  NAND2_X1   g02091(.A1(new_n2214_), .A2(new_n2205_), .ZN(new_n2285_));
  AND2_X2    g02092(.A1(new_n2285_), .A2(new_n2284_), .Z(new_n2286_));
  XOR2_X1    g02093(.A1(new_n2286_), .A2(new_n2223_), .Z(new_n2287_));
  XNOR2_X1   g02094(.A1(new_n2287_), .A2(new_n2283_), .ZN(new_n2288_));
  XOR2_X1    g02095(.A1(new_n2288_), .A2(new_n2271_), .Z(new_n2289_));
  NAND2_X1   g02096(.A1(new_n2226_), .A2(new_n2197_), .ZN(new_n2290_));
  OAI21_X1   g02097(.A1(new_n2172_), .A2(new_n2227_), .B(new_n2290_), .ZN(new_n2291_));
  NAND2_X1   g02098(.A1(new_n2185_), .A2(new_n2195_), .ZN(new_n2292_));
  NAND2_X1   g02099(.A1(new_n2196_), .A2(new_n2175_), .ZN(new_n2293_));
  NAND2_X1   g02100(.A1(new_n2293_), .A2(new_n2292_), .ZN(new_n2294_));
  NAND2_X1   g02101(.A1(new_n2059_), .A2(new_n2071_), .ZN(new_n2295_));
  NAND2_X1   g02102(.A1(new_n2136_), .A2(new_n2111_), .ZN(new_n2296_));
  NAND2_X1   g02103(.A1(new_n2296_), .A2(new_n2295_), .ZN(new_n2297_));
  NAND2_X1   g02104(.A1(new_n2215_), .A2(new_n2207_), .ZN(new_n2298_));
  OAI21_X1   g02105(.A1(new_n2216_), .A2(new_n2225_), .B(new_n2298_), .ZN(new_n2299_));
  XOR2_X1    g02106(.A1(new_n2299_), .A2(new_n2297_), .Z(new_n2300_));
  XOR2_X1    g02107(.A1(new_n2300_), .A2(new_n2294_), .Z(new_n2301_));
  XOR2_X1    g02108(.A1(new_n2291_), .A2(new_n2301_), .Z(new_n2302_));
  XOR2_X1    g02109(.A1(new_n2302_), .A2(new_n2289_), .Z(new_n2303_));
  NAND2_X1   g02110(.A1(new_n2147_), .A2(new_n2137_), .ZN(new_n2304_));
  NAND2_X1   g02111(.A1(new_n2135_), .A2(new_n2148_), .ZN(new_n2305_));
  NAND2_X1   g02112(.A1(new_n2305_), .A2(new_n2304_), .ZN(new_n2306_));
  NAND2_X1   g02113(.A1(new_n2153_), .A2(new_n2156_), .ZN(new_n2307_));
  NAND2_X1   g02114(.A1(new_n2157_), .A2(new_n2152_), .ZN(new_n2308_));
  NAND2_X1   g02115(.A1(new_n2308_), .A2(new_n2307_), .ZN(new_n2309_));
  NOR2_X1    g02116(.A1(new_n2146_), .A2(new_n2142_), .ZN(new_n2310_));
  NOR2_X1    g02117(.A1(new_n982_), .A2(new_n2138_), .ZN(new_n2311_));
  INV_X1     g02118(.I(new_n2311_), .ZN(new_n2312_));
  NAND2_X1   g02119(.A1(\a[10] ), .A2(\a[23] ), .ZN(new_n2313_));
  NAND2_X1   g02120(.A1(new_n2312_), .A2(new_n2313_), .ZN(new_n2314_));
  INV_X1     g02121(.I(new_n2314_), .ZN(new_n2315_));
  NOR2_X1    g02122(.A1(new_n194_), .A2(new_n2200_), .ZN(new_n2316_));
  XOR2_X1    g02123(.A1(new_n2316_), .A2(new_n1023_), .Z(new_n2317_));
  NOR2_X1    g02124(.A1(new_n2312_), .A2(new_n2313_), .ZN(new_n2318_));
  NOR2_X1    g02125(.A1(new_n2315_), .A2(new_n2318_), .ZN(new_n2319_));
  INV_X1     g02126(.I(new_n2317_), .ZN(new_n2320_));
  AOI21_X1   g02127(.A1(new_n2320_), .A2(new_n2314_), .B(new_n2318_), .ZN(new_n2321_));
  INV_X1     g02128(.I(new_n2321_), .ZN(new_n2322_));
  OAI22_X1   g02129(.A1(new_n2322_), .A2(new_n2315_), .B1(new_n2317_), .B2(new_n2319_), .ZN(new_n2323_));
  NOR2_X1    g02130(.A1(new_n767_), .A2(new_n1376_), .ZN(new_n2324_));
  AOI22_X1   g02131(.A1(new_n763_), .A2(new_n1381_), .B1(new_n1378_), .B2(new_n762_), .ZN(new_n2325_));
  NOR2_X1    g02132(.A1(new_n2324_), .A2(new_n2325_), .ZN(new_n2326_));
  NAND2_X1   g02133(.A1(\a[12] ), .A2(\a[21] ), .ZN(new_n2327_));
  AOI22_X1   g02134(.A1(\a[13] ), .A2(\a[20] ), .B1(\a[14] ), .B2(\a[19] ), .ZN(new_n2328_));
  NOR2_X1    g02135(.A1(new_n2326_), .A2(new_n2324_), .ZN(new_n2329_));
  INV_X1     g02136(.I(new_n2329_), .ZN(new_n2330_));
  OAI22_X1   g02137(.A1(new_n2330_), .A2(new_n2328_), .B1(new_n2326_), .B2(new_n2327_), .ZN(new_n2331_));
  XNOR2_X1   g02138(.A1(new_n2323_), .A2(new_n2331_), .ZN(new_n2332_));
  XOR2_X1    g02139(.A1(new_n2332_), .A2(new_n2310_), .Z(new_n2333_));
  XOR2_X1    g02140(.A1(new_n2309_), .A2(new_n2333_), .Z(new_n2334_));
  XOR2_X1    g02141(.A1(new_n2334_), .A2(new_n2306_), .Z(new_n2335_));
  INV_X1     g02142(.I(new_n2335_), .ZN(new_n2336_));
  NOR2_X1    g02143(.A1(new_n2166_), .A2(new_n2162_), .ZN(new_n2337_));
  XOR2_X1    g02144(.A1(new_n2337_), .A2(new_n2336_), .Z(new_n2338_));
  INV_X1     g02145(.I(new_n2338_), .ZN(new_n2339_));
  NOR2_X1    g02146(.A1(new_n2339_), .A2(new_n2303_), .ZN(new_n2340_));
  INV_X1     g02147(.I(new_n2340_), .ZN(new_n2341_));
  NAND2_X1   g02148(.A1(new_n2339_), .A2(new_n2303_), .ZN(new_n2342_));
  AND2_X2    g02149(.A1(new_n2341_), .A2(new_n2342_), .Z(new_n2343_));
  INV_X1     g02150(.I(new_n2343_), .ZN(new_n2344_));
  NOR2_X1    g02151(.A1(new_n2235_), .A2(new_n2231_), .ZN(new_n2345_));
  NOR2_X1    g02152(.A1(new_n2344_), .A2(new_n2345_), .ZN(new_n2346_));
  NOR3_X1    g02153(.A1(new_n2343_), .A2(new_n2231_), .A3(new_n2235_), .ZN(new_n2347_));
  NOR2_X1    g02154(.A1(new_n2346_), .A2(new_n2347_), .ZN(new_n2348_));
  XOR2_X1    g02155(.A1(new_n2244_), .A2(new_n2348_), .Z(\asquared[34] ));
  AOI21_X1   g02156(.A1(new_n2243_), .A2(new_n2239_), .B(new_n2347_), .ZN(new_n2350_));
  NOR2_X1    g02157(.A1(new_n2350_), .A2(new_n2346_), .ZN(new_n2351_));
  NOR2_X1    g02158(.A1(new_n2337_), .A2(new_n2336_), .ZN(new_n2352_));
  NOR2_X1    g02159(.A1(new_n2340_), .A2(new_n2352_), .ZN(new_n2353_));
  NAND2_X1   g02160(.A1(new_n2309_), .A2(new_n2333_), .ZN(new_n2354_));
  NAND2_X1   g02161(.A1(new_n2334_), .A2(new_n2306_), .ZN(new_n2355_));
  NAND2_X1   g02162(.A1(new_n2355_), .A2(new_n2354_), .ZN(new_n2356_));
  XOR2_X1    g02163(.A1(new_n2280_), .A2(new_n2262_), .Z(new_n2357_));
  XOR2_X1    g02164(.A1(new_n2357_), .A2(new_n2252_), .Z(new_n2358_));
  NAND2_X1   g02165(.A1(new_n2263_), .A2(new_n2253_), .ZN(new_n2359_));
  INV_X1     g02166(.I(new_n2264_), .ZN(new_n2360_));
  NAND2_X1   g02167(.A1(new_n2360_), .A2(new_n2270_), .ZN(new_n2361_));
  NAND2_X1   g02168(.A1(new_n2361_), .A2(new_n2359_), .ZN(new_n2362_));
  NAND2_X1   g02169(.A1(\a[1] ), .A2(\a[33] ), .ZN(new_n2363_));
  NOR2_X1    g02170(.A1(new_n1429_), .A2(new_n2363_), .ZN(new_n2364_));
  INV_X1     g02171(.I(new_n2364_), .ZN(new_n2365_));
  NAND2_X1   g02172(.A1(new_n1429_), .A2(new_n2363_), .ZN(new_n2366_));
  NAND2_X1   g02173(.A1(new_n2365_), .A2(new_n2366_), .ZN(new_n2367_));
  INV_X1     g02174(.I(new_n2316_), .ZN(new_n2368_));
  NOR2_X1    g02175(.A1(new_n2368_), .A2(new_n1023_), .ZN(new_n2369_));
  XNOR2_X1   g02176(.A1(new_n2367_), .A2(new_n2369_), .ZN(new_n2370_));
  XOR2_X1    g02177(.A1(new_n2370_), .A2(new_n2269_), .Z(new_n2371_));
  XOR2_X1    g02178(.A1(new_n2362_), .A2(new_n2371_), .Z(new_n2372_));
  NAND2_X1   g02179(.A1(new_n2372_), .A2(new_n2358_), .ZN(new_n2373_));
  OR2_X2     g02180(.A1(new_n2372_), .A2(new_n2358_), .Z(new_n2374_));
  AND2_X2    g02181(.A1(new_n2374_), .A2(new_n2373_), .Z(new_n2375_));
  INV_X1     g02182(.I(new_n2375_), .ZN(new_n2376_));
  NAND2_X1   g02183(.A1(new_n2323_), .A2(new_n2331_), .ZN(new_n2377_));
  OAI21_X1   g02184(.A1(new_n2310_), .A2(new_n2332_), .B(new_n2377_), .ZN(new_n2378_));
  NOR2_X1    g02185(.A1(new_n2322_), .A2(new_n2330_), .ZN(new_n2379_));
  NOR2_X1    g02186(.A1(new_n2321_), .A2(new_n2329_), .ZN(new_n2380_));
  NOR2_X1    g02187(.A1(new_n2379_), .A2(new_n2380_), .ZN(new_n2381_));
  AOI22_X1   g02188(.A1(\a[11] ), .A2(\a[23] ), .B1(\a[12] ), .B2(\a[22] ), .ZN(new_n2382_));
  NOR2_X1    g02189(.A1(new_n197_), .A2(new_n2200_), .ZN(new_n2383_));
  INV_X1     g02190(.I(new_n2383_), .ZN(new_n2384_));
  INV_X1     g02191(.I(new_n1767_), .ZN(new_n2385_));
  NOR2_X1    g02192(.A1(new_n2385_), .A2(new_n619_), .ZN(new_n2386_));
  NOR3_X1    g02193(.A1(new_n2386_), .A2(new_n2382_), .A3(new_n2384_), .ZN(new_n2387_));
  NOR2_X1    g02194(.A1(new_n2387_), .A2(new_n2386_), .ZN(new_n2388_));
  INV_X1     g02195(.I(new_n2388_), .ZN(new_n2389_));
  OAI22_X1   g02196(.A1(new_n2389_), .A2(new_n2382_), .B1(new_n2384_), .B2(new_n2387_), .ZN(new_n2390_));
  XOR2_X1    g02197(.A1(new_n2381_), .A2(new_n2390_), .Z(new_n2391_));
  XOR2_X1    g02198(.A1(new_n2378_), .A2(new_n2391_), .Z(new_n2392_));
  INV_X1     g02199(.I(new_n2392_), .ZN(new_n2393_));
  NAND4_X1   g02200(.A1(\a[5] ), .A2(\a[9] ), .A3(\a[25] ), .A4(\a[29] ), .ZN(new_n2394_));
  NOR4_X1    g02201(.A1(new_n253_), .A2(new_n417_), .A3(new_n1357_), .A4(new_n1814_), .ZN(new_n2395_));
  NOR2_X1    g02202(.A1(new_n1779_), .A2(new_n539_), .ZN(new_n2396_));
  OAI21_X1   g02203(.A1(new_n2396_), .A2(new_n2395_), .B(new_n2394_), .ZN(new_n2397_));
  NAND3_X1   g02204(.A1(new_n2397_), .A2(\a[10] ), .A3(\a[24] ), .ZN(new_n2398_));
  NAND2_X1   g02205(.A1(new_n2397_), .A2(new_n2394_), .ZN(new_n2399_));
  AOI22_X1   g02206(.A1(\a[5] ), .A2(\a[29] ), .B1(\a[9] ), .B2(\a[25] ), .ZN(new_n2400_));
  OAI21_X1   g02207(.A1(new_n2399_), .A2(new_n2400_), .B(new_n2398_), .ZN(new_n2401_));
  OAI22_X1   g02208(.A1(new_n767_), .A2(new_n1382_), .B1(new_n1379_), .B2(new_n836_), .ZN(new_n2402_));
  OAI21_X1   g02209(.A1(new_n1173_), .A2(new_n1376_), .B(new_n2402_), .ZN(new_n2403_));
  NAND3_X1   g02210(.A1(new_n2403_), .A2(\a[13] ), .A3(\a[21] ), .ZN(new_n2404_));
  AOI22_X1   g02211(.A1(\a[14] ), .A2(\a[20] ), .B1(\a[15] ), .B2(\a[19] ), .ZN(new_n2405_));
  NOR2_X1    g02212(.A1(new_n1173_), .A2(new_n1376_), .ZN(new_n2406_));
  NOR2_X1    g02213(.A1(new_n2402_), .A2(new_n2406_), .ZN(new_n2407_));
  INV_X1     g02214(.I(new_n2407_), .ZN(new_n2408_));
  OAI21_X1   g02215(.A1(new_n2405_), .A2(new_n2408_), .B(new_n2404_), .ZN(new_n2409_));
  XNOR2_X1   g02216(.A1(new_n2409_), .A2(new_n2401_), .ZN(new_n2410_));
  NAND2_X1   g02217(.A1(new_n2103_), .A2(new_n479_), .ZN(new_n2411_));
  NOR2_X1    g02218(.A1(new_n1566_), .A2(new_n1718_), .ZN(new_n2412_));
  NAND2_X1   g02219(.A1(new_n2412_), .A2(new_n645_), .ZN(new_n2413_));
  AOI22_X1   g02220(.A1(new_n2411_), .A2(new_n2413_), .B1(new_n693_), .B2(new_n1971_), .ZN(new_n2414_));
  NAND2_X1   g02221(.A1(\a[6] ), .A2(\a[28] ), .ZN(new_n2415_));
  AOI22_X1   g02222(.A1(\a[7] ), .A2(\a[27] ), .B1(\a[8] ), .B2(\a[26] ), .ZN(new_n2416_));
  NAND2_X1   g02223(.A1(new_n1971_), .A2(new_n693_), .ZN(new_n2417_));
  NAND3_X1   g02224(.A1(new_n2417_), .A2(new_n2411_), .A3(new_n2413_), .ZN(new_n2418_));
  OAI22_X1   g02225(.A1(new_n2414_), .A2(new_n2415_), .B1(new_n2418_), .B2(new_n2416_), .ZN(new_n2419_));
  XOR2_X1    g02226(.A1(new_n2410_), .A2(new_n2419_), .Z(new_n2420_));
  NOR2_X1    g02227(.A1(new_n2393_), .A2(new_n2420_), .ZN(new_n2421_));
  NAND2_X1   g02228(.A1(new_n2393_), .A2(new_n2420_), .ZN(new_n2422_));
  INV_X1     g02229(.I(new_n2422_), .ZN(new_n2423_));
  NOR3_X1    g02230(.A1(new_n2376_), .A2(new_n2421_), .A3(new_n2423_), .ZN(new_n2424_));
  NOR2_X1    g02231(.A1(new_n2424_), .A2(new_n2376_), .ZN(new_n2425_));
  NOR3_X1    g02232(.A1(new_n2375_), .A2(new_n2421_), .A3(new_n2423_), .ZN(new_n2426_));
  NOR2_X1    g02233(.A1(new_n2425_), .A2(new_n2426_), .ZN(new_n2427_));
  XOR2_X1    g02234(.A1(new_n2427_), .A2(new_n2356_), .Z(new_n2428_));
  NOR2_X1    g02235(.A1(new_n2291_), .A2(new_n2301_), .ZN(new_n2429_));
  NAND2_X1   g02236(.A1(new_n2291_), .A2(new_n2301_), .ZN(new_n2430_));
  OAI21_X1   g02237(.A1(new_n2289_), .A2(new_n2429_), .B(new_n2430_), .ZN(new_n2431_));
  NAND2_X1   g02238(.A1(new_n2272_), .A2(new_n2282_), .ZN(new_n2432_));
  OAI21_X1   g02239(.A1(new_n2183_), .A2(new_n2192_), .B(new_n2432_), .ZN(new_n2433_));
  NAND2_X1   g02240(.A1(new_n2286_), .A2(new_n2223_), .ZN(new_n2434_));
  NAND2_X1   g02241(.A1(new_n2434_), .A2(new_n2285_), .ZN(new_n2435_));
  OAI22_X1   g02242(.A1(new_n2030_), .A2(new_n595_), .B1(new_n202_), .B2(new_n2051_), .ZN(new_n2436_));
  NOR2_X1    g02243(.A1(new_n2030_), .A2(new_n2051_), .ZN(new_n2437_));
  INV_X1     g02244(.I(new_n2437_), .ZN(new_n2438_));
  NOR2_X1    g02245(.A1(new_n2438_), .A2(new_n370_), .ZN(new_n2439_));
  INV_X1     g02246(.I(new_n2439_), .ZN(new_n2440_));
  NAND3_X1   g02247(.A1(new_n2440_), .A2(new_n2436_), .A3(\a[34] ), .ZN(new_n2441_));
  INV_X1     g02248(.I(\a[34] ), .ZN(new_n2442_));
  AOI22_X1   g02249(.A1(\a[3] ), .A2(\a[31] ), .B1(\a[4] ), .B2(\a[30] ), .ZN(new_n2443_));
  OAI22_X1   g02250(.A1(new_n2439_), .A2(new_n2443_), .B1(new_n196_), .B2(new_n2442_), .ZN(new_n2444_));
  NAND2_X1   g02251(.A1(new_n2441_), .A2(new_n2444_), .ZN(new_n2445_));
  XNOR2_X1   g02252(.A1(new_n2435_), .A2(new_n2445_), .ZN(new_n2446_));
  XOR2_X1    g02253(.A1(new_n2446_), .A2(new_n2433_), .Z(new_n2447_));
  INV_X1     g02254(.I(new_n2271_), .ZN(new_n2448_));
  INV_X1     g02255(.I(new_n2287_), .ZN(new_n2449_));
  NOR2_X1    g02256(.A1(new_n2449_), .A2(new_n2283_), .ZN(new_n2450_));
  AOI21_X1   g02257(.A1(new_n2288_), .A2(new_n2448_), .B(new_n2450_), .ZN(new_n2451_));
  INV_X1     g02258(.I(new_n2451_), .ZN(new_n2452_));
  NAND2_X1   g02259(.A1(new_n2299_), .A2(new_n2297_), .ZN(new_n2453_));
  NAND2_X1   g02260(.A1(new_n2300_), .A2(new_n2294_), .ZN(new_n2454_));
  NAND2_X1   g02261(.A1(new_n2454_), .A2(new_n2453_), .ZN(new_n2455_));
  XOR2_X1    g02262(.A1(new_n2455_), .A2(new_n2452_), .Z(new_n2456_));
  XOR2_X1    g02263(.A1(new_n2456_), .A2(new_n2447_), .Z(new_n2457_));
  NOR2_X1    g02264(.A1(new_n2457_), .A2(new_n2431_), .ZN(new_n2458_));
  NAND2_X1   g02265(.A1(new_n2457_), .A2(new_n2431_), .ZN(new_n2459_));
  INV_X1     g02266(.I(new_n2459_), .ZN(new_n2460_));
  NOR2_X1    g02267(.A1(new_n2460_), .A2(new_n2458_), .ZN(new_n2461_));
  INV_X1     g02268(.I(new_n2461_), .ZN(new_n2462_));
  XOR2_X1    g02269(.A1(new_n2428_), .A2(new_n2462_), .Z(new_n2463_));
  INV_X1     g02270(.I(new_n2463_), .ZN(new_n2464_));
  NOR2_X1    g02271(.A1(new_n2353_), .A2(new_n2464_), .ZN(new_n2465_));
  INV_X1     g02272(.I(new_n2465_), .ZN(new_n2466_));
  NAND2_X1   g02273(.A1(new_n2353_), .A2(new_n2464_), .ZN(new_n2467_));
  NAND2_X1   g02274(.A1(new_n2466_), .A2(new_n2467_), .ZN(new_n2468_));
  INV_X1     g02275(.I(new_n2346_), .ZN(new_n2469_));
  INV_X1     g02276(.I(new_n2006_), .ZN(new_n2470_));
  INV_X1     g02277(.I(new_n1907_), .ZN(new_n2471_));
  INV_X1     g02278(.I(new_n1516_), .ZN(new_n2472_));
  OAI21_X1   g02279(.A1(new_n1417_), .A2(new_n1410_), .B(new_n1514_), .ZN(new_n2473_));
  INV_X1     g02280(.I(new_n1607_), .ZN(new_n2474_));
  AOI21_X1   g02281(.A1(new_n2473_), .A2(new_n2472_), .B(new_n2474_), .ZN(new_n2475_));
  INV_X1     g02282(.I(new_n1694_), .ZN(new_n2476_));
  OAI21_X1   g02283(.A1(new_n2475_), .A2(new_n1608_), .B(new_n2476_), .ZN(new_n2477_));
  INV_X1     g02284(.I(new_n1796_), .ZN(new_n2478_));
  AOI21_X1   g02285(.A1(new_n2477_), .A2(new_n1695_), .B(new_n2478_), .ZN(new_n2479_));
  INV_X1     g02286(.I(new_n1908_), .ZN(new_n2480_));
  OAI21_X1   g02287(.A1(new_n2479_), .A2(new_n1794_), .B(new_n2480_), .ZN(new_n2481_));
  AOI21_X1   g02288(.A1(new_n2481_), .A2(new_n2471_), .B(new_n2004_), .ZN(new_n2482_));
  INV_X1     g02289(.I(new_n2126_), .ZN(new_n2483_));
  OAI21_X1   g02290(.A1(new_n2482_), .A2(new_n2470_), .B(new_n2483_), .ZN(new_n2484_));
  INV_X1     g02291(.I(new_n2240_), .ZN(new_n2485_));
  AOI21_X1   g02292(.A1(new_n2484_), .A2(new_n2124_), .B(new_n2485_), .ZN(new_n2486_));
  INV_X1     g02293(.I(new_n2347_), .ZN(new_n2487_));
  OAI21_X1   g02294(.A1(new_n2486_), .A2(new_n2238_), .B(new_n2487_), .ZN(new_n2488_));
  INV_X1     g02295(.I(new_n2467_), .ZN(new_n2489_));
  AOI21_X1   g02296(.A1(new_n2488_), .A2(new_n2469_), .B(new_n2489_), .ZN(new_n2490_));
  AOI22_X1   g02297(.A1(new_n2490_), .A2(new_n2466_), .B1(new_n2351_), .B2(new_n2468_), .ZN(\asquared[35] ));
  OAI21_X1   g02298(.A1(new_n2350_), .A2(new_n2346_), .B(new_n2467_), .ZN(new_n2492_));
  NAND2_X1   g02299(.A1(new_n2492_), .A2(new_n2466_), .ZN(new_n2493_));
  NOR2_X1    g02300(.A1(new_n2428_), .A2(new_n2462_), .ZN(new_n2494_));
  NOR2_X1    g02301(.A1(new_n2494_), .A2(new_n2460_), .ZN(new_n2495_));
  NAND2_X1   g02302(.A1(new_n2455_), .A2(new_n2452_), .ZN(new_n2496_));
  NAND2_X1   g02303(.A1(new_n2456_), .A2(new_n2447_), .ZN(new_n2497_));
  NAND2_X1   g02304(.A1(new_n2497_), .A2(new_n2496_), .ZN(new_n2498_));
  NAND2_X1   g02305(.A1(new_n2441_), .A2(new_n2440_), .ZN(new_n2499_));
  XOR2_X1    g02306(.A1(new_n2388_), .A2(new_n2407_), .Z(new_n2500_));
  XOR2_X1    g02307(.A1(new_n2500_), .A2(new_n2499_), .Z(new_n2501_));
  NAND2_X1   g02308(.A1(new_n2409_), .A2(new_n2401_), .ZN(new_n2502_));
  INV_X1     g02309(.I(new_n2410_), .ZN(new_n2503_));
  NAND2_X1   g02310(.A1(new_n2503_), .A2(new_n2419_), .ZN(new_n2504_));
  NAND2_X1   g02311(.A1(new_n2504_), .A2(new_n2502_), .ZN(new_n2505_));
  NOR2_X1    g02312(.A1(new_n194_), .A2(new_n2442_), .ZN(new_n2506_));
  NOR2_X1    g02313(.A1(new_n955_), .A2(new_n2442_), .ZN(new_n2507_));
  INV_X1     g02314(.I(new_n2507_), .ZN(new_n2508_));
  OAI21_X1   g02315(.A1(\a[18] ), .A2(new_n2506_), .B(new_n2508_), .ZN(new_n2509_));
  XNOR2_X1   g02316(.A1(new_n2418_), .A2(new_n2509_), .ZN(new_n2510_));
  XOR2_X1    g02317(.A1(new_n2510_), .A2(new_n2399_), .Z(new_n2511_));
  XOR2_X1    g02318(.A1(new_n2505_), .A2(new_n2511_), .Z(new_n2512_));
  XOR2_X1    g02319(.A1(new_n2512_), .A2(new_n2501_), .Z(new_n2513_));
  XOR2_X1    g02320(.A1(new_n2498_), .A2(new_n2513_), .Z(new_n2514_));
  AOI22_X1   g02321(.A1(\a[11] ), .A2(\a[24] ), .B1(\a[12] ), .B2(\a[23] ), .ZN(new_n2515_));
  NOR2_X1    g02322(.A1(new_n225_), .A2(new_n2200_), .ZN(new_n2516_));
  NOR2_X1    g02323(.A1(new_n1529_), .A2(new_n619_), .ZN(new_n2517_));
  OAI21_X1   g02324(.A1(new_n2517_), .A2(new_n2515_), .B(new_n2516_), .ZN(new_n2518_));
  INV_X1     g02325(.I(new_n2515_), .ZN(new_n2519_));
  AOI21_X1   g02326(.A1(new_n2516_), .A2(new_n2519_), .B(new_n2517_), .ZN(new_n2520_));
  INV_X1     g02327(.I(new_n2520_), .ZN(new_n2521_));
  OAI21_X1   g02328(.A1(new_n2521_), .A2(new_n2515_), .B(new_n2518_), .ZN(new_n2522_));
  AOI22_X1   g02329(.A1(\a[0] ), .A2(\a[35] ), .B1(\a[2] ), .B2(\a[33] ), .ZN(new_n2523_));
  INV_X1     g02330(.I(\a[35] ), .ZN(new_n2524_));
  NOR2_X1    g02331(.A1(new_n2274_), .A2(new_n2524_), .ZN(new_n2525_));
  INV_X1     g02332(.I(new_n2525_), .ZN(new_n2526_));
  NOR2_X1    g02333(.A1(new_n2526_), .A2(new_n412_), .ZN(new_n2527_));
  NOR2_X1    g02334(.A1(new_n2365_), .A2(new_n2523_), .ZN(new_n2528_));
  NOR2_X1    g02335(.A1(new_n2528_), .A2(new_n2527_), .ZN(new_n2529_));
  INV_X1     g02336(.I(new_n2529_), .ZN(new_n2530_));
  OAI21_X1   g02337(.A1(new_n2523_), .A2(new_n2527_), .B(new_n2364_), .ZN(new_n2531_));
  OAI21_X1   g02338(.A1(new_n2530_), .A2(new_n2523_), .B(new_n2531_), .ZN(new_n2532_));
  XOR2_X1    g02339(.A1(new_n2532_), .A2(new_n2522_), .Z(new_n2533_));
  NAND2_X1   g02340(.A1(new_n760_), .A2(new_n1452_), .ZN(new_n2534_));
  NAND2_X1   g02341(.A1(new_n1552_), .A2(new_n1101_), .ZN(new_n2535_));
  AOI22_X1   g02342(.A1(new_n2534_), .A2(new_n2535_), .B1(new_n897_), .B2(new_n1381_), .ZN(new_n2536_));
  NAND2_X1   g02343(.A1(\a[13] ), .A2(\a[22] ), .ZN(new_n2537_));
  AOI22_X1   g02344(.A1(\a[14] ), .A2(\a[21] ), .B1(\a[15] ), .B2(\a[20] ), .ZN(new_n2538_));
  NAND2_X1   g02345(.A1(new_n897_), .A2(new_n1381_), .ZN(new_n2539_));
  NAND3_X1   g02346(.A1(new_n2539_), .A2(new_n2534_), .A3(new_n2535_), .ZN(new_n2540_));
  OAI22_X1   g02347(.A1(new_n2536_), .A2(new_n2537_), .B1(new_n2540_), .B2(new_n2538_), .ZN(new_n2541_));
  XNOR2_X1   g02348(.A1(new_n2533_), .A2(new_n2541_), .ZN(new_n2542_));
  INV_X1     g02349(.I(new_n2542_), .ZN(new_n2543_));
  NAND3_X1   g02350(.A1(new_n2435_), .A2(new_n2441_), .A3(new_n2444_), .ZN(new_n2544_));
  NAND2_X1   g02351(.A1(new_n2446_), .A2(new_n2433_), .ZN(new_n2545_));
  NAND2_X1   g02352(.A1(new_n2545_), .A2(new_n2544_), .ZN(new_n2546_));
  AOI21_X1   g02353(.A1(\a[16] ), .A2(\a[19] ), .B(new_n1027_), .ZN(new_n2547_));
  NOR2_X1    g02354(.A1(new_n422_), .A2(new_n1718_), .ZN(new_n2548_));
  NOR3_X1    g02355(.A1(new_n1275_), .A2(new_n742_), .A3(new_n979_), .ZN(new_n2549_));
  OAI21_X1   g02356(.A1(new_n2549_), .A2(new_n2547_), .B(new_n2548_), .ZN(new_n2550_));
  INV_X1     g02357(.I(new_n2547_), .ZN(new_n2551_));
  AOI21_X1   g02358(.A1(new_n2551_), .A2(new_n2548_), .B(new_n2549_), .ZN(new_n2552_));
  INV_X1     g02359(.I(new_n2552_), .ZN(new_n2553_));
  OAI21_X1   g02360(.A1(new_n2553_), .A2(new_n2547_), .B(new_n2550_), .ZN(new_n2554_));
  NAND2_X1   g02361(.A1(\a[27] ), .A2(\a[30] ), .ZN(new_n2555_));
  OAI22_X1   g02362(.A1(new_n2255_), .A2(new_n371_), .B1(new_n352_), .B2(new_n2555_), .ZN(new_n2556_));
  OAI21_X1   g02363(.A1(new_n643_), .A2(new_n1816_), .B(new_n2556_), .ZN(new_n2557_));
  NAND3_X1   g02364(.A1(new_n2557_), .A2(\a[5] ), .A3(\a[30] ), .ZN(new_n2558_));
  AOI22_X1   g02365(.A1(\a[6] ), .A2(\a[29] ), .B1(\a[8] ), .B2(\a[27] ), .ZN(new_n2559_));
  NOR2_X1    g02366(.A1(new_n1816_), .A2(new_n643_), .ZN(new_n2560_));
  NOR2_X1    g02367(.A1(new_n2556_), .A2(new_n2560_), .ZN(new_n2561_));
  INV_X1     g02368(.I(new_n2561_), .ZN(new_n2562_));
  OAI21_X1   g02369(.A1(new_n2559_), .A2(new_n2562_), .B(new_n2558_), .ZN(new_n2563_));
  XNOR2_X1   g02370(.A1(new_n2563_), .A2(new_n2554_), .ZN(new_n2564_));
  AOI22_X1   g02371(.A1(\a[9] ), .A2(\a[26] ), .B1(\a[10] ), .B2(\a[25] ), .ZN(new_n2565_));
  NOR2_X1    g02372(.A1(new_n290_), .A2(new_n2051_), .ZN(new_n2566_));
  INV_X1     g02373(.I(new_n2566_), .ZN(new_n2567_));
  NOR2_X1    g02374(.A1(new_n2177_), .A2(new_n539_), .ZN(new_n2568_));
  NOR3_X1    g02375(.A1(new_n2568_), .A2(new_n2565_), .A3(new_n2567_), .ZN(new_n2569_));
  NOR2_X1    g02376(.A1(new_n2569_), .A2(new_n2568_), .ZN(new_n2570_));
  INV_X1     g02377(.I(new_n2570_), .ZN(new_n2571_));
  OAI22_X1   g02378(.A1(new_n2571_), .A2(new_n2565_), .B1(new_n2567_), .B2(new_n2569_), .ZN(new_n2572_));
  INV_X1     g02379(.I(new_n2572_), .ZN(new_n2573_));
  XOR2_X1    g02380(.A1(new_n2564_), .A2(new_n2573_), .Z(new_n2574_));
  NOR2_X1    g02381(.A1(new_n2546_), .A2(new_n2574_), .ZN(new_n2575_));
  NAND2_X1   g02382(.A1(new_n2546_), .A2(new_n2574_), .ZN(new_n2576_));
  INV_X1     g02383(.I(new_n2576_), .ZN(new_n2577_));
  NOR2_X1    g02384(.A1(new_n2577_), .A2(new_n2575_), .ZN(new_n2578_));
  NAND2_X1   g02385(.A1(new_n2578_), .A2(new_n2543_), .ZN(new_n2579_));
  INV_X1     g02386(.I(new_n2579_), .ZN(new_n2580_));
  NOR2_X1    g02387(.A1(new_n2578_), .A2(new_n2543_), .ZN(new_n2581_));
  NOR2_X1    g02388(.A1(new_n2580_), .A2(new_n2581_), .ZN(new_n2582_));
  XNOR2_X1   g02389(.A1(new_n2514_), .A2(new_n2582_), .ZN(new_n2583_));
  INV_X1     g02390(.I(new_n2583_), .ZN(new_n2584_));
  INV_X1     g02391(.I(new_n2424_), .ZN(new_n2585_));
  OAI21_X1   g02392(.A1(new_n2425_), .A2(new_n2426_), .B(new_n2356_), .ZN(new_n2586_));
  NAND2_X1   g02393(.A1(new_n2586_), .A2(new_n2585_), .ZN(new_n2587_));
  NAND2_X1   g02394(.A1(new_n2378_), .A2(new_n2391_), .ZN(new_n2588_));
  OAI21_X1   g02395(.A1(new_n2393_), .A2(new_n2420_), .B(new_n2588_), .ZN(new_n2589_));
  NAND2_X1   g02396(.A1(new_n2321_), .A2(new_n2329_), .ZN(new_n2590_));
  AOI21_X1   g02397(.A1(new_n2390_), .A2(new_n2590_), .B(new_n2380_), .ZN(new_n2591_));
  INV_X1     g02398(.I(new_n2591_), .ZN(new_n2592_));
  NAND2_X1   g02399(.A1(new_n2280_), .A2(new_n2262_), .ZN(new_n2593_));
  NAND2_X1   g02400(.A1(new_n2357_), .A2(new_n2252_), .ZN(new_n2594_));
  NAND2_X1   g02401(.A1(new_n2594_), .A2(new_n2593_), .ZN(new_n2595_));
  NAND3_X1   g02402(.A1(new_n2365_), .A2(new_n2366_), .A3(new_n2369_), .ZN(new_n2596_));
  NAND2_X1   g02403(.A1(new_n2370_), .A2(new_n2269_), .ZN(new_n2597_));
  NAND2_X1   g02404(.A1(new_n2597_), .A2(new_n2596_), .ZN(new_n2598_));
  XOR2_X1    g02405(.A1(new_n2595_), .A2(new_n2598_), .Z(new_n2599_));
  XOR2_X1    g02406(.A1(new_n2599_), .A2(new_n2592_), .Z(new_n2600_));
  NAND2_X1   g02407(.A1(new_n2362_), .A2(new_n2371_), .ZN(new_n2601_));
  NAND2_X1   g02408(.A1(new_n2373_), .A2(new_n2601_), .ZN(new_n2602_));
  XOR2_X1    g02409(.A1(new_n2602_), .A2(new_n2600_), .Z(new_n2603_));
  XOR2_X1    g02410(.A1(new_n2603_), .A2(new_n2589_), .Z(new_n2604_));
  NOR2_X1    g02411(.A1(new_n2587_), .A2(new_n2604_), .ZN(new_n2605_));
  NAND2_X1   g02412(.A1(new_n2587_), .A2(new_n2604_), .ZN(new_n2606_));
  INV_X1     g02413(.I(new_n2606_), .ZN(new_n2607_));
  NOR2_X1    g02414(.A1(new_n2607_), .A2(new_n2605_), .ZN(new_n2608_));
  NAND2_X1   g02415(.A1(new_n2584_), .A2(new_n2608_), .ZN(new_n2609_));
  INV_X1     g02416(.I(new_n2609_), .ZN(new_n2610_));
  NOR2_X1    g02417(.A1(new_n2584_), .A2(new_n2608_), .ZN(new_n2611_));
  NOR2_X1    g02418(.A1(new_n2610_), .A2(new_n2611_), .ZN(new_n2612_));
  INV_X1     g02419(.I(new_n2612_), .ZN(new_n2613_));
  NOR2_X1    g02420(.A1(new_n2613_), .A2(new_n2495_), .ZN(new_n2614_));
  NAND2_X1   g02421(.A1(new_n2613_), .A2(new_n2495_), .ZN(new_n2615_));
  INV_X1     g02422(.I(new_n2615_), .ZN(new_n2616_));
  NOR2_X1    g02423(.A1(new_n2616_), .A2(new_n2614_), .ZN(new_n2617_));
  XOR2_X1    g02424(.A1(new_n2493_), .A2(new_n2617_), .Z(\asquared[36] ));
  AOI21_X1   g02425(.A1(new_n2492_), .A2(new_n2466_), .B(new_n2616_), .ZN(new_n2619_));
  NOR2_X1    g02426(.A1(new_n2619_), .A2(new_n2614_), .ZN(new_n2620_));
  NOR2_X1    g02427(.A1(new_n2610_), .A2(new_n2607_), .ZN(new_n2621_));
  INV_X1     g02428(.I(new_n2621_), .ZN(new_n2622_));
  NAND2_X1   g02429(.A1(new_n2595_), .A2(new_n2598_), .ZN(new_n2623_));
  NAND2_X1   g02430(.A1(new_n2599_), .A2(new_n2592_), .ZN(new_n2624_));
  NAND2_X1   g02431(.A1(new_n2624_), .A2(new_n2623_), .ZN(new_n2625_));
  INV_X1     g02432(.I(\a[36] ), .ZN(new_n2626_));
  NOR2_X1    g02433(.A1(new_n196_), .A2(new_n2626_), .ZN(new_n2627_));
  XOR2_X1    g02434(.A1(new_n2507_), .A2(new_n2627_), .Z(new_n2628_));
  NOR2_X1    g02435(.A1(new_n1023_), .A2(new_n979_), .ZN(new_n2629_));
  NAND2_X1   g02436(.A1(\a[1] ), .A2(\a[35] ), .ZN(new_n2630_));
  XNOR2_X1   g02437(.A1(new_n2629_), .A2(new_n2630_), .ZN(new_n2631_));
  XOR2_X1    g02438(.A1(new_n2628_), .A2(new_n2631_), .Z(new_n2632_));
  AOI22_X1   g02439(.A1(\a[4] ), .A2(\a[32] ), .B1(\a[11] ), .B2(\a[25] ), .ZN(new_n2633_));
  NOR4_X1    g02440(.A1(new_n290_), .A2(new_n513_), .A3(new_n1441_), .A4(new_n2200_), .ZN(new_n2634_));
  INV_X1     g02441(.I(new_n2634_), .ZN(new_n2635_));
  NOR2_X1    g02442(.A1(new_n2200_), .A2(new_n2274_), .ZN(new_n2636_));
  INV_X1     g02443(.I(new_n2636_), .ZN(new_n2637_));
  NOR2_X1    g02444(.A1(new_n225_), .A2(new_n2274_), .ZN(new_n2638_));
  NAND3_X1   g02445(.A1(new_n2638_), .A2(\a[11] ), .A3(\a[25] ), .ZN(new_n2639_));
  OAI21_X1   g02446(.A1(new_n370_), .A2(new_n2637_), .B(new_n2639_), .ZN(new_n2640_));
  NAND2_X1   g02447(.A1(new_n2640_), .A2(new_n2635_), .ZN(new_n2641_));
  NAND2_X1   g02448(.A1(new_n2641_), .A2(new_n2635_), .ZN(new_n2642_));
  NAND2_X1   g02449(.A1(new_n2641_), .A2(new_n2638_), .ZN(new_n2643_));
  OAI21_X1   g02450(.A1(new_n2633_), .A2(new_n2642_), .B(new_n2643_), .ZN(new_n2644_));
  NOR2_X1    g02451(.A1(new_n1382_), .A2(new_n893_), .ZN(new_n2645_));
  NOR2_X1    g02452(.A1(new_n1173_), .A2(new_n1456_), .ZN(new_n2646_));
  INV_X1     g02453(.I(new_n1552_), .ZN(new_n2647_));
  NOR2_X1    g02454(.A1(new_n2028_), .A2(new_n2647_), .ZN(new_n2648_));
  NOR2_X1    g02455(.A1(new_n2646_), .A2(new_n2648_), .ZN(new_n2649_));
  NOR2_X1    g02456(.A1(new_n2649_), .A2(new_n2645_), .ZN(new_n2650_));
  NAND2_X1   g02457(.A1(\a[14] ), .A2(\a[22] ), .ZN(new_n2651_));
  AOI22_X1   g02458(.A1(\a[15] ), .A2(\a[21] ), .B1(\a[16] ), .B2(\a[20] ), .ZN(new_n2652_));
  NOR2_X1    g02459(.A1(new_n2650_), .A2(new_n2645_), .ZN(new_n2653_));
  INV_X1     g02460(.I(new_n2653_), .ZN(new_n2654_));
  OAI22_X1   g02461(.A1(new_n2654_), .A2(new_n2652_), .B1(new_n2650_), .B2(new_n2651_), .ZN(new_n2655_));
  XOR2_X1    g02462(.A1(new_n2655_), .A2(new_n2644_), .Z(new_n2656_));
  XOR2_X1    g02463(.A1(new_n2656_), .A2(new_n2632_), .Z(new_n2657_));
  XOR2_X1    g02464(.A1(new_n2625_), .A2(new_n2657_), .Z(new_n2658_));
  NOR4_X1    g02465(.A1(new_n253_), .A2(new_n403_), .A3(new_n1750_), .A4(new_n2051_), .ZN(new_n2659_));
  INV_X1     g02466(.I(new_n2055_), .ZN(new_n2660_));
  NOR3_X1    g02467(.A1(new_n2660_), .A2(new_n253_), .A3(new_n1566_), .ZN(new_n2661_));
  NOR2_X1    g02468(.A1(new_n1972_), .A2(new_n539_), .ZN(new_n2662_));
  NOR2_X1    g02469(.A1(new_n2661_), .A2(new_n2662_), .ZN(new_n2663_));
  NOR2_X1    g02470(.A1(new_n2663_), .A2(new_n2659_), .ZN(new_n2664_));
  NAND2_X1   g02471(.A1(\a[10] ), .A2(\a[26] ), .ZN(new_n2665_));
  NOR2_X1    g02472(.A1(new_n2664_), .A2(new_n2659_), .ZN(new_n2666_));
  INV_X1     g02473(.I(new_n2666_), .ZN(new_n2667_));
  AOI22_X1   g02474(.A1(\a[5] ), .A2(\a[31] ), .B1(\a[9] ), .B2(\a[27] ), .ZN(new_n2668_));
  OAI22_X1   g02475(.A1(new_n2667_), .A2(new_n2668_), .B1(new_n2664_), .B2(new_n2665_), .ZN(new_n2669_));
  AOI22_X1   g02476(.A1(\a[12] ), .A2(\a[24] ), .B1(\a[13] ), .B2(\a[23] ), .ZN(new_n2670_));
  INV_X1     g02477(.I(new_n2670_), .ZN(new_n2671_));
  NOR2_X1    g02478(.A1(new_n1265_), .A2(new_n1529_), .ZN(new_n2672_));
  NOR2_X1    g02479(.A1(new_n197_), .A2(new_n2442_), .ZN(new_n2673_));
  AOI21_X1   g02480(.A1(new_n2671_), .A2(new_n2673_), .B(new_n2672_), .ZN(new_n2674_));
  INV_X1     g02481(.I(new_n2674_), .ZN(new_n2675_));
  OAI21_X1   g02482(.A1(new_n2672_), .A2(new_n2670_), .B(new_n2673_), .ZN(new_n2676_));
  OAI21_X1   g02483(.A1(new_n2675_), .A2(new_n2670_), .B(new_n2676_), .ZN(new_n2677_));
  XOR2_X1    g02484(.A1(new_n2669_), .A2(new_n2677_), .Z(new_n2678_));
  INV_X1     g02485(.I(new_n2105_), .ZN(new_n2679_));
  NOR2_X1    g02486(.A1(new_n2679_), .A2(new_n415_), .ZN(new_n2680_));
  NOR2_X1    g02487(.A1(new_n1718_), .A2(new_n2030_), .ZN(new_n2681_));
  AOI22_X1   g02488(.A1(new_n645_), .A2(new_n2681_), .B1(new_n2254_), .B2(new_n479_), .ZN(new_n2682_));
  NOR2_X1    g02489(.A1(new_n2680_), .A2(new_n2682_), .ZN(new_n2683_));
  NAND2_X1   g02490(.A1(\a[6] ), .A2(\a[30] ), .ZN(new_n2684_));
  AOI22_X1   g02491(.A1(\a[7] ), .A2(\a[29] ), .B1(\a[8] ), .B2(\a[28] ), .ZN(new_n2685_));
  NOR2_X1    g02492(.A1(new_n2683_), .A2(new_n2680_), .ZN(new_n2686_));
  INV_X1     g02493(.I(new_n2686_), .ZN(new_n2687_));
  OAI22_X1   g02494(.A1(new_n2687_), .A2(new_n2685_), .B1(new_n2683_), .B2(new_n2684_), .ZN(new_n2688_));
  XOR2_X1    g02495(.A1(new_n2678_), .A2(new_n2688_), .Z(new_n2689_));
  XNOR2_X1   g02496(.A1(new_n2658_), .A2(new_n2689_), .ZN(new_n2690_));
  NAND2_X1   g02497(.A1(new_n2602_), .A2(new_n2600_), .ZN(new_n2691_));
  NAND2_X1   g02498(.A1(new_n2603_), .A2(new_n2589_), .ZN(new_n2692_));
  NAND2_X1   g02499(.A1(new_n2692_), .A2(new_n2691_), .ZN(new_n2693_));
  XOR2_X1    g02500(.A1(new_n2570_), .A2(new_n2561_), .Z(new_n2694_));
  XOR2_X1    g02501(.A1(new_n2694_), .A2(new_n2553_), .Z(new_n2695_));
  NAND2_X1   g02502(.A1(new_n2563_), .A2(new_n2554_), .ZN(new_n2696_));
  OAI21_X1   g02503(.A1(new_n2564_), .A2(new_n2573_), .B(new_n2696_), .ZN(new_n2697_));
  XNOR2_X1   g02504(.A1(new_n2520_), .A2(new_n2540_), .ZN(new_n2698_));
  XOR2_X1    g02505(.A1(new_n2698_), .A2(new_n2530_), .Z(new_n2699_));
  XOR2_X1    g02506(.A1(new_n2697_), .A2(new_n2699_), .Z(new_n2700_));
  XOR2_X1    g02507(.A1(new_n2700_), .A2(new_n2695_), .Z(new_n2701_));
  INV_X1     g02508(.I(new_n2701_), .ZN(new_n2702_));
  NAND2_X1   g02509(.A1(new_n2693_), .A2(new_n2702_), .ZN(new_n2703_));
  NOR2_X1    g02510(.A1(new_n2693_), .A2(new_n2702_), .ZN(new_n2704_));
  INV_X1     g02511(.I(new_n2704_), .ZN(new_n2705_));
  AOI21_X1   g02512(.A1(new_n2705_), .A2(new_n2703_), .B(new_n2690_), .ZN(new_n2706_));
  INV_X1     g02513(.I(new_n2706_), .ZN(new_n2707_));
  NAND3_X1   g02514(.A1(new_n2705_), .A2(new_n2690_), .A3(new_n2703_), .ZN(new_n2708_));
  NAND2_X1   g02515(.A1(new_n2707_), .A2(new_n2708_), .ZN(new_n2709_));
  NAND2_X1   g02516(.A1(new_n2498_), .A2(new_n2513_), .ZN(new_n2710_));
  NAND2_X1   g02517(.A1(new_n2514_), .A2(new_n2582_), .ZN(new_n2711_));
  NAND2_X1   g02518(.A1(new_n2711_), .A2(new_n2710_), .ZN(new_n2712_));
  NOR2_X1    g02519(.A1(new_n2580_), .A2(new_n2577_), .ZN(new_n2713_));
  NAND2_X1   g02520(.A1(new_n2532_), .A2(new_n2522_), .ZN(new_n2714_));
  NAND2_X1   g02521(.A1(new_n2533_), .A2(new_n2541_), .ZN(new_n2715_));
  NAND2_X1   g02522(.A1(new_n2715_), .A2(new_n2714_), .ZN(new_n2716_));
  NAND2_X1   g02523(.A1(new_n2500_), .A2(new_n2499_), .ZN(new_n2717_));
  OAI21_X1   g02524(.A1(new_n2388_), .A2(new_n2407_), .B(new_n2717_), .ZN(new_n2718_));
  INV_X1     g02525(.I(new_n2509_), .ZN(new_n2719_));
  NAND2_X1   g02526(.A1(new_n2719_), .A2(new_n2418_), .ZN(new_n2720_));
  NAND2_X1   g02527(.A1(new_n2510_), .A2(new_n2399_), .ZN(new_n2721_));
  NAND2_X1   g02528(.A1(new_n2721_), .A2(new_n2720_), .ZN(new_n2722_));
  XOR2_X1    g02529(.A1(new_n2718_), .A2(new_n2722_), .Z(new_n2723_));
  XOR2_X1    g02530(.A1(new_n2723_), .A2(new_n2716_), .Z(new_n2724_));
  NAND2_X1   g02531(.A1(new_n2505_), .A2(new_n2511_), .ZN(new_n2725_));
  NAND2_X1   g02532(.A1(new_n2512_), .A2(new_n2501_), .ZN(new_n2726_));
  NAND2_X1   g02533(.A1(new_n2726_), .A2(new_n2725_), .ZN(new_n2727_));
  XOR2_X1    g02534(.A1(new_n2727_), .A2(new_n2724_), .Z(new_n2728_));
  XNOR2_X1   g02535(.A1(new_n2713_), .A2(new_n2728_), .ZN(new_n2729_));
  NOR2_X1    g02536(.A1(new_n2712_), .A2(new_n2729_), .ZN(new_n2730_));
  NAND2_X1   g02537(.A1(new_n2712_), .A2(new_n2729_), .ZN(new_n2731_));
  INV_X1     g02538(.I(new_n2731_), .ZN(new_n2732_));
  NOR2_X1    g02539(.A1(new_n2732_), .A2(new_n2730_), .ZN(new_n2733_));
  XNOR2_X1   g02540(.A1(new_n2733_), .A2(new_n2709_), .ZN(new_n2734_));
  NOR2_X1    g02541(.A1(new_n2734_), .A2(new_n2622_), .ZN(new_n2735_));
  INV_X1     g02542(.I(new_n2735_), .ZN(new_n2736_));
  NAND2_X1   g02543(.A1(new_n2734_), .A2(new_n2622_), .ZN(new_n2737_));
  NAND2_X1   g02544(.A1(new_n2736_), .A2(new_n2737_), .ZN(new_n2738_));
  XOR2_X1    g02545(.A1(new_n2620_), .A2(new_n2738_), .Z(\asquared[37] ));
  OAI21_X1   g02546(.A1(new_n2619_), .A2(new_n2614_), .B(new_n2736_), .ZN(new_n2740_));
  NAND2_X1   g02547(.A1(new_n2740_), .A2(new_n2737_), .ZN(new_n2741_));
  AOI22_X1   g02548(.A1(\a[2] ), .A2(\a[35] ), .B1(\a[3] ), .B2(\a[34] ), .ZN(new_n2742_));
  NOR2_X1    g02549(.A1(new_n742_), .A2(new_n1220_), .ZN(new_n2743_));
  INV_X1     g02550(.I(new_n2743_), .ZN(new_n2744_));
  NOR2_X1    g02551(.A1(new_n2442_), .A2(new_n2524_), .ZN(new_n2745_));
  INV_X1     g02552(.I(new_n2745_), .ZN(new_n2746_));
  NOR2_X1    g02553(.A1(new_n2746_), .A2(new_n246_), .ZN(new_n2747_));
  NOR3_X1    g02554(.A1(new_n2747_), .A2(new_n2742_), .A3(new_n2744_), .ZN(new_n2748_));
  NOR2_X1    g02555(.A1(new_n2748_), .A2(new_n2747_), .ZN(new_n2749_));
  INV_X1     g02556(.I(new_n2749_), .ZN(new_n2750_));
  OAI22_X1   g02557(.A1(new_n2750_), .A2(new_n2742_), .B1(new_n2744_), .B2(new_n2748_), .ZN(new_n2751_));
  INV_X1     g02558(.I(\a[37] ), .ZN(new_n2752_));
  AOI22_X1   g02559(.A1(\a[25] ), .A2(new_n537_), .B1(new_n980_), .B2(\a[33] ), .ZN(new_n2753_));
  NAND2_X1   g02560(.A1(\a[25] ), .A2(\a[33] ), .ZN(new_n2754_));
  NOR2_X1    g02561(.A1(new_n758_), .A2(new_n2754_), .ZN(new_n2755_));
  NOR3_X1    g02562(.A1(new_n2753_), .A2(new_n2752_), .A3(new_n2755_), .ZN(new_n2756_));
  NAND2_X1   g02563(.A1(\a[0] ), .A2(\a[37] ), .ZN(new_n2757_));
  NOR2_X1    g02564(.A1(new_n2756_), .A2(new_n2755_), .ZN(new_n2758_));
  INV_X1     g02565(.I(new_n2758_), .ZN(new_n2759_));
  AOI22_X1   g02566(.A1(\a[4] ), .A2(\a[33] ), .B1(\a[12] ), .B2(\a[25] ), .ZN(new_n2760_));
  OAI22_X1   g02567(.A1(new_n2759_), .A2(new_n2760_), .B1(new_n2756_), .B2(new_n2757_), .ZN(new_n2761_));
  XNOR2_X1   g02568(.A1(new_n2751_), .A2(new_n2761_), .ZN(new_n2762_));
  NAND2_X1   g02569(.A1(\a[9] ), .A2(\a[28] ), .ZN(new_n2763_));
  NOR2_X1    g02570(.A1(new_n2438_), .A2(new_n374_), .ZN(new_n2764_));
  NAND4_X1   g02571(.A1(\a[6] ), .A2(\a[9] ), .A3(\a[28] ), .A4(\a[31] ), .ZN(new_n2765_));
  NAND2_X1   g02572(.A1(new_n2681_), .A2(new_n1290_), .ZN(new_n2766_));
  AOI21_X1   g02573(.A1(new_n2765_), .A2(new_n2766_), .B(new_n2764_), .ZN(new_n2767_));
  AOI22_X1   g02574(.A1(\a[6] ), .A2(\a[31] ), .B1(\a[7] ), .B2(\a[30] ), .ZN(new_n2768_));
  NOR2_X1    g02575(.A1(new_n2767_), .A2(new_n2764_), .ZN(new_n2769_));
  INV_X1     g02576(.I(new_n2769_), .ZN(new_n2770_));
  OAI22_X1   g02577(.A1(new_n2770_), .A2(new_n2768_), .B1(new_n2763_), .B2(new_n2767_), .ZN(new_n2771_));
  XOR2_X1    g02578(.A1(new_n2762_), .A2(new_n2771_), .Z(new_n2772_));
  NAND2_X1   g02579(.A1(new_n2718_), .A2(new_n2722_), .ZN(new_n2773_));
  NAND2_X1   g02580(.A1(new_n2723_), .A2(new_n2716_), .ZN(new_n2774_));
  NAND2_X1   g02581(.A1(new_n2774_), .A2(new_n2773_), .ZN(new_n2775_));
  NAND2_X1   g02582(.A1(new_n2521_), .A2(new_n2540_), .ZN(new_n2776_));
  NAND2_X1   g02583(.A1(new_n2698_), .A2(new_n2530_), .ZN(new_n2777_));
  NAND2_X1   g02584(.A1(new_n2777_), .A2(new_n2776_), .ZN(new_n2778_));
  NAND2_X1   g02585(.A1(\a[10] ), .A2(\a[32] ), .ZN(new_n2779_));
  NOR3_X1    g02586(.A1(new_n2779_), .A2(new_n253_), .A3(new_n1750_), .ZN(new_n2780_));
  INV_X1     g02587(.I(new_n2780_), .ZN(new_n2781_));
  NOR2_X1    g02588(.A1(new_n1566_), .A2(new_n2200_), .ZN(new_n2782_));
  NAND2_X1   g02589(.A1(new_n2782_), .A2(new_n744_), .ZN(new_n2783_));
  OAI21_X1   g02590(.A1(new_n1264_), .A2(new_n1972_), .B(new_n2783_), .ZN(new_n2784_));
  NAND2_X1   g02591(.A1(new_n2784_), .A2(new_n2781_), .ZN(new_n2785_));
  NAND3_X1   g02592(.A1(new_n2785_), .A2(\a[11] ), .A3(\a[26] ), .ZN(new_n2786_));
  AOI22_X1   g02593(.A1(\a[5] ), .A2(\a[32] ), .B1(\a[10] ), .B2(\a[27] ), .ZN(new_n2787_));
  NAND2_X1   g02594(.A1(new_n2785_), .A2(new_n2781_), .ZN(new_n2788_));
  OAI21_X1   g02595(.A1(new_n2787_), .A2(new_n2788_), .B(new_n2786_), .ZN(new_n2789_));
  NAND2_X1   g02596(.A1(new_n1092_), .A2(new_n1276_), .ZN(new_n2790_));
  INV_X1     g02597(.I(new_n2790_), .ZN(new_n2791_));
  NOR2_X1    g02598(.A1(new_n1275_), .A2(new_n1376_), .ZN(new_n2792_));
  INV_X1     g02599(.I(new_n2792_), .ZN(new_n2793_));
  NOR2_X1    g02600(.A1(new_n355_), .A2(new_n1814_), .ZN(new_n2794_));
  INV_X1     g02601(.I(new_n2794_), .ZN(new_n2795_));
  OAI21_X1   g02602(.A1(new_n2791_), .A2(new_n2795_), .B(new_n2793_), .ZN(new_n2796_));
  NOR2_X1    g02603(.A1(new_n2796_), .A2(new_n2791_), .ZN(new_n2797_));
  AOI21_X1   g02604(.A1(new_n2793_), .A2(new_n2790_), .B(new_n2795_), .ZN(new_n2798_));
  NOR2_X1    g02605(.A1(new_n2797_), .A2(new_n2798_), .ZN(new_n2799_));
  XNOR2_X1   g02606(.A1(new_n2799_), .A2(new_n2789_), .ZN(new_n2800_));
  XOR2_X1    g02607(.A1(new_n2800_), .A2(new_n2778_), .Z(new_n2801_));
  XOR2_X1    g02608(.A1(new_n2775_), .A2(new_n2801_), .Z(new_n2802_));
  XOR2_X1    g02609(.A1(new_n2802_), .A2(new_n2772_), .Z(new_n2803_));
  NAND2_X1   g02610(.A1(new_n2727_), .A2(new_n2724_), .ZN(new_n2804_));
  INV_X1     g02611(.I(new_n2728_), .ZN(new_n2805_));
  OAI21_X1   g02612(.A1(new_n2805_), .A2(new_n2713_), .B(new_n2804_), .ZN(new_n2806_));
  NAND2_X1   g02613(.A1(new_n2507_), .A2(new_n2627_), .ZN(new_n2807_));
  NAND2_X1   g02614(.A1(new_n2628_), .A2(new_n2631_), .ZN(new_n2808_));
  NAND2_X1   g02615(.A1(new_n2808_), .A2(new_n2807_), .ZN(new_n2809_));
  XNOR2_X1   g02616(.A1(new_n2666_), .A2(new_n2809_), .ZN(new_n2810_));
  NOR2_X1    g02617(.A1(new_n1173_), .A2(new_n2385_), .ZN(new_n2811_));
  AOI22_X1   g02618(.A1(new_n760_), .A2(new_n1528_), .B1(new_n1879_), .B2(new_n1101_), .ZN(new_n2812_));
  NOR2_X1    g02619(.A1(new_n2811_), .A2(new_n2812_), .ZN(new_n2813_));
  NAND2_X1   g02620(.A1(\a[13] ), .A2(\a[24] ), .ZN(new_n2814_));
  AOI22_X1   g02621(.A1(\a[14] ), .A2(\a[23] ), .B1(\a[15] ), .B2(\a[22] ), .ZN(new_n2815_));
  NOR2_X1    g02622(.A1(new_n2813_), .A2(new_n2811_), .ZN(new_n2816_));
  INV_X1     g02623(.I(new_n2816_), .ZN(new_n2817_));
  OAI22_X1   g02624(.A1(new_n2817_), .A2(new_n2815_), .B1(new_n2813_), .B2(new_n2814_), .ZN(new_n2818_));
  XNOR2_X1   g02625(.A1(new_n2810_), .A2(new_n2818_), .ZN(new_n2819_));
  NOR2_X1    g02626(.A1(new_n2654_), .A2(new_n2642_), .ZN(new_n2820_));
  NAND2_X1   g02627(.A1(new_n2654_), .A2(new_n2642_), .ZN(new_n2821_));
  INV_X1     g02628(.I(new_n2821_), .ZN(new_n2822_));
  NOR2_X1    g02629(.A1(new_n2822_), .A2(new_n2820_), .ZN(new_n2823_));
  NOR2_X1    g02630(.A1(new_n2823_), .A2(new_n2675_), .ZN(new_n2824_));
  INV_X1     g02631(.I(new_n2823_), .ZN(new_n2825_));
  NOR2_X1    g02632(.A1(new_n2825_), .A2(new_n2674_), .ZN(new_n2826_));
  NOR2_X1    g02633(.A1(new_n2826_), .A2(new_n2824_), .ZN(new_n2827_));
  NAND2_X1   g02634(.A1(new_n2655_), .A2(new_n2644_), .ZN(new_n2828_));
  NAND2_X1   g02635(.A1(new_n2656_), .A2(new_n2632_), .ZN(new_n2829_));
  NAND2_X1   g02636(.A1(new_n2829_), .A2(new_n2828_), .ZN(new_n2830_));
  XOR2_X1    g02637(.A1(new_n2830_), .A2(new_n2827_), .Z(new_n2831_));
  XOR2_X1    g02638(.A1(new_n2831_), .A2(new_n2819_), .Z(new_n2832_));
  INV_X1     g02639(.I(new_n2832_), .ZN(new_n2833_));
  XOR2_X1    g02640(.A1(new_n2806_), .A2(new_n2833_), .Z(new_n2834_));
  INV_X1     g02641(.I(new_n2834_), .ZN(new_n2835_));
  OR2_X2     g02642(.A1(new_n2835_), .A2(new_n2803_), .Z(new_n2836_));
  NAND2_X1   g02643(.A1(new_n2835_), .A2(new_n2803_), .ZN(new_n2837_));
  AND2_X2    g02644(.A1(new_n2836_), .A2(new_n2837_), .Z(new_n2838_));
  INV_X1     g02645(.I(new_n2838_), .ZN(new_n2839_));
  NAND2_X1   g02646(.A1(new_n2693_), .A2(new_n2701_), .ZN(new_n2840_));
  NAND2_X1   g02647(.A1(new_n2707_), .A2(new_n2840_), .ZN(new_n2841_));
  INV_X1     g02648(.I(new_n2841_), .ZN(new_n2842_));
  NAND2_X1   g02649(.A1(new_n2625_), .A2(new_n2657_), .ZN(new_n2843_));
  NAND2_X1   g02650(.A1(new_n2658_), .A2(new_n2689_), .ZN(new_n2844_));
  NAND2_X1   g02651(.A1(new_n2844_), .A2(new_n2843_), .ZN(new_n2845_));
  NAND2_X1   g02652(.A1(new_n2669_), .A2(new_n2677_), .ZN(new_n2846_));
  NAND2_X1   g02653(.A1(new_n2678_), .A2(new_n2688_), .ZN(new_n2847_));
  NAND2_X1   g02654(.A1(new_n2847_), .A2(new_n2846_), .ZN(new_n2848_));
  NAND2_X1   g02655(.A1(new_n2694_), .A2(new_n2553_), .ZN(new_n2849_));
  OAI21_X1   g02656(.A1(new_n2561_), .A2(new_n2570_), .B(new_n2849_), .ZN(new_n2850_));
  INV_X1     g02657(.I(new_n2629_), .ZN(new_n2851_));
  NOR2_X1    g02658(.A1(new_n2851_), .A2(new_n2630_), .ZN(new_n2852_));
  AOI21_X1   g02659(.A1(\a[1] ), .A2(\a[36] ), .B(\a[19] ), .ZN(new_n2853_));
  NOR2_X1    g02660(.A1(new_n1064_), .A2(new_n2626_), .ZN(new_n2854_));
  NOR2_X1    g02661(.A1(new_n2854_), .A2(new_n2853_), .ZN(new_n2855_));
  INV_X1     g02662(.I(new_n2855_), .ZN(new_n2856_));
  NOR2_X1    g02663(.A1(new_n2856_), .A2(new_n2852_), .ZN(new_n2857_));
  INV_X1     g02664(.I(new_n2852_), .ZN(new_n2858_));
  NOR2_X1    g02665(.A1(new_n2855_), .A2(new_n2858_), .ZN(new_n2859_));
  OAI21_X1   g02666(.A1(new_n2859_), .A2(new_n2857_), .B(new_n2687_), .ZN(new_n2860_));
  OR3_X2     g02667(.A1(new_n2687_), .A2(new_n2857_), .A3(new_n2859_), .Z(new_n2861_));
  NAND2_X1   g02668(.A1(new_n2861_), .A2(new_n2860_), .ZN(new_n2862_));
  XNOR2_X1   g02669(.A1(new_n2850_), .A2(new_n2862_), .ZN(new_n2863_));
  XOR2_X1    g02670(.A1(new_n2848_), .A2(new_n2863_), .Z(new_n2864_));
  NAND2_X1   g02671(.A1(new_n2697_), .A2(new_n2699_), .ZN(new_n2865_));
  NAND2_X1   g02672(.A1(new_n2700_), .A2(new_n2695_), .ZN(new_n2866_));
  NAND2_X1   g02673(.A1(new_n2866_), .A2(new_n2865_), .ZN(new_n2867_));
  XOR2_X1    g02674(.A1(new_n2867_), .A2(new_n2864_), .Z(new_n2868_));
  XOR2_X1    g02675(.A1(new_n2845_), .A2(new_n2868_), .Z(new_n2869_));
  NOR2_X1    g02676(.A1(new_n2842_), .A2(new_n2869_), .ZN(new_n2870_));
  INV_X1     g02677(.I(new_n2869_), .ZN(new_n2871_));
  NOR2_X1    g02678(.A1(new_n2841_), .A2(new_n2871_), .ZN(new_n2872_));
  NOR2_X1    g02679(.A1(new_n2870_), .A2(new_n2872_), .ZN(new_n2873_));
  NOR2_X1    g02680(.A1(new_n2839_), .A2(new_n2873_), .ZN(new_n2874_));
  NOR3_X1    g02681(.A1(new_n2838_), .A2(new_n2870_), .A3(new_n2872_), .ZN(new_n2875_));
  NOR2_X1    g02682(.A1(new_n2874_), .A2(new_n2875_), .ZN(new_n2876_));
  INV_X1     g02683(.I(new_n2876_), .ZN(new_n2877_));
  INV_X1     g02684(.I(new_n2733_), .ZN(new_n2878_));
  NOR2_X1    g02685(.A1(new_n2878_), .A2(new_n2709_), .ZN(new_n2879_));
  NOR2_X1    g02686(.A1(new_n2879_), .A2(new_n2732_), .ZN(new_n2880_));
  NOR2_X1    g02687(.A1(new_n2877_), .A2(new_n2880_), .ZN(new_n2881_));
  NAND2_X1   g02688(.A1(new_n2877_), .A2(new_n2880_), .ZN(new_n2882_));
  INV_X1     g02689(.I(new_n2882_), .ZN(new_n2883_));
  NOR2_X1    g02690(.A1(new_n2883_), .A2(new_n2881_), .ZN(new_n2884_));
  XOR2_X1    g02691(.A1(new_n2741_), .A2(new_n2884_), .Z(\asquared[38] ));
  AOI21_X1   g02692(.A1(new_n2740_), .A2(new_n2737_), .B(new_n2883_), .ZN(new_n2886_));
  NOR2_X1    g02693(.A1(new_n2886_), .A2(new_n2881_), .ZN(new_n2887_));
  AOI21_X1   g02694(.A1(new_n2841_), .A2(new_n2869_), .B(new_n2874_), .ZN(new_n2888_));
  NOR2_X1    g02695(.A1(new_n2826_), .A2(new_n2822_), .ZN(new_n2889_));
  NOR2_X1    g02696(.A1(new_n536_), .A2(new_n2442_), .ZN(new_n2890_));
  AOI22_X1   g02697(.A1(new_n1974_), .A2(new_n2890_), .B1(new_n1971_), .B2(new_n1261_), .ZN(new_n2891_));
  NOR4_X1    g02698(.A1(new_n290_), .A2(new_n513_), .A3(new_n1750_), .A4(new_n2442_), .ZN(new_n2892_));
  NOR2_X1    g02699(.A1(new_n2891_), .A2(new_n2892_), .ZN(new_n2893_));
  NAND2_X1   g02700(.A1(\a[12] ), .A2(\a[26] ), .ZN(new_n2894_));
  AOI22_X1   g02701(.A1(\a[4] ), .A2(\a[34] ), .B1(\a[11] ), .B2(\a[27] ), .ZN(new_n2895_));
  INV_X1     g02702(.I(new_n2892_), .ZN(new_n2896_));
  NAND2_X1   g02703(.A1(new_n2891_), .A2(new_n2896_), .ZN(new_n2897_));
  OAI22_X1   g02704(.A1(new_n2893_), .A2(new_n2894_), .B1(new_n2897_), .B2(new_n2895_), .ZN(new_n2898_));
  OAI21_X1   g02705(.A1(new_n2858_), .A2(new_n2856_), .B(new_n2860_), .ZN(new_n2899_));
  XNOR2_X1   g02706(.A1(new_n2899_), .A2(new_n2898_), .ZN(new_n2900_));
  XOR2_X1    g02707(.A1(new_n2889_), .A2(new_n2900_), .Z(new_n2901_));
  NAND3_X1   g02708(.A1(new_n2850_), .A2(new_n2860_), .A3(new_n2861_), .ZN(new_n2902_));
  NAND2_X1   g02709(.A1(new_n2848_), .A2(new_n2863_), .ZN(new_n2903_));
  NAND2_X1   g02710(.A1(new_n2903_), .A2(new_n2902_), .ZN(new_n2904_));
  AOI22_X1   g02711(.A1(\a[13] ), .A2(\a[25] ), .B1(\a[14] ), .B2(\a[24] ), .ZN(new_n2905_));
  NAND2_X1   g02712(.A1(\a[3] ), .A2(\a[35] ), .ZN(new_n2906_));
  NOR2_X1    g02713(.A1(new_n767_), .A2(new_n1779_), .ZN(new_n2907_));
  NOR3_X1    g02714(.A1(new_n2907_), .A2(new_n2905_), .A3(new_n2906_), .ZN(new_n2908_));
  NOR2_X1    g02715(.A1(new_n2908_), .A2(new_n2907_), .ZN(new_n2909_));
  INV_X1     g02716(.I(new_n2909_), .ZN(new_n2910_));
  OAI22_X1   g02717(.A1(new_n2910_), .A2(new_n2905_), .B1(new_n2906_), .B2(new_n2908_), .ZN(new_n2911_));
  AOI22_X1   g02718(.A1(\a[0] ), .A2(\a[38] ), .B1(\a[2] ), .B2(\a[36] ), .ZN(new_n2912_));
  INV_X1     g02719(.I(new_n2912_), .ZN(new_n2913_));
  INV_X1     g02720(.I(\a[38] ), .ZN(new_n2914_));
  NOR2_X1    g02721(.A1(new_n2626_), .A2(new_n2914_), .ZN(new_n2915_));
  INV_X1     g02722(.I(new_n2915_), .ZN(new_n2916_));
  NOR2_X1    g02723(.A1(new_n2916_), .A2(new_n412_), .ZN(new_n2917_));
  AOI21_X1   g02724(.A1(new_n2854_), .A2(new_n2913_), .B(new_n2917_), .ZN(new_n2918_));
  INV_X1     g02725(.I(new_n2918_), .ZN(new_n2919_));
  OAI21_X1   g02726(.A1(new_n2917_), .A2(new_n2912_), .B(new_n2854_), .ZN(new_n2920_));
  OAI21_X1   g02727(.A1(new_n2919_), .A2(new_n2912_), .B(new_n2920_), .ZN(new_n2921_));
  XOR2_X1    g02728(.A1(new_n2921_), .A2(new_n2788_), .Z(new_n2922_));
  XOR2_X1    g02729(.A1(new_n2922_), .A2(new_n2911_), .Z(new_n2923_));
  XOR2_X1    g02730(.A1(new_n2904_), .A2(new_n2923_), .Z(new_n2924_));
  XNOR2_X1   g02731(.A1(new_n2924_), .A2(new_n2901_), .ZN(new_n2925_));
  NAND2_X1   g02732(.A1(new_n2867_), .A2(new_n2864_), .ZN(new_n2926_));
  NAND2_X1   g02733(.A1(new_n2845_), .A2(new_n2868_), .ZN(new_n2927_));
  NAND2_X1   g02734(.A1(new_n2927_), .A2(new_n2926_), .ZN(new_n2928_));
  NAND2_X1   g02735(.A1(\a[1] ), .A2(\a[37] ), .ZN(new_n2929_));
  XNOR2_X1   g02736(.A1(new_n1273_), .A2(new_n2929_), .ZN(new_n2930_));
  XOR2_X1    g02737(.A1(new_n2796_), .A2(new_n2930_), .Z(new_n2931_));
  OR2_X2     g02738(.A1(new_n2931_), .A2(new_n2770_), .Z(new_n2932_));
  NAND2_X1   g02739(.A1(new_n2931_), .A2(new_n2770_), .ZN(new_n2933_));
  AND2_X2    g02740(.A1(new_n2932_), .A2(new_n2933_), .Z(new_n2934_));
  NAND2_X1   g02741(.A1(new_n2751_), .A2(new_n2761_), .ZN(new_n2935_));
  INV_X1     g02742(.I(new_n2762_), .ZN(new_n2936_));
  NAND2_X1   g02743(.A1(new_n2936_), .A2(new_n2771_), .ZN(new_n2937_));
  NAND2_X1   g02744(.A1(new_n2937_), .A2(new_n2935_), .ZN(new_n2938_));
  NAND2_X1   g02745(.A1(new_n2667_), .A2(new_n2809_), .ZN(new_n2939_));
  NAND2_X1   g02746(.A1(new_n2810_), .A2(new_n2818_), .ZN(new_n2940_));
  NAND2_X1   g02747(.A1(new_n2940_), .A2(new_n2939_), .ZN(new_n2941_));
  XOR2_X1    g02748(.A1(new_n2938_), .A2(new_n2941_), .Z(new_n2942_));
  XOR2_X1    g02749(.A1(new_n2942_), .A2(new_n2934_), .Z(new_n2943_));
  XOR2_X1    g02750(.A1(new_n2928_), .A2(new_n2943_), .Z(new_n2944_));
  XNOR2_X1   g02751(.A1(new_n2944_), .A2(new_n2925_), .ZN(new_n2945_));
  NAND2_X1   g02752(.A1(new_n2806_), .A2(new_n2833_), .ZN(new_n2946_));
  NAND2_X1   g02753(.A1(new_n2836_), .A2(new_n2946_), .ZN(new_n2947_));
  NOR2_X1    g02754(.A1(new_n2775_), .A2(new_n2801_), .ZN(new_n2948_));
  NAND2_X1   g02755(.A1(new_n2775_), .A2(new_n2801_), .ZN(new_n2949_));
  OAI21_X1   g02756(.A1(new_n2772_), .A2(new_n2948_), .B(new_n2949_), .ZN(new_n2950_));
  NAND2_X1   g02757(.A1(new_n2830_), .A2(new_n2827_), .ZN(new_n2951_));
  INV_X1     g02758(.I(new_n2831_), .ZN(new_n2952_));
  OAI21_X1   g02759(.A1(new_n2952_), .A2(new_n2819_), .B(new_n2951_), .ZN(new_n2953_));
  XNOR2_X1   g02760(.A1(new_n2953_), .A2(new_n2950_), .ZN(new_n2954_));
  NAND2_X1   g02761(.A1(new_n1024_), .A2(new_n1452_), .ZN(new_n2955_));
  NOR4_X1    g02762(.A1(new_n717_), .A2(new_n1023_), .A3(new_n1220_), .A4(new_n1299_), .ZN(new_n2956_));
  NOR2_X1    g02763(.A1(new_n2385_), .A2(new_n893_), .ZN(new_n2957_));
  OAI21_X1   g02764(.A1(new_n2957_), .A2(new_n2956_), .B(new_n2955_), .ZN(new_n2958_));
  NAND3_X1   g02765(.A1(new_n2958_), .A2(\a[15] ), .A3(\a[23] ), .ZN(new_n2959_));
  AOI22_X1   g02766(.A1(\a[16] ), .A2(\a[22] ), .B1(\a[17] ), .B2(\a[21] ), .ZN(new_n2960_));
  NAND2_X1   g02767(.A1(new_n2958_), .A2(new_n2955_), .ZN(new_n2961_));
  OAI21_X1   g02768(.A1(new_n2960_), .A2(new_n2961_), .B(new_n2959_), .ZN(new_n2962_));
  NOR2_X1    g02769(.A1(new_n367_), .A2(new_n2200_), .ZN(new_n2963_));
  NOR2_X1    g02770(.A1(new_n417_), .A2(new_n1718_), .ZN(new_n2964_));
  NOR2_X1    g02771(.A1(new_n2963_), .A2(new_n2964_), .ZN(new_n2965_));
  NOR2_X1    g02772(.A1(new_n253_), .A2(new_n2274_), .ZN(new_n2966_));
  INV_X1     g02773(.I(new_n2966_), .ZN(new_n2967_));
  NOR2_X1    g02774(.A1(new_n2637_), .A2(new_n371_), .ZN(new_n2968_));
  AOI21_X1   g02775(.A1(new_n2964_), .A2(new_n2966_), .B(new_n2968_), .ZN(new_n2969_));
  AOI21_X1   g02776(.A1(new_n2963_), .A2(new_n2964_), .B(new_n2969_), .ZN(new_n2970_));
  AOI21_X1   g02777(.A1(new_n2963_), .A2(new_n2964_), .B(new_n2970_), .ZN(new_n2971_));
  INV_X1     g02778(.I(new_n2971_), .ZN(new_n2972_));
  OAI22_X1   g02779(.A1(new_n2972_), .A2(new_n2965_), .B1(new_n2967_), .B2(new_n2970_), .ZN(new_n2973_));
  XNOR2_X1   g02780(.A1(new_n2973_), .A2(new_n2962_), .ZN(new_n2974_));
  NAND2_X1   g02781(.A1(new_n467_), .A2(new_n2254_), .ZN(new_n2975_));
  NOR2_X1    g02782(.A1(new_n1814_), .A2(new_n2051_), .ZN(new_n2976_));
  NAND2_X1   g02783(.A1(new_n2976_), .A2(new_n1290_), .ZN(new_n2977_));
  AOI22_X1   g02784(.A1(new_n2975_), .A2(new_n2977_), .B1(new_n693_), .B2(new_n2437_), .ZN(new_n2978_));
  NAND2_X1   g02785(.A1(\a[9] ), .A2(\a[29] ), .ZN(new_n2979_));
  AOI22_X1   g02786(.A1(\a[7] ), .A2(\a[31] ), .B1(\a[8] ), .B2(\a[30] ), .ZN(new_n2980_));
  NAND2_X1   g02787(.A1(new_n2437_), .A2(new_n693_), .ZN(new_n2981_));
  NAND3_X1   g02788(.A1(new_n2981_), .A2(new_n2975_), .A3(new_n2977_), .ZN(new_n2982_));
  OAI22_X1   g02789(.A1(new_n2978_), .A2(new_n2979_), .B1(new_n2982_), .B2(new_n2980_), .ZN(new_n2983_));
  XOR2_X1    g02790(.A1(new_n2974_), .A2(new_n2983_), .Z(new_n2984_));
  INV_X1     g02791(.I(new_n2984_), .ZN(new_n2985_));
  NOR2_X1    g02792(.A1(new_n2750_), .A2(new_n2759_), .ZN(new_n2986_));
  NOR2_X1    g02793(.A1(new_n2749_), .A2(new_n2758_), .ZN(new_n2987_));
  NOR2_X1    g02794(.A1(new_n2986_), .A2(new_n2987_), .ZN(new_n2988_));
  INV_X1     g02795(.I(new_n2988_), .ZN(new_n2989_));
  NOR2_X1    g02796(.A1(new_n2989_), .A2(new_n2816_), .ZN(new_n2990_));
  NOR2_X1    g02797(.A1(new_n2988_), .A2(new_n2817_), .ZN(new_n2991_));
  NOR2_X1    g02798(.A1(new_n2990_), .A2(new_n2991_), .ZN(new_n2992_));
  OAI21_X1   g02799(.A1(new_n2797_), .A2(new_n2798_), .B(new_n2789_), .ZN(new_n2993_));
  NAND2_X1   g02800(.A1(new_n2800_), .A2(new_n2778_), .ZN(new_n2994_));
  NAND2_X1   g02801(.A1(new_n2994_), .A2(new_n2993_), .ZN(new_n2995_));
  NAND2_X1   g02802(.A1(new_n2995_), .A2(new_n2992_), .ZN(new_n2996_));
  INV_X1     g02803(.I(new_n2996_), .ZN(new_n2997_));
  NOR2_X1    g02804(.A1(new_n2995_), .A2(new_n2992_), .ZN(new_n2998_));
  NOR2_X1    g02805(.A1(new_n2997_), .A2(new_n2998_), .ZN(new_n2999_));
  NOR2_X1    g02806(.A1(new_n2985_), .A2(new_n2999_), .ZN(new_n3000_));
  NAND2_X1   g02807(.A1(new_n2985_), .A2(new_n2999_), .ZN(new_n3001_));
  INV_X1     g02808(.I(new_n3001_), .ZN(new_n3002_));
  NOR2_X1    g02809(.A1(new_n3002_), .A2(new_n3000_), .ZN(new_n3003_));
  XNOR2_X1   g02810(.A1(new_n2954_), .A2(new_n3003_), .ZN(new_n3004_));
  NOR2_X1    g02811(.A1(new_n2947_), .A2(new_n3004_), .ZN(new_n3005_));
  NAND2_X1   g02812(.A1(new_n2947_), .A2(new_n3004_), .ZN(new_n3006_));
  INV_X1     g02813(.I(new_n3006_), .ZN(new_n3007_));
  NOR2_X1    g02814(.A1(new_n3007_), .A2(new_n3005_), .ZN(new_n3008_));
  NAND2_X1   g02815(.A1(new_n3008_), .A2(new_n2945_), .ZN(new_n3009_));
  INV_X1     g02816(.I(new_n3009_), .ZN(new_n3010_));
  NOR2_X1    g02817(.A1(new_n3008_), .A2(new_n2945_), .ZN(new_n3011_));
  NOR2_X1    g02818(.A1(new_n3010_), .A2(new_n3011_), .ZN(new_n3012_));
  INV_X1     g02819(.I(new_n3012_), .ZN(new_n3013_));
  NOR2_X1    g02820(.A1(new_n3013_), .A2(new_n2888_), .ZN(new_n3014_));
  INV_X1     g02821(.I(new_n3014_), .ZN(new_n3015_));
  NAND2_X1   g02822(.A1(new_n3013_), .A2(new_n2888_), .ZN(new_n3016_));
  NAND2_X1   g02823(.A1(new_n3015_), .A2(new_n3016_), .ZN(new_n3017_));
  XOR2_X1    g02824(.A1(new_n2887_), .A2(new_n3017_), .Z(\asquared[39] ));
  OAI21_X1   g02825(.A1(new_n2886_), .A2(new_n2881_), .B(new_n3016_), .ZN(new_n3019_));
  NAND2_X1   g02826(.A1(new_n3019_), .A2(new_n3015_), .ZN(new_n3020_));
  NOR2_X1    g02827(.A1(new_n3010_), .A2(new_n3007_), .ZN(new_n3021_));
  INV_X1     g02828(.I(new_n3021_), .ZN(new_n3022_));
  NOR2_X1    g02829(.A1(new_n3002_), .A2(new_n2997_), .ZN(new_n3023_));
  NAND2_X1   g02830(.A1(new_n2938_), .A2(new_n2941_), .ZN(new_n3024_));
  NAND2_X1   g02831(.A1(new_n2942_), .A2(new_n2934_), .ZN(new_n3025_));
  NAND2_X1   g02832(.A1(new_n3025_), .A2(new_n3024_), .ZN(new_n3026_));
  NAND2_X1   g02833(.A1(new_n1528_), .A2(new_n1288_), .ZN(new_n3027_));
  OAI22_X1   g02834(.A1(new_n2028_), .A2(new_n1443_), .B1(new_n1173_), .B2(new_n1779_), .ZN(new_n3028_));
  NAND2_X1   g02835(.A1(new_n3028_), .A2(new_n3027_), .ZN(new_n3029_));
  NAND3_X1   g02836(.A1(new_n3029_), .A2(\a[14] ), .A3(\a[25] ), .ZN(new_n3030_));
  AOI22_X1   g02837(.A1(\a[15] ), .A2(\a[24] ), .B1(\a[16] ), .B2(\a[23] ), .ZN(new_n3031_));
  NAND2_X1   g02838(.A1(new_n3029_), .A2(new_n3027_), .ZN(new_n3032_));
  OAI21_X1   g02839(.A1(new_n3031_), .A2(new_n3032_), .B(new_n3030_), .ZN(new_n3033_));
  NAND4_X1   g02840(.A1(\a[3] ), .A2(\a[13] ), .A3(\a[26] ), .A4(\a[36] ), .ZN(new_n3034_));
  NOR2_X1    g02841(.A1(new_n597_), .A2(new_n2752_), .ZN(new_n3035_));
  NAND2_X1   g02842(.A1(new_n1710_), .A2(new_n3035_), .ZN(new_n3036_));
  NOR2_X1    g02843(.A1(new_n2626_), .A2(new_n2752_), .ZN(new_n3037_));
  INV_X1     g02844(.I(new_n3037_), .ZN(new_n3038_));
  OAI21_X1   g02845(.A1(new_n246_), .A2(new_n3038_), .B(new_n3036_), .ZN(new_n3039_));
  NAND2_X1   g02846(.A1(new_n3039_), .A2(new_n3034_), .ZN(new_n3040_));
  NAND3_X1   g02847(.A1(new_n3040_), .A2(\a[2] ), .A3(\a[37] ), .ZN(new_n3041_));
  NAND2_X1   g02848(.A1(new_n3040_), .A2(new_n3034_), .ZN(new_n3042_));
  AOI22_X1   g02849(.A1(\a[3] ), .A2(\a[36] ), .B1(\a[13] ), .B2(\a[26] ), .ZN(new_n3043_));
  OAI21_X1   g02850(.A1(new_n3042_), .A2(new_n3043_), .B(new_n3041_), .ZN(new_n3044_));
  XNOR2_X1   g02851(.A1(new_n3044_), .A2(new_n3033_), .ZN(new_n3045_));
  NAND2_X1   g02852(.A1(\a[6] ), .A2(\a[33] ), .ZN(new_n3046_));
  NAND4_X1   g02853(.A1(\a[6] ), .A2(\a[9] ), .A3(\a[30] ), .A4(\a[33] ), .ZN(new_n3047_));
  NAND2_X1   g02854(.A1(new_n2636_), .A2(new_n479_), .ZN(new_n3048_));
  AOI22_X1   g02855(.A1(new_n3048_), .A2(new_n3047_), .B1(new_n1290_), .B2(new_n2201_), .ZN(new_n3049_));
  AOI22_X1   g02856(.A1(\a[7] ), .A2(\a[32] ), .B1(\a[9] ), .B2(\a[30] ), .ZN(new_n3050_));
  NAND2_X1   g02857(.A1(new_n2201_), .A2(new_n1290_), .ZN(new_n3051_));
  NAND3_X1   g02858(.A1(new_n3051_), .A2(new_n3048_), .A3(new_n3047_), .ZN(new_n3052_));
  OAI22_X1   g02859(.A1(new_n3049_), .A2(new_n3046_), .B1(new_n3052_), .B2(new_n3050_), .ZN(new_n3053_));
  XOR2_X1    g02860(.A1(new_n3045_), .A2(new_n3053_), .Z(new_n3054_));
  INV_X1     g02861(.I(new_n3054_), .ZN(new_n3055_));
  NOR2_X1    g02862(.A1(new_n3026_), .A2(new_n3055_), .ZN(new_n3056_));
  NAND2_X1   g02863(.A1(new_n3026_), .A2(new_n3055_), .ZN(new_n3057_));
  INV_X1     g02864(.I(new_n3057_), .ZN(new_n3058_));
  NOR2_X1    g02865(.A1(new_n3058_), .A2(new_n3056_), .ZN(new_n3059_));
  XNOR2_X1   g02866(.A1(new_n3059_), .A2(new_n3023_), .ZN(new_n3060_));
  INV_X1     g02867(.I(new_n3060_), .ZN(new_n3061_));
  NAND2_X1   g02868(.A1(new_n2953_), .A2(new_n2950_), .ZN(new_n3062_));
  INV_X1     g02869(.I(new_n3003_), .ZN(new_n3063_));
  OAI21_X1   g02870(.A1(new_n2954_), .A2(new_n3063_), .B(new_n3062_), .ZN(new_n3064_));
  NOR2_X1    g02871(.A1(new_n884_), .A2(new_n1220_), .ZN(new_n3065_));
  NOR2_X1    g02872(.A1(new_n1375_), .A2(new_n3065_), .ZN(new_n3066_));
  INV_X1     g02873(.I(new_n3066_), .ZN(new_n3067_));
  NOR2_X1    g02874(.A1(new_n1382_), .A2(new_n1092_), .ZN(new_n3068_));
  NOR2_X1    g02875(.A1(new_n355_), .A2(new_n2051_), .ZN(new_n3069_));
  AOI21_X1   g02876(.A1(new_n3067_), .A2(new_n3069_), .B(new_n3068_), .ZN(new_n3070_));
  INV_X1     g02877(.I(new_n3070_), .ZN(new_n3071_));
  OAI21_X1   g02878(.A1(new_n3068_), .A2(new_n3066_), .B(new_n3069_), .ZN(new_n3072_));
  OAI21_X1   g02879(.A1(new_n3071_), .A2(new_n3066_), .B(new_n3072_), .ZN(new_n3073_));
  AOI22_X1   g02880(.A1(\a[4] ), .A2(\a[35] ), .B1(\a[12] ), .B2(\a[27] ), .ZN(new_n3074_));
  INV_X1     g02881(.I(new_n3074_), .ZN(new_n3075_));
  NOR4_X1    g02882(.A1(new_n290_), .A2(new_n536_), .A3(new_n1750_), .A4(new_n2524_), .ZN(new_n3076_));
  NOR2_X1    g02883(.A1(new_n1023_), .A2(new_n1175_), .ZN(new_n3077_));
  AOI21_X1   g02884(.A1(new_n3075_), .A2(new_n3077_), .B(new_n3076_), .ZN(new_n3078_));
  INV_X1     g02885(.I(new_n3078_), .ZN(new_n3079_));
  OAI21_X1   g02886(.A1(new_n3076_), .A2(new_n3074_), .B(new_n3077_), .ZN(new_n3080_));
  OAI21_X1   g02887(.A1(new_n3079_), .A2(new_n3074_), .B(new_n3080_), .ZN(new_n3081_));
  XNOR2_X1   g02888(.A1(new_n3073_), .A2(new_n3081_), .ZN(new_n3082_));
  NOR4_X1    g02889(.A1(new_n253_), .A2(new_n417_), .A3(new_n1814_), .A4(new_n2442_), .ZN(new_n3083_));
  NOR2_X1    g02890(.A1(new_n253_), .A2(new_n2442_), .ZN(new_n3084_));
  AOI22_X1   g02891(.A1(new_n747_), .A2(new_n2105_), .B1(new_n1721_), .B2(new_n3084_), .ZN(new_n3085_));
  NOR2_X1    g02892(.A1(new_n3085_), .A2(new_n3083_), .ZN(new_n3086_));
  INV_X1     g02893(.I(new_n3083_), .ZN(new_n3087_));
  NAND2_X1   g02894(.A1(new_n3085_), .A2(new_n3087_), .ZN(new_n3088_));
  AOI21_X1   g02895(.A1(\a[10] ), .A2(\a[29] ), .B(new_n3084_), .ZN(new_n3089_));
  OAI22_X1   g02896(.A1(new_n1722_), .A2(new_n3086_), .B1(new_n3088_), .B2(new_n3089_), .ZN(new_n3090_));
  XOR2_X1    g02897(.A1(new_n3082_), .A2(new_n3090_), .Z(new_n3091_));
  INV_X1     g02898(.I(new_n3091_), .ZN(new_n3092_));
  NAND2_X1   g02899(.A1(new_n2899_), .A2(new_n2898_), .ZN(new_n3093_));
  OAI21_X1   g02900(.A1(new_n2889_), .A2(new_n2900_), .B(new_n3093_), .ZN(new_n3094_));
  XOR2_X1    g02901(.A1(new_n2897_), .A2(new_n2982_), .Z(new_n3095_));
  XNOR2_X1   g02902(.A1(new_n2971_), .A2(new_n3095_), .ZN(new_n3096_));
  NOR2_X1    g02903(.A1(new_n3094_), .A2(new_n3096_), .ZN(new_n3097_));
  NAND2_X1   g02904(.A1(new_n3094_), .A2(new_n3096_), .ZN(new_n3098_));
  INV_X1     g02905(.I(new_n3098_), .ZN(new_n3099_));
  NOR2_X1    g02906(.A1(new_n3099_), .A2(new_n3097_), .ZN(new_n3100_));
  NAND2_X1   g02907(.A1(new_n3100_), .A2(new_n3092_), .ZN(new_n3101_));
  INV_X1     g02908(.I(new_n3101_), .ZN(new_n3102_));
  NOR2_X1    g02909(.A1(new_n3100_), .A2(new_n3092_), .ZN(new_n3103_));
  NOR2_X1    g02910(.A1(new_n3102_), .A2(new_n3103_), .ZN(new_n3104_));
  XNOR2_X1   g02911(.A1(new_n3064_), .A2(new_n3104_), .ZN(new_n3105_));
  XOR2_X1    g02912(.A1(new_n3105_), .A2(new_n3061_), .Z(new_n3106_));
  NAND2_X1   g02913(.A1(new_n2928_), .A2(new_n2943_), .ZN(new_n3107_));
  INV_X1     g02914(.I(new_n2944_), .ZN(new_n3108_));
  OAI21_X1   g02915(.A1(new_n3108_), .A2(new_n2925_), .B(new_n3107_), .ZN(new_n3109_));
  NAND2_X1   g02916(.A1(new_n2904_), .A2(new_n2923_), .ZN(new_n3110_));
  NAND2_X1   g02917(.A1(new_n2924_), .A2(new_n2901_), .ZN(new_n3111_));
  NAND2_X1   g02918(.A1(new_n3111_), .A2(new_n3110_), .ZN(new_n3112_));
  NAND2_X1   g02919(.A1(new_n2796_), .A2(new_n2930_), .ZN(new_n3113_));
  NAND2_X1   g02920(.A1(new_n2933_), .A2(new_n3113_), .ZN(new_n3114_));
  NOR2_X1    g02921(.A1(new_n1281_), .A2(new_n2929_), .ZN(new_n3115_));
  INV_X1     g02922(.I(\a[39] ), .ZN(new_n3116_));
  NOR2_X1    g02923(.A1(new_n196_), .A2(new_n3116_), .ZN(new_n3117_));
  INV_X1     g02924(.I(new_n3117_), .ZN(new_n3118_));
  XOR2_X1    g02925(.A1(new_n3115_), .A2(new_n3118_), .Z(new_n3119_));
  NOR2_X1    g02926(.A1(new_n1137_), .A2(new_n2914_), .ZN(new_n3120_));
  INV_X1     g02927(.I(new_n3120_), .ZN(new_n3121_));
  NOR2_X1    g02928(.A1(new_n194_), .A2(new_n2914_), .ZN(new_n3122_));
  OAI21_X1   g02929(.A1(\a[20] ), .A2(new_n3122_), .B(new_n3121_), .ZN(new_n3123_));
  XNOR2_X1   g02930(.A1(new_n3119_), .A2(new_n3123_), .ZN(new_n3124_));
  INV_X1     g02931(.I(new_n3124_), .ZN(new_n3125_));
  XOR2_X1    g02932(.A1(new_n3114_), .A2(new_n3125_), .Z(new_n3126_));
  OAI21_X1   g02933(.A1(new_n2987_), .A2(new_n2990_), .B(new_n3126_), .ZN(new_n3127_));
  NOR2_X1    g02934(.A1(new_n2990_), .A2(new_n2987_), .ZN(new_n3128_));
  INV_X1     g02935(.I(new_n3126_), .ZN(new_n3129_));
  NAND2_X1   g02936(.A1(new_n3129_), .A2(new_n3128_), .ZN(new_n3130_));
  AND2_X2    g02937(.A1(new_n3130_), .A2(new_n3127_), .Z(new_n3131_));
  XOR2_X1    g02938(.A1(new_n2909_), .A2(new_n2918_), .Z(new_n3132_));
  XOR2_X1    g02939(.A1(new_n3132_), .A2(new_n2961_), .Z(new_n3133_));
  NAND2_X1   g02940(.A1(new_n2973_), .A2(new_n2962_), .ZN(new_n3134_));
  INV_X1     g02941(.I(new_n2974_), .ZN(new_n3135_));
  NAND2_X1   g02942(.A1(new_n3135_), .A2(new_n2983_), .ZN(new_n3136_));
  NAND2_X1   g02943(.A1(new_n3136_), .A2(new_n3134_), .ZN(new_n3137_));
  NAND2_X1   g02944(.A1(new_n2922_), .A2(new_n2911_), .ZN(new_n3138_));
  NAND2_X1   g02945(.A1(new_n2921_), .A2(new_n2788_), .ZN(new_n3139_));
  NAND2_X1   g02946(.A1(new_n3138_), .A2(new_n3139_), .ZN(new_n3140_));
  XOR2_X1    g02947(.A1(new_n3137_), .A2(new_n3140_), .Z(new_n3141_));
  NAND2_X1   g02948(.A1(new_n3141_), .A2(new_n3133_), .ZN(new_n3142_));
  OR2_X2     g02949(.A1(new_n3141_), .A2(new_n3133_), .Z(new_n3143_));
  AND2_X2    g02950(.A1(new_n3143_), .A2(new_n3142_), .Z(new_n3144_));
  XOR2_X1    g02951(.A1(new_n3144_), .A2(new_n3131_), .Z(new_n3145_));
  XOR2_X1    g02952(.A1(new_n3145_), .A2(new_n3112_), .Z(new_n3146_));
  NOR2_X1    g02953(.A1(new_n3146_), .A2(new_n3109_), .ZN(new_n3147_));
  NAND2_X1   g02954(.A1(new_n3146_), .A2(new_n3109_), .ZN(new_n3148_));
  INV_X1     g02955(.I(new_n3148_), .ZN(new_n3149_));
  NOR2_X1    g02956(.A1(new_n3149_), .A2(new_n3147_), .ZN(new_n3150_));
  NOR2_X1    g02957(.A1(new_n3150_), .A2(new_n3106_), .ZN(new_n3151_));
  NAND2_X1   g02958(.A1(new_n3150_), .A2(new_n3106_), .ZN(new_n3152_));
  INV_X1     g02959(.I(new_n3152_), .ZN(new_n3153_));
  NOR2_X1    g02960(.A1(new_n3153_), .A2(new_n3151_), .ZN(new_n3154_));
  NOR2_X1    g02961(.A1(new_n3022_), .A2(new_n3154_), .ZN(new_n3155_));
  NAND2_X1   g02962(.A1(new_n3022_), .A2(new_n3154_), .ZN(new_n3156_));
  INV_X1     g02963(.I(new_n3156_), .ZN(new_n3157_));
  NOR2_X1    g02964(.A1(new_n3157_), .A2(new_n3155_), .ZN(new_n3158_));
  XOR2_X1    g02965(.A1(new_n3020_), .A2(new_n3158_), .Z(\asquared[40] ));
  AOI21_X1   g02966(.A1(new_n3019_), .A2(new_n3015_), .B(new_n3155_), .ZN(new_n3160_));
  NOR2_X1    g02967(.A1(new_n3160_), .A2(new_n3157_), .ZN(new_n3161_));
  NAND2_X1   g02968(.A1(\a[1] ), .A2(\a[39] ), .ZN(new_n3162_));
  NOR2_X1    g02969(.A1(new_n1379_), .A2(new_n3162_), .ZN(new_n3163_));
  INV_X1     g02970(.I(new_n3163_), .ZN(new_n3164_));
  NAND2_X1   g02971(.A1(new_n1379_), .A2(new_n3162_), .ZN(new_n3165_));
  NAND2_X1   g02972(.A1(new_n3164_), .A2(new_n3165_), .ZN(new_n3166_));
  XOR2_X1    g02973(.A1(new_n3166_), .A2(new_n3121_), .Z(new_n3167_));
  XOR2_X1    g02974(.A1(new_n3167_), .A2(new_n3071_), .Z(new_n3168_));
  NAND2_X1   g02975(.A1(new_n3132_), .A2(new_n2961_), .ZN(new_n3169_));
  OAI21_X1   g02976(.A1(new_n2909_), .A2(new_n2918_), .B(new_n3169_), .ZN(new_n3170_));
  NAND2_X1   g02977(.A1(new_n2897_), .A2(new_n2982_), .ZN(new_n3171_));
  NAND2_X1   g02978(.A1(new_n2972_), .A2(new_n3095_), .ZN(new_n3172_));
  NAND2_X1   g02979(.A1(new_n3172_), .A2(new_n3171_), .ZN(new_n3173_));
  XOR2_X1    g02980(.A1(new_n3170_), .A2(new_n3173_), .Z(new_n3174_));
  XOR2_X1    g02981(.A1(new_n3174_), .A2(new_n3168_), .Z(new_n3175_));
  NAND2_X1   g02982(.A1(new_n3137_), .A2(new_n3140_), .ZN(new_n3176_));
  NAND2_X1   g02983(.A1(new_n3142_), .A2(new_n3176_), .ZN(new_n3177_));
  AOI22_X1   g02984(.A1(\a[13] ), .A2(\a[27] ), .B1(\a[14] ), .B2(\a[26] ), .ZN(new_n3178_));
  INV_X1     g02985(.I(new_n3178_), .ZN(new_n3179_));
  NOR2_X1    g02986(.A1(new_n767_), .A2(new_n1972_), .ZN(new_n3180_));
  NOR2_X1    g02987(.A1(new_n225_), .A2(new_n2752_), .ZN(new_n3181_));
  AOI21_X1   g02988(.A1(new_n3179_), .A2(new_n3181_), .B(new_n3180_), .ZN(new_n3182_));
  INV_X1     g02989(.I(new_n3182_), .ZN(new_n3183_));
  OAI21_X1   g02990(.A1(new_n3180_), .A2(new_n3178_), .B(new_n3181_), .ZN(new_n3184_));
  OAI21_X1   g02991(.A1(new_n3183_), .A2(new_n3178_), .B(new_n3184_), .ZN(new_n3185_));
  OAI22_X1   g02992(.A1(new_n893_), .A2(new_n1779_), .B1(new_n1443_), .B2(new_n982_), .ZN(new_n3186_));
  OAI21_X1   g02993(.A1(new_n1428_), .A2(new_n1529_), .B(new_n3186_), .ZN(new_n3187_));
  NAND3_X1   g02994(.A1(new_n3187_), .A2(\a[15] ), .A3(\a[25] ), .ZN(new_n3188_));
  AOI22_X1   g02995(.A1(\a[16] ), .A2(\a[24] ), .B1(\a[17] ), .B2(\a[23] ), .ZN(new_n3189_));
  NOR2_X1    g02996(.A1(new_n1428_), .A2(new_n1529_), .ZN(new_n3190_));
  NOR2_X1    g02997(.A1(new_n3186_), .A2(new_n3190_), .ZN(new_n3191_));
  INV_X1     g02998(.I(new_n3191_), .ZN(new_n3192_));
  OAI21_X1   g02999(.A1(new_n3189_), .A2(new_n3192_), .B(new_n3188_), .ZN(new_n3193_));
  XOR2_X1    g03000(.A1(new_n3193_), .A2(new_n3185_), .Z(new_n3194_));
  NOR4_X1    g03001(.A1(new_n367_), .A2(new_n417_), .A3(new_n2030_), .A4(new_n2442_), .ZN(new_n3195_));
  NAND4_X1   g03002(.A1(\a[6] ), .A2(\a[11] ), .A3(\a[29] ), .A4(\a[34] ), .ZN(new_n3196_));
  NAND2_X1   g03003(.A1(new_n747_), .A2(new_n2254_), .ZN(new_n3197_));
  AOI21_X1   g03004(.A1(new_n3197_), .A2(new_n3196_), .B(new_n3195_), .ZN(new_n3198_));
  NAND2_X1   g03005(.A1(\a[11] ), .A2(\a[29] ), .ZN(new_n3199_));
  OR2_X2     g03006(.A1(new_n3198_), .A2(new_n3195_), .Z(new_n3200_));
  AOI22_X1   g03007(.A1(\a[6] ), .A2(\a[34] ), .B1(\a[10] ), .B2(\a[30] ), .ZN(new_n3201_));
  OAI22_X1   g03008(.A1(new_n3200_), .A2(new_n3201_), .B1(new_n3198_), .B2(new_n3199_), .ZN(new_n3202_));
  XNOR2_X1   g03009(.A1(new_n3194_), .A2(new_n3202_), .ZN(new_n3203_));
  INV_X1     g03010(.I(new_n3203_), .ZN(new_n3204_));
  XOR2_X1    g03011(.A1(new_n3177_), .A2(new_n3204_), .Z(new_n3205_));
  XNOR2_X1   g03012(.A1(new_n3205_), .A2(new_n3175_), .ZN(new_n3206_));
  NAND2_X1   g03013(.A1(new_n3144_), .A2(new_n3131_), .ZN(new_n3207_));
  NAND2_X1   g03014(.A1(new_n3145_), .A2(new_n3112_), .ZN(new_n3208_));
  NAND2_X1   g03015(.A1(new_n3208_), .A2(new_n3207_), .ZN(new_n3209_));
  NOR2_X1    g03016(.A1(new_n2051_), .A2(new_n2200_), .ZN(new_n3210_));
  NAND2_X1   g03017(.A1(new_n467_), .A2(new_n3210_), .ZN(new_n3211_));
  OAI22_X1   g03018(.A1(new_n415_), .A2(new_n2637_), .B1(new_n2276_), .B2(new_n773_), .ZN(new_n3212_));
  NAND2_X1   g03019(.A1(new_n3212_), .A2(new_n3211_), .ZN(new_n3213_));
  NAND3_X1   g03020(.A1(new_n3213_), .A2(\a[7] ), .A3(\a[33] ), .ZN(new_n3214_));
  AOI22_X1   g03021(.A1(\a[8] ), .A2(\a[32] ), .B1(\a[9] ), .B2(\a[31] ), .ZN(new_n3215_));
  NAND2_X1   g03022(.A1(new_n3213_), .A2(new_n3211_), .ZN(new_n3216_));
  OAI21_X1   g03023(.A1(new_n3215_), .A2(new_n3216_), .B(new_n3214_), .ZN(new_n3217_));
  AOI22_X1   g03024(.A1(\a[0] ), .A2(\a[40] ), .B1(\a[2] ), .B2(\a[38] ), .ZN(new_n3218_));
  INV_X1     g03025(.I(new_n3218_), .ZN(new_n3219_));
  NOR2_X1    g03026(.A1(new_n884_), .A2(new_n1175_), .ZN(new_n3220_));
  INV_X1     g03027(.I(\a[40] ), .ZN(new_n3221_));
  NOR2_X1    g03028(.A1(new_n2914_), .A2(new_n3221_), .ZN(new_n3222_));
  INV_X1     g03029(.I(new_n3222_), .ZN(new_n3223_));
  NOR2_X1    g03030(.A1(new_n3223_), .A2(new_n412_), .ZN(new_n3224_));
  AOI21_X1   g03031(.A1(new_n3220_), .A2(new_n3219_), .B(new_n3224_), .ZN(new_n3225_));
  NAND2_X1   g03032(.A1(new_n3225_), .A2(new_n3219_), .ZN(new_n3226_));
  OAI21_X1   g03033(.A1(new_n3224_), .A2(new_n3218_), .B(new_n3220_), .ZN(new_n3227_));
  NAND2_X1   g03034(.A1(new_n3226_), .A2(new_n3227_), .ZN(new_n3228_));
  XNOR2_X1   g03035(.A1(new_n3217_), .A2(new_n3228_), .ZN(new_n3229_));
  NOR4_X1    g03036(.A1(new_n253_), .A2(new_n536_), .A3(new_n1718_), .A4(new_n2524_), .ZN(new_n3230_));
  NOR2_X1    g03037(.A1(new_n536_), .A2(new_n2626_), .ZN(new_n3231_));
  NOR2_X1    g03038(.A1(new_n2524_), .A2(new_n2626_), .ZN(new_n3232_));
  AOI22_X1   g03039(.A1(new_n2186_), .A2(new_n3231_), .B1(new_n3232_), .B2(new_n243_), .ZN(new_n3233_));
  NOR2_X1    g03040(.A1(new_n3233_), .A2(new_n3230_), .ZN(new_n3234_));
  NAND2_X1   g03041(.A1(\a[4] ), .A2(\a[36] ), .ZN(new_n3235_));
  INV_X1     g03042(.I(new_n3230_), .ZN(new_n3236_));
  NAND2_X1   g03043(.A1(new_n3233_), .A2(new_n3236_), .ZN(new_n3237_));
  AOI22_X1   g03044(.A1(\a[5] ), .A2(\a[35] ), .B1(\a[12] ), .B2(\a[28] ), .ZN(new_n3238_));
  OAI22_X1   g03045(.A1(new_n3234_), .A2(new_n3235_), .B1(new_n3237_), .B2(new_n3238_), .ZN(new_n3239_));
  XOR2_X1    g03046(.A1(new_n3229_), .A2(new_n3239_), .Z(new_n3240_));
  INV_X1     g03047(.I(new_n3240_), .ZN(new_n3241_));
  NAND2_X1   g03048(.A1(new_n3114_), .A2(new_n3125_), .ZN(new_n3242_));
  NAND2_X1   g03049(.A1(new_n3127_), .A2(new_n3242_), .ZN(new_n3243_));
  NOR3_X1    g03050(.A1(new_n1281_), .A2(new_n3118_), .A3(new_n2929_), .ZN(new_n3244_));
  NOR2_X1    g03051(.A1(new_n3119_), .A2(new_n3123_), .ZN(new_n3245_));
  NOR2_X1    g03052(.A1(new_n3245_), .A2(new_n3244_), .ZN(new_n3246_));
  XOR2_X1    g03053(.A1(new_n3032_), .A2(new_n3052_), .Z(new_n3247_));
  XNOR2_X1   g03054(.A1(new_n3247_), .A2(new_n3246_), .ZN(new_n3248_));
  NOR2_X1    g03055(.A1(new_n3243_), .A2(new_n3248_), .ZN(new_n3249_));
  NAND2_X1   g03056(.A1(new_n3243_), .A2(new_n3248_), .ZN(new_n3250_));
  INV_X1     g03057(.I(new_n3250_), .ZN(new_n3251_));
  NOR2_X1    g03058(.A1(new_n3251_), .A2(new_n3249_), .ZN(new_n3252_));
  NOR2_X1    g03059(.A1(new_n3252_), .A2(new_n3241_), .ZN(new_n3253_));
  NAND2_X1   g03060(.A1(new_n3252_), .A2(new_n3241_), .ZN(new_n3254_));
  INV_X1     g03061(.I(new_n3254_), .ZN(new_n3255_));
  NOR2_X1    g03062(.A1(new_n3255_), .A2(new_n3253_), .ZN(new_n3256_));
  XOR2_X1    g03063(.A1(new_n3209_), .A2(new_n3256_), .Z(new_n3257_));
  INV_X1     g03064(.I(new_n3257_), .ZN(new_n3258_));
  NAND2_X1   g03065(.A1(new_n3258_), .A2(new_n3206_), .ZN(new_n3259_));
  OR2_X2     g03066(.A1(new_n3258_), .A2(new_n3206_), .Z(new_n3260_));
  AND2_X2    g03067(.A1(new_n3260_), .A2(new_n3259_), .Z(new_n3261_));
  INV_X1     g03068(.I(new_n3261_), .ZN(new_n3262_));
  INV_X1     g03069(.I(new_n3059_), .ZN(new_n3263_));
  NOR2_X1    g03070(.A1(new_n3263_), .A2(new_n3023_), .ZN(new_n3264_));
  NOR2_X1    g03071(.A1(new_n3264_), .A2(new_n3058_), .ZN(new_n3265_));
  XOR2_X1    g03072(.A1(new_n3042_), .A2(new_n3088_), .Z(new_n3266_));
  XOR2_X1    g03073(.A1(new_n3266_), .A2(new_n3079_), .Z(new_n3267_));
  NAND2_X1   g03074(.A1(new_n3044_), .A2(new_n3033_), .ZN(new_n3268_));
  INV_X1     g03075(.I(new_n3045_), .ZN(new_n3269_));
  NAND2_X1   g03076(.A1(new_n3269_), .A2(new_n3053_), .ZN(new_n3270_));
  NAND2_X1   g03077(.A1(new_n3270_), .A2(new_n3268_), .ZN(new_n3271_));
  NAND2_X1   g03078(.A1(new_n3073_), .A2(new_n3081_), .ZN(new_n3272_));
  INV_X1     g03079(.I(new_n3082_), .ZN(new_n3273_));
  NAND2_X1   g03080(.A1(new_n3273_), .A2(new_n3090_), .ZN(new_n3274_));
  NAND2_X1   g03081(.A1(new_n3274_), .A2(new_n3272_), .ZN(new_n3275_));
  XOR2_X1    g03082(.A1(new_n3271_), .A2(new_n3275_), .Z(new_n3276_));
  XOR2_X1    g03083(.A1(new_n3276_), .A2(new_n3267_), .Z(new_n3277_));
  NOR2_X1    g03084(.A1(new_n3102_), .A2(new_n3099_), .ZN(new_n3278_));
  XOR2_X1    g03085(.A1(new_n3278_), .A2(new_n3277_), .Z(new_n3279_));
  NAND2_X1   g03086(.A1(new_n3265_), .A2(new_n3279_), .ZN(new_n3280_));
  NOR2_X1    g03087(.A1(new_n3265_), .A2(new_n3279_), .ZN(new_n3281_));
  INV_X1     g03088(.I(new_n3281_), .ZN(new_n3282_));
  AND2_X2    g03089(.A1(new_n3282_), .A2(new_n3280_), .Z(new_n3283_));
  INV_X1     g03090(.I(new_n3283_), .ZN(new_n3284_));
  NAND2_X1   g03091(.A1(new_n3064_), .A2(new_n3104_), .ZN(new_n3285_));
  OAI21_X1   g03092(.A1(new_n3105_), .A2(new_n3061_), .B(new_n3285_), .ZN(new_n3286_));
  NOR2_X1    g03093(.A1(new_n3284_), .A2(new_n3286_), .ZN(new_n3287_));
  INV_X1     g03094(.I(new_n3286_), .ZN(new_n3288_));
  NOR2_X1    g03095(.A1(new_n3283_), .A2(new_n3288_), .ZN(new_n3289_));
  NOR2_X1    g03096(.A1(new_n3287_), .A2(new_n3289_), .ZN(new_n3290_));
  NOR2_X1    g03097(.A1(new_n3262_), .A2(new_n3290_), .ZN(new_n3291_));
  NOR3_X1    g03098(.A1(new_n3261_), .A2(new_n3287_), .A3(new_n3289_), .ZN(new_n3292_));
  NOR2_X1    g03099(.A1(new_n3291_), .A2(new_n3292_), .ZN(new_n3293_));
  INV_X1     g03100(.I(new_n3293_), .ZN(new_n3294_));
  NOR2_X1    g03101(.A1(new_n3153_), .A2(new_n3149_), .ZN(new_n3295_));
  NOR2_X1    g03102(.A1(new_n3294_), .A2(new_n3295_), .ZN(new_n3296_));
  INV_X1     g03103(.I(new_n3296_), .ZN(new_n3297_));
  NAND2_X1   g03104(.A1(new_n3294_), .A2(new_n3295_), .ZN(new_n3298_));
  NAND2_X1   g03105(.A1(new_n3297_), .A2(new_n3298_), .ZN(new_n3299_));
  INV_X1     g03106(.I(new_n2881_), .ZN(new_n3300_));
  INV_X1     g03107(.I(new_n2737_), .ZN(new_n3301_));
  INV_X1     g03108(.I(new_n2614_), .ZN(new_n3302_));
  OAI21_X1   g03109(.A1(new_n2490_), .A2(new_n2465_), .B(new_n2615_), .ZN(new_n3303_));
  AOI21_X1   g03110(.A1(new_n3303_), .A2(new_n3302_), .B(new_n2735_), .ZN(new_n3304_));
  OAI21_X1   g03111(.A1(new_n3304_), .A2(new_n3301_), .B(new_n2882_), .ZN(new_n3305_));
  INV_X1     g03112(.I(new_n3016_), .ZN(new_n3306_));
  AOI21_X1   g03113(.A1(new_n3305_), .A2(new_n3300_), .B(new_n3306_), .ZN(new_n3307_));
  INV_X1     g03114(.I(new_n3155_), .ZN(new_n3308_));
  OAI21_X1   g03115(.A1(new_n3307_), .A2(new_n3014_), .B(new_n3308_), .ZN(new_n3309_));
  INV_X1     g03116(.I(new_n3298_), .ZN(new_n3310_));
  AOI21_X1   g03117(.A1(new_n3309_), .A2(new_n3156_), .B(new_n3310_), .ZN(new_n3311_));
  AOI22_X1   g03118(.A1(new_n3311_), .A2(new_n3297_), .B1(new_n3161_), .B2(new_n3299_), .ZN(\asquared[41] ));
  OAI21_X1   g03119(.A1(new_n3160_), .A2(new_n3157_), .B(new_n3298_), .ZN(new_n3313_));
  NAND2_X1   g03120(.A1(new_n3313_), .A2(new_n3297_), .ZN(new_n3314_));
  AOI21_X1   g03121(.A1(new_n3283_), .A2(new_n3286_), .B(new_n3291_), .ZN(new_n3315_));
  NAND2_X1   g03122(.A1(new_n3193_), .A2(new_n3185_), .ZN(new_n3316_));
  NAND2_X1   g03123(.A1(new_n3194_), .A2(new_n3202_), .ZN(new_n3317_));
  NAND2_X1   g03124(.A1(new_n3317_), .A2(new_n3316_), .ZN(new_n3318_));
  NAND2_X1   g03125(.A1(new_n3032_), .A2(new_n3052_), .ZN(new_n3319_));
  INV_X1     g03126(.I(new_n3247_), .ZN(new_n3320_));
  OAI21_X1   g03127(.A1(new_n3320_), .A2(new_n3246_), .B(new_n3319_), .ZN(new_n3321_));
  NAND2_X1   g03128(.A1(new_n3042_), .A2(new_n3088_), .ZN(new_n3322_));
  NAND2_X1   g03129(.A1(new_n3266_), .A2(new_n3079_), .ZN(new_n3323_));
  NAND2_X1   g03130(.A1(new_n3323_), .A2(new_n3322_), .ZN(new_n3324_));
  XOR2_X1    g03131(.A1(new_n3321_), .A2(new_n3324_), .Z(new_n3325_));
  XOR2_X1    g03132(.A1(new_n3325_), .A2(new_n3318_), .Z(new_n3326_));
  INV_X1     g03133(.I(\a[41] ), .ZN(new_n3327_));
  NOR2_X1    g03134(.A1(new_n3116_), .A2(new_n3327_), .ZN(new_n3328_));
  INV_X1     g03135(.I(new_n3328_), .ZN(new_n3329_));
  NOR2_X1    g03136(.A1(new_n3329_), .A2(new_n412_), .ZN(new_n3330_));
  AOI22_X1   g03137(.A1(\a[0] ), .A2(\a[41] ), .B1(\a[2] ), .B2(\a[39] ), .ZN(new_n3331_));
  NOR2_X1    g03138(.A1(new_n3330_), .A2(new_n3331_), .ZN(new_n3332_));
  INV_X1     g03139(.I(new_n3332_), .ZN(new_n3333_));
  NOR2_X1    g03140(.A1(new_n3333_), .A2(new_n3164_), .ZN(new_n3334_));
  NOR2_X1    g03141(.A1(new_n3332_), .A2(new_n3163_), .ZN(new_n3335_));
  NOR2_X1    g03142(.A1(new_n3334_), .A2(new_n3335_), .ZN(new_n3336_));
  XOR2_X1    g03143(.A1(new_n3336_), .A2(new_n3237_), .Z(new_n3337_));
  AOI22_X1   g03144(.A1(\a[13] ), .A2(\a[28] ), .B1(\a[15] ), .B2(\a[26] ), .ZN(new_n3338_));
  NOR2_X1    g03145(.A1(new_n225_), .A2(new_n2914_), .ZN(new_n3339_));
  INV_X1     g03146(.I(new_n3339_), .ZN(new_n3340_));
  INV_X1     g03147(.I(new_n2412_), .ZN(new_n3341_));
  NOR2_X1    g03148(.A1(new_n3341_), .A2(new_n836_), .ZN(new_n3342_));
  NOR3_X1    g03149(.A1(new_n3342_), .A2(new_n3338_), .A3(new_n3340_), .ZN(new_n3343_));
  NOR2_X1    g03150(.A1(new_n3343_), .A2(new_n3342_), .ZN(new_n3344_));
  INV_X1     g03151(.I(new_n3344_), .ZN(new_n3345_));
  OAI22_X1   g03152(.A1(new_n3345_), .A2(new_n3338_), .B1(new_n3340_), .B2(new_n3343_), .ZN(new_n3346_));
  XOR2_X1    g03153(.A1(new_n3337_), .A2(new_n3346_), .Z(new_n3347_));
  NAND2_X1   g03154(.A1(new_n3271_), .A2(new_n3275_), .ZN(new_n3348_));
  NAND2_X1   g03155(.A1(new_n3276_), .A2(new_n3267_), .ZN(new_n3349_));
  NAND2_X1   g03156(.A1(new_n3349_), .A2(new_n3348_), .ZN(new_n3350_));
  XOR2_X1    g03157(.A1(new_n3350_), .A2(new_n3347_), .Z(new_n3351_));
  XOR2_X1    g03158(.A1(new_n3351_), .A2(new_n3326_), .Z(new_n3352_));
  INV_X1     g03159(.I(new_n3352_), .ZN(new_n3353_));
  INV_X1     g03160(.I(new_n3277_), .ZN(new_n3354_));
  NOR2_X1    g03161(.A1(new_n3278_), .A2(new_n3354_), .ZN(new_n3355_));
  NOR2_X1    g03162(.A1(new_n3281_), .A2(new_n3355_), .ZN(new_n3356_));
  NOR2_X1    g03163(.A1(new_n1816_), .A2(new_n623_), .ZN(new_n3357_));
  NOR3_X1    g03164(.A1(new_n892_), .A2(new_n1750_), .A3(new_n2752_), .ZN(new_n3358_));
  NAND4_X1   g03165(.A1(\a[4] ), .A2(\a[12] ), .A3(\a[29] ), .A4(\a[37] ), .ZN(new_n3359_));
  OAI21_X1   g03166(.A1(new_n3357_), .A2(new_n3358_), .B(new_n3359_), .ZN(new_n3360_));
  NAND3_X1   g03167(.A1(new_n3360_), .A2(\a[14] ), .A3(\a[27] ), .ZN(new_n3361_));
  AOI22_X1   g03168(.A1(\a[4] ), .A2(\a[37] ), .B1(\a[12] ), .B2(\a[29] ), .ZN(new_n3362_));
  NAND2_X1   g03169(.A1(new_n3360_), .A2(new_n3359_), .ZN(new_n3363_));
  OAI21_X1   g03170(.A1(new_n3362_), .A2(new_n3363_), .B(new_n3361_), .ZN(new_n3364_));
  OAI22_X1   g03171(.A1(new_n1428_), .A2(new_n1779_), .B1(new_n1429_), .B2(new_n1443_), .ZN(new_n3365_));
  OAI21_X1   g03172(.A1(new_n1275_), .A2(new_n1529_), .B(new_n3365_), .ZN(new_n3366_));
  NAND3_X1   g03173(.A1(new_n3366_), .A2(\a[16] ), .A3(\a[25] ), .ZN(new_n3367_));
  AOI22_X1   g03174(.A1(\a[17] ), .A2(\a[24] ), .B1(\a[18] ), .B2(\a[23] ), .ZN(new_n3368_));
  NOR2_X1    g03175(.A1(new_n1275_), .A2(new_n1529_), .ZN(new_n3369_));
  NOR2_X1    g03176(.A1(new_n3365_), .A2(new_n3369_), .ZN(new_n3370_));
  INV_X1     g03177(.I(new_n3370_), .ZN(new_n3371_));
  OAI21_X1   g03178(.A1(new_n3368_), .A2(new_n3371_), .B(new_n3367_), .ZN(new_n3372_));
  XOR2_X1    g03179(.A1(new_n3372_), .A2(new_n3364_), .Z(new_n3373_));
  NOR2_X1    g03180(.A1(new_n2200_), .A2(new_n2442_), .ZN(new_n3374_));
  INV_X1     g03181(.I(new_n3374_), .ZN(new_n3375_));
  NOR2_X1    g03182(.A1(new_n3375_), .A2(new_n773_), .ZN(new_n3376_));
  NAND3_X1   g03183(.A1(new_n2055_), .A2(\a[7] ), .A3(\a[34] ), .ZN(new_n3377_));
  NAND2_X1   g03184(.A1(new_n3210_), .A2(new_n540_), .ZN(new_n3378_));
  AOI21_X1   g03185(.A1(new_n3377_), .A2(new_n3378_), .B(new_n3376_), .ZN(new_n3379_));
  AOI22_X1   g03186(.A1(\a[7] ), .A2(\a[34] ), .B1(\a[9] ), .B2(\a[32] ), .ZN(new_n3380_));
  NOR2_X1    g03187(.A1(new_n3379_), .A2(new_n3376_), .ZN(new_n3381_));
  INV_X1     g03188(.I(new_n3381_), .ZN(new_n3382_));
  OAI22_X1   g03189(.A1(new_n3382_), .A2(new_n3380_), .B1(new_n2660_), .B2(new_n3379_), .ZN(new_n3383_));
  XNOR2_X1   g03190(.A1(new_n3373_), .A2(new_n3383_), .ZN(new_n3384_));
  INV_X1     g03191(.I(new_n3384_), .ZN(new_n3385_));
  NAND2_X1   g03192(.A1(new_n3170_), .A2(new_n3173_), .ZN(new_n3386_));
  NAND2_X1   g03193(.A1(new_n3174_), .A2(new_n3168_), .ZN(new_n3387_));
  NAND2_X1   g03194(.A1(new_n3387_), .A2(new_n3386_), .ZN(new_n3388_));
  NAND2_X1   g03195(.A1(new_n3167_), .A2(new_n3071_), .ZN(new_n3389_));
  OAI21_X1   g03196(.A1(new_n3121_), .A2(new_n3166_), .B(new_n3389_), .ZN(new_n3390_));
  NOR2_X1    g03197(.A1(new_n979_), .A2(new_n1175_), .ZN(new_n3391_));
  NOR2_X1    g03198(.A1(new_n1381_), .A2(new_n3391_), .ZN(new_n3392_));
  NOR2_X1    g03199(.A1(new_n355_), .A2(new_n2274_), .ZN(new_n3393_));
  INV_X1     g03200(.I(new_n3391_), .ZN(new_n3394_));
  NOR2_X1    g03201(.A1(new_n1382_), .A2(new_n3394_), .ZN(new_n3395_));
  OAI21_X1   g03202(.A1(new_n3395_), .A2(new_n3392_), .B(new_n3393_), .ZN(new_n3396_));
  INV_X1     g03203(.I(new_n3392_), .ZN(new_n3397_));
  AOI21_X1   g03204(.A1(new_n3393_), .A2(new_n3397_), .B(new_n3395_), .ZN(new_n3398_));
  INV_X1     g03205(.I(new_n3398_), .ZN(new_n3399_));
  OAI21_X1   g03206(.A1(new_n3399_), .A2(new_n3392_), .B(new_n3396_), .ZN(new_n3400_));
  NOR2_X1    g03207(.A1(new_n2030_), .A2(new_n2524_), .ZN(new_n3401_));
  INV_X1     g03208(.I(new_n3401_), .ZN(new_n3402_));
  NOR2_X1    g03209(.A1(new_n840_), .A2(new_n3402_), .ZN(new_n3403_));
  NOR3_X1    g03210(.A1(new_n515_), .A2(new_n2030_), .A3(new_n2626_), .ZN(new_n3404_));
  INV_X1     g03211(.I(new_n3232_), .ZN(new_n3405_));
  NOR2_X1    g03212(.A1(new_n3405_), .A2(new_n371_), .ZN(new_n3406_));
  NOR2_X1    g03213(.A1(new_n3406_), .A2(new_n3404_), .ZN(new_n3407_));
  NOR2_X1    g03214(.A1(new_n3407_), .A2(new_n3403_), .ZN(new_n3408_));
  NAND2_X1   g03215(.A1(\a[5] ), .A2(\a[36] ), .ZN(new_n3409_));
  AOI22_X1   g03216(.A1(\a[6] ), .A2(\a[35] ), .B1(\a[11] ), .B2(\a[30] ), .ZN(new_n3410_));
  NOR2_X1    g03217(.A1(new_n3408_), .A2(new_n3403_), .ZN(new_n3411_));
  INV_X1     g03218(.I(new_n3411_), .ZN(new_n3412_));
  OAI22_X1   g03219(.A1(new_n3412_), .A2(new_n3410_), .B1(new_n3408_), .B2(new_n3409_), .ZN(new_n3413_));
  XNOR2_X1   g03220(.A1(new_n3413_), .A2(new_n3400_), .ZN(new_n3414_));
  XNOR2_X1   g03221(.A1(new_n3414_), .A2(new_n3390_), .ZN(new_n3415_));
  XOR2_X1    g03222(.A1(new_n3388_), .A2(new_n3415_), .Z(new_n3416_));
  OR2_X2     g03223(.A1(new_n3416_), .A2(new_n3385_), .Z(new_n3417_));
  NAND2_X1   g03224(.A1(new_n3416_), .A2(new_n3385_), .ZN(new_n3418_));
  AND2_X2    g03225(.A1(new_n3417_), .A2(new_n3418_), .Z(new_n3419_));
  NOR2_X1    g03226(.A1(new_n3356_), .A2(new_n3419_), .ZN(new_n3420_));
  INV_X1     g03227(.I(new_n3419_), .ZN(new_n3421_));
  NOR2_X1    g03228(.A1(new_n3356_), .A2(new_n3421_), .ZN(new_n3422_));
  NOR2_X1    g03229(.A1(new_n3422_), .A2(new_n3421_), .ZN(new_n3423_));
  NOR2_X1    g03230(.A1(new_n3423_), .A2(new_n3420_), .ZN(new_n3424_));
  NOR2_X1    g03231(.A1(new_n3424_), .A2(new_n3353_), .ZN(new_n3425_));
  NOR3_X1    g03232(.A1(new_n3423_), .A2(new_n3352_), .A3(new_n3420_), .ZN(new_n3426_));
  NOR2_X1    g03233(.A1(new_n3425_), .A2(new_n3426_), .ZN(new_n3427_));
  NAND2_X1   g03234(.A1(new_n3209_), .A2(new_n3256_), .ZN(new_n3428_));
  NAND2_X1   g03235(.A1(new_n3260_), .A2(new_n3428_), .ZN(new_n3429_));
  NAND2_X1   g03236(.A1(new_n3177_), .A2(new_n3204_), .ZN(new_n3430_));
  NAND2_X1   g03237(.A1(new_n3205_), .A2(new_n3175_), .ZN(new_n3431_));
  NAND2_X1   g03238(.A1(new_n3431_), .A2(new_n3430_), .ZN(new_n3432_));
  NOR2_X1    g03239(.A1(new_n3255_), .A2(new_n3251_), .ZN(new_n3433_));
  NOR2_X1    g03240(.A1(new_n194_), .A2(new_n3221_), .ZN(new_n3434_));
  NAND2_X1   g03241(.A1(new_n1221_), .A2(\a[40] ), .ZN(new_n3435_));
  OAI21_X1   g03242(.A1(\a[21] ), .A2(new_n3434_), .B(new_n3435_), .ZN(new_n3436_));
  INV_X1     g03243(.I(new_n3436_), .ZN(new_n3437_));
  XOR2_X1    g03244(.A1(new_n3216_), .A2(new_n3437_), .Z(new_n3438_));
  XOR2_X1    g03245(.A1(new_n3438_), .A2(new_n3200_), .Z(new_n3439_));
  NAND2_X1   g03246(.A1(new_n3217_), .A2(new_n3228_), .ZN(new_n3440_));
  INV_X1     g03247(.I(new_n3229_), .ZN(new_n3441_));
  NAND2_X1   g03248(.A1(new_n3441_), .A2(new_n3239_), .ZN(new_n3442_));
  NAND2_X1   g03249(.A1(new_n3442_), .A2(new_n3440_), .ZN(new_n3443_));
  XOR2_X1    g03250(.A1(new_n3191_), .A2(new_n3225_), .Z(new_n3444_));
  NOR2_X1    g03251(.A1(new_n3444_), .A2(new_n3183_), .ZN(new_n3445_));
  INV_X1     g03252(.I(new_n3444_), .ZN(new_n3446_));
  NOR2_X1    g03253(.A1(new_n3446_), .A2(new_n3182_), .ZN(new_n3447_));
  NOR2_X1    g03254(.A1(new_n3447_), .A2(new_n3445_), .ZN(new_n3448_));
  XOR2_X1    g03255(.A1(new_n3443_), .A2(new_n3448_), .Z(new_n3449_));
  OR2_X2     g03256(.A1(new_n3449_), .A2(new_n3439_), .Z(new_n3450_));
  NAND2_X1   g03257(.A1(new_n3449_), .A2(new_n3439_), .ZN(new_n3451_));
  AND2_X2    g03258(.A1(new_n3450_), .A2(new_n3451_), .Z(new_n3452_));
  XOR2_X1    g03259(.A1(new_n3433_), .A2(new_n3452_), .Z(new_n3453_));
  XNOR2_X1   g03260(.A1(new_n3453_), .A2(new_n3432_), .ZN(new_n3454_));
  NOR2_X1    g03261(.A1(new_n3429_), .A2(new_n3454_), .ZN(new_n3455_));
  NAND2_X1   g03262(.A1(new_n3429_), .A2(new_n3454_), .ZN(new_n3456_));
  INV_X1     g03263(.I(new_n3456_), .ZN(new_n3457_));
  NOR2_X1    g03264(.A1(new_n3457_), .A2(new_n3455_), .ZN(new_n3458_));
  NAND2_X1   g03265(.A1(new_n3458_), .A2(new_n3427_), .ZN(new_n3459_));
  INV_X1     g03266(.I(new_n3459_), .ZN(new_n3460_));
  NOR2_X1    g03267(.A1(new_n3458_), .A2(new_n3427_), .ZN(new_n3461_));
  NOR2_X1    g03268(.A1(new_n3460_), .A2(new_n3461_), .ZN(new_n3462_));
  INV_X1     g03269(.I(new_n3462_), .ZN(new_n3463_));
  NOR2_X1    g03270(.A1(new_n3463_), .A2(new_n3315_), .ZN(new_n3464_));
  NAND2_X1   g03271(.A1(new_n3463_), .A2(new_n3315_), .ZN(new_n3465_));
  INV_X1     g03272(.I(new_n3465_), .ZN(new_n3466_));
  NOR2_X1    g03273(.A1(new_n3466_), .A2(new_n3464_), .ZN(new_n3467_));
  XOR2_X1    g03274(.A1(new_n3314_), .A2(new_n3467_), .Z(\asquared[42] ));
  AOI21_X1   g03275(.A1(new_n3313_), .A2(new_n3297_), .B(new_n3466_), .ZN(new_n3469_));
  NOR2_X1    g03276(.A1(new_n3469_), .A2(new_n3464_), .ZN(new_n3470_));
  NOR2_X1    g03277(.A1(new_n3460_), .A2(new_n3457_), .ZN(new_n3471_));
  INV_X1     g03278(.I(new_n3471_), .ZN(new_n3472_));
  NOR2_X1    g03279(.A1(new_n3425_), .A2(new_n3422_), .ZN(new_n3473_));
  NAND2_X1   g03280(.A1(new_n3350_), .A2(new_n3347_), .ZN(new_n3474_));
  NAND2_X1   g03281(.A1(new_n3351_), .A2(new_n3326_), .ZN(new_n3475_));
  NAND2_X1   g03282(.A1(new_n3475_), .A2(new_n3474_), .ZN(new_n3476_));
  NAND2_X1   g03283(.A1(new_n3388_), .A2(new_n3415_), .ZN(new_n3477_));
  NAND2_X1   g03284(.A1(new_n3418_), .A2(new_n3477_), .ZN(new_n3478_));
  NAND2_X1   g03285(.A1(new_n3372_), .A2(new_n3364_), .ZN(new_n3479_));
  NAND2_X1   g03286(.A1(new_n3373_), .A2(new_n3383_), .ZN(new_n3480_));
  NAND2_X1   g03287(.A1(new_n3480_), .A2(new_n3479_), .ZN(new_n3481_));
  NOR2_X1    g03288(.A1(new_n3191_), .A2(new_n3225_), .ZN(new_n3482_));
  NOR2_X1    g03289(.A1(new_n3447_), .A2(new_n3482_), .ZN(new_n3483_));
  NAND2_X1   g03290(.A1(new_n3336_), .A2(new_n3237_), .ZN(new_n3484_));
  NAND2_X1   g03291(.A1(new_n3337_), .A2(new_n3346_), .ZN(new_n3485_));
  NAND2_X1   g03292(.A1(new_n3485_), .A2(new_n3484_), .ZN(new_n3486_));
  XNOR2_X1   g03293(.A1(new_n3486_), .A2(new_n3483_), .ZN(new_n3487_));
  XOR2_X1    g03294(.A1(new_n3487_), .A2(new_n3481_), .Z(new_n3488_));
  XOR2_X1    g03295(.A1(new_n3478_), .A2(new_n3488_), .Z(new_n3489_));
  XOR2_X1    g03296(.A1(new_n3476_), .A2(new_n3489_), .Z(new_n3490_));
  INV_X1     g03297(.I(new_n3490_), .ZN(new_n3491_));
  NAND2_X1   g03298(.A1(new_n3473_), .A2(new_n3491_), .ZN(new_n3492_));
  NOR2_X1    g03299(.A1(new_n3473_), .A2(new_n3491_), .ZN(new_n3493_));
  INV_X1     g03300(.I(new_n3493_), .ZN(new_n3494_));
  AND2_X2    g03301(.A1(new_n3494_), .A2(new_n3492_), .Z(new_n3495_));
  NOR2_X1    g03302(.A1(new_n3334_), .A2(new_n3330_), .ZN(new_n3496_));
  NOR2_X1    g03303(.A1(new_n3345_), .A2(new_n3371_), .ZN(new_n3497_));
  NOR2_X1    g03304(.A1(new_n3344_), .A2(new_n3370_), .ZN(new_n3498_));
  NOR2_X1    g03305(.A1(new_n3497_), .A2(new_n3498_), .ZN(new_n3499_));
  XNOR2_X1   g03306(.A1(new_n3499_), .A2(new_n3496_), .ZN(new_n3500_));
  XNOR2_X1   g03307(.A1(new_n3363_), .A2(new_n3398_), .ZN(new_n3501_));
  XOR2_X1    g03308(.A1(new_n3501_), .A2(new_n3412_), .Z(new_n3502_));
  NAND2_X1   g03309(.A1(new_n3413_), .A2(new_n3400_), .ZN(new_n3503_));
  INV_X1     g03310(.I(new_n3414_), .ZN(new_n3504_));
  NAND2_X1   g03311(.A1(new_n3504_), .A2(new_n3390_), .ZN(new_n3505_));
  NAND2_X1   g03312(.A1(new_n3505_), .A2(new_n3503_), .ZN(new_n3506_));
  XOR2_X1    g03313(.A1(new_n3506_), .A2(new_n3502_), .Z(new_n3507_));
  XNOR2_X1   g03314(.A1(new_n3507_), .A2(new_n3500_), .ZN(new_n3508_));
  NAND2_X1   g03315(.A1(new_n3443_), .A2(new_n3448_), .ZN(new_n3509_));
  NAND2_X1   g03316(.A1(new_n3216_), .A2(new_n3437_), .ZN(new_n3510_));
  NAND2_X1   g03317(.A1(new_n3438_), .A2(new_n3200_), .ZN(new_n3511_));
  NAND2_X1   g03318(.A1(new_n3511_), .A2(new_n3510_), .ZN(new_n3512_));
  NAND2_X1   g03319(.A1(\a[0] ), .A2(\a[42] ), .ZN(new_n3513_));
  XOR2_X1    g03320(.A1(new_n3435_), .A2(new_n3513_), .Z(new_n3514_));
  NAND2_X1   g03321(.A1(\a[1] ), .A2(\a[41] ), .ZN(new_n3515_));
  XNOR2_X1   g03322(.A1(new_n1552_), .A2(new_n3515_), .ZN(new_n3516_));
  XOR2_X1    g03323(.A1(new_n3514_), .A2(new_n3516_), .Z(new_n3517_));
  NAND3_X1   g03324(.A1(new_n3035_), .A2(\a[5] ), .A3(\a[29] ), .ZN(new_n3518_));
  NAND2_X1   g03325(.A1(new_n763_), .A2(new_n2254_), .ZN(new_n3519_));
  NOR4_X1    g03326(.A1(new_n253_), .A2(new_n536_), .A3(new_n2030_), .A4(new_n2752_), .ZN(new_n3520_));
  AOI21_X1   g03327(.A1(new_n3519_), .A2(new_n3518_), .B(new_n3520_), .ZN(new_n3521_));
  NAND2_X1   g03328(.A1(\a[13] ), .A2(\a[29] ), .ZN(new_n3522_));
  AOI22_X1   g03329(.A1(\a[5] ), .A2(\a[37] ), .B1(\a[12] ), .B2(\a[30] ), .ZN(new_n3523_));
  OR2_X2     g03330(.A1(new_n3521_), .A2(new_n3520_), .Z(new_n3524_));
  OAI22_X1   g03331(.A1(new_n3524_), .A2(new_n3523_), .B1(new_n3521_), .B2(new_n3522_), .ZN(new_n3525_));
  XOR2_X1    g03332(.A1(new_n3517_), .A2(new_n3525_), .Z(new_n3526_));
  XOR2_X1    g03333(.A1(new_n3512_), .A2(new_n3526_), .Z(new_n3527_));
  INV_X1     g03334(.I(new_n3527_), .ZN(new_n3528_));
  AND3_X2    g03335(.A1(new_n3451_), .A2(new_n3509_), .A3(new_n3528_), .Z(new_n3529_));
  AOI21_X1   g03336(.A1(new_n3451_), .A2(new_n3509_), .B(new_n3528_), .ZN(new_n3530_));
  NOR2_X1    g03337(.A1(new_n3529_), .A2(new_n3530_), .ZN(new_n3531_));
  XNOR2_X1   g03338(.A1(new_n3531_), .A2(new_n3508_), .ZN(new_n3532_));
  INV_X1     g03339(.I(new_n3432_), .ZN(new_n3533_));
  OAI21_X1   g03340(.A1(new_n3255_), .A2(new_n3251_), .B(new_n3452_), .ZN(new_n3534_));
  OAI21_X1   g03341(.A1(new_n3533_), .A2(new_n3453_), .B(new_n3534_), .ZN(new_n3535_));
  NOR2_X1    g03342(.A1(new_n1529_), .A2(new_n1092_), .ZN(new_n3536_));
  NOR2_X1    g03343(.A1(new_n1275_), .A2(new_n1779_), .ZN(new_n3537_));
  NOR2_X1    g03344(.A1(new_n1443_), .A2(new_n2851_), .ZN(new_n3538_));
  NOR2_X1    g03345(.A1(new_n3537_), .A2(new_n3538_), .ZN(new_n3539_));
  NOR2_X1    g03346(.A1(new_n3539_), .A2(new_n3536_), .ZN(new_n3540_));
  NAND2_X1   g03347(.A1(\a[17] ), .A2(\a[25] ), .ZN(new_n3541_));
  AOI22_X1   g03348(.A1(\a[18] ), .A2(\a[24] ), .B1(\a[19] ), .B2(\a[23] ), .ZN(new_n3542_));
  NOR2_X1    g03349(.A1(new_n3540_), .A2(new_n3536_), .ZN(new_n3543_));
  INV_X1     g03350(.I(new_n3543_), .ZN(new_n3544_));
  OAI22_X1   g03351(.A1(new_n3544_), .A2(new_n3542_), .B1(new_n3540_), .B2(new_n3541_), .ZN(new_n3545_));
  NAND4_X1   g03352(.A1(\a[3] ), .A2(\a[16] ), .A3(\a[26] ), .A4(\a[39] ), .ZN(new_n3546_));
  INV_X1     g03353(.I(new_n1710_), .ZN(new_n3547_));
  NOR2_X1    g03354(.A1(new_n742_), .A2(new_n3221_), .ZN(new_n3548_));
  INV_X1     g03355(.I(new_n3548_), .ZN(new_n3549_));
  NOR2_X1    g03356(.A1(new_n3116_), .A2(new_n3221_), .ZN(new_n3550_));
  INV_X1     g03357(.I(new_n3550_), .ZN(new_n3551_));
  OAI22_X1   g03358(.A1(new_n3547_), .A2(new_n3549_), .B1(new_n3551_), .B2(new_n246_), .ZN(new_n3552_));
  NAND2_X1   g03359(.A1(new_n3552_), .A2(new_n3546_), .ZN(new_n3553_));
  NAND3_X1   g03360(.A1(new_n3553_), .A2(\a[2] ), .A3(\a[40] ), .ZN(new_n3554_));
  NAND2_X1   g03361(.A1(new_n3553_), .A2(new_n3546_), .ZN(new_n3555_));
  AOI22_X1   g03362(.A1(\a[3] ), .A2(\a[39] ), .B1(\a[16] ), .B2(\a[26] ), .ZN(new_n3556_));
  OAI21_X1   g03363(.A1(new_n3555_), .A2(new_n3556_), .B(new_n3554_), .ZN(new_n3557_));
  XOR2_X1    g03364(.A1(new_n3545_), .A2(new_n3557_), .Z(new_n3558_));
  INV_X1     g03365(.I(new_n2186_), .ZN(new_n3559_));
  NOR2_X1    g03366(.A1(new_n759_), .A2(new_n2914_), .ZN(new_n3560_));
  INV_X1     g03367(.I(new_n3560_), .ZN(new_n3561_));
  NOR2_X1    g03368(.A1(new_n3559_), .A2(new_n3561_), .ZN(new_n3562_));
  NOR2_X1    g03369(.A1(new_n717_), .A2(new_n2914_), .ZN(new_n3563_));
  NAND3_X1   g03370(.A1(new_n3563_), .A2(\a[4] ), .A3(\a[27] ), .ZN(new_n3564_));
  NAND2_X1   g03371(.A1(new_n897_), .A2(new_n2103_), .ZN(new_n3565_));
  AOI21_X1   g03372(.A1(new_n3565_), .A2(new_n3564_), .B(new_n3562_), .ZN(new_n3566_));
  NAND2_X1   g03373(.A1(\a[15] ), .A2(\a[27] ), .ZN(new_n3567_));
  NOR2_X1    g03374(.A1(new_n3566_), .A2(new_n3562_), .ZN(new_n3568_));
  INV_X1     g03375(.I(new_n3568_), .ZN(new_n3569_));
  AOI22_X1   g03376(.A1(\a[4] ), .A2(\a[38] ), .B1(\a[14] ), .B2(\a[28] ), .ZN(new_n3570_));
  OAI22_X1   g03377(.A1(new_n3569_), .A2(new_n3570_), .B1(new_n3566_), .B2(new_n3567_), .ZN(new_n3571_));
  XNOR2_X1   g03378(.A1(new_n3558_), .A2(new_n3571_), .ZN(new_n3572_));
  INV_X1     g03379(.I(new_n3572_), .ZN(new_n3573_));
  NAND2_X1   g03380(.A1(new_n3321_), .A2(new_n3324_), .ZN(new_n3574_));
  NAND2_X1   g03381(.A1(new_n3325_), .A2(new_n3318_), .ZN(new_n3575_));
  NAND2_X1   g03382(.A1(new_n3575_), .A2(new_n3574_), .ZN(new_n3576_));
  NOR2_X1    g03383(.A1(new_n2274_), .A2(new_n2442_), .ZN(new_n3577_));
  NAND2_X1   g03384(.A1(new_n2636_), .A2(new_n540_), .ZN(new_n3578_));
  NAND2_X1   g03385(.A1(new_n3374_), .A2(new_n1367_), .ZN(new_n3579_));
  AOI22_X1   g03386(.A1(new_n3578_), .A2(new_n3579_), .B1(new_n467_), .B2(new_n3577_), .ZN(new_n3580_));
  AOI22_X1   g03387(.A1(\a[8] ), .A2(\a[34] ), .B1(\a[9] ), .B2(\a[33] ), .ZN(new_n3581_));
  NAND2_X1   g03388(.A1(new_n467_), .A2(new_n3577_), .ZN(new_n3582_));
  NAND3_X1   g03389(.A1(new_n3582_), .A2(new_n3578_), .A3(new_n3579_), .ZN(new_n3583_));
  OAI22_X1   g03390(.A1(new_n3580_), .A2(new_n2779_), .B1(new_n3583_), .B2(new_n3581_), .ZN(new_n3584_));
  NOR2_X1    g03391(.A1(new_n2051_), .A2(new_n2626_), .ZN(new_n3585_));
  INV_X1     g03392(.I(new_n3585_), .ZN(new_n3586_));
  OAI22_X1   g03393(.A1(new_n840_), .A2(new_n3586_), .B1(new_n3405_), .B2(new_n374_), .ZN(new_n3587_));
  NOR2_X1    g03394(.A1(new_n422_), .A2(new_n2524_), .ZN(new_n3588_));
  INV_X1     g03395(.I(new_n3588_), .ZN(new_n3589_));
  NOR2_X1    g03396(.A1(new_n513_), .A2(new_n2051_), .ZN(new_n3590_));
  INV_X1     g03397(.I(new_n3590_), .ZN(new_n3591_));
  NOR2_X1    g03398(.A1(new_n3589_), .A2(new_n3591_), .ZN(new_n3592_));
  INV_X1     g03399(.I(new_n3592_), .ZN(new_n3593_));
  NAND2_X1   g03400(.A1(new_n3593_), .A2(new_n3587_), .ZN(new_n3594_));
  NOR2_X1    g03401(.A1(new_n367_), .A2(new_n2626_), .ZN(new_n3595_));
  NAND2_X1   g03402(.A1(new_n3594_), .A2(new_n3593_), .ZN(new_n3596_));
  AOI21_X1   g03403(.A1(new_n3589_), .A2(new_n3591_), .B(new_n3596_), .ZN(new_n3597_));
  AOI21_X1   g03404(.A1(new_n3594_), .A2(new_n3595_), .B(new_n3597_), .ZN(new_n3598_));
  XOR2_X1    g03405(.A1(new_n3598_), .A2(new_n3382_), .Z(new_n3599_));
  XNOR2_X1   g03406(.A1(new_n3599_), .A2(new_n3584_), .ZN(new_n3600_));
  XOR2_X1    g03407(.A1(new_n3576_), .A2(new_n3600_), .Z(new_n3601_));
  XOR2_X1    g03408(.A1(new_n3601_), .A2(new_n3573_), .Z(new_n3602_));
  XNOR2_X1   g03409(.A1(new_n3535_), .A2(new_n3602_), .ZN(new_n3603_));
  XOR2_X1    g03410(.A1(new_n3603_), .A2(new_n3532_), .Z(new_n3604_));
  XOR2_X1    g03411(.A1(new_n3495_), .A2(new_n3604_), .Z(new_n3605_));
  INV_X1     g03412(.I(new_n3605_), .ZN(new_n3606_));
  NOR2_X1    g03413(.A1(new_n3472_), .A2(new_n3606_), .ZN(new_n3607_));
  INV_X1     g03414(.I(new_n3607_), .ZN(new_n3608_));
  NOR2_X1    g03415(.A1(new_n3471_), .A2(new_n3605_), .ZN(new_n3609_));
  INV_X1     g03416(.I(new_n3609_), .ZN(new_n3610_));
  NAND2_X1   g03417(.A1(new_n3608_), .A2(new_n3610_), .ZN(new_n3611_));
  XOR2_X1    g03418(.A1(new_n3470_), .A2(new_n3611_), .Z(\asquared[43] ));
  OAI21_X1   g03419(.A1(new_n3469_), .A2(new_n3464_), .B(new_n3608_), .ZN(new_n3613_));
  NAND2_X1   g03420(.A1(new_n3613_), .A2(new_n3610_), .ZN(new_n3614_));
  INV_X1     g03421(.I(new_n3495_), .ZN(new_n3615_));
  OAI21_X1   g03422(.A1(new_n3615_), .A2(new_n3604_), .B(new_n3494_), .ZN(new_n3616_));
  INV_X1     g03423(.I(new_n3616_), .ZN(new_n3617_));
  NAND2_X1   g03424(.A1(new_n3517_), .A2(new_n3525_), .ZN(new_n3618_));
  NAND2_X1   g03425(.A1(new_n3512_), .A2(new_n3526_), .ZN(new_n3619_));
  NAND2_X1   g03426(.A1(new_n3619_), .A2(new_n3618_), .ZN(new_n3620_));
  NOR2_X1    g03427(.A1(new_n3569_), .A2(new_n3596_), .ZN(new_n3621_));
  NAND2_X1   g03428(.A1(new_n3569_), .A2(new_n3596_), .ZN(new_n3622_));
  INV_X1     g03429(.I(new_n3622_), .ZN(new_n3623_));
  NOR2_X1    g03430(.A1(new_n3623_), .A2(new_n3621_), .ZN(new_n3624_));
  NAND2_X1   g03431(.A1(new_n3624_), .A2(new_n3544_), .ZN(new_n3625_));
  INV_X1     g03432(.I(new_n3625_), .ZN(new_n3626_));
  NOR2_X1    g03433(.A1(new_n3624_), .A2(new_n3544_), .ZN(new_n3627_));
  NOR2_X1    g03434(.A1(new_n3626_), .A2(new_n3627_), .ZN(new_n3628_));
  NAND2_X1   g03435(.A1(new_n3514_), .A2(new_n3516_), .ZN(new_n3629_));
  OAI21_X1   g03436(.A1(new_n3435_), .A2(new_n3513_), .B(new_n3629_), .ZN(new_n3630_));
  XOR2_X1    g03437(.A1(new_n3555_), .A2(new_n3524_), .Z(new_n3631_));
  XOR2_X1    g03438(.A1(new_n3631_), .A2(new_n3630_), .Z(new_n3632_));
  XOR2_X1    g03439(.A1(new_n3628_), .A2(new_n3632_), .Z(new_n3633_));
  XOR2_X1    g03440(.A1(new_n3633_), .A2(new_n3620_), .Z(new_n3634_));
  INV_X1     g03441(.I(new_n3499_), .ZN(new_n3635_));
  NOR2_X1    g03442(.A1(new_n3635_), .A2(new_n3496_), .ZN(new_n3636_));
  NOR2_X1    g03443(.A1(new_n3636_), .A2(new_n3498_), .ZN(new_n3637_));
  NAND2_X1   g03444(.A1(new_n3399_), .A2(new_n3363_), .ZN(new_n3638_));
  NAND2_X1   g03445(.A1(new_n3501_), .A2(new_n3412_), .ZN(new_n3639_));
  NAND2_X1   g03446(.A1(new_n3639_), .A2(new_n3638_), .ZN(new_n3640_));
  NOR2_X1    g03447(.A1(new_n367_), .A2(new_n2752_), .ZN(new_n3641_));
  NAND3_X1   g03448(.A1(new_n3641_), .A2(\a[11] ), .A3(\a[32] ), .ZN(new_n3642_));
  INV_X1     g03449(.I(new_n3642_), .ZN(new_n3643_));
  NAND4_X1   g03450(.A1(\a[6] ), .A2(\a[12] ), .A3(\a[31] ), .A4(\a[37] ), .ZN(new_n3644_));
  NAND2_X1   g03451(.A1(new_n3210_), .A2(new_n1261_), .ZN(new_n3645_));
  AOI21_X1   g03452(.A1(new_n3645_), .A2(new_n3644_), .B(new_n3643_), .ZN(new_n3646_));
  NAND2_X1   g03453(.A1(\a[12] ), .A2(\a[31] ), .ZN(new_n3647_));
  NOR2_X1    g03454(.A1(new_n3646_), .A2(new_n3643_), .ZN(new_n3648_));
  INV_X1     g03455(.I(new_n3648_), .ZN(new_n3649_));
  AOI21_X1   g03456(.A1(\a[11] ), .A2(\a[32] ), .B(new_n3641_), .ZN(new_n3650_));
  OAI22_X1   g03457(.A1(new_n3649_), .A2(new_n3650_), .B1(new_n3646_), .B2(new_n3647_), .ZN(new_n3651_));
  XNOR2_X1   g03458(.A1(new_n3640_), .A2(new_n3651_), .ZN(new_n3652_));
  XOR2_X1    g03459(.A1(new_n3652_), .A2(new_n3637_), .Z(new_n3653_));
  NAND2_X1   g03460(.A1(new_n3506_), .A2(new_n3502_), .ZN(new_n3654_));
  NAND2_X1   g03461(.A1(new_n3507_), .A2(new_n3500_), .ZN(new_n3655_));
  NAND2_X1   g03462(.A1(new_n3655_), .A2(new_n3654_), .ZN(new_n3656_));
  XOR2_X1    g03463(.A1(new_n3656_), .A2(new_n3653_), .Z(new_n3657_));
  XNOR2_X1   g03464(.A1(new_n3657_), .A2(new_n3634_), .ZN(new_n3658_));
  NAND2_X1   g03465(.A1(new_n3478_), .A2(new_n3488_), .ZN(new_n3659_));
  NAND2_X1   g03466(.A1(new_n3476_), .A2(new_n3489_), .ZN(new_n3660_));
  NAND2_X1   g03467(.A1(new_n3660_), .A2(new_n3659_), .ZN(new_n3661_));
  OAI21_X1   g03468(.A1(new_n3482_), .A2(new_n3447_), .B(new_n3486_), .ZN(new_n3662_));
  NAND2_X1   g03469(.A1(new_n3487_), .A2(new_n3481_), .ZN(new_n3663_));
  NAND2_X1   g03470(.A1(new_n3663_), .A2(new_n3662_), .ZN(new_n3664_));
  NAND4_X1   g03471(.A1(\a[0] ), .A2(\a[3] ), .A3(\a[40] ), .A4(\a[43] ), .ZN(new_n3665_));
  INV_X1     g03472(.I(\a[43] ), .ZN(new_n3666_));
  NOR3_X1    g03473(.A1(new_n3118_), .A2(new_n290_), .A3(new_n3666_), .ZN(new_n3667_));
  NOR2_X1    g03474(.A1(new_n3551_), .A2(new_n370_), .ZN(new_n3668_));
  OAI21_X1   g03475(.A1(new_n3667_), .A2(new_n3668_), .B(new_n3665_), .ZN(new_n3669_));
  NAND3_X1   g03476(.A1(new_n3669_), .A2(\a[4] ), .A3(\a[39] ), .ZN(new_n3670_));
  NAND2_X1   g03477(.A1(new_n3669_), .A2(new_n3665_), .ZN(new_n3671_));
  AOI22_X1   g03478(.A1(\a[0] ), .A2(\a[43] ), .B1(\a[3] ), .B2(\a[40] ), .ZN(new_n3672_));
  OAI21_X1   g03479(.A1(new_n3671_), .A2(new_n3672_), .B(new_n3670_), .ZN(new_n3673_));
  NOR2_X1    g03480(.A1(new_n2189_), .A2(new_n893_), .ZN(new_n3674_));
  NOR2_X1    g03481(.A1(new_n2028_), .A2(new_n1816_), .ZN(new_n3675_));
  NOR2_X1    g03482(.A1(new_n1173_), .A2(new_n2679_), .ZN(new_n3676_));
  NOR2_X1    g03483(.A1(new_n3675_), .A2(new_n3676_), .ZN(new_n3677_));
  NOR2_X1    g03484(.A1(new_n3677_), .A2(new_n3674_), .ZN(new_n3678_));
  NAND2_X1   g03485(.A1(\a[14] ), .A2(\a[29] ), .ZN(new_n3679_));
  AOI22_X1   g03486(.A1(\a[15] ), .A2(\a[28] ), .B1(\a[16] ), .B2(\a[27] ), .ZN(new_n3680_));
  NOR2_X1    g03487(.A1(new_n3678_), .A2(new_n3674_), .ZN(new_n3681_));
  INV_X1     g03488(.I(new_n3681_), .ZN(new_n3682_));
  OAI22_X1   g03489(.A1(new_n3682_), .A2(new_n3680_), .B1(new_n3678_), .B2(new_n3679_), .ZN(new_n3683_));
  XOR2_X1    g03490(.A1(new_n3683_), .A2(new_n3673_), .Z(new_n3684_));
  NAND2_X1   g03491(.A1(new_n1027_), .A2(new_n2176_), .ZN(new_n3685_));
  NAND2_X1   g03492(.A1(new_n2080_), .A2(new_n2629_), .ZN(new_n3686_));
  AOI22_X1   g03493(.A1(new_n3685_), .A2(new_n3686_), .B1(new_n1194_), .B2(new_n1778_), .ZN(new_n3687_));
  NAND2_X1   g03494(.A1(\a[17] ), .A2(\a[26] ), .ZN(new_n3688_));
  AOI22_X1   g03495(.A1(\a[18] ), .A2(\a[25] ), .B1(\a[19] ), .B2(\a[24] ), .ZN(new_n3689_));
  NAND2_X1   g03496(.A1(new_n1778_), .A2(new_n1194_), .ZN(new_n3690_));
  NAND3_X1   g03497(.A1(new_n3685_), .A2(new_n3686_), .A3(new_n3690_), .ZN(new_n3691_));
  OAI22_X1   g03498(.A1(new_n3687_), .A2(new_n3688_), .B1(new_n3691_), .B2(new_n3689_), .ZN(new_n3692_));
  XOR2_X1    g03499(.A1(new_n3684_), .A2(new_n3692_), .Z(new_n3693_));
  NOR2_X1    g03500(.A1(new_n2526_), .A2(new_n413_), .ZN(new_n3694_));
  NOR4_X1    g03501(.A1(new_n422_), .A2(new_n417_), .A3(new_n2274_), .A4(new_n2626_), .ZN(new_n3695_));
  NOR2_X1    g03502(.A1(new_n3405_), .A2(new_n415_), .ZN(new_n3696_));
  NOR2_X1    g03503(.A1(new_n3696_), .A2(new_n3695_), .ZN(new_n3697_));
  NOR2_X1    g03504(.A1(new_n3697_), .A2(new_n3694_), .ZN(new_n3698_));
  NAND2_X1   g03505(.A1(\a[7] ), .A2(\a[36] ), .ZN(new_n3699_));
  AOI22_X1   g03506(.A1(\a[8] ), .A2(\a[35] ), .B1(\a[10] ), .B2(\a[33] ), .ZN(new_n3700_));
  NOR2_X1    g03507(.A1(new_n3698_), .A2(new_n3694_), .ZN(new_n3701_));
  INV_X1     g03508(.I(new_n3701_), .ZN(new_n3702_));
  OAI22_X1   g03509(.A1(new_n3702_), .A2(new_n3700_), .B1(new_n3698_), .B2(new_n3699_), .ZN(new_n3703_));
  AOI21_X1   g03510(.A1(\a[20] ), .A2(\a[23] ), .B(new_n1452_), .ZN(new_n3704_));
  INV_X1     g03511(.I(new_n3704_), .ZN(new_n3705_));
  NOR2_X1    g03512(.A1(new_n1382_), .A2(new_n2385_), .ZN(new_n3706_));
  NOR2_X1    g03513(.A1(new_n403_), .A2(new_n2442_), .ZN(new_n3707_));
  AOI21_X1   g03514(.A1(new_n3705_), .A2(new_n3707_), .B(new_n3706_), .ZN(new_n3708_));
  INV_X1     g03515(.I(new_n3708_), .ZN(new_n3709_));
  OAI21_X1   g03516(.A1(new_n3706_), .A2(new_n3704_), .B(new_n3707_), .ZN(new_n3710_));
  OAI21_X1   g03517(.A1(new_n3709_), .A2(new_n3704_), .B(new_n3710_), .ZN(new_n3711_));
  XNOR2_X1   g03518(.A1(new_n3703_), .A2(new_n3711_), .ZN(new_n3712_));
  NOR2_X1    g03519(.A1(new_n197_), .A2(new_n3327_), .ZN(new_n3713_));
  INV_X1     g03520(.I(new_n3713_), .ZN(new_n3714_));
  AOI22_X1   g03521(.A1(\a[5] ), .A2(\a[38] ), .B1(\a[13] ), .B2(\a[30] ), .ZN(new_n3715_));
  NOR4_X1    g03522(.A1(new_n253_), .A2(new_n597_), .A3(new_n2030_), .A4(new_n2914_), .ZN(new_n3716_));
  NOR3_X1    g03523(.A1(new_n3714_), .A2(new_n3716_), .A3(new_n3715_), .ZN(new_n3717_));
  NOR2_X1    g03524(.A1(new_n3717_), .A2(new_n3716_), .ZN(new_n3718_));
  INV_X1     g03525(.I(new_n3718_), .ZN(new_n3719_));
  OAI22_X1   g03526(.A1(new_n3719_), .A2(new_n3715_), .B1(new_n3714_), .B2(new_n3717_), .ZN(new_n3720_));
  XOR2_X1    g03527(.A1(new_n3712_), .A2(new_n3720_), .Z(new_n3721_));
  XOR2_X1    g03528(.A1(new_n3693_), .A2(new_n3721_), .Z(new_n3722_));
  XNOR2_X1   g03529(.A1(new_n3722_), .A2(new_n3664_), .ZN(new_n3723_));
  XOR2_X1    g03530(.A1(new_n3661_), .A2(new_n3723_), .Z(new_n3724_));
  INV_X1     g03531(.I(new_n3724_), .ZN(new_n3725_));
  NAND2_X1   g03532(.A1(new_n3725_), .A2(new_n3658_), .ZN(new_n3726_));
  OR2_X2     g03533(.A1(new_n3725_), .A2(new_n3658_), .Z(new_n3727_));
  AND2_X2    g03534(.A1(new_n3727_), .A2(new_n3726_), .Z(new_n3728_));
  INV_X1     g03535(.I(new_n3532_), .ZN(new_n3729_));
  NAND2_X1   g03536(.A1(new_n3535_), .A2(new_n3602_), .ZN(new_n3730_));
  OAI21_X1   g03537(.A1(new_n3603_), .A2(new_n3729_), .B(new_n3730_), .ZN(new_n3731_));
  NOR3_X1    g03538(.A1(new_n3508_), .A2(new_n3529_), .A3(new_n3530_), .ZN(new_n3732_));
  NOR2_X1    g03539(.A1(new_n3732_), .A2(new_n3530_), .ZN(new_n3733_));
  NAND2_X1   g03540(.A1(new_n3576_), .A2(new_n3600_), .ZN(new_n3734_));
  NAND2_X1   g03541(.A1(new_n3601_), .A2(new_n3573_), .ZN(new_n3735_));
  NAND2_X1   g03542(.A1(new_n3735_), .A2(new_n3734_), .ZN(new_n3736_));
  NAND2_X1   g03543(.A1(new_n3545_), .A2(new_n3557_), .ZN(new_n3737_));
  NAND2_X1   g03544(.A1(new_n3558_), .A2(new_n3571_), .ZN(new_n3738_));
  NAND2_X1   g03545(.A1(new_n3738_), .A2(new_n3737_), .ZN(new_n3739_));
  INV_X1     g03546(.I(new_n3599_), .ZN(new_n3740_));
  NAND2_X1   g03547(.A1(new_n3740_), .A2(new_n3584_), .ZN(new_n3741_));
  OAI21_X1   g03548(.A1(new_n3381_), .A2(new_n3598_), .B(new_n3741_), .ZN(new_n3742_));
  INV_X1     g03549(.I(new_n3742_), .ZN(new_n3743_));
  NOR2_X1    g03550(.A1(new_n2647_), .A2(new_n3515_), .ZN(new_n3744_));
  AOI21_X1   g03551(.A1(\a[1] ), .A2(\a[42] ), .B(\a[22] ), .ZN(new_n3745_));
  INV_X1     g03552(.I(\a[42] ), .ZN(new_n3746_));
  NOR2_X1    g03553(.A1(new_n1319_), .A2(new_n3746_), .ZN(new_n3747_));
  NOR2_X1    g03554(.A1(new_n3747_), .A2(new_n3745_), .ZN(new_n3748_));
  XOR2_X1    g03555(.A1(new_n3748_), .A2(new_n3744_), .Z(new_n3749_));
  XOR2_X1    g03556(.A1(new_n3749_), .A2(new_n3583_), .Z(new_n3750_));
  NOR2_X1    g03557(.A1(new_n3743_), .A2(new_n3750_), .ZN(new_n3751_));
  INV_X1     g03558(.I(new_n3750_), .ZN(new_n3752_));
  NOR2_X1    g03559(.A1(new_n3742_), .A2(new_n3752_), .ZN(new_n3753_));
  OAI21_X1   g03560(.A1(new_n3751_), .A2(new_n3753_), .B(new_n3739_), .ZN(new_n3754_));
  INV_X1     g03561(.I(new_n3754_), .ZN(new_n3755_));
  NOR3_X1    g03562(.A1(new_n3751_), .A2(new_n3739_), .A3(new_n3753_), .ZN(new_n3756_));
  NOR2_X1    g03563(.A1(new_n3755_), .A2(new_n3756_), .ZN(new_n3757_));
  XNOR2_X1   g03564(.A1(new_n3757_), .A2(new_n3736_), .ZN(new_n3758_));
  XOR2_X1    g03565(.A1(new_n3758_), .A2(new_n3733_), .Z(new_n3759_));
  NAND2_X1   g03566(.A1(new_n3731_), .A2(new_n3759_), .ZN(new_n3760_));
  NAND2_X1   g03567(.A1(new_n3760_), .A2(new_n3731_), .ZN(new_n3761_));
  NAND2_X1   g03568(.A1(new_n3760_), .A2(new_n3759_), .ZN(new_n3762_));
  NAND2_X1   g03569(.A1(new_n3761_), .A2(new_n3762_), .ZN(new_n3763_));
  NAND2_X1   g03570(.A1(new_n3763_), .A2(new_n3728_), .ZN(new_n3764_));
  INV_X1     g03571(.I(new_n3728_), .ZN(new_n3765_));
  NAND3_X1   g03572(.A1(new_n3761_), .A2(new_n3762_), .A3(new_n3765_), .ZN(new_n3766_));
  NAND2_X1   g03573(.A1(new_n3764_), .A2(new_n3766_), .ZN(new_n3767_));
  NOR2_X1    g03574(.A1(new_n3617_), .A2(new_n3767_), .ZN(new_n3768_));
  NAND2_X1   g03575(.A1(new_n3617_), .A2(new_n3767_), .ZN(new_n3769_));
  INV_X1     g03576(.I(new_n3769_), .ZN(new_n3770_));
  NOR2_X1    g03577(.A1(new_n3770_), .A2(new_n3768_), .ZN(new_n3771_));
  XOR2_X1    g03578(.A1(new_n3614_), .A2(new_n3771_), .Z(\asquared[44] ));
  AOI21_X1   g03579(.A1(new_n3613_), .A2(new_n3610_), .B(new_n3770_), .ZN(new_n3773_));
  NOR2_X1    g03580(.A1(new_n3773_), .A2(new_n3768_), .ZN(new_n3774_));
  NAND2_X1   g03581(.A1(new_n3764_), .A2(new_n3760_), .ZN(new_n3775_));
  NAND2_X1   g03582(.A1(new_n3757_), .A2(new_n3736_), .ZN(new_n3776_));
  OAI21_X1   g03583(.A1(new_n3758_), .A2(new_n3733_), .B(new_n3776_), .ZN(new_n3777_));
  OAI21_X1   g03584(.A1(new_n3743_), .A2(new_n3752_), .B(new_n3754_), .ZN(new_n3778_));
  AOI22_X1   g03585(.A1(\a[15] ), .A2(\a[29] ), .B1(\a[17] ), .B2(\a[27] ), .ZN(new_n3779_));
  INV_X1     g03586(.I(new_n3779_), .ZN(new_n3780_));
  NOR2_X1    g03587(.A1(new_n1816_), .A2(new_n982_), .ZN(new_n3781_));
  NOR2_X1    g03588(.A1(new_n225_), .A2(new_n3327_), .ZN(new_n3782_));
  AOI21_X1   g03589(.A1(new_n3780_), .A2(new_n3782_), .B(new_n3781_), .ZN(new_n3783_));
  NAND2_X1   g03590(.A1(new_n3783_), .A2(new_n3780_), .ZN(new_n3784_));
  OAI21_X1   g03591(.A1(new_n3781_), .A2(new_n3779_), .B(new_n3782_), .ZN(new_n3785_));
  NAND2_X1   g03592(.A1(new_n3784_), .A2(new_n3785_), .ZN(new_n3786_));
  NAND2_X1   g03593(.A1(\a[18] ), .A2(\a[26] ), .ZN(new_n3787_));
  NOR2_X1    g03594(.A1(new_n1376_), .A2(new_n1779_), .ZN(new_n3788_));
  NOR2_X1    g03595(.A1(new_n1281_), .A2(new_n2081_), .ZN(new_n3789_));
  NOR2_X1    g03596(.A1(new_n2177_), .A2(new_n1092_), .ZN(new_n3790_));
  NOR2_X1    g03597(.A1(new_n3789_), .A2(new_n3790_), .ZN(new_n3791_));
  NOR2_X1    g03598(.A1(new_n3791_), .A2(new_n3788_), .ZN(new_n3792_));
  AOI22_X1   g03599(.A1(\a[19] ), .A2(\a[25] ), .B1(\a[20] ), .B2(\a[24] ), .ZN(new_n3793_));
  NOR2_X1    g03600(.A1(new_n3792_), .A2(new_n3788_), .ZN(new_n3794_));
  INV_X1     g03601(.I(new_n3794_), .ZN(new_n3795_));
  OAI22_X1   g03602(.A1(new_n3795_), .A2(new_n3793_), .B1(new_n3787_), .B2(new_n3792_), .ZN(new_n3796_));
  XOR2_X1    g03603(.A1(new_n3796_), .A2(new_n3786_), .Z(new_n3797_));
  NAND2_X1   g03604(.A1(\a[6] ), .A2(\a[38] ), .ZN(new_n3798_));
  NOR2_X1    g03605(.A1(new_n513_), .A2(new_n2752_), .ZN(new_n3799_));
  INV_X1     g03606(.I(new_n3799_), .ZN(new_n3800_));
  NOR3_X1    g03607(.A1(new_n3800_), .A2(new_n422_), .A3(new_n2274_), .ZN(new_n3801_));
  NOR2_X1    g03608(.A1(new_n2274_), .A2(new_n2914_), .ZN(new_n3802_));
  NOR2_X1    g03609(.A1(new_n2752_), .A2(new_n2914_), .ZN(new_n3803_));
  AOI22_X1   g03610(.A1(new_n839_), .A2(new_n3802_), .B1(new_n3803_), .B2(new_n479_), .ZN(new_n3804_));
  NOR2_X1    g03611(.A1(new_n3801_), .A2(new_n3804_), .ZN(new_n3805_));
  AOI22_X1   g03612(.A1(\a[7] ), .A2(\a[37] ), .B1(\a[11] ), .B2(\a[33] ), .ZN(new_n3806_));
  INV_X1     g03613(.I(new_n3801_), .ZN(new_n3807_));
  NAND2_X1   g03614(.A1(new_n3807_), .A2(new_n3804_), .ZN(new_n3808_));
  OAI22_X1   g03615(.A1(new_n3808_), .A2(new_n3806_), .B1(new_n3798_), .B2(new_n3805_), .ZN(new_n3809_));
  XOR2_X1    g03616(.A1(new_n3797_), .A2(new_n3809_), .Z(new_n3810_));
  INV_X1     g03617(.I(new_n2681_), .ZN(new_n3811_));
  OAI22_X1   g03618(.A1(new_n2028_), .A2(new_n3811_), .B1(new_n3559_), .B2(new_n3549_), .ZN(new_n3812_));
  NAND4_X1   g03619(.A1(\a[4] ), .A2(\a[14] ), .A3(\a[30] ), .A4(\a[40] ), .ZN(new_n3813_));
  NAND2_X1   g03620(.A1(new_n3812_), .A2(new_n3813_), .ZN(new_n3814_));
  NAND3_X1   g03621(.A1(new_n3814_), .A2(\a[16] ), .A3(\a[28] ), .ZN(new_n3815_));
  AOI22_X1   g03622(.A1(\a[4] ), .A2(\a[40] ), .B1(\a[14] ), .B2(\a[30] ), .ZN(new_n3816_));
  NAND2_X1   g03623(.A1(new_n3814_), .A2(new_n3813_), .ZN(new_n3817_));
  OAI21_X1   g03624(.A1(new_n3816_), .A2(new_n3817_), .B(new_n3815_), .ZN(new_n3818_));
  NOR2_X1    g03625(.A1(new_n355_), .A2(new_n2626_), .ZN(new_n3819_));
  INV_X1     g03626(.I(new_n3819_), .ZN(new_n3820_));
  NOR2_X1    g03627(.A1(new_n2746_), .A2(new_n539_), .ZN(new_n3821_));
  NOR2_X1    g03628(.A1(new_n2442_), .A2(new_n2626_), .ZN(new_n3822_));
  AOI22_X1   g03629(.A1(new_n467_), .A2(new_n3232_), .B1(new_n3822_), .B2(new_n1367_), .ZN(new_n3823_));
  NOR2_X1    g03630(.A1(new_n3821_), .A2(new_n3823_), .ZN(new_n3824_));
  AOI22_X1   g03631(.A1(\a[9] ), .A2(\a[35] ), .B1(\a[10] ), .B2(\a[34] ), .ZN(new_n3825_));
  NOR2_X1    g03632(.A1(new_n3824_), .A2(new_n3821_), .ZN(new_n3826_));
  INV_X1     g03633(.I(new_n3826_), .ZN(new_n3827_));
  OAI22_X1   g03634(.A1(new_n3827_), .A2(new_n3825_), .B1(new_n3820_), .B2(new_n3824_), .ZN(new_n3828_));
  XNOR2_X1   g03635(.A1(new_n3818_), .A2(new_n3828_), .ZN(new_n3829_));
  AOI22_X1   g03636(.A1(\a[12] ), .A2(\a[32] ), .B1(\a[13] ), .B2(\a[31] ), .ZN(new_n3830_));
  NOR2_X1    g03637(.A1(new_n253_), .A2(new_n3116_), .ZN(new_n3831_));
  INV_X1     g03638(.I(new_n3831_), .ZN(new_n3832_));
  INV_X1     g03639(.I(new_n3210_), .ZN(new_n3833_));
  NOR2_X1    g03640(.A1(new_n1265_), .A2(new_n3833_), .ZN(new_n3834_));
  NOR3_X1    g03641(.A1(new_n3834_), .A2(new_n3830_), .A3(new_n3832_), .ZN(new_n3835_));
  NOR2_X1    g03642(.A1(new_n3835_), .A2(new_n3834_), .ZN(new_n3836_));
  INV_X1     g03643(.I(new_n3836_), .ZN(new_n3837_));
  OAI22_X1   g03644(.A1(new_n3837_), .A2(new_n3830_), .B1(new_n3832_), .B2(new_n3835_), .ZN(new_n3838_));
  XOR2_X1    g03645(.A1(new_n3829_), .A2(new_n3838_), .Z(new_n3839_));
  XNOR2_X1   g03646(.A1(new_n3810_), .A2(new_n3839_), .ZN(new_n3840_));
  XOR2_X1    g03647(.A1(new_n3778_), .A2(new_n3840_), .Z(new_n3841_));
  XOR2_X1    g03648(.A1(new_n3777_), .A2(new_n3841_), .Z(new_n3842_));
  NAND2_X1   g03649(.A1(new_n3640_), .A2(new_n3651_), .ZN(new_n3843_));
  OAI21_X1   g03650(.A1(new_n3652_), .A2(new_n3637_), .B(new_n3843_), .ZN(new_n3844_));
  NAND2_X1   g03651(.A1(\a[1] ), .A2(\a[43] ), .ZN(new_n3845_));
  XNOR2_X1   g03652(.A1(new_n1300_), .A2(new_n3845_), .ZN(new_n3846_));
  NOR2_X1    g03653(.A1(new_n3709_), .A2(new_n3846_), .ZN(new_n3847_));
  INV_X1     g03654(.I(new_n3846_), .ZN(new_n3848_));
  NOR2_X1    g03655(.A1(new_n3708_), .A2(new_n3848_), .ZN(new_n3849_));
  NOR2_X1    g03656(.A1(new_n3847_), .A2(new_n3849_), .ZN(new_n3850_));
  INV_X1     g03657(.I(new_n3850_), .ZN(new_n3851_));
  NAND2_X1   g03658(.A1(new_n3851_), .A2(new_n3701_), .ZN(new_n3852_));
  NOR2_X1    g03659(.A1(new_n3851_), .A2(new_n3701_), .ZN(new_n3853_));
  INV_X1     g03660(.I(new_n3853_), .ZN(new_n3854_));
  AND2_X2    g03661(.A1(new_n3854_), .A2(new_n3852_), .Z(new_n3855_));
  XOR2_X1    g03662(.A1(new_n3681_), .A2(new_n3648_), .Z(new_n3856_));
  INV_X1     g03663(.I(new_n3747_), .ZN(new_n3857_));
  AOI22_X1   g03664(.A1(\a[0] ), .A2(\a[44] ), .B1(\a[2] ), .B2(\a[42] ), .ZN(new_n3858_));
  INV_X1     g03665(.I(\a[44] ), .ZN(new_n3859_));
  NOR2_X1    g03666(.A1(new_n3746_), .A2(new_n3859_), .ZN(new_n3860_));
  INV_X1     g03667(.I(new_n3860_), .ZN(new_n3861_));
  NOR2_X1    g03668(.A1(new_n3861_), .A2(new_n412_), .ZN(new_n3862_));
  NOR3_X1    g03669(.A1(new_n3857_), .A2(new_n3862_), .A3(new_n3858_), .ZN(new_n3863_));
  NOR2_X1    g03670(.A1(new_n3863_), .A2(new_n3862_), .ZN(new_n3864_));
  INV_X1     g03671(.I(new_n3864_), .ZN(new_n3865_));
  OAI22_X1   g03672(.A1(new_n3865_), .A2(new_n3858_), .B1(new_n3863_), .B2(new_n3857_), .ZN(new_n3866_));
  XNOR2_X1   g03673(.A1(new_n3856_), .A2(new_n3866_), .ZN(new_n3867_));
  XOR2_X1    g03674(.A1(new_n3855_), .A2(new_n3867_), .Z(new_n3868_));
  XNOR2_X1   g03675(.A1(new_n3868_), .A2(new_n3844_), .ZN(new_n3869_));
  NAND2_X1   g03676(.A1(new_n3628_), .A2(new_n3632_), .ZN(new_n3870_));
  NAND2_X1   g03677(.A1(new_n3633_), .A2(new_n3620_), .ZN(new_n3871_));
  NAND2_X1   g03678(.A1(new_n3871_), .A2(new_n3870_), .ZN(new_n3872_));
  NOR2_X1    g03679(.A1(new_n3626_), .A2(new_n3623_), .ZN(new_n3873_));
  NAND2_X1   g03680(.A1(new_n3555_), .A2(new_n3524_), .ZN(new_n3874_));
  NAND2_X1   g03681(.A1(new_n3631_), .A2(new_n3630_), .ZN(new_n3875_));
  NAND2_X1   g03682(.A1(new_n3875_), .A2(new_n3874_), .ZN(new_n3876_));
  NAND2_X1   g03683(.A1(new_n3748_), .A2(new_n3744_), .ZN(new_n3877_));
  NAND2_X1   g03684(.A1(new_n3749_), .A2(new_n3583_), .ZN(new_n3878_));
  NAND2_X1   g03685(.A1(new_n3878_), .A2(new_n3877_), .ZN(new_n3879_));
  XOR2_X1    g03686(.A1(new_n3876_), .A2(new_n3879_), .Z(new_n3880_));
  XNOR2_X1   g03687(.A1(new_n3880_), .A2(new_n3873_), .ZN(new_n3881_));
  XOR2_X1    g03688(.A1(new_n3872_), .A2(new_n3881_), .Z(new_n3882_));
  XOR2_X1    g03689(.A1(new_n3882_), .A2(new_n3869_), .Z(new_n3883_));
  XNOR2_X1   g03690(.A1(new_n3842_), .A2(new_n3883_), .ZN(new_n3884_));
  INV_X1     g03691(.I(new_n3884_), .ZN(new_n3885_));
  NAND2_X1   g03692(.A1(new_n3661_), .A2(new_n3723_), .ZN(new_n3886_));
  NAND2_X1   g03693(.A1(new_n3727_), .A2(new_n3886_), .ZN(new_n3887_));
  NAND2_X1   g03694(.A1(new_n3656_), .A2(new_n3653_), .ZN(new_n3888_));
  NAND2_X1   g03695(.A1(new_n3657_), .A2(new_n3634_), .ZN(new_n3889_));
  NAND2_X1   g03696(.A1(new_n3889_), .A2(new_n3888_), .ZN(new_n3890_));
  INV_X1     g03697(.I(new_n3722_), .ZN(new_n3891_));
  NAND2_X1   g03698(.A1(new_n3891_), .A2(new_n3664_), .ZN(new_n3892_));
  INV_X1     g03699(.I(new_n3721_), .ZN(new_n3893_));
  NAND2_X1   g03700(.A1(new_n3893_), .A2(new_n3693_), .ZN(new_n3894_));
  NAND2_X1   g03701(.A1(new_n3892_), .A2(new_n3894_), .ZN(new_n3895_));
  XOR2_X1    g03702(.A1(new_n3671_), .A2(new_n3719_), .Z(new_n3896_));
  XOR2_X1    g03703(.A1(new_n3896_), .A2(new_n3691_), .Z(new_n3897_));
  NAND2_X1   g03704(.A1(new_n3703_), .A2(new_n3711_), .ZN(new_n3898_));
  INV_X1     g03705(.I(new_n3720_), .ZN(new_n3899_));
  OAI21_X1   g03706(.A1(new_n3712_), .A2(new_n3899_), .B(new_n3898_), .ZN(new_n3900_));
  NAND2_X1   g03707(.A1(new_n3683_), .A2(new_n3673_), .ZN(new_n3901_));
  NAND2_X1   g03708(.A1(new_n3684_), .A2(new_n3692_), .ZN(new_n3902_));
  NAND2_X1   g03709(.A1(new_n3902_), .A2(new_n3901_), .ZN(new_n3903_));
  XOR2_X1    g03710(.A1(new_n3903_), .A2(new_n3900_), .Z(new_n3904_));
  XOR2_X1    g03711(.A1(new_n3904_), .A2(new_n3897_), .Z(new_n3905_));
  XOR2_X1    g03712(.A1(new_n3895_), .A2(new_n3905_), .Z(new_n3906_));
  XOR2_X1    g03713(.A1(new_n3890_), .A2(new_n3906_), .Z(new_n3907_));
  XOR2_X1    g03714(.A1(new_n3887_), .A2(new_n3907_), .Z(new_n3908_));
  XOR2_X1    g03715(.A1(new_n3908_), .A2(new_n3885_), .Z(new_n3909_));
  NOR2_X1    g03716(.A1(new_n3909_), .A2(new_n3775_), .ZN(new_n3910_));
  INV_X1     g03717(.I(new_n3910_), .ZN(new_n3911_));
  NAND2_X1   g03718(.A1(new_n3909_), .A2(new_n3775_), .ZN(new_n3912_));
  NAND2_X1   g03719(.A1(new_n3911_), .A2(new_n3912_), .ZN(new_n3913_));
  XOR2_X1    g03720(.A1(new_n3774_), .A2(new_n3913_), .Z(\asquared[45] ));
  OAI21_X1   g03721(.A1(new_n3773_), .A2(new_n3768_), .B(new_n3911_), .ZN(new_n3915_));
  NAND2_X1   g03722(.A1(new_n3915_), .A2(new_n3912_), .ZN(new_n3916_));
  NAND2_X1   g03723(.A1(new_n3887_), .A2(new_n3907_), .ZN(new_n3917_));
  NAND2_X1   g03724(.A1(new_n3908_), .A2(new_n3885_), .ZN(new_n3918_));
  NAND2_X1   g03725(.A1(new_n3918_), .A2(new_n3917_), .ZN(new_n3919_));
  INV_X1     g03726(.I(new_n3839_), .ZN(new_n3920_));
  NAND2_X1   g03727(.A1(new_n3920_), .A2(new_n3810_), .ZN(new_n3921_));
  NAND2_X1   g03728(.A1(new_n3778_), .A2(new_n3840_), .ZN(new_n3922_));
  NAND2_X1   g03729(.A1(new_n3922_), .A2(new_n3921_), .ZN(new_n3923_));
  NAND2_X1   g03730(.A1(new_n3872_), .A2(new_n3881_), .ZN(new_n3924_));
  NAND2_X1   g03731(.A1(new_n3882_), .A2(new_n3869_), .ZN(new_n3925_));
  NAND2_X1   g03732(.A1(new_n3925_), .A2(new_n3924_), .ZN(new_n3926_));
  XOR2_X1    g03733(.A1(new_n3923_), .A2(new_n3926_), .Z(new_n3927_));
  NOR2_X1    g03734(.A1(new_n2442_), .A2(new_n3116_), .ZN(new_n3928_));
  INV_X1     g03735(.I(new_n3928_), .ZN(new_n3929_));
  NOR2_X1    g03736(.A1(new_n840_), .A2(new_n3929_), .ZN(new_n3930_));
  NOR3_X1    g03737(.A1(new_n3046_), .A2(new_n536_), .A3(new_n3116_), .ZN(new_n3931_));
  INV_X1     g03738(.I(new_n3577_), .ZN(new_n3932_));
  NOR2_X1    g03739(.A1(new_n3932_), .A2(new_n619_), .ZN(new_n3933_));
  NOR2_X1    g03740(.A1(new_n3933_), .A2(new_n3931_), .ZN(new_n3934_));
  NOR2_X1    g03741(.A1(new_n3934_), .A2(new_n3930_), .ZN(new_n3935_));
  NAND2_X1   g03742(.A1(\a[12] ), .A2(\a[33] ), .ZN(new_n3936_));
  NOR2_X1    g03743(.A1(new_n3935_), .A2(new_n3930_), .ZN(new_n3937_));
  INV_X1     g03744(.I(new_n3937_), .ZN(new_n3938_));
  AOI22_X1   g03745(.A1(\a[6] ), .A2(\a[39] ), .B1(\a[11] ), .B2(\a[34] ), .ZN(new_n3939_));
  OAI22_X1   g03746(.A1(new_n3938_), .A2(new_n3939_), .B1(new_n3935_), .B2(new_n3936_), .ZN(new_n3940_));
  NAND2_X1   g03747(.A1(\a[15] ), .A2(\a[30] ), .ZN(new_n3941_));
  NOR2_X1    g03748(.A1(new_n1428_), .A2(new_n2679_), .ZN(new_n3942_));
  INV_X1     g03749(.I(new_n982_), .ZN(new_n3943_));
  AOI22_X1   g03750(.A1(new_n1288_), .A2(new_n2254_), .B1(new_n2681_), .B2(new_n3943_), .ZN(new_n3944_));
  NOR2_X1    g03751(.A1(new_n3942_), .A2(new_n3944_), .ZN(new_n3945_));
  AOI22_X1   g03752(.A1(\a[16] ), .A2(\a[29] ), .B1(\a[17] ), .B2(\a[28] ), .ZN(new_n3946_));
  NOR2_X1    g03753(.A1(new_n3945_), .A2(new_n3942_), .ZN(new_n3947_));
  INV_X1     g03754(.I(new_n3947_), .ZN(new_n3948_));
  OAI22_X1   g03755(.A1(new_n3948_), .A2(new_n3946_), .B1(new_n3941_), .B2(new_n3945_), .ZN(new_n3949_));
  XOR2_X1    g03756(.A1(new_n3940_), .A2(new_n3949_), .Z(new_n3950_));
  NOR2_X1    g03757(.A1(new_n1301_), .A2(new_n3845_), .ZN(new_n3951_));
  AOI21_X1   g03758(.A1(\a[3] ), .A2(\a[42] ), .B(new_n3951_), .ZN(new_n3952_));
  NOR2_X1    g03759(.A1(new_n1464_), .A2(new_n3859_), .ZN(new_n3953_));
  INV_X1     g03760(.I(new_n3953_), .ZN(new_n3954_));
  NOR2_X1    g03761(.A1(new_n194_), .A2(new_n3859_), .ZN(new_n3955_));
  OAI21_X1   g03762(.A1(\a[23] ), .A2(new_n3955_), .B(new_n3954_), .ZN(new_n3956_));
  NOR4_X1    g03763(.A1(new_n1301_), .A2(new_n225_), .A3(new_n3746_), .A4(new_n3845_), .ZN(new_n3957_));
  NOR3_X1    g03764(.A1(new_n3956_), .A2(new_n3957_), .A3(new_n3952_), .ZN(new_n3958_));
  NOR2_X1    g03765(.A1(new_n3958_), .A2(new_n3957_), .ZN(new_n3959_));
  INV_X1     g03766(.I(new_n3959_), .ZN(new_n3960_));
  OAI22_X1   g03767(.A1(new_n3960_), .A2(new_n3952_), .B1(new_n3956_), .B2(new_n3958_), .ZN(new_n3961_));
  XNOR2_X1   g03768(.A1(new_n3950_), .A2(new_n3961_), .ZN(new_n3962_));
  INV_X1     g03769(.I(new_n3962_), .ZN(new_n3963_));
  NAND2_X1   g03770(.A1(new_n3876_), .A2(new_n3879_), .ZN(new_n3964_));
  INV_X1     g03771(.I(new_n3880_), .ZN(new_n3965_));
  OAI21_X1   g03772(.A1(new_n3965_), .A2(new_n3873_), .B(new_n3964_), .ZN(new_n3966_));
  XOR2_X1    g03773(.A1(new_n3864_), .A2(new_n3783_), .Z(new_n3967_));
  INV_X1     g03774(.I(new_n3967_), .ZN(new_n3968_));
  NOR2_X1    g03775(.A1(new_n3968_), .A2(new_n3794_), .ZN(new_n3969_));
  NOR2_X1    g03776(.A1(new_n3967_), .A2(new_n3795_), .ZN(new_n3970_));
  NOR2_X1    g03777(.A1(new_n3969_), .A2(new_n3970_), .ZN(new_n3971_));
  XOR2_X1    g03778(.A1(new_n3966_), .A2(new_n3971_), .Z(new_n3972_));
  XOR2_X1    g03779(.A1(new_n3972_), .A2(new_n3963_), .Z(new_n3973_));
  XNOR2_X1   g03780(.A1(new_n3927_), .A2(new_n3973_), .ZN(new_n3974_));
  INV_X1     g03781(.I(new_n3974_), .ZN(new_n3975_));
  NAND2_X1   g03782(.A1(new_n3777_), .A2(new_n3841_), .ZN(new_n3976_));
  NAND2_X1   g03783(.A1(new_n3842_), .A2(new_n3883_), .ZN(new_n3977_));
  NAND2_X1   g03784(.A1(new_n3977_), .A2(new_n3976_), .ZN(new_n3978_));
  XOR2_X1    g03785(.A1(new_n3978_), .A2(new_n3975_), .Z(new_n3979_));
  XOR2_X1    g03786(.A1(new_n3817_), .A2(new_n3808_), .Z(new_n3980_));
  XOR2_X1    g03787(.A1(new_n3980_), .A2(new_n3837_), .Z(new_n3981_));
  NAND2_X1   g03788(.A1(new_n3818_), .A2(new_n3828_), .ZN(new_n3982_));
  INV_X1     g03789(.I(new_n3829_), .ZN(new_n3983_));
  NAND2_X1   g03790(.A1(new_n3983_), .A2(new_n3838_), .ZN(new_n3984_));
  NAND2_X1   g03791(.A1(new_n3984_), .A2(new_n3982_), .ZN(new_n3985_));
  NAND2_X1   g03792(.A1(new_n3796_), .A2(new_n3786_), .ZN(new_n3986_));
  NAND2_X1   g03793(.A1(new_n3797_), .A2(new_n3809_), .ZN(new_n3987_));
  NAND2_X1   g03794(.A1(new_n3987_), .A2(new_n3986_), .ZN(new_n3988_));
  XOR2_X1    g03795(.A1(new_n3985_), .A2(new_n3988_), .Z(new_n3989_));
  XOR2_X1    g03796(.A1(new_n3989_), .A2(new_n3981_), .Z(new_n3990_));
  INV_X1     g03797(.I(new_n3855_), .ZN(new_n3991_));
  INV_X1     g03798(.I(new_n3868_), .ZN(new_n3992_));
  NAND2_X1   g03799(.A1(new_n3992_), .A2(new_n3844_), .ZN(new_n3993_));
  OAI21_X1   g03800(.A1(new_n3991_), .A2(new_n3867_), .B(new_n3993_), .ZN(new_n3994_));
  NOR2_X1    g03801(.A1(new_n3853_), .A2(new_n3849_), .ZN(new_n3995_));
  NAND2_X1   g03802(.A1(new_n3856_), .A2(new_n3866_), .ZN(new_n3996_));
  OAI21_X1   g03803(.A1(new_n3648_), .A2(new_n3681_), .B(new_n3996_), .ZN(new_n3997_));
  NAND2_X1   g03804(.A1(new_n3671_), .A2(new_n3719_), .ZN(new_n3998_));
  NAND2_X1   g03805(.A1(new_n3896_), .A2(new_n3691_), .ZN(new_n3999_));
  NAND2_X1   g03806(.A1(new_n3999_), .A2(new_n3998_), .ZN(new_n4000_));
  XOR2_X1    g03807(.A1(new_n3997_), .A2(new_n4000_), .Z(new_n4001_));
  XNOR2_X1   g03808(.A1(new_n4001_), .A2(new_n3995_), .ZN(new_n4002_));
  XOR2_X1    g03809(.A1(new_n3994_), .A2(new_n4002_), .Z(new_n4003_));
  XNOR2_X1   g03810(.A1(new_n4003_), .A2(new_n3990_), .ZN(new_n4004_));
  NAND2_X1   g03811(.A1(new_n3895_), .A2(new_n3905_), .ZN(new_n4005_));
  NAND2_X1   g03812(.A1(new_n3890_), .A2(new_n3906_), .ZN(new_n4006_));
  NAND2_X1   g03813(.A1(new_n4006_), .A2(new_n4005_), .ZN(new_n4007_));
  NOR2_X1    g03814(.A1(new_n1376_), .A2(new_n2177_), .ZN(new_n4008_));
  INV_X1     g03815(.I(new_n4008_), .ZN(new_n4009_));
  INV_X1     g03816(.I(new_n2246_), .ZN(new_n4010_));
  OAI22_X1   g03817(.A1(new_n1281_), .A2(new_n4010_), .B1(new_n1972_), .B2(new_n1092_), .ZN(new_n4011_));
  NAND2_X1   g03818(.A1(new_n4011_), .A2(new_n4009_), .ZN(new_n4012_));
  NAND3_X1   g03819(.A1(new_n4012_), .A2(\a[18] ), .A3(\a[27] ), .ZN(new_n4013_));
  AOI22_X1   g03820(.A1(\a[19] ), .A2(\a[26] ), .B1(\a[20] ), .B2(\a[25] ), .ZN(new_n4014_));
  NAND2_X1   g03821(.A1(new_n4012_), .A2(new_n4009_), .ZN(new_n4015_));
  OAI21_X1   g03822(.A1(new_n4014_), .A2(new_n4015_), .B(new_n4013_), .ZN(new_n4016_));
  XOR2_X1    g03823(.A1(new_n4016_), .A2(new_n3826_), .Z(new_n4017_));
  NOR4_X1    g03824(.A1(new_n253_), .A2(new_n597_), .A3(new_n2200_), .A4(new_n3221_), .ZN(new_n4018_));
  NOR2_X1    g03825(.A1(new_n759_), .A2(new_n3221_), .ZN(new_n4019_));
  NAND3_X1   g03826(.A1(new_n4019_), .A2(\a[5] ), .A3(\a[31] ), .ZN(new_n4020_));
  NAND2_X1   g03827(.A1(new_n760_), .A2(new_n3210_), .ZN(new_n4021_));
  AOI21_X1   g03828(.A1(new_n4021_), .A2(new_n4020_), .B(new_n4018_), .ZN(new_n4022_));
  NAND2_X1   g03829(.A1(\a[14] ), .A2(\a[31] ), .ZN(new_n4023_));
  OR2_X2     g03830(.A1(new_n4022_), .A2(new_n4018_), .Z(new_n4024_));
  AOI22_X1   g03831(.A1(\a[5] ), .A2(\a[40] ), .B1(\a[13] ), .B2(\a[32] ), .ZN(new_n4025_));
  OAI22_X1   g03832(.A1(new_n4024_), .A2(new_n4025_), .B1(new_n4022_), .B2(new_n4023_), .ZN(new_n4026_));
  XNOR2_X1   g03833(.A1(new_n4017_), .A2(new_n4026_), .ZN(new_n4027_));
  NOR2_X1    g03834(.A1(new_n3327_), .A2(new_n3666_), .ZN(new_n4028_));
  NAND2_X1   g03835(.A1(new_n4028_), .A2(new_n252_), .ZN(new_n4029_));
  INV_X1     g03836(.I(\a[45] ), .ZN(new_n4030_));
  NOR2_X1    g03837(.A1(new_n3327_), .A2(new_n4030_), .ZN(new_n4031_));
  INV_X1     g03838(.I(new_n4031_), .ZN(new_n4032_));
  NOR2_X1    g03839(.A1(new_n3666_), .A2(new_n4030_), .ZN(new_n4033_));
  INV_X1     g03840(.I(new_n4033_), .ZN(new_n4034_));
  OAI22_X1   g03841(.A1(new_n412_), .A2(new_n4034_), .B1(new_n4032_), .B2(new_n595_), .ZN(new_n4035_));
  NAND2_X1   g03842(.A1(new_n4035_), .A2(new_n4029_), .ZN(new_n4036_));
  NAND3_X1   g03843(.A1(new_n4036_), .A2(\a[0] ), .A3(\a[45] ), .ZN(new_n4037_));
  AOI22_X1   g03844(.A1(\a[2] ), .A2(\a[43] ), .B1(\a[4] ), .B2(\a[41] ), .ZN(new_n4038_));
  NAND2_X1   g03845(.A1(new_n4036_), .A2(new_n4029_), .ZN(new_n4039_));
  OAI21_X1   g03846(.A1(new_n4038_), .A2(new_n4039_), .B(new_n4037_), .ZN(new_n4040_));
  NAND2_X1   g03847(.A1(\a[7] ), .A2(\a[38] ), .ZN(new_n4041_));
  NAND2_X1   g03848(.A1(new_n2915_), .A2(new_n1290_), .ZN(new_n4042_));
  NAND2_X1   g03849(.A1(new_n3803_), .A2(new_n693_), .ZN(new_n4043_));
  AOI22_X1   g03850(.A1(new_n4042_), .A2(new_n4043_), .B1(new_n467_), .B2(new_n3037_), .ZN(new_n4044_));
  AOI22_X1   g03851(.A1(\a[8] ), .A2(\a[37] ), .B1(\a[9] ), .B2(\a[36] ), .ZN(new_n4045_));
  NAND2_X1   g03852(.A1(new_n467_), .A2(new_n3037_), .ZN(new_n4046_));
  NAND3_X1   g03853(.A1(new_n4046_), .A2(new_n4042_), .A3(new_n4043_), .ZN(new_n4047_));
  OAI22_X1   g03854(.A1(new_n4044_), .A2(new_n4041_), .B1(new_n4047_), .B2(new_n4045_), .ZN(new_n4048_));
  XNOR2_X1   g03855(.A1(new_n4040_), .A2(new_n4048_), .ZN(new_n4049_));
  NAND2_X1   g03856(.A1(new_n2385_), .A2(new_n1665_), .ZN(new_n4050_));
  INV_X1     g03857(.I(new_n4050_), .ZN(new_n4051_));
  NOR2_X1    g03858(.A1(new_n417_), .A2(new_n2524_), .ZN(new_n4052_));
  INV_X1     g03859(.I(new_n4052_), .ZN(new_n4053_));
  NOR2_X1    g03860(.A1(new_n1456_), .A2(new_n1529_), .ZN(new_n4054_));
  NOR3_X1    g03861(.A1(new_n4051_), .A2(new_n4054_), .A3(new_n4053_), .ZN(new_n4055_));
  NOR2_X1    g03862(.A1(new_n4055_), .A2(new_n4054_), .ZN(new_n4056_));
  INV_X1     g03863(.I(new_n4056_), .ZN(new_n4057_));
  OAI22_X1   g03864(.A1(new_n4057_), .A2(new_n4051_), .B1(new_n4053_), .B2(new_n4055_), .ZN(new_n4058_));
  INV_X1     g03865(.I(new_n4058_), .ZN(new_n4059_));
  XOR2_X1    g03866(.A1(new_n4049_), .A2(new_n4059_), .Z(new_n4060_));
  XOR2_X1    g03867(.A1(new_n4027_), .A2(new_n4060_), .Z(new_n4061_));
  NAND2_X1   g03868(.A1(new_n3903_), .A2(new_n3900_), .ZN(new_n4062_));
  NAND2_X1   g03869(.A1(new_n3904_), .A2(new_n3897_), .ZN(new_n4063_));
  NAND2_X1   g03870(.A1(new_n4063_), .A2(new_n4062_), .ZN(new_n4064_));
  XNOR2_X1   g03871(.A1(new_n4064_), .A2(new_n4061_), .ZN(new_n4065_));
  INV_X1     g03872(.I(new_n4065_), .ZN(new_n4066_));
  XOR2_X1    g03873(.A1(new_n4007_), .A2(new_n4066_), .Z(new_n4067_));
  XNOR2_X1   g03874(.A1(new_n4067_), .A2(new_n4004_), .ZN(new_n4068_));
  XOR2_X1    g03875(.A1(new_n3979_), .A2(new_n4068_), .Z(new_n4069_));
  NOR2_X1    g03876(.A1(new_n3919_), .A2(new_n4069_), .ZN(new_n4070_));
  NAND2_X1   g03877(.A1(new_n3919_), .A2(new_n4069_), .ZN(new_n4071_));
  INV_X1     g03878(.I(new_n4071_), .ZN(new_n4072_));
  NOR2_X1    g03879(.A1(new_n4072_), .A2(new_n4070_), .ZN(new_n4073_));
  XOR2_X1    g03880(.A1(new_n3916_), .A2(new_n4073_), .Z(\asquared[46] ));
  AOI21_X1   g03881(.A1(new_n3915_), .A2(new_n3912_), .B(new_n4070_), .ZN(new_n4075_));
  NOR2_X1    g03882(.A1(new_n4075_), .A2(new_n4072_), .ZN(new_n4076_));
  NAND2_X1   g03883(.A1(new_n3978_), .A2(new_n3975_), .ZN(new_n4077_));
  NAND2_X1   g03884(.A1(new_n3979_), .A2(new_n4068_), .ZN(new_n4078_));
  NAND2_X1   g03885(.A1(new_n4078_), .A2(new_n4077_), .ZN(new_n4079_));
  NAND2_X1   g03886(.A1(new_n4007_), .A2(new_n4066_), .ZN(new_n4080_));
  INV_X1     g03887(.I(new_n4067_), .ZN(new_n4081_));
  OAI21_X1   g03888(.A1(new_n4081_), .A2(new_n4004_), .B(new_n4080_), .ZN(new_n4082_));
  NAND2_X1   g03889(.A1(new_n3817_), .A2(new_n3808_), .ZN(new_n4083_));
  NAND2_X1   g03890(.A1(new_n3980_), .A2(new_n3837_), .ZN(new_n4084_));
  NAND2_X1   g03891(.A1(new_n4084_), .A2(new_n4083_), .ZN(new_n4085_));
  AOI22_X1   g03892(.A1(\a[5] ), .A2(\a[41] ), .B1(\a[15] ), .B2(\a[31] ), .ZN(new_n4086_));
  NOR4_X1    g03893(.A1(new_n253_), .A2(new_n717_), .A3(new_n2051_), .A4(new_n3327_), .ZN(new_n4087_));
  NOR3_X1    g03894(.A1(new_n4086_), .A2(new_n197_), .A3(new_n3859_), .ZN(new_n4088_));
  NOR2_X1    g03895(.A1(new_n4088_), .A2(new_n4087_), .ZN(new_n4089_));
  INV_X1     g03896(.I(new_n4089_), .ZN(new_n4090_));
  NOR2_X1    g03897(.A1(new_n197_), .A2(new_n3859_), .ZN(new_n4091_));
  OAI21_X1   g03898(.A1(new_n4087_), .A2(new_n4086_), .B(new_n4091_), .ZN(new_n4092_));
  OAI21_X1   g03899(.A1(new_n4090_), .A2(new_n4086_), .B(new_n4092_), .ZN(new_n4093_));
  NOR2_X1    g03900(.A1(new_n597_), .A2(new_n2274_), .ZN(new_n4094_));
  NOR2_X1    g03901(.A1(new_n367_), .A2(new_n3221_), .ZN(new_n4095_));
  NOR2_X1    g03902(.A1(new_n767_), .A2(new_n2637_), .ZN(new_n4096_));
  AOI21_X1   g03903(.A1(new_n2963_), .A2(new_n4019_), .B(new_n4096_), .ZN(new_n4097_));
  AOI21_X1   g03904(.A1(new_n4094_), .A2(new_n4095_), .B(new_n4097_), .ZN(new_n4098_));
  NAND2_X1   g03905(.A1(\a[14] ), .A2(\a[32] ), .ZN(new_n4099_));
  NAND2_X1   g03906(.A1(new_n4094_), .A2(new_n4095_), .ZN(new_n4100_));
  INV_X1     g03907(.I(new_n4100_), .ZN(new_n4101_));
  NOR2_X1    g03908(.A1(new_n4098_), .A2(new_n4101_), .ZN(new_n4102_));
  INV_X1     g03909(.I(new_n4102_), .ZN(new_n4103_));
  NOR2_X1    g03910(.A1(new_n4094_), .A2(new_n4095_), .ZN(new_n4104_));
  OAI22_X1   g03911(.A1(new_n4103_), .A2(new_n4104_), .B1(new_n4098_), .B2(new_n4099_), .ZN(new_n4105_));
  XOR2_X1    g03912(.A1(new_n4105_), .A2(new_n4093_), .Z(new_n4106_));
  XOR2_X1    g03913(.A1(new_n4106_), .A2(new_n4085_), .Z(new_n4107_));
  NAND2_X1   g03914(.A1(new_n3997_), .A2(new_n4000_), .ZN(new_n4108_));
  INV_X1     g03915(.I(new_n4001_), .ZN(new_n4109_));
  OAI21_X1   g03916(.A1(new_n4109_), .A2(new_n3995_), .B(new_n4108_), .ZN(new_n4110_));
  NOR2_X1    g03917(.A1(new_n4015_), .A2(new_n3948_), .ZN(new_n4111_));
  NAND2_X1   g03918(.A1(new_n4015_), .A2(new_n3948_), .ZN(new_n4112_));
  INV_X1     g03919(.I(new_n4112_), .ZN(new_n4113_));
  NOR2_X1    g03920(.A1(new_n4113_), .A2(new_n4111_), .ZN(new_n4114_));
  NOR2_X1    g03921(.A1(new_n4114_), .A2(new_n3938_), .ZN(new_n4115_));
  NAND2_X1   g03922(.A1(new_n4114_), .A2(new_n3938_), .ZN(new_n4116_));
  INV_X1     g03923(.I(new_n4116_), .ZN(new_n4117_));
  NOR2_X1    g03924(.A1(new_n4117_), .A2(new_n4115_), .ZN(new_n4118_));
  XOR2_X1    g03925(.A1(new_n4110_), .A2(new_n4118_), .Z(new_n4119_));
  XOR2_X1    g03926(.A1(new_n4119_), .A2(new_n4107_), .Z(new_n4120_));
  NAND2_X1   g03927(.A1(new_n3994_), .A2(new_n4002_), .ZN(new_n4121_));
  NAND2_X1   g03928(.A1(new_n4003_), .A2(new_n3990_), .ZN(new_n4122_));
  NAND2_X1   g03929(.A1(new_n4122_), .A2(new_n4121_), .ZN(new_n4123_));
  NAND2_X1   g03930(.A1(new_n4027_), .A2(new_n4060_), .ZN(new_n4124_));
  NAND2_X1   g03931(.A1(new_n4064_), .A2(new_n4061_), .ZN(new_n4125_));
  NAND2_X1   g03932(.A1(new_n4125_), .A2(new_n4124_), .ZN(new_n4126_));
  XOR2_X1    g03933(.A1(new_n4123_), .A2(new_n4126_), .Z(new_n4127_));
  XOR2_X1    g03934(.A1(new_n4127_), .A2(new_n4120_), .Z(new_n4128_));
  NOR2_X1    g03935(.A1(new_n4082_), .A2(new_n4128_), .ZN(new_n4129_));
  NAND2_X1   g03936(.A1(new_n4082_), .A2(new_n4128_), .ZN(new_n4130_));
  INV_X1     g03937(.I(new_n4130_), .ZN(new_n4131_));
  NOR2_X1    g03938(.A1(new_n4131_), .A2(new_n4129_), .ZN(new_n4132_));
  NOR2_X1    g03939(.A1(new_n4079_), .A2(new_n4132_), .ZN(new_n4133_));
  NAND2_X1   g03940(.A1(new_n4079_), .A2(new_n4132_), .ZN(new_n4134_));
  INV_X1     g03941(.I(new_n4134_), .ZN(new_n4135_));
  NOR2_X1    g03942(.A1(new_n4135_), .A2(new_n4133_), .ZN(new_n4136_));
  INV_X1     g03943(.I(new_n4136_), .ZN(new_n4137_));
  NAND2_X1   g03944(.A1(new_n3940_), .A2(new_n3949_), .ZN(new_n4138_));
  NAND2_X1   g03945(.A1(new_n3950_), .A2(new_n3961_), .ZN(new_n4139_));
  NAND2_X1   g03946(.A1(new_n4139_), .A2(new_n4138_), .ZN(new_n4140_));
  NAND2_X1   g03947(.A1(new_n4016_), .A2(new_n3827_), .ZN(new_n4141_));
  INV_X1     g03948(.I(new_n4026_), .ZN(new_n4142_));
  OAI21_X1   g03949(.A1(new_n4017_), .A2(new_n4142_), .B(new_n4141_), .ZN(new_n4143_));
  NAND2_X1   g03950(.A1(new_n4040_), .A2(new_n4048_), .ZN(new_n4144_));
  OAI21_X1   g03951(.A1(new_n4049_), .A2(new_n4059_), .B(new_n4144_), .ZN(new_n4145_));
  NOR2_X1    g03952(.A1(new_n4143_), .A2(new_n4145_), .ZN(new_n4146_));
  NAND2_X1   g03953(.A1(new_n4143_), .A2(new_n4145_), .ZN(new_n4147_));
  INV_X1     g03954(.I(new_n4147_), .ZN(new_n4148_));
  NOR2_X1    g03955(.A1(new_n4148_), .A2(new_n4146_), .ZN(new_n4149_));
  NOR2_X1    g03956(.A1(new_n4149_), .A2(new_n4140_), .ZN(new_n4150_));
  NAND2_X1   g03957(.A1(new_n4149_), .A2(new_n4140_), .ZN(new_n4151_));
  INV_X1     g03958(.I(new_n4151_), .ZN(new_n4152_));
  NOR2_X1    g03959(.A1(new_n4152_), .A2(new_n4150_), .ZN(new_n4153_));
  NAND2_X1   g03960(.A1(new_n3966_), .A2(new_n3971_), .ZN(new_n4154_));
  NAND2_X1   g03961(.A1(new_n3972_), .A2(new_n3963_), .ZN(new_n4155_));
  NAND2_X1   g03962(.A1(new_n4155_), .A2(new_n4154_), .ZN(new_n4156_));
  XOR2_X1    g03963(.A1(new_n4039_), .A2(new_n4024_), .Z(new_n4157_));
  XNOR2_X1   g03964(.A1(new_n4157_), .A2(new_n4047_), .ZN(new_n4158_));
  NOR2_X1    g03965(.A1(new_n3864_), .A2(new_n3783_), .ZN(new_n4159_));
  NOR2_X1    g03966(.A1(new_n3969_), .A2(new_n4159_), .ZN(new_n4160_));
  NAND2_X1   g03967(.A1(\a[1] ), .A2(\a[45] ), .ZN(new_n4161_));
  XOR2_X1    g03968(.A1(new_n1879_), .A2(new_n4161_), .Z(new_n4162_));
  XOR2_X1    g03969(.A1(new_n4162_), .A2(new_n3953_), .Z(new_n4163_));
  OR2_X2     g03970(.A1(new_n4163_), .A2(new_n4056_), .Z(new_n4164_));
  NAND2_X1   g03971(.A1(new_n4163_), .A2(new_n4056_), .ZN(new_n4165_));
  NAND2_X1   g03972(.A1(new_n4164_), .A2(new_n4165_), .ZN(new_n4166_));
  XNOR2_X1   g03973(.A1(new_n4160_), .A2(new_n4166_), .ZN(new_n4167_));
  XOR2_X1    g03974(.A1(new_n4167_), .A2(new_n4158_), .Z(new_n4168_));
  XOR2_X1    g03975(.A1(new_n4156_), .A2(new_n4168_), .Z(new_n4169_));
  XNOR2_X1   g03976(.A1(new_n4169_), .A2(new_n4153_), .ZN(new_n4170_));
  NAND2_X1   g03977(.A1(new_n3927_), .A2(new_n3973_), .ZN(new_n4171_));
  NAND2_X1   g03978(.A1(new_n3923_), .A2(new_n3926_), .ZN(new_n4172_));
  NAND2_X1   g03979(.A1(new_n4171_), .A2(new_n4172_), .ZN(new_n4173_));
  NAND2_X1   g03980(.A1(new_n3985_), .A2(new_n3988_), .ZN(new_n4174_));
  NAND2_X1   g03981(.A1(new_n3989_), .A2(new_n3981_), .ZN(new_n4175_));
  NAND2_X1   g03982(.A1(new_n4175_), .A2(new_n4174_), .ZN(new_n4176_));
  NAND4_X1   g03983(.A1(\a[0] ), .A2(\a[4] ), .A3(\a[42] ), .A4(\a[46] ), .ZN(new_n4177_));
  INV_X1     g03984(.I(\a[46] ), .ZN(new_n4178_));
  NOR4_X1    g03985(.A1(new_n196_), .A2(new_n225_), .A3(new_n3666_), .A4(new_n4178_), .ZN(new_n4179_));
  NOR2_X1    g03986(.A1(new_n3746_), .A2(new_n3666_), .ZN(new_n4180_));
  INV_X1     g03987(.I(new_n4180_), .ZN(new_n4181_));
  NOR2_X1    g03988(.A1(new_n4181_), .A2(new_n370_), .ZN(new_n4182_));
  OAI21_X1   g03989(.A1(new_n4182_), .A2(new_n4179_), .B(new_n4177_), .ZN(new_n4183_));
  NAND3_X1   g03990(.A1(new_n4183_), .A2(\a[3] ), .A3(\a[43] ), .ZN(new_n4184_));
  NAND2_X1   g03991(.A1(new_n4183_), .A2(new_n4177_), .ZN(new_n4185_));
  AOI22_X1   g03992(.A1(\a[0] ), .A2(\a[46] ), .B1(\a[4] ), .B2(\a[42] ), .ZN(new_n4186_));
  OAI21_X1   g03993(.A1(new_n4185_), .A2(new_n4186_), .B(new_n4184_), .ZN(new_n4187_));
  NAND2_X1   g03994(.A1(new_n747_), .A2(new_n3232_), .ZN(new_n4188_));
  NOR2_X1    g03995(.A1(new_n2524_), .A2(new_n2752_), .ZN(new_n4189_));
  INV_X1     g03996(.I(new_n4189_), .ZN(new_n4190_));
  OAI22_X1   g03997(.A1(new_n539_), .A2(new_n3038_), .B1(new_n4190_), .B2(new_n1063_), .ZN(new_n4191_));
  NAND2_X1   g03998(.A1(new_n4191_), .A2(new_n4188_), .ZN(new_n4192_));
  NAND3_X1   g03999(.A1(new_n4192_), .A2(\a[9] ), .A3(\a[37] ), .ZN(new_n4193_));
  AOI22_X1   g04000(.A1(\a[10] ), .A2(\a[36] ), .B1(\a[11] ), .B2(\a[35] ), .ZN(new_n4194_));
  NAND2_X1   g04001(.A1(new_n4192_), .A2(new_n4188_), .ZN(new_n4195_));
  OAI21_X1   g04002(.A1(new_n4194_), .A2(new_n4195_), .B(new_n4193_), .ZN(new_n4196_));
  XNOR2_X1   g04003(.A1(new_n4196_), .A2(new_n4187_), .ZN(new_n4197_));
  OAI22_X1   g04004(.A1(new_n1376_), .A2(new_n1972_), .B1(new_n1379_), .B2(new_n4010_), .ZN(new_n4198_));
  OAI21_X1   g04005(.A1(new_n1382_), .A2(new_n2177_), .B(new_n4198_), .ZN(new_n4199_));
  NAND3_X1   g04006(.A1(new_n4199_), .A2(\a[19] ), .A3(\a[27] ), .ZN(new_n4200_));
  AOI22_X1   g04007(.A1(\a[20] ), .A2(\a[26] ), .B1(\a[21] ), .B2(\a[25] ), .ZN(new_n4201_));
  NOR2_X1    g04008(.A1(new_n1382_), .A2(new_n2177_), .ZN(new_n4202_));
  NOR2_X1    g04009(.A1(new_n4198_), .A2(new_n4202_), .ZN(new_n4203_));
  INV_X1     g04010(.I(new_n4203_), .ZN(new_n4204_));
  OAI21_X1   g04011(.A1(new_n4201_), .A2(new_n4204_), .B(new_n4200_), .ZN(new_n4205_));
  XOR2_X1    g04012(.A1(new_n4197_), .A2(new_n4205_), .Z(new_n4206_));
  INV_X1     g04013(.I(new_n2890_), .ZN(new_n4207_));
  AOI22_X1   g04014(.A1(\a[7] ), .A2(\a[39] ), .B1(\a[8] ), .B2(\a[38] ), .ZN(new_n4208_));
  NOR2_X1    g04015(.A1(new_n2914_), .A2(new_n3116_), .ZN(new_n4209_));
  INV_X1     g04016(.I(new_n4209_), .ZN(new_n4210_));
  NOR2_X1    g04017(.A1(new_n4210_), .A2(new_n415_), .ZN(new_n4211_));
  NOR3_X1    g04018(.A1(new_n4211_), .A2(new_n4207_), .A3(new_n4208_), .ZN(new_n4212_));
  NOR2_X1    g04019(.A1(new_n4212_), .A2(new_n4211_), .ZN(new_n4213_));
  INV_X1     g04020(.I(new_n4213_), .ZN(new_n4214_));
  OAI22_X1   g04021(.A1(new_n4214_), .A2(new_n4208_), .B1(new_n4207_), .B2(new_n4212_), .ZN(new_n4215_));
  NAND2_X1   g04022(.A1(new_n1027_), .A2(new_n2105_), .ZN(new_n4216_));
  OAI22_X1   g04023(.A1(new_n1428_), .A2(new_n2255_), .B1(new_n1429_), .B2(new_n3811_), .ZN(new_n4217_));
  NAND2_X1   g04024(.A1(new_n4217_), .A2(new_n4216_), .ZN(new_n4218_));
  NOR2_X1    g04025(.A1(new_n742_), .A2(new_n2030_), .ZN(new_n4219_));
  AOI22_X1   g04026(.A1(\a[17] ), .A2(\a[29] ), .B1(\a[18] ), .B2(\a[28] ), .ZN(new_n4220_));
  NAND2_X1   g04027(.A1(new_n4218_), .A2(new_n4216_), .ZN(new_n4221_));
  NOR2_X1    g04028(.A1(new_n4221_), .A2(new_n4220_), .ZN(new_n4222_));
  AOI21_X1   g04029(.A1(new_n4218_), .A2(new_n4219_), .B(new_n4222_), .ZN(new_n4223_));
  XNOR2_X1   g04030(.A1(new_n4223_), .A2(new_n3959_), .ZN(new_n4224_));
  XNOR2_X1   g04031(.A1(new_n4224_), .A2(new_n4215_), .ZN(new_n4225_));
  XOR2_X1    g04032(.A1(new_n4225_), .A2(new_n4206_), .Z(new_n4226_));
  INV_X1     g04033(.I(new_n4226_), .ZN(new_n4227_));
  XOR2_X1    g04034(.A1(new_n4176_), .A2(new_n4227_), .Z(new_n4228_));
  XOR2_X1    g04035(.A1(new_n4173_), .A2(new_n4228_), .Z(new_n4229_));
  INV_X1     g04036(.I(new_n4229_), .ZN(new_n4230_));
  OR2_X2     g04037(.A1(new_n4230_), .A2(new_n4170_), .Z(new_n4231_));
  NAND2_X1   g04038(.A1(new_n4230_), .A2(new_n4170_), .ZN(new_n4232_));
  AND2_X2    g04039(.A1(new_n4231_), .A2(new_n4232_), .Z(new_n4233_));
  INV_X1     g04040(.I(new_n4233_), .ZN(new_n4234_));
  NOR2_X1    g04041(.A1(new_n4137_), .A2(new_n4234_), .ZN(new_n4235_));
  INV_X1     g04042(.I(new_n4235_), .ZN(new_n4236_));
  NOR2_X1    g04043(.A1(new_n4136_), .A2(new_n4233_), .ZN(new_n4237_));
  INV_X1     g04044(.I(new_n4237_), .ZN(new_n4238_));
  NAND2_X1   g04045(.A1(new_n4236_), .A2(new_n4238_), .ZN(new_n4239_));
  XOR2_X1    g04046(.A1(new_n4076_), .A2(new_n4239_), .Z(\asquared[47] ));
  OAI21_X1   g04047(.A1(new_n4075_), .A2(new_n4072_), .B(new_n4238_), .ZN(new_n4241_));
  NAND2_X1   g04048(.A1(new_n4241_), .A2(new_n4236_), .ZN(new_n4242_));
  NOR2_X1    g04049(.A1(new_n4135_), .A2(new_n4131_), .ZN(new_n4243_));
  NAND2_X1   g04050(.A1(new_n4123_), .A2(new_n4126_), .ZN(new_n4244_));
  NAND2_X1   g04051(.A1(new_n4127_), .A2(new_n4120_), .ZN(new_n4245_));
  NAND2_X1   g04052(.A1(new_n4245_), .A2(new_n4244_), .ZN(new_n4246_));
  NAND2_X1   g04053(.A1(new_n4156_), .A2(new_n4168_), .ZN(new_n4247_));
  NAND2_X1   g04054(.A1(new_n4169_), .A2(new_n4153_), .ZN(new_n4248_));
  NAND2_X1   g04055(.A1(new_n4248_), .A2(new_n4247_), .ZN(new_n4249_));
  XOR2_X1    g04056(.A1(new_n4246_), .A2(new_n4249_), .Z(new_n4250_));
  NAND2_X1   g04057(.A1(new_n4105_), .A2(new_n4093_), .ZN(new_n4251_));
  NAND2_X1   g04058(.A1(new_n4106_), .A2(new_n4085_), .ZN(new_n4252_));
  NAND2_X1   g04059(.A1(new_n4252_), .A2(new_n4251_), .ZN(new_n4253_));
  NAND2_X1   g04060(.A1(new_n4196_), .A2(new_n4187_), .ZN(new_n4254_));
  INV_X1     g04061(.I(new_n4197_), .ZN(new_n4255_));
  NAND2_X1   g04062(.A1(new_n4255_), .A2(new_n4205_), .ZN(new_n4256_));
  NAND2_X1   g04063(.A1(new_n4256_), .A2(new_n4254_), .ZN(new_n4257_));
  XOR2_X1    g04064(.A1(new_n4203_), .A2(new_n4089_), .Z(new_n4258_));
  XOR2_X1    g04065(.A1(new_n4258_), .A2(new_n4185_), .Z(new_n4259_));
  XOR2_X1    g04066(.A1(new_n4257_), .A2(new_n4259_), .Z(new_n4260_));
  XOR2_X1    g04067(.A1(new_n4260_), .A2(new_n4253_), .Z(new_n4261_));
  NAND2_X1   g04068(.A1(new_n4110_), .A2(new_n4118_), .ZN(new_n4262_));
  NAND2_X1   g04069(.A1(new_n4119_), .A2(new_n4107_), .ZN(new_n4263_));
  NAND2_X1   g04070(.A1(new_n4263_), .A2(new_n4262_), .ZN(new_n4264_));
  NAND2_X1   g04071(.A1(new_n4176_), .A2(new_n4227_), .ZN(new_n4265_));
  INV_X1     g04072(.I(new_n4206_), .ZN(new_n4266_));
  NAND2_X1   g04073(.A1(new_n4225_), .A2(new_n4266_), .ZN(new_n4267_));
  NAND2_X1   g04074(.A1(new_n4265_), .A2(new_n4267_), .ZN(new_n4268_));
  XNOR2_X1   g04075(.A1(new_n4264_), .A2(new_n4268_), .ZN(new_n4269_));
  XNOR2_X1   g04076(.A1(new_n4269_), .A2(new_n4261_), .ZN(new_n4270_));
  XOR2_X1    g04077(.A1(new_n4250_), .A2(new_n4270_), .Z(new_n4271_));
  NAND2_X1   g04078(.A1(new_n4173_), .A2(new_n4228_), .ZN(new_n4272_));
  NAND2_X1   g04079(.A1(new_n4231_), .A2(new_n4272_), .ZN(new_n4273_));
  NOR2_X1    g04080(.A1(new_n4152_), .A2(new_n4148_), .ZN(new_n4274_));
  OAI21_X1   g04081(.A1(new_n3954_), .A2(new_n4162_), .B(new_n4164_), .ZN(new_n4275_));
  NOR2_X1    g04082(.A1(new_n536_), .A2(new_n3221_), .ZN(new_n4276_));
  NAND2_X1   g04083(.A1(new_n3588_), .A2(new_n4276_), .ZN(new_n4277_));
  NAND4_X1   g04084(.A1(\a[7] ), .A2(\a[13] ), .A3(\a[34] ), .A4(\a[40] ), .ZN(new_n4278_));
  OAI21_X1   g04085(.A1(new_n1265_), .A2(new_n2746_), .B(new_n4278_), .ZN(new_n4279_));
  NAND2_X1   g04086(.A1(new_n4279_), .A2(new_n4277_), .ZN(new_n4280_));
  NAND3_X1   g04087(.A1(new_n4280_), .A2(\a[13] ), .A3(\a[34] ), .ZN(new_n4281_));
  AOI22_X1   g04088(.A1(\a[7] ), .A2(\a[40] ), .B1(\a[12] ), .B2(\a[35] ), .ZN(new_n4282_));
  NAND2_X1   g04089(.A1(new_n4280_), .A2(new_n4277_), .ZN(new_n4283_));
  OAI21_X1   g04090(.A1(new_n4282_), .A2(new_n4283_), .B(new_n4281_), .ZN(new_n4284_));
  XOR2_X1    g04091(.A1(new_n4275_), .A2(new_n4284_), .Z(new_n4285_));
  OAI21_X1   g04092(.A1(new_n4113_), .A2(new_n4117_), .B(new_n4285_), .ZN(new_n4286_));
  OR3_X2     g04093(.A1(new_n4285_), .A2(new_n4113_), .A3(new_n4117_), .Z(new_n4287_));
  NAND2_X1   g04094(.A1(new_n4287_), .A2(new_n4286_), .ZN(new_n4288_));
  NOR2_X1    g04095(.A1(new_n4160_), .A2(new_n4166_), .ZN(new_n4289_));
  NOR2_X1    g04096(.A1(new_n4167_), .A2(new_n4158_), .ZN(new_n4290_));
  NOR2_X1    g04097(.A1(new_n4290_), .A2(new_n4289_), .ZN(new_n4291_));
  XOR2_X1    g04098(.A1(new_n4291_), .A2(new_n4288_), .Z(new_n4292_));
  XNOR2_X1   g04099(.A1(new_n4292_), .A2(new_n4274_), .ZN(new_n4293_));
  INV_X1     g04100(.I(new_n4224_), .ZN(new_n4294_));
  NAND2_X1   g04101(.A1(new_n4294_), .A2(new_n4215_), .ZN(new_n4295_));
  OAI21_X1   g04102(.A1(new_n3959_), .A2(new_n4223_), .B(new_n4295_), .ZN(new_n4296_));
  NAND2_X1   g04103(.A1(new_n4039_), .A2(new_n4024_), .ZN(new_n4297_));
  NAND2_X1   g04104(.A1(new_n4157_), .A2(new_n4047_), .ZN(new_n4298_));
  NAND2_X1   g04105(.A1(new_n4298_), .A2(new_n4297_), .ZN(new_n4299_));
  XOR2_X1    g04106(.A1(new_n4296_), .A2(new_n4299_), .Z(new_n4300_));
  NOR3_X1    g04107(.A1(new_n194_), .A2(new_n1357_), .A3(new_n4178_), .ZN(new_n4301_));
  INV_X1     g04108(.I(new_n4301_), .ZN(new_n4302_));
  NOR2_X1    g04109(.A1(new_n194_), .A2(new_n4178_), .ZN(new_n4303_));
  OAI21_X1   g04110(.A1(new_n4303_), .A2(\a[24] ), .B(new_n4302_), .ZN(new_n4304_));
  XOR2_X1    g04111(.A1(new_n4195_), .A2(new_n4304_), .Z(new_n4305_));
  XOR2_X1    g04112(.A1(new_n4305_), .A2(new_n4214_), .Z(new_n4306_));
  INV_X1     g04113(.I(new_n4306_), .ZN(new_n4307_));
  XOR2_X1    g04114(.A1(new_n4300_), .A2(new_n4307_), .Z(new_n4308_));
  AOI22_X1   g04115(.A1(\a[0] ), .A2(\a[47] ), .B1(\a[2] ), .B2(\a[45] ), .ZN(new_n4309_));
  NOR2_X1    g04116(.A1(new_n1880_), .A2(new_n4161_), .ZN(new_n4310_));
  INV_X1     g04117(.I(new_n4309_), .ZN(new_n4311_));
  INV_X1     g04118(.I(\a[47] ), .ZN(new_n4312_));
  NOR2_X1    g04119(.A1(new_n4030_), .A2(new_n4312_), .ZN(new_n4313_));
  INV_X1     g04120(.I(new_n4313_), .ZN(new_n4314_));
  NOR2_X1    g04121(.A1(new_n4314_), .A2(new_n412_), .ZN(new_n4315_));
  AOI21_X1   g04122(.A1(new_n4310_), .A2(new_n4311_), .B(new_n4315_), .ZN(new_n4316_));
  INV_X1     g04123(.I(new_n4316_), .ZN(new_n4317_));
  OAI21_X1   g04124(.A1(new_n4309_), .A2(new_n4315_), .B(new_n4310_), .ZN(new_n4318_));
  OAI21_X1   g04125(.A1(new_n4317_), .A2(new_n4309_), .B(new_n4318_), .ZN(new_n4319_));
  NAND2_X1   g04126(.A1(new_n1024_), .A2(new_n2437_), .ZN(new_n4320_));
  NAND2_X1   g04127(.A1(new_n1025_), .A2(new_n2976_), .ZN(new_n4321_));
  AOI22_X1   g04128(.A1(new_n4320_), .A2(new_n4321_), .B1(new_n1027_), .B2(new_n2254_), .ZN(new_n4322_));
  NOR3_X1    g04129(.A1(new_n4322_), .A2(new_n742_), .A3(new_n2051_), .ZN(new_n4323_));
  AOI22_X1   g04130(.A1(\a[17] ), .A2(\a[30] ), .B1(\a[18] ), .B2(\a[29] ), .ZN(new_n4324_));
  NAND2_X1   g04131(.A1(new_n1027_), .A2(new_n2254_), .ZN(new_n4325_));
  NAND3_X1   g04132(.A1(new_n4325_), .A2(new_n4320_), .A3(new_n4321_), .ZN(new_n4326_));
  NOR2_X1    g04133(.A1(new_n4326_), .A2(new_n4324_), .ZN(new_n4327_));
  NOR2_X1    g04134(.A1(new_n4323_), .A2(new_n4327_), .ZN(new_n4328_));
  XOR2_X1    g04135(.A1(new_n4319_), .A2(new_n4328_), .Z(new_n4329_));
  NAND2_X1   g04136(.A1(new_n1375_), .A2(new_n2103_), .ZN(new_n4330_));
  NAND2_X1   g04137(.A1(new_n1378_), .A2(new_n2412_), .ZN(new_n4331_));
  AOI22_X1   g04138(.A1(new_n4330_), .A2(new_n4331_), .B1(new_n1381_), .B2(new_n1971_), .ZN(new_n4332_));
  NAND2_X1   g04139(.A1(\a[19] ), .A2(\a[28] ), .ZN(new_n4333_));
  AOI22_X1   g04140(.A1(\a[20] ), .A2(\a[27] ), .B1(\a[21] ), .B2(\a[26] ), .ZN(new_n4334_));
  NAND2_X1   g04141(.A1(new_n1381_), .A2(new_n1971_), .ZN(new_n4335_));
  NAND3_X1   g04142(.A1(new_n4335_), .A2(new_n4330_), .A3(new_n4331_), .ZN(new_n4336_));
  OAI22_X1   g04143(.A1(new_n4332_), .A2(new_n4333_), .B1(new_n4336_), .B2(new_n4334_), .ZN(new_n4337_));
  XNOR2_X1   g04144(.A1(new_n4329_), .A2(new_n4337_), .ZN(new_n4338_));
  XNOR2_X1   g04145(.A1(new_n4102_), .A2(new_n4221_), .ZN(new_n4339_));
  NAND4_X1   g04146(.A1(\a[4] ), .A2(\a[15] ), .A3(\a[32] ), .A4(\a[43] ), .ZN(new_n4340_));
  NAND3_X1   g04147(.A1(new_n2516_), .A2(\a[15] ), .A3(\a[44] ), .ZN(new_n4341_));
  NOR2_X1    g04148(.A1(new_n3666_), .A2(new_n3859_), .ZN(new_n4342_));
  INV_X1     g04149(.I(new_n4342_), .ZN(new_n4343_));
  OAI21_X1   g04150(.A1(new_n370_), .A2(new_n4343_), .B(new_n4341_), .ZN(new_n4344_));
  NAND2_X1   g04151(.A1(new_n4344_), .A2(new_n4340_), .ZN(new_n4345_));
  NAND3_X1   g04152(.A1(new_n4345_), .A2(\a[3] ), .A3(\a[44] ), .ZN(new_n4346_));
  NAND2_X1   g04153(.A1(new_n4345_), .A2(new_n4340_), .ZN(new_n4347_));
  AOI22_X1   g04154(.A1(\a[4] ), .A2(\a[43] ), .B1(\a[15] ), .B2(\a[32] ), .ZN(new_n4348_));
  OAI21_X1   g04155(.A1(new_n4347_), .A2(new_n4348_), .B(new_n4346_), .ZN(new_n4349_));
  XOR2_X1    g04156(.A1(new_n4339_), .A2(new_n4349_), .Z(new_n4350_));
  NOR2_X1    g04157(.A1(new_n1175_), .A2(new_n1441_), .ZN(new_n4351_));
  NOR2_X1    g04158(.A1(new_n1528_), .A2(new_n4351_), .ZN(new_n4352_));
  INV_X1     g04159(.I(new_n4352_), .ZN(new_n4353_));
  NOR2_X1    g04160(.A1(new_n2385_), .A2(new_n1779_), .ZN(new_n4354_));
  NOR2_X1    g04161(.A1(new_n417_), .A2(new_n2752_), .ZN(new_n4355_));
  AOI21_X1   g04162(.A1(new_n4353_), .A2(new_n4355_), .B(new_n4354_), .ZN(new_n4356_));
  INV_X1     g04163(.I(new_n4356_), .ZN(new_n4357_));
  OAI21_X1   g04164(.A1(new_n4354_), .A2(new_n4352_), .B(new_n4355_), .ZN(new_n4358_));
  OAI21_X1   g04165(.A1(new_n4357_), .A2(new_n4352_), .B(new_n4358_), .ZN(new_n4359_));
  NOR2_X1    g04166(.A1(new_n2916_), .A2(new_n1063_), .ZN(new_n4360_));
  INV_X1     g04167(.I(new_n4360_), .ZN(new_n4361_));
  NOR3_X1    g04168(.A1(new_n3820_), .A2(new_n513_), .A3(new_n3116_), .ZN(new_n4362_));
  NOR2_X1    g04169(.A1(new_n4210_), .A2(new_n1427_), .ZN(new_n4363_));
  OAI21_X1   g04170(.A1(new_n4362_), .A2(new_n4363_), .B(new_n4361_), .ZN(new_n4364_));
  NAND3_X1   g04171(.A1(new_n4364_), .A2(\a[8] ), .A3(\a[39] ), .ZN(new_n4365_));
  AOI22_X1   g04172(.A1(\a[9] ), .A2(\a[38] ), .B1(\a[11] ), .B2(\a[36] ), .ZN(new_n4366_));
  NAND2_X1   g04173(.A1(new_n4364_), .A2(new_n4361_), .ZN(new_n4367_));
  OAI21_X1   g04174(.A1(new_n4366_), .A2(new_n4367_), .B(new_n4365_), .ZN(new_n4368_));
  XOR2_X1    g04175(.A1(new_n4368_), .A2(new_n4359_), .Z(new_n4369_));
  NOR2_X1    g04176(.A1(new_n2274_), .A2(new_n3327_), .ZN(new_n4370_));
  NAND3_X1   g04177(.A1(new_n2966_), .A2(\a[14] ), .A3(\a[42] ), .ZN(new_n4371_));
  NOR2_X1    g04178(.A1(new_n3327_), .A2(new_n3746_), .ZN(new_n4372_));
  NAND2_X1   g04179(.A1(new_n4372_), .A2(new_n746_), .ZN(new_n4373_));
  AOI22_X1   g04180(.A1(new_n4371_), .A2(new_n4373_), .B1(new_n1053_), .B2(new_n4370_), .ZN(new_n4374_));
  NAND2_X1   g04181(.A1(\a[5] ), .A2(\a[42] ), .ZN(new_n4375_));
  AOI22_X1   g04182(.A1(\a[6] ), .A2(\a[41] ), .B1(\a[14] ), .B2(\a[33] ), .ZN(new_n4376_));
  NAND2_X1   g04183(.A1(new_n1053_), .A2(new_n4370_), .ZN(new_n4377_));
  NAND3_X1   g04184(.A1(new_n4377_), .A2(new_n4371_), .A3(new_n4373_), .ZN(new_n4378_));
  OAI22_X1   g04185(.A1(new_n4374_), .A2(new_n4375_), .B1(new_n4378_), .B2(new_n4376_), .ZN(new_n4379_));
  XOR2_X1    g04186(.A1(new_n4369_), .A2(new_n4379_), .Z(new_n4380_));
  XOR2_X1    g04187(.A1(new_n4380_), .A2(new_n4350_), .Z(new_n4381_));
  XOR2_X1    g04188(.A1(new_n4381_), .A2(new_n4338_), .Z(new_n4382_));
  NAND2_X1   g04189(.A1(new_n4308_), .A2(new_n4382_), .ZN(new_n4383_));
  NAND2_X1   g04190(.A1(new_n4383_), .A2(new_n4308_), .ZN(new_n4384_));
  NAND2_X1   g04191(.A1(new_n4383_), .A2(new_n4382_), .ZN(new_n4385_));
  NAND2_X1   g04192(.A1(new_n4385_), .A2(new_n4384_), .ZN(new_n4386_));
  AOI21_X1   g04193(.A1(new_n4382_), .A2(new_n4383_), .B(new_n4293_), .ZN(new_n4387_));
  AOI22_X1   g04194(.A1(new_n4387_), .A2(new_n4384_), .B1(new_n4386_), .B2(new_n4293_), .ZN(new_n4388_));
  INV_X1     g04195(.I(new_n4388_), .ZN(new_n4389_));
  NOR2_X1    g04196(.A1(new_n4273_), .A2(new_n4389_), .ZN(new_n4390_));
  INV_X1     g04197(.I(new_n4390_), .ZN(new_n4391_));
  NAND2_X1   g04198(.A1(new_n4273_), .A2(new_n4389_), .ZN(new_n4392_));
  NAND2_X1   g04199(.A1(new_n4391_), .A2(new_n4392_), .ZN(new_n4393_));
  INV_X1     g04200(.I(new_n4392_), .ZN(new_n4394_));
  NOR2_X1    g04201(.A1(new_n4394_), .A2(new_n4271_), .ZN(new_n4395_));
  AOI22_X1   g04202(.A1(new_n4395_), .A2(new_n4391_), .B1(new_n4393_), .B2(new_n4271_), .ZN(new_n4396_));
  INV_X1     g04203(.I(new_n4396_), .ZN(new_n4397_));
  NOR2_X1    g04204(.A1(new_n4397_), .A2(new_n4243_), .ZN(new_n4398_));
  NAND2_X1   g04205(.A1(new_n4397_), .A2(new_n4243_), .ZN(new_n4399_));
  INV_X1     g04206(.I(new_n4399_), .ZN(new_n4400_));
  NOR2_X1    g04207(.A1(new_n4400_), .A2(new_n4398_), .ZN(new_n4401_));
  XOR2_X1    g04208(.A1(new_n4242_), .A2(new_n4401_), .Z(\asquared[48] ));
  NAND2_X1   g04209(.A1(new_n4273_), .A2(new_n4388_), .ZN(new_n4403_));
  NAND2_X1   g04210(.A1(new_n4393_), .A2(new_n4271_), .ZN(new_n4404_));
  NAND2_X1   g04211(.A1(new_n4404_), .A2(new_n4403_), .ZN(new_n4405_));
  INV_X1     g04212(.I(new_n4405_), .ZN(new_n4406_));
  XOR2_X1    g04213(.A1(new_n4347_), .A2(new_n4326_), .Z(new_n4407_));
  XOR2_X1    g04214(.A1(new_n4407_), .A2(new_n4317_), .Z(new_n4408_));
  INV_X1     g04215(.I(new_n4408_), .ZN(new_n4409_));
  INV_X1     g04216(.I(new_n4304_), .ZN(new_n4410_));
  NOR2_X1    g04217(.A1(new_n4305_), .A2(new_n4213_), .ZN(new_n4411_));
  AOI21_X1   g04218(.A1(new_n4195_), .A2(new_n4410_), .B(new_n4411_), .ZN(new_n4412_));
  INV_X1     g04219(.I(new_n4319_), .ZN(new_n4413_));
  INV_X1     g04220(.I(new_n4329_), .ZN(new_n4414_));
  NAND2_X1   g04221(.A1(new_n4414_), .A2(new_n4337_), .ZN(new_n4415_));
  OAI21_X1   g04222(.A1(new_n4413_), .A2(new_n4328_), .B(new_n4415_), .ZN(new_n4416_));
  XNOR2_X1   g04223(.A1(new_n4416_), .A2(new_n4412_), .ZN(new_n4417_));
  INV_X1     g04224(.I(new_n4417_), .ZN(new_n4418_));
  NOR2_X1    g04225(.A1(new_n4418_), .A2(new_n4409_), .ZN(new_n4419_));
  INV_X1     g04226(.I(new_n4419_), .ZN(new_n4420_));
  NAND2_X1   g04227(.A1(new_n4418_), .A2(new_n4409_), .ZN(new_n4421_));
  AND2_X2    g04228(.A1(new_n4420_), .A2(new_n4421_), .Z(new_n4422_));
  NAND2_X1   g04229(.A1(new_n4381_), .A2(new_n4338_), .ZN(new_n4423_));
  NAND2_X1   g04230(.A1(new_n4380_), .A2(new_n4350_), .ZN(new_n4424_));
  NAND2_X1   g04231(.A1(new_n4423_), .A2(new_n4424_), .ZN(new_n4425_));
  XNOR2_X1   g04232(.A1(new_n4283_), .A2(new_n4356_), .ZN(new_n4426_));
  NAND2_X1   g04233(.A1(\a[2] ), .A2(\a[16] ), .ZN(new_n4427_));
  NAND2_X1   g04234(.A1(\a[32] ), .A2(\a[46] ), .ZN(new_n4428_));
  NOR2_X1    g04235(.A1(new_n4030_), .A2(new_n4178_), .ZN(new_n4429_));
  INV_X1     g04236(.I(new_n4429_), .ZN(new_n4430_));
  OAI22_X1   g04237(.A1(new_n4430_), .A2(new_n246_), .B1(new_n4427_), .B2(new_n4428_), .ZN(new_n4431_));
  NAND4_X1   g04238(.A1(\a[3] ), .A2(\a[16] ), .A3(\a[32] ), .A4(\a[45] ), .ZN(new_n4432_));
  NAND2_X1   g04239(.A1(new_n4431_), .A2(new_n4432_), .ZN(new_n4433_));
  NAND3_X1   g04240(.A1(new_n4433_), .A2(\a[2] ), .A3(\a[46] ), .ZN(new_n4434_));
  AOI22_X1   g04241(.A1(\a[3] ), .A2(\a[45] ), .B1(\a[16] ), .B2(\a[32] ), .ZN(new_n4435_));
  NAND2_X1   g04242(.A1(new_n4433_), .A2(new_n4432_), .ZN(new_n4436_));
  OAI21_X1   g04243(.A1(new_n4435_), .A2(new_n4436_), .B(new_n4434_), .ZN(new_n4437_));
  XNOR2_X1   g04244(.A1(new_n4426_), .A2(new_n4437_), .ZN(new_n4438_));
  INV_X1     g04245(.I(new_n4438_), .ZN(new_n4439_));
  XOR2_X1    g04246(.A1(new_n4367_), .A2(new_n4336_), .Z(new_n4440_));
  XOR2_X1    g04247(.A1(new_n4440_), .A2(new_n4378_), .Z(new_n4441_));
  NAND2_X1   g04248(.A1(new_n4368_), .A2(new_n4359_), .ZN(new_n4442_));
  NAND2_X1   g04249(.A1(new_n4369_), .A2(new_n4379_), .ZN(new_n4443_));
  NAND2_X1   g04250(.A1(new_n4443_), .A2(new_n4442_), .ZN(new_n4444_));
  XOR2_X1    g04251(.A1(new_n4444_), .A2(new_n4441_), .Z(new_n4445_));
  XOR2_X1    g04252(.A1(new_n4445_), .A2(new_n4439_), .Z(new_n4446_));
  XOR2_X1    g04253(.A1(new_n4425_), .A2(new_n4446_), .Z(new_n4447_));
  OR2_X2     g04254(.A1(new_n4447_), .A2(new_n4422_), .Z(new_n4448_));
  NAND2_X1   g04255(.A1(new_n4447_), .A2(new_n4422_), .ZN(new_n4449_));
  AND2_X2    g04256(.A1(new_n4448_), .A2(new_n4449_), .Z(new_n4450_));
  NAND2_X1   g04257(.A1(new_n4386_), .A2(new_n4293_), .ZN(new_n4451_));
  NAND2_X1   g04258(.A1(new_n4451_), .A2(new_n4383_), .ZN(new_n4452_));
  NAND2_X1   g04259(.A1(new_n4103_), .A2(new_n4221_), .ZN(new_n4453_));
  NAND2_X1   g04260(.A1(new_n4339_), .A2(new_n4349_), .ZN(new_n4454_));
  NAND2_X1   g04261(.A1(new_n4454_), .A2(new_n4453_), .ZN(new_n4455_));
  NAND2_X1   g04262(.A1(new_n4258_), .A2(new_n4185_), .ZN(new_n4456_));
  OAI21_X1   g04263(.A1(new_n4089_), .A2(new_n4203_), .B(new_n4456_), .ZN(new_n4457_));
  NAND2_X1   g04264(.A1(\a[0] ), .A2(\a[48] ), .ZN(new_n4458_));
  XOR2_X1    g04265(.A1(new_n4301_), .A2(new_n4458_), .Z(new_n4459_));
  NAND2_X1   g04266(.A1(\a[1] ), .A2(\a[47] ), .ZN(new_n4460_));
  XOR2_X1    g04267(.A1(new_n1442_), .A2(new_n4460_), .Z(new_n4461_));
  XNOR2_X1   g04268(.A1(new_n4459_), .A2(new_n4461_), .ZN(new_n4462_));
  INV_X1     g04269(.I(new_n4462_), .ZN(new_n4463_));
  XOR2_X1    g04270(.A1(new_n4457_), .A2(new_n4463_), .Z(new_n4464_));
  XOR2_X1    g04271(.A1(new_n4464_), .A2(new_n4455_), .Z(new_n4465_));
  NAND2_X1   g04272(.A1(new_n4257_), .A2(new_n4259_), .ZN(new_n4466_));
  NAND2_X1   g04273(.A1(new_n4260_), .A2(new_n4253_), .ZN(new_n4467_));
  NAND2_X1   g04274(.A1(new_n4467_), .A2(new_n4466_), .ZN(new_n4468_));
  NAND2_X1   g04275(.A1(new_n4296_), .A2(new_n4299_), .ZN(new_n4469_));
  NAND2_X1   g04276(.A1(new_n4300_), .A2(new_n4307_), .ZN(new_n4470_));
  NAND2_X1   g04277(.A1(new_n4470_), .A2(new_n4469_), .ZN(new_n4471_));
  XOR2_X1    g04278(.A1(new_n4471_), .A2(new_n4468_), .Z(new_n4472_));
  NAND2_X1   g04279(.A1(new_n4472_), .A2(new_n4465_), .ZN(new_n4473_));
  OR2_X2     g04280(.A1(new_n4472_), .A2(new_n4465_), .Z(new_n4474_));
  AND2_X2    g04281(.A1(new_n4474_), .A2(new_n4473_), .Z(new_n4475_));
  INV_X1     g04282(.I(new_n4475_), .ZN(new_n4476_));
  NAND2_X1   g04283(.A1(new_n4476_), .A2(new_n4452_), .ZN(new_n4477_));
  NOR2_X1    g04284(.A1(new_n4476_), .A2(new_n4452_), .ZN(new_n4478_));
  INV_X1     g04285(.I(new_n4478_), .ZN(new_n4479_));
  NAND2_X1   g04286(.A1(new_n4479_), .A2(new_n4477_), .ZN(new_n4480_));
  NAND2_X1   g04287(.A1(new_n4480_), .A2(new_n4450_), .ZN(new_n4481_));
  INV_X1     g04288(.I(new_n4450_), .ZN(new_n4482_));
  NAND3_X1   g04289(.A1(new_n4479_), .A2(new_n4482_), .A3(new_n4477_), .ZN(new_n4483_));
  NAND2_X1   g04290(.A1(new_n4481_), .A2(new_n4483_), .ZN(new_n4484_));
  NAND2_X1   g04291(.A1(new_n4246_), .A2(new_n4249_), .ZN(new_n4485_));
  NAND2_X1   g04292(.A1(new_n4250_), .A2(new_n4270_), .ZN(new_n4486_));
  NAND2_X1   g04293(.A1(new_n4264_), .A2(new_n4268_), .ZN(new_n4487_));
  INV_X1     g04294(.I(new_n4269_), .ZN(new_n4488_));
  NAND2_X1   g04295(.A1(new_n4488_), .A2(new_n4261_), .ZN(new_n4489_));
  NAND2_X1   g04296(.A1(new_n4489_), .A2(new_n4487_), .ZN(new_n4490_));
  NOR2_X1    g04297(.A1(new_n4291_), .A2(new_n4288_), .ZN(new_n4491_));
  INV_X1     g04298(.I(new_n4292_), .ZN(new_n4492_));
  NOR2_X1    g04299(.A1(new_n4492_), .A2(new_n4274_), .ZN(new_n4493_));
  NOR2_X1    g04300(.A1(new_n4493_), .A2(new_n4491_), .ZN(new_n4494_));
  NOR2_X1    g04301(.A1(new_n2274_), .A2(new_n3666_), .ZN(new_n4495_));
  NAND2_X1   g04302(.A1(new_n1054_), .A2(new_n4495_), .ZN(new_n4496_));
  NOR4_X1    g04303(.A1(new_n290_), .A2(new_n717_), .A3(new_n2274_), .A4(new_n3859_), .ZN(new_n4497_));
  NOR2_X1    g04304(.A1(new_n4343_), .A2(new_n242_), .ZN(new_n4498_));
  OAI21_X1   g04305(.A1(new_n4498_), .A2(new_n4497_), .B(new_n4496_), .ZN(new_n4499_));
  NAND3_X1   g04306(.A1(new_n4499_), .A2(\a[4] ), .A3(\a[44] ), .ZN(new_n4500_));
  NAND2_X1   g04307(.A1(new_n4499_), .A2(new_n4496_), .ZN(new_n4501_));
  AOI22_X1   g04308(.A1(\a[5] ), .A2(\a[43] ), .B1(\a[15] ), .B2(\a[33] ), .ZN(new_n4502_));
  OAI21_X1   g04309(.A1(new_n4501_), .A2(new_n4502_), .B(new_n4500_), .ZN(new_n4503_));
  NAND2_X1   g04310(.A1(new_n1452_), .A2(new_n1971_), .ZN(new_n4504_));
  OAI22_X1   g04311(.A1(new_n1382_), .A2(new_n2189_), .B1(new_n2647_), .B2(new_n3341_), .ZN(new_n4505_));
  NAND2_X1   g04312(.A1(new_n4505_), .A2(new_n4504_), .ZN(new_n4506_));
  NAND3_X1   g04313(.A1(new_n4506_), .A2(\a[20] ), .A3(\a[28] ), .ZN(new_n4507_));
  AOI22_X1   g04314(.A1(\a[21] ), .A2(\a[27] ), .B1(\a[22] ), .B2(\a[26] ), .ZN(new_n4508_));
  NAND2_X1   g04315(.A1(new_n4506_), .A2(new_n4504_), .ZN(new_n4509_));
  OAI21_X1   g04316(.A1(new_n4508_), .A2(new_n4509_), .B(new_n4507_), .ZN(new_n4510_));
  XNOR2_X1   g04317(.A1(new_n4510_), .A2(new_n4503_), .ZN(new_n4511_));
  NAND2_X1   g04318(.A1(new_n1027_), .A2(new_n2437_), .ZN(new_n4512_));
  NAND2_X1   g04319(.A1(new_n2629_), .A2(new_n2976_), .ZN(new_n4513_));
  AOI22_X1   g04320(.A1(new_n4512_), .A2(new_n4513_), .B1(new_n1194_), .B2(new_n2254_), .ZN(new_n4514_));
  NAND2_X1   g04321(.A1(\a[17] ), .A2(\a[31] ), .ZN(new_n4515_));
  AOI22_X1   g04322(.A1(\a[18] ), .A2(\a[30] ), .B1(\a[19] ), .B2(\a[29] ), .ZN(new_n4516_));
  NAND2_X1   g04323(.A1(new_n2254_), .A2(new_n1194_), .ZN(new_n4517_));
  NAND3_X1   g04324(.A1(new_n4512_), .A2(new_n4513_), .A3(new_n4517_), .ZN(new_n4518_));
  OAI22_X1   g04325(.A1(new_n4514_), .A2(new_n4515_), .B1(new_n4518_), .B2(new_n4516_), .ZN(new_n4519_));
  XOR2_X1    g04326(.A1(new_n4511_), .A2(new_n4519_), .Z(new_n4520_));
  NAND2_X1   g04327(.A1(new_n4275_), .A2(new_n4284_), .ZN(new_n4521_));
  NAND2_X1   g04328(.A1(new_n4286_), .A2(new_n4521_), .ZN(new_n4522_));
  NAND4_X1   g04329(.A1(\a[6] ), .A2(\a[13] ), .A3(\a[35] ), .A4(\a[42] ), .ZN(new_n4523_));
  NOR4_X1    g04330(.A1(new_n367_), .A2(new_n759_), .A3(new_n2442_), .A4(new_n3746_), .ZN(new_n4524_));
  NOR2_X1    g04331(.A1(new_n767_), .A2(new_n2746_), .ZN(new_n4525_));
  OAI21_X1   g04332(.A1(new_n4525_), .A2(new_n4524_), .B(new_n4523_), .ZN(new_n4526_));
  NAND3_X1   g04333(.A1(new_n4526_), .A2(\a[14] ), .A3(\a[34] ), .ZN(new_n4527_));
  NAND2_X1   g04334(.A1(new_n4526_), .A2(new_n4523_), .ZN(new_n4528_));
  AOI22_X1   g04335(.A1(\a[6] ), .A2(\a[42] ), .B1(\a[13] ), .B2(\a[35] ), .ZN(new_n4529_));
  OAI21_X1   g04336(.A1(new_n4528_), .A2(new_n4529_), .B(new_n4527_), .ZN(new_n4530_));
  NOR2_X1    g04337(.A1(new_n422_), .A2(new_n3327_), .ZN(new_n4531_));
  INV_X1     g04338(.I(new_n4531_), .ZN(new_n4532_));
  NAND2_X1   g04339(.A1(new_n3231_), .A2(new_n4531_), .ZN(new_n4533_));
  NOR2_X1    g04340(.A1(new_n3221_), .A2(new_n3327_), .ZN(new_n4534_));
  NAND2_X1   g04341(.A1(new_n4534_), .A2(new_n693_), .ZN(new_n4535_));
  AOI22_X1   g04342(.A1(new_n4533_), .A2(new_n4535_), .B1(new_n3819_), .B2(new_n4276_), .ZN(new_n4536_));
  AOI21_X1   g04343(.A1(\a[8] ), .A2(\a[40] ), .B(new_n3231_), .ZN(new_n4537_));
  NAND2_X1   g04344(.A1(new_n3819_), .A2(new_n4276_), .ZN(new_n4538_));
  NAND3_X1   g04345(.A1(new_n4533_), .A2(new_n4538_), .A3(new_n4535_), .ZN(new_n4539_));
  OAI22_X1   g04346(.A1(new_n4536_), .A2(new_n4532_), .B1(new_n4539_), .B2(new_n4537_), .ZN(new_n4540_));
  XOR2_X1    g04347(.A1(new_n4530_), .A2(new_n4540_), .Z(new_n4541_));
  NOR2_X1    g04348(.A1(new_n403_), .A2(new_n3116_), .ZN(new_n4542_));
  INV_X1     g04349(.I(new_n4542_), .ZN(new_n4543_));
  NAND2_X1   g04350(.A1(new_n4209_), .A2(new_n540_), .ZN(new_n4544_));
  NOR2_X1    g04351(.A1(new_n2752_), .A2(new_n3116_), .ZN(new_n4545_));
  NAND2_X1   g04352(.A1(new_n1060_), .A2(new_n4545_), .ZN(new_n4546_));
  AOI22_X1   g04353(.A1(new_n4546_), .A2(new_n4544_), .B1(new_n747_), .B2(new_n3803_), .ZN(new_n4547_));
  AOI21_X1   g04354(.A1(\a[10] ), .A2(\a[38] ), .B(new_n3799_), .ZN(new_n4548_));
  NAND2_X1   g04355(.A1(new_n747_), .A2(new_n3803_), .ZN(new_n4549_));
  NAND3_X1   g04356(.A1(new_n4549_), .A2(new_n4546_), .A3(new_n4544_), .ZN(new_n4550_));
  OAI22_X1   g04357(.A1(new_n4547_), .A2(new_n4543_), .B1(new_n4550_), .B2(new_n4548_), .ZN(new_n4551_));
  XOR2_X1    g04358(.A1(new_n4541_), .A2(new_n4551_), .Z(new_n4552_));
  XOR2_X1    g04359(.A1(new_n4522_), .A2(new_n4552_), .Z(new_n4553_));
  XOR2_X1    g04360(.A1(new_n4553_), .A2(new_n4520_), .Z(new_n4554_));
  XOR2_X1    g04361(.A1(new_n4494_), .A2(new_n4554_), .Z(new_n4555_));
  NOR2_X1    g04362(.A1(new_n4490_), .A2(new_n4555_), .ZN(new_n4556_));
  NAND2_X1   g04363(.A1(new_n4490_), .A2(new_n4555_), .ZN(new_n4557_));
  INV_X1     g04364(.I(new_n4557_), .ZN(new_n4558_));
  NOR2_X1    g04365(.A1(new_n4558_), .A2(new_n4556_), .ZN(new_n4559_));
  INV_X1     g04366(.I(new_n4559_), .ZN(new_n4560_));
  AND3_X2    g04367(.A1(new_n4486_), .A2(new_n4485_), .A3(new_n4560_), .Z(new_n4561_));
  AOI21_X1   g04368(.A1(new_n4486_), .A2(new_n4485_), .B(new_n4560_), .ZN(new_n4562_));
  NOR2_X1    g04369(.A1(new_n4561_), .A2(new_n4562_), .ZN(new_n4563_));
  XNOR2_X1   g04370(.A1(new_n4563_), .A2(new_n4484_), .ZN(new_n4564_));
  INV_X1     g04371(.I(new_n4564_), .ZN(new_n4565_));
  NOR2_X1    g04372(.A1(new_n4406_), .A2(new_n4565_), .ZN(new_n4566_));
  INV_X1     g04373(.I(new_n4566_), .ZN(new_n4567_));
  AOI21_X1   g04374(.A1(new_n4241_), .A2(new_n4236_), .B(new_n4400_), .ZN(new_n4568_));
  NOR2_X1    g04375(.A1(new_n4568_), .A2(new_n4398_), .ZN(new_n4569_));
  INV_X1     g04376(.I(new_n4398_), .ZN(new_n4570_));
  INV_X1     g04377(.I(new_n3912_), .ZN(new_n4571_));
  INV_X1     g04378(.I(new_n3768_), .ZN(new_n4572_));
  INV_X1     g04379(.I(new_n3464_), .ZN(new_n4573_));
  OAI21_X1   g04380(.A1(new_n3311_), .A2(new_n3296_), .B(new_n3465_), .ZN(new_n4574_));
  AOI21_X1   g04381(.A1(new_n4574_), .A2(new_n4573_), .B(new_n3607_), .ZN(new_n4575_));
  OAI21_X1   g04382(.A1(new_n4575_), .A2(new_n3609_), .B(new_n3769_), .ZN(new_n4576_));
  AOI21_X1   g04383(.A1(new_n4576_), .A2(new_n4572_), .B(new_n3910_), .ZN(new_n4577_));
  INV_X1     g04384(.I(new_n4070_), .ZN(new_n4578_));
  OAI21_X1   g04385(.A1(new_n4577_), .A2(new_n4571_), .B(new_n4578_), .ZN(new_n4579_));
  AOI21_X1   g04386(.A1(new_n4579_), .A2(new_n4071_), .B(new_n4237_), .ZN(new_n4580_));
  OAI21_X1   g04387(.A1(new_n4580_), .A2(new_n4235_), .B(new_n4399_), .ZN(new_n4581_));
  NOR2_X1    g04388(.A1(new_n4405_), .A2(new_n4564_), .ZN(new_n4582_));
  AOI21_X1   g04389(.A1(new_n4581_), .A2(new_n4570_), .B(new_n4582_), .ZN(new_n4583_));
  INV_X1     g04390(.I(new_n4582_), .ZN(new_n4584_));
  NAND2_X1   g04391(.A1(new_n4567_), .A2(new_n4584_), .ZN(new_n4585_));
  AOI22_X1   g04392(.A1(new_n4583_), .A2(new_n4567_), .B1(new_n4569_), .B2(new_n4585_), .ZN(\asquared[49] ));
  OAI21_X1   g04393(.A1(new_n4568_), .A2(new_n4398_), .B(new_n4584_), .ZN(new_n4587_));
  NAND2_X1   g04394(.A1(new_n4587_), .A2(new_n4567_), .ZN(new_n4588_));
  XOR2_X1    g04395(.A1(new_n4436_), .A2(new_n4501_), .Z(new_n4589_));
  XOR2_X1    g04396(.A1(new_n4589_), .A2(new_n4509_), .Z(new_n4590_));
  NAND2_X1   g04397(.A1(new_n4530_), .A2(new_n4540_), .ZN(new_n4591_));
  NAND2_X1   g04398(.A1(new_n4541_), .A2(new_n4551_), .ZN(new_n4592_));
  NAND2_X1   g04399(.A1(new_n4592_), .A2(new_n4591_), .ZN(new_n4593_));
  NOR2_X1    g04400(.A1(new_n1443_), .A2(new_n4460_), .ZN(new_n4594_));
  AOI21_X1   g04401(.A1(\a[1] ), .A2(\a[48] ), .B(\a[25] ), .ZN(new_n4595_));
  INV_X1     g04402(.I(\a[48] ), .ZN(new_n4596_));
  NOR2_X1    g04403(.A1(new_n1593_), .A2(new_n4596_), .ZN(new_n4597_));
  NOR2_X1    g04404(.A1(new_n4597_), .A2(new_n4595_), .ZN(new_n4598_));
  XOR2_X1    g04405(.A1(new_n4598_), .A2(new_n4594_), .Z(new_n4599_));
  XOR2_X1    g04406(.A1(new_n4599_), .A2(new_n4550_), .Z(new_n4600_));
  XOR2_X1    g04407(.A1(new_n4593_), .A2(new_n4600_), .Z(new_n4601_));
  XOR2_X1    g04408(.A1(new_n4601_), .A2(new_n4590_), .Z(new_n4602_));
  NAND2_X1   g04409(.A1(new_n4457_), .A2(new_n4463_), .ZN(new_n4603_));
  NAND2_X1   g04410(.A1(new_n4464_), .A2(new_n4455_), .ZN(new_n4604_));
  NAND2_X1   g04411(.A1(new_n4604_), .A2(new_n4603_), .ZN(new_n4605_));
  NAND2_X1   g04412(.A1(new_n4510_), .A2(new_n4503_), .ZN(new_n4606_));
  INV_X1     g04413(.I(new_n4511_), .ZN(new_n4607_));
  NAND2_X1   g04414(.A1(new_n4607_), .A2(new_n4519_), .ZN(new_n4608_));
  NAND2_X1   g04415(.A1(new_n4608_), .A2(new_n4606_), .ZN(new_n4609_));
  XOR2_X1    g04416(.A1(new_n4528_), .A2(new_n4518_), .Z(new_n4610_));
  XOR2_X1    g04417(.A1(new_n4610_), .A2(new_n4539_), .Z(new_n4611_));
  XOR2_X1    g04418(.A1(new_n4609_), .A2(new_n4611_), .Z(new_n4612_));
  XOR2_X1    g04419(.A1(new_n4612_), .A2(new_n4605_), .Z(new_n4613_));
  NOR2_X1    g04420(.A1(new_n4522_), .A2(new_n4552_), .ZN(new_n4614_));
  NAND2_X1   g04421(.A1(new_n4522_), .A2(new_n4552_), .ZN(new_n4615_));
  OAI21_X1   g04422(.A1(new_n4520_), .A2(new_n4614_), .B(new_n4615_), .ZN(new_n4616_));
  NAND2_X1   g04423(.A1(new_n4613_), .A2(new_n4616_), .ZN(new_n4617_));
  INV_X1     g04424(.I(new_n4617_), .ZN(new_n4618_));
  NOR2_X1    g04425(.A1(new_n4613_), .A2(new_n4616_), .ZN(new_n4619_));
  NOR2_X1    g04426(.A1(new_n4618_), .A2(new_n4619_), .ZN(new_n4620_));
  NOR2_X1    g04427(.A1(new_n4620_), .A2(new_n4602_), .ZN(new_n4621_));
  NAND2_X1   g04428(.A1(new_n4620_), .A2(new_n4602_), .ZN(new_n4622_));
  INV_X1     g04429(.I(new_n4622_), .ZN(new_n4623_));
  NOR2_X1    g04430(.A1(new_n4494_), .A2(new_n4554_), .ZN(new_n4624_));
  NOR2_X1    g04431(.A1(new_n4558_), .A2(new_n4624_), .ZN(new_n4625_));
  NAND2_X1   g04432(.A1(new_n4347_), .A2(new_n4326_), .ZN(new_n4626_));
  NAND2_X1   g04433(.A1(new_n4407_), .A2(new_n4317_), .ZN(new_n4627_));
  NAND2_X1   g04434(.A1(new_n4627_), .A2(new_n4626_), .ZN(new_n4628_));
  NAND2_X1   g04435(.A1(new_n4367_), .A2(new_n4336_), .ZN(new_n4629_));
  NAND2_X1   g04436(.A1(new_n4440_), .A2(new_n4378_), .ZN(new_n4630_));
  NAND2_X1   g04437(.A1(new_n4630_), .A2(new_n4629_), .ZN(new_n4631_));
  NAND2_X1   g04438(.A1(new_n4357_), .A2(new_n4283_), .ZN(new_n4632_));
  NAND2_X1   g04439(.A1(new_n4426_), .A2(new_n4437_), .ZN(new_n4633_));
  NAND2_X1   g04440(.A1(new_n4633_), .A2(new_n4632_), .ZN(new_n4634_));
  XOR2_X1    g04441(.A1(new_n4631_), .A2(new_n4634_), .Z(new_n4635_));
  XOR2_X1    g04442(.A1(new_n4635_), .A2(new_n4628_), .Z(new_n4636_));
  INV_X1     g04443(.I(new_n4636_), .ZN(new_n4637_));
  NAND2_X1   g04444(.A1(new_n4444_), .A2(new_n4441_), .ZN(new_n4638_));
  NAND2_X1   g04445(.A1(new_n4445_), .A2(new_n4439_), .ZN(new_n4639_));
  NAND2_X1   g04446(.A1(new_n4639_), .A2(new_n4638_), .ZN(new_n4640_));
  INV_X1     g04447(.I(new_n4416_), .ZN(new_n4641_));
  NOR2_X1    g04448(.A1(new_n4641_), .A2(new_n4412_), .ZN(new_n4642_));
  NOR2_X1    g04449(.A1(new_n4419_), .A2(new_n4642_), .ZN(new_n4643_));
  XOR2_X1    g04450(.A1(new_n4643_), .A2(new_n4640_), .Z(new_n4644_));
  NOR2_X1    g04451(.A1(new_n4644_), .A2(new_n4637_), .ZN(new_n4645_));
  INV_X1     g04452(.I(new_n4645_), .ZN(new_n4646_));
  NAND2_X1   g04453(.A1(new_n4644_), .A2(new_n4637_), .ZN(new_n4647_));
  AND2_X2    g04454(.A1(new_n4646_), .A2(new_n4647_), .Z(new_n4648_));
  NOR2_X1    g04455(.A1(new_n4625_), .A2(new_n4648_), .ZN(new_n4649_));
  INV_X1     g04456(.I(new_n4648_), .ZN(new_n4650_));
  NOR2_X1    g04457(.A1(new_n4625_), .A2(new_n4650_), .ZN(new_n4651_));
  NOR2_X1    g04458(.A1(new_n4651_), .A2(new_n4650_), .ZN(new_n4652_));
  NOR2_X1    g04459(.A1(new_n4652_), .A2(new_n4649_), .ZN(new_n4653_));
  NOR3_X1    g04460(.A1(new_n4653_), .A2(new_n4621_), .A3(new_n4623_), .ZN(new_n4654_));
  NOR2_X1    g04461(.A1(new_n4623_), .A2(new_n4621_), .ZN(new_n4655_));
  NOR3_X1    g04462(.A1(new_n4652_), .A2(new_n4655_), .A3(new_n4649_), .ZN(new_n4656_));
  NOR2_X1    g04463(.A1(new_n4654_), .A2(new_n4656_), .ZN(new_n4657_));
  NAND2_X1   g04464(.A1(new_n4475_), .A2(new_n4452_), .ZN(new_n4658_));
  NAND2_X1   g04465(.A1(new_n4481_), .A2(new_n4658_), .ZN(new_n4659_));
  NAND2_X1   g04466(.A1(new_n4425_), .A2(new_n4446_), .ZN(new_n4660_));
  NAND2_X1   g04467(.A1(new_n4449_), .A2(new_n4660_), .ZN(new_n4661_));
  NAND2_X1   g04468(.A1(new_n4471_), .A2(new_n4468_), .ZN(new_n4662_));
  NAND2_X1   g04469(.A1(new_n4473_), .A2(new_n4662_), .ZN(new_n4663_));
  NOR2_X1    g04470(.A1(new_n355_), .A2(new_n3327_), .ZN(new_n4664_));
  AOI21_X1   g04471(.A1(\a[7] ), .A2(\a[42] ), .B(new_n4664_), .ZN(new_n4665_));
  INV_X1     g04472(.I(new_n4665_), .ZN(new_n4666_));
  INV_X1     g04473(.I(new_n4372_), .ZN(new_n4667_));
  NOR2_X1    g04474(.A1(new_n4667_), .A2(new_n415_), .ZN(new_n4668_));
  NOR2_X1    g04475(.A1(new_n597_), .A2(new_n2626_), .ZN(new_n4669_));
  AOI21_X1   g04476(.A1(new_n4666_), .A2(new_n4669_), .B(new_n4668_), .ZN(new_n4670_));
  INV_X1     g04477(.I(new_n4670_), .ZN(new_n4671_));
  OAI21_X1   g04478(.A1(new_n4668_), .A2(new_n4665_), .B(new_n4669_), .ZN(new_n4672_));
  OAI21_X1   g04479(.A1(new_n4671_), .A2(new_n4665_), .B(new_n4672_), .ZN(new_n4673_));
  NOR2_X1    g04480(.A1(new_n513_), .A2(new_n2914_), .ZN(new_n4674_));
  NOR2_X1    g04481(.A1(new_n1778_), .A2(new_n2083_), .ZN(new_n4675_));
  NOR2_X1    g04482(.A1(new_n1779_), .A2(new_n2084_), .ZN(new_n4676_));
  OAI21_X1   g04483(.A1(new_n4676_), .A2(new_n4675_), .B(new_n4674_), .ZN(new_n4677_));
  INV_X1     g04484(.I(new_n4675_), .ZN(new_n4678_));
  AOI21_X1   g04485(.A1(new_n4674_), .A2(new_n4678_), .B(new_n4676_), .ZN(new_n4679_));
  NAND2_X1   g04486(.A1(new_n4679_), .A2(new_n4678_), .ZN(new_n4680_));
  NAND2_X1   g04487(.A1(new_n4680_), .A2(new_n4677_), .ZN(new_n4681_));
  XOR2_X1    g04488(.A1(new_n4673_), .A2(new_n4681_), .Z(new_n4682_));
  NOR4_X1    g04489(.A1(new_n367_), .A2(new_n759_), .A3(new_n2524_), .A4(new_n3666_), .ZN(new_n4683_));
  NAND4_X1   g04490(.A1(\a[6] ), .A2(\a[15] ), .A3(\a[34] ), .A4(\a[43] ), .ZN(new_n4684_));
  NAND2_X1   g04491(.A1(new_n897_), .A2(new_n2745_), .ZN(new_n4685_));
  AOI21_X1   g04492(.A1(new_n4685_), .A2(new_n4684_), .B(new_n4683_), .ZN(new_n4686_));
  NAND2_X1   g04493(.A1(\a[15] ), .A2(\a[34] ), .ZN(new_n4687_));
  AOI22_X1   g04494(.A1(\a[6] ), .A2(\a[43] ), .B1(\a[14] ), .B2(\a[35] ), .ZN(new_n4688_));
  NOR2_X1    g04495(.A1(new_n4686_), .A2(new_n4683_), .ZN(new_n4689_));
  INV_X1     g04496(.I(new_n4689_), .ZN(new_n4690_));
  OAI22_X1   g04497(.A1(new_n4690_), .A2(new_n4688_), .B1(new_n4686_), .B2(new_n4687_), .ZN(new_n4691_));
  XOR2_X1    g04498(.A1(new_n4682_), .A2(new_n4691_), .Z(new_n4692_));
  NAND2_X1   g04499(.A1(new_n1025_), .A2(new_n2275_), .ZN(new_n4693_));
  NAND2_X1   g04500(.A1(new_n1024_), .A2(new_n2636_), .ZN(new_n4694_));
  AOI22_X1   g04501(.A1(new_n4693_), .A2(new_n4694_), .B1(new_n1027_), .B2(new_n3210_), .ZN(new_n4695_));
  NAND2_X1   g04502(.A1(\a[16] ), .A2(\a[33] ), .ZN(new_n4696_));
  AOI22_X1   g04503(.A1(\a[17] ), .A2(\a[32] ), .B1(\a[18] ), .B2(\a[31] ), .ZN(new_n4697_));
  NAND2_X1   g04504(.A1(new_n1027_), .A2(new_n3210_), .ZN(new_n4698_));
  NAND3_X1   g04505(.A1(new_n4698_), .A2(new_n4693_), .A3(new_n4694_), .ZN(new_n4699_));
  OAI22_X1   g04506(.A1(new_n4695_), .A2(new_n4696_), .B1(new_n4699_), .B2(new_n4697_), .ZN(new_n4700_));
  OAI22_X1   g04507(.A1(new_n3859_), .A2(new_n229_), .B1(new_n595_), .B2(new_n4030_), .ZN(new_n4701_));
  INV_X1     g04508(.I(\a[49] ), .ZN(new_n4702_));
  NOR2_X1    g04509(.A1(new_n3859_), .A2(new_n4030_), .ZN(new_n4703_));
  INV_X1     g04510(.I(new_n4703_), .ZN(new_n4704_));
  NOR2_X1    g04511(.A1(new_n4704_), .A2(new_n242_), .ZN(new_n4705_));
  NOR2_X1    g04512(.A1(new_n4705_), .A2(new_n4702_), .ZN(new_n4706_));
  NAND2_X1   g04513(.A1(new_n4706_), .A2(new_n4701_), .ZN(new_n4707_));
  NOR2_X1    g04514(.A1(new_n196_), .A2(new_n4702_), .ZN(new_n4708_));
  INV_X1     g04515(.I(new_n4707_), .ZN(new_n4709_));
  NOR2_X1    g04516(.A1(new_n4709_), .A2(new_n4705_), .ZN(new_n4710_));
  OAI22_X1   g04517(.A1(new_n290_), .A2(new_n4030_), .B1(new_n253_), .B2(new_n3859_), .ZN(new_n4711_));
  AOI22_X1   g04518(.A1(new_n4710_), .A2(new_n4711_), .B1(new_n4707_), .B2(new_n4708_), .ZN(new_n4712_));
  NOR2_X1    g04519(.A1(new_n4302_), .A2(new_n4458_), .ZN(new_n4713_));
  NOR2_X1    g04520(.A1(new_n4459_), .A2(new_n4461_), .ZN(new_n4714_));
  NOR2_X1    g04521(.A1(new_n4714_), .A2(new_n4713_), .ZN(new_n4715_));
  XNOR2_X1   g04522(.A1(new_n4712_), .A2(new_n4715_), .ZN(new_n4716_));
  XNOR2_X1   g04523(.A1(new_n4716_), .A2(new_n4700_), .ZN(new_n4717_));
  AOI22_X1   g04524(.A1(\a[2] ), .A2(\a[47] ), .B1(\a[3] ), .B2(\a[46] ), .ZN(new_n4718_));
  INV_X1     g04525(.I(new_n4718_), .ZN(new_n4719_));
  NOR2_X1    g04526(.A1(new_n4178_), .A2(new_n4312_), .ZN(new_n4720_));
  INV_X1     g04527(.I(new_n4720_), .ZN(new_n4721_));
  NOR2_X1    g04528(.A1(new_n4721_), .A2(new_n246_), .ZN(new_n4722_));
  NOR2_X1    g04529(.A1(new_n1175_), .A2(new_n1750_), .ZN(new_n4723_));
  AOI21_X1   g04530(.A1(new_n4719_), .A2(new_n4723_), .B(new_n4722_), .ZN(new_n4724_));
  INV_X1     g04531(.I(new_n4724_), .ZN(new_n4725_));
  OAI21_X1   g04532(.A1(new_n4722_), .A2(new_n4718_), .B(new_n4723_), .ZN(new_n4726_));
  OAI21_X1   g04533(.A1(new_n4725_), .A2(new_n4718_), .B(new_n4726_), .ZN(new_n4727_));
  NOR2_X1    g04534(.A1(new_n1382_), .A2(new_n2679_), .ZN(new_n4728_));
  NOR2_X1    g04535(.A1(new_n1376_), .A2(new_n2255_), .ZN(new_n4729_));
  NOR2_X1    g04536(.A1(new_n1379_), .A2(new_n3811_), .ZN(new_n4730_));
  NOR2_X1    g04537(.A1(new_n4729_), .A2(new_n4730_), .ZN(new_n4731_));
  NOR2_X1    g04538(.A1(new_n4731_), .A2(new_n4728_), .ZN(new_n4732_));
  NAND2_X1   g04539(.A1(\a[19] ), .A2(\a[30] ), .ZN(new_n4733_));
  AOI22_X1   g04540(.A1(\a[20] ), .A2(\a[29] ), .B1(\a[21] ), .B2(\a[28] ), .ZN(new_n4734_));
  NOR2_X1    g04541(.A1(new_n4732_), .A2(new_n4728_), .ZN(new_n4735_));
  INV_X1     g04542(.I(new_n4735_), .ZN(new_n4736_));
  OAI22_X1   g04543(.A1(new_n4736_), .A2(new_n4734_), .B1(new_n4732_), .B2(new_n4733_), .ZN(new_n4737_));
  XNOR2_X1   g04544(.A1(new_n4737_), .A2(new_n4727_), .ZN(new_n4738_));
  INV_X1     g04545(.I(new_n4545_), .ZN(new_n4739_));
  NOR2_X1    g04546(.A1(new_n4739_), .A2(new_n534_), .ZN(new_n4740_));
  NOR2_X1    g04547(.A1(new_n2752_), .A2(new_n3221_), .ZN(new_n4741_));
  NAND3_X1   g04548(.A1(new_n4741_), .A2(\a[9] ), .A3(\a[12] ), .ZN(new_n4742_));
  NAND2_X1   g04549(.A1(new_n3550_), .A2(new_n540_), .ZN(new_n4743_));
  AOI21_X1   g04550(.A1(new_n4742_), .A2(new_n4743_), .B(new_n4740_), .ZN(new_n4744_));
  NAND2_X1   g04551(.A1(\a[9] ), .A2(\a[40] ), .ZN(new_n4745_));
  AOI22_X1   g04552(.A1(\a[10] ), .A2(\a[39] ), .B1(\a[12] ), .B2(\a[37] ), .ZN(new_n4746_));
  NOR2_X1    g04553(.A1(new_n4744_), .A2(new_n4740_), .ZN(new_n4747_));
  INV_X1     g04554(.I(new_n4747_), .ZN(new_n4748_));
  OAI22_X1   g04555(.A1(new_n4748_), .A2(new_n4746_), .B1(new_n4744_), .B2(new_n4745_), .ZN(new_n4749_));
  XOR2_X1    g04556(.A1(new_n4738_), .A2(new_n4749_), .Z(new_n4750_));
  XNOR2_X1   g04557(.A1(new_n4750_), .A2(new_n4717_), .ZN(new_n4751_));
  XOR2_X1    g04558(.A1(new_n4751_), .A2(new_n4692_), .Z(new_n4752_));
  XOR2_X1    g04559(.A1(new_n4663_), .A2(new_n4752_), .Z(new_n4753_));
  XOR2_X1    g04560(.A1(new_n4753_), .A2(new_n4661_), .Z(new_n4754_));
  XOR2_X1    g04561(.A1(new_n4659_), .A2(new_n4754_), .Z(new_n4755_));
  XNOR2_X1   g04562(.A1(new_n4657_), .A2(new_n4755_), .ZN(new_n4756_));
  NOR3_X1    g04563(.A1(new_n4561_), .A2(new_n4484_), .A3(new_n4562_), .ZN(new_n4757_));
  NOR2_X1    g04564(.A1(new_n4757_), .A2(new_n4562_), .ZN(new_n4758_));
  NOR2_X1    g04565(.A1(new_n4756_), .A2(new_n4758_), .ZN(new_n4759_));
  NAND2_X1   g04566(.A1(new_n4756_), .A2(new_n4758_), .ZN(new_n4760_));
  INV_X1     g04567(.I(new_n4760_), .ZN(new_n4761_));
  NOR2_X1    g04568(.A1(new_n4761_), .A2(new_n4759_), .ZN(new_n4762_));
  XOR2_X1    g04569(.A1(new_n4588_), .A2(new_n4762_), .Z(\asquared[50] ));
  AOI21_X1   g04570(.A1(new_n4587_), .A2(new_n4567_), .B(new_n4761_), .ZN(new_n4764_));
  NOR2_X1    g04571(.A1(new_n4764_), .A2(new_n4759_), .ZN(new_n4765_));
  NAND2_X1   g04572(.A1(new_n4659_), .A2(new_n4754_), .ZN(new_n4766_));
  NAND2_X1   g04573(.A1(new_n4657_), .A2(new_n4755_), .ZN(new_n4767_));
  NAND2_X1   g04574(.A1(new_n4767_), .A2(new_n4766_), .ZN(new_n4768_));
  NAND2_X1   g04575(.A1(\a[1] ), .A2(\a[49] ), .ZN(new_n4769_));
  NOR2_X1    g04576(.A1(new_n2081_), .A2(new_n4769_), .ZN(new_n4770_));
  INV_X1     g04577(.I(new_n4770_), .ZN(new_n4771_));
  NAND2_X1   g04578(.A1(new_n2081_), .A2(new_n4769_), .ZN(new_n4772_));
  NAND2_X1   g04579(.A1(new_n4771_), .A2(new_n4772_), .ZN(new_n4773_));
  XOR2_X1    g04580(.A1(new_n4773_), .A2(new_n4679_), .Z(new_n4774_));
  NOR2_X1    g04581(.A1(new_n4774_), .A2(new_n4748_), .ZN(new_n4775_));
  AND2_X2    g04582(.A1(new_n4774_), .A2(new_n4748_), .Z(new_n4776_));
  NOR2_X1    g04583(.A1(new_n4776_), .A2(new_n4775_), .ZN(new_n4777_));
  INV_X1     g04584(.I(new_n4716_), .ZN(new_n4778_));
  NAND2_X1   g04585(.A1(new_n4778_), .A2(new_n4700_), .ZN(new_n4779_));
  OAI21_X1   g04586(.A1(new_n4712_), .A2(new_n4715_), .B(new_n4779_), .ZN(new_n4780_));
  NAND2_X1   g04587(.A1(new_n4737_), .A2(new_n4727_), .ZN(new_n4781_));
  INV_X1     g04588(.I(new_n4738_), .ZN(new_n4782_));
  NAND2_X1   g04589(.A1(new_n4782_), .A2(new_n4749_), .ZN(new_n4783_));
  NAND2_X1   g04590(.A1(new_n4783_), .A2(new_n4781_), .ZN(new_n4784_));
  XOR2_X1    g04591(.A1(new_n4780_), .A2(new_n4784_), .Z(new_n4785_));
  XOR2_X1    g04592(.A1(new_n4785_), .A2(new_n4777_), .Z(new_n4786_));
  NAND2_X1   g04593(.A1(new_n4631_), .A2(new_n4634_), .ZN(new_n4787_));
  NAND2_X1   g04594(.A1(new_n4635_), .A2(new_n4628_), .ZN(new_n4788_));
  NAND2_X1   g04595(.A1(new_n4788_), .A2(new_n4787_), .ZN(new_n4789_));
  NAND2_X1   g04596(.A1(new_n4673_), .A2(new_n4681_), .ZN(new_n4790_));
  NAND2_X1   g04597(.A1(new_n4682_), .A2(new_n4691_), .ZN(new_n4791_));
  NAND2_X1   g04598(.A1(new_n4791_), .A2(new_n4790_), .ZN(new_n4792_));
  XNOR2_X1   g04599(.A1(new_n4735_), .A2(new_n4699_), .ZN(new_n4793_));
  XOR2_X1    g04600(.A1(new_n4793_), .A2(new_n4671_), .Z(new_n4794_));
  XOR2_X1    g04601(.A1(new_n4794_), .A2(new_n4792_), .Z(new_n4795_));
  XOR2_X1    g04602(.A1(new_n4789_), .A2(new_n4795_), .Z(new_n4796_));
  INV_X1     g04603(.I(new_n4717_), .ZN(new_n4797_));
  NAND2_X1   g04604(.A1(new_n4751_), .A2(new_n4692_), .ZN(new_n4798_));
  OAI21_X1   g04605(.A1(new_n4797_), .A2(new_n4750_), .B(new_n4798_), .ZN(new_n4799_));
  XOR2_X1    g04606(.A1(new_n4799_), .A2(new_n4796_), .Z(new_n4800_));
  XNOR2_X1   g04607(.A1(new_n4800_), .A2(new_n4786_), .ZN(new_n4801_));
  NAND2_X1   g04608(.A1(new_n4663_), .A2(new_n4752_), .ZN(new_n4802_));
  NAND2_X1   g04609(.A1(new_n4753_), .A2(new_n4661_), .ZN(new_n4803_));
  NAND2_X1   g04610(.A1(new_n4803_), .A2(new_n4802_), .ZN(new_n4804_));
  XOR2_X1    g04611(.A1(new_n4710_), .A2(new_n4724_), .Z(new_n4805_));
  NOR2_X1    g04612(.A1(new_n4805_), .A2(new_n4690_), .ZN(new_n4806_));
  AND2_X2    g04613(.A1(new_n4805_), .A2(new_n4690_), .Z(new_n4807_));
  NOR2_X1    g04614(.A1(new_n4807_), .A2(new_n4806_), .ZN(new_n4808_));
  INV_X1     g04615(.I(new_n4808_), .ZN(new_n4809_));
  NAND2_X1   g04616(.A1(new_n4528_), .A2(new_n4518_), .ZN(new_n4810_));
  NAND2_X1   g04617(.A1(new_n4610_), .A2(new_n4539_), .ZN(new_n4811_));
  NAND2_X1   g04618(.A1(new_n4811_), .A2(new_n4810_), .ZN(new_n4812_));
  NAND2_X1   g04619(.A1(new_n4436_), .A2(new_n4501_), .ZN(new_n4813_));
  NAND2_X1   g04620(.A1(new_n4589_), .A2(new_n4509_), .ZN(new_n4814_));
  NAND2_X1   g04621(.A1(new_n4814_), .A2(new_n4813_), .ZN(new_n4815_));
  NOR2_X1    g04622(.A1(new_n4815_), .A2(new_n4812_), .ZN(new_n4816_));
  NAND2_X1   g04623(.A1(new_n4815_), .A2(new_n4812_), .ZN(new_n4817_));
  INV_X1     g04624(.I(new_n4817_), .ZN(new_n4818_));
  NOR2_X1    g04625(.A1(new_n4818_), .A2(new_n4816_), .ZN(new_n4819_));
  INV_X1     g04626(.I(new_n4819_), .ZN(new_n4820_));
  NOR2_X1    g04627(.A1(new_n4820_), .A2(new_n4809_), .ZN(new_n4821_));
  INV_X1     g04628(.I(new_n4821_), .ZN(new_n4822_));
  NAND2_X1   g04629(.A1(new_n4820_), .A2(new_n4809_), .ZN(new_n4823_));
  AND2_X2    g04630(.A1(new_n4822_), .A2(new_n4823_), .Z(new_n4824_));
  NAND2_X1   g04631(.A1(new_n4609_), .A2(new_n4611_), .ZN(new_n4825_));
  NAND2_X1   g04632(.A1(new_n4612_), .A2(new_n4605_), .ZN(new_n4826_));
  NAND2_X1   g04633(.A1(new_n4826_), .A2(new_n4825_), .ZN(new_n4827_));
  NAND2_X1   g04634(.A1(new_n4593_), .A2(new_n4600_), .ZN(new_n4828_));
  NAND2_X1   g04635(.A1(new_n4601_), .A2(new_n4590_), .ZN(new_n4829_));
  NAND2_X1   g04636(.A1(new_n4829_), .A2(new_n4828_), .ZN(new_n4830_));
  XOR2_X1    g04637(.A1(new_n4827_), .A2(new_n4830_), .Z(new_n4831_));
  XOR2_X1    g04638(.A1(new_n4831_), .A2(new_n4824_), .Z(new_n4832_));
  XOR2_X1    g04639(.A1(new_n4804_), .A2(new_n4832_), .Z(new_n4833_));
  XNOR2_X1   g04640(.A1(new_n4833_), .A2(new_n4801_), .ZN(new_n4834_));
  INV_X1     g04641(.I(new_n4834_), .ZN(new_n4835_));
  NOR2_X1    g04642(.A1(new_n4654_), .A2(new_n4651_), .ZN(new_n4836_));
  NOR2_X1    g04643(.A1(new_n4623_), .A2(new_n4618_), .ZN(new_n4837_));
  OAI21_X1   g04644(.A1(new_n4642_), .A2(new_n4419_), .B(new_n4640_), .ZN(new_n4838_));
  NAND2_X1   g04645(.A1(new_n4646_), .A2(new_n4838_), .ZN(new_n4839_));
  INV_X1     g04646(.I(new_n4839_), .ZN(new_n4840_));
  NAND2_X1   g04647(.A1(new_n4598_), .A2(new_n4594_), .ZN(new_n4841_));
  NAND2_X1   g04648(.A1(new_n4599_), .A2(new_n4550_), .ZN(new_n4842_));
  NAND2_X1   g04649(.A1(new_n4842_), .A2(new_n4841_), .ZN(new_n4843_));
  NOR2_X1    g04650(.A1(new_n2524_), .A2(new_n4030_), .ZN(new_n4844_));
  NAND2_X1   g04651(.A1(new_n1054_), .A2(new_n4844_), .ZN(new_n4845_));
  INV_X1     g04652(.I(new_n4845_), .ZN(new_n4846_));
  INV_X1     g04653(.I(new_n3084_), .ZN(new_n4847_));
  NOR2_X1    g04654(.A1(new_n742_), .A2(new_n4030_), .ZN(new_n4848_));
  INV_X1     g04655(.I(new_n4848_), .ZN(new_n4849_));
  NOR2_X1    g04656(.A1(new_n4847_), .A2(new_n4849_), .ZN(new_n4850_));
  NOR2_X1    g04657(.A1(new_n2746_), .A2(new_n893_), .ZN(new_n4851_));
  NOR2_X1    g04658(.A1(new_n4850_), .A2(new_n4851_), .ZN(new_n4852_));
  NOR2_X1    g04659(.A1(new_n4852_), .A2(new_n4846_), .ZN(new_n4853_));
  NAND2_X1   g04660(.A1(\a[16] ), .A2(\a[34] ), .ZN(new_n4854_));
  NOR2_X1    g04661(.A1(new_n4853_), .A2(new_n4846_), .ZN(new_n4855_));
  INV_X1     g04662(.I(new_n4855_), .ZN(new_n4856_));
  AOI22_X1   g04663(.A1(\a[5] ), .A2(\a[45] ), .B1(\a[15] ), .B2(\a[35] ), .ZN(new_n4857_));
  OAI22_X1   g04664(.A1(new_n4856_), .A2(new_n4857_), .B1(new_n4853_), .B2(new_n4854_), .ZN(new_n4858_));
  NAND4_X1   g04665(.A1(\a[18] ), .A2(\a[23] ), .A3(\a[27] ), .A4(\a[32] ), .ZN(new_n4859_));
  NOR2_X1    g04666(.A1(new_n1718_), .A2(new_n2200_), .ZN(new_n4860_));
  NAND2_X1   g04667(.A1(new_n3220_), .A2(new_n4860_), .ZN(new_n4861_));
  OAI21_X1   g04668(.A1(new_n2385_), .A2(new_n2189_), .B(new_n4861_), .ZN(new_n4862_));
  NAND2_X1   g04669(.A1(new_n4862_), .A2(new_n4859_), .ZN(new_n4863_));
  NAND3_X1   g04670(.A1(new_n4863_), .A2(\a[22] ), .A3(\a[28] ), .ZN(new_n4864_));
  NAND2_X1   g04671(.A1(new_n4863_), .A2(new_n4859_), .ZN(new_n4865_));
  AOI22_X1   g04672(.A1(\a[18] ), .A2(\a[32] ), .B1(\a[23] ), .B2(\a[27] ), .ZN(new_n4866_));
  OAI21_X1   g04673(.A1(new_n4865_), .A2(new_n4866_), .B(new_n4864_), .ZN(new_n4867_));
  XOR2_X1    g04674(.A1(new_n4858_), .A2(new_n4867_), .Z(new_n4868_));
  XOR2_X1    g04675(.A1(new_n4868_), .A2(new_n4843_), .Z(new_n4869_));
  NAND4_X1   g04676(.A1(\a[7] ), .A2(\a[14] ), .A3(\a[36] ), .A4(\a[43] ), .ZN(new_n4870_));
  NOR2_X1    g04677(.A1(new_n2626_), .A2(new_n3859_), .ZN(new_n4871_));
  NAND2_X1   g04678(.A1(new_n1053_), .A2(new_n4871_), .ZN(new_n4872_));
  OAI21_X1   g04679(.A1(new_n374_), .A2(new_n4343_), .B(new_n4872_), .ZN(new_n4873_));
  NAND2_X1   g04680(.A1(new_n4873_), .A2(new_n4870_), .ZN(new_n4874_));
  NAND3_X1   g04681(.A1(new_n4874_), .A2(\a[6] ), .A3(\a[44] ), .ZN(new_n4875_));
  NAND2_X1   g04682(.A1(new_n4874_), .A2(new_n4870_), .ZN(new_n4876_));
  AOI22_X1   g04683(.A1(\a[7] ), .A2(\a[43] ), .B1(\a[14] ), .B2(\a[36] ), .ZN(new_n4877_));
  OAI21_X1   g04684(.A1(new_n4876_), .A2(new_n4877_), .B(new_n4875_), .ZN(new_n4878_));
  NOR2_X1    g04685(.A1(new_n2752_), .A2(new_n3327_), .ZN(new_n4879_));
  NAND2_X1   g04686(.A1(new_n4879_), .A2(new_n1184_), .ZN(new_n4880_));
  NOR4_X1    g04687(.A1(new_n355_), .A2(new_n597_), .A3(new_n2752_), .A4(new_n3746_), .ZN(new_n4881_));
  NOR2_X1    g04688(.A1(new_n4667_), .A2(new_n1427_), .ZN(new_n4882_));
  OAI21_X1   g04689(.A1(new_n4882_), .A2(new_n4881_), .B(new_n4880_), .ZN(new_n4883_));
  NAND3_X1   g04690(.A1(new_n4883_), .A2(\a[8] ), .A3(\a[42] ), .ZN(new_n4884_));
  NAND2_X1   g04691(.A1(new_n4883_), .A2(new_n4880_), .ZN(new_n4885_));
  AOI21_X1   g04692(.A1(\a[9] ), .A2(\a[41] ), .B(new_n3035_), .ZN(new_n4886_));
  OAI21_X1   g04693(.A1(new_n4885_), .A2(new_n4886_), .B(new_n4884_), .ZN(new_n4887_));
  XNOR2_X1   g04694(.A1(new_n4878_), .A2(new_n4887_), .ZN(new_n4888_));
  NOR2_X1    g04695(.A1(new_n1264_), .A2(new_n3551_), .ZN(new_n4889_));
  AOI22_X1   g04696(.A1(new_n535_), .A2(new_n3222_), .B1(new_n4209_), .B2(new_n1261_), .ZN(new_n4890_));
  NOR2_X1    g04697(.A1(new_n4889_), .A2(new_n4890_), .ZN(new_n4891_));
  NAND2_X1   g04698(.A1(\a[12] ), .A2(\a[38] ), .ZN(new_n4892_));
  NOR2_X1    g04699(.A1(new_n417_), .A2(new_n3221_), .ZN(new_n4893_));
  AOI21_X1   g04700(.A1(\a[11] ), .A2(\a[39] ), .B(new_n4893_), .ZN(new_n4894_));
  NOR2_X1    g04701(.A1(new_n4891_), .A2(new_n4889_), .ZN(new_n4895_));
  INV_X1     g04702(.I(new_n4895_), .ZN(new_n4896_));
  OAI22_X1   g04703(.A1(new_n4896_), .A2(new_n4894_), .B1(new_n4891_), .B2(new_n4892_), .ZN(new_n4897_));
  XOR2_X1    g04704(.A1(new_n4888_), .A2(new_n4897_), .Z(new_n4898_));
  AOI22_X1   g04705(.A1(\a[0] ), .A2(\a[50] ), .B1(\a[2] ), .B2(\a[48] ), .ZN(new_n4899_));
  INV_X1     g04706(.I(new_n4899_), .ZN(new_n4900_));
  INV_X1     g04707(.I(\a[50] ), .ZN(new_n4901_));
  NOR2_X1    g04708(.A1(new_n4596_), .A2(new_n4901_), .ZN(new_n4902_));
  INV_X1     g04709(.I(new_n4902_), .ZN(new_n4903_));
  NOR2_X1    g04710(.A1(new_n4903_), .A2(new_n412_), .ZN(new_n4904_));
  AOI21_X1   g04711(.A1(new_n4597_), .A2(new_n4900_), .B(new_n4904_), .ZN(new_n4905_));
  INV_X1     g04712(.I(new_n4905_), .ZN(new_n4906_));
  OAI21_X1   g04713(.A1(new_n4904_), .A2(new_n4899_), .B(new_n4597_), .ZN(new_n4907_));
  OAI21_X1   g04714(.A1(new_n4906_), .A2(new_n4899_), .B(new_n4907_), .ZN(new_n4908_));
  NOR3_X1    g04715(.A1(new_n1111_), .A2(new_n2274_), .A3(new_n4178_), .ZN(new_n4909_));
  NOR2_X1    g04716(.A1(new_n4721_), .A2(new_n370_), .ZN(new_n4910_));
  INV_X1     g04717(.I(new_n4910_), .ZN(new_n4911_));
  NAND3_X1   g04718(.A1(new_n2638_), .A2(\a[17] ), .A3(\a[47] ), .ZN(new_n4912_));
  AOI21_X1   g04719(.A1(new_n4911_), .A2(new_n4912_), .B(new_n4909_), .ZN(new_n4913_));
  NAND2_X1   g04720(.A1(\a[3] ), .A2(\a[47] ), .ZN(new_n4914_));
  AOI22_X1   g04721(.A1(\a[4] ), .A2(\a[46] ), .B1(\a[17] ), .B2(\a[33] ), .ZN(new_n4915_));
  NOR2_X1    g04722(.A1(new_n4913_), .A2(new_n4909_), .ZN(new_n4916_));
  INV_X1     g04723(.I(new_n4916_), .ZN(new_n4917_));
  OAI22_X1   g04724(.A1(new_n4917_), .A2(new_n4915_), .B1(new_n4913_), .B2(new_n4914_), .ZN(new_n4918_));
  XOR2_X1    g04725(.A1(new_n4918_), .A2(new_n4908_), .Z(new_n4919_));
  NAND2_X1   g04726(.A1(new_n1375_), .A2(new_n2437_), .ZN(new_n4920_));
  NAND2_X1   g04727(.A1(new_n1378_), .A2(new_n2976_), .ZN(new_n4921_));
  AOI22_X1   g04728(.A1(new_n4920_), .A2(new_n4921_), .B1(new_n1381_), .B2(new_n2254_), .ZN(new_n4922_));
  NAND2_X1   g04729(.A1(\a[19] ), .A2(\a[31] ), .ZN(new_n4923_));
  AOI22_X1   g04730(.A1(\a[20] ), .A2(\a[30] ), .B1(\a[21] ), .B2(\a[29] ), .ZN(new_n4924_));
  NAND2_X1   g04731(.A1(new_n1381_), .A2(new_n2254_), .ZN(new_n4925_));
  NAND3_X1   g04732(.A1(new_n4925_), .A2(new_n4920_), .A3(new_n4921_), .ZN(new_n4926_));
  OAI22_X1   g04733(.A1(new_n4922_), .A2(new_n4923_), .B1(new_n4926_), .B2(new_n4924_), .ZN(new_n4927_));
  XNOR2_X1   g04734(.A1(new_n4919_), .A2(new_n4927_), .ZN(new_n4928_));
  XOR2_X1    g04735(.A1(new_n4928_), .A2(new_n4898_), .Z(new_n4929_));
  AND2_X2    g04736(.A1(new_n4929_), .A2(new_n4869_), .Z(new_n4930_));
  NOR2_X1    g04737(.A1(new_n4929_), .A2(new_n4869_), .ZN(new_n4931_));
  NOR2_X1    g04738(.A1(new_n4930_), .A2(new_n4931_), .ZN(new_n4932_));
  NOR2_X1    g04739(.A1(new_n4840_), .A2(new_n4932_), .ZN(new_n4933_));
  INV_X1     g04740(.I(new_n4933_), .ZN(new_n4934_));
  INV_X1     g04741(.I(new_n4932_), .ZN(new_n4935_));
  NOR2_X1    g04742(.A1(new_n4839_), .A2(new_n4935_), .ZN(new_n4936_));
  INV_X1     g04743(.I(new_n4936_), .ZN(new_n4937_));
  AOI21_X1   g04744(.A1(new_n4934_), .A2(new_n4937_), .B(new_n4837_), .ZN(new_n4938_));
  INV_X1     g04745(.I(new_n4938_), .ZN(new_n4939_));
  NAND3_X1   g04746(.A1(new_n4934_), .A2(new_n4937_), .A3(new_n4837_), .ZN(new_n4940_));
  NAND2_X1   g04747(.A1(new_n4939_), .A2(new_n4940_), .ZN(new_n4941_));
  XNOR2_X1   g04748(.A1(new_n4836_), .A2(new_n4941_), .ZN(new_n4942_));
  XOR2_X1    g04749(.A1(new_n4942_), .A2(new_n4835_), .Z(new_n4943_));
  NAND2_X1   g04750(.A1(new_n4943_), .A2(new_n4768_), .ZN(new_n4944_));
  NOR2_X1    g04751(.A1(new_n4943_), .A2(new_n4768_), .ZN(new_n4945_));
  INV_X1     g04752(.I(new_n4945_), .ZN(new_n4946_));
  NAND2_X1   g04753(.A1(new_n4946_), .A2(new_n4944_), .ZN(new_n4947_));
  INV_X1     g04754(.I(new_n4759_), .ZN(new_n4948_));
  OAI21_X1   g04755(.A1(new_n4583_), .A2(new_n4566_), .B(new_n4760_), .ZN(new_n4949_));
  AOI21_X1   g04756(.A1(new_n4949_), .A2(new_n4948_), .B(new_n4945_), .ZN(new_n4950_));
  AOI22_X1   g04757(.A1(new_n4950_), .A2(new_n4944_), .B1(new_n4765_), .B2(new_n4947_), .ZN(\asquared[51] ));
  OAI21_X1   g04758(.A1(new_n4764_), .A2(new_n4759_), .B(new_n4946_), .ZN(new_n4952_));
  NAND2_X1   g04759(.A1(new_n4952_), .A2(new_n4944_), .ZN(new_n4953_));
  XNOR2_X1   g04760(.A1(new_n4916_), .A2(new_n4926_), .ZN(new_n4954_));
  XOR2_X1    g04761(.A1(new_n4954_), .A2(new_n4906_), .Z(new_n4955_));
  NAND2_X1   g04762(.A1(new_n4878_), .A2(new_n4887_), .ZN(new_n4956_));
  INV_X1     g04763(.I(new_n4897_), .ZN(new_n4957_));
  OAI21_X1   g04764(.A1(new_n4888_), .A2(new_n4957_), .B(new_n4956_), .ZN(new_n4958_));
  XOR2_X1    g04765(.A1(new_n4876_), .A2(new_n4885_), .Z(new_n4959_));
  XOR2_X1    g04766(.A1(new_n4959_), .A2(new_n4865_), .Z(new_n4960_));
  NOR2_X1    g04767(.A1(new_n4958_), .A2(new_n4960_), .ZN(new_n4961_));
  NAND2_X1   g04768(.A1(new_n4958_), .A2(new_n4960_), .ZN(new_n4962_));
  INV_X1     g04769(.I(new_n4962_), .ZN(new_n4963_));
  NOR2_X1    g04770(.A1(new_n4963_), .A2(new_n4961_), .ZN(new_n4964_));
  NOR2_X1    g04771(.A1(new_n4964_), .A2(new_n4955_), .ZN(new_n4965_));
  NAND2_X1   g04772(.A1(new_n4964_), .A2(new_n4955_), .ZN(new_n4966_));
  INV_X1     g04773(.I(new_n4966_), .ZN(new_n4967_));
  NOR2_X1    g04774(.A1(new_n4967_), .A2(new_n4965_), .ZN(new_n4968_));
  NOR2_X1    g04775(.A1(new_n4928_), .A2(new_n4898_), .ZN(new_n4969_));
  NOR2_X1    g04776(.A1(new_n4930_), .A2(new_n4969_), .ZN(new_n4970_));
  NOR2_X1    g04777(.A1(new_n4821_), .A2(new_n4818_), .ZN(new_n4971_));
  NAND2_X1   g04778(.A1(new_n4858_), .A2(new_n4867_), .ZN(new_n4972_));
  NAND2_X1   g04779(.A1(new_n4868_), .A2(new_n4843_), .ZN(new_n4973_));
  NAND2_X1   g04780(.A1(new_n4973_), .A2(new_n4972_), .ZN(new_n4974_));
  XOR2_X1    g04781(.A1(new_n4855_), .A2(new_n4895_), .Z(new_n4975_));
  NOR2_X1    g04782(.A1(new_n4312_), .A2(new_n4596_), .ZN(new_n4976_));
  INV_X1     g04783(.I(new_n4976_), .ZN(new_n4977_));
  NOR2_X1    g04784(.A1(new_n4312_), .A2(new_n4702_), .ZN(new_n4978_));
  INV_X1     g04785(.I(new_n4978_), .ZN(new_n4979_));
  NOR2_X1    g04786(.A1(new_n4596_), .A2(new_n4702_), .ZN(new_n4980_));
  INV_X1     g04787(.I(new_n4980_), .ZN(new_n4981_));
  OAI22_X1   g04788(.A1(new_n246_), .A2(new_n4981_), .B1(new_n4979_), .B2(new_n251_), .ZN(new_n4982_));
  OAI21_X1   g04789(.A1(new_n370_), .A2(new_n4977_), .B(new_n4982_), .ZN(new_n4983_));
  NAND3_X1   g04790(.A1(new_n4983_), .A2(\a[2] ), .A3(\a[49] ), .ZN(new_n4984_));
  AOI22_X1   g04791(.A1(\a[3] ), .A2(\a[48] ), .B1(\a[4] ), .B2(\a[47] ), .ZN(new_n4985_));
  NOR2_X1    g04792(.A1(new_n4977_), .A2(new_n370_), .ZN(new_n4986_));
  NOR2_X1    g04793(.A1(new_n4982_), .A2(new_n4986_), .ZN(new_n4987_));
  INV_X1     g04794(.I(new_n4987_), .ZN(new_n4988_));
  OAI21_X1   g04795(.A1(new_n4985_), .A2(new_n4988_), .B(new_n4984_), .ZN(new_n4989_));
  XOR2_X1    g04796(.A1(new_n4975_), .A2(new_n4989_), .Z(new_n4990_));
  XOR2_X1    g04797(.A1(new_n4974_), .A2(new_n4990_), .Z(new_n4991_));
  INV_X1     g04798(.I(new_n4991_), .ZN(new_n4992_));
  XOR2_X1    g04799(.A1(new_n4971_), .A2(new_n4992_), .Z(new_n4993_));
  XNOR2_X1   g04800(.A1(new_n4993_), .A2(new_n4970_), .ZN(new_n4994_));
  XNOR2_X1   g04801(.A1(new_n4994_), .A2(new_n4968_), .ZN(new_n4995_));
  OAI21_X1   g04802(.A1(new_n4840_), .A2(new_n4935_), .B(new_n4939_), .ZN(new_n4996_));
  NAND2_X1   g04803(.A1(new_n4918_), .A2(new_n4908_), .ZN(new_n4997_));
  NAND2_X1   g04804(.A1(new_n4919_), .A2(new_n4927_), .ZN(new_n4998_));
  NAND2_X1   g04805(.A1(new_n4998_), .A2(new_n4997_), .ZN(new_n4999_));
  NOR2_X1    g04806(.A1(new_n4710_), .A2(new_n4724_), .ZN(new_n5000_));
  NOR2_X1    g04807(.A1(new_n4807_), .A2(new_n5000_), .ZN(new_n5001_));
  NOR2_X1    g04808(.A1(new_n4773_), .A2(new_n4679_), .ZN(new_n5002_));
  NOR2_X1    g04809(.A1(new_n4776_), .A2(new_n5002_), .ZN(new_n5003_));
  XOR2_X1    g04810(.A1(new_n5001_), .A2(new_n5003_), .Z(new_n5004_));
  NAND2_X1   g04811(.A1(new_n5004_), .A2(new_n4999_), .ZN(new_n5005_));
  INV_X1     g04812(.I(new_n5005_), .ZN(new_n5006_));
  NOR2_X1    g04813(.A1(new_n5004_), .A2(new_n4999_), .ZN(new_n5007_));
  NOR2_X1    g04814(.A1(new_n5006_), .A2(new_n5007_), .ZN(new_n5008_));
  NAND2_X1   g04815(.A1(new_n4794_), .A2(new_n4792_), .ZN(new_n5009_));
  NAND2_X1   g04816(.A1(new_n4789_), .A2(new_n4795_), .ZN(new_n5010_));
  NAND2_X1   g04817(.A1(new_n5010_), .A2(new_n5009_), .ZN(new_n5011_));
  NAND2_X1   g04818(.A1(new_n4780_), .A2(new_n4784_), .ZN(new_n5012_));
  NAND2_X1   g04819(.A1(new_n4785_), .A2(new_n4777_), .ZN(new_n5013_));
  NAND2_X1   g04820(.A1(new_n5013_), .A2(new_n5012_), .ZN(new_n5014_));
  XOR2_X1    g04821(.A1(new_n5014_), .A2(new_n5011_), .Z(new_n5015_));
  XOR2_X1    g04822(.A1(new_n5015_), .A2(new_n5008_), .Z(new_n5016_));
  XOR2_X1    g04823(.A1(new_n4996_), .A2(new_n5016_), .Z(new_n5017_));
  INV_X1     g04824(.I(new_n5017_), .ZN(new_n5018_));
  NAND2_X1   g04825(.A1(new_n5018_), .A2(new_n4995_), .ZN(new_n5019_));
  OR2_X2     g04826(.A1(new_n5018_), .A2(new_n4995_), .Z(new_n5020_));
  NAND2_X1   g04827(.A1(new_n5020_), .A2(new_n5019_), .ZN(new_n5021_));
  NAND2_X1   g04828(.A1(new_n4804_), .A2(new_n4832_), .ZN(new_n5022_));
  INV_X1     g04829(.I(new_n4833_), .ZN(new_n5023_));
  OAI21_X1   g04830(.A1(new_n5023_), .A2(new_n4801_), .B(new_n5022_), .ZN(new_n5024_));
  NAND2_X1   g04831(.A1(new_n4799_), .A2(new_n4796_), .ZN(new_n5025_));
  NAND2_X1   g04832(.A1(new_n4800_), .A2(new_n4786_), .ZN(new_n5026_));
  NAND2_X1   g04833(.A1(new_n5026_), .A2(new_n5025_), .ZN(new_n5027_));
  NAND2_X1   g04834(.A1(new_n4827_), .A2(new_n4830_), .ZN(new_n5028_));
  NAND2_X1   g04835(.A1(new_n4831_), .A2(new_n4824_), .ZN(new_n5029_));
  NAND2_X1   g04836(.A1(new_n5029_), .A2(new_n5028_), .ZN(new_n5030_));
  NAND2_X1   g04837(.A1(new_n4736_), .A2(new_n4699_), .ZN(new_n5031_));
  NAND2_X1   g04838(.A1(new_n4793_), .A2(new_n4671_), .ZN(new_n5032_));
  NAND2_X1   g04839(.A1(new_n5032_), .A2(new_n5031_), .ZN(new_n5033_));
  NAND2_X1   g04840(.A1(\a[0] ), .A2(\a[51] ), .ZN(new_n5034_));
  XOR2_X1    g04841(.A1(new_n4770_), .A2(new_n5034_), .Z(new_n5035_));
  NAND2_X1   g04842(.A1(\a[1] ), .A2(\a[50] ), .ZN(new_n5036_));
  XOR2_X1    g04843(.A1(new_n5036_), .A2(\a[26] ), .Z(new_n5037_));
  XNOR2_X1   g04844(.A1(new_n5035_), .A2(new_n5037_), .ZN(new_n5038_));
  NOR2_X1    g04845(.A1(new_n1023_), .A2(new_n2442_), .ZN(new_n5039_));
  INV_X1     g04846(.I(new_n5039_), .ZN(new_n5040_));
  AOI22_X1   g04847(.A1(\a[19] ), .A2(\a[32] ), .B1(\a[20] ), .B2(\a[31] ), .ZN(new_n5041_));
  NOR2_X1    g04848(.A1(new_n1376_), .A2(new_n3833_), .ZN(new_n5042_));
  NOR3_X1    g04849(.A1(new_n5042_), .A2(new_n5040_), .A3(new_n5041_), .ZN(new_n5043_));
  NOR2_X1    g04850(.A1(new_n5043_), .A2(new_n5042_), .ZN(new_n5044_));
  INV_X1     g04851(.I(new_n5044_), .ZN(new_n5045_));
  OAI22_X1   g04852(.A1(new_n5045_), .A2(new_n5041_), .B1(new_n5040_), .B2(new_n5043_), .ZN(new_n5046_));
  XOR2_X1    g04853(.A1(new_n5038_), .A2(new_n5046_), .Z(new_n5047_));
  XNOR2_X1   g04854(.A1(new_n5033_), .A2(new_n5047_), .ZN(new_n5048_));
  NOR2_X1    g04855(.A1(new_n597_), .A2(new_n3666_), .ZN(new_n5049_));
  NAND3_X1   g04856(.A1(new_n5049_), .A2(\a[8] ), .A3(\a[38] ), .ZN(new_n5050_));
  NOR3_X1    g04857(.A1(new_n4041_), .A2(new_n597_), .A3(new_n3859_), .ZN(new_n5051_));
  NOR2_X1    g04858(.A1(new_n4343_), .A2(new_n415_), .ZN(new_n5052_));
  OAI21_X1   g04859(.A1(new_n5052_), .A2(new_n5051_), .B(new_n5050_), .ZN(new_n5053_));
  NAND3_X1   g04860(.A1(new_n5053_), .A2(\a[7] ), .A3(\a[44] ), .ZN(new_n5054_));
  NAND2_X1   g04861(.A1(new_n5053_), .A2(new_n5050_), .ZN(new_n5055_));
  AOI22_X1   g04862(.A1(\a[8] ), .A2(\a[43] ), .B1(\a[13] ), .B2(\a[38] ), .ZN(new_n5056_));
  OAI21_X1   g04863(.A1(new_n5055_), .A2(new_n5056_), .B(new_n5054_), .ZN(new_n5057_));
  NOR2_X1    g04864(.A1(new_n403_), .A2(new_n3746_), .ZN(new_n5058_));
  INV_X1     g04865(.I(new_n5058_), .ZN(new_n5059_));
  NOR2_X1    g04866(.A1(new_n3329_), .A2(new_n534_), .ZN(new_n5060_));
  NAND3_X1   g04867(.A1(new_n5058_), .A2(\a[12] ), .A3(\a[39] ), .ZN(new_n5061_));
  NAND2_X1   g04868(.A1(new_n4372_), .A2(new_n540_), .ZN(new_n5062_));
  AOI21_X1   g04869(.A1(new_n5061_), .A2(new_n5062_), .B(new_n5060_), .ZN(new_n5063_));
  AOI22_X1   g04870(.A1(\a[10] ), .A2(\a[41] ), .B1(\a[12] ), .B2(\a[39] ), .ZN(new_n5064_));
  NOR2_X1    g04871(.A1(new_n5063_), .A2(new_n5060_), .ZN(new_n5065_));
  INV_X1     g04872(.I(new_n5065_), .ZN(new_n5066_));
  OAI22_X1   g04873(.A1(new_n5066_), .A2(new_n5064_), .B1(new_n5059_), .B2(new_n5063_), .ZN(new_n5067_));
  XOR2_X1    g04874(.A1(new_n5067_), .A2(new_n5057_), .Z(new_n5068_));
  AOI21_X1   g04875(.A1(\a[24] ), .A2(\a[27] ), .B(new_n2176_), .ZN(new_n5069_));
  NAND2_X1   g04876(.A1(\a[11] ), .A2(\a[40] ), .ZN(new_n5070_));
  NOR2_X1    g04877(.A1(new_n1779_), .A2(new_n1972_), .ZN(new_n5071_));
  NOR3_X1    g04878(.A1(new_n5071_), .A2(new_n5069_), .A3(new_n5070_), .ZN(new_n5072_));
  OAI22_X1   g04879(.A1(new_n5069_), .A2(new_n5070_), .B1(new_n1779_), .B2(new_n1972_), .ZN(new_n5073_));
  OAI22_X1   g04880(.A1(new_n5072_), .A2(new_n5070_), .B1(new_n5073_), .B2(new_n5069_), .ZN(new_n5074_));
  XOR2_X1    g04881(.A1(new_n5068_), .A2(new_n5074_), .Z(new_n5075_));
  NOR2_X1    g04882(.A1(new_n1429_), .A2(new_n2526_), .ZN(new_n5076_));
  NOR4_X1    g04883(.A1(new_n253_), .A2(new_n884_), .A3(new_n2274_), .A4(new_n4178_), .ZN(new_n5077_));
  NAND4_X1   g04884(.A1(\a[5] ), .A2(\a[16] ), .A3(\a[35] ), .A4(\a[46] ), .ZN(new_n5078_));
  OAI21_X1   g04885(.A1(new_n5076_), .A2(new_n5077_), .B(new_n5078_), .ZN(new_n5079_));
  NAND3_X1   g04886(.A1(new_n5079_), .A2(\a[18] ), .A3(\a[33] ), .ZN(new_n5080_));
  AOI22_X1   g04887(.A1(\a[5] ), .A2(\a[46] ), .B1(\a[16] ), .B2(\a[35] ), .ZN(new_n5081_));
  NAND2_X1   g04888(.A1(new_n5079_), .A2(new_n5078_), .ZN(new_n5082_));
  OAI21_X1   g04889(.A1(new_n5081_), .A2(new_n5082_), .B(new_n5080_), .ZN(new_n5083_));
  NAND2_X1   g04890(.A1(new_n1767_), .A2(new_n2105_), .ZN(new_n5084_));
  OAI22_X1   g04891(.A1(new_n1301_), .A2(new_n3811_), .B1(new_n1456_), .B2(new_n2255_), .ZN(new_n5085_));
  NAND2_X1   g04892(.A1(new_n5085_), .A2(new_n5084_), .ZN(new_n5086_));
  NAND3_X1   g04893(.A1(new_n5086_), .A2(\a[21] ), .A3(\a[30] ), .ZN(new_n5087_));
  AOI22_X1   g04894(.A1(\a[22] ), .A2(\a[29] ), .B1(\a[23] ), .B2(\a[28] ), .ZN(new_n5088_));
  NAND2_X1   g04895(.A1(new_n5086_), .A2(new_n5084_), .ZN(new_n5089_));
  OAI21_X1   g04896(.A1(new_n5088_), .A2(new_n5089_), .B(new_n5087_), .ZN(new_n5090_));
  XNOR2_X1   g04897(.A1(new_n5090_), .A2(new_n5083_), .ZN(new_n5091_));
  NAND2_X1   g04898(.A1(\a[15] ), .A2(\a[36] ), .ZN(new_n5092_));
  NOR2_X1    g04899(.A1(new_n2752_), .A2(new_n4030_), .ZN(new_n5093_));
  NAND2_X1   g04900(.A1(new_n1053_), .A2(new_n5093_), .ZN(new_n5094_));
  INV_X1     g04901(.I(new_n5094_), .ZN(new_n5095_));
  NAND4_X1   g04902(.A1(\a[6] ), .A2(\a[15] ), .A3(\a[36] ), .A4(\a[45] ), .ZN(new_n5096_));
  NAND2_X1   g04903(.A1(new_n897_), .A2(new_n3037_), .ZN(new_n5097_));
  AOI21_X1   g04904(.A1(new_n5097_), .A2(new_n5096_), .B(new_n5095_), .ZN(new_n5098_));
  AOI22_X1   g04905(.A1(\a[6] ), .A2(\a[45] ), .B1(\a[14] ), .B2(\a[37] ), .ZN(new_n5099_));
  NOR2_X1    g04906(.A1(new_n5098_), .A2(new_n5095_), .ZN(new_n5100_));
  INV_X1     g04907(.I(new_n5100_), .ZN(new_n5101_));
  OAI22_X1   g04908(.A1(new_n5101_), .A2(new_n5099_), .B1(new_n5092_), .B2(new_n5098_), .ZN(new_n5102_));
  XNOR2_X1   g04909(.A1(new_n5091_), .A2(new_n5102_), .ZN(new_n5103_));
  XOR2_X1    g04910(.A1(new_n5103_), .A2(new_n5075_), .Z(new_n5104_));
  XOR2_X1    g04911(.A1(new_n5104_), .A2(new_n5048_), .Z(new_n5105_));
  NOR2_X1    g04912(.A1(new_n5030_), .A2(new_n5105_), .ZN(new_n5106_));
  NAND2_X1   g04913(.A1(new_n5030_), .A2(new_n5105_), .ZN(new_n5107_));
  INV_X1     g04914(.I(new_n5107_), .ZN(new_n5108_));
  NOR2_X1    g04915(.A1(new_n5108_), .A2(new_n5106_), .ZN(new_n5109_));
  NAND2_X1   g04916(.A1(new_n5109_), .A2(new_n5027_), .ZN(new_n5110_));
  INV_X1     g04917(.I(new_n5110_), .ZN(new_n5111_));
  NOR2_X1    g04918(.A1(new_n5109_), .A2(new_n5027_), .ZN(new_n5112_));
  NOR2_X1    g04919(.A1(new_n5111_), .A2(new_n5112_), .ZN(new_n5113_));
  XOR2_X1    g04920(.A1(new_n5024_), .A2(new_n5113_), .Z(new_n5114_));
  XOR2_X1    g04921(.A1(new_n5021_), .A2(new_n5114_), .Z(new_n5115_));
  NOR2_X1    g04922(.A1(new_n4836_), .A2(new_n4941_), .ZN(new_n5116_));
  NOR2_X1    g04923(.A1(new_n4942_), .A2(new_n4835_), .ZN(new_n5117_));
  NOR2_X1    g04924(.A1(new_n5117_), .A2(new_n5116_), .ZN(new_n5118_));
  NOR2_X1    g04925(.A1(new_n5118_), .A2(new_n5115_), .ZN(new_n5119_));
  NAND2_X1   g04926(.A1(new_n5118_), .A2(new_n5115_), .ZN(new_n5120_));
  INV_X1     g04927(.I(new_n5120_), .ZN(new_n5121_));
  NOR2_X1    g04928(.A1(new_n5121_), .A2(new_n5119_), .ZN(new_n5122_));
  XOR2_X1    g04929(.A1(new_n4953_), .A2(new_n5122_), .Z(\asquared[52] ));
  NAND2_X1   g04930(.A1(new_n5024_), .A2(new_n5113_), .ZN(new_n5124_));
  NAND3_X1   g04931(.A1(new_n5114_), .A2(new_n5020_), .A3(new_n5019_), .ZN(new_n5125_));
  NAND2_X1   g04932(.A1(new_n5125_), .A2(new_n5124_), .ZN(new_n5126_));
  INV_X1     g04933(.I(new_n5126_), .ZN(new_n5127_));
  NOR2_X1    g04934(.A1(new_n5111_), .A2(new_n5108_), .ZN(new_n5128_));
  NAND2_X1   g04935(.A1(new_n5067_), .A2(new_n5057_), .ZN(new_n5129_));
  NAND2_X1   g04936(.A1(new_n5068_), .A2(new_n5074_), .ZN(new_n5130_));
  NAND2_X1   g04937(.A1(new_n5130_), .A2(new_n5129_), .ZN(new_n5131_));
  NAND2_X1   g04938(.A1(new_n4975_), .A2(new_n4989_), .ZN(new_n5132_));
  OAI21_X1   g04939(.A1(new_n4855_), .A2(new_n4895_), .B(new_n5132_), .ZN(new_n5133_));
  NOR2_X1    g04940(.A1(new_n5036_), .A2(new_n1566_), .ZN(new_n5134_));
  INV_X1     g04941(.I(\a[51] ), .ZN(new_n5135_));
  NOR3_X1    g04942(.A1(new_n4010_), .A2(new_n194_), .A3(new_n5135_), .ZN(new_n5136_));
  AOI21_X1   g04943(.A1(\a[1] ), .A2(\a[51] ), .B(new_n2246_), .ZN(new_n5137_));
  NOR2_X1    g04944(.A1(new_n5136_), .A2(new_n5137_), .ZN(new_n5138_));
  XOR2_X1    g04945(.A1(new_n5138_), .A2(new_n5134_), .Z(new_n5139_));
  XOR2_X1    g04946(.A1(new_n5139_), .A2(new_n5073_), .Z(new_n5140_));
  XOR2_X1    g04947(.A1(new_n5133_), .A2(new_n5140_), .Z(new_n5141_));
  XOR2_X1    g04948(.A1(new_n5141_), .A2(new_n5131_), .Z(new_n5142_));
  NAND2_X1   g04949(.A1(new_n4974_), .A2(new_n4990_), .ZN(new_n5143_));
  OAI21_X1   g04950(.A1(new_n4992_), .A2(new_n4971_), .B(new_n5143_), .ZN(new_n5144_));
  NAND2_X1   g04951(.A1(new_n4876_), .A2(new_n4885_), .ZN(new_n5145_));
  NAND2_X1   g04952(.A1(new_n4959_), .A2(new_n4865_), .ZN(new_n5146_));
  NAND2_X1   g04953(.A1(new_n5146_), .A2(new_n5145_), .ZN(new_n5147_));
  NAND2_X1   g04954(.A1(new_n4917_), .A2(new_n4926_), .ZN(new_n5148_));
  NAND2_X1   g04955(.A1(new_n4954_), .A2(new_n4906_), .ZN(new_n5149_));
  NAND2_X1   g04956(.A1(new_n5149_), .A2(new_n5148_), .ZN(new_n5150_));
  AOI22_X1   g04957(.A1(\a[2] ), .A2(\a[50] ), .B1(\a[3] ), .B2(\a[49] ), .ZN(new_n5151_));
  NOR2_X1    g04958(.A1(new_n979_), .A2(new_n2274_), .ZN(new_n5152_));
  INV_X1     g04959(.I(new_n5152_), .ZN(new_n5153_));
  NOR2_X1    g04960(.A1(new_n4702_), .A2(new_n4901_), .ZN(new_n5154_));
  INV_X1     g04961(.I(new_n5154_), .ZN(new_n5155_));
  NOR2_X1    g04962(.A1(new_n5155_), .A2(new_n246_), .ZN(new_n5156_));
  NOR3_X1    g04963(.A1(new_n5156_), .A2(new_n5151_), .A3(new_n5153_), .ZN(new_n5157_));
  NOR2_X1    g04964(.A1(new_n5157_), .A2(new_n5156_), .ZN(new_n5158_));
  INV_X1     g04965(.I(new_n5158_), .ZN(new_n5159_));
  OAI22_X1   g04966(.A1(new_n5159_), .A2(new_n5151_), .B1(new_n5153_), .B2(new_n5157_), .ZN(new_n5160_));
  XOR2_X1    g04967(.A1(new_n5150_), .A2(new_n5160_), .Z(new_n5161_));
  XOR2_X1    g04968(.A1(new_n5161_), .A2(new_n5147_), .Z(new_n5162_));
  XOR2_X1    g04969(.A1(new_n5144_), .A2(new_n5162_), .Z(new_n5163_));
  XOR2_X1    g04970(.A1(new_n5163_), .A2(new_n5142_), .Z(new_n5164_));
  XNOR2_X1   g04971(.A1(new_n5128_), .A2(new_n5164_), .ZN(new_n5165_));
  NOR2_X1    g04972(.A1(new_n5001_), .A2(new_n5003_), .ZN(new_n5166_));
  NOR2_X1    g04973(.A1(new_n5006_), .A2(new_n5166_), .ZN(new_n5167_));
  NOR2_X1    g04974(.A1(new_n4771_), .A2(new_n5034_), .ZN(new_n5168_));
  NOR2_X1    g04975(.A1(new_n5035_), .A2(new_n5037_), .ZN(new_n5169_));
  NOR2_X1    g04976(.A1(new_n5169_), .A2(new_n5168_), .ZN(new_n5170_));
  NAND2_X1   g04977(.A1(new_n5170_), .A2(new_n5065_), .ZN(new_n5171_));
  NOR2_X1    g04978(.A1(new_n5170_), .A2(new_n5065_), .ZN(new_n5172_));
  INV_X1     g04979(.I(new_n5172_), .ZN(new_n5173_));
  AND2_X2    g04980(.A1(new_n5173_), .A2(new_n5171_), .Z(new_n5174_));
  INV_X1     g04981(.I(\a[52] ), .ZN(new_n5175_));
  OAI22_X1   g04982(.A1(new_n2524_), .A2(new_n814_), .B1(new_n595_), .B2(new_n4596_), .ZN(new_n5176_));
  INV_X1     g04983(.I(new_n5176_), .ZN(new_n5177_));
  NOR4_X1    g04984(.A1(new_n290_), .A2(new_n1023_), .A3(new_n2524_), .A4(new_n4596_), .ZN(new_n5178_));
  NOR3_X1    g04985(.A1(new_n5177_), .A2(new_n5175_), .A3(new_n5178_), .ZN(new_n5179_));
  NOR3_X1    g04986(.A1(new_n5179_), .A2(new_n196_), .A3(new_n5175_), .ZN(new_n5180_));
  NOR2_X1    g04987(.A1(new_n5179_), .A2(new_n5178_), .ZN(new_n5181_));
  OAI22_X1   g04988(.A1(new_n290_), .A2(new_n4596_), .B1(new_n1023_), .B2(new_n2524_), .ZN(new_n5182_));
  AOI21_X1   g04989(.A1(new_n5181_), .A2(new_n5182_), .B(new_n5180_), .ZN(new_n5183_));
  XOR2_X1    g04990(.A1(new_n5174_), .A2(new_n5183_), .Z(new_n5184_));
  INV_X1     g04991(.I(new_n5046_), .ZN(new_n5185_));
  INV_X1     g04992(.I(new_n5047_), .ZN(new_n5186_));
  NAND2_X1   g04993(.A1(new_n5186_), .A2(new_n5033_), .ZN(new_n5187_));
  OAI21_X1   g04994(.A1(new_n5038_), .A2(new_n5185_), .B(new_n5187_), .ZN(new_n5188_));
  XNOR2_X1   g04995(.A1(new_n5188_), .A2(new_n5184_), .ZN(new_n5189_));
  XNOR2_X1   g04996(.A1(new_n5167_), .A2(new_n5189_), .ZN(new_n5190_));
  NAND2_X1   g04997(.A1(new_n5104_), .A2(new_n5048_), .ZN(new_n5191_));
  NAND2_X1   g04998(.A1(new_n5103_), .A2(new_n5075_), .ZN(new_n5192_));
  NAND2_X1   g04999(.A1(new_n5191_), .A2(new_n5192_), .ZN(new_n5193_));
  XOR2_X1    g05000(.A1(new_n5082_), .A2(new_n5055_), .Z(new_n5194_));
  XOR2_X1    g05001(.A1(new_n5194_), .A2(new_n5089_), .Z(new_n5195_));
  NOR2_X1    g05002(.A1(new_n5045_), .A2(new_n4988_), .ZN(new_n5196_));
  NOR2_X1    g05003(.A1(new_n5044_), .A2(new_n4987_), .ZN(new_n5197_));
  NOR2_X1    g05004(.A1(new_n5196_), .A2(new_n5197_), .ZN(new_n5198_));
  NOR2_X1    g05005(.A1(new_n5198_), .A2(new_n5101_), .ZN(new_n5199_));
  INV_X1     g05006(.I(new_n5198_), .ZN(new_n5200_));
  NOR2_X1    g05007(.A1(new_n5200_), .A2(new_n5100_), .ZN(new_n5201_));
  NOR2_X1    g05008(.A1(new_n5201_), .A2(new_n5199_), .ZN(new_n5202_));
  NAND2_X1   g05009(.A1(new_n5090_), .A2(new_n5083_), .ZN(new_n5203_));
  INV_X1     g05010(.I(new_n5102_), .ZN(new_n5204_));
  OAI21_X1   g05011(.A1(new_n5091_), .A2(new_n5204_), .B(new_n5203_), .ZN(new_n5205_));
  NAND2_X1   g05012(.A1(new_n5205_), .A2(new_n5202_), .ZN(new_n5206_));
  INV_X1     g05013(.I(new_n5206_), .ZN(new_n5207_));
  NOR2_X1    g05014(.A1(new_n5205_), .A2(new_n5202_), .ZN(new_n5208_));
  NOR2_X1    g05015(.A1(new_n5207_), .A2(new_n5208_), .ZN(new_n5209_));
  NAND2_X1   g05016(.A1(new_n5209_), .A2(new_n5195_), .ZN(new_n5210_));
  INV_X1     g05017(.I(new_n5210_), .ZN(new_n5211_));
  NOR2_X1    g05018(.A1(new_n5209_), .A2(new_n5195_), .ZN(new_n5212_));
  NOR2_X1    g05019(.A1(new_n5211_), .A2(new_n5212_), .ZN(new_n5213_));
  XOR2_X1    g05020(.A1(new_n5193_), .A2(new_n5213_), .Z(new_n5214_));
  XNOR2_X1   g05021(.A1(new_n5190_), .A2(new_n5214_), .ZN(new_n5215_));
  XOR2_X1    g05022(.A1(new_n5165_), .A2(new_n5215_), .Z(new_n5216_));
  INV_X1     g05023(.I(new_n5216_), .ZN(new_n5217_));
  NAND2_X1   g05024(.A1(new_n4996_), .A2(new_n5016_), .ZN(new_n5218_));
  NAND2_X1   g05025(.A1(new_n5020_), .A2(new_n5218_), .ZN(new_n5219_));
  INV_X1     g05026(.I(new_n4993_), .ZN(new_n5220_));
  NOR2_X1    g05027(.A1(new_n5220_), .A2(new_n4970_), .ZN(new_n5221_));
  INV_X1     g05028(.I(new_n5221_), .ZN(new_n5222_));
  NAND2_X1   g05029(.A1(new_n4994_), .A2(new_n4968_), .ZN(new_n5223_));
  NAND2_X1   g05030(.A1(new_n5223_), .A2(new_n5222_), .ZN(new_n5224_));
  NAND2_X1   g05031(.A1(new_n5014_), .A2(new_n5011_), .ZN(new_n5225_));
  NAND2_X1   g05032(.A1(new_n5015_), .A2(new_n5008_), .ZN(new_n5226_));
  NAND2_X1   g05033(.A1(new_n5226_), .A2(new_n5225_), .ZN(new_n5227_));
  NOR2_X1    g05034(.A1(new_n4967_), .A2(new_n4963_), .ZN(new_n5228_));
  NAND2_X1   g05035(.A1(\a[5] ), .A2(\a[47] ), .ZN(new_n5229_));
  NOR3_X1    g05036(.A1(new_n1181_), .A2(new_n2626_), .A3(new_n4178_), .ZN(new_n5230_));
  NAND4_X1   g05037(.A1(\a[5] ), .A2(\a[16] ), .A3(\a[36] ), .A4(\a[47] ), .ZN(new_n5231_));
  NAND2_X1   g05038(.A1(new_n4720_), .A2(new_n746_), .ZN(new_n5232_));
  AOI21_X1   g05039(.A1(new_n5232_), .A2(new_n5231_), .B(new_n5230_), .ZN(new_n5233_));
  AOI22_X1   g05040(.A1(\a[6] ), .A2(\a[46] ), .B1(\a[16] ), .B2(\a[36] ), .ZN(new_n5234_));
  OR2_X2     g05041(.A1(new_n5233_), .A2(new_n5230_), .Z(new_n5235_));
  OAI22_X1   g05042(.A1(new_n5235_), .A2(new_n5234_), .B1(new_n5229_), .B2(new_n5233_), .ZN(new_n5236_));
  NOR2_X1    g05043(.A1(new_n417_), .A2(new_n3746_), .ZN(new_n5237_));
  INV_X1     g05044(.I(new_n5237_), .ZN(new_n5238_));
  NOR2_X1    g05045(.A1(new_n3221_), .A2(new_n3746_), .ZN(new_n5239_));
  AOI22_X1   g05046(.A1(new_n747_), .A2(new_n4372_), .B1(new_n5239_), .B2(new_n535_), .ZN(new_n5240_));
  AOI21_X1   g05047(.A1(new_n1261_), .A2(new_n4534_), .B(new_n5240_), .ZN(new_n5241_));
  AOI21_X1   g05048(.A1(\a[11] ), .A2(\a[41] ), .B(new_n4276_), .ZN(new_n5242_));
  AOI21_X1   g05049(.A1(new_n1261_), .A2(new_n4534_), .B(new_n5241_), .ZN(new_n5243_));
  INV_X1     g05050(.I(new_n5243_), .ZN(new_n5244_));
  OAI22_X1   g05051(.A1(new_n5244_), .A2(new_n5242_), .B1(new_n5238_), .B2(new_n5241_), .ZN(new_n5245_));
  XNOR2_X1   g05052(.A1(new_n5245_), .A2(new_n5236_), .ZN(new_n5246_));
  AOI22_X1   g05053(.A1(\a[7] ), .A2(\a[45] ), .B1(\a[8] ), .B2(\a[44] ), .ZN(new_n5247_));
  NAND2_X1   g05054(.A1(\a[15] ), .A2(\a[37] ), .ZN(new_n5248_));
  NOR2_X1    g05055(.A1(new_n4704_), .A2(new_n415_), .ZN(new_n5249_));
  NOR3_X1    g05056(.A1(new_n5249_), .A2(new_n5247_), .A3(new_n5248_), .ZN(new_n5250_));
  OAI22_X1   g05057(.A1(new_n4704_), .A2(new_n415_), .B1(new_n5247_), .B2(new_n5248_), .ZN(new_n5251_));
  OAI22_X1   g05058(.A1(new_n5250_), .A2(new_n5248_), .B1(new_n5247_), .B2(new_n5251_), .ZN(new_n5252_));
  XOR2_X1    g05059(.A1(new_n5246_), .A2(new_n5252_), .Z(new_n5253_));
  NOR2_X1    g05060(.A1(new_n1529_), .A2(new_n2679_), .ZN(new_n5254_));
  NOR2_X1    g05061(.A1(new_n2385_), .A2(new_n2255_), .ZN(new_n5255_));
  NOR2_X1    g05062(.A1(new_n1880_), .A2(new_n3811_), .ZN(new_n5256_));
  NOR2_X1    g05063(.A1(new_n5255_), .A2(new_n5256_), .ZN(new_n5257_));
  NOR2_X1    g05064(.A1(new_n5257_), .A2(new_n5254_), .ZN(new_n5258_));
  NAND2_X1   g05065(.A1(\a[22] ), .A2(\a[30] ), .ZN(new_n5259_));
  AOI22_X1   g05066(.A1(\a[23] ), .A2(\a[29] ), .B1(\a[24] ), .B2(\a[28] ), .ZN(new_n5260_));
  NOR2_X1    g05067(.A1(new_n5258_), .A2(new_n5254_), .ZN(new_n5261_));
  INV_X1     g05068(.I(new_n5261_), .ZN(new_n5262_));
  OAI22_X1   g05069(.A1(new_n5262_), .A2(new_n5260_), .B1(new_n5258_), .B2(new_n5259_), .ZN(new_n5263_));
  NAND2_X1   g05070(.A1(new_n1381_), .A2(new_n3210_), .ZN(new_n5264_));
  INV_X1     g05071(.I(new_n3065_), .ZN(new_n5265_));
  NOR3_X1    g05072(.A1(new_n5265_), .A2(new_n2051_), .A3(new_n2442_), .ZN(new_n5266_));
  NOR2_X1    g05073(.A1(new_n1281_), .A2(new_n3375_), .ZN(new_n5267_));
  OAI21_X1   g05074(.A1(new_n5266_), .A2(new_n5267_), .B(new_n5264_), .ZN(new_n5268_));
  NAND3_X1   g05075(.A1(new_n5268_), .A2(\a[18] ), .A3(\a[34] ), .ZN(new_n5269_));
  AOI22_X1   g05076(.A1(\a[20] ), .A2(\a[32] ), .B1(\a[21] ), .B2(\a[31] ), .ZN(new_n5270_));
  NAND2_X1   g05077(.A1(new_n5268_), .A2(new_n5264_), .ZN(new_n5271_));
  OAI21_X1   g05078(.A1(new_n5270_), .A2(new_n5271_), .B(new_n5269_), .ZN(new_n5272_));
  XOR2_X1    g05079(.A1(new_n5263_), .A2(new_n5272_), .Z(new_n5273_));
  NAND2_X1   g05080(.A1(new_n4542_), .A2(new_n5049_), .ZN(new_n5274_));
  INV_X1     g05081(.I(new_n5274_), .ZN(new_n5275_));
  NOR2_X1    g05082(.A1(new_n403_), .A2(new_n3666_), .ZN(new_n5276_));
  AOI22_X1   g05083(.A1(new_n760_), .A2(new_n4209_), .B1(new_n3560_), .B2(new_n5276_), .ZN(new_n5277_));
  NOR2_X1    g05084(.A1(new_n5275_), .A2(new_n5277_), .ZN(new_n5278_));
  AOI21_X1   g05085(.A1(\a[13] ), .A2(\a[39] ), .B(new_n5276_), .ZN(new_n5279_));
  NOR2_X1    g05086(.A1(new_n5278_), .A2(new_n5275_), .ZN(new_n5280_));
  INV_X1     g05087(.I(new_n5280_), .ZN(new_n5281_));
  OAI22_X1   g05088(.A1(new_n5281_), .A2(new_n5279_), .B1(new_n3561_), .B2(new_n5278_), .ZN(new_n5282_));
  XOR2_X1    g05089(.A1(new_n5273_), .A2(new_n5282_), .Z(new_n5283_));
  XOR2_X1    g05090(.A1(new_n5283_), .A2(new_n5253_), .Z(new_n5284_));
  XOR2_X1    g05091(.A1(new_n5228_), .A2(new_n5284_), .Z(new_n5285_));
  XOR2_X1    g05092(.A1(new_n5227_), .A2(new_n5285_), .Z(new_n5286_));
  XOR2_X1    g05093(.A1(new_n5286_), .A2(new_n5224_), .Z(new_n5287_));
  NOR2_X1    g05094(.A1(new_n5219_), .A2(new_n5287_), .ZN(new_n5288_));
  NAND2_X1   g05095(.A1(new_n5219_), .A2(new_n5287_), .ZN(new_n5289_));
  INV_X1     g05096(.I(new_n5289_), .ZN(new_n5290_));
  NOR2_X1    g05097(.A1(new_n5290_), .A2(new_n5288_), .ZN(new_n5291_));
  NOR2_X1    g05098(.A1(new_n5291_), .A2(new_n5217_), .ZN(new_n5292_));
  NAND2_X1   g05099(.A1(new_n5291_), .A2(new_n5217_), .ZN(new_n5293_));
  INV_X1     g05100(.I(new_n5293_), .ZN(new_n5294_));
  NOR2_X1    g05101(.A1(new_n5294_), .A2(new_n5292_), .ZN(new_n5295_));
  INV_X1     g05102(.I(new_n5295_), .ZN(new_n5296_));
  NOR2_X1    g05103(.A1(new_n5296_), .A2(new_n5127_), .ZN(new_n5297_));
  INV_X1     g05104(.I(new_n5297_), .ZN(new_n5298_));
  AOI21_X1   g05105(.A1(new_n4952_), .A2(new_n4944_), .B(new_n5121_), .ZN(new_n5299_));
  NOR2_X1    g05106(.A1(new_n5299_), .A2(new_n5119_), .ZN(new_n5300_));
  INV_X1     g05107(.I(new_n5119_), .ZN(new_n5301_));
  INV_X1     g05108(.I(new_n4944_), .ZN(new_n5302_));
  OAI21_X1   g05109(.A1(new_n4950_), .A2(new_n5302_), .B(new_n5120_), .ZN(new_n5303_));
  NOR2_X1    g05110(.A1(new_n5295_), .A2(new_n5126_), .ZN(new_n5304_));
  AOI21_X1   g05111(.A1(new_n5303_), .A2(new_n5301_), .B(new_n5304_), .ZN(new_n5305_));
  INV_X1     g05112(.I(new_n5304_), .ZN(new_n5306_));
  NAND2_X1   g05113(.A1(new_n5298_), .A2(new_n5306_), .ZN(new_n5307_));
  AOI22_X1   g05114(.A1(new_n5305_), .A2(new_n5298_), .B1(new_n5300_), .B2(new_n5307_), .ZN(\asquared[53] ));
  OAI21_X1   g05115(.A1(new_n5299_), .A2(new_n5119_), .B(new_n5306_), .ZN(new_n5309_));
  NAND2_X1   g05116(.A1(new_n5309_), .A2(new_n5298_), .ZN(new_n5310_));
  NOR2_X1    g05117(.A1(new_n5294_), .A2(new_n5290_), .ZN(new_n5311_));
  NAND2_X1   g05118(.A1(new_n5144_), .A2(new_n5162_), .ZN(new_n5312_));
  NAND2_X1   g05119(.A1(new_n5163_), .A2(new_n5142_), .ZN(new_n5313_));
  NAND2_X1   g05120(.A1(new_n5313_), .A2(new_n5312_), .ZN(new_n5314_));
  XOR2_X1    g05121(.A1(new_n5158_), .A2(new_n5181_), .Z(new_n5315_));
  AND2_X2    g05122(.A1(new_n5315_), .A2(new_n5262_), .Z(new_n5316_));
  NOR2_X1    g05123(.A1(new_n5315_), .A2(new_n5262_), .ZN(new_n5317_));
  NOR2_X1    g05124(.A1(new_n5316_), .A2(new_n5317_), .ZN(new_n5318_));
  NAND2_X1   g05125(.A1(new_n5263_), .A2(new_n5272_), .ZN(new_n5319_));
  NAND2_X1   g05126(.A1(new_n5273_), .A2(new_n5282_), .ZN(new_n5320_));
  NAND2_X1   g05127(.A1(new_n5320_), .A2(new_n5319_), .ZN(new_n5321_));
  INV_X1     g05128(.I(new_n5174_), .ZN(new_n5322_));
  OAI21_X1   g05129(.A1(new_n5322_), .A2(new_n5183_), .B(new_n5173_), .ZN(new_n5323_));
  XOR2_X1    g05130(.A1(new_n5321_), .A2(new_n5323_), .Z(new_n5324_));
  XNOR2_X1   g05131(.A1(new_n5324_), .A2(new_n5318_), .ZN(new_n5325_));
  XOR2_X1    g05132(.A1(new_n5235_), .A2(new_n5271_), .Z(new_n5326_));
  XOR2_X1    g05133(.A1(new_n5326_), .A2(new_n5251_), .Z(new_n5327_));
  NAND2_X1   g05134(.A1(new_n5245_), .A2(new_n5236_), .ZN(new_n5328_));
  INV_X1     g05135(.I(new_n5246_), .ZN(new_n5329_));
  NAND2_X1   g05136(.A1(new_n5329_), .A2(new_n5252_), .ZN(new_n5330_));
  NAND2_X1   g05137(.A1(new_n5330_), .A2(new_n5328_), .ZN(new_n5331_));
  NOR2_X1    g05138(.A1(new_n194_), .A2(new_n5175_), .ZN(new_n5332_));
  OAI22_X1   g05139(.A1(new_n1752_), .A2(new_n5175_), .B1(\a[27] ), .B2(new_n5332_), .ZN(new_n5333_));
  XOR2_X1    g05140(.A1(new_n5243_), .A2(new_n5333_), .Z(new_n5334_));
  NOR2_X1    g05141(.A1(new_n5334_), .A2(new_n5281_), .ZN(new_n5335_));
  NAND2_X1   g05142(.A1(new_n5334_), .A2(new_n5281_), .ZN(new_n5336_));
  INV_X1     g05143(.I(new_n5336_), .ZN(new_n5337_));
  NOR2_X1    g05144(.A1(new_n5337_), .A2(new_n5335_), .ZN(new_n5338_));
  XOR2_X1    g05145(.A1(new_n5331_), .A2(new_n5338_), .Z(new_n5339_));
  XNOR2_X1   g05146(.A1(new_n5339_), .A2(new_n5327_), .ZN(new_n5340_));
  XOR2_X1    g05147(.A1(new_n5340_), .A2(new_n5325_), .Z(new_n5341_));
  XOR2_X1    g05148(.A1(new_n5314_), .A2(new_n5341_), .Z(new_n5342_));
  INV_X1     g05149(.I(new_n5253_), .ZN(new_n5343_));
  NAND2_X1   g05150(.A1(new_n5343_), .A2(new_n5283_), .ZN(new_n5344_));
  OAI21_X1   g05151(.A1(new_n5228_), .A2(new_n5284_), .B(new_n5344_), .ZN(new_n5345_));
  INV_X1     g05152(.I(new_n5184_), .ZN(new_n5346_));
  NAND2_X1   g05153(.A1(new_n5346_), .A2(new_n5188_), .ZN(new_n5347_));
  INV_X1     g05154(.I(new_n5189_), .ZN(new_n5348_));
  OAI21_X1   g05155(.A1(new_n5348_), .A2(new_n5167_), .B(new_n5347_), .ZN(new_n5349_));
  NOR2_X1    g05156(.A1(new_n5201_), .A2(new_n5197_), .ZN(new_n5350_));
  NAND2_X1   g05157(.A1(new_n5082_), .A2(new_n5055_), .ZN(new_n5351_));
  NAND2_X1   g05158(.A1(new_n5194_), .A2(new_n5089_), .ZN(new_n5352_));
  NAND2_X1   g05159(.A1(new_n5352_), .A2(new_n5351_), .ZN(new_n5353_));
  NAND2_X1   g05160(.A1(new_n5138_), .A2(new_n5134_), .ZN(new_n5354_));
  NAND2_X1   g05161(.A1(new_n5139_), .A2(new_n5073_), .ZN(new_n5355_));
  NAND2_X1   g05162(.A1(new_n5355_), .A2(new_n5354_), .ZN(new_n5356_));
  XOR2_X1    g05163(.A1(new_n5353_), .A2(new_n5356_), .Z(new_n5357_));
  XNOR2_X1   g05164(.A1(new_n5357_), .A2(new_n5350_), .ZN(new_n5358_));
  XOR2_X1    g05165(.A1(new_n5349_), .A2(new_n5358_), .Z(new_n5359_));
  XOR2_X1    g05166(.A1(new_n5359_), .A2(new_n5345_), .Z(new_n5360_));
  NAND2_X1   g05167(.A1(new_n5227_), .A2(new_n5285_), .ZN(new_n5361_));
  NAND2_X1   g05168(.A1(new_n5286_), .A2(new_n5224_), .ZN(new_n5362_));
  NAND2_X1   g05169(.A1(new_n5362_), .A2(new_n5361_), .ZN(new_n5363_));
  XOR2_X1    g05170(.A1(new_n5363_), .A2(new_n5360_), .Z(new_n5364_));
  XNOR2_X1   g05171(.A1(new_n5364_), .A2(new_n5342_), .ZN(new_n5365_));
  OAI21_X1   g05172(.A1(new_n5111_), .A2(new_n5108_), .B(new_n5164_), .ZN(new_n5366_));
  INV_X1     g05173(.I(new_n5165_), .ZN(new_n5367_));
  OAI21_X1   g05174(.A1(new_n5367_), .A2(new_n5215_), .B(new_n5366_), .ZN(new_n5368_));
  NAND2_X1   g05175(.A1(new_n5193_), .A2(new_n5213_), .ZN(new_n5369_));
  NAND2_X1   g05176(.A1(new_n5190_), .A2(new_n5214_), .ZN(new_n5370_));
  NAND2_X1   g05177(.A1(new_n5370_), .A2(new_n5369_), .ZN(new_n5371_));
  NOR2_X1    g05178(.A1(new_n5211_), .A2(new_n5207_), .ZN(new_n5372_));
  NAND2_X1   g05179(.A1(new_n5133_), .A2(new_n5140_), .ZN(new_n5373_));
  NAND2_X1   g05180(.A1(new_n5141_), .A2(new_n5131_), .ZN(new_n5374_));
  NAND2_X1   g05181(.A1(new_n5374_), .A2(new_n5373_), .ZN(new_n5375_));
  NAND2_X1   g05182(.A1(new_n4028_), .A2(new_n535_), .ZN(new_n5376_));
  INV_X1     g05183(.I(new_n4534_), .ZN(new_n5377_));
  NAND2_X1   g05184(.A1(new_n4893_), .A2(new_n5049_), .ZN(new_n5378_));
  OAI21_X1   g05185(.A1(new_n1265_), .A2(new_n5377_), .B(new_n5378_), .ZN(new_n5379_));
  NAND2_X1   g05186(.A1(new_n5379_), .A2(new_n5376_), .ZN(new_n5380_));
  NAND3_X1   g05187(.A1(new_n5380_), .A2(\a[13] ), .A3(\a[40] ), .ZN(new_n5381_));
  AOI22_X1   g05188(.A1(\a[10] ), .A2(\a[43] ), .B1(\a[12] ), .B2(\a[41] ), .ZN(new_n5382_));
  NAND2_X1   g05189(.A1(new_n5380_), .A2(new_n5376_), .ZN(new_n5383_));
  OAI21_X1   g05190(.A1(new_n5382_), .A2(new_n5383_), .B(new_n5381_), .ZN(new_n5384_));
  NAND2_X1   g05191(.A1(new_n1767_), .A2(new_n2437_), .ZN(new_n5385_));
  NAND2_X1   g05192(.A1(new_n1879_), .A2(new_n2976_), .ZN(new_n5386_));
  AOI22_X1   g05193(.A1(new_n5385_), .A2(new_n5386_), .B1(new_n1528_), .B2(new_n2254_), .ZN(new_n5387_));
  AOI22_X1   g05194(.A1(\a[23] ), .A2(\a[30] ), .B1(\a[24] ), .B2(\a[29] ), .ZN(new_n5388_));
  NAND2_X1   g05195(.A1(new_n1528_), .A2(new_n2254_), .ZN(new_n5389_));
  NAND3_X1   g05196(.A1(new_n5389_), .A2(new_n5385_), .A3(new_n5386_), .ZN(new_n5390_));
  OAI22_X1   g05197(.A1(new_n5387_), .A2(new_n2053_), .B1(new_n5390_), .B2(new_n5388_), .ZN(new_n5391_));
  XNOR2_X1   g05198(.A1(new_n5384_), .A2(new_n5391_), .ZN(new_n5392_));
  AOI21_X1   g05199(.A1(\a[25] ), .A2(\a[28] ), .B(new_n1971_), .ZN(new_n5393_));
  NAND2_X1   g05200(.A1(\a[11] ), .A2(\a[42] ), .ZN(new_n5394_));
  NOR2_X1    g05201(.A1(new_n2189_), .A2(new_n2177_), .ZN(new_n5395_));
  NOR3_X1    g05202(.A1(new_n5395_), .A2(new_n5393_), .A3(new_n5394_), .ZN(new_n5396_));
  OAI22_X1   g05203(.A1(new_n5393_), .A2(new_n5394_), .B1(new_n2189_), .B2(new_n2177_), .ZN(new_n5397_));
  OAI22_X1   g05204(.A1(new_n5396_), .A2(new_n5394_), .B1(new_n5397_), .B2(new_n5393_), .ZN(new_n5398_));
  XOR2_X1    g05205(.A1(new_n5392_), .A2(new_n5398_), .Z(new_n5399_));
  INV_X1     g05206(.I(new_n5399_), .ZN(new_n5400_));
  XOR2_X1    g05207(.A1(new_n5375_), .A2(new_n5400_), .Z(new_n5401_));
  XNOR2_X1   g05208(.A1(new_n5372_), .A2(new_n5401_), .ZN(new_n5402_));
  NOR4_X1    g05209(.A1(new_n355_), .A2(new_n759_), .A3(new_n3116_), .A4(new_n4030_), .ZN(new_n5403_));
  NOR2_X1    g05210(.A1(new_n4704_), .A2(new_n1427_), .ZN(new_n5404_));
  NOR2_X1    g05211(.A1(new_n759_), .A2(new_n3859_), .ZN(new_n5405_));
  NAND2_X1   g05212(.A1(new_n4542_), .A2(new_n5405_), .ZN(new_n5406_));
  OAI21_X1   g05213(.A1(new_n5404_), .A2(new_n5403_), .B(new_n5406_), .ZN(new_n5407_));
  NAND3_X1   g05214(.A1(new_n5407_), .A2(\a[8] ), .A3(\a[45] ), .ZN(new_n5408_));
  AOI22_X1   g05215(.A1(\a[9] ), .A2(\a[44] ), .B1(\a[14] ), .B2(\a[39] ), .ZN(new_n5409_));
  NAND2_X1   g05216(.A1(new_n5407_), .A2(new_n5406_), .ZN(new_n5410_));
  OAI21_X1   g05217(.A1(new_n5409_), .A2(new_n5410_), .B(new_n5408_), .ZN(new_n5411_));
  NOR2_X1    g05218(.A1(new_n422_), .A2(new_n4178_), .ZN(new_n5412_));
  NOR2_X1    g05219(.A1(new_n3563_), .A2(new_n5412_), .ZN(new_n5413_));
  NAND2_X1   g05220(.A1(new_n3563_), .A2(new_n5412_), .ZN(new_n5414_));
  NOR2_X1    g05221(.A1(new_n367_), .A2(new_n4312_), .ZN(new_n5415_));
  NAND2_X1   g05222(.A1(new_n3563_), .A2(new_n5415_), .ZN(new_n5416_));
  OAI21_X1   g05223(.A1(new_n374_), .A2(new_n4721_), .B(new_n5416_), .ZN(new_n5417_));
  NAND2_X1   g05224(.A1(new_n5417_), .A2(new_n5414_), .ZN(new_n5418_));
  NAND2_X1   g05225(.A1(new_n5418_), .A2(new_n5414_), .ZN(new_n5419_));
  NAND2_X1   g05226(.A1(new_n5418_), .A2(new_n5415_), .ZN(new_n5420_));
  OAI21_X1   g05227(.A1(new_n5413_), .A2(new_n5419_), .B(new_n5420_), .ZN(new_n5421_));
  XNOR2_X1   g05228(.A1(new_n5421_), .A2(new_n5411_), .ZN(new_n5422_));
  AOI22_X1   g05229(.A1(\a[5] ), .A2(\a[48] ), .B1(\a[16] ), .B2(\a[37] ), .ZN(new_n5423_));
  INV_X1     g05230(.I(new_n5423_), .ZN(new_n5424_));
  INV_X1     g05231(.I(\a[53] ), .ZN(new_n5425_));
  NOR2_X1    g05232(.A1(new_n196_), .A2(new_n5425_), .ZN(new_n5426_));
  NOR4_X1    g05233(.A1(new_n253_), .A2(new_n742_), .A3(new_n2752_), .A4(new_n4596_), .ZN(new_n5427_));
  INV_X1     g05234(.I(new_n5427_), .ZN(new_n5428_));
  NOR3_X1    g05235(.A1(new_n5423_), .A2(new_n196_), .A3(new_n5425_), .ZN(new_n5429_));
  NAND2_X1   g05236(.A1(new_n5428_), .A2(new_n5429_), .ZN(new_n5430_));
  NOR2_X1    g05237(.A1(new_n5429_), .A2(new_n5427_), .ZN(new_n5431_));
  AOI22_X1   g05238(.A1(new_n5430_), .A2(new_n5426_), .B1(new_n5431_), .B2(new_n5424_), .ZN(new_n5432_));
  XNOR2_X1   g05239(.A1(new_n5422_), .A2(new_n5432_), .ZN(new_n5433_));
  NAND2_X1   g05240(.A1(new_n5150_), .A2(new_n5160_), .ZN(new_n5434_));
  NAND2_X1   g05241(.A1(new_n5161_), .A2(new_n5147_), .ZN(new_n5435_));
  NAND2_X1   g05242(.A1(new_n5435_), .A2(new_n5434_), .ZN(new_n5436_));
  AOI22_X1   g05243(.A1(\a[2] ), .A2(\a[51] ), .B1(\a[3] ), .B2(\a[50] ), .ZN(new_n5437_));
  INV_X1     g05244(.I(new_n5437_), .ZN(new_n5438_));
  NOR2_X1    g05245(.A1(new_n4901_), .A2(new_n5135_), .ZN(new_n5439_));
  INV_X1     g05246(.I(new_n5439_), .ZN(new_n5440_));
  NOR2_X1    g05247(.A1(new_n5440_), .A2(new_n246_), .ZN(new_n5441_));
  AOI21_X1   g05248(.A1(new_n5136_), .A2(new_n5438_), .B(new_n5441_), .ZN(new_n5442_));
  INV_X1     g05249(.I(new_n5442_), .ZN(new_n5443_));
  OAI21_X1   g05250(.A1(new_n5437_), .A2(new_n5441_), .B(new_n5136_), .ZN(new_n5444_));
  OAI21_X1   g05251(.A1(new_n5443_), .A2(new_n5437_), .B(new_n5444_), .ZN(new_n5445_));
  AOI22_X1   g05252(.A1(\a[17] ), .A2(\a[36] ), .B1(\a[18] ), .B2(\a[35] ), .ZN(new_n5446_));
  INV_X1     g05253(.I(new_n5446_), .ZN(new_n5447_));
  NOR2_X1    g05254(.A1(new_n1275_), .A2(new_n3405_), .ZN(new_n5448_));
  NOR2_X1    g05255(.A1(new_n290_), .A2(new_n4702_), .ZN(new_n5449_));
  AOI21_X1   g05256(.A1(new_n5447_), .A2(new_n5449_), .B(new_n5448_), .ZN(new_n5450_));
  INV_X1     g05257(.I(new_n5450_), .ZN(new_n5451_));
  OAI21_X1   g05258(.A1(new_n5448_), .A2(new_n5446_), .B(new_n5449_), .ZN(new_n5452_));
  OAI21_X1   g05259(.A1(new_n5451_), .A2(new_n5446_), .B(new_n5452_), .ZN(new_n5453_));
  XOR2_X1    g05260(.A1(new_n5453_), .A2(new_n5445_), .Z(new_n5454_));
  OAI22_X1   g05261(.A1(new_n1376_), .A2(new_n3932_), .B1(new_n1379_), .B2(new_n3375_), .ZN(new_n5455_));
  OAI21_X1   g05262(.A1(new_n1382_), .A2(new_n2637_), .B(new_n5455_), .ZN(new_n5456_));
  NAND3_X1   g05263(.A1(new_n5456_), .A2(\a[19] ), .A3(\a[34] ), .ZN(new_n5457_));
  AOI22_X1   g05264(.A1(\a[20] ), .A2(\a[33] ), .B1(\a[21] ), .B2(\a[32] ), .ZN(new_n5458_));
  NOR2_X1    g05265(.A1(new_n1382_), .A2(new_n2637_), .ZN(new_n5459_));
  NOR2_X1    g05266(.A1(new_n5455_), .A2(new_n5459_), .ZN(new_n5460_));
  INV_X1     g05267(.I(new_n5460_), .ZN(new_n5461_));
  OAI21_X1   g05268(.A1(new_n5458_), .A2(new_n5461_), .B(new_n5457_), .ZN(new_n5462_));
  XOR2_X1    g05269(.A1(new_n5454_), .A2(new_n5462_), .Z(new_n5463_));
  XOR2_X1    g05270(.A1(new_n5436_), .A2(new_n5463_), .Z(new_n5464_));
  XOR2_X1    g05271(.A1(new_n5464_), .A2(new_n5433_), .Z(new_n5465_));
  XNOR2_X1   g05272(.A1(new_n5402_), .A2(new_n5465_), .ZN(new_n5466_));
  NOR2_X1    g05273(.A1(new_n5466_), .A2(new_n5371_), .ZN(new_n5467_));
  NAND2_X1   g05274(.A1(new_n5466_), .A2(new_n5371_), .ZN(new_n5468_));
  INV_X1     g05275(.I(new_n5468_), .ZN(new_n5469_));
  NOR2_X1    g05276(.A1(new_n5469_), .A2(new_n5467_), .ZN(new_n5470_));
  NOR2_X1    g05277(.A1(new_n5368_), .A2(new_n5470_), .ZN(new_n5471_));
  NAND2_X1   g05278(.A1(new_n5368_), .A2(new_n5470_), .ZN(new_n5472_));
  INV_X1     g05279(.I(new_n5472_), .ZN(new_n5473_));
  NOR2_X1    g05280(.A1(new_n5473_), .A2(new_n5471_), .ZN(new_n5474_));
  XNOR2_X1   g05281(.A1(new_n5474_), .A2(new_n5365_), .ZN(new_n5475_));
  INV_X1     g05282(.I(new_n5475_), .ZN(new_n5476_));
  NOR2_X1    g05283(.A1(new_n5311_), .A2(new_n5476_), .ZN(new_n5477_));
  NAND2_X1   g05284(.A1(new_n5311_), .A2(new_n5476_), .ZN(new_n5478_));
  INV_X1     g05285(.I(new_n5478_), .ZN(new_n5479_));
  NOR2_X1    g05286(.A1(new_n5479_), .A2(new_n5477_), .ZN(new_n5480_));
  XOR2_X1    g05287(.A1(new_n5310_), .A2(new_n5480_), .Z(\asquared[54] ));
  AOI21_X1   g05288(.A1(new_n5309_), .A2(new_n5298_), .B(new_n5479_), .ZN(new_n5482_));
  NOR2_X1    g05289(.A1(new_n5482_), .A2(new_n5477_), .ZN(new_n5483_));
  INV_X1     g05290(.I(new_n5474_), .ZN(new_n5484_));
  NOR2_X1    g05291(.A1(new_n5484_), .A2(new_n5365_), .ZN(new_n5485_));
  NOR2_X1    g05292(.A1(new_n5485_), .A2(new_n5473_), .ZN(new_n5486_));
  INV_X1     g05293(.I(new_n5486_), .ZN(new_n5487_));
  INV_X1     g05294(.I(new_n5402_), .ZN(new_n5488_));
  NOR2_X1    g05295(.A1(new_n5488_), .A2(new_n5465_), .ZN(new_n5489_));
  NOR2_X1    g05296(.A1(new_n5469_), .A2(new_n5489_), .ZN(new_n5490_));
  XNOR2_X1   g05297(.A1(new_n5419_), .A2(new_n5431_), .ZN(new_n5491_));
  XOR2_X1    g05298(.A1(new_n5491_), .A2(new_n5397_), .Z(new_n5492_));
  NAND2_X1   g05299(.A1(new_n5421_), .A2(new_n5411_), .ZN(new_n5493_));
  OAI21_X1   g05300(.A1(new_n5422_), .A2(new_n5432_), .B(new_n5493_), .ZN(new_n5494_));
  XOR2_X1    g05301(.A1(new_n5450_), .A2(new_n5460_), .Z(new_n5495_));
  XOR2_X1    g05302(.A1(new_n5495_), .A2(new_n5390_), .Z(new_n5496_));
  NOR2_X1    g05303(.A1(new_n5494_), .A2(new_n5496_), .ZN(new_n5497_));
  AND2_X2    g05304(.A1(new_n5494_), .A2(new_n5496_), .Z(new_n5498_));
  NOR2_X1    g05305(.A1(new_n5498_), .A2(new_n5497_), .ZN(new_n5499_));
  AND2_X2    g05306(.A1(new_n5499_), .A2(new_n5492_), .Z(new_n5500_));
  NOR2_X1    g05307(.A1(new_n5499_), .A2(new_n5492_), .ZN(new_n5501_));
  NOR2_X1    g05308(.A1(new_n5500_), .A2(new_n5501_), .ZN(new_n5502_));
  NOR2_X1    g05309(.A1(new_n5436_), .A2(new_n5463_), .ZN(new_n5503_));
  NAND2_X1   g05310(.A1(new_n5436_), .A2(new_n5463_), .ZN(new_n5504_));
  OAI21_X1   g05311(.A1(new_n5433_), .A2(new_n5503_), .B(new_n5504_), .ZN(new_n5505_));
  NOR2_X1    g05312(.A1(new_n5243_), .A2(new_n5333_), .ZN(new_n5506_));
  NOR2_X1    g05313(.A1(new_n5337_), .A2(new_n5506_), .ZN(new_n5507_));
  NAND2_X1   g05314(.A1(new_n5235_), .A2(new_n5271_), .ZN(new_n5508_));
  NAND2_X1   g05315(.A1(new_n5326_), .A2(new_n5251_), .ZN(new_n5509_));
  NAND2_X1   g05316(.A1(new_n5509_), .A2(new_n5508_), .ZN(new_n5510_));
  NOR2_X1    g05317(.A1(new_n5158_), .A2(new_n5181_), .ZN(new_n5511_));
  NOR2_X1    g05318(.A1(new_n5316_), .A2(new_n5511_), .ZN(new_n5512_));
  XNOR2_X1   g05319(.A1(new_n5510_), .A2(new_n5512_), .ZN(new_n5513_));
  XNOR2_X1   g05320(.A1(new_n5513_), .A2(new_n5507_), .ZN(new_n5514_));
  XOR2_X1    g05321(.A1(new_n5505_), .A2(new_n5514_), .Z(new_n5515_));
  XOR2_X1    g05322(.A1(new_n5515_), .A2(new_n5502_), .Z(new_n5516_));
  INV_X1     g05323(.I(new_n5516_), .ZN(new_n5517_));
  NAND2_X1   g05324(.A1(new_n5490_), .A2(new_n5517_), .ZN(new_n5518_));
  OAI21_X1   g05325(.A1(new_n5469_), .A2(new_n5489_), .B(new_n5516_), .ZN(new_n5519_));
  AND2_X2    g05326(.A1(new_n5518_), .A2(new_n5519_), .Z(new_n5520_));
  NAND2_X1   g05327(.A1(new_n5439_), .A2(new_n761_), .ZN(new_n5521_));
  NOR2_X1    g05328(.A1(new_n4901_), .A2(new_n5175_), .ZN(new_n5522_));
  INV_X1     g05329(.I(new_n5522_), .ZN(new_n5523_));
  NOR2_X1    g05330(.A1(new_n5135_), .A2(new_n5175_), .ZN(new_n5524_));
  INV_X1     g05331(.I(new_n5524_), .ZN(new_n5525_));
  OAI22_X1   g05332(.A1(new_n246_), .A2(new_n5525_), .B1(new_n5523_), .B2(new_n251_), .ZN(new_n5526_));
  NAND2_X1   g05333(.A1(new_n5526_), .A2(new_n5521_), .ZN(new_n5527_));
  NAND3_X1   g05334(.A1(new_n5527_), .A2(\a[2] ), .A3(\a[52] ), .ZN(new_n5528_));
  AOI22_X1   g05335(.A1(\a[3] ), .A2(\a[51] ), .B1(\a[4] ), .B2(\a[50] ), .ZN(new_n5529_));
  NAND2_X1   g05336(.A1(new_n5527_), .A2(new_n5521_), .ZN(new_n5530_));
  OAI21_X1   g05337(.A1(new_n5529_), .A2(new_n5530_), .B(new_n5528_), .ZN(new_n5531_));
  NOR2_X1    g05338(.A1(new_n422_), .A2(new_n4312_), .ZN(new_n5532_));
  NOR2_X1    g05339(.A1(new_n717_), .A2(new_n3116_), .ZN(new_n5533_));
  INV_X1     g05340(.I(new_n5533_), .ZN(new_n5534_));
  NOR3_X1    g05341(.A1(new_n5534_), .A2(new_n355_), .A3(new_n4178_), .ZN(new_n5535_));
  AOI22_X1   g05342(.A1(new_n5532_), .A2(new_n5533_), .B1(new_n4720_), .B2(new_n693_), .ZN(new_n5536_));
  OAI21_X1   g05343(.A1(new_n5535_), .A2(new_n5536_), .B(new_n5532_), .ZN(new_n5537_));
  AOI21_X1   g05344(.A1(\a[8] ), .A2(\a[46] ), .B(new_n5533_), .ZN(new_n5538_));
  INV_X1     g05345(.I(new_n5535_), .ZN(new_n5539_));
  NAND2_X1   g05346(.A1(new_n5539_), .A2(new_n5536_), .ZN(new_n5540_));
  OAI21_X1   g05347(.A1(new_n5540_), .A2(new_n5538_), .B(new_n5537_), .ZN(new_n5541_));
  XNOR2_X1   g05348(.A1(new_n5531_), .A2(new_n5541_), .ZN(new_n5542_));
  NOR2_X1    g05349(.A1(new_n403_), .A2(new_n4030_), .ZN(new_n5543_));
  INV_X1     g05350(.I(new_n5543_), .ZN(new_n5544_));
  NAND2_X1   g05351(.A1(new_n4019_), .A2(new_n5543_), .ZN(new_n5545_));
  NAND2_X1   g05352(.A1(new_n4703_), .A2(new_n540_), .ZN(new_n5546_));
  AOI22_X1   g05353(.A1(new_n5545_), .A2(new_n5546_), .B1(new_n4893_), .B2(new_n5405_), .ZN(new_n5547_));
  NAND2_X1   g05354(.A1(new_n4893_), .A2(new_n5405_), .ZN(new_n5548_));
  NAND3_X1   g05355(.A1(new_n5548_), .A2(new_n5545_), .A3(new_n5546_), .ZN(new_n5549_));
  AOI21_X1   g05356(.A1(\a[10] ), .A2(\a[44] ), .B(new_n4019_), .ZN(new_n5550_));
  OAI22_X1   g05357(.A1(new_n5547_), .A2(new_n5544_), .B1(new_n5549_), .B2(new_n5550_), .ZN(new_n5551_));
  XOR2_X1    g05358(.A1(new_n5542_), .A2(new_n5551_), .Z(new_n5552_));
  INV_X1     g05359(.I(new_n5552_), .ZN(new_n5553_));
  NOR2_X1    g05360(.A1(new_n1265_), .A2(new_n4667_), .ZN(new_n5554_));
  AOI21_X1   g05361(.A1(new_n834_), .A2(new_n4028_), .B(new_n5554_), .ZN(new_n5555_));
  AOI21_X1   g05362(.A1(new_n1261_), .A2(new_n4180_), .B(new_n5555_), .ZN(new_n5556_));
  NAND2_X1   g05363(.A1(\a[13] ), .A2(\a[41] ), .ZN(new_n5557_));
  AOI22_X1   g05364(.A1(\a[11] ), .A2(\a[43] ), .B1(\a[12] ), .B2(\a[42] ), .ZN(new_n5558_));
  NOR2_X1    g05365(.A1(new_n4181_), .A2(new_n619_), .ZN(new_n5559_));
  NOR2_X1    g05366(.A1(new_n5556_), .A2(new_n5559_), .ZN(new_n5560_));
  INV_X1     g05367(.I(new_n5560_), .ZN(new_n5561_));
  OAI22_X1   g05368(.A1(new_n5561_), .A2(new_n5558_), .B1(new_n5556_), .B2(new_n5557_), .ZN(new_n5562_));
  NAND4_X1   g05369(.A1(\a[5] ), .A2(\a[18] ), .A3(\a[36] ), .A4(\a[49] ), .ZN(new_n5563_));
  INV_X1     g05370(.I(new_n3822_), .ZN(new_n5564_));
  NOR2_X1    g05371(.A1(new_n1043_), .A2(new_n4702_), .ZN(new_n5565_));
  INV_X1     g05372(.I(new_n5565_), .ZN(new_n5566_));
  OAI22_X1   g05373(.A1(new_n1281_), .A2(new_n5564_), .B1(new_n4847_), .B2(new_n5566_), .ZN(new_n5567_));
  NAND2_X1   g05374(.A1(new_n5567_), .A2(new_n5563_), .ZN(new_n5568_));
  NAND3_X1   g05375(.A1(new_n5568_), .A2(\a[20] ), .A3(\a[34] ), .ZN(new_n5569_));
  NAND2_X1   g05376(.A1(new_n5568_), .A2(new_n5563_), .ZN(new_n5570_));
  AOI22_X1   g05377(.A1(\a[5] ), .A2(\a[49] ), .B1(\a[18] ), .B2(\a[36] ), .ZN(new_n5571_));
  OAI21_X1   g05378(.A1(new_n5570_), .A2(new_n5571_), .B(new_n5569_), .ZN(new_n5572_));
  XOR2_X1    g05379(.A1(new_n5562_), .A2(new_n5572_), .Z(new_n5573_));
  NOR2_X1    g05380(.A1(new_n2914_), .A2(new_n4596_), .ZN(new_n5574_));
  NOR2_X1    g05381(.A1(new_n1023_), .A2(new_n4596_), .ZN(new_n5575_));
  NAND2_X1   g05382(.A1(new_n3641_), .A2(new_n5575_), .ZN(new_n5576_));
  NAND2_X1   g05383(.A1(new_n1024_), .A2(new_n3803_), .ZN(new_n5577_));
  AOI22_X1   g05384(.A1(new_n5576_), .A2(new_n5577_), .B1(new_n743_), .B2(new_n5574_), .ZN(new_n5578_));
  NAND2_X1   g05385(.A1(\a[17] ), .A2(\a[37] ), .ZN(new_n5579_));
  AOI22_X1   g05386(.A1(\a[6] ), .A2(\a[48] ), .B1(\a[16] ), .B2(\a[38] ), .ZN(new_n5580_));
  NAND2_X1   g05387(.A1(new_n743_), .A2(new_n5574_), .ZN(new_n5581_));
  NAND3_X1   g05388(.A1(new_n5581_), .A2(new_n5576_), .A3(new_n5577_), .ZN(new_n5582_));
  OAI22_X1   g05389(.A1(new_n5578_), .A2(new_n5579_), .B1(new_n5582_), .B2(new_n5580_), .ZN(new_n5583_));
  XOR2_X1    g05390(.A1(new_n5573_), .A2(new_n5583_), .Z(new_n5584_));
  NAND2_X1   g05391(.A1(new_n5353_), .A2(new_n5356_), .ZN(new_n5585_));
  INV_X1     g05392(.I(new_n5357_), .ZN(new_n5586_));
  OAI21_X1   g05393(.A1(new_n5586_), .A2(new_n5350_), .B(new_n5585_), .ZN(new_n5587_));
  XOR2_X1    g05394(.A1(new_n5584_), .A2(new_n5587_), .Z(new_n5588_));
  XOR2_X1    g05395(.A1(new_n5588_), .A2(new_n5553_), .Z(new_n5589_));
  NAND2_X1   g05396(.A1(new_n5375_), .A2(new_n5400_), .ZN(new_n5590_));
  INV_X1     g05397(.I(new_n5401_), .ZN(new_n5591_));
  OAI21_X1   g05398(.A1(new_n5591_), .A2(new_n5372_), .B(new_n5590_), .ZN(new_n5592_));
  XOR2_X1    g05399(.A1(new_n5410_), .A2(new_n5443_), .Z(new_n5593_));
  XOR2_X1    g05400(.A1(new_n5593_), .A2(new_n5383_), .Z(new_n5594_));
  NAND2_X1   g05401(.A1(new_n5384_), .A2(new_n5391_), .ZN(new_n5595_));
  INV_X1     g05402(.I(new_n5392_), .ZN(new_n5596_));
  NAND2_X1   g05403(.A1(new_n5596_), .A2(new_n5398_), .ZN(new_n5597_));
  NAND2_X1   g05404(.A1(new_n5597_), .A2(new_n5595_), .ZN(new_n5598_));
  NAND2_X1   g05405(.A1(new_n5453_), .A2(new_n5445_), .ZN(new_n5599_));
  NAND2_X1   g05406(.A1(new_n5454_), .A2(new_n5462_), .ZN(new_n5600_));
  NAND2_X1   g05407(.A1(new_n5600_), .A2(new_n5599_), .ZN(new_n5601_));
  XOR2_X1    g05408(.A1(new_n5598_), .A2(new_n5601_), .Z(new_n5602_));
  XOR2_X1    g05409(.A1(new_n5602_), .A2(new_n5594_), .Z(new_n5603_));
  XOR2_X1    g05410(.A1(new_n5592_), .A2(new_n5603_), .Z(new_n5604_));
  XNOR2_X1   g05411(.A1(new_n5604_), .A2(new_n5589_), .ZN(new_n5605_));
  XOR2_X1    g05412(.A1(new_n5520_), .A2(new_n5605_), .Z(new_n5606_));
  NAND2_X1   g05413(.A1(new_n5314_), .A2(new_n5341_), .ZN(new_n5607_));
  OAI21_X1   g05414(.A1(new_n5325_), .A2(new_n5340_), .B(new_n5607_), .ZN(new_n5608_));
  NAND2_X1   g05415(.A1(new_n5349_), .A2(new_n5358_), .ZN(new_n5609_));
  NAND2_X1   g05416(.A1(new_n5359_), .A2(new_n5345_), .ZN(new_n5610_));
  NAND2_X1   g05417(.A1(new_n5610_), .A2(new_n5609_), .ZN(new_n5611_));
  XOR2_X1    g05418(.A1(new_n5608_), .A2(new_n5611_), .Z(new_n5612_));
  NAND2_X1   g05419(.A1(new_n5321_), .A2(new_n5323_), .ZN(new_n5613_));
  NAND2_X1   g05420(.A1(new_n5324_), .A2(new_n5318_), .ZN(new_n5614_));
  NAND2_X1   g05421(.A1(new_n5614_), .A2(new_n5613_), .ZN(new_n5615_));
  NOR2_X1    g05422(.A1(new_n1752_), .A2(new_n5175_), .ZN(new_n5616_));
  INV_X1     g05423(.I(\a[54] ), .ZN(new_n5617_));
  NOR2_X1    g05424(.A1(new_n196_), .A2(new_n5617_), .ZN(new_n5618_));
  XOR2_X1    g05425(.A1(new_n5616_), .A2(new_n5618_), .Z(new_n5619_));
  NAND2_X1   g05426(.A1(\a[1] ), .A2(\a[53] ), .ZN(new_n5620_));
  XNOR2_X1   g05427(.A1(new_n2412_), .A2(new_n5620_), .ZN(new_n5621_));
  XNOR2_X1   g05428(.A1(new_n5619_), .A2(new_n5621_), .ZN(new_n5622_));
  INV_X1     g05429(.I(new_n5622_), .ZN(new_n5623_));
  NAND2_X1   g05430(.A1(new_n1778_), .A2(new_n2254_), .ZN(new_n5624_));
  INV_X1     g05431(.I(new_n2976_), .ZN(new_n5625_));
  OAI22_X1   g05432(.A1(new_n1443_), .A2(new_n5625_), .B1(new_n1529_), .B2(new_n2438_), .ZN(new_n5626_));
  NAND2_X1   g05433(.A1(new_n5626_), .A2(new_n5624_), .ZN(new_n5627_));
  NAND3_X1   g05434(.A1(new_n5627_), .A2(\a[23] ), .A3(\a[31] ), .ZN(new_n5628_));
  AOI22_X1   g05435(.A1(\a[24] ), .A2(\a[30] ), .B1(\a[25] ), .B2(\a[29] ), .ZN(new_n5629_));
  NAND2_X1   g05436(.A1(new_n5627_), .A2(new_n5624_), .ZN(new_n5630_));
  OAI21_X1   g05437(.A1(new_n5629_), .A2(new_n5630_), .B(new_n5628_), .ZN(new_n5631_));
  NAND2_X1   g05438(.A1(new_n1452_), .A2(new_n2636_), .ZN(new_n5632_));
  NOR2_X1    g05439(.A1(new_n2200_), .A2(new_n2524_), .ZN(new_n5633_));
  INV_X1     g05440(.I(new_n5633_), .ZN(new_n5634_));
  OAI22_X1   g05441(.A1(new_n1379_), .A2(new_n2526_), .B1(new_n3394_), .B2(new_n5634_), .ZN(new_n5635_));
  NAND2_X1   g05442(.A1(new_n5635_), .A2(new_n5632_), .ZN(new_n5636_));
  NAND3_X1   g05443(.A1(new_n5636_), .A2(\a[19] ), .A3(\a[35] ), .ZN(new_n5637_));
  AOI22_X1   g05444(.A1(\a[21] ), .A2(\a[33] ), .B1(\a[22] ), .B2(\a[32] ), .ZN(new_n5638_));
  NAND2_X1   g05445(.A1(new_n5636_), .A2(new_n5632_), .ZN(new_n5639_));
  OAI21_X1   g05446(.A1(new_n5638_), .A2(new_n5639_), .B(new_n5637_), .ZN(new_n5640_));
  XNOR2_X1   g05447(.A1(new_n5631_), .A2(new_n5640_), .ZN(new_n5641_));
  XOR2_X1    g05448(.A1(new_n5641_), .A2(new_n5623_), .Z(new_n5642_));
  XOR2_X1    g05449(.A1(new_n5615_), .A2(new_n5642_), .Z(new_n5643_));
  NAND2_X1   g05450(.A1(new_n5331_), .A2(new_n5338_), .ZN(new_n5644_));
  NAND2_X1   g05451(.A1(new_n5339_), .A2(new_n5327_), .ZN(new_n5645_));
  NAND2_X1   g05452(.A1(new_n5645_), .A2(new_n5644_), .ZN(new_n5646_));
  XOR2_X1    g05453(.A1(new_n5643_), .A2(new_n5646_), .Z(new_n5647_));
  XOR2_X1    g05454(.A1(new_n5612_), .A2(new_n5647_), .Z(new_n5648_));
  NAND2_X1   g05455(.A1(new_n5363_), .A2(new_n5360_), .ZN(new_n5649_));
  NAND2_X1   g05456(.A1(new_n5364_), .A2(new_n5342_), .ZN(new_n5650_));
  NAND2_X1   g05457(.A1(new_n5650_), .A2(new_n5649_), .ZN(new_n5651_));
  XOR2_X1    g05458(.A1(new_n5651_), .A2(new_n5648_), .Z(new_n5652_));
  XNOR2_X1   g05459(.A1(new_n5652_), .A2(new_n5606_), .ZN(new_n5653_));
  INV_X1     g05460(.I(new_n5653_), .ZN(new_n5654_));
  NOR2_X1    g05461(.A1(new_n5487_), .A2(new_n5654_), .ZN(new_n5655_));
  INV_X1     g05462(.I(new_n5655_), .ZN(new_n5656_));
  NOR2_X1    g05463(.A1(new_n5486_), .A2(new_n5653_), .ZN(new_n5657_));
  INV_X1     g05464(.I(new_n5657_), .ZN(new_n5658_));
  NAND2_X1   g05465(.A1(new_n5656_), .A2(new_n5658_), .ZN(new_n5659_));
  XOR2_X1    g05466(.A1(new_n5483_), .A2(new_n5659_), .Z(\asquared[55] ));
  OAI21_X1   g05467(.A1(new_n5482_), .A2(new_n5477_), .B(new_n5656_), .ZN(new_n5661_));
  NAND2_X1   g05468(.A1(new_n5661_), .A2(new_n5658_), .ZN(new_n5662_));
  INV_X1     g05469(.I(new_n5642_), .ZN(new_n5663_));
  NAND2_X1   g05470(.A1(new_n5615_), .A2(new_n5663_), .ZN(new_n5664_));
  INV_X1     g05471(.I(new_n5643_), .ZN(new_n5665_));
  NAND2_X1   g05472(.A1(new_n5665_), .A2(new_n5646_), .ZN(new_n5666_));
  NAND2_X1   g05473(.A1(new_n5666_), .A2(new_n5664_), .ZN(new_n5667_));
  XOR2_X1    g05474(.A1(new_n5639_), .A2(new_n5630_), .Z(new_n5668_));
  XOR2_X1    g05475(.A1(new_n5668_), .A2(new_n5582_), .Z(new_n5669_));
  NAND2_X1   g05476(.A1(new_n5562_), .A2(new_n5572_), .ZN(new_n5670_));
  NAND2_X1   g05477(.A1(new_n5573_), .A2(new_n5583_), .ZN(new_n5671_));
  NAND2_X1   g05478(.A1(new_n5671_), .A2(new_n5670_), .ZN(new_n5672_));
  NAND2_X1   g05479(.A1(new_n5531_), .A2(new_n5541_), .ZN(new_n5673_));
  INV_X1     g05480(.I(new_n5542_), .ZN(new_n5674_));
  NAND2_X1   g05481(.A1(new_n5674_), .A2(new_n5551_), .ZN(new_n5675_));
  NAND2_X1   g05482(.A1(new_n5675_), .A2(new_n5673_), .ZN(new_n5676_));
  XOR2_X1    g05483(.A1(new_n5672_), .A2(new_n5676_), .Z(new_n5677_));
  XNOR2_X1   g05484(.A1(new_n5677_), .A2(new_n5669_), .ZN(new_n5678_));
  XOR2_X1    g05485(.A1(new_n5667_), .A2(new_n5678_), .Z(new_n5679_));
  INV_X1     g05486(.I(\a[55] ), .ZN(new_n5680_));
  AOI22_X1   g05487(.A1(\a[51] ), .A2(new_n980_), .B1(new_n533_), .B2(\a[53] ), .ZN(new_n5681_));
  NOR2_X1    g05488(.A1(new_n5135_), .A2(new_n5425_), .ZN(new_n5682_));
  INV_X1     g05489(.I(new_n5682_), .ZN(new_n5683_));
  NOR2_X1    g05490(.A1(new_n5683_), .A2(new_n251_), .ZN(new_n5684_));
  NOR3_X1    g05491(.A1(new_n5684_), .A2(new_n5681_), .A3(new_n5680_), .ZN(new_n5685_));
  NAND2_X1   g05492(.A1(\a[0] ), .A2(\a[55] ), .ZN(new_n5686_));
  NOR2_X1    g05493(.A1(new_n5685_), .A2(new_n5684_), .ZN(new_n5687_));
  INV_X1     g05494(.I(new_n5687_), .ZN(new_n5688_));
  AOI22_X1   g05495(.A1(\a[2] ), .A2(\a[53] ), .B1(\a[4] ), .B2(\a[51] ), .ZN(new_n5689_));
  OAI22_X1   g05496(.A1(new_n5688_), .A2(new_n5689_), .B1(new_n5685_), .B2(new_n5686_), .ZN(new_n5690_));
  NAND2_X1   g05497(.A1(new_n1552_), .A2(new_n2525_), .ZN(new_n5691_));
  NAND2_X1   g05498(.A1(new_n1381_), .A2(new_n2745_), .ZN(new_n5692_));
  AOI22_X1   g05499(.A1(new_n5691_), .A2(new_n5692_), .B1(new_n1452_), .B2(new_n3577_), .ZN(new_n5693_));
  NAND2_X1   g05500(.A1(\a[20] ), .A2(\a[35] ), .ZN(new_n5694_));
  AOI22_X1   g05501(.A1(\a[21] ), .A2(\a[34] ), .B1(\a[22] ), .B2(\a[33] ), .ZN(new_n5695_));
  NAND2_X1   g05502(.A1(new_n1452_), .A2(new_n3577_), .ZN(new_n5696_));
  NAND3_X1   g05503(.A1(new_n5696_), .A2(new_n5691_), .A3(new_n5692_), .ZN(new_n5697_));
  OAI22_X1   g05504(.A1(new_n5693_), .A2(new_n5694_), .B1(new_n5697_), .B2(new_n5695_), .ZN(new_n5698_));
  XOR2_X1    g05505(.A1(new_n5690_), .A2(new_n5698_), .Z(new_n5699_));
  AOI22_X1   g05506(.A1(new_n1442_), .A2(new_n2201_), .B1(new_n1528_), .B2(new_n3210_), .ZN(new_n5700_));
  AOI21_X1   g05507(.A1(new_n1778_), .A2(new_n2437_), .B(new_n5700_), .ZN(new_n5701_));
  NAND2_X1   g05508(.A1(\a[23] ), .A2(\a[32] ), .ZN(new_n5702_));
  AOI22_X1   g05509(.A1(\a[24] ), .A2(\a[31] ), .B1(\a[25] ), .B2(\a[30] ), .ZN(new_n5703_));
  OAI21_X1   g05510(.A1(new_n1779_), .A2(new_n2438_), .B(new_n5700_), .ZN(new_n5704_));
  OAI22_X1   g05511(.A1(new_n5701_), .A2(new_n5702_), .B1(new_n5704_), .B2(new_n5703_), .ZN(new_n5705_));
  XNOR2_X1   g05512(.A1(new_n5699_), .A2(new_n5705_), .ZN(new_n5706_));
  INV_X1     g05513(.I(new_n5706_), .ZN(new_n5707_));
  OAI21_X1   g05514(.A1(new_n5511_), .A2(new_n5316_), .B(new_n5510_), .ZN(new_n5708_));
  INV_X1     g05515(.I(new_n5513_), .ZN(new_n5709_));
  OAI21_X1   g05516(.A1(new_n5709_), .A2(new_n5507_), .B(new_n5708_), .ZN(new_n5710_));
  NOR2_X1    g05517(.A1(new_n536_), .A2(new_n3666_), .ZN(new_n5711_));
  AOI21_X1   g05518(.A1(\a[26] ), .A2(\a[29] ), .B(new_n2103_), .ZN(new_n5712_));
  INV_X1     g05519(.I(new_n5712_), .ZN(new_n5713_));
  NOR3_X1    g05520(.A1(new_n2189_), .A2(new_n1566_), .A3(new_n1814_), .ZN(new_n5714_));
  INV_X1     g05521(.I(new_n5714_), .ZN(new_n5715_));
  NAND3_X1   g05522(.A1(new_n5715_), .A2(new_n5711_), .A3(new_n5713_), .ZN(new_n5716_));
  NAND2_X1   g05523(.A1(new_n5716_), .A2(new_n5715_), .ZN(new_n5717_));
  INV_X1     g05524(.I(new_n5717_), .ZN(new_n5718_));
  AOI22_X1   g05525(.A1(new_n5718_), .A2(new_n5713_), .B1(new_n5711_), .B2(new_n5716_), .ZN(new_n5719_));
  NOR2_X1    g05526(.A1(new_n3861_), .A2(new_n833_), .ZN(new_n5720_));
  NOR3_X1    g05527(.A1(new_n5238_), .A2(new_n597_), .A3(new_n4030_), .ZN(new_n5721_));
  NOR2_X1    g05528(.A1(new_n1264_), .A2(new_n4704_), .ZN(new_n5722_));
  NOR2_X1    g05529(.A1(new_n5721_), .A2(new_n5722_), .ZN(new_n5723_));
  NOR2_X1    g05530(.A1(new_n5723_), .A2(new_n5720_), .ZN(new_n5724_));
  NAND2_X1   g05531(.A1(\a[10] ), .A2(\a[45] ), .ZN(new_n5725_));
  AOI22_X1   g05532(.A1(\a[11] ), .A2(\a[44] ), .B1(\a[13] ), .B2(\a[42] ), .ZN(new_n5726_));
  NOR2_X1    g05533(.A1(new_n5724_), .A2(new_n5720_), .ZN(new_n5727_));
  INV_X1     g05534(.I(new_n5727_), .ZN(new_n5728_));
  OAI22_X1   g05535(.A1(new_n5728_), .A2(new_n5726_), .B1(new_n5724_), .B2(new_n5725_), .ZN(new_n5729_));
  XNOR2_X1   g05536(.A1(new_n5729_), .A2(new_n5719_), .ZN(new_n5730_));
  AOI22_X1   g05537(.A1(\a[7] ), .A2(\a[48] ), .B1(\a[8] ), .B2(\a[47] ), .ZN(new_n5731_));
  NOR2_X1    g05538(.A1(new_n742_), .A2(new_n3116_), .ZN(new_n5732_));
  INV_X1     g05539(.I(new_n5732_), .ZN(new_n5733_));
  NOR2_X1    g05540(.A1(new_n4977_), .A2(new_n415_), .ZN(new_n5734_));
  NOR3_X1    g05541(.A1(new_n5734_), .A2(new_n5731_), .A3(new_n5733_), .ZN(new_n5735_));
  NOR2_X1    g05542(.A1(new_n5735_), .A2(new_n5734_), .ZN(new_n5736_));
  INV_X1     g05543(.I(new_n5736_), .ZN(new_n5737_));
  OAI22_X1   g05544(.A1(new_n5737_), .A2(new_n5731_), .B1(new_n5733_), .B2(new_n5735_), .ZN(new_n5738_));
  XOR2_X1    g05545(.A1(new_n5730_), .A2(new_n5738_), .Z(new_n5739_));
  XOR2_X1    g05546(.A1(new_n5710_), .A2(new_n5739_), .Z(new_n5740_));
  XOR2_X1    g05547(.A1(new_n5740_), .A2(new_n5707_), .Z(new_n5741_));
  XOR2_X1    g05548(.A1(new_n5679_), .A2(new_n5741_), .Z(new_n5742_));
  NOR2_X1    g05549(.A1(new_n5608_), .A2(new_n5611_), .ZN(new_n5743_));
  NAND2_X1   g05550(.A1(new_n5608_), .A2(new_n5611_), .ZN(new_n5744_));
  OAI21_X1   g05551(.A1(new_n5743_), .A2(new_n5647_), .B(new_n5744_), .ZN(new_n5745_));
  NAND2_X1   g05552(.A1(new_n5584_), .A2(new_n5587_), .ZN(new_n5746_));
  NAND2_X1   g05553(.A1(new_n5588_), .A2(new_n5553_), .ZN(new_n5747_));
  NAND2_X1   g05554(.A1(new_n5747_), .A2(new_n5746_), .ZN(new_n5748_));
  NAND2_X1   g05555(.A1(new_n5410_), .A2(new_n5443_), .ZN(new_n5749_));
  NAND2_X1   g05556(.A1(new_n5593_), .A2(new_n5383_), .ZN(new_n5750_));
  NAND2_X1   g05557(.A1(new_n5750_), .A2(new_n5749_), .ZN(new_n5751_));
  INV_X1     g05558(.I(new_n5419_), .ZN(new_n5752_));
  NAND2_X1   g05559(.A1(new_n5491_), .A2(new_n5397_), .ZN(new_n5753_));
  OAI21_X1   g05560(.A1(new_n5752_), .A2(new_n5431_), .B(new_n5753_), .ZN(new_n5754_));
  XOR2_X1    g05561(.A1(new_n5754_), .A2(new_n5751_), .Z(new_n5755_));
  NOR2_X1    g05562(.A1(new_n3341_), .A2(new_n5620_), .ZN(new_n5756_));
  NOR2_X1    g05563(.A1(new_n1718_), .A2(new_n5617_), .ZN(new_n5757_));
  INV_X1     g05564(.I(new_n5757_), .ZN(new_n5758_));
  NOR2_X1    g05565(.A1(new_n5758_), .A2(new_n194_), .ZN(new_n5759_));
  INV_X1     g05566(.I(new_n5759_), .ZN(new_n5760_));
  NOR2_X1    g05567(.A1(new_n194_), .A2(new_n5617_), .ZN(new_n5761_));
  OAI21_X1   g05568(.A1(\a[28] ), .A2(new_n5761_), .B(new_n5760_), .ZN(new_n5762_));
  XOR2_X1    g05569(.A1(new_n5762_), .A2(new_n5756_), .Z(new_n5763_));
  XNOR2_X1   g05570(.A1(new_n5763_), .A2(new_n5560_), .ZN(new_n5764_));
  INV_X1     g05571(.I(new_n5764_), .ZN(new_n5765_));
  XOR2_X1    g05572(.A1(new_n5755_), .A2(new_n5765_), .Z(new_n5766_));
  XOR2_X1    g05573(.A1(new_n5748_), .A2(new_n5766_), .Z(new_n5767_));
  XOR2_X1    g05574(.A1(new_n5530_), .A2(new_n5549_), .Z(new_n5768_));
  XOR2_X1    g05575(.A1(new_n5768_), .A2(new_n5570_), .Z(new_n5769_));
  NAND2_X1   g05576(.A1(new_n5631_), .A2(new_n5640_), .ZN(new_n5770_));
  OAI21_X1   g05577(.A1(new_n5641_), .A2(new_n5622_), .B(new_n5770_), .ZN(new_n5771_));
  NAND2_X1   g05578(.A1(new_n5771_), .A2(new_n5769_), .ZN(new_n5772_));
  INV_X1     g05579(.I(new_n5772_), .ZN(new_n5773_));
  NOR2_X1    g05580(.A1(new_n5771_), .A2(new_n5769_), .ZN(new_n5774_));
  NOR2_X1    g05581(.A1(new_n5773_), .A2(new_n5774_), .ZN(new_n5775_));
  NAND2_X1   g05582(.A1(new_n5616_), .A2(new_n5618_), .ZN(new_n5776_));
  NAND2_X1   g05583(.A1(new_n5619_), .A2(new_n5621_), .ZN(new_n5777_));
  NAND2_X1   g05584(.A1(new_n5777_), .A2(new_n5776_), .ZN(new_n5778_));
  XOR2_X1    g05585(.A1(new_n5778_), .A2(new_n5540_), .Z(new_n5779_));
  AOI22_X1   g05586(.A1(\a[18] ), .A2(\a[37] ), .B1(\a[19] ), .B2(\a[36] ), .ZN(new_n5780_));
  NOR2_X1    g05587(.A1(new_n253_), .A2(new_n4901_), .ZN(new_n5781_));
  INV_X1     g05588(.I(new_n5781_), .ZN(new_n5782_));
  NOR2_X1    g05589(.A1(new_n3038_), .A2(new_n1092_), .ZN(new_n5783_));
  NOR3_X1    g05590(.A1(new_n5783_), .A2(new_n5780_), .A3(new_n5782_), .ZN(new_n5784_));
  NOR2_X1    g05591(.A1(new_n5784_), .A2(new_n5783_), .ZN(new_n5785_));
  INV_X1     g05592(.I(new_n5785_), .ZN(new_n5786_));
  OAI22_X1   g05593(.A1(new_n5786_), .A2(new_n5780_), .B1(new_n5782_), .B2(new_n5784_), .ZN(new_n5787_));
  XNOR2_X1   g05594(.A1(new_n5779_), .A2(new_n5787_), .ZN(new_n5788_));
  XNOR2_X1   g05595(.A1(new_n5775_), .A2(new_n5788_), .ZN(new_n5789_));
  XNOR2_X1   g05596(.A1(new_n5767_), .A2(new_n5789_), .ZN(new_n5790_));
  INV_X1     g05597(.I(new_n5790_), .ZN(new_n5791_));
  XOR2_X1    g05598(.A1(new_n5745_), .A2(new_n5791_), .Z(new_n5792_));
  XNOR2_X1   g05599(.A1(new_n5792_), .A2(new_n5742_), .ZN(new_n5793_));
  INV_X1     g05600(.I(new_n5520_), .ZN(new_n5794_));
  OAI21_X1   g05601(.A1(new_n5794_), .A2(new_n5605_), .B(new_n5519_), .ZN(new_n5795_));
  NAND2_X1   g05602(.A1(new_n5592_), .A2(new_n5603_), .ZN(new_n5796_));
  NAND2_X1   g05603(.A1(new_n5604_), .A2(new_n5589_), .ZN(new_n5797_));
  NAND2_X1   g05604(.A1(new_n5797_), .A2(new_n5796_), .ZN(new_n5798_));
  NAND2_X1   g05605(.A1(new_n5505_), .A2(new_n5514_), .ZN(new_n5799_));
  NAND2_X1   g05606(.A1(new_n5515_), .A2(new_n5502_), .ZN(new_n5800_));
  NAND2_X1   g05607(.A1(new_n5800_), .A2(new_n5799_), .ZN(new_n5801_));
  NOR2_X1    g05608(.A1(new_n5500_), .A2(new_n5498_), .ZN(new_n5802_));
  NAND2_X1   g05609(.A1(new_n5598_), .A2(new_n5601_), .ZN(new_n5803_));
  NAND2_X1   g05610(.A1(new_n5602_), .A2(new_n5594_), .ZN(new_n5804_));
  NAND2_X1   g05611(.A1(new_n5804_), .A2(new_n5803_), .ZN(new_n5805_));
  NAND2_X1   g05612(.A1(new_n5495_), .A2(new_n5390_), .ZN(new_n5806_));
  OAI21_X1   g05613(.A1(new_n5450_), .A2(new_n5460_), .B(new_n5806_), .ZN(new_n5807_));
  AOI22_X1   g05614(.A1(\a[6] ), .A2(\a[49] ), .B1(\a[17] ), .B2(\a[38] ), .ZN(new_n5808_));
  INV_X1     g05615(.I(new_n5808_), .ZN(new_n5809_));
  NOR3_X1    g05616(.A1(new_n3798_), .A2(new_n1023_), .A3(new_n4702_), .ZN(new_n5810_));
  NOR2_X1    g05617(.A1(new_n225_), .A2(new_n5175_), .ZN(new_n5811_));
  AOI21_X1   g05618(.A1(new_n5809_), .A2(new_n5811_), .B(new_n5810_), .ZN(new_n5812_));
  INV_X1     g05619(.I(new_n5812_), .ZN(new_n5813_));
  OAI21_X1   g05620(.A1(new_n5810_), .A2(new_n5808_), .B(new_n5811_), .ZN(new_n5814_));
  OAI21_X1   g05621(.A1(new_n5813_), .A2(new_n5808_), .B(new_n5814_), .ZN(new_n5815_));
  NOR2_X1    g05622(.A1(new_n759_), .A2(new_n3327_), .ZN(new_n5816_));
  NOR2_X1    g05623(.A1(new_n403_), .A2(new_n4178_), .ZN(new_n5817_));
  NAND2_X1   g05624(.A1(new_n5816_), .A2(new_n5817_), .ZN(new_n5818_));
  INV_X1     g05625(.I(new_n5818_), .ZN(new_n5819_));
  INV_X1     g05626(.I(new_n1370_), .ZN(new_n5820_));
  NOR3_X1    g05627(.A1(new_n5820_), .A2(new_n3221_), .A3(new_n4178_), .ZN(new_n5821_));
  NOR2_X1    g05628(.A1(new_n1173_), .A2(new_n5377_), .ZN(new_n5822_));
  NOR2_X1    g05629(.A1(new_n5821_), .A2(new_n5822_), .ZN(new_n5823_));
  NOR2_X1    g05630(.A1(new_n5823_), .A2(new_n5819_), .ZN(new_n5824_));
  NAND2_X1   g05631(.A1(\a[15] ), .A2(\a[40] ), .ZN(new_n5825_));
  NOR2_X1    g05632(.A1(new_n5824_), .A2(new_n5819_), .ZN(new_n5826_));
  OAI21_X1   g05633(.A1(new_n5816_), .A2(new_n5817_), .B(new_n5826_), .ZN(new_n5827_));
  OAI21_X1   g05634(.A1(new_n5824_), .A2(new_n5825_), .B(new_n5827_), .ZN(new_n5828_));
  XNOR2_X1   g05635(.A1(new_n5828_), .A2(new_n5815_), .ZN(new_n5829_));
  XNOR2_X1   g05636(.A1(new_n5829_), .A2(new_n5807_), .ZN(new_n5830_));
  XNOR2_X1   g05637(.A1(new_n5805_), .A2(new_n5830_), .ZN(new_n5831_));
  NAND2_X1   g05638(.A1(new_n5831_), .A2(new_n5802_), .ZN(new_n5832_));
  OR2_X2     g05639(.A1(new_n5831_), .A2(new_n5802_), .Z(new_n5833_));
  NAND2_X1   g05640(.A1(new_n5833_), .A2(new_n5832_), .ZN(new_n5834_));
  XNOR2_X1   g05641(.A1(new_n5834_), .A2(new_n5801_), .ZN(new_n5835_));
  XOR2_X1    g05642(.A1(new_n5835_), .A2(new_n5798_), .Z(new_n5836_));
  XOR2_X1    g05643(.A1(new_n5795_), .A2(new_n5836_), .Z(new_n5837_));
  NAND2_X1   g05644(.A1(new_n5837_), .A2(new_n5793_), .ZN(new_n5838_));
  INV_X1     g05645(.I(new_n5838_), .ZN(new_n5839_));
  NOR2_X1    g05646(.A1(new_n5837_), .A2(new_n5793_), .ZN(new_n5840_));
  NOR2_X1    g05647(.A1(new_n5839_), .A2(new_n5840_), .ZN(new_n5841_));
  INV_X1     g05648(.I(new_n5841_), .ZN(new_n5842_));
  INV_X1     g05649(.I(new_n5648_), .ZN(new_n5843_));
  NAND2_X1   g05650(.A1(new_n5651_), .A2(new_n5843_), .ZN(new_n5844_));
  OAI21_X1   g05651(.A1(new_n5652_), .A2(new_n5606_), .B(new_n5844_), .ZN(new_n5845_));
  INV_X1     g05652(.I(new_n5845_), .ZN(new_n5846_));
  NOR2_X1    g05653(.A1(new_n5842_), .A2(new_n5846_), .ZN(new_n5847_));
  NOR2_X1    g05654(.A1(new_n5841_), .A2(new_n5845_), .ZN(new_n5848_));
  NOR2_X1    g05655(.A1(new_n5847_), .A2(new_n5848_), .ZN(new_n5849_));
  XOR2_X1    g05656(.A1(new_n5662_), .A2(new_n5849_), .Z(\asquared[56] ));
  AOI21_X1   g05657(.A1(new_n5661_), .A2(new_n5658_), .B(new_n5848_), .ZN(new_n5851_));
  NOR2_X1    g05658(.A1(new_n5851_), .A2(new_n5847_), .ZN(new_n5852_));
  NAND2_X1   g05659(.A1(new_n5795_), .A2(new_n5836_), .ZN(new_n5853_));
  NAND2_X1   g05660(.A1(new_n5838_), .A2(new_n5853_), .ZN(new_n5854_));
  INV_X1     g05661(.I(new_n5854_), .ZN(new_n5855_));
  INV_X1     g05662(.I(\a[56] ), .ZN(new_n5856_));
  NOR2_X1    g05663(.A1(new_n5617_), .A2(new_n5856_), .ZN(new_n5857_));
  AOI22_X1   g05664(.A1(\a[0] ), .A2(\a[56] ), .B1(\a[2] ), .B2(\a[54] ), .ZN(new_n5858_));
  AOI21_X1   g05665(.A1(new_n5857_), .A2(new_n533_), .B(new_n5858_), .ZN(new_n5859_));
  XOR2_X1    g05666(.A1(new_n5759_), .A2(new_n5859_), .Z(new_n5860_));
  XNOR2_X1   g05667(.A1(new_n5860_), .A2(new_n5736_), .ZN(new_n5861_));
  NOR2_X1    g05668(.A1(new_n5175_), .A2(new_n5425_), .ZN(new_n5862_));
  NAND2_X1   g05669(.A1(new_n5862_), .A2(new_n761_), .ZN(new_n5863_));
  NAND3_X1   g05670(.A1(new_n1191_), .A2(\a[37] ), .A3(\a[53] ), .ZN(new_n5864_));
  NOR4_X1    g05671(.A1(new_n290_), .A2(new_n979_), .A3(new_n2752_), .A4(new_n5175_), .ZN(new_n5865_));
  AOI21_X1   g05672(.A1(new_n5864_), .A2(new_n5863_), .B(new_n5865_), .ZN(new_n5866_));
  NAND2_X1   g05673(.A1(\a[3] ), .A2(\a[53] ), .ZN(new_n5867_));
  AOI22_X1   g05674(.A1(\a[4] ), .A2(\a[52] ), .B1(\a[19] ), .B2(\a[37] ), .ZN(new_n5868_));
  OR2_X2     g05675(.A1(new_n5866_), .A2(new_n5865_), .Z(new_n5869_));
  OAI22_X1   g05676(.A1(new_n5869_), .A2(new_n5868_), .B1(new_n5866_), .B2(new_n5867_), .ZN(new_n5870_));
  XOR2_X1    g05677(.A1(new_n5861_), .A2(new_n5870_), .Z(new_n5871_));
  NAND2_X1   g05678(.A1(new_n2176_), .A2(new_n2437_), .ZN(new_n5872_));
  OAI22_X1   g05679(.A1(new_n1779_), .A2(new_n3833_), .B1(new_n2081_), .B2(new_n2202_), .ZN(new_n5873_));
  NAND2_X1   g05680(.A1(new_n5873_), .A2(new_n5872_), .ZN(new_n5874_));
  NAND3_X1   g05681(.A1(new_n5874_), .A2(\a[24] ), .A3(\a[32] ), .ZN(new_n5875_));
  AOI22_X1   g05682(.A1(\a[25] ), .A2(\a[31] ), .B1(\a[26] ), .B2(\a[30] ), .ZN(new_n5876_));
  NAND2_X1   g05683(.A1(new_n5874_), .A2(new_n5872_), .ZN(new_n5877_));
  OAI21_X1   g05684(.A1(new_n5876_), .A2(new_n5877_), .B(new_n5875_), .ZN(new_n5878_));
  NAND2_X1   g05685(.A1(new_n1767_), .A2(new_n3577_), .ZN(new_n5879_));
  NOR2_X1    g05686(.A1(new_n2647_), .A2(new_n5564_), .ZN(new_n5880_));
  NOR4_X1    g05687(.A1(new_n1043_), .A2(new_n1299_), .A3(new_n2274_), .A4(new_n2626_), .ZN(new_n5881_));
  OAI21_X1   g05688(.A1(new_n5880_), .A2(new_n5881_), .B(new_n5879_), .ZN(new_n5882_));
  NAND2_X1   g05689(.A1(new_n5882_), .A2(new_n5879_), .ZN(new_n5883_));
  AOI22_X1   g05690(.A1(\a[22] ), .A2(\a[34] ), .B1(\a[23] ), .B2(\a[33] ), .ZN(new_n5884_));
  NAND3_X1   g05691(.A1(new_n5882_), .A2(\a[20] ), .A3(\a[36] ), .ZN(new_n5885_));
  OAI21_X1   g05692(.A1(new_n5883_), .A2(new_n5884_), .B(new_n5885_), .ZN(new_n5886_));
  XOR2_X1    g05693(.A1(new_n5878_), .A2(new_n5886_), .Z(new_n5887_));
  NOR2_X1    g05694(.A1(new_n759_), .A2(new_n4178_), .ZN(new_n5888_));
  INV_X1     g05695(.I(new_n5888_), .ZN(new_n5889_));
  NAND2_X1   g05696(.A1(\a[14] ), .A2(\a[47] ), .ZN(new_n5890_));
  OAI22_X1   g05697(.A1(new_n539_), .A2(new_n4721_), .B1(new_n5059_), .B2(new_n5890_), .ZN(new_n5891_));
  OAI21_X1   g05698(.A1(new_n5238_), .A2(new_n5889_), .B(new_n5891_), .ZN(new_n5892_));
  NAND3_X1   g05699(.A1(new_n5892_), .A2(\a[9] ), .A3(\a[47] ), .ZN(new_n5893_));
  NOR2_X1    g05700(.A1(new_n5238_), .A2(new_n5889_), .ZN(new_n5894_));
  NOR2_X1    g05701(.A1(new_n5891_), .A2(new_n5894_), .ZN(new_n5895_));
  INV_X1     g05702(.I(new_n5895_), .ZN(new_n5896_));
  AOI22_X1   g05703(.A1(\a[10] ), .A2(\a[46] ), .B1(\a[14] ), .B2(\a[42] ), .ZN(new_n5897_));
  OAI21_X1   g05704(.A1(new_n5896_), .A2(new_n5897_), .B(new_n5893_), .ZN(new_n5898_));
  XOR2_X1    g05705(.A1(new_n5887_), .A2(new_n5898_), .Z(new_n5899_));
  NOR2_X1    g05706(.A1(new_n1023_), .A2(new_n4901_), .ZN(new_n5900_));
  NAND3_X1   g05707(.A1(new_n5900_), .A2(\a[6] ), .A3(\a[39] ), .ZN(new_n5901_));
  OAI21_X1   g05708(.A1(new_n374_), .A2(new_n5155_), .B(new_n5901_), .ZN(new_n5902_));
  NAND4_X1   g05709(.A1(\a[7] ), .A2(\a[17] ), .A3(\a[39] ), .A4(\a[49] ), .ZN(new_n5903_));
  NAND2_X1   g05710(.A1(new_n5902_), .A2(new_n5903_), .ZN(new_n5904_));
  NAND3_X1   g05711(.A1(new_n5904_), .A2(\a[6] ), .A3(\a[50] ), .ZN(new_n5905_));
  AOI22_X1   g05712(.A1(\a[7] ), .A2(\a[49] ), .B1(\a[17] ), .B2(\a[39] ), .ZN(new_n5906_));
  NAND2_X1   g05713(.A1(new_n5904_), .A2(new_n5903_), .ZN(new_n5907_));
  OAI21_X1   g05714(.A1(new_n5906_), .A2(new_n5907_), .B(new_n5905_), .ZN(new_n5908_));
  NAND2_X1   g05715(.A1(new_n763_), .A2(new_n4342_), .ZN(new_n5909_));
  OAI22_X1   g05716(.A1(new_n619_), .A2(new_n4704_), .B1(new_n4034_), .B2(new_n833_), .ZN(new_n5910_));
  NAND2_X1   g05717(.A1(new_n5910_), .A2(new_n5909_), .ZN(new_n5911_));
  NAND3_X1   g05718(.A1(new_n5911_), .A2(\a[11] ), .A3(\a[45] ), .ZN(new_n5912_));
  AOI21_X1   g05719(.A1(\a[12] ), .A2(\a[44] ), .B(new_n5049_), .ZN(new_n5913_));
  NAND2_X1   g05720(.A1(new_n5911_), .A2(new_n5909_), .ZN(new_n5914_));
  OAI21_X1   g05721(.A1(new_n5913_), .A2(new_n5914_), .B(new_n5912_), .ZN(new_n5915_));
  XOR2_X1    g05722(.A1(new_n5908_), .A2(new_n5915_), .Z(new_n5916_));
  NOR2_X1    g05723(.A1(new_n717_), .A2(new_n4596_), .ZN(new_n5917_));
  NOR2_X1    g05724(.A1(new_n3221_), .A2(new_n4596_), .ZN(new_n5918_));
  NAND3_X1   g05725(.A1(new_n5918_), .A2(\a[8] ), .A3(\a[16] ), .ZN(new_n5919_));
  NAND2_X1   g05726(.A1(new_n4534_), .A2(new_n1288_), .ZN(new_n5920_));
  AOI22_X1   g05727(.A1(new_n5919_), .A2(new_n5920_), .B1(new_n4664_), .B2(new_n5917_), .ZN(new_n5921_));
  NAND2_X1   g05728(.A1(new_n4664_), .A2(new_n5917_), .ZN(new_n5922_));
  NAND3_X1   g05729(.A1(new_n5922_), .A2(new_n5919_), .A3(new_n5920_), .ZN(new_n5923_));
  AOI22_X1   g05730(.A1(\a[8] ), .A2(\a[48] ), .B1(\a[15] ), .B2(\a[41] ), .ZN(new_n5924_));
  OAI22_X1   g05731(.A1(new_n5921_), .A2(new_n3549_), .B1(new_n5923_), .B2(new_n5924_), .ZN(new_n5925_));
  XOR2_X1    g05732(.A1(new_n5916_), .A2(new_n5925_), .Z(new_n5926_));
  XOR2_X1    g05733(.A1(new_n5926_), .A2(new_n5899_), .Z(new_n5927_));
  XOR2_X1    g05734(.A1(new_n5927_), .A2(new_n5871_), .Z(new_n5928_));
  NAND2_X1   g05735(.A1(new_n5805_), .A2(new_n5830_), .ZN(new_n5929_));
  NAND2_X1   g05736(.A1(new_n5833_), .A2(new_n5929_), .ZN(new_n5930_));
  XOR2_X1    g05737(.A1(new_n5704_), .A2(new_n5697_), .Z(new_n5931_));
  XOR2_X1    g05738(.A1(new_n5931_), .A2(new_n5813_), .Z(new_n5932_));
  INV_X1     g05739(.I(new_n5719_), .ZN(new_n5933_));
  NAND2_X1   g05740(.A1(new_n5933_), .A2(new_n5729_), .ZN(new_n5934_));
  NAND2_X1   g05741(.A1(new_n5730_), .A2(new_n5738_), .ZN(new_n5935_));
  NAND2_X1   g05742(.A1(new_n5935_), .A2(new_n5934_), .ZN(new_n5936_));
  NAND2_X1   g05743(.A1(\a[1] ), .A2(\a[55] ), .ZN(new_n5937_));
  NOR2_X1    g05744(.A1(new_n1816_), .A2(new_n5937_), .ZN(new_n5938_));
  INV_X1     g05745(.I(new_n5938_), .ZN(new_n5939_));
  NAND2_X1   g05746(.A1(new_n1816_), .A2(new_n5937_), .ZN(new_n5940_));
  AND2_X2    g05747(.A1(new_n5939_), .A2(new_n5940_), .Z(new_n5941_));
  NOR2_X1    g05748(.A1(new_n5718_), .A2(new_n5941_), .ZN(new_n5942_));
  INV_X1     g05749(.I(new_n5941_), .ZN(new_n5943_));
  NOR2_X1    g05750(.A1(new_n5943_), .A2(new_n5717_), .ZN(new_n5944_));
  OAI21_X1   g05751(.A1(new_n5942_), .A2(new_n5944_), .B(new_n5728_), .ZN(new_n5945_));
  INV_X1     g05752(.I(new_n5945_), .ZN(new_n5946_));
  NOR3_X1    g05753(.A1(new_n5942_), .A2(new_n5728_), .A3(new_n5944_), .ZN(new_n5947_));
  NOR2_X1    g05754(.A1(new_n5946_), .A2(new_n5947_), .ZN(new_n5948_));
  XOR2_X1    g05755(.A1(new_n5936_), .A2(new_n5948_), .Z(new_n5949_));
  XOR2_X1    g05756(.A1(new_n5949_), .A2(new_n5932_), .Z(new_n5950_));
  XOR2_X1    g05757(.A1(new_n5930_), .A2(new_n5950_), .Z(new_n5951_));
  XNOR2_X1   g05758(.A1(new_n5951_), .A2(new_n5928_), .ZN(new_n5952_));
  AOI21_X1   g05759(.A1(new_n5799_), .A2(new_n5800_), .B(new_n5834_), .ZN(new_n5953_));
  AOI21_X1   g05760(.A1(new_n5835_), .A2(new_n5798_), .B(new_n5953_), .ZN(new_n5954_));
  NAND2_X1   g05761(.A1(new_n5754_), .A2(new_n5751_), .ZN(new_n5955_));
  NAND2_X1   g05762(.A1(new_n5755_), .A2(new_n5765_), .ZN(new_n5956_));
  NAND2_X1   g05763(.A1(new_n5956_), .A2(new_n5955_), .ZN(new_n5957_));
  NOR2_X1    g05764(.A1(new_n5688_), .A2(new_n5786_), .ZN(new_n5958_));
  NOR2_X1    g05765(.A1(new_n5687_), .A2(new_n5785_), .ZN(new_n5959_));
  NOR2_X1    g05766(.A1(new_n5958_), .A2(new_n5959_), .ZN(new_n5960_));
  XNOR2_X1   g05767(.A1(new_n5960_), .A2(new_n5826_), .ZN(new_n5961_));
  NAND2_X1   g05768(.A1(new_n5828_), .A2(new_n5815_), .ZN(new_n5962_));
  INV_X1     g05769(.I(new_n5829_), .ZN(new_n5963_));
  NAND2_X1   g05770(.A1(new_n5963_), .A2(new_n5807_), .ZN(new_n5964_));
  NAND2_X1   g05771(.A1(new_n5964_), .A2(new_n5962_), .ZN(new_n5965_));
  XOR2_X1    g05772(.A1(new_n5965_), .A2(new_n5961_), .Z(new_n5966_));
  XOR2_X1    g05773(.A1(new_n5966_), .A2(new_n5957_), .Z(new_n5967_));
  INV_X1     g05774(.I(new_n5967_), .ZN(new_n5968_));
  NAND2_X1   g05775(.A1(new_n5690_), .A2(new_n5698_), .ZN(new_n5969_));
  NAND2_X1   g05776(.A1(new_n5699_), .A2(new_n5705_), .ZN(new_n5970_));
  NAND2_X1   g05777(.A1(new_n5970_), .A2(new_n5969_), .ZN(new_n5971_));
  NAND2_X1   g05778(.A1(new_n5639_), .A2(new_n5630_), .ZN(new_n5972_));
  NAND2_X1   g05779(.A1(new_n5668_), .A2(new_n5582_), .ZN(new_n5973_));
  NAND2_X1   g05780(.A1(new_n5973_), .A2(new_n5972_), .ZN(new_n5974_));
  NAND2_X1   g05781(.A1(new_n5778_), .A2(new_n5540_), .ZN(new_n5975_));
  NAND2_X1   g05782(.A1(new_n5779_), .A2(new_n5787_), .ZN(new_n5976_));
  NAND2_X1   g05783(.A1(new_n5976_), .A2(new_n5975_), .ZN(new_n5977_));
  NOR2_X1    g05784(.A1(new_n5977_), .A2(new_n5974_), .ZN(new_n5978_));
  NAND2_X1   g05785(.A1(new_n5977_), .A2(new_n5974_), .ZN(new_n5979_));
  INV_X1     g05786(.I(new_n5979_), .ZN(new_n5980_));
  NOR2_X1    g05787(.A1(new_n5980_), .A2(new_n5978_), .ZN(new_n5981_));
  NOR2_X1    g05788(.A1(new_n5981_), .A2(new_n5971_), .ZN(new_n5982_));
  NAND2_X1   g05789(.A1(new_n5981_), .A2(new_n5971_), .ZN(new_n5983_));
  INV_X1     g05790(.I(new_n5983_), .ZN(new_n5984_));
  NOR2_X1    g05791(.A1(new_n5984_), .A2(new_n5982_), .ZN(new_n5985_));
  NAND2_X1   g05792(.A1(new_n5710_), .A2(new_n5739_), .ZN(new_n5986_));
  NAND2_X1   g05793(.A1(new_n5740_), .A2(new_n5707_), .ZN(new_n5987_));
  NAND2_X1   g05794(.A1(new_n5987_), .A2(new_n5986_), .ZN(new_n5988_));
  NAND2_X1   g05795(.A1(new_n5988_), .A2(new_n5985_), .ZN(new_n5989_));
  NAND2_X1   g05796(.A1(new_n5989_), .A2(new_n5985_), .ZN(new_n5990_));
  NAND2_X1   g05797(.A1(new_n5989_), .A2(new_n5988_), .ZN(new_n5991_));
  AOI21_X1   g05798(.A1(new_n5990_), .A2(new_n5991_), .B(new_n5968_), .ZN(new_n5992_));
  INV_X1     g05799(.I(new_n5992_), .ZN(new_n5993_));
  NAND3_X1   g05800(.A1(new_n5990_), .A2(new_n5991_), .A3(new_n5968_), .ZN(new_n5994_));
  NAND2_X1   g05801(.A1(new_n5993_), .A2(new_n5994_), .ZN(new_n5995_));
  XNOR2_X1   g05802(.A1(new_n5954_), .A2(new_n5995_), .ZN(new_n5996_));
  XNOR2_X1   g05803(.A1(new_n5996_), .A2(new_n5952_), .ZN(new_n5997_));
  NAND2_X1   g05804(.A1(new_n5745_), .A2(new_n5791_), .ZN(new_n5998_));
  INV_X1     g05805(.I(new_n5792_), .ZN(new_n5999_));
  OAI21_X1   g05806(.A1(new_n5999_), .A2(new_n5742_), .B(new_n5998_), .ZN(new_n6000_));
  AOI21_X1   g05807(.A1(new_n5666_), .A2(new_n5664_), .B(new_n5678_), .ZN(new_n6001_));
  INV_X1     g05808(.I(new_n5741_), .ZN(new_n6002_));
  NOR2_X1    g05809(.A1(new_n5679_), .A2(new_n6002_), .ZN(new_n6003_));
  OAI21_X1   g05810(.A1(new_n5788_), .A2(new_n5774_), .B(new_n5772_), .ZN(new_n6004_));
  NAND2_X1   g05811(.A1(new_n5672_), .A2(new_n5676_), .ZN(new_n6005_));
  NAND2_X1   g05812(.A1(new_n5677_), .A2(new_n5669_), .ZN(new_n6006_));
  NAND2_X1   g05813(.A1(new_n6006_), .A2(new_n6005_), .ZN(new_n6007_));
  NAND2_X1   g05814(.A1(new_n5530_), .A2(new_n5549_), .ZN(new_n6008_));
  NAND2_X1   g05815(.A1(new_n5768_), .A2(new_n5570_), .ZN(new_n6009_));
  NAND2_X1   g05816(.A1(new_n6009_), .A2(new_n6008_), .ZN(new_n6010_));
  INV_X1     g05817(.I(new_n5762_), .ZN(new_n6011_));
  NOR2_X1    g05818(.A1(new_n5763_), .A2(new_n5560_), .ZN(new_n6012_));
  AOI21_X1   g05819(.A1(new_n5756_), .A2(new_n6011_), .B(new_n6012_), .ZN(new_n6013_));
  AOI22_X1   g05820(.A1(\a[5] ), .A2(\a[51] ), .B1(\a[18] ), .B2(\a[38] ), .ZN(new_n6014_));
  INV_X1     g05821(.I(new_n6014_), .ZN(new_n6015_));
  NOR2_X1    g05822(.A1(new_n1220_), .A2(new_n2524_), .ZN(new_n6016_));
  NOR4_X1    g05823(.A1(new_n253_), .A2(new_n884_), .A3(new_n2914_), .A4(new_n5135_), .ZN(new_n6017_));
  INV_X1     g05824(.I(new_n6017_), .ZN(new_n6018_));
  NOR3_X1    g05825(.A1(new_n6014_), .A2(new_n1220_), .A3(new_n2524_), .ZN(new_n6019_));
  NAND2_X1   g05826(.A1(new_n6018_), .A2(new_n6019_), .ZN(new_n6020_));
  NOR2_X1    g05827(.A1(new_n6019_), .A2(new_n6017_), .ZN(new_n6021_));
  AOI22_X1   g05828(.A1(new_n6020_), .A2(new_n6016_), .B1(new_n6021_), .B2(new_n6015_), .ZN(new_n6022_));
  XNOR2_X1   g05829(.A1(new_n6013_), .A2(new_n6022_), .ZN(new_n6023_));
  XNOR2_X1   g05830(.A1(new_n6023_), .A2(new_n6010_), .ZN(new_n6024_));
  XOR2_X1    g05831(.A1(new_n6007_), .A2(new_n6024_), .Z(new_n6025_));
  XOR2_X1    g05832(.A1(new_n6025_), .A2(new_n6004_), .Z(new_n6026_));
  NAND2_X1   g05833(.A1(new_n5748_), .A2(new_n5766_), .ZN(new_n6027_));
  NAND2_X1   g05834(.A1(new_n5767_), .A2(new_n5789_), .ZN(new_n6028_));
  NAND2_X1   g05835(.A1(new_n6028_), .A2(new_n6027_), .ZN(new_n6029_));
  XOR2_X1    g05836(.A1(new_n6029_), .A2(new_n6026_), .Z(new_n6030_));
  OR3_X2     g05837(.A1(new_n6003_), .A2(new_n6001_), .A3(new_n6030_), .Z(new_n6031_));
  OAI21_X1   g05838(.A1(new_n6003_), .A2(new_n6001_), .B(new_n6030_), .ZN(new_n6032_));
  AND2_X2    g05839(.A1(new_n6031_), .A2(new_n6032_), .Z(new_n6033_));
  INV_X1     g05840(.I(new_n6033_), .ZN(new_n6034_));
  NAND2_X1   g05841(.A1(new_n6000_), .A2(new_n6034_), .ZN(new_n6035_));
  NOR2_X1    g05842(.A1(new_n6000_), .A2(new_n6034_), .ZN(new_n6036_));
  INV_X1     g05843(.I(new_n6036_), .ZN(new_n6037_));
  AOI21_X1   g05844(.A1(new_n6037_), .A2(new_n6035_), .B(new_n5997_), .ZN(new_n6038_));
  INV_X1     g05845(.I(new_n6038_), .ZN(new_n6039_));
  NAND3_X1   g05846(.A1(new_n6037_), .A2(new_n5997_), .A3(new_n6035_), .ZN(new_n6040_));
  NAND2_X1   g05847(.A1(new_n6039_), .A2(new_n6040_), .ZN(new_n6041_));
  NOR2_X1    g05848(.A1(new_n5855_), .A2(new_n6041_), .ZN(new_n6042_));
  INV_X1     g05849(.I(new_n6042_), .ZN(new_n6043_));
  NAND2_X1   g05850(.A1(new_n5855_), .A2(new_n6041_), .ZN(new_n6044_));
  NAND2_X1   g05851(.A1(new_n6043_), .A2(new_n6044_), .ZN(new_n6045_));
  XOR2_X1    g05852(.A1(new_n5852_), .A2(new_n6045_), .Z(\asquared[57] ));
  OAI21_X1   g05853(.A1(new_n5851_), .A2(new_n5847_), .B(new_n6044_), .ZN(new_n6047_));
  NAND2_X1   g05854(.A1(new_n6047_), .A2(new_n6043_), .ZN(new_n6048_));
  NAND2_X1   g05855(.A1(new_n6000_), .A2(new_n6033_), .ZN(new_n6049_));
  NAND2_X1   g05856(.A1(new_n6039_), .A2(new_n6049_), .ZN(new_n6050_));
  NAND2_X1   g05857(.A1(new_n6029_), .A2(new_n6026_), .ZN(new_n6051_));
  NAND2_X1   g05858(.A1(new_n6032_), .A2(new_n6051_), .ZN(new_n6052_));
  NAND2_X1   g05859(.A1(new_n5908_), .A2(new_n5915_), .ZN(new_n6053_));
  NAND2_X1   g05860(.A1(new_n5916_), .A2(new_n5925_), .ZN(new_n6054_));
  NAND2_X1   g05861(.A1(new_n6054_), .A2(new_n6053_), .ZN(new_n6055_));
  XOR2_X1    g05862(.A1(new_n5877_), .A2(new_n5923_), .Z(new_n6056_));
  XOR2_X1    g05863(.A1(new_n6056_), .A2(new_n5907_), .Z(new_n6057_));
  INV_X1     g05864(.I(new_n5857_), .ZN(new_n6058_));
  OAI22_X1   g05865(.A1(new_n5760_), .A2(new_n5858_), .B1(new_n412_), .B2(new_n6058_), .ZN(new_n6059_));
  XOR2_X1    g05866(.A1(new_n5869_), .A2(new_n5883_), .Z(new_n6060_));
  XOR2_X1    g05867(.A1(new_n6060_), .A2(new_n6059_), .Z(new_n6061_));
  NAND2_X1   g05868(.A1(new_n6057_), .A2(new_n6061_), .ZN(new_n6062_));
  INV_X1     g05869(.I(new_n6062_), .ZN(new_n6063_));
  NOR2_X1    g05870(.A1(new_n6057_), .A2(new_n6061_), .ZN(new_n6064_));
  NOR2_X1    g05871(.A1(new_n6063_), .A2(new_n6064_), .ZN(new_n6065_));
  NOR2_X1    g05872(.A1(new_n6065_), .A2(new_n6055_), .ZN(new_n6066_));
  NAND2_X1   g05873(.A1(new_n6065_), .A2(new_n6055_), .ZN(new_n6067_));
  INV_X1     g05874(.I(new_n6067_), .ZN(new_n6068_));
  NOR2_X1    g05875(.A1(new_n6068_), .A2(new_n6066_), .ZN(new_n6069_));
  NAND2_X1   g05876(.A1(new_n5878_), .A2(new_n5886_), .ZN(new_n6070_));
  NAND2_X1   g05877(.A1(new_n5887_), .A2(new_n5898_), .ZN(new_n6071_));
  NAND2_X1   g05878(.A1(new_n6071_), .A2(new_n6070_), .ZN(new_n6072_));
  AOI21_X1   g05879(.A1(new_n5717_), .A2(new_n5941_), .B(new_n5946_), .ZN(new_n6073_));
  NAND2_X1   g05880(.A1(new_n5737_), .A2(new_n5860_), .ZN(new_n6074_));
  NAND2_X1   g05881(.A1(new_n5861_), .A2(new_n5870_), .ZN(new_n6075_));
  NAND2_X1   g05882(.A1(new_n6075_), .A2(new_n6074_), .ZN(new_n6076_));
  INV_X1     g05883(.I(new_n6076_), .ZN(new_n6077_));
  XOR2_X1    g05884(.A1(new_n6073_), .A2(new_n6077_), .Z(new_n6078_));
  NOR2_X1    g05885(.A1(new_n6078_), .A2(new_n6072_), .ZN(new_n6079_));
  NAND2_X1   g05886(.A1(new_n6078_), .A2(new_n6072_), .ZN(new_n6080_));
  INV_X1     g05887(.I(new_n6080_), .ZN(new_n6081_));
  NOR2_X1    g05888(.A1(new_n6081_), .A2(new_n6079_), .ZN(new_n6082_));
  NAND2_X1   g05889(.A1(new_n5927_), .A2(new_n5871_), .ZN(new_n6083_));
  NAND2_X1   g05890(.A1(new_n5926_), .A2(new_n5899_), .ZN(new_n6084_));
  NAND2_X1   g05891(.A1(new_n6083_), .A2(new_n6084_), .ZN(new_n6085_));
  XOR2_X1    g05892(.A1(new_n6085_), .A2(new_n6082_), .Z(new_n6086_));
  XOR2_X1    g05893(.A1(new_n6086_), .A2(new_n6069_), .Z(new_n6087_));
  XOR2_X1    g05894(.A1(new_n6052_), .A2(new_n6087_), .Z(new_n6088_));
  NOR2_X1    g05895(.A1(new_n5984_), .A2(new_n5980_), .ZN(new_n6089_));
  NAND2_X1   g05896(.A1(new_n2679_), .A2(new_n2555_), .ZN(new_n6090_));
  INV_X1     g05897(.I(new_n6090_), .ZN(new_n6091_));
  NOR2_X1    g05898(.A1(new_n2189_), .A2(new_n2255_), .ZN(new_n6092_));
  INV_X1     g05899(.I(new_n6092_), .ZN(new_n6093_));
  NOR2_X1    g05900(.A1(new_n536_), .A2(new_n4030_), .ZN(new_n6094_));
  INV_X1     g05901(.I(new_n6094_), .ZN(new_n6095_));
  OAI21_X1   g05902(.A1(new_n6091_), .A2(new_n6095_), .B(new_n6093_), .ZN(new_n6096_));
  NOR2_X1    g05903(.A1(new_n6096_), .A2(new_n6091_), .ZN(new_n6097_));
  AOI21_X1   g05904(.A1(new_n6093_), .A2(new_n6090_), .B(new_n6095_), .ZN(new_n6098_));
  NOR2_X1    g05905(.A1(new_n6097_), .A2(new_n6098_), .ZN(new_n6099_));
  NOR2_X1    g05906(.A1(new_n3859_), .A2(new_n4178_), .ZN(new_n6100_));
  INV_X1     g05907(.I(new_n6100_), .ZN(new_n6101_));
  NOR2_X1    g05908(.A1(new_n6101_), .A2(new_n833_), .ZN(new_n6102_));
  NOR3_X1    g05909(.A1(new_n5889_), .A2(new_n513_), .A3(new_n3666_), .ZN(new_n6103_));
  NOR2_X1    g05910(.A1(new_n767_), .A2(new_n4343_), .ZN(new_n6104_));
  NOR2_X1    g05911(.A1(new_n6103_), .A2(new_n6104_), .ZN(new_n6105_));
  NOR2_X1    g05912(.A1(new_n6105_), .A2(new_n6102_), .ZN(new_n6106_));
  NAND2_X1   g05913(.A1(\a[14] ), .A2(\a[43] ), .ZN(new_n6107_));
  AOI22_X1   g05914(.A1(\a[11] ), .A2(\a[46] ), .B1(\a[13] ), .B2(\a[44] ), .ZN(new_n6108_));
  NOR2_X1    g05915(.A1(new_n6106_), .A2(new_n6102_), .ZN(new_n6109_));
  INV_X1     g05916(.I(new_n6109_), .ZN(new_n6110_));
  OAI22_X1   g05917(.A1(new_n6110_), .A2(new_n6108_), .B1(new_n6106_), .B2(new_n6107_), .ZN(new_n6111_));
  XNOR2_X1   g05918(.A1(new_n6111_), .A2(new_n6099_), .ZN(new_n6112_));
  NOR2_X1    g05919(.A1(new_n1023_), .A2(new_n5135_), .ZN(new_n6113_));
  NOR2_X1    g05920(.A1(new_n3116_), .A2(new_n5135_), .ZN(new_n6114_));
  NAND3_X1   g05921(.A1(new_n6114_), .A2(\a[6] ), .A3(\a[18] ), .ZN(new_n6115_));
  NAND2_X1   g05922(.A1(new_n1027_), .A2(new_n3550_), .ZN(new_n6116_));
  AOI22_X1   g05923(.A1(new_n6116_), .A2(new_n6115_), .B1(new_n4095_), .B2(new_n6113_), .ZN(new_n6117_));
  NAND2_X1   g05924(.A1(\a[18] ), .A2(\a[39] ), .ZN(new_n6118_));
  AOI22_X1   g05925(.A1(\a[6] ), .A2(\a[51] ), .B1(\a[17] ), .B2(\a[40] ), .ZN(new_n6119_));
  NAND2_X1   g05926(.A1(new_n4095_), .A2(new_n6113_), .ZN(new_n6120_));
  NAND3_X1   g05927(.A1(new_n6120_), .A2(new_n6116_), .A3(new_n6115_), .ZN(new_n6121_));
  OAI22_X1   g05928(.A1(new_n6117_), .A2(new_n6118_), .B1(new_n6121_), .B2(new_n6119_), .ZN(new_n6122_));
  XOR2_X1    g05929(.A1(new_n6112_), .A2(new_n6122_), .Z(new_n6123_));
  NOR2_X1    g05930(.A1(new_n5425_), .A2(new_n5680_), .ZN(new_n6124_));
  INV_X1     g05931(.I(new_n6124_), .ZN(new_n6125_));
  NOR2_X1    g05932(.A1(new_n5425_), .A2(new_n5617_), .ZN(new_n6126_));
  INV_X1     g05933(.I(new_n6126_), .ZN(new_n6127_));
  NOR2_X1    g05934(.A1(new_n5617_), .A2(new_n5680_), .ZN(new_n6128_));
  INV_X1     g05935(.I(new_n6128_), .ZN(new_n6129_));
  OAI22_X1   g05936(.A1(new_n246_), .A2(new_n6129_), .B1(new_n6127_), .B2(new_n370_), .ZN(new_n6130_));
  OAI21_X1   g05937(.A1(new_n251_), .A2(new_n6125_), .B(new_n6130_), .ZN(new_n6131_));
  NAND3_X1   g05938(.A1(new_n6131_), .A2(\a[3] ), .A3(\a[54] ), .ZN(new_n6132_));
  AOI22_X1   g05939(.A1(\a[2] ), .A2(\a[55] ), .B1(\a[4] ), .B2(\a[53] ), .ZN(new_n6133_));
  NOR2_X1    g05940(.A1(new_n6125_), .A2(new_n251_), .ZN(new_n6134_));
  NOR2_X1    g05941(.A1(new_n6130_), .A2(new_n6134_), .ZN(new_n6135_));
  INV_X1     g05942(.I(new_n6135_), .ZN(new_n6136_));
  OAI21_X1   g05943(.A1(new_n6133_), .A2(new_n6136_), .B(new_n6132_), .ZN(new_n6137_));
  AOI22_X1   g05944(.A1(\a[19] ), .A2(\a[38] ), .B1(\a[20] ), .B2(\a[37] ), .ZN(new_n6138_));
  INV_X1     g05945(.I(new_n6138_), .ZN(new_n6139_));
  INV_X1     g05946(.I(new_n3803_), .ZN(new_n6140_));
  NOR2_X1    g05947(.A1(new_n1376_), .A2(new_n6140_), .ZN(new_n6141_));
  NOR2_X1    g05948(.A1(new_n253_), .A2(new_n5175_), .ZN(new_n6142_));
  AOI21_X1   g05949(.A1(new_n6139_), .A2(new_n6142_), .B(new_n6141_), .ZN(new_n6143_));
  NAND2_X1   g05950(.A1(new_n6143_), .A2(new_n6139_), .ZN(new_n6144_));
  OAI21_X1   g05951(.A1(new_n6141_), .A2(new_n6138_), .B(new_n6142_), .ZN(new_n6145_));
  NAND2_X1   g05952(.A1(new_n6144_), .A2(new_n6145_), .ZN(new_n6146_));
  XNOR2_X1   g05953(.A1(new_n6137_), .A2(new_n6146_), .ZN(new_n6147_));
  AOI22_X1   g05954(.A1(\a[9] ), .A2(\a[48] ), .B1(\a[10] ), .B2(\a[47] ), .ZN(new_n6148_));
  NOR2_X1    g05955(.A1(new_n717_), .A2(new_n3746_), .ZN(new_n6149_));
  INV_X1     g05956(.I(new_n6149_), .ZN(new_n6150_));
  NOR2_X1    g05957(.A1(new_n4977_), .A2(new_n539_), .ZN(new_n6151_));
  NOR3_X1    g05958(.A1(new_n6151_), .A2(new_n6148_), .A3(new_n6150_), .ZN(new_n6152_));
  NOR2_X1    g05959(.A1(new_n6152_), .A2(new_n6151_), .ZN(new_n6153_));
  INV_X1     g05960(.I(new_n6153_), .ZN(new_n6154_));
  OAI22_X1   g05961(.A1(new_n6154_), .A2(new_n6148_), .B1(new_n6150_), .B2(new_n6152_), .ZN(new_n6155_));
  XOR2_X1    g05962(.A1(new_n6147_), .A2(new_n6155_), .Z(new_n6156_));
  XOR2_X1    g05963(.A1(new_n6123_), .A2(new_n6156_), .Z(new_n6157_));
  XOR2_X1    g05964(.A1(new_n6089_), .A2(new_n6157_), .Z(new_n6158_));
  NAND2_X1   g05965(.A1(new_n6007_), .A2(new_n6024_), .ZN(new_n6159_));
  NAND2_X1   g05966(.A1(new_n6025_), .A2(new_n6004_), .ZN(new_n6160_));
  NAND2_X1   g05967(.A1(new_n6160_), .A2(new_n6159_), .ZN(new_n6161_));
  NAND3_X1   g05968(.A1(new_n4664_), .A2(\a[16] ), .A3(\a[49] ), .ZN(new_n6162_));
  NOR3_X1    g05969(.A1(new_n4532_), .A2(new_n742_), .A3(new_n4901_), .ZN(new_n6163_));
  NOR2_X1    g05970(.A1(new_n5155_), .A2(new_n415_), .ZN(new_n6164_));
  OAI21_X1   g05971(.A1(new_n6163_), .A2(new_n6164_), .B(new_n6162_), .ZN(new_n6165_));
  NAND3_X1   g05972(.A1(new_n6165_), .A2(\a[7] ), .A3(\a[50] ), .ZN(new_n6166_));
  NAND2_X1   g05973(.A1(new_n6165_), .A2(new_n6162_), .ZN(new_n6167_));
  AOI22_X1   g05974(.A1(\a[8] ), .A2(\a[49] ), .B1(\a[16] ), .B2(\a[41] ), .ZN(new_n6168_));
  OAI21_X1   g05975(.A1(new_n6167_), .A2(new_n6168_), .B(new_n6166_), .ZN(new_n6169_));
  NOR2_X1    g05976(.A1(new_n2385_), .A2(new_n2746_), .ZN(new_n6170_));
  NOR2_X1    g05977(.A1(new_n1456_), .A2(new_n3405_), .ZN(new_n6171_));
  NOR2_X1    g05978(.A1(new_n1301_), .A2(new_n5564_), .ZN(new_n6172_));
  NOR2_X1    g05979(.A1(new_n6171_), .A2(new_n6172_), .ZN(new_n6173_));
  NOR2_X1    g05980(.A1(new_n6173_), .A2(new_n6170_), .ZN(new_n6174_));
  NAND2_X1   g05981(.A1(\a[21] ), .A2(\a[36] ), .ZN(new_n6175_));
  AOI22_X1   g05982(.A1(\a[22] ), .A2(\a[35] ), .B1(\a[23] ), .B2(\a[34] ), .ZN(new_n6176_));
  NOR2_X1    g05983(.A1(new_n6174_), .A2(new_n6170_), .ZN(new_n6177_));
  INV_X1     g05984(.I(new_n6177_), .ZN(new_n6178_));
  OAI22_X1   g05985(.A1(new_n6178_), .A2(new_n6176_), .B1(new_n6174_), .B2(new_n6175_), .ZN(new_n6179_));
  XOR2_X1    g05986(.A1(new_n6179_), .A2(new_n6169_), .Z(new_n6180_));
  OAI22_X1   g05987(.A1(new_n1779_), .A2(new_n2637_), .B1(new_n2081_), .B2(new_n2276_), .ZN(new_n6181_));
  OAI21_X1   g05988(.A1(new_n2177_), .A2(new_n3833_), .B(new_n6181_), .ZN(new_n6182_));
  NAND3_X1   g05989(.A1(new_n6182_), .A2(\a[24] ), .A3(\a[33] ), .ZN(new_n6183_));
  AOI22_X1   g05990(.A1(\a[25] ), .A2(\a[32] ), .B1(\a[26] ), .B2(\a[31] ), .ZN(new_n6184_));
  NOR2_X1    g05991(.A1(new_n2177_), .A2(new_n3833_), .ZN(new_n6185_));
  NOR2_X1    g05992(.A1(new_n6181_), .A2(new_n6185_), .ZN(new_n6186_));
  INV_X1     g05993(.I(new_n6186_), .ZN(new_n6187_));
  OAI21_X1   g05994(.A1(new_n6184_), .A2(new_n6187_), .B(new_n6183_), .ZN(new_n6188_));
  XNOR2_X1   g05995(.A1(new_n6180_), .A2(new_n6188_), .ZN(new_n6189_));
  INV_X1     g05996(.I(new_n6189_), .ZN(new_n6190_));
  INV_X1     g05997(.I(new_n6023_), .ZN(new_n6191_));
  NAND2_X1   g05998(.A1(new_n6191_), .A2(new_n6010_), .ZN(new_n6192_));
  OAI21_X1   g05999(.A1(new_n6013_), .A2(new_n6022_), .B(new_n6192_), .ZN(new_n6193_));
  XOR2_X1    g06000(.A1(new_n5895_), .A2(new_n6021_), .Z(new_n6194_));
  XOR2_X1    g06001(.A1(new_n6194_), .A2(new_n5914_), .Z(new_n6195_));
  NOR2_X1    g06002(.A1(new_n6193_), .A2(new_n6195_), .ZN(new_n6196_));
  NAND2_X1   g06003(.A1(new_n6193_), .A2(new_n6195_), .ZN(new_n6197_));
  INV_X1     g06004(.I(new_n6197_), .ZN(new_n6198_));
  NOR2_X1    g06005(.A1(new_n6198_), .A2(new_n6196_), .ZN(new_n6199_));
  NAND2_X1   g06006(.A1(new_n6199_), .A2(new_n6190_), .ZN(new_n6200_));
  INV_X1     g06007(.I(new_n6200_), .ZN(new_n6201_));
  NOR2_X1    g06008(.A1(new_n6199_), .A2(new_n6190_), .ZN(new_n6202_));
  NOR2_X1    g06009(.A1(new_n6201_), .A2(new_n6202_), .ZN(new_n6203_));
  XOR2_X1    g06010(.A1(new_n6161_), .A2(new_n6203_), .Z(new_n6204_));
  XNOR2_X1   g06011(.A1(new_n6204_), .A2(new_n6158_), .ZN(new_n6205_));
  XOR2_X1    g06012(.A1(new_n6088_), .A2(new_n6205_), .Z(new_n6206_));
  INV_X1     g06013(.I(new_n6206_), .ZN(new_n6207_));
  NOR2_X1    g06014(.A1(new_n5954_), .A2(new_n5995_), .ZN(new_n6208_));
  NOR2_X1    g06015(.A1(new_n5996_), .A2(new_n5952_), .ZN(new_n6209_));
  NOR2_X1    g06016(.A1(new_n6209_), .A2(new_n6208_), .ZN(new_n6210_));
  NAND2_X1   g06017(.A1(new_n5930_), .A2(new_n5950_), .ZN(new_n6211_));
  NAND2_X1   g06018(.A1(new_n5951_), .A2(new_n5928_), .ZN(new_n6212_));
  NAND2_X1   g06019(.A1(new_n6212_), .A2(new_n6211_), .ZN(new_n6213_));
  NAND2_X1   g06020(.A1(new_n5993_), .A2(new_n5989_), .ZN(new_n6214_));
  INV_X1     g06021(.I(new_n5960_), .ZN(new_n6215_));
  NOR2_X1    g06022(.A1(new_n6215_), .A2(new_n5826_), .ZN(new_n6216_));
  NOR2_X1    g06023(.A1(new_n6216_), .A2(new_n5959_), .ZN(new_n6217_));
  NAND2_X1   g06024(.A1(new_n5704_), .A2(new_n5697_), .ZN(new_n6218_));
  NAND2_X1   g06025(.A1(new_n5931_), .A2(new_n5813_), .ZN(new_n6219_));
  NAND2_X1   g06026(.A1(new_n6219_), .A2(new_n6218_), .ZN(new_n6220_));
  NAND2_X1   g06027(.A1(\a[0] ), .A2(\a[57] ), .ZN(new_n6221_));
  XOR2_X1    g06028(.A1(new_n5938_), .A2(new_n6221_), .Z(new_n6222_));
  NAND2_X1   g06029(.A1(\a[1] ), .A2(\a[56] ), .ZN(new_n6223_));
  XOR2_X1    g06030(.A1(new_n6223_), .A2(\a[29] ), .Z(new_n6224_));
  XNOR2_X1   g06031(.A1(new_n6222_), .A2(new_n6224_), .ZN(new_n6225_));
  XNOR2_X1   g06032(.A1(new_n6220_), .A2(new_n6225_), .ZN(new_n6226_));
  INV_X1     g06033(.I(new_n6226_), .ZN(new_n6227_));
  NAND2_X1   g06034(.A1(new_n6227_), .A2(new_n6217_), .ZN(new_n6228_));
  OAI21_X1   g06035(.A1(new_n5959_), .A2(new_n6216_), .B(new_n6226_), .ZN(new_n6229_));
  AND2_X2    g06036(.A1(new_n6228_), .A2(new_n6229_), .Z(new_n6230_));
  NAND2_X1   g06037(.A1(new_n5965_), .A2(new_n5961_), .ZN(new_n6231_));
  NAND2_X1   g06038(.A1(new_n5966_), .A2(new_n5957_), .ZN(new_n6232_));
  NAND2_X1   g06039(.A1(new_n6232_), .A2(new_n6231_), .ZN(new_n6233_));
  NAND2_X1   g06040(.A1(new_n5936_), .A2(new_n5948_), .ZN(new_n6234_));
  NAND2_X1   g06041(.A1(new_n5949_), .A2(new_n5932_), .ZN(new_n6235_));
  NAND2_X1   g06042(.A1(new_n6235_), .A2(new_n6234_), .ZN(new_n6236_));
  XOR2_X1    g06043(.A1(new_n6233_), .A2(new_n6236_), .Z(new_n6237_));
  XOR2_X1    g06044(.A1(new_n6237_), .A2(new_n6230_), .Z(new_n6238_));
  NOR2_X1    g06045(.A1(new_n6214_), .A2(new_n6238_), .ZN(new_n6239_));
  NAND2_X1   g06046(.A1(new_n6214_), .A2(new_n6238_), .ZN(new_n6240_));
  INV_X1     g06047(.I(new_n6240_), .ZN(new_n6241_));
  NOR2_X1    g06048(.A1(new_n6241_), .A2(new_n6239_), .ZN(new_n6242_));
  NOR2_X1    g06049(.A1(new_n6242_), .A2(new_n6213_), .ZN(new_n6243_));
  NAND2_X1   g06050(.A1(new_n6242_), .A2(new_n6213_), .ZN(new_n6244_));
  INV_X1     g06051(.I(new_n6244_), .ZN(new_n6245_));
  NOR2_X1    g06052(.A1(new_n6245_), .A2(new_n6243_), .ZN(new_n6246_));
  NOR2_X1    g06053(.A1(new_n6210_), .A2(new_n6246_), .ZN(new_n6247_));
  INV_X1     g06054(.I(new_n6246_), .ZN(new_n6248_));
  NOR2_X1    g06055(.A1(new_n6248_), .A2(new_n6210_), .ZN(new_n6249_));
  NOR2_X1    g06056(.A1(new_n6249_), .A2(new_n6248_), .ZN(new_n6250_));
  OAI21_X1   g06057(.A1(new_n6247_), .A2(new_n6250_), .B(new_n6207_), .ZN(new_n6251_));
  INV_X1     g06058(.I(new_n6251_), .ZN(new_n6252_));
  NOR3_X1    g06059(.A1(new_n6207_), .A2(new_n6250_), .A3(new_n6247_), .ZN(new_n6253_));
  NOR2_X1    g06060(.A1(new_n6252_), .A2(new_n6253_), .ZN(new_n6254_));
  NOR2_X1    g06061(.A1(new_n6254_), .A2(new_n6050_), .ZN(new_n6255_));
  NAND2_X1   g06062(.A1(new_n6254_), .A2(new_n6050_), .ZN(new_n6256_));
  INV_X1     g06063(.I(new_n6256_), .ZN(new_n6257_));
  NOR2_X1    g06064(.A1(new_n6257_), .A2(new_n6255_), .ZN(new_n6258_));
  XOR2_X1    g06065(.A1(new_n6048_), .A2(new_n6258_), .Z(\asquared[58] ));
  AOI21_X1   g06066(.A1(new_n6047_), .A2(new_n6043_), .B(new_n6255_), .ZN(new_n6260_));
  NOR2_X1    g06067(.A1(new_n6260_), .A2(new_n6257_), .ZN(new_n6261_));
  NOR2_X1    g06068(.A1(new_n6252_), .A2(new_n6249_), .ZN(new_n6262_));
  NOR2_X1    g06069(.A1(new_n6245_), .A2(new_n6241_), .ZN(new_n6263_));
  NAND2_X1   g06070(.A1(new_n6179_), .A2(new_n6169_), .ZN(new_n6264_));
  NAND2_X1   g06071(.A1(new_n6180_), .A2(new_n6188_), .ZN(new_n6265_));
  NAND2_X1   g06072(.A1(new_n6265_), .A2(new_n6264_), .ZN(new_n6266_));
  XOR2_X1    g06073(.A1(new_n6135_), .A2(new_n6143_), .Z(new_n6267_));
  NOR2_X1    g06074(.A1(new_n6267_), .A2(new_n6110_), .ZN(new_n6268_));
  INV_X1     g06075(.I(new_n6267_), .ZN(new_n6269_));
  NOR2_X1    g06076(.A1(new_n6269_), .A2(new_n6109_), .ZN(new_n6270_));
  NOR2_X1    g06077(.A1(new_n6270_), .A2(new_n6268_), .ZN(new_n6271_));
  NOR2_X1    g06078(.A1(new_n6154_), .A2(new_n6187_), .ZN(new_n6272_));
  NOR2_X1    g06079(.A1(new_n6153_), .A2(new_n6186_), .ZN(new_n6273_));
  NOR2_X1    g06080(.A1(new_n6272_), .A2(new_n6273_), .ZN(new_n6274_));
  NOR2_X1    g06081(.A1(new_n6274_), .A2(new_n6178_), .ZN(new_n6275_));
  INV_X1     g06082(.I(new_n6274_), .ZN(new_n6276_));
  NOR2_X1    g06083(.A1(new_n6276_), .A2(new_n6177_), .ZN(new_n6277_));
  NOR2_X1    g06084(.A1(new_n6277_), .A2(new_n6275_), .ZN(new_n6278_));
  NAND2_X1   g06085(.A1(new_n6278_), .A2(new_n6271_), .ZN(new_n6279_));
  INV_X1     g06086(.I(new_n6279_), .ZN(new_n6280_));
  NOR2_X1    g06087(.A1(new_n6278_), .A2(new_n6271_), .ZN(new_n6281_));
  NOR2_X1    g06088(.A1(new_n6280_), .A2(new_n6281_), .ZN(new_n6282_));
  NOR2_X1    g06089(.A1(new_n6282_), .A2(new_n6266_), .ZN(new_n6283_));
  NAND2_X1   g06090(.A1(new_n6282_), .A2(new_n6266_), .ZN(new_n6284_));
  INV_X1     g06091(.I(new_n6284_), .ZN(new_n6285_));
  NOR2_X1    g06092(.A1(new_n6285_), .A2(new_n6283_), .ZN(new_n6286_));
  INV_X1     g06093(.I(new_n6156_), .ZN(new_n6287_));
  NAND2_X1   g06094(.A1(new_n6123_), .A2(new_n6287_), .ZN(new_n6288_));
  OAI21_X1   g06095(.A1(new_n6089_), .A2(new_n6157_), .B(new_n6288_), .ZN(new_n6289_));
  OAI21_X1   g06096(.A1(new_n6097_), .A2(new_n6098_), .B(new_n6111_), .ZN(new_n6290_));
  NAND2_X1   g06097(.A1(new_n6112_), .A2(new_n6122_), .ZN(new_n6291_));
  NAND2_X1   g06098(.A1(new_n6291_), .A2(new_n6290_), .ZN(new_n6292_));
  NAND2_X1   g06099(.A1(new_n6137_), .A2(new_n6146_), .ZN(new_n6293_));
  INV_X1     g06100(.I(new_n6155_), .ZN(new_n6294_));
  OAI21_X1   g06101(.A1(new_n6147_), .A2(new_n6294_), .B(new_n6293_), .ZN(new_n6295_));
  INV_X1     g06102(.I(new_n6295_), .ZN(new_n6296_));
  NOR2_X1    g06103(.A1(new_n6223_), .A2(new_n1814_), .ZN(new_n6297_));
  INV_X1     g06104(.I(\a[57] ), .ZN(new_n6298_));
  NOR3_X1    g06105(.A1(new_n3811_), .A2(new_n194_), .A3(new_n6298_), .ZN(new_n6299_));
  AOI21_X1   g06106(.A1(\a[1] ), .A2(\a[57] ), .B(new_n2681_), .ZN(new_n6300_));
  NOR2_X1    g06107(.A1(new_n6299_), .A2(new_n6300_), .ZN(new_n6301_));
  XOR2_X1    g06108(.A1(new_n6301_), .A2(new_n6297_), .Z(new_n6302_));
  XOR2_X1    g06109(.A1(new_n6302_), .A2(new_n6096_), .Z(new_n6303_));
  NOR2_X1    g06110(.A1(new_n6296_), .A2(new_n6303_), .ZN(new_n6304_));
  INV_X1     g06111(.I(new_n6303_), .ZN(new_n6305_));
  NOR2_X1    g06112(.A1(new_n6295_), .A2(new_n6305_), .ZN(new_n6306_));
  OAI21_X1   g06113(.A1(new_n6304_), .A2(new_n6306_), .B(new_n6292_), .ZN(new_n6307_));
  INV_X1     g06114(.I(new_n6307_), .ZN(new_n6308_));
  NOR3_X1    g06115(.A1(new_n6304_), .A2(new_n6292_), .A3(new_n6306_), .ZN(new_n6309_));
  NOR2_X1    g06116(.A1(new_n6308_), .A2(new_n6309_), .ZN(new_n6310_));
  XOR2_X1    g06117(.A1(new_n6289_), .A2(new_n6310_), .Z(new_n6311_));
  XOR2_X1    g06118(.A1(new_n6311_), .A2(new_n6286_), .Z(new_n6312_));
  XNOR2_X1   g06119(.A1(new_n6263_), .A2(new_n6312_), .ZN(new_n6313_));
  NOR2_X1    g06120(.A1(new_n6073_), .A2(new_n6077_), .ZN(new_n6314_));
  NOR2_X1    g06121(.A1(new_n6081_), .A2(new_n6314_), .ZN(new_n6315_));
  INV_X1     g06122(.I(\a[58] ), .ZN(new_n6316_));
  NOR2_X1    g06123(.A1(new_n5856_), .A2(new_n6316_), .ZN(new_n6317_));
  INV_X1     g06124(.I(new_n6317_), .ZN(new_n6318_));
  OAI22_X1   g06125(.A1(new_n412_), .A2(new_n6318_), .B1(new_n6058_), .B2(new_n251_), .ZN(new_n6319_));
  NOR2_X1    g06126(.A1(new_n290_), .A2(new_n5617_), .ZN(new_n6320_));
  NOR2_X1    g06127(.A1(new_n196_), .A2(new_n6316_), .ZN(new_n6321_));
  NAND2_X1   g06128(.A1(new_n6320_), .A2(new_n6321_), .ZN(new_n6322_));
  NAND2_X1   g06129(.A1(new_n6319_), .A2(new_n6322_), .ZN(new_n6323_));
  NAND3_X1   g06130(.A1(new_n6323_), .A2(\a[2] ), .A3(\a[56] ), .ZN(new_n6324_));
  NOR2_X1    g06131(.A1(new_n6320_), .A2(new_n6321_), .ZN(new_n6325_));
  NAND2_X1   g06132(.A1(new_n6323_), .A2(new_n6322_), .ZN(new_n6326_));
  OAI21_X1   g06133(.A1(new_n6325_), .A2(new_n6326_), .B(new_n6324_), .ZN(new_n6327_));
  AOI22_X1   g06134(.A1(\a[20] ), .A2(\a[38] ), .B1(\a[21] ), .B2(\a[37] ), .ZN(new_n6328_));
  INV_X1     g06135(.I(new_n6328_), .ZN(new_n6329_));
  NOR2_X1    g06136(.A1(new_n1382_), .A2(new_n6140_), .ZN(new_n6330_));
  NOR2_X1    g06137(.A1(new_n253_), .A2(new_n5425_), .ZN(new_n6331_));
  AOI21_X1   g06138(.A1(new_n6329_), .A2(new_n6331_), .B(new_n6330_), .ZN(new_n6332_));
  NAND2_X1   g06139(.A1(new_n6332_), .A2(new_n6329_), .ZN(new_n6333_));
  OAI21_X1   g06140(.A1(new_n6330_), .A2(new_n6328_), .B(new_n6331_), .ZN(new_n6334_));
  NAND2_X1   g06141(.A1(new_n6333_), .A2(new_n6334_), .ZN(new_n6335_));
  XOR2_X1    g06142(.A1(new_n6327_), .A2(new_n6335_), .Z(new_n6336_));
  NOR2_X1    g06143(.A1(new_n3746_), .A2(new_n4702_), .ZN(new_n6337_));
  INV_X1     g06144(.I(new_n6337_), .ZN(new_n6338_));
  NOR2_X1    g06145(.A1(new_n6338_), .A2(new_n798_), .ZN(new_n6339_));
  NOR2_X1    g06146(.A1(new_n1023_), .A2(new_n4702_), .ZN(new_n6340_));
  NAND3_X1   g06147(.A1(new_n6340_), .A2(\a[9] ), .A3(\a[41] ), .ZN(new_n6341_));
  NAND2_X1   g06148(.A1(new_n1024_), .A2(new_n4372_), .ZN(new_n6342_));
  AOI21_X1   g06149(.A1(new_n6342_), .A2(new_n6341_), .B(new_n6339_), .ZN(new_n6343_));
  NAND2_X1   g06150(.A1(\a[17] ), .A2(\a[41] ), .ZN(new_n6344_));
  AOI22_X1   g06151(.A1(\a[9] ), .A2(\a[49] ), .B1(\a[16] ), .B2(\a[42] ), .ZN(new_n6345_));
  OR2_X2     g06152(.A1(new_n6343_), .A2(new_n6339_), .Z(new_n6346_));
  OAI22_X1   g06153(.A1(new_n6346_), .A2(new_n6345_), .B1(new_n6343_), .B2(new_n6344_), .ZN(new_n6347_));
  XOR2_X1    g06154(.A1(new_n6336_), .A2(new_n6347_), .Z(new_n6348_));
  AOI22_X1   g06155(.A1(\a[7] ), .A2(\a[51] ), .B1(\a[8] ), .B2(\a[50] ), .ZN(new_n6349_));
  NOR2_X1    g06156(.A1(new_n884_), .A2(new_n3221_), .ZN(new_n6350_));
  INV_X1     g06157(.I(new_n6350_), .ZN(new_n6351_));
  OAI22_X1   g06158(.A1(new_n415_), .A2(new_n5440_), .B1(new_n6351_), .B2(new_n6349_), .ZN(new_n6352_));
  NOR2_X1    g06159(.A1(new_n5440_), .A2(new_n415_), .ZN(new_n6353_));
  OAI21_X1   g06160(.A1(new_n6353_), .A2(new_n6349_), .B(new_n6350_), .ZN(new_n6354_));
  OAI21_X1   g06161(.A1(new_n6352_), .A2(new_n6349_), .B(new_n6354_), .ZN(new_n6355_));
  OAI22_X1   g06162(.A1(new_n2385_), .A2(new_n3405_), .B1(new_n1880_), .B2(new_n5564_), .ZN(new_n6356_));
  OAI21_X1   g06163(.A1(new_n1529_), .A2(new_n2746_), .B(new_n6356_), .ZN(new_n6357_));
  NAND3_X1   g06164(.A1(new_n6357_), .A2(\a[22] ), .A3(\a[36] ), .ZN(new_n6358_));
  AOI22_X1   g06165(.A1(\a[23] ), .A2(\a[35] ), .B1(\a[24] ), .B2(\a[34] ), .ZN(new_n6359_));
  NOR2_X1    g06166(.A1(new_n1529_), .A2(new_n2746_), .ZN(new_n6360_));
  NOR2_X1    g06167(.A1(new_n6356_), .A2(new_n6360_), .ZN(new_n6361_));
  INV_X1     g06168(.I(new_n6361_), .ZN(new_n6362_));
  OAI21_X1   g06169(.A1(new_n6359_), .A2(new_n6362_), .B(new_n6358_), .ZN(new_n6363_));
  XOR2_X1    g06170(.A1(new_n6363_), .A2(new_n6355_), .Z(new_n6364_));
  NOR2_X1    g06171(.A1(new_n1972_), .A2(new_n3833_), .ZN(new_n6365_));
  AOI22_X1   g06172(.A1(new_n2176_), .A2(new_n2636_), .B1(new_n2246_), .B2(new_n2275_), .ZN(new_n6366_));
  NOR2_X1    g06173(.A1(new_n6365_), .A2(new_n6366_), .ZN(new_n6367_));
  AOI21_X1   g06174(.A1(\a[27] ), .A2(\a[31] ), .B(new_n2782_), .ZN(new_n6368_));
  NOR2_X1    g06175(.A1(new_n6367_), .A2(new_n6365_), .ZN(new_n6369_));
  INV_X1     g06176(.I(new_n6369_), .ZN(new_n6370_));
  OAI22_X1   g06177(.A1(new_n6370_), .A2(new_n6368_), .B1(new_n2754_), .B2(new_n6367_), .ZN(new_n6371_));
  XOR2_X1    g06178(.A1(new_n6364_), .A2(new_n6371_), .Z(new_n6372_));
  XNOR2_X1   g06179(.A1(new_n6372_), .A2(new_n6348_), .ZN(new_n6373_));
  XOR2_X1    g06180(.A1(new_n6315_), .A2(new_n6373_), .Z(new_n6374_));
  NAND2_X1   g06181(.A1(new_n6233_), .A2(new_n6236_), .ZN(new_n6375_));
  NAND2_X1   g06182(.A1(new_n6237_), .A2(new_n6230_), .ZN(new_n6376_));
  NAND2_X1   g06183(.A1(new_n6376_), .A2(new_n6375_), .ZN(new_n6377_));
  NAND3_X1   g06184(.A1(new_n832_), .A2(\a[43] ), .A3(\a[47] ), .ZN(new_n6378_));
  INV_X1     g06185(.I(new_n5917_), .ZN(new_n6379_));
  NOR3_X1    g06186(.A1(new_n6379_), .A2(new_n417_), .A3(new_n3666_), .ZN(new_n6380_));
  NOR2_X1    g06187(.A1(new_n1264_), .A2(new_n4977_), .ZN(new_n6381_));
  OAI21_X1   g06188(.A1(new_n6380_), .A2(new_n6381_), .B(new_n6378_), .ZN(new_n6382_));
  NAND3_X1   g06189(.A1(new_n6382_), .A2(\a[10] ), .A3(\a[48] ), .ZN(new_n6383_));
  NAND2_X1   g06190(.A1(new_n6382_), .A2(new_n6378_), .ZN(new_n6384_));
  NOR2_X1    g06191(.A1(new_n513_), .A2(new_n4312_), .ZN(new_n6385_));
  AOI21_X1   g06192(.A1(\a[15] ), .A2(\a[43] ), .B(new_n6385_), .ZN(new_n6386_));
  OAI21_X1   g06193(.A1(new_n6384_), .A2(new_n6386_), .B(new_n6383_), .ZN(new_n6387_));
  INV_X1     g06194(.I(new_n5405_), .ZN(new_n6388_));
  NAND2_X1   g06195(.A1(new_n760_), .A2(new_n4703_), .ZN(new_n6389_));
  NAND2_X1   g06196(.A1(new_n6100_), .A2(new_n762_), .ZN(new_n6390_));
  AOI22_X1   g06197(.A1(new_n6389_), .A2(new_n6390_), .B1(new_n763_), .B2(new_n4429_), .ZN(new_n6391_));
  AOI22_X1   g06198(.A1(\a[12] ), .A2(\a[46] ), .B1(\a[13] ), .B2(\a[45] ), .ZN(new_n6392_));
  NAND2_X1   g06199(.A1(new_n763_), .A2(new_n4429_), .ZN(new_n6393_));
  NAND3_X1   g06200(.A1(new_n6393_), .A2(new_n6389_), .A3(new_n6390_), .ZN(new_n6394_));
  OAI22_X1   g06201(.A1(new_n6391_), .A2(new_n6388_), .B1(new_n6394_), .B2(new_n6392_), .ZN(new_n6395_));
  XOR2_X1    g06202(.A1(new_n6387_), .A2(new_n6395_), .Z(new_n6396_));
  NOR2_X1    g06203(.A1(new_n225_), .A2(new_n5680_), .ZN(new_n6397_));
  INV_X1     g06204(.I(new_n6397_), .ZN(new_n6398_));
  AOI22_X1   g06205(.A1(\a[6] ), .A2(\a[52] ), .B1(\a[19] ), .B2(\a[39] ), .ZN(new_n6399_));
  NOR4_X1    g06206(.A1(new_n367_), .A2(new_n979_), .A3(new_n3116_), .A4(new_n5175_), .ZN(new_n6400_));
  NOR3_X1    g06207(.A1(new_n6398_), .A2(new_n6400_), .A3(new_n6399_), .ZN(new_n6401_));
  NOR2_X1    g06208(.A1(new_n6401_), .A2(new_n6400_), .ZN(new_n6402_));
  INV_X1     g06209(.I(new_n6402_), .ZN(new_n6403_));
  OAI22_X1   g06210(.A1(new_n6403_), .A2(new_n6399_), .B1(new_n6398_), .B2(new_n6401_), .ZN(new_n6404_));
  XNOR2_X1   g06211(.A1(new_n6396_), .A2(new_n6404_), .ZN(new_n6405_));
  INV_X1     g06212(.I(new_n6405_), .ZN(new_n6406_));
  INV_X1     g06213(.I(new_n6225_), .ZN(new_n6407_));
  NAND2_X1   g06214(.A1(new_n6407_), .A2(new_n6220_), .ZN(new_n6408_));
  NAND2_X1   g06215(.A1(new_n6229_), .A2(new_n6408_), .ZN(new_n6409_));
  NOR2_X1    g06216(.A1(new_n5939_), .A2(new_n6221_), .ZN(new_n6410_));
  NOR2_X1    g06217(.A1(new_n6222_), .A2(new_n6224_), .ZN(new_n6411_));
  NOR2_X1    g06218(.A1(new_n6411_), .A2(new_n6410_), .ZN(new_n6412_));
  XOR2_X1    g06219(.A1(new_n6167_), .A2(new_n6121_), .Z(new_n6413_));
  XNOR2_X1   g06220(.A1(new_n6413_), .A2(new_n6412_), .ZN(new_n6414_));
  NOR2_X1    g06221(.A1(new_n6409_), .A2(new_n6414_), .ZN(new_n6415_));
  NAND2_X1   g06222(.A1(new_n6409_), .A2(new_n6414_), .ZN(new_n6416_));
  INV_X1     g06223(.I(new_n6416_), .ZN(new_n6417_));
  NOR2_X1    g06224(.A1(new_n6417_), .A2(new_n6415_), .ZN(new_n6418_));
  NAND2_X1   g06225(.A1(new_n6418_), .A2(new_n6406_), .ZN(new_n6419_));
  INV_X1     g06226(.I(new_n6419_), .ZN(new_n6420_));
  NOR2_X1    g06227(.A1(new_n6418_), .A2(new_n6406_), .ZN(new_n6421_));
  NOR2_X1    g06228(.A1(new_n6420_), .A2(new_n6421_), .ZN(new_n6422_));
  XOR2_X1    g06229(.A1(new_n6377_), .A2(new_n6422_), .Z(new_n6423_));
  XNOR2_X1   g06230(.A1(new_n6423_), .A2(new_n6374_), .ZN(new_n6424_));
  XOR2_X1    g06231(.A1(new_n6313_), .A2(new_n6424_), .Z(new_n6425_));
  INV_X1     g06232(.I(new_n6425_), .ZN(new_n6426_));
  NAND2_X1   g06233(.A1(new_n6052_), .A2(new_n6087_), .ZN(new_n6427_));
  INV_X1     g06234(.I(new_n6088_), .ZN(new_n6428_));
  OAI21_X1   g06235(.A1(new_n6428_), .A2(new_n6205_), .B(new_n6427_), .ZN(new_n6429_));
  AND2_X2    g06236(.A1(new_n6161_), .A2(new_n6203_), .Z(new_n6430_));
  AOI21_X1   g06237(.A1(new_n6204_), .A2(new_n6158_), .B(new_n6430_), .ZN(new_n6431_));
  NAND2_X1   g06238(.A1(new_n6085_), .A2(new_n6082_), .ZN(new_n6432_));
  NAND2_X1   g06239(.A1(new_n6086_), .A2(new_n6069_), .ZN(new_n6433_));
  NAND2_X1   g06240(.A1(new_n6433_), .A2(new_n6432_), .ZN(new_n6434_));
  NOR2_X1    g06241(.A1(new_n6201_), .A2(new_n6198_), .ZN(new_n6435_));
  NOR2_X1    g06242(.A1(new_n6068_), .A2(new_n6063_), .ZN(new_n6436_));
  NAND2_X1   g06243(.A1(new_n5877_), .A2(new_n5923_), .ZN(new_n6437_));
  NAND2_X1   g06244(.A1(new_n6056_), .A2(new_n5907_), .ZN(new_n6438_));
  NAND2_X1   g06245(.A1(new_n6438_), .A2(new_n6437_), .ZN(new_n6439_));
  NAND2_X1   g06246(.A1(new_n6194_), .A2(new_n5914_), .ZN(new_n6440_));
  OAI21_X1   g06247(.A1(new_n5895_), .A2(new_n6021_), .B(new_n6440_), .ZN(new_n6441_));
  NAND2_X1   g06248(.A1(new_n5869_), .A2(new_n5883_), .ZN(new_n6442_));
  NAND2_X1   g06249(.A1(new_n6060_), .A2(new_n6059_), .ZN(new_n6443_));
  NAND2_X1   g06250(.A1(new_n6443_), .A2(new_n6442_), .ZN(new_n6444_));
  XOR2_X1    g06251(.A1(new_n6444_), .A2(new_n6441_), .Z(new_n6445_));
  XNOR2_X1   g06252(.A1(new_n6445_), .A2(new_n6439_), .ZN(new_n6446_));
  XOR2_X1    g06253(.A1(new_n6436_), .A2(new_n6446_), .Z(new_n6447_));
  INV_X1     g06254(.I(new_n6447_), .ZN(new_n6448_));
  XOR2_X1    g06255(.A1(new_n6435_), .A2(new_n6448_), .Z(new_n6449_));
  XNOR2_X1   g06256(.A1(new_n6449_), .A2(new_n6434_), .ZN(new_n6450_));
  XOR2_X1    g06257(.A1(new_n6431_), .A2(new_n6450_), .Z(new_n6451_));
  NOR2_X1    g06258(.A1(new_n6429_), .A2(new_n6451_), .ZN(new_n6452_));
  NAND2_X1   g06259(.A1(new_n6429_), .A2(new_n6451_), .ZN(new_n6453_));
  INV_X1     g06260(.I(new_n6453_), .ZN(new_n6454_));
  NOR2_X1    g06261(.A1(new_n6454_), .A2(new_n6452_), .ZN(new_n6455_));
  NOR2_X1    g06262(.A1(new_n6426_), .A2(new_n6455_), .ZN(new_n6456_));
  NAND2_X1   g06263(.A1(new_n6426_), .A2(new_n6455_), .ZN(new_n6457_));
  INV_X1     g06264(.I(new_n6457_), .ZN(new_n6458_));
  NOR2_X1    g06265(.A1(new_n6458_), .A2(new_n6456_), .ZN(new_n6459_));
  INV_X1     g06266(.I(new_n6459_), .ZN(new_n6460_));
  NOR2_X1    g06267(.A1(new_n6460_), .A2(new_n6262_), .ZN(new_n6461_));
  INV_X1     g06268(.I(new_n6461_), .ZN(new_n6462_));
  NAND2_X1   g06269(.A1(new_n6460_), .A2(new_n6262_), .ZN(new_n6463_));
  NAND2_X1   g06270(.A1(new_n6462_), .A2(new_n6463_), .ZN(new_n6464_));
  INV_X1     g06271(.I(new_n5847_), .ZN(new_n6465_));
  INV_X1     g06272(.I(new_n5477_), .ZN(new_n6466_));
  OAI21_X1   g06273(.A1(new_n5305_), .A2(new_n5297_), .B(new_n5478_), .ZN(new_n6467_));
  AOI21_X1   g06274(.A1(new_n6467_), .A2(new_n6466_), .B(new_n5655_), .ZN(new_n6468_));
  INV_X1     g06275(.I(new_n5848_), .ZN(new_n6469_));
  OAI21_X1   g06276(.A1(new_n6468_), .A2(new_n5657_), .B(new_n6469_), .ZN(new_n6470_));
  INV_X1     g06277(.I(new_n6044_), .ZN(new_n6471_));
  AOI21_X1   g06278(.A1(new_n6470_), .A2(new_n6465_), .B(new_n6471_), .ZN(new_n6472_));
  INV_X1     g06279(.I(new_n6255_), .ZN(new_n6473_));
  OAI21_X1   g06280(.A1(new_n6472_), .A2(new_n6042_), .B(new_n6473_), .ZN(new_n6474_));
  INV_X1     g06281(.I(new_n6463_), .ZN(new_n6475_));
  AOI21_X1   g06282(.A1(new_n6474_), .A2(new_n6256_), .B(new_n6475_), .ZN(new_n6476_));
  AOI22_X1   g06283(.A1(new_n6476_), .A2(new_n6462_), .B1(new_n6261_), .B2(new_n6464_), .ZN(\asquared[59] ));
  OAI21_X1   g06284(.A1(new_n6260_), .A2(new_n6257_), .B(new_n6463_), .ZN(new_n6478_));
  NAND2_X1   g06285(.A1(new_n6478_), .A2(new_n6462_), .ZN(new_n6479_));
  NOR2_X1    g06286(.A1(new_n6436_), .A2(new_n6446_), .ZN(new_n6480_));
  NOR2_X1    g06287(.A1(new_n6435_), .A2(new_n6448_), .ZN(new_n6481_));
  NOR2_X1    g06288(.A1(new_n6481_), .A2(new_n6480_), .ZN(new_n6482_));
  OAI21_X1   g06289(.A1(new_n6296_), .A2(new_n6305_), .B(new_n6307_), .ZN(new_n6483_));
  NOR4_X1    g06290(.A1(new_n253_), .A2(new_n979_), .A3(new_n3221_), .A4(new_n5617_), .ZN(new_n6484_));
  NAND4_X1   g06291(.A1(\a[4] ), .A2(\a[19] ), .A3(\a[40] ), .A4(\a[55] ), .ZN(new_n6485_));
  NAND2_X1   g06292(.A1(new_n6128_), .A2(new_n243_), .ZN(new_n6486_));
  AOI21_X1   g06293(.A1(new_n6486_), .A2(new_n6485_), .B(new_n6484_), .ZN(new_n6487_));
  NAND2_X1   g06294(.A1(\a[4] ), .A2(\a[55] ), .ZN(new_n6488_));
  OR2_X2     g06295(.A1(new_n6487_), .A2(new_n6484_), .Z(new_n6489_));
  AOI22_X1   g06296(.A1(\a[5] ), .A2(\a[54] ), .B1(\a[19] ), .B2(\a[40] ), .ZN(new_n6490_));
  OAI22_X1   g06297(.A1(new_n6489_), .A2(new_n6490_), .B1(new_n6487_), .B2(new_n6488_), .ZN(new_n6491_));
  AOI22_X1   g06298(.A1(\a[2] ), .A2(\a[57] ), .B1(\a[3] ), .B2(\a[56] ), .ZN(new_n6492_));
  INV_X1     g06299(.I(new_n6299_), .ZN(new_n6493_));
  NOR2_X1    g06300(.A1(new_n5856_), .A2(new_n6298_), .ZN(new_n6494_));
  NAND2_X1   g06301(.A1(new_n6494_), .A2(new_n256_), .ZN(new_n6495_));
  OAI21_X1   g06302(.A1(new_n6493_), .A2(new_n6492_), .B(new_n6495_), .ZN(new_n6496_));
  NOR2_X1    g06303(.A1(new_n6496_), .A2(new_n6492_), .ZN(new_n6497_));
  INV_X1     g06304(.I(new_n6492_), .ZN(new_n6498_));
  AOI21_X1   g06305(.A1(new_n6498_), .A2(new_n6495_), .B(new_n6493_), .ZN(new_n6499_));
  NOR2_X1    g06306(.A1(new_n6497_), .A2(new_n6499_), .ZN(new_n6500_));
  XOR2_X1    g06307(.A1(new_n6500_), .A2(new_n6370_), .Z(new_n6501_));
  XNOR2_X1   g06308(.A1(new_n6501_), .A2(new_n6491_), .ZN(new_n6502_));
  AOI21_X1   g06309(.A1(\a[28] ), .A2(\a[31] ), .B(new_n2254_), .ZN(new_n6503_));
  INV_X1     g06310(.I(new_n6503_), .ZN(new_n6504_));
  NOR3_X1    g06311(.A1(new_n2255_), .A2(new_n1718_), .A3(new_n2051_), .ZN(new_n6505_));
  NOR2_X1    g06312(.A1(new_n597_), .A2(new_n4178_), .ZN(new_n6506_));
  AOI21_X1   g06313(.A1(new_n6504_), .A2(new_n6506_), .B(new_n6505_), .ZN(new_n6507_));
  INV_X1     g06314(.I(new_n6507_), .ZN(new_n6508_));
  OAI21_X1   g06315(.A1(new_n6505_), .A2(new_n6503_), .B(new_n6506_), .ZN(new_n6509_));
  OAI21_X1   g06316(.A1(new_n6508_), .A2(new_n6503_), .B(new_n6509_), .ZN(new_n6510_));
  NOR2_X1    g06317(.A1(new_n4314_), .A2(new_n623_), .ZN(new_n6511_));
  NAND3_X1   g06318(.A1(new_n1482_), .A2(\a[45] ), .A3(\a[48] ), .ZN(new_n6512_));
  NOR2_X1    g06319(.A1(new_n4977_), .A2(new_n619_), .ZN(new_n6513_));
  INV_X1     g06320(.I(new_n6513_), .ZN(new_n6514_));
  AOI21_X1   g06321(.A1(new_n6514_), .A2(new_n6512_), .B(new_n6511_), .ZN(new_n6515_));
  NAND2_X1   g06322(.A1(\a[11] ), .A2(\a[48] ), .ZN(new_n6516_));
  AOI22_X1   g06323(.A1(\a[12] ), .A2(\a[47] ), .B1(\a[14] ), .B2(\a[45] ), .ZN(new_n6517_));
  NOR2_X1    g06324(.A1(new_n6515_), .A2(new_n6511_), .ZN(new_n6518_));
  INV_X1     g06325(.I(new_n6518_), .ZN(new_n6519_));
  OAI22_X1   g06326(.A1(new_n6519_), .A2(new_n6517_), .B1(new_n6515_), .B2(new_n6516_), .ZN(new_n6520_));
  XOR2_X1    g06327(.A1(new_n6520_), .A2(new_n6510_), .Z(new_n6521_));
  AOI22_X1   g06328(.A1(\a[16] ), .A2(\a[43] ), .B1(\a[17] ), .B2(\a[42] ), .ZN(new_n6522_));
  NAND2_X1   g06329(.A1(\a[8] ), .A2(\a[51] ), .ZN(new_n6523_));
  NOR2_X1    g06330(.A1(new_n1428_), .A2(new_n4181_), .ZN(new_n6524_));
  NOR3_X1    g06331(.A1(new_n6524_), .A2(new_n6522_), .A3(new_n6523_), .ZN(new_n6525_));
  NOR2_X1    g06332(.A1(new_n6525_), .A2(new_n6524_), .ZN(new_n6526_));
  INV_X1     g06333(.I(new_n6526_), .ZN(new_n6527_));
  OAI22_X1   g06334(.A1(new_n6527_), .A2(new_n6522_), .B1(new_n6523_), .B2(new_n6525_), .ZN(new_n6528_));
  XOR2_X1    g06335(.A1(new_n6521_), .A2(new_n6528_), .Z(new_n6529_));
  XOR2_X1    g06336(.A1(new_n6529_), .A2(new_n6502_), .Z(new_n6530_));
  XNOR2_X1   g06337(.A1(new_n6483_), .A2(new_n6530_), .ZN(new_n6531_));
  XOR2_X1    g06338(.A1(new_n6482_), .A2(new_n6531_), .Z(new_n6532_));
  NAND2_X1   g06339(.A1(new_n1452_), .A2(new_n3803_), .ZN(new_n6533_));
  OAI22_X1   g06340(.A1(new_n1382_), .A2(new_n4210_), .B1(new_n2647_), .B2(new_n4739_), .ZN(new_n6534_));
  NAND2_X1   g06341(.A1(new_n6534_), .A2(new_n6533_), .ZN(new_n6535_));
  NAND3_X1   g06342(.A1(new_n6535_), .A2(\a[20] ), .A3(\a[39] ), .ZN(new_n6536_));
  AOI22_X1   g06343(.A1(\a[21] ), .A2(\a[38] ), .B1(\a[22] ), .B2(\a[37] ), .ZN(new_n6537_));
  NAND2_X1   g06344(.A1(new_n6535_), .A2(new_n6533_), .ZN(new_n6538_));
  OAI21_X1   g06345(.A1(new_n6537_), .A2(new_n6538_), .B(new_n6536_), .ZN(new_n6539_));
  NAND2_X1   g06346(.A1(new_n1778_), .A2(new_n2745_), .ZN(new_n6540_));
  OAI22_X1   g06347(.A1(new_n1443_), .A2(new_n5564_), .B1(new_n1529_), .B2(new_n3405_), .ZN(new_n6541_));
  NAND2_X1   g06348(.A1(new_n6541_), .A2(new_n6540_), .ZN(new_n6542_));
  NAND3_X1   g06349(.A1(new_n6542_), .A2(\a[23] ), .A3(\a[36] ), .ZN(new_n6543_));
  AOI22_X1   g06350(.A1(\a[24] ), .A2(\a[35] ), .B1(\a[25] ), .B2(\a[34] ), .ZN(new_n6544_));
  NAND2_X1   g06351(.A1(new_n6542_), .A2(new_n6540_), .ZN(new_n6545_));
  OAI21_X1   g06352(.A1(new_n6544_), .A2(new_n6545_), .B(new_n6543_), .ZN(new_n6546_));
  XNOR2_X1   g06353(.A1(new_n6539_), .A2(new_n6546_), .ZN(new_n6547_));
  INV_X1     g06354(.I(\a[59] ), .ZN(new_n6548_));
  NOR3_X1    g06355(.A1(new_n1659_), .A2(new_n2200_), .A3(new_n6548_), .ZN(new_n6549_));
  NAND4_X1   g06356(.A1(\a[0] ), .A2(\a[26] ), .A3(\a[33] ), .A4(\a[59] ), .ZN(new_n6550_));
  NAND2_X1   g06357(.A1(new_n1971_), .A2(new_n2636_), .ZN(new_n6551_));
  AOI21_X1   g06358(.A1(new_n6551_), .A2(new_n6550_), .B(new_n6549_), .ZN(new_n6552_));
  NAND2_X1   g06359(.A1(\a[26] ), .A2(\a[33] ), .ZN(new_n6553_));
  OR2_X2     g06360(.A1(new_n6552_), .A2(new_n6549_), .Z(new_n6554_));
  AOI22_X1   g06361(.A1(\a[0] ), .A2(\a[59] ), .B1(\a[27] ), .B2(\a[32] ), .ZN(new_n6555_));
  OAI22_X1   g06362(.A1(new_n6554_), .A2(new_n6555_), .B1(new_n6552_), .B2(new_n6553_), .ZN(new_n6556_));
  XOR2_X1    g06363(.A1(new_n6547_), .A2(new_n6556_), .Z(new_n6557_));
  NAND2_X1   g06364(.A1(new_n6301_), .A2(new_n6297_), .ZN(new_n6558_));
  NAND2_X1   g06365(.A1(new_n6302_), .A2(new_n6096_), .ZN(new_n6559_));
  NAND2_X1   g06366(.A1(new_n6559_), .A2(new_n6558_), .ZN(new_n6560_));
  NOR2_X1    g06367(.A1(new_n884_), .A2(new_n5175_), .ZN(new_n6561_));
  INV_X1     g06368(.I(new_n6561_), .ZN(new_n6562_));
  INV_X1     g06369(.I(new_n5862_), .ZN(new_n6563_));
  NAND4_X1   g06370(.A1(\a[6] ), .A2(\a[18] ), .A3(\a[41] ), .A4(\a[53] ), .ZN(new_n6564_));
  OAI21_X1   g06371(.A1(new_n6563_), .A2(new_n374_), .B(new_n6564_), .ZN(new_n6565_));
  OAI21_X1   g06372(.A1(new_n4532_), .A2(new_n6562_), .B(new_n6565_), .ZN(new_n6566_));
  NAND3_X1   g06373(.A1(new_n6566_), .A2(\a[6] ), .A3(\a[53] ), .ZN(new_n6567_));
  NOR2_X1    g06374(.A1(new_n4532_), .A2(new_n6562_), .ZN(new_n6568_));
  NOR2_X1    g06375(.A1(new_n6565_), .A2(new_n6568_), .ZN(new_n6569_));
  INV_X1     g06376(.I(new_n6569_), .ZN(new_n6570_));
  AOI22_X1   g06377(.A1(\a[7] ), .A2(\a[52] ), .B1(\a[18] ), .B2(\a[41] ), .ZN(new_n6571_));
  OAI21_X1   g06378(.A1(new_n6570_), .A2(new_n6571_), .B(new_n6567_), .ZN(new_n6572_));
  NOR2_X1    g06379(.A1(new_n3859_), .A2(new_n4702_), .ZN(new_n6573_));
  NAND2_X1   g06380(.A1(new_n6573_), .A2(new_n1439_), .ZN(new_n6574_));
  NOR3_X1    g06381(.A1(new_n5820_), .A2(new_n3859_), .A3(new_n4901_), .ZN(new_n6575_));
  NOR2_X1    g06382(.A1(new_n5155_), .A2(new_n539_), .ZN(new_n6576_));
  OAI21_X1   g06383(.A1(new_n6575_), .A2(new_n6576_), .B(new_n6574_), .ZN(new_n6577_));
  NAND3_X1   g06384(.A1(new_n6577_), .A2(\a[9] ), .A3(\a[50] ), .ZN(new_n6578_));
  NAND2_X1   g06385(.A1(new_n6577_), .A2(new_n6574_), .ZN(new_n6579_));
  AOI22_X1   g06386(.A1(\a[10] ), .A2(\a[49] ), .B1(\a[15] ), .B2(\a[44] ), .ZN(new_n6580_));
  OAI21_X1   g06387(.A1(new_n6579_), .A2(new_n6580_), .B(new_n6578_), .ZN(new_n6581_));
  XOR2_X1    g06388(.A1(new_n6572_), .A2(new_n6581_), .Z(new_n6582_));
  XOR2_X1    g06389(.A1(new_n6582_), .A2(new_n6560_), .Z(new_n6583_));
  NAND2_X1   g06390(.A1(new_n6444_), .A2(new_n6441_), .ZN(new_n6584_));
  NAND2_X1   g06391(.A1(new_n6445_), .A2(new_n6439_), .ZN(new_n6585_));
  NAND2_X1   g06392(.A1(new_n6585_), .A2(new_n6584_), .ZN(new_n6586_));
  NAND2_X1   g06393(.A1(new_n6586_), .A2(new_n6583_), .ZN(new_n6587_));
  INV_X1     g06394(.I(new_n6587_), .ZN(new_n6588_));
  NOR2_X1    g06395(.A1(new_n6586_), .A2(new_n6583_), .ZN(new_n6589_));
  NOR2_X1    g06396(.A1(new_n6588_), .A2(new_n6589_), .ZN(new_n6590_));
  XOR2_X1    g06397(.A1(new_n6590_), .A2(new_n6557_), .Z(new_n6591_));
  XOR2_X1    g06398(.A1(new_n6532_), .A2(new_n6591_), .Z(new_n6592_));
  NAND2_X1   g06399(.A1(new_n6449_), .A2(new_n6434_), .ZN(new_n6593_));
  OAI21_X1   g06400(.A1(new_n6431_), .A2(new_n6450_), .B(new_n6593_), .ZN(new_n6594_));
  NAND2_X1   g06401(.A1(new_n6327_), .A2(new_n6335_), .ZN(new_n6595_));
  NAND2_X1   g06402(.A1(new_n6336_), .A2(new_n6347_), .ZN(new_n6596_));
  NAND2_X1   g06403(.A1(new_n6596_), .A2(new_n6595_), .ZN(new_n6597_));
  NAND2_X1   g06404(.A1(new_n6387_), .A2(new_n6395_), .ZN(new_n6598_));
  NAND2_X1   g06405(.A1(new_n6396_), .A2(new_n6404_), .ZN(new_n6599_));
  NAND2_X1   g06406(.A1(new_n6599_), .A2(new_n6598_), .ZN(new_n6600_));
  NAND2_X1   g06407(.A1(new_n6363_), .A2(new_n6355_), .ZN(new_n6601_));
  NAND2_X1   g06408(.A1(new_n6364_), .A2(new_n6371_), .ZN(new_n6602_));
  NAND2_X1   g06409(.A1(new_n6602_), .A2(new_n6601_), .ZN(new_n6603_));
  XOR2_X1    g06410(.A1(new_n6603_), .A2(new_n6600_), .Z(new_n6604_));
  NAND2_X1   g06411(.A1(new_n6604_), .A2(new_n6597_), .ZN(new_n6605_));
  OR2_X2     g06412(.A1(new_n6604_), .A2(new_n6597_), .Z(new_n6606_));
  AND2_X2    g06413(.A1(new_n6606_), .A2(new_n6605_), .Z(new_n6607_));
  INV_X1     g06414(.I(new_n6607_), .ZN(new_n6608_));
  NAND2_X1   g06415(.A1(new_n6372_), .A2(new_n6348_), .ZN(new_n6609_));
  OAI21_X1   g06416(.A1(new_n6315_), .A2(new_n6373_), .B(new_n6609_), .ZN(new_n6610_));
  INV_X1     g06417(.I(new_n6610_), .ZN(new_n6611_));
  XOR2_X1    g06418(.A1(new_n6326_), .A2(new_n6403_), .Z(new_n6612_));
  XOR2_X1    g06419(.A1(new_n6612_), .A2(new_n6346_), .Z(new_n6613_));
  XOR2_X1    g06420(.A1(new_n6361_), .A2(new_n6332_), .Z(new_n6614_));
  XOR2_X1    g06421(.A1(new_n6614_), .A2(new_n6352_), .Z(new_n6615_));
  NOR2_X1    g06422(.A1(new_n194_), .A2(new_n6316_), .ZN(new_n6616_));
  NOR2_X1    g06423(.A1(new_n2032_), .A2(new_n6316_), .ZN(new_n6617_));
  INV_X1     g06424(.I(new_n6617_), .ZN(new_n6618_));
  OAI21_X1   g06425(.A1(\a[30] ), .A2(new_n6616_), .B(new_n6618_), .ZN(new_n6619_));
  XNOR2_X1   g06426(.A1(new_n6619_), .A2(new_n6394_), .ZN(new_n6620_));
  XOR2_X1    g06427(.A1(new_n6620_), .A2(new_n6384_), .Z(new_n6621_));
  NAND2_X1   g06428(.A1(new_n6621_), .A2(new_n6615_), .ZN(new_n6622_));
  NAND2_X1   g06429(.A1(new_n6622_), .A2(new_n6615_), .ZN(new_n6623_));
  NAND2_X1   g06430(.A1(new_n6622_), .A2(new_n6621_), .ZN(new_n6624_));
  NAND2_X1   g06431(.A1(new_n6623_), .A2(new_n6624_), .ZN(new_n6625_));
  NAND2_X1   g06432(.A1(new_n6625_), .A2(new_n6613_), .ZN(new_n6626_));
  INV_X1     g06433(.I(new_n6613_), .ZN(new_n6627_));
  NAND3_X1   g06434(.A1(new_n6623_), .A2(new_n6624_), .A3(new_n6627_), .ZN(new_n6628_));
  NAND2_X1   g06435(.A1(new_n6626_), .A2(new_n6628_), .ZN(new_n6629_));
  INV_X1     g06436(.I(new_n6629_), .ZN(new_n6630_));
  NOR2_X1    g06437(.A1(new_n6611_), .A2(new_n6630_), .ZN(new_n6631_));
  INV_X1     g06438(.I(new_n6631_), .ZN(new_n6632_));
  NOR2_X1    g06439(.A1(new_n6610_), .A2(new_n6629_), .ZN(new_n6633_));
  INV_X1     g06440(.I(new_n6633_), .ZN(new_n6634_));
  AOI21_X1   g06441(.A1(new_n6632_), .A2(new_n6634_), .B(new_n6608_), .ZN(new_n6635_));
  NOR3_X1    g06442(.A1(new_n6631_), .A2(new_n6633_), .A3(new_n6607_), .ZN(new_n6636_));
  NOR2_X1    g06443(.A1(new_n6635_), .A2(new_n6636_), .ZN(new_n6637_));
  XOR2_X1    g06444(.A1(new_n6594_), .A2(new_n6637_), .Z(new_n6638_));
  INV_X1     g06445(.I(new_n6638_), .ZN(new_n6639_));
  NAND2_X1   g06446(.A1(new_n6639_), .A2(new_n6592_), .ZN(new_n6640_));
  OR2_X2     g06447(.A1(new_n6639_), .A2(new_n6592_), .Z(new_n6641_));
  NAND2_X1   g06448(.A1(new_n6641_), .A2(new_n6640_), .ZN(new_n6642_));
  OAI21_X1   g06449(.A1(new_n6245_), .A2(new_n6241_), .B(new_n6312_), .ZN(new_n6643_));
  INV_X1     g06450(.I(new_n6313_), .ZN(new_n6644_));
  OAI21_X1   g06451(.A1(new_n6644_), .A2(new_n6424_), .B(new_n6643_), .ZN(new_n6645_));
  NAND2_X1   g06452(.A1(new_n6377_), .A2(new_n6422_), .ZN(new_n6646_));
  NAND2_X1   g06453(.A1(new_n6423_), .A2(new_n6374_), .ZN(new_n6647_));
  NAND2_X1   g06454(.A1(new_n6647_), .A2(new_n6646_), .ZN(new_n6648_));
  NAND2_X1   g06455(.A1(new_n6289_), .A2(new_n6310_), .ZN(new_n6649_));
  NAND2_X1   g06456(.A1(new_n6311_), .A2(new_n6286_), .ZN(new_n6650_));
  NAND2_X1   g06457(.A1(new_n6650_), .A2(new_n6649_), .ZN(new_n6651_));
  NOR2_X1    g06458(.A1(new_n6420_), .A2(new_n6417_), .ZN(new_n6652_));
  NOR2_X1    g06459(.A1(new_n6285_), .A2(new_n6280_), .ZN(new_n6653_));
  NOR2_X1    g06460(.A1(new_n6277_), .A2(new_n6273_), .ZN(new_n6654_));
  NAND2_X1   g06461(.A1(new_n6167_), .A2(new_n6121_), .ZN(new_n6655_));
  INV_X1     g06462(.I(new_n6413_), .ZN(new_n6656_));
  OAI21_X1   g06463(.A1(new_n6656_), .A2(new_n6412_), .B(new_n6655_), .ZN(new_n6657_));
  NOR2_X1    g06464(.A1(new_n6135_), .A2(new_n6143_), .ZN(new_n6658_));
  NOR2_X1    g06465(.A1(new_n6270_), .A2(new_n6658_), .ZN(new_n6659_));
  XNOR2_X1   g06466(.A1(new_n6659_), .A2(new_n6657_), .ZN(new_n6660_));
  XNOR2_X1   g06467(.A1(new_n6660_), .A2(new_n6654_), .ZN(new_n6661_));
  INV_X1     g06468(.I(new_n6661_), .ZN(new_n6662_));
  XOR2_X1    g06469(.A1(new_n6653_), .A2(new_n6662_), .Z(new_n6663_));
  XNOR2_X1   g06470(.A1(new_n6652_), .A2(new_n6663_), .ZN(new_n6664_));
  XOR2_X1    g06471(.A1(new_n6651_), .A2(new_n6664_), .Z(new_n6665_));
  XOR2_X1    g06472(.A1(new_n6648_), .A2(new_n6665_), .Z(new_n6666_));
  NOR2_X1    g06473(.A1(new_n6645_), .A2(new_n6666_), .ZN(new_n6667_));
  NAND2_X1   g06474(.A1(new_n6645_), .A2(new_n6666_), .ZN(new_n6668_));
  INV_X1     g06475(.I(new_n6668_), .ZN(new_n6669_));
  NOR2_X1    g06476(.A1(new_n6669_), .A2(new_n6667_), .ZN(new_n6670_));
  XNOR2_X1   g06477(.A1(new_n6670_), .A2(new_n6642_), .ZN(new_n6671_));
  NOR2_X1    g06478(.A1(new_n6458_), .A2(new_n6454_), .ZN(new_n6672_));
  INV_X1     g06479(.I(new_n6672_), .ZN(new_n6673_));
  NOR2_X1    g06480(.A1(new_n6671_), .A2(new_n6673_), .ZN(new_n6674_));
  NAND2_X1   g06481(.A1(new_n6671_), .A2(new_n6673_), .ZN(new_n6675_));
  INV_X1     g06482(.I(new_n6675_), .ZN(new_n6676_));
  NOR2_X1    g06483(.A1(new_n6676_), .A2(new_n6674_), .ZN(new_n6677_));
  XOR2_X1    g06484(.A1(new_n6479_), .A2(new_n6677_), .Z(\asquared[60] ));
  AOI21_X1   g06485(.A1(new_n6478_), .A2(new_n6462_), .B(new_n6674_), .ZN(new_n6679_));
  NOR2_X1    g06486(.A1(new_n6679_), .A2(new_n6676_), .ZN(new_n6680_));
  NAND2_X1   g06487(.A1(new_n6651_), .A2(new_n6664_), .ZN(new_n6681_));
  NAND2_X1   g06488(.A1(new_n6648_), .A2(new_n6665_), .ZN(new_n6682_));
  NAND2_X1   g06489(.A1(new_n6682_), .A2(new_n6681_), .ZN(new_n6683_));
  NAND2_X1   g06490(.A1(new_n6520_), .A2(new_n6510_), .ZN(new_n6684_));
  NAND2_X1   g06491(.A1(new_n6521_), .A2(new_n6528_), .ZN(new_n6685_));
  NAND2_X1   g06492(.A1(new_n6685_), .A2(new_n6684_), .ZN(new_n6686_));
  NAND2_X1   g06493(.A1(new_n6526_), .A2(new_n6569_), .ZN(new_n6687_));
  NAND2_X1   g06494(.A1(new_n6527_), .A2(new_n6570_), .ZN(new_n6688_));
  AND2_X2    g06495(.A1(new_n6688_), .A2(new_n6687_), .Z(new_n6689_));
  XOR2_X1    g06496(.A1(new_n6689_), .A2(new_n6508_), .Z(new_n6690_));
  NAND2_X1   g06497(.A1(new_n6539_), .A2(new_n6546_), .ZN(new_n6691_));
  INV_X1     g06498(.I(new_n6547_), .ZN(new_n6692_));
  NAND2_X1   g06499(.A1(new_n6692_), .A2(new_n6556_), .ZN(new_n6693_));
  NAND2_X1   g06500(.A1(new_n6693_), .A2(new_n6691_), .ZN(new_n6694_));
  XOR2_X1    g06501(.A1(new_n6694_), .A2(new_n6690_), .Z(new_n6695_));
  XOR2_X1    g06502(.A1(new_n6695_), .A2(new_n6686_), .Z(new_n6696_));
  NAND2_X1   g06503(.A1(new_n6529_), .A2(new_n6502_), .ZN(new_n6697_));
  NAND2_X1   g06504(.A1(new_n6483_), .A2(new_n6530_), .ZN(new_n6698_));
  NAND2_X1   g06505(.A1(new_n6698_), .A2(new_n6697_), .ZN(new_n6699_));
  NAND2_X1   g06506(.A1(new_n6572_), .A2(new_n6581_), .ZN(new_n6700_));
  NAND2_X1   g06507(.A1(new_n6582_), .A2(new_n6560_), .ZN(new_n6701_));
  NAND2_X1   g06508(.A1(new_n6701_), .A2(new_n6700_), .ZN(new_n6702_));
  INV_X1     g06509(.I(new_n6702_), .ZN(new_n6703_));
  XOR2_X1    g06510(.A1(new_n6538_), .A2(new_n6489_), .Z(new_n6704_));
  XOR2_X1    g06511(.A1(new_n6704_), .A2(new_n6545_), .Z(new_n6705_));
  XOR2_X1    g06512(.A1(new_n6554_), .A2(new_n6496_), .Z(new_n6706_));
  XOR2_X1    g06513(.A1(new_n6706_), .A2(new_n6579_), .Z(new_n6707_));
  XNOR2_X1   g06514(.A1(new_n6705_), .A2(new_n6707_), .ZN(new_n6708_));
  XOR2_X1    g06515(.A1(new_n6708_), .A2(new_n6703_), .Z(new_n6709_));
  NAND2_X1   g06516(.A1(new_n6699_), .A2(new_n6709_), .ZN(new_n6710_));
  NAND2_X1   g06517(.A1(new_n6710_), .A2(new_n6699_), .ZN(new_n6711_));
  NAND2_X1   g06518(.A1(new_n6710_), .A2(new_n6709_), .ZN(new_n6712_));
  NAND2_X1   g06519(.A1(new_n6711_), .A2(new_n6712_), .ZN(new_n6713_));
  NAND2_X1   g06520(.A1(new_n6713_), .A2(new_n6696_), .ZN(new_n6714_));
  INV_X1     g06521(.I(new_n6696_), .ZN(new_n6715_));
  NAND3_X1   g06522(.A1(new_n6711_), .A2(new_n6712_), .A3(new_n6715_), .ZN(new_n6716_));
  NAND2_X1   g06523(.A1(new_n6714_), .A2(new_n6716_), .ZN(new_n6717_));
  NOR2_X1    g06524(.A1(new_n6683_), .A2(new_n6717_), .ZN(new_n6718_));
  INV_X1     g06525(.I(new_n6619_), .ZN(new_n6719_));
  NAND2_X1   g06526(.A1(new_n6719_), .A2(new_n6394_), .ZN(new_n6720_));
  NAND2_X1   g06527(.A1(new_n6620_), .A2(new_n6384_), .ZN(new_n6721_));
  NAND2_X1   g06528(.A1(new_n6721_), .A2(new_n6720_), .ZN(new_n6722_));
  INV_X1     g06529(.I(\a[60] ), .ZN(new_n6723_));
  NOR2_X1    g06530(.A1(new_n196_), .A2(new_n6723_), .ZN(new_n6724_));
  XOR2_X1    g06531(.A1(new_n6617_), .A2(new_n6724_), .Z(new_n6725_));
  NOR2_X1    g06532(.A1(new_n194_), .A2(new_n6548_), .ZN(new_n6726_));
  XOR2_X1    g06533(.A1(new_n2976_), .A2(new_n6726_), .Z(new_n6727_));
  XOR2_X1    g06534(.A1(new_n6725_), .A2(new_n6727_), .Z(new_n6728_));
  NAND2_X1   g06535(.A1(new_n2103_), .A2(new_n2636_), .ZN(new_n6729_));
  NOR2_X1    g06536(.A1(new_n1750_), .A2(new_n2752_), .ZN(new_n6730_));
  NAND3_X1   g06537(.A1(new_n6730_), .A2(\a[23] ), .A3(\a[33] ), .ZN(new_n6731_));
  NAND3_X1   g06538(.A1(new_n4860_), .A2(\a[23] ), .A3(\a[37] ), .ZN(new_n6732_));
  INV_X1     g06539(.I(new_n6732_), .ZN(new_n6733_));
  AOI21_X1   g06540(.A1(new_n6729_), .A2(new_n6731_), .B(new_n6733_), .ZN(new_n6734_));
  NAND2_X1   g06541(.A1(\a[27] ), .A2(\a[33] ), .ZN(new_n6735_));
  AOI21_X1   g06542(.A1(\a[23] ), .A2(\a[37] ), .B(new_n4860_), .ZN(new_n6736_));
  NOR2_X1    g06543(.A1(new_n6734_), .A2(new_n6733_), .ZN(new_n6737_));
  INV_X1     g06544(.I(new_n6737_), .ZN(new_n6738_));
  OAI22_X1   g06545(.A1(new_n6738_), .A2(new_n6736_), .B1(new_n6734_), .B2(new_n6735_), .ZN(new_n6739_));
  XOR2_X1    g06546(.A1(new_n6728_), .A2(new_n6739_), .Z(new_n6740_));
  XNOR2_X1   g06547(.A1(new_n6740_), .A2(new_n6722_), .ZN(new_n6741_));
  NAND2_X1   g06548(.A1(new_n760_), .A2(new_n4720_), .ZN(new_n6742_));
  NOR2_X1    g06549(.A1(new_n4178_), .A2(new_n4596_), .ZN(new_n6743_));
  NAND2_X1   g06550(.A1(new_n6743_), .A2(new_n762_), .ZN(new_n6744_));
  AOI22_X1   g06551(.A1(new_n6742_), .A2(new_n6744_), .B1(new_n763_), .B2(new_n4976_), .ZN(new_n6745_));
  AOI22_X1   g06552(.A1(\a[12] ), .A2(\a[48] ), .B1(\a[13] ), .B2(\a[47] ), .ZN(new_n6746_));
  NAND2_X1   g06553(.A1(new_n763_), .A2(new_n4976_), .ZN(new_n6747_));
  NAND3_X1   g06554(.A1(new_n6747_), .A2(new_n6742_), .A3(new_n6744_), .ZN(new_n6748_));
  OAI22_X1   g06555(.A1(new_n6745_), .A2(new_n5889_), .B1(new_n6748_), .B2(new_n6746_), .ZN(new_n6749_));
  NAND4_X1   g06556(.A1(\a[8] ), .A2(\a[18] ), .A3(\a[42] ), .A4(\a[52] ), .ZN(new_n6750_));
  NOR4_X1    g06557(.A1(new_n422_), .A2(new_n884_), .A3(new_n3746_), .A4(new_n5425_), .ZN(new_n6751_));
  NOR2_X1    g06558(.A1(new_n6563_), .A2(new_n415_), .ZN(new_n6752_));
  OAI21_X1   g06559(.A1(new_n6752_), .A2(new_n6751_), .B(new_n6750_), .ZN(new_n6753_));
  NAND3_X1   g06560(.A1(new_n6753_), .A2(\a[7] ), .A3(\a[53] ), .ZN(new_n6754_));
  NAND2_X1   g06561(.A1(new_n6753_), .A2(new_n6750_), .ZN(new_n6755_));
  AOI22_X1   g06562(.A1(\a[8] ), .A2(\a[52] ), .B1(\a[18] ), .B2(\a[42] ), .ZN(new_n6756_));
  OAI21_X1   g06563(.A1(new_n6755_), .A2(new_n6756_), .B(new_n6754_), .ZN(new_n6757_));
  XNOR2_X1   g06564(.A1(new_n6757_), .A2(new_n6749_), .ZN(new_n6758_));
  NAND4_X1   g06565(.A1(\a[5] ), .A2(\a[19] ), .A3(\a[41] ), .A4(\a[55] ), .ZN(new_n6759_));
  NAND2_X1   g06566(.A1(new_n6128_), .A2(new_n746_), .ZN(new_n6760_));
  NOR4_X1    g06567(.A1(new_n367_), .A2(new_n979_), .A3(new_n3327_), .A4(new_n5617_), .ZN(new_n6761_));
  AOI21_X1   g06568(.A1(new_n6760_), .A2(new_n6759_), .B(new_n6761_), .ZN(new_n6762_));
  NAND2_X1   g06569(.A1(\a[5] ), .A2(\a[55] ), .ZN(new_n6763_));
  AOI22_X1   g06570(.A1(\a[6] ), .A2(\a[54] ), .B1(\a[19] ), .B2(\a[41] ), .ZN(new_n6764_));
  OR2_X2     g06571(.A1(new_n6762_), .A2(new_n6761_), .Z(new_n6765_));
  OAI22_X1   g06572(.A1(new_n6765_), .A2(new_n6764_), .B1(new_n6762_), .B2(new_n6763_), .ZN(new_n6766_));
  XOR2_X1    g06573(.A1(new_n6758_), .A2(new_n6766_), .Z(new_n6767_));
  XOR2_X1    g06574(.A1(new_n6741_), .A2(new_n6767_), .Z(new_n6768_));
  INV_X1     g06575(.I(new_n6768_), .ZN(new_n6769_));
  AND3_X2    g06576(.A1(new_n6769_), .A2(new_n6622_), .A3(new_n6626_), .Z(new_n6770_));
  AOI21_X1   g06577(.A1(new_n6622_), .A2(new_n6626_), .B(new_n6769_), .ZN(new_n6771_));
  NOR2_X1    g06578(.A1(new_n6770_), .A2(new_n6771_), .ZN(new_n6772_));
  NOR2_X1    g06579(.A1(new_n6653_), .A2(new_n6662_), .ZN(new_n6773_));
  INV_X1     g06580(.I(new_n6663_), .ZN(new_n6774_));
  NOR2_X1    g06581(.A1(new_n6774_), .A2(new_n6652_), .ZN(new_n6775_));
  NOR2_X1    g06582(.A1(new_n6775_), .A2(new_n6773_), .ZN(new_n6776_));
  NOR2_X1    g06583(.A1(new_n4030_), .A2(new_n4702_), .ZN(new_n6777_));
  INV_X1     g06584(.I(new_n6777_), .ZN(new_n6778_));
  NOR3_X1    g06585(.A1(new_n6778_), .A2(new_n513_), .A3(new_n717_), .ZN(new_n6779_));
  NAND3_X1   g06586(.A1(new_n1439_), .A2(\a[45] ), .A3(\a[50] ), .ZN(new_n6780_));
  NAND2_X1   g06587(.A1(new_n747_), .A2(new_n5154_), .ZN(new_n6781_));
  AOI21_X1   g06588(.A1(new_n6781_), .A2(new_n6780_), .B(new_n6779_), .ZN(new_n6782_));
  NAND2_X1   g06589(.A1(\a[10] ), .A2(\a[50] ), .ZN(new_n6783_));
  AOI22_X1   g06590(.A1(\a[11] ), .A2(\a[49] ), .B1(\a[15] ), .B2(\a[45] ), .ZN(new_n6784_));
  OR2_X2     g06591(.A1(new_n6782_), .A2(new_n6779_), .Z(new_n6785_));
  OAI22_X1   g06592(.A1(new_n6785_), .A2(new_n6784_), .B1(new_n6782_), .B2(new_n6783_), .ZN(new_n6786_));
  NOR3_X1    g06593(.A1(new_n798_), .A2(new_n3859_), .A3(new_n5135_), .ZN(new_n6787_));
  INV_X1     g06594(.I(new_n6787_), .ZN(new_n6788_));
  INV_X1     g06595(.I(new_n5276_), .ZN(new_n6789_));
  INV_X1     g06596(.I(new_n6113_), .ZN(new_n6790_));
  OAI22_X1   g06597(.A1(new_n1428_), .A2(new_n4343_), .B1(new_n6789_), .B2(new_n6790_), .ZN(new_n6791_));
  NAND2_X1   g06598(.A1(new_n6791_), .A2(new_n6788_), .ZN(new_n6792_));
  NAND3_X1   g06599(.A1(new_n6792_), .A2(\a[17] ), .A3(\a[43] ), .ZN(new_n6793_));
  AOI22_X1   g06600(.A1(\a[9] ), .A2(\a[51] ), .B1(\a[16] ), .B2(\a[44] ), .ZN(new_n6794_));
  NAND2_X1   g06601(.A1(new_n6792_), .A2(new_n6788_), .ZN(new_n6795_));
  OAI21_X1   g06602(.A1(new_n6794_), .A2(new_n6795_), .B(new_n6793_), .ZN(new_n6796_));
  XOR2_X1    g06603(.A1(new_n6796_), .A2(new_n6519_), .Z(new_n6797_));
  XOR2_X1    g06604(.A1(new_n6797_), .A2(new_n6786_), .Z(new_n6798_));
  OAI21_X1   g06605(.A1(new_n6658_), .A2(new_n6270_), .B(new_n6657_), .ZN(new_n6799_));
  INV_X1     g06606(.I(new_n6660_), .ZN(new_n6800_));
  OAI21_X1   g06607(.A1(new_n6800_), .A2(new_n6654_), .B(new_n6799_), .ZN(new_n6801_));
  NAND2_X1   g06608(.A1(new_n6494_), .A2(new_n761_), .ZN(new_n6802_));
  NOR2_X1    g06609(.A1(new_n6298_), .A2(new_n6316_), .ZN(new_n6803_));
  INV_X1     g06610(.I(new_n6803_), .ZN(new_n6804_));
  OAI22_X1   g06611(.A1(new_n246_), .A2(new_n6804_), .B1(new_n6318_), .B2(new_n251_), .ZN(new_n6805_));
  NAND2_X1   g06612(.A1(new_n6805_), .A2(new_n6802_), .ZN(new_n6806_));
  NAND3_X1   g06613(.A1(new_n6806_), .A2(\a[2] ), .A3(\a[58] ), .ZN(new_n6807_));
  AOI22_X1   g06614(.A1(\a[3] ), .A2(\a[57] ), .B1(\a[4] ), .B2(\a[56] ), .ZN(new_n6808_));
  NAND2_X1   g06615(.A1(new_n6806_), .A2(new_n6802_), .ZN(new_n6809_));
  OAI21_X1   g06616(.A1(new_n6808_), .A2(new_n6809_), .B(new_n6807_), .ZN(new_n6810_));
  NOR2_X1    g06617(.A1(new_n1456_), .A2(new_n4210_), .ZN(new_n6811_));
  NOR2_X1    g06618(.A1(new_n2647_), .A2(new_n3223_), .ZN(new_n6812_));
  NOR2_X1    g06619(.A1(new_n1382_), .A2(new_n3551_), .ZN(new_n6813_));
  NOR2_X1    g06620(.A1(new_n6812_), .A2(new_n6813_), .ZN(new_n6814_));
  NOR2_X1    g06621(.A1(new_n6814_), .A2(new_n6811_), .ZN(new_n6815_));
  NAND2_X1   g06622(.A1(\a[20] ), .A2(\a[40] ), .ZN(new_n6816_));
  AOI22_X1   g06623(.A1(\a[21] ), .A2(\a[39] ), .B1(\a[22] ), .B2(\a[38] ), .ZN(new_n6817_));
  NOR2_X1    g06624(.A1(new_n6815_), .A2(new_n6811_), .ZN(new_n6818_));
  INV_X1     g06625(.I(new_n6818_), .ZN(new_n6819_));
  OAI22_X1   g06626(.A1(new_n6819_), .A2(new_n6817_), .B1(new_n6815_), .B2(new_n6816_), .ZN(new_n6820_));
  XOR2_X1    g06627(.A1(new_n6820_), .A2(new_n6810_), .Z(new_n6821_));
  NOR2_X1    g06628(.A1(new_n2177_), .A2(new_n2746_), .ZN(new_n6822_));
  AOI22_X1   g06629(.A1(new_n1778_), .A2(new_n3232_), .B1(new_n2080_), .B2(new_n3822_), .ZN(new_n6823_));
  NOR2_X1    g06630(.A1(new_n6822_), .A2(new_n6823_), .ZN(new_n6824_));
  NAND2_X1   g06631(.A1(\a[24] ), .A2(\a[36] ), .ZN(new_n6825_));
  AOI22_X1   g06632(.A1(\a[25] ), .A2(\a[35] ), .B1(\a[26] ), .B2(\a[34] ), .ZN(new_n6826_));
  NOR2_X1    g06633(.A1(new_n6824_), .A2(new_n6822_), .ZN(new_n6827_));
  INV_X1     g06634(.I(new_n6827_), .ZN(new_n6828_));
  OAI22_X1   g06635(.A1(new_n6828_), .A2(new_n6826_), .B1(new_n6824_), .B2(new_n6825_), .ZN(new_n6829_));
  XOR2_X1    g06636(.A1(new_n6821_), .A2(new_n6829_), .Z(new_n6830_));
  XOR2_X1    g06637(.A1(new_n6801_), .A2(new_n6830_), .Z(new_n6831_));
  XNOR2_X1   g06638(.A1(new_n6831_), .A2(new_n6798_), .ZN(new_n6832_));
  XNOR2_X1   g06639(.A1(new_n6776_), .A2(new_n6832_), .ZN(new_n6833_));
  XOR2_X1    g06640(.A1(new_n6833_), .A2(new_n6772_), .Z(new_n6834_));
  INV_X1     g06641(.I(new_n6834_), .ZN(new_n6835_));
  NAND2_X1   g06642(.A1(new_n6683_), .A2(new_n6717_), .ZN(new_n6836_));
  INV_X1     g06643(.I(new_n6836_), .ZN(new_n6837_));
  OAI21_X1   g06644(.A1(new_n6837_), .A2(new_n6718_), .B(new_n6835_), .ZN(new_n6838_));
  NAND2_X1   g06645(.A1(new_n6836_), .A2(new_n6834_), .ZN(new_n6839_));
  OAI21_X1   g06646(.A1(new_n6718_), .A2(new_n6839_), .B(new_n6838_), .ZN(new_n6840_));
  NAND2_X1   g06647(.A1(new_n6594_), .A2(new_n6637_), .ZN(new_n6841_));
  NAND2_X1   g06648(.A1(new_n6641_), .A2(new_n6841_), .ZN(new_n6842_));
  NOR2_X1    g06649(.A1(new_n6482_), .A2(new_n6531_), .ZN(new_n6843_));
  INV_X1     g06650(.I(new_n6532_), .ZN(new_n6844_));
  NOR2_X1    g06651(.A1(new_n6844_), .A2(new_n6591_), .ZN(new_n6845_));
  NOR2_X1    g06652(.A1(new_n6845_), .A2(new_n6843_), .ZN(new_n6846_));
  INV_X1     g06653(.I(new_n6635_), .ZN(new_n6847_));
  OAI21_X1   g06654(.A1(new_n6611_), .A2(new_n6629_), .B(new_n6847_), .ZN(new_n6848_));
  INV_X1     g06655(.I(new_n6590_), .ZN(new_n6849_));
  NOR2_X1    g06656(.A1(new_n6849_), .A2(new_n6557_), .ZN(new_n6850_));
  NOR2_X1    g06657(.A1(new_n6850_), .A2(new_n6588_), .ZN(new_n6851_));
  INV_X1     g06658(.I(new_n6501_), .ZN(new_n6852_));
  NAND2_X1   g06659(.A1(new_n6852_), .A2(new_n6491_), .ZN(new_n6853_));
  OAI21_X1   g06660(.A1(new_n6369_), .A2(new_n6500_), .B(new_n6853_), .ZN(new_n6854_));
  NAND2_X1   g06661(.A1(new_n6326_), .A2(new_n6403_), .ZN(new_n6855_));
  NAND2_X1   g06662(.A1(new_n6612_), .A2(new_n6346_), .ZN(new_n6856_));
  NAND2_X1   g06663(.A1(new_n6856_), .A2(new_n6855_), .ZN(new_n6857_));
  NAND2_X1   g06664(.A1(new_n6614_), .A2(new_n6352_), .ZN(new_n6858_));
  OAI21_X1   g06665(.A1(new_n6332_), .A2(new_n6361_), .B(new_n6858_), .ZN(new_n6859_));
  XOR2_X1    g06666(.A1(new_n6857_), .A2(new_n6859_), .Z(new_n6860_));
  XOR2_X1    g06667(.A1(new_n6854_), .A2(new_n6860_), .Z(new_n6861_));
  NAND2_X1   g06668(.A1(new_n6603_), .A2(new_n6600_), .ZN(new_n6862_));
  NAND2_X1   g06669(.A1(new_n6605_), .A2(new_n6862_), .ZN(new_n6863_));
  XOR2_X1    g06670(.A1(new_n6863_), .A2(new_n6861_), .Z(new_n6864_));
  INV_X1     g06671(.I(new_n6864_), .ZN(new_n6865_));
  XOR2_X1    g06672(.A1(new_n6851_), .A2(new_n6865_), .Z(new_n6866_));
  XOR2_X1    g06673(.A1(new_n6848_), .A2(new_n6866_), .Z(new_n6867_));
  XNOR2_X1   g06674(.A1(new_n6867_), .A2(new_n6846_), .ZN(new_n6868_));
  NOR2_X1    g06675(.A1(new_n6842_), .A2(new_n6868_), .ZN(new_n6869_));
  NAND2_X1   g06676(.A1(new_n6842_), .A2(new_n6868_), .ZN(new_n6870_));
  INV_X1     g06677(.I(new_n6870_), .ZN(new_n6871_));
  NOR2_X1    g06678(.A1(new_n6871_), .A2(new_n6869_), .ZN(new_n6872_));
  XNOR2_X1   g06679(.A1(new_n6872_), .A2(new_n6840_), .ZN(new_n6873_));
  INV_X1     g06680(.I(new_n6873_), .ZN(new_n6874_));
  INV_X1     g06681(.I(new_n6670_), .ZN(new_n6875_));
  NOR2_X1    g06682(.A1(new_n6875_), .A2(new_n6642_), .ZN(new_n6876_));
  NOR2_X1    g06683(.A1(new_n6876_), .A2(new_n6669_), .ZN(new_n6877_));
  NOR2_X1    g06684(.A1(new_n6877_), .A2(new_n6874_), .ZN(new_n6878_));
  INV_X1     g06685(.I(new_n6878_), .ZN(new_n6879_));
  NAND2_X1   g06686(.A1(new_n6877_), .A2(new_n6874_), .ZN(new_n6880_));
  NAND2_X1   g06687(.A1(new_n6879_), .A2(new_n6880_), .ZN(new_n6881_));
  XOR2_X1    g06688(.A1(new_n6680_), .A2(new_n6881_), .Z(\asquared[61] ));
  OAI21_X1   g06689(.A1(new_n6679_), .A2(new_n6676_), .B(new_n6880_), .ZN(new_n6883_));
  NAND2_X1   g06690(.A1(new_n6883_), .A2(new_n6879_), .ZN(new_n6884_));
  INV_X1     g06691(.I(new_n6872_), .ZN(new_n6885_));
  NOR2_X1    g06692(.A1(new_n6885_), .A2(new_n6840_), .ZN(new_n6886_));
  NOR2_X1    g06693(.A1(new_n6886_), .A2(new_n6871_), .ZN(new_n6887_));
  INV_X1     g06694(.I(new_n6887_), .ZN(new_n6888_));
  NAND2_X1   g06695(.A1(new_n6714_), .A2(new_n6710_), .ZN(new_n6889_));
  NAND2_X1   g06696(.A1(new_n6863_), .A2(new_n6861_), .ZN(new_n6890_));
  OAI21_X1   g06697(.A1(new_n6865_), .A2(new_n6851_), .B(new_n6890_), .ZN(new_n6891_));
  NOR2_X1    g06698(.A1(new_n253_), .A2(new_n6548_), .ZN(new_n6892_));
  INV_X1     g06699(.I(new_n6892_), .ZN(new_n6893_));
  NOR3_X1    g06700(.A1(new_n6893_), .A2(new_n197_), .A3(new_n5856_), .ZN(new_n6894_));
  INV_X1     g06701(.I(new_n6894_), .ZN(new_n6895_));
  NAND4_X1   g06702(.A1(\a[0] ), .A2(\a[5] ), .A3(\a[56] ), .A4(\a[61] ), .ZN(new_n6896_));
  INV_X1     g06703(.I(\a[61] ), .ZN(new_n6897_));
  NOR2_X1    g06704(.A1(new_n6548_), .A2(new_n6897_), .ZN(new_n6898_));
  INV_X1     g06705(.I(new_n6898_), .ZN(new_n6899_));
  OAI21_X1   g06706(.A1(new_n6899_), .A2(new_n412_), .B(new_n6896_), .ZN(new_n6900_));
  NAND2_X1   g06707(.A1(new_n6895_), .A2(new_n6900_), .ZN(new_n6901_));
  NAND3_X1   g06708(.A1(new_n6901_), .A2(\a[0] ), .A3(\a[61] ), .ZN(new_n6902_));
  AOI22_X1   g06709(.A1(\a[2] ), .A2(\a[59] ), .B1(\a[5] ), .B2(\a[56] ), .ZN(new_n6903_));
  NOR2_X1    g06710(.A1(new_n6894_), .A2(new_n6900_), .ZN(new_n6904_));
  INV_X1     g06711(.I(new_n6904_), .ZN(new_n6905_));
  OAI21_X1   g06712(.A1(new_n6903_), .A2(new_n6905_), .B(new_n6902_), .ZN(new_n6906_));
  AOI22_X1   g06713(.A1(\a[20] ), .A2(\a[41] ), .B1(\a[21] ), .B2(\a[40] ), .ZN(new_n6907_));
  INV_X1     g06714(.I(new_n6907_), .ZN(new_n6908_));
  NOR2_X1    g06715(.A1(new_n1382_), .A2(new_n5377_), .ZN(new_n6909_));
  NOR2_X1    g06716(.A1(new_n367_), .A2(new_n5680_), .ZN(new_n6910_));
  AOI21_X1   g06717(.A1(new_n6908_), .A2(new_n6910_), .B(new_n6909_), .ZN(new_n6911_));
  NAND2_X1   g06718(.A1(new_n6911_), .A2(new_n6908_), .ZN(new_n6912_));
  OAI21_X1   g06719(.A1(new_n6909_), .A2(new_n6907_), .B(new_n6910_), .ZN(new_n6913_));
  NAND2_X1   g06720(.A1(new_n6912_), .A2(new_n6913_), .ZN(new_n6914_));
  XNOR2_X1   g06721(.A1(new_n6906_), .A2(new_n6914_), .ZN(new_n6915_));
  NOR2_X1    g06722(.A1(new_n2626_), .A2(new_n3116_), .ZN(new_n6916_));
  NAND2_X1   g06723(.A1(new_n4351_), .A2(new_n6916_), .ZN(new_n6917_));
  NAND2_X1   g06724(.A1(new_n1879_), .A2(new_n4545_), .ZN(new_n6918_));
  AOI22_X1   g06725(.A1(new_n6917_), .A2(new_n6918_), .B1(new_n1778_), .B2(new_n3037_), .ZN(new_n6919_));
  NAND2_X1   g06726(.A1(\a[22] ), .A2(\a[39] ), .ZN(new_n6920_));
  AOI22_X1   g06727(.A1(\a[24] ), .A2(\a[37] ), .B1(\a[25] ), .B2(\a[36] ), .ZN(new_n6921_));
  NAND2_X1   g06728(.A1(new_n1778_), .A2(new_n3037_), .ZN(new_n6922_));
  NAND3_X1   g06729(.A1(new_n6922_), .A2(new_n6917_), .A3(new_n6918_), .ZN(new_n6923_));
  OAI22_X1   g06730(.A1(new_n6919_), .A2(new_n6920_), .B1(new_n6923_), .B2(new_n6921_), .ZN(new_n6924_));
  XOR2_X1    g06731(.A1(new_n6915_), .A2(new_n6924_), .Z(new_n6925_));
  INV_X1     g06732(.I(new_n6925_), .ZN(new_n6926_));
  NAND2_X1   g06733(.A1(new_n6857_), .A2(new_n6859_), .ZN(new_n6927_));
  NAND2_X1   g06734(.A1(new_n6854_), .A2(new_n6860_), .ZN(new_n6928_));
  NAND2_X1   g06735(.A1(new_n6928_), .A2(new_n6927_), .ZN(new_n6929_));
  NOR2_X1    g06736(.A1(new_n4178_), .A2(new_n5135_), .ZN(new_n6930_));
  INV_X1     g06737(.I(new_n6930_), .ZN(new_n6931_));
  NOR2_X1    g06738(.A1(new_n6931_), .A2(new_n710_), .ZN(new_n6932_));
  NAND3_X1   g06739(.A1(new_n4848_), .A2(\a[10] ), .A3(\a[51] ), .ZN(new_n6933_));
  NAND2_X1   g06740(.A1(new_n4429_), .A2(new_n1288_), .ZN(new_n6934_));
  AOI21_X1   g06741(.A1(new_n6934_), .A2(new_n6933_), .B(new_n6932_), .ZN(new_n6935_));
  AOI22_X1   g06742(.A1(\a[10] ), .A2(\a[51] ), .B1(\a[15] ), .B2(\a[46] ), .ZN(new_n6936_));
  OR2_X2     g06743(.A1(new_n6935_), .A2(new_n6932_), .Z(new_n6937_));
  OAI22_X1   g06744(.A1(new_n6937_), .A2(new_n6936_), .B1(new_n4849_), .B2(new_n6935_), .ZN(new_n6938_));
  NOR2_X1    g06745(.A1(new_n4979_), .A2(new_n623_), .ZN(new_n6939_));
  NOR2_X1    g06746(.A1(new_n5155_), .A2(new_n619_), .ZN(new_n6940_));
  NOR2_X1    g06747(.A1(new_n759_), .A2(new_n4901_), .ZN(new_n6941_));
  INV_X1     g06748(.I(new_n6941_), .ZN(new_n6942_));
  NOR3_X1    g06749(.A1(new_n6942_), .A2(new_n513_), .A3(new_n4312_), .ZN(new_n6943_));
  NOR2_X1    g06750(.A1(new_n6943_), .A2(new_n6940_), .ZN(new_n6944_));
  NOR2_X1    g06751(.A1(new_n6944_), .A2(new_n6939_), .ZN(new_n6945_));
  NAND2_X1   g06752(.A1(\a[11] ), .A2(\a[50] ), .ZN(new_n6946_));
  AOI22_X1   g06753(.A1(\a[12] ), .A2(\a[49] ), .B1(\a[14] ), .B2(\a[47] ), .ZN(new_n6947_));
  NOR2_X1    g06754(.A1(new_n6945_), .A2(new_n6939_), .ZN(new_n6948_));
  INV_X1     g06755(.I(new_n6948_), .ZN(new_n6949_));
  OAI22_X1   g06756(.A1(new_n6949_), .A2(new_n6947_), .B1(new_n6945_), .B2(new_n6946_), .ZN(new_n6950_));
  XOR2_X1    g06757(.A1(new_n6950_), .A2(new_n6938_), .Z(new_n6951_));
  AOI21_X1   g06758(.A1(\a[29] ), .A2(\a[32] ), .B(new_n2437_), .ZN(new_n6952_));
  NOR2_X1    g06759(.A1(new_n597_), .A2(new_n4596_), .ZN(new_n6953_));
  INV_X1     g06760(.I(new_n6953_), .ZN(new_n6954_));
  NOR2_X1    g06761(.A1(new_n2255_), .A2(new_n3833_), .ZN(new_n6955_));
  NOR3_X1    g06762(.A1(new_n6955_), .A2(new_n6952_), .A3(new_n6954_), .ZN(new_n6956_));
  NOR2_X1    g06763(.A1(new_n6956_), .A2(new_n6955_), .ZN(new_n6957_));
  INV_X1     g06764(.I(new_n6957_), .ZN(new_n6958_));
  OAI22_X1   g06765(.A1(new_n6958_), .A2(new_n6952_), .B1(new_n6954_), .B2(new_n6956_), .ZN(new_n6959_));
  XNOR2_X1   g06766(.A1(new_n6951_), .A2(new_n6959_), .ZN(new_n6960_));
  INV_X1     g06767(.I(new_n6960_), .ZN(new_n6961_));
  XOR2_X1    g06768(.A1(new_n6929_), .A2(new_n6961_), .Z(new_n6962_));
  XOR2_X1    g06769(.A1(new_n6962_), .A2(new_n6926_), .Z(new_n6963_));
  XOR2_X1    g06770(.A1(new_n6891_), .A2(new_n6963_), .Z(new_n6964_));
  XOR2_X1    g06771(.A1(new_n6964_), .A2(new_n6889_), .Z(new_n6965_));
  NAND2_X1   g06772(.A1(new_n6848_), .A2(new_n6866_), .ZN(new_n6966_));
  INV_X1     g06773(.I(new_n6867_), .ZN(new_n6967_));
  OAI21_X1   g06774(.A1(new_n6967_), .A2(new_n6846_), .B(new_n6966_), .ZN(new_n6968_));
  NOR2_X1    g06775(.A1(new_n6741_), .A2(new_n6767_), .ZN(new_n6969_));
  NOR2_X1    g06776(.A1(new_n6771_), .A2(new_n6969_), .ZN(new_n6970_));
  NAND2_X1   g06777(.A1(new_n6728_), .A2(new_n6739_), .ZN(new_n6971_));
  NAND2_X1   g06778(.A1(new_n6740_), .A2(new_n6722_), .ZN(new_n6972_));
  NAND2_X1   g06779(.A1(new_n6972_), .A2(new_n6971_), .ZN(new_n6973_));
  NAND2_X1   g06780(.A1(new_n6617_), .A2(new_n6724_), .ZN(new_n6974_));
  NAND2_X1   g06781(.A1(new_n6725_), .A2(new_n6727_), .ZN(new_n6975_));
  NAND2_X1   g06782(.A1(new_n6975_), .A2(new_n6974_), .ZN(new_n6976_));
  XOR2_X1    g06783(.A1(new_n6795_), .A2(new_n6755_), .Z(new_n6977_));
  XOR2_X1    g06784(.A1(new_n6977_), .A2(new_n6976_), .Z(new_n6978_));
  NAND2_X1   g06785(.A1(new_n6757_), .A2(new_n6749_), .ZN(new_n6979_));
  INV_X1     g06786(.I(new_n6758_), .ZN(new_n6980_));
  NAND2_X1   g06787(.A1(new_n6980_), .A2(new_n6766_), .ZN(new_n6981_));
  NAND2_X1   g06788(.A1(new_n6981_), .A2(new_n6979_), .ZN(new_n6982_));
  XOR2_X1    g06789(.A1(new_n6982_), .A2(new_n6978_), .Z(new_n6983_));
  XOR2_X1    g06790(.A1(new_n6983_), .A2(new_n6973_), .Z(new_n6984_));
  NAND2_X1   g06791(.A1(new_n6820_), .A2(new_n6810_), .ZN(new_n6985_));
  NAND2_X1   g06792(.A1(new_n6821_), .A2(new_n6829_), .ZN(new_n6986_));
  NAND2_X1   g06793(.A1(new_n6986_), .A2(new_n6985_), .ZN(new_n6987_));
  XOR2_X1    g06794(.A1(new_n6809_), .A2(new_n6765_), .Z(new_n6988_));
  XOR2_X1    g06795(.A1(new_n6988_), .A2(new_n6785_), .Z(new_n6989_));
  NOR2_X1    g06796(.A1(new_n6738_), .A2(new_n6828_), .ZN(new_n6990_));
  NOR2_X1    g06797(.A1(new_n6737_), .A2(new_n6827_), .ZN(new_n6991_));
  NOR2_X1    g06798(.A1(new_n6990_), .A2(new_n6991_), .ZN(new_n6992_));
  NAND2_X1   g06799(.A1(new_n6992_), .A2(new_n6819_), .ZN(new_n6993_));
  INV_X1     g06800(.I(new_n6993_), .ZN(new_n6994_));
  NOR2_X1    g06801(.A1(new_n6992_), .A2(new_n6819_), .ZN(new_n6995_));
  NOR2_X1    g06802(.A1(new_n6994_), .A2(new_n6995_), .ZN(new_n6996_));
  XOR2_X1    g06803(.A1(new_n6996_), .A2(new_n6989_), .Z(new_n6997_));
  XOR2_X1    g06804(.A1(new_n6997_), .A2(new_n6987_), .Z(new_n6998_));
  NOR2_X1    g06805(.A1(new_n6984_), .A2(new_n6998_), .ZN(new_n6999_));
  NAND2_X1   g06806(.A1(new_n6984_), .A2(new_n6998_), .ZN(new_n7000_));
  INV_X1     g06807(.I(new_n7000_), .ZN(new_n7001_));
  NOR3_X1    g06808(.A1(new_n7001_), .A2(new_n6970_), .A3(new_n6999_), .ZN(new_n7002_));
  OAI21_X1   g06809(.A1(new_n6970_), .A2(new_n6999_), .B(new_n7000_), .ZN(new_n7003_));
  OAI22_X1   g06810(.A1(new_n7002_), .A2(new_n6970_), .B1(new_n7003_), .B2(new_n6999_), .ZN(new_n7004_));
  XOR2_X1    g06811(.A1(new_n6968_), .A2(new_n7004_), .Z(new_n7005_));
  XOR2_X1    g06812(.A1(new_n7005_), .A2(new_n6965_), .Z(new_n7006_));
  NAND3_X1   g06813(.A1(new_n6683_), .A2(new_n6714_), .A3(new_n6716_), .ZN(new_n7007_));
  NAND2_X1   g06814(.A1(new_n6838_), .A2(new_n7007_), .ZN(new_n7008_));
  NOR2_X1    g06815(.A1(new_n6776_), .A2(new_n6832_), .ZN(new_n7009_));
  INV_X1     g06816(.I(new_n6833_), .ZN(new_n7010_));
  AOI21_X1   g06817(.A1(new_n7010_), .A2(new_n6772_), .B(new_n7009_), .ZN(new_n7011_));
  NOR2_X1    g06818(.A1(new_n3859_), .A2(new_n5175_), .ZN(new_n7012_));
  INV_X1     g06819(.I(new_n7012_), .ZN(new_n7013_));
  NOR2_X1    g06820(.A1(new_n1543_), .A2(new_n7013_), .ZN(new_n7014_));
  INV_X1     g06821(.I(new_n7014_), .ZN(new_n7015_));
  OAI22_X1   g06822(.A1(new_n1275_), .A2(new_n4343_), .B1(new_n6789_), .B2(new_n6562_), .ZN(new_n7016_));
  NAND2_X1   g06823(.A1(new_n7015_), .A2(new_n7016_), .ZN(new_n7017_));
  NAND3_X1   g06824(.A1(new_n7017_), .A2(\a[18] ), .A3(\a[43] ), .ZN(new_n7018_));
  AOI22_X1   g06825(.A1(\a[9] ), .A2(\a[52] ), .B1(\a[17] ), .B2(\a[44] ), .ZN(new_n7019_));
  NAND2_X1   g06826(.A1(new_n7017_), .A2(new_n7015_), .ZN(new_n7020_));
  OAI21_X1   g06827(.A1(new_n7019_), .A2(new_n7020_), .B(new_n7018_), .ZN(new_n7021_));
  AOI22_X1   g06828(.A1(\a[7] ), .A2(\a[54] ), .B1(\a[8] ), .B2(\a[53] ), .ZN(new_n7022_));
  INV_X1     g06829(.I(new_n7022_), .ZN(new_n7023_));
  NOR2_X1    g06830(.A1(new_n6127_), .A2(new_n415_), .ZN(new_n7024_));
  NOR2_X1    g06831(.A1(new_n979_), .A2(new_n3746_), .ZN(new_n7025_));
  AOI21_X1   g06832(.A1(new_n7023_), .A2(new_n7025_), .B(new_n7024_), .ZN(new_n7026_));
  INV_X1     g06833(.I(new_n7026_), .ZN(new_n7027_));
  OAI21_X1   g06834(.A1(new_n7024_), .A2(new_n7022_), .B(new_n7025_), .ZN(new_n7028_));
  OAI21_X1   g06835(.A1(new_n7027_), .A2(new_n7022_), .B(new_n7028_), .ZN(new_n7029_));
  XOR2_X1    g06836(.A1(new_n7021_), .A2(new_n7029_), .Z(new_n7030_));
  OAI22_X1   g06837(.A1(new_n1972_), .A2(new_n2746_), .B1(new_n3341_), .B2(new_n2526_), .ZN(new_n7031_));
  OAI21_X1   g06838(.A1(new_n2189_), .A2(new_n3932_), .B(new_n7031_), .ZN(new_n7032_));
  NAND3_X1   g06839(.A1(new_n7032_), .A2(\a[26] ), .A3(\a[35] ), .ZN(new_n7033_));
  AOI22_X1   g06840(.A1(\a[27] ), .A2(\a[34] ), .B1(\a[28] ), .B2(\a[33] ), .ZN(new_n7034_));
  NOR2_X1    g06841(.A1(new_n2189_), .A2(new_n3932_), .ZN(new_n7035_));
  NOR2_X1    g06842(.A1(new_n7031_), .A2(new_n7035_), .ZN(new_n7036_));
  INV_X1     g06843(.I(new_n7036_), .ZN(new_n7037_));
  OAI21_X1   g06844(.A1(new_n7034_), .A2(new_n7037_), .B(new_n7033_), .ZN(new_n7038_));
  XOR2_X1    g06845(.A1(new_n7030_), .A2(new_n7038_), .Z(new_n7039_));
  NAND2_X1   g06846(.A1(new_n6705_), .A2(new_n6707_), .ZN(new_n7040_));
  OAI21_X1   g06847(.A1(new_n6708_), .A2(new_n6703_), .B(new_n7040_), .ZN(new_n7041_));
  XOR2_X1    g06848(.A1(new_n7041_), .A2(new_n7039_), .Z(new_n7042_));
  NAND2_X1   g06849(.A1(new_n6694_), .A2(new_n6690_), .ZN(new_n7043_));
  NAND2_X1   g06850(.A1(new_n6695_), .A2(new_n6686_), .ZN(new_n7044_));
  NAND2_X1   g06851(.A1(new_n7044_), .A2(new_n7043_), .ZN(new_n7045_));
  XNOR2_X1   g06852(.A1(new_n7045_), .A2(new_n7042_), .ZN(new_n7046_));
  NAND2_X1   g06853(.A1(new_n6801_), .A2(new_n6830_), .ZN(new_n7047_));
  NAND2_X1   g06854(.A1(new_n6831_), .A2(new_n6798_), .ZN(new_n7048_));
  NAND2_X1   g06855(.A1(new_n7048_), .A2(new_n7047_), .ZN(new_n7049_));
  NAND2_X1   g06856(.A1(new_n6689_), .A2(new_n6508_), .ZN(new_n7050_));
  NAND2_X1   g06857(.A1(new_n7050_), .A2(new_n6688_), .ZN(new_n7051_));
  AOI22_X1   g06858(.A1(\a[3] ), .A2(\a[58] ), .B1(\a[4] ), .B2(\a[57] ), .ZN(new_n7052_));
  NOR2_X1    g06859(.A1(new_n1299_), .A2(new_n2914_), .ZN(new_n7053_));
  INV_X1     g06860(.I(new_n7053_), .ZN(new_n7054_));
  NOR2_X1    g06861(.A1(new_n6804_), .A2(new_n370_), .ZN(new_n7055_));
  NOR3_X1    g06862(.A1(new_n7055_), .A2(new_n7052_), .A3(new_n7054_), .ZN(new_n7056_));
  NOR2_X1    g06863(.A1(new_n7056_), .A2(new_n7055_), .ZN(new_n7057_));
  INV_X1     g06864(.I(new_n7057_), .ZN(new_n7058_));
  OAI22_X1   g06865(.A1(new_n7058_), .A2(new_n7052_), .B1(new_n7054_), .B2(new_n7056_), .ZN(new_n7059_));
  XOR2_X1    g06866(.A1(new_n7051_), .A2(new_n7059_), .Z(new_n7060_));
  NAND2_X1   g06867(.A1(new_n6554_), .A2(new_n6496_), .ZN(new_n7061_));
  NAND2_X1   g06868(.A1(new_n6706_), .A2(new_n6579_), .ZN(new_n7062_));
  NAND2_X1   g06869(.A1(new_n7062_), .A2(new_n7061_), .ZN(new_n7063_));
  XNOR2_X1   g06870(.A1(new_n7060_), .A2(new_n7063_), .ZN(new_n7064_));
  NAND2_X1   g06871(.A1(new_n6797_), .A2(new_n6786_), .ZN(new_n7065_));
  NAND2_X1   g06872(.A1(new_n6796_), .A2(new_n6519_), .ZN(new_n7066_));
  NAND2_X1   g06873(.A1(new_n7065_), .A2(new_n7066_), .ZN(new_n7067_));
  NAND2_X1   g06874(.A1(new_n6538_), .A2(new_n6489_), .ZN(new_n7068_));
  NAND2_X1   g06875(.A1(new_n6704_), .A2(new_n6545_), .ZN(new_n7069_));
  NAND2_X1   g06876(.A1(new_n7069_), .A2(new_n7068_), .ZN(new_n7070_));
  INV_X1     g06877(.I(new_n6726_), .ZN(new_n7071_));
  NOR2_X1    g06878(.A1(new_n5625_), .A2(new_n7071_), .ZN(new_n7072_));
  NOR2_X1    g06879(.A1(new_n194_), .A2(new_n6723_), .ZN(new_n7073_));
  INV_X1     g06880(.I(new_n7073_), .ZN(new_n7074_));
  NAND2_X1   g06881(.A1(new_n7074_), .A2(new_n2051_), .ZN(new_n7075_));
  NOR2_X1    g06882(.A1(new_n7074_), .A2(new_n2051_), .ZN(new_n7076_));
  INV_X1     g06883(.I(new_n7076_), .ZN(new_n7077_));
  AND2_X2    g06884(.A1(new_n7077_), .A2(new_n7075_), .Z(new_n7078_));
  XOR2_X1    g06885(.A1(new_n7078_), .A2(new_n7072_), .Z(new_n7079_));
  XOR2_X1    g06886(.A1(new_n7079_), .A2(new_n6748_), .Z(new_n7080_));
  XOR2_X1    g06887(.A1(new_n7080_), .A2(new_n7070_), .Z(new_n7081_));
  XOR2_X1    g06888(.A1(new_n7081_), .A2(new_n7067_), .Z(new_n7082_));
  NOR2_X1    g06889(.A1(new_n7064_), .A2(new_n7082_), .ZN(new_n7083_));
  AND2_X2    g06890(.A1(new_n7064_), .A2(new_n7082_), .Z(new_n7084_));
  OAI21_X1   g06891(.A1(new_n7083_), .A2(new_n7084_), .B(new_n7049_), .ZN(new_n7085_));
  INV_X1     g06892(.I(new_n7085_), .ZN(new_n7086_));
  NOR3_X1    g06893(.A1(new_n7049_), .A2(new_n7083_), .A3(new_n7084_), .ZN(new_n7087_));
  NOR2_X1    g06894(.A1(new_n7086_), .A2(new_n7087_), .ZN(new_n7088_));
  XOR2_X1    g06895(.A1(new_n7088_), .A2(new_n7046_), .Z(new_n7089_));
  XOR2_X1    g06896(.A1(new_n7011_), .A2(new_n7089_), .Z(new_n7090_));
  NAND2_X1   g06897(.A1(new_n7008_), .A2(new_n7090_), .ZN(new_n7091_));
  NAND2_X1   g06898(.A1(new_n7091_), .A2(new_n7008_), .ZN(new_n7092_));
  NAND2_X1   g06899(.A1(new_n7091_), .A2(new_n7090_), .ZN(new_n7093_));
  NAND2_X1   g06900(.A1(new_n7092_), .A2(new_n7093_), .ZN(new_n7094_));
  NAND2_X1   g06901(.A1(new_n7094_), .A2(new_n7006_), .ZN(new_n7095_));
  INV_X1     g06902(.I(new_n7006_), .ZN(new_n7096_));
  NAND3_X1   g06903(.A1(new_n7096_), .A2(new_n7092_), .A3(new_n7093_), .ZN(new_n7097_));
  NAND2_X1   g06904(.A1(new_n7095_), .A2(new_n7097_), .ZN(new_n7098_));
  INV_X1     g06905(.I(new_n7098_), .ZN(new_n7099_));
  NOR2_X1    g06906(.A1(new_n6888_), .A2(new_n7099_), .ZN(new_n7100_));
  NOR2_X1    g06907(.A1(new_n6887_), .A2(new_n7098_), .ZN(new_n7101_));
  NOR2_X1    g06908(.A1(new_n7100_), .A2(new_n7101_), .ZN(new_n7102_));
  XOR2_X1    g06909(.A1(new_n6884_), .A2(new_n7102_), .Z(\asquared[62] ));
  AOI21_X1   g06910(.A1(new_n6883_), .A2(new_n6879_), .B(new_n7100_), .ZN(new_n7104_));
  NOR2_X1    g06911(.A1(new_n7104_), .A2(new_n7101_), .ZN(new_n7105_));
  NAND2_X1   g06912(.A1(new_n7095_), .A2(new_n7091_), .ZN(new_n7106_));
  INV_X1     g06913(.I(new_n7082_), .ZN(new_n7107_));
  OAI21_X1   g06914(.A1(new_n7064_), .A2(new_n7107_), .B(new_n7085_), .ZN(new_n7108_));
  AOI22_X1   g06915(.A1(\a[8] ), .A2(\a[54] ), .B1(\a[18] ), .B2(\a[44] ), .ZN(new_n7109_));
  NAND4_X1   g06916(.A1(\a[8] ), .A2(\a[18] ), .A3(\a[44] ), .A4(\a[54] ), .ZN(new_n7110_));
  NOR4_X1    g06917(.A1(new_n355_), .A2(new_n979_), .A3(new_n3666_), .A4(new_n5617_), .ZN(new_n7111_));
  NOR2_X1    g06918(.A1(new_n4343_), .A2(new_n1092_), .ZN(new_n7112_));
  OAI21_X1   g06919(.A1(new_n7112_), .A2(new_n7111_), .B(new_n7110_), .ZN(new_n7113_));
  NAND2_X1   g06920(.A1(new_n7113_), .A2(new_n7110_), .ZN(new_n7114_));
  NAND3_X1   g06921(.A1(new_n7113_), .A2(\a[19] ), .A3(\a[43] ), .ZN(new_n7115_));
  OAI21_X1   g06922(.A1(new_n7109_), .A2(new_n7114_), .B(new_n7115_), .ZN(new_n7116_));
  NAND2_X1   g06923(.A1(new_n2105_), .A2(new_n3577_), .ZN(new_n7117_));
  OAI22_X1   g06924(.A1(new_n1816_), .A2(new_n2526_), .B1(new_n2189_), .B2(new_n2746_), .ZN(new_n7118_));
  NAND2_X1   g06925(.A1(new_n7118_), .A2(new_n7117_), .ZN(new_n7119_));
  NAND3_X1   g06926(.A1(new_n7119_), .A2(\a[27] ), .A3(\a[35] ), .ZN(new_n7120_));
  AOI22_X1   g06927(.A1(\a[28] ), .A2(\a[34] ), .B1(\a[29] ), .B2(\a[33] ), .ZN(new_n7121_));
  NAND2_X1   g06928(.A1(new_n7119_), .A2(new_n7117_), .ZN(new_n7122_));
  OAI21_X1   g06929(.A1(new_n7121_), .A2(new_n7122_), .B(new_n7120_), .ZN(new_n7123_));
  XNOR2_X1   g06930(.A1(new_n7123_), .A2(new_n7116_), .ZN(new_n7124_));
  OAI22_X1   g06931(.A1(new_n2385_), .A2(new_n3551_), .B1(new_n1880_), .B2(new_n3223_), .ZN(new_n7125_));
  OAI21_X1   g06932(.A1(new_n1529_), .A2(new_n4210_), .B(new_n7125_), .ZN(new_n7126_));
  NAND3_X1   g06933(.A1(new_n7126_), .A2(\a[22] ), .A3(\a[40] ), .ZN(new_n7127_));
  AOI22_X1   g06934(.A1(\a[23] ), .A2(\a[39] ), .B1(\a[24] ), .B2(\a[38] ), .ZN(new_n7128_));
  NOR2_X1    g06935(.A1(new_n1529_), .A2(new_n4210_), .ZN(new_n7129_));
  NOR2_X1    g06936(.A1(new_n7125_), .A2(new_n7129_), .ZN(new_n7130_));
  INV_X1     g06937(.I(new_n7130_), .ZN(new_n7131_));
  OAI21_X1   g06938(.A1(new_n7128_), .A2(new_n7131_), .B(new_n7127_), .ZN(new_n7132_));
  XOR2_X1    g06939(.A1(new_n7124_), .A2(new_n7132_), .Z(new_n7133_));
  AOI22_X1   g06940(.A1(\a[25] ), .A2(\a[37] ), .B1(\a[26] ), .B2(\a[36] ), .ZN(new_n7134_));
  INV_X1     g06941(.I(new_n7134_), .ZN(new_n7135_));
  NOR2_X1    g06942(.A1(new_n2177_), .A2(new_n3038_), .ZN(new_n7136_));
  NOR2_X1    g06943(.A1(new_n1220_), .A2(new_n3327_), .ZN(new_n7137_));
  AOI21_X1   g06944(.A1(new_n7135_), .A2(new_n7137_), .B(new_n7136_), .ZN(new_n7138_));
  NAND2_X1   g06945(.A1(new_n7138_), .A2(new_n7135_), .ZN(new_n7139_));
  OAI21_X1   g06946(.A1(new_n7136_), .A2(new_n7134_), .B(new_n7137_), .ZN(new_n7140_));
  NAND2_X1   g06947(.A1(new_n7139_), .A2(new_n7140_), .ZN(new_n7141_));
  AOI22_X1   g06948(.A1(\a[0] ), .A2(\a[62] ), .B1(\a[2] ), .B2(\a[60] ), .ZN(new_n7142_));
  INV_X1     g06949(.I(new_n7142_), .ZN(new_n7143_));
  INV_X1     g06950(.I(\a[62] ), .ZN(new_n7144_));
  NOR2_X1    g06951(.A1(new_n6723_), .A2(new_n7144_), .ZN(new_n7145_));
  INV_X1     g06952(.I(new_n7145_), .ZN(new_n7146_));
  NOR2_X1    g06953(.A1(new_n7146_), .A2(new_n412_), .ZN(new_n7147_));
  AOI21_X1   g06954(.A1(new_n7076_), .A2(new_n7143_), .B(new_n7147_), .ZN(new_n7148_));
  NAND2_X1   g06955(.A1(new_n7148_), .A2(new_n7143_), .ZN(new_n7149_));
  OAI21_X1   g06956(.A1(new_n7142_), .A2(new_n7147_), .B(new_n7076_), .ZN(new_n7150_));
  NAND2_X1   g06957(.A1(new_n7149_), .A2(new_n7150_), .ZN(new_n7151_));
  XOR2_X1    g06958(.A1(new_n7141_), .A2(new_n7151_), .Z(new_n7152_));
  NOR4_X1    g06959(.A1(new_n417_), .A2(new_n1023_), .A3(new_n4030_), .A4(new_n5175_), .ZN(new_n7153_));
  NAND3_X1   g06960(.A1(new_n5543_), .A2(\a[17] ), .A3(\a[53] ), .ZN(new_n7154_));
  NAND2_X1   g06961(.A1(new_n5862_), .A2(new_n540_), .ZN(new_n7155_));
  AOI21_X1   g06962(.A1(new_n7154_), .A2(new_n7155_), .B(new_n7153_), .ZN(new_n7156_));
  NAND2_X1   g06963(.A1(\a[9] ), .A2(\a[53] ), .ZN(new_n7157_));
  OR2_X2     g06964(.A1(new_n7156_), .A2(new_n7153_), .Z(new_n7158_));
  AOI22_X1   g06965(.A1(\a[10] ), .A2(\a[52] ), .B1(\a[17] ), .B2(\a[45] ), .ZN(new_n7159_));
  OAI22_X1   g06966(.A1(new_n7158_), .A2(new_n7159_), .B1(new_n7156_), .B2(new_n7157_), .ZN(new_n7160_));
  XNOR2_X1   g06967(.A1(new_n7152_), .A2(new_n7160_), .ZN(new_n7161_));
  NOR2_X1    g06968(.A1(new_n4312_), .A2(new_n5135_), .ZN(new_n7162_));
  NAND2_X1   g06969(.A1(new_n832_), .A2(new_n7162_), .ZN(new_n7163_));
  INV_X1     g06970(.I(new_n7163_), .ZN(new_n7164_));
  NOR2_X1    g06971(.A1(new_n1734_), .A2(new_n6931_), .ZN(new_n7165_));
  NOR2_X1    g06972(.A1(new_n4721_), .A2(new_n893_), .ZN(new_n7166_));
  NOR2_X1    g06973(.A1(new_n7165_), .A2(new_n7166_), .ZN(new_n7167_));
  NOR2_X1    g06974(.A1(new_n7167_), .A2(new_n7164_), .ZN(new_n7168_));
  NAND2_X1   g06975(.A1(\a[16] ), .A2(\a[46] ), .ZN(new_n7169_));
  AOI22_X1   g06976(.A1(\a[11] ), .A2(\a[51] ), .B1(\a[15] ), .B2(\a[47] ), .ZN(new_n7170_));
  NOR2_X1    g06977(.A1(new_n7168_), .A2(new_n7164_), .ZN(new_n7171_));
  INV_X1     g06978(.I(new_n7171_), .ZN(new_n7172_));
  OAI22_X1   g06979(.A1(new_n7172_), .A2(new_n7170_), .B1(new_n7168_), .B2(new_n7169_), .ZN(new_n7173_));
  NAND2_X1   g06980(.A1(new_n760_), .A2(new_n4980_), .ZN(new_n7174_));
  OAI22_X1   g06981(.A1(new_n1265_), .A2(new_n5155_), .B1(new_n4903_), .B2(new_n623_), .ZN(new_n7175_));
  NAND2_X1   g06982(.A1(new_n7175_), .A2(new_n7174_), .ZN(new_n7176_));
  NAND3_X1   g06983(.A1(new_n7176_), .A2(\a[12] ), .A3(\a[50] ), .ZN(new_n7177_));
  AOI22_X1   g06984(.A1(\a[13] ), .A2(\a[49] ), .B1(\a[14] ), .B2(\a[48] ), .ZN(new_n7178_));
  NAND2_X1   g06985(.A1(new_n7176_), .A2(new_n7174_), .ZN(new_n7179_));
  OAI21_X1   g06986(.A1(new_n7178_), .A2(new_n7179_), .B(new_n7177_), .ZN(new_n7180_));
  XOR2_X1    g06987(.A1(new_n7173_), .A2(new_n7180_), .Z(new_n7181_));
  AOI22_X1   g06988(.A1(\a[6] ), .A2(\a[56] ), .B1(\a[7] ), .B2(\a[55] ), .ZN(new_n7182_));
  NAND2_X1   g06989(.A1(\a[20] ), .A2(\a[42] ), .ZN(new_n7183_));
  NOR2_X1    g06990(.A1(new_n5680_), .A2(new_n5856_), .ZN(new_n7184_));
  INV_X1     g06991(.I(new_n7184_), .ZN(new_n7185_));
  NOR2_X1    g06992(.A1(new_n7185_), .A2(new_n374_), .ZN(new_n7186_));
  NOR3_X1    g06993(.A1(new_n7186_), .A2(new_n7182_), .A3(new_n7183_), .ZN(new_n7187_));
  NOR2_X1    g06994(.A1(new_n7187_), .A2(new_n7186_), .ZN(new_n7188_));
  INV_X1     g06995(.I(new_n7188_), .ZN(new_n7189_));
  OAI22_X1   g06996(.A1(new_n7189_), .A2(new_n7182_), .B1(new_n7183_), .B2(new_n7187_), .ZN(new_n7190_));
  XOR2_X1    g06997(.A1(new_n7181_), .A2(new_n7190_), .Z(new_n7191_));
  XOR2_X1    g06998(.A1(new_n7191_), .A2(new_n7161_), .Z(new_n7192_));
  XOR2_X1    g06999(.A1(new_n7192_), .A2(new_n7133_), .Z(new_n7193_));
  XOR2_X1    g07000(.A1(new_n7108_), .A2(new_n7193_), .Z(new_n7194_));
  XNOR2_X1   g07001(.A1(new_n7194_), .A2(new_n7003_), .ZN(new_n7195_));
  INV_X1     g07002(.I(new_n7046_), .ZN(new_n7196_));
  NOR2_X1    g07003(.A1(new_n7011_), .A2(new_n7089_), .ZN(new_n7197_));
  AOI21_X1   g07004(.A1(new_n7196_), .A2(new_n7088_), .B(new_n7197_), .ZN(new_n7198_));
  NAND2_X1   g07005(.A1(new_n7051_), .A2(new_n7059_), .ZN(new_n7199_));
  NAND2_X1   g07006(.A1(new_n7060_), .A2(new_n7063_), .ZN(new_n7200_));
  NAND2_X1   g07007(.A1(new_n7200_), .A2(new_n7199_), .ZN(new_n7201_));
  XOR2_X1    g07008(.A1(new_n6937_), .A2(new_n7020_), .Z(new_n7202_));
  NOR2_X1    g07009(.A1(new_n6298_), .A2(new_n6548_), .ZN(new_n7203_));
  INV_X1     g07010(.I(new_n7203_), .ZN(new_n7204_));
  NOR2_X1    g07011(.A1(new_n6316_), .A2(new_n6548_), .ZN(new_n7205_));
  INV_X1     g07012(.I(new_n7205_), .ZN(new_n7206_));
  OAI22_X1   g07013(.A1(new_n370_), .A2(new_n7206_), .B1(new_n7204_), .B2(new_n318_), .ZN(new_n7207_));
  OAI21_X1   g07014(.A1(new_n242_), .A2(new_n6804_), .B(new_n7207_), .ZN(new_n7208_));
  NAND3_X1   g07015(.A1(new_n7208_), .A2(\a[3] ), .A3(\a[59] ), .ZN(new_n7209_));
  AOI22_X1   g07016(.A1(\a[4] ), .A2(\a[58] ), .B1(\a[5] ), .B2(\a[57] ), .ZN(new_n7210_));
  NOR2_X1    g07017(.A1(new_n6804_), .A2(new_n242_), .ZN(new_n7211_));
  NOR2_X1    g07018(.A1(new_n7207_), .A2(new_n7211_), .ZN(new_n7212_));
  INV_X1     g07019(.I(new_n7212_), .ZN(new_n7213_));
  OAI21_X1   g07020(.A1(new_n7210_), .A2(new_n7213_), .B(new_n7209_), .ZN(new_n7214_));
  XNOR2_X1   g07021(.A1(new_n7202_), .A2(new_n7214_), .ZN(new_n7215_));
  NAND2_X1   g07022(.A1(new_n7021_), .A2(new_n7029_), .ZN(new_n7216_));
  NAND2_X1   g07023(.A1(new_n7030_), .A2(new_n7038_), .ZN(new_n7217_));
  NAND2_X1   g07024(.A1(new_n7217_), .A2(new_n7216_), .ZN(new_n7218_));
  XNOR2_X1   g07025(.A1(new_n7218_), .A2(new_n7215_), .ZN(new_n7219_));
  XOR2_X1    g07026(.A1(new_n7201_), .A2(new_n7219_), .Z(new_n7220_));
  INV_X1     g07027(.I(new_n7220_), .ZN(new_n7221_));
  NAND2_X1   g07028(.A1(new_n6929_), .A2(new_n6961_), .ZN(new_n7222_));
  NAND2_X1   g07029(.A1(new_n6962_), .A2(new_n6926_), .ZN(new_n7223_));
  NAND2_X1   g07030(.A1(new_n7223_), .A2(new_n7222_), .ZN(new_n7224_));
  NAND2_X1   g07031(.A1(new_n6795_), .A2(new_n6755_), .ZN(new_n7225_));
  NAND2_X1   g07032(.A1(new_n6977_), .A2(new_n6976_), .ZN(new_n7226_));
  NAND2_X1   g07033(.A1(new_n7226_), .A2(new_n7225_), .ZN(new_n7227_));
  INV_X1     g07034(.I(new_n7072_), .ZN(new_n7228_));
  INV_X1     g07035(.I(new_n7078_), .ZN(new_n7229_));
  NAND2_X1   g07036(.A1(new_n7079_), .A2(new_n6748_), .ZN(new_n7230_));
  OAI21_X1   g07037(.A1(new_n7228_), .A2(new_n7229_), .B(new_n7230_), .ZN(new_n7231_));
  XOR2_X1    g07038(.A1(new_n7231_), .A2(new_n7227_), .Z(new_n7232_));
  OAI21_X1   g07039(.A1(new_n6991_), .A2(new_n6994_), .B(new_n7232_), .ZN(new_n7233_));
  NOR2_X1    g07040(.A1(new_n6994_), .A2(new_n6991_), .ZN(new_n7234_));
  INV_X1     g07041(.I(new_n7232_), .ZN(new_n7235_));
  NAND2_X1   g07042(.A1(new_n7235_), .A2(new_n7234_), .ZN(new_n7236_));
  AND2_X2    g07043(.A1(new_n7236_), .A2(new_n7233_), .Z(new_n7237_));
  INV_X1     g07044(.I(new_n7237_), .ZN(new_n7238_));
  NAND2_X1   g07045(.A1(new_n7224_), .A2(new_n7238_), .ZN(new_n7239_));
  NOR2_X1    g07046(.A1(new_n7224_), .A2(new_n7238_), .ZN(new_n7240_));
  INV_X1     g07047(.I(new_n7240_), .ZN(new_n7241_));
  AOI21_X1   g07048(.A1(new_n7241_), .A2(new_n7239_), .B(new_n7221_), .ZN(new_n7242_));
  INV_X1     g07049(.I(new_n7242_), .ZN(new_n7243_));
  NAND3_X1   g07050(.A1(new_n7241_), .A2(new_n7221_), .A3(new_n7239_), .ZN(new_n7244_));
  NAND2_X1   g07051(.A1(new_n7243_), .A2(new_n7244_), .ZN(new_n7245_));
  XOR2_X1    g07052(.A1(new_n7198_), .A2(new_n7245_), .Z(new_n7246_));
  XNOR2_X1   g07053(.A1(new_n7246_), .A2(new_n7195_), .ZN(new_n7247_));
  NAND2_X1   g07054(.A1(new_n7041_), .A2(new_n7039_), .ZN(new_n7248_));
  NAND2_X1   g07055(.A1(new_n7045_), .A2(new_n7042_), .ZN(new_n7249_));
  NAND2_X1   g07056(.A1(new_n7249_), .A2(new_n7248_), .ZN(new_n7250_));
  NAND2_X1   g07057(.A1(new_n6950_), .A2(new_n6938_), .ZN(new_n7251_));
  NAND2_X1   g07058(.A1(new_n6951_), .A2(new_n6959_), .ZN(new_n7252_));
  NAND2_X1   g07059(.A1(new_n7252_), .A2(new_n7251_), .ZN(new_n7253_));
  NAND2_X1   g07060(.A1(new_n6809_), .A2(new_n6765_), .ZN(new_n7254_));
  NAND2_X1   g07061(.A1(new_n6988_), .A2(new_n6785_), .ZN(new_n7255_));
  NAND2_X1   g07062(.A1(new_n7255_), .A2(new_n7254_), .ZN(new_n7256_));
  NAND2_X1   g07063(.A1(new_n6906_), .A2(new_n6914_), .ZN(new_n7257_));
  INV_X1     g07064(.I(new_n6915_), .ZN(new_n7258_));
  NAND2_X1   g07065(.A1(new_n7258_), .A2(new_n6924_), .ZN(new_n7259_));
  NAND2_X1   g07066(.A1(new_n7259_), .A2(new_n7257_), .ZN(new_n7260_));
  XOR2_X1    g07067(.A1(new_n7260_), .A2(new_n7256_), .Z(new_n7261_));
  XOR2_X1    g07068(.A1(new_n7261_), .A2(new_n7253_), .Z(new_n7262_));
  XOR2_X1    g07069(.A1(new_n6911_), .A2(new_n6904_), .Z(new_n7263_));
  INV_X1     g07070(.I(new_n7263_), .ZN(new_n7264_));
  NAND2_X1   g07071(.A1(new_n7264_), .A2(new_n7026_), .ZN(new_n7265_));
  NOR2_X1    g07072(.A1(new_n7264_), .A2(new_n7026_), .ZN(new_n7266_));
  INV_X1     g07073(.I(new_n7266_), .ZN(new_n7267_));
  AND2_X2    g07074(.A1(new_n7267_), .A2(new_n7265_), .Z(new_n7268_));
  XOR2_X1    g07075(.A1(new_n7057_), .A2(new_n7036_), .Z(new_n7269_));
  XOR2_X1    g07076(.A1(new_n7269_), .A2(new_n6923_), .Z(new_n7270_));
  NAND2_X1   g07077(.A1(\a[1] ), .A2(\a[61] ), .ZN(new_n7271_));
  XNOR2_X1   g07078(.A1(new_n2201_), .A2(new_n7271_), .ZN(new_n7272_));
  NOR2_X1    g07079(.A1(new_n6958_), .A2(new_n7272_), .ZN(new_n7273_));
  INV_X1     g07080(.I(new_n7272_), .ZN(new_n7274_));
  NOR2_X1    g07081(.A1(new_n6957_), .A2(new_n7274_), .ZN(new_n7275_));
  NOR2_X1    g07082(.A1(new_n7273_), .A2(new_n7275_), .ZN(new_n7276_));
  INV_X1     g07083(.I(new_n7276_), .ZN(new_n7277_));
  NAND2_X1   g07084(.A1(new_n7277_), .A2(new_n6948_), .ZN(new_n7278_));
  NOR2_X1    g07085(.A1(new_n7277_), .A2(new_n6948_), .ZN(new_n7279_));
  INV_X1     g07086(.I(new_n7279_), .ZN(new_n7280_));
  AND2_X2    g07087(.A1(new_n7280_), .A2(new_n7278_), .Z(new_n7281_));
  XNOR2_X1   g07088(.A1(new_n7281_), .A2(new_n7270_), .ZN(new_n7282_));
  XOR2_X1    g07089(.A1(new_n7282_), .A2(new_n7268_), .Z(new_n7283_));
  XOR2_X1    g07090(.A1(new_n7262_), .A2(new_n7283_), .Z(new_n7284_));
  XOR2_X1    g07091(.A1(new_n7284_), .A2(new_n7250_), .Z(new_n7285_));
  NAND2_X1   g07092(.A1(new_n6891_), .A2(new_n6963_), .ZN(new_n7286_));
  NAND2_X1   g07093(.A1(new_n6964_), .A2(new_n6889_), .ZN(new_n7287_));
  NAND2_X1   g07094(.A1(new_n7287_), .A2(new_n7286_), .ZN(new_n7288_));
  NAND2_X1   g07095(.A1(new_n6982_), .A2(new_n6978_), .ZN(new_n7289_));
  NAND2_X1   g07096(.A1(new_n6983_), .A2(new_n6973_), .ZN(new_n7290_));
  NAND2_X1   g07097(.A1(new_n7290_), .A2(new_n7289_), .ZN(new_n7291_));
  NAND2_X1   g07098(.A1(new_n6996_), .A2(new_n6989_), .ZN(new_n7292_));
  NAND2_X1   g07099(.A1(new_n6997_), .A2(new_n6987_), .ZN(new_n7293_));
  NAND2_X1   g07100(.A1(new_n7293_), .A2(new_n7292_), .ZN(new_n7294_));
  NAND2_X1   g07101(.A1(new_n7080_), .A2(new_n7070_), .ZN(new_n7295_));
  NAND2_X1   g07102(.A1(new_n7081_), .A2(new_n7067_), .ZN(new_n7296_));
  NAND2_X1   g07103(.A1(new_n7296_), .A2(new_n7295_), .ZN(new_n7297_));
  XOR2_X1    g07104(.A1(new_n7294_), .A2(new_n7297_), .Z(new_n7298_));
  XOR2_X1    g07105(.A1(new_n7298_), .A2(new_n7291_), .Z(new_n7299_));
  XNOR2_X1   g07106(.A1(new_n7288_), .A2(new_n7299_), .ZN(new_n7300_));
  XOR2_X1    g07107(.A1(new_n7300_), .A2(new_n7285_), .Z(new_n7301_));
  NAND2_X1   g07108(.A1(new_n6968_), .A2(new_n7004_), .ZN(new_n7302_));
  NAND2_X1   g07109(.A1(new_n7005_), .A2(new_n6965_), .ZN(new_n7303_));
  NAND2_X1   g07110(.A1(new_n7303_), .A2(new_n7302_), .ZN(new_n7304_));
  NAND2_X1   g07111(.A1(new_n7304_), .A2(new_n7301_), .ZN(new_n7305_));
  NAND2_X1   g07112(.A1(new_n7305_), .A2(new_n7301_), .ZN(new_n7306_));
  NAND2_X1   g07113(.A1(new_n7305_), .A2(new_n7304_), .ZN(new_n7307_));
  NAND2_X1   g07114(.A1(new_n7307_), .A2(new_n7306_), .ZN(new_n7308_));
  AOI21_X1   g07115(.A1(new_n7305_), .A2(new_n7304_), .B(new_n7247_), .ZN(new_n7309_));
  AOI22_X1   g07116(.A1(new_n7308_), .A2(new_n7247_), .B1(new_n7306_), .B2(new_n7309_), .ZN(new_n7310_));
  NAND2_X1   g07117(.A1(new_n7310_), .A2(new_n7106_), .ZN(new_n7311_));
  NOR2_X1    g07118(.A1(new_n7310_), .A2(new_n7106_), .ZN(new_n7312_));
  INV_X1     g07119(.I(new_n7312_), .ZN(new_n7313_));
  NAND2_X1   g07120(.A1(new_n7313_), .A2(new_n7311_), .ZN(new_n7314_));
  INV_X1     g07121(.I(new_n7101_), .ZN(new_n7315_));
  INV_X1     g07122(.I(new_n6674_), .ZN(new_n7316_));
  OAI21_X1   g07123(.A1(new_n6476_), .A2(new_n6461_), .B(new_n7316_), .ZN(new_n7317_));
  INV_X1     g07124(.I(new_n6880_), .ZN(new_n7318_));
  AOI21_X1   g07125(.A1(new_n7317_), .A2(new_n6675_), .B(new_n7318_), .ZN(new_n7319_));
  INV_X1     g07126(.I(new_n7100_), .ZN(new_n7320_));
  OAI21_X1   g07127(.A1(new_n7319_), .A2(new_n6878_), .B(new_n7320_), .ZN(new_n7321_));
  AOI21_X1   g07128(.A1(new_n7321_), .A2(new_n7315_), .B(new_n7312_), .ZN(new_n7322_));
  AOI22_X1   g07129(.A1(new_n7322_), .A2(new_n7311_), .B1(new_n7105_), .B2(new_n7314_), .ZN(\asquared[63] ));
  OAI21_X1   g07130(.A1(new_n7104_), .A2(new_n7101_), .B(new_n7313_), .ZN(new_n7324_));
  NAND2_X1   g07131(.A1(new_n7324_), .A2(new_n7311_), .ZN(new_n7325_));
  NAND2_X1   g07132(.A1(new_n7308_), .A2(new_n7247_), .ZN(new_n7326_));
  NAND2_X1   g07133(.A1(new_n7326_), .A2(new_n7305_), .ZN(new_n7327_));
  NAND2_X1   g07134(.A1(new_n7288_), .A2(new_n7299_), .ZN(new_n7328_));
  OAI21_X1   g07135(.A1(new_n7300_), .A2(new_n7285_), .B(new_n7328_), .ZN(new_n7329_));
  NAND2_X1   g07136(.A1(new_n7294_), .A2(new_n7297_), .ZN(new_n7330_));
  NAND2_X1   g07137(.A1(new_n7298_), .A2(new_n7291_), .ZN(new_n7331_));
  NAND2_X1   g07138(.A1(new_n7331_), .A2(new_n7330_), .ZN(new_n7332_));
  NAND2_X1   g07139(.A1(new_n7231_), .A2(new_n7227_), .ZN(new_n7333_));
  NAND2_X1   g07140(.A1(new_n7233_), .A2(new_n7333_), .ZN(new_n7334_));
  NAND2_X1   g07141(.A1(new_n7141_), .A2(new_n7151_), .ZN(new_n7335_));
  NAND2_X1   g07142(.A1(new_n7152_), .A2(new_n7160_), .ZN(new_n7336_));
  NAND2_X1   g07143(.A1(new_n7336_), .A2(new_n7335_), .ZN(new_n7337_));
  XOR2_X1    g07144(.A1(new_n7334_), .A2(new_n7337_), .Z(new_n7338_));
  NAND3_X1   g07145(.A1(new_n2201_), .A2(\a[1] ), .A3(\a[61] ), .ZN(new_n7339_));
  NAND2_X1   g07146(.A1(\a[0] ), .A2(\a[63] ), .ZN(new_n7340_));
  XNOR2_X1   g07147(.A1(new_n7339_), .A2(new_n7340_), .ZN(new_n7341_));
  INV_X1     g07148(.I(new_n7341_), .ZN(new_n7342_));
  NOR2_X1    g07149(.A1(new_n2368_), .A2(new_n7144_), .ZN(new_n7343_));
  NOR2_X1    g07150(.A1(new_n7343_), .A2(new_n194_), .ZN(new_n7344_));
  INV_X1     g07151(.I(new_n7344_), .ZN(new_n7345_));
  OAI22_X1   g07152(.A1(new_n7345_), .A2(new_n7144_), .B1(new_n2200_), .B2(new_n7343_), .ZN(new_n7346_));
  XOR2_X1    g07153(.A1(new_n7346_), .A2(new_n7342_), .Z(new_n7347_));
  NAND2_X1   g07154(.A1(new_n2176_), .A2(new_n3803_), .ZN(new_n7348_));
  OAI22_X1   g07155(.A1(new_n1779_), .A2(new_n4210_), .B1(new_n2081_), .B2(new_n4739_), .ZN(new_n7349_));
  NAND2_X1   g07156(.A1(new_n7349_), .A2(new_n7348_), .ZN(new_n7350_));
  NAND3_X1   g07157(.A1(new_n7350_), .A2(\a[24] ), .A3(\a[39] ), .ZN(new_n7351_));
  AOI22_X1   g07158(.A1(\a[25] ), .A2(\a[38] ), .B1(\a[26] ), .B2(\a[37] ), .ZN(new_n7352_));
  NAND2_X1   g07159(.A1(new_n7350_), .A2(new_n7348_), .ZN(new_n7353_));
  OAI21_X1   g07160(.A1(new_n7352_), .A2(new_n7353_), .B(new_n7351_), .ZN(new_n7354_));
  NAND2_X1   g07161(.A1(new_n2105_), .A2(new_n2745_), .ZN(new_n7355_));
  OAI22_X1   g07162(.A1(new_n1816_), .A2(new_n5564_), .B1(new_n2189_), .B2(new_n3405_), .ZN(new_n7356_));
  NAND2_X1   g07163(.A1(new_n7356_), .A2(new_n7355_), .ZN(new_n7357_));
  NAND3_X1   g07164(.A1(new_n7357_), .A2(\a[27] ), .A3(\a[36] ), .ZN(new_n7358_));
  AOI22_X1   g07165(.A1(\a[28] ), .A2(\a[35] ), .B1(\a[29] ), .B2(\a[34] ), .ZN(new_n7359_));
  NAND2_X1   g07166(.A1(new_n7357_), .A2(new_n7355_), .ZN(new_n7360_));
  OAI21_X1   g07167(.A1(new_n7359_), .A2(new_n7360_), .B(new_n7358_), .ZN(new_n7361_));
  XOR2_X1    g07168(.A1(new_n7354_), .A2(new_n7361_), .Z(new_n7362_));
  XOR2_X1    g07169(.A1(new_n7362_), .A2(new_n7347_), .Z(new_n7363_));
  XNOR2_X1   g07170(.A1(new_n7338_), .A2(new_n7363_), .ZN(new_n7364_));
  NAND2_X1   g07171(.A1(new_n7173_), .A2(new_n7180_), .ZN(new_n7365_));
  NAND2_X1   g07172(.A1(new_n7181_), .A2(new_n7190_), .ZN(new_n7366_));
  NAND2_X1   g07173(.A1(new_n7366_), .A2(new_n7365_), .ZN(new_n7367_));
  XOR2_X1    g07174(.A1(new_n7122_), .A2(new_n7158_), .Z(new_n7368_));
  XOR2_X1    g07175(.A1(new_n7368_), .A2(new_n7114_), .Z(new_n7369_));
  NAND2_X1   g07176(.A1(new_n7123_), .A2(new_n7116_), .ZN(new_n7370_));
  INV_X1     g07177(.I(new_n7124_), .ZN(new_n7371_));
  NAND2_X1   g07178(.A1(new_n7371_), .A2(new_n7132_), .ZN(new_n7372_));
  NAND2_X1   g07179(.A1(new_n7372_), .A2(new_n7370_), .ZN(new_n7373_));
  XOR2_X1    g07180(.A1(new_n7373_), .A2(new_n7369_), .Z(new_n7374_));
  XOR2_X1    g07181(.A1(new_n7374_), .A2(new_n7367_), .Z(new_n7375_));
  INV_X1     g07182(.I(new_n7375_), .ZN(new_n7376_));
  XOR2_X1    g07183(.A1(new_n7364_), .A2(new_n7376_), .Z(new_n7377_));
  XOR2_X1    g07184(.A1(new_n7377_), .A2(new_n7332_), .Z(new_n7378_));
  XOR2_X1    g07185(.A1(new_n7329_), .A2(new_n7378_), .Z(new_n7379_));
  INV_X1     g07186(.I(new_n7283_), .ZN(new_n7380_));
  NAND2_X1   g07187(.A1(new_n7380_), .A2(new_n7262_), .ZN(new_n7381_));
  INV_X1     g07188(.I(new_n7284_), .ZN(new_n7382_));
  NAND2_X1   g07189(.A1(new_n7382_), .A2(new_n7250_), .ZN(new_n7383_));
  NAND2_X1   g07190(.A1(new_n7383_), .A2(new_n7381_), .ZN(new_n7384_));
  NAND2_X1   g07191(.A1(new_n7224_), .A2(new_n7237_), .ZN(new_n7385_));
  NAND2_X1   g07192(.A1(new_n7243_), .A2(new_n7385_), .ZN(new_n7386_));
  NAND3_X1   g07193(.A1(new_n1628_), .A2(\a[47] ), .A3(\a[52] ), .ZN(new_n7387_));
  NOR4_X1    g07194(.A1(new_n417_), .A2(new_n742_), .A3(new_n4312_), .A4(new_n5425_), .ZN(new_n7388_));
  NOR2_X1    g07195(.A1(new_n1264_), .A2(new_n6563_), .ZN(new_n7389_));
  OAI21_X1   g07196(.A1(new_n7389_), .A2(new_n7388_), .B(new_n7387_), .ZN(new_n7390_));
  NAND3_X1   g07197(.A1(new_n7390_), .A2(\a[10] ), .A3(\a[53] ), .ZN(new_n7391_));
  NAND2_X1   g07198(.A1(new_n7390_), .A2(new_n7387_), .ZN(new_n7392_));
  AOI22_X1   g07199(.A1(\a[11] ), .A2(\a[52] ), .B1(\a[16] ), .B2(\a[47] ), .ZN(new_n7393_));
  OAI21_X1   g07200(.A1(new_n7392_), .A2(new_n7393_), .B(new_n7391_), .ZN(new_n7394_));
  NOR2_X1    g07201(.A1(new_n4178_), .A2(new_n5617_), .ZN(new_n7395_));
  INV_X1     g07202(.I(new_n7395_), .ZN(new_n7396_));
  NAND2_X1   g07203(.A1(\a[18] ), .A2(\a[54] ), .ZN(new_n7397_));
  OAI22_X1   g07204(.A1(new_n1275_), .A2(new_n4430_), .B1(new_n5544_), .B2(new_n7397_), .ZN(new_n7398_));
  OAI21_X1   g07205(.A1(new_n1543_), .A2(new_n7396_), .B(new_n7398_), .ZN(new_n7399_));
  NAND3_X1   g07206(.A1(new_n7399_), .A2(\a[18] ), .A3(\a[45] ), .ZN(new_n7400_));
  AOI22_X1   g07207(.A1(\a[9] ), .A2(\a[54] ), .B1(\a[17] ), .B2(\a[46] ), .ZN(new_n7401_));
  NOR2_X1    g07208(.A1(new_n1543_), .A2(new_n7396_), .ZN(new_n7402_));
  NOR2_X1    g07209(.A1(new_n7398_), .A2(new_n7402_), .ZN(new_n7403_));
  INV_X1     g07210(.I(new_n7403_), .ZN(new_n7404_));
  OAI21_X1   g07211(.A1(new_n7401_), .A2(new_n7404_), .B(new_n7400_), .ZN(new_n7405_));
  XOR2_X1    g07212(.A1(new_n7405_), .A2(new_n7394_), .Z(new_n7406_));
  NAND3_X1   g07213(.A1(new_n5917_), .A2(\a[12] ), .A3(\a[51] ), .ZN(new_n7407_));
  NAND2_X1   g07214(.A1(new_n4902_), .A2(new_n1101_), .ZN(new_n7408_));
  AOI22_X1   g07215(.A1(new_n7407_), .A2(new_n7408_), .B1(new_n763_), .B2(new_n5439_), .ZN(new_n7409_));
  AOI22_X1   g07216(.A1(\a[12] ), .A2(\a[51] ), .B1(\a[13] ), .B2(\a[50] ), .ZN(new_n7410_));
  NAND2_X1   g07217(.A1(new_n763_), .A2(new_n5439_), .ZN(new_n7411_));
  NAND3_X1   g07218(.A1(new_n7411_), .A2(new_n7407_), .A3(new_n7408_), .ZN(new_n7412_));
  OAI22_X1   g07219(.A1(new_n7409_), .A2(new_n6379_), .B1(new_n7412_), .B2(new_n7410_), .ZN(new_n7413_));
  XOR2_X1    g07220(.A1(new_n7406_), .A2(new_n7413_), .Z(new_n7414_));
  AOI22_X1   g07221(.A1(\a[6] ), .A2(\a[57] ), .B1(\a[20] ), .B2(\a[43] ), .ZN(new_n7415_));
  NOR4_X1    g07222(.A1(new_n367_), .A2(new_n1043_), .A3(new_n3666_), .A4(new_n6298_), .ZN(new_n7416_));
  NOR3_X1    g07223(.A1(new_n7415_), .A2(new_n1299_), .A3(new_n3221_), .ZN(new_n7417_));
  NOR2_X1    g07224(.A1(new_n7417_), .A2(new_n7416_), .ZN(new_n7418_));
  INV_X1     g07225(.I(new_n7418_), .ZN(new_n7419_));
  NOR2_X1    g07226(.A1(new_n1299_), .A2(new_n3221_), .ZN(new_n7420_));
  OAI21_X1   g07227(.A1(new_n7416_), .A2(new_n7415_), .B(new_n7420_), .ZN(new_n7421_));
  OAI21_X1   g07228(.A1(new_n7419_), .A2(new_n7415_), .B(new_n7421_), .ZN(new_n7422_));
  NOR2_X1    g07229(.A1(new_n2030_), .A2(new_n2274_), .ZN(new_n7423_));
  NOR2_X1    g07230(.A1(new_n3210_), .A2(new_n7423_), .ZN(new_n7424_));
  NOR2_X1    g07231(.A1(new_n759_), .A2(new_n4702_), .ZN(new_n7425_));
  INV_X1     g07232(.I(new_n7423_), .ZN(new_n7426_));
  NOR2_X1    g07233(.A1(new_n3833_), .A2(new_n7426_), .ZN(new_n7427_));
  OAI21_X1   g07234(.A1(new_n7427_), .A2(new_n7424_), .B(new_n7425_), .ZN(new_n7428_));
  INV_X1     g07235(.I(new_n7424_), .ZN(new_n7429_));
  AOI21_X1   g07236(.A1(new_n7425_), .A2(new_n7429_), .B(new_n7427_), .ZN(new_n7430_));
  INV_X1     g07237(.I(new_n7430_), .ZN(new_n7431_));
  OAI21_X1   g07238(.A1(new_n7431_), .A2(new_n7424_), .B(new_n7428_), .ZN(new_n7432_));
  XNOR2_X1   g07239(.A1(new_n7432_), .A2(new_n7422_), .ZN(new_n7433_));
  NOR3_X1    g07240(.A1(new_n1637_), .A2(new_n3859_), .A3(new_n5680_), .ZN(new_n7434_));
  NAND3_X1   g07241(.A1(new_n1533_), .A2(\a[44] ), .A3(\a[56] ), .ZN(new_n7435_));
  NAND2_X1   g07242(.A1(new_n7184_), .A2(new_n693_), .ZN(new_n7436_));
  AOI21_X1   g07243(.A1(new_n7435_), .A2(new_n7436_), .B(new_n7434_), .ZN(new_n7437_));
  NAND2_X1   g07244(.A1(\a[7] ), .A2(\a[56] ), .ZN(new_n7438_));
  NOR2_X1    g07245(.A1(new_n7437_), .A2(new_n7434_), .ZN(new_n7439_));
  INV_X1     g07246(.I(new_n7439_), .ZN(new_n7440_));
  AOI22_X1   g07247(.A1(\a[8] ), .A2(\a[55] ), .B1(\a[19] ), .B2(\a[44] ), .ZN(new_n7441_));
  OAI22_X1   g07248(.A1(new_n7440_), .A2(new_n7441_), .B1(new_n7437_), .B2(new_n7438_), .ZN(new_n7442_));
  XOR2_X1    g07249(.A1(new_n7433_), .A2(new_n7442_), .Z(new_n7443_));
  AOI22_X1   g07250(.A1(\a[21] ), .A2(\a[42] ), .B1(\a[22] ), .B2(\a[41] ), .ZN(new_n7444_));
  NAND2_X1   g07251(.A1(\a[5] ), .A2(\a[58] ), .ZN(new_n7445_));
  NOR2_X1    g07252(.A1(new_n1456_), .A2(new_n4667_), .ZN(new_n7446_));
  NOR3_X1    g07253(.A1(new_n7446_), .A2(new_n7444_), .A3(new_n7445_), .ZN(new_n7447_));
  NOR2_X1    g07254(.A1(new_n7447_), .A2(new_n7446_), .ZN(new_n7448_));
  INV_X1     g07255(.I(new_n7448_), .ZN(new_n7449_));
  OAI22_X1   g07256(.A1(new_n7449_), .A2(new_n7444_), .B1(new_n7445_), .B2(new_n7447_), .ZN(new_n7450_));
  NOR2_X1    g07257(.A1(new_n6548_), .A2(new_n6723_), .ZN(new_n7451_));
  INV_X1     g07258(.I(new_n7451_), .ZN(new_n7452_));
  NOR2_X1    g07259(.A1(new_n6723_), .A2(new_n6897_), .ZN(new_n7453_));
  INV_X1     g07260(.I(new_n7453_), .ZN(new_n7454_));
  OAI22_X1   g07261(.A1(new_n246_), .A2(new_n7454_), .B1(new_n6899_), .B2(new_n251_), .ZN(new_n7455_));
  OAI21_X1   g07262(.A1(new_n370_), .A2(new_n7452_), .B(new_n7455_), .ZN(new_n7456_));
  NAND3_X1   g07263(.A1(new_n7456_), .A2(\a[2] ), .A3(\a[61] ), .ZN(new_n7457_));
  AOI22_X1   g07264(.A1(\a[3] ), .A2(\a[60] ), .B1(\a[4] ), .B2(\a[59] ), .ZN(new_n7458_));
  NOR2_X1    g07265(.A1(new_n7452_), .A2(new_n370_), .ZN(new_n7459_));
  NOR2_X1    g07266(.A1(new_n7455_), .A2(new_n7459_), .ZN(new_n7460_));
  INV_X1     g07267(.I(new_n7460_), .ZN(new_n7461_));
  OAI21_X1   g07268(.A1(new_n7458_), .A2(new_n7461_), .B(new_n7457_), .ZN(new_n7462_));
  XOR2_X1    g07269(.A1(new_n7462_), .A2(new_n7172_), .Z(new_n7463_));
  XOR2_X1    g07270(.A1(new_n7463_), .A2(new_n7450_), .Z(new_n7464_));
  XNOR2_X1   g07271(.A1(new_n7464_), .A2(new_n7443_), .ZN(new_n7465_));
  XOR2_X1    g07272(.A1(new_n7465_), .A2(new_n7414_), .Z(new_n7466_));
  XNOR2_X1   g07273(.A1(new_n7386_), .A2(new_n7466_), .ZN(new_n7467_));
  XOR2_X1    g07274(.A1(new_n7467_), .A2(new_n7384_), .Z(new_n7468_));
  XOR2_X1    g07275(.A1(new_n7379_), .A2(new_n7468_), .Z(new_n7469_));
  INV_X1     g07276(.I(new_n7469_), .ZN(new_n7470_));
  OR2_X2     g07277(.A1(new_n7198_), .A2(new_n7245_), .Z(new_n7471_));
  INV_X1     g07278(.I(new_n7246_), .ZN(new_n7472_));
  OAI21_X1   g07279(.A1(new_n7472_), .A2(new_n7195_), .B(new_n7471_), .ZN(new_n7473_));
  NAND2_X1   g07280(.A1(new_n7108_), .A2(new_n7193_), .ZN(new_n7474_));
  NAND2_X1   g07281(.A1(new_n7194_), .A2(new_n7003_), .ZN(new_n7475_));
  NAND2_X1   g07282(.A1(new_n7475_), .A2(new_n7474_), .ZN(new_n7476_));
  INV_X1     g07283(.I(new_n7476_), .ZN(new_n7477_));
  INV_X1     g07284(.I(new_n7215_), .ZN(new_n7478_));
  NAND2_X1   g07285(.A1(new_n7478_), .A2(new_n7218_), .ZN(new_n7479_));
  NAND2_X1   g07286(.A1(new_n7201_), .A2(new_n7219_), .ZN(new_n7480_));
  NAND2_X1   g07287(.A1(new_n7480_), .A2(new_n7479_), .ZN(new_n7481_));
  AND2_X2    g07288(.A1(new_n7281_), .A2(new_n7270_), .Z(new_n7482_));
  INV_X1     g07289(.I(new_n7268_), .ZN(new_n7483_));
  NOR2_X1    g07290(.A1(new_n7282_), .A2(new_n7483_), .ZN(new_n7484_));
  NOR2_X1    g07291(.A1(new_n7484_), .A2(new_n7482_), .ZN(new_n7485_));
  NAND2_X1   g07292(.A1(new_n7260_), .A2(new_n7256_), .ZN(new_n7486_));
  NAND2_X1   g07293(.A1(new_n7261_), .A2(new_n7253_), .ZN(new_n7487_));
  NAND2_X1   g07294(.A1(new_n7487_), .A2(new_n7486_), .ZN(new_n7488_));
  XNOR2_X1   g07295(.A1(new_n7488_), .A2(new_n7485_), .ZN(new_n7489_));
  XOR2_X1    g07296(.A1(new_n7489_), .A2(new_n7481_), .Z(new_n7490_));
  XOR2_X1    g07297(.A1(new_n7188_), .A2(new_n7130_), .Z(new_n7491_));
  XOR2_X1    g07298(.A1(new_n7491_), .A2(new_n7179_), .Z(new_n7492_));
  INV_X1     g07299(.I(new_n7492_), .ZN(new_n7493_));
  XOR2_X1    g07300(.A1(new_n7212_), .A2(new_n7138_), .Z(new_n7494_));
  XNOR2_X1   g07301(.A1(new_n7494_), .A2(new_n7148_), .ZN(new_n7495_));
  NOR2_X1    g07302(.A1(new_n6911_), .A2(new_n6904_), .ZN(new_n7496_));
  NOR2_X1    g07303(.A1(new_n7266_), .A2(new_n7496_), .ZN(new_n7497_));
  XNOR2_X1   g07304(.A1(new_n7495_), .A2(new_n7497_), .ZN(new_n7498_));
  INV_X1     g07305(.I(new_n7498_), .ZN(new_n7499_));
  NOR2_X1    g07306(.A1(new_n7499_), .A2(new_n7493_), .ZN(new_n7500_));
  INV_X1     g07307(.I(new_n7500_), .ZN(new_n7501_));
  NAND2_X1   g07308(.A1(new_n7499_), .A2(new_n7493_), .ZN(new_n7502_));
  AND2_X2    g07309(.A1(new_n7501_), .A2(new_n7502_), .Z(new_n7503_));
  NOR2_X1    g07310(.A1(new_n7279_), .A2(new_n7275_), .ZN(new_n7504_));
  NAND2_X1   g07311(.A1(new_n6937_), .A2(new_n7020_), .ZN(new_n7505_));
  NAND2_X1   g07312(.A1(new_n7202_), .A2(new_n7214_), .ZN(new_n7506_));
  NAND2_X1   g07313(.A1(new_n7506_), .A2(new_n7505_), .ZN(new_n7507_));
  NAND2_X1   g07314(.A1(new_n7269_), .A2(new_n6923_), .ZN(new_n7508_));
  OAI21_X1   g07315(.A1(new_n7036_), .A2(new_n7057_), .B(new_n7508_), .ZN(new_n7509_));
  XOR2_X1    g07316(.A1(new_n7507_), .A2(new_n7509_), .Z(new_n7510_));
  XNOR2_X1   g07317(.A1(new_n7510_), .A2(new_n7504_), .ZN(new_n7511_));
  INV_X1     g07318(.I(new_n7161_), .ZN(new_n7512_));
  NAND2_X1   g07319(.A1(new_n7191_), .A2(new_n7512_), .ZN(new_n7513_));
  OAI21_X1   g07320(.A1(new_n7192_), .A2(new_n7133_), .B(new_n7513_), .ZN(new_n7514_));
  XOR2_X1    g07321(.A1(new_n7514_), .A2(new_n7511_), .Z(new_n7515_));
  OR2_X2     g07322(.A1(new_n7515_), .A2(new_n7503_), .Z(new_n7516_));
  NAND2_X1   g07323(.A1(new_n7515_), .A2(new_n7503_), .ZN(new_n7517_));
  AND2_X2    g07324(.A1(new_n7516_), .A2(new_n7517_), .Z(new_n7518_));
  NOR2_X1    g07325(.A1(new_n7518_), .A2(new_n7490_), .ZN(new_n7519_));
  AND2_X2    g07326(.A1(new_n7518_), .A2(new_n7490_), .Z(new_n7520_));
  NOR3_X1    g07327(.A1(new_n7477_), .A2(new_n7520_), .A3(new_n7519_), .ZN(new_n7521_));
  NOR2_X1    g07328(.A1(new_n7521_), .A2(new_n7520_), .ZN(new_n7522_));
  INV_X1     g07329(.I(new_n7522_), .ZN(new_n7523_));
  OAI22_X1   g07330(.A1(new_n7523_), .A2(new_n7519_), .B1(new_n7477_), .B2(new_n7521_), .ZN(new_n7524_));
  NOR2_X1    g07331(.A1(new_n7473_), .A2(new_n7524_), .ZN(new_n7525_));
  NAND2_X1   g07332(.A1(new_n7473_), .A2(new_n7524_), .ZN(new_n7526_));
  INV_X1     g07333(.I(new_n7526_), .ZN(new_n7527_));
  NOR2_X1    g07334(.A1(new_n7527_), .A2(new_n7525_), .ZN(new_n7528_));
  NAND2_X1   g07335(.A1(new_n7528_), .A2(new_n7470_), .ZN(new_n7529_));
  INV_X1     g07336(.I(new_n7529_), .ZN(new_n7530_));
  NOR2_X1    g07337(.A1(new_n7528_), .A2(new_n7470_), .ZN(new_n7531_));
  NOR2_X1    g07338(.A1(new_n7530_), .A2(new_n7531_), .ZN(new_n7532_));
  NOR2_X1    g07339(.A1(new_n7327_), .A2(new_n7532_), .ZN(new_n7533_));
  NAND2_X1   g07340(.A1(new_n7327_), .A2(new_n7532_), .ZN(new_n7534_));
  INV_X1     g07341(.I(new_n7534_), .ZN(new_n7535_));
  NOR2_X1    g07342(.A1(new_n7535_), .A2(new_n7533_), .ZN(new_n7536_));
  XOR2_X1    g07343(.A1(new_n7325_), .A2(new_n7536_), .Z(\asquared[64] ));
  NAND2_X1   g07344(.A1(new_n7514_), .A2(new_n7511_), .ZN(new_n7538_));
  NAND2_X1   g07345(.A1(new_n7517_), .A2(new_n7538_), .ZN(new_n7539_));
  NAND3_X1   g07346(.A1(new_n5532_), .A2(\a[17] ), .A3(\a[57] ), .ZN(new_n7540_));
  NAND2_X1   g07347(.A1(\a[17] ), .A2(\a[58] ), .ZN(new_n7541_));
  NOR3_X1    g07348(.A1(new_n7541_), .A2(new_n367_), .A3(new_n4312_), .ZN(new_n7542_));
  NOR2_X1    g07349(.A1(new_n6804_), .A2(new_n374_), .ZN(new_n7543_));
  OAI21_X1   g07350(.A1(new_n7543_), .A2(new_n7542_), .B(new_n7540_), .ZN(new_n7544_));
  NAND3_X1   g07351(.A1(new_n7544_), .A2(\a[6] ), .A3(\a[58] ), .ZN(new_n7545_));
  NAND2_X1   g07352(.A1(new_n7544_), .A2(new_n7540_), .ZN(new_n7546_));
  AOI22_X1   g07353(.A1(\a[7] ), .A2(\a[57] ), .B1(\a[17] ), .B2(\a[47] ), .ZN(new_n7547_));
  OAI21_X1   g07354(.A1(new_n7546_), .A2(new_n7547_), .B(new_n7545_), .ZN(new_n7548_));
  NAND2_X1   g07355(.A1(new_n1452_), .A2(new_n4180_), .ZN(new_n7549_));
  OAI22_X1   g07356(.A1(new_n1382_), .A2(new_n4343_), .B1(new_n2647_), .B2(new_n3861_), .ZN(new_n7550_));
  NAND2_X1   g07357(.A1(new_n7550_), .A2(new_n7549_), .ZN(new_n7551_));
  NAND3_X1   g07358(.A1(new_n7551_), .A2(\a[20] ), .A3(\a[44] ), .ZN(new_n7552_));
  AOI22_X1   g07359(.A1(\a[21] ), .A2(\a[43] ), .B1(\a[22] ), .B2(\a[42] ), .ZN(new_n7553_));
  NAND2_X1   g07360(.A1(new_n7551_), .A2(new_n7549_), .ZN(new_n7554_));
  OAI21_X1   g07361(.A1(new_n7553_), .A2(new_n7554_), .B(new_n7552_), .ZN(new_n7555_));
  XOR2_X1    g07362(.A1(new_n7555_), .A2(new_n7548_), .Z(new_n7556_));
  NAND2_X1   g07363(.A1(new_n1442_), .A2(new_n3328_), .ZN(new_n7557_));
  NAND2_X1   g07364(.A1(new_n1528_), .A2(new_n4534_), .ZN(new_n7558_));
  AOI22_X1   g07365(.A1(new_n7557_), .A2(new_n7558_), .B1(new_n1778_), .B2(new_n3550_), .ZN(new_n7559_));
  NAND2_X1   g07366(.A1(\a[23] ), .A2(\a[41] ), .ZN(new_n7560_));
  AOI22_X1   g07367(.A1(\a[24] ), .A2(\a[40] ), .B1(\a[25] ), .B2(\a[39] ), .ZN(new_n7561_));
  NAND2_X1   g07368(.A1(new_n1778_), .A2(new_n3550_), .ZN(new_n7562_));
  NAND3_X1   g07369(.A1(new_n7562_), .A2(new_n7557_), .A3(new_n7558_), .ZN(new_n7563_));
  OAI22_X1   g07370(.A1(new_n7559_), .A2(new_n7560_), .B1(new_n7563_), .B2(new_n7561_), .ZN(new_n7564_));
  XNOR2_X1   g07371(.A1(new_n7556_), .A2(new_n7564_), .ZN(new_n7565_));
  INV_X1     g07372(.I(new_n7565_), .ZN(new_n7566_));
  AOI22_X1   g07373(.A1(\a[8] ), .A2(\a[56] ), .B1(\a[16] ), .B2(\a[48] ), .ZN(new_n7567_));
  NOR3_X1    g07374(.A1(new_n1365_), .A2(new_n4596_), .A3(new_n5856_), .ZN(new_n7568_));
  INV_X1     g07375(.I(new_n7568_), .ZN(new_n7569_));
  NOR2_X1    g07376(.A1(new_n1566_), .A2(new_n2914_), .ZN(new_n7570_));
  INV_X1     g07377(.I(new_n7570_), .ZN(new_n7571_));
  OAI21_X1   g07378(.A1(new_n7567_), .A2(new_n7571_), .B(new_n7569_), .ZN(new_n7572_));
  OAI21_X1   g07379(.A1(new_n7568_), .A2(new_n7567_), .B(new_n7570_), .ZN(new_n7573_));
  OAI21_X1   g07380(.A1(new_n7572_), .A2(new_n7567_), .B(new_n7573_), .ZN(new_n7574_));
  NOR2_X1    g07381(.A1(new_n2679_), .A2(new_n3405_), .ZN(new_n7575_));
  INV_X1     g07382(.I(new_n7575_), .ZN(new_n7576_));
  OAI22_X1   g07383(.A1(new_n1816_), .A2(new_n4190_), .B1(new_n2189_), .B2(new_n3038_), .ZN(new_n7577_));
  NAND2_X1   g07384(.A1(new_n7577_), .A2(new_n7576_), .ZN(new_n7578_));
  NAND2_X1   g07385(.A1(new_n7578_), .A2(new_n6730_), .ZN(new_n7579_));
  AOI22_X1   g07386(.A1(\a[28] ), .A2(\a[36] ), .B1(\a[29] ), .B2(\a[35] ), .ZN(new_n7580_));
  NAND2_X1   g07387(.A1(new_n7578_), .A2(new_n7576_), .ZN(new_n7581_));
  OAI21_X1   g07388(.A1(new_n7580_), .A2(new_n7581_), .B(new_n7579_), .ZN(new_n7582_));
  XOR2_X1    g07389(.A1(new_n7582_), .A2(new_n7574_), .Z(new_n7583_));
  AOI21_X1   g07390(.A1(\a[30] ), .A2(\a[34] ), .B(new_n2275_), .ZN(new_n7584_));
  OAI22_X1   g07391(.A1(new_n7584_), .A2(new_n6942_), .B1(new_n2438_), .B2(new_n3932_), .ZN(new_n7585_));
  NOR2_X1    g07392(.A1(new_n2438_), .A2(new_n3932_), .ZN(new_n7586_));
  OAI21_X1   g07393(.A1(new_n7586_), .A2(new_n7584_), .B(new_n6941_), .ZN(new_n7587_));
  OAI21_X1   g07394(.A1(new_n7584_), .A2(new_n7585_), .B(new_n7587_), .ZN(new_n7588_));
  XOR2_X1    g07395(.A1(new_n7583_), .A2(new_n7588_), .Z(new_n7589_));
  NOR2_X1    g07396(.A1(new_n6897_), .A2(new_n7144_), .ZN(new_n7590_));
  INV_X1     g07397(.I(new_n7590_), .ZN(new_n7591_));
  OAI22_X1   g07398(.A1(new_n246_), .A2(new_n7591_), .B1(new_n7146_), .B2(new_n251_), .ZN(new_n7592_));
  OAI21_X1   g07399(.A1(new_n370_), .A2(new_n7454_), .B(new_n7592_), .ZN(new_n7593_));
  NAND3_X1   g07400(.A1(new_n7593_), .A2(\a[2] ), .A3(\a[62] ), .ZN(new_n7594_));
  AOI22_X1   g07401(.A1(\a[3] ), .A2(\a[61] ), .B1(\a[4] ), .B2(\a[60] ), .ZN(new_n7595_));
  NOR2_X1    g07402(.A1(new_n7454_), .A2(new_n370_), .ZN(new_n7596_));
  NOR2_X1    g07403(.A1(new_n7592_), .A2(new_n7596_), .ZN(new_n7597_));
  INV_X1     g07404(.I(new_n7597_), .ZN(new_n7598_));
  OAI21_X1   g07405(.A1(new_n7595_), .A2(new_n7598_), .B(new_n7594_), .ZN(new_n7599_));
  NOR2_X1    g07406(.A1(new_n7339_), .A2(new_n7340_), .ZN(new_n7600_));
  AOI21_X1   g07407(.A1(new_n7346_), .A2(new_n7342_), .B(new_n7600_), .ZN(new_n7601_));
  AOI22_X1   g07408(.A1(\a[18] ), .A2(\a[46] ), .B1(\a[19] ), .B2(\a[45] ), .ZN(new_n7602_));
  NOR2_X1    g07409(.A1(new_n4430_), .A2(new_n1092_), .ZN(new_n7603_));
  OAI21_X1   g07410(.A1(new_n7603_), .A2(new_n7602_), .B(new_n6892_), .ZN(new_n7604_));
  INV_X1     g07411(.I(new_n7602_), .ZN(new_n7605_));
  AOI21_X1   g07412(.A1(new_n6892_), .A2(new_n7605_), .B(new_n7603_), .ZN(new_n7606_));
  INV_X1     g07413(.I(new_n7606_), .ZN(new_n7607_));
  OAI21_X1   g07414(.A1(new_n7607_), .A2(new_n7602_), .B(new_n7604_), .ZN(new_n7608_));
  INV_X1     g07415(.I(new_n7608_), .ZN(new_n7609_));
  XOR2_X1    g07416(.A1(new_n7601_), .A2(new_n7609_), .Z(new_n7610_));
  XOR2_X1    g07417(.A1(new_n7610_), .A2(new_n7599_), .Z(new_n7611_));
  XOR2_X1    g07418(.A1(new_n7589_), .A2(new_n7611_), .Z(new_n7612_));
  XOR2_X1    g07419(.A1(new_n7612_), .A2(new_n7566_), .Z(new_n7613_));
  XOR2_X1    g07420(.A1(new_n7539_), .A2(new_n7613_), .Z(new_n7614_));
  NOR2_X1    g07421(.A1(new_n7212_), .A2(new_n7138_), .ZN(new_n7615_));
  INV_X1     g07422(.I(new_n7494_), .ZN(new_n7616_));
  NOR2_X1    g07423(.A1(new_n7616_), .A2(new_n7148_), .ZN(new_n7617_));
  NOR2_X1    g07424(.A1(new_n7617_), .A2(new_n7615_), .ZN(new_n7618_));
  NAND2_X1   g07425(.A1(new_n7491_), .A2(new_n7179_), .ZN(new_n7619_));
  OAI21_X1   g07426(.A1(new_n7130_), .A2(new_n7188_), .B(new_n7619_), .ZN(new_n7620_));
  NAND2_X1   g07427(.A1(new_n7122_), .A2(new_n7158_), .ZN(new_n7621_));
  NAND2_X1   g07428(.A1(new_n7368_), .A2(new_n7114_), .ZN(new_n7622_));
  NAND2_X1   g07429(.A1(new_n7622_), .A2(new_n7621_), .ZN(new_n7623_));
  XOR2_X1    g07430(.A1(new_n7623_), .A2(new_n7620_), .Z(new_n7624_));
  XNOR2_X1   g07431(.A1(new_n7624_), .A2(new_n7618_), .ZN(new_n7625_));
  INV_X1     g07432(.I(new_n7625_), .ZN(new_n7626_));
  INV_X1     g07433(.I(new_n7495_), .ZN(new_n7627_));
  NOR2_X1    g07434(.A1(new_n7627_), .A2(new_n7497_), .ZN(new_n7628_));
  NOR2_X1    g07435(.A1(new_n7500_), .A2(new_n7628_), .ZN(new_n7629_));
  NAND2_X1   g07436(.A1(new_n7373_), .A2(new_n7369_), .ZN(new_n7630_));
  NAND2_X1   g07437(.A1(new_n7374_), .A2(new_n7367_), .ZN(new_n7631_));
  NAND2_X1   g07438(.A1(new_n7631_), .A2(new_n7630_), .ZN(new_n7632_));
  XOR2_X1    g07439(.A1(new_n7632_), .A2(new_n7629_), .Z(new_n7633_));
  XOR2_X1    g07440(.A1(new_n7633_), .A2(new_n7626_), .Z(new_n7634_));
  XNOR2_X1   g07441(.A1(new_n7614_), .A2(new_n7634_), .ZN(new_n7635_));
  NAND2_X1   g07442(.A1(new_n7507_), .A2(new_n7509_), .ZN(new_n7636_));
  INV_X1     g07443(.I(new_n7510_), .ZN(new_n7637_));
  OAI21_X1   g07444(.A1(new_n7637_), .A2(new_n7504_), .B(new_n7636_), .ZN(new_n7638_));
  NAND2_X1   g07445(.A1(new_n7463_), .A2(new_n7450_), .ZN(new_n7639_));
  NAND2_X1   g07446(.A1(new_n7462_), .A2(new_n7172_), .ZN(new_n7640_));
  NAND2_X1   g07447(.A1(new_n7639_), .A2(new_n7640_), .ZN(new_n7641_));
  XOR2_X1    g07448(.A1(new_n7638_), .A2(new_n7641_), .Z(new_n7642_));
  INV_X1     g07449(.I(\a[63] ), .ZN(new_n7643_));
  NOR2_X1    g07450(.A1(new_n7144_), .A2(new_n7643_), .ZN(new_n7644_));
  NAND2_X1   g07451(.A1(new_n2316_), .A2(new_n7644_), .ZN(new_n7645_));
  NAND2_X1   g07452(.A1(new_n7343_), .A2(new_n7645_), .ZN(new_n7646_));
  OAI21_X1   g07453(.A1(new_n7345_), .A2(new_n7643_), .B(new_n7646_), .ZN(new_n7647_));
  XOR2_X1    g07454(.A1(new_n7647_), .A2(new_n7431_), .Z(new_n7648_));
  NAND2_X1   g07455(.A1(new_n5862_), .A2(new_n1261_), .ZN(new_n7649_));
  OAI22_X1   g07456(.A1(new_n1265_), .A2(new_n5525_), .B1(new_n5683_), .B2(new_n833_), .ZN(new_n7650_));
  NAND2_X1   g07457(.A1(new_n7650_), .A2(new_n7649_), .ZN(new_n7651_));
  NAND3_X1   g07458(.A1(new_n7651_), .A2(\a[13] ), .A3(\a[51] ), .ZN(new_n7652_));
  AOI22_X1   g07459(.A1(\a[11] ), .A2(\a[53] ), .B1(\a[12] ), .B2(\a[52] ), .ZN(new_n7653_));
  NAND2_X1   g07460(.A1(new_n7651_), .A2(new_n7649_), .ZN(new_n7654_));
  OAI21_X1   g07461(.A1(new_n7653_), .A2(new_n7654_), .B(new_n7652_), .ZN(new_n7655_));
  NOR2_X1    g07462(.A1(new_n717_), .A2(new_n4702_), .ZN(new_n7656_));
  NAND3_X1   g07463(.A1(new_n7656_), .A2(\a[10] ), .A3(\a[54] ), .ZN(new_n7657_));
  NOR2_X1    g07464(.A1(new_n4702_), .A2(new_n5680_), .ZN(new_n7658_));
  INV_X1     g07465(.I(new_n7658_), .ZN(new_n7659_));
  OAI22_X1   g07466(.A1(new_n5820_), .A2(new_n7659_), .B1(new_n6129_), .B2(new_n539_), .ZN(new_n7660_));
  NAND2_X1   g07467(.A1(new_n7660_), .A2(new_n7657_), .ZN(new_n7661_));
  NAND3_X1   g07468(.A1(new_n7661_), .A2(\a[9] ), .A3(\a[55] ), .ZN(new_n7662_));
  NAND2_X1   g07469(.A1(new_n7661_), .A2(new_n7657_), .ZN(new_n7663_));
  AOI21_X1   g07470(.A1(\a[10] ), .A2(\a[54] ), .B(new_n7656_), .ZN(new_n7664_));
  OAI21_X1   g07471(.A1(new_n7663_), .A2(new_n7664_), .B(new_n7662_), .ZN(new_n7665_));
  XOR2_X1    g07472(.A1(new_n7655_), .A2(new_n7665_), .Z(new_n7666_));
  XNOR2_X1   g07473(.A1(new_n7666_), .A2(new_n7648_), .ZN(new_n7667_));
  XOR2_X1    g07474(.A1(new_n7642_), .A2(new_n7667_), .Z(new_n7668_));
  INV_X1     g07475(.I(new_n7668_), .ZN(new_n7669_));
  OAI21_X1   g07476(.A1(new_n7482_), .A2(new_n7484_), .B(new_n7488_), .ZN(new_n7670_));
  NAND2_X1   g07477(.A1(new_n7489_), .A2(new_n7481_), .ZN(new_n7671_));
  NAND2_X1   g07478(.A1(new_n7671_), .A2(new_n7670_), .ZN(new_n7672_));
  NAND2_X1   g07479(.A1(new_n7405_), .A2(new_n7394_), .ZN(new_n7673_));
  NAND2_X1   g07480(.A1(new_n7406_), .A2(new_n7413_), .ZN(new_n7674_));
  NAND2_X1   g07481(.A1(new_n7674_), .A2(new_n7673_), .ZN(new_n7675_));
  NAND2_X1   g07482(.A1(new_n7432_), .A2(new_n7422_), .ZN(new_n7676_));
  INV_X1     g07483(.I(new_n7433_), .ZN(new_n7677_));
  NAND2_X1   g07484(.A1(new_n7677_), .A2(new_n7442_), .ZN(new_n7678_));
  NAND2_X1   g07485(.A1(new_n7678_), .A2(new_n7676_), .ZN(new_n7679_));
  XOR2_X1    g07486(.A1(new_n7353_), .A2(new_n7412_), .Z(new_n7680_));
  XOR2_X1    g07487(.A1(new_n7680_), .A2(new_n7392_), .Z(new_n7681_));
  XOR2_X1    g07488(.A1(new_n7679_), .A2(new_n7681_), .Z(new_n7682_));
  XOR2_X1    g07489(.A1(new_n7682_), .A2(new_n7675_), .Z(new_n7683_));
  XOR2_X1    g07490(.A1(new_n7672_), .A2(new_n7683_), .Z(new_n7684_));
  XOR2_X1    g07491(.A1(new_n7684_), .A2(new_n7669_), .Z(new_n7685_));
  XNOR2_X1   g07492(.A1(new_n7522_), .A2(new_n7685_), .ZN(new_n7686_));
  XNOR2_X1   g07493(.A1(new_n7686_), .A2(new_n7635_), .ZN(new_n7687_));
  INV_X1     g07494(.I(new_n7687_), .ZN(new_n7688_));
  NAND2_X1   g07495(.A1(new_n7329_), .A2(new_n7378_), .ZN(new_n7689_));
  INV_X1     g07496(.I(new_n7379_), .ZN(new_n7690_));
  OAI21_X1   g07497(.A1(new_n7690_), .A2(new_n7468_), .B(new_n7689_), .ZN(new_n7691_));
  NAND2_X1   g07498(.A1(new_n7386_), .A2(new_n7466_), .ZN(new_n7692_));
  INV_X1     g07499(.I(new_n7467_), .ZN(new_n7693_));
  NAND2_X1   g07500(.A1(new_n7693_), .A2(new_n7384_), .ZN(new_n7694_));
  NAND2_X1   g07501(.A1(new_n7694_), .A2(new_n7692_), .ZN(new_n7695_));
  NAND2_X1   g07502(.A1(new_n7377_), .A2(new_n7332_), .ZN(new_n7696_));
  OAI21_X1   g07503(.A1(new_n7364_), .A2(new_n7376_), .B(new_n7696_), .ZN(new_n7697_));
  NAND2_X1   g07504(.A1(new_n7354_), .A2(new_n7361_), .ZN(new_n7698_));
  INV_X1     g07505(.I(new_n7698_), .ZN(new_n7699_));
  AOI21_X1   g07506(.A1(new_n7362_), .A2(new_n7347_), .B(new_n7699_), .ZN(new_n7700_));
  XOR2_X1    g07507(.A1(new_n7403_), .A2(new_n7418_), .Z(new_n7701_));
  XOR2_X1    g07508(.A1(new_n7701_), .A2(new_n7360_), .Z(new_n7702_));
  NOR2_X1    g07509(.A1(new_n7449_), .A2(new_n7461_), .ZN(new_n7703_));
  NOR2_X1    g07510(.A1(new_n7448_), .A2(new_n7460_), .ZN(new_n7704_));
  NOR2_X1    g07511(.A1(new_n7703_), .A2(new_n7704_), .ZN(new_n7705_));
  NOR2_X1    g07512(.A1(new_n7705_), .A2(new_n7440_), .ZN(new_n7706_));
  INV_X1     g07513(.I(new_n7705_), .ZN(new_n7707_));
  NOR2_X1    g07514(.A1(new_n7707_), .A2(new_n7439_), .ZN(new_n7708_));
  NOR2_X1    g07515(.A1(new_n7708_), .A2(new_n7706_), .ZN(new_n7709_));
  NAND2_X1   g07516(.A1(new_n7709_), .A2(new_n7702_), .ZN(new_n7710_));
  INV_X1     g07517(.I(new_n7710_), .ZN(new_n7711_));
  NOR2_X1    g07518(.A1(new_n7709_), .A2(new_n7702_), .ZN(new_n7712_));
  NOR2_X1    g07519(.A1(new_n7711_), .A2(new_n7712_), .ZN(new_n7713_));
  INV_X1     g07520(.I(new_n7713_), .ZN(new_n7714_));
  NOR2_X1    g07521(.A1(new_n7714_), .A2(new_n7700_), .ZN(new_n7715_));
  INV_X1     g07522(.I(new_n7715_), .ZN(new_n7716_));
  NAND2_X1   g07523(.A1(new_n7714_), .A2(new_n7700_), .ZN(new_n7717_));
  AND2_X2    g07524(.A1(new_n7716_), .A2(new_n7717_), .Z(new_n7718_));
  INV_X1     g07525(.I(new_n7464_), .ZN(new_n7719_));
  NAND2_X1   g07526(.A1(new_n7465_), .A2(new_n7414_), .ZN(new_n7720_));
  OAI21_X1   g07527(.A1(new_n7443_), .A2(new_n7719_), .B(new_n7720_), .ZN(new_n7721_));
  NAND2_X1   g07528(.A1(new_n7334_), .A2(new_n7337_), .ZN(new_n7722_));
  NAND2_X1   g07529(.A1(new_n7338_), .A2(new_n7363_), .ZN(new_n7723_));
  NAND2_X1   g07530(.A1(new_n7723_), .A2(new_n7722_), .ZN(new_n7724_));
  XOR2_X1    g07531(.A1(new_n7724_), .A2(new_n7721_), .Z(new_n7725_));
  XOR2_X1    g07532(.A1(new_n7725_), .A2(new_n7718_), .Z(new_n7726_));
  XNOR2_X1   g07533(.A1(new_n7697_), .A2(new_n7726_), .ZN(new_n7727_));
  XOR2_X1    g07534(.A1(new_n7695_), .A2(new_n7727_), .Z(new_n7728_));
  XOR2_X1    g07535(.A1(new_n7691_), .A2(new_n7728_), .Z(new_n7729_));
  XOR2_X1    g07536(.A1(new_n7729_), .A2(new_n7688_), .Z(new_n7730_));
  INV_X1     g07537(.I(new_n7730_), .ZN(new_n7731_));
  NOR2_X1    g07538(.A1(new_n7530_), .A2(new_n7527_), .ZN(new_n7732_));
  NOR2_X1    g07539(.A1(new_n7731_), .A2(new_n7732_), .ZN(new_n7733_));
  INV_X1     g07540(.I(new_n7733_), .ZN(new_n7734_));
  AOI21_X1   g07541(.A1(new_n7324_), .A2(new_n7311_), .B(new_n7533_), .ZN(new_n7735_));
  NOR2_X1    g07542(.A1(new_n7735_), .A2(new_n7535_), .ZN(new_n7736_));
  INV_X1     g07543(.I(new_n7311_), .ZN(new_n7737_));
  INV_X1     g07544(.I(new_n7533_), .ZN(new_n7738_));
  OAI21_X1   g07545(.A1(new_n7322_), .A2(new_n7737_), .B(new_n7738_), .ZN(new_n7739_));
  NAND2_X1   g07546(.A1(new_n7731_), .A2(new_n7732_), .ZN(new_n7740_));
  INV_X1     g07547(.I(new_n7740_), .ZN(new_n7741_));
  AOI21_X1   g07548(.A1(new_n7739_), .A2(new_n7534_), .B(new_n7741_), .ZN(new_n7742_));
  NAND2_X1   g07549(.A1(new_n7734_), .A2(new_n7740_), .ZN(new_n7743_));
  AOI22_X1   g07550(.A1(new_n7742_), .A2(new_n7734_), .B1(new_n7736_), .B2(new_n7743_), .ZN(\asquared[65] ));
  OAI21_X1   g07551(.A1(new_n7735_), .A2(new_n7535_), .B(new_n7740_), .ZN(new_n7745_));
  NAND2_X1   g07552(.A1(new_n7745_), .A2(new_n7734_), .ZN(new_n7746_));
  NAND4_X1   g07553(.A1(\a[10] ), .A2(\a[20] ), .A3(\a[45] ), .A4(\a[55] ), .ZN(new_n7747_));
  NOR2_X1    g07554(.A1(new_n1043_), .A2(new_n5856_), .ZN(new_n7748_));
  INV_X1     g07555(.I(new_n7748_), .ZN(new_n7749_));
  OAI22_X1   g07556(.A1(new_n5544_), .A2(new_n7749_), .B1(new_n7185_), .B2(new_n539_), .ZN(new_n7750_));
  NAND2_X1   g07557(.A1(new_n7750_), .A2(new_n7747_), .ZN(new_n7751_));
  NAND3_X1   g07558(.A1(new_n7751_), .A2(\a[9] ), .A3(\a[56] ), .ZN(new_n7752_));
  NAND2_X1   g07559(.A1(new_n7751_), .A2(new_n7747_), .ZN(new_n7753_));
  AOI22_X1   g07560(.A1(\a[10] ), .A2(\a[55] ), .B1(\a[20] ), .B2(\a[45] ), .ZN(new_n7754_));
  OAI21_X1   g07561(.A1(new_n7753_), .A2(new_n7754_), .B(new_n7752_), .ZN(new_n7755_));
  NAND2_X1   g07562(.A1(new_n1778_), .A2(new_n4534_), .ZN(new_n7756_));
  INV_X1     g07563(.I(new_n5239_), .ZN(new_n7757_));
  OAI22_X1   g07564(.A1(new_n1443_), .A2(new_n7757_), .B1(new_n1529_), .B2(new_n4667_), .ZN(new_n7758_));
  NAND2_X1   g07565(.A1(new_n7758_), .A2(new_n7756_), .ZN(new_n7759_));
  NAND3_X1   g07566(.A1(new_n7759_), .A2(\a[23] ), .A3(\a[42] ), .ZN(new_n7760_));
  AOI22_X1   g07567(.A1(\a[24] ), .A2(\a[41] ), .B1(\a[25] ), .B2(\a[40] ), .ZN(new_n7761_));
  NAND2_X1   g07568(.A1(new_n7759_), .A2(new_n7756_), .ZN(new_n7762_));
  OAI21_X1   g07569(.A1(new_n7761_), .A2(new_n7762_), .B(new_n7760_), .ZN(new_n7763_));
  XOR2_X1    g07570(.A1(new_n7763_), .A2(new_n7755_), .Z(new_n7764_));
  NAND2_X1   g07571(.A1(new_n1971_), .A2(new_n4209_), .ZN(new_n7765_));
  NAND2_X1   g07572(.A1(new_n2412_), .A2(new_n4545_), .ZN(new_n7766_));
  AOI22_X1   g07573(.A1(new_n7765_), .A2(new_n7766_), .B1(new_n2103_), .B2(new_n3803_), .ZN(new_n7767_));
  NAND2_X1   g07574(.A1(\a[26] ), .A2(\a[39] ), .ZN(new_n7768_));
  AOI22_X1   g07575(.A1(\a[27] ), .A2(\a[38] ), .B1(\a[28] ), .B2(\a[37] ), .ZN(new_n7769_));
  NAND2_X1   g07576(.A1(new_n2103_), .A2(new_n3803_), .ZN(new_n7770_));
  NAND3_X1   g07577(.A1(new_n7770_), .A2(new_n7765_), .A3(new_n7766_), .ZN(new_n7771_));
  OAI22_X1   g07578(.A1(new_n7767_), .A2(new_n7768_), .B1(new_n7771_), .B2(new_n7769_), .ZN(new_n7772_));
  XNOR2_X1   g07579(.A1(new_n7764_), .A2(new_n7772_), .ZN(new_n7773_));
  NOR2_X1    g07580(.A1(new_n3833_), .A2(new_n3932_), .ZN(new_n7774_));
  NOR2_X1    g07581(.A1(new_n2438_), .A2(new_n2746_), .ZN(new_n7775_));
  NOR2_X1    g07582(.A1(new_n2637_), .A2(new_n3402_), .ZN(new_n7776_));
  NOR2_X1    g07583(.A1(new_n7775_), .A2(new_n7776_), .ZN(new_n7777_));
  NOR2_X1    g07584(.A1(new_n7777_), .A2(new_n7774_), .ZN(new_n7778_));
  AOI21_X1   g07585(.A1(\a[31] ), .A2(\a[34] ), .B(new_n2636_), .ZN(new_n7779_));
  NOR2_X1    g07586(.A1(new_n7778_), .A2(new_n7774_), .ZN(new_n7780_));
  INV_X1     g07587(.I(new_n7780_), .ZN(new_n7781_));
  OAI22_X1   g07588(.A1(new_n7781_), .A2(new_n7779_), .B1(new_n3402_), .B2(new_n7778_), .ZN(new_n7782_));
  AOI22_X1   g07589(.A1(\a[11] ), .A2(\a[54] ), .B1(\a[19] ), .B2(\a[46] ), .ZN(new_n7783_));
  NOR4_X1    g07590(.A1(new_n513_), .A2(new_n979_), .A3(new_n4178_), .A4(new_n5617_), .ZN(new_n7784_));
  INV_X1     g07591(.I(new_n7784_), .ZN(new_n7785_));
  NOR2_X1    g07592(.A1(new_n1814_), .A2(new_n2626_), .ZN(new_n7786_));
  INV_X1     g07593(.I(new_n7786_), .ZN(new_n7787_));
  OAI21_X1   g07594(.A1(new_n7783_), .A2(new_n7787_), .B(new_n7785_), .ZN(new_n7788_));
  OAI21_X1   g07595(.A1(new_n7784_), .A2(new_n7783_), .B(new_n7786_), .ZN(new_n7789_));
  OAI21_X1   g07596(.A1(new_n7788_), .A2(new_n7783_), .B(new_n7789_), .ZN(new_n7790_));
  XNOR2_X1   g07597(.A1(new_n7782_), .A2(new_n7790_), .ZN(new_n7791_));
  INV_X1     g07598(.I(new_n5575_), .ZN(new_n7792_));
  AOI21_X1   g07599(.A1(\a[3] ), .A2(\a[62] ), .B(\a[33] ), .ZN(new_n7793_));
  NOR3_X1    g07600(.A1(new_n225_), .A2(new_n2274_), .A3(new_n7144_), .ZN(new_n7794_));
  NOR3_X1    g07601(.A1(new_n7792_), .A2(new_n7793_), .A3(new_n7794_), .ZN(new_n7795_));
  NOR2_X1    g07602(.A1(new_n7795_), .A2(new_n7794_), .ZN(new_n7796_));
  INV_X1     g07603(.I(new_n7796_), .ZN(new_n7797_));
  OAI22_X1   g07604(.A1(new_n7797_), .A2(new_n7793_), .B1(new_n7792_), .B2(new_n7795_), .ZN(new_n7798_));
  XOR2_X1    g07605(.A1(new_n7791_), .A2(new_n7798_), .Z(new_n7799_));
  NOR2_X1    g07606(.A1(new_n6316_), .A2(new_n6723_), .ZN(new_n7800_));
  INV_X1     g07607(.I(new_n7800_), .ZN(new_n7801_));
  OAI22_X1   g07608(.A1(new_n373_), .A2(new_n7801_), .B1(new_n7452_), .B2(new_n371_), .ZN(new_n7802_));
  OAI21_X1   g07609(.A1(new_n374_), .A2(new_n7206_), .B(new_n7802_), .ZN(new_n7803_));
  NAND3_X1   g07610(.A1(new_n7803_), .A2(\a[5] ), .A3(\a[60] ), .ZN(new_n7804_));
  AOI22_X1   g07611(.A1(\a[6] ), .A2(\a[59] ), .B1(\a[7] ), .B2(\a[58] ), .ZN(new_n7805_));
  NOR2_X1    g07612(.A1(new_n7206_), .A2(new_n374_), .ZN(new_n7806_));
  NOR2_X1    g07613(.A1(new_n7802_), .A2(new_n7806_), .ZN(new_n7807_));
  INV_X1     g07614(.I(new_n7807_), .ZN(new_n7808_));
  OAI21_X1   g07615(.A1(new_n7805_), .A2(new_n7808_), .B(new_n7804_), .ZN(new_n7809_));
  INV_X1     g07616(.I(new_n7809_), .ZN(new_n7810_));
  AOI22_X1   g07617(.A1(\a[21] ), .A2(\a[44] ), .B1(\a[22] ), .B2(\a[43] ), .ZN(new_n7811_));
  NOR2_X1    g07618(.A1(new_n355_), .A2(new_n6298_), .ZN(new_n7812_));
  INV_X1     g07619(.I(new_n7812_), .ZN(new_n7813_));
  NOR2_X1    g07620(.A1(new_n1456_), .A2(new_n4343_), .ZN(new_n7814_));
  NOR3_X1    g07621(.A1(new_n7814_), .A2(new_n7811_), .A3(new_n7813_), .ZN(new_n7815_));
  NOR2_X1    g07622(.A1(new_n7815_), .A2(new_n7814_), .ZN(new_n7816_));
  INV_X1     g07623(.I(new_n7816_), .ZN(new_n7817_));
  OAI22_X1   g07624(.A1(new_n7817_), .A2(new_n7811_), .B1(new_n7813_), .B2(new_n7815_), .ZN(new_n7818_));
  NAND2_X1   g07625(.A1(new_n7647_), .A2(new_n7431_), .ZN(new_n7819_));
  NAND2_X1   g07626(.A1(new_n7819_), .A2(new_n7645_), .ZN(new_n7820_));
  XNOR2_X1   g07627(.A1(new_n7820_), .A2(new_n7818_), .ZN(new_n7821_));
  OR2_X2     g07628(.A1(new_n7821_), .A2(new_n7810_), .Z(new_n7822_));
  NAND2_X1   g07629(.A1(new_n7821_), .A2(new_n7810_), .ZN(new_n7823_));
  NAND2_X1   g07630(.A1(new_n7822_), .A2(new_n7823_), .ZN(new_n7824_));
  XNOR2_X1   g07631(.A1(new_n7799_), .A2(new_n7824_), .ZN(new_n7825_));
  XOR2_X1    g07632(.A1(new_n7825_), .A2(new_n7773_), .Z(new_n7826_));
  NAND2_X1   g07633(.A1(new_n7724_), .A2(new_n7721_), .ZN(new_n7827_));
  NAND2_X1   g07634(.A1(new_n7725_), .A2(new_n7718_), .ZN(new_n7828_));
  NAND2_X1   g07635(.A1(new_n7828_), .A2(new_n7827_), .ZN(new_n7829_));
  XOR2_X1    g07636(.A1(new_n7829_), .A2(new_n7826_), .Z(new_n7830_));
  NOR2_X1    g07637(.A1(new_n7708_), .A2(new_n7704_), .ZN(new_n7831_));
  NAND2_X1   g07638(.A1(new_n7353_), .A2(new_n7412_), .ZN(new_n7832_));
  NAND2_X1   g07639(.A1(new_n7680_), .A2(new_n7392_), .ZN(new_n7833_));
  NAND2_X1   g07640(.A1(new_n7833_), .A2(new_n7832_), .ZN(new_n7834_));
  NAND2_X1   g07641(.A1(new_n7701_), .A2(new_n7360_), .ZN(new_n7835_));
  OAI21_X1   g07642(.A1(new_n7403_), .A2(new_n7418_), .B(new_n7835_), .ZN(new_n7836_));
  XOR2_X1    g07643(.A1(new_n7834_), .A2(new_n7836_), .Z(new_n7837_));
  XNOR2_X1   g07644(.A1(new_n7837_), .A2(new_n7831_), .ZN(new_n7838_));
  NAND2_X1   g07645(.A1(new_n7679_), .A2(new_n7681_), .ZN(new_n7839_));
  NAND2_X1   g07646(.A1(new_n7682_), .A2(new_n7675_), .ZN(new_n7840_));
  NAND2_X1   g07647(.A1(new_n7840_), .A2(new_n7839_), .ZN(new_n7841_));
  NOR2_X1    g07648(.A1(new_n7715_), .A2(new_n7711_), .ZN(new_n7842_));
  XNOR2_X1   g07649(.A1(new_n7842_), .A2(new_n7841_), .ZN(new_n7843_));
  XOR2_X1    g07650(.A1(new_n7843_), .A2(new_n7838_), .Z(new_n7844_));
  XNOR2_X1   g07651(.A1(new_n7830_), .A2(new_n7844_), .ZN(new_n7845_));
  NAND2_X1   g07652(.A1(new_n7623_), .A2(new_n7620_), .ZN(new_n7846_));
  INV_X1     g07653(.I(new_n7624_), .ZN(new_n7847_));
  OAI21_X1   g07654(.A1(new_n7847_), .A2(new_n7618_), .B(new_n7846_), .ZN(new_n7848_));
  NAND2_X1   g07655(.A1(new_n7610_), .A2(new_n7599_), .ZN(new_n7849_));
  OAI21_X1   g07656(.A1(new_n7601_), .A2(new_n7609_), .B(new_n7849_), .ZN(new_n7850_));
  XOR2_X1    g07657(.A1(new_n7848_), .A2(new_n7850_), .Z(new_n7851_));
  NOR2_X1    g07658(.A1(new_n6897_), .A2(new_n7643_), .ZN(new_n7852_));
  NAND2_X1   g07659(.A1(\a[4] ), .A2(\a[61] ), .ZN(new_n7853_));
  NAND2_X1   g07660(.A1(\a[2] ), .A2(\a[63] ), .ZN(new_n7854_));
  AOI22_X1   g07661(.A1(new_n7852_), .A2(new_n252_), .B1(new_n7853_), .B2(new_n7854_), .ZN(new_n7855_));
  XOR2_X1    g07662(.A1(new_n7585_), .A2(new_n7855_), .Z(new_n7856_));
  NAND4_X1   g07663(.A1(\a[13] ), .A2(\a[18] ), .A3(\a[47] ), .A4(\a[52] ), .ZN(new_n7857_));
  NOR4_X1    g07664(.A1(new_n536_), .A2(new_n884_), .A3(new_n4312_), .A4(new_n5425_), .ZN(new_n7858_));
  NOR2_X1    g07665(.A1(new_n1265_), .A2(new_n6563_), .ZN(new_n7859_));
  OAI21_X1   g07666(.A1(new_n7859_), .A2(new_n7858_), .B(new_n7857_), .ZN(new_n7860_));
  NAND3_X1   g07667(.A1(new_n7860_), .A2(\a[12] ), .A3(\a[53] ), .ZN(new_n7861_));
  NAND2_X1   g07668(.A1(new_n7860_), .A2(new_n7857_), .ZN(new_n7862_));
  AOI22_X1   g07669(.A1(\a[13] ), .A2(\a[52] ), .B1(\a[18] ), .B2(\a[47] ), .ZN(new_n7863_));
  OAI21_X1   g07670(.A1(new_n7862_), .A2(new_n7863_), .B(new_n7861_), .ZN(new_n7864_));
  NAND2_X1   g07671(.A1(\a[16] ), .A2(\a[49] ), .ZN(new_n7865_));
  NAND2_X1   g07672(.A1(new_n5154_), .A2(new_n1288_), .ZN(new_n7866_));
  NOR2_X1    g07673(.A1(new_n4702_), .A2(new_n5135_), .ZN(new_n7867_));
  NAND2_X1   g07674(.A1(new_n895_), .A2(new_n7867_), .ZN(new_n7868_));
  AOI22_X1   g07675(.A1(new_n7868_), .A2(new_n7866_), .B1(new_n897_), .B2(new_n5439_), .ZN(new_n7869_));
  AOI22_X1   g07676(.A1(\a[14] ), .A2(\a[51] ), .B1(\a[15] ), .B2(\a[50] ), .ZN(new_n7870_));
  NAND2_X1   g07677(.A1(new_n897_), .A2(new_n5439_), .ZN(new_n7871_));
  NAND3_X1   g07678(.A1(new_n7871_), .A2(new_n7868_), .A3(new_n7866_), .ZN(new_n7872_));
  OAI22_X1   g07679(.A1(new_n7869_), .A2(new_n7865_), .B1(new_n7872_), .B2(new_n7870_), .ZN(new_n7873_));
  XOR2_X1    g07680(.A1(new_n7864_), .A2(new_n7873_), .Z(new_n7874_));
  XNOR2_X1   g07681(.A1(new_n7874_), .A2(new_n7856_), .ZN(new_n7875_));
  XOR2_X1    g07682(.A1(new_n7851_), .A2(new_n7875_), .Z(new_n7876_));
  NAND2_X1   g07683(.A1(new_n7555_), .A2(new_n7548_), .ZN(new_n7877_));
  NAND2_X1   g07684(.A1(new_n7556_), .A2(new_n7564_), .ZN(new_n7878_));
  NAND2_X1   g07685(.A1(new_n7878_), .A2(new_n7877_), .ZN(new_n7879_));
  XOR2_X1    g07686(.A1(new_n7581_), .A2(new_n7554_), .Z(new_n7880_));
  XOR2_X1    g07687(.A1(new_n7880_), .A2(new_n7654_), .Z(new_n7881_));
  NAND2_X1   g07688(.A1(new_n7582_), .A2(new_n7574_), .ZN(new_n7882_));
  NAND2_X1   g07689(.A1(new_n7583_), .A2(new_n7588_), .ZN(new_n7883_));
  NAND2_X1   g07690(.A1(new_n7883_), .A2(new_n7882_), .ZN(new_n7884_));
  XOR2_X1    g07691(.A1(new_n7884_), .A2(new_n7881_), .Z(new_n7885_));
  XOR2_X1    g07692(.A1(new_n7885_), .A2(new_n7879_), .Z(new_n7886_));
  OAI21_X1   g07693(.A1(new_n7500_), .A2(new_n7628_), .B(new_n7632_), .ZN(new_n7887_));
  OAI21_X1   g07694(.A1(new_n7633_), .A2(new_n7626_), .B(new_n7887_), .ZN(new_n7888_));
  XNOR2_X1   g07695(.A1(new_n7888_), .A2(new_n7886_), .ZN(new_n7889_));
  XNOR2_X1   g07696(.A1(new_n7889_), .A2(new_n7876_), .ZN(new_n7890_));
  NAND2_X1   g07697(.A1(new_n7697_), .A2(new_n7726_), .ZN(new_n7891_));
  INV_X1     g07698(.I(new_n7727_), .ZN(new_n7892_));
  NAND2_X1   g07699(.A1(new_n7695_), .A2(new_n7892_), .ZN(new_n7893_));
  NAND2_X1   g07700(.A1(new_n7893_), .A2(new_n7891_), .ZN(new_n7894_));
  XOR2_X1    g07701(.A1(new_n7894_), .A2(new_n7890_), .Z(new_n7895_));
  XNOR2_X1   g07702(.A1(new_n7895_), .A2(new_n7845_), .ZN(new_n7896_));
  INV_X1     g07703(.I(new_n7896_), .ZN(new_n7897_));
  NAND2_X1   g07704(.A1(new_n7523_), .A2(new_n7685_), .ZN(new_n7898_));
  INV_X1     g07705(.I(new_n7686_), .ZN(new_n7899_));
  OAI21_X1   g07706(.A1(new_n7899_), .A2(new_n7635_), .B(new_n7898_), .ZN(new_n7900_));
  NAND2_X1   g07707(.A1(new_n7539_), .A2(new_n7613_), .ZN(new_n7901_));
  NAND2_X1   g07708(.A1(new_n7614_), .A2(new_n7634_), .ZN(new_n7902_));
  NAND2_X1   g07709(.A1(new_n7902_), .A2(new_n7901_), .ZN(new_n7903_));
  NAND2_X1   g07710(.A1(new_n7672_), .A2(new_n7683_), .ZN(new_n7904_));
  NAND2_X1   g07711(.A1(new_n7684_), .A2(new_n7669_), .ZN(new_n7905_));
  NAND2_X1   g07712(.A1(new_n7905_), .A2(new_n7904_), .ZN(new_n7906_));
  NAND2_X1   g07713(.A1(new_n7655_), .A2(new_n7665_), .ZN(new_n7907_));
  INV_X1     g07714(.I(new_n7907_), .ZN(new_n7908_));
  AOI21_X1   g07715(.A1(new_n7666_), .A2(new_n7648_), .B(new_n7908_), .ZN(new_n7909_));
  XOR2_X1    g07716(.A1(new_n7663_), .A2(new_n7563_), .Z(new_n7910_));
  XOR2_X1    g07717(.A1(new_n7910_), .A2(new_n7546_), .Z(new_n7911_));
  XOR2_X1    g07718(.A1(new_n7597_), .A2(new_n7606_), .Z(new_n7912_));
  XOR2_X1    g07719(.A1(new_n7912_), .A2(new_n7572_), .Z(new_n7913_));
  NAND2_X1   g07720(.A1(new_n7911_), .A2(new_n7913_), .ZN(new_n7914_));
  INV_X1     g07721(.I(new_n7914_), .ZN(new_n7915_));
  NOR2_X1    g07722(.A1(new_n7911_), .A2(new_n7913_), .ZN(new_n7916_));
  NOR2_X1    g07723(.A1(new_n7915_), .A2(new_n7916_), .ZN(new_n7917_));
  INV_X1     g07724(.I(new_n7917_), .ZN(new_n7918_));
  NAND2_X1   g07725(.A1(new_n7918_), .A2(new_n7909_), .ZN(new_n7919_));
  NOR2_X1    g07726(.A1(new_n7918_), .A2(new_n7909_), .ZN(new_n7920_));
  INV_X1     g07727(.I(new_n7920_), .ZN(new_n7921_));
  AND2_X2    g07728(.A1(new_n7921_), .A2(new_n7919_), .Z(new_n7922_));
  NAND2_X1   g07729(.A1(new_n7612_), .A2(new_n7566_), .ZN(new_n7923_));
  NAND2_X1   g07730(.A1(new_n7589_), .A2(new_n7611_), .ZN(new_n7924_));
  NAND2_X1   g07731(.A1(new_n7923_), .A2(new_n7924_), .ZN(new_n7925_));
  NOR2_X1    g07732(.A1(new_n7638_), .A2(new_n7641_), .ZN(new_n7926_));
  NAND2_X1   g07733(.A1(new_n7638_), .A2(new_n7641_), .ZN(new_n7927_));
  OAI21_X1   g07734(.A1(new_n7926_), .A2(new_n7667_), .B(new_n7927_), .ZN(new_n7928_));
  XOR2_X1    g07735(.A1(new_n7928_), .A2(new_n7925_), .Z(new_n7929_));
  XOR2_X1    g07736(.A1(new_n7929_), .A2(new_n7922_), .Z(new_n7930_));
  XOR2_X1    g07737(.A1(new_n7906_), .A2(new_n7930_), .Z(new_n7931_));
  XOR2_X1    g07738(.A1(new_n7931_), .A2(new_n7903_), .Z(new_n7932_));
  NOR2_X1    g07739(.A1(new_n7900_), .A2(new_n7932_), .ZN(new_n7933_));
  NAND2_X1   g07740(.A1(new_n7900_), .A2(new_n7932_), .ZN(new_n7934_));
  INV_X1     g07741(.I(new_n7934_), .ZN(new_n7935_));
  NOR2_X1    g07742(.A1(new_n7935_), .A2(new_n7933_), .ZN(new_n7936_));
  NOR2_X1    g07743(.A1(new_n7897_), .A2(new_n7936_), .ZN(new_n7937_));
  NAND2_X1   g07744(.A1(new_n7897_), .A2(new_n7936_), .ZN(new_n7938_));
  INV_X1     g07745(.I(new_n7938_), .ZN(new_n7939_));
  NOR2_X1    g07746(.A1(new_n7939_), .A2(new_n7937_), .ZN(new_n7940_));
  INV_X1     g07747(.I(new_n7728_), .ZN(new_n7941_));
  NAND2_X1   g07748(.A1(new_n7691_), .A2(new_n7941_), .ZN(new_n7942_));
  OAI21_X1   g07749(.A1(new_n7688_), .A2(new_n7729_), .B(new_n7942_), .ZN(new_n7943_));
  NOR2_X1    g07750(.A1(new_n7940_), .A2(new_n7943_), .ZN(new_n7944_));
  NAND2_X1   g07751(.A1(new_n7940_), .A2(new_n7943_), .ZN(new_n7945_));
  INV_X1     g07752(.I(new_n7945_), .ZN(new_n7946_));
  NOR2_X1    g07753(.A1(new_n7946_), .A2(new_n7944_), .ZN(new_n7947_));
  XOR2_X1    g07754(.A1(new_n7746_), .A2(new_n7947_), .Z(\asquared[66] ));
  AOI21_X1   g07755(.A1(new_n7745_), .A2(new_n7734_), .B(new_n7944_), .ZN(new_n7949_));
  NOR2_X1    g07756(.A1(new_n7949_), .A2(new_n7946_), .ZN(new_n7950_));
  NOR2_X1    g07757(.A1(new_n7939_), .A2(new_n7935_), .ZN(new_n7951_));
  INV_X1     g07758(.I(new_n7951_), .ZN(new_n7952_));
  NAND2_X1   g07759(.A1(new_n7843_), .A2(new_n7838_), .ZN(new_n7953_));
  OAI21_X1   g07760(.A1(new_n7715_), .A2(new_n7711_), .B(new_n7841_), .ZN(new_n7954_));
  NAND2_X1   g07761(.A1(new_n7953_), .A2(new_n7954_), .ZN(new_n7955_));
  NAND2_X1   g07762(.A1(new_n7834_), .A2(new_n7836_), .ZN(new_n7956_));
  INV_X1     g07763(.I(new_n7837_), .ZN(new_n7957_));
  OAI21_X1   g07764(.A1(new_n7957_), .A2(new_n7831_), .B(new_n7956_), .ZN(new_n7958_));
  INV_X1     g07765(.I(new_n7852_), .ZN(new_n7959_));
  NAND2_X1   g07766(.A1(new_n7585_), .A2(new_n7855_), .ZN(new_n7960_));
  OAI21_X1   g07767(.A1(new_n251_), .A2(new_n7959_), .B(new_n7960_), .ZN(new_n7961_));
  XOR2_X1    g07768(.A1(new_n7961_), .A2(new_n7771_), .Z(new_n7962_));
  NAND2_X1   g07769(.A1(new_n7451_), .A2(new_n479_), .ZN(new_n7963_));
  NAND2_X1   g07770(.A1(new_n7800_), .A2(new_n645_), .ZN(new_n7964_));
  AOI22_X1   g07771(.A1(new_n7963_), .A2(new_n7964_), .B1(new_n693_), .B2(new_n7205_), .ZN(new_n7965_));
  NAND2_X1   g07772(.A1(\a[6] ), .A2(\a[60] ), .ZN(new_n7966_));
  AOI22_X1   g07773(.A1(\a[7] ), .A2(\a[59] ), .B1(\a[8] ), .B2(\a[58] ), .ZN(new_n7967_));
  NAND2_X1   g07774(.A1(new_n7205_), .A2(new_n693_), .ZN(new_n7968_));
  NAND3_X1   g07775(.A1(new_n7968_), .A2(new_n7963_), .A3(new_n7964_), .ZN(new_n7969_));
  OAI22_X1   g07776(.A1(new_n7965_), .A2(new_n7966_), .B1(new_n7969_), .B2(new_n7967_), .ZN(new_n7970_));
  XNOR2_X1   g07777(.A1(new_n7962_), .A2(new_n7970_), .ZN(new_n7971_));
  NAND2_X1   g07778(.A1(new_n7864_), .A2(new_n7873_), .ZN(new_n7972_));
  NAND2_X1   g07779(.A1(new_n7874_), .A2(new_n7856_), .ZN(new_n7973_));
  NAND2_X1   g07780(.A1(new_n7973_), .A2(new_n7972_), .ZN(new_n7974_));
  XOR2_X1    g07781(.A1(new_n7971_), .A2(new_n7974_), .Z(new_n7975_));
  XNOR2_X1   g07782(.A1(new_n7958_), .A2(new_n7975_), .ZN(new_n7976_));
  XOR2_X1    g07783(.A1(new_n7780_), .A2(new_n7796_), .Z(new_n7977_));
  XOR2_X1    g07784(.A1(new_n7977_), .A2(new_n7872_), .Z(new_n7978_));
  XOR2_X1    g07785(.A1(new_n7816_), .A2(new_n7807_), .Z(new_n7979_));
  XOR2_X1    g07786(.A1(new_n7979_), .A2(new_n7788_), .Z(new_n7980_));
  NAND2_X1   g07787(.A1(new_n7782_), .A2(new_n7790_), .ZN(new_n7981_));
  INV_X1     g07788(.I(new_n7798_), .ZN(new_n7982_));
  OAI21_X1   g07789(.A1(new_n7791_), .A2(new_n7982_), .B(new_n7981_), .ZN(new_n7983_));
  XOR2_X1    g07790(.A1(new_n7983_), .A2(new_n7980_), .Z(new_n7984_));
  XNOR2_X1   g07791(.A1(new_n7984_), .A2(new_n7978_), .ZN(new_n7985_));
  XNOR2_X1   g07792(.A1(new_n7985_), .A2(new_n7976_), .ZN(new_n7986_));
  NOR2_X1    g07793(.A1(new_n7955_), .A2(new_n7986_), .ZN(new_n7987_));
  NAND2_X1   g07794(.A1(new_n7955_), .A2(new_n7986_), .ZN(new_n7988_));
  INV_X1     g07795(.I(new_n7988_), .ZN(new_n7989_));
  NOR2_X1    g07796(.A1(new_n7989_), .A2(new_n7987_), .ZN(new_n7990_));
  INV_X1     g07797(.I(new_n7990_), .ZN(new_n7991_));
  NAND2_X1   g07798(.A1(new_n7888_), .A2(new_n7886_), .ZN(new_n7992_));
  OAI21_X1   g07799(.A1(new_n7889_), .A2(new_n7876_), .B(new_n7992_), .ZN(new_n7993_));
  NAND2_X1   g07800(.A1(new_n7763_), .A2(new_n7755_), .ZN(new_n7994_));
  NAND2_X1   g07801(.A1(new_n7764_), .A2(new_n7772_), .ZN(new_n7995_));
  NAND2_X1   g07802(.A1(new_n7995_), .A2(new_n7994_), .ZN(new_n7996_));
  XOR2_X1    g07803(.A1(new_n7753_), .A2(new_n7862_), .Z(new_n7997_));
  XOR2_X1    g07804(.A1(new_n7997_), .A2(new_n7762_), .Z(new_n7998_));
  NAND2_X1   g07805(.A1(new_n7820_), .A2(new_n7818_), .ZN(new_n7999_));
  NAND2_X1   g07806(.A1(new_n7822_), .A2(new_n7999_), .ZN(new_n8000_));
  NAND2_X1   g07807(.A1(new_n8000_), .A2(new_n7998_), .ZN(new_n8001_));
  INV_X1     g07808(.I(new_n8001_), .ZN(new_n8002_));
  NOR2_X1    g07809(.A1(new_n8000_), .A2(new_n7998_), .ZN(new_n8003_));
  NOR2_X1    g07810(.A1(new_n8002_), .A2(new_n8003_), .ZN(new_n8004_));
  NOR2_X1    g07811(.A1(new_n8004_), .A2(new_n7996_), .ZN(new_n8005_));
  NAND2_X1   g07812(.A1(new_n8004_), .A2(new_n7996_), .ZN(new_n8006_));
  INV_X1     g07813(.I(new_n8006_), .ZN(new_n8007_));
  NOR2_X1    g07814(.A1(new_n8007_), .A2(new_n8005_), .ZN(new_n8008_));
  OR2_X2     g07815(.A1(new_n7799_), .A2(new_n7824_), .Z(new_n8009_));
  OAI21_X1   g07816(.A1(new_n7825_), .A2(new_n7773_), .B(new_n8009_), .ZN(new_n8010_));
  NOR2_X1    g07817(.A1(new_n7848_), .A2(new_n7850_), .ZN(new_n8011_));
  NAND2_X1   g07818(.A1(new_n7848_), .A2(new_n7850_), .ZN(new_n8012_));
  OAI21_X1   g07819(.A1(new_n8011_), .A2(new_n7875_), .B(new_n8012_), .ZN(new_n8013_));
  NOR2_X1    g07820(.A1(new_n8010_), .A2(new_n8013_), .ZN(new_n8014_));
  NAND2_X1   g07821(.A1(new_n8010_), .A2(new_n8013_), .ZN(new_n8015_));
  INV_X1     g07822(.I(new_n8015_), .ZN(new_n8016_));
  NOR2_X1    g07823(.A1(new_n8016_), .A2(new_n8014_), .ZN(new_n8017_));
  NAND2_X1   g07824(.A1(new_n8017_), .A2(new_n8008_), .ZN(new_n8018_));
  INV_X1     g07825(.I(new_n8018_), .ZN(new_n8019_));
  NOR2_X1    g07826(.A1(new_n8017_), .A2(new_n8008_), .ZN(new_n8020_));
  NOR2_X1    g07827(.A1(new_n8019_), .A2(new_n8020_), .ZN(new_n8021_));
  XNOR2_X1   g07828(.A1(new_n7993_), .A2(new_n8021_), .ZN(new_n8022_));
  XOR2_X1    g07829(.A1(new_n8022_), .A2(new_n7991_), .Z(new_n8023_));
  INV_X1     g07830(.I(new_n7890_), .ZN(new_n8024_));
  NAND2_X1   g07831(.A1(new_n7894_), .A2(new_n8024_), .ZN(new_n8025_));
  OAI21_X1   g07832(.A1(new_n7895_), .A2(new_n7845_), .B(new_n8025_), .ZN(new_n8026_));
  XOR2_X1    g07833(.A1(new_n8026_), .A2(new_n8023_), .Z(new_n8027_));
  NAND2_X1   g07834(.A1(new_n7581_), .A2(new_n7554_), .ZN(new_n8028_));
  NAND2_X1   g07835(.A1(new_n7880_), .A2(new_n7654_), .ZN(new_n8029_));
  NAND2_X1   g07836(.A1(new_n8029_), .A2(new_n8028_), .ZN(new_n8030_));
  NAND2_X1   g07837(.A1(new_n7663_), .A2(new_n7563_), .ZN(new_n8031_));
  NAND2_X1   g07838(.A1(new_n7910_), .A2(new_n7546_), .ZN(new_n8032_));
  NAND2_X1   g07839(.A1(new_n8032_), .A2(new_n8031_), .ZN(new_n8033_));
  NAND2_X1   g07840(.A1(new_n7912_), .A2(new_n7572_), .ZN(new_n8034_));
  OAI21_X1   g07841(.A1(new_n7597_), .A2(new_n7606_), .B(new_n8034_), .ZN(new_n8035_));
  XOR2_X1    g07842(.A1(new_n8033_), .A2(new_n8035_), .Z(new_n8036_));
  XOR2_X1    g07843(.A1(new_n8036_), .A2(new_n8030_), .Z(new_n8037_));
  INV_X1     g07844(.I(new_n8037_), .ZN(new_n8038_));
  NOR2_X1    g07845(.A1(new_n7920_), .A2(new_n7915_), .ZN(new_n8039_));
  NAND2_X1   g07846(.A1(new_n7884_), .A2(new_n7881_), .ZN(new_n8040_));
  NAND2_X1   g07847(.A1(new_n7885_), .A2(new_n7879_), .ZN(new_n8041_));
  NAND2_X1   g07848(.A1(new_n8041_), .A2(new_n8040_), .ZN(new_n8042_));
  XOR2_X1    g07849(.A1(new_n8042_), .A2(new_n8039_), .Z(new_n8043_));
  XOR2_X1    g07850(.A1(new_n8043_), .A2(new_n8038_), .Z(new_n8044_));
  NAND2_X1   g07851(.A1(new_n7928_), .A2(new_n7925_), .ZN(new_n8045_));
  NAND2_X1   g07852(.A1(new_n7929_), .A2(new_n7922_), .ZN(new_n8046_));
  NAND2_X1   g07853(.A1(new_n8046_), .A2(new_n8045_), .ZN(new_n8047_));
  NAND2_X1   g07854(.A1(new_n7590_), .A2(new_n243_), .ZN(new_n8048_));
  INV_X1     g07855(.I(new_n7644_), .ZN(new_n8049_));
  OAI22_X1   g07856(.A1(new_n370_), .A2(new_n8049_), .B1(new_n7959_), .B2(new_n318_), .ZN(new_n8050_));
  NAND2_X1   g07857(.A1(new_n8050_), .A2(new_n8048_), .ZN(new_n8051_));
  NAND3_X1   g07858(.A1(new_n8051_), .A2(\a[3] ), .A3(\a[63] ), .ZN(new_n8052_));
  AOI22_X1   g07859(.A1(\a[4] ), .A2(\a[62] ), .B1(\a[5] ), .B2(\a[61] ), .ZN(new_n8053_));
  NAND2_X1   g07860(.A1(new_n8051_), .A2(new_n8048_), .ZN(new_n8054_));
  OAI21_X1   g07861(.A1(new_n8053_), .A2(new_n8054_), .B(new_n8052_), .ZN(new_n8055_));
  NAND2_X1   g07862(.A1(new_n2105_), .A2(new_n3803_), .ZN(new_n8056_));
  OAI22_X1   g07863(.A1(new_n1816_), .A2(new_n4739_), .B1(new_n2189_), .B2(new_n4210_), .ZN(new_n8057_));
  NAND2_X1   g07864(.A1(new_n8057_), .A2(new_n8056_), .ZN(new_n8058_));
  NAND3_X1   g07865(.A1(new_n8058_), .A2(\a[27] ), .A3(\a[39] ), .ZN(new_n8059_));
  AOI22_X1   g07866(.A1(\a[28] ), .A2(\a[38] ), .B1(\a[29] ), .B2(\a[37] ), .ZN(new_n8060_));
  NAND2_X1   g07867(.A1(new_n8058_), .A2(new_n8056_), .ZN(new_n8061_));
  OAI21_X1   g07868(.A1(new_n8060_), .A2(new_n8061_), .B(new_n8059_), .ZN(new_n8062_));
  XOR2_X1    g07869(.A1(new_n8062_), .A2(new_n8055_), .Z(new_n8063_));
  NOR4_X1    g07870(.A1(new_n536_), .A2(new_n979_), .A3(new_n4312_), .A4(new_n5617_), .ZN(new_n8064_));
  INV_X1     g07871(.I(new_n8064_), .ZN(new_n8065_));
  NAND3_X1   g07872(.A1(new_n6385_), .A2(\a[19] ), .A3(\a[55] ), .ZN(new_n8066_));
  OAI21_X1   g07873(.A1(new_n619_), .A2(new_n6129_), .B(new_n8066_), .ZN(new_n8067_));
  NAND2_X1   g07874(.A1(new_n8067_), .A2(new_n8065_), .ZN(new_n8068_));
  NAND3_X1   g07875(.A1(new_n8068_), .A2(\a[11] ), .A3(\a[55] ), .ZN(new_n8069_));
  NOR2_X1    g07876(.A1(new_n8067_), .A2(new_n8064_), .ZN(new_n8070_));
  INV_X1     g07877(.I(new_n8070_), .ZN(new_n8071_));
  AOI22_X1   g07878(.A1(\a[12] ), .A2(\a[54] ), .B1(\a[19] ), .B2(\a[47] ), .ZN(new_n8072_));
  OAI21_X1   g07879(.A1(new_n8071_), .A2(new_n8072_), .B(new_n8069_), .ZN(new_n8073_));
  XNOR2_X1   g07880(.A1(new_n8063_), .A2(new_n8073_), .ZN(new_n8074_));
  NOR2_X1    g07881(.A1(new_n1357_), .A2(new_n6298_), .ZN(new_n8075_));
  INV_X1     g07882(.I(new_n8075_), .ZN(new_n8076_));
  INV_X1     g07883(.I(new_n2191_), .ZN(new_n8077_));
  NAND2_X1   g07884(.A1(\a[43] ), .A2(\a[57] ), .ZN(new_n8078_));
  OAI22_X1   g07885(.A1(new_n1529_), .A2(new_n4181_), .B1(new_n8077_), .B2(new_n8078_), .ZN(new_n8079_));
  OAI21_X1   g07886(.A1(new_n5059_), .A2(new_n8076_), .B(new_n8079_), .ZN(new_n8080_));
  NAND3_X1   g07887(.A1(new_n8080_), .A2(\a[23] ), .A3(\a[43] ), .ZN(new_n8081_));
  AOI22_X1   g07888(.A1(\a[9] ), .A2(\a[57] ), .B1(\a[24] ), .B2(\a[42] ), .ZN(new_n8082_));
  NOR2_X1    g07889(.A1(new_n5059_), .A2(new_n8076_), .ZN(new_n8083_));
  NOR2_X1    g07890(.A1(new_n8079_), .A2(new_n8083_), .ZN(new_n8084_));
  INV_X1     g07891(.I(new_n8084_), .ZN(new_n8085_));
  OAI21_X1   g07892(.A1(new_n8082_), .A2(new_n8085_), .B(new_n8081_), .ZN(new_n8086_));
  NAND2_X1   g07893(.A1(new_n1452_), .A2(new_n4703_), .ZN(new_n8087_));
  OAI22_X1   g07894(.A1(new_n1382_), .A2(new_n4430_), .B1(new_n2647_), .B2(new_n6101_), .ZN(new_n8088_));
  NAND2_X1   g07895(.A1(new_n8088_), .A2(new_n8087_), .ZN(new_n8089_));
  NAND3_X1   g07896(.A1(new_n8089_), .A2(\a[20] ), .A3(\a[46] ), .ZN(new_n8090_));
  AOI22_X1   g07897(.A1(\a[21] ), .A2(\a[45] ), .B1(\a[22] ), .B2(\a[44] ), .ZN(new_n8091_));
  NAND2_X1   g07898(.A1(new_n8089_), .A2(new_n8087_), .ZN(new_n8092_));
  OAI21_X1   g07899(.A1(new_n8091_), .A2(new_n8092_), .B(new_n8090_), .ZN(new_n8093_));
  XNOR2_X1   g07900(.A1(new_n8086_), .A2(new_n8093_), .ZN(new_n8094_));
  AOI22_X1   g07901(.A1(\a[25] ), .A2(\a[41] ), .B1(\a[26] ), .B2(\a[40] ), .ZN(new_n8095_));
  NOR2_X1    g07902(.A1(new_n417_), .A2(new_n5856_), .ZN(new_n8096_));
  INV_X1     g07903(.I(new_n8096_), .ZN(new_n8097_));
  NOR2_X1    g07904(.A1(new_n2177_), .A2(new_n5377_), .ZN(new_n8098_));
  NOR3_X1    g07905(.A1(new_n8098_), .A2(new_n8095_), .A3(new_n8097_), .ZN(new_n8099_));
  NOR2_X1    g07906(.A1(new_n8099_), .A2(new_n8098_), .ZN(new_n8100_));
  INV_X1     g07907(.I(new_n8100_), .ZN(new_n8101_));
  OAI22_X1   g07908(.A1(new_n8101_), .A2(new_n8095_), .B1(new_n8097_), .B2(new_n8099_), .ZN(new_n8102_));
  XOR2_X1    g07909(.A1(new_n8094_), .A2(new_n8102_), .Z(new_n8103_));
  AOI22_X1   g07910(.A1(\a[13] ), .A2(\a[53] ), .B1(\a[15] ), .B2(\a[51] ), .ZN(new_n8104_));
  INV_X1     g07911(.I(new_n8104_), .ZN(new_n8105_));
  NOR2_X1    g07912(.A1(new_n5683_), .A2(new_n836_), .ZN(new_n8106_));
  NOR2_X1    g07913(.A1(new_n884_), .A2(new_n4596_), .ZN(new_n8107_));
  AOI21_X1   g07914(.A1(new_n8105_), .A2(new_n8107_), .B(new_n8106_), .ZN(new_n8108_));
  INV_X1     g07915(.I(new_n8108_), .ZN(new_n8109_));
  OAI21_X1   g07916(.A1(new_n8106_), .A2(new_n8104_), .B(new_n8107_), .ZN(new_n8110_));
  OAI21_X1   g07917(.A1(new_n8109_), .A2(new_n8104_), .B(new_n8110_), .ZN(new_n8111_));
  AOI22_X1   g07918(.A1(\a[30] ), .A2(\a[36] ), .B1(\a[31] ), .B2(\a[35] ), .ZN(new_n8112_));
  INV_X1     g07919(.I(new_n8112_), .ZN(new_n8113_));
  NOR2_X1    g07920(.A1(new_n2438_), .A2(new_n3405_), .ZN(new_n8114_));
  NOR2_X1    g07921(.A1(new_n759_), .A2(new_n5175_), .ZN(new_n8115_));
  AOI21_X1   g07922(.A1(new_n8113_), .A2(new_n8115_), .B(new_n8114_), .ZN(new_n8116_));
  INV_X1     g07923(.I(new_n8116_), .ZN(new_n8117_));
  OAI21_X1   g07924(.A1(new_n8114_), .A2(new_n8112_), .B(new_n8115_), .ZN(new_n8118_));
  OAI21_X1   g07925(.A1(new_n8117_), .A2(new_n8112_), .B(new_n8118_), .ZN(new_n8119_));
  XNOR2_X1   g07926(.A1(new_n8119_), .A2(new_n8111_), .ZN(new_n8120_));
  AOI21_X1   g07927(.A1(\a[16] ), .A2(\a[50] ), .B(new_n6340_), .ZN(new_n8121_));
  NOR2_X1    g07928(.A1(new_n1428_), .A2(new_n5155_), .ZN(new_n8122_));
  NOR3_X1    g07929(.A1(new_n8122_), .A2(new_n3375_), .A3(new_n8121_), .ZN(new_n8123_));
  NOR2_X1    g07930(.A1(new_n8123_), .A2(new_n8122_), .ZN(new_n8124_));
  INV_X1     g07931(.I(new_n8124_), .ZN(new_n8125_));
  OAI22_X1   g07932(.A1(new_n8125_), .A2(new_n8121_), .B1(new_n3375_), .B2(new_n8123_), .ZN(new_n8126_));
  XOR2_X1    g07933(.A1(new_n8120_), .A2(new_n8126_), .Z(new_n8127_));
  XNOR2_X1   g07934(.A1(new_n8103_), .A2(new_n8127_), .ZN(new_n8128_));
  XOR2_X1    g07935(.A1(new_n8128_), .A2(new_n8074_), .Z(new_n8129_));
  XOR2_X1    g07936(.A1(new_n8047_), .A2(new_n8129_), .Z(new_n8130_));
  XNOR2_X1   g07937(.A1(new_n8130_), .A2(new_n8044_), .ZN(new_n8131_));
  NAND2_X1   g07938(.A1(new_n7906_), .A2(new_n7930_), .ZN(new_n8132_));
  NAND2_X1   g07939(.A1(new_n7931_), .A2(new_n7903_), .ZN(new_n8133_));
  NAND2_X1   g07940(.A1(new_n8133_), .A2(new_n8132_), .ZN(new_n8134_));
  NAND2_X1   g07941(.A1(new_n7829_), .A2(new_n7826_), .ZN(new_n8135_));
  NAND2_X1   g07942(.A1(new_n7830_), .A2(new_n7844_), .ZN(new_n8136_));
  NAND2_X1   g07943(.A1(new_n8136_), .A2(new_n8135_), .ZN(new_n8137_));
  XNOR2_X1   g07944(.A1(new_n8134_), .A2(new_n8137_), .ZN(new_n8138_));
  XOR2_X1    g07945(.A1(new_n8138_), .A2(new_n8131_), .Z(new_n8139_));
  XNOR2_X1   g07946(.A1(new_n8027_), .A2(new_n8139_), .ZN(new_n8140_));
  INV_X1     g07947(.I(new_n8140_), .ZN(new_n8141_));
  NOR2_X1    g07948(.A1(new_n8141_), .A2(new_n7952_), .ZN(new_n8142_));
  INV_X1     g07949(.I(new_n8142_), .ZN(new_n8143_));
  NOR2_X1    g07950(.A1(new_n8140_), .A2(new_n7951_), .ZN(new_n8144_));
  INV_X1     g07951(.I(new_n8144_), .ZN(new_n8145_));
  NAND2_X1   g07952(.A1(new_n8143_), .A2(new_n8145_), .ZN(new_n8146_));
  XOR2_X1    g07953(.A1(new_n7950_), .A2(new_n8146_), .Z(\asquared[67] ));
  OAI21_X1   g07954(.A1(new_n7949_), .A2(new_n7946_), .B(new_n8143_), .ZN(new_n8148_));
  NAND2_X1   g07955(.A1(new_n8148_), .A2(new_n8145_), .ZN(new_n8149_));
  NAND2_X1   g07956(.A1(new_n8026_), .A2(new_n8023_), .ZN(new_n8150_));
  NAND2_X1   g07957(.A1(new_n8027_), .A2(new_n8139_), .ZN(new_n8151_));
  NAND2_X1   g07958(.A1(new_n8151_), .A2(new_n8150_), .ZN(new_n8152_));
  NAND2_X1   g07959(.A1(new_n8134_), .A2(new_n8137_), .ZN(new_n8153_));
  OAI21_X1   g07960(.A1(new_n8138_), .A2(new_n8131_), .B(new_n8153_), .ZN(new_n8154_));
  NAND2_X1   g07961(.A1(new_n8033_), .A2(new_n8035_), .ZN(new_n8155_));
  NAND2_X1   g07962(.A1(new_n8036_), .A2(new_n8030_), .ZN(new_n8156_));
  NAND2_X1   g07963(.A1(new_n8156_), .A2(new_n8155_), .ZN(new_n8157_));
  XOR2_X1    g07964(.A1(new_n8070_), .A2(new_n8108_), .Z(new_n8158_));
  NAND2_X1   g07965(.A1(new_n6385_), .A2(new_n7748_), .ZN(new_n8159_));
  NOR4_X1    g07966(.A1(new_n417_), .A2(new_n1043_), .A3(new_n4312_), .A4(new_n6298_), .ZN(new_n8160_));
  INV_X1     g07967(.I(new_n6494_), .ZN(new_n8161_));
  NOR2_X1    g07968(.A1(new_n1264_), .A2(new_n8161_), .ZN(new_n8162_));
  OAI21_X1   g07969(.A1(new_n8162_), .A2(new_n8160_), .B(new_n8159_), .ZN(new_n8163_));
  NAND3_X1   g07970(.A1(new_n8163_), .A2(\a[10] ), .A3(\a[57] ), .ZN(new_n8164_));
  AOI22_X1   g07971(.A1(\a[11] ), .A2(\a[56] ), .B1(\a[20] ), .B2(\a[47] ), .ZN(new_n8165_));
  NAND2_X1   g07972(.A1(new_n8163_), .A2(new_n8159_), .ZN(new_n8166_));
  OAI21_X1   g07973(.A1(new_n8165_), .A2(new_n8166_), .B(new_n8164_), .ZN(new_n8167_));
  XOR2_X1    g07974(.A1(new_n8158_), .A2(new_n8167_), .Z(new_n8168_));
  NAND2_X1   g07975(.A1(new_n8119_), .A2(new_n8111_), .ZN(new_n8169_));
  INV_X1     g07976(.I(new_n8126_), .ZN(new_n8170_));
  OAI21_X1   g07977(.A1(new_n8120_), .A2(new_n8170_), .B(new_n8169_), .ZN(new_n8171_));
  XOR2_X1    g07978(.A1(new_n8171_), .A2(new_n8168_), .Z(new_n8172_));
  XOR2_X1    g07979(.A1(new_n8157_), .A2(new_n8172_), .Z(new_n8173_));
  OR2_X2     g07980(.A1(new_n8103_), .A2(new_n8127_), .Z(new_n8174_));
  OAI21_X1   g07981(.A1(new_n8128_), .A2(new_n8074_), .B(new_n8174_), .ZN(new_n8175_));
  INV_X1     g07982(.I(new_n7971_), .ZN(new_n8176_));
  NAND2_X1   g07983(.A1(new_n8176_), .A2(new_n7974_), .ZN(new_n8177_));
  INV_X1     g07984(.I(new_n7975_), .ZN(new_n8178_));
  NAND2_X1   g07985(.A1(new_n8178_), .A2(new_n7958_), .ZN(new_n8179_));
  NAND2_X1   g07986(.A1(new_n8179_), .A2(new_n8177_), .ZN(new_n8180_));
  XOR2_X1    g07987(.A1(new_n8180_), .A2(new_n8175_), .Z(new_n8181_));
  XOR2_X1    g07988(.A1(new_n8181_), .A2(new_n8173_), .Z(new_n8182_));
  INV_X1     g07989(.I(new_n7976_), .ZN(new_n8183_));
  NOR2_X1    g07990(.A1(new_n8183_), .A2(new_n7985_), .ZN(new_n8184_));
  NOR2_X1    g07991(.A1(new_n7989_), .A2(new_n8184_), .ZN(new_n8185_));
  OAI21_X1   g07992(.A1(new_n7915_), .A2(new_n7920_), .B(new_n8042_), .ZN(new_n8186_));
  OAI21_X1   g07993(.A1(new_n8043_), .A2(new_n8038_), .B(new_n8186_), .ZN(new_n8187_));
  NAND2_X1   g07994(.A1(new_n8062_), .A2(new_n8055_), .ZN(new_n8188_));
  NAND2_X1   g07995(.A1(new_n8063_), .A2(new_n8073_), .ZN(new_n8189_));
  NAND2_X1   g07996(.A1(new_n8189_), .A2(new_n8188_), .ZN(new_n8190_));
  NAND2_X1   g07997(.A1(new_n8086_), .A2(new_n8093_), .ZN(new_n8191_));
  INV_X1     g07998(.I(new_n8102_), .ZN(new_n8192_));
  OAI21_X1   g07999(.A1(new_n8094_), .A2(new_n8192_), .B(new_n8191_), .ZN(new_n8193_));
  NAND2_X1   g08000(.A1(new_n7961_), .A2(new_n7771_), .ZN(new_n8194_));
  NAND2_X1   g08001(.A1(new_n7962_), .A2(new_n7970_), .ZN(new_n8195_));
  NAND2_X1   g08002(.A1(new_n8195_), .A2(new_n8194_), .ZN(new_n8196_));
  XOR2_X1    g08003(.A1(new_n8193_), .A2(new_n8196_), .Z(new_n8197_));
  XOR2_X1    g08004(.A1(new_n8197_), .A2(new_n8190_), .Z(new_n8198_));
  XOR2_X1    g08005(.A1(new_n8054_), .A2(new_n7969_), .Z(new_n8199_));
  XOR2_X1    g08006(.A1(new_n8199_), .A2(new_n8061_), .Z(new_n8200_));
  XOR2_X1    g08007(.A1(new_n8100_), .A2(new_n8084_), .Z(new_n8201_));
  XOR2_X1    g08008(.A1(new_n8201_), .A2(new_n8092_), .Z(new_n8202_));
  NOR2_X1    g08009(.A1(new_n367_), .A2(new_n6897_), .ZN(new_n8203_));
  XNOR2_X1   g08010(.A1(new_n8124_), .A2(new_n8203_), .ZN(new_n8204_));
  XOR2_X1    g08011(.A1(new_n8204_), .A2(new_n8117_), .Z(new_n8205_));
  XOR2_X1    g08012(.A1(new_n8205_), .A2(new_n8202_), .Z(new_n8206_));
  XNOR2_X1   g08013(.A1(new_n8206_), .A2(new_n8200_), .ZN(new_n8207_));
  XNOR2_X1   g08014(.A1(new_n8198_), .A2(new_n8207_), .ZN(new_n8208_));
  NOR2_X1    g08015(.A1(new_n8187_), .A2(new_n8208_), .ZN(new_n8209_));
  NAND2_X1   g08016(.A1(new_n8187_), .A2(new_n8208_), .ZN(new_n8210_));
  INV_X1     g08017(.I(new_n8210_), .ZN(new_n8211_));
  NOR2_X1    g08018(.A1(new_n8211_), .A2(new_n8209_), .ZN(new_n8212_));
  INV_X1     g08019(.I(new_n8212_), .ZN(new_n8213_));
  XOR2_X1    g08020(.A1(new_n8185_), .A2(new_n8213_), .Z(new_n8214_));
  NOR2_X1    g08021(.A1(new_n8214_), .A2(new_n8182_), .ZN(new_n8215_));
  NAND2_X1   g08022(.A1(new_n8214_), .A2(new_n8182_), .ZN(new_n8216_));
  INV_X1     g08023(.I(new_n8216_), .ZN(new_n8217_));
  NOR2_X1    g08024(.A1(new_n8217_), .A2(new_n8215_), .ZN(new_n8218_));
  XOR2_X1    g08025(.A1(new_n8154_), .A2(new_n8218_), .Z(new_n8219_));
  INV_X1     g08026(.I(new_n8219_), .ZN(new_n8220_));
  NAND2_X1   g08027(.A1(new_n7993_), .A2(new_n8021_), .ZN(new_n8221_));
  OAI21_X1   g08028(.A1(new_n8022_), .A2(new_n7991_), .B(new_n8221_), .ZN(new_n8222_));
  NAND2_X1   g08029(.A1(new_n8047_), .A2(new_n8129_), .ZN(new_n8223_));
  NAND2_X1   g08030(.A1(new_n8130_), .A2(new_n8044_), .ZN(new_n8224_));
  NAND2_X1   g08031(.A1(new_n8224_), .A2(new_n8223_), .ZN(new_n8225_));
  XNOR2_X1   g08032(.A1(new_n8222_), .A2(new_n8225_), .ZN(new_n8226_));
  NAND2_X1   g08033(.A1(new_n7977_), .A2(new_n7872_), .ZN(new_n8227_));
  OAI21_X1   g08034(.A1(new_n7780_), .A2(new_n7796_), .B(new_n8227_), .ZN(new_n8228_));
  NAND2_X1   g08035(.A1(new_n7753_), .A2(new_n7862_), .ZN(new_n8229_));
  NAND2_X1   g08036(.A1(new_n7997_), .A2(new_n7762_), .ZN(new_n8230_));
  NAND2_X1   g08037(.A1(new_n8230_), .A2(new_n8229_), .ZN(new_n8231_));
  NAND2_X1   g08038(.A1(new_n7979_), .A2(new_n7788_), .ZN(new_n8232_));
  OAI21_X1   g08039(.A1(new_n7807_), .A2(new_n7816_), .B(new_n8232_), .ZN(new_n8233_));
  XOR2_X1    g08040(.A1(new_n8233_), .A2(new_n8231_), .Z(new_n8234_));
  XOR2_X1    g08041(.A1(new_n8234_), .A2(new_n8228_), .Z(new_n8235_));
  NOR2_X1    g08042(.A1(new_n8007_), .A2(new_n8002_), .ZN(new_n8236_));
  INV_X1     g08043(.I(new_n8236_), .ZN(new_n8237_));
  NAND2_X1   g08044(.A1(new_n7983_), .A2(new_n7980_), .ZN(new_n8238_));
  NAND2_X1   g08045(.A1(new_n7984_), .A2(new_n7978_), .ZN(new_n8239_));
  NAND2_X1   g08046(.A1(new_n8239_), .A2(new_n8238_), .ZN(new_n8240_));
  NOR2_X1    g08047(.A1(new_n8237_), .A2(new_n8240_), .ZN(new_n8241_));
  NAND2_X1   g08048(.A1(new_n8237_), .A2(new_n8240_), .ZN(new_n8242_));
  INV_X1     g08049(.I(new_n8242_), .ZN(new_n8243_));
  NOR2_X1    g08050(.A1(new_n8243_), .A2(new_n8241_), .ZN(new_n8244_));
  NAND2_X1   g08051(.A1(new_n8244_), .A2(new_n8235_), .ZN(new_n8245_));
  INV_X1     g08052(.I(new_n8245_), .ZN(new_n8246_));
  NOR2_X1    g08053(.A1(new_n8244_), .A2(new_n8235_), .ZN(new_n8247_));
  NOR2_X1    g08054(.A1(new_n8246_), .A2(new_n8247_), .ZN(new_n8248_));
  NOR2_X1    g08055(.A1(new_n8019_), .A2(new_n8016_), .ZN(new_n8249_));
  NOR2_X1    g08056(.A1(new_n4596_), .A2(new_n5425_), .ZN(new_n8250_));
  AOI22_X1   g08057(.A1(\a[14] ), .A2(new_n8250_), .B1(new_n4902_), .B2(\a[17] ), .ZN(new_n8251_));
  NOR4_X1    g08058(.A1(new_n759_), .A2(new_n1023_), .A3(new_n4901_), .A4(new_n5425_), .ZN(new_n8252_));
  NOR3_X1    g08059(.A1(new_n8251_), .A2(new_n979_), .A3(new_n8252_), .ZN(new_n8253_));
  NAND2_X1   g08060(.A1(\a[19] ), .A2(\a[48] ), .ZN(new_n8254_));
  NOR2_X1    g08061(.A1(new_n759_), .A2(new_n5425_), .ZN(new_n8255_));
  NOR2_X1    g08062(.A1(new_n8253_), .A2(new_n8252_), .ZN(new_n8256_));
  OAI21_X1   g08063(.A1(new_n5900_), .A2(new_n8255_), .B(new_n8256_), .ZN(new_n8257_));
  OAI21_X1   g08064(.A1(new_n8253_), .A2(new_n8254_), .B(new_n8257_), .ZN(new_n8258_));
  NAND4_X1   g08065(.A1(\a[21] ), .A2(\a[25] ), .A3(\a[42] ), .A4(\a[46] ), .ZN(new_n8259_));
  NAND2_X1   g08066(.A1(new_n2176_), .A2(new_n4372_), .ZN(new_n8260_));
  NOR4_X1    g08067(.A1(new_n1220_), .A2(new_n1566_), .A3(new_n3327_), .A4(new_n4178_), .ZN(new_n8261_));
  AOI21_X1   g08068(.A1(new_n8260_), .A2(new_n8259_), .B(new_n8261_), .ZN(new_n8262_));
  NAND2_X1   g08069(.A1(\a[25] ), .A2(\a[42] ), .ZN(new_n8263_));
  AOI22_X1   g08070(.A1(\a[21] ), .A2(\a[46] ), .B1(\a[26] ), .B2(\a[41] ), .ZN(new_n8264_));
  NOR2_X1    g08071(.A1(new_n8262_), .A2(new_n8261_), .ZN(new_n8265_));
  INV_X1     g08072(.I(new_n8265_), .ZN(new_n8266_));
  OAI22_X1   g08073(.A1(new_n8266_), .A2(new_n8264_), .B1(new_n8262_), .B2(new_n8263_), .ZN(new_n8267_));
  XNOR2_X1   g08074(.A1(new_n8258_), .A2(new_n8267_), .ZN(new_n8268_));
  AOI22_X1   g08075(.A1(\a[27] ), .A2(\a[40] ), .B1(\a[28] ), .B2(\a[39] ), .ZN(new_n8269_));
  NOR2_X1    g08076(.A1(new_n290_), .A2(new_n7643_), .ZN(new_n8270_));
  INV_X1     g08077(.I(new_n8270_), .ZN(new_n8271_));
  NOR2_X1    g08078(.A1(new_n2189_), .A2(new_n3551_), .ZN(new_n8272_));
  NOR3_X1    g08079(.A1(new_n8272_), .A2(new_n8269_), .A3(new_n8271_), .ZN(new_n8273_));
  NOR2_X1    g08080(.A1(new_n8273_), .A2(new_n8272_), .ZN(new_n8274_));
  INV_X1     g08081(.I(new_n8274_), .ZN(new_n8275_));
  OAI22_X1   g08082(.A1(new_n8275_), .A2(new_n8269_), .B1(new_n8271_), .B2(new_n8273_), .ZN(new_n8276_));
  INV_X1     g08083(.I(new_n8276_), .ZN(new_n8277_));
  XOR2_X1    g08084(.A1(new_n8268_), .A2(new_n8277_), .Z(new_n8278_));
  NAND2_X1   g08085(.A1(new_n467_), .A2(new_n7205_), .ZN(new_n8279_));
  OAI22_X1   g08086(.A1(new_n415_), .A2(new_n7452_), .B1(new_n7801_), .B2(new_n773_), .ZN(new_n8280_));
  NAND2_X1   g08087(.A1(new_n8280_), .A2(new_n8279_), .ZN(new_n8281_));
  NAND3_X1   g08088(.A1(new_n8281_), .A2(\a[7] ), .A3(\a[60] ), .ZN(new_n8282_));
  AOI22_X1   g08089(.A1(\a[8] ), .A2(\a[59] ), .B1(\a[9] ), .B2(\a[58] ), .ZN(new_n8283_));
  NAND2_X1   g08090(.A1(new_n8281_), .A2(new_n8279_), .ZN(new_n8284_));
  OAI21_X1   g08091(.A1(new_n8283_), .A2(new_n8284_), .B(new_n8282_), .ZN(new_n8285_));
  NAND2_X1   g08092(.A1(new_n1528_), .A2(new_n4342_), .ZN(new_n8286_));
  OAI22_X1   g08093(.A1(new_n2385_), .A2(new_n4704_), .B1(new_n1880_), .B2(new_n4034_), .ZN(new_n8287_));
  NAND2_X1   g08094(.A1(new_n8287_), .A2(new_n8286_), .ZN(new_n8288_));
  NAND3_X1   g08095(.A1(new_n8288_), .A2(\a[22] ), .A3(\a[45] ), .ZN(new_n8289_));
  AOI22_X1   g08096(.A1(\a[23] ), .A2(\a[44] ), .B1(\a[24] ), .B2(\a[43] ), .ZN(new_n8290_));
  NAND2_X1   g08097(.A1(new_n8288_), .A2(new_n8286_), .ZN(new_n8291_));
  OAI21_X1   g08098(.A1(new_n8290_), .A2(new_n8291_), .B(new_n8289_), .ZN(new_n8292_));
  XOR2_X1    g08099(.A1(new_n8292_), .A2(new_n8285_), .Z(new_n8293_));
  NAND4_X1   g08100(.A1(\a[15] ), .A2(\a[30] ), .A3(\a[37] ), .A4(\a[52] ), .ZN(new_n8294_));
  NAND2_X1   g08101(.A1(new_n5524_), .A2(new_n1288_), .ZN(new_n8295_));
  NOR4_X1    g08102(.A1(new_n742_), .A2(new_n2030_), .A3(new_n2752_), .A4(new_n5135_), .ZN(new_n8296_));
  AOI21_X1   g08103(.A1(new_n8295_), .A2(new_n8294_), .B(new_n8296_), .ZN(new_n8297_));
  NAND2_X1   g08104(.A1(\a[15] ), .A2(\a[52] ), .ZN(new_n8298_));
  AOI22_X1   g08105(.A1(\a[16] ), .A2(\a[51] ), .B1(\a[30] ), .B2(\a[37] ), .ZN(new_n8299_));
  NOR2_X1    g08106(.A1(new_n8297_), .A2(new_n8296_), .ZN(new_n8300_));
  INV_X1     g08107(.I(new_n8300_), .ZN(new_n8301_));
  OAI22_X1   g08108(.A1(new_n8301_), .A2(new_n8299_), .B1(new_n8297_), .B2(new_n8298_), .ZN(new_n8302_));
  XNOR2_X1   g08109(.A1(new_n8293_), .A2(new_n8302_), .ZN(new_n8303_));
  AOI21_X1   g08110(.A1(\a[5] ), .A2(\a[62] ), .B(\a[34] ), .ZN(new_n8304_));
  NOR2_X1    g08111(.A1(new_n884_), .A2(new_n4702_), .ZN(new_n8305_));
  INV_X1     g08112(.I(new_n8305_), .ZN(new_n8306_));
  NOR2_X1    g08113(.A1(new_n4847_), .A2(new_n7144_), .ZN(new_n8307_));
  NOR3_X1    g08114(.A1(new_n8307_), .A2(new_n8304_), .A3(new_n8306_), .ZN(new_n8308_));
  NOR2_X1    g08115(.A1(new_n8308_), .A2(new_n8307_), .ZN(new_n8309_));
  INV_X1     g08116(.I(new_n8309_), .ZN(new_n8310_));
  OAI22_X1   g08117(.A1(new_n8310_), .A2(new_n8304_), .B1(new_n8306_), .B2(new_n8308_), .ZN(new_n8311_));
  OAI22_X1   g08118(.A1(new_n3833_), .A2(new_n3405_), .B1(new_n3932_), .B2(new_n3586_), .ZN(new_n8312_));
  OAI21_X1   g08119(.A1(new_n2637_), .A2(new_n2746_), .B(new_n8312_), .ZN(new_n8313_));
  NAND2_X1   g08120(.A1(new_n8313_), .A2(new_n3585_), .ZN(new_n8314_));
  AOI21_X1   g08121(.A1(new_n2636_), .A2(new_n2745_), .B(new_n8312_), .ZN(new_n8315_));
  OAI21_X1   g08122(.A1(new_n3577_), .A2(new_n5633_), .B(new_n8315_), .ZN(new_n8316_));
  NAND2_X1   g08123(.A1(new_n8316_), .A2(new_n8314_), .ZN(new_n8317_));
  XNOR2_X1   g08124(.A1(new_n8317_), .A2(new_n8311_), .ZN(new_n8318_));
  AOI22_X1   g08125(.A1(\a[12] ), .A2(\a[55] ), .B1(\a[13] ), .B2(\a[54] ), .ZN(new_n8319_));
  NOR2_X1    g08126(.A1(new_n1814_), .A2(new_n2914_), .ZN(new_n8320_));
  INV_X1     g08127(.I(new_n8320_), .ZN(new_n8321_));
  NOR2_X1    g08128(.A1(new_n1265_), .A2(new_n6129_), .ZN(new_n8322_));
  NOR3_X1    g08129(.A1(new_n8322_), .A2(new_n8319_), .A3(new_n8321_), .ZN(new_n8323_));
  NOR2_X1    g08130(.A1(new_n8323_), .A2(new_n8322_), .ZN(new_n8324_));
  INV_X1     g08131(.I(new_n8324_), .ZN(new_n8325_));
  OAI22_X1   g08132(.A1(new_n8325_), .A2(new_n8319_), .B1(new_n8321_), .B2(new_n8323_), .ZN(new_n8326_));
  XOR2_X1    g08133(.A1(new_n8318_), .A2(new_n8326_), .Z(new_n8327_));
  XOR2_X1    g08134(.A1(new_n8327_), .A2(new_n8303_), .Z(new_n8328_));
  XOR2_X1    g08135(.A1(new_n8328_), .A2(new_n8278_), .Z(new_n8329_));
  INV_X1     g08136(.I(new_n8329_), .ZN(new_n8330_));
  XOR2_X1    g08137(.A1(new_n8249_), .A2(new_n8330_), .Z(new_n8331_));
  XNOR2_X1   g08138(.A1(new_n8331_), .A2(new_n8248_), .ZN(new_n8332_));
  OR2_X2     g08139(.A1(new_n8226_), .A2(new_n8332_), .Z(new_n8333_));
  NAND2_X1   g08140(.A1(new_n8226_), .A2(new_n8332_), .ZN(new_n8334_));
  NAND3_X1   g08141(.A1(new_n8219_), .A2(new_n8333_), .A3(new_n8334_), .ZN(new_n8335_));
  INV_X1     g08142(.I(new_n8335_), .ZN(new_n8336_));
  NAND2_X1   g08143(.A1(new_n8333_), .A2(new_n8334_), .ZN(new_n8337_));
  AOI21_X1   g08144(.A1(new_n8220_), .A2(new_n8337_), .B(new_n8336_), .ZN(new_n8338_));
  NAND2_X1   g08145(.A1(new_n8338_), .A2(new_n8152_), .ZN(new_n8339_));
  INV_X1     g08146(.I(new_n8339_), .ZN(new_n8340_));
  NOR2_X1    g08147(.A1(new_n8338_), .A2(new_n8152_), .ZN(new_n8341_));
  NOR2_X1    g08148(.A1(new_n8340_), .A2(new_n8341_), .ZN(new_n8342_));
  XOR2_X1    g08149(.A1(new_n8149_), .A2(new_n8342_), .Z(\asquared[68] ));
  AOI21_X1   g08150(.A1(new_n8148_), .A2(new_n8145_), .B(new_n8341_), .ZN(new_n8344_));
  NOR2_X1    g08151(.A1(new_n8344_), .A2(new_n8340_), .ZN(new_n8345_));
  NOR2_X1    g08152(.A1(new_n8185_), .A2(new_n8213_), .ZN(new_n8346_));
  NOR2_X1    g08153(.A1(new_n8217_), .A2(new_n8346_), .ZN(new_n8347_));
  NAND2_X1   g08154(.A1(new_n8331_), .A2(new_n8248_), .ZN(new_n8348_));
  OAI21_X1   g08155(.A1(new_n8249_), .A2(new_n8330_), .B(new_n8348_), .ZN(new_n8349_));
  NAND2_X1   g08156(.A1(new_n8180_), .A2(new_n8175_), .ZN(new_n8350_));
  NAND2_X1   g08157(.A1(new_n8181_), .A2(new_n8173_), .ZN(new_n8351_));
  NAND2_X1   g08158(.A1(new_n8351_), .A2(new_n8350_), .ZN(new_n8352_));
  NAND2_X1   g08159(.A1(new_n8171_), .A2(new_n8168_), .ZN(new_n8353_));
  NAND2_X1   g08160(.A1(new_n8157_), .A2(new_n8172_), .ZN(new_n8354_));
  NAND2_X1   g08161(.A1(new_n8354_), .A2(new_n8353_), .ZN(new_n8355_));
  NAND2_X1   g08162(.A1(new_n8193_), .A2(new_n8196_), .ZN(new_n8356_));
  NAND2_X1   g08163(.A1(new_n8197_), .A2(new_n8190_), .ZN(new_n8357_));
  NAND2_X1   g08164(.A1(new_n8357_), .A2(new_n8356_), .ZN(new_n8358_));
  NAND2_X1   g08165(.A1(new_n8205_), .A2(new_n8202_), .ZN(new_n8359_));
  NAND2_X1   g08166(.A1(new_n8206_), .A2(new_n8200_), .ZN(new_n8360_));
  NAND2_X1   g08167(.A1(new_n8360_), .A2(new_n8359_), .ZN(new_n8361_));
  XOR2_X1    g08168(.A1(new_n8358_), .A2(new_n8361_), .Z(new_n8362_));
  XOR2_X1    g08169(.A1(new_n8362_), .A2(new_n8355_), .Z(new_n8363_));
  OAI22_X1   g08170(.A1(new_n1063_), .A2(new_n7204_), .B1(new_n7206_), .B2(new_n539_), .ZN(new_n8364_));
  OAI21_X1   g08171(.A1(new_n1264_), .A2(new_n6804_), .B(new_n8364_), .ZN(new_n8365_));
  NAND3_X1   g08172(.A1(new_n8365_), .A2(\a[9] ), .A3(\a[59] ), .ZN(new_n8366_));
  AOI22_X1   g08173(.A1(\a[10] ), .A2(\a[58] ), .B1(\a[11] ), .B2(\a[57] ), .ZN(new_n8367_));
  NOR2_X1    g08174(.A1(new_n1264_), .A2(new_n6804_), .ZN(new_n8368_));
  NOR2_X1    g08175(.A1(new_n8364_), .A2(new_n8368_), .ZN(new_n8369_));
  INV_X1     g08176(.I(new_n8369_), .ZN(new_n8370_));
  OAI21_X1   g08177(.A1(new_n8367_), .A2(new_n8370_), .B(new_n8366_), .ZN(new_n8371_));
  NAND2_X1   g08178(.A1(new_n2105_), .A2(new_n3550_), .ZN(new_n8372_));
  OAI22_X1   g08179(.A1(new_n1816_), .A2(new_n3329_), .B1(new_n2189_), .B2(new_n5377_), .ZN(new_n8373_));
  NAND2_X1   g08180(.A1(new_n8373_), .A2(new_n8372_), .ZN(new_n8374_));
  NAND3_X1   g08181(.A1(new_n8374_), .A2(\a[27] ), .A3(\a[41] ), .ZN(new_n8375_));
  AOI22_X1   g08182(.A1(\a[28] ), .A2(\a[40] ), .B1(\a[29] ), .B2(\a[39] ), .ZN(new_n8376_));
  NAND2_X1   g08183(.A1(new_n8374_), .A2(new_n8372_), .ZN(new_n8377_));
  OAI21_X1   g08184(.A1(new_n8376_), .A2(new_n8377_), .B(new_n8375_), .ZN(new_n8378_));
  XNOR2_X1   g08185(.A1(new_n8371_), .A2(new_n8378_), .ZN(new_n8379_));
  AOI22_X1   g08186(.A1(\a[5] ), .A2(\a[63] ), .B1(\a[6] ), .B2(\a[62] ), .ZN(new_n8380_));
  NOR2_X1    g08187(.A1(new_n1220_), .A2(new_n4312_), .ZN(new_n8381_));
  INV_X1     g08188(.I(new_n8381_), .ZN(new_n8382_));
  NOR2_X1    g08189(.A1(new_n8049_), .A2(new_n371_), .ZN(new_n8383_));
  NOR3_X1    g08190(.A1(new_n8383_), .A2(new_n8380_), .A3(new_n8382_), .ZN(new_n8384_));
  NOR2_X1    g08191(.A1(new_n8384_), .A2(new_n8383_), .ZN(new_n8385_));
  INV_X1     g08192(.I(new_n8385_), .ZN(new_n8386_));
  OAI22_X1   g08193(.A1(new_n8386_), .A2(new_n8380_), .B1(new_n8382_), .B2(new_n8384_), .ZN(new_n8387_));
  INV_X1     g08194(.I(new_n8387_), .ZN(new_n8388_));
  XOR2_X1    g08195(.A1(new_n8379_), .A2(new_n8388_), .Z(new_n8389_));
  AOI22_X1   g08196(.A1(\a[18] ), .A2(\a[50] ), .B1(\a[19] ), .B2(\a[49] ), .ZN(new_n8390_));
  INV_X1     g08197(.I(new_n8390_), .ZN(new_n8391_));
  NOR2_X1    g08198(.A1(new_n5155_), .A2(new_n1092_), .ZN(new_n8392_));
  OR3_X2     g08199(.A1(new_n8392_), .A2(new_n2526_), .A3(new_n8390_), .Z(new_n8393_));
  AOI21_X1   g08200(.A1(new_n2525_), .A2(new_n8391_), .B(new_n8392_), .ZN(new_n8394_));
  AOI22_X1   g08201(.A1(new_n8393_), .A2(new_n2525_), .B1(new_n8394_), .B2(new_n8391_), .ZN(new_n8395_));
  INV_X1     g08202(.I(new_n8395_), .ZN(new_n8396_));
  NOR2_X1    g08203(.A1(new_n3038_), .A2(new_n3833_), .ZN(new_n8397_));
  NOR2_X1    g08204(.A1(new_n2202_), .A2(new_n2916_), .ZN(new_n8398_));
  NOR2_X1    g08205(.A1(new_n2438_), .A2(new_n6140_), .ZN(new_n8399_));
  NOR2_X1    g08206(.A1(new_n8398_), .A2(new_n8399_), .ZN(new_n8400_));
  NOR2_X1    g08207(.A1(new_n8400_), .A2(new_n8397_), .ZN(new_n8401_));
  NAND2_X1   g08208(.A1(\a[30] ), .A2(\a[38] ), .ZN(new_n8402_));
  AOI22_X1   g08209(.A1(\a[31] ), .A2(\a[37] ), .B1(\a[32] ), .B2(\a[36] ), .ZN(new_n8403_));
  NOR2_X1    g08210(.A1(new_n8401_), .A2(new_n8397_), .ZN(new_n8404_));
  INV_X1     g08211(.I(new_n8404_), .ZN(new_n8405_));
  OAI22_X1   g08212(.A1(new_n8405_), .A2(new_n8403_), .B1(new_n8401_), .B2(new_n8402_), .ZN(new_n8406_));
  XOR2_X1    g08213(.A1(new_n8406_), .A2(new_n8396_), .Z(new_n8407_));
  NOR2_X1    g08214(.A1(new_n536_), .A2(new_n5856_), .ZN(new_n8408_));
  INV_X1     g08215(.I(new_n8408_), .ZN(new_n8409_));
  NOR3_X1    g08216(.A1(new_n6790_), .A2(new_n597_), .A3(new_n5680_), .ZN(new_n8410_));
  AOI22_X1   g08217(.A1(new_n763_), .A2(new_n7184_), .B1(new_n6113_), .B2(new_n8408_), .ZN(new_n8411_));
  NOR2_X1    g08218(.A1(new_n8410_), .A2(new_n8411_), .ZN(new_n8412_));
  AOI21_X1   g08219(.A1(\a[13] ), .A2(\a[55] ), .B(new_n6113_), .ZN(new_n8413_));
  INV_X1     g08220(.I(new_n8410_), .ZN(new_n8414_));
  NAND2_X1   g08221(.A1(new_n8414_), .A2(new_n8411_), .ZN(new_n8415_));
  OAI22_X1   g08222(.A1(new_n8415_), .A2(new_n8413_), .B1(new_n8409_), .B2(new_n8412_), .ZN(new_n8416_));
  XOR2_X1    g08223(.A1(new_n8407_), .A2(new_n8416_), .Z(new_n8417_));
  NOR2_X1    g08224(.A1(new_n6563_), .A2(new_n893_), .ZN(new_n8418_));
  NOR2_X1    g08225(.A1(new_n1173_), .A2(new_n6127_), .ZN(new_n8419_));
  NOR2_X1    g08226(.A1(new_n5175_), .A2(new_n5617_), .ZN(new_n8420_));
  INV_X1     g08227(.I(new_n8420_), .ZN(new_n8421_));
  NOR2_X1    g08228(.A1(new_n2028_), .A2(new_n8421_), .ZN(new_n8422_));
  NOR2_X1    g08229(.A1(new_n8419_), .A2(new_n8422_), .ZN(new_n8423_));
  NOR2_X1    g08230(.A1(new_n8423_), .A2(new_n8418_), .ZN(new_n8424_));
  NAND2_X1   g08231(.A1(\a[14] ), .A2(\a[54] ), .ZN(new_n8425_));
  AOI22_X1   g08232(.A1(\a[15] ), .A2(\a[53] ), .B1(\a[16] ), .B2(\a[52] ), .ZN(new_n8426_));
  NOR2_X1    g08233(.A1(new_n8424_), .A2(new_n8418_), .ZN(new_n8427_));
  INV_X1     g08234(.I(new_n8427_), .ZN(new_n8428_));
  OAI22_X1   g08235(.A1(new_n8428_), .A2(new_n8426_), .B1(new_n8424_), .B2(new_n8425_), .ZN(new_n8429_));
  AOI22_X1   g08236(.A1(\a[22] ), .A2(\a[46] ), .B1(\a[23] ), .B2(\a[45] ), .ZN(new_n8430_));
  NOR2_X1    g08237(.A1(new_n1043_), .A2(new_n4596_), .ZN(new_n8431_));
  NOR2_X1    g08238(.A1(new_n2385_), .A2(new_n4430_), .ZN(new_n8432_));
  OAI21_X1   g08239(.A1(new_n8432_), .A2(new_n8430_), .B(new_n8431_), .ZN(new_n8433_));
  INV_X1     g08240(.I(new_n8431_), .ZN(new_n8434_));
  OAI22_X1   g08241(.A1(new_n2385_), .A2(new_n4430_), .B1(new_n8434_), .B2(new_n8430_), .ZN(new_n8435_));
  OAI21_X1   g08242(.A1(new_n8430_), .A2(new_n8435_), .B(new_n8433_), .ZN(new_n8436_));
  XOR2_X1    g08243(.A1(new_n8429_), .A2(new_n8436_), .Z(new_n8437_));
  NAND2_X1   g08244(.A1(new_n2080_), .A2(new_n3860_), .ZN(new_n8438_));
  NAND2_X1   g08245(.A1(new_n1778_), .A2(new_n4342_), .ZN(new_n8439_));
  AOI22_X1   g08246(.A1(new_n8438_), .A2(new_n8439_), .B1(new_n2176_), .B2(new_n4180_), .ZN(new_n8440_));
  NAND2_X1   g08247(.A1(\a[24] ), .A2(\a[44] ), .ZN(new_n8441_));
  AOI22_X1   g08248(.A1(\a[25] ), .A2(\a[43] ), .B1(\a[26] ), .B2(\a[42] ), .ZN(new_n8442_));
  NAND2_X1   g08249(.A1(new_n2176_), .A2(new_n4180_), .ZN(new_n8443_));
  NAND3_X1   g08250(.A1(new_n8443_), .A2(new_n8438_), .A3(new_n8439_), .ZN(new_n8444_));
  OAI22_X1   g08251(.A1(new_n8440_), .A2(new_n8441_), .B1(new_n8444_), .B2(new_n8442_), .ZN(new_n8445_));
  XOR2_X1    g08252(.A1(new_n8437_), .A2(new_n8445_), .Z(new_n8446_));
  XOR2_X1    g08253(.A1(new_n8417_), .A2(new_n8446_), .Z(new_n8447_));
  XOR2_X1    g08254(.A1(new_n8447_), .A2(new_n8389_), .Z(new_n8448_));
  XOR2_X1    g08255(.A1(new_n8363_), .A2(new_n8448_), .Z(new_n8449_));
  XOR2_X1    g08256(.A1(new_n8449_), .A2(new_n8352_), .Z(new_n8450_));
  NOR2_X1    g08257(.A1(new_n8349_), .A2(new_n8450_), .ZN(new_n8451_));
  NAND2_X1   g08258(.A1(new_n8349_), .A2(new_n8450_), .ZN(new_n8452_));
  INV_X1     g08259(.I(new_n8452_), .ZN(new_n8453_));
  NOR2_X1    g08260(.A1(new_n8453_), .A2(new_n8451_), .ZN(new_n8454_));
  INV_X1     g08261(.I(new_n8454_), .ZN(new_n8455_));
  NAND2_X1   g08262(.A1(new_n8455_), .A2(new_n8347_), .ZN(new_n8456_));
  NOR2_X1    g08263(.A1(new_n8455_), .A2(new_n8347_), .ZN(new_n8457_));
  INV_X1     g08264(.I(new_n8457_), .ZN(new_n8458_));
  AND2_X2    g08265(.A1(new_n8458_), .A2(new_n8456_), .Z(new_n8459_));
  NOR2_X1    g08266(.A1(new_n8246_), .A2(new_n8243_), .ZN(new_n8460_));
  NAND2_X1   g08267(.A1(new_n8233_), .A2(new_n8231_), .ZN(new_n8461_));
  NAND2_X1   g08268(.A1(new_n8234_), .A2(new_n8228_), .ZN(new_n8462_));
  NAND2_X1   g08269(.A1(new_n8462_), .A2(new_n8461_), .ZN(new_n8463_));
  XOR2_X1    g08270(.A1(new_n8291_), .A2(new_n8166_), .Z(new_n8464_));
  XOR2_X1    g08271(.A1(new_n8464_), .A2(new_n8284_), .Z(new_n8465_));
  XOR2_X1    g08272(.A1(new_n8274_), .A2(new_n8315_), .Z(new_n8466_));
  NOR2_X1    g08273(.A1(new_n8466_), .A2(new_n8301_), .ZN(new_n8467_));
  AND2_X2    g08274(.A1(new_n8466_), .A2(new_n8301_), .Z(new_n8468_));
  NOR2_X1    g08275(.A1(new_n8468_), .A2(new_n8467_), .ZN(new_n8469_));
  XNOR2_X1   g08276(.A1(new_n8465_), .A2(new_n8469_), .ZN(new_n8470_));
  XNOR2_X1   g08277(.A1(new_n8463_), .A2(new_n8470_), .ZN(new_n8471_));
  XOR2_X1    g08278(.A1(new_n8256_), .A2(new_n8265_), .Z(new_n8472_));
  AND2_X2    g08279(.A1(new_n8472_), .A2(new_n8325_), .Z(new_n8473_));
  NOR2_X1    g08280(.A1(new_n8472_), .A2(new_n8325_), .ZN(new_n8474_));
  NOR2_X1    g08281(.A1(new_n8473_), .A2(new_n8474_), .ZN(new_n8475_));
  NAND2_X1   g08282(.A1(new_n8258_), .A2(new_n8267_), .ZN(new_n8476_));
  OAI21_X1   g08283(.A1(new_n8268_), .A2(new_n8277_), .B(new_n8476_), .ZN(new_n8477_));
  NAND2_X1   g08284(.A1(new_n8317_), .A2(new_n8311_), .ZN(new_n8478_));
  INV_X1     g08285(.I(new_n8318_), .ZN(new_n8479_));
  NAND2_X1   g08286(.A1(new_n8479_), .A2(new_n8326_), .ZN(new_n8480_));
  NAND2_X1   g08287(.A1(new_n8480_), .A2(new_n8478_), .ZN(new_n8481_));
  XOR2_X1    g08288(.A1(new_n8481_), .A2(new_n8477_), .Z(new_n8482_));
  XOR2_X1    g08289(.A1(new_n8482_), .A2(new_n8475_), .Z(new_n8483_));
  XNOR2_X1   g08290(.A1(new_n8483_), .A2(new_n8471_), .ZN(new_n8484_));
  NAND2_X1   g08291(.A1(new_n8460_), .A2(new_n8484_), .ZN(new_n8485_));
  OR2_X2     g08292(.A1(new_n8460_), .A2(new_n8484_), .Z(new_n8486_));
  AND2_X2    g08293(.A1(new_n8486_), .A2(new_n8485_), .Z(new_n8487_));
  INV_X1     g08294(.I(new_n8198_), .ZN(new_n8488_));
  NOR2_X1    g08295(.A1(new_n8488_), .A2(new_n8207_), .ZN(new_n8489_));
  NOR2_X1    g08296(.A1(new_n8211_), .A2(new_n8489_), .ZN(new_n8490_));
  NAND2_X1   g08297(.A1(new_n8328_), .A2(new_n8278_), .ZN(new_n8491_));
  OAI21_X1   g08298(.A1(new_n8303_), .A2(new_n8327_), .B(new_n8491_), .ZN(new_n8492_));
  NAND2_X1   g08299(.A1(new_n8292_), .A2(new_n8285_), .ZN(new_n8493_));
  NAND2_X1   g08300(.A1(new_n8293_), .A2(new_n8302_), .ZN(new_n8494_));
  NAND2_X1   g08301(.A1(new_n8494_), .A2(new_n8493_), .ZN(new_n8495_));
  NAND2_X1   g08302(.A1(new_n8158_), .A2(new_n8167_), .ZN(new_n8496_));
  OAI21_X1   g08303(.A1(new_n8070_), .A2(new_n8108_), .B(new_n8496_), .ZN(new_n8497_));
  NAND2_X1   g08304(.A1(new_n8201_), .A2(new_n8092_), .ZN(new_n8498_));
  OAI21_X1   g08305(.A1(new_n8084_), .A2(new_n8100_), .B(new_n8498_), .ZN(new_n8499_));
  XOR2_X1    g08306(.A1(new_n8499_), .A2(new_n8497_), .Z(new_n8500_));
  XOR2_X1    g08307(.A1(new_n8500_), .A2(new_n8495_), .Z(new_n8501_));
  NAND2_X1   g08308(.A1(new_n8054_), .A2(new_n7969_), .ZN(new_n8502_));
  NAND2_X1   g08309(.A1(new_n8199_), .A2(new_n8061_), .ZN(new_n8503_));
  NAND2_X1   g08310(.A1(new_n8503_), .A2(new_n8502_), .ZN(new_n8504_));
  NAND2_X1   g08311(.A1(new_n8125_), .A2(new_n8203_), .ZN(new_n8505_));
  NAND2_X1   g08312(.A1(new_n8204_), .A2(new_n8117_), .ZN(new_n8506_));
  NAND2_X1   g08313(.A1(new_n8506_), .A2(new_n8505_), .ZN(new_n8507_));
  NOR2_X1    g08314(.A1(new_n7454_), .A2(new_n415_), .ZN(new_n8508_));
  INV_X1     g08315(.I(new_n8508_), .ZN(new_n8509_));
  NOR2_X1    g08316(.A1(new_n355_), .A2(new_n6723_), .ZN(new_n8510_));
  NOR2_X1    g08317(.A1(new_n422_), .A2(new_n6897_), .ZN(new_n8511_));
  OAI21_X1   g08318(.A1(new_n8510_), .A2(new_n8511_), .B(new_n8509_), .ZN(new_n8512_));
  XNOR2_X1   g08319(.A1(new_n8512_), .A2(new_n8309_), .ZN(new_n8513_));
  INV_X1     g08320(.I(new_n8513_), .ZN(new_n8514_));
  XOR2_X1    g08321(.A1(new_n8507_), .A2(new_n8514_), .Z(new_n8515_));
  XOR2_X1    g08322(.A1(new_n8515_), .A2(new_n8504_), .Z(new_n8516_));
  XOR2_X1    g08323(.A1(new_n8501_), .A2(new_n8516_), .Z(new_n8517_));
  XOR2_X1    g08324(.A1(new_n8517_), .A2(new_n8492_), .Z(new_n8518_));
  XOR2_X1    g08325(.A1(new_n8490_), .A2(new_n8518_), .Z(new_n8519_));
  XOR2_X1    g08326(.A1(new_n8487_), .A2(new_n8519_), .Z(new_n8520_));
  NAND2_X1   g08327(.A1(new_n8222_), .A2(new_n8225_), .ZN(new_n8521_));
  NAND2_X1   g08328(.A1(new_n8333_), .A2(new_n8521_), .ZN(new_n8522_));
  XOR2_X1    g08329(.A1(new_n8522_), .A2(new_n8520_), .Z(new_n8523_));
  XOR2_X1    g08330(.A1(new_n8523_), .A2(new_n8459_), .Z(new_n8524_));
  INV_X1     g08331(.I(new_n8524_), .ZN(new_n8525_));
  NAND2_X1   g08332(.A1(new_n8154_), .A2(new_n8218_), .ZN(new_n8526_));
  NAND2_X1   g08333(.A1(new_n8335_), .A2(new_n8526_), .ZN(new_n8527_));
  NOR2_X1    g08334(.A1(new_n8525_), .A2(new_n8527_), .ZN(new_n8528_));
  INV_X1     g08335(.I(new_n8528_), .ZN(new_n8529_));
  NAND2_X1   g08336(.A1(new_n8525_), .A2(new_n8527_), .ZN(new_n8530_));
  NAND2_X1   g08337(.A1(new_n8529_), .A2(new_n8530_), .ZN(new_n8531_));
  XOR2_X1    g08338(.A1(new_n8345_), .A2(new_n8531_), .Z(\asquared[69] ));
  OAI21_X1   g08339(.A1(new_n8344_), .A2(new_n8340_), .B(new_n8529_), .ZN(new_n8533_));
  NAND2_X1   g08340(.A1(new_n8533_), .A2(new_n8530_), .ZN(new_n8534_));
  NOR2_X1    g08341(.A1(new_n8457_), .A2(new_n8453_), .ZN(new_n8535_));
  NAND2_X1   g08342(.A1(new_n8358_), .A2(new_n8361_), .ZN(new_n8536_));
  NAND2_X1   g08343(.A1(new_n8362_), .A2(new_n8355_), .ZN(new_n8537_));
  NAND2_X1   g08344(.A1(new_n8537_), .A2(new_n8536_), .ZN(new_n8538_));
  NAND2_X1   g08345(.A1(new_n8507_), .A2(new_n8514_), .ZN(new_n8539_));
  NAND2_X1   g08346(.A1(new_n8515_), .A2(new_n8504_), .ZN(new_n8540_));
  NAND2_X1   g08347(.A1(new_n8540_), .A2(new_n8539_), .ZN(new_n8541_));
  NAND2_X1   g08348(.A1(new_n8406_), .A2(new_n8396_), .ZN(new_n8542_));
  NAND2_X1   g08349(.A1(new_n8407_), .A2(new_n8416_), .ZN(new_n8543_));
  NAND2_X1   g08350(.A1(new_n8543_), .A2(new_n8542_), .ZN(new_n8544_));
  NAND2_X1   g08351(.A1(new_n8429_), .A2(new_n8436_), .ZN(new_n8545_));
  NAND2_X1   g08352(.A1(new_n8437_), .A2(new_n8445_), .ZN(new_n8546_));
  NAND2_X1   g08353(.A1(new_n8546_), .A2(new_n8545_), .ZN(new_n8547_));
  XOR2_X1    g08354(.A1(new_n8544_), .A2(new_n8547_), .Z(new_n8548_));
  XOR2_X1    g08355(.A1(new_n8548_), .A2(new_n8541_), .Z(new_n8549_));
  XOR2_X1    g08356(.A1(new_n8385_), .A2(new_n8369_), .Z(new_n8550_));
  XOR2_X1    g08357(.A1(new_n8550_), .A2(new_n8435_), .Z(new_n8551_));
  XOR2_X1    g08358(.A1(new_n8404_), .A2(new_n8394_), .Z(new_n8552_));
  XOR2_X1    g08359(.A1(new_n8552_), .A2(new_n8428_), .Z(new_n8553_));
  NAND2_X1   g08360(.A1(new_n8371_), .A2(new_n8378_), .ZN(new_n8554_));
  OAI21_X1   g08361(.A1(new_n8379_), .A2(new_n8388_), .B(new_n8554_), .ZN(new_n8555_));
  XOR2_X1    g08362(.A1(new_n8555_), .A2(new_n8553_), .Z(new_n8556_));
  XOR2_X1    g08363(.A1(new_n8556_), .A2(new_n8551_), .Z(new_n8557_));
  XOR2_X1    g08364(.A1(new_n8549_), .A2(new_n8557_), .Z(new_n8558_));
  XOR2_X1    g08365(.A1(new_n8558_), .A2(new_n8538_), .Z(new_n8559_));
  NAND2_X1   g08366(.A1(new_n8483_), .A2(new_n8471_), .ZN(new_n8560_));
  NAND2_X1   g08367(.A1(new_n8486_), .A2(new_n8560_), .ZN(new_n8561_));
  NAND2_X1   g08368(.A1(new_n8447_), .A2(new_n8389_), .ZN(new_n8562_));
  NAND2_X1   g08369(.A1(new_n8417_), .A2(new_n8446_), .ZN(new_n8563_));
  NAND2_X1   g08370(.A1(new_n8562_), .A2(new_n8563_), .ZN(new_n8564_));
  INV_X1     g08371(.I(new_n8463_), .ZN(new_n8565_));
  NAND2_X1   g08372(.A1(new_n8465_), .A2(new_n8469_), .ZN(new_n8566_));
  OAI21_X1   g08373(.A1(new_n8565_), .A2(new_n8470_), .B(new_n8566_), .ZN(new_n8567_));
  XOR2_X1    g08374(.A1(new_n8415_), .A2(new_n8444_), .Z(new_n8568_));
  XOR2_X1    g08375(.A1(new_n8568_), .A2(new_n8377_), .Z(new_n8569_));
  NOR2_X1    g08376(.A1(new_n8274_), .A2(new_n8315_), .ZN(new_n8570_));
  NOR2_X1    g08377(.A1(new_n8468_), .A2(new_n8570_), .ZN(new_n8571_));
  NOR2_X1    g08378(.A1(new_n8256_), .A2(new_n8265_), .ZN(new_n8572_));
  NOR2_X1    g08379(.A1(new_n8473_), .A2(new_n8572_), .ZN(new_n8573_));
  XOR2_X1    g08380(.A1(new_n8571_), .A2(new_n8573_), .Z(new_n8574_));
  XOR2_X1    g08381(.A1(new_n8574_), .A2(new_n8569_), .Z(new_n8575_));
  NOR2_X1    g08382(.A1(new_n8567_), .A2(new_n8575_), .ZN(new_n8576_));
  NAND2_X1   g08383(.A1(new_n8567_), .A2(new_n8575_), .ZN(new_n8577_));
  INV_X1     g08384(.I(new_n8577_), .ZN(new_n8578_));
  NOR2_X1    g08385(.A1(new_n8578_), .A2(new_n8576_), .ZN(new_n8579_));
  NOR2_X1    g08386(.A1(new_n8579_), .A2(new_n8564_), .ZN(new_n8580_));
  NAND2_X1   g08387(.A1(new_n8579_), .A2(new_n8564_), .ZN(new_n8581_));
  INV_X1     g08388(.I(new_n8581_), .ZN(new_n8582_));
  NOR2_X1    g08389(.A1(new_n8582_), .A2(new_n8580_), .ZN(new_n8583_));
  XOR2_X1    g08390(.A1(new_n8561_), .A2(new_n8583_), .Z(new_n8584_));
  XOR2_X1    g08391(.A1(new_n8584_), .A2(new_n8559_), .Z(new_n8585_));
  XOR2_X1    g08392(.A1(new_n8535_), .A2(new_n8585_), .Z(new_n8586_));
  NAND2_X1   g08393(.A1(new_n8481_), .A2(new_n8477_), .ZN(new_n8587_));
  NAND2_X1   g08394(.A1(new_n8482_), .A2(new_n8475_), .ZN(new_n8588_));
  NAND2_X1   g08395(.A1(new_n8588_), .A2(new_n8587_), .ZN(new_n8589_));
  NAND2_X1   g08396(.A1(new_n8291_), .A2(new_n8166_), .ZN(new_n8590_));
  NAND2_X1   g08397(.A1(new_n8464_), .A2(new_n8284_), .ZN(new_n8591_));
  NAND2_X1   g08398(.A1(new_n8591_), .A2(new_n8590_), .ZN(new_n8592_));
  NAND2_X1   g08399(.A1(new_n1027_), .A2(new_n5524_), .ZN(new_n8593_));
  OAI22_X1   g08400(.A1(new_n2851_), .A2(new_n5523_), .B1(new_n5440_), .B2(new_n1092_), .ZN(new_n8594_));
  NAND2_X1   g08401(.A1(new_n8594_), .A2(new_n8593_), .ZN(new_n8595_));
  NAND3_X1   g08402(.A1(new_n8595_), .A2(\a[19] ), .A3(\a[50] ), .ZN(new_n8596_));
  AOI22_X1   g08403(.A1(\a[17] ), .A2(\a[52] ), .B1(\a[18] ), .B2(\a[51] ), .ZN(new_n8597_));
  NAND2_X1   g08404(.A1(new_n8595_), .A2(new_n8593_), .ZN(new_n8598_));
  OAI21_X1   g08405(.A1(new_n8597_), .A2(new_n8598_), .B(new_n8596_), .ZN(new_n8599_));
  OAI22_X1   g08406(.A1(new_n2679_), .A2(new_n5377_), .B1(new_n3811_), .B2(new_n3329_), .ZN(new_n8600_));
  OAI21_X1   g08407(.A1(new_n2255_), .A2(new_n3551_), .B(new_n8600_), .ZN(new_n8601_));
  NAND3_X1   g08408(.A1(new_n8601_), .A2(\a[28] ), .A3(\a[41] ), .ZN(new_n8602_));
  AOI22_X1   g08409(.A1(\a[29] ), .A2(\a[40] ), .B1(\a[30] ), .B2(\a[39] ), .ZN(new_n8603_));
  NOR2_X1    g08410(.A1(new_n2255_), .A2(new_n3551_), .ZN(new_n8604_));
  NOR2_X1    g08411(.A1(new_n8600_), .A2(new_n8604_), .ZN(new_n8605_));
  INV_X1     g08412(.I(new_n8605_), .ZN(new_n8606_));
  OAI21_X1   g08413(.A1(new_n8603_), .A2(new_n8606_), .B(new_n8602_), .ZN(new_n8607_));
  XOR2_X1    g08414(.A1(new_n8607_), .A2(new_n8599_), .Z(new_n8608_));
  XOR2_X1    g08415(.A1(new_n8608_), .A2(new_n8592_), .Z(new_n8609_));
  INV_X1     g08416(.I(new_n8609_), .ZN(new_n8610_));
  NOR2_X1    g08417(.A1(new_n2637_), .A2(new_n3038_), .ZN(new_n8611_));
  AOI22_X1   g08418(.A1(new_n2275_), .A2(new_n2915_), .B1(new_n3210_), .B2(new_n3803_), .ZN(new_n8612_));
  NOR2_X1    g08419(.A1(new_n8611_), .A2(new_n8612_), .ZN(new_n8613_));
  NOR3_X1    g08420(.A1(new_n8613_), .A2(new_n2051_), .A3(new_n2914_), .ZN(new_n8614_));
  AOI22_X1   g08421(.A1(\a[32] ), .A2(\a[37] ), .B1(\a[33] ), .B2(\a[36] ), .ZN(new_n8615_));
  NOR2_X1    g08422(.A1(new_n8613_), .A2(new_n8611_), .ZN(new_n8616_));
  INV_X1     g08423(.I(new_n8616_), .ZN(new_n8617_));
  NOR2_X1    g08424(.A1(new_n8617_), .A2(new_n8615_), .ZN(new_n8618_));
  NOR2_X1    g08425(.A1(new_n8618_), .A2(new_n8614_), .ZN(new_n8619_));
  AOI21_X1   g08426(.A1(\a[7] ), .A2(\a[62] ), .B(\a[35] ), .ZN(new_n8620_));
  NOR2_X1    g08427(.A1(new_n3589_), .A2(new_n7144_), .ZN(new_n8621_));
  NOR2_X1    g08428(.A1(new_n8621_), .A2(new_n2746_), .ZN(new_n8622_));
  NOR2_X1    g08429(.A1(new_n8621_), .A2(new_n2745_), .ZN(new_n8623_));
  INV_X1     g08430(.I(new_n8623_), .ZN(new_n8624_));
  OAI22_X1   g08431(.A1(new_n8624_), .A2(new_n8620_), .B1(new_n2746_), .B2(new_n8622_), .ZN(new_n8625_));
  INV_X1     g08432(.I(new_n8625_), .ZN(new_n8626_));
  XOR2_X1    g08433(.A1(new_n8619_), .A2(new_n8626_), .Z(new_n8627_));
  NOR2_X1    g08434(.A1(new_n1043_), .A2(new_n5617_), .ZN(new_n8628_));
  NAND2_X1   g08435(.A1(new_n7656_), .A2(new_n8628_), .ZN(new_n8629_));
  NAND2_X1   g08436(.A1(new_n6126_), .A2(new_n1288_), .ZN(new_n8630_));
  NAND3_X1   g08437(.A1(new_n5565_), .A2(\a[16] ), .A3(\a[53] ), .ZN(new_n8631_));
  INV_X1     g08438(.I(new_n8631_), .ZN(new_n8632_));
  AOI21_X1   g08439(.A1(new_n8629_), .A2(new_n8630_), .B(new_n8632_), .ZN(new_n8633_));
  NAND2_X1   g08440(.A1(\a[15] ), .A2(\a[54] ), .ZN(new_n8634_));
  AOI21_X1   g08441(.A1(\a[16] ), .A2(\a[53] ), .B(new_n5565_), .ZN(new_n8635_));
  NAND3_X1   g08442(.A1(new_n8629_), .A2(new_n8631_), .A3(new_n8630_), .ZN(new_n8636_));
  OAI22_X1   g08443(.A1(new_n8633_), .A2(new_n8634_), .B1(new_n8636_), .B2(new_n8635_), .ZN(new_n8637_));
  XNOR2_X1   g08444(.A1(new_n8627_), .A2(new_n8637_), .ZN(new_n8638_));
  NOR2_X1    g08445(.A1(new_n8610_), .A2(new_n8638_), .ZN(new_n8639_));
  INV_X1     g08446(.I(new_n8639_), .ZN(new_n8640_));
  NAND2_X1   g08447(.A1(new_n8610_), .A2(new_n8638_), .ZN(new_n8641_));
  NAND3_X1   g08448(.A1(new_n8589_), .A2(new_n8640_), .A3(new_n8641_), .ZN(new_n8642_));
  NAND2_X1   g08449(.A1(new_n8642_), .A2(new_n8589_), .ZN(new_n8643_));
  NAND3_X1   g08450(.A1(new_n8642_), .A2(new_n8640_), .A3(new_n8641_), .ZN(new_n8644_));
  NAND2_X1   g08451(.A1(new_n8644_), .A2(new_n8643_), .ZN(new_n8645_));
  NAND2_X1   g08452(.A1(new_n8501_), .A2(new_n8516_), .ZN(new_n8646_));
  NAND2_X1   g08453(.A1(new_n8517_), .A2(new_n8492_), .ZN(new_n8647_));
  NAND2_X1   g08454(.A1(new_n8647_), .A2(new_n8646_), .ZN(new_n8648_));
  XOR2_X1    g08455(.A1(new_n8645_), .A2(new_n8648_), .Z(new_n8649_));
  AOI22_X1   g08456(.A1(\a[21] ), .A2(\a[48] ), .B1(\a[22] ), .B2(\a[47] ), .ZN(new_n8650_));
  NOR2_X1    g08457(.A1(new_n759_), .A2(new_n5680_), .ZN(new_n8651_));
  INV_X1     g08458(.I(new_n8651_), .ZN(new_n8652_));
  NOR2_X1    g08459(.A1(new_n1456_), .A2(new_n4977_), .ZN(new_n8653_));
  NOR3_X1    g08460(.A1(new_n8653_), .A2(new_n8650_), .A3(new_n8652_), .ZN(new_n8654_));
  NOR2_X1    g08461(.A1(new_n8654_), .A2(new_n8653_), .ZN(new_n8655_));
  INV_X1     g08462(.I(new_n8655_), .ZN(new_n8656_));
  OAI22_X1   g08463(.A1(new_n8656_), .A2(new_n8650_), .B1(new_n8652_), .B2(new_n8654_), .ZN(new_n8657_));
  NOR2_X1    g08464(.A1(new_n1265_), .A2(new_n8161_), .ZN(new_n8658_));
  AOI22_X1   g08465(.A1(new_n1261_), .A2(new_n6803_), .B1(new_n6317_), .B2(new_n834_), .ZN(new_n8659_));
  NOR2_X1    g08466(.A1(new_n8658_), .A2(new_n8659_), .ZN(new_n8660_));
  NOR3_X1    g08467(.A1(new_n8660_), .A2(new_n513_), .A3(new_n6316_), .ZN(new_n8661_));
  AOI22_X1   g08468(.A1(\a[12] ), .A2(\a[57] ), .B1(\a[13] ), .B2(\a[56] ), .ZN(new_n8662_));
  NOR2_X1    g08469(.A1(new_n8660_), .A2(new_n8658_), .ZN(new_n8663_));
  INV_X1     g08470(.I(new_n8663_), .ZN(new_n8664_));
  NOR2_X1    g08471(.A1(new_n8664_), .A2(new_n8662_), .ZN(new_n8665_));
  NOR2_X1    g08472(.A1(new_n8665_), .A2(new_n8661_), .ZN(new_n8666_));
  OAI21_X1   g08473(.A1(new_n8512_), .A2(new_n8309_), .B(new_n8509_), .ZN(new_n8667_));
  XOR2_X1    g08474(.A1(new_n8666_), .A2(new_n8667_), .Z(new_n8668_));
  XNOR2_X1   g08475(.A1(new_n8668_), .A2(new_n8657_), .ZN(new_n8669_));
  NAND2_X1   g08476(.A1(new_n8499_), .A2(new_n8497_), .ZN(new_n8670_));
  NAND2_X1   g08477(.A1(new_n8500_), .A2(new_n8495_), .ZN(new_n8671_));
  NAND2_X1   g08478(.A1(new_n8671_), .A2(new_n8670_), .ZN(new_n8672_));
  NOR2_X1    g08479(.A1(new_n7452_), .A2(new_n539_), .ZN(new_n8673_));
  INV_X1     g08480(.I(new_n8673_), .ZN(new_n8674_));
  OAI22_X1   g08481(.A1(new_n413_), .A2(new_n6899_), .B1(new_n7454_), .B2(new_n1427_), .ZN(new_n8675_));
  NAND2_X1   g08482(.A1(new_n8675_), .A2(new_n8674_), .ZN(new_n8676_));
  NAND3_X1   g08483(.A1(new_n8676_), .A2(\a[8] ), .A3(\a[61] ), .ZN(new_n8677_));
  AOI22_X1   g08484(.A1(\a[9] ), .A2(\a[60] ), .B1(\a[10] ), .B2(\a[59] ), .ZN(new_n8678_));
  NAND2_X1   g08485(.A1(new_n8676_), .A2(new_n8674_), .ZN(new_n8679_));
  OAI21_X1   g08486(.A1(new_n8678_), .A2(new_n8679_), .B(new_n8677_), .ZN(new_n8680_));
  NOR2_X1    g08487(.A1(new_n1779_), .A2(new_n4704_), .ZN(new_n8681_));
  NOR2_X1    g08488(.A1(new_n1529_), .A2(new_n4430_), .ZN(new_n8682_));
  NOR2_X1    g08489(.A1(new_n1443_), .A2(new_n6101_), .ZN(new_n8683_));
  NOR2_X1    g08490(.A1(new_n8682_), .A2(new_n8683_), .ZN(new_n8684_));
  NOR2_X1    g08491(.A1(new_n8684_), .A2(new_n8681_), .ZN(new_n8685_));
  NAND2_X1   g08492(.A1(\a[23] ), .A2(\a[46] ), .ZN(new_n8686_));
  AOI22_X1   g08493(.A1(\a[24] ), .A2(\a[45] ), .B1(\a[25] ), .B2(\a[44] ), .ZN(new_n8687_));
  NOR2_X1    g08494(.A1(new_n8685_), .A2(new_n8681_), .ZN(new_n8688_));
  INV_X1     g08495(.I(new_n8688_), .ZN(new_n8689_));
  OAI22_X1   g08496(.A1(new_n8689_), .A2(new_n8687_), .B1(new_n8685_), .B2(new_n8686_), .ZN(new_n8690_));
  XNOR2_X1   g08497(.A1(new_n8690_), .A2(new_n8680_), .ZN(new_n8691_));
  AOI22_X1   g08498(.A1(\a[26] ), .A2(\a[43] ), .B1(\a[27] ), .B2(\a[42] ), .ZN(new_n8692_));
  NOR2_X1    g08499(.A1(new_n367_), .A2(new_n7643_), .ZN(new_n8693_));
  INV_X1     g08500(.I(new_n8693_), .ZN(new_n8694_));
  NOR2_X1    g08501(.A1(new_n1972_), .A2(new_n4181_), .ZN(new_n8695_));
  NOR3_X1    g08502(.A1(new_n8695_), .A2(new_n8692_), .A3(new_n8694_), .ZN(new_n8696_));
  NOR2_X1    g08503(.A1(new_n8696_), .A2(new_n8695_), .ZN(new_n8697_));
  INV_X1     g08504(.I(new_n8697_), .ZN(new_n8698_));
  OAI22_X1   g08505(.A1(new_n8698_), .A2(new_n8692_), .B1(new_n8694_), .B2(new_n8696_), .ZN(new_n8699_));
  INV_X1     g08506(.I(new_n8699_), .ZN(new_n8700_));
  XOR2_X1    g08507(.A1(new_n8691_), .A2(new_n8700_), .Z(new_n8701_));
  XOR2_X1    g08508(.A1(new_n8672_), .A2(new_n8701_), .Z(new_n8702_));
  XOR2_X1    g08509(.A1(new_n8702_), .A2(new_n8669_), .Z(new_n8703_));
  XNOR2_X1   g08510(.A1(new_n8649_), .A2(new_n8703_), .ZN(new_n8704_));
  INV_X1     g08511(.I(new_n8518_), .ZN(new_n8705_));
  NOR2_X1    g08512(.A1(new_n8490_), .A2(new_n8705_), .ZN(new_n8706_));
  INV_X1     g08513(.I(new_n8487_), .ZN(new_n8707_));
  NOR2_X1    g08514(.A1(new_n8707_), .A2(new_n8519_), .ZN(new_n8708_));
  NOR2_X1    g08515(.A1(new_n8708_), .A2(new_n8706_), .ZN(new_n8709_));
  NAND2_X1   g08516(.A1(new_n8363_), .A2(new_n8448_), .ZN(new_n8710_));
  NAND2_X1   g08517(.A1(new_n8449_), .A2(new_n8352_), .ZN(new_n8711_));
  NAND2_X1   g08518(.A1(new_n8711_), .A2(new_n8710_), .ZN(new_n8712_));
  XNOR2_X1   g08519(.A1(new_n8709_), .A2(new_n8712_), .ZN(new_n8713_));
  INV_X1     g08520(.I(new_n8713_), .ZN(new_n8714_));
  OR2_X2     g08521(.A1(new_n8714_), .A2(new_n8704_), .Z(new_n8715_));
  NAND2_X1   g08522(.A1(new_n8714_), .A2(new_n8704_), .ZN(new_n8716_));
  AND2_X2    g08523(.A1(new_n8715_), .A2(new_n8716_), .Z(new_n8717_));
  XOR2_X1    g08524(.A1(new_n8717_), .A2(new_n8586_), .Z(new_n8718_));
  INV_X1     g08525(.I(new_n8718_), .ZN(new_n8719_));
  INV_X1     g08526(.I(new_n8459_), .ZN(new_n8720_));
  INV_X1     g08527(.I(new_n8520_), .ZN(new_n8721_));
  NAND2_X1   g08528(.A1(new_n8522_), .A2(new_n8721_), .ZN(new_n8722_));
  OAI21_X1   g08529(.A1(new_n8523_), .A2(new_n8720_), .B(new_n8722_), .ZN(new_n8723_));
  NOR2_X1    g08530(.A1(new_n8719_), .A2(new_n8723_), .ZN(new_n8724_));
  NAND2_X1   g08531(.A1(new_n8719_), .A2(new_n8723_), .ZN(new_n8725_));
  INV_X1     g08532(.I(new_n8725_), .ZN(new_n8726_));
  NOR2_X1    g08533(.A1(new_n8726_), .A2(new_n8724_), .ZN(new_n8727_));
  XOR2_X1    g08534(.A1(new_n8534_), .A2(new_n8727_), .Z(\asquared[70] ));
  OAI21_X1   g08535(.A1(new_n8457_), .A2(new_n8453_), .B(new_n8585_), .ZN(new_n8729_));
  INV_X1     g08536(.I(new_n8717_), .ZN(new_n8730_));
  OAI21_X1   g08537(.A1(new_n8730_), .A2(new_n8586_), .B(new_n8729_), .ZN(new_n8731_));
  INV_X1     g08538(.I(new_n8731_), .ZN(new_n8732_));
  NOR2_X1    g08539(.A1(new_n8582_), .A2(new_n8578_), .ZN(new_n8733_));
  NAND2_X1   g08540(.A1(new_n747_), .A2(new_n7451_), .ZN(new_n8734_));
  OAI22_X1   g08541(.A1(new_n539_), .A2(new_n7454_), .B1(new_n6899_), .B2(new_n1063_), .ZN(new_n8735_));
  NAND2_X1   g08542(.A1(new_n8735_), .A2(new_n8734_), .ZN(new_n8736_));
  NAND3_X1   g08543(.A1(new_n8736_), .A2(\a[9] ), .A3(\a[61] ), .ZN(new_n8737_));
  AOI22_X1   g08544(.A1(\a[10] ), .A2(\a[60] ), .B1(\a[11] ), .B2(\a[59] ), .ZN(new_n8738_));
  NAND2_X1   g08545(.A1(new_n8736_), .A2(new_n8734_), .ZN(new_n8739_));
  OAI21_X1   g08546(.A1(new_n8738_), .A2(new_n8739_), .B(new_n8737_), .ZN(new_n8740_));
  NOR2_X1    g08547(.A1(new_n1428_), .A2(new_n6127_), .ZN(new_n8741_));
  AOI22_X1   g08548(.A1(new_n1025_), .A2(new_n8420_), .B1(new_n1027_), .B2(new_n5862_), .ZN(new_n8742_));
  NOR2_X1    g08549(.A1(new_n8741_), .A2(new_n8742_), .ZN(new_n8743_));
  AOI22_X1   g08550(.A1(\a[16] ), .A2(\a[54] ), .B1(\a[17] ), .B2(\a[53] ), .ZN(new_n8744_));
  NOR2_X1    g08551(.A1(new_n8743_), .A2(new_n8741_), .ZN(new_n8745_));
  INV_X1     g08552(.I(new_n8745_), .ZN(new_n8746_));
  OAI22_X1   g08553(.A1(new_n8746_), .A2(new_n8744_), .B1(new_n6562_), .B2(new_n8743_), .ZN(new_n8747_));
  XNOR2_X1   g08554(.A1(new_n8747_), .A2(new_n8740_), .ZN(new_n8748_));
  NAND4_X1   g08555(.A1(\a[12] ), .A2(\a[24] ), .A3(\a[46] ), .A4(\a[58] ), .ZN(new_n8749_));
  NAND2_X1   g08556(.A1(new_n763_), .A2(new_n6803_), .ZN(new_n8750_));
  AOI22_X1   g08557(.A1(new_n8750_), .A2(new_n8749_), .B1(new_n6506_), .B2(new_n8075_), .ZN(new_n8751_));
  NAND2_X1   g08558(.A1(\a[12] ), .A2(\a[58] ), .ZN(new_n8752_));
  NAND2_X1   g08559(.A1(new_n6506_), .A2(new_n8075_), .ZN(new_n8753_));
  NAND3_X1   g08560(.A1(new_n8753_), .A2(new_n8750_), .A3(new_n8749_), .ZN(new_n8754_));
  AOI22_X1   g08561(.A1(\a[13] ), .A2(\a[57] ), .B1(\a[24] ), .B2(\a[46] ), .ZN(new_n8755_));
  OAI22_X1   g08562(.A1(new_n8751_), .A2(new_n8752_), .B1(new_n8754_), .B2(new_n8755_), .ZN(new_n8756_));
  XOR2_X1    g08563(.A1(new_n8748_), .A2(new_n8756_), .Z(new_n8757_));
  INV_X1     g08564(.I(new_n8757_), .ZN(new_n8758_));
  XOR2_X1    g08565(.A1(new_n8598_), .A2(new_n8636_), .Z(new_n8759_));
  NOR2_X1    g08566(.A1(new_n3038_), .A2(new_n3932_), .ZN(new_n8760_));
  INV_X1     g08567(.I(new_n8760_), .ZN(new_n8761_));
  NOR4_X1    g08568(.A1(new_n2200_), .A2(new_n2442_), .A3(new_n2626_), .A4(new_n2914_), .ZN(new_n8762_));
  NOR2_X1    g08569(.A1(new_n2637_), .A2(new_n6140_), .ZN(new_n8763_));
  OAI21_X1   g08570(.A1(new_n8762_), .A2(new_n8763_), .B(new_n8761_), .ZN(new_n8764_));
  NAND2_X1   g08571(.A1(new_n8764_), .A2(new_n8761_), .ZN(new_n8765_));
  AOI21_X1   g08572(.A1(\a[33] ), .A2(\a[37] ), .B(new_n3822_), .ZN(new_n8766_));
  NAND3_X1   g08573(.A1(new_n8764_), .A2(\a[32] ), .A3(\a[38] ), .ZN(new_n8767_));
  OAI21_X1   g08574(.A1(new_n8765_), .A2(new_n8766_), .B(new_n8767_), .ZN(new_n8768_));
  XOR2_X1    g08575(.A1(new_n8759_), .A2(new_n8768_), .Z(new_n8769_));
  NAND2_X1   g08576(.A1(new_n8574_), .A2(new_n8569_), .ZN(new_n8770_));
  OAI21_X1   g08577(.A1(new_n8571_), .A2(new_n8573_), .B(new_n8770_), .ZN(new_n8771_));
  XOR2_X1    g08578(.A1(new_n8771_), .A2(new_n8769_), .Z(new_n8772_));
  XOR2_X1    g08579(.A1(new_n8772_), .A2(new_n8758_), .Z(new_n8773_));
  INV_X1     g08580(.I(new_n8773_), .ZN(new_n8774_));
  NAND2_X1   g08581(.A1(new_n8733_), .A2(new_n8774_), .ZN(new_n8775_));
  NOR2_X1    g08582(.A1(new_n8733_), .A2(new_n8774_), .ZN(new_n8776_));
  INV_X1     g08583(.I(new_n8776_), .ZN(new_n8777_));
  AND2_X2    g08584(.A1(new_n8777_), .A2(new_n8775_), .Z(new_n8778_));
  NAND2_X1   g08585(.A1(new_n8555_), .A2(new_n8553_), .ZN(new_n8779_));
  NAND2_X1   g08586(.A1(new_n8556_), .A2(new_n8551_), .ZN(new_n8780_));
  NAND2_X1   g08587(.A1(new_n8780_), .A2(new_n8779_), .ZN(new_n8781_));
  NAND2_X1   g08588(.A1(new_n8552_), .A2(new_n8428_), .ZN(new_n8782_));
  OAI21_X1   g08589(.A1(new_n8394_), .A2(new_n8404_), .B(new_n8782_), .ZN(new_n8783_));
  OAI22_X1   g08590(.A1(new_n2255_), .A2(new_n5377_), .B1(new_n5625_), .B2(new_n3329_), .ZN(new_n8784_));
  OAI21_X1   g08591(.A1(new_n2438_), .A2(new_n3551_), .B(new_n8784_), .ZN(new_n8785_));
  NAND3_X1   g08592(.A1(new_n8785_), .A2(\a[29] ), .A3(\a[41] ), .ZN(new_n8786_));
  AOI22_X1   g08593(.A1(\a[30] ), .A2(\a[40] ), .B1(\a[31] ), .B2(\a[39] ), .ZN(new_n8787_));
  NOR2_X1    g08594(.A1(new_n2438_), .A2(new_n3551_), .ZN(new_n8788_));
  NOR2_X1    g08595(.A1(new_n8784_), .A2(new_n8788_), .ZN(new_n8789_));
  INV_X1     g08596(.I(new_n8789_), .ZN(new_n8790_));
  OAI21_X1   g08597(.A1(new_n8787_), .A2(new_n8790_), .B(new_n8786_), .ZN(new_n8791_));
  AOI22_X1   g08598(.A1(\a[7] ), .A2(\a[63] ), .B1(\a[23] ), .B2(\a[47] ), .ZN(new_n8792_));
  INV_X1     g08599(.I(new_n8792_), .ZN(new_n8793_));
  NOR4_X1    g08600(.A1(new_n422_), .A2(new_n1299_), .A3(new_n4312_), .A4(new_n7643_), .ZN(new_n8794_));
  NOR2_X1    g08601(.A1(new_n1718_), .A2(new_n3746_), .ZN(new_n8795_));
  AOI21_X1   g08602(.A1(new_n8793_), .A2(new_n8795_), .B(new_n8794_), .ZN(new_n8796_));
  INV_X1     g08603(.I(new_n8796_), .ZN(new_n8797_));
  OAI21_X1   g08604(.A1(new_n8794_), .A2(new_n8792_), .B(new_n8795_), .ZN(new_n8798_));
  OAI21_X1   g08605(.A1(new_n8797_), .A2(new_n8792_), .B(new_n8798_), .ZN(new_n8799_));
  XOR2_X1    g08606(.A1(new_n8791_), .A2(new_n8799_), .Z(new_n8800_));
  XOR2_X1    g08607(.A1(new_n8783_), .A2(new_n8800_), .Z(new_n8801_));
  INV_X1     g08608(.I(new_n8801_), .ZN(new_n8802_));
  AOI22_X1   g08609(.A1(\a[14] ), .A2(\a[56] ), .B1(\a[15] ), .B2(\a[55] ), .ZN(new_n8803_));
  INV_X1     g08610(.I(new_n8803_), .ZN(new_n8804_));
  NOR2_X1    g08611(.A1(new_n1173_), .A2(new_n7185_), .ZN(new_n8805_));
  NOR2_X1    g08612(.A1(new_n1175_), .A2(new_n4596_), .ZN(new_n8806_));
  AOI21_X1   g08613(.A1(new_n8804_), .A2(new_n8806_), .B(new_n8805_), .ZN(new_n8807_));
  NAND2_X1   g08614(.A1(new_n8807_), .A2(new_n8804_), .ZN(new_n8808_));
  OAI21_X1   g08615(.A1(new_n8805_), .A2(new_n8803_), .B(new_n8806_), .ZN(new_n8809_));
  NAND2_X1   g08616(.A1(new_n8808_), .A2(new_n8809_), .ZN(new_n8810_));
  NOR2_X1    g08617(.A1(new_n1972_), .A2(new_n4343_), .ZN(new_n8811_));
  NOR2_X1    g08618(.A1(new_n4010_), .A2(new_n4034_), .ZN(new_n8812_));
  NOR2_X1    g08619(.A1(new_n2177_), .A2(new_n4704_), .ZN(new_n8813_));
  NOR2_X1    g08620(.A1(new_n8812_), .A2(new_n8813_), .ZN(new_n8814_));
  NOR2_X1    g08621(.A1(new_n8814_), .A2(new_n8811_), .ZN(new_n8815_));
  NAND2_X1   g08622(.A1(\a[25] ), .A2(\a[45] ), .ZN(new_n8816_));
  AOI22_X1   g08623(.A1(\a[26] ), .A2(\a[44] ), .B1(\a[27] ), .B2(\a[43] ), .ZN(new_n8817_));
  NOR2_X1    g08624(.A1(new_n8815_), .A2(new_n8811_), .ZN(new_n8818_));
  INV_X1     g08625(.I(new_n8818_), .ZN(new_n8819_));
  OAI22_X1   g08626(.A1(new_n8819_), .A2(new_n8817_), .B1(new_n8815_), .B2(new_n8816_), .ZN(new_n8820_));
  XOR2_X1    g08627(.A1(new_n8820_), .A2(new_n8810_), .Z(new_n8821_));
  NOR2_X1    g08628(.A1(new_n1376_), .A2(new_n5440_), .ZN(new_n8822_));
  AOI22_X1   g08629(.A1(new_n1378_), .A2(new_n7867_), .B1(new_n1381_), .B2(new_n5154_), .ZN(new_n8823_));
  NOR2_X1    g08630(.A1(new_n8822_), .A2(new_n8823_), .ZN(new_n8824_));
  NAND2_X1   g08631(.A1(\a[21] ), .A2(\a[49] ), .ZN(new_n8825_));
  AOI22_X1   g08632(.A1(\a[19] ), .A2(\a[51] ), .B1(\a[20] ), .B2(\a[50] ), .ZN(new_n8826_));
  NOR2_X1    g08633(.A1(new_n8824_), .A2(new_n8822_), .ZN(new_n8827_));
  INV_X1     g08634(.I(new_n8827_), .ZN(new_n8828_));
  OAI22_X1   g08635(.A1(new_n8828_), .A2(new_n8826_), .B1(new_n8824_), .B2(new_n8825_), .ZN(new_n8829_));
  XNOR2_X1   g08636(.A1(new_n8821_), .A2(new_n8829_), .ZN(new_n8830_));
  NAND2_X1   g08637(.A1(new_n8802_), .A2(new_n8830_), .ZN(new_n8831_));
  NOR2_X1    g08638(.A1(new_n8802_), .A2(new_n8830_), .ZN(new_n8832_));
  INV_X1     g08639(.I(new_n8832_), .ZN(new_n8833_));
  NAND3_X1   g08640(.A1(new_n8833_), .A2(new_n8781_), .A3(new_n8831_), .ZN(new_n8834_));
  NAND2_X1   g08641(.A1(new_n8834_), .A2(new_n8833_), .ZN(new_n8835_));
  INV_X1     g08642(.I(new_n8835_), .ZN(new_n8836_));
  AOI22_X1   g08643(.A1(new_n8836_), .A2(new_n8831_), .B1(new_n8781_), .B2(new_n8834_), .ZN(new_n8837_));
  XOR2_X1    g08644(.A1(new_n8778_), .A2(new_n8837_), .Z(new_n8838_));
  NAND2_X1   g08645(.A1(new_n8561_), .A2(new_n8583_), .ZN(new_n8839_));
  NAND2_X1   g08646(.A1(new_n8584_), .A2(new_n8559_), .ZN(new_n8840_));
  NAND2_X1   g08647(.A1(new_n8840_), .A2(new_n8839_), .ZN(new_n8841_));
  NAND2_X1   g08648(.A1(new_n8607_), .A2(new_n8599_), .ZN(new_n8842_));
  NAND2_X1   g08649(.A1(new_n8608_), .A2(new_n8592_), .ZN(new_n8843_));
  NAND2_X1   g08650(.A1(new_n8843_), .A2(new_n8842_), .ZN(new_n8844_));
  NOR2_X1    g08651(.A1(new_n8698_), .A2(new_n8606_), .ZN(new_n8845_));
  NOR2_X1    g08652(.A1(new_n8697_), .A2(new_n8605_), .ZN(new_n8846_));
  NOR2_X1    g08653(.A1(new_n8845_), .A2(new_n8846_), .ZN(new_n8847_));
  INV_X1     g08654(.I(new_n8847_), .ZN(new_n8848_));
  NOR2_X1    g08655(.A1(new_n8848_), .A2(new_n8688_), .ZN(new_n8849_));
  INV_X1     g08656(.I(new_n8849_), .ZN(new_n8850_));
  NAND2_X1   g08657(.A1(new_n8848_), .A2(new_n8688_), .ZN(new_n8851_));
  AND2_X2    g08658(.A1(new_n8850_), .A2(new_n8851_), .Z(new_n8852_));
  AOI21_X1   g08659(.A1(\a[8] ), .A2(\a[62] ), .B(new_n8624_), .ZN(new_n8853_));
  INV_X1     g08660(.I(new_n8853_), .ZN(new_n8854_));
  NOR3_X1    g08661(.A1(new_n8623_), .A2(new_n355_), .A3(new_n7144_), .ZN(new_n8855_));
  INV_X1     g08662(.I(new_n8855_), .ZN(new_n8856_));
  NAND3_X1   g08663(.A1(new_n8854_), .A2(new_n8617_), .A3(new_n8856_), .ZN(new_n8857_));
  NAND2_X1   g08664(.A1(new_n8857_), .A2(new_n8856_), .ZN(new_n8858_));
  INV_X1     g08665(.I(new_n8858_), .ZN(new_n8859_));
  AOI22_X1   g08666(.A1(new_n8859_), .A2(new_n8854_), .B1(new_n8617_), .B2(new_n8857_), .ZN(new_n8860_));
  XOR2_X1    g08667(.A1(new_n8852_), .A2(new_n8860_), .Z(new_n8861_));
  XNOR2_X1   g08668(.A1(new_n8861_), .A2(new_n8844_), .ZN(new_n8862_));
  NAND2_X1   g08669(.A1(new_n8642_), .A2(new_n8640_), .ZN(new_n8863_));
  NAND2_X1   g08670(.A1(new_n8627_), .A2(new_n8637_), .ZN(new_n8864_));
  OAI21_X1   g08671(.A1(new_n8619_), .A2(new_n8626_), .B(new_n8864_), .ZN(new_n8865_));
  NAND2_X1   g08672(.A1(new_n8690_), .A2(new_n8680_), .ZN(new_n8866_));
  OAI21_X1   g08673(.A1(new_n8691_), .A2(new_n8700_), .B(new_n8866_), .ZN(new_n8867_));
  INV_X1     g08674(.I(new_n8667_), .ZN(new_n8868_));
  INV_X1     g08675(.I(new_n8668_), .ZN(new_n8869_));
  NAND2_X1   g08676(.A1(new_n8869_), .A2(new_n8657_), .ZN(new_n8870_));
  OAI21_X1   g08677(.A1(new_n8666_), .A2(new_n8868_), .B(new_n8870_), .ZN(new_n8871_));
  XOR2_X1    g08678(.A1(new_n8871_), .A2(new_n8867_), .Z(new_n8872_));
  XOR2_X1    g08679(.A1(new_n8872_), .A2(new_n8865_), .Z(new_n8873_));
  XOR2_X1    g08680(.A1(new_n8863_), .A2(new_n8873_), .Z(new_n8874_));
  XOR2_X1    g08681(.A1(new_n8874_), .A2(new_n8862_), .Z(new_n8875_));
  XNOR2_X1   g08682(.A1(new_n8841_), .A2(new_n8875_), .ZN(new_n8876_));
  XNOR2_X1   g08683(.A1(new_n8876_), .A2(new_n8838_), .ZN(new_n8877_));
  INV_X1     g08684(.I(new_n8877_), .ZN(new_n8878_));
  OAI21_X1   g08685(.A1(new_n8708_), .A2(new_n8706_), .B(new_n8712_), .ZN(new_n8879_));
  NAND2_X1   g08686(.A1(new_n8715_), .A2(new_n8879_), .ZN(new_n8880_));
  NAND2_X1   g08687(.A1(new_n8645_), .A2(new_n8648_), .ZN(new_n8881_));
  NAND2_X1   g08688(.A1(new_n8649_), .A2(new_n8703_), .ZN(new_n8882_));
  NAND2_X1   g08689(.A1(new_n8882_), .A2(new_n8881_), .ZN(new_n8883_));
  NAND2_X1   g08690(.A1(new_n8549_), .A2(new_n8557_), .ZN(new_n8884_));
  NAND2_X1   g08691(.A1(new_n8558_), .A2(new_n8538_), .ZN(new_n8885_));
  NAND2_X1   g08692(.A1(new_n8885_), .A2(new_n8884_), .ZN(new_n8886_));
  NAND2_X1   g08693(.A1(new_n8672_), .A2(new_n8701_), .ZN(new_n8887_));
  NAND2_X1   g08694(.A1(new_n8702_), .A2(new_n8669_), .ZN(new_n8888_));
  NAND2_X1   g08695(.A1(new_n8888_), .A2(new_n8887_), .ZN(new_n8889_));
  NAND2_X1   g08696(.A1(new_n8544_), .A2(new_n8547_), .ZN(new_n8890_));
  NAND2_X1   g08697(.A1(new_n8548_), .A2(new_n8541_), .ZN(new_n8891_));
  NAND2_X1   g08698(.A1(new_n8891_), .A2(new_n8890_), .ZN(new_n8892_));
  NOR2_X1    g08699(.A1(new_n8664_), .A2(new_n8679_), .ZN(new_n8893_));
  NAND2_X1   g08700(.A1(new_n8664_), .A2(new_n8679_), .ZN(new_n8894_));
  INV_X1     g08701(.I(new_n8894_), .ZN(new_n8895_));
  NOR2_X1    g08702(.A1(new_n8895_), .A2(new_n8893_), .ZN(new_n8896_));
  INV_X1     g08703(.I(new_n8896_), .ZN(new_n8897_));
  NOR2_X1    g08704(.A1(new_n8897_), .A2(new_n8655_), .ZN(new_n8898_));
  NOR2_X1    g08705(.A1(new_n8896_), .A2(new_n8656_), .ZN(new_n8899_));
  NOR2_X1    g08706(.A1(new_n8898_), .A2(new_n8899_), .ZN(new_n8900_));
  NAND2_X1   g08707(.A1(new_n8550_), .A2(new_n8435_), .ZN(new_n8901_));
  OAI21_X1   g08708(.A1(new_n8369_), .A2(new_n8385_), .B(new_n8901_), .ZN(new_n8902_));
  NAND2_X1   g08709(.A1(new_n8415_), .A2(new_n8444_), .ZN(new_n8903_));
  NAND2_X1   g08710(.A1(new_n8568_), .A2(new_n8377_), .ZN(new_n8904_));
  NAND2_X1   g08711(.A1(new_n8904_), .A2(new_n8903_), .ZN(new_n8905_));
  XOR2_X1    g08712(.A1(new_n8902_), .A2(new_n8905_), .Z(new_n8906_));
  XOR2_X1    g08713(.A1(new_n8906_), .A2(new_n8900_), .Z(new_n8907_));
  XOR2_X1    g08714(.A1(new_n8892_), .A2(new_n8907_), .Z(new_n8908_));
  XOR2_X1    g08715(.A1(new_n8908_), .A2(new_n8889_), .Z(new_n8909_));
  XOR2_X1    g08716(.A1(new_n8886_), .A2(new_n8909_), .Z(new_n8910_));
  XOR2_X1    g08717(.A1(new_n8910_), .A2(new_n8883_), .Z(new_n8911_));
  NAND2_X1   g08718(.A1(new_n8880_), .A2(new_n8911_), .ZN(new_n8912_));
  NAND2_X1   g08719(.A1(new_n8912_), .A2(new_n8880_), .ZN(new_n8913_));
  NAND2_X1   g08720(.A1(new_n8912_), .A2(new_n8911_), .ZN(new_n8914_));
  NAND2_X1   g08721(.A1(new_n8913_), .A2(new_n8914_), .ZN(new_n8915_));
  NAND2_X1   g08722(.A1(new_n8915_), .A2(new_n8878_), .ZN(new_n8916_));
  NAND3_X1   g08723(.A1(new_n8913_), .A2(new_n8914_), .A3(new_n8877_), .ZN(new_n8917_));
  NAND2_X1   g08724(.A1(new_n8916_), .A2(new_n8917_), .ZN(new_n8918_));
  NOR2_X1    g08725(.A1(new_n8918_), .A2(new_n8732_), .ZN(new_n8919_));
  INV_X1     g08726(.I(new_n8919_), .ZN(new_n8920_));
  AOI21_X1   g08727(.A1(new_n8533_), .A2(new_n8530_), .B(new_n8724_), .ZN(new_n8921_));
  NOR2_X1    g08728(.A1(new_n8921_), .A2(new_n8726_), .ZN(new_n8922_));
  INV_X1     g08729(.I(new_n8530_), .ZN(new_n8923_));
  INV_X1     g08730(.I(new_n7944_), .ZN(new_n8924_));
  OAI21_X1   g08731(.A1(new_n7742_), .A2(new_n7733_), .B(new_n8924_), .ZN(new_n8925_));
  AOI21_X1   g08732(.A1(new_n8925_), .A2(new_n7945_), .B(new_n8142_), .ZN(new_n8926_));
  INV_X1     g08733(.I(new_n8341_), .ZN(new_n8927_));
  OAI21_X1   g08734(.A1(new_n8926_), .A2(new_n8144_), .B(new_n8927_), .ZN(new_n8928_));
  AOI21_X1   g08735(.A1(new_n8928_), .A2(new_n8339_), .B(new_n8528_), .ZN(new_n8929_));
  INV_X1     g08736(.I(new_n8724_), .ZN(new_n8930_));
  OAI21_X1   g08737(.A1(new_n8929_), .A2(new_n8923_), .B(new_n8930_), .ZN(new_n8931_));
  NAND2_X1   g08738(.A1(new_n8918_), .A2(new_n8732_), .ZN(new_n8932_));
  INV_X1     g08739(.I(new_n8932_), .ZN(new_n8933_));
  AOI21_X1   g08740(.A1(new_n8931_), .A2(new_n8725_), .B(new_n8933_), .ZN(new_n8934_));
  NAND2_X1   g08741(.A1(new_n8920_), .A2(new_n8932_), .ZN(new_n8935_));
  AOI22_X1   g08742(.A1(new_n8934_), .A2(new_n8920_), .B1(new_n8922_), .B2(new_n8935_), .ZN(\asquared[71] ));
  OAI21_X1   g08743(.A1(new_n8921_), .A2(new_n8726_), .B(new_n8932_), .ZN(new_n8937_));
  NAND2_X1   g08744(.A1(new_n8937_), .A2(new_n8920_), .ZN(new_n8938_));
  NAND2_X1   g08745(.A1(new_n8916_), .A2(new_n8912_), .ZN(new_n8939_));
  INV_X1     g08746(.I(new_n8939_), .ZN(new_n8940_));
  NAND2_X1   g08747(.A1(new_n8871_), .A2(new_n8867_), .ZN(new_n8941_));
  NAND2_X1   g08748(.A1(new_n8872_), .A2(new_n8865_), .ZN(new_n8942_));
  NAND2_X1   g08749(.A1(new_n8942_), .A2(new_n8941_), .ZN(new_n8943_));
  NOR2_X1    g08750(.A1(new_n1265_), .A2(new_n7206_), .ZN(new_n8944_));
  INV_X1     g08751(.I(new_n8944_), .ZN(new_n8945_));
  NOR2_X1    g08752(.A1(new_n597_), .A2(new_n6316_), .ZN(new_n8946_));
  NOR2_X1    g08753(.A1(new_n536_), .A2(new_n6548_), .ZN(new_n8947_));
  OAI21_X1   g08754(.A1(new_n8946_), .A2(new_n8947_), .B(new_n8945_), .ZN(new_n8948_));
  XOR2_X1    g08755(.A1(new_n8948_), .A2(new_n8827_), .Z(new_n8949_));
  NAND2_X1   g08756(.A1(new_n7184_), .A2(new_n1288_), .ZN(new_n8950_));
  NOR2_X1    g08757(.A1(new_n5680_), .A2(new_n6298_), .ZN(new_n8951_));
  INV_X1     g08758(.I(new_n8951_), .ZN(new_n8952_));
  OAI22_X1   g08759(.A1(new_n2028_), .A2(new_n8952_), .B1(new_n1173_), .B2(new_n8161_), .ZN(new_n8953_));
  NAND2_X1   g08760(.A1(new_n8953_), .A2(new_n8950_), .ZN(new_n8954_));
  NAND3_X1   g08761(.A1(new_n8954_), .A2(\a[14] ), .A3(\a[57] ), .ZN(new_n8955_));
  AOI22_X1   g08762(.A1(\a[15] ), .A2(\a[56] ), .B1(\a[16] ), .B2(\a[55] ), .ZN(new_n8956_));
  NAND2_X1   g08763(.A1(new_n8954_), .A2(new_n8950_), .ZN(new_n8957_));
  OAI21_X1   g08764(.A1(new_n8956_), .A2(new_n8957_), .B(new_n8955_), .ZN(new_n8958_));
  NAND2_X1   g08765(.A1(new_n2176_), .A2(new_n4429_), .ZN(new_n8959_));
  OAI22_X1   g08766(.A1(new_n1779_), .A2(new_n4721_), .B1(new_n2081_), .B2(new_n4314_), .ZN(new_n8960_));
  NAND2_X1   g08767(.A1(new_n8960_), .A2(new_n8959_), .ZN(new_n8961_));
  NAND3_X1   g08768(.A1(new_n8961_), .A2(\a[24] ), .A3(\a[47] ), .ZN(new_n8962_));
  AOI22_X1   g08769(.A1(\a[25] ), .A2(\a[46] ), .B1(\a[26] ), .B2(\a[45] ), .ZN(new_n8963_));
  NAND2_X1   g08770(.A1(new_n8961_), .A2(new_n8959_), .ZN(new_n8964_));
  OAI21_X1   g08771(.A1(new_n8963_), .A2(new_n8964_), .B(new_n8962_), .ZN(new_n8965_));
  XOR2_X1    g08772(.A1(new_n8958_), .A2(new_n8965_), .Z(new_n8966_));
  XOR2_X1    g08773(.A1(new_n8966_), .A2(new_n8949_), .Z(new_n8967_));
  OAI22_X1   g08774(.A1(new_n1816_), .A2(new_n3861_), .B1(new_n2189_), .B2(new_n4343_), .ZN(new_n8968_));
  OAI21_X1   g08775(.A1(new_n2679_), .A2(new_n4181_), .B(new_n8968_), .ZN(new_n8969_));
  NAND3_X1   g08776(.A1(new_n8969_), .A2(\a[27] ), .A3(\a[44] ), .ZN(new_n8970_));
  AOI22_X1   g08777(.A1(\a[28] ), .A2(\a[43] ), .B1(\a[29] ), .B2(\a[42] ), .ZN(new_n8971_));
  NOR2_X1    g08778(.A1(new_n2679_), .A2(new_n4181_), .ZN(new_n8972_));
  NOR2_X1    g08779(.A1(new_n8968_), .A2(new_n8972_), .ZN(new_n8973_));
  INV_X1     g08780(.I(new_n8973_), .ZN(new_n8974_));
  OAI21_X1   g08781(.A1(new_n8971_), .A2(new_n8974_), .B(new_n8970_), .ZN(new_n8975_));
  NAND2_X1   g08782(.A1(new_n3210_), .A2(new_n3550_), .ZN(new_n8976_));
  OAI22_X1   g08783(.A1(new_n2202_), .A2(new_n3329_), .B1(new_n2438_), .B2(new_n5377_), .ZN(new_n8977_));
  NAND2_X1   g08784(.A1(new_n8977_), .A2(new_n8976_), .ZN(new_n8978_));
  NAND3_X1   g08785(.A1(new_n8978_), .A2(\a[30] ), .A3(\a[41] ), .ZN(new_n8979_));
  AOI22_X1   g08786(.A1(\a[31] ), .A2(\a[40] ), .B1(\a[32] ), .B2(\a[39] ), .ZN(new_n8980_));
  NAND2_X1   g08787(.A1(new_n8978_), .A2(new_n8976_), .ZN(new_n8981_));
  OAI21_X1   g08788(.A1(new_n8980_), .A2(new_n8981_), .B(new_n8979_), .ZN(new_n8982_));
  XNOR2_X1   g08789(.A1(new_n8975_), .A2(new_n8982_), .ZN(new_n8983_));
  AOI22_X1   g08790(.A1(\a[17] ), .A2(\a[54] ), .B1(\a[18] ), .B2(\a[53] ), .ZN(new_n8984_));
  NOR2_X1    g08791(.A1(new_n1299_), .A2(new_n4596_), .ZN(new_n8985_));
  INV_X1     g08792(.I(new_n8985_), .ZN(new_n8986_));
  NOR2_X1    g08793(.A1(new_n1275_), .A2(new_n6127_), .ZN(new_n8987_));
  NOR3_X1    g08794(.A1(new_n8987_), .A2(new_n8984_), .A3(new_n8986_), .ZN(new_n8988_));
  NOR2_X1    g08795(.A1(new_n8988_), .A2(new_n8987_), .ZN(new_n8989_));
  INV_X1     g08796(.I(new_n8989_), .ZN(new_n8990_));
  OAI22_X1   g08797(.A1(new_n8990_), .A2(new_n8984_), .B1(new_n8986_), .B2(new_n8988_), .ZN(new_n8991_));
  XOR2_X1    g08798(.A1(new_n8983_), .A2(new_n8991_), .Z(new_n8992_));
  XNOR2_X1   g08799(.A1(new_n8992_), .A2(new_n8967_), .ZN(new_n8993_));
  XOR2_X1    g08800(.A1(new_n8943_), .A2(new_n8993_), .Z(new_n8994_));
  NAND2_X1   g08801(.A1(new_n8892_), .A2(new_n8907_), .ZN(new_n8995_));
  NAND2_X1   g08802(.A1(new_n8908_), .A2(new_n8889_), .ZN(new_n8996_));
  NAND2_X1   g08803(.A1(new_n8996_), .A2(new_n8995_), .ZN(new_n8997_));
  AOI21_X1   g08804(.A1(\a[9] ), .A2(\a[62] ), .B(\a[36] ), .ZN(new_n8998_));
  NAND2_X1   g08805(.A1(\a[22] ), .A2(\a[49] ), .ZN(new_n8999_));
  NAND2_X1   g08806(.A1(\a[36] ), .A2(\a[62] ), .ZN(new_n9000_));
  NOR2_X1    g08807(.A1(new_n9000_), .A2(new_n403_), .ZN(new_n9001_));
  NOR3_X1    g08808(.A1(new_n9001_), .A2(new_n8998_), .A3(new_n8999_), .ZN(new_n9002_));
  OAI22_X1   g08809(.A1(new_n8998_), .A2(new_n8999_), .B1(new_n9000_), .B2(new_n403_), .ZN(new_n9003_));
  OAI22_X1   g08810(.A1(new_n9002_), .A2(new_n8999_), .B1(new_n8998_), .B2(new_n9003_), .ZN(new_n9004_));
  NOR2_X1    g08811(.A1(new_n1376_), .A2(new_n5525_), .ZN(new_n9005_));
  INV_X1     g08812(.I(new_n9005_), .ZN(new_n9006_));
  OAI22_X1   g08813(.A1(new_n1379_), .A2(new_n5523_), .B1(new_n1382_), .B2(new_n5440_), .ZN(new_n9007_));
  NAND2_X1   g08814(.A1(new_n9006_), .A2(new_n9007_), .ZN(new_n9008_));
  NAND3_X1   g08815(.A1(new_n9008_), .A2(\a[21] ), .A3(\a[50] ), .ZN(new_n9009_));
  AOI22_X1   g08816(.A1(\a[19] ), .A2(\a[52] ), .B1(\a[20] ), .B2(\a[51] ), .ZN(new_n9010_));
  NAND2_X1   g08817(.A1(new_n9008_), .A2(new_n9006_), .ZN(new_n9011_));
  OAI21_X1   g08818(.A1(new_n9010_), .A2(new_n9011_), .B(new_n9009_), .ZN(new_n9012_));
  XOR2_X1    g08819(.A1(new_n9012_), .A2(new_n9004_), .Z(new_n9013_));
  INV_X1     g08820(.I(new_n3802_), .ZN(new_n9014_));
  NOR2_X1    g08821(.A1(new_n2442_), .A2(new_n2752_), .ZN(new_n9015_));
  NAND2_X1   g08822(.A1(new_n3577_), .A2(new_n3803_), .ZN(new_n9016_));
  NAND2_X1   g08823(.A1(new_n3232_), .A2(new_n3802_), .ZN(new_n9017_));
  AOI22_X1   g08824(.A1(new_n9016_), .A2(new_n9017_), .B1(new_n3232_), .B2(new_n9015_), .ZN(new_n9018_));
  NOR2_X1    g08825(.A1(new_n3232_), .A2(new_n9015_), .ZN(new_n9019_));
  NAND2_X1   g08826(.A1(new_n3232_), .A2(new_n9015_), .ZN(new_n9020_));
  NAND3_X1   g08827(.A1(new_n9020_), .A2(new_n9016_), .A3(new_n9017_), .ZN(new_n9021_));
  OAI22_X1   g08828(.A1(new_n9018_), .A2(new_n9014_), .B1(new_n9021_), .B2(new_n9019_), .ZN(new_n9022_));
  XOR2_X1    g08829(.A1(new_n9013_), .A2(new_n9022_), .Z(new_n9023_));
  NAND2_X1   g08830(.A1(new_n8902_), .A2(new_n8905_), .ZN(new_n9024_));
  NAND2_X1   g08831(.A1(new_n8906_), .A2(new_n8900_), .ZN(new_n9025_));
  NAND2_X1   g08832(.A1(new_n9025_), .A2(new_n9024_), .ZN(new_n9026_));
  XOR2_X1    g08833(.A1(new_n8765_), .A2(new_n8746_), .Z(new_n9027_));
  NAND2_X1   g08834(.A1(new_n7852_), .A2(new_n1367_), .ZN(new_n9028_));
  NOR2_X1    g08835(.A1(new_n1264_), .A2(new_n7454_), .ZN(new_n9029_));
  NOR2_X1    g08836(.A1(new_n6723_), .A2(new_n7643_), .ZN(new_n9030_));
  INV_X1     g08837(.I(new_n9030_), .ZN(new_n9031_));
  NOR3_X1    g08838(.A1(new_n9031_), .A2(new_n355_), .A3(new_n513_), .ZN(new_n9032_));
  OAI21_X1   g08839(.A1(new_n9032_), .A2(new_n9029_), .B(new_n9028_), .ZN(new_n9033_));
  NAND3_X1   g08840(.A1(new_n9033_), .A2(\a[11] ), .A3(\a[60] ), .ZN(new_n9034_));
  AOI22_X1   g08841(.A1(\a[8] ), .A2(\a[63] ), .B1(\a[10] ), .B2(\a[61] ), .ZN(new_n9035_));
  NAND2_X1   g08842(.A1(new_n9033_), .A2(new_n9028_), .ZN(new_n9036_));
  OAI21_X1   g08843(.A1(new_n9035_), .A2(new_n9036_), .B(new_n9034_), .ZN(new_n9037_));
  XOR2_X1    g08844(.A1(new_n9027_), .A2(new_n9037_), .Z(new_n9038_));
  XOR2_X1    g08845(.A1(new_n9026_), .A2(new_n9038_), .Z(new_n9039_));
  XOR2_X1    g08846(.A1(new_n9039_), .A2(new_n9023_), .Z(new_n9040_));
  XOR2_X1    g08847(.A1(new_n8997_), .A2(new_n9040_), .Z(new_n9041_));
  XNOR2_X1   g08848(.A1(new_n9041_), .A2(new_n8994_), .ZN(new_n9042_));
  NAND2_X1   g08849(.A1(new_n8886_), .A2(new_n8909_), .ZN(new_n9043_));
  NAND2_X1   g08850(.A1(new_n8910_), .A2(new_n8883_), .ZN(new_n9044_));
  NAND2_X1   g08851(.A1(new_n9044_), .A2(new_n9043_), .ZN(new_n9045_));
  NAND2_X1   g08852(.A1(new_n8791_), .A2(new_n8799_), .ZN(new_n9046_));
  NAND2_X1   g08853(.A1(new_n8783_), .A2(new_n8800_), .ZN(new_n9047_));
  NAND2_X1   g08854(.A1(new_n9047_), .A2(new_n9046_), .ZN(new_n9048_));
  XOR2_X1    g08855(.A1(new_n8739_), .A2(new_n8754_), .Z(new_n9049_));
  XOR2_X1    g08856(.A1(new_n9049_), .A2(new_n8819_), .Z(new_n9050_));
  XOR2_X1    g08857(.A1(new_n8789_), .A2(new_n8807_), .Z(new_n9051_));
  INV_X1     g08858(.I(new_n9051_), .ZN(new_n9052_));
  NOR2_X1    g08859(.A1(new_n9052_), .A2(new_n8796_), .ZN(new_n9053_));
  NOR2_X1    g08860(.A1(new_n9051_), .A2(new_n8797_), .ZN(new_n9054_));
  NOR2_X1    g08861(.A1(new_n9053_), .A2(new_n9054_), .ZN(new_n9055_));
  XOR2_X1    g08862(.A1(new_n9050_), .A2(new_n9055_), .Z(new_n9056_));
  XOR2_X1    g08863(.A1(new_n9056_), .A2(new_n9048_), .Z(new_n9057_));
  NAND2_X1   g08864(.A1(new_n8820_), .A2(new_n8810_), .ZN(new_n9058_));
  NAND2_X1   g08865(.A1(new_n8821_), .A2(new_n8829_), .ZN(new_n9059_));
  NAND2_X1   g08866(.A1(new_n9059_), .A2(new_n9058_), .ZN(new_n9060_));
  NAND2_X1   g08867(.A1(new_n8747_), .A2(new_n8740_), .ZN(new_n9061_));
  INV_X1     g08868(.I(new_n8756_), .ZN(new_n9062_));
  OAI21_X1   g08869(.A1(new_n8748_), .A2(new_n9062_), .B(new_n9061_), .ZN(new_n9063_));
  NOR2_X1    g08870(.A1(new_n8898_), .A2(new_n8895_), .ZN(new_n9064_));
  INV_X1     g08871(.I(new_n9064_), .ZN(new_n9065_));
  NOR2_X1    g08872(.A1(new_n9065_), .A2(new_n9063_), .ZN(new_n9066_));
  NAND2_X1   g08873(.A1(new_n9065_), .A2(new_n9063_), .ZN(new_n9067_));
  INV_X1     g08874(.I(new_n9067_), .ZN(new_n9068_));
  NOR2_X1    g08875(.A1(new_n9068_), .A2(new_n9066_), .ZN(new_n9069_));
  NAND2_X1   g08876(.A1(new_n9069_), .A2(new_n9060_), .ZN(new_n9070_));
  INV_X1     g08877(.I(new_n9070_), .ZN(new_n9071_));
  NOR2_X1    g08878(.A1(new_n9069_), .A2(new_n9060_), .ZN(new_n9072_));
  NOR2_X1    g08879(.A1(new_n9071_), .A2(new_n9072_), .ZN(new_n9073_));
  INV_X1     g08880(.I(new_n9073_), .ZN(new_n9074_));
  NOR2_X1    g08881(.A1(new_n8836_), .A2(new_n9074_), .ZN(new_n9075_));
  NOR2_X1    g08882(.A1(new_n8835_), .A2(new_n9073_), .ZN(new_n9076_));
  NOR2_X1    g08883(.A1(new_n9075_), .A2(new_n9076_), .ZN(new_n9077_));
  NOR2_X1    g08884(.A1(new_n9077_), .A2(new_n9057_), .ZN(new_n9078_));
  NAND2_X1   g08885(.A1(new_n9077_), .A2(new_n9057_), .ZN(new_n9079_));
  INV_X1     g08886(.I(new_n9079_), .ZN(new_n9080_));
  NOR2_X1    g08887(.A1(new_n9080_), .A2(new_n9078_), .ZN(new_n9081_));
  XOR2_X1    g08888(.A1(new_n9045_), .A2(new_n9081_), .Z(new_n9082_));
  XNOR2_X1   g08889(.A1(new_n9082_), .A2(new_n9042_), .ZN(new_n9083_));
  NAND2_X1   g08890(.A1(new_n8841_), .A2(new_n8875_), .ZN(new_n9084_));
  OAI21_X1   g08891(.A1(new_n8876_), .A2(new_n8838_), .B(new_n9084_), .ZN(new_n9085_));
  INV_X1     g08892(.I(new_n8778_), .ZN(new_n9086_));
  OAI21_X1   g08893(.A1(new_n9086_), .A2(new_n8837_), .B(new_n8777_), .ZN(new_n9087_));
  NAND2_X1   g08894(.A1(new_n8771_), .A2(new_n8769_), .ZN(new_n9088_));
  NAND2_X1   g08895(.A1(new_n8772_), .A2(new_n8758_), .ZN(new_n9089_));
  NAND2_X1   g08896(.A1(new_n9089_), .A2(new_n9088_), .ZN(new_n9090_));
  NOR2_X1    g08897(.A1(new_n8849_), .A2(new_n8846_), .ZN(new_n9091_));
  NAND2_X1   g08898(.A1(new_n8598_), .A2(new_n8636_), .ZN(new_n9092_));
  NAND2_X1   g08899(.A1(new_n8759_), .A2(new_n8768_), .ZN(new_n9093_));
  NAND2_X1   g08900(.A1(new_n9093_), .A2(new_n9092_), .ZN(new_n9094_));
  XOR2_X1    g08901(.A1(new_n9094_), .A2(new_n8858_), .Z(new_n9095_));
  XNOR2_X1   g08902(.A1(new_n9095_), .A2(new_n9091_), .ZN(new_n9096_));
  INV_X1     g08903(.I(new_n8852_), .ZN(new_n9097_));
  INV_X1     g08904(.I(new_n8861_), .ZN(new_n9098_));
  NAND2_X1   g08905(.A1(new_n9098_), .A2(new_n8844_), .ZN(new_n9099_));
  OAI21_X1   g08906(.A1(new_n9097_), .A2(new_n8860_), .B(new_n9099_), .ZN(new_n9100_));
  XOR2_X1    g08907(.A1(new_n9100_), .A2(new_n9096_), .Z(new_n9101_));
  XOR2_X1    g08908(.A1(new_n9101_), .A2(new_n9090_), .Z(new_n9102_));
  NAND2_X1   g08909(.A1(new_n8863_), .A2(new_n8873_), .ZN(new_n9103_));
  NAND2_X1   g08910(.A1(new_n8874_), .A2(new_n8862_), .ZN(new_n9104_));
  NAND2_X1   g08911(.A1(new_n9104_), .A2(new_n9103_), .ZN(new_n9105_));
  NAND2_X1   g08912(.A1(new_n9105_), .A2(new_n9102_), .ZN(new_n9106_));
  INV_X1     g08913(.I(new_n9106_), .ZN(new_n9107_));
  NOR2_X1    g08914(.A1(new_n9105_), .A2(new_n9102_), .ZN(new_n9108_));
  NOR2_X1    g08915(.A1(new_n9107_), .A2(new_n9108_), .ZN(new_n9109_));
  NOR2_X1    g08916(.A1(new_n9087_), .A2(new_n9109_), .ZN(new_n9110_));
  AND2_X2    g08917(.A1(new_n9087_), .A2(new_n9109_), .Z(new_n9111_));
  NOR2_X1    g08918(.A1(new_n9111_), .A2(new_n9110_), .ZN(new_n9112_));
  XOR2_X1    g08919(.A1(new_n9085_), .A2(new_n9112_), .Z(new_n9113_));
  XOR2_X1    g08920(.A1(new_n9113_), .A2(new_n9083_), .Z(new_n9114_));
  INV_X1     g08921(.I(new_n9114_), .ZN(new_n9115_));
  NOR2_X1    g08922(.A1(new_n8940_), .A2(new_n9115_), .ZN(new_n9116_));
  NOR2_X1    g08923(.A1(new_n8939_), .A2(new_n9114_), .ZN(new_n9117_));
  NOR2_X1    g08924(.A1(new_n9116_), .A2(new_n9117_), .ZN(new_n9118_));
  XOR2_X1    g08925(.A1(new_n8938_), .A2(new_n9118_), .Z(\asquared[72] ));
  NOR2_X1    g08926(.A1(new_n9111_), .A2(new_n9107_), .ZN(new_n9120_));
  NAND2_X1   g08927(.A1(new_n8958_), .A2(new_n8965_), .ZN(new_n9121_));
  INV_X1     g08928(.I(new_n9121_), .ZN(new_n9122_));
  AOI21_X1   g08929(.A1(new_n8966_), .A2(new_n8949_), .B(new_n9122_), .ZN(new_n9123_));
  XOR2_X1    g08930(.A1(new_n8989_), .A2(new_n8973_), .Z(new_n9124_));
  XOR2_X1    g08931(.A1(new_n9124_), .A2(new_n8981_), .Z(new_n9125_));
  XOR2_X1    g08932(.A1(new_n9021_), .A2(new_n9003_), .Z(new_n9126_));
  XOR2_X1    g08933(.A1(new_n9126_), .A2(new_n9011_), .Z(new_n9127_));
  NAND2_X1   g08934(.A1(new_n9125_), .A2(new_n9127_), .ZN(new_n9128_));
  INV_X1     g08935(.I(new_n9128_), .ZN(new_n9129_));
  NOR2_X1    g08936(.A1(new_n9125_), .A2(new_n9127_), .ZN(new_n9130_));
  NOR2_X1    g08937(.A1(new_n9129_), .A2(new_n9130_), .ZN(new_n9131_));
  XNOR2_X1   g08938(.A1(new_n9131_), .A2(new_n9123_), .ZN(new_n9132_));
  INV_X1     g08939(.I(new_n8992_), .ZN(new_n9133_));
  NAND2_X1   g08940(.A1(new_n9133_), .A2(new_n8967_), .ZN(new_n9134_));
  NAND2_X1   g08941(.A1(new_n8943_), .A2(new_n8993_), .ZN(new_n9135_));
  NAND2_X1   g08942(.A1(new_n9135_), .A2(new_n9134_), .ZN(new_n9136_));
  NAND2_X1   g08943(.A1(new_n9012_), .A2(new_n9004_), .ZN(new_n9137_));
  NAND2_X1   g08944(.A1(new_n9013_), .A2(new_n9022_), .ZN(new_n9138_));
  NAND2_X1   g08945(.A1(new_n9138_), .A2(new_n9137_), .ZN(new_n9139_));
  NAND2_X1   g08946(.A1(new_n8739_), .A2(new_n8754_), .ZN(new_n9140_));
  NAND2_X1   g08947(.A1(new_n9049_), .A2(new_n8819_), .ZN(new_n9141_));
  NAND2_X1   g08948(.A1(new_n9141_), .A2(new_n9140_), .ZN(new_n9142_));
  NAND2_X1   g08949(.A1(new_n8975_), .A2(new_n8982_), .ZN(new_n9143_));
  INV_X1     g08950(.I(new_n8991_), .ZN(new_n9144_));
  OAI21_X1   g08951(.A1(new_n8983_), .A2(new_n9144_), .B(new_n9143_), .ZN(new_n9145_));
  XOR2_X1    g08952(.A1(new_n9145_), .A2(new_n9142_), .Z(new_n9146_));
  XOR2_X1    g08953(.A1(new_n9146_), .A2(new_n9139_), .Z(new_n9147_));
  XOR2_X1    g08954(.A1(new_n9136_), .A2(new_n9147_), .Z(new_n9148_));
  XOR2_X1    g08955(.A1(new_n9148_), .A2(new_n9132_), .Z(new_n9149_));
  XNOR2_X1   g08956(.A1(new_n9120_), .A2(new_n9149_), .ZN(new_n9150_));
  NOR2_X1    g08957(.A1(new_n9071_), .A2(new_n9068_), .ZN(new_n9151_));
  INV_X1     g08958(.I(new_n9151_), .ZN(new_n9152_));
  AOI22_X1   g08959(.A1(\a[16] ), .A2(\a[56] ), .B1(\a[23] ), .B2(\a[49] ), .ZN(new_n9153_));
  INV_X1     g08960(.I(new_n9153_), .ZN(new_n9154_));
  NOR4_X1    g08961(.A1(new_n742_), .A2(new_n1299_), .A3(new_n4702_), .A4(new_n5856_), .ZN(new_n9155_));
  NOR2_X1    g08962(.A1(new_n2200_), .A2(new_n3221_), .ZN(new_n9156_));
  AOI21_X1   g08963(.A1(new_n9154_), .A2(new_n9156_), .B(new_n9155_), .ZN(new_n9157_));
  INV_X1     g08964(.I(new_n9157_), .ZN(new_n9158_));
  OAI21_X1   g08965(.A1(new_n9155_), .A2(new_n9153_), .B(new_n9156_), .ZN(new_n9159_));
  OAI21_X1   g08966(.A1(new_n9158_), .A2(new_n9153_), .B(new_n9159_), .ZN(new_n9160_));
  OAI22_X1   g08967(.A1(new_n1220_), .A2(new_n5135_), .B1(new_n1175_), .B2(new_n4901_), .ZN(new_n9161_));
  NAND2_X1   g08968(.A1(new_n1452_), .A2(new_n5439_), .ZN(new_n9162_));
  NAND3_X1   g08969(.A1(new_n9162_), .A2(new_n4189_), .A3(new_n9161_), .ZN(new_n9163_));
  NAND2_X1   g08970(.A1(new_n9163_), .A2(new_n4189_), .ZN(new_n9164_));
  NAND3_X1   g08971(.A1(new_n9162_), .A2(new_n4190_), .A3(new_n9161_), .ZN(new_n9165_));
  NAND2_X1   g08972(.A1(new_n9164_), .A2(new_n9165_), .ZN(new_n9166_));
  XOR2_X1    g08973(.A1(new_n9166_), .A2(new_n9160_), .Z(new_n9167_));
  NAND2_X1   g08974(.A1(\a[17] ), .A2(\a[55] ), .ZN(new_n9168_));
  NAND4_X1   g08975(.A1(\a[17] ), .A2(\a[20] ), .A3(\a[52] ), .A4(\a[55] ), .ZN(new_n9169_));
  NAND2_X1   g08976(.A1(new_n1027_), .A2(new_n6128_), .ZN(new_n9170_));
  AOI22_X1   g08977(.A1(new_n9170_), .A2(new_n9169_), .B1(new_n1273_), .B2(new_n8420_), .ZN(new_n9171_));
  AOI22_X1   g08978(.A1(\a[18] ), .A2(\a[54] ), .B1(\a[20] ), .B2(\a[52] ), .ZN(new_n9172_));
  NAND2_X1   g08979(.A1(new_n1273_), .A2(new_n8420_), .ZN(new_n9173_));
  NAND3_X1   g08980(.A1(new_n9173_), .A2(new_n9170_), .A3(new_n9169_), .ZN(new_n9174_));
  OAI22_X1   g08981(.A1(new_n9171_), .A2(new_n9168_), .B1(new_n9174_), .B2(new_n9172_), .ZN(new_n9175_));
  XNOR2_X1   g08982(.A1(new_n9167_), .A2(new_n9175_), .ZN(new_n9176_));
  OAI22_X1   g08983(.A1(new_n539_), .A2(new_n8049_), .B1(new_n7959_), .B2(new_n1063_), .ZN(new_n9177_));
  OAI21_X1   g08984(.A1(new_n1264_), .A2(new_n7591_), .B(new_n9177_), .ZN(new_n9178_));
  NAND3_X1   g08985(.A1(new_n9178_), .A2(\a[9] ), .A3(\a[63] ), .ZN(new_n9179_));
  AOI22_X1   g08986(.A1(\a[10] ), .A2(\a[62] ), .B1(\a[11] ), .B2(\a[61] ), .ZN(new_n9180_));
  NOR2_X1    g08987(.A1(new_n1264_), .A2(new_n7591_), .ZN(new_n9181_));
  NOR2_X1    g08988(.A1(new_n9177_), .A2(new_n9181_), .ZN(new_n9182_));
  INV_X1     g08989(.I(new_n9182_), .ZN(new_n9183_));
  OAI21_X1   g08990(.A1(new_n9180_), .A2(new_n9183_), .B(new_n9179_), .ZN(new_n9184_));
  AOI22_X1   g08991(.A1(\a[24] ), .A2(\a[48] ), .B1(\a[25] ), .B2(\a[47] ), .ZN(new_n9185_));
  NOR2_X1    g08992(.A1(new_n536_), .A2(new_n6723_), .ZN(new_n9186_));
  INV_X1     g08993(.I(new_n9186_), .ZN(new_n9187_));
  NOR2_X1    g08994(.A1(new_n1779_), .A2(new_n4977_), .ZN(new_n9188_));
  NOR3_X1    g08995(.A1(new_n9188_), .A2(new_n9185_), .A3(new_n9187_), .ZN(new_n9189_));
  NOR2_X1    g08996(.A1(new_n9189_), .A2(new_n9188_), .ZN(new_n9190_));
  INV_X1     g08997(.I(new_n9190_), .ZN(new_n9191_));
  OAI22_X1   g08998(.A1(new_n9191_), .A2(new_n9185_), .B1(new_n9187_), .B2(new_n9189_), .ZN(new_n9192_));
  INV_X1     g08999(.I(new_n9192_), .ZN(new_n9193_));
  OAI21_X1   g09000(.A1(new_n8948_), .A2(new_n8827_), .B(new_n8945_), .ZN(new_n9194_));
  NOR2_X1    g09001(.A1(new_n9193_), .A2(new_n9194_), .ZN(new_n9195_));
  INV_X1     g09002(.I(new_n9194_), .ZN(new_n9196_));
  NOR2_X1    g09003(.A1(new_n9192_), .A2(new_n9196_), .ZN(new_n9197_));
  OAI21_X1   g09004(.A1(new_n9195_), .A2(new_n9197_), .B(new_n9184_), .ZN(new_n9198_));
  OR3_X2     g09005(.A1(new_n9195_), .A2(new_n9184_), .A3(new_n9197_), .Z(new_n9199_));
  NAND2_X1   g09006(.A1(new_n9199_), .A2(new_n9198_), .ZN(new_n9200_));
  XOR2_X1    g09007(.A1(new_n9200_), .A2(new_n9176_), .Z(new_n9201_));
  NOR2_X1    g09008(.A1(new_n9152_), .A2(new_n9201_), .ZN(new_n9202_));
  NAND2_X1   g09009(.A1(new_n9152_), .A2(new_n9201_), .ZN(new_n9203_));
  INV_X1     g09010(.I(new_n9203_), .ZN(new_n9204_));
  NOR2_X1    g09011(.A1(new_n9204_), .A2(new_n9202_), .ZN(new_n9205_));
  NAND2_X1   g09012(.A1(new_n9100_), .A2(new_n9096_), .ZN(new_n9206_));
  NAND2_X1   g09013(.A1(new_n9101_), .A2(new_n9090_), .ZN(new_n9207_));
  NAND2_X1   g09014(.A1(new_n9207_), .A2(new_n9206_), .ZN(new_n9208_));
  NAND2_X1   g09015(.A1(new_n897_), .A2(new_n6803_), .ZN(new_n9209_));
  OAI22_X1   g09016(.A1(new_n767_), .A2(new_n7206_), .B1(new_n7204_), .B2(new_n836_), .ZN(new_n9210_));
  NAND2_X1   g09017(.A1(new_n9210_), .A2(new_n9209_), .ZN(new_n9211_));
  NAND3_X1   g09018(.A1(new_n9211_), .A2(\a[13] ), .A3(\a[59] ), .ZN(new_n9212_));
  AOI22_X1   g09019(.A1(\a[14] ), .A2(\a[58] ), .B1(\a[15] ), .B2(\a[57] ), .ZN(new_n9213_));
  NAND2_X1   g09020(.A1(new_n9211_), .A2(new_n9209_), .ZN(new_n9214_));
  OAI21_X1   g09021(.A1(new_n9213_), .A2(new_n9214_), .B(new_n9212_), .ZN(new_n9215_));
  NAND2_X1   g09022(.A1(new_n2103_), .A2(new_n4703_), .ZN(new_n9216_));
  OAI22_X1   g09023(.A1(new_n1972_), .A2(new_n4430_), .B1(new_n3341_), .B2(new_n6101_), .ZN(new_n9217_));
  NAND2_X1   g09024(.A1(new_n9217_), .A2(new_n9216_), .ZN(new_n9218_));
  NAND3_X1   g09025(.A1(new_n9218_), .A2(\a[26] ), .A3(\a[46] ), .ZN(new_n9219_));
  AOI22_X1   g09026(.A1(\a[27] ), .A2(\a[45] ), .B1(\a[28] ), .B2(\a[44] ), .ZN(new_n9220_));
  NAND2_X1   g09027(.A1(new_n9218_), .A2(new_n9216_), .ZN(new_n9221_));
  OAI21_X1   g09028(.A1(new_n9220_), .A2(new_n9221_), .B(new_n9219_), .ZN(new_n9222_));
  XOR2_X1    g09029(.A1(new_n9222_), .A2(new_n9215_), .Z(new_n9223_));
  AOI22_X1   g09030(.A1(\a[33] ), .A2(\a[39] ), .B1(\a[34] ), .B2(\a[38] ), .ZN(new_n9224_));
  NAND2_X1   g09031(.A1(\a[19] ), .A2(\a[53] ), .ZN(new_n9225_));
  NOR2_X1    g09032(.A1(new_n3932_), .A2(new_n4210_), .ZN(new_n9226_));
  NOR3_X1    g09033(.A1(new_n9226_), .A2(new_n9224_), .A3(new_n9225_), .ZN(new_n9227_));
  OAI22_X1   g09034(.A1(new_n3932_), .A2(new_n4210_), .B1(new_n9224_), .B2(new_n9225_), .ZN(new_n9228_));
  OAI22_X1   g09035(.A1(new_n9227_), .A2(new_n9225_), .B1(new_n9224_), .B2(new_n9228_), .ZN(new_n9229_));
  XOR2_X1    g09036(.A1(new_n9223_), .A2(new_n9229_), .Z(new_n9230_));
  NAND2_X1   g09037(.A1(new_n9094_), .A2(new_n8858_), .ZN(new_n9231_));
  INV_X1     g09038(.I(new_n9095_), .ZN(new_n9232_));
  OAI21_X1   g09039(.A1(new_n9232_), .A2(new_n9091_), .B(new_n9231_), .ZN(new_n9233_));
  XOR2_X1    g09040(.A1(new_n8957_), .A2(new_n8964_), .Z(new_n9234_));
  XOR2_X1    g09041(.A1(new_n9234_), .A2(new_n9036_), .Z(new_n9235_));
  XOR2_X1    g09042(.A1(new_n9233_), .A2(new_n9235_), .Z(new_n9236_));
  XOR2_X1    g09043(.A1(new_n9236_), .A2(new_n9230_), .Z(new_n9237_));
  XOR2_X1    g09044(.A1(new_n9208_), .A2(new_n9237_), .Z(new_n9238_));
  XNOR2_X1   g09045(.A1(new_n9238_), .A2(new_n9205_), .ZN(new_n9239_));
  XOR2_X1    g09046(.A1(new_n9150_), .A2(new_n9239_), .Z(new_n9240_));
  INV_X1     g09047(.I(new_n9240_), .ZN(new_n9241_));
  NAND2_X1   g09048(.A1(new_n9045_), .A2(new_n9081_), .ZN(new_n9242_));
  INV_X1     g09049(.I(new_n9082_), .ZN(new_n9243_));
  OAI21_X1   g09050(.A1(new_n9243_), .A2(new_n9042_), .B(new_n9242_), .ZN(new_n9244_));
  NAND2_X1   g09051(.A1(new_n8997_), .A2(new_n9040_), .ZN(new_n9245_));
  NAND2_X1   g09052(.A1(new_n9041_), .A2(new_n8994_), .ZN(new_n9246_));
  NAND2_X1   g09053(.A1(new_n9246_), .A2(new_n9245_), .ZN(new_n9247_));
  NOR2_X1    g09054(.A1(new_n9080_), .A2(new_n9075_), .ZN(new_n9248_));
  NAND2_X1   g09055(.A1(new_n9026_), .A2(new_n9038_), .ZN(new_n9249_));
  NAND2_X1   g09056(.A1(new_n9039_), .A2(new_n9023_), .ZN(new_n9250_));
  NAND2_X1   g09057(.A1(new_n9250_), .A2(new_n9249_), .ZN(new_n9251_));
  NAND2_X1   g09058(.A1(new_n9050_), .A2(new_n9055_), .ZN(new_n9252_));
  NAND2_X1   g09059(.A1(new_n9056_), .A2(new_n9048_), .ZN(new_n9253_));
  NAND2_X1   g09060(.A1(new_n9253_), .A2(new_n9252_), .ZN(new_n9254_));
  NOR2_X1    g09061(.A1(new_n8789_), .A2(new_n8807_), .ZN(new_n9255_));
  NOR2_X1    g09062(.A1(new_n9053_), .A2(new_n9255_), .ZN(new_n9256_));
  NAND2_X1   g09063(.A1(new_n2976_), .A2(new_n4028_), .ZN(new_n9257_));
  NAND2_X1   g09064(.A1(new_n2254_), .A2(new_n4180_), .ZN(new_n9258_));
  AOI22_X1   g09065(.A1(new_n9257_), .A2(new_n9258_), .B1(new_n2437_), .B2(new_n4372_), .ZN(new_n9259_));
  NAND2_X1   g09066(.A1(\a[29] ), .A2(\a[43] ), .ZN(new_n9260_));
  AOI22_X1   g09067(.A1(\a[30] ), .A2(\a[42] ), .B1(\a[31] ), .B2(\a[41] ), .ZN(new_n9261_));
  NAND2_X1   g09068(.A1(new_n2437_), .A2(new_n4372_), .ZN(new_n9262_));
  NAND3_X1   g09069(.A1(new_n9262_), .A2(new_n9257_), .A3(new_n9258_), .ZN(new_n9263_));
  OAI22_X1   g09070(.A1(new_n9259_), .A2(new_n9260_), .B1(new_n9263_), .B2(new_n9261_), .ZN(new_n9264_));
  NAND2_X1   g09071(.A1(new_n8765_), .A2(new_n8746_), .ZN(new_n9265_));
  NAND2_X1   g09072(.A1(new_n9027_), .A2(new_n9037_), .ZN(new_n9266_));
  NAND2_X1   g09073(.A1(new_n9266_), .A2(new_n9265_), .ZN(new_n9267_));
  XNOR2_X1   g09074(.A1(new_n9267_), .A2(new_n9264_), .ZN(new_n9268_));
  XOR2_X1    g09075(.A1(new_n9268_), .A2(new_n9256_), .Z(new_n9269_));
  XOR2_X1    g09076(.A1(new_n9269_), .A2(new_n9254_), .Z(new_n9270_));
  XOR2_X1    g09077(.A1(new_n9251_), .A2(new_n9270_), .Z(new_n9271_));
  INV_X1     g09078(.I(new_n9271_), .ZN(new_n9272_));
  XOR2_X1    g09079(.A1(new_n9248_), .A2(new_n9272_), .Z(new_n9273_));
  XOR2_X1    g09080(.A1(new_n9273_), .A2(new_n9247_), .Z(new_n9274_));
  NOR2_X1    g09081(.A1(new_n9244_), .A2(new_n9274_), .ZN(new_n9275_));
  NAND2_X1   g09082(.A1(new_n9244_), .A2(new_n9274_), .ZN(new_n9276_));
  INV_X1     g09083(.I(new_n9276_), .ZN(new_n9277_));
  NOR2_X1    g09084(.A1(new_n9277_), .A2(new_n9275_), .ZN(new_n9278_));
  NAND2_X1   g09085(.A1(new_n9241_), .A2(new_n9278_), .ZN(new_n9279_));
  INV_X1     g09086(.I(new_n9279_), .ZN(new_n9280_));
  NOR2_X1    g09087(.A1(new_n9241_), .A2(new_n9278_), .ZN(new_n9281_));
  NOR2_X1    g09088(.A1(new_n9280_), .A2(new_n9281_), .ZN(new_n9282_));
  INV_X1     g09089(.I(new_n9282_), .ZN(new_n9283_));
  NAND2_X1   g09090(.A1(new_n9085_), .A2(new_n9112_), .ZN(new_n9284_));
  NAND2_X1   g09091(.A1(new_n9113_), .A2(new_n9083_), .ZN(new_n9285_));
  NAND2_X1   g09092(.A1(new_n9285_), .A2(new_n9284_), .ZN(new_n9286_));
  INV_X1     g09093(.I(new_n9286_), .ZN(new_n9287_));
  NOR2_X1    g09094(.A1(new_n9287_), .A2(new_n9283_), .ZN(new_n9288_));
  INV_X1     g09095(.I(new_n9288_), .ZN(new_n9289_));
  AOI21_X1   g09096(.A1(new_n8937_), .A2(new_n8920_), .B(new_n9117_), .ZN(new_n9290_));
  NOR2_X1    g09097(.A1(new_n9290_), .A2(new_n9116_), .ZN(new_n9291_));
  INV_X1     g09098(.I(new_n9116_), .ZN(new_n9292_));
  INV_X1     g09099(.I(new_n9117_), .ZN(new_n9293_));
  OAI21_X1   g09100(.A1(new_n8934_), .A2(new_n8919_), .B(new_n9293_), .ZN(new_n9294_));
  NOR2_X1    g09101(.A1(new_n9286_), .A2(new_n9282_), .ZN(new_n9295_));
  AOI21_X1   g09102(.A1(new_n9294_), .A2(new_n9292_), .B(new_n9295_), .ZN(new_n9296_));
  INV_X1     g09103(.I(new_n9295_), .ZN(new_n9297_));
  NAND2_X1   g09104(.A1(new_n9289_), .A2(new_n9297_), .ZN(new_n9298_));
  AOI22_X1   g09105(.A1(new_n9296_), .A2(new_n9289_), .B1(new_n9291_), .B2(new_n9298_), .ZN(\asquared[73] ));
  OAI21_X1   g09106(.A1(new_n9290_), .A2(new_n9116_), .B(new_n9297_), .ZN(new_n9300_));
  NAND2_X1   g09107(.A1(new_n9300_), .A2(new_n9289_), .ZN(new_n9301_));
  NOR2_X1    g09108(.A1(new_n9280_), .A2(new_n9277_), .ZN(new_n9302_));
  INV_X1     g09109(.I(new_n9302_), .ZN(new_n9303_));
  NAND2_X1   g09110(.A1(new_n9273_), .A2(new_n9247_), .ZN(new_n9304_));
  OAI21_X1   g09111(.A1(new_n9248_), .A2(new_n9272_), .B(new_n9304_), .ZN(new_n9305_));
  NAND2_X1   g09112(.A1(new_n9166_), .A2(new_n9160_), .ZN(new_n9306_));
  NAND2_X1   g09113(.A1(new_n9167_), .A2(new_n9175_), .ZN(new_n9307_));
  NAND2_X1   g09114(.A1(new_n9307_), .A2(new_n9306_), .ZN(new_n9308_));
  XOR2_X1    g09115(.A1(new_n9190_), .A2(new_n9182_), .Z(new_n9309_));
  XOR2_X1    g09116(.A1(new_n9309_), .A2(new_n9174_), .Z(new_n9310_));
  NAND2_X1   g09117(.A1(new_n9163_), .A2(new_n9162_), .ZN(new_n9311_));
  NOR2_X1    g09118(.A1(new_n597_), .A2(new_n6723_), .ZN(new_n9312_));
  XOR2_X1    g09119(.A1(new_n9311_), .A2(new_n9312_), .Z(new_n9313_));
  XOR2_X1    g09120(.A1(new_n9313_), .A2(new_n9228_), .Z(new_n9314_));
  XOR2_X1    g09121(.A1(new_n9310_), .A2(new_n9314_), .Z(new_n9315_));
  XOR2_X1    g09122(.A1(new_n9315_), .A2(new_n9308_), .Z(new_n9316_));
  NOR2_X1    g09123(.A1(new_n9200_), .A2(new_n9176_), .ZN(new_n9317_));
  NOR2_X1    g09124(.A1(new_n9204_), .A2(new_n9317_), .ZN(new_n9318_));
  NAND2_X1   g09125(.A1(new_n9222_), .A2(new_n9215_), .ZN(new_n9319_));
  NAND2_X1   g09126(.A1(new_n9223_), .A2(new_n9229_), .ZN(new_n9320_));
  NAND2_X1   g09127(.A1(new_n9320_), .A2(new_n9319_), .ZN(new_n9321_));
  OAI21_X1   g09128(.A1(new_n9193_), .A2(new_n9196_), .B(new_n9198_), .ZN(new_n9322_));
  NAND2_X1   g09129(.A1(new_n9021_), .A2(new_n9003_), .ZN(new_n9323_));
  NAND2_X1   g09130(.A1(new_n9126_), .A2(new_n9011_), .ZN(new_n9324_));
  NAND2_X1   g09131(.A1(new_n9324_), .A2(new_n9323_), .ZN(new_n9325_));
  XOR2_X1    g09132(.A1(new_n9322_), .A2(new_n9325_), .Z(new_n9326_));
  XOR2_X1    g09133(.A1(new_n9326_), .A2(new_n9321_), .Z(new_n9327_));
  INV_X1     g09134(.I(new_n9327_), .ZN(new_n9328_));
  NAND2_X1   g09135(.A1(new_n9318_), .A2(new_n9328_), .ZN(new_n9329_));
  OAI21_X1   g09136(.A1(new_n9204_), .A2(new_n9317_), .B(new_n9327_), .ZN(new_n9330_));
  AND2_X2    g09137(.A1(new_n9329_), .A2(new_n9330_), .Z(new_n9331_));
  XOR2_X1    g09138(.A1(new_n9331_), .A2(new_n9316_), .Z(new_n9332_));
  XOR2_X1    g09139(.A1(new_n9305_), .A2(new_n9332_), .Z(new_n9333_));
  NAND2_X1   g09140(.A1(new_n9145_), .A2(new_n9142_), .ZN(new_n9334_));
  NAND2_X1   g09141(.A1(new_n9146_), .A2(new_n9139_), .ZN(new_n9335_));
  NAND2_X1   g09142(.A1(new_n9335_), .A2(new_n9334_), .ZN(new_n9336_));
  AOI22_X1   g09143(.A1(\a[26] ), .A2(\a[47] ), .B1(\a[27] ), .B2(\a[46] ), .ZN(new_n9337_));
  INV_X1     g09144(.I(new_n9337_), .ZN(new_n9338_));
  NOR2_X1    g09145(.A1(new_n1972_), .A2(new_n4721_), .ZN(new_n9339_));
  NOR2_X1    g09146(.A1(new_n1023_), .A2(new_n5856_), .ZN(new_n9340_));
  AOI21_X1   g09147(.A1(new_n9338_), .A2(new_n9340_), .B(new_n9339_), .ZN(new_n9341_));
  NAND2_X1   g09148(.A1(new_n9341_), .A2(new_n9338_), .ZN(new_n9342_));
  OAI21_X1   g09149(.A1(new_n9339_), .A2(new_n9337_), .B(new_n9340_), .ZN(new_n9343_));
  NAND2_X1   g09150(.A1(new_n9342_), .A2(new_n9343_), .ZN(new_n9344_));
  XOR2_X1    g09151(.A1(new_n9344_), .A2(new_n9158_), .Z(new_n9345_));
  NOR2_X1    g09152(.A1(new_n6804_), .A2(new_n893_), .ZN(new_n9346_));
  AOI22_X1   g09153(.A1(new_n895_), .A2(new_n7203_), .B1(new_n897_), .B2(new_n7205_), .ZN(new_n9347_));
  NOR2_X1    g09154(.A1(new_n9347_), .A2(new_n9346_), .ZN(new_n9348_));
  NAND2_X1   g09155(.A1(\a[14] ), .A2(\a[59] ), .ZN(new_n9349_));
  AOI22_X1   g09156(.A1(\a[15] ), .A2(\a[58] ), .B1(\a[16] ), .B2(\a[57] ), .ZN(new_n9350_));
  NOR2_X1    g09157(.A1(new_n9348_), .A2(new_n9346_), .ZN(new_n9351_));
  INV_X1     g09158(.I(new_n9351_), .ZN(new_n9352_));
  OAI22_X1   g09159(.A1(new_n9352_), .A2(new_n9350_), .B1(new_n9348_), .B2(new_n9349_), .ZN(new_n9353_));
  XNOR2_X1   g09160(.A1(new_n9345_), .A2(new_n9353_), .ZN(new_n9354_));
  AOI21_X1   g09161(.A1(\a[11] ), .A2(\a[62] ), .B(\a[37] ), .ZN(new_n9355_));
  NAND2_X1   g09162(.A1(\a[23] ), .A2(\a[50] ), .ZN(new_n9356_));
  NOR2_X1    g09163(.A1(new_n3800_), .A2(new_n7144_), .ZN(new_n9357_));
  NOR3_X1    g09164(.A1(new_n9357_), .A2(new_n9355_), .A3(new_n9356_), .ZN(new_n9358_));
  OAI22_X1   g09165(.A1(new_n3800_), .A2(new_n7144_), .B1(new_n9355_), .B2(new_n9356_), .ZN(new_n9359_));
  OAI22_X1   g09166(.A1(new_n9358_), .A2(new_n9356_), .B1(new_n9355_), .B2(new_n9359_), .ZN(new_n9360_));
  NOR4_X1    g09167(.A1(new_n979_), .A2(new_n1357_), .A3(new_n4702_), .A4(new_n5617_), .ZN(new_n9361_));
  INV_X1     g09168(.I(new_n9361_), .ZN(new_n9362_));
  NOR3_X1    g09169(.A1(new_n7659_), .A2(new_n884_), .A3(new_n1357_), .ZN(new_n9363_));
  NOR2_X1    g09170(.A1(new_n6129_), .A2(new_n1092_), .ZN(new_n9364_));
  OAI21_X1   g09171(.A1(new_n9363_), .A2(new_n9364_), .B(new_n9362_), .ZN(new_n9365_));
  NAND3_X1   g09172(.A1(new_n9365_), .A2(\a[18] ), .A3(\a[55] ), .ZN(new_n9366_));
  NAND2_X1   g09173(.A1(new_n9365_), .A2(new_n9362_), .ZN(new_n9367_));
  AOI22_X1   g09174(.A1(\a[19] ), .A2(\a[54] ), .B1(\a[24] ), .B2(\a[49] ), .ZN(new_n9368_));
  OAI21_X1   g09175(.A1(new_n9367_), .A2(new_n9368_), .B(new_n9366_), .ZN(new_n9369_));
  XNOR2_X1   g09176(.A1(new_n9369_), .A2(new_n9360_), .ZN(new_n9370_));
  AOI22_X1   g09177(.A1(new_n1452_), .A2(new_n5524_), .B1(new_n1552_), .B2(new_n5682_), .ZN(new_n9371_));
  AOI21_X1   g09178(.A1(new_n1381_), .A2(new_n5862_), .B(new_n9371_), .ZN(new_n9372_));
  NAND2_X1   g09179(.A1(\a[22] ), .A2(\a[51] ), .ZN(new_n9373_));
  AOI22_X1   g09180(.A1(\a[20] ), .A2(\a[53] ), .B1(\a[21] ), .B2(\a[52] ), .ZN(new_n9374_));
  OAI21_X1   g09181(.A1(new_n1382_), .A2(new_n6563_), .B(new_n9371_), .ZN(new_n9375_));
  OAI22_X1   g09182(.A1(new_n9372_), .A2(new_n9373_), .B1(new_n9375_), .B2(new_n9374_), .ZN(new_n9376_));
  XOR2_X1    g09183(.A1(new_n9370_), .A2(new_n9376_), .Z(new_n9377_));
  XOR2_X1    g09184(.A1(new_n9377_), .A2(new_n9354_), .Z(new_n9378_));
  XOR2_X1    g09185(.A1(new_n9336_), .A2(new_n9378_), .Z(new_n9379_));
  NAND2_X1   g09186(.A1(new_n9269_), .A2(new_n9254_), .ZN(new_n9380_));
  NAND2_X1   g09187(.A1(new_n9251_), .A2(new_n9270_), .ZN(new_n9381_));
  NAND2_X1   g09188(.A1(new_n9381_), .A2(new_n9380_), .ZN(new_n9382_));
  AOI22_X1   g09189(.A1(\a[10] ), .A2(\a[63] ), .B1(\a[12] ), .B2(\a[61] ), .ZN(new_n9383_));
  NOR2_X1    g09190(.A1(new_n1441_), .A2(new_n4596_), .ZN(new_n9384_));
  INV_X1     g09191(.I(new_n9384_), .ZN(new_n9385_));
  OAI22_X1   g09192(.A1(new_n534_), .A2(new_n7959_), .B1(new_n9385_), .B2(new_n9383_), .ZN(new_n9386_));
  NOR2_X1    g09193(.A1(new_n7959_), .A2(new_n534_), .ZN(new_n9387_));
  OAI21_X1   g09194(.A1(new_n9387_), .A2(new_n9383_), .B(new_n9384_), .ZN(new_n9388_));
  OAI21_X1   g09195(.A1(new_n9386_), .A2(new_n9383_), .B(new_n9388_), .ZN(new_n9389_));
  OAI22_X1   g09196(.A1(new_n2679_), .A2(new_n4704_), .B1(new_n3811_), .B2(new_n4034_), .ZN(new_n9390_));
  OAI21_X1   g09197(.A1(new_n2255_), .A2(new_n4343_), .B(new_n9390_), .ZN(new_n9391_));
  NAND3_X1   g09198(.A1(new_n9391_), .A2(\a[28] ), .A3(\a[45] ), .ZN(new_n9392_));
  AOI22_X1   g09199(.A1(\a[29] ), .A2(\a[44] ), .B1(\a[30] ), .B2(\a[43] ), .ZN(new_n9393_));
  NOR2_X1    g09200(.A1(new_n2255_), .A2(new_n4343_), .ZN(new_n9394_));
  NOR2_X1    g09201(.A1(new_n9390_), .A2(new_n9394_), .ZN(new_n9395_));
  INV_X1     g09202(.I(new_n9395_), .ZN(new_n9396_));
  OAI21_X1   g09203(.A1(new_n9393_), .A2(new_n9396_), .B(new_n9392_), .ZN(new_n9397_));
  XNOR2_X1   g09204(.A1(new_n9397_), .A2(new_n9389_), .ZN(new_n9398_));
  NOR2_X1    g09205(.A1(new_n3405_), .A2(new_n6140_), .ZN(new_n9399_));
  AOI22_X1   g09206(.A1(new_n2745_), .A2(new_n4209_), .B1(new_n3037_), .B2(new_n3928_), .ZN(new_n9400_));
  NOR2_X1    g09207(.A1(new_n9399_), .A2(new_n9400_), .ZN(new_n9401_));
  AOI21_X1   g09208(.A1(\a[35] ), .A2(\a[38] ), .B(new_n3037_), .ZN(new_n9402_));
  NOR2_X1    g09209(.A1(new_n9401_), .A2(new_n9399_), .ZN(new_n9403_));
  INV_X1     g09210(.I(new_n9403_), .ZN(new_n9404_));
  OAI22_X1   g09211(.A1(new_n9404_), .A2(new_n9402_), .B1(new_n3929_), .B2(new_n9401_), .ZN(new_n9405_));
  XOR2_X1    g09212(.A1(new_n9398_), .A2(new_n9405_), .Z(new_n9406_));
  INV_X1     g09213(.I(new_n9406_), .ZN(new_n9407_));
  NAND2_X1   g09214(.A1(new_n9267_), .A2(new_n9264_), .ZN(new_n9408_));
  OAI21_X1   g09215(.A1(new_n9268_), .A2(new_n9256_), .B(new_n9408_), .ZN(new_n9409_));
  XOR2_X1    g09216(.A1(new_n9221_), .A2(new_n9214_), .Z(new_n9410_));
  XOR2_X1    g09217(.A1(new_n9410_), .A2(new_n9263_), .Z(new_n9411_));
  XOR2_X1    g09218(.A1(new_n9409_), .A2(new_n9411_), .Z(new_n9412_));
  XOR2_X1    g09219(.A1(new_n9412_), .A2(new_n9407_), .Z(new_n9413_));
  XOR2_X1    g09220(.A1(new_n9382_), .A2(new_n9413_), .Z(new_n9414_));
  XNOR2_X1   g09221(.A1(new_n9414_), .A2(new_n9379_), .ZN(new_n9415_));
  XOR2_X1    g09222(.A1(new_n9333_), .A2(new_n9415_), .Z(new_n9416_));
  INV_X1     g09223(.I(new_n9416_), .ZN(new_n9417_));
  OAI21_X1   g09224(.A1(new_n9111_), .A2(new_n9107_), .B(new_n9149_), .ZN(new_n9418_));
  INV_X1     g09225(.I(new_n9150_), .ZN(new_n9419_));
  OAI21_X1   g09226(.A1(new_n9419_), .A2(new_n9239_), .B(new_n9418_), .ZN(new_n9420_));
  NAND2_X1   g09227(.A1(new_n9208_), .A2(new_n9237_), .ZN(new_n9421_));
  NAND2_X1   g09228(.A1(new_n9238_), .A2(new_n9205_), .ZN(new_n9422_));
  NAND2_X1   g09229(.A1(new_n9422_), .A2(new_n9421_), .ZN(new_n9423_));
  NAND2_X1   g09230(.A1(new_n9233_), .A2(new_n9235_), .ZN(new_n9424_));
  NAND2_X1   g09231(.A1(new_n9236_), .A2(new_n9230_), .ZN(new_n9425_));
  NAND2_X1   g09232(.A1(new_n9425_), .A2(new_n9424_), .ZN(new_n9426_));
  INV_X1     g09233(.I(new_n9131_), .ZN(new_n9427_));
  NOR2_X1    g09234(.A1(new_n9427_), .A2(new_n9123_), .ZN(new_n9428_));
  NOR2_X1    g09235(.A1(new_n9428_), .A2(new_n9129_), .ZN(new_n9429_));
  NAND2_X1   g09236(.A1(new_n9124_), .A2(new_n8981_), .ZN(new_n9430_));
  OAI21_X1   g09237(.A1(new_n8973_), .A2(new_n8989_), .B(new_n9430_), .ZN(new_n9431_));
  NOR2_X1    g09238(.A1(new_n2637_), .A2(new_n5377_), .ZN(new_n9432_));
  AOI22_X1   g09239(.A1(new_n2275_), .A2(new_n5239_), .B1(new_n3210_), .B2(new_n4372_), .ZN(new_n9433_));
  NOR2_X1    g09240(.A1(new_n9432_), .A2(new_n9433_), .ZN(new_n9434_));
  NAND2_X1   g09241(.A1(\a[31] ), .A2(\a[42] ), .ZN(new_n9435_));
  AOI22_X1   g09242(.A1(\a[32] ), .A2(\a[41] ), .B1(\a[33] ), .B2(\a[40] ), .ZN(new_n9436_));
  NOR2_X1    g09243(.A1(new_n9434_), .A2(new_n9432_), .ZN(new_n9437_));
  INV_X1     g09244(.I(new_n9437_), .ZN(new_n9438_));
  OAI22_X1   g09245(.A1(new_n9438_), .A2(new_n9436_), .B1(new_n9434_), .B2(new_n9435_), .ZN(new_n9439_));
  NAND2_X1   g09246(.A1(new_n8957_), .A2(new_n8964_), .ZN(new_n9440_));
  NAND2_X1   g09247(.A1(new_n9234_), .A2(new_n9036_), .ZN(new_n9441_));
  NAND2_X1   g09248(.A1(new_n9441_), .A2(new_n9440_), .ZN(new_n9442_));
  XOR2_X1    g09249(.A1(new_n9442_), .A2(new_n9439_), .Z(new_n9443_));
  XOR2_X1    g09250(.A1(new_n9443_), .A2(new_n9431_), .Z(new_n9444_));
  INV_X1     g09251(.I(new_n9444_), .ZN(new_n9445_));
  XOR2_X1    g09252(.A1(new_n9429_), .A2(new_n9445_), .Z(new_n9446_));
  XOR2_X1    g09253(.A1(new_n9426_), .A2(new_n9446_), .Z(new_n9447_));
  NAND2_X1   g09254(.A1(new_n9136_), .A2(new_n9147_), .ZN(new_n9448_));
  NAND2_X1   g09255(.A1(new_n9148_), .A2(new_n9132_), .ZN(new_n9449_));
  NAND2_X1   g09256(.A1(new_n9449_), .A2(new_n9448_), .ZN(new_n9450_));
  XOR2_X1    g09257(.A1(new_n9450_), .A2(new_n9447_), .Z(new_n9451_));
  XOR2_X1    g09258(.A1(new_n9423_), .A2(new_n9451_), .Z(new_n9452_));
  NOR2_X1    g09259(.A1(new_n9420_), .A2(new_n9452_), .ZN(new_n9453_));
  NAND2_X1   g09260(.A1(new_n9420_), .A2(new_n9452_), .ZN(new_n9454_));
  INV_X1     g09261(.I(new_n9454_), .ZN(new_n9455_));
  NOR2_X1    g09262(.A1(new_n9455_), .A2(new_n9453_), .ZN(new_n9456_));
  NAND2_X1   g09263(.A1(new_n9456_), .A2(new_n9417_), .ZN(new_n9457_));
  INV_X1     g09264(.I(new_n9457_), .ZN(new_n9458_));
  NOR2_X1    g09265(.A1(new_n9456_), .A2(new_n9417_), .ZN(new_n9459_));
  NOR2_X1    g09266(.A1(new_n9458_), .A2(new_n9459_), .ZN(new_n9460_));
  NOR2_X1    g09267(.A1(new_n9460_), .A2(new_n9303_), .ZN(new_n9461_));
  NAND2_X1   g09268(.A1(new_n9460_), .A2(new_n9303_), .ZN(new_n9462_));
  INV_X1     g09269(.I(new_n9462_), .ZN(new_n9463_));
  NOR2_X1    g09270(.A1(new_n9463_), .A2(new_n9461_), .ZN(new_n9464_));
  XOR2_X1    g09271(.A1(new_n9301_), .A2(new_n9464_), .Z(\asquared[74] ));
  AOI21_X1   g09272(.A1(new_n9300_), .A2(new_n9289_), .B(new_n9461_), .ZN(new_n9466_));
  NOR2_X1    g09273(.A1(new_n9466_), .A2(new_n9463_), .ZN(new_n9467_));
  NOR2_X1    g09274(.A1(new_n9458_), .A2(new_n9455_), .ZN(new_n9468_));
  NAND2_X1   g09275(.A1(new_n9426_), .A2(new_n9446_), .ZN(new_n9469_));
  OAI21_X1   g09276(.A1(new_n9429_), .A2(new_n9445_), .B(new_n9469_), .ZN(new_n9470_));
  XOR2_X1    g09277(.A1(new_n9395_), .A2(new_n9341_), .Z(new_n9471_));
  INV_X1     g09278(.I(new_n9471_), .ZN(new_n9472_));
  NAND2_X1   g09279(.A1(new_n9472_), .A2(new_n9351_), .ZN(new_n9473_));
  NOR2_X1    g09280(.A1(new_n9472_), .A2(new_n9351_), .ZN(new_n9474_));
  INV_X1     g09281(.I(new_n9474_), .ZN(new_n9475_));
  AND2_X2    g09282(.A1(new_n9475_), .A2(new_n9473_), .Z(new_n9476_));
  XOR2_X1    g09283(.A1(new_n9367_), .A2(new_n9375_), .Z(new_n9477_));
  XOR2_X1    g09284(.A1(new_n9477_), .A2(new_n9386_), .Z(new_n9478_));
  NAND2_X1   g09285(.A1(new_n9397_), .A2(new_n9389_), .ZN(new_n9479_));
  INV_X1     g09286(.I(new_n9398_), .ZN(new_n9480_));
  NAND2_X1   g09287(.A1(new_n9480_), .A2(new_n9405_), .ZN(new_n9481_));
  NAND2_X1   g09288(.A1(new_n9481_), .A2(new_n9479_), .ZN(new_n9482_));
  XOR2_X1    g09289(.A1(new_n9482_), .A2(new_n9478_), .Z(new_n9483_));
  XOR2_X1    g09290(.A1(new_n9483_), .A2(new_n9476_), .Z(new_n9484_));
  XOR2_X1    g09291(.A1(new_n9470_), .A2(new_n9484_), .Z(new_n9485_));
  NAND2_X1   g09292(.A1(new_n9221_), .A2(new_n9214_), .ZN(new_n9486_));
  NAND2_X1   g09293(.A1(new_n9410_), .A2(new_n9263_), .ZN(new_n9487_));
  NAND2_X1   g09294(.A1(new_n9487_), .A2(new_n9486_), .ZN(new_n9488_));
  NAND2_X1   g09295(.A1(\a[13] ), .A2(\a[61] ), .ZN(new_n9489_));
  NAND2_X1   g09296(.A1(\a[12] ), .A2(\a[62] ), .ZN(new_n9490_));
  AOI22_X1   g09297(.A1(new_n763_), .A2(new_n7590_), .B1(new_n9489_), .B2(new_n9490_), .ZN(new_n9491_));
  XOR2_X1    g09298(.A1(new_n9359_), .A2(new_n9491_), .Z(new_n9492_));
  NAND4_X1   g09299(.A1(\a[17] ), .A2(\a[29] ), .A3(\a[45] ), .A4(\a[57] ), .ZN(new_n9493_));
  NAND2_X1   g09300(.A1(new_n2254_), .A2(new_n4703_), .ZN(new_n9494_));
  NOR4_X1    g09301(.A1(new_n1023_), .A2(new_n2030_), .A3(new_n3859_), .A4(new_n6298_), .ZN(new_n9495_));
  AOI21_X1   g09302(.A1(new_n9494_), .A2(new_n9493_), .B(new_n9495_), .ZN(new_n9496_));
  NAND2_X1   g09303(.A1(\a[29] ), .A2(\a[45] ), .ZN(new_n9497_));
  AOI22_X1   g09304(.A1(\a[17] ), .A2(\a[57] ), .B1(\a[30] ), .B2(\a[44] ), .ZN(new_n9498_));
  OR2_X2     g09305(.A1(new_n9496_), .A2(new_n9495_), .Z(new_n9499_));
  OAI22_X1   g09306(.A1(new_n9499_), .A2(new_n9498_), .B1(new_n9496_), .B2(new_n9497_), .ZN(new_n9500_));
  XOR2_X1    g09307(.A1(new_n9500_), .A2(new_n9492_), .Z(new_n9501_));
  XOR2_X1    g09308(.A1(new_n9488_), .A2(new_n9501_), .Z(new_n9502_));
  AOI22_X1   g09309(.A1(\a[31] ), .A2(\a[43] ), .B1(\a[32] ), .B2(\a[42] ), .ZN(new_n9503_));
  INV_X1     g09310(.I(new_n9503_), .ZN(new_n9504_));
  NOR2_X1    g09311(.A1(new_n3833_), .A2(new_n4181_), .ZN(new_n9505_));
  NOR2_X1    g09312(.A1(new_n513_), .A2(new_n7643_), .ZN(new_n9506_));
  AOI21_X1   g09313(.A1(new_n9504_), .A2(new_n9506_), .B(new_n9505_), .ZN(new_n9507_));
  INV_X1     g09314(.I(new_n9507_), .ZN(new_n9508_));
  OAI21_X1   g09315(.A1(new_n9505_), .A2(new_n9503_), .B(new_n9506_), .ZN(new_n9509_));
  OAI21_X1   g09316(.A1(new_n9508_), .A2(new_n9503_), .B(new_n9509_), .ZN(new_n9510_));
  AOI22_X1   g09317(.A1(\a[18] ), .A2(\a[56] ), .B1(\a[25] ), .B2(\a[49] ), .ZN(new_n9511_));
  NOR3_X1    g09318(.A1(new_n8306_), .A2(new_n1441_), .A3(new_n5856_), .ZN(new_n9512_));
  NOR3_X1    g09319(.A1(new_n9511_), .A2(new_n2274_), .A3(new_n3327_), .ZN(new_n9513_));
  NOR2_X1    g09320(.A1(new_n9512_), .A2(new_n9513_), .ZN(new_n9514_));
  INV_X1     g09321(.I(new_n9514_), .ZN(new_n9515_));
  OAI21_X1   g09322(.A1(new_n9512_), .A2(new_n9511_), .B(new_n4370_), .ZN(new_n9516_));
  OAI21_X1   g09323(.A1(new_n9515_), .A2(new_n9511_), .B(new_n9516_), .ZN(new_n9517_));
  XNOR2_X1   g09324(.A1(new_n9510_), .A2(new_n9517_), .ZN(new_n9518_));
  NAND2_X1   g09325(.A1(new_n1971_), .A2(new_n4976_), .ZN(new_n9519_));
  NAND2_X1   g09326(.A1(new_n2412_), .A2(new_n6743_), .ZN(new_n9520_));
  AOI22_X1   g09327(.A1(new_n9519_), .A2(new_n9520_), .B1(new_n2103_), .B2(new_n4720_), .ZN(new_n9521_));
  NAND2_X1   g09328(.A1(\a[26] ), .A2(\a[48] ), .ZN(new_n9522_));
  AOI22_X1   g09329(.A1(\a[27] ), .A2(\a[47] ), .B1(\a[28] ), .B2(\a[46] ), .ZN(new_n9523_));
  NAND2_X1   g09330(.A1(new_n2103_), .A2(new_n4720_), .ZN(new_n9524_));
  NAND3_X1   g09331(.A1(new_n9524_), .A2(new_n9519_), .A3(new_n9520_), .ZN(new_n9525_));
  OAI22_X1   g09332(.A1(new_n9521_), .A2(new_n9522_), .B1(new_n9525_), .B2(new_n9523_), .ZN(new_n9526_));
  XOR2_X1    g09333(.A1(new_n9518_), .A2(new_n9526_), .Z(new_n9527_));
  NOR2_X1    g09334(.A1(new_n1379_), .A2(new_n6125_), .ZN(new_n9528_));
  NOR2_X1    g09335(.A1(new_n1456_), .A2(new_n6563_), .ZN(new_n9529_));
  NOR3_X1    g09336(.A1(new_n3394_), .A2(new_n5175_), .A3(new_n5680_), .ZN(new_n9530_));
  NOR2_X1    g09337(.A1(new_n9530_), .A2(new_n9529_), .ZN(new_n9531_));
  NOR2_X1    g09338(.A1(new_n9531_), .A2(new_n9528_), .ZN(new_n9532_));
  NAND2_X1   g09339(.A1(\a[22] ), .A2(\a[52] ), .ZN(new_n9533_));
  AOI22_X1   g09340(.A1(\a[19] ), .A2(\a[55] ), .B1(\a[21] ), .B2(\a[53] ), .ZN(new_n9534_));
  NOR2_X1    g09341(.A1(new_n9532_), .A2(new_n9528_), .ZN(new_n9535_));
  INV_X1     g09342(.I(new_n9535_), .ZN(new_n9536_));
  OAI22_X1   g09343(.A1(new_n9536_), .A2(new_n9534_), .B1(new_n9532_), .B2(new_n9533_), .ZN(new_n9537_));
  AOI22_X1   g09344(.A1(\a[34] ), .A2(\a[40] ), .B1(\a[35] ), .B2(\a[39] ), .ZN(new_n9538_));
  NOR2_X1    g09345(.A1(new_n2746_), .A2(new_n3551_), .ZN(new_n9539_));
  OAI21_X1   g09346(.A1(new_n9539_), .A2(new_n9538_), .B(new_n8628_), .ZN(new_n9540_));
  INV_X1     g09347(.I(new_n9538_), .ZN(new_n9541_));
  AOI21_X1   g09348(.A1(new_n8628_), .A2(new_n9541_), .B(new_n9539_), .ZN(new_n9542_));
  INV_X1     g09349(.I(new_n9542_), .ZN(new_n9543_));
  OAI21_X1   g09350(.A1(new_n9543_), .A2(new_n9538_), .B(new_n9540_), .ZN(new_n9544_));
  XNOR2_X1   g09351(.A1(new_n9537_), .A2(new_n9544_), .ZN(new_n9545_));
  AOI22_X1   g09352(.A1(\a[23] ), .A2(\a[51] ), .B1(\a[24] ), .B2(\a[50] ), .ZN(new_n9546_));
  NOR2_X1    g09353(.A1(new_n1529_), .A2(new_n5440_), .ZN(new_n9547_));
  NOR3_X1    g09354(.A1(new_n9547_), .A2(new_n2916_), .A3(new_n9546_), .ZN(new_n9548_));
  NOR2_X1    g09355(.A1(new_n9548_), .A2(new_n9547_), .ZN(new_n9549_));
  INV_X1     g09356(.I(new_n9549_), .ZN(new_n9550_));
  OAI22_X1   g09357(.A1(new_n9550_), .A2(new_n9546_), .B1(new_n2916_), .B2(new_n9548_), .ZN(new_n9551_));
  XOR2_X1    g09358(.A1(new_n9545_), .A2(new_n9551_), .Z(new_n9552_));
  XNOR2_X1   g09359(.A1(new_n9552_), .A2(new_n9527_), .ZN(new_n9553_));
  XOR2_X1    g09360(.A1(new_n9553_), .A2(new_n9502_), .Z(new_n9554_));
  XOR2_X1    g09361(.A1(new_n9485_), .A2(new_n9554_), .Z(new_n9555_));
  NAND2_X1   g09362(.A1(new_n9450_), .A2(new_n9447_), .ZN(new_n9556_));
  NAND2_X1   g09363(.A1(new_n9423_), .A2(new_n9451_), .ZN(new_n9557_));
  NAND2_X1   g09364(.A1(new_n9557_), .A2(new_n9556_), .ZN(new_n9558_));
  NAND2_X1   g09365(.A1(new_n9442_), .A2(new_n9439_), .ZN(new_n9559_));
  NAND2_X1   g09366(.A1(new_n9443_), .A2(new_n9431_), .ZN(new_n9560_));
  NAND2_X1   g09367(.A1(new_n9560_), .A2(new_n9559_), .ZN(new_n9561_));
  NAND2_X1   g09368(.A1(new_n9369_), .A2(new_n9360_), .ZN(new_n9562_));
  INV_X1     g09369(.I(new_n9376_), .ZN(new_n9563_));
  OAI21_X1   g09370(.A1(new_n9370_), .A2(new_n9563_), .B(new_n9562_), .ZN(new_n9564_));
  XOR2_X1    g09371(.A1(new_n9403_), .A2(new_n9437_), .Z(new_n9565_));
  NAND2_X1   g09372(.A1(new_n7205_), .A2(new_n1288_), .ZN(new_n9566_));
  OAI22_X1   g09373(.A1(new_n2028_), .A2(new_n7801_), .B1(new_n1173_), .B2(new_n7452_), .ZN(new_n9567_));
  NAND2_X1   g09374(.A1(new_n9567_), .A2(new_n9566_), .ZN(new_n9568_));
  NAND3_X1   g09375(.A1(new_n9568_), .A2(\a[14] ), .A3(\a[60] ), .ZN(new_n9569_));
  AOI22_X1   g09376(.A1(\a[15] ), .A2(\a[59] ), .B1(\a[16] ), .B2(\a[58] ), .ZN(new_n9570_));
  NAND2_X1   g09377(.A1(new_n9568_), .A2(new_n9566_), .ZN(new_n9571_));
  OAI21_X1   g09378(.A1(new_n9570_), .A2(new_n9571_), .B(new_n9569_), .ZN(new_n9572_));
  XNOR2_X1   g09379(.A1(new_n9565_), .A2(new_n9572_), .ZN(new_n9573_));
  INV_X1     g09380(.I(new_n9573_), .ZN(new_n9574_));
  NOR2_X1    g09381(.A1(new_n9574_), .A2(new_n9564_), .ZN(new_n9575_));
  NAND2_X1   g09382(.A1(new_n9574_), .A2(new_n9564_), .ZN(new_n9576_));
  INV_X1     g09383(.I(new_n9576_), .ZN(new_n9577_));
  NOR2_X1    g09384(.A1(new_n9577_), .A2(new_n9575_), .ZN(new_n9578_));
  NAND2_X1   g09385(.A1(new_n9561_), .A2(new_n9578_), .ZN(new_n9579_));
  INV_X1     g09386(.I(new_n9579_), .ZN(new_n9580_));
  NOR2_X1    g09387(.A1(new_n9561_), .A2(new_n9578_), .ZN(new_n9581_));
  NOR2_X1    g09388(.A1(new_n9580_), .A2(new_n9581_), .ZN(new_n9582_));
  NAND2_X1   g09389(.A1(new_n9336_), .A2(new_n9378_), .ZN(new_n9583_));
  OAI21_X1   g09390(.A1(new_n9354_), .A2(new_n9377_), .B(new_n9583_), .ZN(new_n9584_));
  NAND2_X1   g09391(.A1(new_n9409_), .A2(new_n9411_), .ZN(new_n9585_));
  NAND2_X1   g09392(.A1(new_n9412_), .A2(new_n9407_), .ZN(new_n9586_));
  NAND2_X1   g09393(.A1(new_n9586_), .A2(new_n9585_), .ZN(new_n9587_));
  XOR2_X1    g09394(.A1(new_n9587_), .A2(new_n9584_), .Z(new_n9588_));
  XOR2_X1    g09395(.A1(new_n9588_), .A2(new_n9582_), .Z(new_n9589_));
  XNOR2_X1   g09396(.A1(new_n9558_), .A2(new_n9589_), .ZN(new_n9590_));
  XNOR2_X1   g09397(.A1(new_n9590_), .A2(new_n9555_), .ZN(new_n9591_));
  INV_X1     g09398(.I(new_n9591_), .ZN(new_n9592_));
  NAND2_X1   g09399(.A1(new_n9305_), .A2(new_n9332_), .ZN(new_n9593_));
  INV_X1     g09400(.I(new_n9333_), .ZN(new_n9594_));
  OAI21_X1   g09401(.A1(new_n9594_), .A2(new_n9415_), .B(new_n9593_), .ZN(new_n9595_));
  NAND2_X1   g09402(.A1(new_n9382_), .A2(new_n9413_), .ZN(new_n9596_));
  NAND2_X1   g09403(.A1(new_n9414_), .A2(new_n9379_), .ZN(new_n9597_));
  NAND2_X1   g09404(.A1(new_n9597_), .A2(new_n9596_), .ZN(new_n9598_));
  NAND2_X1   g09405(.A1(new_n9331_), .A2(new_n9316_), .ZN(new_n9599_));
  NAND2_X1   g09406(.A1(new_n9599_), .A2(new_n9330_), .ZN(new_n9600_));
  NAND2_X1   g09407(.A1(new_n9344_), .A2(new_n9158_), .ZN(new_n9601_));
  NAND2_X1   g09408(.A1(new_n9345_), .A2(new_n9353_), .ZN(new_n9602_));
  NAND2_X1   g09409(.A1(new_n9602_), .A2(new_n9601_), .ZN(new_n9603_));
  NAND2_X1   g09410(.A1(new_n9309_), .A2(new_n9174_), .ZN(new_n9604_));
  OAI21_X1   g09411(.A1(new_n9182_), .A2(new_n9190_), .B(new_n9604_), .ZN(new_n9605_));
  NAND2_X1   g09412(.A1(new_n9311_), .A2(new_n9312_), .ZN(new_n9606_));
  NAND2_X1   g09413(.A1(new_n9313_), .A2(new_n9228_), .ZN(new_n9607_));
  NAND2_X1   g09414(.A1(new_n9607_), .A2(new_n9606_), .ZN(new_n9608_));
  XOR2_X1    g09415(.A1(new_n9605_), .A2(new_n9608_), .Z(new_n9609_));
  NAND2_X1   g09416(.A1(new_n9609_), .A2(new_n9603_), .ZN(new_n9610_));
  OR2_X2     g09417(.A1(new_n9609_), .A2(new_n9603_), .Z(new_n9611_));
  AND2_X2    g09418(.A1(new_n9611_), .A2(new_n9610_), .Z(new_n9612_));
  NAND2_X1   g09419(.A1(new_n9310_), .A2(new_n9314_), .ZN(new_n9613_));
  NAND2_X1   g09420(.A1(new_n9315_), .A2(new_n9308_), .ZN(new_n9614_));
  NAND2_X1   g09421(.A1(new_n9614_), .A2(new_n9613_), .ZN(new_n9615_));
  NAND2_X1   g09422(.A1(new_n9322_), .A2(new_n9325_), .ZN(new_n9616_));
  NAND2_X1   g09423(.A1(new_n9326_), .A2(new_n9321_), .ZN(new_n9617_));
  NAND2_X1   g09424(.A1(new_n9617_), .A2(new_n9616_), .ZN(new_n9618_));
  XOR2_X1    g09425(.A1(new_n9618_), .A2(new_n9615_), .Z(new_n9619_));
  XOR2_X1    g09426(.A1(new_n9619_), .A2(new_n9612_), .Z(new_n9620_));
  XOR2_X1    g09427(.A1(new_n9600_), .A2(new_n9620_), .Z(new_n9621_));
  XOR2_X1    g09428(.A1(new_n9621_), .A2(new_n9598_), .Z(new_n9622_));
  NOR2_X1    g09429(.A1(new_n9595_), .A2(new_n9622_), .ZN(new_n9623_));
  NAND2_X1   g09430(.A1(new_n9595_), .A2(new_n9622_), .ZN(new_n9624_));
  INV_X1     g09431(.I(new_n9624_), .ZN(new_n9625_));
  NOR2_X1    g09432(.A1(new_n9625_), .A2(new_n9623_), .ZN(new_n9626_));
  NOR2_X1    g09433(.A1(new_n9626_), .A2(new_n9592_), .ZN(new_n9627_));
  NAND2_X1   g09434(.A1(new_n9626_), .A2(new_n9592_), .ZN(new_n9628_));
  INV_X1     g09435(.I(new_n9628_), .ZN(new_n9629_));
  NOR2_X1    g09436(.A1(new_n9629_), .A2(new_n9627_), .ZN(new_n9630_));
  INV_X1     g09437(.I(new_n9630_), .ZN(new_n9631_));
  NOR2_X1    g09438(.A1(new_n9468_), .A2(new_n9631_), .ZN(new_n9632_));
  INV_X1     g09439(.I(new_n9632_), .ZN(new_n9633_));
  NAND2_X1   g09440(.A1(new_n9468_), .A2(new_n9631_), .ZN(new_n9634_));
  NAND2_X1   g09441(.A1(new_n9633_), .A2(new_n9634_), .ZN(new_n9635_));
  XOR2_X1    g09442(.A1(new_n9467_), .A2(new_n9635_), .Z(\asquared[75] ));
  OAI21_X1   g09443(.A1(new_n9466_), .A2(new_n9463_), .B(new_n9634_), .ZN(new_n9637_));
  NAND2_X1   g09444(.A1(new_n9637_), .A2(new_n9633_), .ZN(new_n9638_));
  NOR2_X1    g09445(.A1(new_n9629_), .A2(new_n9625_), .ZN(new_n9639_));
  INV_X1     g09446(.I(new_n9639_), .ZN(new_n9640_));
  NAND2_X1   g09447(.A1(new_n9618_), .A2(new_n9615_), .ZN(new_n9641_));
  NAND2_X1   g09448(.A1(new_n9619_), .A2(new_n9612_), .ZN(new_n9642_));
  NAND2_X1   g09449(.A1(new_n9642_), .A2(new_n9641_), .ZN(new_n9643_));
  XOR2_X1    g09450(.A1(new_n9499_), .A2(new_n9525_), .Z(new_n9644_));
  XOR2_X1    g09451(.A1(new_n9644_), .A2(new_n9571_), .Z(new_n9645_));
  NAND2_X1   g09452(.A1(new_n9537_), .A2(new_n9544_), .ZN(new_n9646_));
  INV_X1     g09453(.I(new_n9551_), .ZN(new_n9647_));
  OAI21_X1   g09454(.A1(new_n9545_), .A2(new_n9647_), .B(new_n9646_), .ZN(new_n9648_));
  NAND2_X1   g09455(.A1(new_n9510_), .A2(new_n9517_), .ZN(new_n9649_));
  INV_X1     g09456(.I(new_n9518_), .ZN(new_n9650_));
  NAND2_X1   g09457(.A1(new_n9650_), .A2(new_n9526_), .ZN(new_n9651_));
  NAND2_X1   g09458(.A1(new_n9651_), .A2(new_n9649_), .ZN(new_n9652_));
  XOR2_X1    g09459(.A1(new_n9648_), .A2(new_n9652_), .Z(new_n9653_));
  XOR2_X1    g09460(.A1(new_n9653_), .A2(new_n9645_), .Z(new_n9654_));
  XOR2_X1    g09461(.A1(new_n9643_), .A2(new_n9654_), .Z(new_n9655_));
  NOR2_X1    g09462(.A1(new_n4702_), .A2(new_n6298_), .ZN(new_n9656_));
  INV_X1     g09463(.I(new_n9656_), .ZN(new_n9657_));
  NOR2_X1    g09464(.A1(new_n9657_), .A2(new_n3787_), .ZN(new_n9658_));
  NOR2_X1    g09465(.A1(new_n1566_), .A2(new_n6316_), .ZN(new_n9659_));
  AOI22_X1   g09466(.A1(new_n1027_), .A2(new_n6803_), .B1(new_n6340_), .B2(new_n9659_), .ZN(new_n9660_));
  NOR2_X1    g09467(.A1(new_n9660_), .A2(new_n9658_), .ZN(new_n9661_));
  OAI21_X1   g09468(.A1(new_n3787_), .A2(new_n9657_), .B(new_n9660_), .ZN(new_n9662_));
  AOI22_X1   g09469(.A1(\a[18] ), .A2(\a[57] ), .B1(\a[26] ), .B2(\a[49] ), .ZN(new_n9663_));
  OAI22_X1   g09470(.A1(new_n9662_), .A2(new_n9663_), .B1(new_n9661_), .B2(new_n7541_), .ZN(new_n9664_));
  NAND2_X1   g09471(.A1(new_n7451_), .A2(new_n1288_), .ZN(new_n9665_));
  OAI22_X1   g09472(.A1(new_n2028_), .A2(new_n6899_), .B1(new_n1173_), .B2(new_n7454_), .ZN(new_n9666_));
  NAND2_X1   g09473(.A1(new_n9666_), .A2(new_n9665_), .ZN(new_n9667_));
  NAND3_X1   g09474(.A1(new_n9667_), .A2(\a[14] ), .A3(\a[61] ), .ZN(new_n9668_));
  AOI22_X1   g09475(.A1(\a[15] ), .A2(\a[60] ), .B1(\a[16] ), .B2(\a[59] ), .ZN(new_n9669_));
  NAND2_X1   g09476(.A1(new_n9667_), .A2(new_n9665_), .ZN(new_n9670_));
  OAI21_X1   g09477(.A1(new_n9669_), .A2(new_n9670_), .B(new_n9668_), .ZN(new_n9671_));
  XNOR2_X1   g09478(.A1(new_n9671_), .A2(new_n9664_), .ZN(new_n9672_));
  INV_X1     g09479(.I(new_n6743_), .ZN(new_n9673_));
  OAI22_X1   g09480(.A1(new_n1816_), .A2(new_n9673_), .B1(new_n2189_), .B2(new_n4977_), .ZN(new_n9674_));
  OAI21_X1   g09481(.A1(new_n2679_), .A2(new_n4721_), .B(new_n9674_), .ZN(new_n9675_));
  NAND3_X1   g09482(.A1(new_n9675_), .A2(\a[27] ), .A3(\a[48] ), .ZN(new_n9676_));
  AOI22_X1   g09483(.A1(\a[28] ), .A2(\a[47] ), .B1(\a[29] ), .B2(\a[46] ), .ZN(new_n9677_));
  NOR2_X1    g09484(.A1(new_n2679_), .A2(new_n4721_), .ZN(new_n9678_));
  NOR2_X1    g09485(.A1(new_n9674_), .A2(new_n9678_), .ZN(new_n9679_));
  INV_X1     g09486(.I(new_n9679_), .ZN(new_n9680_));
  OAI21_X1   g09487(.A1(new_n9677_), .A2(new_n9680_), .B(new_n9676_), .ZN(new_n9681_));
  XOR2_X1    g09488(.A1(new_n9672_), .A2(new_n9681_), .Z(new_n9682_));
  INV_X1     g09489(.I(new_n9682_), .ZN(new_n9683_));
  NAND2_X1   g09490(.A1(new_n9605_), .A2(new_n9608_), .ZN(new_n9684_));
  NAND2_X1   g09491(.A1(new_n9610_), .A2(new_n9684_), .ZN(new_n9685_));
  AOI22_X1   g09492(.A1(\a[12] ), .A2(\a[63] ), .B1(\a[19] ), .B2(\a[56] ), .ZN(new_n9686_));
  INV_X1     g09493(.I(new_n9686_), .ZN(new_n9687_));
  NOR2_X1    g09494(.A1(new_n979_), .A2(new_n7643_), .ZN(new_n9688_));
  INV_X1     g09495(.I(new_n9688_), .ZN(new_n9689_));
  NOR2_X1    g09496(.A1(new_n8409_), .A2(new_n9689_), .ZN(new_n9690_));
  NOR2_X1    g09497(.A1(new_n2030_), .A2(new_n4030_), .ZN(new_n9691_));
  AOI21_X1   g09498(.A1(new_n9687_), .A2(new_n9691_), .B(new_n9690_), .ZN(new_n9692_));
  INV_X1     g09499(.I(new_n9692_), .ZN(new_n9693_));
  OAI21_X1   g09500(.A1(new_n9690_), .A2(new_n9686_), .B(new_n9691_), .ZN(new_n9694_));
  OAI21_X1   g09501(.A1(new_n9693_), .A2(new_n9686_), .B(new_n9694_), .ZN(new_n9695_));
  NOR2_X1    g09502(.A1(new_n1299_), .A2(new_n5175_), .ZN(new_n9696_));
  INV_X1     g09503(.I(new_n6916_), .ZN(new_n9697_));
  OAI21_X1   g09504(.A1(new_n2524_), .A2(new_n3221_), .B(new_n9697_), .ZN(new_n9698_));
  NAND2_X1   g09505(.A1(new_n3232_), .A2(new_n3550_), .ZN(new_n9699_));
  NAND3_X1   g09506(.A1(new_n9698_), .A2(new_n9696_), .A3(new_n9699_), .ZN(new_n9700_));
  NAND2_X1   g09507(.A1(new_n9700_), .A2(new_n9696_), .ZN(new_n9701_));
  NAND3_X1   g09508(.A1(new_n9700_), .A2(new_n9698_), .A3(new_n9699_), .ZN(new_n9702_));
  NAND2_X1   g09509(.A1(new_n9702_), .A2(new_n9701_), .ZN(new_n9703_));
  XNOR2_X1   g09510(.A1(new_n9703_), .A2(new_n9695_), .ZN(new_n9704_));
  NAND2_X1   g09511(.A1(\a[38] ), .A2(\a[62] ), .ZN(new_n9705_));
  NOR2_X1    g09512(.A1(new_n9705_), .A2(new_n597_), .ZN(new_n9706_));
  NOR2_X1    g09513(.A1(new_n6140_), .A2(new_n9706_), .ZN(new_n9707_));
  AOI21_X1   g09514(.A1(\a[13] ), .A2(\a[62] ), .B(\a[38] ), .ZN(new_n9708_));
  NOR2_X1    g09515(.A1(new_n9706_), .A2(new_n3803_), .ZN(new_n9709_));
  INV_X1     g09516(.I(new_n9709_), .ZN(new_n9710_));
  OAI22_X1   g09517(.A1(new_n9710_), .A2(new_n9708_), .B1(new_n9707_), .B2(new_n6140_), .ZN(new_n9711_));
  XOR2_X1    g09518(.A1(new_n9704_), .A2(new_n9711_), .Z(new_n9712_));
  INV_X1     g09519(.I(new_n9712_), .ZN(new_n9713_));
  XOR2_X1    g09520(.A1(new_n9685_), .A2(new_n9713_), .Z(new_n9714_));
  XOR2_X1    g09521(.A1(new_n9714_), .A2(new_n9683_), .Z(new_n9715_));
  XNOR2_X1   g09522(.A1(new_n9655_), .A2(new_n9715_), .ZN(new_n9716_));
  NAND2_X1   g09523(.A1(new_n9600_), .A2(new_n9620_), .ZN(new_n9717_));
  NAND2_X1   g09524(.A1(new_n9621_), .A2(new_n9598_), .ZN(new_n9718_));
  NAND2_X1   g09525(.A1(new_n9718_), .A2(new_n9717_), .ZN(new_n9719_));
  NAND2_X1   g09526(.A1(new_n9500_), .A2(new_n9492_), .ZN(new_n9720_));
  NAND2_X1   g09527(.A1(new_n9488_), .A2(new_n9501_), .ZN(new_n9721_));
  NAND2_X1   g09528(.A1(new_n9721_), .A2(new_n9720_), .ZN(new_n9722_));
  XOR2_X1    g09529(.A1(new_n9549_), .A2(new_n9542_), .Z(new_n9723_));
  XOR2_X1    g09530(.A1(new_n9723_), .A2(new_n9536_), .Z(new_n9724_));
  INV_X1     g09531(.I(new_n9724_), .ZN(new_n9725_));
  NAND2_X1   g09532(.A1(new_n9359_), .A2(new_n9491_), .ZN(new_n9726_));
  OAI21_X1   g09533(.A1(new_n1265_), .A2(new_n7591_), .B(new_n9726_), .ZN(new_n9727_));
  XOR2_X1    g09534(.A1(new_n9507_), .A2(new_n9514_), .Z(new_n9728_));
  XOR2_X1    g09535(.A1(new_n9728_), .A2(new_n9727_), .Z(new_n9729_));
  INV_X1     g09536(.I(new_n9729_), .ZN(new_n9730_));
  NOR2_X1    g09537(.A1(new_n9725_), .A2(new_n9730_), .ZN(new_n9731_));
  NOR2_X1    g09538(.A1(new_n9724_), .A2(new_n9729_), .ZN(new_n9732_));
  NOR2_X1    g09539(.A1(new_n9731_), .A2(new_n9732_), .ZN(new_n9733_));
  NOR2_X1    g09540(.A1(new_n9733_), .A2(new_n9722_), .ZN(new_n9734_));
  NAND2_X1   g09541(.A1(new_n9733_), .A2(new_n9722_), .ZN(new_n9735_));
  INV_X1     g09542(.I(new_n9735_), .ZN(new_n9736_));
  NOR2_X1    g09543(.A1(new_n9736_), .A2(new_n9734_), .ZN(new_n9737_));
  NOR2_X1    g09544(.A1(new_n9395_), .A2(new_n9341_), .ZN(new_n9738_));
  NOR2_X1    g09545(.A1(new_n9474_), .A2(new_n9738_), .ZN(new_n9739_));
  NAND2_X1   g09546(.A1(new_n9367_), .A2(new_n9375_), .ZN(new_n9740_));
  NAND2_X1   g09547(.A1(new_n9477_), .A2(new_n9386_), .ZN(new_n9741_));
  NAND2_X1   g09548(.A1(new_n9741_), .A2(new_n9740_), .ZN(new_n9742_));
  NAND2_X1   g09549(.A1(new_n9565_), .A2(new_n9572_), .ZN(new_n9743_));
  OAI21_X1   g09550(.A1(new_n9403_), .A2(new_n9437_), .B(new_n9743_), .ZN(new_n9744_));
  XOR2_X1    g09551(.A1(new_n9744_), .A2(new_n9742_), .Z(new_n9745_));
  XNOR2_X1   g09552(.A1(new_n9745_), .A2(new_n9739_), .ZN(new_n9746_));
  INV_X1     g09553(.I(new_n9746_), .ZN(new_n9747_));
  INV_X1     g09554(.I(new_n9553_), .ZN(new_n9748_));
  NOR2_X1    g09555(.A1(new_n9552_), .A2(new_n9527_), .ZN(new_n9749_));
  AOI21_X1   g09556(.A1(new_n9748_), .A2(new_n9502_), .B(new_n9749_), .ZN(new_n9750_));
  XOR2_X1    g09557(.A1(new_n9750_), .A2(new_n9747_), .Z(new_n9751_));
  NOR2_X1    g09558(.A1(new_n9751_), .A2(new_n9737_), .ZN(new_n9752_));
  NAND2_X1   g09559(.A1(new_n9751_), .A2(new_n9737_), .ZN(new_n9753_));
  INV_X1     g09560(.I(new_n9753_), .ZN(new_n9754_));
  NOR2_X1    g09561(.A1(new_n9754_), .A2(new_n9752_), .ZN(new_n9755_));
  XOR2_X1    g09562(.A1(new_n9719_), .A2(new_n9755_), .Z(new_n9756_));
  INV_X1     g09563(.I(new_n9756_), .ZN(new_n9757_));
  OR2_X2     g09564(.A1(new_n9757_), .A2(new_n9716_), .Z(new_n9758_));
  NAND2_X1   g09565(.A1(new_n9757_), .A2(new_n9716_), .ZN(new_n9759_));
  NAND2_X1   g09566(.A1(new_n9758_), .A2(new_n9759_), .ZN(new_n9760_));
  NAND2_X1   g09567(.A1(new_n9470_), .A2(new_n9484_), .ZN(new_n9761_));
  INV_X1     g09568(.I(new_n9485_), .ZN(new_n9762_));
  OAI21_X1   g09569(.A1(new_n9762_), .A2(new_n9554_), .B(new_n9761_), .ZN(new_n9763_));
  NAND2_X1   g09570(.A1(new_n9482_), .A2(new_n9478_), .ZN(new_n9764_));
  NAND2_X1   g09571(.A1(new_n9483_), .A2(new_n9476_), .ZN(new_n9765_));
  NAND2_X1   g09572(.A1(new_n9765_), .A2(new_n9764_), .ZN(new_n9766_));
  NOR2_X1    g09573(.A1(new_n2637_), .A2(new_n4181_), .ZN(new_n9767_));
  NOR2_X1    g09574(.A1(new_n2276_), .A2(new_n3861_), .ZN(new_n9768_));
  NOR2_X1    g09575(.A1(new_n3833_), .A2(new_n4343_), .ZN(new_n9769_));
  NOR2_X1    g09576(.A1(new_n9768_), .A2(new_n9769_), .ZN(new_n9770_));
  NOR2_X1    g09577(.A1(new_n9770_), .A2(new_n9767_), .ZN(new_n9771_));
  NAND2_X1   g09578(.A1(\a[31] ), .A2(\a[44] ), .ZN(new_n9772_));
  AOI22_X1   g09579(.A1(\a[32] ), .A2(\a[43] ), .B1(\a[33] ), .B2(\a[42] ), .ZN(new_n9773_));
  NOR2_X1    g09580(.A1(new_n9771_), .A2(new_n9767_), .ZN(new_n9774_));
  INV_X1     g09581(.I(new_n9774_), .ZN(new_n9775_));
  OAI22_X1   g09582(.A1(new_n9775_), .A2(new_n9773_), .B1(new_n9771_), .B2(new_n9772_), .ZN(new_n9776_));
  AOI22_X1   g09583(.A1(\a[20] ), .A2(\a[55] ), .B1(\a[25] ), .B2(\a[50] ), .ZN(new_n9777_));
  NOR4_X1    g09584(.A1(new_n1043_), .A2(new_n1441_), .A3(new_n4901_), .A4(new_n5680_), .ZN(new_n9778_));
  NOR3_X1    g09585(.A1(new_n9777_), .A2(new_n2442_), .A3(new_n3327_), .ZN(new_n9779_));
  NOR2_X1    g09586(.A1(new_n9779_), .A2(new_n9778_), .ZN(new_n9780_));
  INV_X1     g09587(.I(new_n9780_), .ZN(new_n9781_));
  NOR2_X1    g09588(.A1(new_n2442_), .A2(new_n3327_), .ZN(new_n9782_));
  OAI21_X1   g09589(.A1(new_n9778_), .A2(new_n9777_), .B(new_n9782_), .ZN(new_n9783_));
  OAI21_X1   g09590(.A1(new_n9781_), .A2(new_n9777_), .B(new_n9783_), .ZN(new_n9784_));
  XNOR2_X1   g09591(.A1(new_n9776_), .A2(new_n9784_), .ZN(new_n9785_));
  NOR2_X1    g09592(.A1(new_n1880_), .A2(new_n5683_), .ZN(new_n9786_));
  NAND4_X1   g09593(.A1(\a[21] ), .A2(\a[24] ), .A3(\a[51] ), .A4(\a[54] ), .ZN(new_n9787_));
  NAND2_X1   g09594(.A1(new_n1452_), .A2(new_n6126_), .ZN(new_n9788_));
  AOI21_X1   g09595(.A1(new_n9787_), .A2(new_n9788_), .B(new_n9786_), .ZN(new_n9789_));
  NAND2_X1   g09596(.A1(\a[21] ), .A2(\a[54] ), .ZN(new_n9790_));
  AOI22_X1   g09597(.A1(\a[22] ), .A2(\a[53] ), .B1(\a[24] ), .B2(\a[51] ), .ZN(new_n9791_));
  NOR2_X1    g09598(.A1(new_n9789_), .A2(new_n9786_), .ZN(new_n9792_));
  INV_X1     g09599(.I(new_n9792_), .ZN(new_n9793_));
  OAI22_X1   g09600(.A1(new_n9793_), .A2(new_n9791_), .B1(new_n9789_), .B2(new_n9790_), .ZN(new_n9794_));
  XOR2_X1    g09601(.A1(new_n9785_), .A2(new_n9794_), .Z(new_n9795_));
  XOR2_X1    g09602(.A1(new_n9766_), .A2(new_n9795_), .Z(new_n9796_));
  NOR2_X1    g09603(.A1(new_n9580_), .A2(new_n9577_), .ZN(new_n9797_));
  XNOR2_X1   g09604(.A1(new_n9796_), .A2(new_n9797_), .ZN(new_n9798_));
  NAND2_X1   g09605(.A1(new_n9587_), .A2(new_n9584_), .ZN(new_n9799_));
  NAND2_X1   g09606(.A1(new_n9588_), .A2(new_n9582_), .ZN(new_n9800_));
  NAND2_X1   g09607(.A1(new_n9800_), .A2(new_n9799_), .ZN(new_n9801_));
  XOR2_X1    g09608(.A1(new_n9801_), .A2(new_n9798_), .Z(new_n9802_));
  XNOR2_X1   g09609(.A1(new_n9802_), .A2(new_n9763_), .ZN(new_n9803_));
  NAND2_X1   g09610(.A1(new_n9558_), .A2(new_n9589_), .ZN(new_n9804_));
  OAI21_X1   g09611(.A1(new_n9590_), .A2(new_n9555_), .B(new_n9804_), .ZN(new_n9805_));
  XOR2_X1    g09612(.A1(new_n9805_), .A2(new_n9803_), .Z(new_n9806_));
  INV_X1     g09613(.I(new_n9806_), .ZN(new_n9807_));
  XOR2_X1    g09614(.A1(new_n9760_), .A2(new_n9807_), .Z(new_n9808_));
  NOR2_X1    g09615(.A1(new_n9640_), .A2(new_n9808_), .ZN(new_n9809_));
  NAND2_X1   g09616(.A1(new_n9640_), .A2(new_n9808_), .ZN(new_n9810_));
  INV_X1     g09617(.I(new_n9810_), .ZN(new_n9811_));
  NOR2_X1    g09618(.A1(new_n9811_), .A2(new_n9809_), .ZN(new_n9812_));
  XOR2_X1    g09619(.A1(new_n9638_), .A2(new_n9812_), .Z(\asquared[76] ));
  AOI21_X1   g09620(.A1(new_n9637_), .A2(new_n9633_), .B(new_n9809_), .ZN(new_n9814_));
  NOR2_X1    g09621(.A1(new_n9814_), .A2(new_n9811_), .ZN(new_n9815_));
  NAND2_X1   g09622(.A1(new_n9719_), .A2(new_n9755_), .ZN(new_n9816_));
  NAND2_X1   g09623(.A1(new_n9758_), .A2(new_n9816_), .ZN(new_n9817_));
  NAND2_X1   g09624(.A1(new_n9643_), .A2(new_n9654_), .ZN(new_n9818_));
  NAND2_X1   g09625(.A1(new_n9655_), .A2(new_n9715_), .ZN(new_n9819_));
  NAND2_X1   g09626(.A1(new_n9819_), .A2(new_n9818_), .ZN(new_n9820_));
  NOR2_X1    g09627(.A1(new_n9750_), .A2(new_n9747_), .ZN(new_n9821_));
  NOR2_X1    g09628(.A1(new_n9754_), .A2(new_n9821_), .ZN(new_n9822_));
  NOR2_X1    g09629(.A1(new_n9736_), .A2(new_n9731_), .ZN(new_n9823_));
  NAND2_X1   g09630(.A1(new_n9648_), .A2(new_n9652_), .ZN(new_n9824_));
  NAND2_X1   g09631(.A1(new_n9653_), .A2(new_n9645_), .ZN(new_n9825_));
  NAND2_X1   g09632(.A1(new_n9825_), .A2(new_n9824_), .ZN(new_n9826_));
  AOI22_X1   g09633(.A1(\a[19] ), .A2(\a[57] ), .B1(\a[23] ), .B2(\a[53] ), .ZN(new_n9827_));
  INV_X1     g09634(.I(new_n9827_), .ZN(new_n9828_));
  NOR4_X1    g09635(.A1(new_n979_), .A2(new_n1299_), .A3(new_n5425_), .A4(new_n6298_), .ZN(new_n9829_));
  AOI21_X1   g09636(.A1(new_n4495_), .A2(new_n9828_), .B(new_n9829_), .ZN(new_n9830_));
  INV_X1     g09637(.I(new_n9830_), .ZN(new_n9831_));
  OAI21_X1   g09638(.A1(new_n9829_), .A2(new_n9827_), .B(new_n4495_), .ZN(new_n9832_));
  OAI21_X1   g09639(.A1(new_n9831_), .A2(new_n9827_), .B(new_n9832_), .ZN(new_n9833_));
  AOI22_X1   g09640(.A1(\a[31] ), .A2(\a[45] ), .B1(\a[32] ), .B2(\a[44] ), .ZN(new_n9834_));
  INV_X1     g09641(.I(new_n9834_), .ZN(new_n9835_));
  NOR2_X1    g09642(.A1(new_n3833_), .A2(new_n4704_), .ZN(new_n9836_));
  NOR2_X1    g09643(.A1(new_n597_), .A2(new_n7643_), .ZN(new_n9837_));
  AOI21_X1   g09644(.A1(new_n9835_), .A2(new_n9837_), .B(new_n9836_), .ZN(new_n9838_));
  INV_X1     g09645(.I(new_n9838_), .ZN(new_n9839_));
  OAI21_X1   g09646(.A1(new_n9836_), .A2(new_n9834_), .B(new_n9837_), .ZN(new_n9840_));
  OAI21_X1   g09647(.A1(new_n9839_), .A2(new_n9834_), .B(new_n9840_), .ZN(new_n9841_));
  XOR2_X1    g09648(.A1(new_n9841_), .A2(new_n9833_), .Z(new_n9842_));
  NAND2_X1   g09649(.A1(new_n1552_), .A2(new_n5857_), .ZN(new_n9843_));
  NAND2_X1   g09650(.A1(new_n1381_), .A2(new_n7184_), .ZN(new_n9844_));
  AOI22_X1   g09651(.A1(new_n9843_), .A2(new_n9844_), .B1(new_n1452_), .B2(new_n6128_), .ZN(new_n9845_));
  AOI22_X1   g09652(.A1(\a[21] ), .A2(\a[55] ), .B1(\a[22] ), .B2(\a[54] ), .ZN(new_n9846_));
  NAND2_X1   g09653(.A1(new_n1452_), .A2(new_n6128_), .ZN(new_n9847_));
  NAND3_X1   g09654(.A1(new_n9847_), .A2(new_n9843_), .A3(new_n9844_), .ZN(new_n9848_));
  OAI22_X1   g09655(.A1(new_n9845_), .A2(new_n7749_), .B1(new_n9848_), .B2(new_n9846_), .ZN(new_n9849_));
  XOR2_X1    g09656(.A1(new_n9842_), .A2(new_n9849_), .Z(new_n9850_));
  XOR2_X1    g09657(.A1(new_n9826_), .A2(new_n9850_), .Z(new_n9851_));
  XOR2_X1    g09658(.A1(new_n9851_), .A2(new_n9823_), .Z(new_n9852_));
  XOR2_X1    g09659(.A1(new_n9822_), .A2(new_n9852_), .Z(new_n9853_));
  NOR2_X1    g09660(.A1(new_n9853_), .A2(new_n9820_), .ZN(new_n9854_));
  NAND2_X1   g09661(.A1(new_n9853_), .A2(new_n9820_), .ZN(new_n9855_));
  INV_X1     g09662(.I(new_n9855_), .ZN(new_n9856_));
  NOR2_X1    g09663(.A1(new_n9856_), .A2(new_n9854_), .ZN(new_n9857_));
  XOR2_X1    g09664(.A1(new_n9817_), .A2(new_n9857_), .Z(new_n9858_));
  INV_X1     g09665(.I(new_n9795_), .ZN(new_n9859_));
  NAND2_X1   g09666(.A1(new_n9766_), .A2(new_n9859_), .ZN(new_n9860_));
  OAI21_X1   g09667(.A1(new_n9796_), .A2(new_n9797_), .B(new_n9860_), .ZN(new_n9861_));
  XOR2_X1    g09668(.A1(new_n9670_), .A2(new_n9662_), .Z(new_n9862_));
  XOR2_X1    g09669(.A1(new_n9862_), .A2(new_n9775_), .Z(new_n9863_));
  NAND2_X1   g09670(.A1(new_n9671_), .A2(new_n9664_), .ZN(new_n9864_));
  INV_X1     g09671(.I(new_n9672_), .ZN(new_n9865_));
  NAND2_X1   g09672(.A1(new_n9865_), .A2(new_n9681_), .ZN(new_n9866_));
  NAND2_X1   g09673(.A1(new_n9866_), .A2(new_n9864_), .ZN(new_n9867_));
  NAND2_X1   g09674(.A1(new_n9703_), .A2(new_n9695_), .ZN(new_n9868_));
  INV_X1     g09675(.I(new_n9711_), .ZN(new_n9869_));
  OAI21_X1   g09676(.A1(new_n9704_), .A2(new_n9869_), .B(new_n9868_), .ZN(new_n9870_));
  XOR2_X1    g09677(.A1(new_n9867_), .A2(new_n9870_), .Z(new_n9871_));
  XOR2_X1    g09678(.A1(new_n9871_), .A2(new_n9863_), .Z(new_n9872_));
  XOR2_X1    g09679(.A1(new_n9861_), .A2(new_n9872_), .Z(new_n9873_));
  AOI22_X1   g09680(.A1(\a[26] ), .A2(\a[50] ), .B1(\a[27] ), .B2(\a[49] ), .ZN(new_n9874_));
  NOR2_X1    g09681(.A1(new_n884_), .A2(new_n6316_), .ZN(new_n9875_));
  INV_X1     g09682(.I(new_n9875_), .ZN(new_n9876_));
  NOR2_X1    g09683(.A1(new_n1972_), .A2(new_n5155_), .ZN(new_n9877_));
  NOR3_X1    g09684(.A1(new_n9877_), .A2(new_n9874_), .A3(new_n9876_), .ZN(new_n9878_));
  NOR2_X1    g09685(.A1(new_n9878_), .A2(new_n9877_), .ZN(new_n9879_));
  INV_X1     g09686(.I(new_n9879_), .ZN(new_n9880_));
  OAI22_X1   g09687(.A1(new_n9880_), .A2(new_n9874_), .B1(new_n9876_), .B2(new_n9878_), .ZN(new_n9881_));
  INV_X1     g09688(.I(new_n9881_), .ZN(new_n9882_));
  OAI22_X1   g09689(.A1(new_n893_), .A2(new_n7454_), .B1(new_n6899_), .B2(new_n982_), .ZN(new_n9883_));
  OAI21_X1   g09690(.A1(new_n1428_), .A2(new_n7452_), .B(new_n9883_), .ZN(new_n9884_));
  NAND3_X1   g09691(.A1(new_n9884_), .A2(\a[15] ), .A3(\a[61] ), .ZN(new_n9885_));
  AOI22_X1   g09692(.A1(\a[16] ), .A2(\a[60] ), .B1(\a[17] ), .B2(\a[59] ), .ZN(new_n9886_));
  NOR2_X1    g09693(.A1(new_n1428_), .A2(new_n7452_), .ZN(new_n9887_));
  NOR2_X1    g09694(.A1(new_n9883_), .A2(new_n9887_), .ZN(new_n9888_));
  INV_X1     g09695(.I(new_n9888_), .ZN(new_n9889_));
  OAI21_X1   g09696(.A1(new_n9886_), .A2(new_n9889_), .B(new_n9885_), .ZN(new_n9890_));
  XOR2_X1    g09697(.A1(new_n9890_), .A2(new_n9792_), .Z(new_n9891_));
  NOR2_X1    g09698(.A1(new_n9891_), .A2(new_n9882_), .ZN(new_n9892_));
  INV_X1     g09699(.I(new_n9892_), .ZN(new_n9893_));
  NAND2_X1   g09700(.A1(new_n9891_), .A2(new_n9882_), .ZN(new_n9894_));
  AND2_X2    g09701(.A1(new_n9893_), .A2(new_n9894_), .Z(new_n9895_));
  NAND2_X1   g09702(.A1(new_n9744_), .A2(new_n9742_), .ZN(new_n9896_));
  INV_X1     g09703(.I(new_n9745_), .ZN(new_n9897_));
  OAI21_X1   g09704(.A1(new_n9897_), .A2(new_n9739_), .B(new_n9896_), .ZN(new_n9898_));
  NAND2_X1   g09705(.A1(new_n2254_), .A2(new_n4720_), .ZN(new_n9899_));
  OAI22_X1   g09706(.A1(new_n2679_), .A2(new_n4977_), .B1(new_n3811_), .B2(new_n9673_), .ZN(new_n9900_));
  NAND2_X1   g09707(.A1(new_n9900_), .A2(new_n9899_), .ZN(new_n9901_));
  NAND3_X1   g09708(.A1(new_n9901_), .A2(\a[28] ), .A3(\a[48] ), .ZN(new_n9902_));
  AOI22_X1   g09709(.A1(\a[29] ), .A2(\a[47] ), .B1(\a[30] ), .B2(\a[46] ), .ZN(new_n9903_));
  NAND2_X1   g09710(.A1(new_n9901_), .A2(new_n9899_), .ZN(new_n9904_));
  OAI21_X1   g09711(.A1(new_n9903_), .A2(new_n9904_), .B(new_n9902_), .ZN(new_n9905_));
  NAND2_X1   g09712(.A1(new_n3232_), .A2(new_n4534_), .ZN(new_n9906_));
  OAI22_X1   g09713(.A1(new_n2746_), .A2(new_n4667_), .B1(new_n5564_), .B2(new_n7757_), .ZN(new_n9907_));
  NAND2_X1   g09714(.A1(new_n9907_), .A2(new_n9906_), .ZN(new_n9908_));
  NAND3_X1   g09715(.A1(new_n9908_), .A2(\a[34] ), .A3(\a[42] ), .ZN(new_n9909_));
  AOI22_X1   g09716(.A1(\a[35] ), .A2(\a[41] ), .B1(\a[36] ), .B2(\a[40] ), .ZN(new_n9910_));
  NAND2_X1   g09717(.A1(new_n9908_), .A2(new_n9906_), .ZN(new_n9911_));
  OAI21_X1   g09718(.A1(new_n9910_), .A2(new_n9911_), .B(new_n9909_), .ZN(new_n9912_));
  XOR2_X1    g09719(.A1(new_n9905_), .A2(new_n9912_), .Z(new_n9913_));
  AOI22_X1   g09720(.A1(\a[24] ), .A2(\a[52] ), .B1(\a[25] ), .B2(\a[51] ), .ZN(new_n9914_));
  OAI21_X1   g09721(.A1(new_n1779_), .A2(new_n5525_), .B(new_n4545_), .ZN(new_n9915_));
  NOR2_X1    g09722(.A1(new_n9915_), .A2(new_n9914_), .ZN(new_n9916_));
  AOI21_X1   g09723(.A1(new_n1778_), .A2(new_n5524_), .B(new_n9916_), .ZN(new_n9917_));
  INV_X1     g09724(.I(new_n9917_), .ZN(new_n9918_));
  OAI22_X1   g09725(.A1(new_n9918_), .A2(new_n9914_), .B1(new_n4739_), .B2(new_n9916_), .ZN(new_n9919_));
  XNOR2_X1   g09726(.A1(new_n9913_), .A2(new_n9919_), .ZN(new_n9920_));
  INV_X1     g09727(.I(new_n9920_), .ZN(new_n9921_));
  XOR2_X1    g09728(.A1(new_n9898_), .A2(new_n9921_), .Z(new_n9922_));
  XOR2_X1    g09729(.A1(new_n9922_), .A2(new_n9895_), .Z(new_n9923_));
  XNOR2_X1   g09730(.A1(new_n9873_), .A2(new_n9923_), .ZN(new_n9924_));
  INV_X1     g09731(.I(new_n9798_), .ZN(new_n9925_));
  NAND2_X1   g09732(.A1(new_n9925_), .A2(new_n9801_), .ZN(new_n9926_));
  INV_X1     g09733(.I(new_n9802_), .ZN(new_n9927_));
  NAND2_X1   g09734(.A1(new_n9927_), .A2(new_n9763_), .ZN(new_n9928_));
  NAND2_X1   g09735(.A1(new_n9928_), .A2(new_n9926_), .ZN(new_n9929_));
  NAND2_X1   g09736(.A1(new_n9685_), .A2(new_n9713_), .ZN(new_n9930_));
  NAND2_X1   g09737(.A1(new_n9714_), .A2(new_n9683_), .ZN(new_n9931_));
  NAND2_X1   g09738(.A1(new_n9931_), .A2(new_n9930_), .ZN(new_n9932_));
  NAND2_X1   g09739(.A1(new_n9723_), .A2(new_n9536_), .ZN(new_n9933_));
  OAI21_X1   g09740(.A1(new_n9542_), .A2(new_n9549_), .B(new_n9933_), .ZN(new_n9934_));
  NAND2_X1   g09741(.A1(new_n9728_), .A2(new_n9727_), .ZN(new_n9935_));
  OAI21_X1   g09742(.A1(new_n9507_), .A2(new_n9514_), .B(new_n9935_), .ZN(new_n9936_));
  NAND2_X1   g09743(.A1(new_n9499_), .A2(new_n9525_), .ZN(new_n9937_));
  NAND2_X1   g09744(.A1(new_n9644_), .A2(new_n9571_), .ZN(new_n9938_));
  NAND2_X1   g09745(.A1(new_n9938_), .A2(new_n9937_), .ZN(new_n9939_));
  XOR2_X1    g09746(.A1(new_n9939_), .A2(new_n9936_), .Z(new_n9940_));
  XOR2_X1    g09747(.A1(new_n9940_), .A2(new_n9934_), .Z(new_n9941_));
  NOR2_X1    g09748(.A1(new_n9932_), .A2(new_n9941_), .ZN(new_n9942_));
  NAND2_X1   g09749(.A1(new_n9932_), .A2(new_n9941_), .ZN(new_n9943_));
  INV_X1     g09750(.I(new_n9943_), .ZN(new_n9944_));
  NOR2_X1    g09751(.A1(new_n9944_), .A2(new_n9942_), .ZN(new_n9945_));
  NAND2_X1   g09752(.A1(new_n9700_), .A2(new_n9699_), .ZN(new_n9946_));
  AOI21_X1   g09753(.A1(\a[14] ), .A2(\a[62] ), .B(new_n9710_), .ZN(new_n9947_));
  INV_X1     g09754(.I(new_n9947_), .ZN(new_n9948_));
  NOR3_X1    g09755(.A1(new_n9709_), .A2(new_n759_), .A3(new_n7144_), .ZN(new_n9949_));
  INV_X1     g09756(.I(new_n9949_), .ZN(new_n9950_));
  NAND3_X1   g09757(.A1(new_n9946_), .A2(new_n9948_), .A3(new_n9950_), .ZN(new_n9951_));
  NAND2_X1   g09758(.A1(new_n9951_), .A2(new_n9950_), .ZN(new_n9952_));
  INV_X1     g09759(.I(new_n9952_), .ZN(new_n9953_));
  AOI22_X1   g09760(.A1(new_n9953_), .A2(new_n9948_), .B1(new_n9946_), .B2(new_n9951_), .ZN(new_n9954_));
  INV_X1     g09761(.I(new_n9954_), .ZN(new_n9955_));
  NAND2_X1   g09762(.A1(new_n9776_), .A2(new_n9784_), .ZN(new_n9956_));
  INV_X1     g09763(.I(new_n9785_), .ZN(new_n9957_));
  NAND2_X1   g09764(.A1(new_n9957_), .A2(new_n9794_), .ZN(new_n9958_));
  NAND2_X1   g09765(.A1(new_n9958_), .A2(new_n9956_), .ZN(new_n9959_));
  XOR2_X1    g09766(.A1(new_n9959_), .A2(new_n9955_), .Z(new_n9960_));
  NOR2_X1    g09767(.A1(new_n9680_), .A2(new_n9781_), .ZN(new_n9961_));
  NOR2_X1    g09768(.A1(new_n9679_), .A2(new_n9780_), .ZN(new_n9962_));
  NOR2_X1    g09769(.A1(new_n9961_), .A2(new_n9962_), .ZN(new_n9963_));
  NOR2_X1    g09770(.A1(new_n9963_), .A2(new_n9693_), .ZN(new_n9964_));
  NAND2_X1   g09771(.A1(new_n9963_), .A2(new_n9693_), .ZN(new_n9965_));
  INV_X1     g09772(.I(new_n9965_), .ZN(new_n9966_));
  NOR2_X1    g09773(.A1(new_n9966_), .A2(new_n9964_), .ZN(new_n9967_));
  XNOR2_X1   g09774(.A1(new_n9960_), .A2(new_n9967_), .ZN(new_n9968_));
  XOR2_X1    g09775(.A1(new_n9945_), .A2(new_n9968_), .Z(new_n9969_));
  XOR2_X1    g09776(.A1(new_n9929_), .A2(new_n9969_), .Z(new_n9970_));
  XOR2_X1    g09777(.A1(new_n9970_), .A2(new_n9924_), .Z(new_n9971_));
  XOR2_X1    g09778(.A1(new_n9858_), .A2(new_n9971_), .Z(new_n9972_));
  NAND2_X1   g09779(.A1(new_n9805_), .A2(new_n9803_), .ZN(new_n9973_));
  OAI21_X1   g09780(.A1(new_n9760_), .A2(new_n9807_), .B(new_n9973_), .ZN(new_n9974_));
  NOR2_X1    g09781(.A1(new_n9972_), .A2(new_n9974_), .ZN(new_n9975_));
  INV_X1     g09782(.I(new_n9975_), .ZN(new_n9976_));
  NAND2_X1   g09783(.A1(new_n9972_), .A2(new_n9974_), .ZN(new_n9977_));
  NAND2_X1   g09784(.A1(new_n9976_), .A2(new_n9977_), .ZN(new_n9978_));
  XOR2_X1    g09785(.A1(new_n9815_), .A2(new_n9978_), .Z(\asquared[77] ));
  OAI21_X1   g09786(.A1(new_n9814_), .A2(new_n9811_), .B(new_n9976_), .ZN(new_n9980_));
  NAND2_X1   g09787(.A1(new_n9980_), .A2(new_n9977_), .ZN(new_n9981_));
  NAND2_X1   g09788(.A1(new_n9817_), .A2(new_n9857_), .ZN(new_n9982_));
  NAND2_X1   g09789(.A1(new_n9858_), .A2(new_n9971_), .ZN(new_n9983_));
  NAND2_X1   g09790(.A1(new_n9983_), .A2(new_n9982_), .ZN(new_n9984_));
  INV_X1     g09791(.I(new_n9969_), .ZN(new_n9985_));
  NAND2_X1   g09792(.A1(new_n9929_), .A2(new_n9985_), .ZN(new_n9986_));
  OAI21_X1   g09793(.A1(new_n9970_), .A2(new_n9924_), .B(new_n9986_), .ZN(new_n9987_));
  NAND2_X1   g09794(.A1(new_n9861_), .A2(new_n9872_), .ZN(new_n9988_));
  NAND2_X1   g09795(.A1(new_n9873_), .A2(new_n9923_), .ZN(new_n9989_));
  NAND2_X1   g09796(.A1(new_n9989_), .A2(new_n9988_), .ZN(new_n9990_));
  OAI21_X1   g09797(.A1(new_n9942_), .A2(new_n9968_), .B(new_n9943_), .ZN(new_n9991_));
  NAND2_X1   g09798(.A1(new_n9959_), .A2(new_n9955_), .ZN(new_n9992_));
  NAND2_X1   g09799(.A1(new_n9960_), .A2(new_n9967_), .ZN(new_n9993_));
  NAND2_X1   g09800(.A1(new_n9993_), .A2(new_n9992_), .ZN(new_n9994_));
  AOI22_X1   g09801(.A1(\a[22] ), .A2(\a[55] ), .B1(\a[26] ), .B2(\a[51] ), .ZN(new_n9995_));
  NOR4_X1    g09802(.A1(new_n1175_), .A2(new_n1566_), .A3(new_n5135_), .A4(new_n5680_), .ZN(new_n9996_));
  NOR3_X1    g09803(.A1(new_n9995_), .A2(new_n2442_), .A3(new_n3666_), .ZN(new_n9997_));
  NOR2_X1    g09804(.A1(new_n9997_), .A2(new_n9996_), .ZN(new_n9998_));
  INV_X1     g09805(.I(new_n9998_), .ZN(new_n9999_));
  NOR2_X1    g09806(.A1(new_n2442_), .A2(new_n3666_), .ZN(new_n10000_));
  OAI21_X1   g09807(.A1(new_n9996_), .A2(new_n9995_), .B(new_n10000_), .ZN(new_n10001_));
  OAI21_X1   g09808(.A1(new_n9999_), .A2(new_n9995_), .B(new_n10001_), .ZN(new_n10002_));
  NOR2_X1    g09809(.A1(new_n1529_), .A2(new_n6127_), .ZN(new_n10003_));
  NOR2_X1    g09810(.A1(new_n1779_), .A2(new_n6563_), .ZN(new_n10004_));
  NOR2_X1    g09811(.A1(new_n1443_), .A2(new_n8421_), .ZN(new_n10005_));
  NOR2_X1    g09812(.A1(new_n10004_), .A2(new_n10005_), .ZN(new_n10006_));
  NOR2_X1    g09813(.A1(new_n10006_), .A2(new_n10003_), .ZN(new_n10007_));
  NAND2_X1   g09814(.A1(\a[25] ), .A2(\a[52] ), .ZN(new_n10008_));
  AOI22_X1   g09815(.A1(\a[23] ), .A2(\a[54] ), .B1(\a[24] ), .B2(\a[53] ), .ZN(new_n10009_));
  NOR2_X1    g09816(.A1(new_n10007_), .A2(new_n10003_), .ZN(new_n10010_));
  INV_X1     g09817(.I(new_n10010_), .ZN(new_n10011_));
  OAI22_X1   g09818(.A1(new_n10011_), .A2(new_n10009_), .B1(new_n10007_), .B2(new_n10008_), .ZN(new_n10012_));
  XOR2_X1    g09819(.A1(new_n10012_), .A2(new_n10002_), .Z(new_n10013_));
  AOI22_X1   g09820(.A1(\a[32] ), .A2(\a[45] ), .B1(\a[33] ), .B2(\a[44] ), .ZN(new_n10014_));
  NAND2_X1   g09821(.A1(\a[16] ), .A2(\a[61] ), .ZN(new_n10015_));
  NOR2_X1    g09822(.A1(new_n2637_), .A2(new_n4704_), .ZN(new_n10016_));
  NOR3_X1    g09823(.A1(new_n10016_), .A2(new_n10014_), .A3(new_n10015_), .ZN(new_n10017_));
  OAI22_X1   g09824(.A1(new_n2637_), .A2(new_n4704_), .B1(new_n10014_), .B2(new_n10015_), .ZN(new_n10018_));
  OAI22_X1   g09825(.A1(new_n10017_), .A2(new_n10015_), .B1(new_n10014_), .B2(new_n10018_), .ZN(new_n10019_));
  XNOR2_X1   g09826(.A1(new_n10013_), .A2(new_n10019_), .ZN(new_n10020_));
  NAND2_X1   g09827(.A1(new_n9867_), .A2(new_n9870_), .ZN(new_n10021_));
  NAND2_X1   g09828(.A1(new_n9871_), .A2(new_n9863_), .ZN(new_n10022_));
  NAND2_X1   g09829(.A1(new_n10022_), .A2(new_n10021_), .ZN(new_n10023_));
  NOR2_X1    g09830(.A1(new_n10023_), .A2(new_n10020_), .ZN(new_n10024_));
  INV_X1     g09831(.I(new_n10024_), .ZN(new_n10025_));
  NAND2_X1   g09832(.A1(new_n10023_), .A2(new_n10020_), .ZN(new_n10026_));
  NAND2_X1   g09833(.A1(new_n10025_), .A2(new_n10026_), .ZN(new_n10027_));
  NAND2_X1   g09834(.A1(new_n10027_), .A2(new_n9994_), .ZN(new_n10028_));
  NAND4_X1   g09835(.A1(new_n10025_), .A2(new_n9992_), .A3(new_n9993_), .A4(new_n10026_), .ZN(new_n10029_));
  AOI21_X1   g09836(.A1(new_n10028_), .A2(new_n10029_), .B(new_n9991_), .ZN(new_n10030_));
  NAND3_X1   g09837(.A1(new_n9991_), .A2(new_n10028_), .A3(new_n10029_), .ZN(new_n10031_));
  INV_X1     g09838(.I(new_n10031_), .ZN(new_n10032_));
  NOR2_X1    g09839(.A1(new_n10032_), .A2(new_n10030_), .ZN(new_n10033_));
  XOR2_X1    g09840(.A1(new_n9990_), .A2(new_n10033_), .Z(new_n10034_));
  XOR2_X1    g09841(.A1(new_n9987_), .A2(new_n10034_), .Z(new_n10035_));
  NOR2_X1    g09842(.A1(new_n9826_), .A2(new_n9850_), .ZN(new_n10036_));
  NAND2_X1   g09843(.A1(new_n9826_), .A2(new_n9850_), .ZN(new_n10037_));
  OAI21_X1   g09844(.A1(new_n9823_), .A2(new_n10036_), .B(new_n10037_), .ZN(new_n10038_));
  NAND2_X1   g09845(.A1(new_n9905_), .A2(new_n9912_), .ZN(new_n10039_));
  NAND2_X1   g09846(.A1(new_n9913_), .A2(new_n9919_), .ZN(new_n10040_));
  NAND2_X1   g09847(.A1(new_n10040_), .A2(new_n10039_), .ZN(new_n10041_));
  NAND2_X1   g09848(.A1(new_n9890_), .A2(new_n9793_), .ZN(new_n10042_));
  NAND2_X1   g09849(.A1(new_n9893_), .A2(new_n10042_), .ZN(new_n10043_));
  NOR2_X1    g09850(.A1(new_n10043_), .A2(new_n9952_), .ZN(new_n10044_));
  NAND2_X1   g09851(.A1(new_n10043_), .A2(new_n9952_), .ZN(new_n10045_));
  INV_X1     g09852(.I(new_n10045_), .ZN(new_n10046_));
  NOR2_X1    g09853(.A1(new_n10046_), .A2(new_n10044_), .ZN(new_n10047_));
  NAND2_X1   g09854(.A1(new_n10047_), .A2(new_n10041_), .ZN(new_n10048_));
  INV_X1     g09855(.I(new_n10048_), .ZN(new_n10049_));
  NOR2_X1    g09856(.A1(new_n10047_), .A2(new_n10041_), .ZN(new_n10050_));
  NOR2_X1    g09857(.A1(new_n10049_), .A2(new_n10050_), .ZN(new_n10051_));
  XOR2_X1    g09858(.A1(new_n10038_), .A2(new_n10051_), .Z(new_n10052_));
  NAND2_X1   g09859(.A1(new_n1815_), .A2(new_n4902_), .ZN(new_n10053_));
  NAND2_X1   g09860(.A1(new_n2103_), .A2(new_n5154_), .ZN(new_n10054_));
  AOI22_X1   g09861(.A1(new_n10053_), .A2(new_n10054_), .B1(new_n2105_), .B2(new_n4980_), .ZN(new_n10055_));
  NAND2_X1   g09862(.A1(\a[27] ), .A2(\a[50] ), .ZN(new_n10056_));
  AOI22_X1   g09863(.A1(\a[28] ), .A2(\a[49] ), .B1(\a[29] ), .B2(\a[48] ), .ZN(new_n10057_));
  NAND2_X1   g09864(.A1(new_n2105_), .A2(new_n4980_), .ZN(new_n10058_));
  NAND3_X1   g09865(.A1(new_n10058_), .A2(new_n10053_), .A3(new_n10054_), .ZN(new_n10059_));
  OAI22_X1   g09866(.A1(new_n10055_), .A2(new_n10056_), .B1(new_n10059_), .B2(new_n10057_), .ZN(new_n10060_));
  OAI22_X1   g09867(.A1(new_n1376_), .A2(new_n6804_), .B1(new_n1379_), .B2(new_n6318_), .ZN(new_n10061_));
  OAI21_X1   g09868(.A1(new_n1382_), .A2(new_n8161_), .B(new_n10061_), .ZN(new_n10062_));
  NAND3_X1   g09869(.A1(new_n10062_), .A2(\a[19] ), .A3(\a[58] ), .ZN(new_n10063_));
  AOI22_X1   g09870(.A1(\a[20] ), .A2(\a[57] ), .B1(\a[21] ), .B2(\a[56] ), .ZN(new_n10064_));
  NOR2_X1    g09871(.A1(new_n1382_), .A2(new_n8161_), .ZN(new_n10065_));
  NOR2_X1    g09872(.A1(new_n10061_), .A2(new_n10065_), .ZN(new_n10066_));
  INV_X1     g09873(.I(new_n10066_), .ZN(new_n10067_));
  OAI21_X1   g09874(.A1(new_n10064_), .A2(new_n10067_), .B(new_n10063_), .ZN(new_n10068_));
  XNOR2_X1   g09875(.A1(new_n10068_), .A2(new_n9911_), .ZN(new_n10069_));
  XNOR2_X1   g09876(.A1(new_n10069_), .A2(new_n10060_), .ZN(new_n10070_));
  NOR2_X1    g09877(.A1(new_n2051_), .A2(new_n7643_), .ZN(new_n10071_));
  NAND2_X1   g09878(.A1(new_n5888_), .A2(new_n10071_), .ZN(new_n10072_));
  NOR4_X1    g09879(.A1(new_n759_), .A2(new_n2030_), .A3(new_n4312_), .A4(new_n7643_), .ZN(new_n10073_));
  NOR2_X1    g09880(.A1(new_n2438_), .A2(new_n4721_), .ZN(new_n10074_));
  OAI21_X1   g09881(.A1(new_n10074_), .A2(new_n10073_), .B(new_n10072_), .ZN(new_n10075_));
  NAND3_X1   g09882(.A1(new_n10075_), .A2(\a[30] ), .A3(\a[47] ), .ZN(new_n10076_));
  AOI22_X1   g09883(.A1(\a[14] ), .A2(\a[63] ), .B1(\a[31] ), .B2(\a[46] ), .ZN(new_n10077_));
  NAND2_X1   g09884(.A1(new_n10075_), .A2(new_n10072_), .ZN(new_n10078_));
  OAI21_X1   g09885(.A1(new_n10077_), .A2(new_n10078_), .B(new_n10076_), .ZN(new_n10079_));
  NAND2_X1   g09886(.A1(new_n3037_), .A2(new_n4534_), .ZN(new_n10080_));
  OAI22_X1   g09887(.A1(new_n3405_), .A2(new_n4667_), .B1(new_n4190_), .B2(new_n7757_), .ZN(new_n10081_));
  NAND2_X1   g09888(.A1(new_n10081_), .A2(new_n10080_), .ZN(new_n10082_));
  NAND3_X1   g09889(.A1(new_n10082_), .A2(\a[35] ), .A3(\a[42] ), .ZN(new_n10083_));
  AOI21_X1   g09890(.A1(\a[36] ), .A2(\a[41] ), .B(new_n4741_), .ZN(new_n10084_));
  NAND2_X1   g09891(.A1(new_n10082_), .A2(new_n10080_), .ZN(new_n10085_));
  OAI21_X1   g09892(.A1(new_n10084_), .A2(new_n10085_), .B(new_n10083_), .ZN(new_n10086_));
  XNOR2_X1   g09893(.A1(new_n10086_), .A2(new_n10079_), .ZN(new_n10087_));
  AOI21_X1   g09894(.A1(\a[15] ), .A2(\a[62] ), .B(\a[39] ), .ZN(new_n10088_));
  NOR2_X1    g09895(.A1(new_n5534_), .A2(new_n7144_), .ZN(new_n10089_));
  NOR2_X1    g09896(.A1(new_n10089_), .A2(new_n4209_), .ZN(new_n10090_));
  INV_X1     g09897(.I(new_n10090_), .ZN(new_n10091_));
  NAND2_X1   g09898(.A1(new_n10089_), .A2(new_n4209_), .ZN(new_n10092_));
  OAI21_X1   g09899(.A1(new_n10091_), .A2(new_n10088_), .B(new_n10092_), .ZN(new_n10093_));
  INV_X1     g09900(.I(new_n10093_), .ZN(new_n10094_));
  XOR2_X1    g09901(.A1(new_n10087_), .A2(new_n10094_), .Z(new_n10095_));
  NAND2_X1   g09902(.A1(new_n9939_), .A2(new_n9936_), .ZN(new_n10096_));
  NAND2_X1   g09903(.A1(new_n9940_), .A2(new_n9934_), .ZN(new_n10097_));
  NAND2_X1   g09904(.A1(new_n10097_), .A2(new_n10096_), .ZN(new_n10098_));
  XOR2_X1    g09905(.A1(new_n10098_), .A2(new_n10095_), .Z(new_n10099_));
  XOR2_X1    g09906(.A1(new_n10099_), .A2(new_n10070_), .Z(new_n10100_));
  XNOR2_X1   g09907(.A1(new_n10052_), .A2(new_n10100_), .ZN(new_n10101_));
  NOR2_X1    g09908(.A1(new_n9822_), .A2(new_n9852_), .ZN(new_n10102_));
  NOR2_X1    g09909(.A1(new_n9856_), .A2(new_n10102_), .ZN(new_n10103_));
  XOR2_X1    g09910(.A1(new_n9904_), .A2(new_n9848_), .Z(new_n10104_));
  XOR2_X1    g09911(.A1(new_n10104_), .A2(new_n9839_), .Z(new_n10105_));
  NOR2_X1    g09912(.A1(new_n9880_), .A2(new_n9889_), .ZN(new_n10106_));
  NOR2_X1    g09913(.A1(new_n9879_), .A2(new_n9888_), .ZN(new_n10107_));
  NOR2_X1    g09914(.A1(new_n10106_), .A2(new_n10107_), .ZN(new_n10108_));
  NAND2_X1   g09915(.A1(new_n10108_), .A2(new_n9831_), .ZN(new_n10109_));
  INV_X1     g09916(.I(new_n10109_), .ZN(new_n10110_));
  NOR2_X1    g09917(.A1(new_n10108_), .A2(new_n9831_), .ZN(new_n10111_));
  NOR2_X1    g09918(.A1(new_n10110_), .A2(new_n10111_), .ZN(new_n10112_));
  NAND2_X1   g09919(.A1(new_n9841_), .A2(new_n9833_), .ZN(new_n10113_));
  NAND2_X1   g09920(.A1(new_n9842_), .A2(new_n9849_), .ZN(new_n10114_));
  NAND2_X1   g09921(.A1(new_n10114_), .A2(new_n10113_), .ZN(new_n10115_));
  XOR2_X1    g09922(.A1(new_n10115_), .A2(new_n10112_), .Z(new_n10116_));
  XOR2_X1    g09923(.A1(new_n10116_), .A2(new_n10105_), .Z(new_n10117_));
  NAND2_X1   g09924(.A1(new_n9898_), .A2(new_n9921_), .ZN(new_n10118_));
  NAND2_X1   g09925(.A1(new_n9922_), .A2(new_n9895_), .ZN(new_n10119_));
  NAND2_X1   g09926(.A1(new_n10119_), .A2(new_n10118_), .ZN(new_n10120_));
  NOR2_X1    g09927(.A1(new_n9966_), .A2(new_n9962_), .ZN(new_n10121_));
  NAND2_X1   g09928(.A1(new_n9670_), .A2(new_n9662_), .ZN(new_n10122_));
  NAND2_X1   g09929(.A1(new_n9862_), .A2(new_n9775_), .ZN(new_n10123_));
  NAND2_X1   g09930(.A1(new_n10123_), .A2(new_n10122_), .ZN(new_n10124_));
  NOR2_X1    g09931(.A1(new_n1275_), .A2(new_n7452_), .ZN(new_n10125_));
  INV_X1     g09932(.I(new_n10125_), .ZN(new_n10126_));
  NOR2_X1    g09933(.A1(new_n884_), .A2(new_n6548_), .ZN(new_n10127_));
  NOR2_X1    g09934(.A1(new_n1023_), .A2(new_n6723_), .ZN(new_n10128_));
  OAI21_X1   g09935(.A1(new_n10127_), .A2(new_n10128_), .B(new_n10126_), .ZN(new_n10129_));
  XNOR2_X1   g09936(.A1(new_n9917_), .A2(new_n10129_), .ZN(new_n10130_));
  INV_X1     g09937(.I(new_n10130_), .ZN(new_n10131_));
  XOR2_X1    g09938(.A1(new_n10124_), .A2(new_n10131_), .Z(new_n10132_));
  XNOR2_X1   g09939(.A1(new_n10132_), .A2(new_n10121_), .ZN(new_n10133_));
  XOR2_X1    g09940(.A1(new_n10120_), .A2(new_n10133_), .Z(new_n10134_));
  OR2_X2     g09941(.A1(new_n10134_), .A2(new_n10117_), .Z(new_n10135_));
  NAND2_X1   g09942(.A1(new_n10134_), .A2(new_n10117_), .ZN(new_n10136_));
  AND2_X2    g09943(.A1(new_n10135_), .A2(new_n10136_), .Z(new_n10137_));
  INV_X1     g09944(.I(new_n10137_), .ZN(new_n10138_));
  XOR2_X1    g09945(.A1(new_n10103_), .A2(new_n10138_), .Z(new_n10139_));
  XNOR2_X1   g09946(.A1(new_n10139_), .A2(new_n10101_), .ZN(new_n10140_));
  XOR2_X1    g09947(.A1(new_n10035_), .A2(new_n10140_), .Z(new_n10141_));
  NOR2_X1    g09948(.A1(new_n9984_), .A2(new_n10141_), .ZN(new_n10142_));
  NAND2_X1   g09949(.A1(new_n9984_), .A2(new_n10141_), .ZN(new_n10143_));
  INV_X1     g09950(.I(new_n10143_), .ZN(new_n10144_));
  NOR2_X1    g09951(.A1(new_n10144_), .A2(new_n10142_), .ZN(new_n10145_));
  XOR2_X1    g09952(.A1(new_n9981_), .A2(new_n10145_), .Z(\asquared[78] ));
  AOI21_X1   g09953(.A1(new_n9980_), .A2(new_n9977_), .B(new_n10142_), .ZN(new_n10147_));
  NOR2_X1    g09954(.A1(new_n10147_), .A2(new_n10144_), .ZN(new_n10148_));
  NAND2_X1   g09955(.A1(new_n9987_), .A2(new_n10034_), .ZN(new_n10149_));
  NAND2_X1   g09956(.A1(new_n10035_), .A2(new_n10140_), .ZN(new_n10150_));
  NAND2_X1   g09957(.A1(new_n10150_), .A2(new_n10149_), .ZN(new_n10151_));
  OAI21_X1   g09958(.A1(new_n9856_), .A2(new_n10102_), .B(new_n10137_), .ZN(new_n10152_));
  INV_X1     g09959(.I(new_n10139_), .ZN(new_n10153_));
  OAI21_X1   g09960(.A1(new_n10153_), .A2(new_n10101_), .B(new_n10152_), .ZN(new_n10154_));
  NAND2_X1   g09961(.A1(new_n10038_), .A2(new_n10051_), .ZN(new_n10155_));
  NAND2_X1   g09962(.A1(new_n10052_), .A2(new_n10100_), .ZN(new_n10156_));
  NAND2_X1   g09963(.A1(new_n10120_), .A2(new_n10133_), .ZN(new_n10157_));
  NOR2_X1    g09964(.A1(new_n10049_), .A2(new_n10046_), .ZN(new_n10158_));
  NAND2_X1   g09965(.A1(new_n1378_), .A2(new_n7203_), .ZN(new_n10159_));
  NOR3_X1    g09966(.A1(new_n5265_), .A2(new_n6298_), .A3(new_n6723_), .ZN(new_n10160_));
  NOR2_X1    g09967(.A1(new_n7452_), .A2(new_n1092_), .ZN(new_n10161_));
  OAI21_X1   g09968(.A1(new_n10160_), .A2(new_n10161_), .B(new_n10159_), .ZN(new_n10162_));
  NAND3_X1   g09969(.A1(new_n10162_), .A2(\a[18] ), .A3(\a[60] ), .ZN(new_n10163_));
  AOI22_X1   g09970(.A1(\a[19] ), .A2(\a[59] ), .B1(\a[21] ), .B2(\a[57] ), .ZN(new_n10164_));
  NAND2_X1   g09971(.A1(new_n10162_), .A2(new_n10159_), .ZN(new_n10165_));
  OAI21_X1   g09972(.A1(new_n10164_), .A2(new_n10165_), .B(new_n10163_), .ZN(new_n10166_));
  NAND2_X1   g09973(.A1(new_n2105_), .A2(new_n5154_), .ZN(new_n10167_));
  INV_X1     g09974(.I(new_n7867_), .ZN(new_n10168_));
  OAI22_X1   g09975(.A1(new_n1816_), .A2(new_n10168_), .B1(new_n2189_), .B2(new_n5440_), .ZN(new_n10169_));
  NAND2_X1   g09976(.A1(new_n10169_), .A2(new_n10167_), .ZN(new_n10170_));
  NAND3_X1   g09977(.A1(new_n10170_), .A2(\a[27] ), .A3(\a[51] ), .ZN(new_n10171_));
  AOI22_X1   g09978(.A1(\a[28] ), .A2(\a[50] ), .B1(\a[29] ), .B2(\a[49] ), .ZN(new_n10172_));
  NAND2_X1   g09979(.A1(new_n10170_), .A2(new_n10167_), .ZN(new_n10173_));
  OAI21_X1   g09980(.A1(new_n10172_), .A2(new_n10173_), .B(new_n10171_), .ZN(new_n10174_));
  XOR2_X1    g09981(.A1(new_n10174_), .A2(new_n10166_), .Z(new_n10175_));
  OAI22_X1   g09982(.A1(new_n893_), .A2(new_n8049_), .B1(new_n7959_), .B2(new_n982_), .ZN(new_n10176_));
  OAI21_X1   g09983(.A1(new_n1428_), .A2(new_n7591_), .B(new_n10176_), .ZN(new_n10177_));
  NAND3_X1   g09984(.A1(new_n10177_), .A2(\a[15] ), .A3(\a[63] ), .ZN(new_n10178_));
  AOI22_X1   g09985(.A1(\a[16] ), .A2(\a[62] ), .B1(\a[17] ), .B2(\a[61] ), .ZN(new_n10179_));
  NOR2_X1    g09986(.A1(new_n1428_), .A2(new_n7591_), .ZN(new_n10180_));
  NOR2_X1    g09987(.A1(new_n10176_), .A2(new_n10180_), .ZN(new_n10181_));
  INV_X1     g09988(.I(new_n10181_), .ZN(new_n10182_));
  OAI21_X1   g09989(.A1(new_n10179_), .A2(new_n10182_), .B(new_n10178_), .ZN(new_n10183_));
  XNOR2_X1   g09990(.A1(new_n10175_), .A2(new_n10183_), .ZN(new_n10184_));
  AOI22_X1   g09991(.A1(\a[30] ), .A2(\a[48] ), .B1(\a[31] ), .B2(\a[47] ), .ZN(new_n10185_));
  INV_X1     g09992(.I(new_n10185_), .ZN(new_n10186_));
  NOR2_X1    g09993(.A1(new_n2438_), .A2(new_n4977_), .ZN(new_n10187_));
  NOR2_X1    g09994(.A1(new_n1043_), .A2(new_n6316_), .ZN(new_n10188_));
  AOI21_X1   g09995(.A1(new_n10186_), .A2(new_n10188_), .B(new_n10187_), .ZN(new_n10189_));
  INV_X1     g09996(.I(new_n10189_), .ZN(new_n10190_));
  OAI21_X1   g09997(.A1(new_n10187_), .A2(new_n10185_), .B(new_n10188_), .ZN(new_n10191_));
  OAI21_X1   g09998(.A1(new_n10190_), .A2(new_n10185_), .B(new_n10191_), .ZN(new_n10192_));
  NOR2_X1    g09999(.A1(new_n3932_), .A2(new_n4704_), .ZN(new_n10193_));
  NOR2_X1    g10000(.A1(new_n2637_), .A2(new_n4430_), .ZN(new_n10194_));
  NOR2_X1    g10001(.A1(new_n3375_), .A2(new_n6101_), .ZN(new_n10195_));
  NOR2_X1    g10002(.A1(new_n10194_), .A2(new_n10195_), .ZN(new_n10196_));
  NOR2_X1    g10003(.A1(new_n10196_), .A2(new_n10193_), .ZN(new_n10197_));
  AOI22_X1   g10004(.A1(\a[33] ), .A2(\a[45] ), .B1(\a[34] ), .B2(\a[44] ), .ZN(new_n10198_));
  NOR2_X1    g10005(.A1(new_n10197_), .A2(new_n10193_), .ZN(new_n10199_));
  INV_X1     g10006(.I(new_n10199_), .ZN(new_n10200_));
  OAI22_X1   g10007(.A1(new_n10200_), .A2(new_n10198_), .B1(new_n4428_), .B2(new_n10197_), .ZN(new_n10201_));
  XOR2_X1    g10008(.A1(new_n10201_), .A2(new_n10192_), .Z(new_n10202_));
  NAND3_X1   g10009(.A1(new_n4351_), .A2(\a[53] ), .A3(\a[56] ), .ZN(new_n10203_));
  NAND2_X1   g10010(.A1(new_n1778_), .A2(new_n6126_), .ZN(new_n10204_));
  AOI22_X1   g10011(.A1(new_n10204_), .A2(new_n10203_), .B1(new_n1879_), .B2(new_n5857_), .ZN(new_n10205_));
  NAND2_X1   g10012(.A1(\a[25] ), .A2(\a[53] ), .ZN(new_n10206_));
  AOI22_X1   g10013(.A1(\a[22] ), .A2(\a[56] ), .B1(\a[24] ), .B2(\a[54] ), .ZN(new_n10207_));
  NAND2_X1   g10014(.A1(new_n1879_), .A2(new_n5857_), .ZN(new_n10208_));
  NAND3_X1   g10015(.A1(new_n10208_), .A2(new_n10204_), .A3(new_n10203_), .ZN(new_n10209_));
  OAI22_X1   g10016(.A1(new_n10205_), .A2(new_n10206_), .B1(new_n10209_), .B2(new_n10207_), .ZN(new_n10210_));
  XNOR2_X1   g10017(.A1(new_n10202_), .A2(new_n10210_), .ZN(new_n10211_));
  XNOR2_X1   g10018(.A1(new_n10211_), .A2(new_n10184_), .ZN(new_n10212_));
  NAND2_X1   g10019(.A1(new_n10158_), .A2(new_n10212_), .ZN(new_n10213_));
  NOR2_X1    g10020(.A1(new_n10158_), .A2(new_n10212_), .ZN(new_n10214_));
  INV_X1     g10021(.I(new_n10214_), .ZN(new_n10215_));
  AND2_X2    g10022(.A1(new_n10215_), .A2(new_n10213_), .Z(new_n10216_));
  INV_X1     g10023(.I(new_n10216_), .ZN(new_n10217_));
  AND3_X2    g10024(.A1(new_n10217_), .A2(new_n10157_), .A3(new_n10136_), .Z(new_n10218_));
  AOI21_X1   g10025(.A1(new_n10136_), .A2(new_n10157_), .B(new_n10217_), .ZN(new_n10219_));
  NOR2_X1    g10026(.A1(new_n10218_), .A2(new_n10219_), .ZN(new_n10220_));
  INV_X1     g10027(.I(new_n10220_), .ZN(new_n10221_));
  AND3_X2    g10028(.A1(new_n10221_), .A2(new_n10155_), .A3(new_n10156_), .Z(new_n10222_));
  AOI21_X1   g10029(.A1(new_n10155_), .A2(new_n10156_), .B(new_n10221_), .ZN(new_n10223_));
  NOR2_X1    g10030(.A1(new_n10222_), .A2(new_n10223_), .ZN(new_n10224_));
  XOR2_X1    g10031(.A1(new_n10154_), .A2(new_n10224_), .Z(new_n10225_));
  NAND2_X1   g10032(.A1(new_n10098_), .A2(new_n10095_), .ZN(new_n10226_));
  NAND2_X1   g10033(.A1(new_n10099_), .A2(new_n10070_), .ZN(new_n10227_));
  NAND2_X1   g10034(.A1(new_n10227_), .A2(new_n10226_), .ZN(new_n10228_));
  INV_X1     g10035(.I(new_n10020_), .ZN(new_n10229_));
  NAND2_X1   g10036(.A1(new_n10023_), .A2(new_n10229_), .ZN(new_n10230_));
  NAND2_X1   g10037(.A1(new_n10028_), .A2(new_n10230_), .ZN(new_n10231_));
  XOR2_X1    g10038(.A1(new_n10231_), .A2(new_n10228_), .Z(new_n10232_));
  NAND2_X1   g10039(.A1(new_n9904_), .A2(new_n9848_), .ZN(new_n10233_));
  NAND2_X1   g10040(.A1(new_n10104_), .A2(new_n9839_), .ZN(new_n10234_));
  NAND2_X1   g10041(.A1(new_n10234_), .A2(new_n10233_), .ZN(new_n10235_));
  AOI22_X1   g10042(.A1(\a[35] ), .A2(\a[43] ), .B1(\a[36] ), .B2(\a[42] ), .ZN(new_n10236_));
  INV_X1     g10043(.I(new_n10236_), .ZN(new_n10237_));
  NOR2_X1    g10044(.A1(new_n3405_), .A2(new_n4181_), .ZN(new_n10238_));
  NOR2_X1    g10045(.A1(new_n1299_), .A2(new_n5680_), .ZN(new_n10239_));
  AOI21_X1   g10046(.A1(new_n10237_), .A2(new_n10239_), .B(new_n10238_), .ZN(new_n10240_));
  INV_X1     g10047(.I(new_n10240_), .ZN(new_n10241_));
  OAI21_X1   g10048(.A1(new_n10238_), .A2(new_n10236_), .B(new_n10239_), .ZN(new_n10242_));
  OAI21_X1   g10049(.A1(new_n10241_), .A2(new_n10236_), .B(new_n10242_), .ZN(new_n10243_));
  INV_X1     g10050(.I(new_n4879_), .ZN(new_n10244_));
  NAND2_X1   g10051(.A1(new_n3803_), .A2(new_n4534_), .ZN(new_n10245_));
  NOR2_X1    g10052(.A1(new_n1566_), .A2(new_n5175_), .ZN(new_n10246_));
  NAND2_X1   g10053(.A1(new_n4879_), .A2(new_n10246_), .ZN(new_n10247_));
  NOR3_X1    g10054(.A1(new_n3223_), .A2(new_n1566_), .A3(new_n5175_), .ZN(new_n10248_));
  AOI21_X1   g10055(.A1(new_n10245_), .A2(new_n10247_), .B(new_n10248_), .ZN(new_n10249_));
  NAND2_X1   g10056(.A1(new_n10245_), .A2(new_n10247_), .ZN(new_n10250_));
  NOR2_X1    g10057(.A1(new_n10250_), .A2(new_n10248_), .ZN(new_n10251_));
  OAI21_X1   g10058(.A1(new_n3222_), .A2(new_n10246_), .B(new_n10251_), .ZN(new_n10252_));
  OAI21_X1   g10059(.A1(new_n10244_), .A2(new_n10249_), .B(new_n10252_), .ZN(new_n10253_));
  XNOR2_X1   g10060(.A1(new_n10253_), .A2(new_n10243_), .ZN(new_n10254_));
  XNOR2_X1   g10061(.A1(new_n10235_), .A2(new_n10254_), .ZN(new_n10255_));
  NAND2_X1   g10062(.A1(new_n10124_), .A2(new_n10131_), .ZN(new_n10256_));
  INV_X1     g10063(.I(new_n10132_), .ZN(new_n10257_));
  OAI21_X1   g10064(.A1(new_n10257_), .A2(new_n10121_), .B(new_n10256_), .ZN(new_n10258_));
  OAI21_X1   g10065(.A1(new_n9917_), .A2(new_n10129_), .B(new_n10126_), .ZN(new_n10259_));
  XOR2_X1    g10066(.A1(new_n10066_), .A2(new_n9998_), .Z(new_n10260_));
  XOR2_X1    g10067(.A1(new_n10260_), .A2(new_n10259_), .Z(new_n10261_));
  NOR2_X1    g10068(.A1(new_n10258_), .A2(new_n10261_), .ZN(new_n10262_));
  NAND2_X1   g10069(.A1(new_n10258_), .A2(new_n10261_), .ZN(new_n10263_));
  INV_X1     g10070(.I(new_n10263_), .ZN(new_n10264_));
  NOR2_X1    g10071(.A1(new_n10264_), .A2(new_n10262_), .ZN(new_n10265_));
  NAND2_X1   g10072(.A1(new_n10265_), .A2(new_n10255_), .ZN(new_n10266_));
  INV_X1     g10073(.I(new_n10266_), .ZN(new_n10267_));
  NOR2_X1    g10074(.A1(new_n10265_), .A2(new_n10255_), .ZN(new_n10268_));
  NOR2_X1    g10075(.A1(new_n10267_), .A2(new_n10268_), .ZN(new_n10269_));
  XNOR2_X1   g10076(.A1(new_n10232_), .A2(new_n10269_), .ZN(new_n10270_));
  NAND2_X1   g10077(.A1(new_n9990_), .A2(new_n10033_), .ZN(new_n10271_));
  NAND2_X1   g10078(.A1(new_n10271_), .A2(new_n10031_), .ZN(new_n10272_));
  XOR2_X1    g10079(.A1(new_n10085_), .A2(new_n10091_), .Z(new_n10273_));
  XOR2_X1    g10080(.A1(new_n10273_), .A2(new_n10011_), .Z(new_n10274_));
  INV_X1     g10081(.I(new_n10274_), .ZN(new_n10275_));
  XOR2_X1    g10082(.A1(new_n10078_), .A2(new_n10059_), .Z(new_n10276_));
  XOR2_X1    g10083(.A1(new_n10276_), .A2(new_n10018_), .Z(new_n10277_));
  NOR2_X1    g10084(.A1(new_n10110_), .A2(new_n10107_), .ZN(new_n10278_));
  XNOR2_X1   g10085(.A1(new_n10278_), .A2(new_n10277_), .ZN(new_n10279_));
  INV_X1     g10086(.I(new_n10279_), .ZN(new_n10280_));
  NOR2_X1    g10087(.A1(new_n10280_), .A2(new_n10275_), .ZN(new_n10281_));
  INV_X1     g10088(.I(new_n10281_), .ZN(new_n10282_));
  NAND2_X1   g10089(.A1(new_n10280_), .A2(new_n10275_), .ZN(new_n10283_));
  AND2_X2    g10090(.A1(new_n10282_), .A2(new_n10283_), .Z(new_n10284_));
  NAND2_X1   g10091(.A1(new_n10012_), .A2(new_n10002_), .ZN(new_n10285_));
  NAND2_X1   g10092(.A1(new_n10013_), .A2(new_n10019_), .ZN(new_n10286_));
  NAND2_X1   g10093(.A1(new_n10286_), .A2(new_n10285_), .ZN(new_n10287_));
  NAND2_X1   g10094(.A1(new_n10086_), .A2(new_n10079_), .ZN(new_n10288_));
  OAI21_X1   g10095(.A1(new_n10087_), .A2(new_n10094_), .B(new_n10288_), .ZN(new_n10289_));
  INV_X1     g10096(.I(new_n10069_), .ZN(new_n10290_));
  NAND2_X1   g10097(.A1(new_n10290_), .A2(new_n10060_), .ZN(new_n10291_));
  NAND2_X1   g10098(.A1(new_n10068_), .A2(new_n9911_), .ZN(new_n10292_));
  NAND2_X1   g10099(.A1(new_n10291_), .A2(new_n10292_), .ZN(new_n10293_));
  XOR2_X1    g10100(.A1(new_n10293_), .A2(new_n10289_), .Z(new_n10294_));
  XOR2_X1    g10101(.A1(new_n10294_), .A2(new_n10287_), .Z(new_n10295_));
  NAND2_X1   g10102(.A1(new_n10115_), .A2(new_n10112_), .ZN(new_n10296_));
  NAND2_X1   g10103(.A1(new_n10116_), .A2(new_n10105_), .ZN(new_n10297_));
  NAND2_X1   g10104(.A1(new_n10297_), .A2(new_n10296_), .ZN(new_n10298_));
  XOR2_X1    g10105(.A1(new_n10295_), .A2(new_n10298_), .Z(new_n10299_));
  NAND2_X1   g10106(.A1(new_n10299_), .A2(new_n10284_), .ZN(new_n10300_));
  OR2_X2     g10107(.A1(new_n10299_), .A2(new_n10284_), .Z(new_n10301_));
  AND2_X2    g10108(.A1(new_n10301_), .A2(new_n10300_), .Z(new_n10302_));
  XOR2_X1    g10109(.A1(new_n10272_), .A2(new_n10302_), .Z(new_n10303_));
  XNOR2_X1   g10110(.A1(new_n10303_), .A2(new_n10270_), .ZN(new_n10304_));
  XNOR2_X1   g10111(.A1(new_n10225_), .A2(new_n10304_), .ZN(new_n10305_));
  INV_X1     g10112(.I(new_n10305_), .ZN(new_n10306_));
  NOR2_X1    g10113(.A1(new_n10306_), .A2(new_n10151_), .ZN(new_n10307_));
  INV_X1     g10114(.I(new_n10307_), .ZN(new_n10308_));
  NAND2_X1   g10115(.A1(new_n10306_), .A2(new_n10151_), .ZN(new_n10309_));
  NAND2_X1   g10116(.A1(new_n10308_), .A2(new_n10309_), .ZN(new_n10310_));
  XOR2_X1    g10117(.A1(new_n10148_), .A2(new_n10310_), .Z(\asquared[79] ));
  OAI21_X1   g10118(.A1(new_n10147_), .A2(new_n10144_), .B(new_n10308_), .ZN(new_n10312_));
  NAND2_X1   g10119(.A1(new_n10312_), .A2(new_n10309_), .ZN(new_n10313_));
  NAND2_X1   g10120(.A1(new_n10154_), .A2(new_n10224_), .ZN(new_n10314_));
  NAND2_X1   g10121(.A1(new_n10225_), .A2(new_n10304_), .ZN(new_n10315_));
  NAND2_X1   g10122(.A1(new_n10315_), .A2(new_n10314_), .ZN(new_n10316_));
  NOR2_X1    g10123(.A1(new_n10223_), .A2(new_n10219_), .ZN(new_n10317_));
  NAND2_X1   g10124(.A1(new_n10231_), .A2(new_n10228_), .ZN(new_n10318_));
  NAND2_X1   g10125(.A1(new_n10232_), .A2(new_n10269_), .ZN(new_n10319_));
  NAND2_X1   g10126(.A1(new_n10319_), .A2(new_n10318_), .ZN(new_n10320_));
  NAND2_X1   g10127(.A1(new_n10201_), .A2(new_n10192_), .ZN(new_n10321_));
  NAND2_X1   g10128(.A1(new_n10202_), .A2(new_n10210_), .ZN(new_n10322_));
  NAND2_X1   g10129(.A1(new_n10322_), .A2(new_n10321_), .ZN(new_n10323_));
  NOR2_X1    g10130(.A1(new_n884_), .A2(new_n6897_), .ZN(new_n10324_));
  INV_X1     g10131(.I(new_n10324_), .ZN(new_n10325_));
  XOR2_X1    g10132(.A1(new_n10251_), .A2(new_n10325_), .Z(new_n10326_));
  NOR2_X1    g10133(.A1(new_n10326_), .A2(new_n10241_), .ZN(new_n10327_));
  INV_X1     g10134(.I(new_n10326_), .ZN(new_n10328_));
  NOR2_X1    g10135(.A1(new_n10328_), .A2(new_n10240_), .ZN(new_n10329_));
  NOR2_X1    g10136(.A1(new_n10329_), .A2(new_n10327_), .ZN(new_n10330_));
  XOR2_X1    g10137(.A1(new_n10189_), .A2(new_n10181_), .Z(new_n10331_));
  XOR2_X1    g10138(.A1(new_n10331_), .A2(new_n10200_), .Z(new_n10332_));
  NAND2_X1   g10139(.A1(new_n10332_), .A2(new_n10330_), .ZN(new_n10333_));
  INV_X1     g10140(.I(new_n10333_), .ZN(new_n10334_));
  NOR2_X1    g10141(.A1(new_n10332_), .A2(new_n10330_), .ZN(new_n10335_));
  NOR2_X1    g10142(.A1(new_n10334_), .A2(new_n10335_), .ZN(new_n10336_));
  NOR2_X1    g10143(.A1(new_n10323_), .A2(new_n10336_), .ZN(new_n10337_));
  NAND2_X1   g10144(.A1(new_n10323_), .A2(new_n10336_), .ZN(new_n10338_));
  INV_X1     g10145(.I(new_n10338_), .ZN(new_n10339_));
  NOR2_X1    g10146(.A1(new_n10339_), .A2(new_n10337_), .ZN(new_n10340_));
  OAI21_X1   g10147(.A1(new_n10184_), .A2(new_n10211_), .B(new_n10215_), .ZN(new_n10341_));
  NAND2_X1   g10148(.A1(new_n10260_), .A2(new_n10259_), .ZN(new_n10342_));
  OAI21_X1   g10149(.A1(new_n9998_), .A2(new_n10066_), .B(new_n10342_), .ZN(new_n10343_));
  AOI22_X1   g10150(.A1(\a[34] ), .A2(\a[45] ), .B1(\a[35] ), .B2(\a[44] ), .ZN(new_n10344_));
  INV_X1     g10151(.I(new_n10344_), .ZN(new_n10345_));
  NOR2_X1    g10152(.A1(new_n2746_), .A2(new_n4704_), .ZN(new_n10346_));
  NOR2_X1    g10153(.A1(new_n742_), .A2(new_n7643_), .ZN(new_n10347_));
  AOI21_X1   g10154(.A1(new_n10345_), .A2(new_n10347_), .B(new_n10346_), .ZN(new_n10348_));
  NAND2_X1   g10155(.A1(new_n10348_), .A2(new_n10345_), .ZN(new_n10349_));
  OAI21_X1   g10156(.A1(new_n10346_), .A2(new_n10344_), .B(new_n10347_), .ZN(new_n10350_));
  NAND2_X1   g10157(.A1(new_n10349_), .A2(new_n10350_), .ZN(new_n10351_));
  AOI22_X1   g10158(.A1(\a[23] ), .A2(\a[56] ), .B1(\a[27] ), .B2(\a[52] ), .ZN(new_n10352_));
  INV_X1     g10159(.I(new_n10352_), .ZN(new_n10353_));
  NOR2_X1    g10160(.A1(new_n1750_), .A2(new_n5856_), .ZN(new_n10354_));
  NAND2_X1   g10161(.A1(new_n9696_), .A2(new_n10354_), .ZN(new_n10355_));
  INV_X1     g10162(.I(new_n10355_), .ZN(new_n10356_));
  NOR2_X1    g10163(.A1(new_n2626_), .A2(new_n3666_), .ZN(new_n10357_));
  AOI21_X1   g10164(.A1(new_n10353_), .A2(new_n10357_), .B(new_n10356_), .ZN(new_n10358_));
  NAND2_X1   g10165(.A1(new_n10358_), .A2(new_n10353_), .ZN(new_n10359_));
  OAI21_X1   g10166(.A1(new_n10356_), .A2(new_n10352_), .B(new_n10357_), .ZN(new_n10360_));
  NAND2_X1   g10167(.A1(new_n10359_), .A2(new_n10360_), .ZN(new_n10361_));
  XNOR2_X1   g10168(.A1(new_n10351_), .A2(new_n10361_), .ZN(new_n10362_));
  INV_X1     g10169(.I(new_n10362_), .ZN(new_n10363_));
  NAND2_X1   g10170(.A1(new_n10363_), .A2(new_n10343_), .ZN(new_n10364_));
  INV_X1     g10171(.I(new_n10364_), .ZN(new_n10365_));
  NOR2_X1    g10172(.A1(new_n10363_), .A2(new_n10343_), .ZN(new_n10366_));
  NOR2_X1    g10173(.A1(new_n10365_), .A2(new_n10366_), .ZN(new_n10367_));
  XOR2_X1    g10174(.A1(new_n10173_), .A2(new_n10165_), .Z(new_n10368_));
  XOR2_X1    g10175(.A1(new_n10368_), .A2(new_n10209_), .Z(new_n10369_));
  NAND2_X1   g10176(.A1(new_n10253_), .A2(new_n10243_), .ZN(new_n10370_));
  INV_X1     g10177(.I(new_n10254_), .ZN(new_n10371_));
  NAND2_X1   g10178(.A1(new_n10371_), .A2(new_n10235_), .ZN(new_n10372_));
  NAND2_X1   g10179(.A1(new_n10372_), .A2(new_n10370_), .ZN(new_n10373_));
  AND2_X2    g10180(.A1(new_n10373_), .A2(new_n10369_), .Z(new_n10374_));
  NOR2_X1    g10181(.A1(new_n10373_), .A2(new_n10369_), .ZN(new_n10375_));
  NOR2_X1    g10182(.A1(new_n10374_), .A2(new_n10375_), .ZN(new_n10376_));
  NOR2_X1    g10183(.A1(new_n10376_), .A2(new_n10367_), .ZN(new_n10377_));
  NOR4_X1    g10184(.A1(new_n10375_), .A2(new_n10365_), .A3(new_n10374_), .A4(new_n10366_), .ZN(new_n10378_));
  NOR2_X1    g10185(.A1(new_n10377_), .A2(new_n10378_), .ZN(new_n10379_));
  NOR2_X1    g10186(.A1(new_n10341_), .A2(new_n10379_), .ZN(new_n10380_));
  NAND2_X1   g10187(.A1(new_n10341_), .A2(new_n10379_), .ZN(new_n10381_));
  INV_X1     g10188(.I(new_n10381_), .ZN(new_n10382_));
  NOR2_X1    g10189(.A1(new_n10382_), .A2(new_n10380_), .ZN(new_n10383_));
  NOR2_X1    g10190(.A1(new_n10383_), .A2(new_n10340_), .ZN(new_n10384_));
  NAND2_X1   g10191(.A1(new_n10383_), .A2(new_n10340_), .ZN(new_n10385_));
  INV_X1     g10192(.I(new_n10385_), .ZN(new_n10386_));
  NOR2_X1    g10193(.A1(new_n10386_), .A2(new_n10384_), .ZN(new_n10387_));
  XOR2_X1    g10194(.A1(new_n10387_), .A2(new_n10320_), .Z(new_n10388_));
  XNOR2_X1   g10195(.A1(new_n10317_), .A2(new_n10388_), .ZN(new_n10389_));
  INV_X1     g10196(.I(new_n10389_), .ZN(new_n10390_));
  NAND2_X1   g10197(.A1(new_n10272_), .A2(new_n10302_), .ZN(new_n10391_));
  INV_X1     g10198(.I(new_n10303_), .ZN(new_n10392_));
  OAI21_X1   g10199(.A1(new_n10392_), .A2(new_n10270_), .B(new_n10391_), .ZN(new_n10393_));
  NOR2_X1    g10200(.A1(new_n10267_), .A2(new_n10264_), .ZN(new_n10394_));
  NAND2_X1   g10201(.A1(new_n10174_), .A2(new_n10166_), .ZN(new_n10395_));
  NAND2_X1   g10202(.A1(new_n10175_), .A2(new_n10183_), .ZN(new_n10396_));
  NAND2_X1   g10203(.A1(new_n10396_), .A2(new_n10395_), .ZN(new_n10397_));
  NAND2_X1   g10204(.A1(new_n10078_), .A2(new_n10059_), .ZN(new_n10398_));
  NAND2_X1   g10205(.A1(new_n10276_), .A2(new_n10018_), .ZN(new_n10399_));
  NAND2_X1   g10206(.A1(new_n10399_), .A2(new_n10398_), .ZN(new_n10400_));
  NAND2_X1   g10207(.A1(new_n10085_), .A2(new_n10091_), .ZN(new_n10401_));
  NAND2_X1   g10208(.A1(new_n10273_), .A2(new_n10011_), .ZN(new_n10402_));
  NAND2_X1   g10209(.A1(new_n10402_), .A2(new_n10401_), .ZN(new_n10403_));
  XOR2_X1    g10210(.A1(new_n10403_), .A2(new_n10400_), .Z(new_n10404_));
  XOR2_X1    g10211(.A1(new_n10404_), .A2(new_n10397_), .Z(new_n10405_));
  NAND2_X1   g10212(.A1(new_n10293_), .A2(new_n10289_), .ZN(new_n10406_));
  NAND2_X1   g10213(.A1(new_n10294_), .A2(new_n10287_), .ZN(new_n10407_));
  NAND2_X1   g10214(.A1(new_n10407_), .A2(new_n10406_), .ZN(new_n10408_));
  XOR2_X1    g10215(.A1(new_n10408_), .A2(new_n10405_), .Z(new_n10409_));
  XOR2_X1    g10216(.A1(new_n10394_), .A2(new_n10409_), .Z(new_n10410_));
  INV_X1     g10217(.I(new_n10277_), .ZN(new_n10411_));
  NOR2_X1    g10218(.A1(new_n10411_), .A2(new_n10278_), .ZN(new_n10412_));
  NOR2_X1    g10219(.A1(new_n10281_), .A2(new_n10412_), .ZN(new_n10413_));
  NAND2_X1   g10220(.A1(\a[37] ), .A2(\a[42] ), .ZN(new_n10414_));
  NAND3_X1   g10221(.A1(new_n3550_), .A2(\a[37] ), .A3(\a[42] ), .ZN(new_n10415_));
  NAND2_X1   g10222(.A1(new_n3803_), .A2(new_n4372_), .ZN(new_n10416_));
  AOI22_X1   g10223(.A1(new_n10416_), .A2(new_n10415_), .B1(new_n4209_), .B2(new_n4534_), .ZN(new_n10417_));
  NAND2_X1   g10224(.A1(new_n4209_), .A2(new_n4534_), .ZN(new_n10418_));
  NAND3_X1   g10225(.A1(new_n10418_), .A2(new_n10416_), .A3(new_n10415_), .ZN(new_n10419_));
  AOI21_X1   g10226(.A1(\a[38] ), .A2(\a[41] ), .B(new_n3550_), .ZN(new_n10420_));
  OAI22_X1   g10227(.A1(new_n10417_), .A2(new_n10414_), .B1(new_n10419_), .B2(new_n10420_), .ZN(new_n10421_));
  OAI22_X1   g10228(.A1(new_n1779_), .A2(new_n6129_), .B1(new_n2081_), .B2(new_n6125_), .ZN(new_n10422_));
  OAI21_X1   g10229(.A1(new_n2177_), .A2(new_n6127_), .B(new_n10422_), .ZN(new_n10423_));
  NAND3_X1   g10230(.A1(new_n10423_), .A2(\a[24] ), .A3(\a[55] ), .ZN(new_n10424_));
  AOI22_X1   g10231(.A1(\a[25] ), .A2(\a[54] ), .B1(\a[26] ), .B2(\a[53] ), .ZN(new_n10425_));
  NOR2_X1    g10232(.A1(new_n2177_), .A2(new_n6127_), .ZN(new_n10426_));
  NOR2_X1    g10233(.A1(new_n10422_), .A2(new_n10426_), .ZN(new_n10427_));
  INV_X1     g10234(.I(new_n10427_), .ZN(new_n10428_));
  OAI21_X1   g10235(.A1(new_n10425_), .A2(new_n10428_), .B(new_n10424_), .ZN(new_n10429_));
  XNOR2_X1   g10236(.A1(new_n10429_), .A2(new_n10421_), .ZN(new_n10430_));
  AOI21_X1   g10237(.A1(\a[17] ), .A2(\a[62] ), .B(\a[40] ), .ZN(new_n10431_));
  NOR2_X1    g10238(.A1(new_n1718_), .A2(new_n5135_), .ZN(new_n10432_));
  INV_X1     g10239(.I(new_n10432_), .ZN(new_n10433_));
  NOR2_X1    g10240(.A1(new_n3221_), .A2(new_n7144_), .ZN(new_n10434_));
  INV_X1     g10241(.I(new_n10434_), .ZN(new_n10435_));
  NOR2_X1    g10242(.A1(new_n10435_), .A2(new_n1023_), .ZN(new_n10436_));
  NOR3_X1    g10243(.A1(new_n10436_), .A2(new_n10431_), .A3(new_n10433_), .ZN(new_n10437_));
  NOR2_X1    g10244(.A1(new_n10437_), .A2(new_n10436_), .ZN(new_n10438_));
  INV_X1     g10245(.I(new_n10438_), .ZN(new_n10439_));
  OAI22_X1   g10246(.A1(new_n10439_), .A2(new_n10431_), .B1(new_n10433_), .B2(new_n10437_), .ZN(new_n10440_));
  XOR2_X1    g10247(.A1(new_n10430_), .A2(new_n10440_), .Z(new_n10441_));
  OAI22_X1   g10248(.A1(new_n1376_), .A2(new_n7452_), .B1(new_n1379_), .B2(new_n7801_), .ZN(new_n10442_));
  OAI21_X1   g10249(.A1(new_n1382_), .A2(new_n7206_), .B(new_n10442_), .ZN(new_n10443_));
  NAND3_X1   g10250(.A1(new_n10443_), .A2(\a[19] ), .A3(\a[60] ), .ZN(new_n10444_));
  AOI22_X1   g10251(.A1(\a[20] ), .A2(\a[59] ), .B1(\a[21] ), .B2(\a[58] ), .ZN(new_n10445_));
  NOR2_X1    g10252(.A1(new_n1382_), .A2(new_n7206_), .ZN(new_n10446_));
  NOR2_X1    g10253(.A1(new_n10442_), .A2(new_n10446_), .ZN(new_n10447_));
  INV_X1     g10254(.I(new_n10447_), .ZN(new_n10448_));
  OAI21_X1   g10255(.A1(new_n10445_), .A2(new_n10448_), .B(new_n10444_), .ZN(new_n10449_));
  AOI22_X1   g10256(.A1(\a[29] ), .A2(\a[50] ), .B1(\a[30] ), .B2(\a[49] ), .ZN(new_n10450_));
  INV_X1     g10257(.I(new_n10450_), .ZN(new_n10451_));
  NOR2_X1    g10258(.A1(new_n2255_), .A2(new_n5155_), .ZN(new_n10452_));
  NOR2_X1    g10259(.A1(new_n1175_), .A2(new_n6298_), .ZN(new_n10453_));
  AOI21_X1   g10260(.A1(new_n10451_), .A2(new_n10453_), .B(new_n10452_), .ZN(new_n10454_));
  INV_X1     g10261(.I(new_n10454_), .ZN(new_n10455_));
  OAI21_X1   g10262(.A1(new_n10452_), .A2(new_n10450_), .B(new_n10453_), .ZN(new_n10456_));
  OAI21_X1   g10263(.A1(new_n10455_), .A2(new_n10450_), .B(new_n10456_), .ZN(new_n10457_));
  XNOR2_X1   g10264(.A1(new_n10449_), .A2(new_n10457_), .ZN(new_n10458_));
  NOR2_X1    g10265(.A1(new_n2637_), .A2(new_n4721_), .ZN(new_n10459_));
  AOI22_X1   g10266(.A1(new_n2275_), .A2(new_n6743_), .B1(new_n3210_), .B2(new_n4976_), .ZN(new_n10460_));
  NOR2_X1    g10267(.A1(new_n10459_), .A2(new_n10460_), .ZN(new_n10461_));
  NAND2_X1   g10268(.A1(\a[31] ), .A2(\a[48] ), .ZN(new_n10462_));
  AOI22_X1   g10269(.A1(\a[32] ), .A2(\a[47] ), .B1(\a[33] ), .B2(\a[46] ), .ZN(new_n10463_));
  NOR2_X1    g10270(.A1(new_n10461_), .A2(new_n10459_), .ZN(new_n10464_));
  INV_X1     g10271(.I(new_n10464_), .ZN(new_n10465_));
  OAI22_X1   g10272(.A1(new_n10465_), .A2(new_n10463_), .B1(new_n10461_), .B2(new_n10462_), .ZN(new_n10466_));
  XOR2_X1    g10273(.A1(new_n10458_), .A2(new_n10466_), .Z(new_n10467_));
  XOR2_X1    g10274(.A1(new_n10441_), .A2(new_n10467_), .Z(new_n10468_));
  XNOR2_X1   g10275(.A1(new_n10413_), .A2(new_n10468_), .ZN(new_n10469_));
  NAND2_X1   g10276(.A1(new_n10295_), .A2(new_n10298_), .ZN(new_n10470_));
  NAND2_X1   g10277(.A1(new_n10300_), .A2(new_n10470_), .ZN(new_n10471_));
  XOR2_X1    g10278(.A1(new_n10471_), .A2(new_n10469_), .Z(new_n10472_));
  INV_X1     g10279(.I(new_n10472_), .ZN(new_n10473_));
  OR2_X2     g10280(.A1(new_n10473_), .A2(new_n10410_), .Z(new_n10474_));
  NAND2_X1   g10281(.A1(new_n10473_), .A2(new_n10410_), .ZN(new_n10475_));
  AND2_X2    g10282(.A1(new_n10474_), .A2(new_n10475_), .Z(new_n10476_));
  INV_X1     g10283(.I(new_n10476_), .ZN(new_n10477_));
  NAND2_X1   g10284(.A1(new_n10393_), .A2(new_n10477_), .ZN(new_n10478_));
  NOR2_X1    g10285(.A1(new_n10393_), .A2(new_n10477_), .ZN(new_n10479_));
  INV_X1     g10286(.I(new_n10479_), .ZN(new_n10480_));
  AOI21_X1   g10287(.A1(new_n10480_), .A2(new_n10478_), .B(new_n10390_), .ZN(new_n10481_));
  INV_X1     g10288(.I(new_n10481_), .ZN(new_n10482_));
  NAND3_X1   g10289(.A1(new_n10480_), .A2(new_n10390_), .A3(new_n10478_), .ZN(new_n10483_));
  NAND2_X1   g10290(.A1(new_n10482_), .A2(new_n10483_), .ZN(new_n10484_));
  INV_X1     g10291(.I(new_n10484_), .ZN(new_n10485_));
  NOR2_X1    g10292(.A1(new_n10316_), .A2(new_n10485_), .ZN(new_n10486_));
  NAND2_X1   g10293(.A1(new_n10316_), .A2(new_n10485_), .ZN(new_n10487_));
  INV_X1     g10294(.I(new_n10487_), .ZN(new_n10488_));
  NOR2_X1    g10295(.A1(new_n10488_), .A2(new_n10486_), .ZN(new_n10489_));
  XOR2_X1    g10296(.A1(new_n10313_), .A2(new_n10489_), .Z(\asquared[80] ));
  AOI21_X1   g10297(.A1(new_n10312_), .A2(new_n10309_), .B(new_n10486_), .ZN(new_n10491_));
  NOR2_X1    g10298(.A1(new_n10491_), .A2(new_n10488_), .ZN(new_n10492_));
  NAND2_X1   g10299(.A1(new_n10393_), .A2(new_n10476_), .ZN(new_n10493_));
  NAND2_X1   g10300(.A1(new_n10482_), .A2(new_n10493_), .ZN(new_n10494_));
  NAND2_X1   g10301(.A1(new_n10471_), .A2(new_n10469_), .ZN(new_n10495_));
  NAND2_X1   g10302(.A1(new_n10474_), .A2(new_n10495_), .ZN(new_n10496_));
  NOR2_X1    g10303(.A1(new_n10251_), .A2(new_n10325_), .ZN(new_n10497_));
  NOR2_X1    g10304(.A1(new_n10329_), .A2(new_n10497_), .ZN(new_n10498_));
  NAND2_X1   g10305(.A1(new_n10173_), .A2(new_n10165_), .ZN(new_n10499_));
  NAND2_X1   g10306(.A1(new_n10368_), .A2(new_n10209_), .ZN(new_n10500_));
  NAND2_X1   g10307(.A1(new_n10500_), .A2(new_n10499_), .ZN(new_n10501_));
  NAND2_X1   g10308(.A1(new_n10331_), .A2(new_n10200_), .ZN(new_n10502_));
  OAI21_X1   g10309(.A1(new_n10181_), .A2(new_n10189_), .B(new_n10502_), .ZN(new_n10503_));
  XOR2_X1    g10310(.A1(new_n10501_), .A2(new_n10503_), .Z(new_n10504_));
  XNOR2_X1   g10311(.A1(new_n10504_), .A2(new_n10498_), .ZN(new_n10505_));
  INV_X1     g10312(.I(new_n10505_), .ZN(new_n10506_));
  NOR2_X1    g10313(.A1(new_n10378_), .A2(new_n10374_), .ZN(new_n10507_));
  NOR2_X1    g10314(.A1(new_n10339_), .A2(new_n10334_), .ZN(new_n10508_));
  XNOR2_X1   g10315(.A1(new_n10507_), .A2(new_n10508_), .ZN(new_n10509_));
  XOR2_X1    g10316(.A1(new_n10509_), .A2(new_n10506_), .Z(new_n10510_));
  NAND2_X1   g10317(.A1(new_n10447_), .A2(new_n10454_), .ZN(new_n10511_));
  NAND2_X1   g10318(.A1(new_n10448_), .A2(new_n10455_), .ZN(new_n10512_));
  AND2_X2    g10319(.A1(new_n10512_), .A2(new_n10511_), .Z(new_n10513_));
  XOR2_X1    g10320(.A1(new_n10513_), .A2(new_n10465_), .Z(new_n10514_));
  NAND2_X1   g10321(.A1(new_n10429_), .A2(new_n10421_), .ZN(new_n10515_));
  INV_X1     g10322(.I(new_n10440_), .ZN(new_n10516_));
  OAI21_X1   g10323(.A1(new_n10430_), .A2(new_n10516_), .B(new_n10515_), .ZN(new_n10517_));
  NAND2_X1   g10324(.A1(new_n10449_), .A2(new_n10457_), .ZN(new_n10518_));
  INV_X1     g10325(.I(new_n10466_), .ZN(new_n10519_));
  OAI21_X1   g10326(.A1(new_n10458_), .A2(new_n10519_), .B(new_n10518_), .ZN(new_n10520_));
  NOR2_X1    g10327(.A1(new_n10517_), .A2(new_n10520_), .ZN(new_n10521_));
  NAND2_X1   g10328(.A1(new_n10517_), .A2(new_n10520_), .ZN(new_n10522_));
  INV_X1     g10329(.I(new_n10522_), .ZN(new_n10523_));
  NOR2_X1    g10330(.A1(new_n10523_), .A2(new_n10521_), .ZN(new_n10524_));
  NAND2_X1   g10331(.A1(new_n10524_), .A2(new_n10514_), .ZN(new_n10525_));
  INV_X1     g10332(.I(new_n10525_), .ZN(new_n10526_));
  NOR2_X1    g10333(.A1(new_n10524_), .A2(new_n10514_), .ZN(new_n10527_));
  NOR2_X1    g10334(.A1(new_n10526_), .A2(new_n10527_), .ZN(new_n10528_));
  NOR2_X1    g10335(.A1(new_n10441_), .A2(new_n10467_), .ZN(new_n10529_));
  INV_X1     g10336(.I(new_n10468_), .ZN(new_n10530_));
  NOR2_X1    g10337(.A1(new_n10530_), .A2(new_n10413_), .ZN(new_n10531_));
  NOR2_X1    g10338(.A1(new_n10531_), .A2(new_n10529_), .ZN(new_n10532_));
  NAND2_X1   g10339(.A1(new_n10403_), .A2(new_n10400_), .ZN(new_n10533_));
  NAND2_X1   g10340(.A1(new_n10404_), .A2(new_n10397_), .ZN(new_n10534_));
  NAND2_X1   g10341(.A1(new_n10534_), .A2(new_n10533_), .ZN(new_n10535_));
  NAND2_X1   g10342(.A1(new_n10351_), .A2(new_n10361_), .ZN(new_n10536_));
  NAND2_X1   g10343(.A1(new_n10364_), .A2(new_n10536_), .ZN(new_n10537_));
  XOR2_X1    g10344(.A1(new_n10427_), .A2(new_n10348_), .Z(new_n10538_));
  XNOR2_X1   g10345(.A1(new_n10538_), .A2(new_n10358_), .ZN(new_n10539_));
  NOR2_X1    g10346(.A1(new_n10537_), .A2(new_n10539_), .ZN(new_n10540_));
  NAND2_X1   g10347(.A1(new_n10537_), .A2(new_n10539_), .ZN(new_n10541_));
  INV_X1     g10348(.I(new_n10541_), .ZN(new_n10542_));
  NOR2_X1    g10349(.A1(new_n10542_), .A2(new_n10540_), .ZN(new_n10543_));
  NOR2_X1    g10350(.A1(new_n10543_), .A2(new_n10535_), .ZN(new_n10544_));
  NAND2_X1   g10351(.A1(new_n10543_), .A2(new_n10535_), .ZN(new_n10545_));
  INV_X1     g10352(.I(new_n10545_), .ZN(new_n10546_));
  NOR2_X1    g10353(.A1(new_n10546_), .A2(new_n10544_), .ZN(new_n10547_));
  INV_X1     g10354(.I(new_n10547_), .ZN(new_n10548_));
  XOR2_X1    g10355(.A1(new_n10532_), .A2(new_n10548_), .Z(new_n10549_));
  NAND2_X1   g10356(.A1(new_n10549_), .A2(new_n10528_), .ZN(new_n10550_));
  INV_X1     g10357(.I(new_n10550_), .ZN(new_n10551_));
  NOR2_X1    g10358(.A1(new_n10549_), .A2(new_n10528_), .ZN(new_n10552_));
  NOR2_X1    g10359(.A1(new_n10551_), .A2(new_n10552_), .ZN(new_n10553_));
  XNOR2_X1   g10360(.A1(new_n10553_), .A2(new_n10510_), .ZN(new_n10554_));
  INV_X1     g10361(.I(new_n10554_), .ZN(new_n10555_));
  XOR2_X1    g10362(.A1(new_n10496_), .A2(new_n10555_), .Z(new_n10556_));
  NAND2_X1   g10363(.A1(new_n10387_), .A2(new_n10320_), .ZN(new_n10557_));
  INV_X1     g10364(.I(new_n10388_), .ZN(new_n10558_));
  OAI21_X1   g10365(.A1(new_n10558_), .A2(new_n10317_), .B(new_n10557_), .ZN(new_n10559_));
  NOR2_X1    g10366(.A1(new_n10386_), .A2(new_n10382_), .ZN(new_n10560_));
  INV_X1     g10367(.I(new_n10560_), .ZN(new_n10561_));
  NAND2_X1   g10368(.A1(new_n10408_), .A2(new_n10405_), .ZN(new_n10562_));
  NOR2_X1    g10369(.A1(new_n10408_), .A2(new_n10405_), .ZN(new_n10563_));
  OAI21_X1   g10370(.A1(new_n10394_), .A2(new_n10563_), .B(new_n10562_), .ZN(new_n10564_));
  NAND2_X1   g10371(.A1(new_n7590_), .A2(new_n1194_), .ZN(new_n10565_));
  NOR2_X1    g10372(.A1(new_n979_), .A2(new_n6897_), .ZN(new_n10566_));
  NOR2_X1    g10373(.A1(new_n884_), .A2(new_n7144_), .ZN(new_n10567_));
  OAI21_X1   g10374(.A1(new_n10566_), .A2(new_n10567_), .B(new_n10565_), .ZN(new_n10568_));
  XNOR2_X1   g10375(.A1(new_n10438_), .A2(new_n10568_), .ZN(new_n10569_));
  AOI22_X1   g10376(.A1(\a[17] ), .A2(\a[63] ), .B1(\a[29] ), .B2(\a[51] ), .ZN(new_n10570_));
  INV_X1     g10377(.I(new_n10570_), .ZN(new_n10571_));
  NOR2_X1    g10378(.A1(new_n1814_), .A2(new_n7643_), .ZN(new_n10572_));
  NAND2_X1   g10379(.A1(new_n6113_), .A2(new_n10572_), .ZN(new_n10573_));
  INV_X1     g10380(.I(new_n10573_), .ZN(new_n10574_));
  NOR2_X1    g10381(.A1(new_n2274_), .A2(new_n4312_), .ZN(new_n10575_));
  AOI21_X1   g10382(.A1(new_n10571_), .A2(new_n10575_), .B(new_n10574_), .ZN(new_n10576_));
  INV_X1     g10383(.I(new_n10576_), .ZN(new_n10577_));
  OAI21_X1   g10384(.A1(new_n10574_), .A2(new_n10570_), .B(new_n10575_), .ZN(new_n10578_));
  OAI21_X1   g10385(.A1(new_n10577_), .A2(new_n10570_), .B(new_n10578_), .ZN(new_n10579_));
  NOR2_X1    g10386(.A1(new_n3405_), .A2(new_n4704_), .ZN(new_n10580_));
  NOR2_X1    g10387(.A1(new_n2746_), .A2(new_n4430_), .ZN(new_n10581_));
  NOR2_X1    g10388(.A1(new_n5564_), .A2(new_n6101_), .ZN(new_n10582_));
  NOR2_X1    g10389(.A1(new_n10581_), .A2(new_n10582_), .ZN(new_n10583_));
  NOR2_X1    g10390(.A1(new_n10583_), .A2(new_n10580_), .ZN(new_n10584_));
  NAND2_X1   g10391(.A1(\a[34] ), .A2(\a[46] ), .ZN(new_n10585_));
  NOR2_X1    g10392(.A1(new_n4844_), .A2(new_n4871_), .ZN(new_n10586_));
  NOR2_X1    g10393(.A1(new_n10584_), .A2(new_n10580_), .ZN(new_n10587_));
  INV_X1     g10394(.I(new_n10587_), .ZN(new_n10588_));
  OAI22_X1   g10395(.A1(new_n10588_), .A2(new_n10586_), .B1(new_n10584_), .B2(new_n10585_), .ZN(new_n10589_));
  XNOR2_X1   g10396(.A1(new_n10589_), .A2(new_n10579_), .ZN(new_n10590_));
  XNOR2_X1   g10397(.A1(new_n10590_), .A2(new_n10569_), .ZN(new_n10591_));
  NOR2_X1    g10398(.A1(new_n1456_), .A2(new_n7206_), .ZN(new_n10592_));
  INV_X1     g10399(.I(new_n10592_), .ZN(new_n10593_));
  OAI22_X1   g10400(.A1(new_n1220_), .A2(new_n6548_), .B1(new_n1175_), .B2(new_n6316_), .ZN(new_n10594_));
  AOI22_X1   g10401(.A1(new_n10593_), .A2(new_n10594_), .B1(\a[20] ), .B2(\a[60] ), .ZN(new_n10595_));
  OAI22_X1   g10402(.A1(new_n1382_), .A2(new_n7452_), .B1(new_n2647_), .B2(new_n7801_), .ZN(new_n10596_));
  NAND2_X1   g10403(.A1(new_n10596_), .A2(new_n10593_), .ZN(new_n10597_));
  INV_X1     g10404(.I(new_n10597_), .ZN(new_n10598_));
  NOR2_X1    g10405(.A1(new_n10598_), .A2(new_n10595_), .ZN(new_n10599_));
  XOR2_X1    g10406(.A1(new_n10599_), .A2(new_n10419_), .Z(new_n10600_));
  OAI22_X1   g10407(.A1(new_n2202_), .A2(new_n4903_), .B1(new_n2438_), .B2(new_n5155_), .ZN(new_n10601_));
  OAI21_X1   g10408(.A1(new_n3833_), .A2(new_n4981_), .B(new_n10601_), .ZN(new_n10602_));
  NAND3_X1   g10409(.A1(new_n10602_), .A2(\a[30] ), .A3(\a[50] ), .ZN(new_n10603_));
  AOI22_X1   g10410(.A1(\a[31] ), .A2(\a[49] ), .B1(\a[32] ), .B2(\a[48] ), .ZN(new_n10604_));
  NOR2_X1    g10411(.A1(new_n3833_), .A2(new_n4981_), .ZN(new_n10605_));
  NOR2_X1    g10412(.A1(new_n10601_), .A2(new_n10605_), .ZN(new_n10606_));
  INV_X1     g10413(.I(new_n10606_), .ZN(new_n10607_));
  OAI21_X1   g10414(.A1(new_n10604_), .A2(new_n10607_), .B(new_n10603_), .ZN(new_n10608_));
  XNOR2_X1   g10415(.A1(new_n10600_), .A2(new_n10608_), .ZN(new_n10609_));
  NOR2_X1    g10416(.A1(new_n2081_), .A2(new_n6058_), .ZN(new_n10610_));
  NOR2_X1    g10417(.A1(new_n5617_), .A2(new_n6298_), .ZN(new_n10611_));
  INV_X1     g10418(.I(new_n10611_), .ZN(new_n10612_));
  NOR2_X1    g10419(.A1(new_n2084_), .A2(new_n10612_), .ZN(new_n10613_));
  NOR2_X1    g10420(.A1(new_n1529_), .A2(new_n8161_), .ZN(new_n10614_));
  NOR2_X1    g10421(.A1(new_n10613_), .A2(new_n10614_), .ZN(new_n10615_));
  NOR2_X1    g10422(.A1(new_n10615_), .A2(new_n10610_), .ZN(new_n10616_));
  NAND2_X1   g10423(.A1(\a[23] ), .A2(\a[57] ), .ZN(new_n10617_));
  AOI22_X1   g10424(.A1(\a[24] ), .A2(\a[56] ), .B1(\a[26] ), .B2(\a[54] ), .ZN(new_n10618_));
  NOR2_X1    g10425(.A1(new_n10616_), .A2(new_n10610_), .ZN(new_n10619_));
  INV_X1     g10426(.I(new_n10619_), .ZN(new_n10620_));
  OAI22_X1   g10427(.A1(new_n10620_), .A2(new_n10618_), .B1(new_n10616_), .B2(new_n10617_), .ZN(new_n10621_));
  AOI22_X1   g10428(.A1(\a[37] ), .A2(\a[43] ), .B1(\a[38] ), .B2(\a[42] ), .ZN(new_n10622_));
  NOR2_X1    g10429(.A1(new_n1441_), .A2(new_n5680_), .ZN(new_n10623_));
  INV_X1     g10430(.I(new_n10623_), .ZN(new_n10624_));
  OAI22_X1   g10431(.A1(new_n6140_), .A2(new_n4181_), .B1(new_n10624_), .B2(new_n10622_), .ZN(new_n10625_));
  NOR2_X1    g10432(.A1(new_n6140_), .A2(new_n4181_), .ZN(new_n10626_));
  OAI21_X1   g10433(.A1(new_n10626_), .A2(new_n10622_), .B(new_n10623_), .ZN(new_n10627_));
  OAI21_X1   g10434(.A1(new_n10625_), .A2(new_n10622_), .B(new_n10627_), .ZN(new_n10628_));
  XNOR2_X1   g10435(.A1(new_n10621_), .A2(new_n10628_), .ZN(new_n10629_));
  AOI22_X1   g10436(.A1(\a[27] ), .A2(\a[53] ), .B1(\a[28] ), .B2(\a[52] ), .ZN(new_n10630_));
  NOR2_X1    g10437(.A1(new_n2189_), .A2(new_n6563_), .ZN(new_n10631_));
  NOR3_X1    g10438(.A1(new_n10631_), .A2(new_n3329_), .A3(new_n10630_), .ZN(new_n10632_));
  NOR2_X1    g10439(.A1(new_n10632_), .A2(new_n10631_), .ZN(new_n10633_));
  INV_X1     g10440(.I(new_n10633_), .ZN(new_n10634_));
  OAI22_X1   g10441(.A1(new_n10634_), .A2(new_n10630_), .B1(new_n3329_), .B2(new_n10632_), .ZN(new_n10635_));
  XOR2_X1    g10442(.A1(new_n10629_), .A2(new_n10635_), .Z(new_n10636_));
  XNOR2_X1   g10443(.A1(new_n10636_), .A2(new_n10609_), .ZN(new_n10637_));
  XOR2_X1    g10444(.A1(new_n10637_), .A2(new_n10591_), .Z(new_n10638_));
  NOR2_X1    g10445(.A1(new_n10564_), .A2(new_n10638_), .ZN(new_n10639_));
  NAND2_X1   g10446(.A1(new_n10564_), .A2(new_n10638_), .ZN(new_n10640_));
  INV_X1     g10447(.I(new_n10640_), .ZN(new_n10641_));
  NOR2_X1    g10448(.A1(new_n10641_), .A2(new_n10639_), .ZN(new_n10642_));
  NOR2_X1    g10449(.A1(new_n10561_), .A2(new_n10642_), .ZN(new_n10643_));
  NAND2_X1   g10450(.A1(new_n10561_), .A2(new_n10642_), .ZN(new_n10644_));
  INV_X1     g10451(.I(new_n10644_), .ZN(new_n10645_));
  NOR2_X1    g10452(.A1(new_n10645_), .A2(new_n10643_), .ZN(new_n10646_));
  XOR2_X1    g10453(.A1(new_n10559_), .A2(new_n10646_), .Z(new_n10647_));
  XOR2_X1    g10454(.A1(new_n10647_), .A2(new_n10556_), .Z(new_n10648_));
  NAND2_X1   g10455(.A1(new_n10494_), .A2(new_n10648_), .ZN(new_n10649_));
  NOR2_X1    g10456(.A1(new_n10494_), .A2(new_n10648_), .ZN(new_n10650_));
  INV_X1     g10457(.I(new_n10650_), .ZN(new_n10651_));
  NAND2_X1   g10458(.A1(new_n10651_), .A2(new_n10649_), .ZN(new_n10652_));
  INV_X1     g10459(.I(new_n10309_), .ZN(new_n10653_));
  INV_X1     g10460(.I(new_n9977_), .ZN(new_n10654_));
  INV_X1     g10461(.I(new_n9461_), .ZN(new_n10655_));
  OAI21_X1   g10462(.A1(new_n9296_), .A2(new_n9288_), .B(new_n10655_), .ZN(new_n10656_));
  INV_X1     g10463(.I(new_n9634_), .ZN(new_n10657_));
  AOI21_X1   g10464(.A1(new_n10656_), .A2(new_n9462_), .B(new_n10657_), .ZN(new_n10658_));
  INV_X1     g10465(.I(new_n9809_), .ZN(new_n10659_));
  OAI21_X1   g10466(.A1(new_n10658_), .A2(new_n9632_), .B(new_n10659_), .ZN(new_n10660_));
  AOI21_X1   g10467(.A1(new_n10660_), .A2(new_n9810_), .B(new_n9975_), .ZN(new_n10661_));
  INV_X1     g10468(.I(new_n10142_), .ZN(new_n10662_));
  OAI21_X1   g10469(.A1(new_n10661_), .A2(new_n10654_), .B(new_n10662_), .ZN(new_n10663_));
  AOI21_X1   g10470(.A1(new_n10663_), .A2(new_n10143_), .B(new_n10307_), .ZN(new_n10664_));
  INV_X1     g10471(.I(new_n10486_), .ZN(new_n10665_));
  OAI21_X1   g10472(.A1(new_n10664_), .A2(new_n10653_), .B(new_n10665_), .ZN(new_n10666_));
  AOI21_X1   g10473(.A1(new_n10666_), .A2(new_n10487_), .B(new_n10650_), .ZN(new_n10667_));
  AOI22_X1   g10474(.A1(new_n10667_), .A2(new_n10649_), .B1(new_n10492_), .B2(new_n10652_), .ZN(\asquared[81] ));
  OAI21_X1   g10475(.A1(new_n10491_), .A2(new_n10488_), .B(new_n10651_), .ZN(new_n10669_));
  NAND2_X1   g10476(.A1(new_n10669_), .A2(new_n10649_), .ZN(new_n10670_));
  NAND2_X1   g10477(.A1(new_n10553_), .A2(new_n10510_), .ZN(new_n10671_));
  NAND2_X1   g10478(.A1(new_n10496_), .A2(new_n10555_), .ZN(new_n10672_));
  NAND2_X1   g10479(.A1(new_n10672_), .A2(new_n10671_), .ZN(new_n10673_));
  NOR2_X1    g10480(.A1(new_n10532_), .A2(new_n10548_), .ZN(new_n10674_));
  NOR2_X1    g10481(.A1(new_n10551_), .A2(new_n10674_), .ZN(new_n10675_));
  OAI22_X1   g10482(.A1(new_n1281_), .A2(new_n7959_), .B1(new_n5265_), .B2(new_n9031_), .ZN(new_n10676_));
  NAND2_X1   g10483(.A1(new_n1381_), .A2(new_n7453_), .ZN(new_n10677_));
  NAND2_X1   g10484(.A1(new_n10676_), .A2(new_n10677_), .ZN(new_n10678_));
  NAND3_X1   g10485(.A1(new_n10678_), .A2(\a[18] ), .A3(\a[63] ), .ZN(new_n10679_));
  AOI22_X1   g10486(.A1(\a[20] ), .A2(\a[61] ), .B1(\a[21] ), .B2(\a[60] ), .ZN(new_n10680_));
  NAND2_X1   g10487(.A1(new_n10678_), .A2(new_n10677_), .ZN(new_n10681_));
  OAI21_X1   g10488(.A1(new_n10680_), .A2(new_n10681_), .B(new_n10679_), .ZN(new_n10682_));
  NAND2_X1   g10489(.A1(\a[35] ), .A2(\a[46] ), .ZN(new_n10683_));
  NAND4_X1   g10490(.A1(\a[35] ), .A2(\a[37] ), .A3(\a[44] ), .A4(\a[46] ), .ZN(new_n10684_));
  NAND2_X1   g10491(.A1(new_n3232_), .A2(new_n4429_), .ZN(new_n10685_));
  AOI22_X1   g10492(.A1(new_n10685_), .A2(new_n10684_), .B1(new_n3037_), .B2(new_n4703_), .ZN(new_n10686_));
  AOI22_X1   g10493(.A1(\a[36] ), .A2(\a[45] ), .B1(\a[37] ), .B2(\a[44] ), .ZN(new_n10687_));
  NAND2_X1   g10494(.A1(new_n3037_), .A2(new_n4703_), .ZN(new_n10688_));
  NAND3_X1   g10495(.A1(new_n10688_), .A2(new_n10685_), .A3(new_n10684_), .ZN(new_n10689_));
  OAI22_X1   g10496(.A1(new_n10686_), .A2(new_n10683_), .B1(new_n10689_), .B2(new_n10687_), .ZN(new_n10690_));
  XNOR2_X1   g10497(.A1(new_n10682_), .A2(new_n10690_), .ZN(new_n10691_));
  AOI22_X1   g10498(.A1(\a[29] ), .A2(new_n10246_), .B1(new_n2412_), .B2(\a[53] ), .ZN(new_n10692_));
  INV_X1     g10499(.I(new_n10692_), .ZN(new_n10693_));
  AOI21_X1   g10500(.A1(new_n2105_), .A2(new_n5862_), .B(new_n5680_), .ZN(new_n10694_));
  NAND2_X1   g10501(.A1(new_n10693_), .A2(new_n10694_), .ZN(new_n10695_));
  OAI21_X1   g10502(.A1(new_n2679_), .A2(new_n6563_), .B(new_n10695_), .ZN(new_n10696_));
  INV_X1     g10503(.I(new_n10696_), .ZN(new_n10697_));
  OAI22_X1   g10504(.A1(new_n1718_), .A2(new_n5425_), .B1(new_n1814_), .B2(new_n5175_), .ZN(new_n10698_));
  NOR2_X1    g10505(.A1(new_n1566_), .A2(new_n5680_), .ZN(new_n10699_));
  AOI22_X1   g10506(.A1(new_n10697_), .A2(new_n10698_), .B1(new_n10695_), .B2(new_n10699_), .ZN(new_n10700_));
  XNOR2_X1   g10507(.A1(new_n10691_), .A2(new_n10700_), .ZN(new_n10701_));
  INV_X1     g10508(.I(new_n10701_), .ZN(new_n10702_));
  NAND2_X1   g10509(.A1(new_n10501_), .A2(new_n10503_), .ZN(new_n10703_));
  INV_X1     g10510(.I(new_n10504_), .ZN(new_n10704_));
  OAI21_X1   g10511(.A1(new_n10704_), .A2(new_n10498_), .B(new_n10703_), .ZN(new_n10705_));
  NOR3_X1    g10512(.A1(new_n979_), .A2(new_n3327_), .A3(new_n7144_), .ZN(new_n10706_));
  NAND2_X1   g10513(.A1(new_n10706_), .A2(new_n4534_), .ZN(new_n10707_));
  AOI21_X1   g10514(.A1(\a[19] ), .A2(\a[62] ), .B(\a[41] ), .ZN(new_n10708_));
  NOR2_X1    g10515(.A1(new_n10706_), .A2(new_n4534_), .ZN(new_n10709_));
  INV_X1     g10516(.I(new_n10709_), .ZN(new_n10710_));
  OAI21_X1   g10517(.A1(new_n10710_), .A2(new_n10708_), .B(new_n10707_), .ZN(new_n10711_));
  NOR2_X1    g10518(.A1(new_n1443_), .A2(new_n6318_), .ZN(new_n10712_));
  INV_X1     g10519(.I(new_n10712_), .ZN(new_n10713_));
  NOR2_X1    g10520(.A1(new_n5856_), .A2(new_n6548_), .ZN(new_n10714_));
  INV_X1     g10521(.I(new_n10714_), .ZN(new_n10715_));
  NOR3_X1    g10522(.A1(new_n10715_), .A2(new_n1175_), .A3(new_n1441_), .ZN(new_n10716_));
  NOR2_X1    g10523(.A1(new_n2385_), .A2(new_n7206_), .ZN(new_n10717_));
  OAI21_X1   g10524(.A1(new_n10716_), .A2(new_n10717_), .B(new_n10713_), .ZN(new_n10718_));
  NAND3_X1   g10525(.A1(new_n10718_), .A2(\a[22] ), .A3(\a[59] ), .ZN(new_n10719_));
  AOI22_X1   g10526(.A1(\a[23] ), .A2(\a[58] ), .B1(\a[25] ), .B2(\a[56] ), .ZN(new_n10720_));
  NAND2_X1   g10527(.A1(new_n10718_), .A2(new_n10713_), .ZN(new_n10721_));
  OAI21_X1   g10528(.A1(new_n10720_), .A2(new_n10721_), .B(new_n10719_), .ZN(new_n10722_));
  XNOR2_X1   g10529(.A1(new_n10722_), .A2(new_n10711_), .ZN(new_n10723_));
  AOI22_X1   g10530(.A1(\a[33] ), .A2(\a[48] ), .B1(\a[34] ), .B2(\a[47] ), .ZN(new_n10724_));
  NOR2_X1    g10531(.A1(new_n3932_), .A2(new_n4977_), .ZN(new_n10725_));
  NOR3_X1    g10532(.A1(new_n10725_), .A2(new_n8076_), .A3(new_n10724_), .ZN(new_n10726_));
  NOR2_X1    g10533(.A1(new_n10726_), .A2(new_n10725_), .ZN(new_n10727_));
  INV_X1     g10534(.I(new_n10727_), .ZN(new_n10728_));
  OAI22_X1   g10535(.A1(new_n10728_), .A2(new_n10724_), .B1(new_n8076_), .B2(new_n10726_), .ZN(new_n10729_));
  INV_X1     g10536(.I(new_n10729_), .ZN(new_n10730_));
  XOR2_X1    g10537(.A1(new_n10723_), .A2(new_n10730_), .Z(new_n10731_));
  XOR2_X1    g10538(.A1(new_n10705_), .A2(new_n10731_), .Z(new_n10732_));
  XOR2_X1    g10539(.A1(new_n10732_), .A2(new_n10702_), .Z(new_n10733_));
  NOR2_X1    g10540(.A1(new_n10509_), .A2(new_n10506_), .ZN(new_n10734_));
  INV_X1     g10541(.I(new_n10734_), .ZN(new_n10735_));
  OAI21_X1   g10542(.A1(new_n10507_), .A2(new_n10508_), .B(new_n10735_), .ZN(new_n10736_));
  XNOR2_X1   g10543(.A1(new_n10736_), .A2(new_n10733_), .ZN(new_n10737_));
  XNOR2_X1   g10544(.A1(new_n10737_), .A2(new_n10675_), .ZN(new_n10738_));
  XOR2_X1    g10545(.A1(new_n10673_), .A2(new_n10738_), .Z(new_n10739_));
  XNOR2_X1   g10546(.A1(new_n10633_), .A2(new_n10625_), .ZN(new_n10740_));
  XOR2_X1    g10547(.A1(new_n10740_), .A2(new_n10620_), .Z(new_n10741_));
  NAND2_X1   g10548(.A1(new_n10621_), .A2(new_n10628_), .ZN(new_n10742_));
  INV_X1     g10549(.I(new_n10635_), .ZN(new_n10743_));
  OAI21_X1   g10550(.A1(new_n10629_), .A2(new_n10743_), .B(new_n10742_), .ZN(new_n10744_));
  NAND2_X1   g10551(.A1(new_n10599_), .A2(new_n10419_), .ZN(new_n10745_));
  NAND2_X1   g10552(.A1(new_n10600_), .A2(new_n10608_), .ZN(new_n10746_));
  NAND2_X1   g10553(.A1(new_n10746_), .A2(new_n10745_), .ZN(new_n10747_));
  XOR2_X1    g10554(.A1(new_n10744_), .A2(new_n10747_), .Z(new_n10748_));
  XOR2_X1    g10555(.A1(new_n10748_), .A2(new_n10741_), .Z(new_n10749_));
  INV_X1     g10556(.I(new_n10749_), .ZN(new_n10750_));
  NOR2_X1    g10557(.A1(new_n10636_), .A2(new_n10609_), .ZN(new_n10751_));
  INV_X1     g10558(.I(new_n10751_), .ZN(new_n10752_));
  OAI21_X1   g10559(.A1(new_n10637_), .A2(new_n10591_), .B(new_n10752_), .ZN(new_n10753_));
  OAI21_X1   g10560(.A1(new_n10438_), .A2(new_n10568_), .B(new_n10565_), .ZN(new_n10754_));
  XNOR2_X1   g10561(.A1(new_n10754_), .A2(new_n10587_), .ZN(new_n10755_));
  NAND2_X1   g10562(.A1(new_n2437_), .A2(new_n5439_), .ZN(new_n10756_));
  NAND2_X1   g10563(.A1(new_n2201_), .A2(new_n7867_), .ZN(new_n10757_));
  AOI22_X1   g10564(.A1(new_n10756_), .A2(new_n10757_), .B1(new_n3210_), .B2(new_n5154_), .ZN(new_n10758_));
  NAND2_X1   g10565(.A1(\a[30] ), .A2(\a[51] ), .ZN(new_n10759_));
  AOI22_X1   g10566(.A1(\a[31] ), .A2(\a[50] ), .B1(\a[32] ), .B2(\a[49] ), .ZN(new_n10760_));
  NAND2_X1   g10567(.A1(new_n3210_), .A2(new_n5154_), .ZN(new_n10761_));
  NAND3_X1   g10568(.A1(new_n10761_), .A2(new_n10756_), .A3(new_n10757_), .ZN(new_n10762_));
  OAI22_X1   g10569(.A1(new_n10758_), .A2(new_n10759_), .B1(new_n10762_), .B2(new_n10760_), .ZN(new_n10763_));
  XNOR2_X1   g10570(.A1(new_n10755_), .A2(new_n10763_), .ZN(new_n10764_));
  NOR2_X1    g10571(.A1(new_n10596_), .A2(new_n10592_), .ZN(new_n10765_));
  NAND2_X1   g10572(.A1(new_n10606_), .A2(new_n10576_), .ZN(new_n10766_));
  NAND2_X1   g10573(.A1(new_n10607_), .A2(new_n10577_), .ZN(new_n10767_));
  AND2_X2    g10574(.A1(new_n10767_), .A2(new_n10766_), .Z(new_n10768_));
  XNOR2_X1   g10575(.A1(new_n10768_), .A2(new_n10765_), .ZN(new_n10769_));
  NAND2_X1   g10576(.A1(new_n10589_), .A2(new_n10579_), .ZN(new_n10770_));
  OAI21_X1   g10577(.A1(new_n10590_), .A2(new_n10569_), .B(new_n10770_), .ZN(new_n10771_));
  XNOR2_X1   g10578(.A1(new_n10771_), .A2(new_n10769_), .ZN(new_n10772_));
  XNOR2_X1   g10579(.A1(new_n10772_), .A2(new_n10764_), .ZN(new_n10773_));
  XNOR2_X1   g10580(.A1(new_n10773_), .A2(new_n10753_), .ZN(new_n10774_));
  INV_X1     g10581(.I(new_n10774_), .ZN(new_n10775_));
  NOR2_X1    g10582(.A1(new_n10775_), .A2(new_n10750_), .ZN(new_n10776_));
  INV_X1     g10583(.I(new_n10776_), .ZN(new_n10777_));
  NAND2_X1   g10584(.A1(new_n10775_), .A2(new_n10750_), .ZN(new_n10778_));
  AND2_X2    g10585(.A1(new_n10777_), .A2(new_n10778_), .Z(new_n10779_));
  NOR2_X1    g10586(.A1(new_n10645_), .A2(new_n10641_), .ZN(new_n10780_));
  NOR2_X1    g10587(.A1(new_n10427_), .A2(new_n10348_), .ZN(new_n10781_));
  INV_X1     g10588(.I(new_n10538_), .ZN(new_n10782_));
  NOR2_X1    g10589(.A1(new_n10782_), .A2(new_n10358_), .ZN(new_n10783_));
  NOR2_X1    g10590(.A1(new_n10783_), .A2(new_n10781_), .ZN(new_n10784_));
  NOR2_X1    g10591(.A1(new_n1750_), .A2(new_n5617_), .ZN(new_n10785_));
  INV_X1     g10592(.I(new_n10785_), .ZN(new_n10786_));
  AOI22_X1   g10593(.A1(\a[38] ), .A2(\a[43] ), .B1(\a[39] ), .B2(\a[42] ), .ZN(new_n10787_));
  NOR2_X1    g10594(.A1(new_n4181_), .A2(new_n4210_), .ZN(new_n10788_));
  NOR3_X1    g10595(.A1(new_n10788_), .A2(new_n10786_), .A3(new_n10787_), .ZN(new_n10789_));
  NOR2_X1    g10596(.A1(new_n10789_), .A2(new_n10788_), .ZN(new_n10790_));
  INV_X1     g10597(.I(new_n10790_), .ZN(new_n10791_));
  OAI22_X1   g10598(.A1(new_n10791_), .A2(new_n10787_), .B1(new_n10786_), .B2(new_n10789_), .ZN(new_n10792_));
  NAND2_X1   g10599(.A1(new_n10513_), .A2(new_n10465_), .ZN(new_n10793_));
  NAND2_X1   g10600(.A1(new_n10793_), .A2(new_n10512_), .ZN(new_n10794_));
  XNOR2_X1   g10601(.A1(new_n10794_), .A2(new_n10792_), .ZN(new_n10795_));
  XOR2_X1    g10602(.A1(new_n10795_), .A2(new_n10784_), .Z(new_n10796_));
  INV_X1     g10603(.I(new_n10796_), .ZN(new_n10797_));
  NOR2_X1    g10604(.A1(new_n10526_), .A2(new_n10523_), .ZN(new_n10798_));
  NOR2_X1    g10605(.A1(new_n10546_), .A2(new_n10542_), .ZN(new_n10799_));
  XNOR2_X1   g10606(.A1(new_n10799_), .A2(new_n10798_), .ZN(new_n10800_));
  NOR2_X1    g10607(.A1(new_n10800_), .A2(new_n10797_), .ZN(new_n10801_));
  INV_X1     g10608(.I(new_n10801_), .ZN(new_n10802_));
  NAND2_X1   g10609(.A1(new_n10800_), .A2(new_n10797_), .ZN(new_n10803_));
  AND2_X2    g10610(.A1(new_n10802_), .A2(new_n10803_), .Z(new_n10804_));
  XOR2_X1    g10611(.A1(new_n10780_), .A2(new_n10804_), .Z(new_n10805_));
  XOR2_X1    g10612(.A1(new_n10805_), .A2(new_n10779_), .Z(new_n10806_));
  XOR2_X1    g10613(.A1(new_n10806_), .A2(new_n10739_), .Z(new_n10807_));
  NAND2_X1   g10614(.A1(new_n10559_), .A2(new_n10646_), .ZN(new_n10808_));
  NAND2_X1   g10615(.A1(new_n10647_), .A2(new_n10556_), .ZN(new_n10809_));
  NAND2_X1   g10616(.A1(new_n10809_), .A2(new_n10808_), .ZN(new_n10810_));
  NOR2_X1    g10617(.A1(new_n10807_), .A2(new_n10810_), .ZN(new_n10811_));
  NAND2_X1   g10618(.A1(new_n10807_), .A2(new_n10810_), .ZN(new_n10812_));
  INV_X1     g10619(.I(new_n10812_), .ZN(new_n10813_));
  NOR2_X1    g10620(.A1(new_n10813_), .A2(new_n10811_), .ZN(new_n10814_));
  XOR2_X1    g10621(.A1(new_n10670_), .A2(new_n10814_), .Z(\asquared[82] ));
  AOI21_X1   g10622(.A1(new_n10669_), .A2(new_n10649_), .B(new_n10811_), .ZN(new_n10816_));
  NOR2_X1    g10623(.A1(new_n10816_), .A2(new_n10813_), .ZN(new_n10817_));
  INV_X1     g10624(.I(new_n10804_), .ZN(new_n10818_));
  NOR2_X1    g10625(.A1(new_n10780_), .A2(new_n10818_), .ZN(new_n10819_));
  INV_X1     g10626(.I(new_n10805_), .ZN(new_n10820_));
  AOI21_X1   g10627(.A1(new_n10820_), .A2(new_n10779_), .B(new_n10819_), .ZN(new_n10821_));
  INV_X1     g10628(.I(new_n10753_), .ZN(new_n10822_));
  NOR2_X1    g10629(.A1(new_n10822_), .A2(new_n10773_), .ZN(new_n10823_));
  NOR2_X1    g10630(.A1(new_n10776_), .A2(new_n10823_), .ZN(new_n10824_));
  OAI21_X1   g10631(.A1(new_n10798_), .A2(new_n10799_), .B(new_n10802_), .ZN(new_n10825_));
  OAI22_X1   g10632(.A1(new_n1814_), .A2(new_n5425_), .B1(new_n2030_), .B2(new_n5175_), .ZN(new_n10826_));
  NAND2_X1   g10633(.A1(new_n2254_), .A2(new_n5862_), .ZN(new_n10827_));
  NAND3_X1   g10634(.A1(new_n10827_), .A2(new_n5239_), .A3(new_n10826_), .ZN(new_n10828_));
  NAND2_X1   g10635(.A1(new_n10828_), .A2(new_n5239_), .ZN(new_n10829_));
  NAND2_X1   g10636(.A1(new_n10828_), .A2(new_n10827_), .ZN(new_n10830_));
  INV_X1     g10637(.I(new_n10830_), .ZN(new_n10831_));
  NAND2_X1   g10638(.A1(new_n10831_), .A2(new_n10826_), .ZN(new_n10832_));
  NAND2_X1   g10639(.A1(new_n10832_), .A2(new_n10829_), .ZN(new_n10833_));
  AOI22_X1   g10640(.A1(\a[38] ), .A2(\a[44] ), .B1(\a[39] ), .B2(\a[43] ), .ZN(new_n10834_));
  INV_X1     g10641(.I(new_n10834_), .ZN(new_n10835_));
  NOR2_X1    g10642(.A1(new_n4210_), .A2(new_n4343_), .ZN(new_n10836_));
  NOR2_X1    g10643(.A1(new_n1566_), .A2(new_n5856_), .ZN(new_n10837_));
  AOI21_X1   g10644(.A1(new_n10835_), .A2(new_n10837_), .B(new_n10836_), .ZN(new_n10838_));
  INV_X1     g10645(.I(new_n10838_), .ZN(new_n10839_));
  OAI21_X1   g10646(.A1(new_n10836_), .A2(new_n10834_), .B(new_n10837_), .ZN(new_n10840_));
  OAI21_X1   g10647(.A1(new_n10839_), .A2(new_n10834_), .B(new_n10840_), .ZN(new_n10841_));
  XNOR2_X1   g10648(.A1(new_n10833_), .A2(new_n10841_), .ZN(new_n10842_));
  NAND3_X1   g10649(.A1(new_n4844_), .A2(\a[37] ), .A3(\a[47] ), .ZN(new_n10843_));
  NAND2_X1   g10650(.A1(new_n3232_), .A2(new_n4720_), .ZN(new_n10844_));
  AOI22_X1   g10651(.A1(new_n10844_), .A2(new_n10843_), .B1(new_n3037_), .B2(new_n4429_), .ZN(new_n10845_));
  NAND2_X1   g10652(.A1(\a[35] ), .A2(\a[47] ), .ZN(new_n10846_));
  AOI21_X1   g10653(.A1(\a[36] ), .A2(\a[46] ), .B(new_n5093_), .ZN(new_n10847_));
  NAND2_X1   g10654(.A1(new_n3037_), .A2(new_n4429_), .ZN(new_n10848_));
  NAND3_X1   g10655(.A1(new_n10848_), .A2(new_n10844_), .A3(new_n10843_), .ZN(new_n10849_));
  OAI22_X1   g10656(.A1(new_n10845_), .A2(new_n10846_), .B1(new_n10849_), .B2(new_n10847_), .ZN(new_n10850_));
  XOR2_X1    g10657(.A1(new_n10842_), .A2(new_n10850_), .Z(new_n10851_));
  INV_X1     g10658(.I(new_n10851_), .ZN(new_n10852_));
  NAND2_X1   g10659(.A1(new_n10794_), .A2(new_n10792_), .ZN(new_n10853_));
  OAI21_X1   g10660(.A1(new_n10795_), .A2(new_n10784_), .B(new_n10853_), .ZN(new_n10854_));
  NOR4_X1    g10661(.A1(new_n1043_), .A2(new_n2051_), .A3(new_n5135_), .A4(new_n7144_), .ZN(new_n10855_));
  NOR2_X1    g10662(.A1(new_n1382_), .A2(new_n7591_), .ZN(new_n10856_));
  NAND4_X1   g10663(.A1(\a[21] ), .A2(\a[31] ), .A3(\a[51] ), .A4(\a[61] ), .ZN(new_n10857_));
  OAI21_X1   g10664(.A1(new_n10856_), .A2(new_n10855_), .B(new_n10857_), .ZN(new_n10858_));
  NAND3_X1   g10665(.A1(new_n10858_), .A2(\a[20] ), .A3(\a[62] ), .ZN(new_n10859_));
  AOI22_X1   g10666(.A1(\a[21] ), .A2(\a[61] ), .B1(\a[31] ), .B2(\a[51] ), .ZN(new_n10860_));
  NAND2_X1   g10667(.A1(new_n10858_), .A2(new_n10857_), .ZN(new_n10861_));
  OAI21_X1   g10668(.A1(new_n10860_), .A2(new_n10861_), .B(new_n10859_), .ZN(new_n10862_));
  NAND2_X1   g10669(.A1(new_n3577_), .A2(new_n4980_), .ZN(new_n10863_));
  OAI22_X1   g10670(.A1(new_n2637_), .A2(new_n5155_), .B1(new_n3375_), .B2(new_n4903_), .ZN(new_n10864_));
  NAND2_X1   g10671(.A1(new_n10864_), .A2(new_n10863_), .ZN(new_n10865_));
  NAND3_X1   g10672(.A1(new_n10865_), .A2(\a[32] ), .A3(\a[50] ), .ZN(new_n10866_));
  AOI22_X1   g10673(.A1(\a[33] ), .A2(\a[49] ), .B1(\a[34] ), .B2(\a[48] ), .ZN(new_n10867_));
  NAND2_X1   g10674(.A1(new_n10865_), .A2(new_n10863_), .ZN(new_n10868_));
  OAI21_X1   g10675(.A1(new_n10867_), .A2(new_n10868_), .B(new_n10866_), .ZN(new_n10869_));
  XOR2_X1    g10676(.A1(new_n10869_), .A2(new_n10862_), .Z(new_n10870_));
  NAND2_X1   g10677(.A1(new_n1767_), .A2(new_n7451_), .ZN(new_n10871_));
  NAND2_X1   g10678(.A1(new_n1879_), .A2(new_n7800_), .ZN(new_n10872_));
  AOI22_X1   g10679(.A1(new_n10871_), .A2(new_n10872_), .B1(new_n1528_), .B2(new_n7205_), .ZN(new_n10873_));
  NAND2_X1   g10680(.A1(\a[22] ), .A2(\a[60] ), .ZN(new_n10874_));
  AOI22_X1   g10681(.A1(\a[23] ), .A2(\a[59] ), .B1(\a[24] ), .B2(\a[58] ), .ZN(new_n10875_));
  NAND2_X1   g10682(.A1(new_n1528_), .A2(new_n7205_), .ZN(new_n10876_));
  NAND3_X1   g10683(.A1(new_n10876_), .A2(new_n10871_), .A3(new_n10872_), .ZN(new_n10877_));
  OAI22_X1   g10684(.A1(new_n10873_), .A2(new_n10874_), .B1(new_n10877_), .B2(new_n10875_), .ZN(new_n10878_));
  XNOR2_X1   g10685(.A1(new_n10870_), .A2(new_n10878_), .ZN(new_n10879_));
  INV_X1     g10686(.I(new_n10879_), .ZN(new_n10880_));
  XOR2_X1    g10687(.A1(new_n10854_), .A2(new_n10880_), .Z(new_n10881_));
  XOR2_X1    g10688(.A1(new_n10881_), .A2(new_n10852_), .Z(new_n10882_));
  XNOR2_X1   g10689(.A1(new_n10825_), .A2(new_n10882_), .ZN(new_n10883_));
  XNOR2_X1   g10690(.A1(new_n10883_), .A2(new_n10824_), .ZN(new_n10884_));
  XNOR2_X1   g10691(.A1(new_n10821_), .A2(new_n10884_), .ZN(new_n10885_));
  NOR2_X1    g10692(.A1(new_n10710_), .A2(new_n9688_), .ZN(new_n10886_));
  NOR2_X1    g10693(.A1(new_n10709_), .A2(new_n9689_), .ZN(new_n10887_));
  NOR2_X1    g10694(.A1(new_n10886_), .A2(new_n10887_), .ZN(new_n10888_));
  NOR2_X1    g10695(.A1(new_n10791_), .A2(new_n10888_), .ZN(new_n10889_));
  INV_X1     g10696(.I(new_n10888_), .ZN(new_n10890_));
  NOR2_X1    g10697(.A1(new_n10890_), .A2(new_n10790_), .ZN(new_n10891_));
  NOR2_X1    g10698(.A1(new_n10889_), .A2(new_n10891_), .ZN(new_n10892_));
  NAND2_X1   g10699(.A1(new_n10722_), .A2(new_n10711_), .ZN(new_n10893_));
  OAI21_X1   g10700(.A1(new_n10723_), .A2(new_n10730_), .B(new_n10893_), .ZN(new_n10894_));
  NAND2_X1   g10701(.A1(new_n10588_), .A2(new_n10754_), .ZN(new_n10895_));
  NAND2_X1   g10702(.A1(new_n10755_), .A2(new_n10763_), .ZN(new_n10896_));
  NAND2_X1   g10703(.A1(new_n10896_), .A2(new_n10895_), .ZN(new_n10897_));
  NOR2_X1    g10704(.A1(new_n10894_), .A2(new_n10897_), .ZN(new_n10898_));
  NAND2_X1   g10705(.A1(new_n10894_), .A2(new_n10897_), .ZN(new_n10899_));
  INV_X1     g10706(.I(new_n10899_), .ZN(new_n10900_));
  NOR2_X1    g10707(.A1(new_n10900_), .A2(new_n10898_), .ZN(new_n10901_));
  NAND2_X1   g10708(.A1(new_n10901_), .A2(new_n10892_), .ZN(new_n10902_));
  INV_X1     g10709(.I(new_n10902_), .ZN(new_n10903_));
  NOR2_X1    g10710(.A1(new_n10901_), .A2(new_n10892_), .ZN(new_n10904_));
  NOR2_X1    g10711(.A1(new_n10903_), .A2(new_n10904_), .ZN(new_n10905_));
  INV_X1     g10712(.I(new_n10905_), .ZN(new_n10906_));
  NAND2_X1   g10713(.A1(new_n10705_), .A2(new_n10731_), .ZN(new_n10907_));
  NAND2_X1   g10714(.A1(new_n10732_), .A2(new_n10702_), .ZN(new_n10908_));
  NAND2_X1   g10715(.A1(new_n10908_), .A2(new_n10907_), .ZN(new_n10909_));
  XNOR2_X1   g10716(.A1(new_n10727_), .A2(new_n10762_), .ZN(new_n10910_));
  XOR2_X1    g10717(.A1(new_n10910_), .A2(new_n10696_), .Z(new_n10911_));
  NAND2_X1   g10718(.A1(new_n10682_), .A2(new_n10690_), .ZN(new_n10912_));
  OAI21_X1   g10719(.A1(new_n10691_), .A2(new_n10700_), .B(new_n10912_), .ZN(new_n10913_));
  XOR2_X1    g10720(.A1(new_n10721_), .A2(new_n10681_), .Z(new_n10914_));
  XOR2_X1    g10721(.A1(new_n10914_), .A2(new_n10689_), .Z(new_n10915_));
  XOR2_X1    g10722(.A1(new_n10915_), .A2(new_n10913_), .Z(new_n10916_));
  XNOR2_X1   g10723(.A1(new_n10916_), .A2(new_n10911_), .ZN(new_n10917_));
  XOR2_X1    g10724(.A1(new_n10909_), .A2(new_n10917_), .Z(new_n10918_));
  XOR2_X1    g10725(.A1(new_n10918_), .A2(new_n10906_), .Z(new_n10919_));
  NOR2_X1    g10726(.A1(new_n10737_), .A2(new_n10675_), .ZN(new_n10920_));
  AOI21_X1   g10727(.A1(new_n10733_), .A2(new_n10736_), .B(new_n10920_), .ZN(new_n10921_));
  NAND2_X1   g10728(.A1(new_n10634_), .A2(new_n10625_), .ZN(new_n10922_));
  NAND2_X1   g10729(.A1(new_n10740_), .A2(new_n10620_), .ZN(new_n10923_));
  NAND2_X1   g10730(.A1(new_n10923_), .A2(new_n10922_), .ZN(new_n10924_));
  INV_X1     g10731(.I(new_n10768_), .ZN(new_n10925_));
  OAI21_X1   g10732(.A1(new_n10925_), .A2(new_n10765_), .B(new_n10767_), .ZN(new_n10926_));
  NAND3_X1   g10733(.A1(new_n5757_), .A2(\a[25] ), .A3(\a[57] ), .ZN(new_n10927_));
  NAND2_X1   g10734(.A1(new_n2103_), .A2(new_n6128_), .ZN(new_n10928_));
  AOI22_X1   g10735(.A1(new_n10928_), .A2(new_n10927_), .B1(new_n2246_), .B2(new_n8951_), .ZN(new_n10929_));
  AOI22_X1   g10736(.A1(\a[25] ), .A2(\a[57] ), .B1(\a[27] ), .B2(\a[55] ), .ZN(new_n10930_));
  NAND2_X1   g10737(.A1(new_n2246_), .A2(new_n8951_), .ZN(new_n10931_));
  NAND3_X1   g10738(.A1(new_n10931_), .A2(new_n10928_), .A3(new_n10927_), .ZN(new_n10932_));
  OAI22_X1   g10739(.A1(new_n10929_), .A2(new_n5758_), .B1(new_n10932_), .B2(new_n10930_), .ZN(new_n10933_));
  XNOR2_X1   g10740(.A1(new_n10926_), .A2(new_n10933_), .ZN(new_n10934_));
  XNOR2_X1   g10741(.A1(new_n10934_), .A2(new_n10924_), .ZN(new_n10935_));
  NAND2_X1   g10742(.A1(new_n10744_), .A2(new_n10747_), .ZN(new_n10936_));
  NAND2_X1   g10743(.A1(new_n10748_), .A2(new_n10741_), .ZN(new_n10937_));
  NAND2_X1   g10744(.A1(new_n10937_), .A2(new_n10936_), .ZN(new_n10938_));
  NAND2_X1   g10745(.A1(new_n10771_), .A2(new_n10769_), .ZN(new_n10939_));
  OAI21_X1   g10746(.A1(new_n10772_), .A2(new_n10764_), .B(new_n10939_), .ZN(new_n10940_));
  XOR2_X1    g10747(.A1(new_n10938_), .A2(new_n10940_), .Z(new_n10941_));
  XOR2_X1    g10748(.A1(new_n10941_), .A2(new_n10935_), .Z(new_n10942_));
  XOR2_X1    g10749(.A1(new_n10921_), .A2(new_n10942_), .Z(new_n10943_));
  XOR2_X1    g10750(.A1(new_n10943_), .A2(new_n10919_), .Z(new_n10944_));
  XNOR2_X1   g10751(.A1(new_n10885_), .A2(new_n10944_), .ZN(new_n10945_));
  INV_X1     g10752(.I(new_n10945_), .ZN(new_n10946_));
  INV_X1     g10753(.I(new_n10738_), .ZN(new_n10947_));
  NAND2_X1   g10754(.A1(new_n10673_), .A2(new_n10947_), .ZN(new_n10948_));
  OAI21_X1   g10755(.A1(new_n10806_), .A2(new_n10739_), .B(new_n10948_), .ZN(new_n10949_));
  NOR2_X1    g10756(.A1(new_n10946_), .A2(new_n10949_), .ZN(new_n10950_));
  INV_X1     g10757(.I(new_n10950_), .ZN(new_n10951_));
  NAND2_X1   g10758(.A1(new_n10946_), .A2(new_n10949_), .ZN(new_n10952_));
  NAND2_X1   g10759(.A1(new_n10951_), .A2(new_n10952_), .ZN(new_n10953_));
  XOR2_X1    g10760(.A1(new_n10817_), .A2(new_n10953_), .Z(\asquared[83] ));
  OAI21_X1   g10761(.A1(new_n10816_), .A2(new_n10813_), .B(new_n10951_), .ZN(new_n10955_));
  NAND2_X1   g10762(.A1(new_n10955_), .A2(new_n10952_), .ZN(new_n10956_));
  NOR2_X1    g10763(.A1(new_n10821_), .A2(new_n10884_), .ZN(new_n10957_));
  NOR2_X1    g10764(.A1(new_n10885_), .A2(new_n10944_), .ZN(new_n10958_));
  NOR2_X1    g10765(.A1(new_n10958_), .A2(new_n10957_), .ZN(new_n10959_));
  INV_X1     g10766(.I(new_n10959_), .ZN(new_n10960_));
  INV_X1     g10767(.I(new_n10942_), .ZN(new_n10961_));
  NOR2_X1    g10768(.A1(new_n10921_), .A2(new_n10961_), .ZN(new_n10962_));
  INV_X1     g10769(.I(new_n10943_), .ZN(new_n10963_));
  AOI21_X1   g10770(.A1(new_n10963_), .A2(new_n10919_), .B(new_n10962_), .ZN(new_n10964_));
  AOI21_X1   g10771(.A1(new_n10908_), .A2(new_n10907_), .B(new_n10917_), .ZN(new_n10965_));
  NOR2_X1    g10772(.A1(new_n10918_), .A2(new_n10906_), .ZN(new_n10966_));
  NOR2_X1    g10773(.A1(new_n10966_), .A2(new_n10965_), .ZN(new_n10967_));
  NAND2_X1   g10774(.A1(new_n10938_), .A2(new_n10940_), .ZN(new_n10968_));
  NAND2_X1   g10775(.A1(new_n10941_), .A2(new_n10935_), .ZN(new_n10969_));
  NAND2_X1   g10776(.A1(new_n10969_), .A2(new_n10968_), .ZN(new_n10970_));
  NOR2_X1    g10777(.A1(new_n5135_), .A2(new_n6298_), .ZN(new_n10971_));
  NAND2_X1   g10778(.A1(new_n2782_), .A2(new_n10971_), .ZN(new_n10972_));
  NOR4_X1    g10779(.A1(new_n1441_), .A2(new_n2200_), .A3(new_n5135_), .A4(new_n6316_), .ZN(new_n10973_));
  NOR2_X1    g10780(.A1(new_n2177_), .A2(new_n6804_), .ZN(new_n10974_));
  OAI21_X1   g10781(.A1(new_n10974_), .A2(new_n10973_), .B(new_n10972_), .ZN(new_n10975_));
  NAND3_X1   g10782(.A1(new_n10975_), .A2(\a[25] ), .A3(\a[58] ), .ZN(new_n10976_));
  AOI22_X1   g10783(.A1(\a[26] ), .A2(\a[57] ), .B1(\a[32] ), .B2(\a[51] ), .ZN(new_n10977_));
  NAND2_X1   g10784(.A1(new_n10975_), .A2(new_n10972_), .ZN(new_n10978_));
  OAI21_X1   g10785(.A1(new_n10977_), .A2(new_n10978_), .B(new_n10976_), .ZN(new_n10979_));
  NAND2_X1   g10786(.A1(new_n3803_), .A2(new_n4429_), .ZN(new_n10980_));
  OAI22_X1   g10787(.A1(new_n2916_), .A2(new_n4314_), .B1(new_n3038_), .B2(new_n4721_), .ZN(new_n10981_));
  NAND2_X1   g10788(.A1(new_n10981_), .A2(new_n10980_), .ZN(new_n10982_));
  NAND3_X1   g10789(.A1(new_n10982_), .A2(\a[36] ), .A3(\a[47] ), .ZN(new_n10983_));
  AOI22_X1   g10790(.A1(\a[37] ), .A2(\a[46] ), .B1(\a[38] ), .B2(\a[45] ), .ZN(new_n10984_));
  NAND2_X1   g10791(.A1(new_n10982_), .A2(new_n10980_), .ZN(new_n10985_));
  OAI21_X1   g10792(.A1(new_n10984_), .A2(new_n10985_), .B(new_n10983_), .ZN(new_n10986_));
  XOR2_X1    g10793(.A1(new_n10986_), .A2(new_n10979_), .Z(new_n10987_));
  INV_X1     g10794(.I(new_n10354_), .ZN(new_n10988_));
  AOI22_X1   g10795(.A1(\a[20] ), .A2(\a[63] ), .B1(\a[22] ), .B2(\a[61] ), .ZN(new_n10989_));
  NOR2_X1    g10796(.A1(new_n2647_), .A2(new_n7959_), .ZN(new_n10990_));
  NOR3_X1    g10797(.A1(new_n10990_), .A2(new_n10988_), .A3(new_n10989_), .ZN(new_n10991_));
  NOR2_X1    g10798(.A1(new_n10991_), .A2(new_n10990_), .ZN(new_n10992_));
  INV_X1     g10799(.I(new_n10992_), .ZN(new_n10993_));
  OAI22_X1   g10800(.A1(new_n10993_), .A2(new_n10989_), .B1(new_n10988_), .B2(new_n10991_), .ZN(new_n10994_));
  XNOR2_X1   g10801(.A1(new_n10987_), .A2(new_n10994_), .ZN(new_n10995_));
  INV_X1     g10802(.I(new_n10995_), .ZN(new_n10996_));
  NAND2_X1   g10803(.A1(new_n10926_), .A2(new_n10933_), .ZN(new_n10997_));
  INV_X1     g10804(.I(new_n10934_), .ZN(new_n10998_));
  NAND2_X1   g10805(.A1(new_n10998_), .A2(new_n10924_), .ZN(new_n10999_));
  NAND2_X1   g10806(.A1(new_n10999_), .A2(new_n10997_), .ZN(new_n11000_));
  NAND4_X1   g10807(.A1(\a[21] ), .A2(\a[41] ), .A3(\a[42] ), .A4(\a[62] ), .ZN(new_n11001_));
  AOI21_X1   g10808(.A1(\a[21] ), .A2(\a[62] ), .B(\a[42] ), .ZN(new_n11002_));
  NAND3_X1   g10809(.A1(\a[21] ), .A2(\a[42] ), .A3(\a[62] ), .ZN(new_n11003_));
  NAND2_X1   g10810(.A1(new_n4667_), .A2(new_n11003_), .ZN(new_n11004_));
  OAI21_X1   g10811(.A1(new_n11004_), .A2(new_n11002_), .B(new_n11001_), .ZN(new_n11005_));
  AOI22_X1   g10812(.A1(\a[39] ), .A2(\a[44] ), .B1(\a[40] ), .B2(\a[43] ), .ZN(new_n11006_));
  NOR2_X1    g10813(.A1(new_n1814_), .A2(new_n5617_), .ZN(new_n11007_));
  INV_X1     g10814(.I(new_n11007_), .ZN(new_n11008_));
  OAI22_X1   g10815(.A1(new_n3551_), .A2(new_n4343_), .B1(new_n11008_), .B2(new_n11006_), .ZN(new_n11009_));
  NOR2_X1    g10816(.A1(new_n3551_), .A2(new_n4343_), .ZN(new_n11010_));
  OAI21_X1   g10817(.A1(new_n11010_), .A2(new_n11006_), .B(new_n11007_), .ZN(new_n11011_));
  OAI21_X1   g10818(.A1(new_n11009_), .A2(new_n11006_), .B(new_n11011_), .ZN(new_n11012_));
  XOR2_X1    g10819(.A1(new_n11012_), .A2(new_n11005_), .Z(new_n11013_));
  AOI22_X1   g10820(.A1(new_n2525_), .A2(new_n4902_), .B1(new_n3577_), .B2(new_n5154_), .ZN(new_n11014_));
  AOI21_X1   g10821(.A1(new_n2745_), .A2(new_n4980_), .B(new_n11014_), .ZN(new_n11015_));
  NAND2_X1   g10822(.A1(\a[33] ), .A2(\a[50] ), .ZN(new_n11016_));
  AOI22_X1   g10823(.A1(\a[34] ), .A2(\a[49] ), .B1(\a[35] ), .B2(\a[48] ), .ZN(new_n11017_));
  OAI21_X1   g10824(.A1(new_n2746_), .A2(new_n4981_), .B(new_n11014_), .ZN(new_n11018_));
  OAI22_X1   g10825(.A1(new_n11015_), .A2(new_n11016_), .B1(new_n11018_), .B2(new_n11017_), .ZN(new_n11019_));
  XNOR2_X1   g10826(.A1(new_n11013_), .A2(new_n11019_), .ZN(new_n11020_));
  INV_X1     g10827(.I(new_n11020_), .ZN(new_n11021_));
  XOR2_X1    g10828(.A1(new_n11000_), .A2(new_n11021_), .Z(new_n11022_));
  XOR2_X1    g10829(.A1(new_n11022_), .A2(new_n10996_), .Z(new_n11023_));
  XOR2_X1    g10830(.A1(new_n10970_), .A2(new_n11023_), .Z(new_n11024_));
  XNOR2_X1   g10831(.A1(new_n11024_), .A2(new_n10967_), .ZN(new_n11025_));
  INV_X1     g10832(.I(new_n11025_), .ZN(new_n11026_));
  NAND2_X1   g10833(.A1(new_n10964_), .A2(new_n11026_), .ZN(new_n11027_));
  NOR2_X1    g10834(.A1(new_n10964_), .A2(new_n11026_), .ZN(new_n11028_));
  INV_X1     g10835(.I(new_n11028_), .ZN(new_n11029_));
  AND2_X2    g10836(.A1(new_n11029_), .A2(new_n11027_), .Z(new_n11030_));
  NAND2_X1   g10837(.A1(new_n10915_), .A2(new_n10913_), .ZN(new_n11031_));
  NAND2_X1   g10838(.A1(new_n10916_), .A2(new_n10911_), .ZN(new_n11032_));
  NAND2_X1   g10839(.A1(new_n11032_), .A2(new_n11031_), .ZN(new_n11033_));
  NAND2_X1   g10840(.A1(new_n10854_), .A2(new_n10880_), .ZN(new_n11034_));
  NAND2_X1   g10841(.A1(new_n10881_), .A2(new_n10852_), .ZN(new_n11035_));
  NAND2_X1   g10842(.A1(new_n11035_), .A2(new_n11034_), .ZN(new_n11036_));
  XOR2_X1    g10843(.A1(new_n11036_), .A2(new_n11033_), .Z(new_n11037_));
  XOR2_X1    g10844(.A1(new_n10877_), .A2(new_n10849_), .Z(new_n11038_));
  XOR2_X1    g10845(.A1(new_n11038_), .A2(new_n10839_), .Z(new_n11039_));
  XOR2_X1    g10846(.A1(new_n10868_), .A2(new_n10861_), .Z(new_n11040_));
  XOR2_X1    g10847(.A1(new_n11040_), .A2(new_n10932_), .Z(new_n11041_));
  NAND2_X1   g10848(.A1(new_n10833_), .A2(new_n10841_), .ZN(new_n11042_));
  INV_X1     g10849(.I(new_n10842_), .ZN(new_n11043_));
  NAND2_X1   g10850(.A1(new_n11043_), .A2(new_n10850_), .ZN(new_n11044_));
  NAND2_X1   g10851(.A1(new_n11044_), .A2(new_n11042_), .ZN(new_n11045_));
  XOR2_X1    g10852(.A1(new_n11045_), .A2(new_n11041_), .Z(new_n11046_));
  XOR2_X1    g10853(.A1(new_n11046_), .A2(new_n11039_), .Z(new_n11047_));
  XNOR2_X1   g10854(.A1(new_n11037_), .A2(new_n11047_), .ZN(new_n11048_));
  NAND2_X1   g10855(.A1(new_n10825_), .A2(new_n10882_), .ZN(new_n11049_));
  OAI21_X1   g10856(.A1(new_n10883_), .A2(new_n10824_), .B(new_n11049_), .ZN(new_n11050_));
  NAND2_X1   g10857(.A1(new_n10869_), .A2(new_n10862_), .ZN(new_n11051_));
  NAND2_X1   g10858(.A1(new_n10870_), .A2(new_n10878_), .ZN(new_n11052_));
  NAND2_X1   g10859(.A1(new_n11052_), .A2(new_n11051_), .ZN(new_n11053_));
  NAND2_X1   g10860(.A1(new_n10728_), .A2(new_n10762_), .ZN(new_n11054_));
  NAND2_X1   g10861(.A1(new_n10910_), .A2(new_n10696_), .ZN(new_n11055_));
  NAND2_X1   g10862(.A1(new_n11055_), .A2(new_n11054_), .ZN(new_n11056_));
  NAND2_X1   g10863(.A1(new_n10721_), .A2(new_n10681_), .ZN(new_n11057_));
  NAND2_X1   g10864(.A1(new_n10914_), .A2(new_n10689_), .ZN(new_n11058_));
  NAND2_X1   g10865(.A1(new_n11058_), .A2(new_n11057_), .ZN(new_n11059_));
  XOR2_X1    g10866(.A1(new_n11059_), .A2(new_n11056_), .Z(new_n11060_));
  XOR2_X1    g10867(.A1(new_n11060_), .A2(new_n11053_), .Z(new_n11061_));
  NOR2_X1    g10868(.A1(new_n10903_), .A2(new_n10900_), .ZN(new_n11062_));
  NOR2_X1    g10869(.A1(new_n10891_), .A2(new_n10887_), .ZN(new_n11063_));
  NAND4_X1   g10870(.A1(\a[28] ), .A2(\a[31] ), .A3(\a[52] ), .A4(\a[55] ), .ZN(new_n11064_));
  NAND2_X1   g10871(.A1(new_n2437_), .A2(new_n5862_), .ZN(new_n11065_));
  AOI22_X1   g10872(.A1(new_n11065_), .A2(new_n11064_), .B1(new_n2681_), .B2(new_n6124_), .ZN(new_n11066_));
  NAND2_X1   g10873(.A1(\a[31] ), .A2(\a[52] ), .ZN(new_n11067_));
  AOI22_X1   g10874(.A1(\a[28] ), .A2(\a[55] ), .B1(\a[30] ), .B2(\a[53] ), .ZN(new_n11068_));
  NAND2_X1   g10875(.A1(new_n2681_), .A2(new_n6124_), .ZN(new_n11069_));
  NAND3_X1   g10876(.A1(new_n11069_), .A2(new_n11065_), .A3(new_n11064_), .ZN(new_n11070_));
  OAI22_X1   g10877(.A1(new_n11066_), .A2(new_n11067_), .B1(new_n11070_), .B2(new_n11068_), .ZN(new_n11071_));
  NOR2_X1    g10878(.A1(new_n1529_), .A2(new_n7452_), .ZN(new_n11072_));
  INV_X1     g10879(.I(new_n11072_), .ZN(new_n11073_));
  NOR2_X1    g10880(.A1(new_n1357_), .A2(new_n6548_), .ZN(new_n11074_));
  NOR2_X1    g10881(.A1(new_n1299_), .A2(new_n6723_), .ZN(new_n11075_));
  OAI21_X1   g10882(.A1(new_n11074_), .A2(new_n11075_), .B(new_n11073_), .ZN(new_n11076_));
  XOR2_X1    g10883(.A1(new_n11076_), .A2(new_n10830_), .Z(new_n11077_));
  XOR2_X1    g10884(.A1(new_n11077_), .A2(new_n11071_), .Z(new_n11078_));
  XOR2_X1    g10885(.A1(new_n11078_), .A2(new_n11063_), .Z(new_n11079_));
  INV_X1     g10886(.I(new_n11079_), .ZN(new_n11080_));
  XOR2_X1    g10887(.A1(new_n11062_), .A2(new_n11080_), .Z(new_n11081_));
  NAND2_X1   g10888(.A1(new_n11081_), .A2(new_n11061_), .ZN(new_n11082_));
  INV_X1     g10889(.I(new_n11082_), .ZN(new_n11083_));
  NOR2_X1    g10890(.A1(new_n11081_), .A2(new_n11061_), .ZN(new_n11084_));
  NOR2_X1    g10891(.A1(new_n11083_), .A2(new_n11084_), .ZN(new_n11085_));
  XOR2_X1    g10892(.A1(new_n11050_), .A2(new_n11085_), .Z(new_n11086_));
  XOR2_X1    g10893(.A1(new_n11086_), .A2(new_n11048_), .Z(new_n11087_));
  XOR2_X1    g10894(.A1(new_n11030_), .A2(new_n11087_), .Z(new_n11088_));
  INV_X1     g10895(.I(new_n11088_), .ZN(new_n11089_));
  NOR2_X1    g10896(.A1(new_n10960_), .A2(new_n11089_), .ZN(new_n11090_));
  NOR2_X1    g10897(.A1(new_n10959_), .A2(new_n11088_), .ZN(new_n11091_));
  NOR2_X1    g10898(.A1(new_n11090_), .A2(new_n11091_), .ZN(new_n11092_));
  XOR2_X1    g10899(.A1(new_n10956_), .A2(new_n11092_), .Z(\asquared[84] ));
  AOI21_X1   g10900(.A1(new_n10955_), .A2(new_n10952_), .B(new_n11090_), .ZN(new_n11094_));
  NOR2_X1    g10901(.A1(new_n11094_), .A2(new_n11091_), .ZN(new_n11095_));
  INV_X1     g10902(.I(new_n11030_), .ZN(new_n11096_));
  OAI21_X1   g10903(.A1(new_n11096_), .A2(new_n11087_), .B(new_n11029_), .ZN(new_n11097_));
  NAND2_X1   g10904(.A1(new_n11000_), .A2(new_n11021_), .ZN(new_n11098_));
  NAND2_X1   g10905(.A1(new_n11022_), .A2(new_n10996_), .ZN(new_n11099_));
  NAND2_X1   g10906(.A1(new_n11099_), .A2(new_n11098_), .ZN(new_n11100_));
  NAND2_X1   g10907(.A1(new_n11045_), .A2(new_n11041_), .ZN(new_n11101_));
  NAND2_X1   g10908(.A1(new_n11046_), .A2(new_n11039_), .ZN(new_n11102_));
  NAND2_X1   g10909(.A1(new_n11102_), .A2(new_n11101_), .ZN(new_n11103_));
  XOR2_X1    g10910(.A1(new_n11100_), .A2(new_n11103_), .Z(new_n11104_));
  XOR2_X1    g10911(.A1(new_n11009_), .A2(new_n11004_), .Z(new_n11105_));
  XOR2_X1    g10912(.A1(new_n11105_), .A2(new_n11070_), .Z(new_n11106_));
  NAND2_X1   g10913(.A1(new_n10986_), .A2(new_n10979_), .ZN(new_n11107_));
  NAND2_X1   g10914(.A1(new_n10987_), .A2(new_n10994_), .ZN(new_n11108_));
  NAND2_X1   g10915(.A1(new_n11108_), .A2(new_n11107_), .ZN(new_n11109_));
  NAND2_X1   g10916(.A1(new_n11012_), .A2(new_n11005_), .ZN(new_n11110_));
  NAND2_X1   g10917(.A1(new_n11013_), .A2(new_n11019_), .ZN(new_n11111_));
  NAND2_X1   g10918(.A1(new_n11111_), .A2(new_n11110_), .ZN(new_n11112_));
  XOR2_X1    g10919(.A1(new_n11109_), .A2(new_n11112_), .Z(new_n11113_));
  XOR2_X1    g10920(.A1(new_n11113_), .A2(new_n11106_), .Z(new_n11114_));
  XNOR2_X1   g10921(.A1(new_n11104_), .A2(new_n11114_), .ZN(new_n11115_));
  NAND2_X1   g10922(.A1(new_n10970_), .A2(new_n11023_), .ZN(new_n11116_));
  INV_X1     g10923(.I(new_n11024_), .ZN(new_n11117_));
  OAI21_X1   g10924(.A1(new_n11117_), .A2(new_n10967_), .B(new_n11116_), .ZN(new_n11118_));
  NAND2_X1   g10925(.A1(new_n11036_), .A2(new_n11033_), .ZN(new_n11119_));
  NAND2_X1   g10926(.A1(new_n11037_), .A2(new_n11047_), .ZN(new_n11120_));
  NAND2_X1   g10927(.A1(new_n11120_), .A2(new_n11119_), .ZN(new_n11121_));
  XOR2_X1    g10928(.A1(new_n11118_), .A2(new_n11121_), .Z(new_n11122_));
  INV_X1     g10929(.I(new_n11122_), .ZN(new_n11123_));
  OR2_X2     g10930(.A1(new_n11123_), .A2(new_n11115_), .Z(new_n11124_));
  NAND2_X1   g10931(.A1(new_n11123_), .A2(new_n11115_), .ZN(new_n11125_));
  AND2_X2    g10932(.A1(new_n11124_), .A2(new_n11125_), .Z(new_n11126_));
  NAND2_X1   g10933(.A1(new_n11050_), .A2(new_n11085_), .ZN(new_n11127_));
  INV_X1     g10934(.I(new_n11086_), .ZN(new_n11128_));
  OAI21_X1   g10935(.A1(new_n11128_), .A2(new_n11048_), .B(new_n11127_), .ZN(new_n11129_));
  XOR2_X1    g10936(.A1(new_n10985_), .A2(new_n11018_), .Z(new_n11130_));
  XOR2_X1    g10937(.A1(new_n11130_), .A2(new_n10978_), .Z(new_n11131_));
  NAND2_X1   g10938(.A1(new_n10868_), .A2(new_n10861_), .ZN(new_n11132_));
  NAND2_X1   g10939(.A1(new_n11040_), .A2(new_n10932_), .ZN(new_n11133_));
  NAND2_X1   g10940(.A1(new_n11133_), .A2(new_n11132_), .ZN(new_n11134_));
  NAND2_X1   g10941(.A1(new_n10877_), .A2(new_n10849_), .ZN(new_n11135_));
  NAND2_X1   g10942(.A1(new_n11038_), .A2(new_n10839_), .ZN(new_n11136_));
  NAND2_X1   g10943(.A1(new_n11136_), .A2(new_n11135_), .ZN(new_n11137_));
  XOR2_X1    g10944(.A1(new_n11134_), .A2(new_n11137_), .Z(new_n11138_));
  XOR2_X1    g10945(.A1(new_n11138_), .A2(new_n11131_), .Z(new_n11139_));
  NOR2_X1    g10946(.A1(new_n2914_), .A2(new_n5856_), .ZN(new_n11140_));
  INV_X1     g10947(.I(new_n11140_), .ZN(new_n11141_));
  NOR3_X1    g10948(.A1(new_n11141_), .A2(new_n1718_), .A3(new_n4178_), .ZN(new_n11142_));
  NOR2_X1    g10949(.A1(new_n2679_), .A2(new_n7185_), .ZN(new_n11143_));
  NAND4_X1   g10950(.A1(\a[29] ), .A2(\a[38] ), .A3(\a[46] ), .A4(\a[55] ), .ZN(new_n11144_));
  OAI21_X1   g10951(.A1(new_n11142_), .A2(new_n11143_), .B(new_n11144_), .ZN(new_n11145_));
  NAND3_X1   g10952(.A1(new_n11145_), .A2(\a[28] ), .A3(\a[56] ), .ZN(new_n11146_));
  AOI22_X1   g10953(.A1(\a[29] ), .A2(\a[55] ), .B1(\a[38] ), .B2(\a[46] ), .ZN(new_n11147_));
  NAND2_X1   g10954(.A1(new_n11145_), .A2(new_n11144_), .ZN(new_n11148_));
  OAI21_X1   g10955(.A1(new_n11147_), .A2(new_n11148_), .B(new_n11146_), .ZN(new_n11149_));
  NAND2_X1   g10956(.A1(new_n4342_), .A2(new_n4534_), .ZN(new_n11150_));
  OAI22_X1   g10957(.A1(new_n3329_), .A2(new_n4034_), .B1(new_n3551_), .B2(new_n4704_), .ZN(new_n11151_));
  NAND2_X1   g10958(.A1(new_n11151_), .A2(new_n11150_), .ZN(new_n11152_));
  NAND3_X1   g10959(.A1(new_n11152_), .A2(\a[39] ), .A3(\a[45] ), .ZN(new_n11153_));
  AOI21_X1   g10960(.A1(\a[40] ), .A2(\a[44] ), .B(new_n4028_), .ZN(new_n11154_));
  NAND2_X1   g10961(.A1(new_n11152_), .A2(new_n11150_), .ZN(new_n11155_));
  OAI21_X1   g10962(.A1(new_n11154_), .A2(new_n11155_), .B(new_n11153_), .ZN(new_n11156_));
  XNOR2_X1   g10963(.A1(new_n11156_), .A2(new_n11149_), .ZN(new_n11157_));
  NAND2_X1   g10964(.A1(\a[37] ), .A2(\a[47] ), .ZN(new_n11158_));
  AOI22_X1   g10965(.A1(\a[27] ), .A2(\a[57] ), .B1(\a[30] ), .B2(\a[54] ), .ZN(new_n11159_));
  NOR2_X1    g10966(.A1(new_n2030_), .A2(new_n6298_), .ZN(new_n11160_));
  NAND2_X1   g10967(.A1(new_n10785_), .A2(new_n11160_), .ZN(new_n11161_));
  INV_X1     g10968(.I(new_n11161_), .ZN(new_n11162_));
  NOR3_X1    g10969(.A1(new_n11162_), .A2(new_n11158_), .A3(new_n11159_), .ZN(new_n11163_));
  OAI21_X1   g10970(.A1(new_n11158_), .A2(new_n11159_), .B(new_n11161_), .ZN(new_n11164_));
  OAI22_X1   g10971(.A1(new_n11163_), .A2(new_n11158_), .B1(new_n11159_), .B2(new_n11164_), .ZN(new_n11165_));
  XOR2_X1    g10972(.A1(new_n11157_), .A2(new_n11165_), .Z(new_n11166_));
  NOR2_X1    g10973(.A1(new_n2385_), .A2(new_n7591_), .ZN(new_n11167_));
  NOR2_X1    g10974(.A1(new_n1456_), .A2(new_n8049_), .ZN(new_n11168_));
  NOR2_X1    g10975(.A1(new_n1301_), .A2(new_n7959_), .ZN(new_n11169_));
  NOR2_X1    g10976(.A1(new_n11168_), .A2(new_n11169_), .ZN(new_n11170_));
  NOR2_X1    g10977(.A1(new_n11170_), .A2(new_n11167_), .ZN(new_n11171_));
  NAND2_X1   g10978(.A1(\a[21] ), .A2(\a[63] ), .ZN(new_n11172_));
  AOI22_X1   g10979(.A1(\a[22] ), .A2(\a[62] ), .B1(\a[23] ), .B2(\a[61] ), .ZN(new_n11173_));
  NOR2_X1    g10980(.A1(new_n11171_), .A2(new_n11167_), .ZN(new_n11174_));
  INV_X1     g10981(.I(new_n11174_), .ZN(new_n11175_));
  OAI22_X1   g10982(.A1(new_n11175_), .A2(new_n11173_), .B1(new_n11171_), .B2(new_n11172_), .ZN(new_n11176_));
  AOI22_X1   g10983(.A1(\a[24] ), .A2(\a[60] ), .B1(\a[25] ), .B2(\a[59] ), .ZN(new_n11177_));
  INV_X1     g10984(.I(new_n11177_), .ZN(new_n11178_));
  NOR2_X1    g10985(.A1(new_n1779_), .A2(new_n7452_), .ZN(new_n11179_));
  NOR2_X1    g10986(.A1(new_n2274_), .A2(new_n5135_), .ZN(new_n11180_));
  AOI21_X1   g10987(.A1(new_n11178_), .A2(new_n11180_), .B(new_n11179_), .ZN(new_n11181_));
  INV_X1     g10988(.I(new_n11181_), .ZN(new_n11182_));
  OAI21_X1   g10989(.A1(new_n11179_), .A2(new_n11177_), .B(new_n11180_), .ZN(new_n11183_));
  OAI21_X1   g10990(.A1(new_n11182_), .A2(new_n11177_), .B(new_n11183_), .ZN(new_n11184_));
  XNOR2_X1   g10991(.A1(new_n11176_), .A2(new_n11184_), .ZN(new_n11185_));
  NOR2_X1    g10992(.A1(new_n3405_), .A2(new_n4981_), .ZN(new_n11186_));
  AOI22_X1   g10993(.A1(new_n2745_), .A2(new_n5154_), .B1(new_n3822_), .B2(new_n4902_), .ZN(new_n11187_));
  NOR2_X1    g10994(.A1(new_n11186_), .A2(new_n11187_), .ZN(new_n11188_));
  NAND2_X1   g10995(.A1(\a[34] ), .A2(\a[50] ), .ZN(new_n11189_));
  AOI22_X1   g10996(.A1(\a[35] ), .A2(\a[49] ), .B1(\a[36] ), .B2(\a[48] ), .ZN(new_n11190_));
  NOR2_X1    g10997(.A1(new_n11188_), .A2(new_n11186_), .ZN(new_n11191_));
  INV_X1     g10998(.I(new_n11191_), .ZN(new_n11192_));
  OAI22_X1   g10999(.A1(new_n11192_), .A2(new_n11190_), .B1(new_n11188_), .B2(new_n11189_), .ZN(new_n11193_));
  XOR2_X1    g11000(.A1(new_n11185_), .A2(new_n11193_), .Z(new_n11194_));
  XNOR2_X1   g11001(.A1(new_n11194_), .A2(new_n11166_), .ZN(new_n11195_));
  XOR2_X1    g11002(.A1(new_n11195_), .A2(new_n11139_), .Z(new_n11196_));
  INV_X1     g11003(.I(new_n11196_), .ZN(new_n11197_));
  NAND2_X1   g11004(.A1(new_n11059_), .A2(new_n11056_), .ZN(new_n11198_));
  NAND2_X1   g11005(.A1(new_n11060_), .A2(new_n11053_), .ZN(new_n11199_));
  NAND2_X1   g11006(.A1(new_n11199_), .A2(new_n11198_), .ZN(new_n11200_));
  INV_X1     g11007(.I(new_n11071_), .ZN(new_n11201_));
  NOR2_X1    g11008(.A1(new_n11078_), .A2(new_n11063_), .ZN(new_n11202_));
  INV_X1     g11009(.I(new_n11202_), .ZN(new_n11203_));
  OAI21_X1   g11010(.A1(new_n11201_), .A2(new_n11077_), .B(new_n11203_), .ZN(new_n11204_));
  OAI21_X1   g11011(.A1(new_n11076_), .A2(new_n10831_), .B(new_n11073_), .ZN(new_n11205_));
  NAND2_X1   g11012(.A1(new_n11205_), .A2(new_n10993_), .ZN(new_n11206_));
  INV_X1     g11013(.I(new_n11206_), .ZN(new_n11207_));
  NOR2_X1    g11014(.A1(new_n11205_), .A2(new_n10993_), .ZN(new_n11208_));
  NOR2_X1    g11015(.A1(new_n11207_), .A2(new_n11208_), .ZN(new_n11209_));
  INV_X1     g11016(.I(new_n9659_), .ZN(new_n11210_));
  AOI22_X1   g11017(.A1(\a[31] ), .A2(\a[53] ), .B1(\a[32] ), .B2(\a[52] ), .ZN(new_n11211_));
  NOR2_X1    g11018(.A1(new_n3833_), .A2(new_n6563_), .ZN(new_n11212_));
  NOR3_X1    g11019(.A1(new_n11212_), .A2(new_n11210_), .A3(new_n11211_), .ZN(new_n11213_));
  NOR2_X1    g11020(.A1(new_n11213_), .A2(new_n11212_), .ZN(new_n11214_));
  INV_X1     g11021(.I(new_n11214_), .ZN(new_n11215_));
  OAI22_X1   g11022(.A1(new_n11215_), .A2(new_n11211_), .B1(new_n11210_), .B2(new_n11213_), .ZN(new_n11216_));
  INV_X1     g11023(.I(new_n11216_), .ZN(new_n11217_));
  XOR2_X1    g11024(.A1(new_n11209_), .A2(new_n11217_), .Z(new_n11218_));
  INV_X1     g11025(.I(new_n11218_), .ZN(new_n11219_));
  XOR2_X1    g11026(.A1(new_n11204_), .A2(new_n11219_), .Z(new_n11220_));
  XOR2_X1    g11027(.A1(new_n11220_), .A2(new_n11200_), .Z(new_n11221_));
  INV_X1     g11028(.I(new_n11221_), .ZN(new_n11222_));
  NOR2_X1    g11029(.A1(new_n11062_), .A2(new_n11080_), .ZN(new_n11223_));
  NOR2_X1    g11030(.A1(new_n11083_), .A2(new_n11223_), .ZN(new_n11224_));
  XOR2_X1    g11031(.A1(new_n11224_), .A2(new_n11222_), .Z(new_n11225_));
  NOR2_X1    g11032(.A1(new_n11225_), .A2(new_n11197_), .ZN(new_n11226_));
  AND2_X2    g11033(.A1(new_n11225_), .A2(new_n11197_), .Z(new_n11227_));
  NOR2_X1    g11034(.A1(new_n11227_), .A2(new_n11226_), .ZN(new_n11228_));
  XNOR2_X1   g11035(.A1(new_n11129_), .A2(new_n11228_), .ZN(new_n11229_));
  XOR2_X1    g11036(.A1(new_n11229_), .A2(new_n11126_), .Z(new_n11230_));
  INV_X1     g11037(.I(new_n11230_), .ZN(new_n11231_));
  NOR2_X1    g11038(.A1(new_n11097_), .A2(new_n11231_), .ZN(new_n11232_));
  INV_X1     g11039(.I(new_n11232_), .ZN(new_n11233_));
  NAND2_X1   g11040(.A1(new_n11097_), .A2(new_n11231_), .ZN(new_n11234_));
  NAND2_X1   g11041(.A1(new_n11233_), .A2(new_n11234_), .ZN(new_n11235_));
  XOR2_X1    g11042(.A1(new_n11095_), .A2(new_n11235_), .Z(\asquared[85] ));
  OAI21_X1   g11043(.A1(new_n11094_), .A2(new_n11091_), .B(new_n11233_), .ZN(new_n11237_));
  NAND2_X1   g11044(.A1(new_n11237_), .A2(new_n11234_), .ZN(new_n11238_));
  INV_X1     g11045(.I(new_n11126_), .ZN(new_n11239_));
  NAND2_X1   g11046(.A1(new_n11129_), .A2(new_n11228_), .ZN(new_n11240_));
  OAI21_X1   g11047(.A1(new_n11229_), .A2(new_n11239_), .B(new_n11240_), .ZN(new_n11241_));
  NOR2_X1    g11048(.A1(new_n11224_), .A2(new_n11222_), .ZN(new_n11242_));
  NAND2_X1   g11049(.A1(new_n11100_), .A2(new_n11103_), .ZN(new_n11243_));
  NAND2_X1   g11050(.A1(new_n11104_), .A2(new_n11114_), .ZN(new_n11244_));
  NAND2_X1   g11051(.A1(new_n11244_), .A2(new_n11243_), .ZN(new_n11245_));
  INV_X1     g11052(.I(new_n11139_), .ZN(new_n11246_));
  NOR2_X1    g11053(.A1(new_n11195_), .A2(new_n11246_), .ZN(new_n11247_));
  NOR2_X1    g11054(.A1(new_n11194_), .A2(new_n11166_), .ZN(new_n11248_));
  NAND2_X1   g11055(.A1(new_n11204_), .A2(new_n11219_), .ZN(new_n11249_));
  NAND2_X1   g11056(.A1(new_n11220_), .A2(new_n11200_), .ZN(new_n11250_));
  NAND2_X1   g11057(.A1(new_n11250_), .A2(new_n11249_), .ZN(new_n11251_));
  AOI21_X1   g11058(.A1(new_n11209_), .A2(new_n11216_), .B(new_n11207_), .ZN(new_n11252_));
  NAND2_X1   g11059(.A1(new_n11009_), .A2(new_n11004_), .ZN(new_n11253_));
  NAND2_X1   g11060(.A1(new_n11105_), .A2(new_n11070_), .ZN(new_n11254_));
  NAND2_X1   g11061(.A1(new_n11254_), .A2(new_n11253_), .ZN(new_n11255_));
  NAND2_X1   g11062(.A1(new_n10985_), .A2(new_n11018_), .ZN(new_n11256_));
  NAND2_X1   g11063(.A1(new_n11130_), .A2(new_n10978_), .ZN(new_n11257_));
  NAND2_X1   g11064(.A1(new_n11257_), .A2(new_n11256_), .ZN(new_n11258_));
  NOR2_X1    g11065(.A1(new_n11258_), .A2(new_n11255_), .ZN(new_n11259_));
  NAND2_X1   g11066(.A1(new_n11258_), .A2(new_n11255_), .ZN(new_n11260_));
  INV_X1     g11067(.I(new_n11260_), .ZN(new_n11261_));
  NOR2_X1    g11068(.A1(new_n11261_), .A2(new_n11259_), .ZN(new_n11262_));
  XNOR2_X1   g11069(.A1(new_n11262_), .A2(new_n11252_), .ZN(new_n11263_));
  XOR2_X1    g11070(.A1(new_n11251_), .A2(new_n11263_), .Z(new_n11264_));
  OAI21_X1   g11071(.A1(new_n11247_), .A2(new_n11248_), .B(new_n11264_), .ZN(new_n11265_));
  OR3_X2     g11072(.A1(new_n11264_), .A2(new_n11247_), .A3(new_n11248_), .Z(new_n11266_));
  NAND2_X1   g11073(.A1(new_n11266_), .A2(new_n11265_), .ZN(new_n11267_));
  XNOR2_X1   g11074(.A1(new_n11245_), .A2(new_n11267_), .ZN(new_n11268_));
  OR3_X2     g11075(.A1(new_n11268_), .A2(new_n11242_), .A3(new_n11227_), .Z(new_n11269_));
  OAI21_X1   g11076(.A1(new_n11227_), .A2(new_n11242_), .B(new_n11268_), .ZN(new_n11270_));
  AND2_X2    g11077(.A1(new_n11269_), .A2(new_n11270_), .Z(new_n11271_));
  INV_X1     g11078(.I(new_n11271_), .ZN(new_n11272_));
  NAND2_X1   g11079(.A1(new_n11109_), .A2(new_n11112_), .ZN(new_n11273_));
  NAND2_X1   g11080(.A1(new_n11113_), .A2(new_n11106_), .ZN(new_n11274_));
  NAND2_X1   g11081(.A1(new_n11274_), .A2(new_n11273_), .ZN(new_n11275_));
  AOI22_X1   g11082(.A1(\a[22] ), .A2(\a[63] ), .B1(\a[28] ), .B2(\a[57] ), .ZN(new_n11276_));
  INV_X1     g11083(.I(new_n11276_), .ZN(new_n11277_));
  NOR4_X1    g11084(.A1(new_n1175_), .A2(new_n1718_), .A3(new_n6298_), .A4(new_n7643_), .ZN(new_n11278_));
  NOR2_X1    g11085(.A1(new_n2524_), .A2(new_n4901_), .ZN(new_n11279_));
  AOI21_X1   g11086(.A1(new_n11277_), .A2(new_n11279_), .B(new_n11278_), .ZN(new_n11280_));
  INV_X1     g11087(.I(new_n11280_), .ZN(new_n11281_));
  OAI21_X1   g11088(.A1(new_n11278_), .A2(new_n11276_), .B(new_n11279_), .ZN(new_n11282_));
  OAI21_X1   g11089(.A1(new_n11281_), .A2(new_n11276_), .B(new_n11282_), .ZN(new_n11283_));
  NOR2_X1    g11090(.A1(new_n3932_), .A2(new_n5525_), .ZN(new_n11284_));
  NOR2_X1    g11091(.A1(new_n3375_), .A2(new_n5683_), .ZN(new_n11285_));
  NOR2_X1    g11092(.A1(new_n2637_), .A2(new_n6563_), .ZN(new_n11286_));
  NOR2_X1    g11093(.A1(new_n11285_), .A2(new_n11286_), .ZN(new_n11287_));
  NOR2_X1    g11094(.A1(new_n11287_), .A2(new_n11284_), .ZN(new_n11288_));
  NAND2_X1   g11095(.A1(\a[32] ), .A2(\a[53] ), .ZN(new_n11289_));
  AOI22_X1   g11096(.A1(\a[33] ), .A2(\a[52] ), .B1(\a[34] ), .B2(\a[51] ), .ZN(new_n11290_));
  NOR2_X1    g11097(.A1(new_n11288_), .A2(new_n11284_), .ZN(new_n11291_));
  INV_X1     g11098(.I(new_n11291_), .ZN(new_n11292_));
  OAI22_X1   g11099(.A1(new_n11292_), .A2(new_n11290_), .B1(new_n11288_), .B2(new_n11289_), .ZN(new_n11293_));
  XNOR2_X1   g11100(.A1(new_n11293_), .A2(new_n11283_), .ZN(new_n11294_));
  NOR2_X1    g11101(.A1(new_n5377_), .A2(new_n4704_), .ZN(new_n11295_));
  AOI22_X1   g11102(.A1(new_n3328_), .A2(new_n6100_), .B1(new_n3550_), .B2(new_n4429_), .ZN(new_n11296_));
  NOR2_X1    g11103(.A1(new_n11295_), .A2(new_n11296_), .ZN(new_n11297_));
  NAND2_X1   g11104(.A1(\a[39] ), .A2(\a[46] ), .ZN(new_n11298_));
  AOI22_X1   g11105(.A1(\a[40] ), .A2(\a[45] ), .B1(\a[41] ), .B2(\a[44] ), .ZN(new_n11299_));
  NOR2_X1    g11106(.A1(new_n11297_), .A2(new_n11295_), .ZN(new_n11300_));
  INV_X1     g11107(.I(new_n11300_), .ZN(new_n11301_));
  OAI22_X1   g11108(.A1(new_n11301_), .A2(new_n11299_), .B1(new_n11297_), .B2(new_n11298_), .ZN(new_n11302_));
  XOR2_X1    g11109(.A1(new_n11294_), .A2(new_n11302_), .Z(new_n11303_));
  NOR3_X1    g11110(.A1(new_n1299_), .A2(new_n3666_), .A3(new_n7144_), .ZN(new_n11304_));
  NAND2_X1   g11111(.A1(new_n11304_), .A2(new_n4180_), .ZN(new_n11305_));
  AOI21_X1   g11112(.A1(\a[23] ), .A2(\a[62] ), .B(\a[43] ), .ZN(new_n11306_));
  OR2_X2     g11113(.A1(new_n11304_), .A2(new_n4180_), .Z(new_n11307_));
  OAI21_X1   g11114(.A1(new_n11307_), .A2(new_n11306_), .B(new_n11305_), .ZN(new_n11308_));
  NOR2_X1    g11115(.A1(new_n6140_), .A2(new_n4977_), .ZN(new_n11309_));
  INV_X1     g11116(.I(new_n11309_), .ZN(new_n11310_));
  OAI22_X1   g11117(.A1(new_n2916_), .A2(new_n4979_), .B1(new_n3038_), .B2(new_n4981_), .ZN(new_n11311_));
  NAND2_X1   g11118(.A1(new_n11310_), .A2(new_n11311_), .ZN(new_n11312_));
  NAND3_X1   g11119(.A1(new_n11312_), .A2(\a[36] ), .A3(\a[49] ), .ZN(new_n11313_));
  AOI22_X1   g11120(.A1(\a[37] ), .A2(\a[48] ), .B1(\a[38] ), .B2(\a[47] ), .ZN(new_n11314_));
  NAND2_X1   g11121(.A1(new_n11312_), .A2(new_n11310_), .ZN(new_n11315_));
  OAI21_X1   g11122(.A1(new_n11314_), .A2(new_n11315_), .B(new_n11313_), .ZN(new_n11316_));
  XOR2_X1    g11123(.A1(new_n11316_), .A2(new_n11308_), .Z(new_n11317_));
  NOR2_X1    g11124(.A1(new_n2438_), .A2(new_n6129_), .ZN(new_n11318_));
  AOI22_X1   g11125(.A1(new_n2254_), .A2(new_n7184_), .B1(new_n2976_), .B2(new_n5857_), .ZN(new_n11319_));
  NOR2_X1    g11126(.A1(new_n11318_), .A2(new_n11319_), .ZN(new_n11320_));
  NAND2_X1   g11127(.A1(\a[29] ), .A2(\a[56] ), .ZN(new_n11321_));
  AOI22_X1   g11128(.A1(\a[30] ), .A2(\a[55] ), .B1(\a[31] ), .B2(\a[54] ), .ZN(new_n11322_));
  NOR2_X1    g11129(.A1(new_n11320_), .A2(new_n11318_), .ZN(new_n11323_));
  INV_X1     g11130(.I(new_n11323_), .ZN(new_n11324_));
  OAI22_X1   g11131(.A1(new_n11324_), .A2(new_n11322_), .B1(new_n11320_), .B2(new_n11321_), .ZN(new_n11325_));
  XNOR2_X1   g11132(.A1(new_n11317_), .A2(new_n11325_), .ZN(new_n11326_));
  XOR2_X1    g11133(.A1(new_n11303_), .A2(new_n11326_), .Z(new_n11327_));
  NOR2_X1    g11134(.A1(new_n11275_), .A2(new_n11327_), .ZN(new_n11328_));
  NAND2_X1   g11135(.A1(new_n11275_), .A2(new_n11327_), .ZN(new_n11329_));
  INV_X1     g11136(.I(new_n11329_), .ZN(new_n11330_));
  NOR2_X1    g11137(.A1(new_n11330_), .A2(new_n11328_), .ZN(new_n11331_));
  NAND2_X1   g11138(.A1(new_n11134_), .A2(new_n11137_), .ZN(new_n11332_));
  NAND2_X1   g11139(.A1(new_n11138_), .A2(new_n11131_), .ZN(new_n11333_));
  NAND2_X1   g11140(.A1(new_n11333_), .A2(new_n11332_), .ZN(new_n11334_));
  NOR2_X1    g11141(.A1(new_n1357_), .A2(new_n6897_), .ZN(new_n11335_));
  XOR2_X1    g11142(.A1(new_n11155_), .A2(new_n11335_), .Z(new_n11336_));
  XOR2_X1    g11143(.A1(new_n11336_), .A2(new_n11148_), .Z(new_n11337_));
  XNOR2_X1   g11144(.A1(new_n11214_), .A2(new_n11164_), .ZN(new_n11338_));
  NAND2_X1   g11145(.A1(new_n1971_), .A2(new_n7205_), .ZN(new_n11339_));
  OAI22_X1   g11146(.A1(new_n2177_), .A2(new_n7452_), .B1(new_n4010_), .B2(new_n7801_), .ZN(new_n11340_));
  NAND2_X1   g11147(.A1(new_n11340_), .A2(new_n11339_), .ZN(new_n11341_));
  NAND3_X1   g11148(.A1(new_n11341_), .A2(\a[25] ), .A3(\a[60] ), .ZN(new_n11342_));
  AOI22_X1   g11149(.A1(\a[26] ), .A2(\a[59] ), .B1(\a[27] ), .B2(\a[58] ), .ZN(new_n11343_));
  NAND2_X1   g11150(.A1(new_n11341_), .A2(new_n11339_), .ZN(new_n11344_));
  OAI21_X1   g11151(.A1(new_n11343_), .A2(new_n11344_), .B(new_n11342_), .ZN(new_n11345_));
  XOR2_X1    g11152(.A1(new_n11338_), .A2(new_n11345_), .Z(new_n11346_));
  NAND2_X1   g11153(.A1(new_n11337_), .A2(new_n11346_), .ZN(new_n11347_));
  OR2_X2     g11154(.A1(new_n11337_), .A2(new_n11346_), .Z(new_n11348_));
  NAND2_X1   g11155(.A1(new_n11348_), .A2(new_n11347_), .ZN(new_n11349_));
  NAND2_X1   g11156(.A1(new_n11334_), .A2(new_n11349_), .ZN(new_n11350_));
  INV_X1     g11157(.I(new_n11347_), .ZN(new_n11351_));
  AOI21_X1   g11158(.A1(new_n11334_), .A2(new_n11348_), .B(new_n11351_), .ZN(new_n11352_));
  NAND2_X1   g11159(.A1(new_n11352_), .A2(new_n11348_), .ZN(new_n11353_));
  NAND2_X1   g11160(.A1(new_n11353_), .A2(new_n11350_), .ZN(new_n11354_));
  NOR2_X1    g11161(.A1(new_n11175_), .A2(new_n11192_), .ZN(new_n11355_));
  NOR2_X1    g11162(.A1(new_n11174_), .A2(new_n11191_), .ZN(new_n11356_));
  NOR2_X1    g11163(.A1(new_n11355_), .A2(new_n11356_), .ZN(new_n11357_));
  INV_X1     g11164(.I(new_n11357_), .ZN(new_n11358_));
  NOR2_X1    g11165(.A1(new_n11358_), .A2(new_n11181_), .ZN(new_n11359_));
  NOR2_X1    g11166(.A1(new_n11357_), .A2(new_n11182_), .ZN(new_n11360_));
  NOR2_X1    g11167(.A1(new_n11359_), .A2(new_n11360_), .ZN(new_n11361_));
  NAND2_X1   g11168(.A1(new_n11156_), .A2(new_n11149_), .ZN(new_n11362_));
  INV_X1     g11169(.I(new_n11157_), .ZN(new_n11363_));
  NAND2_X1   g11170(.A1(new_n11363_), .A2(new_n11165_), .ZN(new_n11364_));
  NAND2_X1   g11171(.A1(new_n11364_), .A2(new_n11362_), .ZN(new_n11365_));
  NAND2_X1   g11172(.A1(new_n11176_), .A2(new_n11184_), .ZN(new_n11366_));
  INV_X1     g11173(.I(new_n11185_), .ZN(new_n11367_));
  NAND2_X1   g11174(.A1(new_n11367_), .A2(new_n11193_), .ZN(new_n11368_));
  NAND2_X1   g11175(.A1(new_n11368_), .A2(new_n11366_), .ZN(new_n11369_));
  XOR2_X1    g11176(.A1(new_n11369_), .A2(new_n11365_), .Z(new_n11370_));
  XOR2_X1    g11177(.A1(new_n11370_), .A2(new_n11361_), .Z(new_n11371_));
  XNOR2_X1   g11178(.A1(new_n11371_), .A2(new_n11354_), .ZN(new_n11372_));
  XOR2_X1    g11179(.A1(new_n11372_), .A2(new_n11331_), .Z(new_n11373_));
  NAND2_X1   g11180(.A1(new_n11118_), .A2(new_n11121_), .ZN(new_n11374_));
  NAND2_X1   g11181(.A1(new_n11124_), .A2(new_n11374_), .ZN(new_n11375_));
  XOR2_X1    g11182(.A1(new_n11375_), .A2(new_n11373_), .Z(new_n11376_));
  XOR2_X1    g11183(.A1(new_n11376_), .A2(new_n11272_), .Z(new_n11377_));
  NOR2_X1    g11184(.A1(new_n11377_), .A2(new_n11241_), .ZN(new_n11378_));
  NAND2_X1   g11185(.A1(new_n11377_), .A2(new_n11241_), .ZN(new_n11379_));
  INV_X1     g11186(.I(new_n11379_), .ZN(new_n11380_));
  NOR2_X1    g11187(.A1(new_n11380_), .A2(new_n11378_), .ZN(new_n11381_));
  XOR2_X1    g11188(.A1(new_n11238_), .A2(new_n11381_), .Z(\asquared[86] ));
  AOI21_X1   g11189(.A1(new_n11237_), .A2(new_n11234_), .B(new_n11378_), .ZN(new_n11383_));
  NOR2_X1    g11190(.A1(new_n11383_), .A2(new_n11380_), .ZN(new_n11384_));
  INV_X1     g11191(.I(new_n11373_), .ZN(new_n11385_));
  NAND2_X1   g11192(.A1(new_n11375_), .A2(new_n11385_), .ZN(new_n11386_));
  OAI21_X1   g11193(.A1(new_n11376_), .A2(new_n11272_), .B(new_n11386_), .ZN(new_n11387_));
  OAI21_X1   g11194(.A1(new_n11303_), .A2(new_n11326_), .B(new_n11329_), .ZN(new_n11388_));
  NOR2_X1    g11195(.A1(new_n11359_), .A2(new_n11356_), .ZN(new_n11389_));
  NAND2_X1   g11196(.A1(new_n11155_), .A2(new_n11335_), .ZN(new_n11390_));
  NAND2_X1   g11197(.A1(new_n11336_), .A2(new_n11148_), .ZN(new_n11391_));
  NAND2_X1   g11198(.A1(new_n11391_), .A2(new_n11390_), .ZN(new_n11392_));
  NAND2_X1   g11199(.A1(\a[25] ), .A2(\a[61] ), .ZN(new_n11393_));
  NAND2_X1   g11200(.A1(\a[24] ), .A2(\a[62] ), .ZN(new_n11394_));
  AOI22_X1   g11201(.A1(new_n1778_), .A2(new_n7590_), .B1(new_n11393_), .B2(new_n11394_), .ZN(new_n11395_));
  XOR2_X1    g11202(.A1(new_n11307_), .A2(new_n11395_), .Z(new_n11396_));
  NOR2_X1    g11203(.A1(new_n11392_), .A2(new_n11396_), .ZN(new_n11397_));
  NAND2_X1   g11204(.A1(new_n11392_), .A2(new_n11396_), .ZN(new_n11398_));
  INV_X1     g11205(.I(new_n11398_), .ZN(new_n11399_));
  NOR2_X1    g11206(.A1(new_n11399_), .A2(new_n11397_), .ZN(new_n11400_));
  XOR2_X1    g11207(.A1(new_n11400_), .A2(new_n11389_), .Z(new_n11401_));
  XOR2_X1    g11208(.A1(new_n11352_), .A2(new_n11401_), .Z(new_n11402_));
  XNOR2_X1   g11209(.A1(new_n11388_), .A2(new_n11402_), .ZN(new_n11403_));
  INV_X1     g11210(.I(new_n11331_), .ZN(new_n11404_));
  NAND2_X1   g11211(.A1(new_n11371_), .A2(new_n11354_), .ZN(new_n11405_));
  OAI21_X1   g11212(.A1(new_n11372_), .A2(new_n11404_), .B(new_n11405_), .ZN(new_n11406_));
  NAND2_X1   g11213(.A1(new_n11251_), .A2(new_n11263_), .ZN(new_n11407_));
  NAND2_X1   g11214(.A1(new_n11265_), .A2(new_n11407_), .ZN(new_n11408_));
  XOR2_X1    g11215(.A1(new_n11408_), .A2(new_n11406_), .Z(new_n11409_));
  XNOR2_X1   g11216(.A1(new_n11409_), .A2(new_n11403_), .ZN(new_n11410_));
  NAND2_X1   g11217(.A1(new_n11369_), .A2(new_n11365_), .ZN(new_n11411_));
  NAND2_X1   g11218(.A1(new_n11370_), .A2(new_n11361_), .ZN(new_n11412_));
  NAND2_X1   g11219(.A1(new_n11412_), .A2(new_n11411_), .ZN(new_n11413_));
  AOI22_X1   g11220(.A1(\a[36] ), .A2(\a[50] ), .B1(\a[37] ), .B2(\a[49] ), .ZN(new_n11414_));
  INV_X1     g11221(.I(new_n11414_), .ZN(new_n11415_));
  NOR2_X1    g11222(.A1(new_n3038_), .A2(new_n5155_), .ZN(new_n11416_));
  NOR2_X1    g11223(.A1(new_n1299_), .A2(new_n7643_), .ZN(new_n11417_));
  AOI21_X1   g11224(.A1(new_n11415_), .A2(new_n11417_), .B(new_n11416_), .ZN(new_n11418_));
  INV_X1     g11225(.I(new_n11418_), .ZN(new_n11419_));
  OAI21_X1   g11226(.A1(new_n11416_), .A2(new_n11414_), .B(new_n11417_), .ZN(new_n11420_));
  OAI21_X1   g11227(.A1(new_n11419_), .A2(new_n11414_), .B(new_n11420_), .ZN(new_n11421_));
  NOR2_X1    g11228(.A1(new_n2746_), .A2(new_n5525_), .ZN(new_n11422_));
  NOR2_X1    g11229(.A1(new_n2526_), .A2(new_n5683_), .ZN(new_n11423_));
  NOR2_X1    g11230(.A1(new_n3932_), .A2(new_n6563_), .ZN(new_n11424_));
  NOR2_X1    g11231(.A1(new_n11423_), .A2(new_n11424_), .ZN(new_n11425_));
  NOR2_X1    g11232(.A1(new_n11425_), .A2(new_n11422_), .ZN(new_n11426_));
  NAND2_X1   g11233(.A1(\a[33] ), .A2(\a[53] ), .ZN(new_n11427_));
  AOI22_X1   g11234(.A1(\a[34] ), .A2(\a[52] ), .B1(\a[35] ), .B2(\a[51] ), .ZN(new_n11428_));
  NOR2_X1    g11235(.A1(new_n11426_), .A2(new_n11422_), .ZN(new_n11429_));
  INV_X1     g11236(.I(new_n11429_), .ZN(new_n11430_));
  OAI22_X1   g11237(.A1(new_n11430_), .A2(new_n11428_), .B1(new_n11426_), .B2(new_n11427_), .ZN(new_n11431_));
  XNOR2_X1   g11238(.A1(new_n11431_), .A2(new_n11421_), .ZN(new_n11432_));
  INV_X1     g11239(.I(new_n5574_), .ZN(new_n11433_));
  AOI22_X1   g11240(.A1(\a[29] ), .A2(\a[57] ), .B1(\a[31] ), .B2(\a[55] ), .ZN(new_n11434_));
  NOR2_X1    g11241(.A1(new_n5625_), .A2(new_n8952_), .ZN(new_n11435_));
  NOR3_X1    g11242(.A1(new_n11435_), .A2(new_n11433_), .A3(new_n11434_), .ZN(new_n11436_));
  NOR2_X1    g11243(.A1(new_n11436_), .A2(new_n11435_), .ZN(new_n11437_));
  INV_X1     g11244(.I(new_n11437_), .ZN(new_n11438_));
  OAI22_X1   g11245(.A1(new_n11438_), .A2(new_n11434_), .B1(new_n11433_), .B2(new_n11436_), .ZN(new_n11439_));
  INV_X1     g11246(.I(new_n11439_), .ZN(new_n11440_));
  XOR2_X1    g11247(.A1(new_n11432_), .A2(new_n11440_), .Z(new_n11441_));
  NOR2_X1    g11248(.A1(new_n2189_), .A2(new_n7206_), .ZN(new_n11442_));
  INV_X1     g11249(.I(new_n11442_), .ZN(new_n11443_));
  OAI22_X1   g11250(.A1(new_n1972_), .A2(new_n7452_), .B1(new_n3341_), .B2(new_n7801_), .ZN(new_n11444_));
  NAND2_X1   g11251(.A1(new_n11444_), .A2(new_n11443_), .ZN(new_n11445_));
  NAND3_X1   g11252(.A1(new_n11445_), .A2(\a[26] ), .A3(\a[60] ), .ZN(new_n11446_));
  AOI22_X1   g11253(.A1(\a[27] ), .A2(\a[59] ), .B1(\a[28] ), .B2(\a[58] ), .ZN(new_n11447_));
  NAND2_X1   g11254(.A1(new_n11445_), .A2(new_n11443_), .ZN(new_n11448_));
  OAI21_X1   g11255(.A1(new_n11447_), .A2(new_n11448_), .B(new_n11446_), .ZN(new_n11449_));
  NOR2_X1    g11256(.A1(new_n2200_), .A2(new_n5617_), .ZN(new_n11450_));
  INV_X1     g11257(.I(new_n11450_), .ZN(new_n11451_));
  OAI22_X1   g11258(.A1(new_n4032_), .A2(new_n11451_), .B1(new_n4667_), .B2(new_n4704_), .ZN(new_n11452_));
  NOR2_X1    g11259(.A1(new_n3861_), .A2(new_n11451_), .ZN(new_n11453_));
  INV_X1     g11260(.I(new_n11453_), .ZN(new_n11454_));
  AND2_X2    g11261(.A1(new_n11454_), .A2(new_n11452_), .Z(new_n11455_));
  NOR2_X1    g11262(.A1(new_n3860_), .A2(new_n11450_), .ZN(new_n11456_));
  NOR2_X1    g11263(.A1(new_n11452_), .A2(new_n11453_), .ZN(new_n11457_));
  INV_X1     g11264(.I(new_n11457_), .ZN(new_n11458_));
  OAI22_X1   g11265(.A1(new_n4032_), .A2(new_n11455_), .B1(new_n11458_), .B2(new_n11456_), .ZN(new_n11459_));
  XOR2_X1    g11266(.A1(new_n11449_), .A2(new_n11459_), .Z(new_n11460_));
  AOI22_X1   g11267(.A1(\a[39] ), .A2(\a[47] ), .B1(\a[40] ), .B2(\a[46] ), .ZN(new_n11461_));
  NAND2_X1   g11268(.A1(\a[30] ), .A2(\a[56] ), .ZN(new_n11462_));
  NOR2_X1    g11269(.A1(new_n3551_), .A2(new_n4721_), .ZN(new_n11463_));
  NOR3_X1    g11270(.A1(new_n11463_), .A2(new_n11461_), .A3(new_n11462_), .ZN(new_n11464_));
  NOR2_X1    g11271(.A1(new_n11464_), .A2(new_n11463_), .ZN(new_n11465_));
  INV_X1     g11272(.I(new_n11465_), .ZN(new_n11466_));
  OAI22_X1   g11273(.A1(new_n11466_), .A2(new_n11461_), .B1(new_n11462_), .B2(new_n11464_), .ZN(new_n11467_));
  XNOR2_X1   g11274(.A1(new_n11460_), .A2(new_n11467_), .ZN(new_n11468_));
  INV_X1     g11275(.I(new_n11468_), .ZN(new_n11469_));
  XOR2_X1    g11276(.A1(new_n11441_), .A2(new_n11469_), .Z(new_n11470_));
  XOR2_X1    g11277(.A1(new_n11413_), .A2(new_n11470_), .Z(new_n11471_));
  OAI21_X1   g11278(.A1(new_n11252_), .A2(new_n11259_), .B(new_n11260_), .ZN(new_n11472_));
  INV_X1     g11279(.I(new_n11472_), .ZN(new_n11473_));
  NOR2_X1    g11280(.A1(new_n11301_), .A2(new_n11324_), .ZN(new_n11474_));
  NOR2_X1    g11281(.A1(new_n11300_), .A2(new_n11323_), .ZN(new_n11475_));
  NOR2_X1    g11282(.A1(new_n11474_), .A2(new_n11475_), .ZN(new_n11476_));
  NAND2_X1   g11283(.A1(new_n11476_), .A2(new_n11315_), .ZN(new_n11477_));
  INV_X1     g11284(.I(new_n11477_), .ZN(new_n11478_));
  NOR2_X1    g11285(.A1(new_n11476_), .A2(new_n11315_), .ZN(new_n11479_));
  NOR2_X1    g11286(.A1(new_n11478_), .A2(new_n11479_), .ZN(new_n11480_));
  XNOR2_X1   g11287(.A1(new_n11291_), .A2(new_n11344_), .ZN(new_n11481_));
  XOR2_X1    g11288(.A1(new_n11481_), .A2(new_n11281_), .Z(new_n11482_));
  XNOR2_X1   g11289(.A1(new_n11482_), .A2(new_n11480_), .ZN(new_n11483_));
  XOR2_X1    g11290(.A1(new_n11483_), .A2(new_n11473_), .Z(new_n11484_));
  INV_X1     g11291(.I(new_n11484_), .ZN(new_n11485_));
  NAND2_X1   g11292(.A1(new_n11316_), .A2(new_n11308_), .ZN(new_n11486_));
  NAND2_X1   g11293(.A1(new_n11317_), .A2(new_n11325_), .ZN(new_n11487_));
  NAND2_X1   g11294(.A1(new_n11487_), .A2(new_n11486_), .ZN(new_n11488_));
  NAND2_X1   g11295(.A1(new_n11215_), .A2(new_n11164_), .ZN(new_n11489_));
  NAND2_X1   g11296(.A1(new_n11338_), .A2(new_n11345_), .ZN(new_n11490_));
  NAND2_X1   g11297(.A1(new_n11490_), .A2(new_n11489_), .ZN(new_n11491_));
  NAND2_X1   g11298(.A1(new_n11293_), .A2(new_n11283_), .ZN(new_n11492_));
  INV_X1     g11299(.I(new_n11294_), .ZN(new_n11493_));
  NAND2_X1   g11300(.A1(new_n11493_), .A2(new_n11302_), .ZN(new_n11494_));
  NAND2_X1   g11301(.A1(new_n11494_), .A2(new_n11492_), .ZN(new_n11495_));
  XOR2_X1    g11302(.A1(new_n11495_), .A2(new_n11491_), .Z(new_n11496_));
  XOR2_X1    g11303(.A1(new_n11496_), .A2(new_n11488_), .Z(new_n11497_));
  INV_X1     g11304(.I(new_n11497_), .ZN(new_n11498_));
  NOR2_X1    g11305(.A1(new_n11498_), .A2(new_n11485_), .ZN(new_n11499_));
  NOR2_X1    g11306(.A1(new_n11497_), .A2(new_n11484_), .ZN(new_n11500_));
  NOR2_X1    g11307(.A1(new_n11499_), .A2(new_n11500_), .ZN(new_n11501_));
  NAND2_X1   g11308(.A1(new_n11501_), .A2(new_n11471_), .ZN(new_n11502_));
  INV_X1     g11309(.I(new_n11502_), .ZN(new_n11503_));
  NOR2_X1    g11310(.A1(new_n11501_), .A2(new_n11471_), .ZN(new_n11504_));
  NOR2_X1    g11311(.A1(new_n11503_), .A2(new_n11504_), .ZN(new_n11505_));
  INV_X1     g11312(.I(new_n11245_), .ZN(new_n11506_));
  OAI21_X1   g11313(.A1(new_n11506_), .A2(new_n11267_), .B(new_n11270_), .ZN(new_n11507_));
  NAND2_X1   g11314(.A1(new_n11507_), .A2(new_n11505_), .ZN(new_n11508_));
  NAND2_X1   g11315(.A1(new_n11508_), .A2(new_n11505_), .ZN(new_n11509_));
  NAND2_X1   g11316(.A1(new_n11508_), .A2(new_n11507_), .ZN(new_n11510_));
  NAND2_X1   g11317(.A1(new_n11510_), .A2(new_n11509_), .ZN(new_n11511_));
  AOI21_X1   g11318(.A1(new_n11508_), .A2(new_n11507_), .B(new_n11410_), .ZN(new_n11512_));
  AOI22_X1   g11319(.A1(new_n11511_), .A2(new_n11410_), .B1(new_n11509_), .B2(new_n11512_), .ZN(new_n11513_));
  NAND2_X1   g11320(.A1(new_n11387_), .A2(new_n11513_), .ZN(new_n11514_));
  NOR2_X1    g11321(.A1(new_n11387_), .A2(new_n11513_), .ZN(new_n11515_));
  INV_X1     g11322(.I(new_n11515_), .ZN(new_n11516_));
  NAND2_X1   g11323(.A1(new_n11516_), .A2(new_n11514_), .ZN(new_n11517_));
  INV_X1     g11324(.I(new_n11234_), .ZN(new_n11518_));
  INV_X1     g11325(.I(new_n11091_), .ZN(new_n11519_));
  INV_X1     g11326(.I(new_n10952_), .ZN(new_n11520_));
  INV_X1     g11327(.I(new_n10649_), .ZN(new_n11521_));
  INV_X1     g11328(.I(new_n10811_), .ZN(new_n11522_));
  OAI21_X1   g11329(.A1(new_n10667_), .A2(new_n11521_), .B(new_n11522_), .ZN(new_n11523_));
  AOI21_X1   g11330(.A1(new_n11523_), .A2(new_n10812_), .B(new_n10950_), .ZN(new_n11524_));
  INV_X1     g11331(.I(new_n11090_), .ZN(new_n11525_));
  OAI21_X1   g11332(.A1(new_n11524_), .A2(new_n11520_), .B(new_n11525_), .ZN(new_n11526_));
  AOI21_X1   g11333(.A1(new_n11526_), .A2(new_n11519_), .B(new_n11232_), .ZN(new_n11527_));
  INV_X1     g11334(.I(new_n11378_), .ZN(new_n11528_));
  OAI21_X1   g11335(.A1(new_n11527_), .A2(new_n11518_), .B(new_n11528_), .ZN(new_n11529_));
  AOI21_X1   g11336(.A1(new_n11529_), .A2(new_n11379_), .B(new_n11515_), .ZN(new_n11530_));
  AOI22_X1   g11337(.A1(new_n11530_), .A2(new_n11514_), .B1(new_n11384_), .B2(new_n11517_), .ZN(\asquared[87] ));
  OAI21_X1   g11338(.A1(new_n11383_), .A2(new_n11380_), .B(new_n11516_), .ZN(new_n11532_));
  NAND2_X1   g11339(.A1(new_n11532_), .A2(new_n11514_), .ZN(new_n11533_));
  NAND2_X1   g11340(.A1(new_n11511_), .A2(new_n11410_), .ZN(new_n11534_));
  NAND2_X1   g11341(.A1(new_n11534_), .A2(new_n11508_), .ZN(new_n11535_));
  NOR2_X1    g11342(.A1(new_n11503_), .A2(new_n11499_), .ZN(new_n11536_));
  NAND2_X1   g11343(.A1(new_n3232_), .A2(new_n5524_), .ZN(new_n11537_));
  NAND4_X1   g11344(.A1(\a[29] ), .A2(\a[35] ), .A3(\a[52] ), .A4(\a[58] ), .ZN(new_n11538_));
  NOR4_X1    g11345(.A1(new_n1814_), .A2(new_n2626_), .A3(new_n5135_), .A4(new_n6316_), .ZN(new_n11539_));
  AOI21_X1   g11346(.A1(new_n11537_), .A2(new_n11538_), .B(new_n11539_), .ZN(new_n11540_));
  NAND2_X1   g11347(.A1(\a[35] ), .A2(\a[52] ), .ZN(new_n11541_));
  AOI22_X1   g11348(.A1(\a[29] ), .A2(\a[58] ), .B1(\a[36] ), .B2(\a[51] ), .ZN(new_n11542_));
  NAND2_X1   g11349(.A1(new_n11537_), .A2(new_n11538_), .ZN(new_n11543_));
  NOR2_X1    g11350(.A1(new_n11543_), .A2(new_n11539_), .ZN(new_n11544_));
  INV_X1     g11351(.I(new_n11544_), .ZN(new_n11545_));
  OAI22_X1   g11352(.A1(new_n11545_), .A2(new_n11542_), .B1(new_n11540_), .B2(new_n11541_), .ZN(new_n11546_));
  NOR2_X1    g11353(.A1(new_n2442_), .A2(new_n5425_), .ZN(new_n11547_));
  NAND2_X1   g11354(.A1(new_n11160_), .A2(new_n11547_), .ZN(new_n11548_));
  INV_X1     g11355(.I(new_n11548_), .ZN(new_n11549_));
  NOR2_X1    g11356(.A1(new_n2442_), .A2(new_n6548_), .ZN(new_n11550_));
  INV_X1     g11357(.I(new_n11550_), .ZN(new_n11551_));
  NOR3_X1    g11358(.A1(new_n11551_), .A2(new_n1718_), .A3(new_n5425_), .ZN(new_n11552_));
  NOR2_X1    g11359(.A1(new_n3811_), .A2(new_n7204_), .ZN(new_n11553_));
  NOR2_X1    g11360(.A1(new_n11552_), .A2(new_n11553_), .ZN(new_n11554_));
  NOR2_X1    g11361(.A1(new_n11554_), .A2(new_n11549_), .ZN(new_n11555_));
  NAND2_X1   g11362(.A1(\a[28] ), .A2(\a[59] ), .ZN(new_n11556_));
  NOR2_X1    g11363(.A1(new_n11555_), .A2(new_n11549_), .ZN(new_n11557_));
  INV_X1     g11364(.I(new_n11557_), .ZN(new_n11558_));
  NOR2_X1    g11365(.A1(new_n11160_), .A2(new_n11547_), .ZN(new_n11559_));
  OAI22_X1   g11366(.A1(new_n11558_), .A2(new_n11559_), .B1(new_n11555_), .B2(new_n11556_), .ZN(new_n11560_));
  NAND2_X1   g11367(.A1(new_n11307_), .A2(new_n11395_), .ZN(new_n11561_));
  OAI21_X1   g11368(.A1(new_n1779_), .A2(new_n7591_), .B(new_n11561_), .ZN(new_n11562_));
  XNOR2_X1   g11369(.A1(new_n11560_), .A2(new_n11562_), .ZN(new_n11563_));
  INV_X1     g11370(.I(new_n11563_), .ZN(new_n11564_));
  NOR2_X1    g11371(.A1(new_n11564_), .A2(new_n11546_), .ZN(new_n11565_));
  NAND2_X1   g11372(.A1(new_n11564_), .A2(new_n11546_), .ZN(new_n11566_));
  INV_X1     g11373(.I(new_n11566_), .ZN(new_n11567_));
  NOR2_X1    g11374(.A1(new_n11567_), .A2(new_n11565_), .ZN(new_n11568_));
  NAND2_X1   g11375(.A1(new_n11292_), .A2(new_n11344_), .ZN(new_n11569_));
  NAND2_X1   g11376(.A1(new_n11481_), .A2(new_n11281_), .ZN(new_n11570_));
  NAND2_X1   g11377(.A1(new_n11570_), .A2(new_n11569_), .ZN(new_n11571_));
  AOI22_X1   g11378(.A1(\a[31] ), .A2(\a[56] ), .B1(\a[33] ), .B2(\a[54] ), .ZN(new_n11572_));
  INV_X1     g11379(.I(new_n11572_), .ZN(new_n11573_));
  NOR2_X1    g11380(.A1(new_n2276_), .A2(new_n6058_), .ZN(new_n11574_));
  NOR2_X1    g11381(.A1(new_n3221_), .A2(new_n4312_), .ZN(new_n11575_));
  AOI21_X1   g11382(.A1(new_n11573_), .A2(new_n11575_), .B(new_n11574_), .ZN(new_n11576_));
  NAND2_X1   g11383(.A1(new_n11576_), .A2(new_n11573_), .ZN(new_n11577_));
  OAI21_X1   g11384(.A1(new_n11574_), .A2(new_n11572_), .B(new_n11575_), .ZN(new_n11578_));
  NAND2_X1   g11385(.A1(new_n11577_), .A2(new_n11578_), .ZN(new_n11579_));
  NOR2_X1    g11386(.A1(new_n3859_), .A2(new_n7144_), .ZN(new_n11580_));
  INV_X1     g11387(.I(new_n11580_), .ZN(new_n11581_));
  NOR3_X1    g11388(.A1(new_n4343_), .A2(new_n11581_), .A3(new_n1441_), .ZN(new_n11582_));
  AOI21_X1   g11389(.A1(\a[25] ), .A2(\a[62] ), .B(\a[44] ), .ZN(new_n11583_));
  NOR2_X1    g11390(.A1(new_n11581_), .A2(new_n1441_), .ZN(new_n11584_));
  NOR2_X1    g11391(.A1(new_n11584_), .A2(new_n4342_), .ZN(new_n11585_));
  INV_X1     g11392(.I(new_n11585_), .ZN(new_n11586_));
  NOR2_X1    g11393(.A1(new_n11586_), .A2(new_n11583_), .ZN(new_n11587_));
  NOR2_X1    g11394(.A1(new_n11587_), .A2(new_n11582_), .ZN(new_n11588_));
  XNOR2_X1   g11395(.A1(new_n11588_), .A2(new_n11579_), .ZN(new_n11589_));
  AND2_X2    g11396(.A1(new_n11571_), .A2(new_n11589_), .Z(new_n11590_));
  NOR2_X1    g11397(.A1(new_n11571_), .A2(new_n11589_), .ZN(new_n11591_));
  NOR2_X1    g11398(.A1(new_n11590_), .A2(new_n11591_), .ZN(new_n11592_));
  NAND2_X1   g11399(.A1(new_n1971_), .A2(new_n7453_), .ZN(new_n11593_));
  NOR3_X1    g11400(.A1(new_n9031_), .A2(new_n1357_), .A3(new_n1750_), .ZN(new_n11594_));
  NOR2_X1    g11401(.A1(new_n2081_), .A2(new_n7959_), .ZN(new_n11595_));
  OAI21_X1   g11402(.A1(new_n11594_), .A2(new_n11595_), .B(new_n11593_), .ZN(new_n11596_));
  NAND3_X1   g11403(.A1(new_n11596_), .A2(\a[24] ), .A3(\a[63] ), .ZN(new_n11597_));
  AOI22_X1   g11404(.A1(\a[26] ), .A2(\a[61] ), .B1(\a[27] ), .B2(\a[60] ), .ZN(new_n11598_));
  NAND2_X1   g11405(.A1(new_n11596_), .A2(new_n11593_), .ZN(new_n11599_));
  OAI21_X1   g11406(.A1(new_n11598_), .A2(new_n11599_), .B(new_n11597_), .ZN(new_n11600_));
  NAND2_X1   g11407(.A1(new_n4209_), .A2(new_n4980_), .ZN(new_n11601_));
  OAI22_X1   g11408(.A1(new_n6140_), .A2(new_n5155_), .B1(new_n4739_), .B2(new_n4903_), .ZN(new_n11602_));
  NAND2_X1   g11409(.A1(new_n11602_), .A2(new_n11601_), .ZN(new_n11603_));
  NAND3_X1   g11410(.A1(new_n11603_), .A2(\a[37] ), .A3(\a[50] ), .ZN(new_n11604_));
  AOI22_X1   g11411(.A1(\a[38] ), .A2(\a[49] ), .B1(\a[39] ), .B2(\a[48] ), .ZN(new_n11605_));
  NAND2_X1   g11412(.A1(new_n11603_), .A2(new_n11601_), .ZN(new_n11606_));
  OAI21_X1   g11413(.A1(new_n11605_), .A2(new_n11606_), .B(new_n11604_), .ZN(new_n11607_));
  XOR2_X1    g11414(.A1(new_n11607_), .A2(new_n11600_), .Z(new_n11608_));
  AOI22_X1   g11415(.A1(\a[41] ), .A2(\a[46] ), .B1(\a[42] ), .B2(\a[45] ), .ZN(new_n11609_));
  NAND2_X1   g11416(.A1(\a[32] ), .A2(\a[55] ), .ZN(new_n11610_));
  NOR2_X1    g11417(.A1(new_n4667_), .A2(new_n4430_), .ZN(new_n11611_));
  NOR3_X1    g11418(.A1(new_n11611_), .A2(new_n11609_), .A3(new_n11610_), .ZN(new_n11612_));
  OAI22_X1   g11419(.A1(new_n4667_), .A2(new_n4430_), .B1(new_n11609_), .B2(new_n11610_), .ZN(new_n11613_));
  OAI22_X1   g11420(.A1(new_n11612_), .A2(new_n11610_), .B1(new_n11609_), .B2(new_n11613_), .ZN(new_n11614_));
  XOR2_X1    g11421(.A1(new_n11608_), .A2(new_n11614_), .Z(new_n11615_));
  XOR2_X1    g11422(.A1(new_n11592_), .A2(new_n11615_), .Z(new_n11616_));
  XOR2_X1    g11423(.A1(new_n11616_), .A2(new_n11568_), .Z(new_n11617_));
  INV_X1     g11424(.I(new_n11617_), .ZN(new_n11618_));
  XOR2_X1    g11425(.A1(new_n11536_), .A2(new_n11618_), .Z(new_n11619_));
  INV_X1     g11426(.I(new_n11400_), .ZN(new_n11620_));
  NOR2_X1    g11427(.A1(new_n11620_), .A2(new_n11389_), .ZN(new_n11621_));
  NOR2_X1    g11428(.A1(new_n11621_), .A2(new_n11399_), .ZN(new_n11622_));
  INV_X1     g11429(.I(new_n11622_), .ZN(new_n11623_));
  NAND2_X1   g11430(.A1(new_n11465_), .A2(new_n11457_), .ZN(new_n11624_));
  NAND2_X1   g11431(.A1(new_n11466_), .A2(new_n11458_), .ZN(new_n11625_));
  AND2_X2    g11432(.A1(new_n11625_), .A2(new_n11624_), .Z(new_n11626_));
  XOR2_X1    g11433(.A1(new_n11626_), .A2(new_n11438_), .Z(new_n11627_));
  NOR2_X1    g11434(.A1(new_n11430_), .A2(new_n11448_), .ZN(new_n11628_));
  NAND2_X1   g11435(.A1(new_n11430_), .A2(new_n11448_), .ZN(new_n11629_));
  INV_X1     g11436(.I(new_n11629_), .ZN(new_n11630_));
  NOR2_X1    g11437(.A1(new_n11630_), .A2(new_n11628_), .ZN(new_n11631_));
  NOR2_X1    g11438(.A1(new_n11631_), .A2(new_n11419_), .ZN(new_n11632_));
  INV_X1     g11439(.I(new_n11631_), .ZN(new_n11633_));
  NOR2_X1    g11440(.A1(new_n11633_), .A2(new_n11418_), .ZN(new_n11634_));
  NOR2_X1    g11441(.A1(new_n11634_), .A2(new_n11632_), .ZN(new_n11635_));
  NAND2_X1   g11442(.A1(new_n11635_), .A2(new_n11627_), .ZN(new_n11636_));
  INV_X1     g11443(.I(new_n11636_), .ZN(new_n11637_));
  NOR2_X1    g11444(.A1(new_n11635_), .A2(new_n11627_), .ZN(new_n11638_));
  NOR2_X1    g11445(.A1(new_n11637_), .A2(new_n11638_), .ZN(new_n11639_));
  NOR2_X1    g11446(.A1(new_n11623_), .A2(new_n11639_), .ZN(new_n11640_));
  NAND2_X1   g11447(.A1(new_n11623_), .A2(new_n11639_), .ZN(new_n11641_));
  INV_X1     g11448(.I(new_n11641_), .ZN(new_n11642_));
  NOR2_X1    g11449(.A1(new_n11642_), .A2(new_n11640_), .ZN(new_n11643_));
  NAND2_X1   g11450(.A1(new_n11482_), .A2(new_n11480_), .ZN(new_n11644_));
  OAI21_X1   g11451(.A1(new_n11483_), .A2(new_n11473_), .B(new_n11644_), .ZN(new_n11645_));
  NAND2_X1   g11452(.A1(new_n11495_), .A2(new_n11491_), .ZN(new_n11646_));
  NAND2_X1   g11453(.A1(new_n11496_), .A2(new_n11488_), .ZN(new_n11647_));
  NAND2_X1   g11454(.A1(new_n11647_), .A2(new_n11646_), .ZN(new_n11648_));
  XOR2_X1    g11455(.A1(new_n11648_), .A2(new_n11645_), .Z(new_n11649_));
  XOR2_X1    g11456(.A1(new_n11649_), .A2(new_n11643_), .Z(new_n11650_));
  XNOR2_X1   g11457(.A1(new_n11619_), .A2(new_n11650_), .ZN(new_n11651_));
  NAND2_X1   g11458(.A1(new_n11388_), .A2(new_n11402_), .ZN(new_n11652_));
  OAI21_X1   g11459(.A1(new_n11352_), .A2(new_n11401_), .B(new_n11652_), .ZN(new_n11653_));
  NAND2_X1   g11460(.A1(new_n11441_), .A2(new_n11469_), .ZN(new_n11654_));
  NAND2_X1   g11461(.A1(new_n11413_), .A2(new_n11470_), .ZN(new_n11655_));
  NAND2_X1   g11462(.A1(new_n11655_), .A2(new_n11654_), .ZN(new_n11656_));
  NAND2_X1   g11463(.A1(new_n11449_), .A2(new_n11459_), .ZN(new_n11657_));
  NAND2_X1   g11464(.A1(new_n11460_), .A2(new_n11467_), .ZN(new_n11658_));
  NAND2_X1   g11465(.A1(new_n11658_), .A2(new_n11657_), .ZN(new_n11659_));
  NOR2_X1    g11466(.A1(new_n11478_), .A2(new_n11475_), .ZN(new_n11660_));
  INV_X1     g11467(.I(new_n11660_), .ZN(new_n11661_));
  NAND2_X1   g11468(.A1(new_n11431_), .A2(new_n11421_), .ZN(new_n11662_));
  OAI21_X1   g11469(.A1(new_n11432_), .A2(new_n11440_), .B(new_n11662_), .ZN(new_n11663_));
  NOR2_X1    g11470(.A1(new_n11663_), .A2(new_n11661_), .ZN(new_n11664_));
  NAND2_X1   g11471(.A1(new_n11663_), .A2(new_n11661_), .ZN(new_n11665_));
  INV_X1     g11472(.I(new_n11665_), .ZN(new_n11666_));
  NOR2_X1    g11473(.A1(new_n11666_), .A2(new_n11664_), .ZN(new_n11667_));
  NAND2_X1   g11474(.A1(new_n11667_), .A2(new_n11659_), .ZN(new_n11668_));
  INV_X1     g11475(.I(new_n11668_), .ZN(new_n11669_));
  NOR2_X1    g11476(.A1(new_n11667_), .A2(new_n11659_), .ZN(new_n11670_));
  NOR2_X1    g11477(.A1(new_n11669_), .A2(new_n11670_), .ZN(new_n11671_));
  XOR2_X1    g11478(.A1(new_n11656_), .A2(new_n11671_), .Z(new_n11672_));
  XOR2_X1    g11479(.A1(new_n11672_), .A2(new_n11653_), .Z(new_n11673_));
  NAND2_X1   g11480(.A1(new_n11408_), .A2(new_n11406_), .ZN(new_n11674_));
  INV_X1     g11481(.I(new_n11409_), .ZN(new_n11675_));
  OAI21_X1   g11482(.A1(new_n11675_), .A2(new_n11403_), .B(new_n11674_), .ZN(new_n11676_));
  XNOR2_X1   g11483(.A1(new_n11676_), .A2(new_n11673_), .ZN(new_n11677_));
  XOR2_X1    g11484(.A1(new_n11677_), .A2(new_n11651_), .Z(new_n11678_));
  NOR2_X1    g11485(.A1(new_n11535_), .A2(new_n11678_), .ZN(new_n11679_));
  NAND2_X1   g11486(.A1(new_n11535_), .A2(new_n11678_), .ZN(new_n11680_));
  INV_X1     g11487(.I(new_n11680_), .ZN(new_n11681_));
  NOR2_X1    g11488(.A1(new_n11681_), .A2(new_n11679_), .ZN(new_n11682_));
  XOR2_X1    g11489(.A1(new_n11533_), .A2(new_n11682_), .Z(\asquared[88] ));
  AOI21_X1   g11490(.A1(new_n11532_), .A2(new_n11514_), .B(new_n11679_), .ZN(new_n11684_));
  NOR2_X1    g11491(.A1(new_n11684_), .A2(new_n11681_), .ZN(new_n11685_));
  NAND2_X1   g11492(.A1(new_n11619_), .A2(new_n11650_), .ZN(new_n11686_));
  OAI21_X1   g11493(.A1(new_n11536_), .A2(new_n11618_), .B(new_n11686_), .ZN(new_n11687_));
  NAND2_X1   g11494(.A1(new_n11648_), .A2(new_n11645_), .ZN(new_n11688_));
  NAND2_X1   g11495(.A1(new_n11649_), .A2(new_n11643_), .ZN(new_n11689_));
  NAND2_X1   g11496(.A1(new_n11689_), .A2(new_n11688_), .ZN(new_n11690_));
  NAND2_X1   g11497(.A1(new_n11607_), .A2(new_n11600_), .ZN(new_n11691_));
  NAND2_X1   g11498(.A1(new_n11608_), .A2(new_n11614_), .ZN(new_n11692_));
  NAND2_X1   g11499(.A1(new_n11692_), .A2(new_n11691_), .ZN(new_n11693_));
  AOI21_X1   g11500(.A1(new_n11560_), .A2(new_n11562_), .B(new_n11567_), .ZN(new_n11694_));
  NOR2_X1    g11501(.A1(new_n11634_), .A2(new_n11630_), .ZN(new_n11695_));
  XOR2_X1    g11502(.A1(new_n11694_), .A2(new_n11695_), .Z(new_n11696_));
  NAND2_X1   g11503(.A1(new_n11696_), .A2(new_n11693_), .ZN(new_n11697_));
  INV_X1     g11504(.I(new_n11697_), .ZN(new_n11698_));
  NOR2_X1    g11505(.A1(new_n11696_), .A2(new_n11693_), .ZN(new_n11699_));
  NOR2_X1    g11506(.A1(new_n11698_), .A2(new_n11699_), .ZN(new_n11700_));
  NAND2_X1   g11507(.A1(new_n11592_), .A2(new_n11615_), .ZN(new_n11701_));
  NAND2_X1   g11508(.A1(new_n11616_), .A2(new_n11568_), .ZN(new_n11702_));
  NAND2_X1   g11509(.A1(new_n11702_), .A2(new_n11701_), .ZN(new_n11703_));
  XOR2_X1    g11510(.A1(new_n11700_), .A2(new_n11703_), .Z(new_n11704_));
  XOR2_X1    g11511(.A1(new_n11704_), .A2(new_n11690_), .Z(new_n11705_));
  NOR2_X1    g11512(.A1(new_n11687_), .A2(new_n11705_), .ZN(new_n11706_));
  NAND2_X1   g11513(.A1(new_n11687_), .A2(new_n11705_), .ZN(new_n11707_));
  INV_X1     g11514(.I(new_n11707_), .ZN(new_n11708_));
  NOR2_X1    g11515(.A1(new_n11708_), .A2(new_n11706_), .ZN(new_n11709_));
  XNOR2_X1   g11516(.A1(new_n11557_), .A2(new_n11599_), .ZN(new_n11710_));
  XOR2_X1    g11517(.A1(new_n11710_), .A2(new_n11606_), .Z(new_n11711_));
  INV_X1     g11518(.I(new_n11588_), .ZN(new_n11712_));
  AOI21_X1   g11519(.A1(new_n11579_), .A2(new_n11712_), .B(new_n11590_), .ZN(new_n11713_));
  XOR2_X1    g11520(.A1(new_n11576_), .A2(new_n11544_), .Z(new_n11714_));
  AOI22_X1   g11521(.A1(\a[33] ), .A2(\a[55] ), .B1(\a[34] ), .B2(\a[54] ), .ZN(new_n11715_));
  NOR2_X1    g11522(.A1(new_n3932_), .A2(new_n6129_), .ZN(new_n11716_));
  NOR3_X1    g11523(.A1(new_n11716_), .A2(new_n4034_), .A3(new_n11715_), .ZN(new_n11717_));
  NOR2_X1    g11524(.A1(new_n11717_), .A2(new_n11716_), .ZN(new_n11718_));
  INV_X1     g11525(.I(new_n11718_), .ZN(new_n11719_));
  OAI22_X1   g11526(.A1(new_n11719_), .A2(new_n11715_), .B1(new_n4034_), .B2(new_n11717_), .ZN(new_n11720_));
  XNOR2_X1   g11527(.A1(new_n11720_), .A2(new_n11714_), .ZN(new_n11721_));
  XOR2_X1    g11528(.A1(new_n11713_), .A2(new_n11721_), .Z(new_n11722_));
  XNOR2_X1   g11529(.A1(new_n11722_), .A2(new_n11711_), .ZN(new_n11723_));
  NOR2_X1    g11530(.A1(new_n11642_), .A2(new_n11637_), .ZN(new_n11724_));
  NOR2_X1    g11531(.A1(new_n11669_), .A2(new_n11666_), .ZN(new_n11725_));
  XOR2_X1    g11532(.A1(new_n11724_), .A2(new_n11725_), .Z(new_n11726_));
  XNOR2_X1   g11533(.A1(new_n11726_), .A2(new_n11723_), .ZN(new_n11727_));
  NAND2_X1   g11534(.A1(new_n11626_), .A2(new_n11438_), .ZN(new_n11728_));
  NAND2_X1   g11535(.A1(new_n11728_), .A2(new_n11625_), .ZN(new_n11729_));
  AOI22_X1   g11536(.A1(\a[38] ), .A2(\a[50] ), .B1(\a[39] ), .B2(\a[49] ), .ZN(new_n11730_));
  INV_X1     g11537(.I(new_n11730_), .ZN(new_n11731_));
  NOR2_X1    g11538(.A1(new_n4210_), .A2(new_n5155_), .ZN(new_n11732_));
  NOR2_X1    g11539(.A1(new_n1814_), .A2(new_n6548_), .ZN(new_n11733_));
  AOI21_X1   g11540(.A1(new_n11731_), .A2(new_n11733_), .B(new_n11732_), .ZN(new_n11734_));
  NAND2_X1   g11541(.A1(new_n11734_), .A2(new_n11731_), .ZN(new_n11735_));
  OAI21_X1   g11542(.A1(new_n11732_), .A2(new_n11730_), .B(new_n11733_), .ZN(new_n11736_));
  NAND2_X1   g11543(.A1(new_n11735_), .A2(new_n11736_), .ZN(new_n11737_));
  AOI22_X1   g11544(.A1(\a[30] ), .A2(\a[58] ), .B1(\a[32] ), .B2(\a[56] ), .ZN(new_n11738_));
  NOR2_X1    g11545(.A1(new_n2202_), .A2(new_n6318_), .ZN(new_n11739_));
  OAI21_X1   g11546(.A1(new_n11739_), .A2(new_n11738_), .B(new_n5918_), .ZN(new_n11740_));
  INV_X1     g11547(.I(new_n11738_), .ZN(new_n11741_));
  AOI21_X1   g11548(.A1(new_n5918_), .A2(new_n11741_), .B(new_n11739_), .ZN(new_n11742_));
  INV_X1     g11549(.I(new_n11742_), .ZN(new_n11743_));
  OAI21_X1   g11550(.A1(new_n11743_), .A2(new_n11738_), .B(new_n11740_), .ZN(new_n11744_));
  XNOR2_X1   g11551(.A1(new_n11744_), .A2(new_n11737_), .ZN(new_n11745_));
  INV_X1     g11552(.I(new_n11745_), .ZN(new_n11746_));
  XOR2_X1    g11553(.A1(new_n11729_), .A2(new_n11746_), .Z(new_n11747_));
  AOI21_X1   g11554(.A1(\a[25] ), .A2(\a[63] ), .B(new_n11586_), .ZN(new_n11748_));
  NOR3_X1    g11555(.A1(new_n11585_), .A2(new_n1441_), .A3(new_n7643_), .ZN(new_n11749_));
  NOR2_X1    g11556(.A1(new_n11748_), .A2(new_n11749_), .ZN(new_n11750_));
  XOR2_X1    g11557(.A1(new_n11750_), .A2(new_n11613_), .Z(new_n11751_));
  AND2_X2    g11558(.A1(new_n11747_), .A2(new_n11751_), .Z(new_n11752_));
  NOR2_X1    g11559(.A1(new_n11747_), .A2(new_n11751_), .ZN(new_n11753_));
  NOR2_X1    g11560(.A1(new_n11752_), .A2(new_n11753_), .ZN(new_n11754_));
  NOR2_X1    g11561(.A1(new_n2189_), .A2(new_n7454_), .ZN(new_n11755_));
  NOR2_X1    g11562(.A1(new_n3341_), .A2(new_n7146_), .ZN(new_n11756_));
  NOR2_X1    g11563(.A1(new_n1972_), .A2(new_n7591_), .ZN(new_n11757_));
  NOR2_X1    g11564(.A1(new_n11756_), .A2(new_n11757_), .ZN(new_n11758_));
  NOR2_X1    g11565(.A1(new_n11758_), .A2(new_n11755_), .ZN(new_n11759_));
  NAND2_X1   g11566(.A1(\a[26] ), .A2(\a[62] ), .ZN(new_n11760_));
  AOI22_X1   g11567(.A1(\a[27] ), .A2(\a[61] ), .B1(\a[28] ), .B2(\a[60] ), .ZN(new_n11761_));
  NOR2_X1    g11568(.A1(new_n11759_), .A2(new_n11755_), .ZN(new_n11762_));
  INV_X1     g11569(.I(new_n11762_), .ZN(new_n11763_));
  OAI22_X1   g11570(.A1(new_n11763_), .A2(new_n11761_), .B1(new_n11759_), .B2(new_n11760_), .ZN(new_n11764_));
  AOI22_X1   g11571(.A1(\a[41] ), .A2(\a[47] ), .B1(\a[42] ), .B2(\a[46] ), .ZN(new_n11765_));
  INV_X1     g11572(.I(new_n11765_), .ZN(new_n11766_));
  NOR2_X1    g11573(.A1(new_n4667_), .A2(new_n4721_), .ZN(new_n11767_));
  NOR2_X1    g11574(.A1(new_n2051_), .A2(new_n6298_), .ZN(new_n11768_));
  AOI21_X1   g11575(.A1(new_n11766_), .A2(new_n11768_), .B(new_n11767_), .ZN(new_n11769_));
  NAND2_X1   g11576(.A1(new_n11769_), .A2(new_n11766_), .ZN(new_n11770_));
  OAI21_X1   g11577(.A1(new_n11767_), .A2(new_n11765_), .B(new_n11768_), .ZN(new_n11771_));
  NAND2_X1   g11578(.A1(new_n11770_), .A2(new_n11771_), .ZN(new_n11772_));
  XNOR2_X1   g11579(.A1(new_n11764_), .A2(new_n11772_), .ZN(new_n11773_));
  NAND2_X1   g11580(.A1(new_n4189_), .A2(new_n5682_), .ZN(new_n11774_));
  NAND2_X1   g11581(.A1(new_n3232_), .A2(new_n5862_), .ZN(new_n11775_));
  AOI22_X1   g11582(.A1(new_n11774_), .A2(new_n11775_), .B1(new_n3037_), .B2(new_n5524_), .ZN(new_n11776_));
  NAND2_X1   g11583(.A1(\a[35] ), .A2(\a[53] ), .ZN(new_n11777_));
  AOI22_X1   g11584(.A1(\a[36] ), .A2(\a[52] ), .B1(\a[37] ), .B2(\a[51] ), .ZN(new_n11778_));
  NAND2_X1   g11585(.A1(new_n3037_), .A2(new_n5524_), .ZN(new_n11779_));
  NAND3_X1   g11586(.A1(new_n11779_), .A2(new_n11774_), .A3(new_n11775_), .ZN(new_n11780_));
  OAI22_X1   g11587(.A1(new_n11776_), .A2(new_n11777_), .B1(new_n11780_), .B2(new_n11778_), .ZN(new_n11781_));
  XOR2_X1    g11588(.A1(new_n11773_), .A2(new_n11781_), .Z(new_n11782_));
  XOR2_X1    g11589(.A1(new_n11754_), .A2(new_n11782_), .Z(new_n11783_));
  NAND2_X1   g11590(.A1(new_n11656_), .A2(new_n11671_), .ZN(new_n11784_));
  NAND2_X1   g11591(.A1(new_n11672_), .A2(new_n11653_), .ZN(new_n11785_));
  NAND2_X1   g11592(.A1(new_n11785_), .A2(new_n11784_), .ZN(new_n11786_));
  XOR2_X1    g11593(.A1(new_n11786_), .A2(new_n11783_), .Z(new_n11787_));
  XOR2_X1    g11594(.A1(new_n11787_), .A2(new_n11727_), .Z(new_n11788_));
  XNOR2_X1   g11595(.A1(new_n11709_), .A2(new_n11788_), .ZN(new_n11789_));
  NAND2_X1   g11596(.A1(new_n11676_), .A2(new_n11673_), .ZN(new_n11790_));
  OAI21_X1   g11597(.A1(new_n11677_), .A2(new_n11651_), .B(new_n11790_), .ZN(new_n11791_));
  NOR2_X1    g11598(.A1(new_n11789_), .A2(new_n11791_), .ZN(new_n11792_));
  INV_X1     g11599(.I(new_n11792_), .ZN(new_n11793_));
  NAND2_X1   g11600(.A1(new_n11789_), .A2(new_n11791_), .ZN(new_n11794_));
  NAND2_X1   g11601(.A1(new_n11793_), .A2(new_n11794_), .ZN(new_n11795_));
  XOR2_X1    g11602(.A1(new_n11685_), .A2(new_n11795_), .Z(\asquared[89] ));
  OAI21_X1   g11603(.A1(new_n11684_), .A2(new_n11681_), .B(new_n11793_), .ZN(new_n11797_));
  NAND2_X1   g11604(.A1(new_n11797_), .A2(new_n11794_), .ZN(new_n11798_));
  OAI21_X1   g11605(.A1(new_n11706_), .A2(new_n11788_), .B(new_n11707_), .ZN(new_n11799_));
  INV_X1     g11606(.I(new_n11799_), .ZN(new_n11800_));
  AOI22_X1   g11607(.A1(\a[33] ), .A2(\a[56] ), .B1(\a[35] ), .B2(\a[54] ), .ZN(new_n11801_));
  INV_X1     g11608(.I(new_n11801_), .ZN(new_n11802_));
  NOR2_X1    g11609(.A1(new_n2526_), .A2(new_n6058_), .ZN(new_n11803_));
  NOR2_X1    g11610(.A1(new_n3327_), .A2(new_n4596_), .ZN(new_n11804_));
  AOI21_X1   g11611(.A1(new_n11802_), .A2(new_n11804_), .B(new_n11803_), .ZN(new_n11805_));
  INV_X1     g11612(.I(new_n11805_), .ZN(new_n11806_));
  OAI21_X1   g11613(.A1(new_n11803_), .A2(new_n11801_), .B(new_n11804_), .ZN(new_n11807_));
  OAI21_X1   g11614(.A1(new_n11806_), .A2(new_n11801_), .B(new_n11807_), .ZN(new_n11808_));
  NOR2_X1    g11615(.A1(new_n6140_), .A2(new_n5525_), .ZN(new_n11809_));
  NOR2_X1    g11616(.A1(new_n2916_), .A2(new_n5683_), .ZN(new_n11810_));
  NOR2_X1    g11617(.A1(new_n3038_), .A2(new_n6563_), .ZN(new_n11811_));
  NOR2_X1    g11618(.A1(new_n11810_), .A2(new_n11811_), .ZN(new_n11812_));
  NOR2_X1    g11619(.A1(new_n11812_), .A2(new_n11809_), .ZN(new_n11813_));
  NAND2_X1   g11620(.A1(\a[36] ), .A2(\a[53] ), .ZN(new_n11814_));
  AOI22_X1   g11621(.A1(\a[37] ), .A2(\a[52] ), .B1(\a[38] ), .B2(\a[51] ), .ZN(new_n11815_));
  NOR2_X1    g11622(.A1(new_n11813_), .A2(new_n11809_), .ZN(new_n11816_));
  INV_X1     g11623(.I(new_n11816_), .ZN(new_n11817_));
  OAI22_X1   g11624(.A1(new_n11817_), .A2(new_n11815_), .B1(new_n11813_), .B2(new_n11814_), .ZN(new_n11818_));
  XOR2_X1    g11625(.A1(new_n11818_), .A2(new_n11808_), .Z(new_n11819_));
  NAND2_X1   g11626(.A1(new_n2201_), .A2(new_n7203_), .ZN(new_n11820_));
  NAND2_X1   g11627(.A1(new_n2437_), .A2(new_n7205_), .ZN(new_n11821_));
  AOI22_X1   g11628(.A1(new_n11820_), .A2(new_n11821_), .B1(new_n3210_), .B2(new_n6803_), .ZN(new_n11822_));
  NAND2_X1   g11629(.A1(\a[30] ), .A2(\a[59] ), .ZN(new_n11823_));
  AOI22_X1   g11630(.A1(\a[31] ), .A2(\a[58] ), .B1(\a[32] ), .B2(\a[57] ), .ZN(new_n11824_));
  NAND2_X1   g11631(.A1(new_n3210_), .A2(new_n6803_), .ZN(new_n11825_));
  NAND3_X1   g11632(.A1(new_n11825_), .A2(new_n11820_), .A3(new_n11821_), .ZN(new_n11826_));
  OAI22_X1   g11633(.A1(new_n11822_), .A2(new_n11823_), .B1(new_n11826_), .B2(new_n11824_), .ZN(new_n11827_));
  XOR2_X1    g11634(.A1(new_n11819_), .A2(new_n11827_), .Z(new_n11828_));
  XNOR2_X1   g11635(.A1(new_n11762_), .A2(new_n11780_), .ZN(new_n11829_));
  XOR2_X1    g11636(.A1(new_n11829_), .A2(new_n11743_), .Z(new_n11830_));
  NOR2_X1    g11637(.A1(new_n2679_), .A2(new_n7454_), .ZN(new_n11831_));
  INV_X1     g11638(.I(new_n11831_), .ZN(new_n11832_));
  NOR2_X1    g11639(.A1(new_n1814_), .A2(new_n6723_), .ZN(new_n11833_));
  NOR2_X1    g11640(.A1(new_n1718_), .A2(new_n6897_), .ZN(new_n11834_));
  OAI21_X1   g11641(.A1(new_n11833_), .A2(new_n11834_), .B(new_n11832_), .ZN(new_n11835_));
  XNOR2_X1   g11642(.A1(new_n11835_), .A2(new_n11718_), .ZN(new_n11836_));
  NOR3_X1    g11643(.A1(new_n1750_), .A2(new_n4030_), .A3(new_n7144_), .ZN(new_n11837_));
  NAND2_X1   g11644(.A1(new_n11837_), .A2(new_n4703_), .ZN(new_n11838_));
  AOI21_X1   g11645(.A1(\a[27] ), .A2(\a[62] ), .B(\a[45] ), .ZN(new_n11839_));
  NOR2_X1    g11646(.A1(new_n11837_), .A2(new_n4703_), .ZN(new_n11840_));
  INV_X1     g11647(.I(new_n11840_), .ZN(new_n11841_));
  OAI21_X1   g11648(.A1(new_n11841_), .A2(new_n11839_), .B(new_n11838_), .ZN(new_n11842_));
  AOI22_X1   g11649(.A1(\a[42] ), .A2(\a[47] ), .B1(\a[43] ), .B2(\a[46] ), .ZN(new_n11843_));
  NOR2_X1    g11650(.A1(new_n2442_), .A2(new_n5680_), .ZN(new_n11844_));
  INV_X1     g11651(.I(new_n11844_), .ZN(new_n11845_));
  OAI22_X1   g11652(.A1(new_n4181_), .A2(new_n4721_), .B1(new_n11845_), .B2(new_n11843_), .ZN(new_n11846_));
  NOR2_X1    g11653(.A1(new_n4181_), .A2(new_n4721_), .ZN(new_n11847_));
  OAI21_X1   g11654(.A1(new_n11847_), .A2(new_n11843_), .B(new_n11844_), .ZN(new_n11848_));
  OAI21_X1   g11655(.A1(new_n11846_), .A2(new_n11843_), .B(new_n11848_), .ZN(new_n11849_));
  XOR2_X1    g11656(.A1(new_n11849_), .A2(new_n11842_), .Z(new_n11850_));
  XOR2_X1    g11657(.A1(new_n11850_), .A2(new_n11836_), .Z(new_n11851_));
  XNOR2_X1   g11658(.A1(new_n11830_), .A2(new_n11851_), .ZN(new_n11852_));
  XNOR2_X1   g11659(.A1(new_n11852_), .A2(new_n11828_), .ZN(new_n11853_));
  NAND2_X1   g11660(.A1(new_n11700_), .A2(new_n11703_), .ZN(new_n11854_));
  NAND2_X1   g11661(.A1(new_n11704_), .A2(new_n11690_), .ZN(new_n11855_));
  NAND2_X1   g11662(.A1(new_n11855_), .A2(new_n11854_), .ZN(new_n11856_));
  XOR2_X1    g11663(.A1(new_n11856_), .A2(new_n11853_), .Z(new_n11857_));
  NAND2_X1   g11664(.A1(new_n11722_), .A2(new_n11711_), .ZN(new_n11858_));
  OAI21_X1   g11665(.A1(new_n11713_), .A2(new_n11721_), .B(new_n11858_), .ZN(new_n11859_));
  NOR2_X1    g11666(.A1(new_n11694_), .A2(new_n11695_), .ZN(new_n11860_));
  NOR2_X1    g11667(.A1(new_n11698_), .A2(new_n11860_), .ZN(new_n11861_));
  NAND2_X1   g11668(.A1(new_n11576_), .A2(new_n11544_), .ZN(new_n11862_));
  NOR2_X1    g11669(.A1(new_n11576_), .A2(new_n11544_), .ZN(new_n11863_));
  AOI21_X1   g11670(.A1(new_n11720_), .A2(new_n11862_), .B(new_n11863_), .ZN(new_n11864_));
  INV_X1     g11671(.I(new_n11864_), .ZN(new_n11865_));
  NAND2_X1   g11672(.A1(new_n11558_), .A2(new_n11599_), .ZN(new_n11866_));
  NAND2_X1   g11673(.A1(new_n11710_), .A2(new_n11606_), .ZN(new_n11867_));
  NAND2_X1   g11674(.A1(new_n11867_), .A2(new_n11866_), .ZN(new_n11868_));
  INV_X1     g11675(.I(new_n11749_), .ZN(new_n11869_));
  NAND2_X1   g11676(.A1(new_n11750_), .A2(new_n11613_), .ZN(new_n11870_));
  NAND2_X1   g11677(.A1(new_n11870_), .A2(new_n11869_), .ZN(new_n11871_));
  XOR2_X1    g11678(.A1(new_n11868_), .A2(new_n11871_), .Z(new_n11872_));
  XOR2_X1    g11679(.A1(new_n11872_), .A2(new_n11865_), .Z(new_n11873_));
  INV_X1     g11680(.I(new_n11873_), .ZN(new_n11874_));
  XOR2_X1    g11681(.A1(new_n11861_), .A2(new_n11874_), .Z(new_n11875_));
  NOR2_X1    g11682(.A1(new_n11875_), .A2(new_n11859_), .ZN(new_n11876_));
  NAND2_X1   g11683(.A1(new_n11875_), .A2(new_n11859_), .ZN(new_n11877_));
  INV_X1     g11684(.I(new_n11877_), .ZN(new_n11878_));
  NOR2_X1    g11685(.A1(new_n11878_), .A2(new_n11876_), .ZN(new_n11879_));
  XOR2_X1    g11686(.A1(new_n11857_), .A2(new_n11879_), .Z(new_n11880_));
  INV_X1     g11687(.I(new_n11880_), .ZN(new_n11881_));
  INV_X1     g11688(.I(new_n11727_), .ZN(new_n11882_));
  INV_X1     g11689(.I(new_n11783_), .ZN(new_n11883_));
  NAND2_X1   g11690(.A1(new_n11786_), .A2(new_n11883_), .ZN(new_n11884_));
  OAI21_X1   g11691(.A1(new_n11787_), .A2(new_n11882_), .B(new_n11884_), .ZN(new_n11885_));
  NOR2_X1    g11692(.A1(new_n11724_), .A2(new_n11725_), .ZN(new_n11886_));
  INV_X1     g11693(.I(new_n11726_), .ZN(new_n11887_));
  NOR2_X1    g11694(.A1(new_n11887_), .A2(new_n11723_), .ZN(new_n11888_));
  NOR2_X1    g11695(.A1(new_n11888_), .A2(new_n11886_), .ZN(new_n11889_));
  NOR3_X1    g11696(.A1(new_n11752_), .A2(new_n11753_), .A3(new_n11782_), .ZN(new_n11890_));
  NOR2_X1    g11697(.A1(new_n11890_), .A2(new_n11752_), .ZN(new_n11891_));
  XOR2_X1    g11698(.A1(new_n11734_), .A2(new_n11769_), .Z(new_n11892_));
  AOI22_X1   g11699(.A1(\a[39] ), .A2(\a[50] ), .B1(\a[40] ), .B2(\a[49] ), .ZN(new_n11893_));
  NOR2_X1    g11700(.A1(new_n1566_), .A2(new_n7643_), .ZN(new_n11894_));
  INV_X1     g11701(.I(new_n11894_), .ZN(new_n11895_));
  NOR2_X1    g11702(.A1(new_n3551_), .A2(new_n5155_), .ZN(new_n11896_));
  NOR3_X1    g11703(.A1(new_n11896_), .A2(new_n11893_), .A3(new_n11895_), .ZN(new_n11897_));
  NOR2_X1    g11704(.A1(new_n11897_), .A2(new_n11896_), .ZN(new_n11898_));
  INV_X1     g11705(.I(new_n11898_), .ZN(new_n11899_));
  OAI22_X1   g11706(.A1(new_n11899_), .A2(new_n11893_), .B1(new_n11895_), .B2(new_n11897_), .ZN(new_n11900_));
  XNOR2_X1   g11707(.A1(new_n11900_), .A2(new_n11892_), .ZN(new_n11901_));
  INV_X1     g11708(.I(new_n11901_), .ZN(new_n11902_));
  NAND2_X1   g11709(.A1(new_n11744_), .A2(new_n11737_), .ZN(new_n11903_));
  NAND2_X1   g11710(.A1(new_n11729_), .A2(new_n11746_), .ZN(new_n11904_));
  NAND2_X1   g11711(.A1(new_n11904_), .A2(new_n11903_), .ZN(new_n11905_));
  NAND2_X1   g11712(.A1(new_n11764_), .A2(new_n11772_), .ZN(new_n11906_));
  INV_X1     g11713(.I(new_n11773_), .ZN(new_n11907_));
  NAND2_X1   g11714(.A1(new_n11907_), .A2(new_n11781_), .ZN(new_n11908_));
  NAND2_X1   g11715(.A1(new_n11908_), .A2(new_n11906_), .ZN(new_n11909_));
  XOR2_X1    g11716(.A1(new_n11909_), .A2(new_n11905_), .Z(new_n11910_));
  XOR2_X1    g11717(.A1(new_n11910_), .A2(new_n11902_), .Z(new_n11911_));
  XOR2_X1    g11718(.A1(new_n11911_), .A2(new_n11891_), .Z(new_n11912_));
  XOR2_X1    g11719(.A1(new_n11889_), .A2(new_n11912_), .Z(new_n11913_));
  NAND2_X1   g11720(.A1(new_n11885_), .A2(new_n11913_), .ZN(new_n11914_));
  NAND2_X1   g11721(.A1(new_n11914_), .A2(new_n11885_), .ZN(new_n11915_));
  NAND2_X1   g11722(.A1(new_n11914_), .A2(new_n11913_), .ZN(new_n11916_));
  NAND2_X1   g11723(.A1(new_n11915_), .A2(new_n11916_), .ZN(new_n11917_));
  NAND2_X1   g11724(.A1(new_n11917_), .A2(new_n11881_), .ZN(new_n11918_));
  NAND3_X1   g11725(.A1(new_n11915_), .A2(new_n11916_), .A3(new_n11880_), .ZN(new_n11919_));
  NAND2_X1   g11726(.A1(new_n11918_), .A2(new_n11919_), .ZN(new_n11920_));
  NOR2_X1    g11727(.A1(new_n11920_), .A2(new_n11800_), .ZN(new_n11921_));
  NAND2_X1   g11728(.A1(new_n11920_), .A2(new_n11800_), .ZN(new_n11922_));
  INV_X1     g11729(.I(new_n11922_), .ZN(new_n11923_));
  NOR2_X1    g11730(.A1(new_n11923_), .A2(new_n11921_), .ZN(new_n11924_));
  XOR2_X1    g11731(.A1(new_n11798_), .A2(new_n11924_), .Z(\asquared[90] ));
  AOI21_X1   g11732(.A1(new_n11797_), .A2(new_n11794_), .B(new_n11923_), .ZN(new_n11926_));
  NOR2_X1    g11733(.A1(new_n11926_), .A2(new_n11921_), .ZN(new_n11927_));
  NAND2_X1   g11734(.A1(new_n11918_), .A2(new_n11914_), .ZN(new_n11928_));
  INV_X1     g11735(.I(new_n11911_), .ZN(new_n11929_));
  NOR2_X1    g11736(.A1(new_n11929_), .A2(new_n11891_), .ZN(new_n11930_));
  NOR2_X1    g11737(.A1(new_n11889_), .A2(new_n11912_), .ZN(new_n11931_));
  NOR2_X1    g11738(.A1(new_n11931_), .A2(new_n11930_), .ZN(new_n11932_));
  NAND2_X1   g11739(.A1(new_n3577_), .A2(new_n6494_), .ZN(new_n11933_));
  OAI22_X1   g11740(.A1(new_n2526_), .A2(new_n8952_), .B1(new_n2746_), .B2(new_n7185_), .ZN(new_n11934_));
  NAND2_X1   g11741(.A1(new_n11934_), .A2(new_n11933_), .ZN(new_n11935_));
  NAND3_X1   g11742(.A1(new_n11935_), .A2(\a[35] ), .A3(\a[55] ), .ZN(new_n11936_));
  AOI22_X1   g11743(.A1(\a[33] ), .A2(\a[57] ), .B1(\a[34] ), .B2(\a[56] ), .ZN(new_n11937_));
  NAND2_X1   g11744(.A1(new_n11935_), .A2(new_n11933_), .ZN(new_n11938_));
  OAI21_X1   g11745(.A1(new_n11937_), .A2(new_n11938_), .B(new_n11936_), .ZN(new_n11939_));
  NOR2_X1    g11746(.A1(new_n6140_), .A2(new_n6563_), .ZN(new_n11940_));
  NOR2_X1    g11747(.A1(new_n3038_), .A2(new_n6127_), .ZN(new_n11941_));
  NOR2_X1    g11748(.A1(new_n2916_), .A2(new_n8421_), .ZN(new_n11942_));
  NOR2_X1    g11749(.A1(new_n11941_), .A2(new_n11942_), .ZN(new_n11943_));
  NOR2_X1    g11750(.A1(new_n11943_), .A2(new_n11940_), .ZN(new_n11944_));
  NOR3_X1    g11751(.A1(new_n11944_), .A2(new_n2626_), .A3(new_n5617_), .ZN(new_n11945_));
  AOI22_X1   g11752(.A1(\a[37] ), .A2(\a[53] ), .B1(\a[38] ), .B2(\a[52] ), .ZN(new_n11946_));
  NOR3_X1    g11753(.A1(new_n11944_), .A2(new_n11940_), .A3(new_n11946_), .ZN(new_n11947_));
  NOR2_X1    g11754(.A1(new_n11947_), .A2(new_n11945_), .ZN(new_n11948_));
  XOR2_X1    g11755(.A1(new_n11948_), .A2(new_n11939_), .Z(new_n11949_));
  NAND2_X1   g11756(.A1(new_n4180_), .A2(new_n4976_), .ZN(new_n11950_));
  NAND2_X1   g11757(.A1(new_n3860_), .A2(new_n6743_), .ZN(new_n11951_));
  AOI22_X1   g11758(.A1(new_n11950_), .A2(new_n11951_), .B1(new_n4342_), .B2(new_n4720_), .ZN(new_n11952_));
  NAND2_X1   g11759(.A1(new_n4342_), .A2(new_n4720_), .ZN(new_n11953_));
  NAND3_X1   g11760(.A1(new_n11953_), .A2(new_n11950_), .A3(new_n11951_), .ZN(new_n11954_));
  AOI21_X1   g11761(.A1(\a[43] ), .A2(\a[47] ), .B(new_n6100_), .ZN(new_n11955_));
  NAND2_X1   g11762(.A1(\a[42] ), .A2(\a[48] ), .ZN(new_n11956_));
  OAI22_X1   g11763(.A1(new_n11952_), .A2(new_n11956_), .B1(new_n11954_), .B2(new_n11955_), .ZN(new_n11957_));
  XOR2_X1    g11764(.A1(new_n11949_), .A2(new_n11957_), .Z(new_n11958_));
  INV_X1     g11765(.I(new_n11958_), .ZN(new_n11959_));
  NAND2_X1   g11766(.A1(new_n11868_), .A2(new_n11871_), .ZN(new_n11960_));
  NAND2_X1   g11767(.A1(new_n11872_), .A2(new_n11865_), .ZN(new_n11961_));
  NAND2_X1   g11768(.A1(new_n11961_), .A2(new_n11960_), .ZN(new_n11962_));
  XNOR2_X1   g11769(.A1(new_n11816_), .A2(new_n11826_), .ZN(new_n11963_));
  XOR2_X1    g11770(.A1(new_n11963_), .A2(new_n11899_), .Z(new_n11964_));
  XOR2_X1    g11771(.A1(new_n11962_), .A2(new_n11964_), .Z(new_n11965_));
  XOR2_X1    g11772(.A1(new_n11965_), .A2(new_n11959_), .Z(new_n11966_));
  XOR2_X1    g11773(.A1(new_n11932_), .A2(new_n11966_), .Z(new_n11967_));
  NAND2_X1   g11774(.A1(new_n11909_), .A2(new_n11905_), .ZN(new_n11968_));
  NAND2_X1   g11775(.A1(new_n11910_), .A2(new_n11902_), .ZN(new_n11969_));
  NAND2_X1   g11776(.A1(new_n11969_), .A2(new_n11968_), .ZN(new_n11970_));
  NOR2_X1    g11777(.A1(new_n2679_), .A2(new_n7591_), .ZN(new_n11971_));
  AOI22_X1   g11778(.A1(new_n1815_), .A2(new_n7852_), .B1(new_n2103_), .B2(new_n7644_), .ZN(new_n11972_));
  NOR2_X1    g11779(.A1(new_n11971_), .A2(new_n11972_), .ZN(new_n11973_));
  NAND2_X1   g11780(.A1(\a[27] ), .A2(\a[63] ), .ZN(new_n11974_));
  AOI22_X1   g11781(.A1(\a[28] ), .A2(\a[62] ), .B1(\a[29] ), .B2(\a[61] ), .ZN(new_n11975_));
  NOR2_X1    g11782(.A1(new_n11973_), .A2(new_n11971_), .ZN(new_n11976_));
  INV_X1     g11783(.I(new_n11976_), .ZN(new_n11977_));
  OAI22_X1   g11784(.A1(new_n11977_), .A2(new_n11975_), .B1(new_n11973_), .B2(new_n11974_), .ZN(new_n11978_));
  OAI21_X1   g11785(.A1(new_n11835_), .A2(new_n11718_), .B(new_n11832_), .ZN(new_n11979_));
  INV_X1     g11786(.I(new_n11979_), .ZN(new_n11980_));
  NOR2_X1    g11787(.A1(new_n3833_), .A2(new_n7206_), .ZN(new_n11981_));
  AOI22_X1   g11788(.A1(\a[31] ), .A2(\a[59] ), .B1(\a[32] ), .B2(\a[58] ), .ZN(new_n11982_));
  OAI22_X1   g11789(.A1(new_n11981_), .A2(new_n11982_), .B1(new_n2030_), .B2(new_n6723_), .ZN(new_n11983_));
  OAI22_X1   g11790(.A1(new_n2202_), .A2(new_n7801_), .B1(new_n2438_), .B2(new_n7452_), .ZN(new_n11984_));
  OAI21_X1   g11791(.A1(new_n3833_), .A2(new_n7206_), .B(new_n11984_), .ZN(new_n11985_));
  NAND2_X1   g11792(.A1(new_n11985_), .A2(new_n11983_), .ZN(new_n11986_));
  NOR2_X1    g11793(.A1(new_n11980_), .A2(new_n11986_), .ZN(new_n11987_));
  NOR2_X1    g11794(.A1(new_n11987_), .A2(new_n11980_), .ZN(new_n11988_));
  NOR2_X1    g11795(.A1(new_n11979_), .A2(new_n11986_), .ZN(new_n11989_));
  OAI21_X1   g11796(.A1(new_n11988_), .A2(new_n11989_), .B(new_n11978_), .ZN(new_n11990_));
  INV_X1     g11797(.I(new_n11990_), .ZN(new_n11991_));
  NOR3_X1    g11798(.A1(new_n11988_), .A2(new_n11978_), .A3(new_n11989_), .ZN(new_n11992_));
  NOR2_X1    g11799(.A1(new_n11991_), .A2(new_n11992_), .ZN(new_n11993_));
  NAND2_X1   g11800(.A1(new_n11900_), .A2(new_n11892_), .ZN(new_n11994_));
  OAI21_X1   g11801(.A1(new_n11734_), .A2(new_n11769_), .B(new_n11994_), .ZN(new_n11995_));
  INV_X1     g11802(.I(new_n11995_), .ZN(new_n11996_));
  INV_X1     g11803(.I(new_n6114_), .ZN(new_n11997_));
  NOR2_X1    g11804(.A1(new_n5377_), .A2(new_n5155_), .ZN(new_n11998_));
  AOI22_X1   g11805(.A1(new_n3328_), .A2(new_n7867_), .B1(new_n3550_), .B2(new_n5439_), .ZN(new_n11999_));
  NOR2_X1    g11806(.A1(new_n11998_), .A2(new_n11999_), .ZN(new_n12000_));
  AOI22_X1   g11807(.A1(\a[40] ), .A2(\a[50] ), .B1(\a[41] ), .B2(\a[49] ), .ZN(new_n12001_));
  NOR2_X1    g11808(.A1(new_n12000_), .A2(new_n11998_), .ZN(new_n12002_));
  INV_X1     g11809(.I(new_n12002_), .ZN(new_n12003_));
  OAI22_X1   g11810(.A1(new_n12003_), .A2(new_n12001_), .B1(new_n11997_), .B2(new_n12000_), .ZN(new_n12004_));
  NAND2_X1   g11811(.A1(new_n11763_), .A2(new_n11780_), .ZN(new_n12005_));
  NAND2_X1   g11812(.A1(new_n11829_), .A2(new_n11743_), .ZN(new_n12006_));
  NAND2_X1   g11813(.A1(new_n12006_), .A2(new_n12005_), .ZN(new_n12007_));
  XNOR2_X1   g11814(.A1(new_n12007_), .A2(new_n12004_), .ZN(new_n12008_));
  XOR2_X1    g11815(.A1(new_n12008_), .A2(new_n11996_), .Z(new_n12009_));
  XOR2_X1    g11816(.A1(new_n12009_), .A2(new_n11993_), .Z(new_n12010_));
  XNOR2_X1   g11817(.A1(new_n12010_), .A2(new_n11970_), .ZN(new_n12011_));
  XNOR2_X1   g11818(.A1(new_n11967_), .A2(new_n12011_), .ZN(new_n12012_));
  INV_X1     g11819(.I(new_n12012_), .ZN(new_n12013_));
  INV_X1     g11820(.I(new_n11853_), .ZN(new_n12014_));
  NAND2_X1   g11821(.A1(new_n11856_), .A2(new_n12014_), .ZN(new_n12015_));
  INV_X1     g11822(.I(new_n11857_), .ZN(new_n12016_));
  NAND2_X1   g11823(.A1(new_n12016_), .A2(new_n11879_), .ZN(new_n12017_));
  NAND2_X1   g11824(.A1(new_n12017_), .A2(new_n12015_), .ZN(new_n12018_));
  NOR2_X1    g11825(.A1(new_n11861_), .A2(new_n11874_), .ZN(new_n12019_));
  NOR2_X1    g11826(.A1(new_n11878_), .A2(new_n12019_), .ZN(new_n12020_));
  INV_X1     g11827(.I(new_n12020_), .ZN(new_n12021_));
  INV_X1     g11828(.I(new_n11830_), .ZN(new_n12022_));
  NAND2_X1   g11829(.A1(new_n11852_), .A2(new_n11828_), .ZN(new_n12023_));
  OAI21_X1   g11830(.A1(new_n12022_), .A2(new_n11851_), .B(new_n12023_), .ZN(new_n12024_));
  XOR2_X1    g11831(.A1(new_n11846_), .A2(new_n11841_), .Z(new_n12025_));
  OR2_X2     g11832(.A1(new_n12025_), .A2(new_n11806_), .Z(new_n12026_));
  NAND2_X1   g11833(.A1(new_n12025_), .A2(new_n11806_), .ZN(new_n12027_));
  AND2_X2    g11834(.A1(new_n12026_), .A2(new_n12027_), .Z(new_n12028_));
  NAND2_X1   g11835(.A1(new_n11849_), .A2(new_n11842_), .ZN(new_n12029_));
  INV_X1     g11836(.I(new_n11836_), .ZN(new_n12030_));
  NAND2_X1   g11837(.A1(new_n12030_), .A2(new_n11850_), .ZN(new_n12031_));
  NAND2_X1   g11838(.A1(new_n12031_), .A2(new_n12029_), .ZN(new_n12032_));
  NAND2_X1   g11839(.A1(new_n11818_), .A2(new_n11808_), .ZN(new_n12033_));
  NAND2_X1   g11840(.A1(new_n11819_), .A2(new_n11827_), .ZN(new_n12034_));
  NAND2_X1   g11841(.A1(new_n12034_), .A2(new_n12033_), .ZN(new_n12035_));
  XOR2_X1    g11842(.A1(new_n12035_), .A2(new_n12032_), .Z(new_n12036_));
  XOR2_X1    g11843(.A1(new_n12036_), .A2(new_n12028_), .Z(new_n12037_));
  NOR2_X1    g11844(.A1(new_n12037_), .A2(new_n12024_), .ZN(new_n12038_));
  NAND2_X1   g11845(.A1(new_n12037_), .A2(new_n12024_), .ZN(new_n12039_));
  INV_X1     g11846(.I(new_n12039_), .ZN(new_n12040_));
  NOR2_X1    g11847(.A1(new_n12040_), .A2(new_n12038_), .ZN(new_n12041_));
  NOR2_X1    g11848(.A1(new_n12021_), .A2(new_n12041_), .ZN(new_n12042_));
  NAND2_X1   g11849(.A1(new_n12021_), .A2(new_n12041_), .ZN(new_n12043_));
  INV_X1     g11850(.I(new_n12043_), .ZN(new_n12044_));
  NOR2_X1    g11851(.A1(new_n12044_), .A2(new_n12042_), .ZN(new_n12045_));
  XOR2_X1    g11852(.A1(new_n12018_), .A2(new_n12045_), .Z(new_n12046_));
  XOR2_X1    g11853(.A1(new_n12046_), .A2(new_n12013_), .Z(new_n12047_));
  NAND2_X1   g11854(.A1(new_n12047_), .A2(new_n11928_), .ZN(new_n12048_));
  NOR2_X1    g11855(.A1(new_n12047_), .A2(new_n11928_), .ZN(new_n12049_));
  INV_X1     g11856(.I(new_n12049_), .ZN(new_n12050_));
  NAND2_X1   g11857(.A1(new_n12050_), .A2(new_n12048_), .ZN(new_n12051_));
  INV_X1     g11858(.I(new_n11921_), .ZN(new_n12052_));
  INV_X1     g11859(.I(new_n11794_), .ZN(new_n12053_));
  INV_X1     g11860(.I(new_n11514_), .ZN(new_n12054_));
  INV_X1     g11861(.I(new_n11679_), .ZN(new_n12055_));
  OAI21_X1   g11862(.A1(new_n11530_), .A2(new_n12054_), .B(new_n12055_), .ZN(new_n12056_));
  AOI21_X1   g11863(.A1(new_n12056_), .A2(new_n11680_), .B(new_n11792_), .ZN(new_n12057_));
  OAI21_X1   g11864(.A1(new_n12057_), .A2(new_n12053_), .B(new_n11922_), .ZN(new_n12058_));
  AOI21_X1   g11865(.A1(new_n12058_), .A2(new_n12052_), .B(new_n12049_), .ZN(new_n12059_));
  AOI22_X1   g11866(.A1(new_n12059_), .A2(new_n12048_), .B1(new_n11927_), .B2(new_n12051_), .ZN(\asquared[91] ));
  OAI21_X1   g11867(.A1(new_n11926_), .A2(new_n11921_), .B(new_n12050_), .ZN(new_n12061_));
  NAND2_X1   g11868(.A1(new_n12061_), .A2(new_n12048_), .ZN(new_n12062_));
  NAND2_X1   g11869(.A1(new_n12018_), .A2(new_n12045_), .ZN(new_n12063_));
  NAND2_X1   g11870(.A1(new_n12046_), .A2(new_n12013_), .ZN(new_n12064_));
  NAND2_X1   g11871(.A1(new_n12064_), .A2(new_n12063_), .ZN(new_n12065_));
  NOR2_X1    g11872(.A1(new_n12044_), .A2(new_n12040_), .ZN(new_n12066_));
  AOI22_X1   g11873(.A1(\a[40] ), .A2(\a[51] ), .B1(\a[41] ), .B2(\a[50] ), .ZN(new_n12067_));
  INV_X1     g11874(.I(new_n12067_), .ZN(new_n12068_));
  NOR2_X1    g11875(.A1(new_n5377_), .A2(new_n5440_), .ZN(new_n12069_));
  NOR2_X1    g11876(.A1(new_n1718_), .A2(new_n7643_), .ZN(new_n12070_));
  AOI21_X1   g11877(.A1(new_n12068_), .A2(new_n12070_), .B(new_n12069_), .ZN(new_n12071_));
  INV_X1     g11878(.I(new_n12071_), .ZN(new_n12072_));
  OAI21_X1   g11879(.A1(new_n12069_), .A2(new_n12067_), .B(new_n12070_), .ZN(new_n12073_));
  OAI21_X1   g11880(.A1(new_n12072_), .A2(new_n12067_), .B(new_n12073_), .ZN(new_n12074_));
  AOI22_X1   g11881(.A1(\a[43] ), .A2(\a[48] ), .B1(\a[44] ), .B2(\a[47] ), .ZN(new_n12075_));
  INV_X1     g11882(.I(new_n12075_), .ZN(new_n12076_));
  NOR2_X1    g11883(.A1(new_n4343_), .A2(new_n4977_), .ZN(new_n12077_));
  NOR2_X1    g11884(.A1(new_n2524_), .A2(new_n5856_), .ZN(new_n12078_));
  AOI21_X1   g11885(.A1(new_n12076_), .A2(new_n12078_), .B(new_n12077_), .ZN(new_n12079_));
  INV_X1     g11886(.I(new_n12079_), .ZN(new_n12080_));
  OAI21_X1   g11887(.A1(new_n12077_), .A2(new_n12075_), .B(new_n12078_), .ZN(new_n12081_));
  OAI21_X1   g11888(.A1(new_n12080_), .A2(new_n12075_), .B(new_n12081_), .ZN(new_n12082_));
  XOR2_X1    g11889(.A1(new_n12074_), .A2(new_n12082_), .Z(new_n12083_));
  NOR3_X1    g11890(.A1(new_n1814_), .A2(new_n4178_), .A3(new_n7144_), .ZN(new_n12084_));
  NAND2_X1   g11891(.A1(new_n12084_), .A2(new_n4429_), .ZN(new_n12085_));
  AOI21_X1   g11892(.A1(\a[29] ), .A2(\a[62] ), .B(\a[46] ), .ZN(new_n12086_));
  OR2_X2     g11893(.A1(new_n12084_), .A2(new_n4429_), .Z(new_n12087_));
  OAI21_X1   g11894(.A1(new_n12087_), .A2(new_n12086_), .B(new_n12085_), .ZN(new_n12088_));
  XNOR2_X1   g11895(.A1(new_n12083_), .A2(new_n12088_), .ZN(new_n12089_));
  INV_X1     g11896(.I(new_n12089_), .ZN(new_n12090_));
  NAND2_X1   g11897(.A1(new_n12007_), .A2(new_n12004_), .ZN(new_n12091_));
  OAI21_X1   g11898(.A1(new_n12008_), .A2(new_n11996_), .B(new_n12091_), .ZN(new_n12092_));
  NOR2_X1    g11899(.A1(new_n11984_), .A2(new_n11981_), .ZN(new_n12093_));
  NOR2_X1    g11900(.A1(new_n11944_), .A2(new_n11940_), .ZN(new_n12094_));
  XOR2_X1    g11901(.A1(new_n12094_), .A2(new_n11976_), .Z(new_n12095_));
  XNOR2_X1   g11902(.A1(new_n12095_), .A2(new_n12093_), .ZN(new_n12096_));
  NOR2_X1    g11903(.A1(new_n12092_), .A2(new_n12096_), .ZN(new_n12097_));
  NAND2_X1   g11904(.A1(new_n12092_), .A2(new_n12096_), .ZN(new_n12098_));
  INV_X1     g11905(.I(new_n12098_), .ZN(new_n12099_));
  NOR2_X1    g11906(.A1(new_n12099_), .A2(new_n12097_), .ZN(new_n12100_));
  NOR2_X1    g11907(.A1(new_n12100_), .A2(new_n12090_), .ZN(new_n12101_));
  NAND2_X1   g11908(.A1(new_n12100_), .A2(new_n12090_), .ZN(new_n12102_));
  INV_X1     g11909(.I(new_n12102_), .ZN(new_n12103_));
  NOR2_X1    g11910(.A1(new_n12103_), .A2(new_n12101_), .ZN(new_n12104_));
  INV_X1     g11911(.I(new_n12104_), .ZN(new_n12105_));
  XOR2_X1    g11912(.A1(new_n12066_), .A2(new_n12105_), .Z(new_n12106_));
  NAND2_X1   g11913(.A1(new_n11817_), .A2(new_n11826_), .ZN(new_n12107_));
  NAND2_X1   g11914(.A1(new_n11963_), .A2(new_n11899_), .ZN(new_n12108_));
  NAND2_X1   g11915(.A1(new_n12108_), .A2(new_n12107_), .ZN(new_n12109_));
  AOI22_X1   g11916(.A1(\a[34] ), .A2(\a[57] ), .B1(\a[36] ), .B2(\a[55] ), .ZN(new_n12110_));
  NOR2_X1    g11917(.A1(new_n5564_), .A2(new_n8952_), .ZN(new_n12111_));
  NOR3_X1    g11918(.A1(new_n12111_), .A2(new_n6338_), .A3(new_n12110_), .ZN(new_n12112_));
  NOR2_X1    g11919(.A1(new_n12112_), .A2(new_n12111_), .ZN(new_n12113_));
  INV_X1     g11920(.I(new_n12113_), .ZN(new_n12114_));
  OAI22_X1   g11921(.A1(new_n12114_), .A2(new_n12110_), .B1(new_n6338_), .B2(new_n12112_), .ZN(new_n12115_));
  NAND2_X1   g11922(.A1(new_n11846_), .A2(new_n11841_), .ZN(new_n12116_));
  NAND2_X1   g11923(.A1(new_n12027_), .A2(new_n12116_), .ZN(new_n12117_));
  XOR2_X1    g11924(.A1(new_n12117_), .A2(new_n12115_), .Z(new_n12118_));
  XOR2_X1    g11925(.A1(new_n12109_), .A2(new_n12118_), .Z(new_n12119_));
  INV_X1     g11926(.I(new_n12119_), .ZN(new_n12120_));
  NAND2_X1   g11927(.A1(new_n12035_), .A2(new_n12032_), .ZN(new_n12121_));
  NAND2_X1   g11928(.A1(new_n12036_), .A2(new_n12028_), .ZN(new_n12122_));
  NAND2_X1   g11929(.A1(new_n12122_), .A2(new_n12121_), .ZN(new_n12123_));
  NOR2_X1    g11930(.A1(new_n4210_), .A2(new_n6563_), .ZN(new_n12124_));
  INV_X1     g11931(.I(new_n12124_), .ZN(new_n12125_));
  OAI22_X1   g11932(.A1(new_n6140_), .A2(new_n6127_), .B1(new_n4739_), .B2(new_n8421_), .ZN(new_n12126_));
  NAND2_X1   g11933(.A1(new_n12126_), .A2(new_n12125_), .ZN(new_n12127_));
  NAND3_X1   g11934(.A1(new_n12127_), .A2(\a[37] ), .A3(\a[54] ), .ZN(new_n12128_));
  AOI22_X1   g11935(.A1(\a[38] ), .A2(\a[53] ), .B1(\a[39] ), .B2(\a[52] ), .ZN(new_n12129_));
  NAND2_X1   g11936(.A1(new_n12127_), .A2(new_n12125_), .ZN(new_n12130_));
  OAI21_X1   g11937(.A1(new_n12129_), .A2(new_n12130_), .B(new_n12128_), .ZN(new_n12131_));
  XOR2_X1    g11938(.A1(new_n12131_), .A2(new_n12002_), .Z(new_n12132_));
  NAND2_X1   g11939(.A1(new_n3210_), .A2(new_n7451_), .ZN(new_n12133_));
  NAND2_X1   g11940(.A1(new_n2275_), .A2(new_n7800_), .ZN(new_n12134_));
  AOI22_X1   g11941(.A1(new_n12133_), .A2(new_n12134_), .B1(new_n2636_), .B2(new_n7205_), .ZN(new_n12135_));
  NAND2_X1   g11942(.A1(\a[31] ), .A2(\a[60] ), .ZN(new_n12136_));
  AOI22_X1   g11943(.A1(\a[32] ), .A2(\a[59] ), .B1(\a[33] ), .B2(\a[58] ), .ZN(new_n12137_));
  NAND2_X1   g11944(.A1(new_n2636_), .A2(new_n7205_), .ZN(new_n12138_));
  NAND3_X1   g11945(.A1(new_n12138_), .A2(new_n12133_), .A3(new_n12134_), .ZN(new_n12139_));
  OAI22_X1   g11946(.A1(new_n12135_), .A2(new_n12136_), .B1(new_n12139_), .B2(new_n12137_), .ZN(new_n12140_));
  XOR2_X1    g11947(.A1(new_n12132_), .A2(new_n12140_), .Z(new_n12141_));
  XOR2_X1    g11948(.A1(new_n12123_), .A2(new_n12141_), .Z(new_n12142_));
  XOR2_X1    g11949(.A1(new_n12142_), .A2(new_n12120_), .Z(new_n12143_));
  XOR2_X1    g11950(.A1(new_n12106_), .A2(new_n12143_), .Z(new_n12144_));
  INV_X1     g11951(.I(new_n11966_), .ZN(new_n12145_));
  NOR2_X1    g11952(.A1(new_n11932_), .A2(new_n12145_), .ZN(new_n12146_));
  NOR2_X1    g11953(.A1(new_n11967_), .A2(new_n12011_), .ZN(new_n12147_));
  NOR2_X1    g11954(.A1(new_n12147_), .A2(new_n12146_), .ZN(new_n12148_));
  NAND2_X1   g11955(.A1(new_n12009_), .A2(new_n11993_), .ZN(new_n12149_));
  NAND2_X1   g11956(.A1(new_n12010_), .A2(new_n11970_), .ZN(new_n12150_));
  NAND2_X1   g11957(.A1(new_n12150_), .A2(new_n12149_), .ZN(new_n12151_));
  NAND2_X1   g11958(.A1(new_n11962_), .A2(new_n11964_), .ZN(new_n12152_));
  NAND2_X1   g11959(.A1(new_n11965_), .A2(new_n11959_), .ZN(new_n12153_));
  NAND2_X1   g11960(.A1(new_n12153_), .A2(new_n12152_), .ZN(new_n12154_));
  NOR2_X1    g11961(.A1(new_n2030_), .A2(new_n6897_), .ZN(new_n12155_));
  XOR2_X1    g11962(.A1(new_n11954_), .A2(new_n12155_), .Z(new_n12156_));
  XOR2_X1    g11963(.A1(new_n12156_), .A2(new_n11938_), .Z(new_n12157_));
  OAI21_X1   g11964(.A1(new_n11945_), .A2(new_n11947_), .B(new_n11939_), .ZN(new_n12158_));
  INV_X1     g11965(.I(new_n11957_), .ZN(new_n12159_));
  OAI21_X1   g11966(.A1(new_n11949_), .A2(new_n12159_), .B(new_n12158_), .ZN(new_n12160_));
  NOR2_X1    g11967(.A1(new_n11991_), .A2(new_n11987_), .ZN(new_n12161_));
  INV_X1     g11968(.I(new_n12161_), .ZN(new_n12162_));
  NOR2_X1    g11969(.A1(new_n12162_), .A2(new_n12160_), .ZN(new_n12163_));
  NAND2_X1   g11970(.A1(new_n12162_), .A2(new_n12160_), .ZN(new_n12164_));
  INV_X1     g11971(.I(new_n12164_), .ZN(new_n12165_));
  NOR2_X1    g11972(.A1(new_n12165_), .A2(new_n12163_), .ZN(new_n12166_));
  NAND2_X1   g11973(.A1(new_n12166_), .A2(new_n12157_), .ZN(new_n12167_));
  INV_X1     g11974(.I(new_n12167_), .ZN(new_n12168_));
  NOR2_X1    g11975(.A1(new_n12166_), .A2(new_n12157_), .ZN(new_n12169_));
  NOR2_X1    g11976(.A1(new_n12168_), .A2(new_n12169_), .ZN(new_n12170_));
  XNOR2_X1   g11977(.A1(new_n12154_), .A2(new_n12170_), .ZN(new_n12171_));
  XOR2_X1    g11978(.A1(new_n12171_), .A2(new_n12151_), .Z(new_n12172_));
  XOR2_X1    g11979(.A1(new_n12148_), .A2(new_n12172_), .Z(new_n12173_));
  XOR2_X1    g11980(.A1(new_n12144_), .A2(new_n12173_), .Z(new_n12174_));
  NOR2_X1    g11981(.A1(new_n12174_), .A2(new_n12065_), .ZN(new_n12175_));
  NAND2_X1   g11982(.A1(new_n12174_), .A2(new_n12065_), .ZN(new_n12176_));
  INV_X1     g11983(.I(new_n12176_), .ZN(new_n12177_));
  NOR2_X1    g11984(.A1(new_n12177_), .A2(new_n12175_), .ZN(new_n12178_));
  XOR2_X1    g11985(.A1(new_n12062_), .A2(new_n12178_), .Z(\asquared[92] ));
  AOI21_X1   g11986(.A1(new_n12061_), .A2(new_n12048_), .B(new_n12175_), .ZN(new_n12180_));
  NOR2_X1    g11987(.A1(new_n12180_), .A2(new_n12177_), .ZN(new_n12181_));
  INV_X1     g11988(.I(new_n12151_), .ZN(new_n12182_));
  NAND2_X1   g11989(.A1(new_n12154_), .A2(new_n12170_), .ZN(new_n12183_));
  OAI21_X1   g11990(.A1(new_n12171_), .A2(new_n12182_), .B(new_n12183_), .ZN(new_n12184_));
  NOR2_X1    g11991(.A1(new_n12168_), .A2(new_n12165_), .ZN(new_n12185_));
  NOR2_X1    g11992(.A1(new_n4704_), .A2(new_n4977_), .ZN(new_n12186_));
  NOR2_X1    g11993(.A1(new_n4034_), .A2(new_n4979_), .ZN(new_n12187_));
  NOR2_X1    g11994(.A1(new_n4343_), .A2(new_n4981_), .ZN(new_n12188_));
  NOR2_X1    g11995(.A1(new_n12187_), .A2(new_n12188_), .ZN(new_n12189_));
  NOR2_X1    g11996(.A1(new_n12189_), .A2(new_n12186_), .ZN(new_n12190_));
  NOR2_X1    g11997(.A1(new_n12190_), .A2(new_n12186_), .ZN(new_n12191_));
  INV_X1     g11998(.I(new_n12191_), .ZN(new_n12192_));
  AOI21_X1   g11999(.A1(\a[44] ), .A2(\a[48] ), .B(new_n4313_), .ZN(new_n12193_));
  NAND2_X1   g12000(.A1(\a[43] ), .A2(\a[49] ), .ZN(new_n12194_));
  OAI22_X1   g12001(.A1(new_n12192_), .A2(new_n12193_), .B1(new_n12190_), .B2(new_n12194_), .ZN(new_n12195_));
  AOI22_X1   g12002(.A1(\a[35] ), .A2(\a[57] ), .B1(\a[42] ), .B2(\a[50] ), .ZN(new_n12196_));
  NAND4_X1   g12003(.A1(\a[35] ), .A2(\a[42] ), .A3(\a[50] ), .A4(\a[57] ), .ZN(new_n12197_));
  NOR2_X1    g12004(.A1(new_n2746_), .A2(new_n6804_), .ZN(new_n12198_));
  NOR4_X1    g12005(.A1(new_n2442_), .A2(new_n3746_), .A3(new_n4901_), .A4(new_n6316_), .ZN(new_n12199_));
  OAI21_X1   g12006(.A1(new_n12198_), .A2(new_n12199_), .B(new_n12197_), .ZN(new_n12200_));
  NAND2_X1   g12007(.A1(new_n12200_), .A2(new_n12197_), .ZN(new_n12201_));
  NAND3_X1   g12008(.A1(new_n12200_), .A2(\a[34] ), .A3(\a[58] ), .ZN(new_n12202_));
  OAI21_X1   g12009(.A1(new_n12196_), .A2(new_n12201_), .B(new_n12202_), .ZN(new_n12203_));
  XOR2_X1    g12010(.A1(new_n12195_), .A2(new_n12203_), .Z(new_n12204_));
  AOI21_X1   g12011(.A1(\a[33] ), .A2(\a[59] ), .B(new_n10572_), .ZN(new_n12205_));
  NAND2_X1   g12012(.A1(\a[36] ), .A2(\a[56] ), .ZN(new_n12206_));
  NAND3_X1   g12013(.A1(new_n10572_), .A2(\a[33] ), .A3(\a[59] ), .ZN(new_n12207_));
  INV_X1     g12014(.I(new_n12207_), .ZN(new_n12208_));
  NOR3_X1    g12015(.A1(new_n12208_), .A2(new_n12205_), .A3(new_n12206_), .ZN(new_n12209_));
  NOR2_X1    g12016(.A1(new_n12209_), .A2(new_n12208_), .ZN(new_n12210_));
  INV_X1     g12017(.I(new_n12210_), .ZN(new_n12211_));
  OAI22_X1   g12018(.A1(new_n12211_), .A2(new_n12205_), .B1(new_n12206_), .B2(new_n12209_), .ZN(new_n12212_));
  XNOR2_X1   g12019(.A1(new_n12204_), .A2(new_n12212_), .ZN(new_n12213_));
  NAND2_X1   g12020(.A1(new_n11954_), .A2(new_n12155_), .ZN(new_n12214_));
  NAND2_X1   g12021(.A1(new_n12156_), .A2(new_n11938_), .ZN(new_n12215_));
  NAND2_X1   g12022(.A1(new_n12215_), .A2(new_n12214_), .ZN(new_n12216_));
  NAND2_X1   g12023(.A1(\a[31] ), .A2(\a[61] ), .ZN(new_n12217_));
  NAND2_X1   g12024(.A1(\a[30] ), .A2(\a[62] ), .ZN(new_n12218_));
  AOI22_X1   g12025(.A1(new_n2437_), .A2(new_n7590_), .B1(new_n12217_), .B2(new_n12218_), .ZN(new_n12219_));
  XNOR2_X1   g12026(.A1(new_n12087_), .A2(new_n12219_), .ZN(new_n12220_));
  NAND2_X1   g12027(.A1(new_n3328_), .A2(new_n5682_), .ZN(new_n12221_));
  NAND2_X1   g12028(.A1(new_n3550_), .A2(new_n5862_), .ZN(new_n12222_));
  AOI22_X1   g12029(.A1(new_n12221_), .A2(new_n12222_), .B1(new_n4534_), .B2(new_n5524_), .ZN(new_n12223_));
  NAND2_X1   g12030(.A1(\a[39] ), .A2(\a[53] ), .ZN(new_n12224_));
  AOI22_X1   g12031(.A1(\a[40] ), .A2(\a[52] ), .B1(\a[41] ), .B2(\a[51] ), .ZN(new_n12225_));
  NAND2_X1   g12032(.A1(new_n4534_), .A2(new_n5524_), .ZN(new_n12226_));
  NAND3_X1   g12033(.A1(new_n12226_), .A2(new_n12221_), .A3(new_n12222_), .ZN(new_n12227_));
  OAI22_X1   g12034(.A1(new_n12223_), .A2(new_n12224_), .B1(new_n12227_), .B2(new_n12225_), .ZN(new_n12228_));
  XNOR2_X1   g12035(.A1(new_n12220_), .A2(new_n12228_), .ZN(new_n12229_));
  XOR2_X1    g12036(.A1(new_n12229_), .A2(new_n12216_), .Z(new_n12230_));
  INV_X1     g12037(.I(new_n12230_), .ZN(new_n12231_));
  NAND2_X1   g12038(.A1(new_n12213_), .A2(new_n12231_), .ZN(new_n12232_));
  OR2_X2     g12039(.A1(new_n12213_), .A2(new_n12231_), .Z(new_n12233_));
  NAND2_X1   g12040(.A1(new_n12233_), .A2(new_n12232_), .ZN(new_n12234_));
  XOR2_X1    g12041(.A1(new_n12185_), .A2(new_n12234_), .Z(new_n12235_));
  INV_X1     g12042(.I(new_n12141_), .ZN(new_n12236_));
  NAND2_X1   g12043(.A1(new_n12123_), .A2(new_n12236_), .ZN(new_n12237_));
  OAI21_X1   g12044(.A1(new_n12142_), .A2(new_n12120_), .B(new_n12237_), .ZN(new_n12238_));
  XOR2_X1    g12045(.A1(new_n12235_), .A2(new_n12238_), .Z(new_n12239_));
  XOR2_X1    g12046(.A1(new_n12239_), .A2(new_n12184_), .Z(new_n12240_));
  NAND2_X1   g12047(.A1(new_n12106_), .A2(new_n12143_), .ZN(new_n12241_));
  OAI21_X1   g12048(.A1(new_n12066_), .A2(new_n12105_), .B(new_n12241_), .ZN(new_n12242_));
  NAND2_X1   g12049(.A1(new_n12074_), .A2(new_n12082_), .ZN(new_n12243_));
  NAND2_X1   g12050(.A1(new_n12083_), .A2(new_n12088_), .ZN(new_n12244_));
  NAND2_X1   g12051(.A1(new_n12244_), .A2(new_n12243_), .ZN(new_n12245_));
  NAND2_X1   g12052(.A1(new_n12131_), .A2(new_n12003_), .ZN(new_n12246_));
  INV_X1     g12053(.I(new_n12140_), .ZN(new_n12247_));
  OAI21_X1   g12054(.A1(new_n12132_), .A2(new_n12247_), .B(new_n12246_), .ZN(new_n12248_));
  NOR2_X1    g12055(.A1(new_n12094_), .A2(new_n11976_), .ZN(new_n12249_));
  INV_X1     g12056(.I(new_n12095_), .ZN(new_n12250_));
  NOR2_X1    g12057(.A1(new_n12250_), .A2(new_n12093_), .ZN(new_n12251_));
  NOR2_X1    g12058(.A1(new_n12251_), .A2(new_n12249_), .ZN(new_n12252_));
  INV_X1     g12059(.I(new_n12252_), .ZN(new_n12253_));
  NOR2_X1    g12060(.A1(new_n12253_), .A2(new_n12248_), .ZN(new_n12254_));
  NAND2_X1   g12061(.A1(new_n12253_), .A2(new_n12248_), .ZN(new_n12255_));
  INV_X1     g12062(.I(new_n12255_), .ZN(new_n12256_));
  NOR2_X1    g12063(.A1(new_n12256_), .A2(new_n12254_), .ZN(new_n12257_));
  NAND2_X1   g12064(.A1(new_n12257_), .A2(new_n12245_), .ZN(new_n12258_));
  INV_X1     g12065(.I(new_n12258_), .ZN(new_n12259_));
  NOR2_X1    g12066(.A1(new_n12257_), .A2(new_n12245_), .ZN(new_n12260_));
  NOR2_X1    g12067(.A1(new_n12259_), .A2(new_n12260_), .ZN(new_n12261_));
  NOR2_X1    g12068(.A1(new_n12103_), .A2(new_n12099_), .ZN(new_n12262_));
  NAND2_X1   g12069(.A1(new_n12117_), .A2(new_n12115_), .ZN(new_n12263_));
  NAND2_X1   g12070(.A1(new_n12109_), .A2(new_n12118_), .ZN(new_n12264_));
  NAND2_X1   g12071(.A1(new_n12264_), .A2(new_n12263_), .ZN(new_n12265_));
  XOR2_X1    g12072(.A1(new_n12130_), .A2(new_n12139_), .Z(new_n12266_));
  XOR2_X1    g12073(.A1(new_n12266_), .A2(new_n12072_), .Z(new_n12267_));
  XOR2_X1    g12074(.A1(new_n12113_), .A2(new_n12079_), .Z(new_n12268_));
  NAND2_X1   g12075(.A1(\a[32] ), .A2(\a[60] ), .ZN(new_n12269_));
  AOI22_X1   g12076(.A1(\a[37] ), .A2(\a[55] ), .B1(\a[38] ), .B2(\a[54] ), .ZN(new_n12270_));
  NOR2_X1    g12077(.A1(new_n6140_), .A2(new_n6129_), .ZN(new_n12271_));
  NOR3_X1    g12078(.A1(new_n12271_), .A2(new_n12269_), .A3(new_n12270_), .ZN(new_n12272_));
  NOR2_X1    g12079(.A1(new_n12272_), .A2(new_n12271_), .ZN(new_n12273_));
  INV_X1     g12080(.I(new_n12273_), .ZN(new_n12274_));
  OAI22_X1   g12081(.A1(new_n12274_), .A2(new_n12270_), .B1(new_n12269_), .B2(new_n12272_), .ZN(new_n12275_));
  XNOR2_X1   g12082(.A1(new_n12268_), .A2(new_n12275_), .ZN(new_n12276_));
  XNOR2_X1   g12083(.A1(new_n12267_), .A2(new_n12276_), .ZN(new_n12277_));
  NOR2_X1    g12084(.A1(new_n12277_), .A2(new_n12265_), .ZN(new_n12278_));
  NAND2_X1   g12085(.A1(new_n12277_), .A2(new_n12265_), .ZN(new_n12279_));
  INV_X1     g12086(.I(new_n12279_), .ZN(new_n12280_));
  NOR2_X1    g12087(.A1(new_n12280_), .A2(new_n12278_), .ZN(new_n12281_));
  INV_X1     g12088(.I(new_n12281_), .ZN(new_n12282_));
  XOR2_X1    g12089(.A1(new_n12262_), .A2(new_n12282_), .Z(new_n12283_));
  NOR2_X1    g12090(.A1(new_n12283_), .A2(new_n12261_), .ZN(new_n12284_));
  NAND2_X1   g12091(.A1(new_n12283_), .A2(new_n12261_), .ZN(new_n12285_));
  INV_X1     g12092(.I(new_n12285_), .ZN(new_n12286_));
  NOR2_X1    g12093(.A1(new_n12286_), .A2(new_n12284_), .ZN(new_n12287_));
  XOR2_X1    g12094(.A1(new_n12242_), .A2(new_n12287_), .Z(new_n12288_));
  XNOR2_X1   g12095(.A1(new_n12288_), .A2(new_n12240_), .ZN(new_n12289_));
  NOR2_X1    g12096(.A1(new_n12148_), .A2(new_n12172_), .ZN(new_n12290_));
  AOI21_X1   g12097(.A1(new_n12144_), .A2(new_n12173_), .B(new_n12290_), .ZN(new_n12291_));
  NOR2_X1    g12098(.A1(new_n12289_), .A2(new_n12291_), .ZN(new_n12292_));
  INV_X1     g12099(.I(new_n12292_), .ZN(new_n12293_));
  NAND2_X1   g12100(.A1(new_n12289_), .A2(new_n12291_), .ZN(new_n12294_));
  NAND2_X1   g12101(.A1(new_n12293_), .A2(new_n12294_), .ZN(new_n12295_));
  INV_X1     g12102(.I(new_n12048_), .ZN(new_n12296_));
  INV_X1     g12103(.I(new_n12175_), .ZN(new_n12297_));
  OAI21_X1   g12104(.A1(new_n12059_), .A2(new_n12296_), .B(new_n12297_), .ZN(new_n12298_));
  INV_X1     g12105(.I(new_n12294_), .ZN(new_n12299_));
  AOI21_X1   g12106(.A1(new_n12298_), .A2(new_n12176_), .B(new_n12299_), .ZN(new_n12300_));
  AOI22_X1   g12107(.A1(new_n12300_), .A2(new_n12293_), .B1(new_n12181_), .B2(new_n12295_), .ZN(\asquared[93] ));
  OAI21_X1   g12108(.A1(new_n12180_), .A2(new_n12177_), .B(new_n12294_), .ZN(new_n12302_));
  NAND2_X1   g12109(.A1(new_n12302_), .A2(new_n12293_), .ZN(new_n12303_));
  NAND2_X1   g12110(.A1(new_n12242_), .A2(new_n12287_), .ZN(new_n12304_));
  NAND2_X1   g12111(.A1(new_n12288_), .A2(new_n12240_), .ZN(new_n12305_));
  NAND2_X1   g12112(.A1(new_n12305_), .A2(new_n12304_), .ZN(new_n12306_));
  NOR2_X1    g12113(.A1(new_n12262_), .A2(new_n12282_), .ZN(new_n12307_));
  NOR2_X1    g12114(.A1(new_n12286_), .A2(new_n12307_), .ZN(new_n12308_));
  OAI21_X1   g12115(.A1(new_n12185_), .A2(new_n12234_), .B(new_n12233_), .ZN(new_n12309_));
  NOR2_X1    g12116(.A1(new_n12259_), .A2(new_n12256_), .ZN(new_n12310_));
  NOR3_X1    g12117(.A1(new_n11433_), .A2(new_n4030_), .A3(new_n5680_), .ZN(new_n12311_));
  NAND3_X1   g12118(.A1(new_n5093_), .A2(\a[48] ), .A3(\a[56] ), .ZN(new_n12312_));
  NOR2_X1    g12119(.A1(new_n6140_), .A2(new_n7185_), .ZN(new_n12313_));
  INV_X1     g12120(.I(new_n12313_), .ZN(new_n12314_));
  AOI21_X1   g12121(.A1(new_n12314_), .A2(new_n12312_), .B(new_n12311_), .ZN(new_n12315_));
  NAND2_X1   g12122(.A1(\a[37] ), .A2(\a[56] ), .ZN(new_n12316_));
  NOR2_X1    g12123(.A1(new_n12315_), .A2(new_n12311_), .ZN(new_n12317_));
  INV_X1     g12124(.I(new_n12317_), .ZN(new_n12318_));
  AOI22_X1   g12125(.A1(\a[38] ), .A2(\a[55] ), .B1(\a[45] ), .B2(\a[48] ), .ZN(new_n12319_));
  OAI22_X1   g12126(.A1(new_n12318_), .A2(new_n12319_), .B1(new_n12315_), .B2(new_n12316_), .ZN(new_n12320_));
  NAND2_X1   g12127(.A1(new_n4342_), .A2(new_n5154_), .ZN(new_n12321_));
  OAI22_X1   g12128(.A1(new_n3861_), .A2(new_n10168_), .B1(new_n4181_), .B2(new_n5440_), .ZN(new_n12322_));
  NAND2_X1   g12129(.A1(new_n12322_), .A2(new_n12321_), .ZN(new_n12323_));
  NAND3_X1   g12130(.A1(new_n12323_), .A2(\a[42] ), .A3(\a[51] ), .ZN(new_n12324_));
  AOI21_X1   g12131(.A1(\a[43] ), .A2(\a[50] ), .B(new_n6573_), .ZN(new_n12325_));
  NAND2_X1   g12132(.A1(new_n12323_), .A2(new_n12321_), .ZN(new_n12326_));
  OAI21_X1   g12133(.A1(new_n12325_), .A2(new_n12326_), .B(new_n12324_), .ZN(new_n12327_));
  XOR2_X1    g12134(.A1(new_n12320_), .A2(new_n12327_), .Z(new_n12328_));
  NOR3_X1    g12135(.A1(new_n2051_), .A2(new_n4312_), .A3(new_n7144_), .ZN(new_n12329_));
  NAND2_X1   g12136(.A1(new_n12329_), .A2(new_n4720_), .ZN(new_n12330_));
  AOI21_X1   g12137(.A1(\a[31] ), .A2(\a[62] ), .B(\a[47] ), .ZN(new_n12331_));
  NOR2_X1    g12138(.A1(new_n12329_), .A2(new_n4720_), .ZN(new_n12332_));
  INV_X1     g12139(.I(new_n12332_), .ZN(new_n12333_));
  OAI21_X1   g12140(.A1(new_n12333_), .A2(new_n12331_), .B(new_n12330_), .ZN(new_n12334_));
  XNOR2_X1   g12141(.A1(new_n12328_), .A2(new_n12334_), .ZN(new_n12335_));
  NAND2_X1   g12142(.A1(\a[35] ), .A2(\a[58] ), .ZN(new_n12336_));
  NOR2_X1    g12143(.A1(new_n9697_), .A2(new_n10612_), .ZN(new_n12337_));
  NAND4_X1   g12144(.A1(\a[35] ), .A2(\a[39] ), .A3(\a[54] ), .A4(\a[58] ), .ZN(new_n12338_));
  NAND2_X1   g12145(.A1(new_n3232_), .A2(new_n6803_), .ZN(new_n12339_));
  AOI21_X1   g12146(.A1(new_n12339_), .A2(new_n12338_), .B(new_n12337_), .ZN(new_n12340_));
  AOI22_X1   g12147(.A1(\a[36] ), .A2(\a[57] ), .B1(\a[39] ), .B2(\a[54] ), .ZN(new_n12341_));
  NOR2_X1    g12148(.A1(new_n12340_), .A2(new_n12337_), .ZN(new_n12342_));
  INV_X1     g12149(.I(new_n12342_), .ZN(new_n12343_));
  OAI22_X1   g12150(.A1(new_n12343_), .A2(new_n12341_), .B1(new_n12336_), .B2(new_n12340_), .ZN(new_n12344_));
  NOR2_X1    g12151(.A1(new_n2637_), .A2(new_n7454_), .ZN(new_n12345_));
  INV_X1     g12152(.I(new_n12345_), .ZN(new_n12346_));
  OAI22_X1   g12153(.A1(new_n2202_), .A2(new_n7959_), .B1(new_n7426_), .B2(new_n9031_), .ZN(new_n12347_));
  NAND2_X1   g12154(.A1(new_n12347_), .A2(new_n12346_), .ZN(new_n12348_));
  NAND3_X1   g12155(.A1(new_n12348_), .A2(\a[30] ), .A3(\a[63] ), .ZN(new_n12349_));
  AOI22_X1   g12156(.A1(\a[32] ), .A2(\a[61] ), .B1(\a[33] ), .B2(\a[60] ), .ZN(new_n12350_));
  NAND2_X1   g12157(.A1(new_n12348_), .A2(new_n12346_), .ZN(new_n12351_));
  OAI21_X1   g12158(.A1(new_n12350_), .A2(new_n12351_), .B(new_n12349_), .ZN(new_n12352_));
  XOR2_X1    g12159(.A1(new_n12344_), .A2(new_n12352_), .Z(new_n12353_));
  AOI22_X1   g12160(.A1(\a[40] ), .A2(\a[53] ), .B1(\a[41] ), .B2(\a[52] ), .ZN(new_n12354_));
  OAI21_X1   g12161(.A1(new_n5377_), .A2(new_n6563_), .B(new_n11550_), .ZN(new_n12355_));
  NOR2_X1    g12162(.A1(new_n12355_), .A2(new_n12354_), .ZN(new_n12356_));
  AOI21_X1   g12163(.A1(new_n4534_), .A2(new_n5862_), .B(new_n12356_), .ZN(new_n12357_));
  INV_X1     g12164(.I(new_n12357_), .ZN(new_n12358_));
  OAI22_X1   g12165(.A1(new_n12358_), .A2(new_n12354_), .B1(new_n11551_), .B2(new_n12356_), .ZN(new_n12359_));
  XNOR2_X1   g12166(.A1(new_n12353_), .A2(new_n12359_), .ZN(new_n12360_));
  XOR2_X1    g12167(.A1(new_n12335_), .A2(new_n12360_), .Z(new_n12361_));
  INV_X1     g12168(.I(new_n12361_), .ZN(new_n12362_));
  XOR2_X1    g12169(.A1(new_n12310_), .A2(new_n12362_), .Z(new_n12363_));
  XNOR2_X1   g12170(.A1(new_n12363_), .A2(new_n12309_), .ZN(new_n12364_));
  OR2_X2     g12171(.A1(new_n12308_), .A2(new_n12364_), .Z(new_n12365_));
  NAND2_X1   g12172(.A1(new_n12308_), .A2(new_n12364_), .ZN(new_n12366_));
  AND2_X2    g12173(.A1(new_n12365_), .A2(new_n12366_), .Z(new_n12367_));
  NAND2_X1   g12174(.A1(new_n12235_), .A2(new_n12238_), .ZN(new_n12368_));
  NAND2_X1   g12175(.A1(new_n12239_), .A2(new_n12184_), .ZN(new_n12369_));
  INV_X1     g12176(.I(new_n12228_), .ZN(new_n12370_));
  NAND2_X1   g12177(.A1(new_n12229_), .A2(new_n12216_), .ZN(new_n12371_));
  OAI21_X1   g12178(.A1(new_n12220_), .A2(new_n12370_), .B(new_n12371_), .ZN(new_n12372_));
  XNOR2_X1   g12179(.A1(new_n12191_), .A2(new_n12201_), .ZN(new_n12373_));
  XOR2_X1    g12180(.A1(new_n12373_), .A2(new_n12227_), .Z(new_n12374_));
  NAND2_X1   g12181(.A1(new_n12087_), .A2(new_n12219_), .ZN(new_n12375_));
  OAI21_X1   g12182(.A1(new_n2438_), .A2(new_n7591_), .B(new_n12375_), .ZN(new_n12376_));
  XOR2_X1    g12183(.A1(new_n12273_), .A2(new_n12210_), .Z(new_n12377_));
  XOR2_X1    g12184(.A1(new_n12377_), .A2(new_n12376_), .Z(new_n12378_));
  NAND2_X1   g12185(.A1(new_n12374_), .A2(new_n12378_), .ZN(new_n12379_));
  INV_X1     g12186(.I(new_n12379_), .ZN(new_n12380_));
  NOR2_X1    g12187(.A1(new_n12374_), .A2(new_n12378_), .ZN(new_n12381_));
  NOR2_X1    g12188(.A1(new_n12380_), .A2(new_n12381_), .ZN(new_n12382_));
  NOR2_X1    g12189(.A1(new_n12382_), .A2(new_n12372_), .ZN(new_n12383_));
  NAND2_X1   g12190(.A1(new_n12382_), .A2(new_n12372_), .ZN(new_n12384_));
  INV_X1     g12191(.I(new_n12384_), .ZN(new_n12385_));
  NOR2_X1    g12192(.A1(new_n12385_), .A2(new_n12383_), .ZN(new_n12386_));
  NAND2_X1   g12193(.A1(new_n12195_), .A2(new_n12203_), .ZN(new_n12387_));
  NAND2_X1   g12194(.A1(new_n12204_), .A2(new_n12212_), .ZN(new_n12388_));
  NAND2_X1   g12195(.A1(new_n12388_), .A2(new_n12387_), .ZN(new_n12389_));
  NAND2_X1   g12196(.A1(new_n12268_), .A2(new_n12275_), .ZN(new_n12390_));
  OAI21_X1   g12197(.A1(new_n12079_), .A2(new_n12113_), .B(new_n12390_), .ZN(new_n12391_));
  NAND2_X1   g12198(.A1(new_n12130_), .A2(new_n12139_), .ZN(new_n12392_));
  NAND2_X1   g12199(.A1(new_n12266_), .A2(new_n12072_), .ZN(new_n12393_));
  NAND2_X1   g12200(.A1(new_n12393_), .A2(new_n12392_), .ZN(new_n12394_));
  XOR2_X1    g12201(.A1(new_n12394_), .A2(new_n12391_), .Z(new_n12395_));
  XOR2_X1    g12202(.A1(new_n12395_), .A2(new_n12389_), .Z(new_n12396_));
  INV_X1     g12203(.I(new_n12396_), .ZN(new_n12397_));
  INV_X1     g12204(.I(new_n12267_), .ZN(new_n12398_));
  NOR2_X1    g12205(.A1(new_n12398_), .A2(new_n12276_), .ZN(new_n12399_));
  NOR2_X1    g12206(.A1(new_n12280_), .A2(new_n12399_), .ZN(new_n12400_));
  XOR2_X1    g12207(.A1(new_n12400_), .A2(new_n12397_), .Z(new_n12401_));
  NOR2_X1    g12208(.A1(new_n12401_), .A2(new_n12386_), .ZN(new_n12402_));
  NAND2_X1   g12209(.A1(new_n12401_), .A2(new_n12386_), .ZN(new_n12403_));
  INV_X1     g12210(.I(new_n12403_), .ZN(new_n12404_));
  NOR2_X1    g12211(.A1(new_n12404_), .A2(new_n12402_), .ZN(new_n12405_));
  INV_X1     g12212(.I(new_n12405_), .ZN(new_n12406_));
  AND3_X2    g12213(.A1(new_n12369_), .A2(new_n12368_), .A3(new_n12406_), .Z(new_n12407_));
  AOI21_X1   g12214(.A1(new_n12369_), .A2(new_n12368_), .B(new_n12406_), .ZN(new_n12408_));
  NOR2_X1    g12215(.A1(new_n12407_), .A2(new_n12408_), .ZN(new_n12409_));
  AND2_X2    g12216(.A1(new_n12367_), .A2(new_n12409_), .Z(new_n12410_));
  NOR2_X1    g12217(.A1(new_n12367_), .A2(new_n12409_), .ZN(new_n12411_));
  NOR2_X1    g12218(.A1(new_n12410_), .A2(new_n12411_), .ZN(new_n12412_));
  NOR2_X1    g12219(.A1(new_n12306_), .A2(new_n12412_), .ZN(new_n12413_));
  NAND2_X1   g12220(.A1(new_n12306_), .A2(new_n12412_), .ZN(new_n12414_));
  INV_X1     g12221(.I(new_n12414_), .ZN(new_n12415_));
  NOR2_X1    g12222(.A1(new_n12415_), .A2(new_n12413_), .ZN(new_n12416_));
  XOR2_X1    g12223(.A1(new_n12303_), .A2(new_n12416_), .Z(\asquared[94] ));
  AOI21_X1   g12224(.A1(new_n12302_), .A2(new_n12293_), .B(new_n12413_), .ZN(new_n12418_));
  NOR2_X1    g12225(.A1(new_n12418_), .A2(new_n12415_), .ZN(new_n12419_));
  NOR2_X1    g12226(.A1(new_n12400_), .A2(new_n12397_), .ZN(new_n12420_));
  NOR2_X1    g12227(.A1(new_n12404_), .A2(new_n12420_), .ZN(new_n12421_));
  NOR2_X1    g12228(.A1(new_n12343_), .A2(new_n12351_), .ZN(new_n12422_));
  NAND2_X1   g12229(.A1(new_n12343_), .A2(new_n12351_), .ZN(new_n12423_));
  INV_X1     g12230(.I(new_n12423_), .ZN(new_n12424_));
  NOR2_X1    g12231(.A1(new_n12424_), .A2(new_n12422_), .ZN(new_n12425_));
  INV_X1     g12232(.I(new_n12425_), .ZN(new_n12426_));
  NOR2_X1    g12233(.A1(new_n12426_), .A2(new_n12357_), .ZN(new_n12427_));
  INV_X1     g12234(.I(new_n12427_), .ZN(new_n12428_));
  NAND2_X1   g12235(.A1(new_n12426_), .A2(new_n12357_), .ZN(new_n12429_));
  AND2_X2    g12236(.A1(new_n12428_), .A2(new_n12429_), .Z(new_n12430_));
  NAND2_X1   g12237(.A1(new_n12320_), .A2(new_n12327_), .ZN(new_n12431_));
  NAND2_X1   g12238(.A1(new_n12328_), .A2(new_n12334_), .ZN(new_n12432_));
  NAND2_X1   g12239(.A1(new_n12432_), .A2(new_n12431_), .ZN(new_n12433_));
  NOR2_X1    g12240(.A1(new_n12333_), .A2(new_n10071_), .ZN(new_n12434_));
  NAND2_X1   g12241(.A1(new_n12333_), .A2(new_n10071_), .ZN(new_n12435_));
  INV_X1     g12242(.I(new_n12435_), .ZN(new_n12436_));
  NOR2_X1    g12243(.A1(new_n12436_), .A2(new_n12434_), .ZN(new_n12437_));
  NOR2_X1    g12244(.A1(new_n12318_), .A2(new_n12437_), .ZN(new_n12438_));
  NAND2_X1   g12245(.A1(new_n12318_), .A2(new_n12437_), .ZN(new_n12439_));
  INV_X1     g12246(.I(new_n12439_), .ZN(new_n12440_));
  NOR2_X1    g12247(.A1(new_n12440_), .A2(new_n12438_), .ZN(new_n12441_));
  XOR2_X1    g12248(.A1(new_n12433_), .A2(new_n12441_), .Z(new_n12442_));
  OR2_X2     g12249(.A1(new_n12442_), .A2(new_n12430_), .Z(new_n12443_));
  NAND2_X1   g12250(.A1(new_n12442_), .A2(new_n12430_), .ZN(new_n12444_));
  AND2_X2    g12251(.A1(new_n12443_), .A2(new_n12444_), .Z(new_n12445_));
  INV_X1     g12252(.I(new_n12445_), .ZN(new_n12446_));
  XOR2_X1    g12253(.A1(new_n12421_), .A2(new_n12446_), .Z(new_n12447_));
  NOR4_X1    g12254(.A1(new_n2442_), .A2(new_n3116_), .A3(new_n5680_), .A4(new_n6723_), .ZN(new_n12448_));
  NAND3_X1   g12255(.A1(new_n9015_), .A2(\a[57] ), .A3(\a[60] ), .ZN(new_n12449_));
  NAND2_X1   g12256(.A1(new_n4545_), .A2(new_n8951_), .ZN(new_n12450_));
  AOI21_X1   g12257(.A1(new_n12450_), .A2(new_n12449_), .B(new_n12448_), .ZN(new_n12451_));
  NAND2_X1   g12258(.A1(\a[37] ), .A2(\a[57] ), .ZN(new_n12452_));
  OR2_X2     g12259(.A1(new_n12451_), .A2(new_n12448_), .Z(new_n12453_));
  AOI22_X1   g12260(.A1(\a[34] ), .A2(\a[60] ), .B1(\a[39] ), .B2(\a[55] ), .ZN(new_n12454_));
  OAI22_X1   g12261(.A1(new_n12453_), .A2(new_n12454_), .B1(new_n12451_), .B2(new_n12452_), .ZN(new_n12455_));
  NOR2_X1    g12262(.A1(new_n2526_), .A2(new_n6899_), .ZN(new_n12456_));
  INV_X1     g12263(.I(new_n12456_), .ZN(new_n12457_));
  NOR2_X1    g12264(.A1(new_n6548_), .A2(new_n7144_), .ZN(new_n12458_));
  INV_X1     g12265(.I(new_n12458_), .ZN(new_n12459_));
  OAI22_X1   g12266(.A1(new_n2637_), .A2(new_n7591_), .B1(new_n5634_), .B2(new_n12459_), .ZN(new_n12460_));
  NAND2_X1   g12267(.A1(new_n12457_), .A2(new_n12460_), .ZN(new_n12461_));
  NAND3_X1   g12268(.A1(new_n12461_), .A2(\a[32] ), .A3(\a[62] ), .ZN(new_n12462_));
  AOI22_X1   g12269(.A1(\a[33] ), .A2(\a[61] ), .B1(\a[35] ), .B2(\a[59] ), .ZN(new_n12463_));
  NAND2_X1   g12270(.A1(new_n12461_), .A2(new_n12457_), .ZN(new_n12464_));
  OAI21_X1   g12271(.A1(new_n12463_), .A2(new_n12464_), .B(new_n12462_), .ZN(new_n12465_));
  XNOR2_X1   g12272(.A1(new_n12465_), .A2(new_n12326_), .ZN(new_n12466_));
  XNOR2_X1   g12273(.A1(new_n12466_), .A2(new_n12455_), .ZN(new_n12467_));
  NAND2_X1   g12274(.A1(new_n12394_), .A2(new_n12391_), .ZN(new_n12468_));
  NAND2_X1   g12275(.A1(new_n12395_), .A2(new_n12389_), .ZN(new_n12469_));
  NAND2_X1   g12276(.A1(new_n12469_), .A2(new_n12468_), .ZN(new_n12470_));
  AOI22_X1   g12277(.A1(\a[43] ), .A2(\a[51] ), .B1(\a[44] ), .B2(\a[50] ), .ZN(new_n12471_));
  INV_X1     g12278(.I(new_n12471_), .ZN(new_n12472_));
  NOR2_X1    g12279(.A1(new_n4343_), .A2(new_n5440_), .ZN(new_n12473_));
  NOR2_X1    g12280(.A1(new_n2626_), .A2(new_n6316_), .ZN(new_n12474_));
  AOI21_X1   g12281(.A1(new_n12472_), .A2(new_n12474_), .B(new_n12473_), .ZN(new_n12475_));
  INV_X1     g12282(.I(new_n12475_), .ZN(new_n12476_));
  OAI21_X1   g12283(.A1(new_n12473_), .A2(new_n12471_), .B(new_n12474_), .ZN(new_n12477_));
  OAI21_X1   g12284(.A1(new_n12476_), .A2(new_n12471_), .B(new_n12477_), .ZN(new_n12478_));
  NOR2_X1    g12285(.A1(new_n4667_), .A2(new_n6563_), .ZN(new_n12479_));
  NOR2_X1    g12286(.A1(new_n5377_), .A2(new_n6127_), .ZN(new_n12480_));
  NOR2_X1    g12287(.A1(new_n7757_), .A2(new_n8421_), .ZN(new_n12481_));
  NOR2_X1    g12288(.A1(new_n12480_), .A2(new_n12481_), .ZN(new_n12482_));
  NOR2_X1    g12289(.A1(new_n12482_), .A2(new_n12479_), .ZN(new_n12483_));
  NAND2_X1   g12290(.A1(\a[40] ), .A2(\a[54] ), .ZN(new_n12484_));
  AOI22_X1   g12291(.A1(\a[41] ), .A2(\a[53] ), .B1(\a[42] ), .B2(\a[52] ), .ZN(new_n12485_));
  NOR2_X1    g12292(.A1(new_n12483_), .A2(new_n12479_), .ZN(new_n12486_));
  INV_X1     g12293(.I(new_n12486_), .ZN(new_n12487_));
  OAI22_X1   g12294(.A1(new_n12487_), .A2(new_n12485_), .B1(new_n12483_), .B2(new_n12484_), .ZN(new_n12488_));
  XNOR2_X1   g12295(.A1(new_n12488_), .A2(new_n12478_), .ZN(new_n12489_));
  AOI22_X1   g12296(.A1(new_n4429_), .A2(new_n4980_), .B1(new_n6777_), .B2(new_n11140_), .ZN(new_n12490_));
  NOR2_X1    g12297(.A1(new_n9673_), .A2(new_n11141_), .ZN(new_n12491_));
  NOR2_X1    g12298(.A1(new_n12491_), .A2(new_n12490_), .ZN(new_n12492_));
  NOR2_X1    g12299(.A1(new_n12492_), .A2(new_n12491_), .ZN(new_n12493_));
  OAI21_X1   g12300(.A1(new_n6743_), .A2(new_n11140_), .B(new_n12493_), .ZN(new_n12494_));
  OAI21_X1   g12301(.A1(new_n6778_), .A2(new_n12492_), .B(new_n12494_), .ZN(new_n12495_));
  XOR2_X1    g12302(.A1(new_n12489_), .A2(new_n12495_), .Z(new_n12496_));
  INV_X1     g12303(.I(new_n12496_), .ZN(new_n12497_));
  NOR2_X1    g12304(.A1(new_n12470_), .A2(new_n12497_), .ZN(new_n12498_));
  NAND2_X1   g12305(.A1(new_n12470_), .A2(new_n12497_), .ZN(new_n12499_));
  INV_X1     g12306(.I(new_n12499_), .ZN(new_n12500_));
  NOR2_X1    g12307(.A1(new_n12500_), .A2(new_n12498_), .ZN(new_n12501_));
  NAND2_X1   g12308(.A1(new_n12501_), .A2(new_n12467_), .ZN(new_n12502_));
  INV_X1     g12309(.I(new_n12502_), .ZN(new_n12503_));
  NOR2_X1    g12310(.A1(new_n12501_), .A2(new_n12467_), .ZN(new_n12504_));
  NOR2_X1    g12311(.A1(new_n12503_), .A2(new_n12504_), .ZN(new_n12505_));
  XNOR2_X1   g12312(.A1(new_n12447_), .A2(new_n12505_), .ZN(new_n12506_));
  NAND2_X1   g12313(.A1(new_n12363_), .A2(new_n12309_), .ZN(new_n12507_));
  NAND2_X1   g12314(.A1(new_n12365_), .A2(new_n12507_), .ZN(new_n12508_));
  NOR2_X1    g12315(.A1(new_n12335_), .A2(new_n12360_), .ZN(new_n12509_));
  NOR2_X1    g12316(.A1(new_n12310_), .A2(new_n12362_), .ZN(new_n12510_));
  NOR2_X1    g12317(.A1(new_n12510_), .A2(new_n12509_), .ZN(new_n12511_));
  NAND2_X1   g12318(.A1(new_n12344_), .A2(new_n12352_), .ZN(new_n12512_));
  NAND2_X1   g12319(.A1(new_n12353_), .A2(new_n12359_), .ZN(new_n12513_));
  NAND2_X1   g12320(.A1(new_n12513_), .A2(new_n12512_), .ZN(new_n12514_));
  NAND2_X1   g12321(.A1(new_n12377_), .A2(new_n12376_), .ZN(new_n12515_));
  OAI21_X1   g12322(.A1(new_n12210_), .A2(new_n12273_), .B(new_n12515_), .ZN(new_n12516_));
  NAND2_X1   g12323(.A1(new_n12192_), .A2(new_n12201_), .ZN(new_n12517_));
  NAND2_X1   g12324(.A1(new_n12373_), .A2(new_n12227_), .ZN(new_n12518_));
  NAND2_X1   g12325(.A1(new_n12518_), .A2(new_n12517_), .ZN(new_n12519_));
  XOR2_X1    g12326(.A1(new_n12519_), .A2(new_n12516_), .Z(new_n12520_));
  XOR2_X1    g12327(.A1(new_n12520_), .A2(new_n12514_), .Z(new_n12521_));
  INV_X1     g12328(.I(new_n12521_), .ZN(new_n12522_));
  NOR2_X1    g12329(.A1(new_n12385_), .A2(new_n12380_), .ZN(new_n12523_));
  NOR2_X1    g12330(.A1(new_n12523_), .A2(new_n12522_), .ZN(new_n12524_));
  INV_X1     g12331(.I(new_n12524_), .ZN(new_n12525_));
  NAND2_X1   g12332(.A1(new_n12523_), .A2(new_n12522_), .ZN(new_n12526_));
  AND2_X2    g12333(.A1(new_n12525_), .A2(new_n12526_), .Z(new_n12527_));
  XNOR2_X1   g12334(.A1(new_n12527_), .A2(new_n12511_), .ZN(new_n12528_));
  XOR2_X1    g12335(.A1(new_n12508_), .A2(new_n12528_), .Z(new_n12529_));
  XOR2_X1    g12336(.A1(new_n12529_), .A2(new_n12506_), .Z(new_n12530_));
  NOR2_X1    g12337(.A1(new_n12410_), .A2(new_n12408_), .ZN(new_n12531_));
  NOR2_X1    g12338(.A1(new_n12530_), .A2(new_n12531_), .ZN(new_n12532_));
  INV_X1     g12339(.I(new_n12532_), .ZN(new_n12533_));
  NAND2_X1   g12340(.A1(new_n12530_), .A2(new_n12531_), .ZN(new_n12534_));
  NAND2_X1   g12341(.A1(new_n12533_), .A2(new_n12534_), .ZN(new_n12535_));
  XOR2_X1    g12342(.A1(new_n12419_), .A2(new_n12535_), .Z(\asquared[95] ));
  OAI21_X1   g12343(.A1(new_n12418_), .A2(new_n12415_), .B(new_n12534_), .ZN(new_n12537_));
  NAND2_X1   g12344(.A1(new_n12537_), .A2(new_n12533_), .ZN(new_n12538_));
  NAND2_X1   g12345(.A1(new_n12447_), .A2(new_n12505_), .ZN(new_n12539_));
  OAI21_X1   g12346(.A1(new_n12421_), .A2(new_n12446_), .B(new_n12539_), .ZN(new_n12540_));
  NOR2_X1    g12347(.A1(new_n12503_), .A2(new_n12500_), .ZN(new_n12541_));
  NAND2_X1   g12348(.A1(new_n12433_), .A2(new_n12441_), .ZN(new_n12542_));
  NAND2_X1   g12349(.A1(new_n12444_), .A2(new_n12542_), .ZN(new_n12543_));
  NOR2_X1    g12350(.A1(new_n12427_), .A2(new_n12424_), .ZN(new_n12544_));
  NOR2_X1    g12351(.A1(new_n12440_), .A2(new_n12436_), .ZN(new_n12545_));
  NOR2_X1    g12352(.A1(new_n3405_), .A2(new_n7452_), .ZN(new_n12546_));
  INV_X1     g12353(.I(new_n12546_), .ZN(new_n12547_));
  NOR2_X1    g12354(.A1(new_n2626_), .A2(new_n6548_), .ZN(new_n12548_));
  NOR2_X1    g12355(.A1(new_n2524_), .A2(new_n6723_), .ZN(new_n12549_));
  OAI21_X1   g12356(.A1(new_n12548_), .A2(new_n12549_), .B(new_n12547_), .ZN(new_n12550_));
  XNOR2_X1   g12357(.A1(new_n12550_), .A2(new_n12493_), .ZN(new_n12551_));
  XOR2_X1    g12358(.A1(new_n12545_), .A2(new_n12551_), .Z(new_n12552_));
  XNOR2_X1   g12359(.A1(new_n12552_), .A2(new_n12544_), .ZN(new_n12553_));
  XNOR2_X1   g12360(.A1(new_n12543_), .A2(new_n12553_), .ZN(new_n12554_));
  XOR2_X1    g12361(.A1(new_n12541_), .A2(new_n12554_), .Z(new_n12555_));
  NOR2_X1    g12362(.A1(new_n12540_), .A2(new_n12555_), .ZN(new_n12556_));
  NAND2_X1   g12363(.A1(new_n12540_), .A2(new_n12555_), .ZN(new_n12557_));
  INV_X1     g12364(.I(new_n12557_), .ZN(new_n12558_));
  NOR2_X1    g12365(.A1(new_n12558_), .A2(new_n12556_), .ZN(new_n12559_));
  NAND2_X1   g12366(.A1(new_n12519_), .A2(new_n12516_), .ZN(new_n12560_));
  NAND2_X1   g12367(.A1(new_n12520_), .A2(new_n12514_), .ZN(new_n12561_));
  NAND2_X1   g12368(.A1(new_n12561_), .A2(new_n12560_), .ZN(new_n12562_));
  NOR3_X1    g12369(.A1(new_n2274_), .A2(new_n4596_), .A3(new_n7144_), .ZN(new_n12563_));
  NAND2_X1   g12370(.A1(new_n12563_), .A2(new_n4976_), .ZN(new_n12564_));
  AOI21_X1   g12371(.A1(\a[33] ), .A2(\a[62] ), .B(\a[48] ), .ZN(new_n12565_));
  NOR2_X1    g12372(.A1(new_n12563_), .A2(new_n4976_), .ZN(new_n12566_));
  INV_X1     g12373(.I(new_n12566_), .ZN(new_n12567_));
  OAI21_X1   g12374(.A1(new_n12567_), .A2(new_n12565_), .B(new_n12564_), .ZN(new_n12568_));
  AOI22_X1   g12375(.A1(\a[45] ), .A2(\a[50] ), .B1(\a[46] ), .B2(\a[49] ), .ZN(new_n12569_));
  NOR2_X1    g12376(.A1(new_n3116_), .A2(new_n5856_), .ZN(new_n12570_));
  NOR2_X1    g12377(.A1(new_n4430_), .A2(new_n5155_), .ZN(new_n12571_));
  OAI21_X1   g12378(.A1(new_n12571_), .A2(new_n12569_), .B(new_n12570_), .ZN(new_n12572_));
  INV_X1     g12379(.I(new_n12569_), .ZN(new_n12573_));
  AOI21_X1   g12380(.A1(new_n12570_), .A2(new_n12573_), .B(new_n12571_), .ZN(new_n12574_));
  INV_X1     g12381(.I(new_n12574_), .ZN(new_n12575_));
  OAI21_X1   g12382(.A1(new_n12575_), .A2(new_n12569_), .B(new_n12572_), .ZN(new_n12576_));
  XNOR2_X1   g12383(.A1(new_n12576_), .A2(new_n12568_), .ZN(new_n12577_));
  NAND2_X1   g12384(.A1(new_n3860_), .A2(new_n5682_), .ZN(new_n12578_));
  NAND2_X1   g12385(.A1(new_n4180_), .A2(new_n5862_), .ZN(new_n12579_));
  AOI22_X1   g12386(.A1(new_n12578_), .A2(new_n12579_), .B1(new_n4342_), .B2(new_n5524_), .ZN(new_n12580_));
  NAND2_X1   g12387(.A1(\a[42] ), .A2(\a[53] ), .ZN(new_n12581_));
  AOI22_X1   g12388(.A1(\a[43] ), .A2(\a[52] ), .B1(\a[44] ), .B2(\a[51] ), .ZN(new_n12582_));
  NAND2_X1   g12389(.A1(new_n4342_), .A2(new_n5524_), .ZN(new_n12583_));
  NAND3_X1   g12390(.A1(new_n12583_), .A2(new_n12578_), .A3(new_n12579_), .ZN(new_n12584_));
  OAI22_X1   g12391(.A1(new_n12580_), .A2(new_n12581_), .B1(new_n12584_), .B2(new_n12582_), .ZN(new_n12585_));
  XOR2_X1    g12392(.A1(new_n12577_), .A2(new_n12585_), .Z(new_n12586_));
  INV_X1     g12393(.I(new_n12586_), .ZN(new_n12587_));
  XOR2_X1    g12394(.A1(new_n12562_), .A2(new_n12587_), .Z(new_n12588_));
  INV_X1     g12395(.I(new_n4741_), .ZN(new_n12589_));
  NAND2_X1   g12396(.A1(\a[55] ), .A2(\a[58] ), .ZN(new_n12590_));
  OAI22_X1   g12397(.A1(new_n6140_), .A2(new_n6804_), .B1(new_n12589_), .B2(new_n12590_), .ZN(new_n12591_));
  OAI21_X1   g12398(.A1(new_n3223_), .A2(new_n8952_), .B(new_n12591_), .ZN(new_n12592_));
  NAND3_X1   g12399(.A1(new_n12592_), .A2(\a[37] ), .A3(\a[58] ), .ZN(new_n12593_));
  AOI22_X1   g12400(.A1(\a[38] ), .A2(\a[57] ), .B1(\a[40] ), .B2(\a[55] ), .ZN(new_n12594_));
  NOR2_X1    g12401(.A1(new_n3223_), .A2(new_n8952_), .ZN(new_n12595_));
  NOR2_X1    g12402(.A1(new_n12591_), .A2(new_n12595_), .ZN(new_n12596_));
  INV_X1     g12403(.I(new_n12596_), .ZN(new_n12597_));
  OAI21_X1   g12404(.A1(new_n12594_), .A2(new_n12597_), .B(new_n12593_), .ZN(new_n12598_));
  XOR2_X1    g12405(.A1(new_n12598_), .A2(new_n12475_), .Z(new_n12599_));
  AOI22_X1   g12406(.A1(\a[32] ), .A2(\a[63] ), .B1(\a[34] ), .B2(\a[61] ), .ZN(new_n12600_));
  NOR2_X1    g12407(.A1(new_n3327_), .A2(new_n5617_), .ZN(new_n12601_));
  INV_X1     g12408(.I(new_n12601_), .ZN(new_n12602_));
  NOR2_X1    g12409(.A1(new_n3375_), .A2(new_n7959_), .ZN(new_n12603_));
  NOR3_X1    g12410(.A1(new_n12603_), .A2(new_n12600_), .A3(new_n12602_), .ZN(new_n12604_));
  NOR2_X1    g12411(.A1(new_n12604_), .A2(new_n12603_), .ZN(new_n12605_));
  INV_X1     g12412(.I(new_n12605_), .ZN(new_n12606_));
  OAI22_X1   g12413(.A1(new_n12606_), .A2(new_n12600_), .B1(new_n12602_), .B2(new_n12604_), .ZN(new_n12607_));
  XOR2_X1    g12414(.A1(new_n12599_), .A2(new_n12607_), .Z(new_n12608_));
  XOR2_X1    g12415(.A1(new_n12588_), .A2(new_n12608_), .Z(new_n12609_));
  INV_X1     g12416(.I(new_n12527_), .ZN(new_n12610_));
  OAI21_X1   g12417(.A1(new_n12610_), .A2(new_n12511_), .B(new_n12525_), .ZN(new_n12611_));
  XOR2_X1    g12418(.A1(new_n12464_), .A2(new_n12453_), .Z(new_n12612_));
  XOR2_X1    g12419(.A1(new_n12612_), .A2(new_n12487_), .Z(new_n12613_));
  INV_X1     g12420(.I(new_n12466_), .ZN(new_n12614_));
  NAND2_X1   g12421(.A1(new_n12614_), .A2(new_n12455_), .ZN(new_n12615_));
  NAND2_X1   g12422(.A1(new_n12465_), .A2(new_n12326_), .ZN(new_n12616_));
  NAND2_X1   g12423(.A1(new_n12615_), .A2(new_n12616_), .ZN(new_n12617_));
  NAND2_X1   g12424(.A1(new_n12488_), .A2(new_n12478_), .ZN(new_n12618_));
  INV_X1     g12425(.I(new_n12489_), .ZN(new_n12619_));
  NAND2_X1   g12426(.A1(new_n12619_), .A2(new_n12495_), .ZN(new_n12620_));
  NAND2_X1   g12427(.A1(new_n12620_), .A2(new_n12618_), .ZN(new_n12621_));
  XOR2_X1    g12428(.A1(new_n12621_), .A2(new_n12617_), .Z(new_n12622_));
  NAND2_X1   g12429(.A1(new_n12622_), .A2(new_n12613_), .ZN(new_n12623_));
  OR2_X2     g12430(.A1(new_n12622_), .A2(new_n12613_), .Z(new_n12624_));
  AND2_X2    g12431(.A1(new_n12624_), .A2(new_n12623_), .Z(new_n12625_));
  OR2_X2     g12432(.A1(new_n12611_), .A2(new_n12625_), .Z(new_n12626_));
  NAND2_X1   g12433(.A1(new_n12611_), .A2(new_n12625_), .ZN(new_n12627_));
  AND2_X2    g12434(.A1(new_n12626_), .A2(new_n12627_), .Z(new_n12628_));
  XOR2_X1    g12435(.A1(new_n12628_), .A2(new_n12609_), .Z(new_n12629_));
  XOR2_X1    g12436(.A1(new_n12559_), .A2(new_n12629_), .Z(new_n12630_));
  INV_X1     g12437(.I(new_n12630_), .ZN(new_n12631_));
  NOR2_X1    g12438(.A1(new_n12508_), .A2(new_n12528_), .ZN(new_n12632_));
  NAND2_X1   g12439(.A1(new_n12508_), .A2(new_n12528_), .ZN(new_n12633_));
  OAI21_X1   g12440(.A1(new_n12506_), .A2(new_n12632_), .B(new_n12633_), .ZN(new_n12634_));
  NOR2_X1    g12441(.A1(new_n12631_), .A2(new_n12634_), .ZN(new_n12635_));
  NAND2_X1   g12442(.A1(new_n12631_), .A2(new_n12634_), .ZN(new_n12636_));
  INV_X1     g12443(.I(new_n12636_), .ZN(new_n12637_));
  NOR2_X1    g12444(.A1(new_n12637_), .A2(new_n12635_), .ZN(new_n12638_));
  XOR2_X1    g12445(.A1(new_n12538_), .A2(new_n12638_), .Z(\asquared[96] ));
  AOI21_X1   g12446(.A1(new_n12537_), .A2(new_n12533_), .B(new_n12635_), .ZN(new_n12640_));
  NOR2_X1    g12447(.A1(new_n12640_), .A2(new_n12637_), .ZN(new_n12641_));
  NAND2_X1   g12448(.A1(new_n12464_), .A2(new_n12453_), .ZN(new_n12642_));
  NAND2_X1   g12449(.A1(new_n12612_), .A2(new_n12487_), .ZN(new_n12643_));
  NAND2_X1   g12450(.A1(new_n12643_), .A2(new_n12642_), .ZN(new_n12644_));
  NAND2_X1   g12451(.A1(\a[41] ), .A2(\a[55] ), .ZN(new_n12645_));
  NOR2_X1    g12452(.A1(new_n4181_), .A2(new_n6127_), .ZN(new_n12646_));
  NOR2_X1    g12453(.A1(new_n3666_), .A2(new_n5425_), .ZN(new_n12647_));
  NAND3_X1   g12454(.A1(new_n12647_), .A2(\a[41] ), .A3(\a[55] ), .ZN(new_n12648_));
  NAND2_X1   g12455(.A1(new_n4372_), .A2(new_n6128_), .ZN(new_n12649_));
  AOI21_X1   g12456(.A1(new_n12648_), .A2(new_n12649_), .B(new_n12646_), .ZN(new_n12650_));
  AOI21_X1   g12457(.A1(\a[42] ), .A2(\a[54] ), .B(new_n12647_), .ZN(new_n12651_));
  NOR2_X1    g12458(.A1(new_n12650_), .A2(new_n12646_), .ZN(new_n12652_));
  INV_X1     g12459(.I(new_n12652_), .ZN(new_n12653_));
  OAI22_X1   g12460(.A1(new_n12653_), .A2(new_n12651_), .B1(new_n12645_), .B2(new_n12650_), .ZN(new_n12654_));
  NAND2_X1   g12461(.A1(new_n2745_), .A2(new_n7590_), .ZN(new_n12655_));
  OAI22_X1   g12462(.A1(new_n2526_), .A2(new_n7959_), .B1(new_n3932_), .B2(new_n8049_), .ZN(new_n12656_));
  NAND2_X1   g12463(.A1(new_n12656_), .A2(new_n12655_), .ZN(new_n12657_));
  NAND3_X1   g12464(.A1(new_n12657_), .A2(\a[33] ), .A3(\a[63] ), .ZN(new_n12658_));
  AOI22_X1   g12465(.A1(\a[34] ), .A2(\a[62] ), .B1(\a[35] ), .B2(\a[61] ), .ZN(new_n12659_));
  NAND2_X1   g12466(.A1(new_n12657_), .A2(new_n12655_), .ZN(new_n12660_));
  OAI21_X1   g12467(.A1(new_n12659_), .A2(new_n12660_), .B(new_n12658_), .ZN(new_n12661_));
  XNOR2_X1   g12468(.A1(new_n12654_), .A2(new_n12661_), .ZN(new_n12662_));
  XNOR2_X1   g12469(.A1(new_n12662_), .A2(new_n12644_), .ZN(new_n12663_));
  INV_X1     g12470(.I(new_n12544_), .ZN(new_n12664_));
  NOR2_X1    g12471(.A1(new_n12545_), .A2(new_n12551_), .ZN(new_n12665_));
  AOI21_X1   g12472(.A1(new_n12664_), .A2(new_n12552_), .B(new_n12665_), .ZN(new_n12666_));
  OAI21_X1   g12473(.A1(new_n12550_), .A2(new_n12493_), .B(new_n12547_), .ZN(new_n12667_));
  NOR2_X1    g12474(.A1(new_n12606_), .A2(new_n12597_), .ZN(new_n12668_));
  NOR2_X1    g12475(.A1(new_n12605_), .A2(new_n12596_), .ZN(new_n12669_));
  NOR2_X1    g12476(.A1(new_n12668_), .A2(new_n12669_), .ZN(new_n12670_));
  XNOR2_X1   g12477(.A1(new_n12670_), .A2(new_n12667_), .ZN(new_n12671_));
  XOR2_X1    g12478(.A1(new_n12666_), .A2(new_n12671_), .Z(new_n12672_));
  XNOR2_X1   g12479(.A1(new_n12672_), .A2(new_n12663_), .ZN(new_n12673_));
  NAND2_X1   g12480(.A1(new_n12543_), .A2(new_n12553_), .ZN(new_n12674_));
  OAI21_X1   g12481(.A1(new_n12541_), .A2(new_n12554_), .B(new_n12674_), .ZN(new_n12675_));
  XOR2_X1    g12482(.A1(new_n12574_), .A2(new_n12566_), .Z(new_n12676_));
  XOR2_X1    g12483(.A1(new_n12676_), .A2(new_n12584_), .Z(new_n12677_));
  NAND2_X1   g12484(.A1(new_n12598_), .A2(new_n12476_), .ZN(new_n12678_));
  INV_X1     g12485(.I(new_n12607_), .ZN(new_n12679_));
  OAI21_X1   g12486(.A1(new_n12599_), .A2(new_n12679_), .B(new_n12678_), .ZN(new_n12680_));
  NAND2_X1   g12487(.A1(new_n12576_), .A2(new_n12568_), .ZN(new_n12681_));
  INV_X1     g12488(.I(new_n12585_), .ZN(new_n12682_));
  OAI21_X1   g12489(.A1(new_n12577_), .A2(new_n12682_), .B(new_n12681_), .ZN(new_n12683_));
  NOR2_X1    g12490(.A1(new_n12680_), .A2(new_n12683_), .ZN(new_n12684_));
  NAND2_X1   g12491(.A1(new_n12680_), .A2(new_n12683_), .ZN(new_n12685_));
  INV_X1     g12492(.I(new_n12685_), .ZN(new_n12686_));
  NOR2_X1    g12493(.A1(new_n12686_), .A2(new_n12684_), .ZN(new_n12687_));
  NAND2_X1   g12494(.A1(new_n12687_), .A2(new_n12677_), .ZN(new_n12688_));
  INV_X1     g12495(.I(new_n12688_), .ZN(new_n12689_));
  NOR2_X1    g12496(.A1(new_n12687_), .A2(new_n12677_), .ZN(new_n12690_));
  NOR2_X1    g12497(.A1(new_n12689_), .A2(new_n12690_), .ZN(new_n12691_));
  XOR2_X1    g12498(.A1(new_n12675_), .A2(new_n12691_), .Z(new_n12692_));
  INV_X1     g12499(.I(new_n12692_), .ZN(new_n12693_));
  OR2_X2     g12500(.A1(new_n12693_), .A2(new_n12673_), .Z(new_n12694_));
  NAND2_X1   g12501(.A1(new_n12693_), .A2(new_n12673_), .ZN(new_n12695_));
  AND2_X2    g12502(.A1(new_n12694_), .A2(new_n12695_), .Z(new_n12696_));
  INV_X1     g12503(.I(new_n12628_), .ZN(new_n12697_));
  OAI21_X1   g12504(.A1(new_n12697_), .A2(new_n12609_), .B(new_n12627_), .ZN(new_n12698_));
  NOR2_X1    g12505(.A1(new_n12589_), .A2(new_n10715_), .ZN(new_n12699_));
  INV_X1     g12506(.I(new_n12699_), .ZN(new_n12700_));
  NOR3_X1    g12507(.A1(new_n12206_), .A2(new_n3221_), .A3(new_n6723_), .ZN(new_n12701_));
  NOR2_X1    g12508(.A1(new_n3038_), .A2(new_n7452_), .ZN(new_n12702_));
  OAI21_X1   g12509(.A1(new_n12701_), .A2(new_n12702_), .B(new_n12700_), .ZN(new_n12703_));
  NAND3_X1   g12510(.A1(new_n12703_), .A2(\a[36] ), .A3(\a[60] ), .ZN(new_n12704_));
  NAND2_X1   g12511(.A1(new_n12703_), .A2(new_n12700_), .ZN(new_n12705_));
  AOI22_X1   g12512(.A1(\a[37] ), .A2(\a[59] ), .B1(\a[40] ), .B2(\a[56] ), .ZN(new_n12706_));
  OAI21_X1   g12513(.A1(new_n12705_), .A2(new_n12706_), .B(new_n12704_), .ZN(new_n12707_));
  AOI22_X1   g12514(.A1(\a[38] ), .A2(\a[58] ), .B1(\a[39] ), .B2(\a[57] ), .ZN(new_n12708_));
  NOR2_X1    g12515(.A1(new_n4210_), .A2(new_n6804_), .ZN(new_n12709_));
  OAI21_X1   g12516(.A1(new_n12709_), .A2(new_n12708_), .B(new_n7012_), .ZN(new_n12710_));
  INV_X1     g12517(.I(new_n12708_), .ZN(new_n12711_));
  AOI21_X1   g12518(.A1(new_n7012_), .A2(new_n12711_), .B(new_n12709_), .ZN(new_n12712_));
  INV_X1     g12519(.I(new_n12712_), .ZN(new_n12713_));
  OAI21_X1   g12520(.A1(new_n12713_), .A2(new_n12708_), .B(new_n12710_), .ZN(new_n12714_));
  XOR2_X1    g12521(.A1(new_n12707_), .A2(new_n12714_), .Z(new_n12715_));
  NAND2_X1   g12522(.A1(\a[45] ), .A2(\a[51] ), .ZN(new_n12716_));
  NAND3_X1   g12523(.A1(new_n4978_), .A2(\a[45] ), .A3(\a[51] ), .ZN(new_n12717_));
  NAND2_X1   g12524(.A1(new_n4429_), .A2(new_n5439_), .ZN(new_n12718_));
  AOI22_X1   g12525(.A1(new_n12718_), .A2(new_n12717_), .B1(new_n4720_), .B2(new_n5154_), .ZN(new_n12719_));
  NAND2_X1   g12526(.A1(new_n4720_), .A2(new_n5154_), .ZN(new_n12720_));
  NAND3_X1   g12527(.A1(new_n12720_), .A2(new_n12718_), .A3(new_n12717_), .ZN(new_n12721_));
  AOI21_X1   g12528(.A1(\a[46] ), .A2(\a[50] ), .B(new_n4978_), .ZN(new_n12722_));
  OAI22_X1   g12529(.A1(new_n12719_), .A2(new_n12716_), .B1(new_n12721_), .B2(new_n12722_), .ZN(new_n12723_));
  XOR2_X1    g12530(.A1(new_n12715_), .A2(new_n12723_), .Z(new_n12724_));
  NAND2_X1   g12531(.A1(new_n12621_), .A2(new_n12617_), .ZN(new_n12725_));
  NAND2_X1   g12532(.A1(new_n12623_), .A2(new_n12725_), .ZN(new_n12726_));
  XOR2_X1    g12533(.A1(new_n12726_), .A2(new_n12724_), .Z(new_n12727_));
  NAND2_X1   g12534(.A1(new_n12562_), .A2(new_n12587_), .ZN(new_n12728_));
  INV_X1     g12535(.I(new_n12588_), .ZN(new_n12729_));
  OAI21_X1   g12536(.A1(new_n12729_), .A2(new_n12608_), .B(new_n12728_), .ZN(new_n12730_));
  XNOR2_X1   g12537(.A1(new_n12727_), .A2(new_n12730_), .ZN(new_n12731_));
  NAND2_X1   g12538(.A1(new_n12698_), .A2(new_n12731_), .ZN(new_n12732_));
  NOR2_X1    g12539(.A1(new_n12698_), .A2(new_n12731_), .ZN(new_n12733_));
  INV_X1     g12540(.I(new_n12733_), .ZN(new_n12734_));
  NAND2_X1   g12541(.A1(new_n12734_), .A2(new_n12732_), .ZN(new_n12735_));
  NAND2_X1   g12542(.A1(new_n12735_), .A2(new_n12696_), .ZN(new_n12736_));
  INV_X1     g12543(.I(new_n12696_), .ZN(new_n12737_));
  NAND3_X1   g12544(.A1(new_n12734_), .A2(new_n12737_), .A3(new_n12732_), .ZN(new_n12738_));
  NAND2_X1   g12545(.A1(new_n12736_), .A2(new_n12738_), .ZN(new_n12739_));
  OAI21_X1   g12546(.A1(new_n12629_), .A2(new_n12556_), .B(new_n12557_), .ZN(new_n12740_));
  INV_X1     g12547(.I(new_n12740_), .ZN(new_n12741_));
  NOR2_X1    g12548(.A1(new_n12739_), .A2(new_n12741_), .ZN(new_n12742_));
  INV_X1     g12549(.I(new_n12742_), .ZN(new_n12743_));
  NAND2_X1   g12550(.A1(new_n12739_), .A2(new_n12741_), .ZN(new_n12744_));
  NAND2_X1   g12551(.A1(new_n12743_), .A2(new_n12744_), .ZN(new_n12745_));
  INV_X1     g12552(.I(new_n12413_), .ZN(new_n12746_));
  OAI21_X1   g12553(.A1(new_n12300_), .A2(new_n12292_), .B(new_n12746_), .ZN(new_n12747_));
  INV_X1     g12554(.I(new_n12534_), .ZN(new_n12748_));
  AOI21_X1   g12555(.A1(new_n12747_), .A2(new_n12414_), .B(new_n12748_), .ZN(new_n12749_));
  INV_X1     g12556(.I(new_n12635_), .ZN(new_n12750_));
  OAI21_X1   g12557(.A1(new_n12749_), .A2(new_n12532_), .B(new_n12750_), .ZN(new_n12751_));
  INV_X1     g12558(.I(new_n12744_), .ZN(new_n12752_));
  AOI21_X1   g12559(.A1(new_n12751_), .A2(new_n12636_), .B(new_n12752_), .ZN(new_n12753_));
  AOI22_X1   g12560(.A1(new_n12753_), .A2(new_n12743_), .B1(new_n12641_), .B2(new_n12745_), .ZN(\asquared[97] ));
  OAI21_X1   g12561(.A1(new_n12640_), .A2(new_n12637_), .B(new_n12744_), .ZN(new_n12755_));
  NAND2_X1   g12562(.A1(new_n12755_), .A2(new_n12743_), .ZN(new_n12756_));
  INV_X1     g12563(.I(new_n12731_), .ZN(new_n12757_));
  NAND2_X1   g12564(.A1(new_n12698_), .A2(new_n12757_), .ZN(new_n12758_));
  NAND2_X1   g12565(.A1(new_n12736_), .A2(new_n12758_), .ZN(new_n12759_));
  NAND2_X1   g12566(.A1(new_n12726_), .A2(new_n12724_), .ZN(new_n12760_));
  NAND2_X1   g12567(.A1(new_n12727_), .A2(new_n12730_), .ZN(new_n12761_));
  NAND2_X1   g12568(.A1(new_n12761_), .A2(new_n12760_), .ZN(new_n12762_));
  NOR2_X1    g12569(.A1(new_n2626_), .A2(new_n6897_), .ZN(new_n12763_));
  XOR2_X1    g12570(.A1(new_n12721_), .A2(new_n12763_), .Z(new_n12764_));
  XOR2_X1    g12571(.A1(new_n12764_), .A2(new_n12713_), .Z(new_n12765_));
  NAND2_X1   g12572(.A1(new_n12707_), .A2(new_n12714_), .ZN(new_n12766_));
  NAND2_X1   g12573(.A1(new_n12715_), .A2(new_n12723_), .ZN(new_n12767_));
  NAND2_X1   g12574(.A1(new_n12767_), .A2(new_n12766_), .ZN(new_n12768_));
  NAND2_X1   g12575(.A1(new_n12670_), .A2(new_n12667_), .ZN(new_n12769_));
  OAI21_X1   g12576(.A1(new_n12596_), .A2(new_n12605_), .B(new_n12769_), .ZN(new_n12770_));
  XOR2_X1    g12577(.A1(new_n12768_), .A2(new_n12770_), .Z(new_n12771_));
  XOR2_X1    g12578(.A1(new_n12771_), .A2(new_n12765_), .Z(new_n12772_));
  NAND2_X1   g12579(.A1(new_n12676_), .A2(new_n12584_), .ZN(new_n12773_));
  OAI21_X1   g12580(.A1(new_n12566_), .A2(new_n12574_), .B(new_n12773_), .ZN(new_n12774_));
  AOI21_X1   g12581(.A1(\a[47] ), .A2(\a[50] ), .B(new_n6930_), .ZN(new_n12775_));
  INV_X1     g12582(.I(new_n12775_), .ZN(new_n12776_));
  NOR2_X1    g12583(.A1(new_n4721_), .A2(new_n5440_), .ZN(new_n12777_));
  NOR2_X1    g12584(.A1(new_n3221_), .A2(new_n6298_), .ZN(new_n12778_));
  AOI21_X1   g12585(.A1(new_n12776_), .A2(new_n12778_), .B(new_n12777_), .ZN(new_n12779_));
  INV_X1     g12586(.I(new_n12779_), .ZN(new_n12780_));
  OAI21_X1   g12587(.A1(new_n12777_), .A2(new_n12775_), .B(new_n12778_), .ZN(new_n12781_));
  OAI21_X1   g12588(.A1(new_n12780_), .A2(new_n12775_), .B(new_n12781_), .ZN(new_n12782_));
  NOR4_X1    g12589(.A1(new_n2524_), .A2(new_n4596_), .A3(new_n4702_), .A4(new_n7144_), .ZN(new_n12783_));
  NOR3_X1    g12590(.A1(new_n2524_), .A2(new_n4702_), .A3(new_n7144_), .ZN(new_n12784_));
  AOI21_X1   g12591(.A1(\a[35] ), .A2(\a[62] ), .B(\a[49] ), .ZN(new_n12785_));
  NOR3_X1    g12592(.A1(new_n12784_), .A2(new_n4980_), .A3(new_n12785_), .ZN(new_n12786_));
  NOR2_X1    g12593(.A1(new_n12786_), .A2(new_n12783_), .ZN(new_n12787_));
  XOR2_X1    g12594(.A1(new_n12782_), .A2(new_n12787_), .Z(new_n12788_));
  XNOR2_X1   g12595(.A1(new_n12774_), .A2(new_n12788_), .ZN(new_n12789_));
  NAND2_X1   g12596(.A1(new_n12654_), .A2(new_n12661_), .ZN(new_n12790_));
  INV_X1     g12597(.I(new_n12662_), .ZN(new_n12791_));
  NAND2_X1   g12598(.A1(new_n12791_), .A2(new_n12644_), .ZN(new_n12792_));
  NAND2_X1   g12599(.A1(new_n12792_), .A2(new_n12790_), .ZN(new_n12793_));
  XOR2_X1    g12600(.A1(new_n12705_), .A2(new_n12660_), .Z(new_n12794_));
  XOR2_X1    g12601(.A1(new_n12794_), .A2(new_n12653_), .Z(new_n12795_));
  NOR2_X1    g12602(.A1(new_n12793_), .A2(new_n12795_), .ZN(new_n12796_));
  NAND2_X1   g12603(.A1(new_n12793_), .A2(new_n12795_), .ZN(new_n12797_));
  INV_X1     g12604(.I(new_n12797_), .ZN(new_n12798_));
  NOR2_X1    g12605(.A1(new_n12798_), .A2(new_n12796_), .ZN(new_n12799_));
  NAND2_X1   g12606(.A1(new_n12799_), .A2(new_n12789_), .ZN(new_n12800_));
  INV_X1     g12607(.I(new_n12800_), .ZN(new_n12801_));
  NOR2_X1    g12608(.A1(new_n12799_), .A2(new_n12789_), .ZN(new_n12802_));
  NOR2_X1    g12609(.A1(new_n12801_), .A2(new_n12802_), .ZN(new_n12803_));
  XOR2_X1    g12610(.A1(new_n12803_), .A2(new_n12772_), .Z(new_n12804_));
  XOR2_X1    g12611(.A1(new_n12762_), .A2(new_n12804_), .Z(new_n12805_));
  NAND2_X1   g12612(.A1(new_n12675_), .A2(new_n12691_), .ZN(new_n12806_));
  NAND2_X1   g12613(.A1(new_n12694_), .A2(new_n12806_), .ZN(new_n12807_));
  NOR2_X1    g12614(.A1(new_n12689_), .A2(new_n12686_), .ZN(new_n12808_));
  AOI22_X1   g12615(.A1(\a[34] ), .A2(\a[63] ), .B1(\a[42] ), .B2(\a[55] ), .ZN(new_n12809_));
  NAND4_X1   g12616(.A1(\a[34] ), .A2(\a[42] ), .A3(\a[55] ), .A4(\a[63] ), .ZN(new_n12810_));
  NOR2_X1    g12617(.A1(new_n4667_), .A2(new_n7185_), .ZN(new_n12811_));
  NOR4_X1    g12618(.A1(new_n2442_), .A2(new_n3327_), .A3(new_n5856_), .A4(new_n7643_), .ZN(new_n12812_));
  OAI21_X1   g12619(.A1(new_n12811_), .A2(new_n12812_), .B(new_n12810_), .ZN(new_n12813_));
  NAND2_X1   g12620(.A1(new_n12813_), .A2(new_n12810_), .ZN(new_n12814_));
  NAND3_X1   g12621(.A1(new_n12813_), .A2(\a[41] ), .A3(\a[56] ), .ZN(new_n12815_));
  OAI21_X1   g12622(.A1(new_n12809_), .A2(new_n12814_), .B(new_n12815_), .ZN(new_n12816_));
  NAND2_X1   g12623(.A1(new_n4209_), .A2(new_n7205_), .ZN(new_n12817_));
  OAI22_X1   g12624(.A1(new_n6140_), .A2(new_n7452_), .B1(new_n4739_), .B2(new_n7801_), .ZN(new_n12818_));
  NAND2_X1   g12625(.A1(new_n12818_), .A2(new_n12817_), .ZN(new_n12819_));
  NAND3_X1   g12626(.A1(new_n12819_), .A2(\a[37] ), .A3(\a[60] ), .ZN(new_n12820_));
  AOI22_X1   g12627(.A1(\a[38] ), .A2(\a[59] ), .B1(\a[39] ), .B2(\a[58] ), .ZN(new_n12821_));
  NAND2_X1   g12628(.A1(new_n12819_), .A2(new_n12817_), .ZN(new_n12822_));
  OAI21_X1   g12629(.A1(new_n12821_), .A2(new_n12822_), .B(new_n12820_), .ZN(new_n12823_));
  XOR2_X1    g12630(.A1(new_n12823_), .A2(new_n12816_), .Z(new_n12824_));
  NOR2_X1    g12631(.A1(new_n4704_), .A2(new_n6563_), .ZN(new_n12825_));
  AOI22_X1   g12632(.A1(new_n4033_), .A2(new_n8420_), .B1(new_n4342_), .B2(new_n6126_), .ZN(new_n12826_));
  NOR2_X1    g12633(.A1(new_n12825_), .A2(new_n12826_), .ZN(new_n12827_));
  NAND2_X1   g12634(.A1(\a[43] ), .A2(\a[54] ), .ZN(new_n12828_));
  AOI22_X1   g12635(.A1(\a[44] ), .A2(\a[53] ), .B1(\a[45] ), .B2(\a[52] ), .ZN(new_n12829_));
  NOR2_X1    g12636(.A1(new_n12827_), .A2(new_n12825_), .ZN(new_n12830_));
  INV_X1     g12637(.I(new_n12830_), .ZN(new_n12831_));
  OAI22_X1   g12638(.A1(new_n12831_), .A2(new_n12829_), .B1(new_n12827_), .B2(new_n12828_), .ZN(new_n12832_));
  XNOR2_X1   g12639(.A1(new_n12824_), .A2(new_n12832_), .ZN(new_n12833_));
  XOR2_X1    g12640(.A1(new_n12808_), .A2(new_n12833_), .Z(new_n12834_));
  NAND2_X1   g12641(.A1(new_n12672_), .A2(new_n12663_), .ZN(new_n12835_));
  OAI21_X1   g12642(.A1(new_n12666_), .A2(new_n12671_), .B(new_n12835_), .ZN(new_n12836_));
  XNOR2_X1   g12643(.A1(new_n12834_), .A2(new_n12836_), .ZN(new_n12837_));
  INV_X1     g12644(.I(new_n12837_), .ZN(new_n12838_));
  NOR2_X1    g12645(.A1(new_n12807_), .A2(new_n12838_), .ZN(new_n12839_));
  NAND2_X1   g12646(.A1(new_n12807_), .A2(new_n12838_), .ZN(new_n12840_));
  INV_X1     g12647(.I(new_n12840_), .ZN(new_n12841_));
  NOR2_X1    g12648(.A1(new_n12841_), .A2(new_n12839_), .ZN(new_n12842_));
  NAND2_X1   g12649(.A1(new_n12842_), .A2(new_n12805_), .ZN(new_n12843_));
  INV_X1     g12650(.I(new_n12843_), .ZN(new_n12844_));
  NOR2_X1    g12651(.A1(new_n12842_), .A2(new_n12805_), .ZN(new_n12845_));
  NOR2_X1    g12652(.A1(new_n12844_), .A2(new_n12845_), .ZN(new_n12846_));
  NOR2_X1    g12653(.A1(new_n12846_), .A2(new_n12759_), .ZN(new_n12847_));
  NAND2_X1   g12654(.A1(new_n12846_), .A2(new_n12759_), .ZN(new_n12848_));
  INV_X1     g12655(.I(new_n12848_), .ZN(new_n12849_));
  NOR2_X1    g12656(.A1(new_n12849_), .A2(new_n12847_), .ZN(new_n12850_));
  XOR2_X1    g12657(.A1(new_n12756_), .A2(new_n12850_), .Z(\asquared[98] ));
  AOI21_X1   g12658(.A1(new_n12755_), .A2(new_n12743_), .B(new_n12847_), .ZN(new_n12852_));
  NOR2_X1    g12659(.A1(new_n12852_), .A2(new_n12849_), .ZN(new_n12853_));
  NOR2_X1    g12660(.A1(new_n12844_), .A2(new_n12841_), .ZN(new_n12854_));
  NAND2_X1   g12661(.A1(new_n12834_), .A2(new_n12836_), .ZN(new_n12855_));
  OAI21_X1   g12662(.A1(new_n12808_), .A2(new_n12833_), .B(new_n12855_), .ZN(new_n12856_));
  INV_X1     g12663(.I(new_n12782_), .ZN(new_n12857_));
  INV_X1     g12664(.I(new_n12788_), .ZN(new_n12858_));
  NAND2_X1   g12665(.A1(new_n12858_), .A2(new_n12774_), .ZN(new_n12859_));
  OAI21_X1   g12666(.A1(new_n12857_), .A2(new_n12787_), .B(new_n12859_), .ZN(new_n12860_));
  XOR2_X1    g12667(.A1(new_n12822_), .A2(new_n12814_), .Z(new_n12861_));
  XOR2_X1    g12668(.A1(new_n12861_), .A2(new_n12831_), .Z(new_n12862_));
  NOR2_X1    g12669(.A1(new_n12860_), .A2(new_n12862_), .ZN(new_n12863_));
  NAND2_X1   g12670(.A1(new_n12860_), .A2(new_n12862_), .ZN(new_n12864_));
  INV_X1     g12671(.I(new_n12864_), .ZN(new_n12865_));
  NOR2_X1    g12672(.A1(new_n12865_), .A2(new_n12863_), .ZN(new_n12866_));
  NOR2_X1    g12673(.A1(new_n12784_), .A2(new_n4980_), .ZN(new_n12867_));
  NAND2_X1   g12674(.A1(new_n3037_), .A2(new_n7590_), .ZN(new_n12868_));
  OAI21_X1   g12675(.A1(new_n2752_), .A2(new_n6897_), .B(new_n9000_), .ZN(new_n12869_));
  NAND2_X1   g12676(.A1(new_n12868_), .A2(new_n12869_), .ZN(new_n12870_));
  NAND2_X1   g12677(.A1(new_n12870_), .A2(new_n12867_), .ZN(new_n12871_));
  NOR2_X1    g12678(.A1(new_n12870_), .A2(new_n12867_), .ZN(new_n12872_));
  INV_X1     g12679(.I(new_n12872_), .ZN(new_n12873_));
  AND2_X2    g12680(.A1(new_n12873_), .A2(new_n12871_), .Z(new_n12874_));
  NOR2_X1    g12681(.A1(new_n4977_), .A2(new_n5440_), .ZN(new_n12875_));
  NAND4_X1   g12682(.A1(\a[46] ), .A2(\a[48] ), .A3(\a[50] ), .A4(\a[52] ), .ZN(new_n12876_));
  OAI21_X1   g12683(.A1(new_n4721_), .A2(new_n5525_), .B(new_n12876_), .ZN(new_n12877_));
  NOR2_X1    g12684(.A1(new_n12877_), .A2(new_n12875_), .ZN(new_n12878_));
  OAI21_X1   g12685(.A1(new_n4902_), .A2(new_n7162_), .B(new_n12878_), .ZN(new_n12879_));
  OAI21_X1   g12686(.A1(new_n4977_), .A2(new_n5440_), .B(new_n12877_), .ZN(new_n12880_));
  NAND3_X1   g12687(.A1(new_n12880_), .A2(\a[46] ), .A3(\a[52] ), .ZN(new_n12881_));
  NAND2_X1   g12688(.A1(new_n12881_), .A2(new_n12879_), .ZN(new_n12882_));
  AOI22_X1   g12689(.A1(\a[39] ), .A2(\a[59] ), .B1(\a[40] ), .B2(\a[58] ), .ZN(new_n12883_));
  INV_X1     g12690(.I(new_n12883_), .ZN(new_n12884_));
  NOR2_X1    g12691(.A1(new_n3551_), .A2(new_n7206_), .ZN(new_n12885_));
  NOR2_X1    g12692(.A1(new_n4030_), .A2(new_n5425_), .ZN(new_n12886_));
  AOI21_X1   g12693(.A1(new_n12884_), .A2(new_n12886_), .B(new_n12885_), .ZN(new_n12887_));
  INV_X1     g12694(.I(new_n12887_), .ZN(new_n12888_));
  OAI21_X1   g12695(.A1(new_n12885_), .A2(new_n12883_), .B(new_n12886_), .ZN(new_n12889_));
  OAI21_X1   g12696(.A1(new_n12888_), .A2(new_n12883_), .B(new_n12889_), .ZN(new_n12890_));
  XNOR2_X1   g12697(.A1(new_n12882_), .A2(new_n12890_), .ZN(new_n12891_));
  XOR2_X1    g12698(.A1(new_n12891_), .A2(new_n12874_), .Z(new_n12892_));
  XOR2_X1    g12699(.A1(new_n12866_), .A2(new_n12892_), .Z(new_n12893_));
  INV_X1     g12700(.I(new_n12893_), .ZN(new_n12894_));
  NAND2_X1   g12701(.A1(new_n12823_), .A2(new_n12816_), .ZN(new_n12895_));
  NAND2_X1   g12702(.A1(new_n12824_), .A2(new_n12832_), .ZN(new_n12896_));
  NAND2_X1   g12703(.A1(new_n12896_), .A2(new_n12895_), .ZN(new_n12897_));
  NAND2_X1   g12704(.A1(new_n12705_), .A2(new_n12660_), .ZN(new_n12898_));
  NAND2_X1   g12705(.A1(new_n12794_), .A2(new_n12653_), .ZN(new_n12899_));
  NAND2_X1   g12706(.A1(new_n12899_), .A2(new_n12898_), .ZN(new_n12900_));
  NAND2_X1   g12707(.A1(new_n12721_), .A2(new_n12763_), .ZN(new_n12901_));
  NAND2_X1   g12708(.A1(new_n12764_), .A2(new_n12713_), .ZN(new_n12902_));
  NAND2_X1   g12709(.A1(new_n12902_), .A2(new_n12901_), .ZN(new_n12903_));
  XOR2_X1    g12710(.A1(new_n12900_), .A2(new_n12903_), .Z(new_n12904_));
  XOR2_X1    g12711(.A1(new_n12904_), .A2(new_n12897_), .Z(new_n12905_));
  NOR2_X1    g12712(.A1(new_n12894_), .A2(new_n12905_), .ZN(new_n12906_));
  INV_X1     g12713(.I(new_n12906_), .ZN(new_n12907_));
  NAND2_X1   g12714(.A1(new_n12894_), .A2(new_n12905_), .ZN(new_n12908_));
  NAND3_X1   g12715(.A1(new_n12856_), .A2(new_n12907_), .A3(new_n12908_), .ZN(new_n12909_));
  NAND2_X1   g12716(.A1(new_n12909_), .A2(new_n12908_), .ZN(new_n12910_));
  INV_X1     g12717(.I(new_n12910_), .ZN(new_n12911_));
  AOI22_X1   g12718(.A1(new_n12911_), .A2(new_n12907_), .B1(new_n12856_), .B2(new_n12909_), .ZN(new_n12912_));
  INV_X1     g12719(.I(new_n12912_), .ZN(new_n12913_));
  NAND2_X1   g12720(.A1(new_n12803_), .A2(new_n12772_), .ZN(new_n12914_));
  NAND2_X1   g12721(.A1(new_n12762_), .A2(new_n12804_), .ZN(new_n12915_));
  NAND2_X1   g12722(.A1(new_n12915_), .A2(new_n12914_), .ZN(new_n12916_));
  NOR2_X1    g12723(.A1(new_n12801_), .A2(new_n12798_), .ZN(new_n12917_));
  INV_X1     g12724(.I(new_n12917_), .ZN(new_n12918_));
  NOR2_X1    g12725(.A1(new_n4343_), .A2(new_n6129_), .ZN(new_n12919_));
  AOI22_X1   g12726(.A1(\a[43] ), .A2(\a[55] ), .B1(\a[44] ), .B2(\a[54] ), .ZN(new_n12920_));
  NOR2_X1    g12727(.A1(new_n12919_), .A2(new_n12920_), .ZN(new_n12921_));
  INV_X1     g12728(.I(new_n12921_), .ZN(new_n12922_));
  NOR2_X1    g12729(.A1(new_n2524_), .A2(new_n7643_), .ZN(new_n12923_));
  INV_X1     g12730(.I(new_n12923_), .ZN(new_n12924_));
  NOR2_X1    g12731(.A1(new_n12922_), .A2(new_n12924_), .ZN(new_n12925_));
  NOR2_X1    g12732(.A1(new_n12921_), .A2(new_n12923_), .ZN(new_n12926_));
  NOR2_X1    g12733(.A1(new_n12925_), .A2(new_n12926_), .ZN(new_n12927_));
  NOR2_X1    g12734(.A1(new_n12927_), .A2(new_n12780_), .ZN(new_n12928_));
  INV_X1     g12735(.I(new_n12927_), .ZN(new_n12929_));
  NOR2_X1    g12736(.A1(new_n12929_), .A2(new_n12779_), .ZN(new_n12930_));
  NOR2_X1    g12737(.A1(new_n12930_), .A2(new_n12928_), .ZN(new_n12931_));
  NOR2_X1    g12738(.A1(new_n2914_), .A2(new_n6723_), .ZN(new_n12932_));
  INV_X1     g12739(.I(new_n12932_), .ZN(new_n12933_));
  AOI22_X1   g12740(.A1(\a[41] ), .A2(\a[57] ), .B1(\a[42] ), .B2(\a[56] ), .ZN(new_n12934_));
  NOR2_X1    g12741(.A1(new_n4667_), .A2(new_n8161_), .ZN(new_n12935_));
  NOR3_X1    g12742(.A1(new_n12935_), .A2(new_n12933_), .A3(new_n12934_), .ZN(new_n12936_));
  NOR2_X1    g12743(.A1(new_n12936_), .A2(new_n12935_), .ZN(new_n12937_));
  INV_X1     g12744(.I(new_n12937_), .ZN(new_n12938_));
  OAI22_X1   g12745(.A1(new_n12938_), .A2(new_n12934_), .B1(new_n12933_), .B2(new_n12936_), .ZN(new_n12939_));
  INV_X1     g12746(.I(new_n12939_), .ZN(new_n12940_));
  XOR2_X1    g12747(.A1(new_n12931_), .A2(new_n12940_), .Z(new_n12941_));
  NAND2_X1   g12748(.A1(new_n12768_), .A2(new_n12770_), .ZN(new_n12942_));
  NAND2_X1   g12749(.A1(new_n12771_), .A2(new_n12765_), .ZN(new_n12943_));
  NAND2_X1   g12750(.A1(new_n12943_), .A2(new_n12942_), .ZN(new_n12944_));
  NOR2_X1    g12751(.A1(new_n12944_), .A2(new_n12941_), .ZN(new_n12945_));
  NAND2_X1   g12752(.A1(new_n12944_), .A2(new_n12941_), .ZN(new_n12946_));
  INV_X1     g12753(.I(new_n12946_), .ZN(new_n12947_));
  OAI21_X1   g12754(.A1(new_n12945_), .A2(new_n12947_), .B(new_n12918_), .ZN(new_n12948_));
  INV_X1     g12755(.I(new_n12948_), .ZN(new_n12949_));
  NOR3_X1    g12756(.A1(new_n12918_), .A2(new_n12945_), .A3(new_n12947_), .ZN(new_n12950_));
  NOR2_X1    g12757(.A1(new_n12949_), .A2(new_n12950_), .ZN(new_n12951_));
  NAND2_X1   g12758(.A1(new_n12916_), .A2(new_n12951_), .ZN(new_n12952_));
  NAND2_X1   g12759(.A1(new_n12952_), .A2(new_n12916_), .ZN(new_n12953_));
  NAND2_X1   g12760(.A1(new_n12952_), .A2(new_n12951_), .ZN(new_n12954_));
  NAND2_X1   g12761(.A1(new_n12953_), .A2(new_n12954_), .ZN(new_n12955_));
  NAND2_X1   g12762(.A1(new_n12955_), .A2(new_n12913_), .ZN(new_n12956_));
  NAND3_X1   g12763(.A1(new_n12953_), .A2(new_n12954_), .A3(new_n12912_), .ZN(new_n12957_));
  NAND2_X1   g12764(.A1(new_n12956_), .A2(new_n12957_), .ZN(new_n12958_));
  NOR2_X1    g12765(.A1(new_n12854_), .A2(new_n12958_), .ZN(new_n12959_));
  INV_X1     g12766(.I(new_n12959_), .ZN(new_n12960_));
  NAND2_X1   g12767(.A1(new_n12854_), .A2(new_n12958_), .ZN(new_n12961_));
  NAND2_X1   g12768(.A1(new_n12960_), .A2(new_n12961_), .ZN(new_n12962_));
  XOR2_X1    g12769(.A1(new_n12853_), .A2(new_n12962_), .Z(\asquared[99] ));
  OAI21_X1   g12770(.A1(new_n12852_), .A2(new_n12849_), .B(new_n12961_), .ZN(new_n12964_));
  NAND2_X1   g12771(.A1(new_n12964_), .A2(new_n12960_), .ZN(new_n12965_));
  INV_X1     g12772(.I(new_n12941_), .ZN(new_n12966_));
  NAND2_X1   g12773(.A1(new_n12944_), .A2(new_n12966_), .ZN(new_n12967_));
  NAND2_X1   g12774(.A1(new_n12948_), .A2(new_n12967_), .ZN(new_n12968_));
  NAND2_X1   g12775(.A1(new_n12873_), .A2(new_n12868_), .ZN(new_n12969_));
  XNOR2_X1   g12776(.A1(new_n12969_), .A2(new_n12937_), .ZN(new_n12970_));
  NAND2_X1   g12777(.A1(new_n6916_), .A2(new_n9030_), .ZN(new_n12971_));
  NAND2_X1   g12778(.A1(new_n2915_), .A2(new_n7852_), .ZN(new_n12972_));
  AOI22_X1   g12779(.A1(new_n12971_), .A2(new_n12972_), .B1(new_n4209_), .B2(new_n7453_), .ZN(new_n12973_));
  NAND2_X1   g12780(.A1(\a[36] ), .A2(\a[63] ), .ZN(new_n12974_));
  AOI22_X1   g12781(.A1(\a[38] ), .A2(\a[61] ), .B1(\a[39] ), .B2(\a[60] ), .ZN(new_n12975_));
  NAND2_X1   g12782(.A1(new_n4209_), .A2(new_n7453_), .ZN(new_n12976_));
  NAND3_X1   g12783(.A1(new_n12971_), .A2(new_n12972_), .A3(new_n12976_), .ZN(new_n12977_));
  OAI22_X1   g12784(.A1(new_n12973_), .A2(new_n12974_), .B1(new_n12977_), .B2(new_n12975_), .ZN(new_n12978_));
  XNOR2_X1   g12785(.A1(new_n12970_), .A2(new_n12978_), .ZN(new_n12979_));
  INV_X1     g12786(.I(new_n12874_), .ZN(new_n12980_));
  NAND2_X1   g12787(.A1(new_n12882_), .A2(new_n12890_), .ZN(new_n12981_));
  OAI21_X1   g12788(.A1(new_n12891_), .A2(new_n12980_), .B(new_n12981_), .ZN(new_n12982_));
  NOR2_X1    g12789(.A1(new_n12925_), .A2(new_n12919_), .ZN(new_n12983_));
  NAND2_X1   g12790(.A1(new_n12887_), .A2(new_n12878_), .ZN(new_n12984_));
  OAI21_X1   g12791(.A1(new_n12875_), .A2(new_n12877_), .B(new_n12888_), .ZN(new_n12985_));
  AND2_X2    g12792(.A1(new_n12985_), .A2(new_n12984_), .Z(new_n12986_));
  XNOR2_X1   g12793(.A1(new_n12986_), .A2(new_n12983_), .ZN(new_n12987_));
  NOR2_X1    g12794(.A1(new_n12987_), .A2(new_n12982_), .ZN(new_n12988_));
  NAND2_X1   g12795(.A1(new_n12987_), .A2(new_n12982_), .ZN(new_n12989_));
  INV_X1     g12796(.I(new_n12989_), .ZN(new_n12990_));
  NOR2_X1    g12797(.A1(new_n12990_), .A2(new_n12988_), .ZN(new_n12991_));
  XOR2_X1    g12798(.A1(new_n12991_), .A2(new_n12979_), .Z(new_n12992_));
  INV_X1     g12799(.I(new_n12992_), .ZN(new_n12993_));
  AOI21_X1   g12800(.A1(new_n12931_), .A2(new_n12939_), .B(new_n12930_), .ZN(new_n12994_));
  NOR2_X1    g12801(.A1(new_n4901_), .A2(new_n7144_), .ZN(new_n12995_));
  INV_X1     g12802(.I(new_n12995_), .ZN(new_n12996_));
  NOR2_X1    g12803(.A1(new_n12996_), .A2(new_n2752_), .ZN(new_n12997_));
  NAND2_X1   g12804(.A1(new_n12997_), .A2(new_n5154_), .ZN(new_n12998_));
  AOI21_X1   g12805(.A1(\a[37] ), .A2(\a[62] ), .B(\a[50] ), .ZN(new_n12999_));
  NOR2_X1    g12806(.A1(new_n12997_), .A2(new_n5154_), .ZN(new_n13000_));
  INV_X1     g12807(.I(new_n13000_), .ZN(new_n13001_));
  OAI21_X1   g12808(.A1(new_n13001_), .A2(new_n12999_), .B(new_n12998_), .ZN(new_n13002_));
  NAND2_X1   g12809(.A1(new_n12822_), .A2(new_n12814_), .ZN(new_n13003_));
  NAND2_X1   g12810(.A1(new_n12861_), .A2(new_n12831_), .ZN(new_n13004_));
  NAND2_X1   g12811(.A1(new_n13004_), .A2(new_n13003_), .ZN(new_n13005_));
  XNOR2_X1   g12812(.A1(new_n13005_), .A2(new_n13002_), .ZN(new_n13006_));
  XOR2_X1    g12813(.A1(new_n13006_), .A2(new_n12994_), .Z(new_n13007_));
  NOR2_X1    g12814(.A1(new_n12993_), .A2(new_n13007_), .ZN(new_n13008_));
  NAND2_X1   g12815(.A1(new_n12993_), .A2(new_n13007_), .ZN(new_n13009_));
  INV_X1     g12816(.I(new_n13009_), .ZN(new_n13010_));
  NOR2_X1    g12817(.A1(new_n13010_), .A2(new_n13008_), .ZN(new_n13011_));
  NOR2_X1    g12818(.A1(new_n12968_), .A2(new_n13011_), .ZN(new_n13012_));
  NAND2_X1   g12819(.A1(new_n12968_), .A2(new_n13011_), .ZN(new_n13013_));
  INV_X1     g12820(.I(new_n13013_), .ZN(new_n13014_));
  NOR2_X1    g12821(.A1(new_n13014_), .A2(new_n13012_), .ZN(new_n13015_));
  OAI21_X1   g12822(.A1(new_n12863_), .A2(new_n12892_), .B(new_n12864_), .ZN(new_n13016_));
  NAND2_X1   g12823(.A1(new_n12900_), .A2(new_n12903_), .ZN(new_n13017_));
  NAND2_X1   g12824(.A1(new_n12904_), .A2(new_n12897_), .ZN(new_n13018_));
  NAND2_X1   g12825(.A1(new_n13018_), .A2(new_n13017_), .ZN(new_n13019_));
  NOR4_X1    g12826(.A1(new_n3221_), .A2(new_n3859_), .A3(new_n5680_), .A4(new_n6548_), .ZN(new_n13020_));
  NOR2_X1    g12827(.A1(new_n5377_), .A2(new_n7206_), .ZN(new_n13021_));
  NOR2_X1    g12828(.A1(new_n13021_), .A2(new_n13020_), .ZN(new_n13022_));
  NOR2_X1    g12829(.A1(new_n3859_), .A2(new_n5680_), .ZN(new_n13023_));
  NOR2_X1    g12830(.A1(new_n3327_), .A2(new_n6316_), .ZN(new_n13024_));
  NAND2_X1   g12831(.A1(new_n13023_), .A2(new_n13024_), .ZN(new_n13025_));
  INV_X1     g12832(.I(new_n13025_), .ZN(new_n13026_));
  NOR2_X1    g12833(.A1(new_n13022_), .A2(new_n13026_), .ZN(new_n13027_));
  NOR3_X1    g12834(.A1(new_n13027_), .A2(new_n3221_), .A3(new_n6548_), .ZN(new_n13028_));
  INV_X1     g12835(.I(new_n13028_), .ZN(new_n13029_));
  NOR2_X1    g12836(.A1(new_n13027_), .A2(new_n13026_), .ZN(new_n13030_));
  OAI21_X1   g12837(.A1(new_n13023_), .A2(new_n13024_), .B(new_n13030_), .ZN(new_n13031_));
  AND2_X2    g12838(.A1(new_n13031_), .A2(new_n13029_), .Z(new_n13032_));
  NAND2_X1   g12839(.A1(new_n4720_), .A2(new_n5862_), .ZN(new_n13033_));
  OAI22_X1   g12840(.A1(new_n4314_), .A2(new_n8421_), .B1(new_n4430_), .B2(new_n6127_), .ZN(new_n13034_));
  NAND2_X1   g12841(.A1(new_n13034_), .A2(new_n13033_), .ZN(new_n13035_));
  NAND3_X1   g12842(.A1(new_n13035_), .A2(\a[45] ), .A3(\a[54] ), .ZN(new_n13036_));
  AOI22_X1   g12843(.A1(\a[46] ), .A2(\a[53] ), .B1(\a[47] ), .B2(\a[52] ), .ZN(new_n13037_));
  NAND2_X1   g12844(.A1(new_n13035_), .A2(new_n13033_), .ZN(new_n13038_));
  OAI21_X1   g12845(.A1(new_n13037_), .A2(new_n13038_), .B(new_n13036_), .ZN(new_n13039_));
  XOR2_X1    g12846(.A1(new_n13032_), .A2(new_n13039_), .Z(new_n13040_));
  NOR2_X1    g12847(.A1(new_n4596_), .A2(new_n5135_), .ZN(new_n13041_));
  INV_X1     g12848(.I(new_n13041_), .ZN(new_n13042_));
  AOI22_X1   g12849(.A1(\a[42] ), .A2(\a[57] ), .B1(\a[43] ), .B2(\a[56] ), .ZN(new_n13043_));
  NOR2_X1    g12850(.A1(new_n4181_), .A2(new_n8161_), .ZN(new_n13044_));
  NOR3_X1    g12851(.A1(new_n13044_), .A2(new_n13042_), .A3(new_n13043_), .ZN(new_n13045_));
  NOR2_X1    g12852(.A1(new_n13045_), .A2(new_n13044_), .ZN(new_n13046_));
  INV_X1     g12853(.I(new_n13046_), .ZN(new_n13047_));
  OAI22_X1   g12854(.A1(new_n13047_), .A2(new_n13043_), .B1(new_n13042_), .B2(new_n13045_), .ZN(new_n13048_));
  XOR2_X1    g12855(.A1(new_n13040_), .A2(new_n13048_), .Z(new_n13049_));
  INV_X1     g12856(.I(new_n13049_), .ZN(new_n13050_));
  XOR2_X1    g12857(.A1(new_n13019_), .A2(new_n13050_), .Z(new_n13051_));
  XOR2_X1    g12858(.A1(new_n13051_), .A2(new_n13016_), .Z(new_n13052_));
  NAND2_X1   g12859(.A1(new_n12911_), .A2(new_n13052_), .ZN(new_n13053_));
  NAND2_X1   g12860(.A1(new_n12910_), .A2(new_n13052_), .ZN(new_n13054_));
  NAND2_X1   g12861(.A1(new_n13054_), .A2(new_n12910_), .ZN(new_n13055_));
  NAND2_X1   g12862(.A1(new_n13055_), .A2(new_n13053_), .ZN(new_n13056_));
  AOI21_X1   g12863(.A1(new_n13054_), .A2(new_n12910_), .B(new_n13015_), .ZN(new_n13057_));
  AOI22_X1   g12864(.A1(new_n13056_), .A2(new_n13015_), .B1(new_n13053_), .B2(new_n13057_), .ZN(new_n13058_));
  NAND2_X1   g12865(.A1(new_n12956_), .A2(new_n12952_), .ZN(new_n13059_));
  NAND2_X1   g12866(.A1(new_n13059_), .A2(new_n13058_), .ZN(new_n13060_));
  INV_X1     g12867(.I(new_n13060_), .ZN(new_n13061_));
  NOR2_X1    g12868(.A1(new_n13059_), .A2(new_n13058_), .ZN(new_n13062_));
  NOR2_X1    g12869(.A1(new_n13061_), .A2(new_n13062_), .ZN(new_n13063_));
  XOR2_X1    g12870(.A1(new_n12965_), .A2(new_n13063_), .Z(\asquared[100] ));
  AOI21_X1   g12871(.A1(new_n12964_), .A2(new_n12960_), .B(new_n13062_), .ZN(new_n13065_));
  NOR2_X1    g12872(.A1(new_n13065_), .A2(new_n13061_), .ZN(new_n13066_));
  NAND2_X1   g12873(.A1(new_n13056_), .A2(new_n13015_), .ZN(new_n13067_));
  NAND2_X1   g12874(.A1(new_n13067_), .A2(new_n13054_), .ZN(new_n13068_));
  AOI21_X1   g12875(.A1(\a[37] ), .A2(\a[63] ), .B(new_n13001_), .ZN(new_n13069_));
  NOR3_X1    g12876(.A1(new_n13000_), .A2(new_n2752_), .A3(new_n7643_), .ZN(new_n13070_));
  NOR2_X1    g12877(.A1(new_n13069_), .A2(new_n13070_), .ZN(new_n13071_));
  NOR2_X1    g12878(.A1(new_n13071_), .A2(new_n13047_), .ZN(new_n13072_));
  INV_X1     g12879(.I(new_n13071_), .ZN(new_n13073_));
  NOR2_X1    g12880(.A1(new_n13073_), .A2(new_n13046_), .ZN(new_n13074_));
  NOR2_X1    g12881(.A1(new_n13074_), .A2(new_n13072_), .ZN(new_n13075_));
  INV_X1     g12882(.I(new_n13030_), .ZN(new_n13076_));
  XOR2_X1    g12883(.A1(new_n13038_), .A2(new_n12977_), .Z(new_n13077_));
  XOR2_X1    g12884(.A1(new_n13077_), .A2(new_n13076_), .Z(new_n13078_));
  INV_X1     g12885(.I(new_n13032_), .ZN(new_n13079_));
  NAND2_X1   g12886(.A1(new_n13079_), .A2(new_n13039_), .ZN(new_n13080_));
  INV_X1     g12887(.I(new_n13048_), .ZN(new_n13081_));
  OAI21_X1   g12888(.A1(new_n13040_), .A2(new_n13081_), .B(new_n13080_), .ZN(new_n13082_));
  NAND2_X1   g12889(.A1(new_n13082_), .A2(new_n13078_), .ZN(new_n13083_));
  INV_X1     g12890(.I(new_n13083_), .ZN(new_n13084_));
  NOR2_X1    g12891(.A1(new_n13082_), .A2(new_n13078_), .ZN(new_n13085_));
  NOR2_X1    g12892(.A1(new_n13084_), .A2(new_n13085_), .ZN(new_n13086_));
  NOR2_X1    g12893(.A1(new_n13086_), .A2(new_n13075_), .ZN(new_n13087_));
  NAND2_X1   g12894(.A1(new_n13086_), .A2(new_n13075_), .ZN(new_n13088_));
  INV_X1     g12895(.I(new_n13088_), .ZN(new_n13089_));
  NOR2_X1    g12896(.A1(new_n13089_), .A2(new_n13087_), .ZN(new_n13090_));
  NAND2_X1   g12897(.A1(new_n13019_), .A2(new_n13050_), .ZN(new_n13091_));
  NAND2_X1   g12898(.A1(new_n13051_), .A2(new_n13016_), .ZN(new_n13092_));
  NAND2_X1   g12899(.A1(new_n13092_), .A2(new_n13091_), .ZN(new_n13093_));
  NAND2_X1   g12900(.A1(new_n12938_), .A2(new_n12969_), .ZN(new_n13094_));
  NAND2_X1   g12901(.A1(new_n12970_), .A2(new_n12978_), .ZN(new_n13095_));
  NAND2_X1   g12902(.A1(new_n13095_), .A2(new_n13094_), .ZN(new_n13096_));
  INV_X1     g12903(.I(new_n12986_), .ZN(new_n13097_));
  OAI21_X1   g12904(.A1(new_n13097_), .A2(new_n12983_), .B(new_n12985_), .ZN(new_n13098_));
  NOR2_X1    g12905(.A1(new_n4981_), .A2(new_n5525_), .ZN(new_n13099_));
  AOI22_X1   g12906(.A1(new_n4976_), .A2(new_n5862_), .B1(new_n4978_), .B2(new_n5682_), .ZN(new_n13100_));
  NOR2_X1    g12907(.A1(new_n13099_), .A2(new_n13100_), .ZN(new_n13101_));
  NOR2_X1    g12908(.A1(new_n13101_), .A2(new_n13099_), .ZN(new_n13102_));
  INV_X1     g12909(.I(new_n13102_), .ZN(new_n13103_));
  AOI21_X1   g12910(.A1(\a[48] ), .A2(\a[52] ), .B(new_n7867_), .ZN(new_n13104_));
  NAND2_X1   g12911(.A1(\a[47] ), .A2(\a[53] ), .ZN(new_n13105_));
  OAI22_X1   g12912(.A1(new_n13103_), .A2(new_n13104_), .B1(new_n13101_), .B2(new_n13105_), .ZN(new_n13106_));
  XNOR2_X1   g12913(.A1(new_n13098_), .A2(new_n13106_), .ZN(new_n13107_));
  XNOR2_X1   g12914(.A1(new_n13107_), .A2(new_n13096_), .ZN(new_n13108_));
  XOR2_X1    g12915(.A1(new_n13093_), .A2(new_n13108_), .Z(new_n13109_));
  OR2_X2     g12916(.A1(new_n13109_), .A2(new_n13090_), .Z(new_n13110_));
  NAND2_X1   g12917(.A1(new_n13109_), .A2(new_n13090_), .ZN(new_n13111_));
  AND2_X2    g12918(.A1(new_n13110_), .A2(new_n13111_), .Z(new_n13112_));
  NOR2_X1    g12919(.A1(new_n13014_), .A2(new_n13010_), .ZN(new_n13113_));
  OAI21_X1   g12920(.A1(new_n12979_), .A2(new_n12988_), .B(new_n12989_), .ZN(new_n13114_));
  OAI22_X1   g12921(.A1(new_n4210_), .A2(new_n7591_), .B1(new_n10435_), .B2(new_n12933_), .ZN(new_n13115_));
  OAI21_X1   g12922(.A1(new_n3551_), .A2(new_n7454_), .B(new_n13115_), .ZN(new_n13116_));
  INV_X1     g12923(.I(new_n13116_), .ZN(new_n13117_));
  AOI22_X1   g12924(.A1(\a[39] ), .A2(\a[61] ), .B1(\a[40] ), .B2(\a[60] ), .ZN(new_n13118_));
  NOR2_X1    g12925(.A1(new_n3551_), .A2(new_n7454_), .ZN(new_n13119_));
  NOR2_X1    g12926(.A1(new_n13115_), .A2(new_n13119_), .ZN(new_n13120_));
  INV_X1     g12927(.I(new_n13120_), .ZN(new_n13121_));
  OAI22_X1   g12928(.A1(new_n13117_), .A2(new_n9705_), .B1(new_n13118_), .B2(new_n13121_), .ZN(new_n13122_));
  NOR2_X1    g12929(.A1(new_n4704_), .A2(new_n7185_), .ZN(new_n13123_));
  AOI22_X1   g12930(.A1(new_n4033_), .A2(new_n8951_), .B1(new_n4342_), .B2(new_n6494_), .ZN(new_n13124_));
  NOR2_X1    g12931(.A1(new_n13123_), .A2(new_n13124_), .ZN(new_n13125_));
  AOI22_X1   g12932(.A1(\a[44] ), .A2(\a[56] ), .B1(\a[45] ), .B2(\a[55] ), .ZN(new_n13126_));
  NOR2_X1    g12933(.A1(new_n13125_), .A2(new_n13123_), .ZN(new_n13127_));
  INV_X1     g12934(.I(new_n13127_), .ZN(new_n13128_));
  OAI22_X1   g12935(.A1(new_n13128_), .A2(new_n13126_), .B1(new_n8078_), .B2(new_n13125_), .ZN(new_n13129_));
  XNOR2_X1   g12936(.A1(new_n13122_), .A2(new_n13129_), .ZN(new_n13130_));
  AOI22_X1   g12937(.A1(\a[41] ), .A2(\a[59] ), .B1(\a[42] ), .B2(\a[58] ), .ZN(new_n13131_));
  NOR2_X1    g12938(.A1(new_n4667_), .A2(new_n7206_), .ZN(new_n13132_));
  NOR3_X1    g12939(.A1(new_n13132_), .A2(new_n7396_), .A3(new_n13131_), .ZN(new_n13133_));
  NOR2_X1    g12940(.A1(new_n13133_), .A2(new_n13132_), .ZN(new_n13134_));
  INV_X1     g12941(.I(new_n13134_), .ZN(new_n13135_));
  OAI22_X1   g12942(.A1(new_n13135_), .A2(new_n13131_), .B1(new_n7396_), .B2(new_n13133_), .ZN(new_n13136_));
  INV_X1     g12943(.I(new_n13136_), .ZN(new_n13137_));
  XOR2_X1    g12944(.A1(new_n13130_), .A2(new_n13137_), .Z(new_n13138_));
  NAND2_X1   g12945(.A1(new_n13005_), .A2(new_n13002_), .ZN(new_n13139_));
  OAI21_X1   g12946(.A1(new_n13006_), .A2(new_n12994_), .B(new_n13139_), .ZN(new_n13140_));
  NOR2_X1    g12947(.A1(new_n13140_), .A2(new_n13138_), .ZN(new_n13141_));
  NAND2_X1   g12948(.A1(new_n13140_), .A2(new_n13138_), .ZN(new_n13142_));
  INV_X1     g12949(.I(new_n13142_), .ZN(new_n13143_));
  NOR2_X1    g12950(.A1(new_n13143_), .A2(new_n13141_), .ZN(new_n13144_));
  NOR2_X1    g12951(.A1(new_n13144_), .A2(new_n13114_), .ZN(new_n13145_));
  NAND2_X1   g12952(.A1(new_n13144_), .A2(new_n13114_), .ZN(new_n13146_));
  INV_X1     g12953(.I(new_n13146_), .ZN(new_n13147_));
  NOR2_X1    g12954(.A1(new_n13147_), .A2(new_n13145_), .ZN(new_n13148_));
  INV_X1     g12955(.I(new_n13148_), .ZN(new_n13149_));
  NAND2_X1   g12956(.A1(new_n13113_), .A2(new_n13149_), .ZN(new_n13150_));
  NOR2_X1    g12957(.A1(new_n13113_), .A2(new_n13149_), .ZN(new_n13151_));
  INV_X1     g12958(.I(new_n13151_), .ZN(new_n13152_));
  AND2_X2    g12959(.A1(new_n13152_), .A2(new_n13150_), .Z(new_n13153_));
  AND2_X2    g12960(.A1(new_n13153_), .A2(new_n13112_), .Z(new_n13154_));
  NOR2_X1    g12961(.A1(new_n13153_), .A2(new_n13112_), .ZN(new_n13155_));
  NOR2_X1    g12962(.A1(new_n13154_), .A2(new_n13155_), .ZN(new_n13156_));
  NAND2_X1   g12963(.A1(new_n13156_), .A2(new_n13068_), .ZN(new_n13157_));
  NOR2_X1    g12964(.A1(new_n13156_), .A2(new_n13068_), .ZN(new_n13158_));
  INV_X1     g12965(.I(new_n13158_), .ZN(new_n13159_));
  NAND2_X1   g12966(.A1(new_n13159_), .A2(new_n13157_), .ZN(new_n13160_));
  INV_X1     g12967(.I(new_n12847_), .ZN(new_n13161_));
  OAI21_X1   g12968(.A1(new_n12753_), .A2(new_n12742_), .B(new_n13161_), .ZN(new_n13162_));
  INV_X1     g12969(.I(new_n12961_), .ZN(new_n13163_));
  AOI21_X1   g12970(.A1(new_n13162_), .A2(new_n12848_), .B(new_n13163_), .ZN(new_n13164_));
  INV_X1     g12971(.I(new_n13062_), .ZN(new_n13165_));
  OAI21_X1   g12972(.A1(new_n13164_), .A2(new_n12959_), .B(new_n13165_), .ZN(new_n13166_));
  AOI21_X1   g12973(.A1(new_n13166_), .A2(new_n13060_), .B(new_n13158_), .ZN(new_n13167_));
  AOI22_X1   g12974(.A1(new_n13167_), .A2(new_n13157_), .B1(new_n13066_), .B2(new_n13160_), .ZN(\asquared[101] ));
  OAI21_X1   g12975(.A1(new_n13065_), .A2(new_n13061_), .B(new_n13159_), .ZN(new_n13169_));
  NAND2_X1   g12976(.A1(new_n13169_), .A2(new_n13157_), .ZN(new_n13170_));
  NOR2_X1    g12977(.A1(new_n13154_), .A2(new_n13151_), .ZN(new_n13171_));
  INV_X1     g12978(.I(new_n13171_), .ZN(new_n13172_));
  NOR2_X1    g12979(.A1(new_n13147_), .A2(new_n13143_), .ZN(new_n13173_));
  NOR2_X1    g12980(.A1(new_n13089_), .A2(new_n13084_), .ZN(new_n13174_));
  XNOR2_X1   g12981(.A1(new_n13173_), .A2(new_n13174_), .ZN(new_n13175_));
  NOR2_X1    g12982(.A1(new_n13135_), .A2(new_n13121_), .ZN(new_n13176_));
  NOR2_X1    g12983(.A1(new_n13134_), .A2(new_n13120_), .ZN(new_n13177_));
  NOR2_X1    g12984(.A1(new_n13176_), .A2(new_n13177_), .ZN(new_n13178_));
  INV_X1     g12985(.I(new_n13178_), .ZN(new_n13179_));
  NOR2_X1    g12986(.A1(new_n13179_), .A2(new_n13127_), .ZN(new_n13180_));
  NOR2_X1    g12987(.A1(new_n13178_), .A2(new_n13128_), .ZN(new_n13181_));
  NOR2_X1    g12988(.A1(new_n13180_), .A2(new_n13181_), .ZN(new_n13182_));
  NAND2_X1   g12989(.A1(new_n13122_), .A2(new_n13129_), .ZN(new_n13183_));
  OAI21_X1   g12990(.A1(new_n13130_), .A2(new_n13137_), .B(new_n13183_), .ZN(new_n13184_));
  NAND2_X1   g12991(.A1(new_n13038_), .A2(new_n12977_), .ZN(new_n13185_));
  NAND2_X1   g12992(.A1(new_n13077_), .A2(new_n13076_), .ZN(new_n13186_));
  NAND2_X1   g12993(.A1(new_n13186_), .A2(new_n13185_), .ZN(new_n13187_));
  XOR2_X1    g12994(.A1(new_n13184_), .A2(new_n13187_), .Z(new_n13188_));
  XOR2_X1    g12995(.A1(new_n13188_), .A2(new_n13182_), .Z(new_n13189_));
  XOR2_X1    g12996(.A1(new_n13175_), .A2(new_n13189_), .Z(new_n13190_));
  INV_X1     g12997(.I(new_n13190_), .ZN(new_n13191_));
  NAND2_X1   g12998(.A1(new_n13093_), .A2(new_n13108_), .ZN(new_n13192_));
  NAND2_X1   g12999(.A1(new_n13111_), .A2(new_n13192_), .ZN(new_n13193_));
  AOI21_X1   g13000(.A1(\a[39] ), .A2(\a[62] ), .B(\a[51] ), .ZN(new_n13194_));
  OAI21_X1   g13001(.A1(new_n7144_), .A2(new_n11997_), .B(new_n5440_), .ZN(new_n13195_));
  NAND3_X1   g13002(.A1(new_n5439_), .A2(new_n6114_), .A3(\a[62] ), .ZN(new_n13196_));
  OAI21_X1   g13003(.A1(new_n13195_), .A2(new_n13194_), .B(new_n13196_), .ZN(new_n13197_));
  NOR2_X1    g13004(.A1(new_n5377_), .A2(new_n7454_), .ZN(new_n13198_));
  INV_X1     g13005(.I(new_n13198_), .ZN(new_n13199_));
  NOR2_X1    g13006(.A1(new_n3327_), .A2(new_n6723_), .ZN(new_n13200_));
  NOR2_X1    g13007(.A1(new_n3221_), .A2(new_n6897_), .ZN(new_n13201_));
  OAI21_X1   g13008(.A1(new_n13200_), .A2(new_n13201_), .B(new_n13199_), .ZN(new_n13202_));
  XNOR2_X1   g13009(.A1(new_n13202_), .A2(new_n13102_), .ZN(new_n13203_));
  XOR2_X1    g13010(.A1(new_n13203_), .A2(new_n13197_), .Z(new_n13204_));
  NOR2_X1    g13011(.A1(new_n13074_), .A2(new_n13070_), .ZN(new_n13205_));
  XNOR2_X1   g13012(.A1(new_n13204_), .A2(new_n13205_), .ZN(new_n13206_));
  INV_X1     g13013(.I(new_n13206_), .ZN(new_n13207_));
  NAND2_X1   g13014(.A1(new_n13098_), .A2(new_n13106_), .ZN(new_n13208_));
  INV_X1     g13015(.I(new_n13107_), .ZN(new_n13209_));
  NAND2_X1   g13016(.A1(new_n13209_), .A2(new_n13096_), .ZN(new_n13210_));
  NAND2_X1   g13017(.A1(new_n13210_), .A2(new_n13208_), .ZN(new_n13211_));
  AOI22_X1   g13018(.A1(\a[46] ), .A2(\a[55] ), .B1(\a[47] ), .B2(\a[54] ), .ZN(new_n13212_));
  NOR2_X1    g13019(.A1(new_n2914_), .A2(new_n7643_), .ZN(new_n13213_));
  INV_X1     g13020(.I(new_n13213_), .ZN(new_n13214_));
  OAI22_X1   g13021(.A1(new_n4721_), .A2(new_n6129_), .B1(new_n13214_), .B2(new_n13212_), .ZN(new_n13215_));
  NOR2_X1    g13022(.A1(new_n4721_), .A2(new_n6129_), .ZN(new_n13216_));
  OAI21_X1   g13023(.A1(new_n13216_), .A2(new_n13212_), .B(new_n13213_), .ZN(new_n13217_));
  OAI21_X1   g13024(.A1(new_n13215_), .A2(new_n13212_), .B(new_n13217_), .ZN(new_n13218_));
  NOR2_X1    g13025(.A1(new_n4034_), .A2(new_n6318_), .ZN(new_n13219_));
  NAND2_X1   g13026(.A1(\a[42] ), .A2(\a[45] ), .ZN(new_n13220_));
  NOR2_X1    g13027(.A1(new_n10715_), .A2(new_n13220_), .ZN(new_n13221_));
  NOR2_X1    g13028(.A1(new_n4181_), .A2(new_n7206_), .ZN(new_n13222_));
  NOR2_X1    g13029(.A1(new_n13222_), .A2(new_n13221_), .ZN(new_n13223_));
  NOR2_X1    g13030(.A1(new_n13223_), .A2(new_n13219_), .ZN(new_n13224_));
  NAND2_X1   g13031(.A1(\a[42] ), .A2(\a[59] ), .ZN(new_n13225_));
  AOI22_X1   g13032(.A1(\a[43] ), .A2(\a[58] ), .B1(\a[45] ), .B2(\a[56] ), .ZN(new_n13226_));
  NOR2_X1    g13033(.A1(new_n13224_), .A2(new_n13219_), .ZN(new_n13227_));
  INV_X1     g13034(.I(new_n13227_), .ZN(new_n13228_));
  OAI22_X1   g13035(.A1(new_n13228_), .A2(new_n13226_), .B1(new_n13224_), .B2(new_n13225_), .ZN(new_n13229_));
  XOR2_X1    g13036(.A1(new_n13229_), .A2(new_n13218_), .Z(new_n13230_));
  INV_X1     g13037(.I(new_n8250_), .ZN(new_n13231_));
  NOR2_X1    g13038(.A1(new_n7013_), .A2(new_n9657_), .ZN(new_n13232_));
  NAND3_X1   g13039(.A1(new_n8250_), .A2(\a[44] ), .A3(\a[57] ), .ZN(new_n13233_));
  NAND2_X1   g13040(.A1(new_n4980_), .A2(new_n5862_), .ZN(new_n13234_));
  AOI21_X1   g13041(.A1(new_n13234_), .A2(new_n13233_), .B(new_n13232_), .ZN(new_n13235_));
  AOI22_X1   g13042(.A1(\a[44] ), .A2(\a[57] ), .B1(\a[49] ), .B2(\a[52] ), .ZN(new_n13236_));
  OR2_X2     g13043(.A1(new_n13235_), .A2(new_n13232_), .Z(new_n13237_));
  OAI22_X1   g13044(.A1(new_n13237_), .A2(new_n13236_), .B1(new_n13231_), .B2(new_n13235_), .ZN(new_n13238_));
  XNOR2_X1   g13045(.A1(new_n13230_), .A2(new_n13238_), .ZN(new_n13239_));
  INV_X1     g13046(.I(new_n13239_), .ZN(new_n13240_));
  XOR2_X1    g13047(.A1(new_n13211_), .A2(new_n13240_), .Z(new_n13241_));
  XOR2_X1    g13048(.A1(new_n13241_), .A2(new_n13207_), .Z(new_n13242_));
  XNOR2_X1   g13049(.A1(new_n13193_), .A2(new_n13242_), .ZN(new_n13243_));
  XOR2_X1    g13050(.A1(new_n13243_), .A2(new_n13191_), .Z(new_n13244_));
  INV_X1     g13051(.I(new_n13244_), .ZN(new_n13245_));
  NOR2_X1    g13052(.A1(new_n13172_), .A2(new_n13245_), .ZN(new_n13246_));
  NOR2_X1    g13053(.A1(new_n13171_), .A2(new_n13244_), .ZN(new_n13247_));
  NOR2_X1    g13054(.A1(new_n13246_), .A2(new_n13247_), .ZN(new_n13248_));
  XOR2_X1    g13055(.A1(new_n13170_), .A2(new_n13248_), .Z(\asquared[102] ));
  NAND2_X1   g13056(.A1(new_n13193_), .A2(new_n13242_), .ZN(new_n13250_));
  OAI21_X1   g13057(.A1(new_n13243_), .A2(new_n13190_), .B(new_n13250_), .ZN(new_n13251_));
  INV_X1     g13058(.I(new_n13251_), .ZN(new_n13252_));
  NAND2_X1   g13059(.A1(new_n13229_), .A2(new_n13218_), .ZN(new_n13253_));
  NAND2_X1   g13060(.A1(new_n13230_), .A2(new_n13238_), .ZN(new_n13254_));
  NAND2_X1   g13061(.A1(new_n13254_), .A2(new_n13253_), .ZN(new_n13255_));
  XOR2_X1    g13062(.A1(new_n13237_), .A2(new_n13195_), .Z(new_n13256_));
  XOR2_X1    g13063(.A1(new_n13256_), .A2(new_n13215_), .Z(new_n13257_));
  NOR2_X1    g13064(.A1(new_n13180_), .A2(new_n13177_), .ZN(new_n13258_));
  INV_X1     g13065(.I(new_n13258_), .ZN(new_n13259_));
  NAND2_X1   g13066(.A1(new_n13259_), .A2(new_n13257_), .ZN(new_n13260_));
  INV_X1     g13067(.I(new_n13260_), .ZN(new_n13261_));
  NOR2_X1    g13068(.A1(new_n13259_), .A2(new_n13257_), .ZN(new_n13262_));
  NOR2_X1    g13069(.A1(new_n13261_), .A2(new_n13262_), .ZN(new_n13263_));
  NOR2_X1    g13070(.A1(new_n13263_), .A2(new_n13255_), .ZN(new_n13264_));
  NAND2_X1   g13071(.A1(new_n13263_), .A2(new_n13255_), .ZN(new_n13265_));
  INV_X1     g13072(.I(new_n13265_), .ZN(new_n13266_));
  NOR2_X1    g13073(.A1(new_n13266_), .A2(new_n13264_), .ZN(new_n13267_));
  INV_X1     g13074(.I(new_n13267_), .ZN(new_n13268_));
  NAND2_X1   g13075(.A1(new_n13184_), .A2(new_n13187_), .ZN(new_n13269_));
  NAND2_X1   g13076(.A1(new_n13188_), .A2(new_n13182_), .ZN(new_n13270_));
  NAND2_X1   g13077(.A1(new_n13270_), .A2(new_n13269_), .ZN(new_n13271_));
  NAND2_X1   g13078(.A1(new_n13211_), .A2(new_n13240_), .ZN(new_n13272_));
  NAND2_X1   g13079(.A1(new_n13241_), .A2(new_n13207_), .ZN(new_n13273_));
  NAND2_X1   g13080(.A1(new_n13273_), .A2(new_n13272_), .ZN(new_n13274_));
  XNOR2_X1   g13081(.A1(new_n13274_), .A2(new_n13271_), .ZN(new_n13275_));
  NAND2_X1   g13082(.A1(new_n13275_), .A2(new_n13268_), .ZN(new_n13276_));
  NOR2_X1    g13083(.A1(new_n13275_), .A2(new_n13268_), .ZN(new_n13277_));
  INV_X1     g13084(.I(new_n13277_), .ZN(new_n13278_));
  AND2_X2    g13085(.A1(new_n13278_), .A2(new_n13276_), .Z(new_n13279_));
  NOR2_X1    g13086(.A1(new_n13173_), .A2(new_n13174_), .ZN(new_n13280_));
  INV_X1     g13087(.I(new_n13175_), .ZN(new_n13281_));
  AOI21_X1   g13088(.A1(new_n13281_), .A2(new_n13189_), .B(new_n13280_), .ZN(new_n13282_));
  NOR2_X1    g13089(.A1(new_n4721_), .A2(new_n7185_), .ZN(new_n13283_));
  NOR2_X1    g13090(.A1(new_n4430_), .A2(new_n8161_), .ZN(new_n13284_));
  NOR2_X1    g13091(.A1(new_n4314_), .A2(new_n8952_), .ZN(new_n13285_));
  NOR2_X1    g13092(.A1(new_n13284_), .A2(new_n13285_), .ZN(new_n13286_));
  NOR2_X1    g13093(.A1(new_n13286_), .A2(new_n13283_), .ZN(new_n13287_));
  NAND2_X1   g13094(.A1(\a[45] ), .A2(\a[57] ), .ZN(new_n13288_));
  AOI22_X1   g13095(.A1(\a[46] ), .A2(\a[56] ), .B1(\a[47] ), .B2(\a[55] ), .ZN(new_n13289_));
  NOR2_X1    g13096(.A1(new_n13287_), .A2(new_n13283_), .ZN(new_n13290_));
  INV_X1     g13097(.I(new_n13290_), .ZN(new_n13291_));
  OAI22_X1   g13098(.A1(new_n13291_), .A2(new_n13289_), .B1(new_n13287_), .B2(new_n13288_), .ZN(new_n13292_));
  AOI22_X1   g13099(.A1(\a[43] ), .A2(\a[59] ), .B1(\a[44] ), .B2(\a[58] ), .ZN(new_n13293_));
  NOR2_X1    g13100(.A1(new_n4343_), .A2(new_n7206_), .ZN(new_n13294_));
  OAI21_X1   g13101(.A1(new_n13294_), .A2(new_n13293_), .B(new_n10434_), .ZN(new_n13295_));
  INV_X1     g13102(.I(new_n13293_), .ZN(new_n13296_));
  AOI21_X1   g13103(.A1(new_n10434_), .A2(new_n13296_), .B(new_n13294_), .ZN(new_n13297_));
  INV_X1     g13104(.I(new_n13297_), .ZN(new_n13298_));
  OAI21_X1   g13105(.A1(new_n13298_), .A2(new_n13293_), .B(new_n13295_), .ZN(new_n13299_));
  XOR2_X1    g13106(.A1(new_n13292_), .A2(new_n13299_), .Z(new_n13300_));
  NAND2_X1   g13107(.A1(new_n4980_), .A2(new_n6126_), .ZN(new_n13301_));
  NAND2_X1   g13108(.A1(new_n4902_), .A2(new_n8420_), .ZN(new_n13302_));
  AOI22_X1   g13109(.A1(new_n13301_), .A2(new_n13302_), .B1(new_n5154_), .B2(new_n5862_), .ZN(new_n13303_));
  NAND2_X1   g13110(.A1(new_n5154_), .A2(new_n5862_), .ZN(new_n13304_));
  NAND3_X1   g13111(.A1(new_n13304_), .A2(new_n13301_), .A3(new_n13302_), .ZN(new_n13305_));
  AOI21_X1   g13112(.A1(\a[49] ), .A2(\a[53] ), .B(new_n5522_), .ZN(new_n13306_));
  NAND2_X1   g13113(.A1(\a[48] ), .A2(\a[54] ), .ZN(new_n13307_));
  OAI22_X1   g13114(.A1(new_n13303_), .A2(new_n13307_), .B1(new_n13305_), .B2(new_n13306_), .ZN(new_n13308_));
  XNOR2_X1   g13115(.A1(new_n13300_), .A2(new_n13308_), .ZN(new_n13309_));
  OAI21_X1   g13116(.A1(new_n13202_), .A2(new_n13102_), .B(new_n13199_), .ZN(new_n13310_));
  NOR2_X1    g13117(.A1(new_n13228_), .A2(new_n13310_), .ZN(new_n13311_));
  INV_X1     g13118(.I(new_n13310_), .ZN(new_n13312_));
  NOR2_X1    g13119(.A1(new_n13312_), .A2(new_n13227_), .ZN(new_n13313_));
  NOR2_X1    g13120(.A1(new_n13313_), .A2(new_n13311_), .ZN(new_n13314_));
  NAND3_X1   g13121(.A1(new_n9030_), .A2(\a[39] ), .A3(\a[42] ), .ZN(new_n13315_));
  NAND2_X1   g13122(.A1(new_n3328_), .A2(new_n7852_), .ZN(new_n13316_));
  AOI22_X1   g13123(.A1(new_n13316_), .A2(new_n13315_), .B1(new_n4372_), .B2(new_n7453_), .ZN(new_n13317_));
  NAND2_X1   g13124(.A1(\a[39] ), .A2(\a[63] ), .ZN(new_n13318_));
  AOI22_X1   g13125(.A1(\a[41] ), .A2(\a[61] ), .B1(\a[42] ), .B2(\a[60] ), .ZN(new_n13319_));
  NAND2_X1   g13126(.A1(new_n4372_), .A2(new_n7453_), .ZN(new_n13320_));
  NAND3_X1   g13127(.A1(new_n13320_), .A2(new_n13316_), .A3(new_n13315_), .ZN(new_n13321_));
  OAI22_X1   g13128(.A1(new_n13317_), .A2(new_n13318_), .B1(new_n13321_), .B2(new_n13319_), .ZN(new_n13322_));
  XOR2_X1    g13129(.A1(new_n13314_), .A2(new_n13322_), .Z(new_n13323_));
  INV_X1     g13130(.I(new_n13203_), .ZN(new_n13324_));
  NAND2_X1   g13131(.A1(new_n13324_), .A2(new_n13197_), .ZN(new_n13325_));
  OAI21_X1   g13132(.A1(new_n13204_), .A2(new_n13205_), .B(new_n13325_), .ZN(new_n13326_));
  XOR2_X1    g13133(.A1(new_n13323_), .A2(new_n13326_), .Z(new_n13327_));
  XNOR2_X1   g13134(.A1(new_n13327_), .A2(new_n13309_), .ZN(new_n13328_));
  XOR2_X1    g13135(.A1(new_n13282_), .A2(new_n13328_), .Z(new_n13329_));
  XOR2_X1    g13136(.A1(new_n13329_), .A2(new_n13279_), .Z(new_n13330_));
  NOR2_X1    g13137(.A1(new_n13330_), .A2(new_n13252_), .ZN(new_n13331_));
  INV_X1     g13138(.I(new_n13331_), .ZN(new_n13332_));
  AOI21_X1   g13139(.A1(new_n13169_), .A2(new_n13157_), .B(new_n13246_), .ZN(new_n13333_));
  NOR2_X1    g13140(.A1(new_n13333_), .A2(new_n13247_), .ZN(new_n13334_));
  INV_X1     g13141(.I(new_n13247_), .ZN(new_n13335_));
  INV_X1     g13142(.I(new_n13157_), .ZN(new_n13336_));
  INV_X1     g13143(.I(new_n13246_), .ZN(new_n13337_));
  OAI21_X1   g13144(.A1(new_n13167_), .A2(new_n13336_), .B(new_n13337_), .ZN(new_n13338_));
  NAND2_X1   g13145(.A1(new_n13330_), .A2(new_n13252_), .ZN(new_n13339_));
  INV_X1     g13146(.I(new_n13339_), .ZN(new_n13340_));
  AOI21_X1   g13147(.A1(new_n13338_), .A2(new_n13335_), .B(new_n13340_), .ZN(new_n13341_));
  NAND2_X1   g13148(.A1(new_n13332_), .A2(new_n13339_), .ZN(new_n13342_));
  AOI22_X1   g13149(.A1(new_n13341_), .A2(new_n13332_), .B1(new_n13334_), .B2(new_n13342_), .ZN(\asquared[103] ));
  OAI21_X1   g13150(.A1(new_n13333_), .A2(new_n13247_), .B(new_n13339_), .ZN(new_n13344_));
  NAND2_X1   g13151(.A1(new_n13344_), .A2(new_n13332_), .ZN(new_n13345_));
  INV_X1     g13152(.I(new_n13328_), .ZN(new_n13346_));
  NOR2_X1    g13153(.A1(new_n13282_), .A2(new_n13346_), .ZN(new_n13347_));
  INV_X1     g13154(.I(new_n13279_), .ZN(new_n13348_));
  NOR2_X1    g13155(.A1(new_n13348_), .A2(new_n13329_), .ZN(new_n13349_));
  NOR2_X1    g13156(.A1(new_n13349_), .A2(new_n13347_), .ZN(new_n13350_));
  INV_X1     g13157(.I(new_n13350_), .ZN(new_n13351_));
  XNOR2_X1   g13158(.A1(new_n13297_), .A2(new_n13321_), .ZN(new_n13352_));
  NAND2_X1   g13159(.A1(new_n4703_), .A2(new_n7205_), .ZN(new_n13353_));
  NOR2_X1    g13160(.A1(new_n3861_), .A2(new_n6899_), .ZN(new_n13354_));
  NOR4_X1    g13161(.A1(new_n3746_), .A2(new_n4030_), .A3(new_n6316_), .A4(new_n6897_), .ZN(new_n13355_));
  OAI21_X1   g13162(.A1(new_n13354_), .A2(new_n13355_), .B(new_n13353_), .ZN(new_n13356_));
  NAND3_X1   g13163(.A1(new_n13356_), .A2(\a[42] ), .A3(\a[61] ), .ZN(new_n13357_));
  NAND2_X1   g13164(.A1(new_n13356_), .A2(new_n13353_), .ZN(new_n13358_));
  AOI22_X1   g13165(.A1(\a[44] ), .A2(\a[59] ), .B1(\a[45] ), .B2(\a[58] ), .ZN(new_n13359_));
  OAI21_X1   g13166(.A1(new_n13358_), .A2(new_n13359_), .B(new_n13357_), .ZN(new_n13360_));
  XNOR2_X1   g13167(.A1(new_n13352_), .A2(new_n13360_), .ZN(new_n13361_));
  NOR2_X1    g13168(.A1(new_n3221_), .A2(new_n7643_), .ZN(new_n13362_));
  XOR2_X1    g13169(.A1(new_n13305_), .A2(new_n13362_), .Z(new_n13363_));
  XNOR2_X1   g13170(.A1(new_n13290_), .A2(new_n13363_), .ZN(new_n13364_));
  INV_X1     g13171(.I(new_n13364_), .ZN(new_n13365_));
  NAND2_X1   g13172(.A1(new_n13361_), .A2(new_n13365_), .ZN(new_n13366_));
  NOR2_X1    g13173(.A1(new_n13361_), .A2(new_n13365_), .ZN(new_n13367_));
  INV_X1     g13174(.I(new_n13367_), .ZN(new_n13368_));
  AND2_X2    g13175(.A1(new_n13368_), .A2(new_n13366_), .Z(new_n13369_));
  AOI22_X1   g13176(.A1(\a[46] ), .A2(\a[57] ), .B1(\a[47] ), .B2(\a[56] ), .ZN(new_n13370_));
  INV_X1     g13177(.I(new_n13370_), .ZN(new_n13371_));
  NOR2_X1    g13178(.A1(new_n4721_), .A2(new_n8161_), .ZN(new_n13372_));
  NOR2_X1    g13179(.A1(new_n3666_), .A2(new_n6723_), .ZN(new_n13373_));
  AOI21_X1   g13180(.A1(new_n13371_), .A2(new_n13373_), .B(new_n13372_), .ZN(new_n13374_));
  INV_X1     g13181(.I(new_n13374_), .ZN(new_n13375_));
  OAI21_X1   g13182(.A1(new_n13372_), .A2(new_n13370_), .B(new_n13373_), .ZN(new_n13376_));
  OAI21_X1   g13183(.A1(new_n13375_), .A2(new_n13370_), .B(new_n13376_), .ZN(new_n13377_));
  OAI22_X1   g13184(.A1(new_n4903_), .A2(new_n6125_), .B1(new_n4981_), .B2(new_n6129_), .ZN(new_n13378_));
  OAI21_X1   g13185(.A1(new_n5155_), .A2(new_n6127_), .B(new_n13378_), .ZN(new_n13379_));
  NAND3_X1   g13186(.A1(new_n13379_), .A2(\a[48] ), .A3(\a[55] ), .ZN(new_n13380_));
  AOI22_X1   g13187(.A1(\a[49] ), .A2(\a[54] ), .B1(\a[50] ), .B2(\a[53] ), .ZN(new_n13381_));
  NOR2_X1    g13188(.A1(new_n5155_), .A2(new_n6127_), .ZN(new_n13382_));
  NOR2_X1    g13189(.A1(new_n13378_), .A2(new_n13382_), .ZN(new_n13383_));
  INV_X1     g13190(.I(new_n13383_), .ZN(new_n13384_));
  OAI21_X1   g13191(.A1(new_n13381_), .A2(new_n13384_), .B(new_n13380_), .ZN(new_n13385_));
  XNOR2_X1   g13192(.A1(new_n13385_), .A2(new_n13377_), .ZN(new_n13386_));
  NOR2_X1    g13193(.A1(new_n3327_), .A2(new_n7144_), .ZN(new_n13387_));
  NOR3_X1    g13194(.A1(new_n13387_), .A2(new_n5135_), .A3(new_n5175_), .ZN(new_n13388_));
  NOR2_X1    g13195(.A1(new_n13387_), .A2(\a[52] ), .ZN(new_n13389_));
  OAI21_X1   g13196(.A1(new_n13387_), .A2(\a[51] ), .B(\a[52] ), .ZN(new_n13390_));
  INV_X1     g13197(.I(new_n13390_), .ZN(new_n13391_));
  OAI22_X1   g13198(.A1(new_n13391_), .A2(new_n13389_), .B1(new_n5525_), .B2(new_n13388_), .ZN(new_n13392_));
  XOR2_X1    g13199(.A1(new_n13386_), .A2(new_n13392_), .Z(new_n13393_));
  XOR2_X1    g13200(.A1(new_n13369_), .A2(new_n13393_), .Z(new_n13394_));
  NAND2_X1   g13201(.A1(new_n13274_), .A2(new_n13271_), .ZN(new_n13395_));
  NAND2_X1   g13202(.A1(new_n13278_), .A2(new_n13395_), .ZN(new_n13396_));
  XOR2_X1    g13203(.A1(new_n13396_), .A2(new_n13394_), .Z(new_n13397_));
  NAND2_X1   g13204(.A1(new_n13292_), .A2(new_n13299_), .ZN(new_n13398_));
  NAND2_X1   g13205(.A1(new_n13300_), .A2(new_n13308_), .ZN(new_n13399_));
  AOI21_X1   g13206(.A1(new_n13314_), .A2(new_n13322_), .B(new_n13313_), .ZN(new_n13400_));
  NAND2_X1   g13207(.A1(new_n13237_), .A2(new_n13195_), .ZN(new_n13401_));
  NAND2_X1   g13208(.A1(new_n13256_), .A2(new_n13215_), .ZN(new_n13402_));
  NAND2_X1   g13209(.A1(new_n13402_), .A2(new_n13401_), .ZN(new_n13403_));
  XNOR2_X1   g13210(.A1(new_n13403_), .A2(new_n13400_), .ZN(new_n13404_));
  INV_X1     g13211(.I(new_n13404_), .ZN(new_n13405_));
  AND3_X2    g13212(.A1(new_n13405_), .A2(new_n13398_), .A3(new_n13399_), .Z(new_n13406_));
  AOI21_X1   g13213(.A1(new_n13398_), .A2(new_n13399_), .B(new_n13405_), .ZN(new_n13407_));
  NOR2_X1    g13214(.A1(new_n13406_), .A2(new_n13407_), .ZN(new_n13408_));
  NOR2_X1    g13215(.A1(new_n13323_), .A2(new_n13326_), .ZN(new_n13409_));
  NAND2_X1   g13216(.A1(new_n13323_), .A2(new_n13326_), .ZN(new_n13410_));
  OAI21_X1   g13217(.A1(new_n13309_), .A2(new_n13409_), .B(new_n13410_), .ZN(new_n13411_));
  NOR2_X1    g13218(.A1(new_n13266_), .A2(new_n13261_), .ZN(new_n13412_));
  XNOR2_X1   g13219(.A1(new_n13412_), .A2(new_n13411_), .ZN(new_n13413_));
  XOR2_X1    g13220(.A1(new_n13413_), .A2(new_n13408_), .Z(new_n13414_));
  XOR2_X1    g13221(.A1(new_n13397_), .A2(new_n13414_), .Z(new_n13415_));
  INV_X1     g13222(.I(new_n13415_), .ZN(new_n13416_));
  NOR2_X1    g13223(.A1(new_n13416_), .A2(new_n13351_), .ZN(new_n13417_));
  NOR2_X1    g13224(.A1(new_n13415_), .A2(new_n13350_), .ZN(new_n13418_));
  NOR2_X1    g13225(.A1(new_n13417_), .A2(new_n13418_), .ZN(new_n13419_));
  XOR2_X1    g13226(.A1(new_n13345_), .A2(new_n13419_), .Z(\asquared[104] ));
  AOI21_X1   g13227(.A1(new_n13344_), .A2(new_n13332_), .B(new_n13417_), .ZN(new_n13421_));
  NOR2_X1    g13228(.A1(new_n13421_), .A2(new_n13418_), .ZN(new_n13422_));
  INV_X1     g13229(.I(new_n13394_), .ZN(new_n13423_));
  NAND2_X1   g13230(.A1(new_n13396_), .A2(new_n13423_), .ZN(new_n13424_));
  INV_X1     g13231(.I(new_n13414_), .ZN(new_n13425_));
  OAI21_X1   g13232(.A1(new_n13397_), .A2(new_n13425_), .B(new_n13424_), .ZN(new_n13426_));
  NAND2_X1   g13233(.A1(new_n13298_), .A2(new_n13321_), .ZN(new_n13427_));
  NAND2_X1   g13234(.A1(new_n13352_), .A2(new_n13360_), .ZN(new_n13428_));
  NAND2_X1   g13235(.A1(new_n13428_), .A2(new_n13427_), .ZN(new_n13429_));
  NAND2_X1   g13236(.A1(new_n13305_), .A2(new_n13362_), .ZN(new_n13430_));
  NAND2_X1   g13237(.A1(new_n13291_), .A2(new_n13363_), .ZN(new_n13431_));
  NAND2_X1   g13238(.A1(new_n13431_), .A2(new_n13430_), .ZN(new_n13432_));
  NOR2_X1    g13239(.A1(new_n4667_), .A2(new_n8049_), .ZN(new_n13433_));
  AOI22_X1   g13240(.A1(\a[41] ), .A2(\a[63] ), .B1(\a[42] ), .B2(\a[62] ), .ZN(new_n13434_));
  NOR2_X1    g13241(.A1(new_n13433_), .A2(new_n13434_), .ZN(new_n13435_));
  INV_X1     g13242(.I(new_n13435_), .ZN(new_n13436_));
  NOR2_X1    g13243(.A1(new_n13436_), .A2(new_n13390_), .ZN(new_n13437_));
  NOR2_X1    g13244(.A1(new_n13435_), .A2(new_n13391_), .ZN(new_n13438_));
  NOR2_X1    g13245(.A1(new_n13437_), .A2(new_n13438_), .ZN(new_n13439_));
  XOR2_X1    g13246(.A1(new_n13432_), .A2(new_n13439_), .Z(new_n13440_));
  XOR2_X1    g13247(.A1(new_n13440_), .A2(new_n13429_), .Z(new_n13441_));
  INV_X1     g13248(.I(new_n13369_), .ZN(new_n13442_));
  OAI21_X1   g13249(.A1(new_n13442_), .A2(new_n13393_), .B(new_n13368_), .ZN(new_n13443_));
  INV_X1     g13250(.I(new_n13443_), .ZN(new_n13444_));
  AOI21_X1   g13251(.A1(new_n13401_), .A2(new_n13402_), .B(new_n13400_), .ZN(new_n13445_));
  NOR2_X1    g13252(.A1(new_n13407_), .A2(new_n13445_), .ZN(new_n13446_));
  XOR2_X1    g13253(.A1(new_n13446_), .A2(new_n13444_), .Z(new_n13447_));
  AND2_X2    g13254(.A1(new_n13447_), .A2(new_n13441_), .Z(new_n13448_));
  NOR2_X1    g13255(.A1(new_n13447_), .A2(new_n13441_), .ZN(new_n13449_));
  NOR2_X1    g13256(.A1(new_n13448_), .A2(new_n13449_), .ZN(new_n13450_));
  OAI21_X1   g13257(.A1(new_n13266_), .A2(new_n13261_), .B(new_n13411_), .ZN(new_n13451_));
  NAND2_X1   g13258(.A1(new_n13413_), .A2(new_n13408_), .ZN(new_n13452_));
  NAND2_X1   g13259(.A1(new_n13452_), .A2(new_n13451_), .ZN(new_n13453_));
  NAND2_X1   g13260(.A1(new_n4033_), .A2(new_n6898_), .ZN(new_n13454_));
  OAI22_X1   g13261(.A1(new_n4343_), .A2(new_n7454_), .B1(new_n4704_), .B2(new_n7452_), .ZN(new_n13455_));
  NAND2_X1   g13262(.A1(new_n13455_), .A2(new_n13454_), .ZN(new_n13456_));
  NAND3_X1   g13263(.A1(new_n13456_), .A2(\a[44] ), .A3(\a[60] ), .ZN(new_n13457_));
  AOI22_X1   g13264(.A1(\a[43] ), .A2(\a[61] ), .B1(\a[45] ), .B2(\a[59] ), .ZN(new_n13458_));
  NAND2_X1   g13265(.A1(new_n13456_), .A2(new_n13454_), .ZN(new_n13459_));
  OAI21_X1   g13266(.A1(new_n13458_), .A2(new_n13459_), .B(new_n13457_), .ZN(new_n13460_));
  NAND2_X1   g13267(.A1(new_n4976_), .A2(new_n6494_), .ZN(new_n13461_));
  NOR4_X1    g13268(.A1(new_n4178_), .A2(new_n4596_), .A3(new_n5856_), .A4(new_n6316_), .ZN(new_n13462_));
  NOR2_X1    g13269(.A1(new_n4721_), .A2(new_n6804_), .ZN(new_n13463_));
  OAI21_X1   g13270(.A1(new_n13463_), .A2(new_n13462_), .B(new_n13461_), .ZN(new_n13464_));
  NAND3_X1   g13271(.A1(new_n13464_), .A2(\a[46] ), .A3(\a[58] ), .ZN(new_n13465_));
  AOI22_X1   g13272(.A1(\a[47] ), .A2(\a[57] ), .B1(\a[48] ), .B2(\a[56] ), .ZN(new_n13466_));
  NAND2_X1   g13273(.A1(new_n13464_), .A2(new_n13461_), .ZN(new_n13467_));
  OAI21_X1   g13274(.A1(new_n13466_), .A2(new_n13467_), .B(new_n13465_), .ZN(new_n13468_));
  XNOR2_X1   g13275(.A1(new_n13460_), .A2(new_n13468_), .ZN(new_n13469_));
  NAND2_X1   g13276(.A1(new_n5154_), .A2(new_n6128_), .ZN(new_n13470_));
  NAND2_X1   g13277(.A1(new_n5682_), .A2(new_n7658_), .ZN(new_n13471_));
  AOI22_X1   g13278(.A1(new_n13470_), .A2(new_n13471_), .B1(new_n5439_), .B2(new_n6126_), .ZN(new_n13472_));
  AOI21_X1   g13279(.A1(\a[50] ), .A2(\a[54] ), .B(new_n5682_), .ZN(new_n13473_));
  NAND2_X1   g13280(.A1(new_n5439_), .A2(new_n6126_), .ZN(new_n13474_));
  NAND3_X1   g13281(.A1(new_n13474_), .A2(new_n13470_), .A3(new_n13471_), .ZN(new_n13475_));
  OAI22_X1   g13282(.A1(new_n13472_), .A2(new_n7659_), .B1(new_n13475_), .B2(new_n13473_), .ZN(new_n13476_));
  XOR2_X1    g13283(.A1(new_n13469_), .A2(new_n13476_), .Z(new_n13477_));
  INV_X1     g13284(.I(new_n13477_), .ZN(new_n13478_));
  XOR2_X1    g13285(.A1(new_n13383_), .A2(new_n13374_), .Z(new_n13479_));
  XOR2_X1    g13286(.A1(new_n13479_), .A2(new_n13358_), .Z(new_n13480_));
  NAND2_X1   g13287(.A1(new_n13385_), .A2(new_n13377_), .ZN(new_n13481_));
  INV_X1     g13288(.I(new_n13392_), .ZN(new_n13482_));
  OAI21_X1   g13289(.A1(new_n13386_), .A2(new_n13482_), .B(new_n13481_), .ZN(new_n13483_));
  NAND2_X1   g13290(.A1(new_n13483_), .A2(new_n13480_), .ZN(new_n13484_));
  INV_X1     g13291(.I(new_n13484_), .ZN(new_n13485_));
  NOR2_X1    g13292(.A1(new_n13483_), .A2(new_n13480_), .ZN(new_n13486_));
  NOR2_X1    g13293(.A1(new_n13485_), .A2(new_n13486_), .ZN(new_n13487_));
  NOR2_X1    g13294(.A1(new_n13487_), .A2(new_n13478_), .ZN(new_n13488_));
  NAND2_X1   g13295(.A1(new_n13487_), .A2(new_n13478_), .ZN(new_n13489_));
  INV_X1     g13296(.I(new_n13489_), .ZN(new_n13490_));
  NOR2_X1    g13297(.A1(new_n13490_), .A2(new_n13488_), .ZN(new_n13491_));
  XOR2_X1    g13298(.A1(new_n13453_), .A2(new_n13491_), .Z(new_n13492_));
  XNOR2_X1   g13299(.A1(new_n13492_), .A2(new_n13450_), .ZN(new_n13493_));
  INV_X1     g13300(.I(new_n13493_), .ZN(new_n13494_));
  NOR2_X1    g13301(.A1(new_n13426_), .A2(new_n13494_), .ZN(new_n13495_));
  INV_X1     g13302(.I(new_n13495_), .ZN(new_n13496_));
  NAND2_X1   g13303(.A1(new_n13426_), .A2(new_n13494_), .ZN(new_n13497_));
  NAND2_X1   g13304(.A1(new_n13496_), .A2(new_n13497_), .ZN(new_n13498_));
  XOR2_X1    g13305(.A1(new_n13422_), .A2(new_n13498_), .Z(\asquared[105] ));
  OAI21_X1   g13306(.A1(new_n13421_), .A2(new_n13418_), .B(new_n13496_), .ZN(new_n13500_));
  NAND2_X1   g13307(.A1(new_n13500_), .A2(new_n13497_), .ZN(new_n13501_));
  NOR2_X1    g13308(.A1(new_n13490_), .A2(new_n13485_), .ZN(new_n13502_));
  NAND2_X1   g13309(.A1(new_n13479_), .A2(new_n13358_), .ZN(new_n13503_));
  OAI21_X1   g13310(.A1(new_n13374_), .A2(new_n13383_), .B(new_n13503_), .ZN(new_n13504_));
  NOR2_X1    g13311(.A1(new_n5440_), .A2(new_n6129_), .ZN(new_n13505_));
  INV_X1     g13312(.I(new_n13505_), .ZN(new_n13506_));
  OAI22_X1   g13313(.A1(new_n5155_), .A2(new_n7185_), .B1(new_n6058_), .B2(new_n10168_), .ZN(new_n13507_));
  NAND2_X1   g13314(.A1(new_n13507_), .A2(new_n13506_), .ZN(new_n13508_));
  NAND3_X1   g13315(.A1(new_n13508_), .A2(\a[49] ), .A3(\a[56] ), .ZN(new_n13509_));
  AOI22_X1   g13316(.A1(\a[50] ), .A2(\a[55] ), .B1(\a[51] ), .B2(\a[54] ), .ZN(new_n13510_));
  NAND2_X1   g13317(.A1(new_n13508_), .A2(new_n13506_), .ZN(new_n13511_));
  OAI21_X1   g13318(.A1(new_n13510_), .A2(new_n13511_), .B(new_n13509_), .ZN(new_n13512_));
  AOI21_X1   g13319(.A1(\a[43] ), .A2(\a[62] ), .B(\a[53] ), .ZN(new_n13513_));
  NAND2_X1   g13320(.A1(new_n12647_), .A2(\a[62] ), .ZN(new_n13514_));
  INV_X1     g13321(.I(new_n13514_), .ZN(new_n13515_));
  NOR2_X1    g13322(.A1(new_n13515_), .A2(new_n5862_), .ZN(new_n13516_));
  INV_X1     g13323(.I(new_n13516_), .ZN(new_n13517_));
  NAND2_X1   g13324(.A1(new_n13515_), .A2(new_n5862_), .ZN(new_n13518_));
  OAI21_X1   g13325(.A1(new_n13517_), .A2(new_n13513_), .B(new_n13518_), .ZN(new_n13519_));
  XNOR2_X1   g13326(.A1(new_n13512_), .A2(new_n13519_), .ZN(new_n13520_));
  XNOR2_X1   g13327(.A1(new_n13520_), .A2(new_n13504_), .ZN(new_n13521_));
  NOR2_X1    g13328(.A1(new_n4977_), .A2(new_n6804_), .ZN(new_n13522_));
  AOI22_X1   g13329(.A1(new_n4720_), .A2(new_n7205_), .B1(new_n6743_), .B2(new_n7203_), .ZN(new_n13523_));
  NOR2_X1    g13330(.A1(new_n13522_), .A2(new_n13523_), .ZN(new_n13524_));
  NAND2_X1   g13331(.A1(\a[46] ), .A2(\a[59] ), .ZN(new_n13525_));
  AOI22_X1   g13332(.A1(\a[47] ), .A2(\a[58] ), .B1(\a[48] ), .B2(\a[57] ), .ZN(new_n13526_));
  NOR2_X1    g13333(.A1(new_n13524_), .A2(new_n13522_), .ZN(new_n13527_));
  INV_X1     g13334(.I(new_n13527_), .ZN(new_n13528_));
  OAI22_X1   g13335(.A1(new_n13528_), .A2(new_n13526_), .B1(new_n13524_), .B2(new_n13525_), .ZN(new_n13529_));
  OAI22_X1   g13336(.A1(new_n3861_), .A2(new_n7959_), .B1(new_n9031_), .B2(new_n13220_), .ZN(new_n13530_));
  NOR2_X1    g13337(.A1(new_n4704_), .A2(new_n7454_), .ZN(new_n13531_));
  INV_X1     g13338(.I(new_n13531_), .ZN(new_n13532_));
  NAND2_X1   g13339(.A1(new_n13532_), .A2(new_n13530_), .ZN(new_n13533_));
  NAND3_X1   g13340(.A1(new_n13533_), .A2(\a[42] ), .A3(\a[63] ), .ZN(new_n13534_));
  AOI22_X1   g13341(.A1(\a[44] ), .A2(\a[61] ), .B1(\a[45] ), .B2(\a[60] ), .ZN(new_n13535_));
  NAND2_X1   g13342(.A1(new_n13533_), .A2(new_n13532_), .ZN(new_n13536_));
  OAI21_X1   g13343(.A1(new_n13535_), .A2(new_n13536_), .B(new_n13534_), .ZN(new_n13537_));
  NOR2_X1    g13344(.A1(new_n13437_), .A2(new_n13433_), .ZN(new_n13538_));
  XOR2_X1    g13345(.A1(new_n13537_), .A2(new_n13538_), .Z(new_n13539_));
  XNOR2_X1   g13346(.A1(new_n13539_), .A2(new_n13529_), .ZN(new_n13540_));
  XNOR2_X1   g13347(.A1(new_n13521_), .A2(new_n13540_), .ZN(new_n13541_));
  XOR2_X1    g13348(.A1(new_n13502_), .A2(new_n13541_), .Z(new_n13542_));
  NAND2_X1   g13349(.A1(new_n13432_), .A2(new_n13439_), .ZN(new_n13543_));
  NAND2_X1   g13350(.A1(new_n13440_), .A2(new_n13429_), .ZN(new_n13544_));
  NAND2_X1   g13351(.A1(new_n13544_), .A2(new_n13543_), .ZN(new_n13545_));
  XOR2_X1    g13352(.A1(new_n13467_), .A2(new_n13475_), .Z(new_n13546_));
  XOR2_X1    g13353(.A1(new_n13546_), .A2(new_n13459_), .Z(new_n13547_));
  NAND2_X1   g13354(.A1(new_n13460_), .A2(new_n13468_), .ZN(new_n13548_));
  INV_X1     g13355(.I(new_n13469_), .ZN(new_n13549_));
  NAND2_X1   g13356(.A1(new_n13549_), .A2(new_n13476_), .ZN(new_n13550_));
  NAND2_X1   g13357(.A1(new_n13550_), .A2(new_n13548_), .ZN(new_n13551_));
  XOR2_X1    g13358(.A1(new_n13551_), .A2(new_n13547_), .Z(new_n13552_));
  XNOR2_X1   g13359(.A1(new_n13552_), .A2(new_n13545_), .ZN(new_n13553_));
  NOR2_X1    g13360(.A1(new_n13446_), .A2(new_n13444_), .ZN(new_n13554_));
  NOR2_X1    g13361(.A1(new_n13448_), .A2(new_n13554_), .ZN(new_n13555_));
  XOR2_X1    g13362(.A1(new_n13555_), .A2(new_n13553_), .Z(new_n13556_));
  XOR2_X1    g13363(.A1(new_n13556_), .A2(new_n13542_), .Z(new_n13557_));
  INV_X1     g13364(.I(new_n13557_), .ZN(new_n13558_));
  NAND2_X1   g13365(.A1(new_n13453_), .A2(new_n13491_), .ZN(new_n13559_));
  NAND2_X1   g13366(.A1(new_n13492_), .A2(new_n13450_), .ZN(new_n13560_));
  NAND2_X1   g13367(.A1(new_n13560_), .A2(new_n13559_), .ZN(new_n13561_));
  INV_X1     g13368(.I(new_n13561_), .ZN(new_n13562_));
  NOR2_X1    g13369(.A1(new_n13558_), .A2(new_n13562_), .ZN(new_n13563_));
  NOR2_X1    g13370(.A1(new_n13557_), .A2(new_n13561_), .ZN(new_n13564_));
  NOR2_X1    g13371(.A1(new_n13563_), .A2(new_n13564_), .ZN(new_n13565_));
  XOR2_X1    g13372(.A1(new_n13501_), .A2(new_n13565_), .Z(\asquared[106] ));
  AOI21_X1   g13373(.A1(new_n13500_), .A2(new_n13497_), .B(new_n13564_), .ZN(new_n13567_));
  NOR2_X1    g13374(.A1(new_n13567_), .A2(new_n13563_), .ZN(new_n13568_));
  NAND2_X1   g13375(.A1(new_n13551_), .A2(new_n13547_), .ZN(new_n13569_));
  NAND2_X1   g13376(.A1(new_n13552_), .A2(new_n13545_), .ZN(new_n13570_));
  NAND2_X1   g13377(.A1(new_n13570_), .A2(new_n13569_), .ZN(new_n13571_));
  NAND2_X1   g13378(.A1(new_n13467_), .A2(new_n13475_), .ZN(new_n13572_));
  NAND2_X1   g13379(.A1(new_n13546_), .A2(new_n13459_), .ZN(new_n13573_));
  NAND2_X1   g13380(.A1(new_n13573_), .A2(new_n13572_), .ZN(new_n13574_));
  NOR2_X1    g13381(.A1(new_n4981_), .A2(new_n6804_), .ZN(new_n13575_));
  NOR2_X1    g13382(.A1(new_n4979_), .A2(new_n7204_), .ZN(new_n13576_));
  NOR2_X1    g13383(.A1(new_n4977_), .A2(new_n7206_), .ZN(new_n13577_));
  NOR2_X1    g13384(.A1(new_n13576_), .A2(new_n13577_), .ZN(new_n13578_));
  NOR2_X1    g13385(.A1(new_n13578_), .A2(new_n13575_), .ZN(new_n13579_));
  NAND2_X1   g13386(.A1(\a[47] ), .A2(\a[59] ), .ZN(new_n13580_));
  AOI21_X1   g13387(.A1(\a[48] ), .A2(\a[58] ), .B(new_n9656_), .ZN(new_n13581_));
  NOR2_X1    g13388(.A1(new_n13579_), .A2(new_n13575_), .ZN(new_n13582_));
  INV_X1     g13389(.I(new_n13582_), .ZN(new_n13583_));
  OAI22_X1   g13390(.A1(new_n13583_), .A2(new_n13581_), .B1(new_n13579_), .B2(new_n13580_), .ZN(new_n13584_));
  NAND2_X1   g13391(.A1(new_n5524_), .A2(new_n6128_), .ZN(new_n13585_));
  OAI22_X1   g13392(.A1(new_n5440_), .A2(new_n7185_), .B1(new_n5523_), .B2(new_n6058_), .ZN(new_n13586_));
  NAND2_X1   g13393(.A1(new_n13586_), .A2(new_n13585_), .ZN(new_n13587_));
  NAND2_X1   g13394(.A1(new_n13587_), .A2(new_n13585_), .ZN(new_n13588_));
  AOI21_X1   g13395(.A1(\a[51] ), .A2(\a[55] ), .B(new_n8420_), .ZN(new_n13589_));
  NAND3_X1   g13396(.A1(new_n13587_), .A2(\a[50] ), .A3(\a[56] ), .ZN(new_n13590_));
  OAI21_X1   g13397(.A1(new_n13588_), .A2(new_n13589_), .B(new_n13590_), .ZN(new_n13591_));
  XOR2_X1    g13398(.A1(new_n13584_), .A2(new_n13591_), .Z(new_n13592_));
  XOR2_X1    g13399(.A1(new_n13592_), .A2(new_n13574_), .Z(new_n13593_));
  INV_X1     g13400(.I(new_n13593_), .ZN(new_n13594_));
  XNOR2_X1   g13401(.A1(new_n13536_), .A2(new_n13527_), .ZN(new_n13595_));
  NOR3_X1    g13402(.A1(new_n11581_), .A2(new_n4178_), .A3(new_n6723_), .ZN(new_n13596_));
  NOR2_X1    g13403(.A1(new_n4704_), .A2(new_n7591_), .ZN(new_n13597_));
  OAI22_X1   g13404(.A1(new_n13596_), .A2(new_n13597_), .B1(new_n4430_), .B2(new_n7454_), .ZN(new_n13598_));
  INV_X1     g13405(.I(new_n13598_), .ZN(new_n13599_));
  AOI22_X1   g13406(.A1(\a[45] ), .A2(\a[61] ), .B1(\a[46] ), .B2(\a[60] ), .ZN(new_n13600_));
  NOR2_X1    g13407(.A1(new_n4430_), .A2(new_n7454_), .ZN(new_n13601_));
  NOR2_X1    g13408(.A1(new_n13599_), .A2(new_n13601_), .ZN(new_n13602_));
  INV_X1     g13409(.I(new_n13602_), .ZN(new_n13603_));
  OAI22_X1   g13410(.A1(new_n13603_), .A2(new_n13600_), .B1(new_n11581_), .B2(new_n13599_), .ZN(new_n13604_));
  XNOR2_X1   g13411(.A1(new_n13604_), .A2(new_n13595_), .ZN(new_n13605_));
  NOR2_X1    g13412(.A1(new_n13594_), .A2(new_n13605_), .ZN(new_n13606_));
  INV_X1     g13413(.I(new_n13606_), .ZN(new_n13607_));
  NAND2_X1   g13414(.A1(new_n13594_), .A2(new_n13605_), .ZN(new_n13608_));
  NAND3_X1   g13415(.A1(new_n13571_), .A2(new_n13607_), .A3(new_n13608_), .ZN(new_n13609_));
  NAND2_X1   g13416(.A1(new_n13609_), .A2(new_n13571_), .ZN(new_n13610_));
  NAND2_X1   g13417(.A1(new_n13609_), .A2(new_n13607_), .ZN(new_n13611_));
  INV_X1     g13418(.I(new_n13611_), .ZN(new_n13612_));
  NAND2_X1   g13419(.A1(new_n13612_), .A2(new_n13608_), .ZN(new_n13613_));
  NAND2_X1   g13420(.A1(new_n13613_), .A2(new_n13610_), .ZN(new_n13614_));
  NAND2_X1   g13421(.A1(new_n13512_), .A2(new_n13519_), .ZN(new_n13615_));
  INV_X1     g13422(.I(new_n13520_), .ZN(new_n13616_));
  NAND2_X1   g13423(.A1(new_n13616_), .A2(new_n13504_), .ZN(new_n13617_));
  NAND2_X1   g13424(.A1(new_n13617_), .A2(new_n13615_), .ZN(new_n13618_));
  INV_X1     g13425(.I(new_n13537_), .ZN(new_n13619_));
  INV_X1     g13426(.I(new_n13539_), .ZN(new_n13620_));
  NAND2_X1   g13427(.A1(new_n13620_), .A2(new_n13529_), .ZN(new_n13621_));
  OAI21_X1   g13428(.A1(new_n13619_), .A2(new_n13538_), .B(new_n13621_), .ZN(new_n13622_));
  NAND2_X1   g13429(.A1(\a[43] ), .A2(\a[63] ), .ZN(new_n13623_));
  XOR2_X1    g13430(.A1(new_n13516_), .A2(new_n13623_), .Z(new_n13624_));
  XOR2_X1    g13431(.A1(new_n13624_), .A2(new_n13511_), .Z(new_n13625_));
  NOR2_X1    g13432(.A1(new_n13622_), .A2(new_n13625_), .ZN(new_n13626_));
  NAND2_X1   g13433(.A1(new_n13622_), .A2(new_n13625_), .ZN(new_n13627_));
  INV_X1     g13434(.I(new_n13627_), .ZN(new_n13628_));
  NOR2_X1    g13435(.A1(new_n13628_), .A2(new_n13626_), .ZN(new_n13629_));
  NOR2_X1    g13436(.A1(new_n13629_), .A2(new_n13618_), .ZN(new_n13630_));
  NAND2_X1   g13437(.A1(new_n13629_), .A2(new_n13618_), .ZN(new_n13631_));
  INV_X1     g13438(.I(new_n13631_), .ZN(new_n13632_));
  NOR2_X1    g13439(.A1(new_n13632_), .A2(new_n13630_), .ZN(new_n13633_));
  INV_X1     g13440(.I(new_n13633_), .ZN(new_n13634_));
  NAND2_X1   g13441(.A1(new_n13521_), .A2(new_n13540_), .ZN(new_n13635_));
  OAI21_X1   g13442(.A1(new_n13502_), .A2(new_n13541_), .B(new_n13635_), .ZN(new_n13636_));
  INV_X1     g13443(.I(new_n13636_), .ZN(new_n13637_));
  NOR2_X1    g13444(.A1(new_n13634_), .A2(new_n13637_), .ZN(new_n13638_));
  NOR2_X1    g13445(.A1(new_n13633_), .A2(new_n13636_), .ZN(new_n13639_));
  NOR2_X1    g13446(.A1(new_n13638_), .A2(new_n13639_), .ZN(new_n13640_));
  XOR2_X1    g13447(.A1(new_n13614_), .A2(new_n13640_), .Z(new_n13641_));
  NAND2_X1   g13448(.A1(new_n13556_), .A2(new_n13542_), .ZN(new_n13642_));
  OAI21_X1   g13449(.A1(new_n13553_), .A2(new_n13555_), .B(new_n13642_), .ZN(new_n13643_));
  NAND2_X1   g13450(.A1(new_n13643_), .A2(new_n13641_), .ZN(new_n13644_));
  NOR2_X1    g13451(.A1(new_n13643_), .A2(new_n13641_), .ZN(new_n13645_));
  INV_X1     g13452(.I(new_n13645_), .ZN(new_n13646_));
  NAND2_X1   g13453(.A1(new_n13646_), .A2(new_n13644_), .ZN(new_n13647_));
  INV_X1     g13454(.I(new_n13563_), .ZN(new_n13648_));
  INV_X1     g13455(.I(new_n13497_), .ZN(new_n13649_));
  INV_X1     g13456(.I(new_n13418_), .ZN(new_n13650_));
  INV_X1     g13457(.I(new_n13417_), .ZN(new_n13651_));
  OAI21_X1   g13458(.A1(new_n13341_), .A2(new_n13331_), .B(new_n13651_), .ZN(new_n13652_));
  AOI21_X1   g13459(.A1(new_n13652_), .A2(new_n13650_), .B(new_n13495_), .ZN(new_n13653_));
  INV_X1     g13460(.I(new_n13564_), .ZN(new_n13654_));
  OAI21_X1   g13461(.A1(new_n13653_), .A2(new_n13649_), .B(new_n13654_), .ZN(new_n13655_));
  AOI21_X1   g13462(.A1(new_n13655_), .A2(new_n13648_), .B(new_n13645_), .ZN(new_n13656_));
  AOI22_X1   g13463(.A1(new_n13656_), .A2(new_n13644_), .B1(new_n13568_), .B2(new_n13647_), .ZN(\asquared[107] ));
  OAI21_X1   g13464(.A1(new_n13567_), .A2(new_n13563_), .B(new_n13646_), .ZN(new_n13658_));
  NAND2_X1   g13465(.A1(new_n13658_), .A2(new_n13644_), .ZN(new_n13659_));
  AOI21_X1   g13466(.A1(new_n13614_), .A2(new_n13640_), .B(new_n13638_), .ZN(new_n13660_));
  NOR2_X1    g13467(.A1(new_n13632_), .A2(new_n13628_), .ZN(new_n13661_));
  XOR2_X1    g13468(.A1(new_n13602_), .A2(new_n13582_), .Z(new_n13662_));
  NAND2_X1   g13469(.A1(\a[59] ), .A2(\a[63] ), .ZN(new_n13663_));
  NOR3_X1    g13470(.A1(new_n13663_), .A2(new_n3859_), .A3(new_n4596_), .ZN(new_n13664_));
  NOR2_X1    g13471(.A1(new_n4981_), .A2(new_n7206_), .ZN(new_n13665_));
  NOR2_X1    g13472(.A1(new_n6316_), .A2(new_n7643_), .ZN(new_n13666_));
  NAND2_X1   g13473(.A1(new_n6573_), .A2(new_n13666_), .ZN(new_n13667_));
  OAI21_X1   g13474(.A1(new_n13665_), .A2(new_n13664_), .B(new_n13667_), .ZN(new_n13668_));
  NAND3_X1   g13475(.A1(new_n13668_), .A2(\a[48] ), .A3(\a[59] ), .ZN(new_n13669_));
  AOI22_X1   g13476(.A1(\a[44] ), .A2(\a[63] ), .B1(\a[49] ), .B2(\a[58] ), .ZN(new_n13670_));
  NAND2_X1   g13477(.A1(new_n13668_), .A2(new_n13667_), .ZN(new_n13671_));
  OAI21_X1   g13478(.A1(new_n13670_), .A2(new_n13671_), .B(new_n13669_), .ZN(new_n13672_));
  XOR2_X1    g13479(.A1(new_n13662_), .A2(new_n13672_), .Z(new_n13673_));
  NAND2_X1   g13480(.A1(\a[47] ), .A2(\a[60] ), .ZN(new_n13674_));
  NAND2_X1   g13481(.A1(\a[46] ), .A2(\a[61] ), .ZN(new_n13675_));
  AOI22_X1   g13482(.A1(new_n4720_), .A2(new_n7453_), .B1(new_n13674_), .B2(new_n13675_), .ZN(new_n13676_));
  XNOR2_X1   g13483(.A1(new_n13588_), .A2(new_n13676_), .ZN(new_n13677_));
  OAI22_X1   g13484(.A1(new_n5440_), .A2(new_n8161_), .B1(new_n5523_), .B2(new_n8952_), .ZN(new_n13678_));
  OAI21_X1   g13485(.A1(new_n5525_), .A2(new_n7185_), .B(new_n13678_), .ZN(new_n13679_));
  NAND3_X1   g13486(.A1(new_n13679_), .A2(\a[50] ), .A3(\a[57] ), .ZN(new_n13680_));
  AOI22_X1   g13487(.A1(\a[51] ), .A2(\a[56] ), .B1(\a[52] ), .B2(\a[55] ), .ZN(new_n13681_));
  NOR2_X1    g13488(.A1(new_n5525_), .A2(new_n7185_), .ZN(new_n13682_));
  NOR2_X1    g13489(.A1(new_n13678_), .A2(new_n13682_), .ZN(new_n13683_));
  INV_X1     g13490(.I(new_n13683_), .ZN(new_n13684_));
  OAI21_X1   g13491(.A1(new_n13681_), .A2(new_n13684_), .B(new_n13680_), .ZN(new_n13685_));
  NOR2_X1    g13492(.A1(new_n4030_), .A2(new_n7144_), .ZN(new_n13686_));
  NAND3_X1   g13493(.A1(new_n13686_), .A2(\a[53] ), .A3(\a[54] ), .ZN(new_n13687_));
  NOR2_X1    g13494(.A1(new_n13686_), .A2(\a[54] ), .ZN(new_n13688_));
  OAI21_X1   g13495(.A1(new_n13686_), .A2(\a[53] ), .B(\a[54] ), .ZN(new_n13689_));
  INV_X1     g13496(.I(new_n13689_), .ZN(new_n13690_));
  OAI21_X1   g13497(.A1(new_n13688_), .A2(new_n13690_), .B(new_n13687_), .ZN(new_n13691_));
  XNOR2_X1   g13498(.A1(new_n13685_), .A2(new_n13691_), .ZN(new_n13692_));
  XNOR2_X1   g13499(.A1(new_n13692_), .A2(new_n13677_), .ZN(new_n13693_));
  XOR2_X1    g13500(.A1(new_n13693_), .A2(new_n13673_), .Z(new_n13694_));
  XOR2_X1    g13501(.A1(new_n13661_), .A2(new_n13694_), .Z(new_n13695_));
  NAND2_X1   g13502(.A1(new_n13584_), .A2(new_n13591_), .ZN(new_n13696_));
  NAND2_X1   g13503(.A1(new_n13592_), .A2(new_n13574_), .ZN(new_n13697_));
  NAND2_X1   g13504(.A1(new_n13697_), .A2(new_n13696_), .ZN(new_n13698_));
  NAND2_X1   g13505(.A1(new_n13528_), .A2(new_n13536_), .ZN(new_n13699_));
  NAND2_X1   g13506(.A1(new_n13604_), .A2(new_n13595_), .ZN(new_n13700_));
  NAND2_X1   g13507(.A1(new_n13700_), .A2(new_n13699_), .ZN(new_n13701_));
  NAND2_X1   g13508(.A1(new_n13624_), .A2(new_n13511_), .ZN(new_n13702_));
  OAI21_X1   g13509(.A1(new_n13516_), .A2(new_n13623_), .B(new_n13702_), .ZN(new_n13703_));
  XOR2_X1    g13510(.A1(new_n13701_), .A2(new_n13703_), .Z(new_n13704_));
  XOR2_X1    g13511(.A1(new_n13704_), .A2(new_n13698_), .Z(new_n13705_));
  NOR2_X1    g13512(.A1(new_n13611_), .A2(new_n13705_), .ZN(new_n13706_));
  INV_X1     g13513(.I(new_n13705_), .ZN(new_n13707_));
  NOR2_X1    g13514(.A1(new_n13612_), .A2(new_n13707_), .ZN(new_n13708_));
  NOR2_X1    g13515(.A1(new_n13708_), .A2(new_n13706_), .ZN(new_n13709_));
  NAND2_X1   g13516(.A1(new_n13709_), .A2(new_n13695_), .ZN(new_n13710_));
  INV_X1     g13517(.I(new_n13710_), .ZN(new_n13711_));
  NOR2_X1    g13518(.A1(new_n13709_), .A2(new_n13695_), .ZN(new_n13712_));
  NOR2_X1    g13519(.A1(new_n13711_), .A2(new_n13712_), .ZN(new_n13713_));
  INV_X1     g13520(.I(new_n13713_), .ZN(new_n13714_));
  NOR2_X1    g13521(.A1(new_n13714_), .A2(new_n13660_), .ZN(new_n13715_));
  NAND2_X1   g13522(.A1(new_n13714_), .A2(new_n13660_), .ZN(new_n13716_));
  INV_X1     g13523(.I(new_n13716_), .ZN(new_n13717_));
  NOR2_X1    g13524(.A1(new_n13717_), .A2(new_n13715_), .ZN(new_n13718_));
  XOR2_X1    g13525(.A1(new_n13659_), .A2(new_n13718_), .Z(\asquared[108] ));
  NOR2_X1    g13526(.A1(new_n13711_), .A2(new_n13708_), .ZN(new_n13720_));
  INV_X1     g13527(.I(new_n13693_), .ZN(new_n13721_));
  NAND2_X1   g13528(.A1(new_n13721_), .A2(new_n13673_), .ZN(new_n13722_));
  OAI21_X1   g13529(.A1(new_n13661_), .A2(new_n13694_), .B(new_n13722_), .ZN(new_n13723_));
  NAND2_X1   g13530(.A1(new_n13662_), .A2(new_n13672_), .ZN(new_n13724_));
  OAI21_X1   g13531(.A1(new_n13582_), .A2(new_n13602_), .B(new_n13724_), .ZN(new_n13725_));
  INV_X1     g13532(.I(new_n10971_), .ZN(new_n13726_));
  NAND2_X1   g13533(.A1(new_n5524_), .A2(new_n6494_), .ZN(new_n13727_));
  NAND2_X1   g13534(.A1(new_n5682_), .A2(new_n8951_), .ZN(new_n13728_));
  AOI22_X1   g13535(.A1(new_n13727_), .A2(new_n13728_), .B1(new_n5862_), .B2(new_n7184_), .ZN(new_n13729_));
  NAND2_X1   g13536(.A1(new_n5862_), .A2(new_n7184_), .ZN(new_n13730_));
  NAND3_X1   g13537(.A1(new_n13730_), .A2(new_n13727_), .A3(new_n13728_), .ZN(new_n13731_));
  AOI21_X1   g13538(.A1(\a[52] ), .A2(\a[56] ), .B(new_n6124_), .ZN(new_n13732_));
  OAI22_X1   g13539(.A1(new_n13729_), .A2(new_n13726_), .B1(new_n13731_), .B2(new_n13732_), .ZN(new_n13733_));
  XOR2_X1    g13540(.A1(new_n13725_), .A2(new_n13733_), .Z(new_n13734_));
  NAND2_X1   g13541(.A1(new_n13685_), .A2(new_n13691_), .ZN(new_n13735_));
  OAI21_X1   g13542(.A1(new_n13692_), .A2(new_n13677_), .B(new_n13735_), .ZN(new_n13736_));
  XNOR2_X1   g13543(.A1(new_n13734_), .A2(new_n13736_), .ZN(new_n13737_));
  INV_X1     g13544(.I(new_n13737_), .ZN(new_n13738_));
  NOR2_X1    g13545(.A1(new_n13723_), .A2(new_n13738_), .ZN(new_n13739_));
  NAND2_X1   g13546(.A1(new_n13723_), .A2(new_n13738_), .ZN(new_n13740_));
  INV_X1     g13547(.I(new_n13740_), .ZN(new_n13741_));
  NOR2_X1    g13548(.A1(new_n13741_), .A2(new_n13739_), .ZN(new_n13742_));
  NAND2_X1   g13549(.A1(new_n4980_), .A2(new_n7451_), .ZN(new_n13743_));
  NAND2_X1   g13550(.A1(new_n4902_), .A2(new_n7800_), .ZN(new_n13744_));
  AOI22_X1   g13551(.A1(new_n13743_), .A2(new_n13744_), .B1(new_n5154_), .B2(new_n7205_), .ZN(new_n13745_));
  NAND2_X1   g13552(.A1(\a[48] ), .A2(\a[60] ), .ZN(new_n13746_));
  AOI22_X1   g13553(.A1(\a[49] ), .A2(\a[59] ), .B1(\a[50] ), .B2(\a[58] ), .ZN(new_n13747_));
  NAND2_X1   g13554(.A1(new_n5154_), .A2(new_n7205_), .ZN(new_n13748_));
  NAND3_X1   g13555(.A1(new_n13748_), .A2(new_n13743_), .A3(new_n13744_), .ZN(new_n13749_));
  OAI22_X1   g13556(.A1(new_n13745_), .A2(new_n13746_), .B1(new_n13749_), .B2(new_n13747_), .ZN(new_n13750_));
  NAND2_X1   g13557(.A1(new_n13588_), .A2(new_n13676_), .ZN(new_n13751_));
  OAI21_X1   g13558(.A1(new_n4721_), .A2(new_n7454_), .B(new_n13751_), .ZN(new_n13752_));
  NOR2_X1    g13559(.A1(new_n4721_), .A2(new_n7591_), .ZN(new_n13753_));
  AOI22_X1   g13560(.A1(new_n4313_), .A2(new_n7852_), .B1(new_n4429_), .B2(new_n7644_), .ZN(new_n13754_));
  NOR2_X1    g13561(.A1(new_n13753_), .A2(new_n13754_), .ZN(new_n13755_));
  NOR3_X1    g13562(.A1(new_n13755_), .A2(new_n4030_), .A3(new_n7643_), .ZN(new_n13756_));
  AOI22_X1   g13563(.A1(\a[46] ), .A2(\a[62] ), .B1(\a[47] ), .B2(\a[61] ), .ZN(new_n13757_));
  NOR2_X1    g13564(.A1(new_n13755_), .A2(new_n13753_), .ZN(new_n13758_));
  INV_X1     g13565(.I(new_n13758_), .ZN(new_n13759_));
  NOR2_X1    g13566(.A1(new_n13759_), .A2(new_n13757_), .ZN(new_n13760_));
  NOR2_X1    g13567(.A1(new_n13760_), .A2(new_n13756_), .ZN(new_n13761_));
  XNOR2_X1   g13568(.A1(new_n13752_), .A2(new_n13761_), .ZN(new_n13762_));
  XOR2_X1    g13569(.A1(new_n13762_), .A2(new_n13750_), .Z(new_n13763_));
  NAND2_X1   g13570(.A1(new_n13701_), .A2(new_n13703_), .ZN(new_n13764_));
  NAND2_X1   g13571(.A1(new_n13704_), .A2(new_n13698_), .ZN(new_n13765_));
  NAND2_X1   g13572(.A1(new_n13765_), .A2(new_n13764_), .ZN(new_n13766_));
  XOR2_X1    g13573(.A1(new_n13683_), .A2(new_n13689_), .Z(new_n13767_));
  XOR2_X1    g13574(.A1(new_n13767_), .A2(new_n13671_), .Z(new_n13768_));
  XOR2_X1    g13575(.A1(new_n13766_), .A2(new_n13768_), .Z(new_n13769_));
  NAND2_X1   g13576(.A1(new_n13769_), .A2(new_n13763_), .ZN(new_n13770_));
  OR2_X2     g13577(.A1(new_n13769_), .A2(new_n13763_), .Z(new_n13771_));
  AND2_X2    g13578(.A1(new_n13771_), .A2(new_n13770_), .Z(new_n13772_));
  XNOR2_X1   g13579(.A1(new_n13742_), .A2(new_n13772_), .ZN(new_n13773_));
  NOR2_X1    g13580(.A1(new_n13773_), .A2(new_n13720_), .ZN(new_n13774_));
  INV_X1     g13581(.I(new_n13774_), .ZN(new_n13775_));
  AOI21_X1   g13582(.A1(new_n13658_), .A2(new_n13644_), .B(new_n13717_), .ZN(new_n13776_));
  NOR2_X1    g13583(.A1(new_n13776_), .A2(new_n13715_), .ZN(new_n13777_));
  INV_X1     g13584(.I(new_n13715_), .ZN(new_n13778_));
  INV_X1     g13585(.I(new_n13644_), .ZN(new_n13779_));
  OAI21_X1   g13586(.A1(new_n13656_), .A2(new_n13779_), .B(new_n13716_), .ZN(new_n13780_));
  NAND2_X1   g13587(.A1(new_n13773_), .A2(new_n13720_), .ZN(new_n13781_));
  INV_X1     g13588(.I(new_n13781_), .ZN(new_n13782_));
  AOI21_X1   g13589(.A1(new_n13780_), .A2(new_n13778_), .B(new_n13782_), .ZN(new_n13783_));
  NAND2_X1   g13590(.A1(new_n13775_), .A2(new_n13781_), .ZN(new_n13784_));
  AOI22_X1   g13591(.A1(new_n13783_), .A2(new_n13775_), .B1(new_n13777_), .B2(new_n13784_), .ZN(\asquared[109] ));
  OAI21_X1   g13592(.A1(new_n13776_), .A2(new_n13715_), .B(new_n13781_), .ZN(new_n13786_));
  NAND2_X1   g13593(.A1(new_n13786_), .A2(new_n13775_), .ZN(new_n13787_));
  NAND2_X1   g13594(.A1(new_n13766_), .A2(new_n13768_), .ZN(new_n13788_));
  NAND2_X1   g13595(.A1(new_n13762_), .A2(new_n13750_), .ZN(new_n13789_));
  OAI21_X1   g13596(.A1(new_n13756_), .A2(new_n13760_), .B(new_n13752_), .ZN(new_n13790_));
  NAND2_X1   g13597(.A1(new_n13789_), .A2(new_n13790_), .ZN(new_n13791_));
  NAND2_X1   g13598(.A1(new_n13767_), .A2(new_n13671_), .ZN(new_n13792_));
  OAI21_X1   g13599(.A1(new_n13683_), .A2(new_n13689_), .B(new_n13792_), .ZN(new_n13793_));
  NOR2_X1    g13600(.A1(new_n4312_), .A2(new_n7144_), .ZN(new_n13794_));
  NAND3_X1   g13601(.A1(new_n13794_), .A2(\a[54] ), .A3(\a[55] ), .ZN(new_n13795_));
  OAI21_X1   g13602(.A1(new_n13794_), .A2(\a[54] ), .B(\a[55] ), .ZN(new_n13796_));
  OAI21_X1   g13603(.A1(\a[55] ), .A2(new_n13794_), .B(new_n13796_), .ZN(new_n13797_));
  NAND2_X1   g13604(.A1(new_n13795_), .A2(new_n13797_), .ZN(new_n13798_));
  XNOR2_X1   g13605(.A1(new_n13793_), .A2(new_n13798_), .ZN(new_n13799_));
  XNOR2_X1   g13606(.A1(new_n13791_), .A2(new_n13799_), .ZN(new_n13800_));
  INV_X1     g13607(.I(new_n13800_), .ZN(new_n13801_));
  AND3_X2    g13608(.A1(new_n13770_), .A2(new_n13788_), .A3(new_n13801_), .Z(new_n13802_));
  AOI21_X1   g13609(.A1(new_n13770_), .A2(new_n13788_), .B(new_n13801_), .ZN(new_n13803_));
  NOR2_X1    g13610(.A1(new_n13802_), .A2(new_n13803_), .ZN(new_n13804_));
  NOR2_X1    g13611(.A1(new_n6563_), .A2(new_n8161_), .ZN(new_n13805_));
  AOI22_X1   g13612(.A1(new_n5524_), .A2(new_n6803_), .B1(new_n5682_), .B2(new_n6317_), .ZN(new_n13806_));
  NOR2_X1    g13613(.A1(new_n13805_), .A2(new_n13806_), .ZN(new_n13807_));
  NAND2_X1   g13614(.A1(\a[51] ), .A2(\a[58] ), .ZN(new_n13808_));
  AOI22_X1   g13615(.A1(\a[52] ), .A2(\a[57] ), .B1(\a[53] ), .B2(\a[56] ), .ZN(new_n13809_));
  NOR2_X1    g13616(.A1(new_n13807_), .A2(new_n13805_), .ZN(new_n13810_));
  INV_X1     g13617(.I(new_n13810_), .ZN(new_n13811_));
  OAI22_X1   g13618(.A1(new_n13811_), .A2(new_n13809_), .B1(new_n13807_), .B2(new_n13808_), .ZN(new_n13812_));
  NOR2_X1    g13619(.A1(new_n5155_), .A2(new_n7452_), .ZN(new_n13813_));
  INV_X1     g13620(.I(new_n13813_), .ZN(new_n13814_));
  OAI22_X1   g13621(.A1(new_n4903_), .A2(new_n6899_), .B1(new_n4981_), .B2(new_n7454_), .ZN(new_n13815_));
  NAND2_X1   g13622(.A1(new_n13815_), .A2(new_n13814_), .ZN(new_n13816_));
  NAND3_X1   g13623(.A1(new_n13816_), .A2(\a[48] ), .A3(\a[61] ), .ZN(new_n13817_));
  AOI22_X1   g13624(.A1(\a[49] ), .A2(\a[60] ), .B1(\a[50] ), .B2(\a[59] ), .ZN(new_n13818_));
  NAND2_X1   g13625(.A1(new_n13816_), .A2(new_n13814_), .ZN(new_n13819_));
  OAI21_X1   g13626(.A1(new_n13818_), .A2(new_n13819_), .B(new_n13817_), .ZN(new_n13820_));
  XOR2_X1    g13627(.A1(new_n13820_), .A2(new_n13758_), .Z(new_n13821_));
  INV_X1     g13628(.I(new_n13821_), .ZN(new_n13822_));
  NAND2_X1   g13629(.A1(new_n13822_), .A2(new_n13812_), .ZN(new_n13823_));
  INV_X1     g13630(.I(new_n13823_), .ZN(new_n13824_));
  NOR2_X1    g13631(.A1(new_n13822_), .A2(new_n13812_), .ZN(new_n13825_));
  NOR2_X1    g13632(.A1(new_n13824_), .A2(new_n13825_), .ZN(new_n13826_));
  NAND2_X1   g13633(.A1(new_n13725_), .A2(new_n13733_), .ZN(new_n13827_));
  NAND2_X1   g13634(.A1(new_n13734_), .A2(new_n13736_), .ZN(new_n13828_));
  NAND2_X1   g13635(.A1(new_n13828_), .A2(new_n13827_), .ZN(new_n13829_));
  NOR2_X1    g13636(.A1(new_n4178_), .A2(new_n7643_), .ZN(new_n13830_));
  XOR2_X1    g13637(.A1(new_n13731_), .A2(new_n13830_), .Z(new_n13831_));
  XOR2_X1    g13638(.A1(new_n13831_), .A2(new_n13749_), .Z(new_n13832_));
  XOR2_X1    g13639(.A1(new_n13829_), .A2(new_n13832_), .Z(new_n13833_));
  XOR2_X1    g13640(.A1(new_n13833_), .A2(new_n13826_), .Z(new_n13834_));
  XNOR2_X1   g13641(.A1(new_n13804_), .A2(new_n13834_), .ZN(new_n13835_));
  INV_X1     g13642(.I(new_n13835_), .ZN(new_n13836_));
  AOI21_X1   g13643(.A1(new_n13742_), .A2(new_n13772_), .B(new_n13741_), .ZN(new_n13837_));
  INV_X1     g13644(.I(new_n13837_), .ZN(new_n13838_));
  NOR2_X1    g13645(.A1(new_n13836_), .A2(new_n13838_), .ZN(new_n13839_));
  NOR2_X1    g13646(.A1(new_n13835_), .A2(new_n13837_), .ZN(new_n13840_));
  NOR2_X1    g13647(.A1(new_n13839_), .A2(new_n13840_), .ZN(new_n13841_));
  XOR2_X1    g13648(.A1(new_n13787_), .A2(new_n13841_), .Z(\asquared[110] ));
  AOI21_X1   g13649(.A1(new_n13786_), .A2(new_n13775_), .B(new_n13839_), .ZN(new_n13843_));
  NOR2_X1    g13650(.A1(new_n13843_), .A2(new_n13840_), .ZN(new_n13844_));
  AOI21_X1   g13651(.A1(new_n13804_), .A2(new_n13834_), .B(new_n13803_), .ZN(new_n13845_));
  NAND2_X1   g13652(.A1(new_n13793_), .A2(new_n13798_), .ZN(new_n13846_));
  INV_X1     g13653(.I(new_n13799_), .ZN(new_n13847_));
  NAND2_X1   g13654(.A1(new_n13847_), .A2(new_n13791_), .ZN(new_n13848_));
  NAND2_X1   g13655(.A1(new_n13848_), .A2(new_n13846_), .ZN(new_n13849_));
  XOR2_X1    g13656(.A1(new_n13819_), .A2(new_n13811_), .Z(new_n13850_));
  NAND2_X1   g13657(.A1(new_n5439_), .A2(new_n7451_), .ZN(new_n13851_));
  OAI22_X1   g13658(.A1(new_n5155_), .A2(new_n7454_), .B1(new_n6899_), .B2(new_n10168_), .ZN(new_n13852_));
  NAND2_X1   g13659(.A1(new_n13852_), .A2(new_n13851_), .ZN(new_n13853_));
  NAND3_X1   g13660(.A1(new_n13853_), .A2(\a[49] ), .A3(\a[61] ), .ZN(new_n13854_));
  AOI22_X1   g13661(.A1(\a[50] ), .A2(\a[60] ), .B1(\a[51] ), .B2(\a[59] ), .ZN(new_n13855_));
  NAND2_X1   g13662(.A1(new_n13853_), .A2(new_n13851_), .ZN(new_n13856_));
  OAI21_X1   g13663(.A1(new_n13855_), .A2(new_n13856_), .B(new_n13854_), .ZN(new_n13857_));
  XNOR2_X1   g13664(.A1(new_n13850_), .A2(new_n13857_), .ZN(new_n13858_));
  INV_X1     g13665(.I(new_n13858_), .ZN(new_n13859_));
  NAND2_X1   g13666(.A1(new_n13820_), .A2(new_n13759_), .ZN(new_n13860_));
  NAND2_X1   g13667(.A1(new_n13823_), .A2(new_n13860_), .ZN(new_n13861_));
  NOR2_X1    g13668(.A1(new_n13861_), .A2(new_n13859_), .ZN(new_n13862_));
  NAND2_X1   g13669(.A1(new_n13861_), .A2(new_n13859_), .ZN(new_n13863_));
  INV_X1     g13670(.I(new_n13863_), .ZN(new_n13864_));
  NOR2_X1    g13671(.A1(new_n13864_), .A2(new_n13862_), .ZN(new_n13865_));
  NOR2_X1    g13672(.A1(new_n13865_), .A2(new_n13849_), .ZN(new_n13866_));
  NAND2_X1   g13673(.A1(new_n13865_), .A2(new_n13849_), .ZN(new_n13867_));
  INV_X1     g13674(.I(new_n13867_), .ZN(new_n13868_));
  NOR2_X1    g13675(.A1(new_n13868_), .A2(new_n13866_), .ZN(new_n13869_));
  NAND2_X1   g13676(.A1(new_n13829_), .A2(new_n13832_), .ZN(new_n13870_));
  NAND2_X1   g13677(.A1(new_n13833_), .A2(new_n13826_), .ZN(new_n13871_));
  NAND2_X1   g13678(.A1(new_n13871_), .A2(new_n13870_), .ZN(new_n13872_));
  NAND2_X1   g13679(.A1(new_n13731_), .A2(new_n13830_), .ZN(new_n13873_));
  NAND2_X1   g13680(.A1(new_n13831_), .A2(new_n13749_), .ZN(new_n13874_));
  NAND2_X1   g13681(.A1(new_n13874_), .A2(new_n13873_), .ZN(new_n13875_));
  AOI22_X1   g13682(.A1(\a[47] ), .A2(\a[63] ), .B1(\a[48] ), .B2(\a[62] ), .ZN(new_n13876_));
  AOI21_X1   g13683(.A1(new_n4976_), .A2(new_n7644_), .B(new_n13876_), .ZN(new_n13877_));
  XOR2_X1    g13684(.A1(new_n13877_), .A2(new_n13796_), .Z(new_n13878_));
  NAND2_X1   g13685(.A1(new_n6126_), .A2(new_n6494_), .ZN(new_n13879_));
  NOR4_X1    g13686(.A1(new_n5175_), .A2(new_n5617_), .A3(new_n5856_), .A4(new_n6316_), .ZN(new_n13880_));
  NOR2_X1    g13687(.A1(new_n6563_), .A2(new_n6804_), .ZN(new_n13881_));
  OAI21_X1   g13688(.A1(new_n13881_), .A2(new_n13880_), .B(new_n13879_), .ZN(new_n13882_));
  NAND2_X1   g13689(.A1(new_n13882_), .A2(new_n13879_), .ZN(new_n13883_));
  AOI21_X1   g13690(.A1(\a[53] ), .A2(\a[57] ), .B(new_n5857_), .ZN(new_n13884_));
  NOR2_X1    g13691(.A1(new_n13883_), .A2(new_n13884_), .ZN(new_n13885_));
  NOR2_X1    g13692(.A1(new_n5175_), .A2(new_n6316_), .ZN(new_n13886_));
  AOI21_X1   g13693(.A1(new_n13882_), .A2(new_n13886_), .B(new_n13885_), .ZN(new_n13887_));
  XOR2_X1    g13694(.A1(new_n13887_), .A2(new_n13878_), .Z(new_n13888_));
  NOR2_X1    g13695(.A1(new_n13888_), .A2(new_n13875_), .ZN(new_n13889_));
  NAND2_X1   g13696(.A1(new_n13888_), .A2(new_n13875_), .ZN(new_n13890_));
  INV_X1     g13697(.I(new_n13890_), .ZN(new_n13891_));
  NOR2_X1    g13698(.A1(new_n13891_), .A2(new_n13889_), .ZN(new_n13892_));
  INV_X1     g13699(.I(new_n13892_), .ZN(new_n13893_));
  NAND2_X1   g13700(.A1(new_n13872_), .A2(new_n13893_), .ZN(new_n13894_));
  NOR2_X1    g13701(.A1(new_n13872_), .A2(new_n13893_), .ZN(new_n13895_));
  INV_X1     g13702(.I(new_n13895_), .ZN(new_n13896_));
  NAND2_X1   g13703(.A1(new_n13896_), .A2(new_n13894_), .ZN(new_n13897_));
  NAND2_X1   g13704(.A1(new_n13897_), .A2(new_n13869_), .ZN(new_n13898_));
  INV_X1     g13705(.I(new_n13869_), .ZN(new_n13899_));
  NAND3_X1   g13706(.A1(new_n13896_), .A2(new_n13899_), .A3(new_n13894_), .ZN(new_n13900_));
  NAND2_X1   g13707(.A1(new_n13898_), .A2(new_n13900_), .ZN(new_n13901_));
  NOR2_X1    g13708(.A1(new_n13901_), .A2(new_n13845_), .ZN(new_n13902_));
  INV_X1     g13709(.I(new_n13902_), .ZN(new_n13903_));
  NAND2_X1   g13710(.A1(new_n13901_), .A2(new_n13845_), .ZN(new_n13904_));
  NAND2_X1   g13711(.A1(new_n13903_), .A2(new_n13904_), .ZN(new_n13905_));
  INV_X1     g13712(.I(new_n13840_), .ZN(new_n13906_));
  INV_X1     g13713(.I(new_n13839_), .ZN(new_n13907_));
  OAI21_X1   g13714(.A1(new_n13783_), .A2(new_n13774_), .B(new_n13907_), .ZN(new_n13908_));
  INV_X1     g13715(.I(new_n13904_), .ZN(new_n13909_));
  AOI21_X1   g13716(.A1(new_n13908_), .A2(new_n13906_), .B(new_n13909_), .ZN(new_n13910_));
  AOI22_X1   g13717(.A1(new_n13910_), .A2(new_n13903_), .B1(new_n13844_), .B2(new_n13905_), .ZN(\asquared[111] ));
  OAI21_X1   g13718(.A1(new_n13843_), .A2(new_n13840_), .B(new_n13904_), .ZN(new_n13912_));
  NAND2_X1   g13719(.A1(new_n13912_), .A2(new_n13903_), .ZN(new_n13913_));
  NAND2_X1   g13720(.A1(new_n13872_), .A2(new_n13892_), .ZN(new_n13914_));
  NAND2_X1   g13721(.A1(new_n13898_), .A2(new_n13914_), .ZN(new_n13915_));
  OAI21_X1   g13722(.A1(new_n13878_), .A2(new_n13887_), .B(new_n13890_), .ZN(new_n13916_));
  OAI22_X1   g13723(.A1(new_n13796_), .A2(new_n13876_), .B1(new_n4977_), .B2(new_n8049_), .ZN(new_n13917_));
  XOR2_X1    g13724(.A1(new_n13856_), .A2(new_n13883_), .Z(new_n13918_));
  XOR2_X1    g13725(.A1(new_n13918_), .A2(new_n13917_), .Z(new_n13919_));
  NAND2_X1   g13726(.A1(new_n13819_), .A2(new_n13811_), .ZN(new_n13920_));
  NAND2_X1   g13727(.A1(new_n13850_), .A2(new_n13857_), .ZN(new_n13921_));
  NAND2_X1   g13728(.A1(new_n13921_), .A2(new_n13920_), .ZN(new_n13922_));
  NAND2_X1   g13729(.A1(new_n13919_), .A2(new_n13922_), .ZN(new_n13923_));
  INV_X1     g13730(.I(new_n13923_), .ZN(new_n13924_));
  NOR2_X1    g13731(.A1(new_n13919_), .A2(new_n13922_), .ZN(new_n13925_));
  NOR2_X1    g13732(.A1(new_n13924_), .A2(new_n13925_), .ZN(new_n13926_));
  NOR2_X1    g13733(.A1(new_n13926_), .A2(new_n13916_), .ZN(new_n13927_));
  NAND2_X1   g13734(.A1(new_n13926_), .A2(new_n13916_), .ZN(new_n13928_));
  INV_X1     g13735(.I(new_n13928_), .ZN(new_n13929_));
  NOR2_X1    g13736(.A1(new_n13929_), .A2(new_n13927_), .ZN(new_n13930_));
  NOR2_X1    g13737(.A1(new_n13868_), .A2(new_n13864_), .ZN(new_n13931_));
  NOR2_X1    g13738(.A1(new_n5856_), .A2(new_n7144_), .ZN(new_n13932_));
  INV_X1     g13739(.I(new_n13932_), .ZN(new_n13933_));
  NOR2_X1    g13740(.A1(new_n13933_), .A2(new_n4702_), .ZN(new_n13934_));
  NAND2_X1   g13741(.A1(new_n13934_), .A2(new_n7184_), .ZN(new_n13935_));
  AOI21_X1   g13742(.A1(\a[49] ), .A2(\a[62] ), .B(\a[56] ), .ZN(new_n13936_));
  NOR2_X1    g13743(.A1(new_n13934_), .A2(new_n7184_), .ZN(new_n13937_));
  INV_X1     g13744(.I(new_n13937_), .ZN(new_n13938_));
  OAI21_X1   g13745(.A1(new_n13938_), .A2(new_n13936_), .B(new_n13935_), .ZN(new_n13939_));
  NOR2_X1    g13746(.A1(new_n5440_), .A2(new_n7454_), .ZN(new_n13940_));
  INV_X1     g13747(.I(new_n13940_), .ZN(new_n13941_));
  OAI22_X1   g13748(.A1(new_n4903_), .A2(new_n7959_), .B1(new_n9031_), .B2(new_n13042_), .ZN(new_n13942_));
  NAND2_X1   g13749(.A1(new_n13941_), .A2(new_n13942_), .ZN(new_n13943_));
  NAND3_X1   g13750(.A1(new_n13943_), .A2(\a[48] ), .A3(\a[63] ), .ZN(new_n13944_));
  AOI22_X1   g13751(.A1(\a[50] ), .A2(\a[61] ), .B1(\a[51] ), .B2(\a[60] ), .ZN(new_n13945_));
  NAND2_X1   g13752(.A1(new_n13943_), .A2(new_n13941_), .ZN(new_n13946_));
  OAI21_X1   g13753(.A1(new_n13945_), .A2(new_n13946_), .B(new_n13944_), .ZN(new_n13947_));
  XNOR2_X1   g13754(.A1(new_n13947_), .A2(new_n13939_), .ZN(new_n13948_));
  NOR2_X1    g13755(.A1(new_n6127_), .A2(new_n6804_), .ZN(new_n13949_));
  AOI22_X1   g13756(.A1(new_n5862_), .A2(new_n7205_), .B1(new_n7203_), .B2(new_n8420_), .ZN(new_n13950_));
  NOR2_X1    g13757(.A1(new_n13949_), .A2(new_n13950_), .ZN(new_n13951_));
  NAND2_X1   g13758(.A1(\a[52] ), .A2(\a[59] ), .ZN(new_n13952_));
  AOI21_X1   g13759(.A1(\a[53] ), .A2(\a[58] ), .B(new_n10611_), .ZN(new_n13953_));
  NOR2_X1    g13760(.A1(new_n13951_), .A2(new_n13949_), .ZN(new_n13954_));
  INV_X1     g13761(.I(new_n13954_), .ZN(new_n13955_));
  OAI22_X1   g13762(.A1(new_n13955_), .A2(new_n13953_), .B1(new_n13951_), .B2(new_n13952_), .ZN(new_n13956_));
  XOR2_X1    g13763(.A1(new_n13948_), .A2(new_n13956_), .Z(new_n13957_));
  XOR2_X1    g13764(.A1(new_n13931_), .A2(new_n13957_), .Z(new_n13958_));
  NAND2_X1   g13765(.A1(new_n13958_), .A2(new_n13930_), .ZN(new_n13959_));
  INV_X1     g13766(.I(new_n13959_), .ZN(new_n13960_));
  NOR2_X1    g13767(.A1(new_n13958_), .A2(new_n13930_), .ZN(new_n13961_));
  NOR2_X1    g13768(.A1(new_n13960_), .A2(new_n13961_), .ZN(new_n13962_));
  NOR2_X1    g13769(.A1(new_n13915_), .A2(new_n13962_), .ZN(new_n13963_));
  NAND2_X1   g13770(.A1(new_n13915_), .A2(new_n13962_), .ZN(new_n13964_));
  INV_X1     g13771(.I(new_n13964_), .ZN(new_n13965_));
  NOR2_X1    g13772(.A1(new_n13965_), .A2(new_n13963_), .ZN(new_n13966_));
  XOR2_X1    g13773(.A1(new_n13913_), .A2(new_n13966_), .Z(\asquared[112] ));
  NOR2_X1    g13774(.A1(new_n13931_), .A2(new_n13957_), .ZN(new_n13968_));
  NOR2_X1    g13775(.A1(new_n13960_), .A2(new_n13968_), .ZN(new_n13969_));
  NOR2_X1    g13776(.A1(new_n13938_), .A2(new_n12995_), .ZN(new_n13970_));
  NOR2_X1    g13777(.A1(new_n13937_), .A2(new_n12996_), .ZN(new_n13971_));
  NOR2_X1    g13778(.A1(new_n13970_), .A2(new_n13971_), .ZN(new_n13972_));
  NOR2_X1    g13779(.A1(new_n13972_), .A2(new_n13955_), .ZN(new_n13973_));
  INV_X1     g13780(.I(new_n13972_), .ZN(new_n13974_));
  NOR2_X1    g13781(.A1(new_n13974_), .A2(new_n13954_), .ZN(new_n13975_));
  NOR2_X1    g13782(.A1(new_n13975_), .A2(new_n13973_), .ZN(new_n13976_));
  NAND2_X1   g13783(.A1(new_n13856_), .A2(new_n13883_), .ZN(new_n13977_));
  NAND2_X1   g13784(.A1(new_n13918_), .A2(new_n13917_), .ZN(new_n13978_));
  NAND2_X1   g13785(.A1(new_n13978_), .A2(new_n13977_), .ZN(new_n13979_));
  NAND2_X1   g13786(.A1(new_n13947_), .A2(new_n13939_), .ZN(new_n13980_));
  INV_X1     g13787(.I(new_n13948_), .ZN(new_n13981_));
  NAND2_X1   g13788(.A1(new_n13981_), .A2(new_n13956_), .ZN(new_n13982_));
  NAND2_X1   g13789(.A1(new_n13982_), .A2(new_n13980_), .ZN(new_n13983_));
  XOR2_X1    g13790(.A1(new_n13983_), .A2(new_n13979_), .Z(new_n13984_));
  XNOR2_X1   g13791(.A1(new_n13984_), .A2(new_n13976_), .ZN(new_n13985_));
  NOR2_X1    g13792(.A1(new_n13929_), .A2(new_n13924_), .ZN(new_n13986_));
  NOR2_X1    g13793(.A1(new_n6129_), .A2(new_n6804_), .ZN(new_n13987_));
  NOR2_X1    g13794(.A1(new_n5680_), .A2(new_n6548_), .ZN(new_n13988_));
  NAND3_X1   g13795(.A1(new_n13988_), .A2(\a[53] ), .A3(\a[57] ), .ZN(new_n13989_));
  NAND2_X1   g13796(.A1(new_n6126_), .A2(new_n7205_), .ZN(new_n13990_));
  AOI21_X1   g13797(.A1(new_n13989_), .A2(new_n13990_), .B(new_n13987_), .ZN(new_n13991_));
  NOR2_X1    g13798(.A1(new_n13991_), .A2(new_n13987_), .ZN(new_n13992_));
  INV_X1     g13799(.I(new_n13992_), .ZN(new_n13993_));
  AOI21_X1   g13800(.A1(\a[54] ), .A2(\a[58] ), .B(new_n8951_), .ZN(new_n13994_));
  NAND2_X1   g13801(.A1(\a[53] ), .A2(\a[59] ), .ZN(new_n13995_));
  OAI22_X1   g13802(.A1(new_n13993_), .A2(new_n13994_), .B1(new_n13991_), .B2(new_n13995_), .ZN(new_n13996_));
  AOI22_X1   g13803(.A1(\a[51] ), .A2(new_n7852_), .B1(new_n9030_), .B2(\a[52] ), .ZN(new_n13997_));
  NOR2_X1    g13804(.A1(new_n5525_), .A2(new_n7454_), .ZN(new_n13998_));
  NOR3_X1    g13805(.A1(new_n13998_), .A2(new_n4702_), .A3(new_n13997_), .ZN(new_n13999_));
  NOR3_X1    g13806(.A1(new_n13999_), .A2(new_n4702_), .A3(new_n7643_), .ZN(new_n14000_));
  NOR2_X1    g13807(.A1(new_n13999_), .A2(new_n13998_), .ZN(new_n14001_));
  AOI22_X1   g13808(.A1(\a[51] ), .A2(\a[61] ), .B1(\a[52] ), .B2(\a[60] ), .ZN(new_n14002_));
  INV_X1     g13809(.I(new_n14002_), .ZN(new_n14003_));
  AOI21_X1   g13810(.A1(new_n14001_), .A2(new_n14003_), .B(new_n14000_), .ZN(new_n14004_));
  XOR2_X1    g13811(.A1(new_n14004_), .A2(new_n13946_), .Z(new_n14005_));
  INV_X1     g13812(.I(new_n14005_), .ZN(new_n14006_));
  NOR2_X1    g13813(.A1(new_n14006_), .A2(new_n13996_), .ZN(new_n14007_));
  NAND2_X1   g13814(.A1(new_n14006_), .A2(new_n13996_), .ZN(new_n14008_));
  INV_X1     g13815(.I(new_n14008_), .ZN(new_n14009_));
  NOR2_X1    g13816(.A1(new_n14009_), .A2(new_n14007_), .ZN(new_n14010_));
  INV_X1     g13817(.I(new_n14010_), .ZN(new_n14011_));
  XOR2_X1    g13818(.A1(new_n13986_), .A2(new_n14011_), .Z(new_n14012_));
  XNOR2_X1   g13819(.A1(new_n14012_), .A2(new_n13985_), .ZN(new_n14013_));
  INV_X1     g13820(.I(new_n14013_), .ZN(new_n14014_));
  NOR2_X1    g13821(.A1(new_n13969_), .A2(new_n14014_), .ZN(new_n14015_));
  INV_X1     g13822(.I(new_n14015_), .ZN(new_n14016_));
  AOI21_X1   g13823(.A1(new_n13912_), .A2(new_n13903_), .B(new_n13963_), .ZN(new_n14017_));
  NOR2_X1    g13824(.A1(new_n14017_), .A2(new_n13965_), .ZN(new_n14018_));
  INV_X1     g13825(.I(new_n13963_), .ZN(new_n14019_));
  OAI21_X1   g13826(.A1(new_n13910_), .A2(new_n13902_), .B(new_n14019_), .ZN(new_n14020_));
  NAND2_X1   g13827(.A1(new_n13969_), .A2(new_n14014_), .ZN(new_n14021_));
  INV_X1     g13828(.I(new_n14021_), .ZN(new_n14022_));
  AOI21_X1   g13829(.A1(new_n14020_), .A2(new_n13964_), .B(new_n14022_), .ZN(new_n14023_));
  NAND2_X1   g13830(.A1(new_n14016_), .A2(new_n14021_), .ZN(new_n14024_));
  AOI22_X1   g13831(.A1(new_n14023_), .A2(new_n14016_), .B1(new_n14018_), .B2(new_n14024_), .ZN(\asquared[113] ));
  OAI21_X1   g13832(.A1(new_n14017_), .A2(new_n13965_), .B(new_n14021_), .ZN(new_n14026_));
  NAND2_X1   g13833(.A1(new_n14026_), .A2(new_n14016_), .ZN(new_n14027_));
  NOR2_X1    g13834(.A1(new_n13986_), .A2(new_n14011_), .ZN(new_n14028_));
  INV_X1     g13835(.I(new_n14012_), .ZN(new_n14029_));
  NOR2_X1    g13836(.A1(new_n14029_), .A2(new_n13985_), .ZN(new_n14030_));
  NOR2_X1    g13837(.A1(new_n14030_), .A2(new_n14028_), .ZN(new_n14031_));
  INV_X1     g13838(.I(new_n14004_), .ZN(new_n14032_));
  AOI21_X1   g13839(.A1(new_n13946_), .A2(new_n14032_), .B(new_n14009_), .ZN(new_n14033_));
  NOR2_X1    g13840(.A1(new_n6563_), .A2(new_n7454_), .ZN(new_n14034_));
  INV_X1     g13841(.I(new_n14034_), .ZN(new_n14035_));
  NOR2_X1    g13842(.A1(new_n5425_), .A2(new_n6723_), .ZN(new_n14036_));
  NOR2_X1    g13843(.A1(new_n5175_), .A2(new_n6897_), .ZN(new_n14037_));
  OAI21_X1   g13844(.A1(new_n14036_), .A2(new_n14037_), .B(new_n14035_), .ZN(new_n14038_));
  XNOR2_X1   g13845(.A1(new_n13992_), .A2(new_n14038_), .ZN(new_n14039_));
  NOR2_X1    g13846(.A1(new_n13975_), .A2(new_n13971_), .ZN(new_n14040_));
  XOR2_X1    g13847(.A1(new_n14040_), .A2(new_n14039_), .Z(new_n14041_));
  XNOR2_X1   g13848(.A1(new_n14041_), .A2(new_n14033_), .ZN(new_n14042_));
  NAND2_X1   g13849(.A1(new_n13983_), .A2(new_n13979_), .ZN(new_n14043_));
  NAND2_X1   g13850(.A1(new_n13984_), .A2(new_n13976_), .ZN(new_n14044_));
  NAND2_X1   g13851(.A1(new_n14044_), .A2(new_n14043_), .ZN(new_n14045_));
  AOI21_X1   g13852(.A1(\a[51] ), .A2(\a[62] ), .B(\a[57] ), .ZN(new_n14046_));
  NOR2_X1    g13853(.A1(new_n13726_), .A2(new_n7144_), .ZN(new_n14047_));
  NOR2_X1    g13854(.A1(new_n14047_), .A2(new_n6494_), .ZN(new_n14048_));
  INV_X1     g13855(.I(new_n14048_), .ZN(new_n14049_));
  NAND2_X1   g13856(.A1(new_n14047_), .A2(new_n6494_), .ZN(new_n14050_));
  OAI21_X1   g13857(.A1(new_n14049_), .A2(new_n14046_), .B(new_n14050_), .ZN(new_n14051_));
  OAI21_X1   g13858(.A1(new_n5617_), .A2(new_n6548_), .B(new_n12590_), .ZN(new_n14052_));
  NOR2_X1    g13859(.A1(new_n4901_), .A2(new_n7643_), .ZN(new_n14053_));
  NOR2_X1    g13860(.A1(new_n6129_), .A2(new_n7206_), .ZN(new_n14054_));
  INV_X1     g13861(.I(new_n14054_), .ZN(new_n14055_));
  NAND3_X1   g13862(.A1(new_n14055_), .A2(new_n14052_), .A3(new_n14053_), .ZN(new_n14056_));
  AOI21_X1   g13863(.A1(new_n14052_), .A2(new_n14053_), .B(new_n14054_), .ZN(new_n14057_));
  AOI22_X1   g13864(.A1(new_n14056_), .A2(new_n14053_), .B1(new_n14052_), .B2(new_n14057_), .ZN(new_n14058_));
  XNOR2_X1   g13865(.A1(new_n14058_), .A2(new_n14001_), .ZN(new_n14059_));
  XNOR2_X1   g13866(.A1(new_n14059_), .A2(new_n14051_), .ZN(new_n14060_));
  NOR2_X1    g13867(.A1(new_n14045_), .A2(new_n14060_), .ZN(new_n14061_));
  NAND2_X1   g13868(.A1(new_n14045_), .A2(new_n14060_), .ZN(new_n14062_));
  INV_X1     g13869(.I(new_n14062_), .ZN(new_n14063_));
  NOR2_X1    g13870(.A1(new_n14063_), .A2(new_n14061_), .ZN(new_n14064_));
  NAND2_X1   g13871(.A1(new_n14064_), .A2(new_n14042_), .ZN(new_n14065_));
  INV_X1     g13872(.I(new_n14065_), .ZN(new_n14066_));
  NOR2_X1    g13873(.A1(new_n14064_), .A2(new_n14042_), .ZN(new_n14067_));
  NOR2_X1    g13874(.A1(new_n14066_), .A2(new_n14067_), .ZN(new_n14068_));
  INV_X1     g13875(.I(new_n14068_), .ZN(new_n14069_));
  NOR2_X1    g13876(.A1(new_n14069_), .A2(new_n14031_), .ZN(new_n14070_));
  NAND2_X1   g13877(.A1(new_n14069_), .A2(new_n14031_), .ZN(new_n14071_));
  INV_X1     g13878(.I(new_n14071_), .ZN(new_n14072_));
  NOR2_X1    g13879(.A1(new_n14072_), .A2(new_n14070_), .ZN(new_n14073_));
  XOR2_X1    g13880(.A1(new_n14027_), .A2(new_n14073_), .Z(\asquared[114] ));
  AOI21_X1   g13881(.A1(new_n14026_), .A2(new_n14016_), .B(new_n14072_), .ZN(new_n14075_));
  NOR2_X1    g13882(.A1(new_n14075_), .A2(new_n14070_), .ZN(new_n14076_));
  NOR2_X1    g13883(.A1(new_n14066_), .A2(new_n14063_), .ZN(new_n14077_));
  INV_X1     g13884(.I(new_n14077_), .ZN(new_n14078_));
  INV_X1     g13885(.I(new_n14059_), .ZN(new_n14079_));
  NAND2_X1   g13886(.A1(new_n14079_), .A2(new_n14051_), .ZN(new_n14080_));
  OAI21_X1   g13887(.A1(new_n14001_), .A2(new_n14058_), .B(new_n14080_), .ZN(new_n14081_));
  NOR2_X1    g13888(.A1(new_n6563_), .A2(new_n7591_), .ZN(new_n14082_));
  NOR2_X1    g13889(.A1(new_n5525_), .A2(new_n8049_), .ZN(new_n14083_));
  NOR2_X1    g13890(.A1(new_n5683_), .A2(new_n7959_), .ZN(new_n14084_));
  NOR2_X1    g13891(.A1(new_n14083_), .A2(new_n14084_), .ZN(new_n14085_));
  NOR2_X1    g13892(.A1(new_n14085_), .A2(new_n14082_), .ZN(new_n14086_));
  NOR3_X1    g13893(.A1(new_n14086_), .A2(new_n5135_), .A3(new_n7643_), .ZN(new_n14087_));
  AOI22_X1   g13894(.A1(\a[52] ), .A2(\a[62] ), .B1(\a[53] ), .B2(\a[61] ), .ZN(new_n14088_));
  NOR3_X1    g13895(.A1(new_n14086_), .A2(new_n14082_), .A3(new_n14088_), .ZN(new_n14089_));
  NOR2_X1    g13896(.A1(new_n14089_), .A2(new_n14087_), .ZN(new_n14090_));
  OAI22_X1   g13897(.A1(new_n6058_), .A2(new_n7801_), .B1(new_n6129_), .B2(new_n7452_), .ZN(new_n14091_));
  AOI21_X1   g13898(.A1(new_n7184_), .A2(new_n7205_), .B(new_n14091_), .ZN(new_n14092_));
  OAI21_X1   g13899(.A1(new_n6317_), .A2(new_n13988_), .B(new_n14092_), .ZN(new_n14093_));
  OAI21_X1   g13900(.A1(new_n7185_), .A2(new_n7206_), .B(new_n14091_), .ZN(new_n14094_));
  NAND3_X1   g13901(.A1(new_n14094_), .A2(\a[54] ), .A3(\a[60] ), .ZN(new_n14095_));
  NAND2_X1   g13902(.A1(new_n14093_), .A2(new_n14095_), .ZN(new_n14096_));
  XOR2_X1    g13903(.A1(new_n14090_), .A2(new_n14096_), .Z(new_n14097_));
  XNOR2_X1   g13904(.A1(new_n14081_), .A2(new_n14097_), .ZN(new_n14098_));
  NOR2_X1    g13905(.A1(new_n14040_), .A2(new_n14039_), .ZN(new_n14099_));
  INV_X1     g13906(.I(new_n14041_), .ZN(new_n14100_));
  NOR2_X1    g13907(.A1(new_n14033_), .A2(new_n14100_), .ZN(new_n14101_));
  NOR2_X1    g13908(.A1(new_n14101_), .A2(new_n14099_), .ZN(new_n14102_));
  OAI21_X1   g13909(.A1(new_n13992_), .A2(new_n14038_), .B(new_n14035_), .ZN(new_n14103_));
  XOR2_X1    g13910(.A1(new_n14057_), .A2(new_n14048_), .Z(new_n14104_));
  NOR2_X1    g13911(.A1(new_n14104_), .A2(new_n14103_), .ZN(new_n14105_));
  NAND2_X1   g13912(.A1(new_n14104_), .A2(new_n14103_), .ZN(new_n14106_));
  INV_X1     g13913(.I(new_n14106_), .ZN(new_n14107_));
  NOR2_X1    g13914(.A1(new_n14107_), .A2(new_n14105_), .ZN(new_n14108_));
  INV_X1     g13915(.I(new_n14108_), .ZN(new_n14109_));
  XOR2_X1    g13916(.A1(new_n14102_), .A2(new_n14109_), .Z(new_n14110_));
  NAND2_X1   g13917(.A1(new_n14110_), .A2(new_n14098_), .ZN(new_n14111_));
  INV_X1     g13918(.I(new_n14111_), .ZN(new_n14112_));
  NOR2_X1    g13919(.A1(new_n14110_), .A2(new_n14098_), .ZN(new_n14113_));
  NOR2_X1    g13920(.A1(new_n14112_), .A2(new_n14113_), .ZN(new_n14114_));
  NAND2_X1   g13921(.A1(new_n14078_), .A2(new_n14114_), .ZN(new_n14115_));
  NOR2_X1    g13922(.A1(new_n14078_), .A2(new_n14114_), .ZN(new_n14116_));
  INV_X1     g13923(.I(new_n14116_), .ZN(new_n14117_));
  NAND2_X1   g13924(.A1(new_n14117_), .A2(new_n14115_), .ZN(new_n14118_));
  INV_X1     g13925(.I(new_n14070_), .ZN(new_n14119_));
  OAI21_X1   g13926(.A1(new_n14023_), .A2(new_n14015_), .B(new_n14071_), .ZN(new_n14120_));
  AOI21_X1   g13927(.A1(new_n14120_), .A2(new_n14119_), .B(new_n14116_), .ZN(new_n14121_));
  AOI22_X1   g13928(.A1(new_n14121_), .A2(new_n14115_), .B1(new_n14076_), .B2(new_n14118_), .ZN(\asquared[115] ));
  OAI21_X1   g13929(.A1(new_n14075_), .A2(new_n14070_), .B(new_n14117_), .ZN(new_n14123_));
  NAND2_X1   g13930(.A1(new_n14123_), .A2(new_n14115_), .ZN(new_n14124_));
  NOR2_X1    g13931(.A1(new_n14102_), .A2(new_n14109_), .ZN(new_n14125_));
  NOR2_X1    g13932(.A1(new_n14112_), .A2(new_n14125_), .ZN(new_n14126_));
  INV_X1     g13933(.I(new_n14126_), .ZN(new_n14127_));
  NOR2_X1    g13934(.A1(new_n14057_), .A2(new_n14048_), .ZN(new_n14128_));
  NOR2_X1    g13935(.A1(new_n14107_), .A2(new_n14128_), .ZN(new_n14129_));
  NOR2_X1    g13936(.A1(new_n7185_), .A2(new_n7452_), .ZN(new_n14130_));
  INV_X1     g13937(.I(new_n14130_), .ZN(new_n14131_));
  OAI22_X1   g13938(.A1(new_n6058_), .A2(new_n6899_), .B1(new_n6129_), .B2(new_n7454_), .ZN(new_n14132_));
  NAND2_X1   g13939(.A1(new_n14132_), .A2(new_n14131_), .ZN(new_n14133_));
  NAND3_X1   g13940(.A1(new_n14133_), .A2(\a[54] ), .A3(\a[61] ), .ZN(new_n14134_));
  AOI21_X1   g13941(.A1(\a[55] ), .A2(\a[60] ), .B(new_n10714_), .ZN(new_n14135_));
  NAND2_X1   g13942(.A1(new_n14133_), .A2(new_n14131_), .ZN(new_n14136_));
  OAI21_X1   g13943(.A1(new_n14135_), .A2(new_n14136_), .B(new_n14134_), .ZN(new_n14137_));
  NAND2_X1   g13944(.A1(\a[53] ), .A2(\a[62] ), .ZN(new_n14138_));
  NAND2_X1   g13945(.A1(new_n14138_), .A2(new_n6316_), .ZN(new_n14139_));
  NOR2_X1    g13946(.A1(new_n14138_), .A2(new_n6316_), .ZN(new_n14140_));
  NOR2_X1    g13947(.A1(new_n6804_), .A2(new_n14140_), .ZN(new_n14141_));
  INV_X1     g13948(.I(new_n14141_), .ZN(new_n14142_));
  NOR2_X1    g13949(.A1(new_n14140_), .A2(new_n6803_), .ZN(new_n14143_));
  AOI22_X1   g13950(.A1(new_n14142_), .A2(new_n6803_), .B1(new_n14139_), .B2(new_n14143_), .ZN(new_n14144_));
  XOR2_X1    g13951(.A1(new_n14137_), .A2(new_n14144_), .Z(new_n14145_));
  XOR2_X1    g13952(.A1(new_n14145_), .A2(new_n14129_), .Z(new_n14146_));
  INV_X1     g13953(.I(new_n14081_), .ZN(new_n14147_));
  OAI21_X1   g13954(.A1(new_n14087_), .A2(new_n14089_), .B(new_n14096_), .ZN(new_n14148_));
  OAI21_X1   g13955(.A1(new_n14147_), .A2(new_n14097_), .B(new_n14148_), .ZN(new_n14149_));
  NOR2_X1    g13956(.A1(new_n14086_), .A2(new_n14082_), .ZN(new_n14150_));
  NOR2_X1    g13957(.A1(new_n5175_), .A2(new_n7643_), .ZN(new_n14151_));
  INV_X1     g13958(.I(new_n14151_), .ZN(new_n14152_));
  XOR2_X1    g13959(.A1(new_n14092_), .A2(new_n14152_), .Z(new_n14153_));
  XNOR2_X1   g13960(.A1(new_n14153_), .A2(new_n14150_), .ZN(new_n14154_));
  NOR2_X1    g13961(.A1(new_n14149_), .A2(new_n14154_), .ZN(new_n14155_));
  NAND2_X1   g13962(.A1(new_n14149_), .A2(new_n14154_), .ZN(new_n14156_));
  INV_X1     g13963(.I(new_n14156_), .ZN(new_n14157_));
  NOR2_X1    g13964(.A1(new_n14157_), .A2(new_n14155_), .ZN(new_n14158_));
  NAND2_X1   g13965(.A1(new_n14158_), .A2(new_n14146_), .ZN(new_n14159_));
  INV_X1     g13966(.I(new_n14159_), .ZN(new_n14160_));
  NOR2_X1    g13967(.A1(new_n14158_), .A2(new_n14146_), .ZN(new_n14161_));
  NOR2_X1    g13968(.A1(new_n14160_), .A2(new_n14161_), .ZN(new_n14162_));
  NOR2_X1    g13969(.A1(new_n14127_), .A2(new_n14162_), .ZN(new_n14163_));
  NAND2_X1   g13970(.A1(new_n14127_), .A2(new_n14162_), .ZN(new_n14164_));
  INV_X1     g13971(.I(new_n14164_), .ZN(new_n14165_));
  NOR2_X1    g13972(.A1(new_n14165_), .A2(new_n14163_), .ZN(new_n14166_));
  XOR2_X1    g13973(.A1(new_n14124_), .A2(new_n14166_), .Z(\asquared[116] ));
  AOI21_X1   g13974(.A1(new_n14123_), .A2(new_n14115_), .B(new_n14163_), .ZN(new_n14168_));
  NOR2_X1    g13975(.A1(new_n14168_), .A2(new_n14165_), .ZN(new_n14169_));
  OAI22_X1   g13976(.A1(new_n6899_), .A2(new_n8952_), .B1(new_n7185_), .B2(new_n7454_), .ZN(new_n14170_));
  OAI21_X1   g13977(.A1(new_n8161_), .A2(new_n7452_), .B(new_n14170_), .ZN(new_n14171_));
  NOR2_X1    g13978(.A1(new_n8161_), .A2(new_n7452_), .ZN(new_n14172_));
  NOR2_X1    g13979(.A1(new_n14170_), .A2(new_n14172_), .ZN(new_n14173_));
  AOI21_X1   g13980(.A1(\a[56] ), .A2(\a[60] ), .B(new_n7203_), .ZN(new_n14174_));
  INV_X1     g13981(.I(new_n14174_), .ZN(new_n14175_));
  NOR2_X1    g13982(.A1(new_n5680_), .A2(new_n6897_), .ZN(new_n14176_));
  AOI22_X1   g13983(.A1(new_n14173_), .A2(new_n14175_), .B1(new_n14171_), .B2(new_n14176_), .ZN(new_n14177_));
  NOR2_X1    g13984(.A1(new_n14177_), .A2(new_n14136_), .ZN(new_n14178_));
  INV_X1     g13985(.I(new_n14178_), .ZN(new_n14179_));
  AND2_X2    g13986(.A1(new_n14177_), .A2(new_n14136_), .Z(new_n14180_));
  INV_X1     g13987(.I(new_n14180_), .ZN(new_n14181_));
  NAND2_X1   g13988(.A1(new_n6126_), .A2(new_n7644_), .ZN(new_n14182_));
  NOR2_X1    g13989(.A1(new_n5617_), .A2(new_n7144_), .ZN(new_n14183_));
  NOR2_X1    g13990(.A1(new_n5425_), .A2(new_n7643_), .ZN(new_n14184_));
  OAI21_X1   g13991(.A1(new_n14183_), .A2(new_n14184_), .B(new_n14182_), .ZN(new_n14185_));
  XNOR2_X1   g13992(.A1(new_n14185_), .A2(new_n14143_), .ZN(new_n14186_));
  AOI21_X1   g13993(.A1(new_n14181_), .A2(new_n14179_), .B(new_n14186_), .ZN(new_n14187_));
  INV_X1     g13994(.I(new_n14187_), .ZN(new_n14188_));
  NAND3_X1   g13995(.A1(new_n14181_), .A2(new_n14179_), .A3(new_n14186_), .ZN(new_n14189_));
  NAND2_X1   g13996(.A1(new_n14188_), .A2(new_n14189_), .ZN(new_n14190_));
  INV_X1     g13997(.I(new_n14190_), .ZN(new_n14191_));
  INV_X1     g13998(.I(new_n14144_), .ZN(new_n14192_));
  NOR2_X1    g13999(.A1(new_n14145_), .A2(new_n14129_), .ZN(new_n14193_));
  AOI21_X1   g14000(.A1(new_n14137_), .A2(new_n14192_), .B(new_n14193_), .ZN(new_n14194_));
  NOR2_X1    g14001(.A1(new_n14092_), .A2(new_n14152_), .ZN(new_n14195_));
  INV_X1     g14002(.I(new_n14153_), .ZN(new_n14196_));
  NOR2_X1    g14003(.A1(new_n14196_), .A2(new_n14150_), .ZN(new_n14197_));
  NOR2_X1    g14004(.A1(new_n14197_), .A2(new_n14195_), .ZN(new_n14198_));
  XOR2_X1    g14005(.A1(new_n14194_), .A2(new_n14198_), .Z(new_n14199_));
  XOR2_X1    g14006(.A1(new_n14199_), .A2(new_n14191_), .Z(new_n14200_));
  NOR2_X1    g14007(.A1(new_n14160_), .A2(new_n14157_), .ZN(new_n14201_));
  INV_X1     g14008(.I(new_n14201_), .ZN(new_n14202_));
  NAND2_X1   g14009(.A1(new_n14202_), .A2(new_n14200_), .ZN(new_n14203_));
  NOR2_X1    g14010(.A1(new_n14202_), .A2(new_n14200_), .ZN(new_n14204_));
  INV_X1     g14011(.I(new_n14204_), .ZN(new_n14205_));
  NAND2_X1   g14012(.A1(new_n14205_), .A2(new_n14203_), .ZN(new_n14206_));
  INV_X1     g14013(.I(new_n14115_), .ZN(new_n14207_));
  INV_X1     g14014(.I(new_n14163_), .ZN(new_n14208_));
  OAI21_X1   g14015(.A1(new_n14121_), .A2(new_n14207_), .B(new_n14208_), .ZN(new_n14209_));
  AOI21_X1   g14016(.A1(new_n14209_), .A2(new_n14164_), .B(new_n14204_), .ZN(new_n14210_));
  AOI22_X1   g14017(.A1(new_n14210_), .A2(new_n14203_), .B1(new_n14169_), .B2(new_n14206_), .ZN(\asquared[117] ));
  OAI21_X1   g14018(.A1(new_n14168_), .A2(new_n14165_), .B(new_n14205_), .ZN(new_n14212_));
  NAND2_X1   g14019(.A1(new_n14212_), .A2(new_n14203_), .ZN(new_n14213_));
  NOR2_X1    g14020(.A1(new_n14194_), .A2(new_n14198_), .ZN(new_n14214_));
  AOI21_X1   g14021(.A1(new_n14199_), .A2(new_n14191_), .B(new_n14214_), .ZN(new_n14215_));
  OAI21_X1   g14022(.A1(new_n14185_), .A2(new_n14143_), .B(new_n14182_), .ZN(new_n14216_));
  XNOR2_X1   g14023(.A1(new_n14216_), .A2(new_n14173_), .ZN(new_n14217_));
  NAND2_X1   g14024(.A1(new_n5857_), .A2(new_n7852_), .ZN(new_n14218_));
  NAND2_X1   g14025(.A1(new_n9030_), .A2(new_n10611_), .ZN(new_n14219_));
  AOI22_X1   g14026(.A1(new_n14218_), .A2(new_n14219_), .B1(new_n6494_), .B2(new_n7453_), .ZN(new_n14220_));
  NAND2_X1   g14027(.A1(\a[54] ), .A2(\a[63] ), .ZN(new_n14221_));
  AOI22_X1   g14028(.A1(\a[56] ), .A2(\a[61] ), .B1(\a[57] ), .B2(\a[60] ), .ZN(new_n14222_));
  NAND2_X1   g14029(.A1(new_n6494_), .A2(new_n7453_), .ZN(new_n14223_));
  NAND3_X1   g14030(.A1(new_n14223_), .A2(new_n14218_), .A3(new_n14219_), .ZN(new_n14224_));
  OAI22_X1   g14031(.A1(new_n14220_), .A2(new_n14221_), .B1(new_n14224_), .B2(new_n14222_), .ZN(new_n14225_));
  XOR2_X1    g14032(.A1(new_n14217_), .A2(new_n14225_), .Z(new_n14226_));
  NOR2_X1    g14033(.A1(new_n12459_), .A2(new_n5680_), .ZN(new_n14227_));
  NAND2_X1   g14034(.A1(new_n14227_), .A2(new_n7205_), .ZN(new_n14228_));
  AOI21_X1   g14035(.A1(\a[55] ), .A2(\a[62] ), .B(\a[59] ), .ZN(new_n14229_));
  NOR2_X1    g14036(.A1(new_n14227_), .A2(new_n7205_), .ZN(new_n14230_));
  INV_X1     g14037(.I(new_n14230_), .ZN(new_n14231_));
  OAI21_X1   g14038(.A1(new_n14231_), .A2(new_n14229_), .B(new_n14228_), .ZN(new_n14232_));
  INV_X1     g14039(.I(new_n14136_), .ZN(new_n14233_));
  OAI21_X1   g14040(.A1(new_n14233_), .A2(new_n14177_), .B(new_n14188_), .ZN(new_n14234_));
  XOR2_X1    g14041(.A1(new_n14234_), .A2(new_n14232_), .Z(new_n14235_));
  XNOR2_X1   g14042(.A1(new_n14235_), .A2(new_n14226_), .ZN(new_n14236_));
  NAND2_X1   g14043(.A1(new_n14236_), .A2(new_n14215_), .ZN(new_n14237_));
  INV_X1     g14044(.I(new_n14237_), .ZN(new_n14238_));
  NOR2_X1    g14045(.A1(new_n14236_), .A2(new_n14215_), .ZN(new_n14239_));
  NOR2_X1    g14046(.A1(new_n14238_), .A2(new_n14239_), .ZN(new_n14240_));
  XOR2_X1    g14047(.A1(new_n14213_), .A2(new_n14240_), .Z(\asquared[118] ));
  AOI21_X1   g14048(.A1(new_n14212_), .A2(new_n14203_), .B(new_n14238_), .ZN(new_n14242_));
  NOR2_X1    g14049(.A1(new_n14242_), .A2(new_n14239_), .ZN(new_n14243_));
  NAND2_X1   g14050(.A1(new_n14234_), .A2(new_n14232_), .ZN(new_n14244_));
  NAND2_X1   g14051(.A1(new_n14235_), .A2(new_n14226_), .ZN(new_n14245_));
  NAND2_X1   g14052(.A1(new_n14245_), .A2(new_n14244_), .ZN(new_n14246_));
  AOI21_X1   g14053(.A1(\a[55] ), .A2(\a[63] ), .B(new_n14231_), .ZN(new_n14247_));
  NOR3_X1    g14054(.A1(new_n14230_), .A2(new_n5680_), .A3(new_n7643_), .ZN(new_n14248_));
  NOR2_X1    g14055(.A1(new_n14247_), .A2(new_n14248_), .ZN(new_n14249_));
  XOR2_X1    g14056(.A1(new_n14249_), .A2(new_n14224_), .Z(new_n14250_));
  OAI21_X1   g14057(.A1(new_n14172_), .A2(new_n14170_), .B(new_n14216_), .ZN(new_n14251_));
  NAND2_X1   g14058(.A1(new_n14217_), .A2(new_n14225_), .ZN(new_n14252_));
  NAND2_X1   g14059(.A1(new_n14252_), .A2(new_n14251_), .ZN(new_n14253_));
  NOR2_X1    g14060(.A1(new_n6804_), .A2(new_n7454_), .ZN(new_n14254_));
  AOI22_X1   g14061(.A1(new_n6494_), .A2(new_n7590_), .B1(new_n7800_), .B2(new_n13932_), .ZN(new_n14255_));
  NOR2_X1    g14062(.A1(new_n14254_), .A2(new_n14255_), .ZN(new_n14256_));
  AOI21_X1   g14063(.A1(\a[57] ), .A2(\a[61] ), .B(new_n7800_), .ZN(new_n14257_));
  NOR2_X1    g14064(.A1(new_n14256_), .A2(new_n14254_), .ZN(new_n14258_));
  INV_X1     g14065(.I(new_n14258_), .ZN(new_n14259_));
  OAI22_X1   g14066(.A1(new_n14259_), .A2(new_n14257_), .B1(new_n13933_), .B2(new_n14256_), .ZN(new_n14260_));
  XNOR2_X1   g14067(.A1(new_n14253_), .A2(new_n14260_), .ZN(new_n14261_));
  XNOR2_X1   g14068(.A1(new_n14261_), .A2(new_n14250_), .ZN(new_n14262_));
  NOR2_X1    g14069(.A1(new_n14246_), .A2(new_n14262_), .ZN(new_n14263_));
  INV_X1     g14070(.I(new_n14263_), .ZN(new_n14264_));
  NAND2_X1   g14071(.A1(new_n14246_), .A2(new_n14262_), .ZN(new_n14265_));
  NAND2_X1   g14072(.A1(new_n14264_), .A2(new_n14265_), .ZN(new_n14266_));
  XOR2_X1    g14073(.A1(new_n14243_), .A2(new_n14266_), .Z(\asquared[119] ));
  OAI21_X1   g14074(.A1(new_n14242_), .A2(new_n14239_), .B(new_n14264_), .ZN(new_n14268_));
  NAND2_X1   g14075(.A1(new_n14268_), .A2(new_n14265_), .ZN(new_n14269_));
  INV_X1     g14076(.I(new_n14248_), .ZN(new_n14270_));
  NAND2_X1   g14077(.A1(new_n14249_), .A2(new_n14224_), .ZN(new_n14271_));
  NAND2_X1   g14078(.A1(new_n14271_), .A2(new_n14270_), .ZN(new_n14272_));
  NOR2_X1    g14079(.A1(new_n7146_), .A2(new_n6298_), .ZN(new_n14273_));
  NAND2_X1   g14080(.A1(new_n14273_), .A2(new_n7451_), .ZN(new_n14274_));
  AOI21_X1   g14081(.A1(\a[57] ), .A2(\a[62] ), .B(\a[60] ), .ZN(new_n14275_));
  NOR2_X1    g14082(.A1(new_n14273_), .A2(new_n7451_), .ZN(new_n14276_));
  INV_X1     g14083(.I(new_n14276_), .ZN(new_n14277_));
  OAI21_X1   g14084(.A1(new_n14277_), .A2(new_n14275_), .B(new_n14274_), .ZN(new_n14278_));
  INV_X1     g14085(.I(new_n14278_), .ZN(new_n14279_));
  NOR2_X1    g14086(.A1(new_n6318_), .A2(new_n7959_), .ZN(new_n14280_));
  INV_X1     g14087(.I(new_n14280_), .ZN(new_n14281_));
  NOR2_X1    g14088(.A1(new_n6316_), .A2(new_n6897_), .ZN(new_n14282_));
  NOR2_X1    g14089(.A1(new_n5856_), .A2(new_n7643_), .ZN(new_n14283_));
  OAI21_X1   g14090(.A1(new_n14282_), .A2(new_n14283_), .B(new_n14281_), .ZN(new_n14284_));
  XNOR2_X1   g14091(.A1(new_n14284_), .A2(new_n14258_), .ZN(new_n14285_));
  XOR2_X1    g14092(.A1(new_n14285_), .A2(new_n14279_), .Z(new_n14286_));
  XOR2_X1    g14093(.A1(new_n14286_), .A2(new_n14272_), .Z(new_n14287_));
  NAND2_X1   g14094(.A1(new_n14253_), .A2(new_n14260_), .ZN(new_n14288_));
  INV_X1     g14095(.I(new_n14261_), .ZN(new_n14289_));
  NAND2_X1   g14096(.A1(new_n14289_), .A2(new_n14250_), .ZN(new_n14290_));
  NAND2_X1   g14097(.A1(new_n14290_), .A2(new_n14288_), .ZN(new_n14291_));
  NOR2_X1    g14098(.A1(new_n14291_), .A2(new_n14287_), .ZN(new_n14292_));
  NAND2_X1   g14099(.A1(new_n14291_), .A2(new_n14287_), .ZN(new_n14293_));
  INV_X1     g14100(.I(new_n14293_), .ZN(new_n14294_));
  NOR2_X1    g14101(.A1(new_n14294_), .A2(new_n14292_), .ZN(new_n14295_));
  XOR2_X1    g14102(.A1(new_n14269_), .A2(new_n14295_), .Z(\asquared[120] ));
  AOI21_X1   g14103(.A1(new_n14268_), .A2(new_n14265_), .B(new_n14292_), .ZN(new_n14297_));
  NOR2_X1    g14104(.A1(new_n14297_), .A2(new_n14294_), .ZN(new_n14298_));
  NAND2_X1   g14105(.A1(new_n6803_), .A2(new_n7644_), .ZN(new_n14299_));
  NAND2_X1   g14106(.A1(new_n7203_), .A2(new_n7852_), .ZN(new_n14300_));
  AOI22_X1   g14107(.A1(new_n14299_), .A2(new_n14300_), .B1(new_n7205_), .B2(new_n7590_), .ZN(new_n14301_));
  NAND2_X1   g14108(.A1(new_n7205_), .A2(new_n7590_), .ZN(new_n14302_));
  NAND3_X1   g14109(.A1(new_n14302_), .A2(new_n14299_), .A3(new_n14300_), .ZN(new_n14303_));
  AOI21_X1   g14110(.A1(\a[58] ), .A2(\a[62] ), .B(new_n6898_), .ZN(new_n14304_));
  NAND2_X1   g14111(.A1(\a[57] ), .A2(\a[63] ), .ZN(new_n14305_));
  OAI22_X1   g14112(.A1(new_n14301_), .A2(new_n14305_), .B1(new_n14303_), .B2(new_n14304_), .ZN(new_n14306_));
  OAI21_X1   g14113(.A1(new_n14284_), .A2(new_n14258_), .B(new_n14281_), .ZN(new_n14307_));
  NOR2_X1    g14114(.A1(new_n14307_), .A2(new_n14277_), .ZN(new_n14308_));
  AND2_X2    g14115(.A1(new_n14307_), .A2(new_n14277_), .Z(new_n14309_));
  NOR2_X1    g14116(.A1(new_n14309_), .A2(new_n14308_), .ZN(new_n14310_));
  NOR2_X1    g14117(.A1(new_n14310_), .A2(new_n14306_), .ZN(new_n14311_));
  AND2_X2    g14118(.A1(new_n14310_), .A2(new_n14306_), .Z(new_n14312_));
  NOR2_X1    g14119(.A1(new_n14312_), .A2(new_n14311_), .ZN(new_n14313_));
  INV_X1     g14120(.I(new_n14313_), .ZN(new_n14314_));
  OR2_X2     g14121(.A1(new_n14285_), .A2(new_n14279_), .Z(new_n14315_));
  NAND2_X1   g14122(.A1(new_n14286_), .A2(new_n14272_), .ZN(new_n14316_));
  NAND2_X1   g14123(.A1(new_n14316_), .A2(new_n14315_), .ZN(new_n14317_));
  INV_X1     g14124(.I(new_n14317_), .ZN(new_n14318_));
  NOR2_X1    g14125(.A1(new_n14318_), .A2(new_n14314_), .ZN(new_n14319_));
  INV_X1     g14126(.I(new_n14319_), .ZN(new_n14320_));
  NOR2_X1    g14127(.A1(new_n14317_), .A2(new_n14313_), .ZN(new_n14321_));
  INV_X1     g14128(.I(new_n14321_), .ZN(new_n14322_));
  NAND2_X1   g14129(.A1(new_n14320_), .A2(new_n14322_), .ZN(new_n14323_));
  INV_X1     g14130(.I(new_n14265_), .ZN(new_n14324_));
  INV_X1     g14131(.I(new_n14239_), .ZN(new_n14325_));
  INV_X1     g14132(.I(new_n14203_), .ZN(new_n14326_));
  OAI21_X1   g14133(.A1(new_n14210_), .A2(new_n14326_), .B(new_n14237_), .ZN(new_n14327_));
  AOI21_X1   g14134(.A1(new_n14327_), .A2(new_n14325_), .B(new_n14263_), .ZN(new_n14328_));
  INV_X1     g14135(.I(new_n14292_), .ZN(new_n14329_));
  OAI21_X1   g14136(.A1(new_n14328_), .A2(new_n14324_), .B(new_n14329_), .ZN(new_n14330_));
  AOI21_X1   g14137(.A1(new_n14330_), .A2(new_n14293_), .B(new_n14321_), .ZN(new_n14331_));
  AOI22_X1   g14138(.A1(new_n14331_), .A2(new_n14320_), .B1(new_n14298_), .B2(new_n14323_), .ZN(\asquared[121] ));
  OAI21_X1   g14139(.A1(new_n14297_), .A2(new_n14294_), .B(new_n14322_), .ZN(new_n14333_));
  NAND2_X1   g14140(.A1(new_n14333_), .A2(new_n14320_), .ZN(new_n14334_));
  NOR2_X1    g14141(.A1(new_n14312_), .A2(new_n14309_), .ZN(new_n14335_));
  NOR2_X1    g14142(.A1(new_n6897_), .A2(\a[60] ), .ZN(new_n14336_));
  XOR2_X1    g14143(.A1(new_n12458_), .A2(new_n14336_), .Z(new_n14337_));
  XOR2_X1    g14144(.A1(new_n14303_), .A2(new_n13666_), .Z(new_n14338_));
  XNOR2_X1   g14145(.A1(new_n14338_), .A2(new_n14337_), .ZN(new_n14339_));
  NAND2_X1   g14146(.A1(new_n14335_), .A2(new_n14339_), .ZN(new_n14340_));
  INV_X1     g14147(.I(new_n14340_), .ZN(new_n14341_));
  NOR2_X1    g14148(.A1(new_n14335_), .A2(new_n14339_), .ZN(new_n14342_));
  NOR2_X1    g14149(.A1(new_n14341_), .A2(new_n14342_), .ZN(new_n14343_));
  XOR2_X1    g14150(.A1(new_n14334_), .A2(new_n14343_), .Z(\asquared[122] ));
  AOI21_X1   g14151(.A1(new_n14333_), .A2(new_n14320_), .B(new_n14341_), .ZN(new_n14345_));
  NOR2_X1    g14152(.A1(new_n14345_), .A2(new_n14342_), .ZN(new_n14346_));
  NAND2_X1   g14153(.A1(new_n14303_), .A2(new_n13666_), .ZN(new_n14347_));
  NAND2_X1   g14154(.A1(new_n14338_), .A2(new_n14337_), .ZN(new_n14348_));
  NAND2_X1   g14155(.A1(new_n14348_), .A2(new_n14347_), .ZN(new_n14349_));
  NAND2_X1   g14156(.A1(new_n7146_), .A2(new_n13663_), .ZN(new_n14350_));
  INV_X1     g14157(.I(new_n14350_), .ZN(new_n14351_));
  OAI21_X1   g14158(.A1(new_n12458_), .A2(\a[60] ), .B(\a[61] ), .ZN(new_n14352_));
  NOR2_X1    g14159(.A1(new_n7452_), .A2(new_n8049_), .ZN(new_n14353_));
  NOR2_X1    g14160(.A1(new_n14351_), .A2(new_n14353_), .ZN(new_n14354_));
  INV_X1     g14161(.I(new_n14352_), .ZN(new_n14355_));
  AOI21_X1   g14162(.A1(new_n14350_), .A2(new_n14355_), .B(new_n14353_), .ZN(new_n14356_));
  INV_X1     g14163(.I(new_n14356_), .ZN(new_n14357_));
  OAI22_X1   g14164(.A1(new_n14357_), .A2(new_n14351_), .B1(new_n14352_), .B2(new_n14354_), .ZN(new_n14358_));
  NAND2_X1   g14165(.A1(new_n14349_), .A2(new_n14358_), .ZN(new_n14359_));
  NOR2_X1    g14166(.A1(new_n14349_), .A2(new_n14358_), .ZN(new_n14360_));
  INV_X1     g14167(.I(new_n14360_), .ZN(new_n14361_));
  NAND2_X1   g14168(.A1(new_n14361_), .A2(new_n14359_), .ZN(new_n14362_));
  INV_X1     g14169(.I(new_n14342_), .ZN(new_n14363_));
  OAI21_X1   g14170(.A1(new_n14331_), .A2(new_n14319_), .B(new_n14340_), .ZN(new_n14364_));
  AOI21_X1   g14171(.A1(new_n14364_), .A2(new_n14363_), .B(new_n14360_), .ZN(new_n14365_));
  AOI22_X1   g14172(.A1(new_n14365_), .A2(new_n14359_), .B1(new_n14346_), .B2(new_n14362_), .ZN(\asquared[123] ));
  OAI21_X1   g14173(.A1(new_n14345_), .A2(new_n14342_), .B(new_n14361_), .ZN(new_n14367_));
  NAND2_X1   g14174(.A1(new_n14367_), .A2(new_n14359_), .ZN(new_n14368_));
  NOR2_X1    g14175(.A1(new_n7144_), .A2(\a[61] ), .ZN(new_n14369_));
  NOR2_X1    g14176(.A1(new_n9030_), .A2(new_n14369_), .ZN(new_n14370_));
  INV_X1     g14177(.I(new_n14369_), .ZN(new_n14371_));
  NOR2_X1    g14178(.A1(new_n9031_), .A2(new_n14371_), .ZN(new_n14372_));
  NOR2_X1    g14179(.A1(new_n14372_), .A2(new_n14370_), .ZN(new_n14373_));
  NOR2_X1    g14180(.A1(new_n14357_), .A2(new_n14373_), .ZN(new_n14374_));
  NAND2_X1   g14181(.A1(new_n14357_), .A2(new_n14373_), .ZN(new_n14375_));
  INV_X1     g14182(.I(new_n14375_), .ZN(new_n14376_));
  NOR2_X1    g14183(.A1(new_n14376_), .A2(new_n14374_), .ZN(new_n14377_));
  XOR2_X1    g14184(.A1(new_n14368_), .A2(new_n14377_), .Z(\asquared[124] ));
  AOI21_X1   g14185(.A1(new_n14367_), .A2(new_n14359_), .B(new_n14374_), .ZN(new_n14379_));
  NOR2_X1    g14186(.A1(new_n14379_), .A2(new_n14376_), .ZN(new_n14380_));
  NOR3_X1    g14187(.A1(new_n14372_), .A2(new_n7590_), .A3(new_n7852_), .ZN(new_n14381_));
  NOR2_X1    g14188(.A1(new_n7959_), .A2(new_n7144_), .ZN(new_n14382_));
  NOR2_X1    g14189(.A1(new_n14381_), .A2(new_n14382_), .ZN(new_n14383_));
  INV_X1     g14190(.I(new_n14383_), .ZN(new_n14384_));
  XOR2_X1    g14191(.A1(new_n14380_), .A2(new_n14384_), .Z(\asquared[125] ));
  NOR2_X1    g14192(.A1(new_n7643_), .A2(\a[62] ), .ZN(new_n14386_));
  INV_X1     g14193(.I(new_n14359_), .ZN(new_n14387_));
  INV_X1     g14194(.I(new_n14374_), .ZN(new_n14388_));
  OAI21_X1   g14195(.A1(new_n14365_), .A2(new_n14387_), .B(new_n14388_), .ZN(new_n14389_));
  AOI21_X1   g14196(.A1(new_n14389_), .A2(new_n14375_), .B(new_n14381_), .ZN(new_n14390_));
  NOR3_X1    g14197(.A1(new_n14390_), .A2(new_n14382_), .A3(new_n14386_), .ZN(new_n14391_));
  INV_X1     g14198(.I(new_n14382_), .ZN(new_n14392_));
  INV_X1     g14199(.I(new_n14386_), .ZN(new_n14393_));
  INV_X1     g14200(.I(new_n14381_), .ZN(new_n14394_));
  OAI21_X1   g14201(.A1(new_n14379_), .A2(new_n14376_), .B(new_n14394_), .ZN(new_n14395_));
  AOI21_X1   g14202(.A1(new_n14395_), .A2(new_n14392_), .B(new_n14393_), .ZN(new_n14396_));
  NOR2_X1    g14203(.A1(new_n14391_), .A2(new_n14396_), .ZN(\asquared[126] ));
  OAI21_X1   g14204(.A1(new_n14390_), .A2(new_n14382_), .B(\a[63] ), .ZN(new_n14398_));
  NAND2_X1   g14205(.A1(new_n14398_), .A2(new_n8049_), .ZN(\asquared[127] ));
  assign     \asquared[1]  = 1'b0;
  BUF_X16    g14206(.I(\a[0] ), .Z(\asquared[0] ));
endmodule


