// Benchmark "i3" written by ABC on Fri Feb 25 15:12:56 2022

module i3 ( 
    \V56(0) , \V28(0) , \V56(1) , \V28(1) , \V56(2) , \V28(2) , \V56(3) ,
    \V28(3) , \V56(4) , \V28(4) , \V56(5) , \V28(5) , \V56(6) , \V28(6) ,
    \V56(7) , \V28(7) , \V56(8) , \V28(8) , \V56(9) , \V28(9) , \V56(10) ,
    \V28(10) , \V56(11) , \V28(11) , \V56(12) , \V28(12) , \V56(13) ,
    \V28(13) , \V56(14) , \V28(14) , \V56(15) , \V28(15) , \V56(16) ,
    \V28(16) , \V56(17) , \V28(17) , \V56(18) , \V28(18) , \V56(19) ,
    \V28(19) , \V56(20) , \V28(20) , \V56(21) , \V28(21) , \V56(22) ,
    \V28(22) , \V56(23) , \V28(23) , \V56(24) , \V28(24) , \V56(25) ,
    \V28(25) , \V56(26) , \V28(26) , \V56(27) , \V28(27) , \V120(0) ,
    \V88(0) , \V120(1) , \V88(1) , \V120(2) , \V88(2) , \V120(3) ,
    \V88(3) , \V120(4) , \V88(4) , \V120(5) , \V88(5) , \V120(6) ,
    \V88(6) , \V120(7) , \V88(7) , \V120(8) , \V88(8) , \V120(9) ,
    \V88(9) , \V120(10) , \V88(10) , \V120(11) , \V88(11) , \V120(12) ,
    \V88(12) , \V120(13) , \V88(13) , \V120(14) , \V88(14) , \V120(15) ,
    \V88(15) , \V120(16) , \V88(16) , \V120(17) , \V88(17) , \V120(18) ,
    \V88(18) , \V120(19) , \V88(19) , \V120(20) , \V88(20) , \V120(21) ,
    \V88(21) , \V120(22) , \V88(22) , \V120(23) , \V88(23) , \V120(24) ,
    \V88(24) , \V120(25) , \V88(25) , \V120(26) , \V88(26) , \V120(27) ,
    \V88(27) , \V120(28) , \V88(28) , \V120(29) , \V88(29) , \V120(30) ,
    \V88(30) , \V120(31) , \V88(31) , \V132(0) , \V126(0) , \V132(1) ,
    \V126(1) , \V132(2) , \V126(2) , \V132(3) , \V126(3) , \V132(4) ,
    \V126(4) , \V132(5) , \V126(5) ,
    \V134(0) , \V134(1) , \V138(0) , \V138(1) , \V138(2) , \V138(3)   );
  input  \V56(0) , \V28(0) , \V56(1) , \V28(1) , \V56(2) , \V28(2) ,
    \V56(3) , \V28(3) , \V56(4) , \V28(4) , \V56(5) , \V28(5) , \V56(6) ,
    \V28(6) , \V56(7) , \V28(7) , \V56(8) , \V28(8) , \V56(9) , \V28(9) ,
    \V56(10) , \V28(10) , \V56(11) , \V28(11) , \V56(12) , \V28(12) ,
    \V56(13) , \V28(13) , \V56(14) , \V28(14) , \V56(15) , \V28(15) ,
    \V56(16) , \V28(16) , \V56(17) , \V28(17) , \V56(18) , \V28(18) ,
    \V56(19) , \V28(19) , \V56(20) , \V28(20) , \V56(21) , \V28(21) ,
    \V56(22) , \V28(22) , \V56(23) , \V28(23) , \V56(24) , \V28(24) ,
    \V56(25) , \V28(25) , \V56(26) , \V28(26) , \V56(27) , \V28(27) ,
    \V120(0) , \V88(0) , \V120(1) , \V88(1) , \V120(2) , \V88(2) ,
    \V120(3) , \V88(3) , \V120(4) , \V88(4) , \V120(5) , \V88(5) ,
    \V120(6) , \V88(6) , \V120(7) , \V88(7) , \V120(8) , \V88(8) ,
    \V120(9) , \V88(9) , \V120(10) , \V88(10) , \V120(11) , \V88(11) ,
    \V120(12) , \V88(12) , \V120(13) , \V88(13) , \V120(14) , \V88(14) ,
    \V120(15) , \V88(15) , \V120(16) , \V88(16) , \V120(17) , \V88(17) ,
    \V120(18) , \V88(18) , \V120(19) , \V88(19) , \V120(20) , \V88(20) ,
    \V120(21) , \V88(21) , \V120(22) , \V88(22) , \V120(23) , \V88(23) ,
    \V120(24) , \V88(24) , \V120(25) , \V88(25) , \V120(26) , \V88(26) ,
    \V120(27) , \V88(27) , \V120(28) , \V88(28) , \V120(29) , \V88(29) ,
    \V120(30) , \V88(30) , \V120(31) , \V88(31) , \V132(0) , \V126(0) ,
    \V132(1) , \V126(1) , \V132(2) , \V126(2) , \V132(3) , \V126(3) ,
    \V132(4) , \V126(4) , \V132(5) , \V126(5) ;
  output \V134(0) , \V134(1) , \V138(0) , \V138(1) , \V138(2) , \V138(3) ;
  wire new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_;
  assign \V134(0)  = \V56(0)  | \V28(0) ;
  assign \V134(1)  = \V56(1)  | \V28(1) ;
  assign new_n141_ = ~\V56(17)  & ~\V28(17) ;
  assign new_n142_ = ~\V56(16)  & ~\V28(16) ;
  assign new_n143_ = ~\V56(14)  & ~\V28(14) ;
  assign new_n144_ = ~\V56(15)  & ~\V28(15) ;
  assign new_n145_ = ~\V56(5)  & ~\V28(5) ;
  assign new_n146_ = ~\V56(4)  & ~\V28(4) ;
  assign new_n147_ = ~\V56(2)  & ~\V28(2) ;
  assign new_n148_ = ~\V56(3)  & ~\V28(3) ;
  assign new_n149_ = ~\V56(8)  & ~\V28(8) ;
  assign new_n150_ = ~\V56(6)  & ~\V28(6) ;
  assign new_n151_ = ~\V56(7)  & ~\V28(7) ;
  assign new_n152_ = ~\V56(9)  & ~\V28(9) ;
  assign new_n153_ = ~\V56(11)  & ~\V28(11) ;
  assign new_n154_ = ~\V56(10)  & ~\V28(10) ;
  assign new_n155_ = ~\V56(12)  & ~\V28(12) ;
  assign new_n156_ = ~\V56(13)  & ~\V28(13) ;
  assign new_n157_ = ~new_n141_ & ~new_n142_;
  assign new_n158_ = ~new_n143_ & new_n157_;
  assign new_n159_ = ~new_n144_ & new_n158_;
  assign new_n160_ = ~new_n145_ & new_n159_;
  assign new_n161_ = ~new_n146_ & new_n160_;
  assign new_n162_ = ~new_n147_ & new_n161_;
  assign new_n163_ = ~new_n148_ & new_n162_;
  assign new_n164_ = ~new_n149_ & new_n163_;
  assign new_n165_ = ~new_n150_ & new_n164_;
  assign new_n166_ = ~new_n151_ & new_n165_;
  assign new_n167_ = ~new_n152_ & new_n166_;
  assign new_n168_ = ~new_n153_ & new_n167_;
  assign new_n169_ = ~new_n154_ & new_n168_;
  assign new_n170_ = ~new_n155_ & new_n169_;
  assign \V138(0)  = ~new_n156_ & new_n170_;
  assign new_n172_ = ~\V120(5)  & ~\V88(5) ;
  assign new_n173_ = ~\V120(4)  & ~\V88(4) ;
  assign new_n174_ = ~\V120(2)  & ~\V88(2) ;
  assign new_n175_ = ~\V120(3)  & ~\V88(3) ;
  assign new_n176_ = ~\V56(21)  & ~\V28(21) ;
  assign new_n177_ = ~\V56(20)  & ~\V28(20) ;
  assign new_n178_ = ~\V56(18)  & ~\V28(18) ;
  assign new_n179_ = ~\V56(19)  & ~\V28(19) ;
  assign new_n180_ = ~\V56(24)  & ~\V28(24) ;
  assign new_n181_ = ~\V56(22)  & ~\V28(22) ;
  assign new_n182_ = ~\V56(23)  & ~\V28(23) ;
  assign new_n183_ = ~\V56(25)  & ~\V28(25) ;
  assign new_n184_ = ~\V56(27)  & ~\V28(27) ;
  assign new_n185_ = ~\V56(26)  & ~\V28(26) ;
  assign new_n186_ = ~\V120(0)  & ~\V88(0) ;
  assign new_n187_ = ~\V120(1)  & ~\V88(1) ;
  assign new_n188_ = ~new_n172_ & ~new_n173_;
  assign new_n189_ = ~new_n174_ & new_n188_;
  assign new_n190_ = ~new_n175_ & new_n189_;
  assign new_n191_ = ~new_n176_ & new_n190_;
  assign new_n192_ = ~new_n177_ & new_n191_;
  assign new_n193_ = ~new_n178_ & new_n192_;
  assign new_n194_ = ~new_n179_ & new_n193_;
  assign new_n195_ = ~new_n180_ & new_n194_;
  assign new_n196_ = ~new_n181_ & new_n195_;
  assign new_n197_ = ~new_n182_ & new_n196_;
  assign new_n198_ = ~new_n183_ & new_n197_;
  assign new_n199_ = ~new_n184_ & new_n198_;
  assign new_n200_ = ~new_n185_ & new_n199_;
  assign new_n201_ = ~new_n186_ & new_n200_;
  assign \V138(1)  = ~new_n187_ & new_n201_;
  assign new_n203_ = ~\V120(21)  & ~\V88(21) ;
  assign new_n204_ = ~\V120(20)  & ~\V88(20) ;
  assign new_n205_ = ~\V120(18)  & ~\V88(18) ;
  assign new_n206_ = ~\V120(19)  & ~\V88(19) ;
  assign new_n207_ = ~\V120(9)  & ~\V88(9) ;
  assign new_n208_ = ~\V120(8)  & ~\V88(8) ;
  assign new_n209_ = ~\V120(6)  & ~\V88(6) ;
  assign new_n210_ = ~\V120(7)  & ~\V88(7) ;
  assign new_n211_ = ~\V120(12)  & ~\V88(12) ;
  assign new_n212_ = ~\V120(10)  & ~\V88(10) ;
  assign new_n213_ = ~\V120(11)  & ~\V88(11) ;
  assign new_n214_ = ~\V120(13)  & ~\V88(13) ;
  assign new_n215_ = ~\V120(15)  & ~\V88(15) ;
  assign new_n216_ = ~\V120(14)  & ~\V88(14) ;
  assign new_n217_ = ~\V120(16)  & ~\V88(16) ;
  assign new_n218_ = ~\V120(17)  & ~\V88(17) ;
  assign new_n219_ = ~new_n203_ & ~new_n204_;
  assign new_n220_ = ~new_n205_ & new_n219_;
  assign new_n221_ = ~new_n206_ & new_n220_;
  assign new_n222_ = ~new_n207_ & new_n221_;
  assign new_n223_ = ~new_n208_ & new_n222_;
  assign new_n224_ = ~new_n209_ & new_n223_;
  assign new_n225_ = ~new_n210_ & new_n224_;
  assign new_n226_ = ~new_n211_ & new_n225_;
  assign new_n227_ = ~new_n212_ & new_n226_;
  assign new_n228_ = ~new_n213_ & new_n227_;
  assign new_n229_ = ~new_n214_ & new_n228_;
  assign new_n230_ = ~new_n215_ & new_n229_;
  assign new_n231_ = ~new_n216_ & new_n230_;
  assign new_n232_ = ~new_n217_ & new_n231_;
  assign \V138(2)  = ~new_n218_ & new_n232_;
  assign new_n234_ = ~\V132(5)  & ~\V126(5) ;
  assign new_n235_ = ~\V132(4)  & ~\V126(4) ;
  assign new_n236_ = ~\V132(2)  & ~\V126(2) ;
  assign new_n237_ = ~\V132(3)  & ~\V126(3) ;
  assign new_n238_ = ~\V120(25)  & ~\V88(25) ;
  assign new_n239_ = ~\V120(24)  & ~\V88(24) ;
  assign new_n240_ = ~\V120(22)  & ~\V88(22) ;
  assign new_n241_ = ~\V120(23)  & ~\V88(23) ;
  assign new_n242_ = ~\V120(28)  & ~\V88(28) ;
  assign new_n243_ = ~\V120(26)  & ~\V88(26) ;
  assign new_n244_ = ~\V120(27)  & ~\V88(27) ;
  assign new_n245_ = ~\V120(29)  & ~\V88(29) ;
  assign new_n246_ = ~\V120(31)  & ~\V88(31) ;
  assign new_n247_ = ~\V120(30)  & ~\V88(30) ;
  assign new_n248_ = ~\V132(0)  & ~\V126(0) ;
  assign new_n249_ = ~\V132(1)  & ~\V126(1) ;
  assign new_n250_ = ~new_n234_ & ~new_n235_;
  assign new_n251_ = ~new_n236_ & new_n250_;
  assign new_n252_ = ~new_n237_ & new_n251_;
  assign new_n253_ = ~new_n238_ & new_n252_;
  assign new_n254_ = ~new_n239_ & new_n253_;
  assign new_n255_ = ~new_n240_ & new_n254_;
  assign new_n256_ = ~new_n241_ & new_n255_;
  assign new_n257_ = ~new_n242_ & new_n256_;
  assign new_n258_ = ~new_n243_ & new_n257_;
  assign new_n259_ = ~new_n244_ & new_n258_;
  assign new_n260_ = ~new_n245_ & new_n259_;
  assign new_n261_ = ~new_n246_ & new_n260_;
  assign new_n262_ = ~new_n247_ & new_n261_;
  assign new_n263_ = ~new_n248_ & new_n262_;
  assign \V138(3)  = ~new_n249_ & new_n263_;
endmodule


