// Benchmark "log2" written by ABC on Tue Sep  5 18:07:10 2023

module log2 ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] ;
  wire new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_,
    new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_,
    new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_,
    new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_,
    new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_,
    new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_,
    new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_,
    new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_,
    new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_,
    new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_,
    new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_,
    new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_,
    new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_,
    new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_,
    new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_,
    new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_,
    new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_,
    new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_,
    new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_,
    new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_,
    new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_,
    new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_,
    new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_,
    new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_,
    new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_,
    new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_,
    new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_,
    new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_,
    new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_,
    new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_,
    new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_,
    new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_,
    new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_,
    new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_,
    new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_,
    new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_,
    new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_,
    new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_,
    new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_,
    new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_,
    new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_,
    new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_,
    new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_,
    new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_,
    new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_,
    new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_,
    new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_,
    new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_,
    new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_,
    new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_,
    new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_,
    new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_,
    new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_,
    new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_,
    new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_,
    new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_,
    new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_,
    new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_,
    new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_,
    new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_,
    new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_,
    new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_,
    new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_,
    new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_,
    new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_,
    new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_, new_n4509_,
    new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_,
    new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_,
    new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_,
    new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_,
    new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_,
    new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_,
    new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_,
    new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_,
    new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_,
    new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_,
    new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_,
    new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_,
    new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_,
    new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_,
    new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_,
    new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_,
    new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_,
    new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_,
    new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_,
    new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_,
    new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_,
    new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_,
    new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_,
    new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_,
    new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_,
    new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_,
    new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_,
    new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_,
    new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_,
    new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_,
    new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_,
    new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_,
    new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_,
    new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_,
    new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_,
    new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_,
    new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_,
    new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_,
    new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_,
    new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_,
    new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_,
    new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_,
    new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_,
    new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_,
    new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_,
    new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_,
    new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_,
    new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_,
    new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_,
    new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_,
    new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_,
    new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_,
    new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_,
    new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_,
    new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_,
    new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_,
    new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_,
    new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_,
    new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_,
    new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_,
    new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_,
    new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_,
    new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_,
    new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_,
    new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_,
    new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_,
    new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_,
    new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_,
    new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_,
    new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_,
    new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_,
    new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_,
    new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_,
    new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_,
    new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_,
    new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_,
    new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_,
    new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_,
    new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_,
    new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_,
    new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_,
    new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_,
    new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_,
    new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_,
    new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_,
    new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_,
    new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_,
    new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_,
    new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_,
    new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_,
    new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_,
    new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_,
    new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_,
    new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_,
    new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_,
    new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_,
    new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_,
    new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_,
    new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_,
    new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_,
    new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_,
    new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_,
    new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_,
    new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_,
    new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_,
    new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_,
    new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_,
    new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_,
    new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_,
    new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_,
    new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_,
    new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_,
    new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_,
    new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_,
    new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_,
    new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_,
    new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_,
    new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_,
    new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_,
    new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_,
    new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_,
    new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_,
    new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_,
    new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_,
    new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_,
    new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_,
    new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_,
    new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_,
    new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_,
    new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_,
    new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_,
    new_n6316_, new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_,
    new_n6322_, new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_,
    new_n6328_, new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_,
    new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_,
    new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_,
    new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_,
    new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_,
    new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_,
    new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_,
    new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_,
    new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_,
    new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_,
    new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_,
    new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_,
    new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_,
    new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_,
    new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_,
    new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_,
    new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_,
    new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_,
    new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_,
    new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_,
    new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_,
    new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_,
    new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_,
    new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_,
    new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_,
    new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_,
    new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_,
    new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_,
    new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_,
    new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_,
    new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_,
    new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_,
    new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_,
    new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_,
    new_n6574_, new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_,
    new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_,
    new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_,
    new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_,
    new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_,
    new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_,
    new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_,
    new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_,
    new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_,
    new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_,
    new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_,
    new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_,
    new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_,
    new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_,
    new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_,
    new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_,
    new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_,
    new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_,
    new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_,
    new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_,
    new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_,
    new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_,
    new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_,
    new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_, new_n6735_,
    new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_, new_n6741_,
    new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_,
    new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_,
    new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_,
    new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_,
    new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_,
    new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_,
    new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_,
    new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_,
    new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_,
    new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_,
    new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_,
    new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_,
    new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_,
    new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_,
    new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_,
    new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_,
    new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_,
    new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_,
    new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_,
    new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6867_,
    new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_,
    new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_,
    new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_,
    new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_,
    new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_,
    new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_,
    new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_,
    new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_,
    new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_,
    new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_,
    new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_,
    new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_,
    new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_,
    new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_, new_n6951_,
    new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_,
    new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_,
    new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_,
    new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_,
    new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_,
    new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_,
    new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_,
    new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_,
    new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_,
    new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_,
    new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_,
    new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_,
    new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_,
    new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_,
    new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_,
    new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_,
    new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_,
    new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_,
    new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_,
    new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_,
    new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_,
    new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_,
    new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_,
    new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_,
    new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_,
    new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_,
    new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_,
    new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_,
    new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_,
    new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7131_,
    new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_,
    new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_,
    new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_,
    new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_,
    new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_,
    new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_, new_n7167_,
    new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_, new_n7173_,
    new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_,
    new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_,
    new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_,
    new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_,
    new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_,
    new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_,
    new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_,
    new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_,
    new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_,
    new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_,
    new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_,
    new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_,
    new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_,
    new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_,
    new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_,
    new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_,
    new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_,
    new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_,
    new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_,
    new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_,
    new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_,
    new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_,
    new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_,
    new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_,
    new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_,
    new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_,
    new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_,
    new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_,
    new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_,
    new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_,
    new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_,
    new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_,
    new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_,
    new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_,
    new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_,
    new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_,
    new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_,
    new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_,
    new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_,
    new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_,
    new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_,
    new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_,
    new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_,
    new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_,
    new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_,
    new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_,
    new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_,
    new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_,
    new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_,
    new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_,
    new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_,
    new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_,
    new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_,
    new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_,
    new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_,
    new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_,
    new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_,
    new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_,
    new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_,
    new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_,
    new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_,
    new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_,
    new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_,
    new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_,
    new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_,
    new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_,
    new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_,
    new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_,
    new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_,
    new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_,
    new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_,
    new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_,
    new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_,
    new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_,
    new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_,
    new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_,
    new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_,
    new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_,
    new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_,
    new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_,
    new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_,
    new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_,
    new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_,
    new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_,
    new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_,
    new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_,
    new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_,
    new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_,
    new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_,
    new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_,
    new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_,
    new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_,
    new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_,
    new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_,
    new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_,
    new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_,
    new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_,
    new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_,
    new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_,
    new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_,
    new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_,
    new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_,
    new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_,
    new_n8398_, new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_,
    new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_,
    new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_,
    new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_,
    new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_,
    new_n8428_, new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_,
    new_n8434_, new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_,
    new_n8440_, new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_,
    new_n8446_, new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_,
    new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_,
    new_n8458_, new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_,
    new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_,
    new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_,
    new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_,
    new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_,
    new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_,
    new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_,
    new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_,
    new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_,
    new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_,
    new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_,
    new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_,
    new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_,
    new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_,
    new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_,
    new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_,
    new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_,
    new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_,
    new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_,
    new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_,
    new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_,
    new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_,
    new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_,
    new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_,
    new_n8632_, new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_,
    new_n8638_, new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_,
    new_n8644_, new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_,
    new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_,
    new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_,
    new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_,
    new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_,
    new_n8674_, new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_,
    new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_,
    new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_,
    new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_,
    new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_,
    new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_,
    new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_,
    new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_,
    new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_,
    new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_,
    new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_,
    new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_,
    new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_,
    new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_,
    new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_,
    new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_,
    new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_,
    new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_,
    new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8824_, new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_,
    new_n8830_, new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_,
    new_n8860_, new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_,
    new_n8866_, new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_,
    new_n8872_, new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_,
    new_n8878_, new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_,
    new_n8884_, new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_,
    new_n8890_, new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_,
    new_n8896_, new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_,
    new_n8902_, new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_,
    new_n8908_, new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_,
    new_n8914_, new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_,
    new_n8920_, new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_,
    new_n8926_, new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_,
    new_n8932_, new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_,
    new_n8938_, new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_,
    new_n8944_, new_n8945_, new_n8946_, new_n8947_, new_n8948_, new_n8949_,
    new_n8950_, new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_,
    new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_,
    new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_,
    new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_,
    new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_,
    new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_,
    new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_,
    new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_,
    new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_,
    new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_,
    new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_,
    new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_,
    new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_,
    new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_,
    new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_,
    new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_,
    new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_,
    new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_,
    new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_,
    new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_,
    new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_,
    new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_,
    new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_,
    new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_,
    new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_,
    new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_,
    new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_,
    new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_,
    new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_,
    new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_,
    new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_,
    new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_,
    new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_,
    new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_,
    new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_,
    new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_,
    new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_,
    new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_,
    new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_,
    new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_,
    new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_,
    new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_,
    new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_,
    new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_,
    new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_,
    new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_,
    new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_,
    new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_,
    new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_,
    new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_,
    new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_,
    new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_,
    new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_,
    new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_,
    new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_,
    new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_,
    new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_,
    new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_,
    new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_,
    new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_,
    new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_,
    new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_,
    new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_,
    new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_,
    new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_,
    new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_,
    new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_,
    new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_,
    new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_,
    new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_,
    new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_,
    new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_,
    new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_,
    new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_,
    new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_,
    new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_,
    new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_,
    new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_,
    new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_,
    new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10439_,
    new_n10440_, new_n10441_, new_n10442_, new_n10443_, new_n10444_,
    new_n10445_, new_n10446_, new_n10447_, new_n10448_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10453_, new_n10454_,
    new_n10455_, new_n10456_, new_n10457_, new_n10458_, new_n10459_,
    new_n10460_, new_n10461_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10868_, new_n10869_,
    new_n10870_, new_n10871_, new_n10872_, new_n10873_, new_n10874_,
    new_n10875_, new_n10876_, new_n10877_, new_n10878_, new_n10879_,
    new_n10880_, new_n10881_, new_n10882_, new_n10883_, new_n10884_,
    new_n10885_, new_n10886_, new_n10887_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10894_,
    new_n10895_, new_n10896_, new_n10897_, new_n10898_, new_n10899_,
    new_n10900_, new_n10901_, new_n10902_, new_n10903_, new_n10904_,
    new_n10905_, new_n10906_, new_n10907_, new_n10908_, new_n10909_,
    new_n10910_, new_n10911_, new_n10912_, new_n10913_, new_n10914_,
    new_n10915_, new_n10916_, new_n10917_, new_n10918_, new_n10919_,
    new_n10920_, new_n10921_, new_n10922_, new_n10923_, new_n10924_,
    new_n10925_, new_n10926_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10933_, new_n10934_,
    new_n10935_, new_n10936_, new_n10937_, new_n10938_, new_n10939_,
    new_n10940_, new_n10941_, new_n10942_, new_n10943_, new_n10944_,
    new_n10945_, new_n10946_, new_n10947_, new_n10948_, new_n10949_,
    new_n10950_, new_n10951_, new_n10952_, new_n10953_, new_n10954_,
    new_n10955_, new_n10956_, new_n10957_, new_n10958_, new_n10959_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10974_,
    new_n10975_, new_n10976_, new_n10977_, new_n10978_, new_n10979_,
    new_n10980_, new_n10981_, new_n10982_, new_n10983_, new_n10984_,
    new_n10985_, new_n10986_, new_n10987_, new_n10988_, new_n10989_,
    new_n10990_, new_n10991_, new_n10992_, new_n10993_, new_n10994_,
    new_n10995_, new_n10996_, new_n10997_, new_n10998_, new_n10999_,
    new_n11000_, new_n11001_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11050_, new_n11051_, new_n11052_, new_n11053_, new_n11054_,
    new_n11055_, new_n11056_, new_n11057_, new_n11058_, new_n11059_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11073_, new_n11074_,
    new_n11075_, new_n11076_, new_n11077_, new_n11078_, new_n11079_,
    new_n11080_, new_n11081_, new_n11082_, new_n11083_, new_n11084_,
    new_n11085_, new_n11086_, new_n11087_, new_n11088_, new_n11089_,
    new_n11090_, new_n11091_, new_n11092_, new_n11093_, new_n11094_,
    new_n11095_, new_n11096_, new_n11097_, new_n11098_, new_n11099_,
    new_n11100_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11106_, new_n11107_, new_n11108_, new_n11109_,
    new_n11110_, new_n11111_, new_n11112_, new_n11113_, new_n11114_,
    new_n11115_, new_n11116_, new_n11117_, new_n11118_, new_n11119_,
    new_n11120_, new_n11121_, new_n11122_, new_n11123_, new_n11124_,
    new_n11125_, new_n11126_, new_n11127_, new_n11128_, new_n11129_,
    new_n11130_, new_n11131_, new_n11132_, new_n11133_, new_n11134_,
    new_n11135_, new_n11136_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11146_, new_n11147_, new_n11148_, new_n11149_,
    new_n11150_, new_n11151_, new_n11152_, new_n11153_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11166_, new_n11167_, new_n11168_, new_n11169_,
    new_n11170_, new_n11171_, new_n11172_, new_n11173_, new_n11174_,
    new_n11175_, new_n11176_, new_n11177_, new_n11178_, new_n11179_,
    new_n11180_, new_n11181_, new_n11182_, new_n11183_, new_n11184_,
    new_n11185_, new_n11186_, new_n11187_, new_n11188_, new_n11189_,
    new_n11190_, new_n11191_, new_n11192_, new_n11193_, new_n11194_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11260_, new_n11261_, new_n11262_, new_n11263_, new_n11264_,
    new_n11265_, new_n11266_, new_n11267_, new_n11268_, new_n11269_,
    new_n11270_, new_n11271_, new_n11272_, new_n11273_, new_n11274_,
    new_n11275_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11286_, new_n11287_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11298_, new_n11299_,
    new_n11300_, new_n11301_, new_n11302_, new_n11303_, new_n11304_,
    new_n11305_, new_n11306_, new_n11307_, new_n11308_, new_n11309_,
    new_n11310_, new_n11311_, new_n11312_, new_n11313_, new_n11314_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11324_,
    new_n11325_, new_n11326_, new_n11327_, new_n11328_, new_n11329_,
    new_n11330_, new_n11331_, new_n11332_, new_n11333_, new_n11334_,
    new_n11335_, new_n11336_, new_n11337_, new_n11338_, new_n11339_,
    new_n11340_, new_n11341_, new_n11342_, new_n11343_, new_n11344_,
    new_n11345_, new_n11346_, new_n11347_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11352_, new_n11353_, new_n11354_,
    new_n11355_, new_n11356_, new_n11357_, new_n11358_, new_n11359_,
    new_n11360_, new_n11361_, new_n11362_, new_n11363_, new_n11364_,
    new_n11365_, new_n11366_, new_n11367_, new_n11368_, new_n11369_,
    new_n11370_, new_n11371_, new_n11372_, new_n11373_, new_n11374_,
    new_n11375_, new_n11376_, new_n11377_, new_n11378_, new_n11379_,
    new_n11380_, new_n11381_, new_n11382_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11528_, new_n11529_,
    new_n11530_, new_n11531_, new_n11532_, new_n11533_, new_n11534_,
    new_n11535_, new_n11536_, new_n11537_, new_n11538_, new_n11539_,
    new_n11540_, new_n11541_, new_n11542_, new_n11543_, new_n11544_,
    new_n11545_, new_n11546_, new_n11547_, new_n11548_, new_n11549_,
    new_n11550_, new_n11551_, new_n11552_, new_n11553_, new_n11554_,
    new_n11555_, new_n11556_, new_n11557_, new_n11558_, new_n11559_,
    new_n11560_, new_n11561_, new_n11562_, new_n11563_, new_n11564_,
    new_n11565_, new_n11566_, new_n11567_, new_n11568_, new_n11569_,
    new_n11570_, new_n11571_, new_n11572_, new_n11573_, new_n11574_,
    new_n11575_, new_n11576_, new_n11577_, new_n11578_, new_n11579_,
    new_n11580_, new_n11581_, new_n11582_, new_n11583_, new_n11584_,
    new_n11585_, new_n11586_, new_n11587_, new_n11588_, new_n11589_,
    new_n11590_, new_n11591_, new_n11592_, new_n11593_, new_n11594_,
    new_n11595_, new_n11596_, new_n11597_, new_n11598_, new_n11599_,
    new_n11600_, new_n11601_, new_n11602_, new_n11603_, new_n11604_,
    new_n11605_, new_n11606_, new_n11607_, new_n11608_, new_n11609_,
    new_n11610_, new_n11611_, new_n11612_, new_n11613_, new_n11614_,
    new_n11615_, new_n11616_, new_n11617_, new_n11618_, new_n11619_,
    new_n11620_, new_n11621_, new_n11622_, new_n11623_, new_n11624_,
    new_n11625_, new_n11626_, new_n11627_, new_n11628_, new_n11629_,
    new_n11630_, new_n11631_, new_n11632_, new_n11633_, new_n11634_,
    new_n11635_, new_n11636_, new_n11637_, new_n11638_, new_n11639_,
    new_n11640_, new_n11641_, new_n11642_, new_n11643_, new_n11644_,
    new_n11645_, new_n11646_, new_n11647_, new_n11648_, new_n11649_,
    new_n11650_, new_n11651_, new_n11652_, new_n11653_, new_n11654_,
    new_n11655_, new_n11656_, new_n11657_, new_n11658_, new_n11659_,
    new_n11660_, new_n11661_, new_n11662_, new_n11663_, new_n11664_,
    new_n11665_, new_n11666_, new_n11667_, new_n11668_, new_n11669_,
    new_n11670_, new_n11671_, new_n11672_, new_n11673_, new_n11674_,
    new_n11675_, new_n11676_, new_n11677_, new_n11678_, new_n11679_,
    new_n11680_, new_n11681_, new_n11682_, new_n11683_, new_n11684_,
    new_n11685_, new_n11686_, new_n11687_, new_n11688_, new_n11689_,
    new_n11690_, new_n11691_, new_n11692_, new_n11693_, new_n11694_,
    new_n11695_, new_n11696_, new_n11697_, new_n11698_, new_n11699_,
    new_n11700_, new_n11701_, new_n11702_, new_n11703_, new_n11704_,
    new_n11705_, new_n11706_, new_n11707_, new_n11708_, new_n11709_,
    new_n11710_, new_n11711_, new_n11712_, new_n11713_, new_n11714_,
    new_n11715_, new_n11716_, new_n11717_, new_n11718_, new_n11719_,
    new_n11720_, new_n11721_, new_n11722_, new_n11723_, new_n11724_,
    new_n11725_, new_n11726_, new_n11727_, new_n11728_, new_n11729_,
    new_n11730_, new_n11731_, new_n11732_, new_n11733_, new_n11734_,
    new_n11735_, new_n11736_, new_n11737_, new_n11738_, new_n11739_,
    new_n11740_, new_n11741_, new_n11742_, new_n11743_, new_n11744_,
    new_n11745_, new_n11746_, new_n11747_, new_n11748_, new_n11749_,
    new_n11750_, new_n11751_, new_n11752_, new_n11753_, new_n11754_,
    new_n11755_, new_n11756_, new_n11757_, new_n11758_, new_n11759_,
    new_n11760_, new_n11761_, new_n11762_, new_n11763_, new_n11764_,
    new_n11765_, new_n11766_, new_n11767_, new_n11768_, new_n11769_,
    new_n11770_, new_n11771_, new_n11772_, new_n11773_, new_n11774_,
    new_n11775_, new_n11776_, new_n11777_, new_n11778_, new_n11779_,
    new_n11780_, new_n11781_, new_n11782_, new_n11783_, new_n11784_,
    new_n11785_, new_n11786_, new_n11787_, new_n11788_, new_n11789_,
    new_n11790_, new_n11791_, new_n11792_, new_n11793_, new_n11794_,
    new_n11795_, new_n11796_, new_n11797_, new_n11798_, new_n11799_,
    new_n11800_, new_n11801_, new_n11802_, new_n11803_, new_n11804_,
    new_n11805_, new_n11806_, new_n11807_, new_n11808_, new_n11809_,
    new_n11810_, new_n11811_, new_n11812_, new_n11813_, new_n11814_,
    new_n11815_, new_n11816_, new_n11817_, new_n11818_, new_n11819_,
    new_n11820_, new_n11821_, new_n11822_, new_n11823_, new_n11824_,
    new_n11825_, new_n11826_, new_n11827_, new_n11828_, new_n11829_,
    new_n11830_, new_n11831_, new_n11832_, new_n11833_, new_n11834_,
    new_n11835_, new_n11836_, new_n11837_, new_n11838_, new_n11839_,
    new_n11840_, new_n11841_, new_n11842_, new_n11843_, new_n11844_,
    new_n11845_, new_n11846_, new_n11847_, new_n11848_, new_n11849_,
    new_n11850_, new_n11851_, new_n11852_, new_n11853_, new_n11854_,
    new_n11855_, new_n11856_, new_n11857_, new_n11858_, new_n11859_,
    new_n11860_, new_n11861_, new_n11862_, new_n11863_, new_n11864_,
    new_n11865_, new_n11866_, new_n11867_, new_n11868_, new_n11869_,
    new_n11870_, new_n11871_, new_n11872_, new_n11873_, new_n11874_,
    new_n11875_, new_n11876_, new_n11877_, new_n11878_, new_n11879_,
    new_n11880_, new_n11881_, new_n11882_, new_n11883_, new_n11884_,
    new_n11885_, new_n11886_, new_n11887_, new_n11888_, new_n11889_,
    new_n11890_, new_n11891_, new_n11892_, new_n11893_, new_n11894_,
    new_n11895_, new_n11896_, new_n11897_, new_n11898_, new_n11899_,
    new_n11900_, new_n11901_, new_n11902_, new_n11903_, new_n11904_,
    new_n11905_, new_n11906_, new_n11907_, new_n11908_, new_n11909_,
    new_n11910_, new_n11911_, new_n11912_, new_n11913_, new_n11914_,
    new_n11915_, new_n11916_, new_n11917_, new_n11918_, new_n11919_,
    new_n11920_, new_n11921_, new_n11922_, new_n11923_, new_n11924_,
    new_n11925_, new_n11926_, new_n11927_, new_n11928_, new_n11929_,
    new_n11930_, new_n11931_, new_n11932_, new_n11933_, new_n11934_,
    new_n11935_, new_n11936_, new_n11937_, new_n11938_, new_n11939_,
    new_n11940_, new_n11941_, new_n11942_, new_n11943_, new_n11944_,
    new_n11945_, new_n11946_, new_n11947_, new_n11948_, new_n11949_,
    new_n11950_, new_n11951_, new_n11952_, new_n11953_, new_n11954_,
    new_n11955_, new_n11956_, new_n11957_, new_n11958_, new_n11959_,
    new_n11960_, new_n11961_, new_n11962_, new_n11963_, new_n11964_,
    new_n11965_, new_n11966_, new_n11967_, new_n11968_, new_n11969_,
    new_n11970_, new_n11971_, new_n11972_, new_n11973_, new_n11974_,
    new_n11975_, new_n11976_, new_n11977_, new_n11978_, new_n11979_,
    new_n11980_, new_n11981_, new_n11982_, new_n11983_, new_n11984_,
    new_n11985_, new_n11986_, new_n11987_, new_n11988_, new_n11989_,
    new_n11990_, new_n11991_, new_n11992_, new_n11993_, new_n11994_,
    new_n11995_, new_n11996_, new_n11997_, new_n11998_, new_n11999_,
    new_n12000_, new_n12001_, new_n12002_, new_n12003_, new_n12004_,
    new_n12005_, new_n12006_, new_n12007_, new_n12008_, new_n12009_,
    new_n12010_, new_n12011_, new_n12012_, new_n12013_, new_n12014_,
    new_n12015_, new_n12016_, new_n12017_, new_n12018_, new_n12019_,
    new_n12020_, new_n12021_, new_n12022_, new_n12023_, new_n12024_,
    new_n12025_, new_n12026_, new_n12027_, new_n12028_, new_n12029_,
    new_n12030_, new_n12031_, new_n12032_, new_n12033_, new_n12034_,
    new_n12035_, new_n12036_, new_n12037_, new_n12038_, new_n12039_,
    new_n12040_, new_n12041_, new_n12042_, new_n12043_, new_n12044_,
    new_n12045_, new_n12046_, new_n12047_, new_n12048_, new_n12049_,
    new_n12050_, new_n12051_, new_n12052_, new_n12053_, new_n12054_,
    new_n12055_, new_n12056_, new_n12057_, new_n12058_, new_n12059_,
    new_n12060_, new_n12061_, new_n12062_, new_n12063_, new_n12064_,
    new_n12065_, new_n12066_, new_n12067_, new_n12068_, new_n12069_,
    new_n12070_, new_n12071_, new_n12072_, new_n12073_, new_n12074_,
    new_n12075_, new_n12076_, new_n12077_, new_n12078_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12084_,
    new_n12085_, new_n12086_, new_n12087_, new_n12088_, new_n12089_,
    new_n12090_, new_n12091_, new_n12092_, new_n12093_, new_n12094_,
    new_n12095_, new_n12096_, new_n12097_, new_n12098_, new_n12099_,
    new_n12100_, new_n12101_, new_n12102_, new_n12103_, new_n12104_,
    new_n12105_, new_n12106_, new_n12107_, new_n12108_, new_n12109_,
    new_n12110_, new_n12111_, new_n12112_, new_n12113_, new_n12114_,
    new_n12115_, new_n12116_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12214_,
    new_n12215_, new_n12216_, new_n12217_, new_n12218_, new_n12219_,
    new_n12220_, new_n12221_, new_n12222_, new_n12223_, new_n12224_,
    new_n12225_, new_n12226_, new_n12227_, new_n12228_, new_n12229_,
    new_n12230_, new_n12231_, new_n12232_, new_n12233_, new_n12234_,
    new_n12235_, new_n12236_, new_n12237_, new_n12238_, new_n12239_,
    new_n12240_, new_n12241_, new_n12242_, new_n12243_, new_n12244_,
    new_n12245_, new_n12246_, new_n12247_, new_n12248_, new_n12249_,
    new_n12250_, new_n12251_, new_n12252_, new_n12253_, new_n12254_,
    new_n12255_, new_n12256_, new_n12257_, new_n12258_, new_n12259_,
    new_n12260_, new_n12261_, new_n12262_, new_n12263_, new_n12264_,
    new_n12265_, new_n12266_, new_n12267_, new_n12268_, new_n12269_,
    new_n12270_, new_n12271_, new_n12272_, new_n12273_, new_n12274_,
    new_n12275_, new_n12276_, new_n12277_, new_n12278_, new_n12279_,
    new_n12280_, new_n12281_, new_n12282_, new_n12283_, new_n12284_,
    new_n12285_, new_n12286_, new_n12287_, new_n12288_, new_n12289_,
    new_n12290_, new_n12291_, new_n12292_, new_n12293_, new_n12294_,
    new_n12295_, new_n12296_, new_n12297_, new_n12298_, new_n12299_,
    new_n12300_, new_n12301_, new_n12302_, new_n12303_, new_n12304_,
    new_n12305_, new_n12306_, new_n12307_, new_n12308_, new_n12309_,
    new_n12310_, new_n12311_, new_n12312_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12561_, new_n12562_, new_n12563_, new_n12564_,
    new_n12565_, new_n12566_, new_n12567_, new_n12568_, new_n12569_,
    new_n12570_, new_n12571_, new_n12572_, new_n12573_, new_n12574_,
    new_n12575_, new_n12576_, new_n12577_, new_n12578_, new_n12579_,
    new_n12580_, new_n12581_, new_n12582_, new_n12583_, new_n12584_,
    new_n12585_, new_n12586_, new_n12587_, new_n12588_, new_n12589_,
    new_n12590_, new_n12591_, new_n12592_, new_n12593_, new_n12594_,
    new_n12595_, new_n12596_, new_n12597_, new_n12598_, new_n12599_,
    new_n12600_, new_n12601_, new_n12602_, new_n12603_, new_n12604_,
    new_n12605_, new_n12606_, new_n12607_, new_n12608_, new_n12609_,
    new_n12610_, new_n12611_, new_n12612_, new_n12613_, new_n12614_,
    new_n12615_, new_n12616_, new_n12617_, new_n12618_, new_n12619_,
    new_n12620_, new_n12621_, new_n12622_, new_n12623_, new_n12624_,
    new_n12625_, new_n12626_, new_n12627_, new_n12628_, new_n12629_,
    new_n12630_, new_n12631_, new_n12632_, new_n12633_, new_n12634_,
    new_n12635_, new_n12636_, new_n12637_, new_n12638_, new_n12639_,
    new_n12640_, new_n12641_, new_n12642_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12649_,
    new_n12650_, new_n12651_, new_n12652_, new_n12653_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12663_, new_n12664_,
    new_n12665_, new_n12666_, new_n12667_, new_n12668_, new_n12669_,
    new_n12670_, new_n12671_, new_n12672_, new_n12673_, new_n12674_,
    new_n12675_, new_n12676_, new_n12677_, new_n12678_, new_n12679_,
    new_n12680_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12687_, new_n12688_, new_n12689_,
    new_n12690_, new_n12691_, new_n12692_, new_n12693_, new_n12694_,
    new_n12695_, new_n12696_, new_n12697_, new_n12698_, new_n12699_,
    new_n12700_, new_n12701_, new_n12702_, new_n12703_, new_n12704_,
    new_n12705_, new_n12706_, new_n12707_, new_n12708_, new_n12709_,
    new_n12710_, new_n12711_, new_n12712_, new_n12713_, new_n12714_,
    new_n12715_, new_n12716_, new_n12717_, new_n12718_, new_n12719_,
    new_n12720_, new_n12721_, new_n12722_, new_n12723_, new_n12724_,
    new_n12725_, new_n12726_, new_n12727_, new_n12728_, new_n12729_,
    new_n12730_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13089_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13096_, new_n13097_, new_n13098_, new_n13099_,
    new_n13100_, new_n13101_, new_n13102_, new_n13103_, new_n13104_,
    new_n13105_, new_n13106_, new_n13107_, new_n13108_, new_n13109_,
    new_n13110_, new_n13111_, new_n13112_, new_n13113_, new_n13114_,
    new_n13115_, new_n13116_, new_n13117_, new_n13118_, new_n13119_,
    new_n13120_, new_n13121_, new_n13122_, new_n13123_, new_n13124_,
    new_n13125_, new_n13126_, new_n13127_, new_n13128_, new_n13129_,
    new_n13130_, new_n13131_, new_n13132_, new_n13133_, new_n13134_,
    new_n13135_, new_n13136_, new_n13137_, new_n13138_, new_n13139_,
    new_n13140_, new_n13141_, new_n13142_, new_n13143_, new_n13144_,
    new_n13145_, new_n13146_, new_n13147_, new_n13148_, new_n13149_,
    new_n13150_, new_n13151_, new_n13152_, new_n13153_, new_n13154_,
    new_n13155_, new_n13156_, new_n13157_, new_n13158_, new_n13159_,
    new_n13160_, new_n13161_, new_n13162_, new_n13163_, new_n13164_,
    new_n13165_, new_n13166_, new_n13167_, new_n13168_, new_n13169_,
    new_n13170_, new_n13171_, new_n13172_, new_n13173_, new_n13174_,
    new_n13175_, new_n13176_, new_n13177_, new_n13178_, new_n13179_,
    new_n13180_, new_n13181_, new_n13182_, new_n13183_, new_n13184_,
    new_n13185_, new_n13186_, new_n13187_, new_n13188_, new_n13189_,
    new_n13190_, new_n13191_, new_n13192_, new_n13193_, new_n13194_,
    new_n13195_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13200_, new_n13201_, new_n13202_, new_n13203_, new_n13204_,
    new_n13205_, new_n13206_, new_n13207_, new_n13208_, new_n13209_,
    new_n13210_, new_n13211_, new_n13212_, new_n13213_, new_n13214_,
    new_n13215_, new_n13216_, new_n13217_, new_n13218_, new_n13219_,
    new_n13220_, new_n13221_, new_n13222_, new_n13223_, new_n13224_,
    new_n13225_, new_n13226_, new_n13227_, new_n13228_, new_n13229_,
    new_n13230_, new_n13231_, new_n13232_, new_n13233_, new_n13234_,
    new_n13235_, new_n13236_, new_n13237_, new_n13238_, new_n13239_,
    new_n13240_, new_n13241_, new_n13242_, new_n13243_, new_n13244_,
    new_n13245_, new_n13246_, new_n13247_, new_n13248_, new_n13249_,
    new_n13250_, new_n13251_, new_n13252_, new_n13253_, new_n13254_,
    new_n13255_, new_n13256_, new_n13257_, new_n13258_, new_n13259_,
    new_n13260_, new_n13261_, new_n13262_, new_n13263_, new_n13264_,
    new_n13265_, new_n13266_, new_n13267_, new_n13268_, new_n13269_,
    new_n13270_, new_n13271_, new_n13272_, new_n13273_, new_n13274_,
    new_n13275_, new_n13276_, new_n13277_, new_n13278_, new_n13279_,
    new_n13280_, new_n13281_, new_n13282_, new_n13283_, new_n13284_,
    new_n13285_, new_n13286_, new_n13287_, new_n13288_, new_n13289_,
    new_n13290_, new_n13291_, new_n13292_, new_n13293_, new_n13294_,
    new_n13295_, new_n13296_, new_n13297_, new_n13298_, new_n13299_,
    new_n13300_, new_n13301_, new_n13302_, new_n13303_, new_n13304_,
    new_n13305_, new_n13306_, new_n13307_, new_n13308_, new_n13309_,
    new_n13310_, new_n13311_, new_n13312_, new_n13313_, new_n13314_,
    new_n13315_, new_n13316_, new_n13317_, new_n13318_, new_n13319_,
    new_n13320_, new_n13321_, new_n13322_, new_n13323_, new_n13324_,
    new_n13325_, new_n13326_, new_n13327_, new_n13328_, new_n13329_,
    new_n13330_, new_n13331_, new_n13332_, new_n13333_, new_n13334_,
    new_n13335_, new_n13336_, new_n13337_, new_n13338_, new_n13339_,
    new_n13340_, new_n13341_, new_n13342_, new_n13343_, new_n13344_,
    new_n13345_, new_n13346_, new_n13347_, new_n13348_, new_n13349_,
    new_n13350_, new_n13351_, new_n13352_, new_n13353_, new_n13354_,
    new_n13355_, new_n13356_, new_n13357_, new_n13358_, new_n13359_,
    new_n13360_, new_n13361_, new_n13362_, new_n13363_, new_n13364_,
    new_n13365_, new_n13366_, new_n13367_, new_n13368_, new_n13369_,
    new_n13370_, new_n13371_, new_n13372_, new_n13373_, new_n13374_,
    new_n13375_, new_n13376_, new_n13377_, new_n13378_, new_n13379_,
    new_n13380_, new_n13381_, new_n13382_, new_n13383_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13396_, new_n13397_, new_n13398_, new_n13399_,
    new_n13400_, new_n13401_, new_n13402_, new_n13403_, new_n13404_,
    new_n13405_, new_n13406_, new_n13407_, new_n13408_, new_n13409_,
    new_n13410_, new_n13411_, new_n13412_, new_n13413_, new_n13414_,
    new_n13415_, new_n13416_, new_n13417_, new_n13418_, new_n13419_,
    new_n13420_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13425_, new_n13426_, new_n13427_, new_n13428_, new_n13429_,
    new_n13430_, new_n13431_, new_n13432_, new_n13433_, new_n13434_,
    new_n13435_, new_n13436_, new_n13437_, new_n13438_, new_n13439_,
    new_n13440_, new_n13441_, new_n13442_, new_n13443_, new_n13444_,
    new_n13445_, new_n13446_, new_n13447_, new_n13448_, new_n13449_,
    new_n13450_, new_n13451_, new_n13452_, new_n13453_, new_n13454_,
    new_n13455_, new_n13456_, new_n13457_, new_n13458_, new_n13459_,
    new_n13460_, new_n13461_, new_n13462_, new_n13463_, new_n13464_,
    new_n13465_, new_n13466_, new_n13467_, new_n13468_, new_n13469_,
    new_n13470_, new_n13471_, new_n13472_, new_n13473_, new_n13474_,
    new_n13475_, new_n13476_, new_n13477_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13487_, new_n13488_, new_n13489_,
    new_n13490_, new_n13491_, new_n13492_, new_n13493_, new_n13494_,
    new_n13495_, new_n13496_, new_n13497_, new_n13498_, new_n13499_,
    new_n13500_, new_n13501_, new_n13502_, new_n13503_, new_n13504_,
    new_n13505_, new_n13506_, new_n13507_, new_n13508_, new_n13509_,
    new_n13510_, new_n13511_, new_n13512_, new_n13513_, new_n13514_,
    new_n13515_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13523_, new_n13524_,
    new_n13525_, new_n13526_, new_n13527_, new_n13528_, new_n13529_,
    new_n13530_, new_n13531_, new_n13532_, new_n13533_, new_n13534_,
    new_n13535_, new_n13536_, new_n13537_, new_n13538_, new_n13539_,
    new_n13540_, new_n13541_, new_n13542_, new_n13543_, new_n13544_,
    new_n13545_, new_n13546_, new_n13547_, new_n13548_, new_n13549_,
    new_n13550_, new_n13551_, new_n13552_, new_n13553_, new_n13554_,
    new_n13555_, new_n13556_, new_n13557_, new_n13558_, new_n13559_,
    new_n13560_, new_n13561_, new_n13562_, new_n13563_, new_n13564_,
    new_n13565_, new_n13566_, new_n13567_, new_n13568_, new_n13569_,
    new_n13570_, new_n13571_, new_n13572_, new_n13573_, new_n13574_,
    new_n13575_, new_n13576_, new_n13577_, new_n13578_, new_n13579_,
    new_n13580_, new_n13581_, new_n13582_, new_n13583_, new_n13584_,
    new_n13585_, new_n13586_, new_n13587_, new_n13588_, new_n13589_,
    new_n13590_, new_n13591_, new_n13592_, new_n13593_, new_n13594_,
    new_n13595_, new_n13596_, new_n13597_, new_n13598_, new_n13599_,
    new_n13600_, new_n13601_, new_n13602_, new_n13603_, new_n13604_,
    new_n13605_, new_n13606_, new_n13607_, new_n13608_, new_n13609_,
    new_n13610_, new_n13611_, new_n13612_, new_n13613_, new_n13614_,
    new_n13615_, new_n13616_, new_n13617_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13627_, new_n13628_, new_n13629_,
    new_n13630_, new_n13631_, new_n13632_, new_n13633_, new_n13634_,
    new_n13635_, new_n13636_, new_n13637_, new_n13638_, new_n13639_,
    new_n13640_, new_n13641_, new_n13642_, new_n13643_, new_n13644_,
    new_n13645_, new_n13646_, new_n13647_, new_n13648_, new_n13649_,
    new_n13650_, new_n13651_, new_n13652_, new_n13653_, new_n13654_,
    new_n13655_, new_n13656_, new_n13657_, new_n13658_, new_n13659_,
    new_n13660_, new_n13661_, new_n13662_, new_n13663_, new_n13664_,
    new_n13665_, new_n13666_, new_n13667_, new_n13668_, new_n13669_,
    new_n13670_, new_n13671_, new_n13672_, new_n13673_, new_n13674_,
    new_n13675_, new_n13676_, new_n13677_, new_n13678_, new_n13679_,
    new_n13680_, new_n13681_, new_n13682_, new_n13683_, new_n13684_,
    new_n13685_, new_n13686_, new_n13687_, new_n13688_, new_n13689_,
    new_n13690_, new_n13691_, new_n13692_, new_n13693_, new_n13694_,
    new_n13695_, new_n13696_, new_n13697_, new_n13698_, new_n13699_,
    new_n13700_, new_n13701_, new_n13702_, new_n13703_, new_n13704_,
    new_n13705_, new_n13706_, new_n13707_, new_n13708_, new_n13709_,
    new_n13710_, new_n13711_, new_n13712_, new_n13713_, new_n13714_,
    new_n13715_, new_n13716_, new_n13717_, new_n13718_, new_n13719_,
    new_n13720_, new_n13721_, new_n13722_, new_n13723_, new_n13724_,
    new_n13725_, new_n13726_, new_n13727_, new_n13728_, new_n13729_,
    new_n13730_, new_n13731_, new_n13732_, new_n13733_, new_n13734_,
    new_n13735_, new_n13736_, new_n13737_, new_n13738_, new_n13739_,
    new_n13740_, new_n13741_, new_n13742_, new_n13743_, new_n13744_,
    new_n13745_, new_n13746_, new_n13747_, new_n13748_, new_n13749_,
    new_n13750_, new_n13751_, new_n13752_, new_n13753_, new_n13754_,
    new_n13755_, new_n13756_, new_n13757_, new_n13758_, new_n13759_,
    new_n13760_, new_n13761_, new_n13762_, new_n13763_, new_n13764_,
    new_n13765_, new_n13766_, new_n13767_, new_n13768_, new_n13769_,
    new_n13770_, new_n13771_, new_n13772_, new_n13773_, new_n13774_,
    new_n13775_, new_n13776_, new_n13777_, new_n13778_, new_n13779_,
    new_n13780_, new_n13781_, new_n13782_, new_n13783_, new_n13784_,
    new_n13785_, new_n13786_, new_n13787_, new_n13788_, new_n13789_,
    new_n13790_, new_n13791_, new_n13792_, new_n13793_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13799_,
    new_n13800_, new_n13801_, new_n13802_, new_n13803_, new_n13804_,
    new_n13805_, new_n13806_, new_n13807_, new_n13808_, new_n13809_,
    new_n13810_, new_n13811_, new_n13812_, new_n13813_, new_n13814_,
    new_n13815_, new_n13816_, new_n13817_, new_n13818_, new_n13819_,
    new_n13820_, new_n13821_, new_n13822_, new_n13823_, new_n13824_,
    new_n13825_, new_n13826_, new_n13827_, new_n13828_, new_n13829_,
    new_n13830_, new_n13831_, new_n13832_, new_n13833_, new_n13834_,
    new_n13835_, new_n13836_, new_n13837_, new_n13838_, new_n13839_,
    new_n13840_, new_n13841_, new_n13842_, new_n13843_, new_n13844_,
    new_n13845_, new_n13846_, new_n13847_, new_n13848_, new_n13849_,
    new_n13850_, new_n13851_, new_n13852_, new_n13853_, new_n13854_,
    new_n13855_, new_n13856_, new_n13857_, new_n13858_, new_n13859_,
    new_n13860_, new_n13861_, new_n13862_, new_n13863_, new_n13864_,
    new_n13865_, new_n13866_, new_n13867_, new_n13868_, new_n13869_,
    new_n13870_, new_n13871_, new_n13872_, new_n13873_, new_n13874_,
    new_n13875_, new_n13876_, new_n13877_, new_n13878_, new_n13879_,
    new_n13880_, new_n13881_, new_n13882_, new_n13883_, new_n13884_,
    new_n13885_, new_n13886_, new_n13887_, new_n13888_, new_n13889_,
    new_n13890_, new_n13891_, new_n13892_, new_n13893_, new_n13894_,
    new_n13895_, new_n13896_, new_n13897_, new_n13898_, new_n13899_,
    new_n13900_, new_n13901_, new_n13902_, new_n13903_, new_n13904_,
    new_n13905_, new_n13906_, new_n13907_, new_n13908_, new_n13909_,
    new_n13910_, new_n13911_, new_n13912_, new_n13913_, new_n13914_,
    new_n13915_, new_n13916_, new_n13917_, new_n13918_, new_n13919_,
    new_n13920_, new_n13921_, new_n13922_, new_n13923_, new_n13924_,
    new_n13925_, new_n13926_, new_n13927_, new_n13928_, new_n13929_,
    new_n13930_, new_n13931_, new_n13932_, new_n13933_, new_n13934_,
    new_n13935_, new_n13936_, new_n13937_, new_n13938_, new_n13939_,
    new_n13940_, new_n13941_, new_n13942_, new_n13943_, new_n13944_,
    new_n13945_, new_n13946_, new_n13947_, new_n13948_, new_n13949_,
    new_n13950_, new_n13951_, new_n13952_, new_n13953_, new_n13954_,
    new_n13955_, new_n13956_, new_n13957_, new_n13958_, new_n13959_,
    new_n13960_, new_n13961_, new_n13962_, new_n13963_, new_n13964_,
    new_n13965_, new_n13966_, new_n13967_, new_n13968_, new_n13969_,
    new_n13970_, new_n13971_, new_n13972_, new_n13973_, new_n13974_,
    new_n13975_, new_n13976_, new_n13977_, new_n13978_, new_n13979_,
    new_n13980_, new_n13981_, new_n13982_, new_n13983_, new_n13984_,
    new_n13985_, new_n13986_, new_n13987_, new_n13988_, new_n13989_,
    new_n13990_, new_n13991_, new_n13992_, new_n13993_, new_n13994_,
    new_n13995_, new_n13996_, new_n13997_, new_n13998_, new_n13999_,
    new_n14000_, new_n14001_, new_n14002_, new_n14003_, new_n14004_,
    new_n14005_, new_n14006_, new_n14007_, new_n14008_, new_n14009_,
    new_n14010_, new_n14011_, new_n14012_, new_n14013_, new_n14014_,
    new_n14015_, new_n14016_, new_n14017_, new_n14018_, new_n14019_,
    new_n14020_, new_n14021_, new_n14022_, new_n14023_, new_n14024_,
    new_n14025_, new_n14026_, new_n14027_, new_n14028_, new_n14029_,
    new_n14030_, new_n14031_, new_n14032_, new_n14033_, new_n14034_,
    new_n14035_, new_n14036_, new_n14037_, new_n14038_, new_n14039_,
    new_n14040_, new_n14041_, new_n14042_, new_n14043_, new_n14044_,
    new_n14045_, new_n14046_, new_n14047_, new_n14048_, new_n14049_,
    new_n14050_, new_n14051_, new_n14052_, new_n14053_, new_n14054_,
    new_n14055_, new_n14056_, new_n14057_, new_n14058_, new_n14059_,
    new_n14060_, new_n14061_, new_n14062_, new_n14063_, new_n14064_,
    new_n14065_, new_n14066_, new_n14067_, new_n14068_, new_n14069_,
    new_n14070_, new_n14071_, new_n14072_, new_n14073_, new_n14074_,
    new_n14075_, new_n14076_, new_n14077_, new_n14078_, new_n14079_,
    new_n14080_, new_n14081_, new_n14082_, new_n14083_, new_n14084_,
    new_n14085_, new_n14086_, new_n14087_, new_n14088_, new_n14089_,
    new_n14090_, new_n14091_, new_n14092_, new_n14093_, new_n14094_,
    new_n14095_, new_n14096_, new_n14097_, new_n14098_, new_n14099_,
    new_n14100_, new_n14101_, new_n14102_, new_n14103_, new_n14104_,
    new_n14105_, new_n14106_, new_n14107_, new_n14108_, new_n14109_,
    new_n14110_, new_n14111_, new_n14112_, new_n14113_, new_n14114_,
    new_n14115_, new_n14116_, new_n14117_, new_n14118_, new_n14119_,
    new_n14120_, new_n14121_, new_n14122_, new_n14123_, new_n14124_,
    new_n14125_, new_n14126_, new_n14127_, new_n14128_, new_n14129_,
    new_n14130_, new_n14131_, new_n14132_, new_n14133_, new_n14134_,
    new_n14135_, new_n14136_, new_n14137_, new_n14138_, new_n14139_,
    new_n14140_, new_n14141_, new_n14142_, new_n14143_, new_n14144_,
    new_n14145_, new_n14146_, new_n14147_, new_n14148_, new_n14149_,
    new_n14150_, new_n14151_, new_n14152_, new_n14153_, new_n14154_,
    new_n14155_, new_n14156_, new_n14157_, new_n14158_, new_n14159_,
    new_n14160_, new_n14161_, new_n14162_, new_n14163_, new_n14164_,
    new_n14165_, new_n14166_, new_n14167_, new_n14168_, new_n14169_,
    new_n14170_, new_n14171_, new_n14172_, new_n14173_, new_n14174_,
    new_n14175_, new_n14176_, new_n14177_, new_n14178_, new_n14179_,
    new_n14180_, new_n14181_, new_n14182_, new_n14183_, new_n14184_,
    new_n14185_, new_n14186_, new_n14187_, new_n14188_, new_n14189_,
    new_n14190_, new_n14191_, new_n14192_, new_n14193_, new_n14194_,
    new_n14195_, new_n14196_, new_n14197_, new_n14198_, new_n14199_,
    new_n14200_, new_n14201_, new_n14202_, new_n14203_, new_n14204_,
    new_n14205_, new_n14206_, new_n14207_, new_n14208_, new_n14209_,
    new_n14210_, new_n14211_, new_n14212_, new_n14213_, new_n14214_,
    new_n14215_, new_n14216_, new_n14217_, new_n14218_, new_n14219_,
    new_n14220_, new_n14221_, new_n14222_, new_n14223_, new_n14224_,
    new_n14225_, new_n14226_, new_n14227_, new_n14228_, new_n14229_,
    new_n14230_, new_n14231_, new_n14232_, new_n14233_, new_n14234_,
    new_n14235_, new_n14236_, new_n14237_, new_n14238_, new_n14239_,
    new_n14240_, new_n14241_, new_n14242_, new_n14243_, new_n14244_,
    new_n14245_, new_n14246_, new_n14247_, new_n14248_, new_n14249_,
    new_n14250_, new_n14251_, new_n14252_, new_n14253_, new_n14254_,
    new_n14255_, new_n14256_, new_n14257_, new_n14258_, new_n14259_,
    new_n14260_, new_n14261_, new_n14262_, new_n14263_, new_n14264_,
    new_n14265_, new_n14266_, new_n14267_, new_n14268_, new_n14269_,
    new_n14270_, new_n14271_, new_n14272_, new_n14273_, new_n14274_,
    new_n14275_, new_n14276_, new_n14277_, new_n14278_, new_n14279_,
    new_n14280_, new_n14281_, new_n14282_, new_n14283_, new_n14284_,
    new_n14285_, new_n14286_, new_n14287_, new_n14288_, new_n14289_,
    new_n14290_, new_n14291_, new_n14292_, new_n14293_, new_n14294_,
    new_n14295_, new_n14296_, new_n14297_, new_n14298_, new_n14299_,
    new_n14300_, new_n14301_, new_n14302_, new_n14303_, new_n14304_,
    new_n14305_, new_n14306_, new_n14307_, new_n14308_, new_n14309_,
    new_n14310_, new_n14311_, new_n14312_, new_n14313_, new_n14314_,
    new_n14315_, new_n14316_, new_n14317_, new_n14318_, new_n14319_,
    new_n14320_, new_n14321_, new_n14322_, new_n14323_, new_n14324_,
    new_n14325_, new_n14326_, new_n14327_, new_n14328_, new_n14329_,
    new_n14330_, new_n14331_, new_n14332_, new_n14333_, new_n14334_,
    new_n14335_, new_n14336_, new_n14337_, new_n14338_, new_n14339_,
    new_n14340_, new_n14341_, new_n14342_, new_n14343_, new_n14344_,
    new_n14345_, new_n14346_, new_n14347_, new_n14348_, new_n14349_,
    new_n14350_, new_n14351_, new_n14352_, new_n14353_, new_n14354_,
    new_n14355_, new_n14356_, new_n14357_, new_n14358_, new_n14359_,
    new_n14360_, new_n14361_, new_n14362_, new_n14363_, new_n14364_,
    new_n14365_, new_n14366_, new_n14367_, new_n14368_, new_n14369_,
    new_n14370_, new_n14371_, new_n14372_, new_n14373_, new_n14374_,
    new_n14375_, new_n14376_, new_n14377_, new_n14378_, new_n14379_,
    new_n14380_, new_n14381_, new_n14382_, new_n14383_, new_n14384_,
    new_n14385_, new_n14386_, new_n14387_, new_n14388_, new_n14389_,
    new_n14390_, new_n14391_, new_n14392_, new_n14393_, new_n14394_,
    new_n14395_, new_n14396_, new_n14397_, new_n14398_, new_n14399_,
    new_n14400_, new_n14401_, new_n14402_, new_n14403_, new_n14404_,
    new_n14405_, new_n14406_, new_n14407_, new_n14408_, new_n14409_,
    new_n14410_, new_n14411_, new_n14412_, new_n14413_, new_n14414_,
    new_n14415_, new_n14416_, new_n14417_, new_n14418_, new_n14419_,
    new_n14420_, new_n14421_, new_n14422_, new_n14423_, new_n14424_,
    new_n14425_, new_n14426_, new_n14427_, new_n14428_, new_n14429_,
    new_n14430_, new_n14431_, new_n14432_, new_n14433_, new_n14434_,
    new_n14435_, new_n14436_, new_n14437_, new_n14438_, new_n14439_,
    new_n14440_, new_n14441_, new_n14442_, new_n14443_, new_n14444_,
    new_n14445_, new_n14446_, new_n14447_, new_n14448_, new_n14449_,
    new_n14450_, new_n14451_, new_n14452_, new_n14453_, new_n14454_,
    new_n14455_, new_n14456_, new_n14457_, new_n14458_, new_n14459_,
    new_n14460_, new_n14461_, new_n14462_, new_n14463_, new_n14464_,
    new_n14465_, new_n14466_, new_n14467_, new_n14468_, new_n14469_,
    new_n14470_, new_n14471_, new_n14472_, new_n14473_, new_n14474_,
    new_n14475_, new_n14476_, new_n14477_, new_n14478_, new_n14479_,
    new_n14480_, new_n14481_, new_n14482_, new_n14483_, new_n14484_,
    new_n14485_, new_n14486_, new_n14487_, new_n14488_, new_n14489_,
    new_n14490_, new_n14491_, new_n14492_, new_n14493_, new_n14494_,
    new_n14495_, new_n14496_, new_n14497_, new_n14498_, new_n14499_,
    new_n14500_, new_n14501_, new_n14502_, new_n14503_, new_n14504_,
    new_n14505_, new_n14506_, new_n14507_, new_n14508_, new_n14509_,
    new_n14510_, new_n14511_, new_n14512_, new_n14513_, new_n14514_,
    new_n14515_, new_n14516_, new_n14517_, new_n14518_, new_n14519_,
    new_n14520_, new_n14521_, new_n14522_, new_n14523_, new_n14524_,
    new_n14525_, new_n14526_, new_n14527_, new_n14528_, new_n14529_,
    new_n14530_, new_n14531_, new_n14532_, new_n14533_, new_n14534_,
    new_n14535_, new_n14536_, new_n14537_, new_n14538_, new_n14539_,
    new_n14540_, new_n14541_, new_n14542_, new_n14543_, new_n14544_,
    new_n14545_, new_n14546_, new_n14547_, new_n14548_, new_n14549_,
    new_n14550_, new_n14551_, new_n14552_, new_n14553_, new_n14554_,
    new_n14555_, new_n14556_, new_n14557_, new_n14558_, new_n14559_,
    new_n14560_, new_n14561_, new_n14562_, new_n14563_, new_n14564_,
    new_n14565_, new_n14566_, new_n14567_, new_n14568_, new_n14569_,
    new_n14570_, new_n14571_, new_n14572_, new_n14573_, new_n14574_,
    new_n14575_, new_n14576_, new_n14577_, new_n14578_, new_n14579_,
    new_n14580_, new_n14581_, new_n14582_, new_n14583_, new_n14584_,
    new_n14585_, new_n14586_, new_n14587_, new_n14588_, new_n14589_,
    new_n14590_, new_n14591_, new_n14592_, new_n14593_, new_n14594_,
    new_n14595_, new_n14596_, new_n14597_, new_n14598_, new_n14599_,
    new_n14600_, new_n14601_, new_n14602_, new_n14603_, new_n14604_,
    new_n14605_, new_n14606_, new_n14607_, new_n14608_, new_n14609_,
    new_n14610_, new_n14611_, new_n14612_, new_n14613_, new_n14614_,
    new_n14615_, new_n14616_, new_n14617_, new_n14618_, new_n14619_,
    new_n14620_, new_n14621_, new_n14622_, new_n14623_, new_n14624_,
    new_n14625_, new_n14626_, new_n14627_, new_n14628_, new_n14629_,
    new_n14630_, new_n14631_, new_n14632_, new_n14633_, new_n14634_,
    new_n14635_, new_n14636_, new_n14637_, new_n14638_, new_n14639_,
    new_n14640_, new_n14641_, new_n14642_, new_n14643_, new_n14644_,
    new_n14645_, new_n14646_, new_n14647_, new_n14648_, new_n14649_,
    new_n14650_, new_n14651_, new_n14652_, new_n14653_, new_n14654_,
    new_n14655_, new_n14656_, new_n14657_, new_n14658_, new_n14659_,
    new_n14660_, new_n14661_, new_n14662_, new_n14663_, new_n14664_,
    new_n14665_, new_n14666_, new_n14667_, new_n14668_, new_n14669_,
    new_n14670_, new_n14671_, new_n14672_, new_n14673_, new_n14674_,
    new_n14675_, new_n14676_, new_n14677_, new_n14678_, new_n14679_,
    new_n14680_, new_n14681_, new_n14682_, new_n14683_, new_n14684_,
    new_n14685_, new_n14686_, new_n14687_, new_n14688_, new_n14689_,
    new_n14690_, new_n14691_, new_n14692_, new_n14693_, new_n14694_,
    new_n14695_, new_n14696_, new_n14697_, new_n14698_, new_n14699_,
    new_n14700_, new_n14701_, new_n14702_, new_n14703_, new_n14704_,
    new_n14705_, new_n14706_, new_n14707_, new_n14708_, new_n14709_,
    new_n14710_, new_n14711_, new_n14712_, new_n14713_, new_n14714_,
    new_n14715_, new_n14716_, new_n14717_, new_n14718_, new_n14719_,
    new_n14720_, new_n14721_, new_n14722_, new_n14723_, new_n14724_,
    new_n14725_, new_n14726_, new_n14727_, new_n14728_, new_n14729_,
    new_n14730_, new_n14731_, new_n14732_, new_n14733_, new_n14734_,
    new_n14735_, new_n14736_, new_n14737_, new_n14738_, new_n14739_,
    new_n14740_, new_n14741_, new_n14742_, new_n14743_, new_n14744_,
    new_n14745_, new_n14746_, new_n14747_, new_n14748_, new_n14749_,
    new_n14750_, new_n14751_, new_n14752_, new_n14753_, new_n14754_,
    new_n14755_, new_n14756_, new_n14757_, new_n14758_, new_n14759_,
    new_n14760_, new_n14761_, new_n14762_, new_n14763_, new_n14764_,
    new_n14765_, new_n14766_, new_n14767_, new_n14768_, new_n14769_,
    new_n14770_, new_n14771_, new_n14772_, new_n14773_, new_n14774_,
    new_n14775_, new_n14776_, new_n14777_, new_n14778_, new_n14779_,
    new_n14780_, new_n14781_, new_n14782_, new_n14783_, new_n14784_,
    new_n14785_, new_n14786_, new_n14787_, new_n14788_, new_n14789_,
    new_n14790_, new_n14791_, new_n14792_, new_n14793_, new_n14794_,
    new_n14795_, new_n14796_, new_n14797_, new_n14798_, new_n14799_,
    new_n14800_, new_n14801_, new_n14802_, new_n14803_, new_n14804_,
    new_n14805_, new_n14806_, new_n14807_, new_n14808_, new_n14809_,
    new_n14810_, new_n14811_, new_n14812_, new_n14813_, new_n14814_,
    new_n14815_, new_n14816_, new_n14817_, new_n14818_, new_n14819_,
    new_n14820_, new_n14821_, new_n14822_, new_n14823_, new_n14824_,
    new_n14825_, new_n14826_, new_n14827_, new_n14828_, new_n14829_,
    new_n14830_, new_n14831_, new_n14832_, new_n14833_, new_n14834_,
    new_n14835_, new_n14836_, new_n14837_, new_n14838_, new_n14839_,
    new_n14840_, new_n14841_, new_n14842_, new_n14843_, new_n14844_,
    new_n14845_, new_n14846_, new_n14847_, new_n14848_, new_n14849_,
    new_n14850_, new_n14851_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14907_, new_n14908_, new_n14909_,
    new_n14910_, new_n14911_, new_n14912_, new_n14913_, new_n14914_,
    new_n14915_, new_n14916_, new_n14917_, new_n14918_, new_n14919_,
    new_n14920_, new_n14921_, new_n14922_, new_n14923_, new_n14924_,
    new_n14925_, new_n14926_, new_n14927_, new_n14928_, new_n14929_,
    new_n14930_, new_n14931_, new_n14932_, new_n14933_, new_n14934_,
    new_n14935_, new_n14936_, new_n14937_, new_n14938_, new_n14939_,
    new_n14940_, new_n14941_, new_n14942_, new_n14943_, new_n14944_,
    new_n14945_, new_n14946_, new_n14947_, new_n14948_, new_n14949_,
    new_n14950_, new_n14951_, new_n14952_, new_n14953_, new_n14954_,
    new_n14955_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14960_, new_n14961_, new_n14962_, new_n14963_, new_n14964_,
    new_n14965_, new_n14966_, new_n14967_, new_n14968_, new_n14969_,
    new_n14970_, new_n14971_, new_n14972_, new_n14973_, new_n14974_,
    new_n14975_, new_n14976_, new_n14977_, new_n14978_, new_n14979_,
    new_n14980_, new_n14981_, new_n14982_, new_n14983_, new_n14984_,
    new_n14985_, new_n14986_, new_n14987_, new_n14988_, new_n14989_,
    new_n14990_, new_n14991_, new_n14992_, new_n14993_, new_n14994_,
    new_n14995_, new_n14996_, new_n14997_, new_n14998_, new_n14999_,
    new_n15000_, new_n15001_, new_n15002_, new_n15003_, new_n15004_,
    new_n15005_, new_n15006_, new_n15007_, new_n15008_, new_n15009_,
    new_n15010_, new_n15011_, new_n15012_, new_n15013_, new_n15014_,
    new_n15015_, new_n15016_, new_n15017_, new_n15018_, new_n15019_,
    new_n15020_, new_n15021_, new_n15022_, new_n15023_, new_n15024_,
    new_n15025_, new_n15026_, new_n15027_, new_n15028_, new_n15029_,
    new_n15030_, new_n15031_, new_n15032_, new_n15033_, new_n15034_,
    new_n15035_, new_n15036_, new_n15037_, new_n15038_, new_n15039_,
    new_n15040_, new_n15041_, new_n15042_, new_n15043_, new_n15044_,
    new_n15045_, new_n15046_, new_n15047_, new_n15048_, new_n15049_,
    new_n15050_, new_n15051_, new_n15052_, new_n15053_, new_n15054_,
    new_n15055_, new_n15056_, new_n15057_, new_n15058_, new_n15059_,
    new_n15060_, new_n15061_, new_n15062_, new_n15063_, new_n15064_,
    new_n15065_, new_n15066_, new_n15067_, new_n15068_, new_n15069_,
    new_n15070_, new_n15071_, new_n15072_, new_n15073_, new_n15074_,
    new_n15075_, new_n15076_, new_n15077_, new_n15078_, new_n15079_,
    new_n15080_, new_n15081_, new_n15082_, new_n15083_, new_n15084_,
    new_n15085_, new_n15086_, new_n15087_, new_n15088_, new_n15089_,
    new_n15090_, new_n15091_, new_n15092_, new_n15093_, new_n15094_,
    new_n15095_, new_n15096_, new_n15097_, new_n15098_, new_n15099_,
    new_n15100_, new_n15101_, new_n15102_, new_n15103_, new_n15104_,
    new_n15105_, new_n15106_, new_n15107_, new_n15108_, new_n15109_,
    new_n15110_, new_n15111_, new_n15112_, new_n15113_, new_n15114_,
    new_n15115_, new_n15116_, new_n15117_, new_n15118_, new_n15119_,
    new_n15120_, new_n15121_, new_n15122_, new_n15123_, new_n15124_,
    new_n15125_, new_n15126_, new_n15127_, new_n15128_, new_n15129_,
    new_n15130_, new_n15131_, new_n15132_, new_n15133_, new_n15134_,
    new_n15135_, new_n15136_, new_n15137_, new_n15138_, new_n15139_,
    new_n15140_, new_n15141_, new_n15142_, new_n15143_, new_n15144_,
    new_n15145_, new_n15146_, new_n15147_, new_n15148_, new_n15149_,
    new_n15150_, new_n15151_, new_n15152_, new_n15153_, new_n15154_,
    new_n15155_, new_n15156_, new_n15157_, new_n15158_, new_n15159_,
    new_n15160_, new_n15161_, new_n15162_, new_n15163_, new_n15164_,
    new_n15165_, new_n15166_, new_n15167_, new_n15168_, new_n15169_,
    new_n15170_, new_n15171_, new_n15172_, new_n15173_, new_n15174_,
    new_n15175_, new_n15176_, new_n15177_, new_n15178_, new_n15179_,
    new_n15180_, new_n15181_, new_n15182_, new_n15183_, new_n15184_,
    new_n15185_, new_n15186_, new_n15187_, new_n15188_, new_n15189_,
    new_n15190_, new_n15191_, new_n15192_, new_n15193_, new_n15194_,
    new_n15195_, new_n15196_, new_n15197_, new_n15198_, new_n15199_,
    new_n15200_, new_n15201_, new_n15202_, new_n15203_, new_n15204_,
    new_n15205_, new_n15206_, new_n15207_, new_n15208_, new_n15209_,
    new_n15210_, new_n15211_, new_n15212_, new_n15213_, new_n15214_,
    new_n15215_, new_n15216_, new_n15217_, new_n15218_, new_n15219_,
    new_n15220_, new_n15221_, new_n15222_, new_n15223_, new_n15224_,
    new_n15225_, new_n15226_, new_n15227_, new_n15228_, new_n15229_,
    new_n15230_, new_n15231_, new_n15232_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15369_,
    new_n15370_, new_n15371_, new_n15372_, new_n15373_, new_n15374_,
    new_n15375_, new_n15376_, new_n15377_, new_n15378_, new_n15379_,
    new_n15380_, new_n15381_, new_n15382_, new_n15383_, new_n15384_,
    new_n15385_, new_n15386_, new_n15387_, new_n15388_, new_n15389_,
    new_n15390_, new_n15391_, new_n15392_, new_n15393_, new_n15394_,
    new_n15395_, new_n15396_, new_n15397_, new_n15398_, new_n15399_,
    new_n15400_, new_n15401_, new_n15402_, new_n15403_, new_n15404_,
    new_n15405_, new_n15406_, new_n15407_, new_n15408_, new_n15409_,
    new_n15410_, new_n15411_, new_n15412_, new_n15413_, new_n15414_,
    new_n15415_, new_n15416_, new_n15417_, new_n15418_, new_n15419_,
    new_n15420_, new_n15421_, new_n15422_, new_n15423_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15428_, new_n15429_,
    new_n15430_, new_n15431_, new_n15432_, new_n15433_, new_n15434_,
    new_n15435_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15469_,
    new_n15470_, new_n15471_, new_n15472_, new_n15473_, new_n15474_,
    new_n15475_, new_n15476_, new_n15477_, new_n15478_, new_n15479_,
    new_n15480_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15488_, new_n15489_,
    new_n15490_, new_n15491_, new_n15492_, new_n15493_, new_n15494_,
    new_n15495_, new_n15496_, new_n15497_, new_n15498_, new_n15499_,
    new_n15500_, new_n15501_, new_n15502_, new_n15503_, new_n15504_,
    new_n15505_, new_n15506_, new_n15507_, new_n15508_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15575_, new_n15576_, new_n15577_, new_n15578_, new_n15579_,
    new_n15580_, new_n15581_, new_n15582_, new_n15583_, new_n15584_,
    new_n15585_, new_n15586_, new_n15587_, new_n15588_, new_n15589_,
    new_n15590_, new_n15591_, new_n15592_, new_n15593_, new_n15594_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15601_, new_n15602_, new_n15603_, new_n15604_,
    new_n15605_, new_n15606_, new_n15607_, new_n15608_, new_n15609_,
    new_n15610_, new_n15611_, new_n15612_, new_n15613_, new_n15614_,
    new_n15615_, new_n15616_, new_n15617_, new_n15618_, new_n15619_,
    new_n15620_, new_n15621_, new_n15622_, new_n15623_, new_n15624_,
    new_n15625_, new_n15626_, new_n15627_, new_n15628_, new_n15629_,
    new_n15630_, new_n15631_, new_n15632_, new_n15633_, new_n15634_,
    new_n15635_, new_n15636_, new_n15637_, new_n15638_, new_n15639_,
    new_n15640_, new_n15641_, new_n15642_, new_n15643_, new_n15644_,
    new_n15645_, new_n15646_, new_n15647_, new_n15648_, new_n15649_,
    new_n15650_, new_n15651_, new_n15652_, new_n15653_, new_n15654_,
    new_n15655_, new_n15656_, new_n15657_, new_n15658_, new_n15659_,
    new_n15660_, new_n15661_, new_n15662_, new_n15663_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15674_,
    new_n15675_, new_n15676_, new_n15677_, new_n15678_, new_n15679_,
    new_n15680_, new_n15681_, new_n15682_, new_n15683_, new_n15684_,
    new_n15685_, new_n15686_, new_n15687_, new_n15688_, new_n15689_,
    new_n15690_, new_n15691_, new_n15692_, new_n15693_, new_n15694_,
    new_n15695_, new_n15696_, new_n15697_, new_n15698_, new_n15699_,
    new_n15700_, new_n15701_, new_n15702_, new_n15703_, new_n15704_,
    new_n15705_, new_n15706_, new_n15707_, new_n15708_, new_n15709_,
    new_n15710_, new_n15711_, new_n15712_, new_n15713_, new_n15714_,
    new_n15715_, new_n15716_, new_n15717_, new_n15718_, new_n15719_,
    new_n15720_, new_n15721_, new_n15722_, new_n15723_, new_n15724_,
    new_n15725_, new_n15726_, new_n15727_, new_n15728_, new_n15729_,
    new_n15730_, new_n15731_, new_n15732_, new_n15733_, new_n15734_,
    new_n15735_, new_n15736_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15755_, new_n15756_, new_n15757_, new_n15758_, new_n15759_,
    new_n15760_, new_n15761_, new_n15762_, new_n15763_, new_n15764_,
    new_n15765_, new_n15766_, new_n15767_, new_n15768_, new_n15769_,
    new_n15770_, new_n15771_, new_n15772_, new_n15773_, new_n15774_,
    new_n15775_, new_n15776_, new_n15777_, new_n15778_, new_n15779_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15786_, new_n15787_, new_n15788_, new_n15789_,
    new_n15790_, new_n15791_, new_n15792_, new_n15793_, new_n15794_,
    new_n15795_, new_n15796_, new_n15797_, new_n15798_, new_n15799_,
    new_n15800_, new_n15801_, new_n15802_, new_n15803_, new_n15804_,
    new_n15805_, new_n15806_, new_n15807_, new_n15808_, new_n15809_,
    new_n15810_, new_n15811_, new_n15812_, new_n15813_, new_n15814_,
    new_n15815_, new_n15816_, new_n15817_, new_n15818_, new_n15819_,
    new_n15820_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15865_, new_n15866_, new_n15867_, new_n15868_, new_n15869_,
    new_n15870_, new_n15871_, new_n15872_, new_n15873_, new_n15874_,
    new_n15875_, new_n15876_, new_n15877_, new_n15878_, new_n15879_,
    new_n15880_, new_n15881_, new_n15882_, new_n15883_, new_n15884_,
    new_n15885_, new_n15886_, new_n15887_, new_n15888_, new_n15889_,
    new_n15890_, new_n15891_, new_n15892_, new_n15893_, new_n15894_,
    new_n15895_, new_n15896_, new_n15897_, new_n15898_, new_n15899_,
    new_n15900_, new_n15901_, new_n15902_, new_n15903_, new_n15904_,
    new_n15905_, new_n15906_, new_n15907_, new_n15908_, new_n15909_,
    new_n15910_, new_n15911_, new_n15912_, new_n15913_, new_n15914_,
    new_n15915_, new_n15916_, new_n15917_, new_n15918_, new_n15919_,
    new_n15920_, new_n15921_, new_n15922_, new_n15923_, new_n15924_,
    new_n15925_, new_n15926_, new_n15927_, new_n15928_, new_n15929_,
    new_n15930_, new_n15931_, new_n15932_, new_n15933_, new_n15934_,
    new_n15935_, new_n15936_, new_n15937_, new_n15938_, new_n15939_,
    new_n15940_, new_n15941_, new_n15942_, new_n15943_, new_n15944_,
    new_n15945_, new_n15946_, new_n15947_, new_n15948_, new_n15949_,
    new_n15950_, new_n15951_, new_n15952_, new_n15953_, new_n15954_,
    new_n15955_, new_n15956_, new_n15957_, new_n15958_, new_n15959_,
    new_n15960_, new_n15961_, new_n15962_, new_n15963_, new_n15964_,
    new_n15965_, new_n15966_, new_n15967_, new_n15968_, new_n15969_,
    new_n15970_, new_n15971_, new_n15972_, new_n15973_, new_n15974_,
    new_n15975_, new_n15976_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15987_, new_n15988_, new_n15989_,
    new_n15990_, new_n15991_, new_n15992_, new_n15993_, new_n15994_,
    new_n15995_, new_n15996_, new_n15997_, new_n15998_, new_n15999_,
    new_n16000_, new_n16001_, new_n16002_, new_n16003_, new_n16004_,
    new_n16005_, new_n16006_, new_n16007_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16012_, new_n16013_, new_n16014_,
    new_n16015_, new_n16016_, new_n16017_, new_n16018_, new_n16019_,
    new_n16020_, new_n16021_, new_n16022_, new_n16023_, new_n16024_,
    new_n16025_, new_n16026_, new_n16027_, new_n16028_, new_n16029_,
    new_n16030_, new_n16031_, new_n16032_, new_n16033_, new_n16034_,
    new_n16035_, new_n16036_, new_n16037_, new_n16038_, new_n16039_,
    new_n16040_, new_n16041_, new_n16042_, new_n16043_, new_n16044_,
    new_n16045_, new_n16046_, new_n16047_, new_n16048_, new_n16049_,
    new_n16050_, new_n16051_, new_n16052_, new_n16053_, new_n16054_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16060_, new_n16061_, new_n16062_, new_n16063_, new_n16064_,
    new_n16065_, new_n16066_, new_n16067_, new_n16068_, new_n16069_,
    new_n16070_, new_n16071_, new_n16072_, new_n16073_, new_n16074_,
    new_n16075_, new_n16076_, new_n16077_, new_n16078_, new_n16079_,
    new_n16080_, new_n16081_, new_n16082_, new_n16083_, new_n16084_,
    new_n16085_, new_n16086_, new_n16087_, new_n16088_, new_n16089_,
    new_n16090_, new_n16091_, new_n16092_, new_n16093_, new_n16094_,
    new_n16095_, new_n16096_, new_n16097_, new_n16098_, new_n16099_,
    new_n16100_, new_n16101_, new_n16102_, new_n16103_, new_n16104_,
    new_n16105_, new_n16106_, new_n16107_, new_n16108_, new_n16109_,
    new_n16110_, new_n16111_, new_n16112_, new_n16113_, new_n16114_,
    new_n16115_, new_n16116_, new_n16117_, new_n16118_, new_n16119_,
    new_n16120_, new_n16121_, new_n16122_, new_n16123_, new_n16124_,
    new_n16125_, new_n16126_, new_n16127_, new_n16128_, new_n16129_,
    new_n16130_, new_n16131_, new_n16132_, new_n16133_, new_n16134_,
    new_n16135_, new_n16136_, new_n16137_, new_n16138_, new_n16139_,
    new_n16140_, new_n16141_, new_n16142_, new_n16143_, new_n16144_,
    new_n16145_, new_n16146_, new_n16147_, new_n16148_, new_n16149_,
    new_n16150_, new_n16151_, new_n16152_, new_n16153_, new_n16154_,
    new_n16155_, new_n16156_, new_n16157_, new_n16158_, new_n16159_,
    new_n16160_, new_n16161_, new_n16162_, new_n16163_, new_n16164_,
    new_n16165_, new_n16166_, new_n16167_, new_n16168_, new_n16169_,
    new_n16170_, new_n16171_, new_n16172_, new_n16173_, new_n16174_,
    new_n16175_, new_n16176_, new_n16177_, new_n16178_, new_n16179_,
    new_n16180_, new_n16181_, new_n16182_, new_n16183_, new_n16184_,
    new_n16185_, new_n16186_, new_n16187_, new_n16188_, new_n16189_,
    new_n16190_, new_n16191_, new_n16192_, new_n16193_, new_n16194_,
    new_n16195_, new_n16196_, new_n16197_, new_n16198_, new_n16199_,
    new_n16200_, new_n16201_, new_n16202_, new_n16203_, new_n16204_,
    new_n16205_, new_n16206_, new_n16207_, new_n16208_, new_n16209_,
    new_n16210_, new_n16211_, new_n16212_, new_n16213_, new_n16214_,
    new_n16215_, new_n16216_, new_n16217_, new_n16218_, new_n16219_,
    new_n16220_, new_n16221_, new_n16222_, new_n16223_, new_n16224_,
    new_n16225_, new_n16226_, new_n16227_, new_n16228_, new_n16229_,
    new_n16230_, new_n16231_, new_n16232_, new_n16233_, new_n16234_,
    new_n16235_, new_n16236_, new_n16237_, new_n16238_, new_n16239_,
    new_n16240_, new_n16241_, new_n16242_, new_n16243_, new_n16244_,
    new_n16245_, new_n16246_, new_n16247_, new_n16248_, new_n16249_,
    new_n16250_, new_n16251_, new_n16252_, new_n16253_, new_n16254_,
    new_n16255_, new_n16256_, new_n16257_, new_n16258_, new_n16259_,
    new_n16260_, new_n16261_, new_n16262_, new_n16263_, new_n16264_,
    new_n16265_, new_n16266_, new_n16267_, new_n16268_, new_n16269_,
    new_n16270_, new_n16271_, new_n16272_, new_n16273_, new_n16274_,
    new_n16275_, new_n16276_, new_n16277_, new_n16278_, new_n16279_,
    new_n16280_, new_n16281_, new_n16282_, new_n16283_, new_n16284_,
    new_n16285_, new_n16286_, new_n16287_, new_n16288_, new_n16289_,
    new_n16290_, new_n16291_, new_n16292_, new_n16293_, new_n16294_,
    new_n16295_, new_n16296_, new_n16297_, new_n16298_, new_n16299_,
    new_n16300_, new_n16301_, new_n16302_, new_n16303_, new_n16304_,
    new_n16305_, new_n16306_, new_n16307_, new_n16308_, new_n16309_,
    new_n16310_, new_n16311_, new_n16312_, new_n16313_, new_n16314_,
    new_n16315_, new_n16316_, new_n16317_, new_n16318_, new_n16319_,
    new_n16320_, new_n16321_, new_n16322_, new_n16323_, new_n16324_,
    new_n16325_, new_n16326_, new_n16327_, new_n16328_, new_n16329_,
    new_n16330_, new_n16331_, new_n16332_, new_n16333_, new_n16334_,
    new_n16335_, new_n16336_, new_n16337_, new_n16338_, new_n16339_,
    new_n16340_, new_n16341_, new_n16342_, new_n16343_, new_n16344_,
    new_n16345_, new_n16346_, new_n16347_, new_n16348_, new_n16349_,
    new_n16350_, new_n16351_, new_n16352_, new_n16353_, new_n16354_,
    new_n16355_, new_n16356_, new_n16357_, new_n16358_, new_n16359_,
    new_n16360_, new_n16361_, new_n16362_, new_n16363_, new_n16364_,
    new_n16365_, new_n16366_, new_n16367_, new_n16368_, new_n16369_,
    new_n16370_, new_n16371_, new_n16372_, new_n16373_, new_n16374_,
    new_n16375_, new_n16376_, new_n16377_, new_n16378_, new_n16379_,
    new_n16380_, new_n16381_, new_n16382_, new_n16383_, new_n16384_,
    new_n16385_, new_n16386_, new_n16387_, new_n16388_, new_n16389_,
    new_n16390_, new_n16391_, new_n16392_, new_n16393_, new_n16394_,
    new_n16395_, new_n16396_, new_n16397_, new_n16398_, new_n16399_,
    new_n16400_, new_n16401_, new_n16402_, new_n16403_, new_n16404_,
    new_n16405_, new_n16406_, new_n16407_, new_n16408_, new_n16409_,
    new_n16410_, new_n16411_, new_n16412_, new_n16413_, new_n16414_,
    new_n16415_, new_n16416_, new_n16417_, new_n16418_, new_n16419_,
    new_n16420_, new_n16421_, new_n16422_, new_n16423_, new_n16424_,
    new_n16425_, new_n16426_, new_n16427_, new_n16428_, new_n16429_,
    new_n16430_, new_n16431_, new_n16432_, new_n16433_, new_n16434_,
    new_n16435_, new_n16436_, new_n16437_, new_n16438_, new_n16439_,
    new_n16440_, new_n16441_, new_n16442_, new_n16443_, new_n16444_,
    new_n16445_, new_n16446_, new_n16447_, new_n16448_, new_n16449_,
    new_n16450_, new_n16451_, new_n16452_, new_n16453_, new_n16454_,
    new_n16455_, new_n16456_, new_n16457_, new_n16458_, new_n16459_,
    new_n16460_, new_n16461_, new_n16462_, new_n16463_, new_n16464_,
    new_n16465_, new_n16466_, new_n16467_, new_n16468_, new_n16469_,
    new_n16470_, new_n16471_, new_n16472_, new_n16473_, new_n16474_,
    new_n16475_, new_n16476_, new_n16477_, new_n16478_, new_n16479_,
    new_n16480_, new_n16481_, new_n16482_, new_n16483_, new_n16484_,
    new_n16485_, new_n16486_, new_n16487_, new_n16488_, new_n16489_,
    new_n16490_, new_n16491_, new_n16492_, new_n16493_, new_n16494_,
    new_n16495_, new_n16496_, new_n16497_, new_n16498_, new_n16499_,
    new_n16500_, new_n16501_, new_n16502_, new_n16503_, new_n16504_,
    new_n16505_, new_n16506_, new_n16507_, new_n16508_, new_n16509_,
    new_n16510_, new_n16511_, new_n16512_, new_n16513_, new_n16514_,
    new_n16515_, new_n16516_, new_n16517_, new_n16518_, new_n16519_,
    new_n16520_, new_n16521_, new_n16522_, new_n16523_, new_n16524_,
    new_n16525_, new_n16526_, new_n16527_, new_n16528_, new_n16529_,
    new_n16530_, new_n16531_, new_n16532_, new_n16533_, new_n16534_,
    new_n16535_, new_n16536_, new_n16537_, new_n16538_, new_n16539_,
    new_n16540_, new_n16541_, new_n16542_, new_n16543_, new_n16544_,
    new_n16545_, new_n16546_, new_n16547_, new_n16548_, new_n16549_,
    new_n16550_, new_n16551_, new_n16552_, new_n16553_, new_n16554_,
    new_n16555_, new_n16556_, new_n16557_, new_n16558_, new_n16559_,
    new_n16560_, new_n16561_, new_n16562_, new_n16563_, new_n16564_,
    new_n16565_, new_n16566_, new_n16567_, new_n16568_, new_n16569_,
    new_n16570_, new_n16571_, new_n16572_, new_n16573_, new_n16574_,
    new_n16575_, new_n16576_, new_n16577_, new_n16578_, new_n16579_,
    new_n16580_, new_n16581_, new_n16582_, new_n16583_, new_n16584_,
    new_n16585_, new_n16586_, new_n16587_, new_n16588_, new_n16589_,
    new_n16590_, new_n16591_, new_n16592_, new_n16593_, new_n16594_,
    new_n16595_, new_n16596_, new_n16597_, new_n16598_, new_n16599_,
    new_n16600_, new_n16601_, new_n16602_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16610_, new_n16611_, new_n16612_, new_n16613_, new_n16614_,
    new_n16615_, new_n16616_, new_n16617_, new_n16618_, new_n16619_,
    new_n16620_, new_n16621_, new_n16622_, new_n16623_, new_n16624_,
    new_n16625_, new_n16626_, new_n16627_, new_n16628_, new_n16629_,
    new_n16630_, new_n16631_, new_n16632_, new_n16633_, new_n16634_,
    new_n16635_, new_n16636_, new_n16637_, new_n16638_, new_n16639_,
    new_n16640_, new_n16641_, new_n16642_, new_n16643_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16650_, new_n16651_, new_n16652_, new_n16653_, new_n16654_,
    new_n16655_, new_n16656_, new_n16657_, new_n16658_, new_n16659_,
    new_n16660_, new_n16661_, new_n16662_, new_n16663_, new_n16664_,
    new_n16665_, new_n16666_, new_n16667_, new_n16668_, new_n16669_,
    new_n16670_, new_n16671_, new_n16672_, new_n16673_, new_n16674_,
    new_n16675_, new_n16676_, new_n16677_, new_n16678_, new_n16679_,
    new_n16680_, new_n16681_, new_n16682_, new_n16683_, new_n16684_,
    new_n16685_, new_n16686_, new_n16687_, new_n16688_, new_n16689_,
    new_n16690_, new_n16691_, new_n16692_, new_n16693_, new_n16694_,
    new_n16695_, new_n16696_, new_n16697_, new_n16698_, new_n16699_,
    new_n16700_, new_n16701_, new_n16702_, new_n16703_, new_n16704_,
    new_n16705_, new_n16706_, new_n16707_, new_n16708_, new_n16709_,
    new_n16710_, new_n16711_, new_n16712_, new_n16713_, new_n16714_,
    new_n16715_, new_n16716_, new_n16717_, new_n16718_, new_n16719_,
    new_n16720_, new_n16721_, new_n16722_, new_n16723_, new_n16724_,
    new_n16725_, new_n16726_, new_n16727_, new_n16728_, new_n16729_,
    new_n16730_, new_n16731_, new_n16732_, new_n16733_, new_n16734_,
    new_n16735_, new_n16736_, new_n16737_, new_n16738_, new_n16739_,
    new_n16740_, new_n16741_, new_n16742_, new_n16743_, new_n16744_,
    new_n16745_, new_n16746_, new_n16747_, new_n16748_, new_n16749_,
    new_n16750_, new_n16751_, new_n16752_, new_n16753_, new_n16754_,
    new_n16755_, new_n16756_, new_n16757_, new_n16758_, new_n16759_,
    new_n16760_, new_n16761_, new_n16762_, new_n16763_, new_n16764_,
    new_n16765_, new_n16766_, new_n16767_, new_n16768_, new_n16769_,
    new_n16770_, new_n16771_, new_n16772_, new_n16773_, new_n16774_,
    new_n16775_, new_n16776_, new_n16777_, new_n16778_, new_n16779_,
    new_n16780_, new_n16781_, new_n16782_, new_n16783_, new_n16784_,
    new_n16785_, new_n16786_, new_n16787_, new_n16788_, new_n16789_,
    new_n16790_, new_n16791_, new_n16792_, new_n16793_, new_n16794_,
    new_n16795_, new_n16796_, new_n16797_, new_n16798_, new_n16799_,
    new_n16800_, new_n16801_, new_n16802_, new_n16803_, new_n16804_,
    new_n16805_, new_n16806_, new_n16807_, new_n16808_, new_n16809_,
    new_n16810_, new_n16811_, new_n16812_, new_n16813_, new_n16814_,
    new_n16815_, new_n16816_, new_n16817_, new_n16818_, new_n16819_,
    new_n16820_, new_n16821_, new_n16822_, new_n16823_, new_n16824_,
    new_n16825_, new_n16826_, new_n16827_, new_n16828_, new_n16829_,
    new_n16830_, new_n16831_, new_n16832_, new_n16833_, new_n16834_,
    new_n16835_, new_n16836_, new_n16837_, new_n16838_, new_n16839_,
    new_n16840_, new_n16841_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16848_, new_n16849_,
    new_n16850_, new_n16851_, new_n16852_, new_n16853_, new_n16854_,
    new_n16855_, new_n16856_, new_n16857_, new_n16858_, new_n16859_,
    new_n16860_, new_n16861_, new_n16862_, new_n16863_, new_n16864_,
    new_n16865_, new_n16866_, new_n16867_, new_n16868_, new_n16869_,
    new_n16870_, new_n16871_, new_n16872_, new_n16873_, new_n16874_,
    new_n16875_, new_n16876_, new_n16877_, new_n16878_, new_n16879_,
    new_n16880_, new_n16881_, new_n16882_, new_n16883_, new_n16884_,
    new_n16885_, new_n16886_, new_n16887_, new_n16888_, new_n16889_,
    new_n16890_, new_n16891_, new_n16892_, new_n16893_, new_n16894_,
    new_n16895_, new_n16896_, new_n16897_, new_n16898_, new_n16899_,
    new_n16900_, new_n16901_, new_n16902_, new_n16903_, new_n16904_,
    new_n16905_, new_n16906_, new_n16907_, new_n16908_, new_n16909_,
    new_n16910_, new_n16911_, new_n16912_, new_n16913_, new_n16914_,
    new_n16915_, new_n16916_, new_n16917_, new_n16918_, new_n16919_,
    new_n16920_, new_n16921_, new_n16922_, new_n16923_, new_n16924_,
    new_n16925_, new_n16926_, new_n16927_, new_n16928_, new_n16929_,
    new_n16930_, new_n16931_, new_n16932_, new_n16933_, new_n16934_,
    new_n16935_, new_n16936_, new_n16937_, new_n16938_, new_n16939_,
    new_n16940_, new_n16941_, new_n16942_, new_n16943_, new_n16944_,
    new_n16945_, new_n16946_, new_n16947_, new_n16948_, new_n16949_,
    new_n16950_, new_n16951_, new_n16952_, new_n16953_, new_n16954_,
    new_n16955_, new_n16956_, new_n16957_, new_n16958_, new_n16959_,
    new_n16960_, new_n16961_, new_n16962_, new_n16963_, new_n16964_,
    new_n16965_, new_n16966_, new_n16967_, new_n16968_, new_n16969_,
    new_n16970_, new_n16971_, new_n16972_, new_n16973_, new_n16974_,
    new_n16975_, new_n16976_, new_n16977_, new_n16978_, new_n16979_,
    new_n16980_, new_n16981_, new_n16982_, new_n16983_, new_n16984_,
    new_n16985_, new_n16986_, new_n16987_, new_n16988_, new_n16989_,
    new_n16990_, new_n16991_, new_n16992_, new_n16993_, new_n16994_,
    new_n16995_, new_n16996_, new_n16997_, new_n16998_, new_n16999_,
    new_n17000_, new_n17001_, new_n17002_, new_n17003_, new_n17004_,
    new_n17005_, new_n17006_, new_n17007_, new_n17008_, new_n17009_,
    new_n17010_, new_n17011_, new_n17012_, new_n17013_, new_n17014_,
    new_n17015_, new_n17016_, new_n17017_, new_n17018_, new_n17019_,
    new_n17020_, new_n17021_, new_n17022_, new_n17023_, new_n17024_,
    new_n17025_, new_n17026_, new_n17027_, new_n17028_, new_n17029_,
    new_n17030_, new_n17031_, new_n17032_, new_n17033_, new_n17034_,
    new_n17035_, new_n17036_, new_n17037_, new_n17038_, new_n17039_,
    new_n17040_, new_n17041_, new_n17042_, new_n17043_, new_n17044_,
    new_n17045_, new_n17046_, new_n17047_, new_n17048_, new_n17049_,
    new_n17050_, new_n17051_, new_n17052_, new_n17053_, new_n17054_,
    new_n17055_, new_n17056_, new_n17057_, new_n17058_, new_n17059_,
    new_n17060_, new_n17061_, new_n17062_, new_n17063_, new_n17064_,
    new_n17065_, new_n17066_, new_n17067_, new_n17068_, new_n17069_,
    new_n17070_, new_n17071_, new_n17072_, new_n17073_, new_n17074_,
    new_n17075_, new_n17076_, new_n17077_, new_n17078_, new_n17079_,
    new_n17080_, new_n17081_, new_n17082_, new_n17083_, new_n17084_,
    new_n17085_, new_n17086_, new_n17087_, new_n17088_, new_n17089_,
    new_n17090_, new_n17091_, new_n17092_, new_n17093_, new_n17094_,
    new_n17095_, new_n17096_, new_n17097_, new_n17098_, new_n17099_,
    new_n17100_, new_n17101_, new_n17102_, new_n17103_, new_n17104_,
    new_n17105_, new_n17106_, new_n17107_, new_n17108_, new_n17109_,
    new_n17110_, new_n17111_, new_n17112_, new_n17113_, new_n17114_,
    new_n17115_, new_n17116_, new_n17117_, new_n17118_, new_n17119_,
    new_n17120_, new_n17121_, new_n17122_, new_n17123_, new_n17124_,
    new_n17125_, new_n17126_, new_n17127_, new_n17128_, new_n17129_,
    new_n17130_, new_n17131_, new_n17132_, new_n17133_, new_n17134_,
    new_n17135_, new_n17136_, new_n17137_, new_n17138_, new_n17139_,
    new_n17140_, new_n17141_, new_n17142_, new_n17143_, new_n17144_,
    new_n17145_, new_n17146_, new_n17147_, new_n17148_, new_n17149_,
    new_n17150_, new_n17151_, new_n17152_, new_n17153_, new_n17154_,
    new_n17155_, new_n17156_, new_n17157_, new_n17158_, new_n17159_,
    new_n17160_, new_n17161_, new_n17162_, new_n17163_, new_n17164_,
    new_n17165_, new_n17166_, new_n17167_, new_n17168_, new_n17169_,
    new_n17170_, new_n17171_, new_n17172_, new_n17173_, new_n17174_,
    new_n17175_, new_n17176_, new_n17177_, new_n17178_, new_n17179_,
    new_n17180_, new_n17181_, new_n17182_, new_n17183_, new_n17184_,
    new_n17185_, new_n17186_, new_n17187_, new_n17188_, new_n17189_,
    new_n17190_, new_n17191_, new_n17192_, new_n17193_, new_n17194_,
    new_n17195_, new_n17196_, new_n17197_, new_n17198_, new_n17199_,
    new_n17200_, new_n17201_, new_n17202_, new_n17203_, new_n17204_,
    new_n17205_, new_n17206_, new_n17207_, new_n17208_, new_n17209_,
    new_n17210_, new_n17211_, new_n17212_, new_n17213_, new_n17214_,
    new_n17215_, new_n17216_, new_n17217_, new_n17218_, new_n17219_,
    new_n17220_, new_n17221_, new_n17222_, new_n17223_, new_n17224_,
    new_n17225_, new_n17226_, new_n17227_, new_n17228_, new_n17229_,
    new_n17230_, new_n17231_, new_n17232_, new_n17233_, new_n17234_,
    new_n17235_, new_n17236_, new_n17237_, new_n17238_, new_n17239_,
    new_n17240_, new_n17241_, new_n17242_, new_n17243_, new_n17244_,
    new_n17245_, new_n17246_, new_n17247_, new_n17248_, new_n17249_,
    new_n17250_, new_n17251_, new_n17252_, new_n17253_, new_n17254_,
    new_n17255_, new_n17256_, new_n17257_, new_n17258_, new_n17259_,
    new_n17260_, new_n17261_, new_n17262_, new_n17263_, new_n17264_,
    new_n17265_, new_n17266_, new_n17267_, new_n17268_, new_n17269_,
    new_n17270_, new_n17271_, new_n17272_, new_n17273_, new_n17274_,
    new_n17275_, new_n17276_, new_n17277_, new_n17278_, new_n17279_,
    new_n17280_, new_n17281_, new_n17282_, new_n17283_, new_n17284_,
    new_n17285_, new_n17286_, new_n17287_, new_n17288_, new_n17289_,
    new_n17290_, new_n17291_, new_n17292_, new_n17293_, new_n17294_,
    new_n17295_, new_n17296_, new_n17297_, new_n17298_, new_n17299_,
    new_n17300_, new_n17301_, new_n17302_, new_n17303_, new_n17304_,
    new_n17305_, new_n17306_, new_n17307_, new_n17308_, new_n17309_,
    new_n17310_, new_n17311_, new_n17312_, new_n17313_, new_n17314_,
    new_n17315_, new_n17316_, new_n17317_, new_n17318_, new_n17319_,
    new_n17320_, new_n17321_, new_n17322_, new_n17323_, new_n17324_,
    new_n17325_, new_n17326_, new_n17327_, new_n17328_, new_n17329_,
    new_n17330_, new_n17331_, new_n17332_, new_n17333_, new_n17334_,
    new_n17335_, new_n17336_, new_n17337_, new_n17338_, new_n17339_,
    new_n17340_, new_n17341_, new_n17342_, new_n17343_, new_n17344_,
    new_n17345_, new_n17346_, new_n17347_, new_n17348_, new_n17349_,
    new_n17350_, new_n17351_, new_n17352_, new_n17353_, new_n17354_,
    new_n17355_, new_n17356_, new_n17357_, new_n17358_, new_n17359_,
    new_n17360_, new_n17361_, new_n17362_, new_n17363_, new_n17364_,
    new_n17365_, new_n17366_, new_n17367_, new_n17368_, new_n17369_,
    new_n17370_, new_n17371_, new_n17372_, new_n17373_, new_n17374_,
    new_n17375_, new_n17376_, new_n17377_, new_n17378_, new_n17379_,
    new_n17380_, new_n17381_, new_n17382_, new_n17383_, new_n17384_,
    new_n17385_, new_n17386_, new_n17387_, new_n17388_, new_n17389_,
    new_n17390_, new_n17391_, new_n17392_, new_n17393_, new_n17394_,
    new_n17395_, new_n17396_, new_n17397_, new_n17398_, new_n17399_,
    new_n17400_, new_n17401_, new_n17402_, new_n17403_, new_n17404_,
    new_n17405_, new_n17406_, new_n17407_, new_n17408_, new_n17409_,
    new_n17410_, new_n17411_, new_n17412_, new_n17413_, new_n17414_,
    new_n17415_, new_n17416_, new_n17417_, new_n17418_, new_n17419_,
    new_n17420_, new_n17421_, new_n17422_, new_n17423_, new_n17424_,
    new_n17425_, new_n17426_, new_n17427_, new_n17428_, new_n17429_,
    new_n17430_, new_n17431_, new_n17432_, new_n17433_, new_n17434_,
    new_n17435_, new_n17436_, new_n17437_, new_n17438_, new_n17439_,
    new_n17440_, new_n17441_, new_n17442_, new_n17443_, new_n17444_,
    new_n17445_, new_n17446_, new_n17447_, new_n17448_, new_n17449_,
    new_n17450_, new_n17451_, new_n17452_, new_n17453_, new_n17454_,
    new_n17455_, new_n17456_, new_n17457_, new_n17458_, new_n17459_,
    new_n17460_, new_n17461_, new_n17462_, new_n17463_, new_n17464_,
    new_n17465_, new_n17466_, new_n17467_, new_n17468_, new_n17469_,
    new_n17470_, new_n17471_, new_n17472_, new_n17473_, new_n17474_,
    new_n17475_, new_n17476_, new_n17477_, new_n17478_, new_n17479_,
    new_n17480_, new_n17481_, new_n17482_, new_n17483_, new_n17484_,
    new_n17485_, new_n17486_, new_n17487_, new_n17488_, new_n17489_,
    new_n17490_, new_n17491_, new_n17492_, new_n17493_, new_n17494_,
    new_n17495_, new_n17496_, new_n17497_, new_n17498_, new_n17499_,
    new_n17500_, new_n17501_, new_n17502_, new_n17503_, new_n17504_,
    new_n17505_, new_n17506_, new_n17507_, new_n17508_, new_n17509_,
    new_n17510_, new_n17511_, new_n17512_, new_n17513_, new_n17514_,
    new_n17515_, new_n17516_, new_n17517_, new_n17518_, new_n17519_,
    new_n17520_, new_n17521_, new_n17522_, new_n17523_, new_n17524_,
    new_n17525_, new_n17526_, new_n17527_, new_n17528_, new_n17529_,
    new_n17530_, new_n17531_, new_n17532_, new_n17533_, new_n17534_,
    new_n17535_, new_n17536_, new_n17537_, new_n17538_, new_n17539_,
    new_n17540_, new_n17541_, new_n17542_, new_n17543_, new_n17544_,
    new_n17545_, new_n17546_, new_n17547_, new_n17548_, new_n17549_,
    new_n17550_, new_n17551_, new_n17552_, new_n17553_, new_n17554_,
    new_n17555_, new_n17556_, new_n17557_, new_n17558_, new_n17559_,
    new_n17560_, new_n17561_, new_n17562_, new_n17563_, new_n17564_,
    new_n17565_, new_n17566_, new_n17567_, new_n17568_, new_n17569_,
    new_n17570_, new_n17571_, new_n17572_, new_n17573_, new_n17574_,
    new_n17575_, new_n17576_, new_n17577_, new_n17578_, new_n17579_,
    new_n17580_, new_n17581_, new_n17582_, new_n17583_, new_n17584_,
    new_n17585_, new_n17586_, new_n17587_, new_n17588_, new_n17589_,
    new_n17590_, new_n17591_, new_n17592_, new_n17593_, new_n17594_,
    new_n17595_, new_n17596_, new_n17597_, new_n17598_, new_n17599_,
    new_n17600_, new_n17601_, new_n17602_, new_n17603_, new_n17604_,
    new_n17605_, new_n17606_, new_n17607_, new_n17608_, new_n17609_,
    new_n17610_, new_n17611_, new_n17612_, new_n17613_, new_n17614_,
    new_n17615_, new_n17616_, new_n17617_, new_n17618_, new_n17619_,
    new_n17620_, new_n17621_, new_n17622_, new_n17623_, new_n17624_,
    new_n17625_, new_n17626_, new_n17627_, new_n17628_, new_n17629_,
    new_n17630_, new_n17631_, new_n17632_, new_n17633_, new_n17634_,
    new_n17635_, new_n17636_, new_n17637_, new_n17638_, new_n17639_,
    new_n17640_, new_n17641_, new_n17642_, new_n17643_, new_n17644_,
    new_n17645_, new_n17646_, new_n17647_, new_n17648_, new_n17649_,
    new_n17650_, new_n17651_, new_n17652_, new_n17653_, new_n17654_,
    new_n17655_, new_n17656_, new_n17657_, new_n17658_, new_n17659_,
    new_n17660_, new_n17661_, new_n17662_, new_n17663_, new_n17664_,
    new_n17665_, new_n17666_, new_n17667_, new_n17668_, new_n17669_,
    new_n17670_, new_n17671_, new_n17672_, new_n17673_, new_n17674_,
    new_n17675_, new_n17676_, new_n17677_, new_n17678_, new_n17679_,
    new_n17680_, new_n17681_, new_n17682_, new_n17683_, new_n17684_,
    new_n17685_, new_n17686_, new_n17687_, new_n17688_, new_n17689_,
    new_n17690_, new_n17691_, new_n17692_, new_n17693_, new_n17694_,
    new_n17695_, new_n17696_, new_n17697_, new_n17698_, new_n17699_,
    new_n17700_, new_n17701_, new_n17702_, new_n17703_, new_n17704_,
    new_n17705_, new_n17706_, new_n17707_, new_n17708_, new_n17709_,
    new_n17710_, new_n17711_, new_n17712_, new_n17713_, new_n17714_,
    new_n17715_, new_n17716_, new_n17717_, new_n17718_, new_n17719_,
    new_n17720_, new_n17721_, new_n17722_, new_n17723_, new_n17724_,
    new_n17725_, new_n17726_, new_n17727_, new_n17728_, new_n17729_,
    new_n17730_, new_n17731_, new_n17732_, new_n17733_, new_n17734_,
    new_n17735_, new_n17736_, new_n17737_, new_n17738_, new_n17739_,
    new_n17740_, new_n17741_, new_n17742_, new_n17743_, new_n17744_,
    new_n17745_, new_n17746_, new_n17747_, new_n17748_, new_n17749_,
    new_n17750_, new_n17751_, new_n17752_, new_n17753_, new_n17754_,
    new_n17755_, new_n17756_, new_n17757_, new_n17758_, new_n17759_,
    new_n17760_, new_n17761_, new_n17762_, new_n17763_, new_n17764_,
    new_n17765_, new_n17766_, new_n17767_, new_n17768_, new_n17769_,
    new_n17770_, new_n17771_, new_n17772_, new_n17773_, new_n17774_,
    new_n17775_, new_n17776_, new_n17777_, new_n17778_, new_n17779_,
    new_n17780_, new_n17781_, new_n17782_, new_n17783_, new_n17784_,
    new_n17785_, new_n17786_, new_n17787_, new_n17788_, new_n17789_,
    new_n17790_, new_n17791_, new_n17792_, new_n17793_, new_n17794_,
    new_n17795_, new_n17796_, new_n17797_, new_n17798_, new_n17799_,
    new_n17800_, new_n17801_, new_n17802_, new_n17803_, new_n17804_,
    new_n17805_, new_n17806_, new_n17807_, new_n17808_, new_n17809_,
    new_n17810_, new_n17811_, new_n17812_, new_n17813_, new_n17814_,
    new_n17815_, new_n17816_, new_n17817_, new_n17818_, new_n17819_,
    new_n17820_, new_n17821_, new_n17822_, new_n17823_, new_n17824_,
    new_n17825_, new_n17826_, new_n17827_, new_n17828_, new_n17829_,
    new_n17830_, new_n17831_, new_n17832_, new_n17833_, new_n17834_,
    new_n17835_, new_n17836_, new_n17837_, new_n17838_, new_n17839_,
    new_n17840_, new_n17841_, new_n17842_, new_n17843_, new_n17844_,
    new_n17845_, new_n17846_, new_n17847_, new_n17848_, new_n17849_,
    new_n17850_, new_n17851_, new_n17852_, new_n17853_, new_n17854_,
    new_n17855_, new_n17856_, new_n17857_, new_n17858_, new_n17859_,
    new_n17860_, new_n17861_, new_n17862_, new_n17863_, new_n17864_,
    new_n17865_, new_n17866_, new_n17867_, new_n17868_, new_n17869_,
    new_n17870_, new_n17871_, new_n17872_, new_n17873_, new_n17874_,
    new_n17875_, new_n17876_, new_n17877_, new_n17878_, new_n17879_,
    new_n17880_, new_n17881_, new_n17882_, new_n17883_, new_n17884_,
    new_n17885_, new_n17886_, new_n17887_, new_n17888_, new_n17889_,
    new_n17890_, new_n17891_, new_n17892_, new_n17893_, new_n17894_,
    new_n17895_, new_n17896_, new_n17897_, new_n17898_, new_n17899_,
    new_n17900_, new_n17901_, new_n17902_, new_n17903_, new_n17904_,
    new_n17905_, new_n17906_, new_n17907_, new_n17908_, new_n17909_,
    new_n17910_, new_n17911_, new_n17912_, new_n17913_, new_n17914_,
    new_n17915_, new_n17916_, new_n17917_, new_n17918_, new_n17919_,
    new_n17920_, new_n17921_, new_n17922_, new_n17923_, new_n17924_,
    new_n17925_, new_n17926_, new_n17927_, new_n17928_, new_n17929_,
    new_n17930_, new_n17931_, new_n17932_, new_n17933_, new_n17934_,
    new_n17935_, new_n17936_, new_n17937_, new_n17938_, new_n17939_,
    new_n17940_, new_n17941_, new_n17942_, new_n17943_, new_n17944_,
    new_n17945_, new_n17946_, new_n17947_, new_n17948_, new_n17949_,
    new_n17950_, new_n17951_, new_n17952_, new_n17953_, new_n17954_,
    new_n17955_, new_n17956_, new_n17957_, new_n17958_, new_n17959_,
    new_n17960_, new_n17961_, new_n17962_, new_n17963_, new_n17964_,
    new_n17965_, new_n17966_, new_n17967_, new_n17968_, new_n17969_,
    new_n17970_, new_n17971_, new_n17972_, new_n17973_, new_n17974_,
    new_n17975_, new_n17976_, new_n17977_, new_n17978_, new_n17979_,
    new_n17980_, new_n17981_, new_n17982_, new_n17983_, new_n17984_,
    new_n17985_, new_n17986_, new_n17987_, new_n17988_, new_n17989_,
    new_n17990_, new_n17991_, new_n17992_, new_n17993_, new_n17994_,
    new_n17995_, new_n17996_, new_n17997_, new_n17998_, new_n17999_,
    new_n18000_, new_n18001_, new_n18002_, new_n18003_, new_n18004_,
    new_n18005_, new_n18006_, new_n18007_, new_n18008_, new_n18009_,
    new_n18010_, new_n18011_, new_n18012_, new_n18013_, new_n18014_,
    new_n18015_, new_n18016_, new_n18017_, new_n18018_, new_n18019_,
    new_n18020_, new_n18021_, new_n18022_, new_n18023_, new_n18024_,
    new_n18025_, new_n18026_, new_n18027_, new_n18028_, new_n18029_,
    new_n18030_, new_n18031_, new_n18032_, new_n18033_, new_n18034_,
    new_n18035_, new_n18036_, new_n18037_, new_n18038_, new_n18039_,
    new_n18040_, new_n18041_, new_n18042_, new_n18043_, new_n18044_,
    new_n18045_, new_n18046_, new_n18047_, new_n18048_, new_n18049_,
    new_n18050_, new_n18051_, new_n18052_, new_n18053_, new_n18054_,
    new_n18055_, new_n18056_, new_n18057_, new_n18058_, new_n18059_,
    new_n18060_, new_n18061_, new_n18062_, new_n18063_, new_n18064_,
    new_n18065_, new_n18066_, new_n18067_, new_n18068_, new_n18069_,
    new_n18070_, new_n18071_, new_n18072_, new_n18073_, new_n18074_,
    new_n18075_, new_n18076_, new_n18077_, new_n18078_, new_n18079_,
    new_n18080_, new_n18081_, new_n18082_, new_n18083_, new_n18084_,
    new_n18085_, new_n18086_, new_n18087_, new_n18088_, new_n18089_,
    new_n18090_, new_n18091_, new_n18092_, new_n18093_, new_n18094_,
    new_n18095_, new_n18096_, new_n18097_, new_n18098_, new_n18099_,
    new_n18100_, new_n18101_, new_n18102_, new_n18103_, new_n18104_,
    new_n18105_, new_n18106_, new_n18107_, new_n18108_, new_n18109_,
    new_n18110_, new_n18111_, new_n18112_, new_n18113_, new_n18114_,
    new_n18115_, new_n18116_, new_n18117_, new_n18118_, new_n18119_,
    new_n18120_, new_n18121_, new_n18122_, new_n18123_, new_n18124_,
    new_n18125_, new_n18126_, new_n18127_, new_n18128_, new_n18129_,
    new_n18130_, new_n18131_, new_n18132_, new_n18133_, new_n18134_,
    new_n18135_, new_n18136_, new_n18137_, new_n18138_, new_n18139_,
    new_n18140_, new_n18141_, new_n18142_, new_n18143_, new_n18144_,
    new_n18145_, new_n18146_, new_n18147_, new_n18148_, new_n18149_,
    new_n18150_, new_n18151_, new_n18152_, new_n18153_, new_n18154_,
    new_n18155_, new_n18156_, new_n18157_, new_n18158_, new_n18159_,
    new_n18160_, new_n18161_, new_n18162_, new_n18163_, new_n18164_,
    new_n18165_, new_n18166_, new_n18167_, new_n18168_, new_n18169_,
    new_n18170_, new_n18171_, new_n18172_, new_n18173_, new_n18174_,
    new_n18175_, new_n18176_, new_n18177_, new_n18178_, new_n18179_,
    new_n18180_, new_n18181_, new_n18182_, new_n18183_, new_n18184_,
    new_n18185_, new_n18186_, new_n18187_, new_n18188_, new_n18189_,
    new_n18190_, new_n18191_, new_n18192_, new_n18193_, new_n18194_,
    new_n18195_, new_n18196_, new_n18197_, new_n18198_, new_n18199_,
    new_n18200_, new_n18201_, new_n18202_, new_n18203_, new_n18204_,
    new_n18205_, new_n18206_, new_n18207_, new_n18208_, new_n18209_,
    new_n18210_, new_n18211_, new_n18212_, new_n18213_, new_n18214_,
    new_n18215_, new_n18216_, new_n18217_, new_n18218_, new_n18219_,
    new_n18220_, new_n18221_, new_n18222_, new_n18223_, new_n18224_,
    new_n18225_, new_n18226_, new_n18227_, new_n18228_, new_n18229_,
    new_n18230_, new_n18231_, new_n18232_, new_n18233_, new_n18234_,
    new_n18235_, new_n18236_, new_n18237_, new_n18238_, new_n18239_,
    new_n18240_, new_n18241_, new_n18242_, new_n18243_, new_n18244_,
    new_n18245_, new_n18246_, new_n18247_, new_n18248_, new_n18249_,
    new_n18250_, new_n18251_, new_n18252_, new_n18253_, new_n18254_,
    new_n18255_, new_n18256_, new_n18257_, new_n18258_, new_n18259_,
    new_n18260_, new_n18261_, new_n18262_, new_n18263_, new_n18264_,
    new_n18265_, new_n18266_, new_n18267_, new_n18268_, new_n18269_,
    new_n18270_, new_n18271_, new_n18272_, new_n18273_, new_n18274_,
    new_n18275_, new_n18276_, new_n18277_, new_n18278_, new_n18279_,
    new_n18280_, new_n18281_, new_n18282_, new_n18283_, new_n18284_,
    new_n18285_, new_n18286_, new_n18287_, new_n18288_, new_n18289_,
    new_n18290_, new_n18291_, new_n18292_, new_n18293_, new_n18294_,
    new_n18295_, new_n18296_, new_n18297_, new_n18298_, new_n18299_,
    new_n18300_, new_n18301_, new_n18302_, new_n18303_, new_n18304_,
    new_n18305_, new_n18306_, new_n18307_, new_n18308_, new_n18309_,
    new_n18310_, new_n18311_, new_n18312_, new_n18313_, new_n18314_,
    new_n18315_, new_n18316_, new_n18317_, new_n18318_, new_n18319_,
    new_n18320_, new_n18321_, new_n18322_, new_n18323_, new_n18324_,
    new_n18325_, new_n18326_, new_n18327_, new_n18328_, new_n18329_,
    new_n18330_, new_n18331_, new_n18332_, new_n18333_, new_n18334_,
    new_n18335_, new_n18336_, new_n18337_, new_n18338_, new_n18339_,
    new_n18340_, new_n18341_, new_n18342_, new_n18343_, new_n18344_,
    new_n18345_, new_n18346_, new_n18347_, new_n18348_, new_n18349_,
    new_n18350_, new_n18351_, new_n18352_, new_n18353_, new_n18354_,
    new_n18355_, new_n18356_, new_n18357_, new_n18358_, new_n18359_,
    new_n18360_, new_n18361_, new_n18362_, new_n18363_, new_n18364_,
    new_n18365_, new_n18366_, new_n18367_, new_n18368_, new_n18369_,
    new_n18370_, new_n18371_, new_n18372_, new_n18373_, new_n18374_,
    new_n18375_, new_n18376_, new_n18377_, new_n18378_, new_n18379_,
    new_n18380_, new_n18381_, new_n18382_, new_n18383_, new_n18384_,
    new_n18385_, new_n18386_, new_n18387_, new_n18388_, new_n18389_,
    new_n18390_, new_n18391_, new_n18392_, new_n18393_, new_n18394_,
    new_n18395_, new_n18396_, new_n18397_, new_n18398_, new_n18399_,
    new_n18400_, new_n18401_, new_n18402_, new_n18403_, new_n18404_,
    new_n18405_, new_n18406_, new_n18407_, new_n18408_, new_n18409_,
    new_n18410_, new_n18411_, new_n18412_, new_n18413_, new_n18414_,
    new_n18415_, new_n18416_, new_n18417_, new_n18418_, new_n18419_,
    new_n18420_, new_n18421_, new_n18422_, new_n18423_, new_n18424_,
    new_n18425_, new_n18426_, new_n18427_, new_n18428_, new_n18429_,
    new_n18430_, new_n18431_, new_n18432_, new_n18433_, new_n18434_,
    new_n18435_, new_n18436_, new_n18437_, new_n18438_, new_n18439_,
    new_n18440_, new_n18441_, new_n18442_, new_n18443_, new_n18444_,
    new_n18445_, new_n18446_, new_n18447_, new_n18448_, new_n18449_,
    new_n18450_, new_n18451_, new_n18452_, new_n18453_, new_n18454_,
    new_n18455_, new_n18456_, new_n18457_, new_n18458_, new_n18459_,
    new_n18460_, new_n18461_, new_n18462_, new_n18463_, new_n18464_,
    new_n18465_, new_n18466_, new_n18467_, new_n18468_, new_n18469_,
    new_n18470_, new_n18471_, new_n18472_, new_n18473_, new_n18474_,
    new_n18475_, new_n18476_, new_n18477_, new_n18478_, new_n18479_,
    new_n18480_, new_n18481_, new_n18482_, new_n18483_, new_n18484_,
    new_n18485_, new_n18486_, new_n18487_, new_n18488_, new_n18489_,
    new_n18490_, new_n18491_, new_n18492_, new_n18493_, new_n18494_,
    new_n18495_, new_n18496_, new_n18497_, new_n18498_, new_n18499_,
    new_n18500_, new_n18501_, new_n18502_, new_n18503_, new_n18504_,
    new_n18505_, new_n18506_, new_n18507_, new_n18508_, new_n18509_,
    new_n18510_, new_n18511_, new_n18512_, new_n18513_, new_n18514_,
    new_n18515_, new_n18516_, new_n18517_, new_n18518_, new_n18519_,
    new_n18520_, new_n18521_, new_n18522_, new_n18523_, new_n18524_,
    new_n18525_, new_n18526_, new_n18527_, new_n18528_, new_n18529_,
    new_n18530_, new_n18531_, new_n18532_, new_n18533_, new_n18534_,
    new_n18535_, new_n18536_, new_n18537_, new_n18538_, new_n18539_,
    new_n18540_, new_n18541_, new_n18542_, new_n18543_, new_n18544_,
    new_n18545_, new_n18546_, new_n18547_, new_n18548_, new_n18549_,
    new_n18550_, new_n18551_, new_n18552_, new_n18553_, new_n18554_,
    new_n18555_, new_n18556_, new_n18557_, new_n18558_, new_n18559_,
    new_n18560_, new_n18561_, new_n18562_, new_n18563_, new_n18564_,
    new_n18565_, new_n18566_, new_n18567_, new_n18568_, new_n18569_,
    new_n18570_, new_n18571_, new_n18572_, new_n18573_, new_n18574_,
    new_n18575_, new_n18576_, new_n18577_, new_n18578_, new_n18579_,
    new_n18580_, new_n18581_, new_n18582_, new_n18583_, new_n18584_,
    new_n18585_, new_n18586_, new_n18587_, new_n18588_, new_n18589_,
    new_n18590_, new_n18591_, new_n18592_, new_n18593_, new_n18594_,
    new_n18595_, new_n18596_, new_n18597_, new_n18598_, new_n18599_,
    new_n18600_, new_n18601_, new_n18602_, new_n18603_, new_n18604_,
    new_n18605_, new_n18606_, new_n18607_, new_n18608_, new_n18609_,
    new_n18610_, new_n18611_, new_n18612_, new_n18613_, new_n18614_,
    new_n18615_, new_n18616_, new_n18617_, new_n18618_, new_n18619_,
    new_n18620_, new_n18621_, new_n18622_, new_n18623_, new_n18624_,
    new_n18625_, new_n18626_, new_n18627_, new_n18628_, new_n18629_,
    new_n18630_, new_n18631_, new_n18632_, new_n18633_, new_n18634_,
    new_n18635_, new_n18636_, new_n18637_, new_n18638_, new_n18639_,
    new_n18640_, new_n18641_, new_n18642_, new_n18643_, new_n18644_,
    new_n18645_, new_n18646_, new_n18647_, new_n18648_, new_n18649_,
    new_n18650_, new_n18651_, new_n18652_, new_n18653_, new_n18654_,
    new_n18655_, new_n18656_, new_n18657_, new_n18658_, new_n18659_,
    new_n18660_, new_n18661_, new_n18662_, new_n18663_, new_n18664_,
    new_n18665_, new_n18666_, new_n18667_, new_n18668_, new_n18669_,
    new_n18670_, new_n18671_, new_n18672_, new_n18673_, new_n18674_,
    new_n18675_, new_n18676_, new_n18677_, new_n18678_, new_n18679_,
    new_n18680_, new_n18681_, new_n18682_, new_n18683_, new_n18684_,
    new_n18685_, new_n18686_, new_n18687_, new_n18688_, new_n18689_,
    new_n18690_, new_n18691_, new_n18692_, new_n18693_, new_n18694_,
    new_n18695_, new_n18696_, new_n18697_, new_n18698_, new_n18699_,
    new_n18700_, new_n18701_, new_n18702_, new_n18703_, new_n18704_,
    new_n18705_, new_n18706_, new_n18707_, new_n18708_, new_n18709_,
    new_n18710_, new_n18711_, new_n18712_, new_n18713_, new_n18714_,
    new_n18715_, new_n18716_, new_n18717_, new_n18718_, new_n18719_,
    new_n18720_, new_n18721_, new_n18722_, new_n18723_, new_n18724_,
    new_n18725_, new_n18726_, new_n18727_, new_n18728_, new_n18729_,
    new_n18730_, new_n18731_, new_n18732_, new_n18733_, new_n18734_,
    new_n18735_, new_n18736_, new_n18737_, new_n18738_, new_n18739_,
    new_n18740_, new_n18741_, new_n18742_, new_n18743_, new_n18744_,
    new_n18745_, new_n18746_, new_n18747_, new_n18748_, new_n18749_,
    new_n18750_, new_n18751_, new_n18752_, new_n18753_, new_n18754_,
    new_n18755_, new_n18756_, new_n18757_, new_n18758_, new_n18759_,
    new_n18760_, new_n18761_, new_n18762_, new_n18763_, new_n18764_,
    new_n18765_, new_n18766_, new_n18767_, new_n18768_, new_n18769_,
    new_n18770_, new_n18771_, new_n18772_, new_n18773_, new_n18774_,
    new_n18775_, new_n18776_, new_n18777_, new_n18778_, new_n18779_,
    new_n18780_, new_n18781_, new_n18782_, new_n18783_, new_n18784_,
    new_n18785_, new_n18786_, new_n18787_, new_n18788_, new_n18789_,
    new_n18790_, new_n18791_, new_n18792_, new_n18793_, new_n18794_,
    new_n18795_, new_n18796_, new_n18797_, new_n18798_, new_n18799_,
    new_n18800_, new_n18801_, new_n18802_, new_n18803_, new_n18804_,
    new_n18805_, new_n18806_, new_n18807_, new_n18808_, new_n18809_,
    new_n18810_, new_n18811_, new_n18812_, new_n18813_, new_n18814_,
    new_n18815_, new_n18816_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18821_, new_n18822_, new_n18823_, new_n18824_,
    new_n18825_, new_n18826_, new_n18827_, new_n18828_, new_n18829_,
    new_n18830_, new_n18831_, new_n18832_, new_n18833_, new_n18834_,
    new_n18835_, new_n18836_, new_n18837_, new_n18838_, new_n18839_,
    new_n18840_, new_n18841_, new_n18842_, new_n18843_, new_n18844_,
    new_n18845_, new_n18846_, new_n18847_, new_n18848_, new_n18849_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18866_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18903_, new_n18904_,
    new_n18905_, new_n18906_, new_n18907_, new_n18908_, new_n18909_,
    new_n18910_, new_n18911_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18917_, new_n18918_, new_n18919_,
    new_n18920_, new_n18921_, new_n18922_, new_n18923_, new_n18924_,
    new_n18925_, new_n18926_, new_n18927_, new_n18928_, new_n18929_,
    new_n18930_, new_n18931_, new_n18932_, new_n18933_, new_n18934_,
    new_n18935_, new_n18936_, new_n18937_, new_n18938_, new_n18939_,
    new_n18940_, new_n18941_, new_n18942_, new_n18943_, new_n18944_,
    new_n18945_, new_n18946_, new_n18947_, new_n18948_, new_n18949_,
    new_n18950_, new_n18951_, new_n18952_, new_n18953_, new_n18954_,
    new_n18955_, new_n18956_, new_n18957_, new_n18958_, new_n18959_,
    new_n18960_, new_n18961_, new_n18962_, new_n18963_, new_n18964_,
    new_n18965_, new_n18966_, new_n18967_, new_n18968_, new_n18969_,
    new_n18970_, new_n18971_, new_n18972_, new_n18973_, new_n18974_,
    new_n18975_, new_n18976_, new_n18977_, new_n18978_, new_n18979_,
    new_n18980_, new_n18981_, new_n18982_, new_n18983_, new_n18984_,
    new_n18985_, new_n18986_, new_n18987_, new_n18988_, new_n18989_,
    new_n18990_, new_n18991_, new_n18992_, new_n18993_, new_n18994_,
    new_n18995_, new_n18996_, new_n18997_, new_n18998_, new_n18999_,
    new_n19000_, new_n19001_, new_n19002_, new_n19003_, new_n19004_,
    new_n19005_, new_n19006_, new_n19007_, new_n19008_, new_n19009_,
    new_n19010_, new_n19011_, new_n19012_, new_n19013_, new_n19014_,
    new_n19015_, new_n19016_, new_n19017_, new_n19018_, new_n19019_,
    new_n19020_, new_n19021_, new_n19022_, new_n19023_, new_n19024_,
    new_n19025_, new_n19026_, new_n19027_, new_n19028_, new_n19029_,
    new_n19030_, new_n19031_, new_n19032_, new_n19033_, new_n19034_,
    new_n19035_, new_n19036_, new_n19037_, new_n19038_, new_n19039_,
    new_n19040_, new_n19041_, new_n19042_, new_n19043_, new_n19044_,
    new_n19045_, new_n19046_, new_n19047_, new_n19048_, new_n19049_,
    new_n19050_, new_n19051_, new_n19052_, new_n19053_, new_n19054_,
    new_n19055_, new_n19056_, new_n19057_, new_n19058_, new_n19059_,
    new_n19060_, new_n19061_, new_n19062_, new_n19063_, new_n19064_,
    new_n19065_, new_n19066_, new_n19067_, new_n19068_, new_n19069_,
    new_n19070_, new_n19071_, new_n19072_, new_n19073_, new_n19074_,
    new_n19075_, new_n19076_, new_n19077_, new_n19078_, new_n19079_,
    new_n19080_, new_n19081_, new_n19082_, new_n19083_, new_n19084_,
    new_n19085_, new_n19086_, new_n19087_, new_n19088_, new_n19089_,
    new_n19090_, new_n19091_, new_n19092_, new_n19093_, new_n19094_,
    new_n19095_, new_n19096_, new_n19097_, new_n19098_, new_n19099_,
    new_n19100_, new_n19101_, new_n19102_, new_n19103_, new_n19104_,
    new_n19105_, new_n19106_, new_n19107_, new_n19108_, new_n19109_,
    new_n19110_, new_n19111_, new_n19112_, new_n19113_, new_n19114_,
    new_n19115_, new_n19116_, new_n19117_, new_n19118_, new_n19119_,
    new_n19120_, new_n19121_, new_n19122_, new_n19123_, new_n19124_,
    new_n19125_, new_n19126_, new_n19127_, new_n19128_, new_n19129_,
    new_n19130_, new_n19131_, new_n19132_, new_n19133_, new_n19134_,
    new_n19135_, new_n19136_, new_n19137_, new_n19138_, new_n19139_,
    new_n19140_, new_n19141_, new_n19142_, new_n19143_, new_n19144_,
    new_n19145_, new_n19146_, new_n19147_, new_n19148_, new_n19149_,
    new_n19150_, new_n19151_, new_n19152_, new_n19153_, new_n19154_,
    new_n19155_, new_n19156_, new_n19157_, new_n19158_, new_n19159_,
    new_n19160_, new_n19161_, new_n19162_, new_n19163_, new_n19164_,
    new_n19165_, new_n19166_, new_n19167_, new_n19168_, new_n19169_,
    new_n19170_, new_n19171_, new_n19172_, new_n19173_, new_n19174_,
    new_n19175_, new_n19176_, new_n19177_, new_n19178_, new_n19179_,
    new_n19180_, new_n19181_, new_n19182_, new_n19183_, new_n19184_,
    new_n19185_, new_n19186_, new_n19187_, new_n19188_, new_n19189_,
    new_n19190_, new_n19191_, new_n19192_, new_n19193_, new_n19194_,
    new_n19195_, new_n19196_, new_n19197_, new_n19198_, new_n19199_,
    new_n19200_, new_n19201_, new_n19202_, new_n19203_, new_n19204_,
    new_n19205_, new_n19206_, new_n19207_, new_n19208_, new_n19209_,
    new_n19210_, new_n19211_, new_n19212_, new_n19213_, new_n19214_,
    new_n19215_, new_n19216_, new_n19217_, new_n19218_, new_n19219_,
    new_n19220_, new_n19221_, new_n19222_, new_n19223_, new_n19224_,
    new_n19225_, new_n19226_, new_n19227_, new_n19228_, new_n19229_,
    new_n19230_, new_n19231_, new_n19232_, new_n19233_, new_n19234_,
    new_n19235_, new_n19236_, new_n19237_, new_n19238_, new_n19239_,
    new_n19240_, new_n19241_, new_n19242_, new_n19243_, new_n19244_,
    new_n19245_, new_n19246_, new_n19247_, new_n19248_, new_n19249_,
    new_n19250_, new_n19251_, new_n19252_, new_n19253_, new_n19254_,
    new_n19255_, new_n19256_, new_n19257_, new_n19258_, new_n19259_,
    new_n19260_, new_n19261_, new_n19262_, new_n19263_, new_n19264_,
    new_n19265_, new_n19266_, new_n19267_, new_n19268_, new_n19269_,
    new_n19270_, new_n19271_, new_n19272_, new_n19273_, new_n19274_,
    new_n19275_, new_n19276_, new_n19277_, new_n19278_, new_n19279_,
    new_n19280_, new_n19281_, new_n19282_, new_n19283_, new_n19284_,
    new_n19285_, new_n19286_, new_n19287_, new_n19288_, new_n19289_,
    new_n19290_, new_n19291_, new_n19292_, new_n19293_, new_n19294_,
    new_n19295_, new_n19296_, new_n19297_, new_n19298_, new_n19299_,
    new_n19300_, new_n19301_, new_n19302_, new_n19303_, new_n19304_,
    new_n19305_, new_n19306_, new_n19307_, new_n19308_, new_n19309_,
    new_n19310_, new_n19311_, new_n19312_, new_n19313_, new_n19314_,
    new_n19315_, new_n19316_, new_n19317_, new_n19318_, new_n19319_,
    new_n19320_, new_n19321_, new_n19322_, new_n19323_, new_n19324_,
    new_n19325_, new_n19326_, new_n19327_, new_n19328_, new_n19329_,
    new_n19330_, new_n19331_, new_n19332_, new_n19333_, new_n19334_,
    new_n19335_, new_n19336_, new_n19337_, new_n19338_, new_n19339_,
    new_n19340_, new_n19341_, new_n19342_, new_n19343_, new_n19344_,
    new_n19345_, new_n19346_, new_n19347_, new_n19348_, new_n19349_,
    new_n19350_, new_n19351_, new_n19352_, new_n19353_, new_n19354_,
    new_n19355_, new_n19356_, new_n19357_, new_n19358_, new_n19359_,
    new_n19360_, new_n19361_, new_n19362_, new_n19363_, new_n19364_,
    new_n19365_, new_n19366_, new_n19367_, new_n19368_, new_n19369_,
    new_n19370_, new_n19371_, new_n19372_, new_n19373_, new_n19374_,
    new_n19375_, new_n19376_, new_n19377_, new_n19378_, new_n19379_,
    new_n19380_, new_n19381_, new_n19382_, new_n19383_, new_n19384_,
    new_n19385_, new_n19386_, new_n19387_, new_n19388_, new_n19389_,
    new_n19390_, new_n19391_, new_n19392_, new_n19393_, new_n19394_,
    new_n19395_, new_n19396_, new_n19397_, new_n19398_, new_n19399_,
    new_n19400_, new_n19401_, new_n19402_, new_n19403_, new_n19404_,
    new_n19405_, new_n19406_, new_n19407_, new_n19408_, new_n19409_,
    new_n19410_, new_n19411_, new_n19412_, new_n19413_, new_n19414_,
    new_n19415_, new_n19416_, new_n19417_, new_n19418_, new_n19419_,
    new_n19420_, new_n19421_, new_n19422_, new_n19423_, new_n19424_,
    new_n19425_, new_n19426_, new_n19427_, new_n19428_, new_n19429_,
    new_n19430_, new_n19431_, new_n19432_, new_n19433_, new_n19434_,
    new_n19435_, new_n19436_, new_n19437_, new_n19438_, new_n19439_,
    new_n19440_, new_n19441_, new_n19442_, new_n19443_, new_n19444_,
    new_n19445_, new_n19446_, new_n19447_, new_n19448_, new_n19449_,
    new_n19450_, new_n19451_, new_n19452_, new_n19453_, new_n19454_,
    new_n19455_, new_n19456_, new_n19457_, new_n19458_, new_n19459_,
    new_n19460_, new_n19461_, new_n19462_, new_n19463_, new_n19464_,
    new_n19465_, new_n19466_, new_n19467_, new_n19468_, new_n19469_,
    new_n19470_, new_n19471_, new_n19472_, new_n19473_, new_n19474_,
    new_n19475_, new_n19476_, new_n19477_, new_n19478_, new_n19479_,
    new_n19480_, new_n19481_, new_n19482_, new_n19483_, new_n19484_,
    new_n19485_, new_n19486_, new_n19487_, new_n19488_, new_n19489_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19514_,
    new_n19515_, new_n19516_, new_n19517_, new_n19518_, new_n19519_,
    new_n19520_, new_n19521_, new_n19522_, new_n19523_, new_n19524_,
    new_n19525_, new_n19526_, new_n19527_, new_n19528_, new_n19529_,
    new_n19530_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19580_, new_n19581_,
    new_n19582_, new_n19583_, new_n19584_, new_n19585_, new_n19586_,
    new_n19587_, new_n19588_, new_n19589_, new_n19590_, new_n19591_,
    new_n19592_, new_n19593_, new_n19594_, new_n19595_, new_n19596_,
    new_n19597_, new_n19598_, new_n19599_, new_n19600_, new_n19601_,
    new_n19602_, new_n19603_, new_n19604_, new_n19605_, new_n19606_,
    new_n19607_, new_n19608_, new_n19609_, new_n19610_, new_n19611_,
    new_n19612_, new_n19613_, new_n19614_, new_n19615_, new_n19616_,
    new_n19617_, new_n19618_, new_n19619_, new_n19620_, new_n19621_,
    new_n19622_, new_n19623_, new_n19624_, new_n19625_, new_n19626_,
    new_n19627_, new_n19628_, new_n19629_, new_n19630_, new_n19631_,
    new_n19632_, new_n19633_, new_n19634_, new_n19635_, new_n19636_,
    new_n19637_, new_n19638_, new_n19639_, new_n19640_, new_n19641_,
    new_n19642_, new_n19643_, new_n19644_, new_n19645_, new_n19646_,
    new_n19647_, new_n19648_, new_n19649_, new_n19650_, new_n19651_,
    new_n19652_, new_n19653_, new_n19654_, new_n19655_, new_n19656_,
    new_n19657_, new_n19658_, new_n19659_, new_n19660_, new_n19661_,
    new_n19662_, new_n19663_, new_n19664_, new_n19665_, new_n19666_,
    new_n19667_, new_n19668_, new_n19669_, new_n19670_, new_n19671_,
    new_n19672_, new_n19673_, new_n19674_, new_n19675_, new_n19676_,
    new_n19677_, new_n19678_, new_n19679_, new_n19680_, new_n19681_,
    new_n19682_, new_n19683_, new_n19684_, new_n19685_, new_n19686_,
    new_n19687_, new_n19688_, new_n19689_, new_n19690_, new_n19691_,
    new_n19692_, new_n19693_, new_n19694_, new_n19695_, new_n19696_,
    new_n19697_, new_n19698_, new_n19699_, new_n19700_, new_n19701_,
    new_n19702_, new_n19703_, new_n19704_, new_n19705_, new_n19706_,
    new_n19707_, new_n19708_, new_n19709_, new_n19710_, new_n19711_,
    new_n19712_, new_n19713_, new_n19714_, new_n19715_, new_n19716_,
    new_n19717_, new_n19718_, new_n19719_, new_n19720_, new_n19721_,
    new_n19722_, new_n19723_, new_n19724_, new_n19725_, new_n19726_,
    new_n19727_, new_n19728_, new_n19729_, new_n19730_, new_n19731_,
    new_n19732_, new_n19733_, new_n19734_, new_n19735_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19804_, new_n19805_, new_n19806_,
    new_n19807_, new_n19808_, new_n19809_, new_n19810_, new_n19811_,
    new_n19812_, new_n19813_, new_n19814_, new_n19815_, new_n19816_,
    new_n19817_, new_n19818_, new_n19819_, new_n19820_, new_n19821_,
    new_n19822_, new_n19823_, new_n19824_, new_n19825_, new_n19826_,
    new_n19827_, new_n19828_, new_n19829_, new_n19830_, new_n19831_,
    new_n19832_, new_n19833_, new_n19834_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19840_, new_n19841_,
    new_n19842_, new_n19843_, new_n19844_, new_n19845_, new_n19846_,
    new_n19847_, new_n19848_, new_n19849_, new_n19850_, new_n19851_,
    new_n19852_, new_n19853_, new_n19854_, new_n19855_, new_n19856_,
    new_n19857_, new_n19858_, new_n19859_, new_n19860_, new_n19861_,
    new_n19862_, new_n19863_, new_n19864_, new_n19865_, new_n19866_,
    new_n19867_, new_n19868_, new_n19869_, new_n19870_, new_n19871_,
    new_n19872_, new_n19873_, new_n19874_, new_n19875_, new_n19876_,
    new_n19877_, new_n19878_, new_n19879_, new_n19880_, new_n19881_,
    new_n19882_, new_n19883_, new_n19884_, new_n19885_, new_n19886_,
    new_n19887_, new_n19888_, new_n19889_, new_n19890_, new_n19891_,
    new_n19892_, new_n19893_, new_n19894_, new_n19895_, new_n19896_,
    new_n19897_, new_n19898_, new_n19899_, new_n19900_, new_n19901_,
    new_n19902_, new_n19903_, new_n19904_, new_n19905_, new_n19906_,
    new_n19907_, new_n19908_, new_n19909_, new_n19910_, new_n19911_,
    new_n19912_, new_n19913_, new_n19914_, new_n19915_, new_n19916_,
    new_n19917_, new_n19918_, new_n19919_, new_n19920_, new_n19921_,
    new_n19922_, new_n19923_, new_n19924_, new_n19925_, new_n19926_,
    new_n19927_, new_n19928_, new_n19929_, new_n19930_, new_n19931_,
    new_n19932_, new_n19933_, new_n19934_, new_n19935_, new_n19936_,
    new_n19937_, new_n19938_, new_n19939_, new_n19940_, new_n19941_,
    new_n19942_, new_n19943_, new_n19944_, new_n19945_, new_n19946_,
    new_n19947_, new_n19948_, new_n19949_, new_n19950_, new_n19951_,
    new_n19952_, new_n19953_, new_n19954_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20127_, new_n20128_, new_n20129_, new_n20130_, new_n20131_,
    new_n20132_, new_n20133_, new_n20134_, new_n20135_, new_n20136_,
    new_n20137_, new_n20138_, new_n20139_, new_n20140_, new_n20141_,
    new_n20142_, new_n20143_, new_n20144_, new_n20145_, new_n20146_,
    new_n20147_, new_n20148_, new_n20149_, new_n20150_, new_n20151_,
    new_n20152_, new_n20153_, new_n20154_, new_n20155_, new_n20156_,
    new_n20157_, new_n20158_, new_n20159_, new_n20160_, new_n20161_,
    new_n20162_, new_n20163_, new_n20164_, new_n20165_, new_n20166_,
    new_n20167_, new_n20168_, new_n20169_, new_n20170_, new_n20171_,
    new_n20172_, new_n20173_, new_n20174_, new_n20175_, new_n20176_,
    new_n20177_, new_n20178_, new_n20179_, new_n20180_, new_n20181_,
    new_n20182_, new_n20183_, new_n20184_, new_n20185_, new_n20186_,
    new_n20187_, new_n20188_, new_n20189_, new_n20190_, new_n20191_,
    new_n20192_, new_n20193_, new_n20194_, new_n20195_, new_n20196_,
    new_n20197_, new_n20198_, new_n20199_, new_n20200_, new_n20201_,
    new_n20202_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20210_, new_n20211_,
    new_n20212_, new_n20213_, new_n20214_, new_n20215_, new_n20216_,
    new_n20217_, new_n20218_, new_n20219_, new_n20220_, new_n20221_,
    new_n20222_, new_n20223_, new_n20224_, new_n20225_, new_n20226_,
    new_n20227_, new_n20228_, new_n20229_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20282_, new_n20283_, new_n20284_, new_n20285_, new_n20286_,
    new_n20287_, new_n20288_, new_n20289_, new_n20290_, new_n20291_,
    new_n20292_, new_n20293_, new_n20294_, new_n20295_, new_n20296_,
    new_n20297_, new_n20298_, new_n20299_, new_n20300_, new_n20301_,
    new_n20302_, new_n20303_, new_n20304_, new_n20305_, new_n20306_,
    new_n20307_, new_n20308_, new_n20309_, new_n20310_, new_n20311_,
    new_n20312_, new_n20313_, new_n20314_, new_n20315_, new_n20316_,
    new_n20317_, new_n20318_, new_n20319_, new_n20320_, new_n20321_,
    new_n20322_, new_n20323_, new_n20324_, new_n20325_, new_n20326_,
    new_n20327_, new_n20328_, new_n20329_, new_n20330_, new_n20331_,
    new_n20332_, new_n20333_, new_n20334_, new_n20335_, new_n20336_,
    new_n20337_, new_n20338_, new_n20339_, new_n20340_, new_n20341_,
    new_n20342_, new_n20343_, new_n20344_, new_n20345_, new_n20346_,
    new_n20347_, new_n20348_, new_n20349_, new_n20350_, new_n20351_,
    new_n20352_, new_n20353_, new_n20354_, new_n20355_, new_n20356_,
    new_n20357_, new_n20358_, new_n20359_, new_n20360_, new_n20361_,
    new_n20362_, new_n20363_, new_n20364_, new_n20365_, new_n20366_,
    new_n20367_, new_n20368_, new_n20369_, new_n20370_, new_n20371_,
    new_n20372_, new_n20373_, new_n20374_, new_n20375_, new_n20376_,
    new_n20377_, new_n20378_, new_n20379_, new_n20380_, new_n20381_,
    new_n20382_, new_n20383_, new_n20384_, new_n20385_, new_n20386_,
    new_n20387_, new_n20388_, new_n20389_, new_n20390_, new_n20391_,
    new_n20392_, new_n20393_, new_n20394_, new_n20395_, new_n20396_,
    new_n20397_, new_n20398_, new_n20399_, new_n20400_, new_n20401_,
    new_n20402_, new_n20403_, new_n20404_, new_n20405_, new_n20406_,
    new_n20407_, new_n20408_, new_n20409_, new_n20410_, new_n20411_,
    new_n20412_, new_n20413_, new_n20414_, new_n20415_, new_n20416_,
    new_n20417_, new_n20418_, new_n20419_, new_n20420_, new_n20421_,
    new_n20422_, new_n20423_, new_n20424_, new_n20425_, new_n20426_,
    new_n20427_, new_n20428_, new_n20429_, new_n20430_, new_n20431_,
    new_n20432_, new_n20433_, new_n20434_, new_n20435_, new_n20436_,
    new_n20437_, new_n20438_, new_n20439_, new_n20440_, new_n20441_,
    new_n20442_, new_n20443_, new_n20444_, new_n20445_, new_n20446_,
    new_n20447_, new_n20448_, new_n20449_, new_n20450_, new_n20451_,
    new_n20452_, new_n20453_, new_n20454_, new_n20455_, new_n20456_,
    new_n20457_, new_n20458_, new_n20459_, new_n20460_, new_n20461_,
    new_n20462_, new_n20463_, new_n20464_, new_n20465_, new_n20466_,
    new_n20467_, new_n20468_, new_n20469_, new_n20470_, new_n20471_,
    new_n20472_, new_n20473_, new_n20474_, new_n20475_, new_n20476_,
    new_n20477_, new_n20478_, new_n20479_, new_n20480_, new_n20481_,
    new_n20482_, new_n20483_, new_n20484_, new_n20485_, new_n20486_,
    new_n20487_, new_n20488_, new_n20489_, new_n20490_, new_n20491_,
    new_n20492_, new_n20493_, new_n20494_, new_n20495_, new_n20496_,
    new_n20497_, new_n20498_, new_n20499_, new_n20500_, new_n20501_,
    new_n20502_, new_n20503_, new_n20504_, new_n20505_, new_n20506_,
    new_n20507_, new_n20508_, new_n20509_, new_n20510_, new_n20511_,
    new_n20512_, new_n20513_, new_n20514_, new_n20515_, new_n20516_,
    new_n20517_, new_n20518_, new_n20519_, new_n20520_, new_n20521_,
    new_n20522_, new_n20523_, new_n20524_, new_n20525_, new_n20526_,
    new_n20527_, new_n20528_, new_n20529_, new_n20530_, new_n20531_,
    new_n20532_, new_n20533_, new_n20534_, new_n20535_, new_n20536_,
    new_n20537_, new_n20538_, new_n20539_, new_n20540_, new_n20541_,
    new_n20542_, new_n20543_, new_n20544_, new_n20545_, new_n20546_,
    new_n20547_, new_n20548_, new_n20549_, new_n20550_, new_n20551_,
    new_n20552_, new_n20553_, new_n20554_, new_n20555_, new_n20556_,
    new_n20557_, new_n20558_, new_n20559_, new_n20560_, new_n20561_,
    new_n20562_, new_n20563_, new_n20564_, new_n20565_, new_n20566_,
    new_n20567_, new_n20568_, new_n20569_, new_n20570_, new_n20571_,
    new_n20572_, new_n20573_, new_n20574_, new_n20575_, new_n20576_,
    new_n20577_, new_n20578_, new_n20579_, new_n20580_, new_n20581_,
    new_n20582_, new_n20583_, new_n20584_, new_n20585_, new_n20586_,
    new_n20587_, new_n20588_, new_n20589_, new_n20590_, new_n20591_,
    new_n20592_, new_n20593_, new_n20594_, new_n20595_, new_n20596_,
    new_n20597_, new_n20598_, new_n20599_, new_n20600_, new_n20601_,
    new_n20602_, new_n20603_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20642_, new_n20643_, new_n20644_, new_n20645_, new_n20646_,
    new_n20647_, new_n20648_, new_n20649_, new_n20650_, new_n20651_,
    new_n20652_, new_n20653_, new_n20654_, new_n20655_, new_n20656_,
    new_n20657_, new_n20658_, new_n20659_, new_n20660_, new_n20661_,
    new_n20662_, new_n20663_, new_n20664_, new_n20665_, new_n20666_,
    new_n20667_, new_n20668_, new_n20669_, new_n20670_, new_n20671_,
    new_n20672_, new_n20673_, new_n20674_, new_n20675_, new_n20676_,
    new_n20677_, new_n20678_, new_n20679_, new_n20680_, new_n20681_,
    new_n20682_, new_n20683_, new_n20684_, new_n20685_, new_n20686_,
    new_n20687_, new_n20688_, new_n20689_, new_n20690_, new_n20691_,
    new_n20692_, new_n20693_, new_n20694_, new_n20695_, new_n20696_,
    new_n20697_, new_n20698_, new_n20699_, new_n20700_, new_n20701_,
    new_n20702_, new_n20703_, new_n20704_, new_n20705_, new_n20706_,
    new_n20707_, new_n20708_, new_n20709_, new_n20710_, new_n20711_,
    new_n20712_, new_n20713_, new_n20714_, new_n20715_, new_n20716_,
    new_n20717_, new_n20718_, new_n20719_, new_n20720_, new_n20721_,
    new_n20722_, new_n20723_, new_n20724_, new_n20725_, new_n20726_,
    new_n20727_, new_n20728_, new_n20729_, new_n20730_, new_n20731_,
    new_n20732_, new_n20733_, new_n20734_, new_n20735_, new_n20736_,
    new_n20737_, new_n20738_, new_n20739_, new_n20740_, new_n20741_,
    new_n20742_, new_n20743_, new_n20744_, new_n20745_, new_n20746_,
    new_n20747_, new_n20748_, new_n20749_, new_n20750_, new_n20751_,
    new_n20752_, new_n20753_, new_n20754_, new_n20755_, new_n20756_,
    new_n20757_, new_n20758_, new_n20759_, new_n20760_, new_n20761_,
    new_n20762_, new_n20763_, new_n20764_, new_n20765_, new_n20766_,
    new_n20767_, new_n20768_, new_n20769_, new_n20770_, new_n20771_,
    new_n20772_, new_n20773_, new_n20774_, new_n20775_, new_n20776_,
    new_n20777_, new_n20778_, new_n20779_, new_n20780_, new_n20781_,
    new_n20782_, new_n20783_, new_n20784_, new_n20785_, new_n20786_,
    new_n20787_, new_n20788_, new_n20789_, new_n20790_, new_n20791_,
    new_n20792_, new_n20793_, new_n20794_, new_n20795_, new_n20796_,
    new_n20797_, new_n20798_, new_n20799_, new_n20800_, new_n20801_,
    new_n20802_, new_n20803_, new_n20804_, new_n20805_, new_n20806_,
    new_n20807_, new_n20808_, new_n20809_, new_n20810_, new_n20811_,
    new_n20812_, new_n20813_, new_n20814_, new_n20815_, new_n20816_,
    new_n20817_, new_n20818_, new_n20819_, new_n20820_, new_n20821_,
    new_n20822_, new_n20823_, new_n20824_, new_n20825_, new_n20826_,
    new_n20827_, new_n20828_, new_n20829_, new_n20830_, new_n20831_,
    new_n20832_, new_n20833_, new_n20834_, new_n20835_, new_n20836_,
    new_n20837_, new_n20838_, new_n20839_, new_n20840_, new_n20841_,
    new_n20842_, new_n20843_, new_n20844_, new_n20845_, new_n20846_,
    new_n20847_, new_n20848_, new_n20849_, new_n20850_, new_n20851_,
    new_n20852_, new_n20853_, new_n20854_, new_n20855_, new_n20856_,
    new_n20857_, new_n20858_, new_n20859_, new_n20860_, new_n20861_,
    new_n20862_, new_n20863_, new_n20864_, new_n20865_, new_n20866_,
    new_n20867_, new_n20868_, new_n20869_, new_n20870_, new_n20871_,
    new_n20872_, new_n20873_, new_n20874_, new_n20875_, new_n20876_,
    new_n20877_, new_n20878_, new_n20879_, new_n20880_, new_n20881_,
    new_n20882_, new_n20883_, new_n20884_, new_n20885_, new_n20886_,
    new_n20887_, new_n20888_, new_n20889_, new_n20890_, new_n20891_,
    new_n20892_, new_n20893_, new_n20894_, new_n20895_, new_n20896_,
    new_n20897_, new_n20898_, new_n20899_, new_n20900_, new_n20901_,
    new_n20902_, new_n20903_, new_n20904_, new_n20905_, new_n20906_,
    new_n20907_, new_n20908_, new_n20909_, new_n20910_, new_n20911_,
    new_n20912_, new_n20913_, new_n20914_, new_n20915_, new_n20916_,
    new_n20917_, new_n20918_, new_n20919_, new_n20920_, new_n20921_,
    new_n20922_, new_n20923_, new_n20924_, new_n20925_, new_n20926_,
    new_n20927_, new_n20928_, new_n20929_, new_n20930_, new_n20931_,
    new_n20932_, new_n20933_, new_n20934_, new_n20935_, new_n20936_,
    new_n20937_, new_n20938_, new_n20939_, new_n20940_, new_n20941_,
    new_n20942_, new_n20943_, new_n20944_, new_n20945_, new_n20946_,
    new_n20947_, new_n20948_, new_n20949_, new_n20950_, new_n20951_,
    new_n20952_, new_n20953_, new_n20954_, new_n20955_, new_n20956_,
    new_n20957_, new_n20958_, new_n20959_, new_n20960_, new_n20961_,
    new_n20962_, new_n20963_, new_n20964_, new_n20965_, new_n20966_,
    new_n20967_, new_n20968_, new_n20969_, new_n20970_, new_n20971_,
    new_n20972_, new_n20973_, new_n20974_, new_n20975_, new_n20976_,
    new_n20977_, new_n20978_, new_n20979_, new_n20980_, new_n20981_,
    new_n20982_, new_n20983_, new_n20984_, new_n20985_, new_n20986_,
    new_n20987_, new_n20988_, new_n20989_, new_n20990_, new_n20991_,
    new_n20992_, new_n20993_, new_n20994_, new_n20995_, new_n20996_,
    new_n20997_, new_n20998_, new_n20999_, new_n21000_, new_n21001_,
    new_n21002_, new_n21003_, new_n21004_, new_n21005_, new_n21006_,
    new_n21007_, new_n21008_, new_n21009_, new_n21010_, new_n21011_,
    new_n21012_, new_n21013_, new_n21014_, new_n21015_, new_n21016_,
    new_n21017_, new_n21018_, new_n21019_, new_n21020_, new_n21021_,
    new_n21022_, new_n21023_, new_n21024_, new_n21025_, new_n21026_,
    new_n21027_, new_n21028_, new_n21029_, new_n21030_, new_n21031_,
    new_n21032_, new_n21033_, new_n21034_, new_n21035_, new_n21036_,
    new_n21037_, new_n21038_, new_n21039_, new_n21040_, new_n21041_,
    new_n21042_, new_n21043_, new_n21044_, new_n21045_, new_n21046_,
    new_n21047_, new_n21048_, new_n21049_, new_n21050_, new_n21051_,
    new_n21052_, new_n21053_, new_n21054_, new_n21055_, new_n21056_,
    new_n21057_, new_n21058_, new_n21059_, new_n21060_, new_n21061_,
    new_n21062_, new_n21063_, new_n21064_, new_n21065_, new_n21066_,
    new_n21067_, new_n21068_, new_n21069_, new_n21070_, new_n21071_,
    new_n21072_, new_n21073_, new_n21074_, new_n21075_, new_n21076_,
    new_n21077_, new_n21078_, new_n21079_, new_n21080_, new_n21081_,
    new_n21082_, new_n21083_, new_n21084_, new_n21085_, new_n21086_,
    new_n21087_, new_n21088_, new_n21089_, new_n21090_, new_n21091_,
    new_n21092_, new_n21093_, new_n21094_, new_n21095_, new_n21096_,
    new_n21097_, new_n21098_, new_n21099_, new_n21100_, new_n21101_,
    new_n21102_, new_n21103_, new_n21104_, new_n21105_, new_n21106_,
    new_n21107_, new_n21108_, new_n21109_, new_n21110_, new_n21111_,
    new_n21112_, new_n21113_, new_n21114_, new_n21115_, new_n21116_,
    new_n21117_, new_n21118_, new_n21119_, new_n21120_, new_n21121_,
    new_n21122_, new_n21123_, new_n21124_, new_n21125_, new_n21126_,
    new_n21127_, new_n21128_, new_n21129_, new_n21130_, new_n21131_,
    new_n21132_, new_n21133_, new_n21134_, new_n21135_, new_n21136_,
    new_n21137_, new_n21138_, new_n21139_, new_n21140_, new_n21141_,
    new_n21142_, new_n21143_, new_n21144_, new_n21145_, new_n21146_,
    new_n21147_, new_n21148_, new_n21149_, new_n21150_, new_n21151_,
    new_n21152_, new_n21153_, new_n21154_, new_n21155_, new_n21156_,
    new_n21157_, new_n21158_, new_n21159_, new_n21160_, new_n21161_,
    new_n21162_, new_n21163_, new_n21164_, new_n21165_, new_n21166_,
    new_n21167_, new_n21168_, new_n21169_, new_n21170_, new_n21171_,
    new_n21172_, new_n21173_, new_n21174_, new_n21175_, new_n21176_,
    new_n21177_, new_n21178_, new_n21179_, new_n21180_, new_n21181_,
    new_n21182_, new_n21183_, new_n21184_, new_n21185_, new_n21186_,
    new_n21187_, new_n21188_, new_n21189_, new_n21190_, new_n21191_,
    new_n21192_, new_n21193_, new_n21194_, new_n21195_, new_n21196_,
    new_n21197_, new_n21198_, new_n21199_, new_n21200_, new_n21201_,
    new_n21202_, new_n21203_, new_n21204_, new_n21205_, new_n21206_,
    new_n21207_, new_n21208_, new_n21209_, new_n21210_, new_n21211_,
    new_n21212_, new_n21213_, new_n21214_, new_n21215_, new_n21216_,
    new_n21217_, new_n21218_, new_n21219_, new_n21220_, new_n21221_,
    new_n21222_, new_n21223_, new_n21224_, new_n21225_, new_n21226_,
    new_n21227_, new_n21228_, new_n21229_, new_n21230_, new_n21231_,
    new_n21232_, new_n21233_, new_n21234_, new_n21235_, new_n21236_,
    new_n21237_, new_n21238_, new_n21239_, new_n21240_, new_n21241_,
    new_n21242_, new_n21243_, new_n21244_, new_n21245_, new_n21246_,
    new_n21247_, new_n21248_, new_n21249_, new_n21250_, new_n21251_,
    new_n21252_, new_n21253_, new_n21254_, new_n21255_, new_n21256_,
    new_n21257_, new_n21258_, new_n21259_, new_n21260_, new_n21261_,
    new_n21262_, new_n21263_, new_n21264_, new_n21265_, new_n21266_,
    new_n21267_, new_n21268_, new_n21269_, new_n21270_, new_n21271_,
    new_n21272_, new_n21273_, new_n21274_, new_n21275_, new_n21276_,
    new_n21277_, new_n21278_, new_n21279_, new_n21280_, new_n21281_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21297_, new_n21298_, new_n21299_, new_n21300_, new_n21301_,
    new_n21302_, new_n21303_, new_n21304_, new_n21305_, new_n21306_,
    new_n21307_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21332_, new_n21333_, new_n21334_, new_n21335_, new_n21336_,
    new_n21337_, new_n21338_, new_n21339_, new_n21340_, new_n21341_,
    new_n21342_, new_n21343_, new_n21344_, new_n21345_, new_n21346_,
    new_n21347_, new_n21348_, new_n21349_, new_n21350_, new_n21351_,
    new_n21352_, new_n21353_, new_n21354_, new_n21355_, new_n21356_,
    new_n21357_, new_n21358_, new_n21359_, new_n21360_, new_n21361_,
    new_n21362_, new_n21363_, new_n21364_, new_n21365_, new_n21366_,
    new_n21367_, new_n21368_, new_n21369_, new_n21370_, new_n21371_,
    new_n21372_, new_n21373_, new_n21374_, new_n21375_, new_n21376_,
    new_n21377_, new_n21378_, new_n21379_, new_n21380_, new_n21381_,
    new_n21382_, new_n21383_, new_n21384_, new_n21385_, new_n21386_,
    new_n21387_, new_n21388_, new_n21389_, new_n21390_, new_n21391_,
    new_n21392_, new_n21393_, new_n21394_, new_n21395_, new_n21396_,
    new_n21397_, new_n21398_, new_n21399_, new_n21400_, new_n21401_,
    new_n21402_, new_n21403_, new_n21404_, new_n21405_, new_n21406_,
    new_n21407_, new_n21408_, new_n21409_, new_n21410_, new_n21411_,
    new_n21412_, new_n21413_, new_n21414_, new_n21415_, new_n21416_,
    new_n21417_, new_n21418_, new_n21419_, new_n21420_, new_n21421_,
    new_n21422_, new_n21423_, new_n21424_, new_n21425_, new_n21426_,
    new_n21427_, new_n21428_, new_n21429_, new_n21430_, new_n21431_,
    new_n21432_, new_n21433_, new_n21434_, new_n21435_, new_n21436_,
    new_n21437_, new_n21438_, new_n21439_, new_n21440_, new_n21441_,
    new_n21442_, new_n21443_, new_n21444_, new_n21445_, new_n21446_,
    new_n21447_, new_n21448_, new_n21449_, new_n21450_, new_n21451_,
    new_n21452_, new_n21453_, new_n21454_, new_n21455_, new_n21456_,
    new_n21457_, new_n21458_, new_n21459_, new_n21460_, new_n21461_,
    new_n21462_, new_n21463_, new_n21464_, new_n21465_, new_n21466_,
    new_n21467_, new_n21468_, new_n21469_, new_n21470_, new_n21471_,
    new_n21472_, new_n21473_, new_n21474_, new_n21475_, new_n21476_,
    new_n21477_, new_n21478_, new_n21479_, new_n21480_, new_n21481_,
    new_n21482_, new_n21483_, new_n21484_, new_n21485_, new_n21486_,
    new_n21487_, new_n21488_, new_n21489_, new_n21490_, new_n21491_,
    new_n21492_, new_n21493_, new_n21494_, new_n21495_, new_n21496_,
    new_n21497_, new_n21498_, new_n21499_, new_n21500_, new_n21501_,
    new_n21502_, new_n21503_, new_n21504_, new_n21505_, new_n21506_,
    new_n21507_, new_n21508_, new_n21509_, new_n21510_, new_n21511_,
    new_n21512_, new_n21513_, new_n21514_, new_n21515_, new_n21516_,
    new_n21517_, new_n21518_, new_n21519_, new_n21520_, new_n21521_,
    new_n21522_, new_n21523_, new_n21524_, new_n21525_, new_n21526_,
    new_n21527_, new_n21528_, new_n21529_, new_n21530_, new_n21531_,
    new_n21532_, new_n21533_, new_n21534_, new_n21535_, new_n21536_,
    new_n21537_, new_n21538_, new_n21539_, new_n21540_, new_n21541_,
    new_n21542_, new_n21543_, new_n21544_, new_n21545_, new_n21546_,
    new_n21547_, new_n21548_, new_n21549_, new_n21550_, new_n21551_,
    new_n21552_, new_n21553_, new_n21554_, new_n21555_, new_n21556_,
    new_n21557_, new_n21558_, new_n21559_, new_n21560_, new_n21561_,
    new_n21562_, new_n21563_, new_n21564_, new_n21565_, new_n21566_,
    new_n21567_, new_n21568_, new_n21569_, new_n21570_, new_n21571_,
    new_n21572_, new_n21573_, new_n21574_, new_n21575_, new_n21576_,
    new_n21577_, new_n21578_, new_n21579_, new_n21580_, new_n21581_,
    new_n21582_, new_n21583_, new_n21584_, new_n21585_, new_n21586_,
    new_n21587_, new_n21588_, new_n21589_, new_n21590_, new_n21591_,
    new_n21592_, new_n21593_, new_n21594_, new_n21595_, new_n21596_,
    new_n21597_, new_n21598_, new_n21599_, new_n21600_, new_n21601_,
    new_n21602_, new_n21603_, new_n21604_, new_n21605_, new_n21606_,
    new_n21607_, new_n21608_, new_n21609_, new_n21610_, new_n21611_,
    new_n21612_, new_n21613_, new_n21614_, new_n21615_, new_n21616_,
    new_n21617_, new_n21618_, new_n21619_, new_n21620_, new_n21621_,
    new_n21622_, new_n21623_, new_n21624_, new_n21625_, new_n21626_,
    new_n21627_, new_n21628_, new_n21629_, new_n21630_, new_n21631_,
    new_n21632_, new_n21633_, new_n21634_, new_n21635_, new_n21636_,
    new_n21637_, new_n21638_, new_n21639_, new_n21640_, new_n21641_,
    new_n21642_, new_n21643_, new_n21644_, new_n21645_, new_n21646_,
    new_n21647_, new_n21648_, new_n21649_, new_n21650_, new_n21651_,
    new_n21652_, new_n21653_, new_n21654_, new_n21655_, new_n21656_,
    new_n21657_, new_n21658_, new_n21659_, new_n21660_, new_n21661_,
    new_n21662_, new_n21663_, new_n21664_, new_n21665_, new_n21666_,
    new_n21667_, new_n21668_, new_n21669_, new_n21670_, new_n21671_,
    new_n21672_, new_n21673_, new_n21674_, new_n21675_, new_n21676_,
    new_n21677_, new_n21678_, new_n21679_, new_n21680_, new_n21681_,
    new_n21682_, new_n21683_, new_n21684_, new_n21685_, new_n21686_,
    new_n21687_, new_n21688_, new_n21689_, new_n21690_, new_n21691_,
    new_n21692_, new_n21693_, new_n21694_, new_n21695_, new_n21696_,
    new_n21697_, new_n21698_, new_n21699_, new_n21700_, new_n21701_,
    new_n21702_, new_n21703_, new_n21704_, new_n21705_, new_n21706_,
    new_n21707_, new_n21708_, new_n21709_, new_n21710_, new_n21711_,
    new_n21712_, new_n21713_, new_n21714_, new_n21715_, new_n21716_,
    new_n21717_, new_n21718_, new_n21719_, new_n21720_, new_n21721_,
    new_n21722_, new_n21723_, new_n21724_, new_n21725_, new_n21726_,
    new_n21727_, new_n21728_, new_n21729_, new_n21730_, new_n21731_,
    new_n21732_, new_n21733_, new_n21734_, new_n21735_, new_n21736_,
    new_n21737_, new_n21738_, new_n21739_, new_n21740_, new_n21741_,
    new_n21742_, new_n21743_, new_n21744_, new_n21745_, new_n21746_,
    new_n21747_, new_n21748_, new_n21749_, new_n21750_, new_n21751_,
    new_n21752_, new_n21753_, new_n21754_, new_n21755_, new_n21756_,
    new_n21757_, new_n21758_, new_n21759_, new_n21760_, new_n21761_,
    new_n21762_, new_n21763_, new_n21764_, new_n21765_, new_n21766_,
    new_n21767_, new_n21768_, new_n21769_, new_n21770_, new_n21771_,
    new_n21772_, new_n21773_, new_n21774_, new_n21775_, new_n21776_,
    new_n21777_, new_n21778_, new_n21779_, new_n21780_, new_n21781_,
    new_n21782_, new_n21783_, new_n21784_, new_n21785_, new_n21786_,
    new_n21787_, new_n21788_, new_n21789_, new_n21790_, new_n21791_,
    new_n21792_, new_n21793_, new_n21794_, new_n21795_, new_n21796_,
    new_n21797_, new_n21798_, new_n21799_, new_n21800_, new_n21801_,
    new_n21802_, new_n21803_, new_n21804_, new_n21805_, new_n21806_,
    new_n21807_, new_n21808_, new_n21809_, new_n21810_, new_n21811_,
    new_n21812_, new_n21813_, new_n21814_, new_n21815_, new_n21816_,
    new_n21817_, new_n21818_, new_n21819_, new_n21820_, new_n21821_,
    new_n21822_, new_n21823_, new_n21824_, new_n21825_, new_n21826_,
    new_n21827_, new_n21828_, new_n21829_, new_n21830_, new_n21831_,
    new_n21832_, new_n21833_, new_n21834_, new_n21835_, new_n21836_,
    new_n21837_, new_n21838_, new_n21839_, new_n21840_, new_n21841_,
    new_n21842_, new_n21843_, new_n21844_, new_n21845_, new_n21846_,
    new_n21847_, new_n21848_, new_n21849_, new_n21850_, new_n21851_,
    new_n21852_, new_n21853_, new_n21854_, new_n21855_, new_n21856_,
    new_n21857_, new_n21858_, new_n21859_, new_n21860_, new_n21861_,
    new_n21862_, new_n21863_, new_n21864_, new_n21865_, new_n21866_,
    new_n21867_, new_n21868_, new_n21869_, new_n21870_, new_n21871_,
    new_n21872_, new_n21873_, new_n21874_, new_n21875_, new_n21876_,
    new_n21877_, new_n21878_, new_n21879_, new_n21880_, new_n21881_,
    new_n21882_, new_n21883_, new_n21884_, new_n21885_, new_n21886_,
    new_n21887_, new_n21888_, new_n21889_, new_n21890_, new_n21891_,
    new_n21892_, new_n21893_, new_n21894_, new_n21895_, new_n21896_,
    new_n21897_, new_n21898_, new_n21899_, new_n21900_, new_n21901_,
    new_n21902_, new_n21903_, new_n21904_, new_n21905_, new_n21906_,
    new_n21907_, new_n21908_, new_n21909_, new_n21910_, new_n21911_,
    new_n21912_, new_n21913_, new_n21914_, new_n21915_, new_n21916_,
    new_n21917_, new_n21918_, new_n21919_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21938_, new_n21939_, new_n21940_, new_n21941_,
    new_n21942_, new_n21943_, new_n21944_, new_n21945_, new_n21946_,
    new_n21947_, new_n21948_, new_n21949_, new_n21950_, new_n21951_,
    new_n21952_, new_n21953_, new_n21954_, new_n21955_, new_n21956_,
    new_n21957_, new_n21958_, new_n21959_, new_n21960_, new_n21961_,
    new_n21962_, new_n21963_, new_n21964_, new_n21965_, new_n21966_,
    new_n21967_, new_n21968_, new_n21969_, new_n21970_, new_n21971_,
    new_n21972_, new_n21973_, new_n21974_, new_n21975_, new_n21976_,
    new_n21977_, new_n21978_, new_n21979_, new_n21980_, new_n21981_,
    new_n21982_, new_n21983_, new_n21984_, new_n21985_, new_n21986_,
    new_n21987_, new_n21988_, new_n21989_, new_n21990_, new_n21991_,
    new_n21992_, new_n21993_, new_n21994_, new_n21995_, new_n21996_,
    new_n21997_, new_n21998_, new_n21999_, new_n22000_, new_n22001_,
    new_n22002_, new_n22003_, new_n22004_, new_n22005_, new_n22006_,
    new_n22007_, new_n22008_, new_n22009_, new_n22010_, new_n22011_,
    new_n22012_, new_n22013_, new_n22014_, new_n22015_, new_n22016_,
    new_n22017_, new_n22018_, new_n22019_, new_n22020_, new_n22021_,
    new_n22022_, new_n22023_, new_n22024_, new_n22025_, new_n22026_,
    new_n22027_, new_n22028_, new_n22029_, new_n22030_, new_n22031_,
    new_n22032_, new_n22033_, new_n22034_, new_n22035_, new_n22036_,
    new_n22037_, new_n22038_, new_n22039_, new_n22040_, new_n22041_,
    new_n22042_, new_n22043_, new_n22044_, new_n22045_, new_n22046_,
    new_n22047_, new_n22048_, new_n22049_, new_n22050_, new_n22051_,
    new_n22052_, new_n22053_, new_n22054_, new_n22055_, new_n22056_,
    new_n22057_, new_n22058_, new_n22059_, new_n22060_, new_n22061_,
    new_n22062_, new_n22063_, new_n22064_, new_n22065_, new_n22066_,
    new_n22067_, new_n22068_, new_n22069_, new_n22070_, new_n22071_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22079_, new_n22080_, new_n22081_,
    new_n22082_, new_n22083_, new_n22084_, new_n22085_, new_n22086_,
    new_n22087_, new_n22088_, new_n22089_, new_n22090_, new_n22091_,
    new_n22092_, new_n22093_, new_n22094_, new_n22095_, new_n22096_,
    new_n22097_, new_n22098_, new_n22099_, new_n22100_, new_n22101_,
    new_n22102_, new_n22103_, new_n22104_, new_n22105_, new_n22106_,
    new_n22107_, new_n22108_, new_n22109_, new_n22110_, new_n22111_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22119_, new_n22120_, new_n22121_,
    new_n22122_, new_n22123_, new_n22124_, new_n22125_, new_n22126_,
    new_n22127_, new_n22128_, new_n22129_, new_n22130_, new_n22131_,
    new_n22132_, new_n22133_, new_n22134_, new_n22135_, new_n22136_,
    new_n22137_, new_n22138_, new_n22139_, new_n22140_, new_n22141_,
    new_n22142_, new_n22143_, new_n22144_, new_n22145_, new_n22146_,
    new_n22147_, new_n22148_, new_n22149_, new_n22150_, new_n22151_,
    new_n22152_, new_n22153_, new_n22154_, new_n22155_, new_n22156_,
    new_n22157_, new_n22158_, new_n22159_, new_n22160_, new_n22161_,
    new_n22162_, new_n22163_, new_n22164_, new_n22165_, new_n22166_,
    new_n22167_, new_n22168_, new_n22169_, new_n22170_, new_n22171_,
    new_n22172_, new_n22173_, new_n22174_, new_n22175_, new_n22176_,
    new_n22177_, new_n22178_, new_n22179_, new_n22180_, new_n22181_,
    new_n22182_, new_n22183_, new_n22184_, new_n22185_, new_n22186_,
    new_n22187_, new_n22188_, new_n22189_, new_n22190_, new_n22191_,
    new_n22192_, new_n22193_, new_n22194_, new_n22195_, new_n22196_,
    new_n22197_, new_n22198_, new_n22199_, new_n22200_, new_n22201_,
    new_n22202_, new_n22203_, new_n22204_, new_n22205_, new_n22206_,
    new_n22207_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22226_,
    new_n22227_, new_n22228_, new_n22229_, new_n22230_, new_n22231_,
    new_n22232_, new_n22233_, new_n22234_, new_n22235_, new_n22236_,
    new_n22237_, new_n22238_, new_n22239_, new_n22240_, new_n22241_,
    new_n22242_, new_n22243_, new_n22244_, new_n22245_, new_n22246_,
    new_n22247_, new_n22248_, new_n22249_, new_n22250_, new_n22251_,
    new_n22252_, new_n22253_, new_n22254_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22261_,
    new_n22262_, new_n22263_, new_n22264_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22269_, new_n22270_, new_n22271_,
    new_n22272_, new_n22273_, new_n22274_, new_n22275_, new_n22276_,
    new_n22277_, new_n22278_, new_n22279_, new_n22280_, new_n22281_,
    new_n22282_, new_n22283_, new_n22284_, new_n22285_, new_n22286_,
    new_n22287_, new_n22288_, new_n22289_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22296_,
    new_n22297_, new_n22298_, new_n22299_, new_n22300_, new_n22301_,
    new_n22302_, new_n22303_, new_n22304_, new_n22305_, new_n22306_,
    new_n22307_, new_n22308_, new_n22309_, new_n22310_, new_n22311_,
    new_n22312_, new_n22313_, new_n22314_, new_n22315_, new_n22316_,
    new_n22317_, new_n22318_, new_n22319_, new_n22320_, new_n22321_,
    new_n22322_, new_n22323_, new_n22324_, new_n22325_, new_n22326_,
    new_n22327_, new_n22328_, new_n22329_, new_n22330_, new_n22331_,
    new_n22332_, new_n22333_, new_n22334_, new_n22335_, new_n22336_,
    new_n22337_, new_n22338_, new_n22339_, new_n22340_, new_n22341_,
    new_n22342_, new_n22343_, new_n22344_, new_n22345_, new_n22346_,
    new_n22347_, new_n22348_, new_n22349_, new_n22350_, new_n22351_,
    new_n22352_, new_n22353_, new_n22354_, new_n22355_, new_n22356_,
    new_n22357_, new_n22358_, new_n22359_, new_n22360_, new_n22361_,
    new_n22362_, new_n22363_, new_n22364_, new_n22365_, new_n22366_,
    new_n22367_, new_n22368_, new_n22369_, new_n22370_, new_n22371_,
    new_n22372_, new_n22373_, new_n22374_, new_n22375_, new_n22376_,
    new_n22377_, new_n22378_, new_n22379_, new_n22380_, new_n22381_,
    new_n22382_, new_n22383_, new_n22384_, new_n22385_, new_n22386_,
    new_n22387_, new_n22388_, new_n22389_, new_n22390_, new_n22391_,
    new_n22392_, new_n22393_, new_n22394_, new_n22395_, new_n22396_,
    new_n22397_, new_n22398_, new_n22399_, new_n22400_, new_n22401_,
    new_n22402_, new_n22403_, new_n22404_, new_n22405_, new_n22406_,
    new_n22407_, new_n22408_, new_n22409_, new_n22410_, new_n22411_,
    new_n22412_, new_n22413_, new_n22414_, new_n22415_, new_n22416_,
    new_n22417_, new_n22418_, new_n22419_, new_n22420_, new_n22421_,
    new_n22422_, new_n22423_, new_n22424_, new_n22425_, new_n22426_,
    new_n22427_, new_n22428_, new_n22429_, new_n22430_, new_n22431_,
    new_n22432_, new_n22433_, new_n22434_, new_n22435_, new_n22436_,
    new_n22437_, new_n22438_, new_n22439_, new_n22440_, new_n22441_,
    new_n22442_, new_n22443_, new_n22444_, new_n22445_, new_n22446_,
    new_n22447_, new_n22448_, new_n22449_, new_n22450_, new_n22451_,
    new_n22452_, new_n22453_, new_n22454_, new_n22455_, new_n22456_,
    new_n22457_, new_n22458_, new_n22459_, new_n22460_, new_n22461_,
    new_n22462_, new_n22463_, new_n22464_, new_n22465_, new_n22466_,
    new_n22467_, new_n22468_, new_n22469_, new_n22470_, new_n22471_,
    new_n22472_, new_n22473_, new_n22474_, new_n22475_, new_n22476_,
    new_n22477_, new_n22478_, new_n22479_, new_n22480_, new_n22481_,
    new_n22482_, new_n22483_, new_n22484_, new_n22485_, new_n22486_,
    new_n22487_, new_n22488_, new_n22489_, new_n22490_, new_n22491_,
    new_n22492_, new_n22493_, new_n22494_, new_n22495_, new_n22496_,
    new_n22497_, new_n22498_, new_n22499_, new_n22500_, new_n22501_,
    new_n22502_, new_n22503_, new_n22504_, new_n22505_, new_n22506_,
    new_n22507_, new_n22508_, new_n22509_, new_n22510_, new_n22511_,
    new_n22512_, new_n22513_, new_n22514_, new_n22515_, new_n22516_,
    new_n22517_, new_n22518_, new_n22519_, new_n22520_, new_n22521_,
    new_n22522_, new_n22523_, new_n22524_, new_n22525_, new_n22526_,
    new_n22527_, new_n22528_, new_n22529_, new_n22530_, new_n22531_,
    new_n22532_, new_n22533_, new_n22534_, new_n22535_, new_n22536_,
    new_n22537_, new_n22538_, new_n22539_, new_n22540_, new_n22541_,
    new_n22542_, new_n22543_, new_n22544_, new_n22545_, new_n22546_,
    new_n22547_, new_n22548_, new_n22549_, new_n22550_, new_n22551_,
    new_n22552_, new_n22553_, new_n22554_, new_n22555_, new_n22556_,
    new_n22557_, new_n22558_, new_n22559_, new_n22560_, new_n22561_,
    new_n22562_, new_n22563_, new_n22564_, new_n22565_, new_n22566_,
    new_n22567_, new_n22568_, new_n22569_, new_n22570_, new_n22571_,
    new_n22572_, new_n22573_, new_n22574_, new_n22575_, new_n22576_,
    new_n22577_, new_n22578_, new_n22579_, new_n22580_, new_n22581_,
    new_n22582_, new_n22583_, new_n22584_, new_n22585_, new_n22586_,
    new_n22587_, new_n22588_, new_n22589_, new_n22590_, new_n22591_,
    new_n22592_, new_n22593_, new_n22594_, new_n22595_, new_n22596_,
    new_n22597_, new_n22598_, new_n22599_, new_n22600_, new_n22601_,
    new_n22602_, new_n22603_, new_n22604_, new_n22605_, new_n22606_,
    new_n22607_, new_n22608_, new_n22609_, new_n22610_, new_n22611_,
    new_n22612_, new_n22613_, new_n22614_, new_n22615_, new_n22616_,
    new_n22617_, new_n22618_, new_n22619_, new_n22620_, new_n22621_,
    new_n22622_, new_n22623_, new_n22624_, new_n22625_, new_n22626_,
    new_n22627_, new_n22628_, new_n22629_, new_n22630_, new_n22631_,
    new_n22632_, new_n22633_, new_n22634_, new_n22635_, new_n22636_,
    new_n22637_, new_n22638_, new_n22639_, new_n22640_, new_n22641_,
    new_n22642_, new_n22643_, new_n22644_, new_n22645_, new_n22646_,
    new_n22647_, new_n22648_, new_n22649_, new_n22650_, new_n22651_,
    new_n22652_, new_n22653_, new_n22654_, new_n22655_, new_n22656_,
    new_n22657_, new_n22658_, new_n22659_, new_n22660_, new_n22661_,
    new_n22662_, new_n22663_, new_n22664_, new_n22665_, new_n22666_,
    new_n22667_, new_n22668_, new_n22669_, new_n22670_, new_n22671_,
    new_n22672_, new_n22673_, new_n22674_, new_n22675_, new_n22676_,
    new_n22677_, new_n22678_, new_n22679_, new_n22680_, new_n22681_,
    new_n22682_, new_n22683_, new_n22684_, new_n22685_, new_n22686_,
    new_n22687_, new_n22688_, new_n22689_, new_n22690_, new_n22691_,
    new_n22692_, new_n22693_, new_n22694_, new_n22695_, new_n22696_,
    new_n22697_, new_n22698_, new_n22699_, new_n22700_, new_n22701_,
    new_n22702_, new_n22703_, new_n22704_, new_n22705_, new_n22706_,
    new_n22707_, new_n22708_, new_n22709_, new_n22710_, new_n22711_,
    new_n22712_, new_n22713_, new_n22714_, new_n22715_, new_n22716_,
    new_n22717_, new_n22718_, new_n22719_, new_n22720_, new_n22721_,
    new_n22722_, new_n22723_, new_n22724_, new_n22725_, new_n22726_,
    new_n22727_, new_n22728_, new_n22729_, new_n22730_, new_n22731_,
    new_n22732_, new_n22733_, new_n22734_, new_n22735_, new_n22736_,
    new_n22737_, new_n22738_, new_n22739_, new_n22740_, new_n22741_,
    new_n22742_, new_n22743_, new_n22744_, new_n22745_, new_n22746_,
    new_n22747_, new_n22748_, new_n22749_, new_n22750_, new_n22751_,
    new_n22752_, new_n22753_, new_n22754_, new_n22755_, new_n22756_,
    new_n22757_, new_n22758_, new_n22759_, new_n22760_, new_n22761_,
    new_n22762_, new_n22763_, new_n22764_, new_n22765_, new_n22766_,
    new_n22767_, new_n22768_, new_n22769_, new_n22770_, new_n22771_,
    new_n22772_, new_n22773_, new_n22774_, new_n22775_, new_n22776_,
    new_n22777_, new_n22778_, new_n22779_, new_n22780_, new_n22781_,
    new_n22782_, new_n22783_, new_n22784_, new_n22785_, new_n22786_,
    new_n22787_, new_n22788_, new_n22789_, new_n22790_, new_n22791_,
    new_n22792_, new_n22793_, new_n22794_, new_n22795_, new_n22796_,
    new_n22797_, new_n22798_, new_n22799_, new_n22800_, new_n22801_,
    new_n22802_, new_n22803_, new_n22804_, new_n22805_, new_n22806_,
    new_n22807_, new_n22808_, new_n22809_, new_n22810_, new_n22811_,
    new_n22812_, new_n22813_, new_n22814_, new_n22815_, new_n22816_,
    new_n22817_, new_n22818_, new_n22819_, new_n22820_, new_n22821_,
    new_n22822_, new_n22823_, new_n22824_, new_n22825_, new_n22826_,
    new_n22827_, new_n22828_, new_n22829_, new_n22830_, new_n22831_,
    new_n22832_, new_n22833_, new_n22834_, new_n22835_, new_n22836_,
    new_n22837_, new_n22838_, new_n22839_, new_n22840_, new_n22841_,
    new_n22842_, new_n22843_, new_n22844_, new_n22845_, new_n22846_,
    new_n22847_, new_n22848_, new_n22849_, new_n22850_, new_n22851_,
    new_n22852_, new_n22853_, new_n22854_, new_n22855_, new_n22856_,
    new_n22857_, new_n22858_, new_n22859_, new_n22860_, new_n22861_,
    new_n22862_, new_n22863_, new_n22864_, new_n22865_, new_n22866_,
    new_n22867_, new_n22868_, new_n22869_, new_n22870_, new_n22871_,
    new_n22872_, new_n22873_, new_n22874_, new_n22875_, new_n22876_,
    new_n22877_, new_n22878_, new_n22879_, new_n22880_, new_n22881_,
    new_n22882_, new_n22883_, new_n22884_, new_n22885_, new_n22886_,
    new_n22887_, new_n22888_, new_n22889_, new_n22890_, new_n22891_,
    new_n22892_, new_n22893_, new_n22894_, new_n22895_, new_n22896_,
    new_n22897_, new_n22898_, new_n22899_, new_n22900_, new_n22901_,
    new_n22902_, new_n22903_, new_n22904_, new_n22905_, new_n22906_,
    new_n22907_, new_n22908_, new_n22909_, new_n22910_, new_n22911_,
    new_n22912_, new_n22913_, new_n22914_, new_n22915_, new_n22916_,
    new_n22917_, new_n22918_, new_n22919_, new_n22920_, new_n22921_,
    new_n22922_, new_n22923_, new_n22924_, new_n22925_, new_n22926_,
    new_n22927_, new_n22928_, new_n22929_, new_n22930_, new_n22931_,
    new_n22932_, new_n22933_, new_n22934_, new_n22935_, new_n22936_,
    new_n22937_, new_n22938_, new_n22939_, new_n22940_, new_n22941_,
    new_n22942_, new_n22943_, new_n22944_, new_n22945_, new_n22946_,
    new_n22947_, new_n22948_, new_n22949_, new_n22950_, new_n22951_,
    new_n22952_, new_n22953_, new_n22954_, new_n22955_, new_n22956_,
    new_n22957_, new_n22958_, new_n22959_, new_n22960_, new_n22961_,
    new_n22962_, new_n22963_, new_n22964_, new_n22965_, new_n22966_,
    new_n22967_, new_n22968_, new_n22969_, new_n22970_, new_n22971_,
    new_n22972_, new_n22973_, new_n22974_, new_n22975_, new_n22976_,
    new_n22977_, new_n22978_, new_n22979_, new_n22980_, new_n22981_,
    new_n22982_, new_n22983_, new_n22984_, new_n22985_, new_n22986_,
    new_n22987_, new_n22988_, new_n22989_, new_n22990_, new_n22991_,
    new_n22992_, new_n22993_, new_n22994_, new_n22995_, new_n22996_,
    new_n22997_, new_n22998_, new_n22999_, new_n23000_, new_n23001_,
    new_n23002_, new_n23003_, new_n23004_, new_n23005_, new_n23006_,
    new_n23007_, new_n23008_, new_n23009_, new_n23010_, new_n23011_,
    new_n23012_, new_n23013_, new_n23014_, new_n23015_, new_n23016_,
    new_n23017_, new_n23018_, new_n23019_, new_n23020_, new_n23021_,
    new_n23022_, new_n23023_, new_n23024_, new_n23025_, new_n23026_,
    new_n23027_, new_n23028_, new_n23029_, new_n23030_, new_n23031_,
    new_n23032_, new_n23033_, new_n23034_, new_n23035_, new_n23036_,
    new_n23037_, new_n23038_, new_n23039_, new_n23040_, new_n23041_,
    new_n23042_, new_n23043_, new_n23044_, new_n23045_, new_n23046_,
    new_n23047_, new_n23048_, new_n23049_, new_n23050_, new_n23051_,
    new_n23052_, new_n23053_, new_n23054_, new_n23055_, new_n23056_,
    new_n23057_, new_n23058_, new_n23059_, new_n23060_, new_n23061_,
    new_n23062_, new_n23063_, new_n23064_, new_n23065_, new_n23066_,
    new_n23067_, new_n23068_, new_n23069_, new_n23070_, new_n23071_,
    new_n23072_, new_n23073_, new_n23074_, new_n23075_, new_n23076_,
    new_n23077_, new_n23078_, new_n23079_, new_n23080_, new_n23081_,
    new_n23082_, new_n23083_, new_n23084_, new_n23085_, new_n23086_,
    new_n23087_, new_n23088_, new_n23089_, new_n23090_, new_n23091_,
    new_n23092_, new_n23093_, new_n23094_, new_n23095_, new_n23096_,
    new_n23097_, new_n23098_, new_n23099_, new_n23100_, new_n23101_,
    new_n23102_, new_n23103_, new_n23104_, new_n23105_, new_n23106_,
    new_n23107_, new_n23108_, new_n23109_, new_n23110_, new_n23111_,
    new_n23112_, new_n23113_, new_n23114_, new_n23115_, new_n23116_,
    new_n23117_, new_n23118_, new_n23119_, new_n23120_, new_n23121_,
    new_n23122_, new_n23123_, new_n23124_, new_n23125_, new_n23126_,
    new_n23127_, new_n23128_, new_n23129_, new_n23130_, new_n23131_,
    new_n23132_, new_n23133_, new_n23134_, new_n23135_, new_n23136_,
    new_n23137_, new_n23138_, new_n23139_, new_n23140_, new_n23141_,
    new_n23142_, new_n23143_, new_n23144_, new_n23145_, new_n23146_,
    new_n23147_, new_n23148_, new_n23149_, new_n23150_, new_n23151_,
    new_n23152_, new_n23153_, new_n23154_, new_n23155_, new_n23156_,
    new_n23157_, new_n23158_, new_n23159_, new_n23160_, new_n23161_,
    new_n23162_, new_n23163_, new_n23164_, new_n23165_, new_n23166_,
    new_n23167_, new_n23168_, new_n23169_, new_n23170_, new_n23171_,
    new_n23172_, new_n23173_, new_n23174_, new_n23175_, new_n23176_,
    new_n23177_, new_n23178_, new_n23179_, new_n23180_, new_n23181_,
    new_n23182_, new_n23183_, new_n23184_, new_n23185_, new_n23186_,
    new_n23187_, new_n23188_, new_n23189_, new_n23190_, new_n23191_,
    new_n23192_, new_n23193_, new_n23194_, new_n23195_, new_n23196_,
    new_n23197_, new_n23198_, new_n23199_, new_n23200_, new_n23201_,
    new_n23202_, new_n23203_, new_n23204_, new_n23205_, new_n23206_,
    new_n23207_, new_n23208_, new_n23209_, new_n23210_, new_n23211_,
    new_n23212_, new_n23213_, new_n23214_, new_n23215_, new_n23216_,
    new_n23217_, new_n23218_, new_n23219_, new_n23220_, new_n23221_,
    new_n23222_, new_n23223_, new_n23224_, new_n23225_, new_n23226_,
    new_n23227_, new_n23228_, new_n23229_, new_n23230_, new_n23231_,
    new_n23232_, new_n23233_, new_n23234_, new_n23235_, new_n23236_,
    new_n23237_, new_n23238_, new_n23239_, new_n23240_, new_n23241_,
    new_n23242_, new_n23243_, new_n23244_, new_n23245_, new_n23246_,
    new_n23247_, new_n23248_, new_n23249_, new_n23250_, new_n23251_,
    new_n23252_, new_n23253_, new_n23254_, new_n23255_, new_n23256_,
    new_n23257_, new_n23258_, new_n23259_, new_n23260_, new_n23261_,
    new_n23262_, new_n23263_, new_n23264_, new_n23265_, new_n23266_,
    new_n23267_, new_n23268_, new_n23269_, new_n23270_, new_n23271_,
    new_n23272_, new_n23273_, new_n23274_, new_n23275_, new_n23276_,
    new_n23277_, new_n23278_, new_n23279_, new_n23280_, new_n23281_,
    new_n23282_, new_n23283_, new_n23284_, new_n23285_, new_n23286_,
    new_n23287_, new_n23288_, new_n23289_, new_n23290_, new_n23291_,
    new_n23292_, new_n23293_, new_n23294_, new_n23295_, new_n23296_,
    new_n23297_, new_n23298_, new_n23299_, new_n23300_, new_n23301_,
    new_n23302_, new_n23303_, new_n23304_, new_n23305_, new_n23306_,
    new_n23307_, new_n23308_, new_n23309_, new_n23310_, new_n23311_,
    new_n23312_, new_n23313_, new_n23314_, new_n23315_, new_n23316_,
    new_n23317_, new_n23318_, new_n23319_, new_n23320_, new_n23321_,
    new_n23322_, new_n23323_, new_n23324_, new_n23325_, new_n23326_,
    new_n23327_, new_n23328_, new_n23329_, new_n23330_, new_n23331_,
    new_n23332_, new_n23333_, new_n23334_, new_n23335_, new_n23336_,
    new_n23337_, new_n23338_, new_n23339_, new_n23340_, new_n23341_,
    new_n23342_, new_n23343_, new_n23344_, new_n23345_, new_n23346_,
    new_n23347_, new_n23348_, new_n23349_, new_n23350_, new_n23351_,
    new_n23352_, new_n23353_, new_n23354_, new_n23355_, new_n23356_,
    new_n23357_, new_n23358_, new_n23359_, new_n23360_, new_n23361_,
    new_n23362_, new_n23363_, new_n23364_, new_n23365_, new_n23366_,
    new_n23367_, new_n23368_, new_n23369_, new_n23370_, new_n23371_,
    new_n23372_, new_n23373_, new_n23374_, new_n23375_, new_n23376_,
    new_n23377_, new_n23378_, new_n23379_, new_n23380_, new_n23381_,
    new_n23382_, new_n23383_, new_n23384_, new_n23385_, new_n23386_,
    new_n23387_, new_n23388_, new_n23389_, new_n23390_, new_n23391_,
    new_n23392_, new_n23393_, new_n23394_, new_n23395_, new_n23396_,
    new_n23397_, new_n23398_, new_n23399_, new_n23400_, new_n23401_,
    new_n23402_, new_n23403_, new_n23404_, new_n23405_, new_n23406_,
    new_n23407_, new_n23408_, new_n23409_, new_n23410_, new_n23411_,
    new_n23412_, new_n23413_, new_n23414_, new_n23415_, new_n23416_,
    new_n23417_, new_n23418_, new_n23419_, new_n23420_, new_n23421_,
    new_n23422_, new_n23423_, new_n23424_, new_n23425_, new_n23426_,
    new_n23427_, new_n23428_, new_n23429_, new_n23430_, new_n23431_,
    new_n23432_, new_n23433_, new_n23434_, new_n23435_, new_n23436_,
    new_n23437_, new_n23438_, new_n23439_, new_n23440_, new_n23441_,
    new_n23442_, new_n23443_, new_n23444_, new_n23445_, new_n23446_,
    new_n23447_, new_n23448_, new_n23449_, new_n23450_, new_n23451_,
    new_n23452_, new_n23453_, new_n23454_, new_n23455_, new_n23456_,
    new_n23457_, new_n23458_, new_n23459_, new_n23460_, new_n23461_,
    new_n23462_, new_n23463_, new_n23464_, new_n23465_, new_n23466_,
    new_n23467_, new_n23468_, new_n23469_, new_n23470_, new_n23471_,
    new_n23472_, new_n23473_, new_n23474_, new_n23475_, new_n23476_,
    new_n23477_, new_n23478_, new_n23479_, new_n23480_, new_n23481_,
    new_n23482_, new_n23483_, new_n23484_, new_n23485_, new_n23486_,
    new_n23487_, new_n23488_, new_n23489_, new_n23490_, new_n23491_,
    new_n23492_, new_n23493_, new_n23494_, new_n23495_, new_n23496_,
    new_n23497_, new_n23498_, new_n23499_, new_n23500_, new_n23501_,
    new_n23502_, new_n23503_, new_n23504_, new_n23505_, new_n23506_,
    new_n23507_, new_n23508_, new_n23509_, new_n23510_, new_n23511_,
    new_n23512_, new_n23513_, new_n23514_, new_n23515_, new_n23516_,
    new_n23517_, new_n23518_, new_n23519_, new_n23520_, new_n23521_,
    new_n23522_, new_n23523_, new_n23524_, new_n23525_, new_n23526_,
    new_n23527_, new_n23528_, new_n23529_, new_n23530_, new_n23531_,
    new_n23532_, new_n23533_, new_n23534_, new_n23535_, new_n23536_,
    new_n23537_, new_n23538_, new_n23539_, new_n23540_, new_n23541_,
    new_n23542_, new_n23543_, new_n23544_, new_n23545_, new_n23546_,
    new_n23547_, new_n23548_, new_n23549_, new_n23550_, new_n23551_,
    new_n23552_, new_n23553_, new_n23554_, new_n23555_, new_n23556_,
    new_n23557_, new_n23558_, new_n23559_, new_n23560_, new_n23561_,
    new_n23562_, new_n23563_, new_n23564_, new_n23565_, new_n23566_,
    new_n23567_, new_n23568_, new_n23569_, new_n23570_, new_n23571_,
    new_n23572_, new_n23573_, new_n23574_, new_n23575_, new_n23576_,
    new_n23577_, new_n23578_, new_n23579_, new_n23580_, new_n23581_,
    new_n23582_, new_n23583_, new_n23584_, new_n23585_, new_n23586_,
    new_n23587_, new_n23588_, new_n23589_, new_n23590_, new_n23591_,
    new_n23592_, new_n23593_, new_n23594_, new_n23595_, new_n23596_,
    new_n23597_, new_n23598_, new_n23599_, new_n23600_, new_n23601_,
    new_n23602_, new_n23603_, new_n23604_, new_n23605_, new_n23606_,
    new_n23607_, new_n23608_, new_n23609_, new_n23610_, new_n23611_,
    new_n23612_, new_n23613_, new_n23614_, new_n23615_, new_n23616_,
    new_n23617_, new_n23618_, new_n23619_, new_n23620_, new_n23621_,
    new_n23622_, new_n23623_, new_n23624_, new_n23625_, new_n23626_,
    new_n23627_, new_n23628_, new_n23629_, new_n23630_, new_n23631_,
    new_n23632_, new_n23633_, new_n23634_, new_n23635_, new_n23636_,
    new_n23637_, new_n23638_, new_n23639_, new_n23640_, new_n23641_,
    new_n23642_, new_n23643_, new_n23644_, new_n23645_, new_n23646_,
    new_n23647_, new_n23648_, new_n23649_, new_n23650_, new_n23651_,
    new_n23652_, new_n23653_, new_n23654_, new_n23655_, new_n23656_,
    new_n23657_, new_n23658_, new_n23659_, new_n23660_, new_n23661_,
    new_n23662_, new_n23663_, new_n23664_, new_n23665_, new_n23666_,
    new_n23667_, new_n23668_, new_n23669_, new_n23670_, new_n23671_,
    new_n23672_, new_n23673_, new_n23674_, new_n23675_, new_n23676_,
    new_n23677_, new_n23678_, new_n23679_, new_n23680_, new_n23681_,
    new_n23682_, new_n23683_, new_n23684_, new_n23685_, new_n23686_,
    new_n23687_, new_n23688_, new_n23689_, new_n23690_, new_n23691_,
    new_n23692_, new_n23693_, new_n23694_, new_n23695_, new_n23696_,
    new_n23697_, new_n23698_, new_n23699_, new_n23700_, new_n23701_,
    new_n23702_, new_n23703_, new_n23704_, new_n23705_, new_n23706_,
    new_n23707_, new_n23708_, new_n23709_, new_n23710_, new_n23711_,
    new_n23712_, new_n23713_, new_n23715_, new_n23716_, new_n23717_,
    new_n23718_, new_n23719_, new_n23720_, new_n23721_, new_n23722_,
    new_n23723_, new_n23724_, new_n23725_, new_n23726_, new_n23727_,
    new_n23728_, new_n23729_, new_n23730_, new_n23731_, new_n23732_,
    new_n23733_, new_n23734_, new_n23735_, new_n23736_, new_n23737_,
    new_n23738_, new_n23739_, new_n23740_, new_n23741_, new_n23742_,
    new_n23743_, new_n23744_, new_n23745_, new_n23746_, new_n23747_,
    new_n23748_, new_n23749_, new_n23750_, new_n23751_, new_n23752_,
    new_n23753_, new_n23754_, new_n23755_, new_n23756_, new_n23757_,
    new_n23758_, new_n23759_, new_n23760_, new_n23761_, new_n23762_,
    new_n23763_, new_n23764_, new_n23765_, new_n23766_, new_n23767_,
    new_n23768_, new_n23769_, new_n23770_, new_n23771_, new_n23772_,
    new_n23773_, new_n23774_, new_n23775_, new_n23776_, new_n23777_,
    new_n23778_, new_n23779_, new_n23780_, new_n23781_, new_n23782_,
    new_n23783_, new_n23784_, new_n23785_, new_n23786_, new_n23787_,
    new_n23788_, new_n23789_, new_n23790_, new_n23791_, new_n23792_,
    new_n23793_, new_n23794_, new_n23795_, new_n23796_, new_n23797_,
    new_n23798_, new_n23799_, new_n23800_, new_n23801_, new_n23802_,
    new_n23803_, new_n23804_, new_n23805_, new_n23806_, new_n23807_,
    new_n23808_, new_n23809_, new_n23810_, new_n23811_, new_n23812_,
    new_n23813_, new_n23814_, new_n23815_, new_n23816_, new_n23817_,
    new_n23818_, new_n23819_, new_n23820_, new_n23821_, new_n23822_,
    new_n23823_, new_n23824_, new_n23825_, new_n23826_, new_n23827_,
    new_n23828_, new_n23829_, new_n23830_, new_n23831_, new_n23832_,
    new_n23833_, new_n23834_, new_n23835_, new_n23836_, new_n23837_,
    new_n23838_, new_n23839_, new_n23840_, new_n23841_, new_n23842_,
    new_n23843_, new_n23844_, new_n23845_, new_n23846_, new_n23847_,
    new_n23848_, new_n23849_, new_n23850_, new_n23851_, new_n23852_,
    new_n23853_, new_n23854_, new_n23855_, new_n23856_, new_n23857_,
    new_n23858_, new_n23859_, new_n23860_, new_n23861_, new_n23862_,
    new_n23863_, new_n23864_, new_n23865_, new_n23866_, new_n23867_,
    new_n23868_, new_n23869_, new_n23870_, new_n23871_, new_n23872_,
    new_n23873_, new_n23874_, new_n23875_, new_n23876_, new_n23877_,
    new_n23878_, new_n23879_, new_n23880_, new_n23881_, new_n23882_,
    new_n23883_, new_n23884_, new_n23885_, new_n23886_, new_n23887_,
    new_n23888_, new_n23889_, new_n23890_, new_n23891_, new_n23892_,
    new_n23893_, new_n23894_, new_n23895_, new_n23896_, new_n23897_,
    new_n23898_, new_n23899_, new_n23900_, new_n23901_, new_n23902_,
    new_n23903_, new_n23904_, new_n23905_, new_n23906_, new_n23907_,
    new_n23908_, new_n23909_, new_n23910_, new_n23911_, new_n23912_,
    new_n23913_, new_n23914_, new_n23915_, new_n23916_, new_n23917_,
    new_n23918_, new_n23919_, new_n23920_, new_n23921_, new_n23922_,
    new_n23923_, new_n23924_, new_n23925_, new_n23926_, new_n23927_,
    new_n23928_, new_n23929_, new_n23930_, new_n23931_, new_n23932_,
    new_n23933_, new_n23934_, new_n23935_, new_n23936_, new_n23937_,
    new_n23938_, new_n23939_, new_n23940_, new_n23941_, new_n23942_,
    new_n23943_, new_n23944_, new_n23945_, new_n23946_, new_n23947_,
    new_n23948_, new_n23949_, new_n23950_, new_n23951_, new_n23952_,
    new_n23953_, new_n23954_, new_n23955_, new_n23956_, new_n23957_,
    new_n23958_, new_n23959_, new_n23960_, new_n23961_, new_n23962_,
    new_n23963_, new_n23964_, new_n23965_, new_n23966_, new_n23967_,
    new_n23968_, new_n23970_, new_n23971_, new_n23972_, new_n23973_,
    new_n23974_, new_n23975_, new_n23976_, new_n23977_, new_n23978_,
    new_n23979_, new_n23980_, new_n23981_, new_n23982_, new_n23983_,
    new_n23984_, new_n23985_, new_n23986_, new_n23987_, new_n23988_,
    new_n23989_, new_n23990_, new_n23991_, new_n23992_, new_n23993_,
    new_n23994_, new_n23995_, new_n23996_, new_n23997_, new_n23998_,
    new_n23999_, new_n24000_, new_n24001_, new_n24002_, new_n24003_,
    new_n24004_, new_n24005_, new_n24006_, new_n24007_, new_n24008_,
    new_n24009_, new_n24010_, new_n24011_, new_n24012_, new_n24013_,
    new_n24014_, new_n24015_, new_n24016_, new_n24017_, new_n24018_,
    new_n24019_, new_n24020_, new_n24021_, new_n24022_, new_n24023_,
    new_n24024_, new_n24025_, new_n24026_, new_n24027_, new_n24028_,
    new_n24029_, new_n24030_, new_n24031_, new_n24032_, new_n24033_,
    new_n24034_, new_n24035_, new_n24036_, new_n24037_, new_n24038_,
    new_n24039_, new_n24040_, new_n24041_, new_n24042_, new_n24043_,
    new_n24044_, new_n24045_, new_n24046_, new_n24047_, new_n24048_,
    new_n24049_, new_n24050_, new_n24051_, new_n24052_, new_n24053_,
    new_n24054_, new_n24055_, new_n24056_, new_n24057_, new_n24058_,
    new_n24059_, new_n24060_, new_n24061_, new_n24062_, new_n24063_,
    new_n24064_, new_n24065_, new_n24066_, new_n24067_, new_n24068_,
    new_n24069_, new_n24070_, new_n24071_, new_n24072_, new_n24073_,
    new_n24074_, new_n24075_, new_n24076_, new_n24077_, new_n24078_,
    new_n24079_, new_n24080_, new_n24081_, new_n24082_, new_n24083_,
    new_n24084_, new_n24085_, new_n24086_, new_n24087_, new_n24088_,
    new_n24089_, new_n24090_, new_n24091_, new_n24092_, new_n24093_,
    new_n24094_, new_n24095_, new_n24096_, new_n24097_, new_n24098_,
    new_n24099_, new_n24100_, new_n24101_, new_n24102_, new_n24103_,
    new_n24104_, new_n24105_, new_n24106_, new_n24107_, new_n24108_,
    new_n24109_, new_n24110_, new_n24111_, new_n24112_, new_n24113_,
    new_n24114_, new_n24115_, new_n24116_, new_n24117_, new_n24118_,
    new_n24119_, new_n24120_, new_n24121_, new_n24122_, new_n24123_,
    new_n24124_, new_n24125_, new_n24126_, new_n24127_, new_n24128_,
    new_n24129_, new_n24130_, new_n24131_, new_n24132_, new_n24133_,
    new_n24134_, new_n24135_, new_n24136_, new_n24137_, new_n24138_,
    new_n24139_, new_n24140_, new_n24141_, new_n24142_, new_n24143_,
    new_n24144_, new_n24145_, new_n24146_, new_n24147_, new_n24148_,
    new_n24149_, new_n24150_, new_n24151_, new_n24152_, new_n24153_,
    new_n24154_, new_n24155_, new_n24156_, new_n24157_, new_n24158_,
    new_n24159_, new_n24160_, new_n24161_, new_n24162_, new_n24163_,
    new_n24164_, new_n24165_, new_n24166_, new_n24167_, new_n24168_,
    new_n24169_, new_n24170_, new_n24171_, new_n24172_, new_n24173_,
    new_n24174_, new_n24175_, new_n24176_, new_n24177_, new_n24178_,
    new_n24179_, new_n24180_, new_n24181_, new_n24183_, new_n24184_,
    new_n24185_, new_n24186_, new_n24187_, new_n24188_, new_n24189_,
    new_n24190_, new_n24191_, new_n24192_, new_n24193_, new_n24194_,
    new_n24195_, new_n24196_, new_n24197_, new_n24198_, new_n24199_,
    new_n24200_, new_n24201_, new_n24202_, new_n24203_, new_n24204_,
    new_n24205_, new_n24206_, new_n24207_, new_n24208_, new_n24209_,
    new_n24210_, new_n24211_, new_n24212_, new_n24213_, new_n24214_,
    new_n24215_, new_n24216_, new_n24217_, new_n24218_, new_n24219_,
    new_n24220_, new_n24221_, new_n24222_, new_n24223_, new_n24224_,
    new_n24225_, new_n24226_, new_n24227_, new_n24228_, new_n24229_,
    new_n24230_, new_n24231_, new_n24232_, new_n24233_, new_n24234_,
    new_n24235_, new_n24236_, new_n24237_, new_n24238_, new_n24239_,
    new_n24240_, new_n24241_, new_n24242_, new_n24243_, new_n24244_,
    new_n24245_, new_n24246_, new_n24247_, new_n24248_, new_n24249_,
    new_n24250_, new_n24251_, new_n24252_, new_n24253_, new_n24254_,
    new_n24255_, new_n24256_, new_n24257_, new_n24258_, new_n24259_,
    new_n24260_, new_n24261_, new_n24262_, new_n24263_, new_n24264_,
    new_n24265_, new_n24266_, new_n24267_, new_n24268_, new_n24269_,
    new_n24270_, new_n24271_, new_n24272_, new_n24273_, new_n24274_,
    new_n24275_, new_n24276_, new_n24277_, new_n24278_, new_n24279_,
    new_n24280_, new_n24281_, new_n24282_, new_n24283_, new_n24284_,
    new_n24285_, new_n24286_, new_n24287_, new_n24288_, new_n24289_,
    new_n24290_, new_n24291_, new_n24292_, new_n24293_, new_n24294_,
    new_n24295_, new_n24296_, new_n24297_, new_n24298_, new_n24299_,
    new_n24300_, new_n24301_, new_n24302_, new_n24303_, new_n24304_,
    new_n24305_, new_n24306_, new_n24307_, new_n24308_, new_n24309_,
    new_n24310_, new_n24311_, new_n24312_, new_n24313_, new_n24314_,
    new_n24315_, new_n24316_, new_n24317_, new_n24318_, new_n24319_,
    new_n24320_, new_n24321_, new_n24322_, new_n24323_, new_n24324_,
    new_n24325_, new_n24326_, new_n24327_, new_n24328_, new_n24329_,
    new_n24330_, new_n24331_, new_n24332_, new_n24333_, new_n24334_,
    new_n24335_, new_n24336_, new_n24337_, new_n24338_, new_n24339_,
    new_n24340_, new_n24341_, new_n24342_, new_n24343_, new_n24344_,
    new_n24345_, new_n24346_, new_n24347_, new_n24348_, new_n24349_,
    new_n24350_, new_n24351_, new_n24352_, new_n24353_, new_n24354_,
    new_n24355_, new_n24356_, new_n24357_, new_n24358_, new_n24359_,
    new_n24360_, new_n24361_, new_n24362_, new_n24363_, new_n24364_,
    new_n24365_, new_n24366_, new_n24367_, new_n24368_, new_n24369_,
    new_n24370_, new_n24371_, new_n24372_, new_n24373_, new_n24374_,
    new_n24375_, new_n24376_, new_n24377_, new_n24378_, new_n24379_,
    new_n24380_, new_n24381_, new_n24382_, new_n24383_, new_n24384_,
    new_n24385_, new_n24386_, new_n24387_, new_n24388_, new_n24389_,
    new_n24390_, new_n24391_, new_n24392_, new_n24393_, new_n24394_,
    new_n24395_, new_n24396_, new_n24397_, new_n24398_, new_n24399_,
    new_n24400_, new_n24401_, new_n24403_, new_n24404_, new_n24405_,
    new_n24406_, new_n24407_, new_n24408_, new_n24409_, new_n24410_,
    new_n24411_, new_n24412_, new_n24413_, new_n24414_, new_n24415_,
    new_n24416_, new_n24417_, new_n24418_, new_n24419_, new_n24420_,
    new_n24421_, new_n24422_, new_n24423_, new_n24424_, new_n24425_,
    new_n24426_, new_n24427_, new_n24428_, new_n24429_, new_n24430_,
    new_n24431_, new_n24432_, new_n24433_, new_n24434_, new_n24435_,
    new_n24436_, new_n24437_, new_n24438_, new_n24439_, new_n24440_,
    new_n24441_, new_n24442_, new_n24443_, new_n24444_, new_n24445_,
    new_n24446_, new_n24447_, new_n24448_, new_n24449_, new_n24450_,
    new_n24451_, new_n24452_, new_n24453_, new_n24454_, new_n24455_,
    new_n24456_, new_n24457_, new_n24458_, new_n24459_, new_n24460_,
    new_n24461_, new_n24462_, new_n24463_, new_n24464_, new_n24465_,
    new_n24466_, new_n24467_, new_n24468_, new_n24469_, new_n24470_,
    new_n24471_, new_n24472_, new_n24473_, new_n24474_, new_n24475_,
    new_n24476_, new_n24477_, new_n24478_, new_n24479_, new_n24480_,
    new_n24481_, new_n24482_, new_n24483_, new_n24484_, new_n24485_,
    new_n24486_, new_n24487_, new_n24488_, new_n24489_, new_n24490_,
    new_n24491_, new_n24492_, new_n24493_, new_n24494_, new_n24495_,
    new_n24496_, new_n24497_, new_n24498_, new_n24499_, new_n24500_,
    new_n24501_, new_n24502_, new_n24503_, new_n24504_, new_n24505_,
    new_n24506_, new_n24507_, new_n24508_, new_n24509_, new_n24510_,
    new_n24511_, new_n24512_, new_n24513_, new_n24514_, new_n24515_,
    new_n24516_, new_n24517_, new_n24518_, new_n24519_, new_n24520_,
    new_n24521_, new_n24522_, new_n24523_, new_n24524_, new_n24525_,
    new_n24526_, new_n24527_, new_n24528_, new_n24529_, new_n24530_,
    new_n24531_, new_n24532_, new_n24533_, new_n24534_, new_n24535_,
    new_n24536_, new_n24537_, new_n24538_, new_n24539_, new_n24540_,
    new_n24541_, new_n24542_, new_n24543_, new_n24544_, new_n24545_,
    new_n24546_, new_n24547_, new_n24548_, new_n24549_, new_n24550_,
    new_n24551_, new_n24552_, new_n24553_, new_n24554_, new_n24555_,
    new_n24556_, new_n24557_, new_n24558_, new_n24559_, new_n24560_,
    new_n24561_, new_n24562_, new_n24563_, new_n24564_, new_n24565_,
    new_n24566_, new_n24567_, new_n24568_, new_n24569_, new_n24570_,
    new_n24571_, new_n24572_, new_n24573_, new_n24574_, new_n24575_,
    new_n24576_, new_n24577_, new_n24578_, new_n24579_, new_n24580_,
    new_n24581_, new_n24582_, new_n24583_, new_n24584_, new_n24585_,
    new_n24586_, new_n24587_, new_n24588_, new_n24589_, new_n24590_,
    new_n24591_, new_n24592_, new_n24593_, new_n24594_, new_n24595_,
    new_n24596_, new_n24597_, new_n24598_, new_n24599_, new_n24600_,
    new_n24601_, new_n24602_, new_n24603_, new_n24604_, new_n24605_,
    new_n24606_, new_n24607_, new_n24608_, new_n24609_, new_n24610_,
    new_n24611_, new_n24612_, new_n24613_, new_n24614_, new_n24615_,
    new_n24616_, new_n24617_, new_n24618_, new_n24619_, new_n24620_,
    new_n24621_, new_n24622_, new_n24623_, new_n24624_, new_n24625_,
    new_n24626_, new_n24627_, new_n24628_, new_n24629_, new_n24630_,
    new_n24631_, new_n24632_, new_n24633_, new_n24634_, new_n24635_,
    new_n24636_, new_n24638_, new_n24639_, new_n24640_, new_n24641_,
    new_n24642_, new_n24643_, new_n24644_, new_n24645_, new_n24646_,
    new_n24647_, new_n24648_, new_n24649_, new_n24650_, new_n24651_,
    new_n24652_, new_n24653_, new_n24654_, new_n24655_, new_n24656_,
    new_n24657_, new_n24658_, new_n24659_, new_n24660_, new_n24661_,
    new_n24662_, new_n24663_, new_n24664_, new_n24665_, new_n24666_,
    new_n24667_, new_n24668_, new_n24669_, new_n24670_, new_n24671_,
    new_n24672_, new_n24673_, new_n24674_, new_n24675_, new_n24676_,
    new_n24677_, new_n24678_, new_n24679_, new_n24680_, new_n24681_,
    new_n24682_, new_n24683_, new_n24684_, new_n24685_, new_n24686_,
    new_n24687_, new_n24688_, new_n24689_, new_n24690_, new_n24691_,
    new_n24692_, new_n24693_, new_n24694_, new_n24695_, new_n24696_,
    new_n24697_, new_n24698_, new_n24699_, new_n24700_, new_n24701_,
    new_n24702_, new_n24703_, new_n24704_, new_n24705_, new_n24706_,
    new_n24707_, new_n24708_, new_n24709_, new_n24710_, new_n24711_,
    new_n24712_, new_n24713_, new_n24714_, new_n24715_, new_n24716_,
    new_n24717_, new_n24718_, new_n24719_, new_n24720_, new_n24721_,
    new_n24722_, new_n24723_, new_n24724_, new_n24725_, new_n24726_,
    new_n24727_, new_n24728_, new_n24729_, new_n24730_, new_n24731_,
    new_n24732_, new_n24733_, new_n24734_, new_n24735_, new_n24736_,
    new_n24737_, new_n24738_, new_n24739_, new_n24740_, new_n24741_,
    new_n24742_, new_n24743_, new_n24744_, new_n24745_, new_n24746_,
    new_n24747_, new_n24748_, new_n24749_, new_n24750_, new_n24751_,
    new_n24752_, new_n24753_, new_n24754_, new_n24755_, new_n24756_,
    new_n24757_, new_n24758_, new_n24759_, new_n24760_, new_n24761_,
    new_n24762_, new_n24763_, new_n24764_, new_n24765_, new_n24766_,
    new_n24767_, new_n24768_, new_n24769_, new_n24770_, new_n24771_,
    new_n24772_, new_n24773_, new_n24774_, new_n24775_, new_n24776_,
    new_n24777_, new_n24778_, new_n24779_, new_n24780_, new_n24781_,
    new_n24782_, new_n24783_, new_n24784_, new_n24785_, new_n24786_,
    new_n24787_, new_n24788_, new_n24789_, new_n24790_, new_n24791_,
    new_n24792_, new_n24793_, new_n24794_, new_n24795_, new_n24796_,
    new_n24797_, new_n24798_, new_n24799_, new_n24800_, new_n24801_,
    new_n24802_, new_n24803_, new_n24804_, new_n24805_, new_n24806_,
    new_n24807_, new_n24808_, new_n24809_, new_n24810_, new_n24811_,
    new_n24812_, new_n24813_, new_n24814_, new_n24815_, new_n24816_,
    new_n24817_, new_n24818_, new_n24819_, new_n24820_, new_n24821_,
    new_n24822_, new_n24823_, new_n24824_, new_n24825_, new_n24826_,
    new_n24827_, new_n24828_, new_n24829_, new_n24830_, new_n24831_,
    new_n24832_, new_n24833_, new_n24834_, new_n24835_, new_n24836_,
    new_n24837_, new_n24838_, new_n24839_, new_n24840_, new_n24841_,
    new_n24842_, new_n24843_, new_n24844_, new_n24846_, new_n24847_,
    new_n24848_, new_n24849_, new_n24850_, new_n24851_, new_n24852_,
    new_n24853_, new_n24854_, new_n24855_, new_n24856_, new_n24857_,
    new_n24858_, new_n24859_, new_n24860_, new_n24861_, new_n24862_,
    new_n24863_, new_n24864_, new_n24865_, new_n24866_, new_n24867_,
    new_n24868_, new_n24869_, new_n24870_, new_n24871_, new_n24872_,
    new_n24873_, new_n24874_, new_n24875_, new_n24876_, new_n24877_,
    new_n24878_, new_n24879_, new_n24880_, new_n24881_, new_n24882_,
    new_n24883_, new_n24884_, new_n24885_, new_n24886_, new_n24887_,
    new_n24888_, new_n24889_, new_n24890_, new_n24891_, new_n24892_,
    new_n24893_, new_n24894_, new_n24895_, new_n24896_, new_n24897_,
    new_n24898_, new_n24899_, new_n24900_, new_n24901_, new_n24902_,
    new_n24903_, new_n24904_, new_n24905_, new_n24906_, new_n24907_,
    new_n24908_, new_n24909_, new_n24910_, new_n24911_, new_n24912_,
    new_n24913_, new_n24914_, new_n24915_, new_n24916_, new_n24917_,
    new_n24918_, new_n24919_, new_n24920_, new_n24921_, new_n24922_,
    new_n24923_, new_n24924_, new_n24925_, new_n24926_, new_n24927_,
    new_n24928_, new_n24929_, new_n24930_, new_n24931_, new_n24932_,
    new_n24933_, new_n24934_, new_n24935_, new_n24936_, new_n24937_,
    new_n24938_, new_n24939_, new_n24940_, new_n24941_, new_n24942_,
    new_n24943_, new_n24944_, new_n24945_, new_n24946_, new_n24947_,
    new_n24948_, new_n24949_, new_n24950_, new_n24951_, new_n24952_,
    new_n24953_, new_n24954_, new_n24955_, new_n24956_, new_n24957_,
    new_n24958_, new_n24959_, new_n24960_, new_n24961_, new_n24962_,
    new_n24963_, new_n24964_, new_n24965_, new_n24966_, new_n24967_,
    new_n24968_, new_n24969_, new_n24970_, new_n24971_, new_n24972_,
    new_n24973_, new_n24974_, new_n24975_, new_n24976_, new_n24977_,
    new_n24978_, new_n24979_, new_n24980_, new_n24981_, new_n24982_,
    new_n24983_, new_n24984_, new_n24985_, new_n24986_, new_n24987_,
    new_n24988_, new_n24989_, new_n24990_, new_n24991_, new_n24992_,
    new_n24993_, new_n24994_, new_n24995_, new_n24996_, new_n24997_,
    new_n24998_, new_n24999_, new_n25000_, new_n25001_, new_n25002_,
    new_n25003_, new_n25004_, new_n25005_, new_n25006_, new_n25007_,
    new_n25008_, new_n25009_, new_n25010_, new_n25011_, new_n25012_,
    new_n25013_, new_n25014_, new_n25015_, new_n25017_, new_n25018_,
    new_n25019_, new_n25020_, new_n25021_, new_n25022_, new_n25023_,
    new_n25024_, new_n25025_, new_n25026_, new_n25027_, new_n25028_,
    new_n25029_, new_n25030_, new_n25031_, new_n25032_, new_n25033_,
    new_n25034_, new_n25035_, new_n25036_, new_n25037_, new_n25038_,
    new_n25039_, new_n25040_, new_n25041_, new_n25042_, new_n25043_,
    new_n25044_, new_n25045_, new_n25046_, new_n25048_, new_n25049_,
    new_n25050_, new_n25051_, new_n25052_, new_n25053_, new_n25054_,
    new_n25055_, new_n25056_, new_n25057_, new_n25058_, new_n25059_,
    new_n25060_, new_n25061_, new_n25062_, new_n25063_, new_n25064_,
    new_n25065_, new_n25066_, new_n25067_, new_n25068_, new_n25069_,
    new_n25070_, new_n25071_, new_n25072_, new_n25073_, new_n25074_,
    new_n25075_, new_n25076_, new_n25077_, new_n25078_, new_n25079_,
    new_n25080_, new_n25081_, new_n25082_, new_n25083_, new_n25084_,
    new_n25085_, new_n25086_, new_n25087_, new_n25088_, new_n25089_,
    new_n25090_, new_n25091_, new_n25092_, new_n25093_, new_n25094_,
    new_n25095_, new_n25096_, new_n25097_, new_n25098_, new_n25099_,
    new_n25100_, new_n25101_, new_n25102_, new_n25103_, new_n25104_,
    new_n25105_, new_n25106_, new_n25107_, new_n25108_, new_n25109_,
    new_n25110_, new_n25111_, new_n25112_, new_n25113_, new_n25114_,
    new_n25115_, new_n25116_, new_n25117_, new_n25118_, new_n25119_,
    new_n25120_, new_n25121_, new_n25122_, new_n25123_, new_n25124_,
    new_n25125_, new_n25126_, new_n25127_, new_n25128_, new_n25129_,
    new_n25130_, new_n25131_, new_n25132_, new_n25133_, new_n25134_,
    new_n25135_, new_n25136_, new_n25137_, new_n25138_, new_n25139_,
    new_n25140_, new_n25141_, new_n25142_, new_n25143_, new_n25144_,
    new_n25145_, new_n25146_, new_n25147_, new_n25148_, new_n25149_,
    new_n25150_, new_n25151_, new_n25152_, new_n25153_, new_n25154_,
    new_n25155_, new_n25156_, new_n25157_, new_n25158_, new_n25159_,
    new_n25160_, new_n25161_, new_n25162_, new_n25163_, new_n25164_,
    new_n25165_, new_n25166_, new_n25167_, new_n25168_, new_n25169_,
    new_n25170_, new_n25171_, new_n25172_, new_n25173_, new_n25174_,
    new_n25175_, new_n25176_, new_n25177_, new_n25178_, new_n25179_,
    new_n25180_, new_n25181_, new_n25182_, new_n25183_, new_n25184_,
    new_n25185_, new_n25186_, new_n25187_, new_n25188_, new_n25189_,
    new_n25190_, new_n25191_, new_n25192_, new_n25193_, new_n25194_,
    new_n25195_, new_n25196_, new_n25197_, new_n25198_, new_n25199_,
    new_n25200_, new_n25201_, new_n25202_, new_n25203_, new_n25204_,
    new_n25205_, new_n25206_, new_n25207_, new_n25208_, new_n25209_,
    new_n25210_, new_n25211_, new_n25212_, new_n25213_, new_n25214_,
    new_n25215_, new_n25216_, new_n25217_, new_n25218_, new_n25219_,
    new_n25220_, new_n25221_, new_n25222_, new_n25223_, new_n25224_,
    new_n25225_, new_n25226_, new_n25227_, new_n25228_, new_n25229_,
    new_n25230_, new_n25231_, new_n25233_, new_n25234_, new_n25235_,
    new_n25236_, new_n25237_, new_n25238_, new_n25239_, new_n25240_,
    new_n25241_, new_n25242_, new_n25243_, new_n25244_, new_n25245_,
    new_n25246_, new_n25247_, new_n25248_, new_n25249_, new_n25250_,
    new_n25251_, new_n25252_, new_n25253_, new_n25254_, new_n25255_,
    new_n25256_, new_n25257_, new_n25258_, new_n25259_, new_n25260_,
    new_n25261_, new_n25262_, new_n25263_, new_n25264_, new_n25265_,
    new_n25266_, new_n25267_, new_n25268_, new_n25269_, new_n25270_,
    new_n25271_, new_n25272_, new_n25273_, new_n25274_, new_n25275_,
    new_n25276_, new_n25277_, new_n25278_, new_n25279_, new_n25280_,
    new_n25281_, new_n25282_, new_n25283_, new_n25284_, new_n25285_,
    new_n25286_, new_n25287_, new_n25288_, new_n25289_, new_n25290_,
    new_n25291_, new_n25292_, new_n25293_, new_n25294_, new_n25295_,
    new_n25296_, new_n25297_, new_n25298_, new_n25299_, new_n25300_,
    new_n25301_, new_n25302_, new_n25303_, new_n25304_, new_n25305_,
    new_n25306_, new_n25307_, new_n25308_, new_n25309_, new_n25310_,
    new_n25311_, new_n25312_, new_n25313_, new_n25314_, new_n25315_,
    new_n25316_, new_n25317_, new_n25318_, new_n25319_, new_n25320_,
    new_n25321_, new_n25322_, new_n25323_, new_n25324_, new_n25325_,
    new_n25326_, new_n25327_, new_n25328_, new_n25329_, new_n25330_,
    new_n25331_, new_n25332_, new_n25333_, new_n25334_, new_n25335_,
    new_n25336_, new_n25337_, new_n25338_, new_n25339_, new_n25340_,
    new_n25341_, new_n25342_, new_n25343_, new_n25344_, new_n25345_,
    new_n25346_, new_n25347_, new_n25348_, new_n25349_, new_n25350_,
    new_n25351_, new_n25352_, new_n25353_, new_n25354_, new_n25355_,
    new_n25356_, new_n25357_, new_n25358_, new_n25359_, new_n25360_,
    new_n25361_, new_n25362_, new_n25363_, new_n25364_, new_n25365_,
    new_n25366_, new_n25367_, new_n25368_, new_n25369_, new_n25370_,
    new_n25371_, new_n25372_, new_n25373_, new_n25374_, new_n25375_,
    new_n25376_, new_n25377_, new_n25378_, new_n25379_, new_n25380_,
    new_n25381_, new_n25382_, new_n25383_, new_n25384_, new_n25385_,
    new_n25386_, new_n25387_, new_n25388_, new_n25389_, new_n25390_,
    new_n25391_, new_n25392_, new_n25393_, new_n25394_, new_n25395_,
    new_n25396_, new_n25397_, new_n25398_, new_n25399_, new_n25400_,
    new_n25401_, new_n25402_, new_n25403_, new_n25404_, new_n25405_,
    new_n25406_, new_n25407_, new_n25408_, new_n25409_, new_n25410_,
    new_n25411_, new_n25412_, new_n25413_, new_n25414_, new_n25415_,
    new_n25416_, new_n25417_, new_n25418_, new_n25419_, new_n25420_,
    new_n25421_, new_n25422_, new_n25423_, new_n25424_, new_n25425_,
    new_n25426_, new_n25427_, new_n25428_, new_n25429_, new_n25430_,
    new_n25431_, new_n25432_, new_n25433_, new_n25434_, new_n25435_,
    new_n25436_, new_n25437_, new_n25438_, new_n25439_, new_n25440_,
    new_n25441_, new_n25442_, new_n25443_, new_n25444_, new_n25445_,
    new_n25447_, new_n25448_, new_n25449_, new_n25450_, new_n25451_,
    new_n25452_, new_n25453_, new_n25454_, new_n25455_, new_n25456_,
    new_n25457_, new_n25458_, new_n25459_, new_n25460_, new_n25461_,
    new_n25462_, new_n25463_, new_n25464_, new_n25465_, new_n25466_,
    new_n25467_, new_n25468_, new_n25469_, new_n25470_, new_n25471_,
    new_n25472_, new_n25473_, new_n25474_, new_n25475_, new_n25476_,
    new_n25477_, new_n25478_, new_n25479_, new_n25480_, new_n25481_,
    new_n25482_, new_n25483_, new_n25484_, new_n25485_, new_n25486_,
    new_n25487_, new_n25488_, new_n25489_, new_n25490_, new_n25491_,
    new_n25492_, new_n25493_, new_n25494_, new_n25495_, new_n25496_,
    new_n25497_, new_n25498_, new_n25499_, new_n25500_, new_n25501_,
    new_n25502_, new_n25503_, new_n25504_, new_n25505_, new_n25506_,
    new_n25507_, new_n25508_, new_n25509_, new_n25510_, new_n25511_,
    new_n25512_, new_n25513_, new_n25514_, new_n25515_, new_n25516_,
    new_n25517_, new_n25518_, new_n25519_, new_n25520_, new_n25521_,
    new_n25522_, new_n25523_, new_n25524_, new_n25525_, new_n25526_,
    new_n25527_, new_n25528_, new_n25529_, new_n25530_, new_n25531_,
    new_n25532_, new_n25533_, new_n25534_, new_n25535_, new_n25536_,
    new_n25537_, new_n25538_, new_n25539_, new_n25540_, new_n25541_,
    new_n25542_, new_n25543_, new_n25544_, new_n25545_, new_n25546_,
    new_n25547_, new_n25548_, new_n25549_, new_n25550_, new_n25551_,
    new_n25552_, new_n25553_, new_n25554_, new_n25555_, new_n25556_,
    new_n25557_, new_n25558_, new_n25559_, new_n25560_, new_n25561_,
    new_n25562_, new_n25563_, new_n25564_, new_n25565_, new_n25566_,
    new_n25567_, new_n25568_, new_n25569_, new_n25570_, new_n25571_,
    new_n25572_, new_n25573_, new_n25574_, new_n25575_, new_n25576_,
    new_n25577_, new_n25578_, new_n25579_, new_n25580_, new_n25581_,
    new_n25582_, new_n25583_, new_n25584_, new_n25585_, new_n25586_,
    new_n25587_, new_n25588_, new_n25589_, new_n25590_, new_n25591_,
    new_n25592_, new_n25593_, new_n25594_, new_n25595_, new_n25596_,
    new_n25597_, new_n25598_, new_n25599_, new_n25600_, new_n25601_,
    new_n25602_, new_n25603_, new_n25604_, new_n25605_, new_n25606_,
    new_n25607_, new_n25608_, new_n25609_, new_n25610_, new_n25611_,
    new_n25612_, new_n25613_, new_n25614_, new_n25615_, new_n25616_,
    new_n25617_, new_n25618_, new_n25619_, new_n25620_, new_n25621_,
    new_n25622_, new_n25623_, new_n25624_, new_n25625_, new_n25626_,
    new_n25627_, new_n25628_, new_n25629_, new_n25630_, new_n25631_,
    new_n25632_, new_n25633_, new_n25634_, new_n25635_, new_n25636_,
    new_n25637_, new_n25638_, new_n25639_, new_n25640_, new_n25641_,
    new_n25642_, new_n25643_, new_n25644_, new_n25645_, new_n25646_,
    new_n25647_, new_n25648_, new_n25649_, new_n25650_, new_n25651_,
    new_n25652_, new_n25653_, new_n25654_, new_n25655_, new_n25656_,
    new_n25657_, new_n25658_, new_n25659_, new_n25660_, new_n25661_,
    new_n25662_, new_n25663_, new_n25664_, new_n25665_, new_n25666_,
    new_n25667_, new_n25668_, new_n25669_, new_n25670_, new_n25671_,
    new_n25672_, new_n25673_, new_n25674_, new_n25675_, new_n25676_,
    new_n25677_, new_n25678_, new_n25679_, new_n25680_, new_n25681_,
    new_n25683_, new_n25684_, new_n25685_, new_n25686_, new_n25687_,
    new_n25688_, new_n25689_, new_n25690_, new_n25691_, new_n25692_,
    new_n25693_, new_n25694_, new_n25695_, new_n25696_, new_n25697_,
    new_n25698_, new_n25699_, new_n25700_, new_n25701_, new_n25702_,
    new_n25703_, new_n25704_, new_n25705_, new_n25706_, new_n25707_,
    new_n25708_, new_n25709_, new_n25710_, new_n25711_, new_n25712_,
    new_n25713_, new_n25714_, new_n25715_, new_n25716_, new_n25717_,
    new_n25718_, new_n25719_, new_n25720_, new_n25721_, new_n25722_,
    new_n25723_, new_n25724_, new_n25725_, new_n25726_, new_n25727_,
    new_n25728_, new_n25729_, new_n25730_, new_n25731_, new_n25732_,
    new_n25733_, new_n25734_, new_n25735_, new_n25736_, new_n25737_,
    new_n25738_, new_n25739_, new_n25740_, new_n25741_, new_n25742_,
    new_n25743_, new_n25744_, new_n25745_, new_n25746_, new_n25747_,
    new_n25748_, new_n25749_, new_n25750_, new_n25751_, new_n25752_,
    new_n25753_, new_n25754_, new_n25755_, new_n25756_, new_n25757_,
    new_n25758_, new_n25759_, new_n25760_, new_n25761_, new_n25762_,
    new_n25763_, new_n25764_, new_n25765_, new_n25766_, new_n25767_,
    new_n25768_, new_n25769_, new_n25770_, new_n25771_, new_n25772_,
    new_n25773_, new_n25774_, new_n25775_, new_n25776_, new_n25777_,
    new_n25778_, new_n25779_, new_n25780_, new_n25781_, new_n25782_,
    new_n25783_, new_n25784_, new_n25785_, new_n25786_, new_n25787_,
    new_n25788_, new_n25789_, new_n25790_, new_n25791_, new_n25792_,
    new_n25793_, new_n25794_, new_n25795_, new_n25796_, new_n25797_,
    new_n25798_, new_n25799_, new_n25800_, new_n25801_, new_n25802_,
    new_n25803_, new_n25804_, new_n25805_, new_n25806_, new_n25807_,
    new_n25808_, new_n25809_, new_n25810_, new_n25811_, new_n25812_,
    new_n25813_, new_n25814_, new_n25815_, new_n25816_, new_n25817_,
    new_n25818_, new_n25819_, new_n25820_, new_n25821_, new_n25822_,
    new_n25823_, new_n25824_, new_n25825_, new_n25826_, new_n25827_,
    new_n25828_, new_n25829_, new_n25830_, new_n25831_, new_n25832_,
    new_n25833_, new_n25834_, new_n25835_, new_n25836_, new_n25837_,
    new_n25838_, new_n25839_, new_n25840_, new_n25841_, new_n25842_,
    new_n25843_, new_n25844_, new_n25845_, new_n25846_, new_n25847_,
    new_n25848_, new_n25849_, new_n25850_, new_n25851_, new_n25852_,
    new_n25853_, new_n25854_, new_n25855_, new_n25856_, new_n25857_,
    new_n25858_, new_n25859_, new_n25860_, new_n25861_, new_n25862_,
    new_n25863_, new_n25864_, new_n25865_, new_n25866_, new_n25867_,
    new_n25868_, new_n25869_, new_n25870_, new_n25871_, new_n25872_,
    new_n25873_, new_n25874_, new_n25875_, new_n25876_, new_n25877_,
    new_n25878_, new_n25879_, new_n25880_, new_n25881_, new_n25882_,
    new_n25883_, new_n25884_, new_n25885_, new_n25886_, new_n25887_,
    new_n25888_, new_n25889_, new_n25890_, new_n25891_, new_n25892_,
    new_n25893_, new_n25894_, new_n25895_, new_n25897_, new_n25898_,
    new_n25899_, new_n25900_, new_n25901_, new_n25902_, new_n25903_,
    new_n25904_, new_n25905_, new_n25906_, new_n25907_, new_n25908_,
    new_n25909_, new_n25910_, new_n25911_, new_n25912_, new_n25913_,
    new_n25914_, new_n25915_, new_n25916_, new_n25917_, new_n25918_,
    new_n25919_, new_n25920_, new_n25921_, new_n25922_, new_n25923_,
    new_n25924_, new_n25925_, new_n25926_, new_n25927_, new_n25928_,
    new_n25929_, new_n25930_, new_n25931_, new_n25932_, new_n25933_,
    new_n25934_, new_n25935_, new_n25936_, new_n25937_, new_n25938_,
    new_n25939_, new_n25940_, new_n25941_, new_n25942_, new_n25943_,
    new_n25944_, new_n25945_, new_n25946_, new_n25947_, new_n25948_,
    new_n25949_, new_n25950_, new_n25951_, new_n25952_, new_n25953_,
    new_n25954_, new_n25955_, new_n25956_, new_n25957_, new_n25958_,
    new_n25959_, new_n25960_, new_n25961_, new_n25962_, new_n25963_,
    new_n25964_, new_n25965_, new_n25966_, new_n25967_, new_n25968_,
    new_n25969_, new_n25970_, new_n25971_, new_n25972_, new_n25973_,
    new_n25974_, new_n25975_, new_n25976_, new_n25977_, new_n25978_,
    new_n25979_, new_n25980_, new_n25981_, new_n25982_, new_n25983_,
    new_n25984_, new_n25985_, new_n25986_, new_n25987_, new_n25988_,
    new_n25989_, new_n25990_, new_n25991_, new_n25992_, new_n25993_,
    new_n25994_, new_n25995_, new_n25996_, new_n25997_, new_n25998_,
    new_n25999_, new_n26000_, new_n26001_, new_n26002_, new_n26003_,
    new_n26004_, new_n26005_, new_n26006_, new_n26007_, new_n26008_,
    new_n26009_, new_n26010_, new_n26011_, new_n26012_, new_n26013_,
    new_n26014_, new_n26015_, new_n26016_, new_n26017_, new_n26018_,
    new_n26019_, new_n26020_, new_n26021_, new_n26022_, new_n26023_,
    new_n26024_, new_n26025_, new_n26026_, new_n26027_, new_n26028_,
    new_n26029_, new_n26030_, new_n26031_, new_n26032_, new_n26033_,
    new_n26034_, new_n26035_, new_n26036_, new_n26037_, new_n26038_,
    new_n26039_, new_n26040_, new_n26041_, new_n26042_, new_n26043_,
    new_n26044_, new_n26045_, new_n26046_, new_n26047_, new_n26048_,
    new_n26049_, new_n26050_, new_n26051_, new_n26052_, new_n26053_,
    new_n26054_, new_n26055_, new_n26056_, new_n26057_, new_n26058_,
    new_n26059_, new_n26060_, new_n26061_, new_n26062_, new_n26063_,
    new_n26064_, new_n26065_, new_n26066_, new_n26067_, new_n26068_,
    new_n26069_, new_n26070_, new_n26071_, new_n26072_, new_n26073_,
    new_n26074_, new_n26075_, new_n26076_, new_n26077_, new_n26078_,
    new_n26079_, new_n26080_, new_n26081_, new_n26082_, new_n26083_,
    new_n26084_, new_n26085_, new_n26086_, new_n26087_, new_n26088_,
    new_n26089_, new_n26090_, new_n26091_, new_n26092_, new_n26093_,
    new_n26094_, new_n26095_, new_n26096_, new_n26097_, new_n26098_,
    new_n26099_, new_n26100_, new_n26101_, new_n26102_, new_n26104_,
    new_n26105_, new_n26106_, new_n26107_, new_n26108_, new_n26109_,
    new_n26110_, new_n26111_, new_n26112_, new_n26113_, new_n26114_,
    new_n26115_, new_n26116_, new_n26117_, new_n26118_, new_n26119_,
    new_n26120_, new_n26121_, new_n26122_, new_n26123_, new_n26124_,
    new_n26125_, new_n26126_, new_n26127_, new_n26128_, new_n26129_,
    new_n26130_, new_n26131_, new_n26132_, new_n26133_, new_n26134_,
    new_n26135_, new_n26136_, new_n26137_, new_n26138_, new_n26139_,
    new_n26140_, new_n26141_, new_n26142_, new_n26143_, new_n26144_,
    new_n26145_, new_n26146_, new_n26147_, new_n26148_, new_n26149_,
    new_n26150_, new_n26151_, new_n26152_, new_n26153_, new_n26154_,
    new_n26155_, new_n26156_, new_n26157_, new_n26158_, new_n26159_,
    new_n26160_, new_n26161_, new_n26162_, new_n26163_, new_n26164_,
    new_n26165_, new_n26166_, new_n26167_, new_n26168_, new_n26169_,
    new_n26170_, new_n26171_, new_n26172_, new_n26173_, new_n26174_,
    new_n26175_, new_n26176_, new_n26177_, new_n26178_, new_n26179_,
    new_n26180_, new_n26181_, new_n26182_, new_n26183_, new_n26184_,
    new_n26185_, new_n26186_, new_n26187_, new_n26188_, new_n26189_,
    new_n26190_, new_n26191_, new_n26192_, new_n26193_, new_n26194_,
    new_n26195_, new_n26196_, new_n26197_, new_n26198_, new_n26199_,
    new_n26200_, new_n26201_, new_n26202_, new_n26203_, new_n26204_,
    new_n26205_, new_n26206_, new_n26207_, new_n26208_, new_n26209_,
    new_n26210_, new_n26211_, new_n26212_, new_n26213_, new_n26214_,
    new_n26215_, new_n26216_, new_n26217_, new_n26218_, new_n26219_,
    new_n26220_, new_n26221_, new_n26222_, new_n26223_, new_n26224_,
    new_n26225_, new_n26226_, new_n26227_, new_n26228_, new_n26229_,
    new_n26230_, new_n26231_, new_n26232_, new_n26233_, new_n26234_,
    new_n26235_, new_n26236_, new_n26237_, new_n26238_, new_n26239_,
    new_n26240_, new_n26241_, new_n26242_, new_n26243_, new_n26244_,
    new_n26245_, new_n26246_, new_n26247_, new_n26248_, new_n26249_,
    new_n26250_, new_n26251_, new_n26252_, new_n26253_, new_n26254_,
    new_n26255_, new_n26256_, new_n26257_, new_n26258_, new_n26259_,
    new_n26260_, new_n26261_, new_n26262_, new_n26263_, new_n26265_,
    new_n26266_, new_n26267_, new_n26268_, new_n26269_, new_n26270_,
    new_n26271_, new_n26272_, new_n26273_, new_n26274_, new_n26275_,
    new_n26276_, new_n26277_, new_n26278_, new_n26279_, new_n26280_,
    new_n26281_, new_n26282_, new_n26283_, new_n26284_, new_n26285_,
    new_n26286_, new_n26287_, new_n26288_, new_n26289_, new_n26290_,
    new_n26291_, new_n26292_, new_n26293_, new_n26294_, new_n26295_,
    new_n26296_, new_n26297_, new_n26298_, new_n26299_, new_n26300_,
    new_n26301_, new_n26302_, new_n26303_, new_n26304_, new_n26305_,
    new_n26306_, new_n26307_, new_n26308_, new_n26309_, new_n26310_,
    new_n26311_, new_n26312_, new_n26313_, new_n26314_, new_n26315_,
    new_n26316_, new_n26317_, new_n26318_, new_n26319_, new_n26320_,
    new_n26321_, new_n26322_, new_n26323_, new_n26324_, new_n26325_,
    new_n26326_, new_n26327_, new_n26328_, new_n26329_, new_n26330_,
    new_n26331_, new_n26332_, new_n26333_, new_n26334_, new_n26335_,
    new_n26336_, new_n26337_, new_n26338_, new_n26339_, new_n26340_,
    new_n26341_, new_n26342_, new_n26343_, new_n26344_, new_n26345_,
    new_n26346_, new_n26347_, new_n26348_, new_n26349_, new_n26350_,
    new_n26351_, new_n26352_, new_n26353_, new_n26354_, new_n26355_,
    new_n26356_, new_n26357_, new_n26358_, new_n26359_, new_n26360_,
    new_n26361_, new_n26362_, new_n26363_, new_n26364_, new_n26365_,
    new_n26366_, new_n26367_, new_n26368_, new_n26369_, new_n26370_,
    new_n26371_, new_n26372_, new_n26373_, new_n26374_, new_n26375_,
    new_n26376_, new_n26377_, new_n26378_, new_n26379_, new_n26380_,
    new_n26381_, new_n26382_, new_n26383_, new_n26384_, new_n26385_,
    new_n26386_, new_n26387_, new_n26388_, new_n26389_, new_n26390_,
    new_n26391_, new_n26392_, new_n26393_, new_n26394_, new_n26395_,
    new_n26396_, new_n26397_, new_n26398_, new_n26399_, new_n26400_,
    new_n26401_, new_n26402_, new_n26403_, new_n26404_, new_n26405_,
    new_n26406_, new_n26407_, new_n26408_, new_n26409_, new_n26410_,
    new_n26411_, new_n26412_, new_n26413_, new_n26414_, new_n26415_,
    new_n26416_, new_n26417_, new_n26418_, new_n26419_, new_n26420_,
    new_n26421_, new_n26422_, new_n26423_, new_n26424_, new_n26425_,
    new_n26426_, new_n26427_, new_n26428_, new_n26429_, new_n26430_,
    new_n26431_, new_n26432_, new_n26433_, new_n26435_, new_n26436_,
    new_n26437_, new_n26438_, new_n26439_, new_n26440_, new_n26441_,
    new_n26442_, new_n26443_, new_n26444_, new_n26445_, new_n26446_,
    new_n26447_, new_n26448_, new_n26449_, new_n26450_, new_n26451_,
    new_n26452_, new_n26453_, new_n26454_, new_n26455_, new_n26456_,
    new_n26457_, new_n26458_, new_n26459_, new_n26460_, new_n26461_,
    new_n26462_, new_n26463_, new_n26464_, new_n26465_, new_n26466_,
    new_n26467_, new_n26468_, new_n26469_, new_n26470_, new_n26471_,
    new_n26472_, new_n26473_, new_n26474_, new_n26475_, new_n26476_,
    new_n26477_, new_n26478_, new_n26479_, new_n26480_, new_n26481_,
    new_n26482_, new_n26483_, new_n26484_, new_n26485_, new_n26486_,
    new_n26487_, new_n26488_, new_n26489_, new_n26490_, new_n26491_,
    new_n26492_, new_n26493_, new_n26494_, new_n26495_, new_n26496_,
    new_n26497_, new_n26498_, new_n26499_, new_n26500_, new_n26501_,
    new_n26502_, new_n26503_, new_n26504_, new_n26505_, new_n26506_,
    new_n26507_, new_n26508_, new_n26509_, new_n26510_, new_n26511_,
    new_n26512_, new_n26513_, new_n26514_, new_n26515_, new_n26516_,
    new_n26517_, new_n26518_, new_n26519_, new_n26520_, new_n26521_,
    new_n26522_, new_n26523_, new_n26524_, new_n26525_, new_n26526_,
    new_n26527_, new_n26528_, new_n26529_, new_n26530_, new_n26531_,
    new_n26532_, new_n26533_, new_n26534_, new_n26535_, new_n26536_,
    new_n26537_, new_n26538_, new_n26539_, new_n26540_, new_n26541_,
    new_n26542_, new_n26543_, new_n26544_, new_n26545_, new_n26546_,
    new_n26547_, new_n26548_, new_n26549_, new_n26550_, new_n26551_,
    new_n26552_, new_n26553_, new_n26554_, new_n26555_, new_n26556_,
    new_n26557_, new_n26558_, new_n26559_, new_n26560_, new_n26561_,
    new_n26562_, new_n26563_, new_n26564_, new_n26565_, new_n26566_,
    new_n26567_, new_n26568_, new_n26569_, new_n26570_, new_n26571_,
    new_n26572_, new_n26573_, new_n26574_, new_n26575_, new_n26576_,
    new_n26577_, new_n26578_, new_n26579_, new_n26580_, new_n26581_,
    new_n26582_, new_n26583_, new_n26584_, new_n26585_, new_n26586_,
    new_n26587_, new_n26588_, new_n26589_, new_n26590_, new_n26591_,
    new_n26592_, new_n26593_, new_n26595_, new_n26596_, new_n26597_,
    new_n26598_, new_n26599_, new_n26600_, new_n26601_, new_n26602_,
    new_n26603_, new_n26604_, new_n26605_, new_n26606_, new_n26607_,
    new_n26608_, new_n26609_, new_n26610_, new_n26611_, new_n26612_,
    new_n26613_, new_n26614_, new_n26615_, new_n26616_, new_n26617_,
    new_n26618_, new_n26619_, new_n26620_, new_n26621_, new_n26622_,
    new_n26623_, new_n26624_, new_n26625_, new_n26626_, new_n26627_,
    new_n26628_, new_n26629_, new_n26630_, new_n26631_, new_n26632_,
    new_n26633_, new_n26634_, new_n26635_, new_n26636_, new_n26637_,
    new_n26638_, new_n26639_, new_n26640_, new_n26641_, new_n26642_,
    new_n26643_, new_n26644_, new_n26645_, new_n26646_, new_n26647_,
    new_n26648_, new_n26649_, new_n26650_, new_n26651_, new_n26652_,
    new_n26653_, new_n26654_, new_n26655_, new_n26656_, new_n26657_,
    new_n26658_, new_n26659_, new_n26660_, new_n26661_, new_n26662_,
    new_n26663_, new_n26664_, new_n26665_, new_n26666_, new_n26667_,
    new_n26668_, new_n26669_, new_n26670_, new_n26671_, new_n26672_,
    new_n26673_, new_n26674_, new_n26675_, new_n26676_, new_n26677_,
    new_n26678_, new_n26679_, new_n26680_, new_n26681_, new_n26682_,
    new_n26683_, new_n26684_, new_n26685_, new_n26686_, new_n26687_,
    new_n26688_, new_n26689_, new_n26690_, new_n26691_, new_n26692_,
    new_n26693_, new_n26694_, new_n26695_, new_n26696_, new_n26697_,
    new_n26698_, new_n26699_, new_n26700_, new_n26701_, new_n26702_,
    new_n26703_, new_n26704_, new_n26705_, new_n26706_, new_n26707_,
    new_n26708_, new_n26709_, new_n26710_, new_n26712_, new_n26713_,
    new_n26714_, new_n26715_, new_n26716_, new_n26717_, new_n26718_,
    new_n26719_, new_n26720_, new_n26721_, new_n26722_, new_n26723_,
    new_n26724_, new_n26725_, new_n26726_, new_n26727_, new_n26728_,
    new_n26729_, new_n26730_, new_n26731_, new_n26732_, new_n26733_,
    new_n26734_, new_n26735_, new_n26736_, new_n26737_, new_n26738_,
    new_n26739_, new_n26740_, new_n26741_, new_n26742_, new_n26743_,
    new_n26744_, new_n26745_, new_n26746_, new_n26747_, new_n26748_,
    new_n26749_, new_n26750_, new_n26751_, new_n26752_, new_n26753_,
    new_n26754_, new_n26755_, new_n26756_, new_n26757_, new_n26758_,
    new_n26759_, new_n26760_, new_n26761_, new_n26762_, new_n26763_,
    new_n26764_, new_n26765_, new_n26766_, new_n26767_, new_n26768_,
    new_n26769_, new_n26770_, new_n26771_, new_n26772_, new_n26773_,
    new_n26774_, new_n26775_, new_n26776_, new_n26777_, new_n26778_,
    new_n26779_, new_n26780_, new_n26781_, new_n26782_, new_n26783_,
    new_n26784_, new_n26785_, new_n26786_, new_n26787_, new_n26788_,
    new_n26789_, new_n26790_, new_n26791_, new_n26792_, new_n26793_,
    new_n26794_, new_n26795_, new_n26796_, new_n26797_, new_n26798_,
    new_n26799_, new_n26800_, new_n26801_, new_n26802_, new_n26803_,
    new_n26804_, new_n26805_, new_n26806_, new_n26807_, new_n26808_,
    new_n26809_, new_n26810_, new_n26811_, new_n26812_, new_n26813_,
    new_n26814_, new_n26815_, new_n26816_, new_n26817_, new_n26818_,
    new_n26819_, new_n26820_, new_n26821_, new_n26822_, new_n26823_,
    new_n26824_, new_n26825_, new_n26826_, new_n26827_, new_n26828_,
    new_n26829_, new_n26830_, new_n26832_, new_n26833_, new_n26834_,
    new_n26835_, new_n26836_, new_n26837_, new_n26838_, new_n26839_,
    new_n26840_, new_n26841_, new_n26842_, new_n26843_, new_n26844_,
    new_n26845_, new_n26846_, new_n26847_, new_n26848_, new_n26849_,
    new_n26850_, new_n26851_, new_n26852_, new_n26853_, new_n26854_,
    new_n26855_, new_n26856_, new_n26857_, new_n26858_, new_n26859_,
    new_n26860_, new_n26861_, new_n26862_, new_n26863_, new_n26864_,
    new_n26865_, new_n26866_, new_n26867_, new_n26868_, new_n26869_,
    new_n26870_, new_n26871_, new_n26872_, new_n26873_, new_n26874_,
    new_n26875_, new_n26876_, new_n26877_, new_n26878_, new_n26879_,
    new_n26880_, new_n26881_, new_n26882_, new_n26883_, new_n26884_,
    new_n26885_, new_n26886_, new_n26887_, new_n26888_, new_n26889_,
    new_n26890_, new_n26891_, new_n26892_, new_n26893_, new_n26894_,
    new_n26895_, new_n26896_, new_n26897_, new_n26898_, new_n26899_,
    new_n26900_, new_n26901_, new_n26902_, new_n26903_, new_n26904_,
    new_n26905_, new_n26906_, new_n26907_, new_n26908_, new_n26909_,
    new_n26910_, new_n26911_, new_n26912_, new_n26913_, new_n26914_,
    new_n26915_, new_n26916_, new_n26917_, new_n26918_, new_n26919_,
    new_n26920_, new_n26921_, new_n26922_, new_n26923_, new_n26924_,
    new_n26925_, new_n26926_, new_n26927_, new_n26928_, new_n26929_,
    new_n26930_, new_n26931_, new_n26932_, new_n26933_, new_n26934_,
    new_n26935_, new_n26936_, new_n26937_, new_n26938_, new_n26939_,
    new_n26940_, new_n26941_, new_n26942_, new_n26943_, new_n26945_,
    new_n26946_, new_n26947_, new_n26948_, new_n26949_, new_n26950_,
    new_n26951_, new_n26952_, new_n26953_, new_n26954_, new_n26955_,
    new_n26956_, new_n26957_, new_n26958_, new_n26959_, new_n26960_,
    new_n26961_, new_n26962_, new_n26963_, new_n26964_, new_n26965_,
    new_n26966_, new_n26967_, new_n26968_, new_n26969_, new_n26970_,
    new_n26971_, new_n26972_, new_n26973_, new_n26974_, new_n26975_,
    new_n26976_, new_n26977_, new_n26978_, new_n26979_, new_n26980_,
    new_n26981_, new_n26982_, new_n26983_, new_n26984_, new_n26985_,
    new_n26986_, new_n26987_, new_n26988_, new_n26989_, new_n26990_,
    new_n26991_, new_n26992_, new_n26993_, new_n26994_, new_n26995_,
    new_n26996_, new_n26997_, new_n26998_, new_n26999_, new_n27000_,
    new_n27001_, new_n27002_, new_n27003_, new_n27004_, new_n27005_,
    new_n27006_, new_n27007_, new_n27008_, new_n27009_, new_n27010_,
    new_n27011_, new_n27012_, new_n27013_, new_n27014_, new_n27015_,
    new_n27016_, new_n27017_, new_n27018_, new_n27019_, new_n27020_,
    new_n27021_, new_n27022_, new_n27023_, new_n27024_, new_n27025_,
    new_n27026_, new_n27027_, new_n27028_, new_n27029_, new_n27030_,
    new_n27031_, new_n27032_, new_n27033_, new_n27034_, new_n27035_,
    new_n27036_, new_n27037_, new_n27038_, new_n27039_, new_n27040_,
    new_n27041_, new_n27042_, new_n27043_, new_n27044_, new_n27045_,
    new_n27046_, new_n27047_, new_n27048_, new_n27049_, new_n27050_,
    new_n27051_, new_n27052_, new_n27053_, new_n27054_, new_n27055_,
    new_n27056_, new_n27057_, new_n27059_, new_n27060_, new_n27061_,
    new_n27062_, new_n27063_, new_n27064_, new_n27065_, new_n27066_,
    new_n27067_, new_n27068_, new_n27069_, new_n27070_, new_n27071_,
    new_n27072_, new_n27073_, new_n27074_, new_n27075_, new_n27076_,
    new_n27077_, new_n27078_, new_n27079_, new_n27080_, new_n27081_,
    new_n27082_, new_n27083_, new_n27084_, new_n27085_, new_n27086_,
    new_n27087_, new_n27088_, new_n27089_, new_n27090_, new_n27091_,
    new_n27092_, new_n27093_, new_n27094_, new_n27095_, new_n27096_,
    new_n27097_, new_n27098_, new_n27099_, new_n27100_, new_n27101_,
    new_n27102_, new_n27103_, new_n27104_, new_n27105_, new_n27106_,
    new_n27107_, new_n27108_, new_n27109_, new_n27110_, new_n27111_,
    new_n27112_, new_n27113_, new_n27114_, new_n27115_, new_n27116_,
    new_n27117_, new_n27118_, new_n27119_, new_n27120_, new_n27121_,
    new_n27122_, new_n27123_, new_n27124_, new_n27125_, new_n27126_,
    new_n27127_, new_n27128_, new_n27129_, new_n27130_, new_n27131_,
    new_n27132_, new_n27133_, new_n27134_, new_n27135_, new_n27136_,
    new_n27137_, new_n27138_, new_n27139_, new_n27140_, new_n27141_,
    new_n27142_, new_n27143_, new_n27144_, new_n27145_, new_n27146_,
    new_n27147_, new_n27148_, new_n27149_, new_n27150_, new_n27151_,
    new_n27152_, new_n27153_, new_n27154_, new_n27155_, new_n27156_,
    new_n27157_, new_n27158_, new_n27159_, new_n27160_, new_n27161_,
    new_n27162_, new_n27163_, new_n27164_, new_n27165_, new_n27166_,
    new_n27167_, new_n27168_, new_n27169_, new_n27170_, new_n27171_,
    new_n27172_, new_n27173_, new_n27174_, new_n27175_, new_n27176_,
    new_n27177_, new_n27178_, new_n27179_, new_n27180_, new_n27181_,
    new_n27182_, new_n27183_, new_n27184_, new_n27185_, new_n27186_,
    new_n27188_, new_n27189_, new_n27190_, new_n27191_, new_n27192_,
    new_n27193_, new_n27194_, new_n27195_, new_n27196_, new_n27197_,
    new_n27198_, new_n27199_, new_n27200_, new_n27201_, new_n27202_,
    new_n27203_, new_n27204_, new_n27205_, new_n27206_, new_n27207_,
    new_n27208_, new_n27209_, new_n27210_, new_n27211_, new_n27212_,
    new_n27213_, new_n27214_, new_n27215_, new_n27216_, new_n27217_,
    new_n27218_, new_n27219_, new_n27220_, new_n27221_, new_n27222_,
    new_n27223_, new_n27224_, new_n27225_, new_n27226_, new_n27227_,
    new_n27228_, new_n27229_, new_n27230_, new_n27231_, new_n27232_,
    new_n27233_, new_n27234_, new_n27235_, new_n27236_, new_n27237_,
    new_n27238_, new_n27239_, new_n27240_, new_n27241_, new_n27242_,
    new_n27243_, new_n27244_, new_n27245_, new_n27246_, new_n27247_,
    new_n27248_, new_n27249_, new_n27250_, new_n27251_, new_n27252_,
    new_n27253_, new_n27254_, new_n27255_, new_n27256_, new_n27257_,
    new_n27258_, new_n27259_, new_n27260_, new_n27261_, new_n27262_,
    new_n27263_, new_n27264_, new_n27265_, new_n27266_, new_n27267_,
    new_n27268_, new_n27269_, new_n27270_, new_n27271_, new_n27272_,
    new_n27273_, new_n27274_, new_n27275_, new_n27276_, new_n27277_,
    new_n27278_, new_n27279_, new_n27280_, new_n27281_, new_n27282_,
    new_n27283_, new_n27284_, new_n27285_, new_n27286_, new_n27287_,
    new_n27288_, new_n27289_, new_n27290_, new_n27291_, new_n27292_,
    new_n27293_, new_n27294_, new_n27295_, new_n27296_, new_n27297_,
    new_n27298_, new_n27299_, new_n27300_, new_n27301_, new_n27302_,
    new_n27303_, new_n27304_, new_n27305_, new_n27306_, new_n27307_,
    new_n27308_, new_n27309_, new_n27311_, new_n27312_, new_n27313_,
    new_n27314_, new_n27315_, new_n27316_, new_n27317_, new_n27318_,
    new_n27319_, new_n27320_, new_n27321_, new_n27322_, new_n27323_,
    new_n27324_, new_n27325_, new_n27326_, new_n27327_, new_n27328_,
    new_n27329_, new_n27330_, new_n27331_, new_n27332_, new_n27333_,
    new_n27334_, new_n27335_, new_n27336_, new_n27337_, new_n27338_,
    new_n27339_, new_n27340_, new_n27341_, new_n27342_, new_n27343_,
    new_n27344_, new_n27345_, new_n27346_, new_n27347_, new_n27348_,
    new_n27349_, new_n27350_, new_n27351_, new_n27352_, new_n27353_,
    new_n27354_, new_n27355_, new_n27356_, new_n27357_, new_n27358_,
    new_n27359_, new_n27360_, new_n27361_, new_n27362_, new_n27363_,
    new_n27364_, new_n27365_, new_n27366_, new_n27367_, new_n27368_,
    new_n27369_, new_n27370_, new_n27371_, new_n27372_, new_n27373_,
    new_n27374_, new_n27375_, new_n27376_, new_n27377_, new_n27378_,
    new_n27379_, new_n27380_, new_n27381_, new_n27382_, new_n27383_,
    new_n27384_, new_n27385_, new_n27386_, new_n27387_, new_n27388_,
    new_n27389_, new_n27390_, new_n27391_, new_n27392_, new_n27393_,
    new_n27394_, new_n27395_, new_n27396_, new_n27397_, new_n27398_,
    new_n27399_, new_n27400_, new_n27401_, new_n27402_, new_n27403_,
    new_n27404_, new_n27405_, new_n27406_, new_n27407_, new_n27408_,
    new_n27409_, new_n27410_, new_n27411_, new_n27412_, new_n27413_,
    new_n27414_, new_n27415_, new_n27416_, new_n27417_, new_n27418_,
    new_n27419_, new_n27420_, new_n27421_, new_n27423_, new_n27424_,
    new_n27425_, new_n27426_, new_n27427_, new_n27428_, new_n27429_,
    new_n27430_, new_n27431_, new_n27432_, new_n27433_, new_n27434_,
    new_n27435_, new_n27436_, new_n27437_, new_n27438_, new_n27439_,
    new_n27440_, new_n27441_, new_n27442_, new_n27443_, new_n27444_,
    new_n27445_, new_n27446_, new_n27447_, new_n27448_, new_n27449_,
    new_n27450_, new_n27451_, new_n27452_, new_n27453_, new_n27454_,
    new_n27455_, new_n27456_, new_n27457_, new_n27458_, new_n27459_,
    new_n27460_, new_n27461_, new_n27462_, new_n27463_, new_n27464_,
    new_n27465_, new_n27466_, new_n27467_, new_n27468_, new_n27469_,
    new_n27470_, new_n27471_, new_n27472_, new_n27473_, new_n27474_,
    new_n27475_, new_n27476_, new_n27477_, new_n27478_, new_n27479_,
    new_n27480_, new_n27481_, new_n27482_, new_n27483_, new_n27484_,
    new_n27485_, new_n27486_, new_n27487_, new_n27488_, new_n27489_,
    new_n27490_, new_n27491_, new_n27492_, new_n27493_, new_n27494_,
    new_n27495_, new_n27496_, new_n27497_, new_n27498_, new_n27499_,
    new_n27500_, new_n27501_, new_n27502_, new_n27503_, new_n27504_,
    new_n27505_, new_n27506_, new_n27507_, new_n27508_, new_n27509_,
    new_n27510_, new_n27511_, new_n27512_, new_n27513_, new_n27514_,
    new_n27515_, new_n27517_, new_n27518_, new_n27519_, new_n27520_,
    new_n27521_, new_n27522_, new_n27523_, new_n27524_, new_n27525_,
    new_n27526_, new_n27527_, new_n27528_, new_n27529_, new_n27530_,
    new_n27531_, new_n27532_, new_n27533_, new_n27534_, new_n27535_,
    new_n27536_, new_n27537_, new_n27538_, new_n27539_, new_n27540_,
    new_n27541_, new_n27542_, new_n27543_, new_n27544_, new_n27545_,
    new_n27546_, new_n27547_, new_n27548_, new_n27549_, new_n27550_,
    new_n27551_, new_n27552_, new_n27553_, new_n27554_, new_n27555_,
    new_n27556_, new_n27557_, new_n27558_, new_n27559_, new_n27560_,
    new_n27561_, new_n27562_, new_n27563_, new_n27564_, new_n27565_,
    new_n27566_, new_n27567_, new_n27568_, new_n27569_, new_n27570_,
    new_n27571_, new_n27572_, new_n27573_, new_n27574_, new_n27575_,
    new_n27576_, new_n27577_, new_n27578_, new_n27579_, new_n27580_,
    new_n27581_, new_n27582_, new_n27583_, new_n27584_, new_n27585_,
    new_n27586_, new_n27587_, new_n27588_, new_n27589_, new_n27590_,
    new_n27591_, new_n27592_, new_n27593_, new_n27594_, new_n27595_,
    new_n27596_, new_n27597_, new_n27598_, new_n27599_, new_n27600_,
    new_n27601_, new_n27602_, new_n27603_, new_n27604_, new_n27605_,
    new_n27606_, new_n27607_, new_n27608_, new_n27609_, new_n27610_,
    new_n27611_, new_n27612_, new_n27613_, new_n27614_, new_n27615_,
    new_n27616_, new_n27617_, new_n27618_, new_n27620_, new_n27621_,
    new_n27622_, new_n27623_, new_n27624_, new_n27625_, new_n27626_,
    new_n27627_, new_n27628_, new_n27629_, new_n27630_, new_n27631_,
    new_n27632_, new_n27633_, new_n27634_, new_n27635_, new_n27636_,
    new_n27637_, new_n27638_, new_n27639_, new_n27640_, new_n27641_,
    new_n27642_, new_n27643_, new_n27644_, new_n27645_, new_n27646_,
    new_n27647_, new_n27648_, new_n27649_, new_n27650_, new_n27651_,
    new_n27652_, new_n27653_, new_n27654_, new_n27655_, new_n27656_,
    new_n27657_, new_n27658_, new_n27659_, new_n27660_, new_n27661_,
    new_n27662_, new_n27663_, new_n27664_, new_n27665_, new_n27666_,
    new_n27667_, new_n27668_, new_n27669_, new_n27670_, new_n27671_,
    new_n27672_, new_n27673_, new_n27674_, new_n27675_, new_n27676_,
    new_n27677_, new_n27678_, new_n27679_, new_n27680_, new_n27681_,
    new_n27682_, new_n27683_, new_n27684_, new_n27685_, new_n27686_,
    new_n27687_, new_n27688_, new_n27689_, new_n27690_, new_n27691_,
    new_n27692_, new_n27693_, new_n27694_, new_n27695_, new_n27696_,
    new_n27697_, new_n27698_, new_n27699_, new_n27700_, new_n27701_,
    new_n27702_, new_n27704_, new_n27705_, new_n27706_, new_n27707_,
    new_n27708_, new_n27709_, new_n27710_, new_n27711_, new_n27712_,
    new_n27713_, new_n27714_, new_n27715_, new_n27716_, new_n27717_,
    new_n27718_, new_n27719_, new_n27720_, new_n27721_, new_n27722_,
    new_n27723_, new_n27724_, new_n27725_, new_n27726_, new_n27727_,
    new_n27728_, new_n27729_, new_n27730_, new_n27731_, new_n27732_,
    new_n27733_, new_n27734_, new_n27735_, new_n27736_, new_n27737_,
    new_n27738_, new_n27739_, new_n27740_, new_n27741_, new_n27742_,
    new_n27743_, new_n27744_, new_n27745_, new_n27746_, new_n27747_,
    new_n27748_, new_n27749_, new_n27750_, new_n27751_, new_n27752_,
    new_n27753_, new_n27754_, new_n27755_, new_n27756_, new_n27757_,
    new_n27758_, new_n27759_, new_n27760_, new_n27761_, new_n27762_,
    new_n27763_, new_n27764_, new_n27765_, new_n27766_, new_n27767_,
    new_n27768_, new_n27769_, new_n27770_, new_n27771_, new_n27772_,
    new_n27773_, new_n27774_, new_n27775_, new_n27776_, new_n27777_,
    new_n27778_, new_n27779_, new_n27780_, new_n27781_, new_n27782_,
    new_n27783_, new_n27784_, new_n27785_, new_n27786_, new_n27787_,
    new_n27788_, new_n27789_, new_n27790_, new_n27791_, new_n27792_,
    new_n27793_, new_n27794_, new_n27795_, new_n27796_, new_n27797_,
    new_n27798_, new_n27799_, new_n27800_, new_n27801_, new_n27802_,
    new_n27803_, new_n27804_, new_n27805_, new_n27806_, new_n27807_,
    new_n27808_, new_n27809_, new_n27810_, new_n27811_, new_n27812_,
    new_n27813_, new_n27814_, new_n27815_, new_n27816_, new_n27818_,
    new_n27819_, new_n27820_, new_n27821_, new_n27822_, new_n27823_,
    new_n27824_, new_n27825_, new_n27826_, new_n27827_, new_n27828_,
    new_n27829_, new_n27830_, new_n27831_, new_n27832_, new_n27833_,
    new_n27834_, new_n27835_, new_n27836_, new_n27837_, new_n27838_,
    new_n27839_, new_n27840_, new_n27841_, new_n27842_, new_n27843_,
    new_n27844_, new_n27845_, new_n27846_, new_n27847_, new_n27848_,
    new_n27849_, new_n27850_, new_n27851_, new_n27852_, new_n27853_,
    new_n27854_, new_n27855_, new_n27856_, new_n27857_, new_n27858_,
    new_n27859_, new_n27860_, new_n27861_, new_n27862_, new_n27863_,
    new_n27864_, new_n27865_, new_n27866_, new_n27867_, new_n27868_,
    new_n27869_, new_n27870_, new_n27871_, new_n27872_, new_n27873_,
    new_n27874_, new_n27875_, new_n27876_, new_n27877_, new_n27878_,
    new_n27879_, new_n27880_, new_n27881_, new_n27882_, new_n27883_,
    new_n27884_, new_n27885_, new_n27886_, new_n27887_, new_n27888_,
    new_n27889_, new_n27890_, new_n27891_, new_n27892_, new_n27893_,
    new_n27894_, new_n27895_, new_n27896_, new_n27897_, new_n27898_,
    new_n27899_, new_n27900_, new_n27901_, new_n27902_, new_n27904_,
    new_n27905_, new_n27906_, new_n27907_, new_n27908_, new_n27909_,
    new_n27910_, new_n27911_, new_n27912_, new_n27913_, new_n27914_,
    new_n27915_, new_n27916_, new_n27917_, new_n27918_, new_n27919_,
    new_n27920_, new_n27921_, new_n27922_, new_n27923_, new_n27924_,
    new_n27925_, new_n27926_, new_n27927_, new_n27928_, new_n27929_,
    new_n27930_, new_n27931_, new_n27932_, new_n27933_, new_n27934_,
    new_n27935_, new_n27936_, new_n27937_, new_n27938_, new_n27939_,
    new_n27940_, new_n27941_, new_n27942_, new_n27943_, new_n27944_,
    new_n27945_, new_n27946_, new_n27947_, new_n27948_, new_n27949_,
    new_n27950_, new_n27951_, new_n27952_, new_n27953_, new_n27954_,
    new_n27955_, new_n27956_, new_n27957_, new_n27958_, new_n27959_,
    new_n27960_, new_n27961_, new_n27962_, new_n27963_, new_n27964_,
    new_n27965_, new_n27966_, new_n27967_, new_n27968_, new_n27969_,
    new_n27970_, new_n27971_, new_n27972_, new_n27973_, new_n27974_,
    new_n27975_, new_n27976_, new_n27977_, new_n27978_, new_n27979_,
    new_n27980_, new_n27981_, new_n27982_, new_n27983_, new_n27984_,
    new_n27985_, new_n27986_, new_n27987_, new_n27988_, new_n27989_,
    new_n27990_, new_n27991_, new_n27992_, new_n27993_, new_n27995_,
    new_n27996_, new_n27997_, new_n27998_, new_n27999_, new_n28000_,
    new_n28001_, new_n28002_, new_n28003_, new_n28004_, new_n28005_,
    new_n28006_, new_n28007_, new_n28008_, new_n28009_, new_n28010_,
    new_n28011_, new_n28012_, new_n28013_, new_n28014_, new_n28015_,
    new_n28016_, new_n28017_, new_n28018_, new_n28019_, new_n28020_,
    new_n28021_, new_n28022_, new_n28023_, new_n28024_, new_n28025_,
    new_n28026_, new_n28027_, new_n28028_, new_n28029_, new_n28030_,
    new_n28031_, new_n28032_, new_n28033_, new_n28034_, new_n28035_,
    new_n28036_, new_n28037_, new_n28038_, new_n28039_, new_n28040_,
    new_n28041_, new_n28042_, new_n28043_, new_n28044_, new_n28045_,
    new_n28046_, new_n28047_, new_n28048_, new_n28049_, new_n28050_,
    new_n28051_, new_n28052_, new_n28053_, new_n28054_, new_n28055_,
    new_n28056_, new_n28057_, new_n28058_, new_n28059_, new_n28060_,
    new_n28061_, new_n28062_, new_n28063_, new_n28064_, new_n28065_,
    new_n28066_, new_n28067_, new_n28068_, new_n28069_, new_n28070_,
    new_n28071_, new_n28072_, new_n28073_, new_n28074_, new_n28075_,
    new_n28076_, new_n28077_, new_n28078_, new_n28079_, new_n28080_,
    new_n28081_, new_n28082_, new_n28083_, new_n28084_, new_n28085_,
    new_n28086_, new_n28087_, new_n28089_, new_n28090_, new_n28091_,
    new_n28092_, new_n28093_, new_n28094_, new_n28095_, new_n28096_,
    new_n28097_, new_n28098_, new_n28099_, new_n28100_, new_n28101_,
    new_n28102_, new_n28103_, new_n28104_, new_n28105_, new_n28106_,
    new_n28107_, new_n28108_, new_n28109_, new_n28110_, new_n28111_,
    new_n28112_, new_n28113_, new_n28114_, new_n28115_, new_n28116_,
    new_n28117_, new_n28118_, new_n28119_, new_n28120_, new_n28121_,
    new_n28122_, new_n28123_, new_n28124_, new_n28125_, new_n28126_,
    new_n28127_, new_n28128_, new_n28129_, new_n28130_, new_n28131_,
    new_n28132_, new_n28133_, new_n28134_, new_n28135_, new_n28136_,
    new_n28137_, new_n28138_, new_n28139_, new_n28140_, new_n28141_,
    new_n28142_, new_n28143_, new_n28144_, new_n28145_, new_n28146_,
    new_n28147_, new_n28148_, new_n28149_, new_n28150_, new_n28151_,
    new_n28152_, new_n28153_, new_n28154_, new_n28155_, new_n28156_,
    new_n28157_, new_n28158_, new_n28159_, new_n28161_, new_n28162_,
    new_n28163_, new_n28164_, new_n28165_, new_n28166_, new_n28167_,
    new_n28168_, new_n28169_, new_n28170_, new_n28171_, new_n28172_,
    new_n28173_, new_n28174_, new_n28175_, new_n28176_, new_n28177_,
    new_n28178_, new_n28179_, new_n28180_, new_n28181_, new_n28182_,
    new_n28183_, new_n28184_, new_n28185_, new_n28186_, new_n28187_,
    new_n28188_, new_n28189_, new_n28190_, new_n28191_, new_n28192_,
    new_n28193_, new_n28194_, new_n28195_, new_n28196_, new_n28197_,
    new_n28198_, new_n28199_, new_n28200_, new_n28201_, new_n28202_,
    new_n28203_, new_n28204_, new_n28205_, new_n28206_, new_n28207_,
    new_n28208_, new_n28209_, new_n28210_, new_n28211_, new_n28212_,
    new_n28213_, new_n28214_, new_n28215_, new_n28217_, new_n28218_,
    new_n28219_, new_n28220_, new_n28221_, new_n28222_, new_n28223_,
    new_n28224_, new_n28225_, new_n28226_, new_n28227_, new_n28228_,
    new_n28229_, new_n28230_, new_n28231_, new_n28232_, new_n28233_,
    new_n28234_, new_n28235_, new_n28236_, new_n28237_, new_n28238_,
    new_n28239_, new_n28240_, new_n28241_, new_n28242_, new_n28243_,
    new_n28244_, new_n28245_, new_n28246_, new_n28247_, new_n28248_,
    new_n28249_, new_n28250_, new_n28251_, new_n28252_, new_n28253_,
    new_n28254_, new_n28255_, new_n28256_;
  INV_X1     g00000(.I(\a[5] ), .ZN(new_n65_));
  NAND4_X1   g00001(.A1(\a[23] ), .A2(\a[24] ), .A3(\a[25] ), .A4(\a[26] ), .ZN(new_n66_));
  INV_X1     g00002(.I(\a[28] ), .ZN(new_n67_));
  INV_X1     g00003(.I(\a[30] ), .ZN(new_n68_));
  NAND4_X1   g00004(.A1(new_n67_), .A2(new_n68_), .A3(\a[27] ), .A4(\a[29] ), .ZN(new_n69_));
  NOR2_X1    g00005(.A1(new_n69_), .A2(new_n66_), .ZN(new_n70_));
  INV_X1     g00006(.I(\a[24] ), .ZN(new_n71_));
  INV_X1     g00007(.I(\a[26] ), .ZN(new_n72_));
  NAND4_X1   g00008(.A1(new_n71_), .A2(new_n72_), .A3(\a[23] ), .A4(\a[25] ), .ZN(new_n73_));
  INV_X1     g00009(.I(\a[29] ), .ZN(new_n74_));
  NAND4_X1   g00010(.A1(new_n67_), .A2(new_n74_), .A3(\a[27] ), .A4(\a[30] ), .ZN(new_n75_));
  NOR2_X1    g00011(.A1(new_n73_), .A2(new_n75_), .ZN(new_n76_));
  NOR4_X1    g00012(.A1(new_n74_), .A2(\a[27] ), .A3(\a[28] ), .A4(\a[30] ), .ZN(new_n77_));
  INV_X1     g00013(.I(\a[25] ), .ZN(new_n78_));
  NOR4_X1    g00014(.A1(new_n71_), .A2(new_n78_), .A3(new_n72_), .A4(\a[23] ), .ZN(new_n79_));
  NAND2_X1   g00015(.A1(new_n79_), .A2(new_n77_), .ZN(new_n80_));
  INV_X1     g00016(.I(new_n80_), .ZN(new_n81_));
  INV_X1     g00017(.I(\a[27] ), .ZN(new_n82_));
  NAND4_X1   g00018(.A1(new_n82_), .A2(new_n68_), .A3(\a[28] ), .A4(\a[29] ), .ZN(new_n83_));
  INV_X1     g00019(.I(\a[23] ), .ZN(new_n84_));
  NAND4_X1   g00020(.A1(new_n84_), .A2(new_n78_), .A3(\a[24] ), .A4(\a[26] ), .ZN(new_n85_));
  NOR2_X1    g00021(.A1(new_n83_), .A2(new_n85_), .ZN(new_n86_));
  NOR4_X1    g00022(.A1(new_n81_), .A2(new_n70_), .A3(new_n76_), .A4(new_n86_), .ZN(new_n87_));
  NAND4_X1   g00023(.A1(new_n84_), .A2(\a[24] ), .A3(\a[25] ), .A4(\a[26] ), .ZN(new_n88_));
  NAND4_X1   g00024(.A1(new_n74_), .A2(new_n68_), .A3(\a[27] ), .A4(\a[28] ), .ZN(new_n89_));
  NOR2_X1    g00025(.A1(new_n89_), .A2(new_n88_), .ZN(new_n90_));
  NAND4_X1   g00026(.A1(new_n67_), .A2(\a[27] ), .A3(\a[29] ), .A4(\a[30] ), .ZN(new_n91_));
  NOR2_X1    g00027(.A1(new_n91_), .A2(new_n66_), .ZN(new_n92_));
  NOR2_X1    g00028(.A1(new_n90_), .A2(new_n92_), .ZN(new_n93_));
  INV_X1     g00029(.I(new_n93_), .ZN(new_n94_));
  NAND4_X1   g00030(.A1(new_n78_), .A2(new_n72_), .A3(\a[23] ), .A4(\a[24] ), .ZN(new_n95_));
  NOR2_X1    g00031(.A1(\a[27] ), .A2(\a[28] ), .ZN(new_n96_));
  NAND3_X1   g00032(.A1(new_n96_), .A2(new_n74_), .A3(\a[30] ), .ZN(new_n97_));
  NOR2_X1    g00033(.A1(new_n97_), .A2(new_n95_), .ZN(new_n98_));
  NOR2_X1    g00034(.A1(new_n78_), .A2(\a[26] ), .ZN(new_n99_));
  NOR2_X1    g00035(.A1(\a[23] ), .A2(\a[24] ), .ZN(new_n100_));
  NAND2_X1   g00036(.A1(new_n99_), .A2(new_n100_), .ZN(new_n101_));
  NOR2_X1    g00037(.A1(new_n101_), .A2(new_n97_), .ZN(new_n102_));
  NOR2_X1    g00038(.A1(new_n102_), .A2(new_n98_), .ZN(new_n103_));
  INV_X1     g00039(.I(new_n103_), .ZN(new_n104_));
  NAND4_X1   g00040(.A1(new_n84_), .A2(new_n71_), .A3(\a[25] ), .A4(\a[26] ), .ZN(new_n105_));
  NOR2_X1    g00041(.A1(new_n75_), .A2(new_n105_), .ZN(new_n106_));
  NOR4_X1    g00042(.A1(new_n87_), .A2(new_n104_), .A3(new_n94_), .A4(new_n106_), .ZN(new_n107_));
  NOR4_X1    g00043(.A1(new_n78_), .A2(\a[23] ), .A3(\a[24] ), .A4(\a[26] ), .ZN(new_n108_));
  AND4_X2    g00044(.A1(\a[27] ), .A2(\a[28] ), .A3(\a[29] ), .A4(\a[30] ), .Z(new_n109_));
  NAND2_X1   g00045(.A1(new_n109_), .A2(new_n108_), .ZN(new_n110_));
  NOR4_X1    g00046(.A1(new_n82_), .A2(new_n67_), .A3(new_n68_), .A4(\a[29] ), .ZN(new_n111_));
  NOR4_X1    g00047(.A1(new_n71_), .A2(new_n78_), .A3(\a[23] ), .A4(\a[26] ), .ZN(new_n112_));
  NAND2_X1   g00048(.A1(new_n111_), .A2(new_n112_), .ZN(new_n113_));
  NAND2_X1   g00049(.A1(new_n113_), .A2(new_n110_), .ZN(new_n114_));
  NAND4_X1   g00050(.A1(new_n71_), .A2(new_n78_), .A3(\a[23] ), .A4(\a[26] ), .ZN(new_n115_));
  NAND4_X1   g00051(.A1(new_n82_), .A2(new_n74_), .A3(\a[28] ), .A4(\a[30] ), .ZN(new_n116_));
  NOR2_X1    g00052(.A1(new_n115_), .A2(new_n116_), .ZN(new_n117_));
  NAND4_X1   g00053(.A1(new_n71_), .A2(new_n78_), .A3(new_n72_), .A4(\a[23] ), .ZN(new_n118_));
  NOR2_X1    g00054(.A1(new_n118_), .A2(new_n75_), .ZN(new_n119_));
  NOR2_X1    g00055(.A1(new_n117_), .A2(new_n119_), .ZN(new_n120_));
  INV_X1     g00056(.I(new_n120_), .ZN(new_n121_));
  NAND4_X1   g00057(.A1(new_n71_), .A2(\a[23] ), .A3(\a[25] ), .A4(\a[26] ), .ZN(new_n122_));
  NAND4_X1   g00058(.A1(new_n82_), .A2(\a[28] ), .A3(\a[29] ), .A4(\a[30] ), .ZN(new_n123_));
  NOR2_X1    g00059(.A1(new_n122_), .A2(new_n123_), .ZN(new_n124_));
  NOR2_X1    g00060(.A1(new_n83_), .A2(new_n66_), .ZN(new_n125_));
  NOR2_X1    g00061(.A1(new_n124_), .A2(new_n125_), .ZN(new_n126_));
  INV_X1     g00062(.I(new_n126_), .ZN(new_n127_));
  NOR3_X1    g00063(.A1(new_n121_), .A2(new_n127_), .A3(new_n114_), .ZN(new_n128_));
  NAND4_X1   g00064(.A1(new_n74_), .A2(\a[27] ), .A3(\a[28] ), .A4(\a[30] ), .ZN(new_n129_));
  NOR2_X1    g00065(.A1(new_n118_), .A2(new_n129_), .ZN(new_n130_));
  NAND4_X1   g00066(.A1(new_n82_), .A2(new_n67_), .A3(\a[29] ), .A4(\a[30] ), .ZN(new_n131_));
  NOR2_X1    g00067(.A1(new_n131_), .A2(new_n66_), .ZN(new_n132_));
  NAND4_X1   g00068(.A1(new_n84_), .A2(new_n72_), .A3(\a[24] ), .A4(\a[25] ), .ZN(new_n133_));
  NAND4_X1   g00069(.A1(new_n67_), .A2(new_n74_), .A3(new_n68_), .A4(\a[27] ), .ZN(new_n134_));
  NOR2_X1    g00070(.A1(new_n134_), .A2(new_n133_), .ZN(new_n135_));
  NOR2_X1    g00071(.A1(new_n105_), .A2(new_n123_), .ZN(new_n136_));
  NOR2_X1    g00072(.A1(new_n118_), .A2(new_n97_), .ZN(new_n137_));
  NOR2_X1    g00073(.A1(new_n137_), .A2(new_n136_), .ZN(new_n138_));
  NOR4_X1    g00074(.A1(new_n71_), .A2(new_n72_), .A3(\a[23] ), .A4(\a[25] ), .ZN(new_n139_));
  NOR4_X1    g00075(.A1(new_n74_), .A2(new_n68_), .A3(\a[27] ), .A4(\a[28] ), .ZN(new_n140_));
  NAND2_X1   g00076(.A1(new_n139_), .A2(new_n140_), .ZN(new_n141_));
  NOR4_X1    g00077(.A1(new_n82_), .A2(new_n68_), .A3(\a[28] ), .A4(\a[29] ), .ZN(new_n142_));
  NOR4_X1    g00078(.A1(new_n72_), .A2(\a[23] ), .A3(\a[24] ), .A4(\a[25] ), .ZN(new_n143_));
  NAND2_X1   g00079(.A1(new_n142_), .A2(new_n143_), .ZN(new_n144_));
  NAND3_X1   g00080(.A1(new_n138_), .A2(new_n141_), .A3(new_n144_), .ZN(new_n145_));
  NOR4_X1    g00081(.A1(new_n145_), .A2(new_n130_), .A3(new_n132_), .A4(new_n135_), .ZN(new_n146_));
  NOR2_X1    g00082(.A1(new_n101_), .A2(new_n131_), .ZN(new_n147_));
  NAND4_X1   g00083(.A1(new_n72_), .A2(\a[23] ), .A3(\a[24] ), .A4(\a[25] ), .ZN(new_n148_));
  NOR2_X1    g00084(.A1(new_n134_), .A2(new_n148_), .ZN(new_n149_));
  NAND4_X1   g00085(.A1(\a[27] ), .A2(\a[28] ), .A3(\a[29] ), .A4(\a[30] ), .ZN(new_n150_));
  NAND4_X1   g00086(.A1(new_n78_), .A2(\a[23] ), .A3(\a[24] ), .A4(\a[26] ), .ZN(new_n151_));
  NOR2_X1    g00087(.A1(new_n151_), .A2(new_n150_), .ZN(new_n152_));
  NOR4_X1    g00088(.A1(\a[23] ), .A2(\a[24] ), .A3(\a[25] ), .A4(\a[26] ), .ZN(new_n153_));
  NOR2_X1    g00089(.A1(new_n123_), .A2(new_n153_), .ZN(new_n154_));
  NOR4_X1    g00090(.A1(new_n147_), .A2(new_n149_), .A3(new_n152_), .A4(new_n154_), .ZN(new_n155_));
  NOR4_X1    g00091(.A1(new_n82_), .A2(new_n67_), .A3(\a[29] ), .A4(\a[30] ), .ZN(new_n156_));
  NAND2_X1   g00092(.A1(new_n156_), .A2(new_n108_), .ZN(new_n157_));
  NOR4_X1    g00093(.A1(new_n84_), .A2(new_n71_), .A3(new_n72_), .A4(\a[25] ), .ZN(new_n158_));
  NOR4_X1    g00094(.A1(new_n82_), .A2(new_n67_), .A3(new_n74_), .A4(\a[30] ), .ZN(new_n159_));
  NAND2_X1   g00095(.A1(new_n158_), .A2(new_n159_), .ZN(new_n160_));
  NAND2_X1   g00096(.A1(new_n160_), .A2(new_n157_), .ZN(new_n161_));
  INV_X1     g00097(.I(new_n161_), .ZN(new_n162_));
  NOR2_X1    g00098(.A1(new_n91_), .A2(new_n153_), .ZN(new_n163_));
  NOR2_X1    g00099(.A1(new_n129_), .A2(new_n151_), .ZN(new_n164_));
  NOR2_X1    g00100(.A1(new_n164_), .A2(new_n163_), .ZN(new_n165_));
  NAND2_X1   g00101(.A1(new_n162_), .A2(new_n165_), .ZN(new_n166_));
  NOR2_X1    g00102(.A1(new_n166_), .A2(new_n155_), .ZN(new_n167_));
  NAND4_X1   g00103(.A1(new_n167_), .A2(new_n107_), .A3(new_n146_), .A4(new_n128_), .ZN(new_n168_));
  NAND4_X1   g00104(.A1(new_n68_), .A2(\a[27] ), .A3(\a[28] ), .A4(\a[29] ), .ZN(new_n169_));
  NOR2_X1    g00105(.A1(new_n122_), .A2(new_n169_), .ZN(new_n170_));
  NAND4_X1   g00106(.A1(new_n82_), .A2(new_n74_), .A3(new_n68_), .A4(\a[28] ), .ZN(new_n171_));
  NOR2_X1    g00107(.A1(new_n171_), .A2(new_n153_), .ZN(new_n172_));
  NOR2_X1    g00108(.A1(new_n171_), .A2(new_n151_), .ZN(new_n173_));
  NOR3_X1    g00109(.A1(new_n172_), .A2(new_n173_), .A3(new_n170_), .ZN(new_n174_));
  NAND3_X1   g00110(.A1(new_n96_), .A2(\a[29] ), .A3(new_n68_), .ZN(new_n175_));
  NAND3_X1   g00111(.A1(new_n100_), .A2(new_n78_), .A3(\a[26] ), .ZN(new_n176_));
  AOI21_X1   g00112(.A1(new_n101_), .A2(new_n176_), .B(new_n175_), .ZN(new_n177_));
  AOI21_X1   g00113(.A1(new_n73_), .A2(new_n148_), .B(new_n169_), .ZN(new_n178_));
  NOR2_X1    g00114(.A1(new_n177_), .A2(new_n178_), .ZN(new_n179_));
  NOR4_X1    g00115(.A1(new_n82_), .A2(new_n74_), .A3(\a[28] ), .A4(\a[30] ), .ZN(new_n180_));
  NAND3_X1   g00116(.A1(new_n100_), .A2(new_n78_), .A3(new_n72_), .ZN(new_n181_));
  NAND2_X1   g00117(.A1(new_n180_), .A2(new_n181_), .ZN(new_n182_));
  NOR2_X1    g00118(.A1(new_n133_), .A2(new_n91_), .ZN(new_n183_));
  INV_X1     g00119(.I(new_n183_), .ZN(new_n184_));
  NOR4_X1    g00120(.A1(new_n67_), .A2(new_n68_), .A3(\a[27] ), .A4(\a[29] ), .ZN(new_n185_));
  NOR4_X1    g00121(.A1(new_n84_), .A2(\a[24] ), .A3(\a[25] ), .A4(\a[26] ), .ZN(new_n186_));
  NAND2_X1   g00122(.A1(new_n185_), .A2(new_n186_), .ZN(new_n187_));
  NAND2_X1   g00123(.A1(new_n180_), .A2(new_n143_), .ZN(new_n188_));
  NAND4_X1   g00124(.A1(new_n184_), .A2(new_n182_), .A3(new_n187_), .A4(new_n188_), .ZN(new_n189_));
  NOR2_X1    g00125(.A1(new_n115_), .A2(new_n91_), .ZN(new_n190_));
  NOR2_X1    g00126(.A1(new_n89_), .A2(new_n151_), .ZN(new_n191_));
  NOR2_X1    g00127(.A1(new_n97_), .A2(new_n88_), .ZN(new_n192_));
  NOR3_X1    g00128(.A1(new_n190_), .A2(new_n192_), .A3(new_n191_), .ZN(new_n193_));
  NAND4_X1   g00129(.A1(new_n189_), .A2(new_n179_), .A3(new_n174_), .A4(new_n193_), .ZN(new_n194_));
  OR2_X2     g00130(.A1(new_n168_), .A2(new_n194_), .Z(new_n195_));
  NOR4_X1    g00131(.A1(new_n67_), .A2(new_n74_), .A3(\a[27] ), .A4(\a[30] ), .ZN(new_n196_));
  NAND2_X1   g00132(.A1(new_n196_), .A2(new_n108_), .ZN(new_n197_));
  NOR2_X1    g00133(.A1(new_n97_), .A2(new_n176_), .ZN(new_n198_));
  INV_X1     g00134(.I(new_n198_), .ZN(new_n199_));
  NAND2_X1   g00135(.A1(new_n199_), .A2(new_n197_), .ZN(new_n200_));
  INV_X1     g00136(.I(new_n200_), .ZN(new_n201_));
  NOR2_X1    g00137(.A1(new_n134_), .A2(new_n73_), .ZN(new_n202_));
  NOR2_X1    g00138(.A1(new_n97_), .A2(new_n105_), .ZN(new_n203_));
  NOR2_X1    g00139(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR4_X1    g00140(.A1(new_n84_), .A2(new_n71_), .A3(new_n78_), .A4(\a[26] ), .ZN(new_n205_));
  NOR4_X1    g00141(.A1(new_n67_), .A2(\a[27] ), .A3(\a[29] ), .A4(\a[30] ), .ZN(new_n206_));
  NAND2_X1   g00142(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1   g00143(.A1(new_n111_), .A2(new_n143_), .ZN(new_n208_));
  NAND3_X1   g00144(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1   g00145(.A1(new_n201_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1    g00146(.A1(new_n171_), .A2(new_n105_), .ZN(new_n211_));
  NOR2_X1    g00147(.A1(new_n118_), .A2(new_n171_), .ZN(new_n212_));
  NOR2_X1    g00148(.A1(new_n118_), .A2(new_n83_), .ZN(new_n213_));
  NOR2_X1    g00149(.A1(new_n69_), .A2(new_n73_), .ZN(new_n214_));
  NOR4_X1    g00150(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  NOR2_X1    g00151(.A1(new_n69_), .A2(new_n122_), .ZN(new_n216_));
  NOR2_X1    g00152(.A1(new_n118_), .A2(new_n175_), .ZN(new_n217_));
  NOR2_X1    g00153(.A1(new_n217_), .A2(new_n216_), .ZN(new_n218_));
  NOR2_X1    g00154(.A1(new_n97_), .A2(new_n85_), .ZN(new_n219_));
  INV_X1     g00155(.I(new_n219_), .ZN(new_n220_));
  NAND2_X1   g00156(.A1(new_n139_), .A2(new_n77_), .ZN(new_n221_));
  NAND2_X1   g00157(.A1(new_n109_), .A2(new_n186_), .ZN(new_n222_));
  NAND4_X1   g00158(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  NOR3_X1    g00159(.A1(new_n210_), .A2(new_n223_), .A3(new_n215_), .ZN(new_n224_));
  NOR2_X1    g00160(.A1(new_n171_), .A2(new_n85_), .ZN(new_n225_));
  NOR2_X1    g00161(.A1(new_n95_), .A2(new_n129_), .ZN(new_n226_));
  NOR2_X1    g00162(.A1(new_n91_), .A2(new_n122_), .ZN(new_n227_));
  NOR3_X1    g00163(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1     g00164(.I(new_n228_), .ZN(new_n229_));
  NOR4_X1    g00165(.A1(new_n78_), .A2(new_n72_), .A3(\a[23] ), .A4(\a[24] ), .ZN(new_n230_));
  NAND2_X1   g00166(.A1(new_n196_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1    g00167(.A1(new_n175_), .A2(new_n151_), .ZN(new_n232_));
  INV_X1     g00168(.I(new_n232_), .ZN(new_n233_));
  NAND2_X1   g00169(.A1(new_n233_), .A2(new_n231_), .ZN(new_n234_));
  NOR2_X1    g00170(.A1(new_n134_), .A2(new_n66_), .ZN(new_n235_));
  NOR2_X1    g00171(.A1(new_n131_), .A2(new_n122_), .ZN(new_n236_));
  NOR3_X1    g00172(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NOR2_X1    g00173(.A1(new_n115_), .A2(new_n131_), .ZN(new_n238_));
  NOR2_X1    g00174(.A1(new_n171_), .A2(new_n73_), .ZN(new_n239_));
  NOR4_X1    g00175(.A1(new_n237_), .A2(new_n229_), .A3(new_n238_), .A4(new_n239_), .ZN(new_n240_));
  NOR2_X1    g00176(.A1(new_n118_), .A2(new_n169_), .ZN(new_n241_));
  NOR2_X1    g00177(.A1(new_n95_), .A2(new_n169_), .ZN(new_n242_));
  NOR2_X1    g00178(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1     g00179(.I(new_n243_), .ZN(new_n244_));
  NOR4_X1    g00180(.A1(new_n84_), .A2(new_n72_), .A3(\a[24] ), .A4(\a[25] ), .ZN(new_n245_));
  NAND2_X1   g00181(.A1(new_n159_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1    g00182(.A1(new_n69_), .A2(new_n95_), .ZN(new_n247_));
  INV_X1     g00183(.I(new_n247_), .ZN(new_n248_));
  NAND2_X1   g00184(.A1(new_n248_), .A2(new_n246_), .ZN(new_n249_));
  NAND2_X1   g00185(.A1(new_n185_), .A2(new_n108_), .ZN(new_n250_));
  INV_X1     g00186(.I(new_n250_), .ZN(new_n251_));
  NOR2_X1    g00187(.A1(new_n134_), .A2(new_n176_), .ZN(new_n252_));
  NOR2_X1    g00188(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1     g00189(.I(new_n253_), .ZN(new_n254_));
  NOR2_X1    g00190(.A1(new_n105_), .A2(new_n131_), .ZN(new_n255_));
  NOR2_X1    g00191(.A1(new_n95_), .A2(new_n123_), .ZN(new_n256_));
  NOR2_X1    g00192(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1     g00193(.I(new_n257_), .ZN(new_n258_));
  NOR4_X1    g00194(.A1(new_n254_), .A2(new_n244_), .A3(new_n258_), .A4(new_n249_), .ZN(new_n259_));
  NOR2_X1    g00195(.A1(new_n134_), .A2(new_n115_), .ZN(new_n260_));
  NOR2_X1    g00196(.A1(new_n105_), .A2(new_n91_), .ZN(new_n261_));
  NOR2_X1    g00197(.A1(new_n105_), .A2(new_n129_), .ZN(new_n262_));
  NOR3_X1    g00198(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NOR2_X1    g00199(.A1(new_n148_), .A2(new_n150_), .ZN(new_n264_));
  NOR4_X1    g00200(.A1(new_n84_), .A2(new_n71_), .A3(\a[25] ), .A4(\a[26] ), .ZN(new_n265_));
  NAND2_X1   g00201(.A1(new_n265_), .A2(new_n109_), .ZN(new_n266_));
  INV_X1     g00202(.I(new_n266_), .ZN(new_n267_));
  NOR2_X1    g00203(.A1(new_n176_), .A2(new_n150_), .ZN(new_n268_));
  NOR3_X1    g00204(.A1(new_n267_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n269_));
  AND4_X2    g00205(.A1(\a[23] ), .A2(\a[24] ), .A3(\a[25] ), .A4(\a[26] ), .Z(new_n270_));
  NAND2_X1   g00206(.A1(new_n142_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1   g00207(.A1(new_n156_), .A2(new_n181_), .ZN(new_n272_));
  NOR4_X1    g00208(.A1(new_n71_), .A2(\a[23] ), .A3(\a[25] ), .A4(\a[26] ), .ZN(new_n273_));
  NAND2_X1   g00209(.A1(new_n77_), .A2(new_n273_), .ZN(new_n274_));
  NOR4_X1    g00210(.A1(new_n67_), .A2(new_n74_), .A3(new_n68_), .A4(\a[27] ), .ZN(new_n275_));
  NAND2_X1   g00211(.A1(new_n275_), .A2(new_n112_), .ZN(new_n276_));
  NAND4_X1   g00212(.A1(new_n271_), .A2(new_n272_), .A3(new_n276_), .A4(new_n274_), .ZN(new_n277_));
  AND3_X2    g00213(.A1(new_n269_), .A2(new_n263_), .A3(new_n277_), .Z(new_n278_));
  NAND4_X1   g00214(.A1(new_n224_), .A2(new_n240_), .A3(new_n259_), .A4(new_n278_), .ZN(new_n279_));
  NOR2_X1    g00215(.A1(new_n169_), .A2(new_n66_), .ZN(new_n280_));
  NOR2_X1    g00216(.A1(new_n176_), .A2(new_n83_), .ZN(new_n281_));
  NOR2_X1    g00217(.A1(new_n134_), .A2(new_n88_), .ZN(new_n282_));
  NOR3_X1    g00218(.A1(new_n281_), .A2(new_n282_), .A3(new_n280_), .ZN(new_n283_));
  NOR4_X1    g00219(.A1(new_n84_), .A2(new_n78_), .A3(\a[24] ), .A4(\a[26] ), .ZN(new_n284_));
  OAI21_X1   g00220(.A1(new_n205_), .A2(new_n284_), .B(new_n77_), .ZN(new_n285_));
  NOR2_X1    g00221(.A1(new_n95_), .A2(new_n91_), .ZN(new_n286_));
  INV_X1     g00222(.I(new_n286_), .ZN(new_n287_));
  NOR2_X1    g00223(.A1(new_n75_), .A2(new_n85_), .ZN(new_n288_));
  NOR2_X1    g00224(.A1(new_n176_), .A2(new_n89_), .ZN(new_n289_));
  NOR2_X1    g00225(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND4_X1   g00226(.A1(new_n283_), .A2(new_n290_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n291_));
  NAND2_X1   g00227(.A1(new_n205_), .A2(new_n140_), .ZN(new_n292_));
  NAND2_X1   g00228(.A1(new_n142_), .A2(new_n265_), .ZN(new_n293_));
  NOR2_X1    g00229(.A1(new_n89_), .A2(new_n95_), .ZN(new_n294_));
  INV_X1     g00230(.I(new_n294_), .ZN(new_n295_));
  NAND3_X1   g00231(.A1(new_n295_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n296_));
  NOR2_X1    g00232(.A1(new_n171_), .A2(new_n66_), .ZN(new_n297_));
  NOR2_X1    g00233(.A1(new_n115_), .A2(new_n129_), .ZN(new_n298_));
  NOR2_X1    g00234(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1     g00235(.I(new_n299_), .ZN(new_n300_));
  NAND2_X1   g00236(.A1(new_n181_), .A2(new_n109_), .ZN(new_n301_));
  NAND2_X1   g00237(.A1(new_n112_), .A2(new_n206_), .ZN(new_n302_));
  NAND3_X1   g00238(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  NOR2_X1    g00239(.A1(new_n133_), .A2(new_n116_), .ZN(new_n304_));
  NOR2_X1    g00240(.A1(new_n83_), .A2(new_n133_), .ZN(new_n305_));
  NOR2_X1    g00241(.A1(new_n89_), .A2(new_n66_), .ZN(new_n306_));
  NOR2_X1    g00242(.A1(new_n97_), .A2(new_n66_), .ZN(new_n307_));
  NOR4_X1    g00243(.A1(new_n304_), .A2(new_n305_), .A3(new_n307_), .A4(new_n306_), .ZN(new_n308_));
  NAND2_X1   g00244(.A1(new_n111_), .A2(new_n181_), .ZN(new_n309_));
  NOR2_X1    g00245(.A1(new_n66_), .A2(new_n150_), .ZN(new_n310_));
  INV_X1     g00246(.I(new_n310_), .ZN(new_n311_));
  NOR2_X1    g00247(.A1(new_n97_), .A2(new_n133_), .ZN(new_n312_));
  INV_X1     g00248(.I(new_n312_), .ZN(new_n313_));
  NAND3_X1   g00249(.A1(new_n313_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n314_));
  NOR4_X1    g00250(.A1(new_n303_), .A2(new_n296_), .A3(new_n314_), .A4(new_n308_), .ZN(new_n315_));
  OAI22_X1   g00251(.A1(new_n69_), .A2(new_n85_), .B1(new_n116_), .B2(new_n88_), .ZN(new_n316_));
  INV_X1     g00252(.I(new_n316_), .ZN(new_n317_));
  NOR4_X1    g00253(.A1(new_n84_), .A2(new_n78_), .A3(new_n72_), .A4(\a[24] ), .ZN(new_n318_));
  NAND2_X1   g00254(.A1(new_n318_), .A2(new_n77_), .ZN(new_n319_));
  NOR2_X1    g00255(.A1(new_n115_), .A2(new_n123_), .ZN(new_n320_));
  INV_X1     g00256(.I(new_n320_), .ZN(new_n321_));
  NAND2_X1   g00257(.A1(new_n79_), .A2(new_n111_), .ZN(new_n322_));
  NAND4_X1   g00258(.A1(new_n317_), .A2(new_n321_), .A3(new_n319_), .A4(new_n322_), .ZN(new_n323_));
  NOR2_X1    g00259(.A1(new_n116_), .A2(new_n151_), .ZN(new_n324_));
  NAND2_X1   g00260(.A1(new_n140_), .A2(new_n186_), .ZN(new_n325_));
  INV_X1     g00261(.I(new_n325_), .ZN(new_n326_));
  NOR2_X1    g00262(.A1(new_n326_), .A2(new_n324_), .ZN(new_n327_));
  INV_X1     g00263(.I(new_n327_), .ZN(new_n328_));
  NOR2_X1    g00264(.A1(new_n88_), .A2(new_n150_), .ZN(new_n329_));
  NOR2_X1    g00265(.A1(new_n89_), .A2(new_n148_), .ZN(new_n330_));
  NOR2_X1    g00266(.A1(new_n330_), .A2(new_n329_), .ZN(new_n331_));
  INV_X1     g00267(.I(new_n331_), .ZN(new_n332_));
  NOR2_X1    g00268(.A1(new_n85_), .A2(new_n123_), .ZN(new_n333_));
  NAND4_X1   g00269(.A1(new_n84_), .A2(new_n78_), .A3(new_n72_), .A4(\a[24] ), .ZN(new_n334_));
  NOR2_X1    g00270(.A1(new_n334_), .A2(new_n123_), .ZN(new_n335_));
  NOR2_X1    g00271(.A1(new_n335_), .A2(new_n333_), .ZN(new_n336_));
  INV_X1     g00272(.I(new_n336_), .ZN(new_n337_));
  NOR4_X1    g00273(.A1(new_n323_), .A2(new_n328_), .A3(new_n332_), .A4(new_n337_), .ZN(new_n338_));
  NAND2_X1   g00274(.A1(new_n315_), .A2(new_n338_), .ZN(new_n339_));
  OR3_X2     g00275(.A1(new_n279_), .A2(new_n291_), .A3(new_n339_), .Z(new_n340_));
  NOR2_X1    g00276(.A1(new_n340_), .A2(new_n195_), .ZN(new_n341_));
  NAND2_X1   g00277(.A1(new_n159_), .A2(new_n112_), .ZN(new_n342_));
  INV_X1     g00278(.I(new_n342_), .ZN(new_n343_));
  NOR2_X1    g00279(.A1(new_n343_), .A2(new_n178_), .ZN(new_n344_));
  NOR2_X1    g00280(.A1(new_n171_), .A2(new_n122_), .ZN(new_n345_));
  NOR4_X1    g00281(.A1(\a[27] ), .A2(\a[28] ), .A3(\a[29] ), .A4(\a[30] ), .ZN(new_n346_));
  NOR2_X1    g00282(.A1(new_n73_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1    g00283(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1   g00284(.A1(new_n186_), .A2(new_n206_), .ZN(new_n349_));
  NOR4_X1    g00285(.A1(new_n82_), .A2(\a[28] ), .A3(\a[29] ), .A4(\a[30] ), .ZN(new_n350_));
  NAND2_X1   g00286(.A1(new_n79_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1    g00287(.A1(new_n85_), .A2(new_n129_), .ZN(new_n352_));
  INV_X1     g00288(.I(new_n352_), .ZN(new_n353_));
  NOR2_X1    g00289(.A1(\a[29] ), .A2(\a[30] ), .ZN(new_n354_));
  NAND2_X1   g00290(.A1(new_n96_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1   g00291(.A1(new_n355_), .A2(new_n143_), .ZN(new_n356_));
  NAND4_X1   g00292(.A1(new_n353_), .A2(new_n349_), .A3(new_n351_), .A4(new_n356_), .ZN(new_n357_));
  INV_X1     g00293(.I(new_n226_), .ZN(new_n358_));
  NOR2_X1    g00294(.A1(new_n69_), .A2(new_n88_), .ZN(new_n359_));
  INV_X1     g00295(.I(new_n359_), .ZN(new_n360_));
  NAND2_X1   g00296(.A1(new_n196_), .A2(new_n265_), .ZN(new_n361_));
  NAND2_X1   g00297(.A1(new_n159_), .A2(new_n108_), .ZN(new_n362_));
  NAND4_X1   g00298(.A1(new_n360_), .A2(new_n358_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  NAND4_X1   g00299(.A1(new_n363_), .A2(new_n357_), .A3(new_n344_), .A4(new_n348_), .ZN(new_n364_));
  INV_X1     g00300(.I(new_n197_), .ZN(new_n365_));
  NOR2_X1    g00301(.A1(new_n69_), .A2(new_n85_), .ZN(new_n366_));
  NOR2_X1    g00302(.A1(new_n118_), .A2(new_n69_), .ZN(new_n367_));
  NOR2_X1    g00303(.A1(new_n367_), .A2(new_n125_), .ZN(new_n368_));
  INV_X1     g00304(.I(new_n368_), .ZN(new_n369_));
  NOR2_X1    g00305(.A1(new_n83_), .A2(new_n88_), .ZN(new_n370_));
  NOR4_X1    g00306(.A1(new_n369_), .A2(new_n365_), .A3(new_n366_), .A4(new_n370_), .ZN(new_n371_));
  INV_X1     g00307(.I(new_n371_), .ZN(new_n372_));
  NAND2_X1   g00308(.A1(new_n275_), .A2(new_n230_), .ZN(new_n373_));
  NOR2_X1    g00309(.A1(new_n88_), .A2(new_n123_), .ZN(new_n374_));
  NOR2_X1    g00310(.A1(new_n374_), .A2(new_n329_), .ZN(new_n375_));
  NOR2_X1    g00311(.A1(new_n122_), .A2(new_n150_), .ZN(new_n376_));
  INV_X1     g00312(.I(new_n376_), .ZN(new_n377_));
  NAND2_X1   g00313(.A1(new_n245_), .A2(new_n109_), .ZN(new_n378_));
  NAND4_X1   g00314(.A1(new_n375_), .A2(new_n373_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  NOR3_X1    g00315(.A1(new_n372_), .A2(new_n364_), .A3(new_n379_), .ZN(new_n380_));
  NOR2_X1    g00316(.A1(new_n176_), .A2(new_n116_), .ZN(new_n381_));
  INV_X1     g00317(.I(new_n381_), .ZN(new_n382_));
  NAND2_X1   g00318(.A1(new_n139_), .A2(new_n350_), .ZN(new_n383_));
  NOR2_X1    g00319(.A1(new_n123_), .A2(new_n148_), .ZN(new_n384_));
  INV_X1     g00320(.I(new_n384_), .ZN(new_n385_));
  NAND4_X1   g00321(.A1(new_n382_), .A2(new_n385_), .A3(new_n311_), .A4(new_n383_), .ZN(new_n386_));
  NOR2_X1    g00322(.A1(new_n75_), .A2(new_n95_), .ZN(new_n387_));
  NOR2_X1    g00323(.A1(new_n116_), .A2(new_n148_), .ZN(new_n388_));
  NOR2_X1    g00324(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1   g00325(.A1(new_n350_), .A2(new_n273_), .ZN(new_n390_));
  NAND2_X1   g00326(.A1(new_n355_), .A2(new_n139_), .ZN(new_n391_));
  NAND4_X1   g00327(.A1(new_n386_), .A2(new_n389_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n392_));
  NAND2_X1   g00328(.A1(new_n318_), .A2(new_n159_), .ZN(new_n393_));
  NAND2_X1   g00329(.A1(new_n156_), .A2(new_n270_), .ZN(new_n394_));
  NAND2_X1   g00330(.A1(new_n245_), .A2(new_n77_), .ZN(new_n395_));
  NOR2_X1    g00331(.A1(new_n175_), .A2(new_n73_), .ZN(new_n396_));
  NOR2_X1    g00332(.A1(new_n129_), .A2(new_n153_), .ZN(new_n397_));
  NOR2_X1    g00333(.A1(new_n175_), .A2(new_n95_), .ZN(new_n398_));
  NOR2_X1    g00334(.A1(new_n398_), .A2(new_n397_), .ZN(new_n399_));
  INV_X1     g00335(.I(new_n399_), .ZN(new_n400_));
  NOR3_X1    g00336(.A1(new_n400_), .A2(new_n130_), .A3(new_n396_), .ZN(new_n401_));
  NAND4_X1   g00337(.A1(new_n401_), .A2(new_n393_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n402_));
  NOR2_X1    g00338(.A1(new_n97_), .A2(new_n115_), .ZN(new_n403_));
  NOR4_X1    g00339(.A1(new_n82_), .A2(new_n74_), .A3(new_n68_), .A4(\a[28] ), .ZN(new_n404_));
  NAND2_X1   g00340(.A1(new_n404_), .A2(new_n143_), .ZN(new_n405_));
  INV_X1     g00341(.I(new_n405_), .ZN(new_n406_));
  NOR4_X1    g00342(.A1(new_n406_), .A2(new_n214_), .A3(new_n288_), .A4(new_n403_), .ZN(new_n407_));
  INV_X1     g00343(.I(new_n190_), .ZN(new_n408_));
  NAND2_X1   g00344(.A1(new_n142_), .A2(new_n108_), .ZN(new_n409_));
  NAND2_X1   g00345(.A1(new_n159_), .A2(new_n181_), .ZN(new_n410_));
  NAND3_X1   g00346(.A1(new_n408_), .A2(new_n410_), .A3(new_n409_), .ZN(new_n411_));
  NOR4_X1    g00347(.A1(new_n402_), .A2(new_n392_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n412_));
  NOR2_X1    g00348(.A1(new_n151_), .A2(new_n169_), .ZN(new_n413_));
  NAND2_X1   g00349(.A1(new_n180_), .A2(new_n273_), .ZN(new_n414_));
  INV_X1     g00350(.I(new_n414_), .ZN(new_n415_));
  NOR3_X1    g00351(.A1(new_n415_), .A2(new_n413_), .A3(new_n191_), .ZN(new_n416_));
  INV_X1     g00352(.I(new_n416_), .ZN(new_n417_));
  NOR2_X1    g00353(.A1(new_n116_), .A2(new_n66_), .ZN(new_n418_));
  NOR2_X1    g00354(.A1(new_n91_), .A2(new_n148_), .ZN(new_n419_));
  NOR2_X1    g00355(.A1(new_n131_), .A2(new_n151_), .ZN(new_n420_));
  NOR4_X1    g00356(.A1(new_n238_), .A2(new_n419_), .A3(new_n420_), .A4(new_n418_), .ZN(new_n421_));
  AOI21_X1   g00357(.A1(new_n85_), .A2(new_n105_), .B(new_n91_), .ZN(new_n422_));
  NAND2_X1   g00358(.A1(new_n230_), .A2(new_n109_), .ZN(new_n423_));
  INV_X1     g00359(.I(new_n423_), .ZN(new_n424_));
  NOR2_X1    g00360(.A1(new_n424_), .A2(new_n304_), .ZN(new_n425_));
  INV_X1     g00361(.I(new_n425_), .ZN(new_n426_));
  NOR4_X1    g00362(.A1(new_n417_), .A2(new_n426_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n427_));
  NOR2_X1    g00363(.A1(new_n116_), .A2(new_n88_), .ZN(new_n428_));
  INV_X1     g00364(.I(new_n428_), .ZN(new_n429_));
  NOR2_X1    g00365(.A1(new_n83_), .A2(new_n153_), .ZN(new_n430_));
  INV_X1     g00366(.I(new_n430_), .ZN(new_n431_));
  NAND2_X1   g00367(.A1(new_n112_), .A2(new_n77_), .ZN(new_n432_));
  NAND4_X1   g00368(.A1(new_n295_), .A2(new_n429_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1   g00369(.A1(new_n111_), .A2(new_n230_), .ZN(new_n434_));
  NAND2_X1   g00370(.A1(new_n156_), .A2(new_n245_), .ZN(new_n435_));
  NAND2_X1   g00371(.A1(new_n79_), .A2(new_n142_), .ZN(new_n436_));
  NOR2_X1    g00372(.A1(new_n97_), .A2(new_n151_), .ZN(new_n437_));
  INV_X1     g00373(.I(new_n437_), .ZN(new_n438_));
  NAND4_X1   g00374(.A1(new_n438_), .A2(new_n434_), .A3(new_n435_), .A4(new_n436_), .ZN(new_n439_));
  NOR4_X1    g00375(.A1(new_n68_), .A2(\a[27] ), .A3(\a[28] ), .A4(\a[29] ), .ZN(new_n440_));
  NAND2_X1   g00376(.A1(new_n265_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1     g00377(.I(new_n333_), .ZN(new_n442_));
  NAND4_X1   g00378(.A1(new_n321_), .A2(new_n442_), .A3(new_n80_), .A4(new_n441_), .ZN(new_n443_));
  AND3_X2    g00379(.A1(new_n433_), .A2(new_n443_), .A3(new_n439_), .Z(new_n444_));
  NAND4_X1   g00380(.A1(new_n412_), .A2(new_n380_), .A3(new_n427_), .A4(new_n444_), .ZN(new_n445_));
  INV_X1     g00381(.I(new_n319_), .ZN(new_n446_));
  NOR2_X1    g00382(.A1(new_n73_), .A2(new_n116_), .ZN(new_n447_));
  NOR3_X1    g00383(.A1(new_n446_), .A2(new_n152_), .A3(new_n447_), .ZN(new_n448_));
  NOR2_X1    g00384(.A1(new_n133_), .A2(new_n123_), .ZN(new_n449_));
  NOR3_X1    g00385(.A1(new_n203_), .A2(new_n449_), .A3(new_n70_), .ZN(new_n450_));
  NAND2_X1   g00386(.A1(new_n111_), .A2(new_n318_), .ZN(new_n451_));
  NAND2_X1   g00387(.A1(new_n451_), .A2(new_n292_), .ZN(new_n452_));
  NOR2_X1    g00388(.A1(new_n176_), .A2(new_n123_), .ZN(new_n453_));
  NOR2_X1    g00389(.A1(new_n453_), .A2(new_n236_), .ZN(new_n454_));
  NAND4_X1   g00390(.A1(new_n448_), .A2(new_n450_), .A3(new_n452_), .A4(new_n454_), .ZN(new_n455_));
  NOR2_X1    g00391(.A1(new_n334_), .A2(new_n346_), .ZN(new_n456_));
  NOR2_X1    g00392(.A1(new_n135_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1     g00393(.I(new_n457_), .ZN(new_n458_));
  NOR2_X1    g00394(.A1(new_n129_), .A2(new_n66_), .ZN(new_n459_));
  NOR2_X1    g00395(.A1(new_n171_), .A2(new_n95_), .ZN(new_n460_));
  NOR4_X1    g00396(.A1(new_n458_), .A2(new_n183_), .A3(new_n459_), .A4(new_n460_), .ZN(new_n461_));
  INV_X1     g00397(.I(new_n461_), .ZN(new_n462_));
  NOR2_X1    g00398(.A1(new_n334_), .A2(new_n175_), .ZN(new_n463_));
  NAND2_X1   g00399(.A1(new_n440_), .A2(new_n273_), .ZN(new_n464_));
  INV_X1     g00400(.I(new_n464_), .ZN(new_n465_));
  NOR2_X1    g00401(.A1(new_n465_), .A2(new_n463_), .ZN(new_n466_));
  NAND2_X1   g00402(.A1(new_n196_), .A2(new_n245_), .ZN(new_n467_));
  NOR2_X1    g00403(.A1(new_n122_), .A2(new_n346_), .ZN(new_n468_));
  INV_X1     g00404(.I(new_n468_), .ZN(new_n469_));
  NOR2_X1    g00405(.A1(new_n72_), .A2(\a[25] ), .ZN(new_n470_));
  NAND3_X1   g00406(.A1(new_n206_), .A2(new_n470_), .A3(new_n100_), .ZN(new_n471_));
  NAND4_X1   g00407(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n472_));
  NOR2_X1    g00408(.A1(new_n86_), .A2(new_n219_), .ZN(new_n473_));
  NOR2_X1    g00409(.A1(new_n83_), .A2(new_n151_), .ZN(new_n474_));
  NOR2_X1    g00410(.A1(new_n73_), .A2(new_n91_), .ZN(new_n475_));
  NOR2_X1    g00411(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1   g00412(.A1(new_n253_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  NOR4_X1    g00413(.A1(new_n462_), .A2(new_n455_), .A3(new_n472_), .A4(new_n477_), .ZN(new_n478_));
  NAND2_X1   g00414(.A1(new_n79_), .A2(new_n156_), .ZN(new_n479_));
  INV_X1     g00415(.I(new_n119_), .ZN(new_n480_));
  INV_X1     g00416(.I(new_n225_), .ZN(new_n481_));
  NOR2_X1    g00417(.A1(new_n89_), .A2(new_n105_), .ZN(new_n482_));
  NOR2_X1    g00418(.A1(new_n482_), .A2(new_n297_), .ZN(new_n483_));
  NAND4_X1   g00419(.A1(new_n483_), .A2(new_n479_), .A3(new_n481_), .A4(new_n480_), .ZN(new_n484_));
  NOR2_X1    g00420(.A1(new_n88_), .A2(new_n129_), .ZN(new_n485_));
  NOR2_X1    g00421(.A1(new_n134_), .A2(new_n105_), .ZN(new_n486_));
  NOR2_X1    g00422(.A1(new_n75_), .A2(new_n151_), .ZN(new_n487_));
  NOR2_X1    g00423(.A1(new_n73_), .A2(new_n83_), .ZN(new_n488_));
  NOR4_X1    g00424(.A1(new_n485_), .A2(new_n486_), .A3(new_n488_), .A4(new_n487_), .ZN(new_n489_));
  NOR2_X1    g00425(.A1(new_n89_), .A2(new_n153_), .ZN(new_n490_));
  NOR2_X1    g00426(.A1(new_n133_), .A2(new_n131_), .ZN(new_n491_));
  NOR3_X1    g00427(.A1(new_n491_), .A2(new_n124_), .A3(new_n490_), .ZN(new_n492_));
  INV_X1     g00428(.I(new_n492_), .ZN(new_n493_));
  NOR3_X1    g00429(.A1(new_n484_), .A2(new_n493_), .A3(new_n489_), .ZN(new_n494_));
  INV_X1     g00430(.I(new_n141_), .ZN(new_n495_));
  NOR2_X1    g00431(.A1(new_n176_), .A2(new_n131_), .ZN(new_n496_));
  NOR4_X1    g00432(.A1(new_n495_), .A2(new_n106_), .A3(new_n289_), .A4(new_n496_), .ZN(new_n497_));
  NOR2_X1    g00433(.A1(new_n69_), .A2(new_n133_), .ZN(new_n498_));
  AOI21_X1   g00434(.A1(new_n69_), .A2(new_n123_), .B(new_n151_), .ZN(new_n499_));
  NOR2_X1    g00435(.A1(new_n499_), .A2(new_n498_), .ZN(new_n500_));
  NAND2_X1   g00436(.A1(new_n142_), .A2(new_n273_), .ZN(new_n501_));
  NAND2_X1   g00437(.A1(new_n156_), .A2(new_n273_), .ZN(new_n502_));
  NAND2_X1   g00438(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR4_X1    g00439(.A1(new_n497_), .A2(new_n102_), .A3(new_n500_), .A4(new_n503_), .ZN(new_n504_));
  NOR2_X1    g00440(.A1(new_n101_), .A2(new_n134_), .ZN(new_n505_));
  NOR2_X1    g00441(.A1(new_n346_), .A2(new_n66_), .ZN(new_n506_));
  NOR2_X1    g00442(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1   g00443(.A1(new_n111_), .A2(new_n273_), .ZN(new_n508_));
  NAND2_X1   g00444(.A1(new_n159_), .A2(new_n230_), .ZN(new_n509_));
  NOR2_X1    g00445(.A1(new_n75_), .A2(new_n122_), .ZN(new_n510_));
  INV_X1     g00446(.I(new_n510_), .ZN(new_n511_));
  NAND2_X1   g00447(.A1(new_n265_), .A2(new_n185_), .ZN(new_n512_));
  NAND4_X1   g00448(.A1(new_n511_), .A2(new_n508_), .A3(new_n509_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1   g00449(.A1(new_n513_), .A2(new_n507_), .ZN(new_n514_));
  NOR2_X1    g00450(.A1(new_n175_), .A2(new_n85_), .ZN(new_n515_));
  NOR2_X1    g00451(.A1(new_n515_), .A2(new_n239_), .ZN(new_n516_));
  NOR2_X1    g00452(.A1(new_n91_), .A2(new_n151_), .ZN(new_n517_));
  NOR2_X1    g00453(.A1(new_n151_), .A2(new_n346_), .ZN(new_n518_));
  NOR2_X1    g00454(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1   g00455(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1   g00456(.A1(new_n284_), .A2(new_n156_), .ZN(new_n521_));
  NAND2_X1   g00457(.A1(new_n139_), .A2(new_n109_), .ZN(new_n522_));
  NAND2_X1   g00458(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1    g00459(.A1(new_n255_), .A2(new_n164_), .ZN(new_n524_));
  INV_X1     g00460(.I(new_n524_), .ZN(new_n525_));
  NOR4_X1    g00461(.A1(new_n514_), .A2(new_n520_), .A3(new_n523_), .A4(new_n525_), .ZN(new_n526_));
  AND3_X2    g00462(.A1(new_n526_), .A2(new_n494_), .A3(new_n504_), .Z(new_n527_));
  NAND2_X1   g00463(.A1(new_n527_), .A2(new_n478_), .ZN(new_n528_));
  NOR2_X1    g00464(.A1(new_n528_), .A2(new_n445_), .ZN(new_n529_));
  NOR2_X1    g00465(.A1(new_n147_), .A2(new_n485_), .ZN(new_n530_));
  NOR2_X1    g00466(.A1(new_n73_), .A2(new_n131_), .ZN(new_n531_));
  NOR4_X1    g00467(.A1(new_n530_), .A2(new_n262_), .A3(new_n459_), .A4(new_n531_), .ZN(new_n532_));
  NAND2_X1   g00468(.A1(new_n464_), .A2(new_n502_), .ZN(new_n533_));
  NOR2_X1    g00469(.A1(new_n101_), .A2(new_n89_), .ZN(new_n534_));
  NOR2_X1    g00470(.A1(new_n75_), .A2(new_n148_), .ZN(new_n535_));
  NOR2_X1    g00471(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1   g00472(.A1(new_n159_), .A2(new_n440_), .B(new_n143_), .ZN(new_n537_));
  NAND2_X1   g00473(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1    g00474(.A1(new_n406_), .A2(new_n312_), .ZN(new_n539_));
  NAND2_X1   g00475(.A1(new_n404_), .A2(new_n139_), .ZN(new_n540_));
  INV_X1     g00476(.I(new_n540_), .ZN(new_n541_));
  NOR2_X1    g00477(.A1(new_n541_), .A2(new_n135_), .ZN(new_n542_));
  NOR2_X1    g00478(.A1(new_n172_), .A2(new_n235_), .ZN(new_n543_));
  OAI22_X1   g00479(.A1(new_n118_), .A2(new_n175_), .B1(new_n89_), .B2(new_n88_), .ZN(new_n544_));
  INV_X1     g00480(.I(new_n544_), .ZN(new_n545_));
  NAND4_X1   g00481(.A1(new_n542_), .A2(new_n539_), .A3(new_n543_), .A4(new_n545_), .ZN(new_n546_));
  NOR3_X1    g00482(.A1(new_n546_), .A2(new_n533_), .A3(new_n538_), .ZN(new_n547_));
  NOR2_X1    g00483(.A1(new_n176_), .A2(new_n69_), .ZN(new_n548_));
  NOR2_X1    g00484(.A1(new_n105_), .A2(new_n116_), .ZN(new_n549_));
  NOR4_X1    g00485(.A1(new_n548_), .A2(new_n549_), .A3(new_n261_), .A4(new_n506_), .ZN(new_n550_));
  NAND2_X1   g00486(.A1(new_n355_), .A2(new_n112_), .ZN(new_n551_));
  NAND2_X1   g00487(.A1(new_n551_), .A2(new_n325_), .ZN(new_n552_));
  NOR2_X1    g00488(.A1(new_n75_), .A2(new_n133_), .ZN(new_n553_));
  NOR2_X1    g00489(.A1(new_n76_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1     g00490(.I(new_n554_), .ZN(new_n555_));
  NOR2_X1    g00491(.A1(new_n116_), .A2(new_n122_), .ZN(new_n556_));
  NOR2_X1    g00492(.A1(new_n556_), .A2(new_n347_), .ZN(new_n557_));
  INV_X1     g00493(.I(new_n557_), .ZN(new_n558_));
  NOR4_X1    g00494(.A1(new_n555_), .A2(new_n558_), .A3(new_n550_), .A4(new_n552_), .ZN(new_n559_));
  NOR2_X1    g00495(.A1(new_n85_), .A2(new_n150_), .ZN(new_n560_));
  NOR2_X1    g00496(.A1(new_n131_), .A2(new_n153_), .ZN(new_n561_));
  NOR4_X1    g00497(.A1(new_n190_), .A2(new_n475_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  INV_X1     g00498(.I(new_n389_), .ZN(new_n563_));
  NAND2_X1   g00499(.A1(new_n245_), .A2(new_n206_), .ZN(new_n564_));
  NAND2_X1   g00500(.A1(new_n378_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1    g00501(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1     g00502(.I(new_n566_), .ZN(new_n567_));
  NAND2_X1   g00503(.A1(new_n205_), .A2(new_n440_), .ZN(new_n568_));
  NAND2_X1   g00504(.A1(new_n568_), .A2(new_n409_), .ZN(new_n569_));
  NOR2_X1    g00505(.A1(new_n569_), .A2(new_n324_), .ZN(new_n570_));
  INV_X1     g00506(.I(new_n570_), .ZN(new_n571_));
  NAND2_X1   g00507(.A1(new_n159_), .A2(new_n284_), .ZN(new_n572_));
  INV_X1     g00508(.I(new_n572_), .ZN(new_n573_));
  NOR2_X1    g00509(.A1(new_n69_), .A2(new_n148_), .ZN(new_n574_));
  NOR2_X1    g00510(.A1(new_n214_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1     g00511(.I(new_n575_), .ZN(new_n576_));
  NOR2_X1    g00512(.A1(new_n175_), .A2(new_n153_), .ZN(new_n577_));
  NOR3_X1    g00513(.A1(new_n576_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1     g00514(.I(new_n578_), .ZN(new_n579_));
  NOR4_X1    g00515(.A1(new_n579_), .A2(new_n567_), .A3(new_n562_), .A4(new_n571_), .ZN(new_n580_));
  NAND4_X1   g00516(.A1(new_n580_), .A2(new_n532_), .A3(new_n547_), .A4(new_n559_), .ZN(new_n581_));
  NOR2_X1    g00517(.A1(new_n176_), .A2(new_n346_), .ZN(new_n582_));
  NOR3_X1    g00518(.A1(new_n343_), .A2(new_n582_), .A3(new_n517_), .ZN(new_n583_));
  NOR2_X1    g00519(.A1(new_n75_), .A2(new_n115_), .ZN(new_n584_));
  NOR4_X1    g00520(.A1(new_n294_), .A2(new_n498_), .A3(new_n584_), .A4(new_n282_), .ZN(new_n585_));
  INV_X1     g00521(.I(new_n585_), .ZN(new_n586_));
  NOR2_X1    g00522(.A1(new_n88_), .A2(new_n91_), .ZN(new_n587_));
  NOR2_X1    g00523(.A1(new_n304_), .A2(new_n587_), .ZN(new_n588_));
  AND3_X2    g00524(.A1(new_n586_), .A2(new_n583_), .A3(new_n588_), .Z(new_n589_));
  NOR2_X1    g00525(.A1(new_n148_), .A2(new_n169_), .ZN(new_n590_));
  NOR2_X1    g00526(.A1(new_n171_), .A2(new_n176_), .ZN(new_n591_));
  NAND2_X1   g00527(.A1(new_n139_), .A2(new_n185_), .ZN(new_n592_));
  INV_X1     g00528(.I(new_n592_), .ZN(new_n593_));
  NOR2_X1    g00529(.A1(new_n153_), .A2(new_n346_), .ZN(new_n594_));
  NOR4_X1    g00530(.A1(new_n593_), .A2(new_n590_), .A3(new_n591_), .A4(new_n594_), .ZN(new_n595_));
  NOR2_X1    g00531(.A1(new_n97_), .A2(new_n73_), .ZN(new_n596_));
  NOR2_X1    g00532(.A1(new_n596_), .A2(new_n419_), .ZN(new_n597_));
  NAND2_X1   g00533(.A1(new_n77_), .A2(new_n143_), .ZN(new_n598_));
  NAND2_X1   g00534(.A1(new_n404_), .A2(new_n318_), .ZN(new_n599_));
  NAND2_X1   g00535(.A1(new_n599_), .A2(new_n598_), .ZN(new_n600_));
  INV_X1     g00536(.I(new_n600_), .ZN(new_n601_));
  INV_X1     g00537(.I(new_n362_), .ZN(new_n602_));
  NOR2_X1    g00538(.A1(new_n83_), .A2(new_n115_), .ZN(new_n603_));
  NOR2_X1    g00539(.A1(new_n69_), .A2(new_n115_), .ZN(new_n604_));
  NOR4_X1    g00540(.A1(new_n98_), .A2(new_n117_), .A3(new_n604_), .A4(new_n183_), .ZN(new_n605_));
  NAND2_X1   g00541(.A1(new_n265_), .A2(new_n140_), .ZN(new_n606_));
  INV_X1     g00542(.I(new_n606_), .ZN(new_n607_));
  NOR4_X1    g00543(.A1(new_n605_), .A2(new_n602_), .A3(new_n603_), .A4(new_n607_), .ZN(new_n608_));
  NAND4_X1   g00544(.A1(new_n608_), .A2(new_n595_), .A3(new_n597_), .A4(new_n601_), .ZN(new_n609_));
  NOR2_X1    g00545(.A1(new_n129_), .A2(new_n122_), .ZN(new_n610_));
  NOR2_X1    g00546(.A1(new_n334_), .A2(new_n131_), .ZN(new_n611_));
  INV_X1     g00547(.I(new_n164_), .ZN(new_n612_));
  NAND2_X1   g00548(.A1(new_n612_), .A2(new_n394_), .ZN(new_n613_));
  NOR4_X1    g00549(.A1(new_n613_), .A2(new_n381_), .A3(new_n610_), .A4(new_n611_), .ZN(new_n614_));
  NOR2_X1    g00550(.A1(new_n176_), .A2(new_n75_), .ZN(new_n615_));
  NOR2_X1    g00551(.A1(new_n102_), .A2(new_n149_), .ZN(new_n616_));
  INV_X1     g00552(.I(new_n616_), .ZN(new_n617_));
  AOI22_X1   g00553(.A1(new_n318_), .A2(new_n77_), .B1(new_n181_), .B2(new_n350_), .ZN(new_n618_));
  NOR3_X1    g00554(.A1(new_n617_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1   g00555(.A1(new_n619_), .A2(new_n614_), .ZN(new_n620_));
  NOR2_X1    g00556(.A1(new_n609_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1   g00557(.A1(new_n621_), .A2(new_n589_), .ZN(new_n622_));
  INV_X1     g00558(.I(new_n622_), .ZN(new_n623_));
  OAI22_X1   g00559(.A1(new_n134_), .A2(new_n85_), .B1(new_n95_), .B2(new_n123_), .ZN(new_n624_));
  NOR2_X1    g00560(.A1(new_n69_), .A2(new_n153_), .ZN(new_n625_));
  NOR2_X1    g00561(.A1(new_n625_), .A2(new_n329_), .ZN(new_n626_));
  NAND2_X1   g00562(.A1(new_n180_), .A2(new_n270_), .ZN(new_n627_));
  INV_X1     g00563(.I(new_n154_), .ZN(new_n628_));
  NAND2_X1   g00564(.A1(new_n628_), .A2(new_n627_), .ZN(new_n629_));
  AOI21_X1   g00565(.A1(new_n118_), .A2(new_n334_), .B(new_n75_), .ZN(new_n630_));
  INV_X1     g00566(.I(new_n630_), .ZN(new_n631_));
  NAND4_X1   g00567(.A1(new_n629_), .A2(new_n624_), .A3(new_n631_), .A4(new_n626_), .ZN(new_n632_));
  NOR2_X1    g00568(.A1(new_n134_), .A2(new_n334_), .ZN(new_n633_));
  NOR2_X1    g00569(.A1(new_n134_), .A2(new_n95_), .ZN(new_n634_));
  NOR3_X1    g00570(.A1(new_n633_), .A2(new_n634_), .A3(new_n518_), .ZN(new_n635_));
  INV_X1     g00571(.I(new_n635_), .ZN(new_n636_));
  NOR2_X1    g00572(.A1(new_n83_), .A2(new_n105_), .ZN(new_n637_));
  NOR2_X1    g00573(.A1(new_n334_), .A2(new_n83_), .ZN(new_n638_));
  NOR4_X1    g00574(.A1(new_n637_), .A2(new_n638_), .A3(new_n352_), .A4(new_n430_), .ZN(new_n639_));
  NOR2_X1    g00575(.A1(new_n115_), .A2(new_n169_), .ZN(new_n640_));
  NOR2_X1    g00576(.A1(new_n640_), .A2(new_n359_), .ZN(new_n641_));
  INV_X1     g00577(.I(new_n641_), .ZN(new_n642_));
  NAND2_X1   g00578(.A1(new_n108_), .A2(new_n206_), .ZN(new_n643_));
  INV_X1     g00579(.I(new_n643_), .ZN(new_n644_));
  NOR4_X1    g00580(.A1(new_n642_), .A2(new_n335_), .A3(new_n456_), .A4(new_n644_), .ZN(new_n645_));
  NOR2_X1    g00581(.A1(new_n152_), .A2(new_n310_), .ZN(new_n646_));
  INV_X1     g00582(.I(new_n646_), .ZN(new_n647_));
  NOR2_X1    g00583(.A1(new_n175_), .A2(new_n133_), .ZN(new_n648_));
  NOR2_X1    g00584(.A1(new_n648_), .A2(new_n376_), .ZN(new_n649_));
  INV_X1     g00585(.I(new_n649_), .ZN(new_n650_));
  NOR2_X1    g00586(.A1(new_n650_), .A2(new_n647_), .ZN(new_n651_));
  NOR2_X1    g00587(.A1(new_n85_), .A2(new_n89_), .ZN(new_n652_));
  NOR2_X1    g00588(.A1(new_n81_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1    g00589(.A1(new_n134_), .A2(new_n151_), .ZN(new_n654_));
  NAND2_X1   g00590(.A1(new_n355_), .A2(new_n230_), .ZN(new_n655_));
  INV_X1     g00591(.I(new_n655_), .ZN(new_n656_));
  NOR2_X1    g00592(.A1(new_n656_), .A2(new_n654_), .ZN(new_n657_));
  NAND4_X1   g00593(.A1(new_n645_), .A2(new_n651_), .A3(new_n653_), .A4(new_n657_), .ZN(new_n658_));
  NOR4_X1    g00594(.A1(new_n658_), .A2(new_n632_), .A3(new_n636_), .A4(new_n639_), .ZN(new_n659_));
  NOR2_X1    g00595(.A1(new_n73_), .A2(new_n123_), .ZN(new_n660_));
  NOR3_X1    g00596(.A1(new_n213_), .A2(new_n447_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1   g00597(.A1(new_n196_), .A2(new_n139_), .ZN(new_n662_));
  NAND2_X1   g00598(.A1(new_n662_), .A2(new_n423_), .ZN(new_n663_));
  INV_X1     g00599(.I(new_n663_), .ZN(new_n664_));
  NAND2_X1   g00600(.A1(new_n355_), .A2(new_n245_), .ZN(new_n665_));
  NOR2_X1    g00601(.A1(new_n101_), .A2(new_n123_), .ZN(new_n666_));
  INV_X1     g00602(.I(new_n666_), .ZN(new_n667_));
  NAND4_X1   g00603(.A1(new_n664_), .A2(new_n661_), .A3(new_n665_), .A4(new_n667_), .ZN(new_n668_));
  NAND2_X1   g00604(.A1(new_n156_), .A2(new_n143_), .ZN(new_n669_));
  NOR2_X1    g00605(.A1(new_n95_), .A2(new_n116_), .ZN(new_n670_));
  NOR2_X1    g00606(.A1(new_n251_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1   g00607(.A1(new_n79_), .A2(new_n206_), .ZN(new_n672_));
  NAND3_X1   g00608(.A1(new_n671_), .A2(new_n669_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1     g00609(.I(new_n673_), .ZN(new_n674_));
  INV_X1     g00610(.I(new_n92_), .ZN(new_n675_));
  NAND2_X1   g00611(.A1(new_n355_), .A2(new_n265_), .ZN(new_n676_));
  NAND2_X1   g00612(.A1(new_n275_), .A2(new_n186_), .ZN(new_n677_));
  NAND3_X1   g00613(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  NOR3_X1    g00614(.A1(new_n674_), .A2(new_n668_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1   g00615(.A1(new_n158_), .A2(new_n196_), .ZN(new_n680_));
  NOR2_X1    g00616(.A1(new_n89_), .A2(new_n115_), .ZN(new_n681_));
  NOR2_X1    g00617(.A1(new_n83_), .A2(new_n122_), .ZN(new_n682_));
  NOR2_X1    g00618(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1    g00619(.A1(new_n175_), .A2(new_n66_), .ZN(new_n684_));
  INV_X1     g00620(.I(new_n684_), .ZN(new_n685_));
  NAND2_X1   g00621(.A1(new_n205_), .A2(new_n77_), .ZN(new_n686_));
  NAND2_X1   g00622(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1     g00623(.I(new_n687_), .ZN(new_n688_));
  NOR2_X1    g00624(.A1(new_n85_), .A2(new_n169_), .ZN(new_n689_));
  INV_X1     g00625(.I(new_n689_), .ZN(new_n690_));
  NAND4_X1   g00626(.A1(new_n688_), .A2(new_n683_), .A3(new_n680_), .A4(new_n690_), .ZN(new_n691_));
  NOR4_X1    g00627(.A1(new_n691_), .A2(new_n345_), .A3(new_n396_), .A4(new_n460_), .ZN(new_n692_));
  NAND4_X1   g00628(.A1(new_n623_), .A2(new_n659_), .A3(new_n679_), .A4(new_n692_), .ZN(new_n693_));
  NOR2_X1    g00629(.A1(new_n693_), .A2(new_n581_), .ZN(new_n694_));
  NOR2_X1    g00630(.A1(new_n97_), .A2(new_n148_), .ZN(new_n695_));
  NOR4_X1    g00631(.A1(new_n465_), .A2(new_n307_), .A3(new_n437_), .A4(new_n695_), .ZN(new_n696_));
  AOI21_X1   g00632(.A1(new_n85_), .A2(new_n95_), .B(new_n83_), .ZN(new_n697_));
  NOR2_X1    g00633(.A1(new_n69_), .A2(new_n105_), .ZN(new_n698_));
  NOR3_X1    g00634(.A1(new_n697_), .A2(new_n420_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1     g00635(.I(new_n699_), .ZN(new_n700_));
  NAND2_X1   g00636(.A1(new_n111_), .A2(new_n205_), .ZN(new_n701_));
  NAND3_X1   g00637(.A1(new_n701_), .A2(new_n246_), .A3(new_n394_), .ZN(new_n702_));
  NOR2_X1    g00638(.A1(new_n175_), .A2(new_n148_), .ZN(new_n703_));
  NOR4_X1    g00639(.A1(new_n214_), .A2(new_n241_), .A3(new_n648_), .A4(new_n703_), .ZN(new_n704_));
  NOR4_X1    g00640(.A1(new_n700_), .A2(new_n696_), .A3(new_n702_), .A4(new_n704_), .ZN(new_n705_));
  NOR2_X1    g00641(.A1(new_n251_), .A2(new_n256_), .ZN(new_n706_));
  NAND2_X1   g00642(.A1(new_n196_), .A2(new_n112_), .ZN(new_n707_));
  NAND2_X1   g00643(.A1(new_n707_), .A2(new_n665_), .ZN(new_n708_));
  NAND2_X1   g00644(.A1(new_n318_), .A2(new_n350_), .ZN(new_n709_));
  NAND4_X1   g00645(.A1(new_n706_), .A2(new_n708_), .A3(new_n353_), .A4(new_n709_), .ZN(new_n710_));
  INV_X1     g00646(.I(new_n710_), .ZN(new_n711_));
  NOR2_X1    g00647(.A1(new_n183_), .A2(new_n428_), .ZN(new_n712_));
  NAND2_X1   g00648(.A1(new_n540_), .A2(new_n271_), .ZN(new_n713_));
  NOR2_X1    g00649(.A1(new_n118_), .A2(new_n134_), .ZN(new_n714_));
  NOR2_X1    g00650(.A1(new_n73_), .A2(new_n150_), .ZN(new_n715_));
  NOR2_X1    g00651(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1     g00652(.I(new_n716_), .ZN(new_n717_));
  NOR2_X1    g00653(.A1(new_n131_), .A2(new_n88_), .ZN(new_n718_));
  NOR2_X1    g00654(.A1(new_n334_), .A2(new_n91_), .ZN(new_n719_));
  NOR2_X1    g00655(.A1(new_n719_), .A2(new_n718_), .ZN(new_n720_));
  NOR2_X1    g00656(.A1(new_n97_), .A2(new_n122_), .ZN(new_n721_));
  NOR2_X1    g00657(.A1(new_n117_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1    g00658(.A1(new_n634_), .A2(new_n297_), .ZN(new_n723_));
  NOR2_X1    g00659(.A1(new_n153_), .A2(new_n150_), .ZN(new_n724_));
  NOR2_X1    g00660(.A1(new_n90_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1   g00661(.A1(new_n722_), .A2(new_n723_), .A3(new_n720_), .A4(new_n725_), .ZN(new_n726_));
  NOR4_X1    g00662(.A1(new_n726_), .A2(new_n712_), .A3(new_n713_), .A4(new_n717_), .ZN(new_n727_));
  NAND3_X1   g00663(.A1(new_n727_), .A2(new_n711_), .A3(new_n705_), .ZN(new_n728_));
  OAI22_X1   g00664(.A1(new_n176_), .A2(new_n75_), .B1(new_n151_), .B2(new_n346_), .ZN(new_n729_));
  INV_X1     g00665(.I(new_n729_), .ZN(new_n730_));
  NOR2_X1    g00666(.A1(new_n169_), .A2(new_n153_), .ZN(new_n731_));
  NOR2_X1    g00667(.A1(new_n97_), .A2(new_n153_), .ZN(new_n732_));
  NOR4_X1    g00668(.A1(new_n147_), .A2(new_n731_), .A3(new_n682_), .A4(new_n732_), .ZN(new_n733_));
  NOR2_X1    g00669(.A1(new_n171_), .A2(new_n115_), .ZN(new_n734_));
  NOR4_X1    g00670(.A1(new_n602_), .A2(new_n288_), .A3(new_n549_), .A4(new_n734_), .ZN(new_n735_));
  NOR2_X1    g00671(.A1(new_n123_), .A2(new_n66_), .ZN(new_n736_));
  NOR4_X1    g00672(.A1(new_n345_), .A2(new_n242_), .A3(new_n560_), .A4(new_n736_), .ZN(new_n737_));
  NOR4_X1    g00673(.A1(new_n735_), .A2(new_n733_), .A3(new_n730_), .A4(new_n737_), .ZN(new_n738_));
  NAND2_X1   g00674(.A1(new_n77_), .A2(new_n108_), .ZN(new_n739_));
  INV_X1     g00675(.I(new_n739_), .ZN(new_n740_));
  NOR2_X1    g00676(.A1(new_n83_), .A2(new_n148_), .ZN(new_n741_));
  NOR4_X1    g00677(.A1(new_n740_), .A2(new_n191_), .A3(new_n403_), .A4(new_n741_), .ZN(new_n742_));
  NOR4_X1    g00678(.A1(new_n76_), .A2(new_n304_), .A3(new_n652_), .A4(new_n152_), .ZN(new_n743_));
  NOR2_X1    g00679(.A1(new_n133_), .A2(new_n150_), .ZN(new_n744_));
  NOR3_X1    g00680(.A1(new_n670_), .A2(new_n136_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1     g00681(.I(new_n745_), .ZN(new_n746_));
  NOR2_X1    g00682(.A1(new_n460_), .A2(new_n574_), .ZN(new_n747_));
  INV_X1     g00683(.I(new_n747_), .ZN(new_n748_));
  NOR2_X1    g00684(.A1(new_n148_), .A2(new_n346_), .ZN(new_n749_));
  NOR4_X1    g00685(.A1(new_n748_), .A2(new_n495_), .A3(new_n633_), .A4(new_n749_), .ZN(new_n750_));
  NOR2_X1    g00686(.A1(new_n118_), .A2(new_n116_), .ZN(new_n751_));
  NOR2_X1    g00687(.A1(new_n171_), .A2(new_n133_), .ZN(new_n752_));
  NOR2_X1    g00688(.A1(new_n118_), .A2(new_n89_), .ZN(new_n753_));
  NOR4_X1    g00689(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .A4(new_n330_), .ZN(new_n754_));
  AOI22_X1   g00690(.A1(new_n404_), .A2(new_n318_), .B1(new_n109_), .B2(new_n186_), .ZN(new_n755_));
  AOI21_X1   g00691(.A1(new_n69_), .A2(new_n97_), .B(new_n95_), .ZN(new_n756_));
  INV_X1     g00692(.I(new_n756_), .ZN(new_n757_));
  NAND4_X1   g00693(.A1(new_n750_), .A2(new_n754_), .A3(new_n755_), .A4(new_n757_), .ZN(new_n758_));
  NOR4_X1    g00694(.A1(new_n758_), .A2(new_n742_), .A3(new_n743_), .A4(new_n746_), .ZN(new_n759_));
  NAND2_X1   g00695(.A1(new_n759_), .A2(new_n738_), .ZN(new_n760_));
  NAND2_X1   g00696(.A1(new_n284_), .A2(new_n77_), .ZN(new_n761_));
  NOR2_X1    g00697(.A1(new_n415_), .A2(new_n282_), .ZN(new_n762_));
  NOR2_X1    g00698(.A1(new_n101_), .A2(new_n346_), .ZN(new_n763_));
  NOR2_X1    g00699(.A1(new_n88_), .A2(new_n346_), .ZN(new_n764_));
  NOR2_X1    g00700(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1    g00701(.A1(new_n607_), .A2(new_n449_), .ZN(new_n766_));
  NAND4_X1   g00702(.A1(new_n766_), .A2(new_n762_), .A3(new_n761_), .A4(new_n765_), .ZN(new_n767_));
  NOR2_X1    g00703(.A1(new_n106_), .A2(new_n216_), .ZN(new_n768_));
  INV_X1     g00704(.I(new_n768_), .ZN(new_n769_));
  NOR2_X1    g00705(.A1(new_n101_), .A2(new_n69_), .ZN(new_n770_));
  NOR4_X1    g00706(.A1(new_n769_), .A2(new_n161_), .A3(new_n596_), .A4(new_n770_), .ZN(new_n771_));
  NOR2_X1    g00707(.A1(new_n105_), .A2(new_n169_), .ZN(new_n772_));
  NAND2_X1   g00708(.A1(new_n79_), .A2(new_n159_), .ZN(new_n773_));
  INV_X1     g00709(.I(new_n773_), .ZN(new_n774_));
  NOR2_X1    g00710(.A1(new_n774_), .A2(new_n772_), .ZN(new_n775_));
  NOR2_X1    g00711(.A1(new_n123_), .A2(new_n151_), .ZN(new_n776_));
  NOR2_X1    g00712(.A1(new_n587_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1     g00713(.I(new_n100_), .ZN(new_n778_));
  NOR4_X1    g00714(.A1(new_n129_), .A2(new_n778_), .A3(new_n78_), .A4(\a[26] ), .ZN(new_n779_));
  NOR2_X1    g00715(.A1(new_n779_), .A2(new_n475_), .ZN(new_n780_));
  INV_X1     g00716(.I(new_n780_), .ZN(new_n781_));
  NOR2_X1    g00717(.A1(new_n133_), .A2(new_n129_), .ZN(new_n782_));
  NOR2_X1    g00718(.A1(new_n89_), .A2(new_n133_), .ZN(new_n783_));
  NOR2_X1    g00719(.A1(new_n783_), .A2(new_n782_), .ZN(new_n784_));
  INV_X1     g00720(.I(new_n784_), .ZN(new_n785_));
  NOR2_X1    g00721(.A1(new_n781_), .A2(new_n785_), .ZN(new_n786_));
  NAND4_X1   g00722(.A1(new_n771_), .A2(new_n786_), .A3(new_n775_), .A4(new_n777_), .ZN(new_n787_));
  INV_X1     g00723(.I(new_n110_), .ZN(new_n788_));
  NOR4_X1    g00724(.A1(new_n788_), .A2(new_n235_), .A3(new_n638_), .A4(new_n190_), .ZN(new_n789_));
  INV_X1     g00725(.I(new_n213_), .ZN(new_n790_));
  NOR2_X1    g00726(.A1(new_n118_), .A2(new_n346_), .ZN(new_n791_));
  NOR2_X1    g00727(.A1(new_n791_), .A2(new_n594_), .ZN(new_n792_));
  NAND3_X1   g00728(.A1(new_n792_), .A2(new_n480_), .A3(new_n790_), .ZN(new_n793_));
  INV_X1     g00729(.I(new_n793_), .ZN(new_n794_));
  NAND2_X1   g00730(.A1(new_n158_), .A2(new_n206_), .ZN(new_n795_));
  NOR2_X1    g00731(.A1(new_n118_), .A2(new_n91_), .ZN(new_n796_));
  INV_X1     g00732(.I(new_n796_), .ZN(new_n797_));
  NAND4_X1   g00733(.A1(new_n797_), .A2(new_n795_), .A3(new_n598_), .A4(new_n342_), .ZN(new_n798_));
  INV_X1     g00734(.I(new_n798_), .ZN(new_n799_));
  NOR3_X1    g00735(.A1(new_n794_), .A2(new_n799_), .A3(new_n789_), .ZN(new_n800_));
  NOR2_X1    g00736(.A1(new_n115_), .A2(new_n150_), .ZN(new_n801_));
  NOR4_X1    g00737(.A1(new_n387_), .A2(new_n491_), .A3(new_n130_), .A4(new_n561_), .ZN(new_n802_));
  NOR4_X1    g00738(.A1(new_n802_), .A2(new_n310_), .A3(new_n801_), .A4(new_n498_), .ZN(new_n803_));
  NOR2_X1    g00739(.A1(new_n131_), .A2(new_n148_), .ZN(new_n804_));
  NOR2_X1    g00740(.A1(new_n804_), .A2(new_n610_), .ZN(new_n805_));
  NOR3_X1    g00741(.A1(new_n805_), .A2(new_n335_), .A3(new_n359_), .ZN(new_n806_));
  NAND2_X1   g00742(.A1(new_n158_), .A2(new_n185_), .ZN(new_n807_));
  NAND2_X1   g00743(.A1(new_n79_), .A2(new_n196_), .ZN(new_n808_));
  NAND2_X1   g00744(.A1(new_n206_), .A2(new_n273_), .ZN(new_n809_));
  NAND4_X1   g00745(.A1(new_n385_), .A2(new_n807_), .A3(new_n808_), .A4(new_n809_), .ZN(new_n810_));
  NAND4_X1   g00746(.A1(new_n800_), .A2(new_n803_), .A3(new_n806_), .A4(new_n810_), .ZN(new_n811_));
  OR4_X2     g00747(.A1(new_n760_), .A2(new_n767_), .A3(new_n787_), .A4(new_n811_), .Z(new_n812_));
  NOR2_X1    g00748(.A1(new_n812_), .A2(new_n728_), .ZN(new_n813_));
  INV_X1     g00749(.I(new_n813_), .ZN(new_n814_));
  INV_X1     g00750(.I(new_n527_), .ZN(new_n815_));
  NOR2_X1    g00751(.A1(new_n212_), .A2(new_n460_), .ZN(new_n816_));
  NOR2_X1    g00752(.A1(new_n334_), .A2(new_n116_), .ZN(new_n817_));
  NOR2_X1    g00753(.A1(new_n817_), .A2(new_n561_), .ZN(new_n818_));
  OAI21_X1   g00754(.A1(new_n158_), .A2(new_n230_), .B(new_n77_), .ZN(new_n819_));
  NOR2_X1    g00755(.A1(new_n98_), .A2(new_n324_), .ZN(new_n820_));
  NAND4_X1   g00756(.A1(new_n816_), .A2(new_n820_), .A3(new_n818_), .A4(new_n819_), .ZN(new_n821_));
  NAND2_X1   g00757(.A1(new_n378_), .A2(new_n395_), .ZN(new_n822_));
  NAND2_X1   g00758(.A1(new_n230_), .A2(new_n440_), .ZN(new_n823_));
  NAND2_X1   g00759(.A1(new_n245_), .A2(new_n440_), .ZN(new_n824_));
  NAND2_X1   g00760(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NOR4_X1    g00761(.A1(new_n822_), .A2(new_n825_), .A3(new_n312_), .A4(new_n335_), .ZN(new_n826_));
  NOR2_X1    g00762(.A1(new_n396_), .A2(new_n749_), .ZN(new_n827_));
  NOR2_X1    g00763(.A1(new_n788_), .A2(new_n227_), .ZN(new_n828_));
  NOR2_X1    g00764(.A1(new_n370_), .A2(new_n594_), .ZN(new_n829_));
  NAND4_X1   g00765(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .A4(new_n829_), .ZN(new_n830_));
  NOR2_X1    g00766(.A1(new_n830_), .A2(new_n821_), .ZN(new_n831_));
  NAND2_X1   g00767(.A1(new_n142_), .A2(new_n181_), .ZN(new_n832_));
  NAND4_X1   g00768(.A1(new_n199_), .A2(new_n739_), .A3(new_n311_), .A4(new_n832_), .ZN(new_n833_));
  NAND2_X1   g00769(.A1(new_n284_), .A2(new_n142_), .ZN(new_n834_));
  NAND2_X1   g00770(.A1(new_n834_), .A2(new_n276_), .ZN(new_n835_));
  INV_X1     g00771(.I(new_n835_), .ZN(new_n836_));
  NOR2_X1    g00772(.A1(new_n83_), .A2(new_n95_), .ZN(new_n837_));
  NOR4_X1    g00773(.A1(new_n602_), .A2(new_n666_), .A3(new_n359_), .A4(new_n837_), .ZN(new_n838_));
  INV_X1     g00774(.I(new_n838_), .ZN(new_n839_));
  NAND2_X1   g00775(.A1(new_n275_), .A2(new_n270_), .ZN(new_n840_));
  NOR2_X1    g00776(.A1(new_n73_), .A2(new_n129_), .ZN(new_n841_));
  INV_X1     g00777(.I(new_n841_), .ZN(new_n842_));
  NAND2_X1   g00778(.A1(new_n270_), .A2(new_n350_), .ZN(new_n843_));
  NAND2_X1   g00779(.A1(new_n467_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1     g00780(.I(new_n844_), .ZN(new_n845_));
  NAND3_X1   g00781(.A1(new_n845_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n846_));
  NAND4_X1   g00782(.A1(new_n846_), .A2(new_n839_), .A3(new_n833_), .A4(new_n836_), .ZN(new_n847_));
  OAI22_X1   g00783(.A1(new_n171_), .A2(new_n176_), .B1(new_n148_), .B2(new_n150_), .ZN(new_n848_));
  NAND2_X1   g00784(.A1(new_n185_), .A2(new_n270_), .ZN(new_n849_));
  NAND2_X1   g00785(.A1(new_n572_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1     g00786(.I(new_n850_), .ZN(new_n851_));
  NOR2_X1    g00787(.A1(new_n446_), .A2(new_n531_), .ZN(new_n852_));
  NAND4_X1   g00788(.A1(new_n851_), .A2(new_n852_), .A3(new_n389_), .A4(new_n848_), .ZN(new_n853_));
  NAND2_X1   g00789(.A1(new_n205_), .A2(new_n180_), .ZN(new_n854_));
  NAND3_X1   g00790(.A1(new_n287_), .A2(new_n854_), .A3(new_n676_), .ZN(new_n855_));
  NAND2_X1   g00791(.A1(new_n159_), .A2(new_n143_), .ZN(new_n856_));
  NAND3_X1   g00792(.A1(new_n80_), .A2(new_n856_), .A3(new_n301_), .ZN(new_n857_));
  NOR4_X1    g00793(.A1(new_n847_), .A2(new_n853_), .A3(new_n855_), .A4(new_n857_), .ZN(new_n858_));
  NOR3_X1    g00794(.A1(new_n437_), .A2(new_n453_), .A3(new_n170_), .ZN(new_n859_));
  NOR3_X1    g00795(.A1(new_n774_), .A2(new_n132_), .A3(new_n192_), .ZN(new_n860_));
  NAND4_X1   g00796(.A1(new_n860_), .A2(new_n657_), .A3(new_n784_), .A4(new_n859_), .ZN(new_n861_));
  INV_X1     g00797(.I(new_n861_), .ZN(new_n862_));
  INV_X1     g00798(.I(new_n218_), .ZN(new_n863_));
  NOR2_X1    g00799(.A1(new_n241_), .A2(new_n92_), .ZN(new_n864_));
  INV_X1     g00800(.I(new_n864_), .ZN(new_n865_));
  INV_X1     g00801(.I(new_n208_), .ZN(new_n866_));
  NOR2_X1    g00802(.A1(new_n334_), .A2(new_n150_), .ZN(new_n867_));
  NOR2_X1    g00803(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1     g00804(.I(new_n868_), .ZN(new_n869_));
  NOR2_X1    g00805(.A1(new_n553_), .A2(new_n721_), .ZN(new_n870_));
  NAND2_X1   g00806(.A1(new_n139_), .A2(new_n156_), .ZN(new_n871_));
  NAND2_X1   g00807(.A1(new_n79_), .A2(new_n140_), .ZN(new_n872_));
  NAND2_X1   g00808(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1     g00809(.I(new_n873_), .ZN(new_n874_));
  NOR2_X1    g00810(.A1(new_n475_), .A2(new_n625_), .ZN(new_n875_));
  NAND4_X1   g00811(.A1(new_n874_), .A2(new_n317_), .A3(new_n870_), .A4(new_n875_), .ZN(new_n876_));
  NOR4_X1    g00812(.A1(new_n876_), .A2(new_n863_), .A3(new_n865_), .A4(new_n869_), .ZN(new_n877_));
  AND2_X2    g00813(.A1(new_n877_), .A2(new_n862_), .Z(new_n878_));
  INV_X1     g00814(.I(new_n597_), .ZN(new_n879_));
  NAND2_X1   g00815(.A1(new_n181_), .A2(new_n77_), .ZN(new_n880_));
  NAND2_X1   g00816(.A1(new_n795_), .A2(new_n880_), .ZN(new_n881_));
  NOR4_X1    g00817(.A1(new_n426_), .A2(new_n879_), .A3(new_n607_), .A4(new_n881_), .ZN(new_n882_));
  INV_X1     g00818(.I(new_n882_), .ZN(new_n883_));
  NOR3_X1    g00819(.A1(new_n734_), .A2(new_n190_), .A3(new_n430_), .ZN(new_n884_));
  INV_X1     g00820(.I(new_n884_), .ZN(new_n885_));
  NOR4_X1    g00821(.A1(new_n751_), .A2(new_n367_), .A3(new_n753_), .A4(new_n640_), .ZN(new_n886_));
  NOR2_X1    g00822(.A1(new_n202_), .A2(new_n637_), .ZN(new_n887_));
  NOR2_X1    g00823(.A1(new_n219_), .A2(new_n791_), .ZN(new_n888_));
  NOR2_X1    g00824(.A1(new_n307_), .A2(new_n741_), .ZN(new_n889_));
  NOR2_X1    g00825(.A1(new_n796_), .A2(new_n684_), .ZN(new_n890_));
  INV_X1     g00826(.I(new_n890_), .ZN(new_n891_));
  NOR4_X1    g00827(.A1(new_n717_), .A2(new_n891_), .A3(new_n552_), .A4(new_n569_), .ZN(new_n892_));
  NAND4_X1   g00828(.A1(new_n892_), .A2(new_n887_), .A3(new_n888_), .A4(new_n889_), .ZN(new_n893_));
  NOR4_X1    g00829(.A1(new_n893_), .A2(new_n883_), .A3(new_n885_), .A4(new_n886_), .ZN(new_n894_));
  NAND4_X1   g00830(.A1(new_n878_), .A2(new_n894_), .A3(new_n831_), .A4(new_n858_), .ZN(new_n895_));
  NOR2_X1    g00831(.A1(new_n895_), .A2(new_n815_), .ZN(new_n896_));
  INV_X1     g00832(.I(new_n896_), .ZN(new_n897_));
  INV_X1     g00833(.I(new_n383_), .ZN(new_n898_));
  NOR2_X1    g00834(.A1(new_n334_), .A2(new_n89_), .ZN(new_n899_));
  NOR2_X1    g00835(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1     g00836(.I(new_n900_), .ZN(new_n901_));
  NOR2_X1    g00837(.A1(new_n69_), .A2(new_n151_), .ZN(new_n902_));
  NOR4_X1    g00838(.A1(new_n901_), .A2(new_n343_), .A3(new_n689_), .A4(new_n902_), .ZN(new_n903_));
  NOR4_X1    g00839(.A1(new_n534_), .A2(new_n260_), .A3(new_n288_), .A4(new_n286_), .ZN(new_n904_));
  INV_X1     g00840(.I(new_n904_), .ZN(new_n905_));
  NOR2_X1    g00841(.A1(new_n101_), .A2(new_n75_), .ZN(new_n906_));
  NOR2_X1    g00842(.A1(new_n593_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1     g00843(.I(new_n907_), .ZN(new_n908_));
  NOR2_X1    g00844(.A1(new_n908_), .A2(new_n670_), .ZN(new_n909_));
  NOR2_X1    g00845(.A1(new_n134_), .A2(new_n153_), .ZN(new_n910_));
  NOR2_X1    g00846(.A1(new_n910_), .A2(new_n370_), .ZN(new_n911_));
  INV_X1     g00847(.I(new_n911_), .ZN(new_n912_));
  INV_X1     g00848(.I(new_n238_), .ZN(new_n913_));
  NAND2_X1   g00849(.A1(new_n913_), .A2(new_n707_), .ZN(new_n914_));
  NOR2_X1    g00850(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  NAND4_X1   g00851(.A1(new_n903_), .A2(new_n905_), .A3(new_n909_), .A4(new_n915_), .ZN(new_n916_));
  NOR4_X1    g00852(.A1(new_n183_), .A2(new_n352_), .A3(new_n791_), .A4(new_n587_), .ZN(new_n917_));
  NOR4_X1    g00853(.A1(new_n602_), .A2(new_n345_), .A3(new_n553_), .A4(new_n268_), .ZN(new_n918_));
  INV_X1     g00854(.I(new_n918_), .ZN(new_n919_));
  NOR4_X1    g00855(.A1(new_n919_), .A2(new_n447_), .A3(new_n576_), .A4(new_n917_), .ZN(new_n920_));
  INV_X1     g00856(.I(new_n920_), .ZN(new_n921_));
  INV_X1     g00857(.I(new_n596_), .ZN(new_n922_));
  NOR2_X1    g00858(.A1(new_n714_), .A2(new_n604_), .ZN(new_n923_));
  NOR2_X1    g00859(.A1(new_n796_), .A2(new_n625_), .ZN(new_n924_));
  NAND4_X1   g00860(.A1(new_n765_), .A2(new_n923_), .A3(new_n924_), .A4(new_n922_), .ZN(new_n925_));
  INV_X1     g00861(.I(new_n925_), .ZN(new_n926_));
  NOR2_X1    g00862(.A1(new_n365_), .A2(new_n772_), .ZN(new_n927_));
  NOR2_X1    g00863(.A1(new_n453_), .A2(new_n330_), .ZN(new_n928_));
  INV_X1     g00864(.I(new_n928_), .ZN(new_n929_));
  NOR2_X1    g00865(.A1(new_n334_), .A2(new_n169_), .ZN(new_n930_));
  NOR2_X1    g00866(.A1(new_n930_), .A2(new_n577_), .ZN(new_n931_));
  INV_X1     g00867(.I(new_n931_), .ZN(new_n932_));
  NOR2_X1    g00868(.A1(new_n932_), .A2(new_n929_), .ZN(new_n933_));
  NAND2_X1   g00869(.A1(new_n284_), .A2(new_n206_), .ZN(new_n934_));
  NAND2_X1   g00870(.A1(new_n221_), .A2(new_n934_), .ZN(new_n935_));
  NOR2_X1    g00871(.A1(new_n611_), .A2(new_n418_), .ZN(new_n936_));
  NOR2_X1    g00872(.A1(new_n85_), .A2(new_n346_), .ZN(new_n937_));
  NOR2_X1    g00873(.A1(new_n517_), .A2(new_n937_), .ZN(new_n938_));
  INV_X1     g00874(.I(new_n938_), .ZN(new_n939_));
  NOR4_X1    g00875(.A1(new_n939_), .A2(new_n805_), .A3(new_n935_), .A4(new_n936_), .ZN(new_n940_));
  NAND4_X1   g00876(.A1(new_n926_), .A2(new_n927_), .A3(new_n940_), .A4(new_n933_), .ZN(new_n941_));
  NOR3_X1    g00877(.A1(new_n916_), .A2(new_n921_), .A3(new_n941_), .ZN(new_n942_));
  INV_X1     g00878(.I(new_n942_), .ZN(new_n943_));
  NOR2_X1    g00879(.A1(new_n175_), .A2(new_n115_), .ZN(new_n944_));
  INV_X1     g00880(.I(new_n551_), .ZN(new_n945_));
  INV_X1     g00881(.I(new_n676_), .ZN(new_n946_));
  NOR2_X1    g00882(.A1(new_n946_), .A2(new_n456_), .ZN(new_n947_));
  INV_X1     g00883(.I(new_n947_), .ZN(new_n948_));
  NOR2_X1    g00884(.A1(new_n948_), .A2(new_n582_), .ZN(new_n949_));
  INV_X1     g00885(.I(new_n949_), .ZN(new_n950_));
  NOR3_X1    g00886(.A1(new_n950_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n951_));
  INV_X1     g00887(.I(new_n951_), .ZN(new_n952_));
  NOR2_X1    g00888(.A1(new_n584_), .A2(new_n92_), .ZN(new_n953_));
  INV_X1     g00889(.I(new_n953_), .ZN(new_n954_));
  NOR2_X1    g00890(.A1(new_n176_), .A2(new_n169_), .ZN(new_n955_));
  NOR2_X1    g00891(.A1(new_n955_), .A2(new_n384_), .ZN(new_n956_));
  NOR2_X1    g00892(.A1(new_n779_), .A2(new_n98_), .ZN(new_n957_));
  INV_X1     g00893(.I(new_n957_), .ZN(new_n958_));
  NOR2_X1    g00894(.A1(new_n232_), .A2(new_n132_), .ZN(new_n959_));
  INV_X1     g00895(.I(new_n959_), .ZN(new_n960_));
  NOR4_X1    g00896(.A1(new_n958_), .A2(new_n954_), .A3(new_n960_), .A4(new_n956_), .ZN(new_n961_));
  NAND2_X1   g00897(.A1(new_n322_), .A2(new_n394_), .ZN(new_n962_));
  NOR2_X1    g00898(.A1(new_n369_), .A2(new_n962_), .ZN(new_n963_));
  NAND4_X1   g00899(.A1(new_n961_), .A2(new_n766_), .A3(new_n828_), .A4(new_n963_), .ZN(new_n964_));
  INV_X1     g00900(.I(new_n753_), .ZN(new_n965_));
  NAND2_X1   g00901(.A1(new_n196_), .A2(new_n273_), .ZN(new_n966_));
  NAND2_X1   g00902(.A1(new_n701_), .A2(new_n966_), .ZN(new_n967_));
  NOR2_X1    g00903(.A1(new_n261_), .A2(new_n320_), .ZN(new_n968_));
  NAND4_X1   g00904(.A1(new_n967_), .A2(new_n968_), .A3(new_n965_), .A4(new_n467_), .ZN(new_n969_));
  NOR3_X1    g00905(.A1(new_n969_), .A2(new_n488_), .A3(new_n565_), .ZN(new_n970_));
  NOR3_X1    g00906(.A1(new_n387_), .A2(new_n719_), .A3(new_n190_), .ZN(new_n971_));
  NOR2_X1    g00907(.A1(new_n697_), .A2(new_n359_), .ZN(new_n972_));
  NOR4_X1    g00908(.A1(new_n656_), .A2(new_n149_), .A3(new_n496_), .A4(new_n770_), .ZN(new_n973_));
  NAND4_X1   g00909(.A1(new_n970_), .A2(new_n971_), .A3(new_n972_), .A4(new_n973_), .ZN(new_n974_));
  NOR3_X1    g00910(.A1(new_n952_), .A2(new_n964_), .A3(new_n974_), .ZN(new_n975_));
  NOR2_X1    g00911(.A1(new_n424_), .A2(new_n211_), .ZN(new_n976_));
  NAND4_X1   g00912(.A1(new_n976_), .A2(new_n507_), .A3(new_n649_), .A4(new_n665_), .ZN(new_n977_));
  NAND2_X1   g00913(.A1(new_n440_), .A2(new_n108_), .ZN(new_n978_));
  INV_X1     g00914(.I(new_n241_), .ZN(new_n979_));
  NAND2_X1   g00915(.A1(new_n156_), .A2(new_n112_), .ZN(new_n980_));
  NAND4_X1   g00916(.A1(new_n979_), .A2(new_n672_), .A3(new_n980_), .A4(new_n978_), .ZN(new_n981_));
  INV_X1     g00917(.I(new_n475_), .ZN(new_n982_));
  NAND2_X1   g00918(.A1(new_n181_), .A2(new_n440_), .ZN(new_n983_));
  NAND2_X1   g00919(.A1(new_n205_), .A2(new_n196_), .ZN(new_n984_));
  NAND2_X1   g00920(.A1(new_n185_), .A2(new_n181_), .ZN(new_n985_));
  NAND4_X1   g00921(.A1(new_n982_), .A2(new_n984_), .A3(new_n985_), .A4(new_n983_), .ZN(new_n986_));
  NOR2_X1    g00922(.A1(new_n633_), .A2(new_n463_), .ZN(new_n987_));
  INV_X1     g00923(.I(new_n987_), .ZN(new_n988_));
  NOR2_X1    g00924(.A1(new_n988_), .A2(new_n154_), .ZN(new_n989_));
  NAND4_X1   g00925(.A1(new_n989_), .A2(new_n283_), .A3(new_n981_), .A4(new_n986_), .ZN(new_n990_));
  NOR2_X1    g00926(.A1(new_n990_), .A2(new_n977_), .ZN(new_n991_));
  NAND2_X1   g00927(.A1(new_n112_), .A2(new_n350_), .ZN(new_n992_));
  NOR2_X1    g00928(.A1(new_n252_), .A2(new_n374_), .ZN(new_n993_));
  INV_X1     g00929(.I(new_n993_), .ZN(new_n994_));
  NOR2_X1    g00930(.A1(new_n752_), .A2(new_n486_), .ZN(new_n995_));
  NOR4_X1    g00931(.A1(new_n994_), .A2(new_n419_), .A3(new_n510_), .A4(new_n995_), .ZN(new_n996_));
  NAND4_X1   g00932(.A1(new_n996_), .A2(new_n113_), .A3(new_n992_), .A4(new_n393_), .ZN(new_n997_));
  INV_X1     g00933(.I(new_n997_), .ZN(new_n998_));
  NAND2_X1   g00934(.A1(new_n404_), .A2(new_n108_), .ZN(new_n999_));
  NOR2_X1    g00935(.A1(new_n541_), .A2(new_n591_), .ZN(new_n1000_));
  NOR2_X1    g00936(.A1(new_n76_), .A2(new_n163_), .ZN(new_n1001_));
  NOR2_X1    g00937(.A1(new_n130_), .A2(new_n736_), .ZN(new_n1002_));
  NAND4_X1   g00938(.A1(new_n1000_), .A2(new_n1001_), .A3(new_n1002_), .A4(new_n999_), .ZN(new_n1003_));
  NOR4_X1    g00939(.A1(new_n326_), .A2(new_n740_), .A3(new_n491_), .A4(new_n556_), .ZN(new_n1004_));
  NOR4_X1    g00940(.A1(new_n406_), .A2(new_n267_), .A3(new_n388_), .A4(new_n684_), .ZN(new_n1005_));
  NOR3_X1    g00941(.A1(new_n1003_), .A2(new_n1004_), .A3(new_n1005_), .ZN(new_n1006_));
  NAND4_X1   g00942(.A1(new_n975_), .A2(new_n991_), .A3(new_n998_), .A4(new_n1006_), .ZN(new_n1007_));
  NOR2_X1    g00943(.A1(new_n1007_), .A2(new_n943_), .ZN(new_n1008_));
  NAND2_X1   g00944(.A1(new_n265_), .A2(new_n350_), .ZN(new_n1009_));
  AND4_X2    g00945(.A1(new_n287_), .A2(new_n820_), .A3(new_n353_), .A4(new_n1009_), .Z(new_n1010_));
  AOI21_X1   g00946(.A1(new_n85_), .A2(new_n105_), .B(new_n150_), .ZN(new_n1011_));
  AOI22_X1   g00947(.A1(new_n205_), .A2(new_n355_), .B1(new_n180_), .B2(new_n230_), .ZN(new_n1012_));
  NOR4_X1    g00948(.A1(new_n251_), .A2(new_n1012_), .A3(new_n260_), .A4(new_n1011_), .ZN(new_n1013_));
  INV_X1     g00949(.I(new_n507_), .ZN(new_n1014_));
  NOR4_X1    g00950(.A1(new_n1014_), .A2(new_n366_), .A3(new_n376_), .A4(new_n430_), .ZN(new_n1015_));
  NAND3_X1   g00951(.A1(new_n1015_), .A2(new_n1010_), .A3(new_n1013_), .ZN(new_n1016_));
  NOR4_X1    g00952(.A1(new_n596_), .A2(new_n782_), .A3(new_n190_), .A4(new_n92_), .ZN(new_n1017_));
  INV_X1     g00953(.I(new_n660_), .ZN(new_n1018_));
  NAND2_X1   g00954(.A1(new_n1018_), .A2(new_n356_), .ZN(new_n1019_));
  INV_X1     g00955(.I(new_n1019_), .ZN(new_n1020_));
  NOR2_X1    g00956(.A1(new_n365_), .A2(new_n370_), .ZN(new_n1021_));
  NAND2_X1   g00957(.A1(new_n1020_), .A2(new_n1021_), .ZN(new_n1022_));
  NOR3_X1    g00958(.A1(new_n515_), .A2(new_n638_), .A3(new_n490_), .ZN(new_n1023_));
  INV_X1     g00959(.I(new_n1023_), .ZN(new_n1024_));
  NAND2_X1   g00960(.A1(new_n230_), .A2(new_n206_), .ZN(new_n1025_));
  INV_X1     g00961(.I(new_n763_), .ZN(new_n1026_));
  NAND2_X1   g00962(.A1(new_n1026_), .A2(new_n1025_), .ZN(new_n1027_));
  NOR3_X1    g00963(.A1(new_n1027_), .A2(new_n573_), .A3(new_n396_), .ZN(new_n1028_));
  NOR4_X1    g00964(.A1(new_n1022_), .A2(new_n1028_), .A3(new_n1017_), .A4(new_n1024_), .ZN(new_n1029_));
  INV_X1     g00965(.I(new_n1029_), .ZN(new_n1030_));
  NOR2_X1    g00966(.A1(new_n171_), .A2(new_n88_), .ZN(new_n1031_));
  NOR4_X1    g00967(.A1(new_n714_), .A2(new_n403_), .A3(new_n1031_), .A4(new_n517_), .ZN(new_n1032_));
  NOR3_X1    g00968(.A1(new_n255_), .A2(new_n447_), .A3(new_n264_), .ZN(new_n1033_));
  INV_X1     g00969(.I(new_n1033_), .ZN(new_n1034_));
  NOR2_X1    g00970(.A1(new_n115_), .A2(new_n346_), .ZN(new_n1035_));
  NOR2_X1    g00971(.A1(new_n359_), .A2(new_n1035_), .ZN(new_n1036_));
  INV_X1     g00972(.I(new_n1036_), .ZN(new_n1037_));
  NOR2_X1    g00973(.A1(new_n496_), .A2(new_n183_), .ZN(new_n1038_));
  INV_X1     g00974(.I(new_n1038_), .ZN(new_n1039_));
  NOR4_X1    g00975(.A1(new_n1034_), .A2(new_n1037_), .A3(new_n1039_), .A4(new_n1032_), .ZN(new_n1040_));
  INV_X1     g00976(.I(new_n1040_), .ZN(new_n1041_));
  NOR3_X1    g00977(.A1(new_n544_), .A2(new_n191_), .A3(new_n482_), .ZN(new_n1042_));
  INV_X1     g00978(.I(new_n875_), .ZN(new_n1043_));
  NOR2_X1    g00979(.A1(new_n289_), .A2(new_n154_), .ZN(new_n1044_));
  INV_X1     g00980(.I(new_n1044_), .ZN(new_n1045_));
  NOR2_X1    g00981(.A1(new_n1043_), .A2(new_n1045_), .ZN(new_n1046_));
  NOR3_X1    g00982(.A1(new_n164_), .A2(new_n282_), .A3(new_n262_), .ZN(new_n1047_));
  INV_X1     g00983(.I(new_n222_), .ZN(new_n1048_));
  NOR3_X1    g00984(.A1(new_n1048_), .A2(new_n689_), .A3(new_n776_), .ZN(new_n1049_));
  NAND4_X1   g00985(.A1(new_n1046_), .A2(new_n1042_), .A3(new_n1047_), .A4(new_n1049_), .ZN(new_n1050_));
  NOR4_X1    g00986(.A1(new_n1030_), .A2(new_n1016_), .A3(new_n1041_), .A4(new_n1050_), .ZN(new_n1051_));
  INV_X1     g00987(.I(new_n1051_), .ZN(new_n1052_));
  AOI22_X1   g00988(.A1(new_n275_), .A2(new_n265_), .B1(new_n139_), .B2(new_n350_), .ZN(new_n1053_));
  AOI22_X1   g00989(.A1(new_n142_), .A2(new_n230_), .B1(new_n139_), .B2(new_n440_), .ZN(new_n1054_));
  AOI21_X1   g00990(.A1(new_n334_), .A2(new_n85_), .B(new_n131_), .ZN(new_n1055_));
  NOR3_X1    g00991(.A1(new_n1053_), .A2(new_n1054_), .A3(new_n1055_), .ZN(new_n1056_));
  NOR3_X1    g00992(.A1(new_n137_), .A2(new_n485_), .A3(new_n682_), .ZN(new_n1057_));
  NAND2_X1   g00993(.A1(new_n159_), .A2(new_n270_), .ZN(new_n1058_));
  NAND2_X1   g00994(.A1(new_n109_), .A2(new_n273_), .ZN(new_n1059_));
  NAND4_X1   g00995(.A1(new_n1058_), .A2(new_n854_), .A3(new_n980_), .A4(new_n1059_), .ZN(new_n1060_));
  NOR3_X1    g00996(.A1(new_n615_), .A2(new_n703_), .A3(new_n70_), .ZN(new_n1061_));
  NAND4_X1   g00997(.A1(new_n1056_), .A2(new_n1057_), .A3(new_n1060_), .A4(new_n1061_), .ZN(new_n1062_));
  NAND2_X1   g00998(.A1(new_n284_), .A2(new_n350_), .ZN(new_n1063_));
  NAND4_X1   g00999(.A1(new_n992_), .A2(new_n1063_), .A3(new_n391_), .A4(new_n471_), .ZN(new_n1064_));
  NAND2_X1   g01000(.A1(new_n205_), .A2(new_n156_), .ZN(new_n1065_));
  NAND2_X1   g01001(.A1(new_n275_), .A2(new_n143_), .ZN(new_n1066_));
  NAND2_X1   g01002(.A1(new_n142_), .A2(new_n112_), .ZN(new_n1067_));
  NAND2_X1   g01003(.A1(new_n111_), .A2(new_n108_), .ZN(new_n1068_));
  NAND4_X1   g01004(.A1(new_n1065_), .A2(new_n1066_), .A3(new_n1067_), .A4(new_n1068_), .ZN(new_n1069_));
  NAND2_X1   g01005(.A1(new_n205_), .A2(new_n142_), .ZN(new_n1070_));
  NAND4_X1   g01006(.A1(new_n662_), .A2(new_n409_), .A3(new_n1070_), .A4(new_n983_), .ZN(new_n1071_));
  NAND3_X1   g01007(.A1(new_n1069_), .A2(new_n1071_), .A3(new_n1064_), .ZN(new_n1072_));
  NOR2_X1    g01008(.A1(new_n129_), .A2(new_n148_), .ZN(new_n1073_));
  NOR3_X1    g01009(.A1(new_n640_), .A2(new_n1073_), .A3(new_n306_), .ZN(new_n1074_));
  NOR2_X1    g01010(.A1(new_n654_), .A2(new_n610_), .ZN(new_n1075_));
  AOI21_X1   g01011(.A1(new_n105_), .A2(new_n176_), .B(new_n83_), .ZN(new_n1076_));
  NOR3_X1    g01012(.A1(new_n1076_), .A2(new_n561_), .A3(new_n744_), .ZN(new_n1077_));
  AOI22_X1   g01013(.A1(new_n142_), .A2(new_n245_), .B1(new_n270_), .B2(new_n109_), .ZN(new_n1078_));
  AOI21_X1   g01014(.A1(new_n115_), .A2(new_n88_), .B(new_n123_), .ZN(new_n1079_));
  NOR2_X1    g01015(.A1(new_n1078_), .A2(new_n1079_), .ZN(new_n1080_));
  NAND4_X1   g01016(.A1(new_n1080_), .A2(new_n1077_), .A3(new_n1074_), .A4(new_n1075_), .ZN(new_n1081_));
  NOR3_X1    g01017(.A1(new_n1062_), .A2(new_n1072_), .A3(new_n1081_), .ZN(new_n1082_));
  NOR4_X1    g01018(.A1(new_n465_), .A2(new_n548_), .A3(new_n345_), .A4(new_n152_), .ZN(new_n1083_));
  INV_X1     g01019(.I(new_n501_), .ZN(new_n1084_));
  NOR4_X1    g01020(.A1(new_n326_), .A2(new_n1084_), .A3(new_n252_), .A4(new_n648_), .ZN(new_n1085_));
  NOR2_X1    g01021(.A1(new_n604_), .A2(new_n731_), .ZN(new_n1086_));
  INV_X1     g01022(.I(new_n1086_), .ZN(new_n1087_));
  INV_X1     g01023(.I(new_n518_), .ZN(new_n1088_));
  NAND2_X1   g01024(.A1(new_n1088_), .A2(new_n509_), .ZN(new_n1089_));
  NOR4_X1    g01025(.A1(new_n1085_), .A2(new_n1083_), .A3(new_n1087_), .A4(new_n1089_), .ZN(new_n1090_));
  NAND2_X1   g01026(.A1(new_n245_), .A2(new_n185_), .ZN(new_n1091_));
  NOR2_X1    g01027(.A1(new_n116_), .A2(new_n153_), .ZN(new_n1092_));
  NOR3_X1    g01028(.A1(new_n132_), .A2(new_n1092_), .A3(new_n397_), .ZN(new_n1093_));
  NAND3_X1   g01029(.A1(new_n1093_), .A2(new_n1091_), .A3(new_n313_), .ZN(new_n1094_));
  NAND2_X1   g01030(.A1(new_n185_), .A2(new_n273_), .ZN(new_n1095_));
  NAND2_X1   g01031(.A1(new_n230_), .A2(new_n77_), .ZN(new_n1096_));
  NAND2_X1   g01032(.A1(new_n1095_), .A2(new_n1096_), .ZN(new_n1097_));
  NAND3_X1   g01033(.A1(new_n852_), .A2(new_n1097_), .A3(new_n511_), .ZN(new_n1098_));
  NOR2_X1    g01034(.A1(new_n1098_), .A2(new_n1094_), .ZN(new_n1099_));
  NAND2_X1   g01035(.A1(new_n79_), .A2(new_n109_), .ZN(new_n1100_));
  NAND2_X1   g01036(.A1(new_n85_), .A2(new_n66_), .ZN(new_n1101_));
  AOI22_X1   g01037(.A1(new_n1100_), .A2(new_n362_), .B1(new_n1101_), .B2(new_n185_), .ZN(new_n1102_));
  AOI22_X1   g01038(.A1(new_n142_), .A2(new_n181_), .B1(new_n270_), .B2(new_n440_), .ZN(new_n1103_));
  NOR3_X1    g01039(.A1(new_n1103_), .A2(new_n801_), .A3(new_n577_), .ZN(new_n1104_));
  NAND2_X1   g01040(.A1(new_n404_), .A2(new_n205_), .ZN(new_n1105_));
  INV_X1     g01041(.I(new_n594_), .ZN(new_n1106_));
  NAND4_X1   g01042(.A1(new_n1106_), .A2(new_n1105_), .A3(new_n871_), .A4(new_n508_), .ZN(new_n1107_));
  AOI21_X1   g01043(.A1(new_n395_), .A2(new_n999_), .B(new_n268_), .ZN(new_n1108_));
  NAND4_X1   g01044(.A1(new_n1104_), .A2(new_n1107_), .A3(new_n1102_), .A4(new_n1108_), .ZN(new_n1109_));
  INV_X1     g01045(.I(new_n422_), .ZN(new_n1110_));
  NOR2_X1    g01046(.A1(new_n656_), .A2(new_n488_), .ZN(new_n1111_));
  NOR2_X1    g01047(.A1(new_n214_), .A2(new_n459_), .ZN(new_n1112_));
  NOR2_X1    g01048(.A1(new_n127_), .A2(new_n1112_), .ZN(new_n1113_));
  NOR4_X1    g01049(.A1(new_n406_), .A2(new_n491_), .A3(new_n930_), .A4(new_n741_), .ZN(new_n1114_));
  NOR2_X1    g01050(.A1(new_n487_), .A2(new_n468_), .ZN(new_n1115_));
  INV_X1     g01051(.I(new_n1115_), .ZN(new_n1116_));
  NOR4_X1    g01052(.A1(new_n1114_), .A2(new_n1116_), .A3(new_n81_), .A4(new_n752_), .ZN(new_n1117_));
  NAND4_X1   g01053(.A1(new_n1117_), .A2(new_n1110_), .A3(new_n1111_), .A4(new_n1113_), .ZN(new_n1118_));
  NOR2_X1    g01054(.A1(new_n1118_), .A2(new_n1109_), .ZN(new_n1119_));
  NAND4_X1   g01055(.A1(new_n1119_), .A2(new_n1082_), .A3(new_n1090_), .A4(new_n1099_), .ZN(new_n1120_));
  NOR2_X1    g01056(.A1(new_n1052_), .A2(new_n1120_), .ZN(new_n1121_));
  INV_X1     g01057(.I(new_n1121_), .ZN(new_n1122_));
  NOR4_X1    g01058(.A1(new_n587_), .A2(new_n841_), .A3(new_n937_), .A4(new_n280_), .ZN(new_n1123_));
  INV_X1     g01059(.I(new_n1123_), .ZN(new_n1124_));
  NOR3_X1    g01060(.A1(new_n225_), .A2(new_n899_), .A3(new_n804_), .ZN(new_n1125_));
  NOR2_X1    g01061(.A1(new_n791_), .A2(new_n1035_), .ZN(new_n1126_));
  NOR2_X1    g01062(.A1(new_n633_), .A2(new_n719_), .ZN(new_n1127_));
  NAND4_X1   g01063(.A1(new_n1124_), .A2(new_n1125_), .A3(new_n1126_), .A4(new_n1127_), .ZN(new_n1128_));
  INV_X1     g01064(.I(new_n459_), .ZN(new_n1129_));
  NOR2_X1    g01065(.A1(new_n695_), .A2(new_n703_), .ZN(new_n1130_));
  NAND4_X1   g01066(.A1(new_n1130_), .A2(new_n383_), .A3(new_n1129_), .A4(new_n966_), .ZN(new_n1131_));
  NOR4_X1    g01067(.A1(new_n593_), .A2(new_n242_), .A3(new_n312_), .A4(new_n660_), .ZN(new_n1132_));
  NOR2_X1    g01068(.A1(new_n247_), .A2(new_n764_), .ZN(new_n1133_));
  INV_X1     g01069(.I(new_n1133_), .ZN(new_n1134_));
  NOR4_X1    g01070(.A1(new_n1132_), .A2(new_n288_), .A3(new_n796_), .A4(new_n1134_), .ZN(new_n1135_));
  INV_X1     g01071(.I(new_n1135_), .ZN(new_n1136_));
  INV_X1     g01072(.I(new_n683_), .ZN(new_n1137_));
  NOR2_X1    g01073(.A1(new_n175_), .A2(new_n105_), .ZN(new_n1138_));
  NOR2_X1    g01074(.A1(new_n817_), .A2(new_n1138_), .ZN(new_n1139_));
  NOR3_X1    g01075(.A1(new_n932_), .A2(new_n1137_), .A3(new_n1139_), .ZN(new_n1140_));
  INV_X1     g01076(.I(new_n1140_), .ZN(new_n1141_));
  NOR4_X1    g01077(.A1(new_n1136_), .A2(new_n1128_), .A3(new_n1131_), .A4(new_n1141_), .ZN(new_n1142_));
  NOR4_X1    g01078(.A1(new_n446_), .A2(new_n211_), .A3(new_n324_), .A4(new_n491_), .ZN(new_n1143_));
  NOR2_X1    g01079(.A1(new_n698_), .A2(new_n867_), .ZN(new_n1144_));
  INV_X1     g01080(.I(new_n1144_), .ZN(new_n1145_));
  NOR2_X1    g01081(.A1(new_n73_), .A2(new_n89_), .ZN(new_n1146_));
  NOR2_X1    g01082(.A1(new_n1146_), .A2(new_n420_), .ZN(new_n1147_));
  NOR3_X1    g01083(.A1(new_n1143_), .A2(new_n1145_), .A3(new_n1147_), .ZN(new_n1148_));
  INV_X1     g01084(.I(new_n775_), .ZN(new_n1149_));
  NOR2_X1    g01085(.A1(new_n666_), .A2(new_n198_), .ZN(new_n1150_));
  INV_X1     g01086(.I(new_n1150_), .ZN(new_n1151_));
  NOR2_X1    g01087(.A1(new_n334_), .A2(new_n129_), .ZN(new_n1152_));
  NOR2_X1    g01088(.A1(new_n294_), .A2(new_n1152_), .ZN(new_n1153_));
  INV_X1     g01089(.I(new_n1153_), .ZN(new_n1154_));
  NOR4_X1    g01090(.A1(new_n1149_), .A2(new_n844_), .A3(new_n1151_), .A4(new_n1154_), .ZN(new_n1155_));
  NOR2_X1    g01091(.A1(new_n498_), .A2(new_n902_), .ZN(new_n1156_));
  INV_X1     g01092(.I(new_n1156_), .ZN(new_n1157_));
  NAND2_X1   g01093(.A1(new_n321_), .A2(new_n311_), .ZN(new_n1158_));
  NOR2_X1    g01094(.A1(new_n1084_), .A2(new_n736_), .ZN(new_n1159_));
  INV_X1     g01095(.I(new_n1159_), .ZN(new_n1160_));
  NAND2_X1   g01096(.A1(new_n377_), .A2(new_n512_), .ZN(new_n1161_));
  NOR4_X1    g01097(.A1(new_n1160_), .A2(new_n1158_), .A3(new_n1157_), .A4(new_n1161_), .ZN(new_n1162_));
  NAND3_X1   g01098(.A1(new_n1155_), .A2(new_n1162_), .A3(new_n1148_), .ZN(new_n1163_));
  INV_X1     g01099(.I(new_n822_), .ZN(new_n1164_));
  NOR2_X1    g01100(.A1(new_n644_), .A2(new_n752_), .ZN(new_n1165_));
  NOR2_X1    g01101(.A1(new_n367_), .A2(new_n227_), .ZN(new_n1166_));
  NOR2_X1    g01102(.A1(new_n75_), .A2(new_n66_), .ZN(new_n1167_));
  NOR2_X1    g01103(.A1(new_n89_), .A2(new_n122_), .ZN(new_n1168_));
  NOR4_X1    g01104(.A1(new_n1031_), .A2(new_n783_), .A3(new_n1168_), .A4(new_n1167_), .ZN(new_n1169_));
  NOR4_X1    g01105(.A1(new_n1169_), .A2(new_n214_), .A3(new_n326_), .A4(new_n837_), .ZN(new_n1170_));
  NAND4_X1   g01106(.A1(new_n1170_), .A2(new_n1164_), .A3(new_n1165_), .A4(new_n1166_), .ZN(new_n1171_));
  AOI22_X1   g01107(.A1(new_n205_), .A2(new_n109_), .B1(new_n143_), .B2(new_n206_), .ZN(new_n1172_));
  NOR2_X1    g01108(.A1(new_n866_), .A2(new_n1172_), .ZN(new_n1173_));
  NOR3_X1    g01109(.A1(new_n345_), .A2(new_n582_), .A3(new_n610_), .ZN(new_n1174_));
  NOR2_X1    g01110(.A1(new_n171_), .A2(new_n148_), .ZN(new_n1175_));
  NOR2_X1    g01111(.A1(new_n553_), .A2(new_n1175_), .ZN(new_n1176_));
  NAND4_X1   g01112(.A1(new_n1173_), .A2(new_n1174_), .A3(new_n669_), .A4(new_n1176_), .ZN(new_n1177_));
  NOR3_X1    g01113(.A1(new_n1163_), .A2(new_n1171_), .A3(new_n1177_), .ZN(new_n1178_));
  NAND2_X1   g01114(.A1(new_n1178_), .A2(new_n1142_), .ZN(new_n1179_));
  NOR2_X1    g01115(.A1(new_n1179_), .A2(new_n168_), .ZN(new_n1180_));
  INV_X1     g01116(.I(new_n1180_), .ZN(new_n1181_));
  NOR3_X1    g01117(.A1(new_n618_), .A2(new_n316_), .A3(new_n670_), .ZN(new_n1182_));
  AOI21_X1   g01118(.A1(new_n97_), .A2(new_n169_), .B(new_n176_), .ZN(new_n1183_));
  AOI21_X1   g01119(.A1(new_n118_), .A2(new_n153_), .B(new_n83_), .ZN(new_n1184_));
  AOI21_X1   g01120(.A1(new_n115_), .A2(new_n148_), .B(new_n131_), .ZN(new_n1185_));
  AOI21_X1   g01121(.A1(new_n89_), .A2(new_n134_), .B(new_n334_), .ZN(new_n1186_));
  NOR4_X1    g01122(.A1(new_n1183_), .A2(new_n1186_), .A3(new_n1184_), .A4(new_n1185_), .ZN(new_n1187_));
  NAND3_X1   g01123(.A1(new_n1013_), .A2(new_n1187_), .A3(new_n1182_), .ZN(new_n1188_));
  NAND2_X1   g01124(.A1(new_n79_), .A2(new_n440_), .ZN(new_n1189_));
  NAND2_X1   g01125(.A1(new_n205_), .A2(new_n185_), .ZN(new_n1190_));
  NAND4_X1   g01126(.A1(new_n479_), .A2(new_n272_), .A3(new_n1190_), .A4(new_n1189_), .ZN(new_n1191_));
  NAND2_X1   g01127(.A1(new_n112_), .A2(new_n185_), .ZN(new_n1192_));
  NAND4_X1   g01128(.A1(new_n823_), .A2(new_n1192_), .A3(new_n807_), .A4(new_n356_), .ZN(new_n1193_));
  NOR2_X1    g01129(.A1(new_n236_), .A2(new_n242_), .ZN(new_n1194_));
  NAND4_X1   g01130(.A1(new_n1191_), .A2(new_n1193_), .A3(new_n643_), .A4(new_n1194_), .ZN(new_n1195_));
  NOR3_X1    g01131(.A1(new_n1188_), .A2(new_n1109_), .A3(new_n1195_), .ZN(new_n1196_));
  INV_X1     g01132(.I(new_n765_), .ZN(new_n1197_));
  INV_X1     g01133(.I(new_n859_), .ZN(new_n1198_));
  AOI22_X1   g01134(.A1(new_n196_), .A2(new_n112_), .B1(new_n181_), .B2(new_n206_), .ZN(new_n1199_));
  INV_X1     g01135(.I(new_n1199_), .ZN(new_n1200_));
  NOR4_X1    g01136(.A1(new_n1198_), .A2(new_n1197_), .A3(new_n1200_), .A4(new_n518_), .ZN(new_n1201_));
  NOR4_X1    g01137(.A1(new_n326_), .A2(new_n211_), .A3(new_n288_), .A4(new_n681_), .ZN(new_n1202_));
  NOR4_X1    g01138(.A1(new_n751_), .A2(new_n703_), .A3(new_n561_), .A4(new_n376_), .ZN(new_n1203_));
  NOR2_X1    g01139(.A1(new_n1202_), .A2(new_n1203_), .ZN(new_n1204_));
  NOR2_X1    g01140(.A1(new_n1146_), .A2(new_n796_), .ZN(new_n1205_));
  INV_X1     g01141(.I(new_n1205_), .ZN(new_n1206_));
  NOR2_X1    g01142(.A1(new_n1206_), .A2(new_n281_), .ZN(new_n1207_));
  NOR3_X1    g01143(.A1(new_n642_), .A2(new_n297_), .A3(new_n607_), .ZN(new_n1208_));
  NAND3_X1   g01144(.A1(new_n1204_), .A2(new_n1208_), .A3(new_n1207_), .ZN(new_n1209_));
  NAND2_X1   g01145(.A1(new_n680_), .A2(new_n598_), .ZN(new_n1210_));
  INV_X1     g01146(.I(new_n1210_), .ZN(new_n1211_));
  NAND2_X1   g01147(.A1(new_n284_), .A2(new_n185_), .ZN(new_n1212_));
  NAND2_X1   g01148(.A1(new_n342_), .A2(new_n1212_), .ZN(new_n1213_));
  INV_X1     g01149(.I(new_n1213_), .ZN(new_n1214_));
  NAND2_X1   g01150(.A1(new_n1214_), .A2(new_n1097_), .ZN(new_n1215_));
  NAND2_X1   g01151(.A1(new_n140_), .A2(new_n108_), .ZN(new_n1216_));
  AOI21_X1   g01152(.A1(new_n385_), .A2(new_n501_), .B(new_n732_), .ZN(new_n1217_));
  NAND4_X1   g01153(.A1(new_n1217_), .A2(new_n536_), .A3(new_n1216_), .A4(new_n287_), .ZN(new_n1218_));
  NOR4_X1    g01154(.A1(new_n1209_), .A2(new_n1211_), .A3(new_n1215_), .A4(new_n1218_), .ZN(new_n1219_));
  NAND2_X1   g01155(.A1(new_n1219_), .A2(new_n1201_), .ZN(new_n1220_));
  INV_X1     g01156(.I(new_n264_), .ZN(new_n1221_));
  INV_X1     g01157(.I(new_n498_), .ZN(new_n1222_));
  NOR3_X1    g01158(.A1(new_n774_), .A2(new_n937_), .A3(new_n660_), .ZN(new_n1223_));
  NAND4_X1   g01159(.A1(new_n1223_), .A2(new_n1221_), .A3(new_n1222_), .A4(new_n701_), .ZN(new_n1224_));
  NOR4_X1    g01160(.A1(new_n217_), .A2(new_n486_), .A3(new_n734_), .A4(new_n282_), .ZN(new_n1225_));
  INV_X1     g01161(.I(new_n1225_), .ZN(new_n1226_));
  NOR3_X1    g01162(.A1(new_n714_), .A2(new_n574_), .A3(new_n776_), .ZN(new_n1227_));
  NAND2_X1   g01163(.A1(new_n1226_), .A2(new_n1227_), .ZN(new_n1228_));
  NOR2_X1    g01164(.A1(new_n788_), .A2(new_n235_), .ZN(new_n1229_));
  INV_X1     g01165(.I(new_n1176_), .ZN(new_n1230_));
  AOI21_X1   g01166(.A1(new_n1229_), .A2(new_n165_), .B(new_n1230_), .ZN(new_n1231_));
  NOR4_X1    g01167(.A1(new_n617_), .A2(new_n637_), .A3(new_n756_), .A4(new_n1168_), .ZN(new_n1232_));
  NAND2_X1   g01168(.A1(new_n1232_), .A2(new_n1231_), .ZN(new_n1233_));
  OR3_X2     g01169(.A1(new_n1233_), .A2(new_n1224_), .A3(new_n1228_), .Z(new_n1234_));
  NOR3_X1    g01170(.A1(new_n837_), .A2(new_n719_), .A3(new_n590_), .ZN(new_n1235_));
  NOR2_X1    g01171(.A1(new_n134_), .A2(new_n122_), .ZN(new_n1236_));
  NOR2_X1    g01172(.A1(new_n463_), .A2(new_n1236_), .ZN(new_n1237_));
  NAND4_X1   g01173(.A1(new_n739_), .A2(new_n840_), .A3(new_n809_), .A4(new_n1059_), .ZN(new_n1238_));
  NAND3_X1   g01174(.A1(new_n1238_), .A2(new_n1235_), .A3(new_n1237_), .ZN(new_n1239_));
  NOR4_X1    g01175(.A1(new_n1220_), .A2(new_n1118_), .A3(new_n1234_), .A4(new_n1239_), .ZN(new_n1240_));
  NAND2_X1   g01176(.A1(new_n1240_), .A2(new_n1196_), .ZN(new_n1241_));
  NOR2_X1    g01177(.A1(new_n721_), .A2(new_n280_), .ZN(new_n1242_));
  INV_X1     g01178(.I(new_n1242_), .ZN(new_n1243_));
  NAND2_X1   g01179(.A1(new_n410_), .A2(new_n676_), .ZN(new_n1244_));
  INV_X1     g01180(.I(new_n1244_), .ZN(new_n1245_));
  NOR2_X1    g01181(.A1(new_n241_), .A2(new_n749_), .ZN(new_n1246_));
  NAND2_X1   g01182(.A1(new_n808_), .A2(new_n394_), .ZN(new_n1247_));
  INV_X1     g01183(.I(new_n1247_), .ZN(new_n1248_));
  NAND2_X1   g01184(.A1(new_n1248_), .A2(new_n1246_), .ZN(new_n1249_));
  NAND3_X1   g01185(.A1(new_n627_), .A2(new_n686_), .A3(new_n144_), .ZN(new_n1250_));
  NOR4_X1    g01186(.A1(new_n202_), .A2(new_n347_), .A3(new_n374_), .A4(new_n1035_), .ZN(new_n1251_));
  OR3_X2     g01187(.A1(new_n1024_), .A2(new_n1250_), .A3(new_n1251_), .Z(new_n1252_));
  NOR4_X1    g01188(.A1(new_n1252_), .A2(new_n1243_), .A3(new_n1245_), .A4(new_n1249_), .ZN(new_n1253_));
  NOR3_X1    g01189(.A1(new_n697_), .A2(new_n117_), .A3(new_n130_), .ZN(new_n1254_));
  INV_X1     g01190(.I(new_n1254_), .ZN(new_n1255_));
  NOR2_X1    g01191(.A1(new_n593_), .A2(new_n930_), .ZN(new_n1256_));
  INV_X1     g01192(.I(new_n1256_), .ZN(new_n1257_));
  NOR2_X1    g01193(.A1(new_n1257_), .A2(new_n236_), .ZN(new_n1258_));
  INV_X1     g01194(.I(new_n1258_), .ZN(new_n1259_));
  NOR4_X1    g01195(.A1(new_n183_), .A2(new_n288_), .A3(new_n298_), .A4(new_n510_), .ZN(new_n1260_));
  NOR4_X1    g01196(.A1(new_n1259_), .A2(new_n1198_), .A3(new_n1255_), .A4(new_n1260_), .ZN(new_n1261_));
  INV_X1     g01197(.I(new_n436_), .ZN(new_n1262_));
  NOR2_X1    g01198(.A1(new_n1262_), .A2(new_n330_), .ZN(new_n1263_));
  INV_X1     g01199(.I(new_n888_), .ZN(new_n1264_));
  NOR2_X1    g01200(.A1(new_n447_), .A2(new_n753_), .ZN(new_n1265_));
  INV_X1     g01201(.I(new_n1265_), .ZN(new_n1266_));
  NOR2_X1    g01202(.A1(new_n1266_), .A2(new_n1264_), .ZN(new_n1267_));
  NOR4_X1    g01203(.A1(new_n198_), .A2(new_n172_), .A3(new_n164_), .A4(new_n715_), .ZN(new_n1268_));
  NOR3_X1    g01204(.A1(new_n337_), .A2(new_n463_), .A3(new_n320_), .ZN(new_n1269_));
  NAND4_X1   g01205(.A1(new_n1267_), .A2(new_n1269_), .A3(new_n1263_), .A4(new_n1268_), .ZN(new_n1270_));
  INV_X1     g01206(.I(new_n1270_), .ZN(new_n1271_));
  NOR4_X1    g01207(.A1(new_n81_), .A2(new_n225_), .A3(new_n456_), .A4(new_n1236_), .ZN(new_n1272_));
  NOR2_X1    g01208(.A1(new_n1272_), .A2(new_n785_), .ZN(new_n1273_));
  INV_X1     g01209(.I(new_n1273_), .ZN(new_n1274_));
  NOR2_X1    g01210(.A1(new_n505_), .A2(new_n217_), .ZN(new_n1275_));
  INV_X1     g01211(.I(new_n1275_), .ZN(new_n1276_));
  NOR3_X1    g01212(.A1(new_n426_), .A2(new_n681_), .A3(new_n1276_), .ZN(new_n1277_));
  INV_X1     g01213(.I(new_n1277_), .ZN(new_n1278_));
  NOR2_X1    g01214(.A1(new_n1278_), .A2(new_n1274_), .ZN(new_n1279_));
  NAND4_X1   g01215(.A1(new_n1261_), .A2(new_n1253_), .A3(new_n1279_), .A4(new_n1271_), .ZN(new_n1280_));
  NOR2_X1    g01216(.A1(new_n400_), .A2(new_n366_), .ZN(new_n1281_));
  NOR2_X1    g01217(.A1(new_n251_), .A2(new_n718_), .ZN(new_n1282_));
  NAND3_X1   g01218(.A1(new_n1282_), .A2(new_n982_), .A3(new_n568_), .ZN(new_n1283_));
  NOR3_X1    g01219(.A1(new_n326_), .A2(new_n488_), .A3(new_n498_), .ZN(new_n1284_));
  AND3_X2    g01220(.A1(new_n1283_), .A2(new_n1281_), .A3(new_n1284_), .Z(new_n1285_));
  NOR4_X1    g01221(.A1(new_n343_), .A2(new_n214_), .A3(new_n239_), .A4(new_n247_), .ZN(new_n1286_));
  NOR3_X1    g01222(.A1(new_n1286_), .A2(new_n633_), .A3(new_n1073_), .ZN(new_n1287_));
  NOR2_X1    g01223(.A1(new_n495_), .A2(new_n1167_), .ZN(new_n1288_));
  INV_X1     g01224(.I(new_n1288_), .ZN(new_n1289_));
  NOR4_X1    g01225(.A1(new_n1289_), .A2(new_n1045_), .A3(new_n76_), .A4(new_n387_), .ZN(new_n1290_));
  NOR3_X1    g01226(.A1(new_n267_), .A2(new_n294_), .A3(new_n763_), .ZN(new_n1291_));
  NOR3_X1    g01227(.A1(new_n136_), .A2(new_n235_), .A3(new_n419_), .ZN(new_n1292_));
  NAND4_X1   g01228(.A1(new_n1291_), .A2(new_n1292_), .A3(new_n246_), .A4(new_n382_), .ZN(new_n1293_));
  NOR3_X1    g01229(.A1(new_n191_), .A2(new_n517_), .A3(new_n430_), .ZN(new_n1294_));
  NAND4_X1   g01230(.A1(new_n667_), .A2(new_n992_), .A3(new_n362_), .A4(new_n842_), .ZN(new_n1295_));
  NOR3_X1    g01231(.A1(new_n406_), .A2(new_n211_), .A3(new_n604_), .ZN(new_n1296_));
  NAND4_X1   g01232(.A1(new_n1295_), .A2(new_n1205_), .A3(new_n1294_), .A4(new_n1296_), .ZN(new_n1297_));
  NOR2_X1    g01233(.A1(new_n1297_), .A2(new_n1293_), .ZN(new_n1298_));
  NAND4_X1   g01234(.A1(new_n1298_), .A2(new_n1285_), .A3(new_n1287_), .A4(new_n1290_), .ZN(new_n1299_));
  NOR4_X1    g01235(.A1(new_n1019_), .A2(new_n305_), .A3(new_n1138_), .A4(new_n822_), .ZN(new_n1300_));
  INV_X1     g01236(.I(new_n1300_), .ZN(new_n1301_));
  NOR4_X1    g01237(.A1(new_n955_), .A2(new_n779_), .A3(new_n587_), .A4(new_n1168_), .ZN(new_n1302_));
  NOR3_X1    g01238(.A1(new_n591_), .A2(new_n173_), .A3(new_n152_), .ZN(new_n1303_));
  INV_X1     g01239(.I(new_n1303_), .ZN(new_n1304_));
  INV_X1     g01240(.I(new_n506_), .ZN(new_n1305_));
  NAND3_X1   g01241(.A1(new_n1305_), .A2(new_n160_), .A3(new_n508_), .ZN(new_n1306_));
  NOR4_X1    g01242(.A1(new_n1301_), .A2(new_n1302_), .A3(new_n1304_), .A4(new_n1306_), .ZN(new_n1307_));
  INV_X1     g01243(.I(new_n1307_), .ZN(new_n1308_));
  NOR4_X1    g01244(.A1(new_n106_), .A2(new_n611_), .A3(new_n190_), .A4(new_n264_), .ZN(new_n1309_));
  INV_X1     g01245(.I(new_n1309_), .ZN(new_n1310_));
  INV_X1     g01246(.I(new_n252_), .ZN(new_n1311_));
  NAND4_X1   g01247(.A1(new_n1311_), .A2(new_n157_), .A3(new_n984_), .A4(new_n999_), .ZN(new_n1312_));
  NAND3_X1   g01248(.A1(new_n1310_), .A2(new_n1312_), .A3(new_n775_), .ZN(new_n1313_));
  NAND2_X1   g01249(.A1(new_n318_), .A2(new_n275_), .ZN(new_n1314_));
  INV_X1     g01250(.I(new_n345_), .ZN(new_n1315_));
  NAND4_X1   g01251(.A1(new_n1315_), .A2(new_n1314_), .A3(new_n391_), .A4(new_n854_), .ZN(new_n1316_));
  NOR4_X1    g01252(.A1(new_n147_), .A2(new_n163_), .A3(new_n670_), .A4(new_n286_), .ZN(new_n1317_));
  NOR2_X1    g01253(.A1(new_n203_), .A2(new_n531_), .ZN(new_n1318_));
  NOR2_X1    g01254(.A1(new_n535_), .A2(new_n1092_), .ZN(new_n1319_));
  NAND4_X1   g01255(.A1(new_n1316_), .A2(new_n1317_), .A3(new_n1318_), .A4(new_n1319_), .ZN(new_n1320_));
  INV_X1     g01256(.I(new_n618_), .ZN(new_n1321_));
  NAND2_X1   g01257(.A1(new_n158_), .A2(new_n350_), .ZN(new_n1322_));
  NAND2_X1   g01258(.A1(new_n451_), .A2(new_n1322_), .ZN(new_n1323_));
  NOR4_X1    g01259(.A1(new_n1323_), .A2(new_n561_), .A3(new_n744_), .A4(new_n1076_), .ZN(new_n1324_));
  NAND2_X1   g01260(.A1(new_n180_), .A2(new_n108_), .ZN(new_n1325_));
  NAND2_X1   g01261(.A1(new_n832_), .A2(new_n1325_), .ZN(new_n1326_));
  NAND2_X1   g01262(.A1(new_n318_), .A2(new_n185_), .ZN(new_n1327_));
  NAND2_X1   g01263(.A1(new_n1327_), .A2(new_n1189_), .ZN(new_n1328_));
  INV_X1     g01264(.I(new_n1328_), .ZN(new_n1329_));
  NAND4_X1   g01265(.A1(new_n1324_), .A2(new_n1321_), .A3(new_n1326_), .A4(new_n1329_), .ZN(new_n1330_));
  OR3_X2     g01266(.A1(new_n1330_), .A2(new_n1313_), .A3(new_n1320_), .Z(new_n1331_));
  OR3_X2     g01267(.A1(new_n1299_), .A2(new_n1308_), .A3(new_n1331_), .Z(new_n1332_));
  NOR2_X1    g01268(.A1(new_n1332_), .A2(new_n1280_), .ZN(new_n1333_));
  INV_X1     g01269(.I(new_n1333_), .ZN(new_n1334_));
  INV_X1     g01270(.I(new_n152_), .ZN(new_n1335_));
  NOR2_X1    g01271(.A1(new_n491_), .A2(new_n268_), .ZN(new_n1336_));
  INV_X1     g01272(.I(new_n1336_), .ZN(new_n1337_));
  NOR2_X1    g01273(.A1(new_n482_), .A2(new_n374_), .ZN(new_n1338_));
  INV_X1     g01274(.I(new_n1338_), .ZN(new_n1339_));
  NOR2_X1    g01275(.A1(new_n136_), .A2(new_n731_), .ZN(new_n1340_));
  INV_X1     g01276(.I(new_n1340_), .ZN(new_n1341_));
  NOR3_X1    g01277(.A1(new_n1337_), .A2(new_n1339_), .A3(new_n1341_), .ZN(new_n1342_));
  NOR2_X1    g01278(.A1(new_n751_), .A2(new_n698_), .ZN(new_n1343_));
  NOR2_X1    g01279(.A1(new_n1343_), .A2(new_n294_), .ZN(new_n1344_));
  NOR2_X1    g01280(.A1(new_n170_), .A2(new_n689_), .ZN(new_n1345_));
  INV_X1     g01281(.I(new_n1345_), .ZN(new_n1346_));
  NOR3_X1    g01282(.A1(new_n1346_), .A2(new_n788_), .A3(new_n719_), .ZN(new_n1347_));
  NAND4_X1   g01283(.A1(new_n1342_), .A2(new_n1347_), .A3(new_n1226_), .A4(new_n1344_), .ZN(new_n1348_));
  NOR3_X1    g01284(.A1(new_n106_), .A2(new_n615_), .A3(new_n1167_), .ZN(new_n1349_));
  NOR3_X1    g01285(.A1(new_n396_), .A2(new_n611_), .A3(new_n397_), .ZN(new_n1350_));
  NOR3_X1    g01286(.A1(new_n267_), .A2(new_n744_), .A3(new_n154_), .ZN(new_n1351_));
  NOR3_X1    g01287(.A1(new_n602_), .A2(new_n226_), .A3(new_n804_), .ZN(new_n1352_));
  NAND4_X1   g01288(.A1(new_n1352_), .A2(new_n1351_), .A3(new_n1349_), .A4(new_n1350_), .ZN(new_n1353_));
  INV_X1     g01289(.I(new_n1076_), .ZN(new_n1354_));
  INV_X1     g01290(.I(new_n677_), .ZN(new_n1355_));
  NOR2_X1    g01291(.A1(new_n1355_), .A2(new_n596_), .ZN(new_n1356_));
  NAND3_X1   g01292(.A1(new_n1329_), .A2(new_n1356_), .A3(new_n1354_), .ZN(new_n1357_));
  NOR2_X1    g01293(.A1(new_n260_), .A2(new_n648_), .ZN(new_n1358_));
  INV_X1     g01294(.I(new_n1358_), .ZN(new_n1359_));
  NOR3_X1    g01295(.A1(new_n1359_), .A2(new_n490_), .A3(new_n867_), .ZN(new_n1360_));
  NAND3_X1   g01296(.A1(new_n1360_), .A2(new_n1165_), .A3(new_n1205_), .ZN(new_n1361_));
  NOR4_X1    g01297(.A1(new_n1348_), .A2(new_n1353_), .A3(new_n1357_), .A4(new_n1361_), .ZN(new_n1362_));
  NAND3_X1   g01298(.A1(new_n1362_), .A2(new_n1335_), .A3(new_n765_), .ZN(new_n1363_));
  INV_X1     g01299(.I(new_n1363_), .ZN(new_n1364_));
  INV_X1     g01300(.I(new_n777_), .ZN(new_n1365_));
  NOR3_X1    g01301(.A1(new_n1365_), .A2(new_n137_), .A3(new_n638_), .ZN(new_n1366_));
  NOR3_X1    g01302(.A1(new_n541_), .A2(new_n1262_), .A3(new_n498_), .ZN(new_n1367_));
  NOR4_X1    g01303(.A1(new_n70_), .A2(new_n352_), .A3(new_n437_), .A4(new_n132_), .ZN(new_n1368_));
  INV_X1     g01304(.I(new_n1368_), .ZN(new_n1369_));
  AOI22_X1   g01305(.A1(new_n180_), .A2(new_n108_), .B1(new_n185_), .B2(new_n143_), .ZN(new_n1370_));
  NOR2_X1    g01306(.A1(new_n1211_), .A2(new_n756_), .ZN(new_n1371_));
  NAND2_X1   g01307(.A1(new_n1371_), .A2(new_n1370_), .ZN(new_n1372_));
  NOR4_X1    g01308(.A1(new_n535_), .A2(new_n841_), .A3(new_n468_), .A4(new_n594_), .ZN(new_n1373_));
  INV_X1     g01309(.I(new_n1373_), .ZN(new_n1374_));
  NOR2_X1    g01310(.A1(new_n607_), .A2(new_n591_), .ZN(new_n1375_));
  NAND3_X1   g01311(.A1(new_n1374_), .A2(new_n543_), .A3(new_n1375_), .ZN(new_n1376_));
  NOR4_X1    g01312(.A1(new_n1372_), .A2(new_n210_), .A3(new_n1098_), .A4(new_n1376_), .ZN(new_n1377_));
  NAND4_X1   g01313(.A1(new_n1377_), .A2(new_n1366_), .A3(new_n1367_), .A4(new_n1369_), .ZN(new_n1378_));
  INV_X1     g01314(.I(new_n725_), .ZN(new_n1379_));
  NOR2_X1    g01315(.A1(new_n1168_), .A2(new_n625_), .ZN(new_n1380_));
  INV_X1     g01316(.I(new_n1380_), .ZN(new_n1381_));
  NAND2_X1   g01317(.A1(new_n999_), .A2(new_n349_), .ZN(new_n1382_));
  NOR4_X1    g01318(.A1(new_n1257_), .A2(new_n1379_), .A3(new_n1381_), .A4(new_n1382_), .ZN(new_n1383_));
  NOR4_X1    g01319(.A1(new_n81_), .A2(new_n252_), .A3(new_n681_), .A4(new_n286_), .ZN(new_n1384_));
  INV_X1     g01320(.I(new_n1384_), .ZN(new_n1385_));
  NAND4_X1   g01321(.A1(new_n141_), .A2(new_n1100_), .A3(new_n985_), .A4(new_n1068_), .ZN(new_n1386_));
  NOR3_X1    g01322(.A1(new_n102_), .A2(new_n488_), .A3(new_n1035_), .ZN(new_n1387_));
  NAND4_X1   g01323(.A1(new_n1383_), .A2(new_n1385_), .A3(new_n1386_), .A4(new_n1387_), .ZN(new_n1388_));
  OAI22_X1   g01324(.A1(new_n73_), .A2(new_n346_), .B1(new_n151_), .B2(new_n169_), .ZN(new_n1389_));
  INV_X1     g01325(.I(new_n1389_), .ZN(new_n1390_));
  NAND2_X1   g01326(.A1(new_n599_), .A2(new_n222_), .ZN(new_n1391_));
  NOR2_X1    g01327(.A1(new_n1391_), .A2(new_n1112_), .ZN(new_n1392_));
  NAND2_X1   g01328(.A1(new_n205_), .A2(new_n355_), .ZN(new_n1393_));
  NAND4_X1   g01329(.A1(new_n377_), .A2(new_n311_), .A3(new_n1393_), .A4(new_n669_), .ZN(new_n1394_));
  NAND2_X1   g01330(.A1(new_n270_), .A2(new_n440_), .ZN(new_n1395_));
  NAND2_X1   g01331(.A1(new_n318_), .A2(new_n196_), .ZN(new_n1396_));
  NAND4_X1   g01332(.A1(new_n434_), .A2(new_n1395_), .A3(new_n1396_), .A4(new_n880_), .ZN(new_n1397_));
  NAND4_X1   g01333(.A1(new_n1392_), .A2(new_n1390_), .A3(new_n1394_), .A4(new_n1397_), .ZN(new_n1398_));
  NOR2_X1    g01334(.A1(new_n225_), .A2(new_n173_), .ZN(new_n1399_));
  NOR4_X1    g01335(.A1(new_n548_), .A2(new_n190_), .A3(new_n654_), .A4(new_n384_), .ZN(new_n1400_));
  INV_X1     g01336(.I(new_n1400_), .ZN(new_n1401_));
  NOR3_X1    g01337(.A1(new_n367_), .A2(new_n335_), .A3(new_n506_), .ZN(new_n1402_));
  NAND2_X1   g01338(.A1(new_n318_), .A2(new_n140_), .ZN(new_n1403_));
  INV_X1     g01339(.I(new_n496_), .ZN(new_n1404_));
  NAND4_X1   g01340(.A1(new_n1404_), .A2(new_n1403_), .A3(new_n1190_), .A4(new_n423_), .ZN(new_n1405_));
  NAND4_X1   g01341(.A1(new_n1401_), .A2(new_n1399_), .A3(new_n1405_), .A4(new_n1402_), .ZN(new_n1406_));
  NOR4_X1    g01342(.A1(new_n1378_), .A2(new_n1388_), .A3(new_n1398_), .A4(new_n1406_), .ZN(new_n1407_));
  NAND2_X1   g01343(.A1(new_n1364_), .A2(new_n1407_), .ZN(new_n1408_));
  INV_X1     g01344(.I(new_n1408_), .ZN(new_n1409_));
  INV_X1     g01345(.I(new_n539_), .ZN(new_n1410_));
  NOR3_X1    g01346(.A1(new_n1410_), .A2(new_n310_), .A3(new_n930_), .ZN(new_n1411_));
  NOR2_X1    g01347(.A1(new_n734_), .A2(new_n149_), .ZN(new_n1412_));
  NAND4_X1   g01348(.A1(new_n1411_), .A2(new_n667_), .A3(new_n1281_), .A4(new_n1412_), .ZN(new_n1413_));
  NOR2_X1    g01349(.A1(new_n945_), .A2(new_n495_), .ZN(new_n1414_));
  INV_X1     g01350(.I(new_n1414_), .ZN(new_n1415_));
  NOR2_X1    g01351(.A1(new_n132_), .A2(new_n280_), .ZN(new_n1416_));
  INV_X1     g01352(.I(new_n1416_), .ZN(new_n1417_));
  NOR4_X1    g01353(.A1(new_n1415_), .A2(new_n1417_), .A3(new_n1343_), .A4(new_n1039_), .ZN(new_n1418_));
  NOR2_X1    g01354(.A1(new_n415_), .A2(new_n638_), .ZN(new_n1419_));
  INV_X1     g01355(.I(new_n1419_), .ZN(new_n1420_));
  NOR3_X1    g01356(.A1(new_n1420_), .A2(new_n125_), .A3(new_n430_), .ZN(new_n1421_));
  NAND4_X1   g01357(.A1(new_n1418_), .A2(new_n775_), .A3(new_n911_), .A4(new_n1421_), .ZN(new_n1422_));
  NOR3_X1    g01358(.A1(new_n687_), .A2(new_n634_), .A3(new_n1213_), .ZN(new_n1423_));
  NOR2_X1    g01359(.A1(new_n374_), .A2(new_n517_), .ZN(new_n1424_));
  INV_X1     g01360(.I(new_n1424_), .ZN(new_n1425_));
  NOR4_X1    g01361(.A1(new_n1425_), .A2(new_n648_), .A3(new_n486_), .A4(new_n644_), .ZN(new_n1426_));
  NAND2_X1   g01362(.A1(new_n1426_), .A2(new_n1423_), .ZN(new_n1427_));
  NOR4_X1    g01363(.A1(new_n1308_), .A2(new_n1413_), .A3(new_n1422_), .A4(new_n1427_), .ZN(new_n1428_));
  INV_X1     g01364(.I(new_n107_), .ZN(new_n1429_));
  NOR3_X1    g01365(.A1(new_n593_), .A2(new_n633_), .A3(new_n791_), .ZN(new_n1430_));
  INV_X1     g01366(.I(new_n1370_), .ZN(new_n1431_));
  NOR2_X1    g01367(.A1(new_n577_), .A2(new_n352_), .ZN(new_n1432_));
  INV_X1     g01368(.I(new_n1432_), .ZN(new_n1433_));
  NOR2_X1    g01369(.A1(new_n603_), .A2(new_n437_), .ZN(new_n1434_));
  NOR4_X1    g01370(.A1(new_n717_), .A2(new_n1433_), .A3(new_n1434_), .A4(new_n1431_), .ZN(new_n1435_));
  NAND2_X1   g01371(.A1(new_n284_), .A2(new_n196_), .ZN(new_n1436_));
  NAND3_X1   g01372(.A1(new_n690_), .A2(new_n1436_), .A3(new_n521_), .ZN(new_n1437_));
  NOR4_X1    g01373(.A1(new_n748_), .A2(new_n1437_), .A3(new_n534_), .A4(new_n456_), .ZN(new_n1438_));
  NAND3_X1   g01374(.A1(new_n1435_), .A2(new_n1438_), .A3(new_n1430_), .ZN(new_n1439_));
  INV_X1     g01375(.I(new_n569_), .ZN(new_n1440_));
  NOR2_X1    g01376(.A1(new_n753_), .A2(new_n1092_), .ZN(new_n1441_));
  NOR3_X1    g01377(.A1(new_n763_), .A2(new_n1236_), .A3(new_n741_), .ZN(new_n1442_));
  NAND4_X1   g01378(.A1(new_n1440_), .A2(new_n1156_), .A3(new_n1442_), .A4(new_n1441_), .ZN(new_n1443_));
  INV_X1     g01379(.I(new_n744_), .ZN(new_n1444_));
  NAND4_X1   g01380(.A1(new_n1444_), .A2(new_n464_), .A3(new_n871_), .A4(new_n840_), .ZN(new_n1445_));
  NAND2_X1   g01381(.A1(new_n180_), .A2(new_n186_), .ZN(new_n1446_));
  NAND4_X1   g01382(.A1(new_n1190_), .A2(new_n849_), .A3(new_n1067_), .A4(new_n1446_), .ZN(new_n1447_));
  NAND2_X1   g01383(.A1(new_n112_), .A2(new_n140_), .ZN(new_n1448_));
  NAND4_X1   g01384(.A1(new_n410_), .A2(new_n1448_), .A3(new_n606_), .A4(new_n1095_), .ZN(new_n1449_));
  NAND3_X1   g01385(.A1(new_n1445_), .A2(new_n1447_), .A3(new_n1449_), .ZN(new_n1450_));
  NOR4_X1    g01386(.A1(new_n1439_), .A2(new_n1429_), .A3(new_n1443_), .A4(new_n1450_), .ZN(new_n1451_));
  NAND2_X1   g01387(.A1(new_n1428_), .A2(new_n1451_), .ZN(new_n1452_));
  NOR2_X1    g01388(.A1(new_n1452_), .A2(new_n279_), .ZN(new_n1453_));
  NAND2_X1   g01389(.A1(new_n140_), .A2(new_n181_), .ZN(new_n1454_));
  NAND3_X1   g01390(.A1(new_n527_), .A2(new_n302_), .A3(new_n1454_), .ZN(new_n1455_));
  NOR2_X1    g01391(.A1(new_n288_), .A2(new_n587_), .ZN(new_n1456_));
  INV_X1     g01392(.I(new_n1456_), .ZN(new_n1457_));
  NOR3_X1    g01393(.A1(new_n785_), .A2(new_n1457_), .A3(new_n594_), .ZN(new_n1458_));
  NAND4_X1   g01394(.A1(new_n321_), .A2(new_n795_), .A3(new_n739_), .A4(new_n984_), .ZN(new_n1459_));
  NOR2_X1    g01395(.A1(new_n367_), .A2(new_n428_), .ZN(new_n1460_));
  INV_X1     g01396(.I(new_n1460_), .ZN(new_n1461_));
  NOR3_X1    g01397(.A1(new_n1461_), .A2(new_n615_), .A3(new_n666_), .ZN(new_n1462_));
  NOR2_X1    g01398(.A1(new_n1433_), .A2(new_n1343_), .ZN(new_n1463_));
  NAND4_X1   g01399(.A1(new_n1458_), .A2(new_n1462_), .A3(new_n1463_), .A4(new_n1459_), .ZN(new_n1464_));
  NAND2_X1   g01400(.A1(new_n355_), .A2(new_n186_), .ZN(new_n1465_));
  NAND4_X1   g01401(.A1(new_n469_), .A2(new_n773_), .A3(new_n871_), .A4(new_n1465_), .ZN(new_n1466_));
  NOR3_X1    g01402(.A1(new_n304_), .A2(new_n236_), .A3(new_n264_), .ZN(new_n1467_));
  NAND2_X1   g01403(.A1(new_n284_), .A2(new_n140_), .ZN(new_n1468_));
  NAND4_X1   g01404(.A1(new_n790_), .A2(new_n1468_), .A3(new_n856_), .A4(new_n809_), .ZN(new_n1469_));
  NAND3_X1   g01405(.A1(new_n1469_), .A2(new_n1466_), .A3(new_n1467_), .ZN(new_n1470_));
  NOR2_X1    g01406(.A1(new_n305_), .A2(new_n1175_), .ZN(new_n1471_));
  NAND2_X1   g01407(.A1(new_n690_), .A2(new_n1025_), .ZN(new_n1472_));
  NAND3_X1   g01408(.A1(new_n947_), .A2(new_n1472_), .A3(new_n1471_), .ZN(new_n1473_));
  NOR3_X1    g01409(.A1(new_n326_), .A2(new_n415_), .A3(new_n460_), .ZN(new_n1474_));
  NAND2_X1   g01410(.A1(new_n1474_), .A2(new_n439_), .ZN(new_n1475_));
  NOR4_X1    g01411(.A1(new_n1464_), .A2(new_n1470_), .A3(new_n1473_), .A4(new_n1475_), .ZN(new_n1476_));
  NOR3_X1    g01412(.A1(new_n954_), .A2(new_n1087_), .A3(new_n1185_), .ZN(new_n1477_));
  NOR3_X1    g01413(.A1(new_n117_), .A2(new_n944_), .A3(new_n286_), .ZN(new_n1478_));
  NOR3_X1    g01414(.A1(new_n1359_), .A2(new_n125_), .A3(new_n267_), .ZN(new_n1479_));
  NAND4_X1   g01415(.A1(new_n1479_), .A2(new_n1477_), .A3(new_n448_), .A4(new_n1478_), .ZN(new_n1480_));
  INV_X1     g01416(.I(new_n1480_), .ZN(new_n1481_));
  NOR4_X1    g01417(.A1(new_n424_), .A2(new_n216_), .A3(new_n430_), .A4(new_n549_), .ZN(new_n1482_));
  NOR3_X1    g01418(.A1(new_n212_), .A2(new_n198_), .A3(new_n256_), .ZN(new_n1483_));
  INV_X1     g01419(.I(new_n1483_), .ZN(new_n1484_));
  NOR4_X1    g01420(.A1(new_n1484_), .A2(new_n1482_), .A3(new_n465_), .A4(new_n634_), .ZN(new_n1485_));
  INV_X1     g01421(.I(new_n473_), .ZN(new_n1486_));
  INV_X1     g01422(.I(new_n720_), .ZN(new_n1487_));
  NOR4_X1    g01423(.A1(new_n1486_), .A2(new_n1487_), .A3(new_n1134_), .A4(new_n565_), .ZN(new_n1488_));
  NAND2_X1   g01424(.A1(new_n205_), .A2(new_n350_), .ZN(new_n1489_));
  NAND4_X1   g01425(.A1(new_n685_), .A2(new_n1489_), .A3(new_n157_), .A4(new_n246_), .ZN(new_n1490_));
  NAND2_X1   g01426(.A1(new_n109_), .A2(new_n143_), .ZN(new_n1491_));
  NAND4_X1   g01427(.A1(new_n1063_), .A2(new_n1491_), .A3(new_n985_), .A4(new_n409_), .ZN(new_n1492_));
  NOR2_X1    g01428(.A1(new_n70_), .A2(new_n154_), .ZN(new_n1493_));
  NAND2_X1   g01429(.A1(new_n140_), .A2(new_n273_), .ZN(new_n1494_));
  NAND2_X1   g01430(.A1(new_n849_), .A2(new_n1494_), .ZN(new_n1495_));
  NAND3_X1   g01431(.A1(new_n1495_), .A2(new_n336_), .A3(new_n761_), .ZN(new_n1496_));
  NOR2_X1    g01432(.A1(new_n1048_), .A2(new_n841_), .ZN(new_n1497_));
  INV_X1     g01433(.I(new_n1497_), .ZN(new_n1498_));
  NAND2_X1   g01434(.A1(new_n1189_), .A2(new_n1325_), .ZN(new_n1499_));
  NOR4_X1    g01435(.A1(new_n1498_), .A2(new_n1496_), .A3(new_n1493_), .A4(new_n1499_), .ZN(new_n1500_));
  AND4_X2    g01436(.A1(new_n1488_), .A2(new_n1500_), .A3(new_n1490_), .A4(new_n1492_), .Z(new_n1501_));
  NAND4_X1   g01437(.A1(new_n1501_), .A2(new_n1476_), .A3(new_n1481_), .A4(new_n1485_), .ZN(new_n1502_));
  NOR2_X1    g01438(.A1(new_n1455_), .A2(new_n1502_), .ZN(new_n1503_));
  INV_X1     g01439(.I(new_n1503_), .ZN(new_n1504_));
  NOR4_X1    g01440(.A1(new_n121_), .A2(new_n906_), .A3(new_n459_), .A4(new_n496_), .ZN(new_n1505_));
  NAND2_X1   g01441(.A1(new_n275_), .A2(new_n265_), .ZN(new_n1506_));
  NAND2_X1   g01442(.A1(new_n1403_), .A2(new_n1506_), .ZN(new_n1507_));
  NOR3_X1    g01443(.A1(new_n1507_), .A2(new_n307_), .A3(new_n656_), .ZN(new_n1508_));
  NOR4_X1    g01444(.A1(new_n1508_), .A2(new_n232_), .A3(new_n329_), .A4(new_n791_), .ZN(new_n1509_));
  NOR2_X1    g01445(.A1(new_n491_), .A2(new_n428_), .ZN(new_n1510_));
  INV_X1     g01446(.I(new_n1510_), .ZN(new_n1511_));
  NOR4_X1    g01447(.A1(new_n1511_), .A2(new_n1434_), .A3(new_n420_), .A4(new_n698_), .ZN(new_n1512_));
  NAND3_X1   g01448(.A1(new_n1509_), .A2(new_n1505_), .A3(new_n1512_), .ZN(new_n1513_));
  NOR2_X1    g01449(.A1(new_n1266_), .A2(new_n749_), .ZN(new_n1514_));
  NOR2_X1    g01450(.A1(new_n548_), .A2(new_n130_), .ZN(new_n1515_));
  NOR2_X1    g01451(.A1(new_n482_), .A2(new_n764_), .ZN(new_n1516_));
  NAND4_X1   g01452(.A1(new_n1514_), .A2(new_n1356_), .A3(new_n1515_), .A4(new_n1516_), .ZN(new_n1517_));
  NOR4_X1    g01453(.A1(new_n945_), .A2(new_n324_), .A3(new_n715_), .A4(new_n902_), .ZN(new_n1518_));
  NOR4_X1    g01454(.A1(new_n1518_), .A2(new_n1048_), .A3(new_n804_), .A4(new_n1262_), .ZN(new_n1519_));
  NOR3_X1    g01455(.A1(new_n515_), .A2(new_n584_), .A3(new_n684_), .ZN(new_n1520_));
  NOR3_X1    g01456(.A1(new_n573_), .A2(new_n946_), .A3(new_n255_), .ZN(new_n1521_));
  NAND3_X1   g01457(.A1(new_n1519_), .A2(new_n1520_), .A3(new_n1521_), .ZN(new_n1522_));
  NOR4_X1    g01458(.A1(new_n1513_), .A2(new_n1522_), .A3(new_n1239_), .A4(new_n1517_), .ZN(new_n1523_));
  NOR4_X1    g01459(.A1(new_n593_), .A2(new_n172_), .A3(new_n226_), .A4(new_n460_), .ZN(new_n1524_));
  NOR4_X1    g01460(.A1(new_n213_), .A2(new_n238_), .A3(new_n281_), .A4(new_n70_), .ZN(new_n1525_));
  NOR2_X1    g01461(.A1(new_n682_), .A2(new_n163_), .ZN(new_n1526_));
  INV_X1     g01462(.I(new_n1526_), .ZN(new_n1527_));
  NOR3_X1    g01463(.A1(new_n1524_), .A2(new_n1525_), .A3(new_n1527_), .ZN(new_n1528_));
  INV_X1     g01464(.I(new_n1528_), .ZN(new_n1529_));
  INV_X1     g01465(.I(new_n288_), .ZN(new_n1530_));
  NOR4_X1    g01466(.A1(new_n91_), .A2(new_n778_), .A3(new_n78_), .A4(\a[26] ), .ZN(new_n1531_));
  NOR3_X1    g01467(.A1(new_n1531_), .A2(new_n591_), .A3(new_n937_), .ZN(new_n1532_));
  NAND4_X1   g01468(.A1(new_n1532_), .A2(new_n1530_), .A3(new_n784_), .A4(new_n540_), .ZN(new_n1533_));
  NOR2_X1    g01469(.A1(new_n901_), .A2(new_n535_), .ZN(new_n1534_));
  NOR4_X1    g01470(.A1(new_n217_), .A2(new_n817_), .A3(new_n268_), .A4(new_n518_), .ZN(new_n1535_));
  INV_X1     g01471(.I(new_n1535_), .ZN(new_n1536_));
  NAND2_X1   g01472(.A1(new_n1534_), .A2(new_n1536_), .ZN(new_n1537_));
  OAI21_X1   g01473(.A1(new_n139_), .A2(new_n230_), .B(new_n109_), .ZN(new_n1538_));
  NAND2_X1   g01474(.A1(new_n377_), .A2(new_n508_), .ZN(new_n1539_));
  NOR4_X1    g01475(.A1(new_n1539_), .A2(new_n192_), .A3(new_n241_), .A4(new_n453_), .ZN(new_n1540_));
  AOI21_X1   g01476(.A1(new_n171_), .A2(new_n129_), .B(new_n151_), .ZN(new_n1541_));
  INV_X1     g01477(.I(new_n1541_), .ZN(new_n1542_));
  NAND4_X1   g01478(.A1(new_n1540_), .A2(new_n768_), .A3(new_n1538_), .A4(new_n1542_), .ZN(new_n1543_));
  NOR4_X1    g01479(.A1(new_n1537_), .A2(new_n1529_), .A3(new_n1543_), .A4(new_n1533_), .ZN(new_n1544_));
  INV_X1     g01480(.I(new_n1544_), .ZN(new_n1545_));
  NOR2_X1    g01481(.A1(new_n1545_), .A2(new_n1299_), .ZN(new_n1546_));
  NAND2_X1   g01482(.A1(new_n1546_), .A2(new_n1523_), .ZN(new_n1547_));
  NAND4_X1   g01483(.A1(new_n1444_), .A2(new_n1335_), .A3(new_n1106_), .A4(new_n669_), .ZN(new_n1548_));
  NOR2_X1    g01484(.A1(new_n633_), .A2(new_n1073_), .ZN(new_n1549_));
  NAND3_X1   g01485(.A1(new_n1549_), .A2(new_n207_), .A3(new_n871_), .ZN(new_n1550_));
  NOR2_X1    g01486(.A1(new_n496_), .A2(new_n577_), .ZN(new_n1551_));
  NAND3_X1   g01487(.A1(new_n1550_), .A2(new_n1548_), .A3(new_n1551_), .ZN(new_n1552_));
  NOR4_X1    g01488(.A1(new_n678_), .A2(new_n782_), .A3(new_n219_), .A4(new_n930_), .ZN(new_n1553_));
  NOR3_X1    g01489(.A1(new_n172_), .A2(new_n255_), .A3(new_n164_), .ZN(new_n1554_));
  NAND3_X1   g01490(.A1(new_n1553_), .A2(new_n1217_), .A3(new_n1554_), .ZN(new_n1555_));
  INV_X1     g01491(.I(new_n214_), .ZN(new_n1556_));
  NAND2_X1   g01492(.A1(new_n180_), .A2(new_n230_), .ZN(new_n1557_));
  NAND4_X1   g01493(.A1(new_n1556_), .A2(new_n436_), .A3(new_n1557_), .A4(new_n1216_), .ZN(new_n1558_));
  NAND3_X1   g01494(.A1(new_n1558_), .A2(new_n521_), .A3(new_n809_), .ZN(new_n1559_));
  NOR2_X1    g01495(.A1(new_n460_), .A2(new_n428_), .ZN(new_n1560_));
  NAND2_X1   g01496(.A1(new_n1088_), .A2(new_n319_), .ZN(new_n1561_));
  INV_X1     g01497(.I(new_n1561_), .ZN(new_n1562_));
  NAND2_X1   g01498(.A1(new_n140_), .A2(new_n270_), .ZN(new_n1563_));
  NAND2_X1   g01499(.A1(new_n292_), .A2(new_n1563_), .ZN(new_n1564_));
  INV_X1     g01500(.I(new_n1564_), .ZN(new_n1565_));
  NAND4_X1   g01501(.A1(new_n1562_), .A2(new_n1565_), .A3(new_n1265_), .A4(new_n1560_), .ZN(new_n1566_));
  NOR4_X1    g01502(.A1(new_n1555_), .A2(new_n1552_), .A3(new_n1566_), .A4(new_n1559_), .ZN(new_n1567_));
  NAND3_X1   g01503(.A1(new_n1567_), .A2(new_n690_), .A3(new_n716_), .ZN(new_n1568_));
  NAND4_X1   g01504(.A1(new_n391_), .A2(new_n849_), .A3(new_n854_), .A4(new_n522_), .ZN(new_n1569_));
  NOR2_X1    g01505(.A1(new_n505_), .A2(new_n136_), .ZN(new_n1570_));
  NAND4_X1   g01506(.A1(new_n1569_), .A2(new_n971_), .A3(new_n1570_), .A4(new_n1315_), .ZN(new_n1571_));
  NAND2_X1   g01507(.A1(new_n318_), .A2(new_n156_), .ZN(new_n1572_));
  NOR2_X1    g01508(.A1(new_n1031_), .A2(new_n485_), .ZN(new_n1573_));
  NAND4_X1   g01509(.A1(new_n1573_), .A2(new_n266_), .A3(new_n511_), .A4(new_n1572_), .ZN(new_n1574_));
  NOR2_X1    g01510(.A1(new_n251_), .A2(new_n396_), .ZN(new_n1575_));
  NOR2_X1    g01511(.A1(new_n774_), .A2(new_n910_), .ZN(new_n1576_));
  NAND4_X1   g01512(.A1(new_n1576_), .A2(new_n723_), .A3(new_n1575_), .A4(new_n768_), .ZN(new_n1577_));
  NOR2_X1    g01513(.A1(new_n463_), .A2(new_n305_), .ZN(new_n1578_));
  NOR2_X1    g01514(.A1(new_n352_), .A2(new_n724_), .ZN(new_n1579_));
  NAND4_X1   g01515(.A1(new_n1288_), .A2(new_n399_), .A3(new_n1578_), .A4(new_n1579_), .ZN(new_n1580_));
  NOR4_X1    g01516(.A1(new_n1577_), .A2(new_n1580_), .A3(new_n1571_), .A4(new_n1574_), .ZN(new_n1581_));
  NAND2_X1   g01517(.A1(new_n142_), .A2(new_n245_), .ZN(new_n1582_));
  NAND4_X1   g01518(.A1(new_n1222_), .A2(new_n1105_), .A3(new_n1582_), .A4(new_n1494_), .ZN(new_n1583_));
  NAND4_X1   g01519(.A1(new_n480_), .A2(new_n434_), .A3(new_n1468_), .A4(new_n1446_), .ZN(new_n1584_));
  NAND2_X1   g01520(.A1(new_n355_), .A2(new_n273_), .ZN(new_n1585_));
  NAND4_X1   g01521(.A1(new_n1100_), .A2(new_n1585_), .A3(new_n680_), .A4(new_n1095_), .ZN(new_n1586_));
  NAND3_X1   g01522(.A1(new_n1583_), .A2(new_n1584_), .A3(new_n1586_), .ZN(new_n1587_));
  OAI22_X1   g01523(.A1(new_n89_), .A2(new_n105_), .B1(new_n88_), .B2(new_n346_), .ZN(new_n1588_));
  NAND2_X1   g01524(.A1(new_n295_), .A2(new_n157_), .ZN(new_n1589_));
  NAND2_X1   g01525(.A1(new_n196_), .A2(new_n143_), .ZN(new_n1590_));
  NAND2_X1   g01526(.A1(new_n272_), .A2(new_n1590_), .ZN(new_n1591_));
  NOR4_X1    g01527(.A1(new_n200_), .A2(new_n1589_), .A3(new_n1591_), .A4(new_n1588_), .ZN(new_n1592_));
  NAND2_X1   g01528(.A1(new_n1592_), .A2(new_n826_), .ZN(new_n1593_));
  NOR2_X1    g01529(.A1(new_n1593_), .A2(new_n1587_), .ZN(new_n1594_));
  NAND2_X1   g01530(.A1(new_n508_), .A2(new_n978_), .ZN(new_n1595_));
  NAND4_X1   g01531(.A1(new_n160_), .A2(new_n362_), .A3(new_n551_), .A4(new_n502_), .ZN(new_n1596_));
  NAND4_X1   g01532(.A1(new_n1596_), .A2(new_n1311_), .A3(new_n1506_), .A4(new_n438_), .ZN(new_n1597_));
  NOR4_X1    g01533(.A1(new_n1597_), .A2(new_n1019_), .A3(new_n1161_), .A4(new_n1595_), .ZN(new_n1598_));
  NOR2_X1    g01534(.A1(new_n212_), .A2(new_n241_), .ZN(new_n1599_));
  NAND3_X1   g01535(.A1(new_n798_), .A2(new_n1165_), .A3(new_n1599_), .ZN(new_n1600_));
  NAND2_X1   g01536(.A1(new_n79_), .A2(new_n404_), .ZN(new_n1601_));
  NAND4_X1   g01537(.A1(new_n1066_), .A2(new_n1601_), .A3(new_n686_), .A4(new_n934_), .ZN(new_n1602_));
  NAND4_X1   g01538(.A1(new_n360_), .A2(new_n627_), .A3(new_n662_), .A4(new_n464_), .ZN(new_n1603_));
  NAND2_X1   g01539(.A1(new_n1603_), .A2(new_n1602_), .ZN(new_n1604_));
  NAND2_X1   g01540(.A1(new_n245_), .A2(new_n350_), .ZN(new_n1605_));
  NAND2_X1   g01541(.A1(new_n1192_), .A2(new_n188_), .ZN(new_n1606_));
  NAND4_X1   g01542(.A1(new_n1606_), .A2(new_n248_), .A3(new_n1605_), .A4(new_n469_), .ZN(new_n1607_));
  NOR2_X1    g01543(.A1(new_n604_), .A2(new_n749_), .ZN(new_n1608_));
  NAND4_X1   g01544(.A1(new_n1110_), .A2(new_n1126_), .A3(new_n1608_), .A4(new_n1002_), .ZN(new_n1609_));
  NOR4_X1    g01545(.A1(new_n1600_), .A2(new_n1604_), .A3(new_n1607_), .A4(new_n1609_), .ZN(new_n1610_));
  NAND4_X1   g01546(.A1(new_n1594_), .A2(new_n1581_), .A3(new_n1598_), .A4(new_n1610_), .ZN(new_n1611_));
  NOR2_X1    g01547(.A1(new_n1568_), .A2(new_n1611_), .ZN(new_n1612_));
  INV_X1     g01548(.I(new_n1612_), .ZN(new_n1613_));
  INV_X1     g01549(.I(new_n348_), .ZN(new_n1614_));
  NOR2_X1    g01550(.A1(new_n1175_), .A2(new_n298_), .ZN(new_n1615_));
  NOR4_X1    g01551(.A1(new_n1614_), .A2(new_n873_), .A3(new_n600_), .A4(new_n1615_), .ZN(new_n1616_));
  NAND4_X1   g01552(.A1(new_n197_), .A2(new_n840_), .A3(new_n436_), .A4(new_n383_), .ZN(new_n1617_));
  NAND2_X1   g01553(.A1(new_n1314_), .A2(new_n809_), .ZN(new_n1618_));
  NOR2_X1    g01554(.A1(new_n534_), .A2(new_n381_), .ZN(new_n1619_));
  NAND2_X1   g01555(.A1(new_n435_), .A2(new_n351_), .ZN(new_n1620_));
  NOR4_X1    g01556(.A1(new_n1619_), .A2(new_n1618_), .A3(new_n1620_), .A4(new_n420_), .ZN(new_n1621_));
  NAND3_X1   g01557(.A1(new_n1616_), .A2(new_n1621_), .A3(new_n1617_), .ZN(new_n1622_));
  NOR3_X1    g01558(.A1(new_n1073_), .A2(new_n518_), .A3(new_n724_), .ZN(new_n1623_));
  NAND4_X1   g01559(.A1(new_n1404_), .A2(new_n302_), .A3(new_n469_), .A4(new_n568_), .ZN(new_n1624_));
  NOR2_X1    g01560(.A1(new_n944_), .A2(new_n590_), .ZN(new_n1625_));
  NAND4_X1   g01561(.A1(new_n1624_), .A2(new_n664_), .A3(new_n1623_), .A4(new_n1625_), .ZN(new_n1626_));
  NOR2_X1    g01562(.A1(new_n582_), .A2(new_n561_), .ZN(new_n1627_));
  INV_X1     g01563(.I(new_n398_), .ZN(new_n1628_));
  NAND2_X1   g01564(.A1(new_n1628_), .A2(new_n934_), .ZN(new_n1629_));
  AOI22_X1   g01565(.A1(new_n142_), .A2(new_n181_), .B1(new_n77_), .B2(new_n273_), .ZN(new_n1630_));
  NOR4_X1    g01566(.A1(new_n1629_), .A2(new_n1247_), .A3(new_n1627_), .A4(new_n1630_), .ZN(new_n1631_));
  INV_X1     g01567(.I(new_n1599_), .ZN(new_n1632_));
  NAND2_X1   g01568(.A1(new_n1111_), .A2(new_n1321_), .ZN(new_n1633_));
  NOR4_X1    g01569(.A1(new_n1633_), .A2(new_n192_), .A3(new_n1152_), .A4(new_n1632_), .ZN(new_n1634_));
  NAND4_X1   g01570(.A1(new_n353_), .A2(new_n393_), .A3(new_n739_), .A4(new_n222_), .ZN(new_n1635_));
  NAND4_X1   g01571(.A1(new_n1634_), .A2(new_n884_), .A3(new_n1631_), .A4(new_n1635_), .ZN(new_n1636_));
  OR3_X2     g01572(.A1(new_n1636_), .A2(new_n1622_), .A3(new_n1626_), .Z(new_n1637_));
  NAND2_X1   g01573(.A1(new_n108_), .A2(new_n350_), .ZN(new_n1638_));
  NAND4_X1   g01574(.A1(new_n480_), .A2(new_n479_), .A3(new_n1638_), .A4(new_n665_), .ZN(new_n1639_));
  NAND3_X1   g01575(.A1(new_n823_), .A2(new_n606_), .A3(new_n409_), .ZN(new_n1640_));
  NOR3_X1    g01576(.A1(new_n1640_), .A2(new_n268_), .A3(new_n796_), .ZN(new_n1641_));
  NAND2_X1   g01577(.A1(new_n1641_), .A2(new_n1639_), .ZN(new_n1642_));
  NAND3_X1   g01578(.A1(new_n1129_), .A2(new_n1572_), .A3(new_n362_), .ZN(new_n1643_));
  INV_X1     g01579(.I(new_n1643_), .ZN(new_n1644_));
  NOR4_X1    g01580(.A1(new_n255_), .A2(new_n312_), .A3(new_n610_), .A4(new_n474_), .ZN(new_n1645_));
  NAND2_X1   g01581(.A1(new_n318_), .A2(new_n180_), .ZN(new_n1646_));
  NAND2_X1   g01582(.A1(new_n230_), .A2(new_n350_), .ZN(new_n1647_));
  NAND3_X1   g01583(.A1(new_n1646_), .A2(new_n843_), .A3(new_n1647_), .ZN(new_n1648_));
  NOR2_X1    g01584(.A1(new_n1645_), .A2(new_n1648_), .ZN(new_n1649_));
  NOR3_X1    g01585(.A1(new_n914_), .A2(new_n772_), .A3(new_n666_), .ZN(new_n1650_));
  NOR4_X1    g01586(.A1(new_n1650_), .A2(new_n247_), .A3(new_n304_), .A4(new_n801_), .ZN(new_n1651_));
  NAND2_X1   g01587(.A1(new_n1530_), .A2(new_n1058_), .ZN(new_n1652_));
  NOR4_X1    g01588(.A1(new_n1359_), .A2(new_n1652_), .A3(new_n114_), .A4(new_n316_), .ZN(new_n1653_));
  NAND4_X1   g01589(.A1(new_n1651_), .A2(new_n1644_), .A3(new_n1649_), .A4(new_n1653_), .ZN(new_n1654_));
  NOR2_X1    g01590(.A1(new_n1654_), .A2(new_n1642_), .ZN(new_n1655_));
  NAND2_X1   g01591(.A1(new_n287_), .A2(new_n980_), .ZN(new_n1656_));
  NOR4_X1    g01592(.A1(new_n1656_), .A2(new_n214_), .A3(new_n456_), .A4(new_n867_), .ZN(new_n1657_));
  INV_X1     g01593(.I(new_n106_), .ZN(new_n1658_));
  NAND3_X1   g01594(.A1(new_n1658_), .A2(new_n1105_), .A3(new_n184_), .ZN(new_n1659_));
  NOR4_X1    g01595(.A1(new_n1659_), .A2(new_n397_), .A3(new_n517_), .A4(new_n1076_), .ZN(new_n1660_));
  NAND3_X1   g01596(.A1(new_n1660_), .A2(new_n1657_), .A3(new_n1423_), .ZN(new_n1661_));
  NAND2_X1   g01597(.A1(new_n284_), .A2(new_n109_), .ZN(new_n1662_));
  NAND3_X1   g01598(.A1(new_n208_), .A2(new_n1662_), .A3(new_n414_), .ZN(new_n1663_));
  NAND2_X1   g01599(.A1(new_n572_), .A2(new_n985_), .ZN(new_n1664_));
  NOR4_X1    g01600(.A1(new_n1663_), .A2(new_n1664_), .A3(new_n329_), .A4(new_n644_), .ZN(new_n1665_));
  NAND2_X1   g01601(.A1(new_n440_), .A2(new_n186_), .ZN(new_n1666_));
  NAND3_X1   g01602(.A1(new_n322_), .A2(new_n1396_), .A3(new_n1666_), .ZN(new_n1667_));
  NOR3_X1    g01603(.A1(new_n135_), .A2(new_n320_), .A3(new_n125_), .ZN(new_n1668_));
  INV_X1     g01604(.I(new_n1668_), .ZN(new_n1669_));
  NOR2_X1    g01605(.A1(new_n1669_), .A2(new_n1667_), .ZN(new_n1670_));
  OAI22_X1   g01606(.A1(new_n334_), .A2(new_n75_), .B1(new_n123_), .B2(new_n148_), .ZN(new_n1671_));
  NAND2_X1   g01607(.A1(new_n1671_), .A2(new_n983_), .ZN(new_n1672_));
  NOR3_X1    g01608(.A1(new_n1672_), .A2(new_n251_), .A3(new_n1434_), .ZN(new_n1673_));
  NOR3_X1    g01609(.A1(new_n713_), .A2(new_n523_), .A3(new_n1541_), .ZN(new_n1674_));
  NAND4_X1   g01610(.A1(new_n1670_), .A2(new_n1665_), .A3(new_n1673_), .A4(new_n1674_), .ZN(new_n1675_));
  NOR2_X1    g01611(.A1(new_n1661_), .A2(new_n1675_), .ZN(new_n1676_));
  NAND2_X1   g01612(.A1(new_n1655_), .A2(new_n1676_), .ZN(new_n1677_));
  NOR2_X1    g01613(.A1(new_n1677_), .A2(new_n1637_), .ZN(new_n1678_));
  OAI22_X1   g01614(.A1(new_n75_), .A2(new_n105_), .B1(new_n97_), .B2(new_n85_), .ZN(new_n1679_));
  NAND4_X1   g01615(.A1(new_n1679_), .A2(new_n624_), .A3(new_n141_), .A4(new_n1494_), .ZN(new_n1680_));
  NOR4_X1    g01616(.A1(new_n783_), .A2(new_n867_), .A3(new_n574_), .A4(new_n280_), .ZN(new_n1681_));
  NOR4_X1    g01617(.A1(new_n1680_), .A2(new_n1667_), .A3(new_n1681_), .A4(new_n1250_), .ZN(new_n1682_));
  NOR4_X1    g01618(.A1(new_n135_), .A2(new_n591_), .A3(new_n202_), .A4(new_n937_), .ZN(new_n1683_));
  NOR4_X1    g01619(.A1(new_n453_), .A2(new_n779_), .A3(new_n553_), .A4(new_n330_), .ZN(new_n1684_));
  NOR4_X1    g01620(.A1(new_n906_), .A2(new_n86_), .A3(new_n535_), .A4(new_n732_), .ZN(new_n1685_));
  NOR3_X1    g01621(.A1(new_n1683_), .A2(new_n1685_), .A3(new_n1684_), .ZN(new_n1686_));
  NOR3_X1    g01622(.A1(new_n702_), .A2(new_n1078_), .A3(new_n1079_), .ZN(new_n1687_));
  NAND4_X1   g01623(.A1(new_n1682_), .A2(new_n1686_), .A3(new_n1324_), .A4(new_n1687_), .ZN(new_n1688_));
  OAI21_X1   g01624(.A1(new_n270_), .A2(new_n139_), .B(new_n185_), .ZN(new_n1689_));
  OAI22_X1   g01625(.A1(new_n101_), .A2(new_n169_), .B1(new_n88_), .B2(new_n150_), .ZN(new_n1690_));
  NAND2_X1   g01626(.A1(new_n1690_), .A2(new_n1689_), .ZN(new_n1691_));
  OAI22_X1   g01627(.A1(new_n66_), .A2(new_n97_), .B1(new_n75_), .B2(new_n153_), .ZN(new_n1692_));
  NAND3_X1   g01628(.A1(new_n1692_), .A2(new_n378_), .A3(new_n880_), .ZN(new_n1693_));
  NOR4_X1    g01629(.A1(new_n652_), .A2(new_n1152_), .A3(new_n419_), .A4(new_n594_), .ZN(new_n1694_));
  OAI21_X1   g01630(.A1(new_n1531_), .A2(new_n944_), .B(new_n1491_), .ZN(new_n1695_));
  NOR4_X1    g01631(.A1(new_n1691_), .A2(new_n1693_), .A3(new_n1694_), .A4(new_n1695_), .ZN(new_n1696_));
  OAI22_X1   g01632(.A1(new_n69_), .A2(new_n105_), .B1(new_n148_), .B2(new_n346_), .ZN(new_n1697_));
  NAND4_X1   g01633(.A1(new_n1697_), .A2(new_n1538_), .A3(new_n250_), .A4(new_n1605_), .ZN(new_n1698_));
  OAI21_X1   g01634(.A1(new_n186_), .A2(new_n181_), .B(new_n196_), .ZN(new_n1699_));
  OAI21_X1   g01635(.A1(new_n205_), .A2(new_n245_), .B(new_n140_), .ZN(new_n1700_));
  OAI21_X1   g01636(.A1(new_n156_), .A2(new_n350_), .B(new_n273_), .ZN(new_n1701_));
  NAND4_X1   g01637(.A1(new_n537_), .A2(new_n1699_), .A3(new_n1700_), .A4(new_n1701_), .ZN(new_n1702_));
  NOR2_X1    g01638(.A1(new_n1702_), .A2(new_n1698_), .ZN(new_n1703_));
  NOR4_X1    g01639(.A1(new_n90_), .A2(new_n192_), .A3(new_n388_), .A4(new_n490_), .ZN(new_n1704_));
  NOR4_X1    g01640(.A1(new_n203_), .A2(new_n304_), .A3(new_n582_), .A4(new_n324_), .ZN(new_n1705_));
  NAND2_X1   g01641(.A1(new_n159_), .A2(new_n265_), .ZN(new_n1706_));
  NAND3_X1   g01642(.A1(new_n1403_), .A2(new_n1706_), .A3(new_n643_), .ZN(new_n1707_));
  NOR3_X1    g01643(.A1(new_n1705_), .A2(new_n1704_), .A3(new_n1707_), .ZN(new_n1708_));
  NAND4_X1   g01644(.A1(new_n1696_), .A2(new_n1703_), .A3(new_n1708_), .A4(new_n1182_), .ZN(new_n1709_));
  INV_X1     g01645(.I(new_n1554_), .ZN(new_n1710_));
  OAI22_X1   g01646(.A1(new_n118_), .A2(new_n129_), .B1(new_n131_), .B2(new_n151_), .ZN(new_n1711_));
  AOI22_X1   g01647(.A1(new_n79_), .A2(new_n206_), .B1(new_n318_), .B2(new_n350_), .ZN(new_n1712_));
  NAND4_X1   g01648(.A1(new_n1712_), .A2(new_n1711_), .A3(new_n373_), .A4(new_n564_), .ZN(new_n1713_));
  NAND3_X1   g01649(.A1(new_n113_), .A2(new_n1489_), .A3(new_n934_), .ZN(new_n1714_));
  NOR4_X1    g01650(.A1(new_n170_), .A2(new_n370_), .A3(new_n721_), .A4(new_n715_), .ZN(new_n1715_));
  NOR4_X1    g01651(.A1(new_n1710_), .A2(new_n1713_), .A3(new_n1714_), .A4(new_n1715_), .ZN(new_n1716_));
  NOR4_X1    g01652(.A1(new_n173_), .A2(new_n92_), .A3(new_n736_), .A4(new_n724_), .ZN(new_n1717_));
  NOR4_X1    g01653(.A1(new_n102_), .A2(new_n98_), .A3(new_n396_), .A4(new_n625_), .ZN(new_n1718_));
  NAND2_X1   g01654(.A1(new_n265_), .A2(new_n206_), .ZN(new_n1719_));
  NAND2_X1   g01655(.A1(new_n1646_), .A2(new_n1719_), .ZN(new_n1720_));
  NOR4_X1    g01656(.A1(new_n1718_), .A2(new_n347_), .A3(new_n1717_), .A4(new_n1720_), .ZN(new_n1721_));
  NAND3_X1   g01657(.A1(new_n1471_), .A2(new_n1516_), .A3(new_n1370_), .ZN(new_n1722_));
  NOR4_X1    g01658(.A1(new_n147_), .A2(new_n154_), .A3(new_n634_), .A4(new_n556_), .ZN(new_n1723_));
  NOR4_X1    g01659(.A1(new_n227_), .A2(new_n463_), .A3(new_n262_), .A4(new_n449_), .ZN(new_n1724_));
  NAND2_X1   g01660(.A1(new_n275_), .A2(new_n158_), .ZN(new_n1725_));
  NAND4_X1   g01661(.A1(new_n160_), .A2(new_n1601_), .A3(new_n1725_), .A4(new_n872_), .ZN(new_n1726_));
  NOR4_X1    g01662(.A1(new_n1722_), .A2(new_n1723_), .A3(new_n1724_), .A4(new_n1726_), .ZN(new_n1727_));
  NAND3_X1   g01663(.A1(new_n1727_), .A2(new_n1716_), .A3(new_n1721_), .ZN(new_n1728_));
  NOR3_X1    g01664(.A1(new_n1728_), .A2(new_n1688_), .A3(new_n1709_), .ZN(new_n1729_));
  NAND2_X1   g01665(.A1(new_n80_), .A2(new_n1063_), .ZN(new_n1730_));
  NOR4_X1    g01666(.A1(new_n552_), .A2(new_n850_), .A3(new_n1499_), .A4(new_n1730_), .ZN(new_n1731_));
  NAND3_X1   g01667(.A1(new_n138_), .A2(new_n790_), .A3(new_n1454_), .ZN(new_n1732_));
  NAND2_X1   g01668(.A1(new_n1358_), .A2(new_n1237_), .ZN(new_n1733_));
  NOR4_X1    g01669(.A1(new_n549_), .A2(new_n256_), .A3(new_n388_), .A4(new_n731_), .ZN(new_n1734_));
  NOR4_X1    g01670(.A1(new_n644_), .A2(new_n264_), .A3(new_n320_), .A4(new_n376_), .ZN(new_n1735_));
  NOR4_X1    g01671(.A1(new_n1733_), .A2(new_n1732_), .A3(new_n1735_), .A4(new_n1734_), .ZN(new_n1736_));
  NAND2_X1   g01672(.A1(new_n1736_), .A2(new_n1731_), .ZN(new_n1737_));
  NOR4_X1    g01673(.A1(new_n569_), .A2(new_n170_), .A3(new_n465_), .A4(new_n437_), .ZN(new_n1738_));
  NOR4_X1    g01674(.A1(new_n135_), .A2(new_n615_), .A3(new_n610_), .A4(new_n306_), .ZN(new_n1739_));
  NOR4_X1    g01675(.A1(new_n1739_), .A2(new_n238_), .A3(new_n638_), .A4(new_n796_), .ZN(new_n1740_));
  NOR4_X1    g01676(.A1(new_n183_), .A2(new_n420_), .A3(new_n488_), .A4(new_n682_), .ZN(new_n1741_));
  NOR4_X1    g01677(.A1(new_n1741_), .A2(new_n247_), .A3(new_n560_), .A4(new_n783_), .ZN(new_n1742_));
  NAND3_X1   g01678(.A1(new_n1742_), .A2(new_n1740_), .A3(new_n1738_), .ZN(new_n1743_));
  NOR3_X1    g01679(.A1(new_n299_), .A2(new_n637_), .A3(new_n282_), .ZN(new_n1744_));
  OAI21_X1   g01680(.A1(new_n139_), .A2(new_n230_), .B(new_n350_), .ZN(new_n1745_));
  NOR4_X1    g01681(.A1(new_n510_), .A2(new_n611_), .A3(new_n684_), .A4(new_n718_), .ZN(new_n1746_));
  NOR4_X1    g01682(.A1(new_n1746_), .A2(new_n468_), .A3(new_n475_), .A4(new_n910_), .ZN(new_n1747_));
  NAND4_X1   g01683(.A1(new_n1747_), .A2(new_n545_), .A3(new_n1744_), .A4(new_n1745_), .ZN(new_n1748_));
  NOR4_X1    g01684(.A1(new_n1737_), .A2(new_n847_), .A3(new_n1748_), .A4(new_n1743_), .ZN(new_n1749_));
  NAND3_X1   g01685(.A1(new_n1010_), .A2(new_n823_), .A3(new_n672_), .ZN(new_n1750_));
  NOR2_X1    g01686(.A1(new_n604_), .A2(new_n190_), .ZN(new_n1751_));
  NAND3_X1   g01687(.A1(new_n722_), .A2(new_n1751_), .A3(new_n348_), .ZN(new_n1752_));
  INV_X1     g01688(.I(new_n374_), .ZN(new_n1753_));
  NAND2_X1   g01689(.A1(new_n1753_), .A2(new_n1646_), .ZN(new_n1754_));
  NAND2_X1   g01690(.A1(new_n1065_), .A2(new_n302_), .ZN(new_n1755_));
  NOR2_X1    g01691(.A1(new_n1754_), .A2(new_n1755_), .ZN(new_n1756_));
  NAND3_X1   g01692(.A1(new_n1756_), .A2(new_n507_), .A3(new_n1156_), .ZN(new_n1757_));
  NAND4_X1   g01693(.A1(new_n221_), .A2(new_n1105_), .A3(new_n1706_), .A4(new_n1465_), .ZN(new_n1758_));
  NAND2_X1   g01694(.A1(new_n196_), .A2(new_n270_), .ZN(new_n1759_));
  NAND4_X1   g01695(.A1(new_n295_), .A2(new_n405_), .A3(new_n854_), .A4(new_n1759_), .ZN(new_n1760_));
  NAND2_X1   g01696(.A1(new_n1760_), .A2(new_n1758_), .ZN(new_n1761_));
  NOR4_X1    g01697(.A1(new_n1750_), .A2(new_n1752_), .A3(new_n1757_), .A4(new_n1761_), .ZN(new_n1762_));
  NAND3_X1   g01698(.A1(new_n1749_), .A2(new_n1567_), .A3(new_n1762_), .ZN(new_n1763_));
  INV_X1     g01699(.I(new_n1763_), .ZN(new_n1764_));
  NOR2_X1    g01700(.A1(new_n281_), .A2(new_n490_), .ZN(new_n1765_));
  NOR2_X1    g01701(.A1(new_n1355_), .A2(new_n261_), .ZN(new_n1766_));
  NAND2_X1   g01702(.A1(new_n1068_), .A2(new_n627_), .ZN(new_n1767_));
  NAND4_X1   g01703(.A1(new_n1766_), .A2(new_n537_), .A3(new_n1765_), .A4(new_n1767_), .ZN(new_n1768_));
  NAND3_X1   g01704(.A1(new_n761_), .A2(new_n405_), .A3(new_n414_), .ZN(new_n1769_));
  OAI21_X1   g01705(.A1(new_n112_), .A2(new_n186_), .B(new_n440_), .ZN(new_n1770_));
  NAND3_X1   g01706(.A1(new_n1770_), .A2(new_n322_), .A3(new_n598_), .ZN(new_n1771_));
  NAND3_X1   g01707(.A1(new_n773_), .A2(new_n293_), .A3(new_n1662_), .ZN(new_n1772_));
  OR4_X2     g01708(.A1(new_n1373_), .A2(new_n1771_), .A3(new_n1772_), .A4(new_n1769_), .Z(new_n1773_));
  NAND3_X1   g01709(.A1(new_n795_), .A2(new_n872_), .A3(new_n1322_), .ZN(new_n1774_));
  NAND4_X1   g01710(.A1(new_n819_), .A2(new_n643_), .A3(new_n1325_), .A4(new_n809_), .ZN(new_n1775_));
  NOR2_X1    g01711(.A1(new_n1775_), .A2(new_n1774_), .ZN(new_n1776_));
  INV_X1     g01712(.I(new_n1776_), .ZN(new_n1777_));
  NOR4_X1    g01713(.A1(new_n1773_), .A2(new_n1642_), .A3(new_n1777_), .A4(new_n1768_), .ZN(new_n1778_));
  AOI21_X1   g01714(.A1(new_n101_), .A2(new_n115_), .B(new_n123_), .ZN(new_n1779_));
  AOI21_X1   g01715(.A1(new_n95_), .A2(new_n153_), .B(new_n123_), .ZN(new_n1780_));
  NOR4_X1    g01716(.A1(new_n1779_), .A2(new_n92_), .A3(new_n1780_), .A4(new_n453_), .ZN(new_n1781_));
  NOR2_X1    g01717(.A1(new_n125_), .A2(new_n937_), .ZN(new_n1782_));
  NOR4_X1    g01718(.A1(new_n712_), .A2(new_n1782_), .A3(new_n618_), .A4(new_n1185_), .ZN(new_n1783_));
  NOR2_X1    g01719(.A1(new_n698_), .A2(new_n510_), .ZN(new_n1784_));
  NOR4_X1    g01720(.A1(new_n1784_), .A2(new_n241_), .A3(new_n734_), .A4(new_n763_), .ZN(new_n1785_));
  NAND4_X1   g01721(.A1(new_n1673_), .A2(new_n1783_), .A3(new_n1785_), .A4(new_n1781_), .ZN(new_n1786_));
  NOR2_X1    g01722(.A1(new_n637_), .A2(new_n124_), .ZN(new_n1787_));
  NOR2_X1    g01723(.A1(new_n590_), .A2(new_n1168_), .ZN(new_n1788_));
  OAI22_X1   g01724(.A1(new_n534_), .A2(new_n381_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n1789_));
  NOR3_X1    g01725(.A1(new_n1789_), .A2(new_n1787_), .A3(new_n1788_), .ZN(new_n1790_));
  NOR4_X1    g01726(.A1(new_n211_), .A2(new_n398_), .A3(new_n531_), .A4(new_n640_), .ZN(new_n1791_));
  NOR4_X1    g01727(.A1(new_n226_), .A2(new_n374_), .A3(new_n163_), .A4(new_n329_), .ZN(new_n1792_));
  NOR2_X1    g01728(.A1(new_n1791_), .A2(new_n1792_), .ZN(new_n1793_));
  NOR4_X1    g01729(.A1(new_n403_), .A2(new_n652_), .A3(new_n306_), .A4(new_n430_), .ZN(new_n1794_));
  NOR4_X1    g01730(.A1(new_n213_), .A2(new_n498_), .A3(new_n136_), .A4(new_n152_), .ZN(new_n1795_));
  NAND2_X1   g01731(.A1(new_n318_), .A2(new_n440_), .ZN(new_n1796_));
  NAND3_X1   g01732(.A1(new_n80_), .A2(new_n351_), .A3(new_n1796_), .ZN(new_n1797_));
  NOR3_X1    g01733(.A1(new_n1794_), .A2(new_n1795_), .A3(new_n1797_), .ZN(new_n1798_));
  NAND3_X1   g01734(.A1(new_n1790_), .A2(new_n1798_), .A3(new_n1793_), .ZN(new_n1799_));
  NOR2_X1    g01735(.A1(new_n1799_), .A2(new_n1786_), .ZN(new_n1800_));
  NOR3_X1    g01736(.A1(new_n788_), .A2(new_n242_), .A3(new_n280_), .ZN(new_n1801_));
  NOR2_X1    g01737(.A1(new_n333_), .A2(new_n475_), .ZN(new_n1802_));
  NOR2_X1    g01738(.A1(new_n1802_), .A2(new_n1054_), .ZN(new_n1803_));
  NOR3_X1    g01739(.A1(new_n604_), .A2(new_n731_), .A3(new_n764_), .ZN(new_n1804_));
  NAND2_X1   g01740(.A1(new_n180_), .A2(new_n139_), .ZN(new_n1805_));
  NAND4_X1   g01741(.A1(new_n1805_), .A2(new_n1327_), .A3(new_n672_), .A4(new_n1095_), .ZN(new_n1806_));
  NAND4_X1   g01742(.A1(new_n1803_), .A2(new_n1801_), .A3(new_n1806_), .A4(new_n1804_), .ZN(new_n1807_));
  AOI21_X1   g01743(.A1(new_n122_), .A2(new_n151_), .B(new_n69_), .ZN(new_n1808_));
  NOR4_X1    g01744(.A1(new_n1808_), .A2(new_n944_), .A3(new_n491_), .A4(new_n560_), .ZN(new_n1809_));
  NOR2_X1    g01745(.A1(new_n147_), .A2(new_n783_), .ZN(new_n1810_));
  NAND4_X1   g01746(.A1(new_n1809_), .A2(new_n1199_), .A3(new_n1810_), .A4(new_n1745_), .ZN(new_n1811_));
  NOR3_X1    g01747(.A1(new_n1398_), .A2(new_n1807_), .A3(new_n1811_), .ZN(new_n1812_));
  NAND3_X1   g01748(.A1(new_n1800_), .A2(new_n1778_), .A3(new_n1812_), .ZN(new_n1813_));
  NOR2_X1    g01749(.A1(new_n465_), .A2(new_n899_), .ZN(new_n1814_));
  NAND3_X1   g01750(.A1(new_n1814_), .A2(new_n761_), .A3(new_n757_), .ZN(new_n1815_));
  INV_X1     g01751(.I(new_n298_), .ZN(new_n1816_));
  NAND2_X1   g01752(.A1(new_n1816_), .A2(new_n207_), .ZN(new_n1817_));
  NAND2_X1   g01753(.A1(new_n1454_), .A2(new_n356_), .ZN(new_n1818_));
  NAND2_X1   g01754(.A1(new_n662_), .A2(new_n856_), .ZN(new_n1819_));
  NAND4_X1   g01755(.A1(new_n1472_), .A2(new_n1817_), .A3(new_n1819_), .A4(new_n1818_), .ZN(new_n1820_));
  NOR4_X1    g01756(.A1(new_n238_), .A2(new_n387_), .A3(new_n320_), .A4(new_n625_), .ZN(new_n1821_));
  NAND3_X1   g01757(.A1(new_n871_), .A2(new_n655_), .A3(new_n809_), .ZN(new_n1822_));
  NOR4_X1    g01758(.A1(new_n1820_), .A2(new_n1815_), .A3(new_n1821_), .A4(new_n1822_), .ZN(new_n1823_));
  NAND4_X1   g01759(.A1(new_n1314_), .A2(new_n1563_), .A3(new_n309_), .A4(new_n390_), .ZN(new_n1824_));
  OAI22_X1   g01760(.A1(new_n129_), .A2(new_n118_), .B1(new_n171_), .B2(new_n122_), .ZN(new_n1825_));
  NOR2_X1    g01761(.A1(new_n837_), .A2(new_n474_), .ZN(new_n1826_));
  NAND4_X1   g01762(.A1(new_n1824_), .A2(new_n729_), .A3(new_n1825_), .A4(new_n1826_), .ZN(new_n1827_));
  NOR3_X1    g01763(.A1(new_n485_), .A2(new_n456_), .A3(new_n125_), .ZN(new_n1828_));
  NAND2_X1   g01764(.A1(new_n205_), .A2(new_n159_), .ZN(new_n1829_));
  NAND4_X1   g01765(.A1(new_n1829_), .A2(new_n572_), .A3(new_n435_), .A4(new_n157_), .ZN(new_n1830_));
  NAND2_X1   g01766(.A1(new_n275_), .A2(new_n273_), .ZN(new_n1831_));
  NAND2_X1   g01767(.A1(new_n158_), .A2(new_n142_), .ZN(new_n1832_));
  NAND4_X1   g01768(.A1(new_n1831_), .A2(new_n1832_), .A3(new_n1468_), .A4(new_n849_), .ZN(new_n1833_));
  NAND3_X1   g01769(.A1(new_n1833_), .A2(new_n1830_), .A3(new_n1828_), .ZN(new_n1834_));
  INV_X1     g01770(.I(new_n1147_), .ZN(new_n1835_));
  NAND2_X1   g01771(.A1(new_n1436_), .A2(new_n823_), .ZN(new_n1836_));
  NAND3_X1   g01772(.A1(new_n1835_), .A2(new_n1767_), .A3(new_n1836_), .ZN(new_n1837_));
  NAND2_X1   g01773(.A1(new_n181_), .A2(new_n350_), .ZN(new_n1838_));
  NOR2_X1    g01774(.A1(new_n76_), .A2(new_n136_), .ZN(new_n1839_));
  NOR2_X1    g01775(.A1(new_n587_), .A2(new_n306_), .ZN(new_n1840_));
  NAND4_X1   g01776(.A1(new_n1839_), .A2(new_n1840_), .A3(new_n1110_), .A4(new_n1838_), .ZN(new_n1841_));
  NOR4_X1    g01777(.A1(new_n1827_), .A2(new_n1837_), .A3(new_n1834_), .A4(new_n1841_), .ZN(new_n1842_));
  NOR2_X1    g01778(.A1(new_n460_), .A2(new_n584_), .ZN(new_n1843_));
  NOR3_X1    g01779(.A1(new_n670_), .A2(new_n191_), .A3(new_n1092_), .ZN(new_n1844_));
  NOR4_X1    g01780(.A1(new_n1630_), .A2(new_n782_), .A3(new_n548_), .A4(new_n801_), .ZN(new_n1845_));
  NAND4_X1   g01781(.A1(new_n1845_), .A2(new_n1173_), .A3(new_n1843_), .A4(new_n1844_), .ZN(new_n1846_));
  NAND4_X1   g01782(.A1(new_n1305_), .A2(new_n1091_), .A3(new_n854_), .A4(new_n432_), .ZN(new_n1847_));
  NOR3_X1    g01783(.A1(new_n553_), .A2(new_n791_), .A3(new_n535_), .ZN(new_n1848_));
  NAND4_X1   g01784(.A1(new_n1847_), .A2(new_n592_), .A3(new_n1848_), .A4(new_n1059_), .ZN(new_n1849_));
  NOR3_X1    g01785(.A1(new_n170_), .A2(new_n772_), .A3(new_n741_), .ZN(new_n1850_));
  NOR3_X1    g01786(.A1(new_n177_), .A2(new_n447_), .A3(new_n1236_), .ZN(new_n1851_));
  NAND4_X1   g01787(.A1(new_n271_), .A2(new_n451_), .A3(new_n272_), .A4(new_n302_), .ZN(new_n1852_));
  NAND2_X1   g01788(.A1(new_n230_), .A2(new_n185_), .ZN(new_n1853_));
  NAND4_X1   g01789(.A1(new_n808_), .A2(new_n701_), .A3(new_n1853_), .A4(new_n1590_), .ZN(new_n1854_));
  NAND4_X1   g01790(.A1(new_n1851_), .A2(new_n1852_), .A3(new_n1854_), .A4(new_n1850_), .ZN(new_n1855_));
  OAI22_X1   g01791(.A1(new_n134_), .A2(new_n148_), .B1(new_n150_), .B2(new_n153_), .ZN(new_n1856_));
  NOR3_X1    g01792(.A1(new_n906_), .A2(new_n695_), .A3(new_n719_), .ZN(new_n1857_));
  AOI21_X1   g01793(.A1(new_n133_), .A2(new_n118_), .B(new_n97_), .ZN(new_n1858_));
  NOR2_X1    g01794(.A1(new_n544_), .A2(new_n1858_), .ZN(new_n1859_));
  NAND4_X1   g01795(.A1(new_n1859_), .A2(new_n1857_), .A3(new_n516_), .A4(new_n1856_), .ZN(new_n1860_));
  NOR4_X1    g01796(.A1(new_n1846_), .A2(new_n1855_), .A3(new_n1849_), .A4(new_n1860_), .ZN(new_n1861_));
  NAND4_X1   g01797(.A1(new_n1861_), .A2(new_n1812_), .A3(new_n1842_), .A4(new_n1823_), .ZN(new_n1862_));
  NAND2_X1   g01798(.A1(new_n1862_), .A2(new_n1729_), .ZN(new_n1863_));
  AOI22_X1   g01799(.A1(new_n140_), .A2(new_n158_), .B1(new_n111_), .B2(new_n186_), .ZN(new_n1864_));
  OAI22_X1   g01800(.A1(new_n88_), .A2(new_n171_), .B1(new_n134_), .B2(new_n122_), .ZN(new_n1865_));
  OAI22_X1   g01801(.A1(new_n171_), .A2(new_n115_), .B1(new_n105_), .B2(new_n123_), .ZN(new_n1866_));
  NOR3_X1    g01802(.A1(new_n1864_), .A2(new_n1865_), .A3(new_n1866_), .ZN(new_n1867_));
  NOR3_X1    g01803(.A1(new_n149_), .A2(new_n239_), .A3(new_n782_), .ZN(new_n1868_));
  NAND4_X1   g01804(.A1(new_n393_), .A2(new_n808_), .A3(new_n1796_), .A4(new_n1662_), .ZN(new_n1869_));
  NAND4_X1   g01805(.A1(new_n1867_), .A2(new_n1554_), .A3(new_n1869_), .A4(new_n1868_), .ZN(new_n1870_));
  NAND4_X1   g01806(.A1(new_n675_), .A2(new_n795_), .A3(new_n840_), .A4(new_n301_), .ZN(new_n1871_));
  NAND4_X1   g01807(.A1(new_n441_), .A2(new_n978_), .A3(new_n182_), .A4(new_n761_), .ZN(new_n1872_));
  NOR2_X1    g01808(.A1(new_n1720_), .A2(new_n347_), .ZN(new_n1873_));
  NAND3_X1   g01809(.A1(new_n1873_), .A2(new_n1871_), .A3(new_n1872_), .ZN(new_n1874_));
  OAI22_X1   g01810(.A1(new_n148_), .A2(new_n171_), .B1(new_n83_), .B2(new_n133_), .ZN(new_n1875_));
  NOR4_X1    g01811(.A1(new_n1875_), .A2(new_n1588_), .A3(new_n770_), .A4(new_n381_), .ZN(new_n1876_));
  NAND4_X1   g01812(.A1(new_n628_), .A2(new_n1216_), .A3(new_n1327_), .A4(new_n1009_), .ZN(new_n1877_));
  NAND4_X1   g01813(.A1(new_n599_), .A2(new_n434_), .A3(new_n276_), .A4(new_n274_), .ZN(new_n1878_));
  NOR4_X1    g01814(.A1(new_n413_), .A2(new_n587_), .A3(new_n718_), .A4(new_n776_), .ZN(new_n1879_));
  NAND4_X1   g01815(.A1(new_n1876_), .A2(new_n1877_), .A3(new_n1878_), .A4(new_n1879_), .ZN(new_n1880_));
  NOR3_X1    g01816(.A1(new_n1880_), .A2(new_n1870_), .A3(new_n1874_), .ZN(new_n1881_));
  NAND3_X1   g01817(.A1(new_n1881_), .A2(new_n1196_), .A3(new_n1082_), .ZN(new_n1882_));
  OAI22_X1   g01818(.A1(new_n69_), .A2(new_n73_), .B1(new_n129_), .B2(new_n66_), .ZN(new_n1883_));
  NAND2_X1   g01819(.A1(new_n755_), .A2(new_n1883_), .ZN(new_n1884_));
  NOR4_X1    g01820(.A1(new_n289_), .A2(new_n376_), .A3(new_n749_), .A4(new_n310_), .ZN(new_n1885_));
  NOR4_X1    g01821(.A1(new_n262_), .A2(new_n307_), .A3(new_n577_), .A4(new_n682_), .ZN(new_n1886_));
  NOR4_X1    g01822(.A1(new_n1886_), .A2(new_n1884_), .A3(new_n1885_), .A4(new_n1389_), .ZN(new_n1887_));
  NAND3_X1   g01823(.A1(new_n1058_), .A2(new_n1706_), .A3(new_n110_), .ZN(new_n1888_));
  OAI22_X1   g01824(.A1(new_n73_), .A2(new_n91_), .B1(new_n85_), .B2(new_n123_), .ZN(new_n1889_));
  NAND2_X1   g01825(.A1(new_n1679_), .A2(new_n1889_), .ZN(new_n1890_));
  NAND2_X1   g01826(.A1(new_n180_), .A2(new_n245_), .ZN(new_n1891_));
  NAND2_X1   g01827(.A1(new_n79_), .A2(new_n355_), .ZN(new_n1892_));
  NAND3_X1   g01828(.A1(new_n410_), .A2(new_n1892_), .A3(new_n1891_), .ZN(new_n1893_));
  NOR4_X1    g01829(.A1(new_n366_), .A2(new_n1031_), .A3(new_n817_), .A4(new_n556_), .ZN(new_n1894_));
  NOR4_X1    g01830(.A1(new_n1890_), .A2(new_n1894_), .A3(new_n1893_), .A4(new_n1888_), .ZN(new_n1895_));
  OAI21_X1   g01831(.A1(new_n318_), .A2(new_n158_), .B(new_n180_), .ZN(new_n1896_));
  NAND4_X1   g01832(.A1(new_n1896_), .A2(new_n395_), .A3(new_n1448_), .A4(new_n522_), .ZN(new_n1897_));
  NAND4_X1   g01833(.A1(new_n1199_), .A2(new_n1216_), .A3(new_n1745_), .A4(new_n980_), .ZN(new_n1898_));
  NOR2_X1    g01834(.A1(new_n1898_), .A2(new_n1897_), .ZN(new_n1899_));
  NAND3_X1   g01835(.A1(new_n1895_), .A2(new_n1887_), .A3(new_n1899_), .ZN(new_n1900_));
  NOR3_X1    g01836(.A1(new_n533_), .A2(new_n396_), .A3(new_n756_), .ZN(new_n1901_));
  NOR2_X1    g01837(.A1(new_n211_), .A2(new_n689_), .ZN(new_n1902_));
  NOR2_X1    g01838(.A1(new_n86_), .A2(new_n955_), .ZN(new_n1903_));
  NOR4_X1    g01839(.A1(new_n1902_), .A2(new_n1615_), .A3(new_n1903_), .A4(new_n1627_), .ZN(new_n1904_));
  NOR2_X1    g01840(.A1(new_n1821_), .A2(new_n1822_), .ZN(new_n1905_));
  NAND3_X1   g01841(.A1(new_n1904_), .A2(new_n1905_), .A3(new_n1901_), .ZN(new_n1906_));
  NOR4_X1    g01842(.A1(new_n633_), .A2(new_n124_), .A3(new_n132_), .A4(new_n397_), .ZN(new_n1907_));
  NAND4_X1   g01843(.A1(new_n1825_), .A2(new_n361_), .A3(new_n729_), .A4(new_n680_), .ZN(new_n1908_));
  NOR2_X1    g01844(.A1(new_n1908_), .A2(new_n1907_), .ZN(new_n1909_));
  NAND3_X1   g01845(.A1(new_n322_), .A2(new_n1759_), .A3(new_n1585_), .ZN(new_n1910_));
  NOR3_X1    g01846(.A1(new_n534_), .A2(new_n178_), .A3(new_n681_), .ZN(new_n1911_));
  NOR4_X1    g01847(.A1(new_n335_), .A2(new_n531_), .A3(new_n487_), .A4(new_n418_), .ZN(new_n1912_));
  NOR3_X1    g01848(.A1(new_n1912_), .A2(new_n1911_), .A3(new_n1910_), .ZN(new_n1913_));
  NOR2_X1    g01849(.A1(new_n779_), .A2(new_n70_), .ZN(new_n1914_));
  NOR2_X1    g01850(.A1(new_n203_), .A2(new_n488_), .ZN(new_n1915_));
  NOR3_X1    g01851(.A1(new_n1914_), .A2(new_n1915_), .A3(new_n1147_), .ZN(new_n1916_));
  NAND3_X1   g01852(.A1(new_n834_), .A2(new_n373_), .A3(new_n1838_), .ZN(new_n1917_));
  NOR4_X1    g01853(.A1(new_n1917_), .A2(new_n306_), .A3(new_n422_), .A4(new_n587_), .ZN(new_n1918_));
  NAND4_X1   g01854(.A1(new_n1909_), .A2(new_n1913_), .A3(new_n1918_), .A4(new_n1916_), .ZN(new_n1919_));
  NAND4_X1   g01855(.A1(new_n848_), .A2(new_n208_), .A3(new_n1582_), .A4(new_n1719_), .ZN(new_n1920_));
  NAND2_X1   g01856(.A1(new_n158_), .A2(new_n156_), .ZN(new_n1921_));
  NAND3_X1   g01857(.A1(new_n1921_), .A2(new_n512_), .A3(new_n985_), .ZN(new_n1922_));
  OAI22_X1   g01858(.A1(new_n334_), .A2(new_n175_), .B1(new_n75_), .B2(new_n153_), .ZN(new_n1923_));
  NAND4_X1   g01859(.A1(new_n1923_), .A2(new_n113_), .A3(new_n188_), .A4(new_n378_), .ZN(new_n1924_));
  NOR3_X1    g01860(.A1(new_n1924_), .A2(new_n1920_), .A3(new_n1922_), .ZN(new_n1925_));
  NOR4_X1    g01861(.A1(new_n117_), .A2(new_n648_), .A3(new_n574_), .A4(new_n506_), .ZN(new_n1926_));
  NAND3_X1   g01862(.A1(new_n1070_), .A2(new_n1067_), .A3(new_n1465_), .ZN(new_n1927_));
  NOR4_X1    g01863(.A1(new_n1926_), .A2(new_n1927_), .A3(new_n593_), .A4(new_n867_), .ZN(new_n1928_));
  NAND3_X1   g01864(.A1(new_n393_), .A2(new_n509_), .A3(new_n984_), .ZN(new_n1929_));
  OAI21_X1   g01865(.A1(new_n108_), .A2(new_n143_), .B(new_n77_), .ZN(new_n1930_));
  NAND3_X1   g01866(.A1(new_n1930_), .A2(new_n1212_), .A3(new_n709_), .ZN(new_n1931_));
  NOR4_X1    g01867(.A1(new_n1167_), .A2(new_n752_), .A3(new_n610_), .A4(new_n490_), .ZN(new_n1932_));
  NOR4_X1    g01868(.A1(new_n281_), .A2(new_n370_), .A3(new_n549_), .A4(new_n1073_), .ZN(new_n1933_));
  NOR4_X1    g01869(.A1(new_n1932_), .A2(new_n1933_), .A3(new_n1929_), .A4(new_n1931_), .ZN(new_n1934_));
  NAND2_X1   g01870(.A1(new_n404_), .A2(new_n273_), .ZN(new_n1935_));
  NAND4_X1   g01871(.A1(new_n1856_), .A2(new_n568_), .A3(new_n1935_), .A4(new_n409_), .ZN(new_n1936_));
  NOR4_X1    g01872(.A1(new_n1936_), .A2(new_n935_), .A3(new_n544_), .A4(new_n1858_), .ZN(new_n1937_));
  NAND4_X1   g01873(.A1(new_n1934_), .A2(new_n1925_), .A3(new_n1937_), .A4(new_n1928_), .ZN(new_n1938_));
  NOR4_X1    g01874(.A1(new_n1938_), .A2(new_n1900_), .A3(new_n1919_), .A4(new_n1906_), .ZN(new_n1939_));
  NAND2_X1   g01875(.A1(new_n1939_), .A2(new_n1882_), .ZN(new_n1940_));
  AOI21_X1   g01876(.A1(new_n1863_), .A2(new_n1940_), .B(new_n1813_), .ZN(new_n1941_));
  NAND2_X1   g01877(.A1(new_n1091_), .A2(new_n978_), .ZN(new_n1942_));
  NAND4_X1   g01878(.A1(new_n1942_), .A2(new_n1025_), .A3(new_n405_), .A4(new_n1468_), .ZN(new_n1943_));
  NOR2_X1    g01879(.A1(new_n149_), .A2(new_n724_), .ZN(new_n1944_));
  NOR2_X1    g01880(.A1(new_n1944_), .A2(new_n1864_), .ZN(new_n1945_));
  AOI22_X1   g01881(.A1(new_n325_), .A2(new_n980_), .B1(new_n1067_), .B2(new_n390_), .ZN(new_n1946_));
  NAND2_X1   g01882(.A1(new_n1945_), .A2(new_n1946_), .ZN(new_n1947_));
  NOR3_X1    g01883(.A1(new_n1947_), .A2(new_n1607_), .A3(new_n1943_), .ZN(new_n1948_));
  NAND2_X1   g01884(.A1(new_n1563_), .A2(new_n441_), .ZN(new_n1949_));
  AOI22_X1   g01885(.A1(new_n1646_), .A2(new_n1838_), .B1(new_n1506_), .B2(new_n222_), .ZN(new_n1950_));
  NAND3_X1   g01886(.A1(new_n1950_), .A2(new_n1210_), .A3(new_n1949_), .ZN(new_n1951_));
  OAI22_X1   g01887(.A1(new_n75_), .A2(new_n115_), .B1(new_n66_), .B2(new_n150_), .ZN(new_n1952_));
  NAND2_X1   g01888(.A1(new_n1829_), .A2(new_n824_), .ZN(new_n1953_));
  AOI21_X1   g01889(.A1(new_n73_), .A2(new_n133_), .B(new_n123_), .ZN(new_n1954_));
  INV_X1     g01890(.I(new_n1954_), .ZN(new_n1955_));
  NAND4_X1   g01891(.A1(new_n1953_), .A2(new_n631_), .A3(new_n1955_), .A4(new_n1952_), .ZN(new_n1956_));
  NOR2_X1    g01892(.A1(new_n1951_), .A2(new_n1956_), .ZN(new_n1957_));
  NAND2_X1   g01893(.A1(new_n385_), .A2(new_n856_), .ZN(new_n1958_));
  NAND4_X1   g01894(.A1(new_n1958_), .A2(new_n967_), .A3(new_n1244_), .A4(new_n1326_), .ZN(new_n1959_));
  INV_X1     g01895(.I(new_n163_), .ZN(new_n1960_));
  NAND2_X1   g01896(.A1(new_n302_), .A2(new_n1647_), .ZN(new_n1961_));
  AOI21_X1   g01897(.A1(new_n176_), .A2(new_n115_), .B(new_n129_), .ZN(new_n1962_));
  INV_X1     g01898(.I(new_n1962_), .ZN(new_n1963_));
  NAND4_X1   g01899(.A1(new_n708_), .A2(new_n1961_), .A3(new_n1963_), .A4(new_n1960_), .ZN(new_n1964_));
  NOR2_X1    g01900(.A1(new_n1959_), .A2(new_n1964_), .ZN(new_n1965_));
  NAND3_X1   g01901(.A1(new_n1948_), .A2(new_n1965_), .A3(new_n1957_), .ZN(new_n1966_));
  INV_X1     g01902(.I(new_n291_), .ZN(new_n1967_));
  NOR2_X1    g01903(.A1(new_n734_), .A2(new_n801_), .ZN(new_n1968_));
  NAND2_X1   g01904(.A1(new_n1968_), .A2(new_n655_), .ZN(new_n1969_));
  NAND2_X1   g01905(.A1(new_n1495_), .A2(new_n992_), .ZN(new_n1970_));
  NOR4_X1    g01906(.A1(new_n268_), .A2(new_n648_), .A3(new_n1031_), .A4(new_n191_), .ZN(new_n1971_));
  NOR4_X1    g01907(.A1(new_n1970_), .A2(new_n1969_), .A3(new_n500_), .A4(new_n1971_), .ZN(new_n1972_));
  NOR4_X1    g01908(.A1(new_n1531_), .A2(new_n226_), .A3(new_n370_), .A4(new_n744_), .ZN(new_n1973_));
  NAND2_X1   g01909(.A1(new_n1396_), .A2(new_n250_), .ZN(new_n1974_));
  NOR3_X1    g01910(.A1(new_n1973_), .A2(new_n190_), .A3(new_n1974_), .ZN(new_n1975_));
  NAND2_X1   g01911(.A1(new_n436_), .A2(new_n423_), .ZN(new_n1976_));
  NOR4_X1    g01912(.A1(new_n161_), .A2(new_n1328_), .A3(new_n1976_), .A4(new_n114_), .ZN(new_n1977_));
  NAND4_X1   g01913(.A1(new_n1972_), .A2(new_n1967_), .A3(new_n1975_), .A4(new_n1977_), .ZN(new_n1978_));
  NOR4_X1    g01914(.A1(new_n1139_), .A2(new_n1343_), .A3(new_n1915_), .A4(new_n1541_), .ZN(new_n1979_));
  NOR4_X1    g01915(.A1(new_n496_), .A2(new_n779_), .A3(new_n549_), .A4(new_n125_), .ZN(new_n1980_));
  NAND3_X1   g01916(.A1(new_n233_), .A2(new_n1706_), .A3(new_n1719_), .ZN(new_n1981_));
  NOR2_X1    g01917(.A1(new_n1981_), .A2(new_n1980_), .ZN(new_n1982_));
  NAND2_X1   g01918(.A1(new_n1979_), .A2(new_n1982_), .ZN(new_n1983_));
  NOR2_X1    g01919(.A1(new_n171_), .A2(new_n334_), .ZN(new_n1984_));
  NOR2_X1    g01920(.A1(new_n1984_), .A2(new_n367_), .ZN(new_n1985_));
  NOR4_X1    g01921(.A1(new_n1985_), .A2(new_n805_), .A3(new_n1493_), .A4(new_n697_), .ZN(new_n1986_));
  NOR2_X1    g01922(.A1(new_n90_), .A2(new_n741_), .ZN(new_n1987_));
  NAND2_X1   g01923(.A1(new_n739_), .A2(new_n349_), .ZN(new_n1988_));
  NOR4_X1    g01924(.A1(new_n530_), .A2(new_n1802_), .A3(new_n1988_), .A4(new_n1987_), .ZN(new_n1989_));
  NOR2_X1    g01925(.A1(new_n753_), .A2(new_n517_), .ZN(new_n1990_));
  NOR2_X1    g01926(.A1(new_n684_), .A2(new_n594_), .ZN(new_n1991_));
  NOR2_X1    g01927(.A1(new_n219_), .A2(new_n235_), .ZN(new_n1992_));
  NOR3_X1    g01928(.A1(new_n1992_), .A2(new_n1990_), .A3(new_n1991_), .ZN(new_n1993_));
  NOR2_X1    g01929(.A1(new_n252_), .A2(new_n1168_), .ZN(new_n1994_));
  NOR2_X1    g01930(.A1(new_n582_), .A2(new_n330_), .ZN(new_n1995_));
  AOI21_X1   g01931(.A1(new_n175_), .A2(new_n116_), .B(new_n95_), .ZN(new_n1996_));
  NOR4_X1    g01932(.A1(new_n1994_), .A2(new_n1995_), .A3(new_n1112_), .A4(new_n1996_), .ZN(new_n1997_));
  NAND4_X1   g01933(.A1(new_n1989_), .A2(new_n1997_), .A3(new_n1986_), .A4(new_n1993_), .ZN(new_n1998_));
  NOR4_X1    g01934(.A1(new_n1966_), .A2(new_n1978_), .A3(new_n1983_), .A4(new_n1998_), .ZN(new_n1999_));
  NOR3_X1    g01935(.A1(new_n1999_), .A2(new_n1882_), .A3(new_n1939_), .ZN(new_n2000_));
  NOR2_X1    g01936(.A1(new_n1941_), .A2(new_n2000_), .ZN(new_n2001_));
  NAND2_X1   g01937(.A1(new_n2001_), .A2(new_n1613_), .ZN(new_n2002_));
  AOI21_X1   g01938(.A1(new_n2002_), .A2(new_n1764_), .B(new_n1729_), .ZN(new_n2003_));
  OAI21_X1   g01939(.A1(new_n2001_), .A2(new_n1613_), .B(new_n1763_), .ZN(new_n2004_));
  INV_X1     g01940(.I(new_n2004_), .ZN(new_n2005_));
  NOR2_X1    g01941(.A1(new_n2003_), .A2(new_n2005_), .ZN(new_n2006_));
  NOR4_X1    g01942(.A1(new_n486_), .A2(new_n130_), .A3(new_n590_), .A4(new_n163_), .ZN(new_n2007_));
  NOR4_X1    g01943(.A1(new_n2007_), .A2(new_n226_), .A3(new_n804_), .A4(new_n602_), .ZN(new_n2008_));
  INV_X1     g01944(.I(new_n2008_), .ZN(new_n2009_));
  NOR4_X1    g01945(.A1(new_n714_), .A2(new_n286_), .A3(new_n517_), .A4(new_n535_), .ZN(new_n2010_));
  NOR2_X1    g01946(.A1(new_n656_), .A2(new_n203_), .ZN(new_n2011_));
  NOR2_X1    g01947(.A1(new_n132_), .A2(new_n749_), .ZN(new_n2012_));
  NOR2_X1    g01948(.A1(new_n173_), .A2(new_n384_), .ZN(new_n2013_));
  NAND4_X1   g01949(.A1(new_n2011_), .A2(new_n1835_), .A3(new_n2012_), .A4(new_n2013_), .ZN(new_n2014_));
  NOR3_X1    g01950(.A1(new_n2009_), .A2(new_n2014_), .A3(new_n2010_), .ZN(new_n2015_));
  NOR4_X1    g01951(.A1(new_n1027_), .A2(new_n712_), .A3(new_n262_), .A4(new_n611_), .ZN(new_n2016_));
  NAND4_X1   g01952(.A1(new_n2016_), .A2(new_n511_), .A3(new_n816_), .A4(new_n1467_), .ZN(new_n2017_));
  NAND4_X1   g01953(.A1(new_n675_), .A2(new_n807_), .A3(new_n1105_), .A4(new_n665_), .ZN(new_n2018_));
  NOR3_X1    g01954(.A1(new_n1589_), .A2(new_n192_), .A3(new_n447_), .ZN(new_n2019_));
  NOR4_X1    g01955(.A1(new_n149_), .A2(new_n297_), .A3(new_n335_), .A4(new_n610_), .ZN(new_n2020_));
  INV_X1     g01956(.I(new_n2020_), .ZN(new_n2021_));
  NOR2_X1    g01957(.A1(new_n282_), .A2(new_n227_), .ZN(new_n2022_));
  INV_X1     g01958(.I(new_n2022_), .ZN(new_n2023_));
  NOR2_X1    g01959(.A1(new_n1365_), .A2(new_n2023_), .ZN(new_n2024_));
  NAND4_X1   g01960(.A1(new_n2024_), .A2(new_n2019_), .A3(new_n2018_), .A4(new_n2021_), .ZN(new_n2025_));
  NOR2_X1    g01961(.A1(new_n563_), .A2(new_n1976_), .ZN(new_n2026_));
  NAND4_X1   g01962(.A1(new_n797_), .A2(new_n144_), .A3(new_n405_), .A4(new_n464_), .ZN(new_n2027_));
  NAND4_X1   g01963(.A1(new_n2026_), .A2(new_n745_), .A3(new_n1064_), .A4(new_n2027_), .ZN(new_n2028_));
  NOR3_X1    g01964(.A1(new_n2017_), .A2(new_n2025_), .A3(new_n2028_), .ZN(new_n2029_));
  NAND2_X1   g01965(.A1(new_n2029_), .A2(new_n2015_), .ZN(new_n2030_));
  NAND2_X1   g01966(.A1(new_n188_), .A2(new_n1325_), .ZN(new_n2031_));
  NOR4_X1    g01967(.A1(new_n2031_), .A2(new_n70_), .A3(new_n305_), .A4(new_n1184_), .ZN(new_n2032_));
  NOR2_X1    g01968(.A1(new_n488_), .A2(new_n682_), .ZN(new_n2033_));
  NAND2_X1   g01969(.A1(new_n1156_), .A2(new_n2033_), .ZN(new_n2034_));
  INV_X1     g01970(.I(new_n2034_), .ZN(new_n2035_));
  NAND4_X1   g01971(.A1(new_n371_), .A2(new_n2035_), .A3(new_n972_), .A4(new_n2032_), .ZN(new_n2036_));
  NOR3_X1    g01972(.A1(new_n2036_), .A2(new_n625_), .A3(new_n515_), .ZN(new_n2037_));
  NOR2_X1    g01973(.A1(new_n531_), .A2(new_n549_), .ZN(new_n2038_));
  INV_X1     g01974(.I(new_n2038_), .ZN(new_n2039_));
  NOR2_X1    g01975(.A1(new_n899_), .A2(new_n333_), .ZN(new_n2040_));
  INV_X1     g01976(.I(new_n2040_), .ZN(new_n2041_));
  INV_X1     g01977(.I(new_n1441_), .ZN(new_n2042_));
  NOR3_X1    g01978(.A1(new_n2039_), .A2(new_n2041_), .A3(new_n2042_), .ZN(new_n2043_));
  NOR3_X1    g01979(.A1(new_n607_), .A2(new_n307_), .A3(new_n561_), .ZN(new_n2044_));
  NOR3_X1    g01980(.A1(new_n530_), .A2(new_n490_), .A3(new_n1152_), .ZN(new_n2045_));
  NOR2_X1    g01981(.A1(new_n751_), .A2(new_n239_), .ZN(new_n2046_));
  INV_X1     g01982(.I(new_n2046_), .ZN(new_n2047_));
  NOR2_X1    g01983(.A1(new_n2047_), .A2(new_n713_), .ZN(new_n2048_));
  NAND4_X1   g01984(.A1(new_n2043_), .A2(new_n2045_), .A3(new_n2048_), .A4(new_n2044_), .ZN(new_n2049_));
  INV_X1     g01985(.I(new_n2049_), .ZN(new_n2050_));
  NAND2_X1   g01986(.A1(new_n851_), .A2(new_n706_), .ZN(new_n2051_));
  NAND2_X1   g01987(.A1(new_n378_), .A2(new_n978_), .ZN(new_n2052_));
  NOR2_X1    g01988(.A1(new_n1994_), .A2(new_n2052_), .ZN(new_n2053_));
  NAND4_X1   g01989(.A1(new_n2053_), .A2(new_n1666_), .A3(new_n824_), .A4(new_n1796_), .ZN(new_n2054_));
  INV_X1     g01990(.I(new_n261_), .ZN(new_n2055_));
  NAND2_X1   g01991(.A1(new_n2055_), .A2(new_n872_), .ZN(new_n2056_));
  NOR4_X1    g01992(.A1(new_n121_), .A2(new_n332_), .A3(new_n2056_), .A4(new_n689_), .ZN(new_n2057_));
  NAND2_X1   g01993(.A1(new_n2057_), .A2(new_n1273_), .ZN(new_n2058_));
  NOR4_X1    g01994(.A1(new_n2058_), .A2(new_n958_), .A3(new_n2051_), .A4(new_n2054_), .ZN(new_n2059_));
  NOR4_X1    g01995(.A1(new_n687_), .A2(new_n306_), .A3(new_n398_), .A4(new_n544_), .ZN(new_n2060_));
  NAND4_X1   g01996(.A1(new_n2060_), .A2(new_n395_), .A3(new_n761_), .A4(new_n880_), .ZN(new_n2061_));
  NOR4_X1    g01997(.A1(new_n288_), .A2(new_n867_), .A3(new_n154_), .A4(new_n280_), .ZN(new_n2062_));
  NAND3_X1   g01998(.A1(new_n1404_), .A2(new_n568_), .A3(new_n1638_), .ZN(new_n2063_));
  NOR2_X1    g01999(.A1(new_n191_), .A2(new_n347_), .ZN(new_n2064_));
  INV_X1     g02000(.I(new_n2064_), .ZN(new_n2065_));
  NAND2_X1   g02001(.A1(new_n1009_), .A2(new_n983_), .ZN(new_n2066_));
  NOR4_X1    g02002(.A1(new_n2063_), .A2(new_n2065_), .A3(new_n2062_), .A4(new_n2066_), .ZN(new_n2067_));
  INV_X1     g02003(.I(new_n2067_), .ZN(new_n2068_));
  NOR2_X1    g02004(.A1(new_n2061_), .A2(new_n2068_), .ZN(new_n2069_));
  NAND4_X1   g02005(.A1(new_n2059_), .A2(new_n2037_), .A3(new_n2050_), .A4(new_n2069_), .ZN(new_n2070_));
  NOR2_X1    g02006(.A1(new_n2070_), .A2(new_n2030_), .ZN(new_n2071_));
  OAI21_X1   g02007(.A1(new_n2006_), .A2(new_n2071_), .B(new_n1678_), .ZN(new_n2072_));
  NAND2_X1   g02008(.A1(new_n2072_), .A2(new_n1613_), .ZN(new_n2073_));
  INV_X1     g02009(.I(new_n1678_), .ZN(new_n2074_));
  NAND2_X1   g02010(.A1(new_n2006_), .A2(new_n2071_), .ZN(new_n2075_));
  NAND2_X1   g02011(.A1(new_n2075_), .A2(new_n2074_), .ZN(new_n2076_));
  NAND2_X1   g02012(.A1(new_n378_), .A2(new_n880_), .ZN(new_n2077_));
  NOR4_X1    g02013(.A1(new_n238_), .A2(new_n670_), .A3(new_n298_), .A4(new_n518_), .ZN(new_n2078_));
  INV_X1     g02014(.I(new_n530_), .ZN(new_n2079_));
  NAND2_X1   g02015(.A1(new_n2079_), .A2(new_n1070_), .ZN(new_n2080_));
  NOR4_X1    g02016(.A1(new_n2080_), .A2(new_n2077_), .A3(new_n1211_), .A4(new_n2078_), .ZN(new_n2081_));
  NOR2_X1    g02017(.A1(new_n666_), .A2(new_n837_), .ZN(new_n2082_));
  INV_X1     g02018(.I(new_n2082_), .ZN(new_n2083_));
  NOR3_X1    g02019(.A1(new_n2083_), .A2(new_n2039_), .A3(new_n1431_), .ZN(new_n2084_));
  NAND4_X1   g02020(.A1(new_n2081_), .A2(new_n1287_), .A3(new_n1509_), .A4(new_n2084_), .ZN(new_n2085_));
  INV_X1     g02021(.I(new_n2085_), .ZN(new_n2086_));
  NOR3_X1    g02022(.A1(new_n825_), .A2(new_n183_), .A3(new_n1865_), .ZN(new_n2087_));
  INV_X1     g02023(.I(new_n2087_), .ZN(new_n2088_));
  NOR3_X1    g02024(.A1(new_n1518_), .A2(new_n124_), .A3(new_n525_), .ZN(new_n2089_));
  INV_X1     g02025(.I(new_n2089_), .ZN(new_n2090_));
  NOR2_X1    g02026(.A1(new_n652_), .A2(new_n1152_), .ZN(new_n2091_));
  INV_X1     g02027(.I(new_n2091_), .ZN(new_n2092_));
  NOR3_X1    g02028(.A1(new_n2092_), .A2(new_n642_), .A3(new_n1011_), .ZN(new_n2093_));
  INV_X1     g02029(.I(new_n2093_), .ZN(new_n2094_));
  INV_X1     g02030(.I(new_n1131_), .ZN(new_n2095_));
  INV_X1     g02031(.I(new_n766_), .ZN(new_n2096_));
  NOR3_X1    g02032(.A1(new_n2096_), .A2(new_n939_), .A3(new_n1266_), .ZN(new_n2097_));
  INV_X1     g02033(.I(new_n1579_), .ZN(new_n2098_));
  NOR4_X1    g02034(.A1(new_n1669_), .A2(new_n2098_), .A3(new_n465_), .A4(new_n783_), .ZN(new_n2099_));
  NAND4_X1   g02035(.A1(new_n2097_), .A2(new_n1015_), .A3(new_n2099_), .A4(new_n2095_), .ZN(new_n2100_));
  NOR4_X1    g02036(.A1(new_n2100_), .A2(new_n2088_), .A3(new_n2090_), .A4(new_n2094_), .ZN(new_n2101_));
  NAND3_X1   g02037(.A1(new_n1364_), .A2(new_n2086_), .A3(new_n2101_), .ZN(new_n2102_));
  INV_X1     g02038(.I(new_n2102_), .ZN(new_n2103_));
  NOR2_X1    g02039(.A1(new_n2103_), .A2(new_n2071_), .ZN(new_n2104_));
  INV_X1     g02040(.I(new_n2104_), .ZN(new_n2105_));
  NAND3_X1   g02041(.A1(new_n2073_), .A2(new_n2076_), .A3(new_n2105_), .ZN(new_n2106_));
  INV_X1     g02042(.I(new_n2071_), .ZN(new_n2107_));
  NOR2_X1    g02043(.A1(new_n2102_), .A2(new_n2107_), .ZN(new_n2108_));
  INV_X1     g02044(.I(new_n2108_), .ZN(new_n2109_));
  NAND2_X1   g02045(.A1(new_n385_), .A2(new_n1647_), .ZN(new_n2110_));
  NAND2_X1   g02046(.A1(new_n1214_), .A2(new_n2012_), .ZN(new_n2111_));
  NOR4_X1    g02047(.A1(new_n1031_), .A2(new_n90_), .A3(new_n125_), .A4(new_n594_), .ZN(new_n2112_));
  INV_X1     g02048(.I(new_n1664_), .ZN(new_n2113_));
  NOR4_X1    g02049(.A1(new_n198_), .A2(new_n106_), .A3(new_n236_), .A4(new_n418_), .ZN(new_n2114_));
  NAND3_X1   g02050(.A1(new_n2113_), .A2(new_n729_), .A3(new_n2114_), .ZN(new_n2115_));
  NOR4_X1    g02051(.A1(new_n2115_), .A2(new_n2110_), .A3(new_n2111_), .A4(new_n2112_), .ZN(new_n2116_));
  NOR4_X1    g02052(.A1(new_n463_), .A2(new_n587_), .A3(new_n1073_), .A4(new_n310_), .ZN(new_n2117_));
  NOR4_X1    g02053(.A1(new_n946_), .A2(new_n1084_), .A3(new_n242_), .A4(new_n460_), .ZN(new_n2118_));
  INV_X1     g02054(.I(new_n255_), .ZN(new_n2119_));
  NAND4_X1   g02055(.A1(new_n913_), .A2(new_n2119_), .A3(new_n358_), .A4(new_n361_), .ZN(new_n2120_));
  NOR3_X1    g02056(.A1(new_n2118_), .A2(new_n2120_), .A3(new_n2117_), .ZN(new_n2121_));
  NOR2_X1    g02057(.A1(new_n656_), .A2(new_n70_), .ZN(new_n2122_));
  NOR2_X1    g02058(.A1(new_n719_), .A2(new_n556_), .ZN(new_n2123_));
  AOI21_X1   g02059(.A1(new_n2122_), .A2(new_n2123_), .B(new_n1037_), .ZN(new_n2124_));
  INV_X1     g02060(.I(new_n825_), .ZN(new_n2125_));
  NAND4_X1   g02061(.A1(new_n2125_), .A2(new_n852_), .A3(new_n1766_), .A4(new_n927_), .ZN(new_n2126_));
  NOR2_X1    g02062(.A1(new_n1278_), .A2(new_n2126_), .ZN(new_n2127_));
  NAND4_X1   g02063(.A1(new_n2127_), .A2(new_n2116_), .A3(new_n2121_), .A4(new_n2124_), .ZN(new_n2128_));
  NAND4_X1   g02064(.A1(new_n667_), .A2(new_n795_), .A3(new_n188_), .A4(new_n592_), .ZN(new_n2129_));
  NOR2_X1    g02065(.A1(new_n1211_), .A2(new_n517_), .ZN(new_n2130_));
  NOR4_X1    g02066(.A1(new_n320_), .A2(new_n420_), .A3(new_n776_), .A4(new_n715_), .ZN(new_n2131_));
  NAND3_X1   g02067(.A1(new_n2130_), .A2(new_n2129_), .A3(new_n2131_), .ZN(new_n2132_));
  NOR4_X1    g02068(.A1(new_n225_), .A2(new_n654_), .A3(new_n449_), .A4(new_n1167_), .ZN(new_n2133_));
  NOR4_X1    g02069(.A1(new_n866_), .A2(new_n288_), .A3(new_n387_), .A4(new_n459_), .ZN(new_n2134_));
  INV_X1     g02070(.I(new_n828_), .ZN(new_n2135_));
  NOR2_X1    g02071(.A1(new_n2135_), .A2(new_n1337_), .ZN(new_n2136_));
  INV_X1     g02072(.I(new_n723_), .ZN(new_n2137_));
  NAND2_X1   g02073(.A1(new_n1853_), .A2(new_n464_), .ZN(new_n2138_));
  NOR4_X1    g02074(.A1(new_n2137_), .A2(new_n781_), .A3(new_n1527_), .A4(new_n2138_), .ZN(new_n2139_));
  NAND3_X1   g02075(.A1(new_n2136_), .A2(new_n2139_), .A3(new_n1516_), .ZN(new_n2140_));
  NOR4_X1    g02076(.A1(new_n2140_), .A2(new_n2132_), .A3(new_n2133_), .A4(new_n2134_), .ZN(new_n2141_));
  NOR2_X1    g02077(.A1(new_n648_), .A2(new_n596_), .ZN(new_n2142_));
  NAND4_X1   g02078(.A1(new_n1248_), .A2(new_n336_), .A3(new_n1796_), .A4(new_n2142_), .ZN(new_n2143_));
  INV_X1     g02079(.I(new_n2143_), .ZN(new_n2144_));
  NOR2_X1    g02080(.A1(new_n770_), .A2(new_n753_), .ZN(new_n2145_));
  INV_X1     g02081(.I(new_n536_), .ZN(new_n2146_));
  NOR2_X1    g02082(.A1(new_n2146_), .A2(new_n523_), .ZN(new_n2147_));
  NOR2_X1    g02083(.A1(new_n326_), .A2(new_n164_), .ZN(new_n2148_));
  INV_X1     g02084(.I(new_n2148_), .ZN(new_n2149_));
  NOR4_X1    g02085(.A1(new_n2149_), .A2(new_n565_), .A3(new_n1262_), .A4(new_n1055_), .ZN(new_n2150_));
  NAND4_X1   g02086(.A1(new_n2144_), .A2(new_n2150_), .A3(new_n2145_), .A4(new_n2147_), .ZN(new_n2151_));
  NAND4_X1   g02087(.A1(new_n292_), .A2(new_n405_), .A3(new_n1572_), .A4(new_n983_), .ZN(new_n2152_));
  NOR3_X1    g02088(.A1(new_n530_), .A2(new_n92_), .A3(new_n415_), .ZN(new_n2153_));
  NOR3_X1    g02089(.A1(new_n76_), .A2(new_n782_), .A3(new_n731_), .ZN(new_n2154_));
  NAND4_X1   g02090(.A1(new_n1598_), .A2(new_n2152_), .A3(new_n2153_), .A4(new_n2154_), .ZN(new_n2155_));
  NOR2_X1    g02091(.A1(new_n2155_), .A2(new_n2151_), .ZN(new_n2156_));
  NAND2_X1   g02092(.A1(new_n2156_), .A2(new_n2141_), .ZN(new_n2157_));
  NOR2_X1    g02093(.A1(new_n2157_), .A2(new_n2128_), .ZN(new_n2158_));
  NOR2_X1    g02094(.A1(new_n2103_), .A2(new_n2158_), .ZN(new_n2159_));
  AOI21_X1   g02095(.A1(new_n2106_), .A2(new_n2109_), .B(new_n2159_), .ZN(new_n2160_));
  INV_X1     g02096(.I(new_n2158_), .ZN(new_n2161_));
  NOR2_X1    g02097(.A1(new_n2161_), .A2(new_n2102_), .ZN(new_n2162_));
  INV_X1     g02098(.I(new_n1520_), .ZN(new_n2163_));
  INV_X1     g02099(.I(new_n1976_), .ZN(new_n2164_));
  NOR2_X1    g02100(.A1(new_n590_), .A2(new_n333_), .ZN(new_n2165_));
  NAND4_X1   g02101(.A1(new_n2164_), .A2(new_n1111_), .A3(new_n887_), .A4(new_n2165_), .ZN(new_n2166_));
  NOR3_X1    g02102(.A1(new_n1175_), .A2(new_n487_), .A3(new_n556_), .ZN(new_n2167_));
  INV_X1     g02103(.I(new_n2167_), .ZN(new_n2168_));
  NOR4_X1    g02104(.A1(new_n648_), .A2(new_n1146_), .A3(new_n474_), .A4(new_n506_), .ZN(new_n2169_));
  NOR4_X1    g02105(.A1(new_n2166_), .A2(new_n2163_), .A3(new_n2168_), .A4(new_n2169_), .ZN(new_n2170_));
  NOR4_X1    g02106(.A1(new_n403_), .A2(new_n779_), .A3(new_n496_), .A4(new_n370_), .ZN(new_n2171_));
  NOR4_X1    g02107(.A1(new_n788_), .A2(new_n534_), .A3(new_n214_), .A4(new_n280_), .ZN(new_n2172_));
  NOR4_X1    g02108(.A1(new_n219_), .A2(new_n419_), .A3(new_n776_), .A4(new_n1092_), .ZN(new_n2173_));
  NOR3_X1    g02109(.A1(new_n2172_), .A2(new_n2171_), .A3(new_n2173_), .ZN(new_n2174_));
  NOR2_X1    g02110(.A1(new_n335_), .A2(new_n320_), .ZN(new_n2175_));
  INV_X1     g02111(.I(new_n2175_), .ZN(new_n2176_));
  NOR4_X1    g02112(.A1(new_n462_), .A2(new_n544_), .A3(new_n1185_), .A4(new_n2176_), .ZN(new_n2177_));
  INV_X1     g02113(.I(new_n482_), .ZN(new_n2178_));
  NAND4_X1   g02114(.A1(new_n2178_), .A2(new_n358_), .A3(new_n361_), .A4(new_n871_), .ZN(new_n2179_));
  NAND3_X1   g02115(.A1(new_n2179_), .A2(new_n1026_), .A3(new_n1419_), .ZN(new_n2180_));
  NOR3_X1    g02116(.A1(new_n835_), .A2(new_n594_), .A3(new_n1858_), .ZN(new_n2181_));
  INV_X1     g02117(.I(new_n2181_), .ZN(new_n2182_));
  NOR2_X1    g02118(.A1(new_n2180_), .A2(new_n2182_), .ZN(new_n2183_));
  NAND4_X1   g02119(.A1(new_n2177_), .A2(new_n2170_), .A3(new_n2174_), .A4(new_n2183_), .ZN(new_n2184_));
  NOR2_X1    g02120(.A1(new_n617_), .A2(new_n1985_), .ZN(new_n2185_));
  NOR4_X1    g02121(.A1(new_n1198_), .A2(new_n81_), .A3(new_n117_), .A4(new_n607_), .ZN(new_n2186_));
  NAND4_X1   g02122(.A1(new_n2186_), .A2(new_n2185_), .A3(new_n1814_), .A4(new_n1804_), .ZN(new_n2187_));
  NOR3_X1    g02123(.A1(new_n753_), .A2(new_n902_), .A3(new_n306_), .ZN(new_n2188_));
  NAND4_X1   g02124(.A1(new_n480_), .A2(new_n1067_), .A3(new_n1662_), .A4(new_n144_), .ZN(new_n2189_));
  NAND3_X1   g02125(.A1(new_n1344_), .A2(new_n2189_), .A3(new_n2188_), .ZN(new_n2190_));
  NOR2_X1    g02126(.A1(new_n247_), .A2(new_n152_), .ZN(new_n2191_));
  NOR2_X1    g02127(.A1(new_n191_), .A2(new_n518_), .ZN(new_n2192_));
  INV_X1     g02128(.I(new_n2192_), .ZN(new_n2193_));
  NOR4_X1    g02129(.A1(new_n244_), .A2(new_n525_), .A3(new_n2193_), .A4(new_n689_), .ZN(new_n2194_));
  NAND4_X1   g02130(.A1(new_n2194_), .A2(new_n852_), .A3(new_n1044_), .A4(new_n2191_), .ZN(new_n2195_));
  NOR3_X1    g02131(.A1(new_n2187_), .A2(new_n2195_), .A3(new_n2190_), .ZN(new_n2196_));
  NAND2_X1   g02132(.A1(new_n2196_), .A2(new_n1581_), .ZN(new_n2197_));
  NOR2_X1    g02133(.A1(new_n2197_), .A2(new_n2184_), .ZN(new_n2198_));
  NOR2_X1    g02134(.A1(new_n2158_), .A2(new_n2198_), .ZN(new_n2199_));
  INV_X1     g02135(.I(new_n2199_), .ZN(new_n2200_));
  OAI21_X1   g02136(.A1(new_n2160_), .A2(new_n2162_), .B(new_n2200_), .ZN(new_n2201_));
  INV_X1     g02137(.I(new_n2198_), .ZN(new_n2202_));
  NOR2_X1    g02138(.A1(new_n2161_), .A2(new_n2202_), .ZN(new_n2203_));
  INV_X1     g02139(.I(new_n2203_), .ZN(new_n2204_));
  NOR2_X1    g02140(.A1(new_n1503_), .A2(new_n2198_), .ZN(new_n2205_));
  AOI21_X1   g02141(.A1(new_n2201_), .A2(new_n2204_), .B(new_n2205_), .ZN(new_n2206_));
  NOR2_X1    g02142(.A1(new_n1504_), .A2(new_n2202_), .ZN(new_n2207_));
  NAND2_X1   g02143(.A1(new_n331_), .A2(new_n1889_), .ZN(new_n2208_));
  NAND4_X1   g02144(.A1(new_n1489_), .A2(new_n362_), .A3(new_n808_), .A4(new_n274_), .ZN(new_n2209_));
  NAND4_X1   g02145(.A1(new_n2209_), .A2(new_n1105_), .A3(new_n677_), .A4(new_n1325_), .ZN(new_n2210_));
  NOR4_X1    g02146(.A1(new_n2210_), .A2(new_n1161_), .A3(new_n1632_), .A4(new_n2208_), .ZN(new_n2211_));
  INV_X1     g02147(.I(new_n2211_), .ZN(new_n2212_));
  INV_X1     g02148(.I(new_n713_), .ZN(new_n2213_));
  NAND4_X1   g02149(.A1(new_n199_), .A2(new_n1222_), .A3(new_n1753_), .A4(new_n1070_), .ZN(new_n2214_));
  NOR4_X1    g02150(.A1(new_n154_), .A2(new_n170_), .A3(new_n306_), .A4(new_n397_), .ZN(new_n2215_));
  NAND4_X1   g02151(.A1(new_n2214_), .A2(new_n2213_), .A3(new_n2192_), .A4(new_n2215_), .ZN(new_n2216_));
  NOR4_X1    g02152(.A1(new_n644_), .A2(new_n106_), .A3(new_n403_), .A4(new_n804_), .ZN(new_n2217_));
  NOR3_X1    g02153(.A1(new_n2217_), .A2(new_n558_), .A3(new_n1627_), .ZN(new_n2218_));
  NOR2_X1    g02154(.A1(new_n515_), .A2(new_n1138_), .ZN(new_n2219_));
  NAND4_X1   g02155(.A1(new_n2218_), .A2(new_n967_), .A3(new_n1075_), .A4(new_n2219_), .ZN(new_n2220_));
  NOR3_X1    g02156(.A1(new_n2212_), .A2(new_n2216_), .A3(new_n2220_), .ZN(new_n2221_));
  NAND3_X1   g02157(.A1(new_n2221_), .A2(new_n992_), .A3(new_n1335_), .ZN(new_n2222_));
  NOR4_X1    g02158(.A1(new_n119_), .A2(new_n202_), .A3(new_n611_), .A4(new_n594_), .ZN(new_n2223_));
  NOR4_X1    g02159(.A1(new_n324_), .A2(new_n398_), .A3(new_n753_), .A4(new_n772_), .ZN(new_n2224_));
  NOR3_X1    g02160(.A1(new_n2223_), .A2(new_n2224_), .A3(new_n1917_), .ZN(new_n2225_));
  NOR4_X1    g02161(.A1(new_n2176_), .A2(new_n132_), .A3(new_n573_), .A4(new_n261_), .ZN(new_n2226_));
  NOR4_X1    g02162(.A1(new_n1014_), .A2(new_n1391_), .A3(new_n995_), .A4(new_n565_), .ZN(new_n2227_));
  NAND4_X1   g02163(.A1(new_n2227_), .A2(new_n1528_), .A3(new_n2226_), .A4(new_n2225_), .ZN(new_n2228_));
  INV_X1     g02164(.I(new_n2228_), .ZN(new_n2229_));
  NOR4_X1    g02165(.A1(new_n615_), .A2(new_n190_), .A3(new_n577_), .A4(new_n776_), .ZN(new_n2230_));
  NOR3_X1    g02166(.A1(new_n2230_), .A2(new_n590_), .A3(new_n447_), .ZN(new_n2231_));
  INV_X1     g02167(.I(new_n1002_), .ZN(new_n2232_));
  NOR2_X1    g02168(.A1(new_n242_), .A2(new_n744_), .ZN(new_n2233_));
  INV_X1     g02169(.I(new_n2233_), .ZN(new_n2234_));
  NOR4_X1    g02170(.A1(new_n767_), .A2(new_n2232_), .A3(new_n1103_), .A4(new_n2234_), .ZN(new_n2235_));
  NOR2_X1    g02171(.A1(new_n453_), .A2(new_n262_), .ZN(new_n2236_));
  NOR2_X1    g02172(.A1(new_n2149_), .A2(new_n1784_), .ZN(new_n2237_));
  NAND3_X1   g02173(.A1(new_n2237_), .A2(new_n1358_), .A3(new_n2236_), .ZN(new_n2238_));
  NAND4_X1   g02174(.A1(new_n184_), .A2(new_n295_), .A3(new_n385_), .A4(new_n436_), .ZN(new_n2239_));
  INV_X1     g02175(.I(new_n297_), .ZN(new_n2240_));
  NAND4_X1   g02176(.A1(new_n2240_), .A2(new_n843_), .A3(new_n1935_), .A4(new_n809_), .ZN(new_n2241_));
  NOR3_X1    g02177(.A1(new_n2238_), .A2(new_n2239_), .A3(new_n2241_), .ZN(new_n2242_));
  INV_X1     g02178(.I(new_n2242_), .ZN(new_n2243_));
  INV_X1     g02179(.I(new_n697_), .ZN(new_n2244_));
  NOR2_X1    g02180(.A1(new_n732_), .A2(new_n430_), .ZN(new_n2245_));
  NAND4_X1   g02181(.A1(new_n688_), .A2(new_n1440_), .A3(new_n2244_), .A4(new_n2245_), .ZN(new_n2246_));
  NOR4_X1    g02182(.A1(new_n102_), .A2(new_n217_), .A3(new_n715_), .A4(new_n718_), .ZN(new_n2247_));
  NAND3_X1   g02183(.A1(new_n287_), .A2(new_n197_), .A3(new_n208_), .ZN(new_n2248_));
  NOR4_X1    g02184(.A1(new_n2243_), .A2(new_n2246_), .A3(new_n2247_), .A4(new_n2248_), .ZN(new_n2249_));
  NAND4_X1   g02185(.A1(new_n2249_), .A2(new_n2229_), .A3(new_n2231_), .A4(new_n2235_), .ZN(new_n2250_));
  NOR2_X1    g02186(.A1(new_n2250_), .A2(new_n2222_), .ZN(new_n2251_));
  NOR3_X1    g02187(.A1(new_n2206_), .A2(new_n2207_), .A3(new_n2251_), .ZN(new_n2252_));
  OAI21_X1   g02188(.A1(new_n2252_), .A2(new_n1547_), .B(new_n1504_), .ZN(new_n2253_));
  NOR2_X1    g02189(.A1(new_n2206_), .A2(new_n2207_), .ZN(new_n2254_));
  INV_X1     g02190(.I(new_n2251_), .ZN(new_n2255_));
  OAI21_X1   g02191(.A1(new_n2254_), .A2(new_n2255_), .B(new_n1547_), .ZN(new_n2256_));
  NOR4_X1    g02192(.A1(new_n2098_), .A2(new_n1200_), .A3(new_n1175_), .A4(new_n388_), .ZN(new_n2257_));
  NAND4_X1   g02193(.A1(new_n393_), .A2(new_n1605_), .A3(new_n1009_), .A4(new_n1325_), .ZN(new_n2258_));
  INV_X1     g02194(.I(new_n1430_), .ZN(new_n2259_));
  NOR2_X1    g02195(.A1(new_n343_), .A2(new_n752_), .ZN(new_n2260_));
  NAND2_X1   g02196(.A1(new_n2260_), .A2(new_n80_), .ZN(new_n2261_));
  NOR2_X1    g02197(.A1(new_n2259_), .A2(new_n2261_), .ZN(new_n2262_));
  NAND4_X1   g02198(.A1(new_n2262_), .A2(new_n1093_), .A3(new_n2257_), .A4(new_n2258_), .ZN(new_n2263_));
  INV_X1     g02199(.I(new_n2263_), .ZN(new_n2264_));
  NOR3_X1    g02200(.A1(new_n328_), .A2(new_n92_), .A3(new_n365_), .ZN(new_n2265_));
  NOR4_X1    g02201(.A1(new_n837_), .A2(new_n487_), .A3(new_n715_), .A4(new_n594_), .ZN(new_n2266_));
  INV_X1     g02202(.I(new_n2266_), .ZN(new_n2267_));
  NAND3_X1   g02203(.A1(new_n2265_), .A2(new_n1521_), .A3(new_n2267_), .ZN(new_n2268_));
  NOR2_X1    g02204(.A1(new_n689_), .A2(new_n1073_), .ZN(new_n2269_));
  INV_X1     g02205(.I(new_n2269_), .ZN(new_n2270_));
  NAND2_X1   g02206(.A1(new_n1599_), .A2(new_n1690_), .ZN(new_n2271_));
  NOR4_X1    g02207(.A1(new_n2268_), .A2(new_n1574_), .A3(new_n2270_), .A4(new_n2271_), .ZN(new_n2272_));
  AND3_X2    g02208(.A1(new_n2272_), .A2(new_n427_), .A3(new_n2264_), .Z(new_n2273_));
  INV_X1     g02209(.I(new_n1995_), .ZN(new_n2274_));
  NOR2_X1    g02210(.A1(new_n345_), .A2(new_n506_), .ZN(new_n2275_));
  NAND3_X1   g02211(.A1(new_n1288_), .A2(new_n2274_), .A3(new_n2275_), .ZN(new_n2276_));
  NOR4_X1    g02212(.A1(new_n656_), .A2(new_n102_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n2277_));
  NAND2_X1   g02213(.A1(new_n922_), .A2(new_n222_), .ZN(new_n2278_));
  NOR4_X1    g02214(.A1(new_n2276_), .A2(new_n560_), .A3(new_n2277_), .A4(new_n2278_), .ZN(new_n2279_));
  NAND2_X1   g02215(.A1(new_n2273_), .A2(new_n2279_), .ZN(new_n2280_));
  INV_X1     g02216(.I(new_n2280_), .ZN(new_n2281_));
  INV_X1     g02217(.I(new_n285_), .ZN(new_n2282_));
  NOR2_X1    g02218(.A1(new_n867_), .A2(new_n124_), .ZN(new_n2283_));
  INV_X1     g02219(.I(new_n2283_), .ZN(new_n2284_));
  NOR4_X1    g02220(.A1(new_n2284_), .A2(new_n1400_), .A3(new_n333_), .A4(new_n841_), .ZN(new_n2285_));
  OR3_X2     g02221(.A1(new_n1539_), .A2(new_n217_), .A3(new_n906_), .Z(new_n2286_));
  NAND4_X1   g02222(.A1(new_n480_), .A2(new_n1530_), .A3(new_n1448_), .A4(new_n665_), .ZN(new_n2287_));
  NAND3_X1   g02223(.A1(new_n2285_), .A2(new_n2286_), .A3(new_n2287_), .ZN(new_n2288_));
  NOR4_X1    g02224(.A1(new_n898_), .A2(new_n648_), .A3(new_n670_), .A4(new_n753_), .ZN(new_n2289_));
  NOR2_X1    g02225(.A1(new_n312_), .A2(new_n549_), .ZN(new_n2290_));
  INV_X1     g02226(.I(new_n2290_), .ZN(new_n2291_));
  NOR4_X1    g02227(.A1(new_n2291_), .A2(new_n297_), .A3(new_n556_), .A4(new_n930_), .ZN(new_n2292_));
  NOR2_X1    g02228(.A1(new_n1043_), .A2(new_n600_), .ZN(new_n2293_));
  NOR2_X1    g02229(.A1(new_n446_), .A2(new_n374_), .ZN(new_n2294_));
  NAND4_X1   g02230(.A1(new_n2292_), .A2(new_n1810_), .A3(new_n2293_), .A4(new_n2294_), .ZN(new_n2295_));
  NOR4_X1    g02231(.A1(new_n2295_), .A2(new_n2282_), .A3(new_n2288_), .A4(new_n2289_), .ZN(new_n2296_));
  NOR3_X1    g02232(.A1(new_n498_), .A2(new_n638_), .A3(new_n764_), .ZN(new_n2297_));
  NOR2_X1    g02233(.A1(new_n403_), .A2(new_n298_), .ZN(new_n2298_));
  NAND4_X1   g02234(.A1(new_n2297_), .A2(new_n1303_), .A3(new_n2298_), .A4(new_n1095_), .ZN(new_n2299_));
  NOR3_X1    g02235(.A1(new_n289_), .A2(new_n307_), .A3(new_n437_), .ZN(new_n2300_));
  NOR4_X1    g02236(.A1(new_n740_), .A2(new_n282_), .A3(new_n553_), .A4(new_n163_), .ZN(new_n2301_));
  NAND4_X1   g02237(.A1(new_n479_), .A2(new_n1829_), .A3(new_n394_), .A4(new_n441_), .ZN(new_n2302_));
  NAND4_X1   g02238(.A1(new_n2019_), .A2(new_n2300_), .A3(new_n2301_), .A4(new_n2302_), .ZN(new_n2303_));
  NAND4_X1   g02239(.A1(new_n469_), .A2(new_n1706_), .A3(new_n502_), .A4(new_n1396_), .ZN(new_n2304_));
  NAND2_X1   g02240(.A1(new_n2304_), .A2(new_n2236_), .ZN(new_n2305_));
  NOR2_X1    g02241(.A1(new_n1531_), .A2(new_n944_), .ZN(new_n2306_));
  INV_X1     g02242(.I(new_n2306_), .ZN(new_n2307_));
  NAND3_X1   g02243(.A1(new_n775_), .A2(new_n2307_), .A3(new_n537_), .ZN(new_n2308_));
  NOR4_X1    g02244(.A1(new_n2303_), .A2(new_n2299_), .A3(new_n2305_), .A4(new_n2308_), .ZN(new_n2309_));
  NAND3_X1   g02245(.A1(new_n2281_), .A2(new_n2296_), .A3(new_n2309_), .ZN(new_n2310_));
  INV_X1     g02246(.I(new_n2310_), .ZN(new_n2311_));
  NOR2_X1    g02247(.A1(new_n2311_), .A2(new_n2251_), .ZN(new_n2312_));
  INV_X1     g02248(.I(new_n2312_), .ZN(new_n2313_));
  NAND3_X1   g02249(.A1(new_n2253_), .A2(new_n2256_), .A3(new_n2313_), .ZN(new_n2314_));
  NOR2_X1    g02250(.A1(new_n2255_), .A2(new_n2310_), .ZN(new_n2315_));
  INV_X1     g02251(.I(new_n2315_), .ZN(new_n2316_));
  NOR4_X1    g02252(.A1(new_n788_), .A2(new_n252_), .A3(new_n654_), .A4(new_n163_), .ZN(new_n2317_));
  NOR4_X1    g02253(.A1(new_n644_), .A2(new_n226_), .A3(new_n906_), .A4(new_n1152_), .ZN(new_n2318_));
  INV_X1     g02254(.I(new_n2318_), .ZN(new_n2319_));
  NOR3_X1    g02255(.A1(new_n2319_), .A2(new_n891_), .A3(new_n2317_), .ZN(new_n2320_));
  NAND2_X1   g02256(.A1(new_n627_), .A2(new_n301_), .ZN(new_n2321_));
  NOR2_X1    g02257(.A1(new_n388_), .A2(new_n1168_), .ZN(new_n2322_));
  INV_X1     g02258(.I(new_n2322_), .ZN(new_n2323_));
  NOR4_X1    g02259(.A1(new_n2323_), .A2(new_n682_), .A3(new_n1915_), .A4(new_n2321_), .ZN(new_n2324_));
  NOR4_X1    g02260(.A1(new_n946_), .A2(new_n268_), .A3(new_n741_), .A4(new_n1092_), .ZN(new_n2325_));
  NOR2_X1    g02261(.A1(new_n648_), .A2(new_n345_), .ZN(new_n2326_));
  AOI21_X1   g02262(.A1(new_n588_), .A2(new_n2326_), .B(new_n2325_), .ZN(new_n2327_));
  INV_X1     g02263(.I(new_n930_), .ZN(new_n2328_));
  NOR2_X1    g02264(.A1(new_n137_), .A2(new_n1236_), .ZN(new_n2329_));
  NAND4_X1   g02265(.A1(new_n2329_), .A2(new_n199_), .A3(new_n2328_), .A4(new_n362_), .ZN(new_n2330_));
  NOR4_X1    g02266(.A1(new_n147_), .A2(new_n298_), .A3(new_n910_), .A4(new_n736_), .ZN(new_n2331_));
  NOR2_X1    g02267(.A1(new_n135_), .A2(new_n213_), .ZN(new_n2332_));
  INV_X1     g02268(.I(new_n2332_), .ZN(new_n2333_));
  NOR3_X1    g02269(.A1(new_n2330_), .A2(new_n2331_), .A3(new_n2333_), .ZN(new_n2334_));
  NAND4_X1   g02270(.A1(new_n2320_), .A2(new_n2324_), .A3(new_n2327_), .A4(new_n2334_), .ZN(new_n2335_));
  NOR4_X1    g02271(.A1(new_n217_), .A2(new_n307_), .A3(new_n136_), .A4(new_n264_), .ZN(new_n2336_));
  NOR2_X1    g02272(.A1(new_n2336_), .A2(new_n1619_), .ZN(new_n2337_));
  INV_X1     g02273(.I(new_n832_), .ZN(new_n2338_));
  NOR2_X1    g02274(.A1(new_n2338_), .A2(new_n225_), .ZN(new_n2339_));
  NOR2_X1    g02275(.A1(new_n1486_), .A2(new_n822_), .ZN(new_n2340_));
  NOR2_X1    g02276(.A1(new_n867_), .A2(new_n329_), .ZN(new_n2341_));
  INV_X1     g02277(.I(new_n2341_), .ZN(new_n2342_));
  NOR4_X1    g02278(.A1(new_n939_), .A2(new_n1511_), .A3(new_n337_), .A4(new_n2342_), .ZN(new_n2343_));
  NAND4_X1   g02279(.A1(new_n2343_), .A2(new_n2337_), .A3(new_n2339_), .A4(new_n2340_), .ZN(new_n2344_));
  NOR3_X1    g02280(.A1(new_n1084_), .A2(new_n577_), .A3(new_n714_), .ZN(new_n2345_));
  NOR3_X1    g02281(.A1(new_n1243_), .A2(new_n132_), .A3(new_n235_), .ZN(new_n2346_));
  NAND4_X1   g02282(.A1(new_n311_), .A2(new_n390_), .A3(new_n665_), .A4(new_n414_), .ZN(new_n2347_));
  NAND4_X1   g02283(.A1(new_n2346_), .A2(new_n2129_), .A3(new_n2345_), .A4(new_n2347_), .ZN(new_n2348_));
  NOR3_X1    g02284(.A1(new_n1030_), .A2(new_n2344_), .A3(new_n2348_), .ZN(new_n2349_));
  NAND2_X1   g02285(.A1(new_n2349_), .A2(new_n2196_), .ZN(new_n2350_));
  NOR2_X1    g02286(.A1(new_n2350_), .A2(new_n2335_), .ZN(new_n2351_));
  NOR2_X1    g02287(.A1(new_n2311_), .A2(new_n2351_), .ZN(new_n2352_));
  AOI21_X1   g02288(.A1(new_n2314_), .A2(new_n2316_), .B(new_n2352_), .ZN(new_n2353_));
  INV_X1     g02289(.I(new_n2351_), .ZN(new_n2354_));
  NOR2_X1    g02290(.A1(new_n2310_), .A2(new_n2354_), .ZN(new_n2355_));
  NOR2_X1    g02291(.A1(new_n1453_), .A2(new_n2351_), .ZN(new_n2356_));
  INV_X1     g02292(.I(new_n2356_), .ZN(new_n2357_));
  OAI21_X1   g02293(.A1(new_n2353_), .A2(new_n2355_), .B(new_n2357_), .ZN(new_n2358_));
  INV_X1     g02294(.I(new_n1453_), .ZN(new_n2359_));
  NOR2_X1    g02295(.A1(new_n2359_), .A2(new_n2354_), .ZN(new_n2360_));
  INV_X1     g02296(.I(new_n2360_), .ZN(new_n2361_));
  NAND2_X1   g02297(.A1(new_n2358_), .A2(new_n2361_), .ZN(new_n2362_));
  AOI21_X1   g02298(.A1(new_n2362_), .A2(new_n1453_), .B(new_n1409_), .ZN(new_n2363_));
  OAI21_X1   g02299(.A1(new_n2363_), .A2(new_n1334_), .B(new_n1241_), .ZN(new_n2364_));
  OAI21_X1   g02300(.A1(new_n2362_), .A2(new_n1453_), .B(new_n1409_), .ZN(new_n2365_));
  NAND2_X1   g02301(.A1(new_n2365_), .A2(new_n1334_), .ZN(new_n2366_));
  INV_X1     g02302(.I(new_n1241_), .ZN(new_n2367_));
  NOR2_X1    g02303(.A1(new_n119_), .A2(new_n262_), .ZN(new_n2368_));
  NAND4_X1   g02304(.A1(new_n1263_), .A2(new_n2368_), .A3(new_n188_), .A4(new_n643_), .ZN(new_n2369_));
  NOR2_X1    g02305(.A1(new_n1420_), .A2(new_n731_), .ZN(new_n2370_));
  NAND4_X1   g02306(.A1(new_n913_), .A2(new_n442_), .A3(new_n309_), .A4(new_n807_), .ZN(new_n2371_));
  NAND4_X1   g02307(.A1(new_n233_), .A2(new_n353_), .A3(new_n1327_), .A4(new_n266_), .ZN(new_n2372_));
  NAND3_X1   g02308(.A1(new_n2370_), .A2(new_n2371_), .A3(new_n2372_), .ZN(new_n2373_));
  NOR2_X1    g02309(.A1(new_n2373_), .A2(new_n2369_), .ZN(new_n2374_));
  INV_X1     g02310(.I(new_n902_), .ZN(new_n2375_));
  NAND2_X1   g02311(.A1(new_n2375_), .A2(new_n1009_), .ZN(new_n2376_));
  NAND2_X1   g02312(.A1(new_n999_), .A2(new_n502_), .ZN(new_n2377_));
  NOR4_X1    g02313(.A1(new_n1774_), .A2(new_n2376_), .A3(new_n2377_), .A4(new_n603_), .ZN(new_n2378_));
  NOR4_X1    g02314(.A1(new_n117_), .A2(new_n183_), .A3(new_n374_), .A4(new_n280_), .ZN(new_n2379_));
  NOR3_X1    g02315(.A1(new_n684_), .A2(new_n190_), .A3(new_n749_), .ZN(new_n2380_));
  INV_X1     g02316(.I(new_n2275_), .ZN(new_n2381_));
  NOR2_X1    g02317(.A1(new_n2381_), .A2(new_n695_), .ZN(new_n2382_));
  NAND2_X1   g02318(.A1(new_n2382_), .A2(new_n2380_), .ZN(new_n2383_));
  NOR4_X1    g02319(.A1(new_n2383_), .A2(new_n191_), .A3(new_n1359_), .A4(new_n2379_), .ZN(new_n2384_));
  NAND4_X1   g02320(.A1(new_n2091_), .A2(new_n349_), .A3(new_n1706_), .A4(new_n1770_), .ZN(new_n2385_));
  NAND4_X1   g02321(.A1(new_n1321_), .A2(new_n1692_), .A3(new_n1126_), .A4(new_n1699_), .ZN(new_n2386_));
  NOR2_X1    g02322(.A1(new_n2386_), .A2(new_n2385_), .ZN(new_n2387_));
  NAND4_X1   g02323(.A1(new_n2374_), .A2(new_n2384_), .A3(new_n2378_), .A4(new_n2387_), .ZN(new_n2388_));
  INV_X1     g02324(.I(new_n2145_), .ZN(new_n2389_));
  NOR2_X1    g02325(.A1(new_n510_), .A2(new_n937_), .ZN(new_n2390_));
  NAND4_X1   g02326(.A1(new_n2390_), .A2(new_n1063_), .A3(new_n1585_), .A4(new_n1891_), .ZN(new_n2391_));
  NAND2_X1   g02327(.A1(new_n870_), .A2(new_n1336_), .ZN(new_n2392_));
  NOR4_X1    g02328(.A1(new_n2009_), .A2(new_n2389_), .A3(new_n2391_), .A4(new_n2392_), .ZN(new_n2393_));
  NOR3_X1    g02329(.A1(new_n615_), .A2(new_n304_), .A3(new_n227_), .ZN(new_n2394_));
  NOR2_X1    g02330(.A1(new_n779_), .A2(new_n216_), .ZN(new_n2395_));
  INV_X1     g02331(.I(new_n2395_), .ZN(new_n2396_));
  NOR3_X1    g02332(.A1(new_n2396_), .A2(new_n495_), .A3(new_n490_), .ZN(new_n2397_));
  NOR2_X1    g02333(.A1(new_n255_), .A2(new_n549_), .ZN(new_n2398_));
  NOR2_X1    g02334(.A1(new_n366_), .A2(new_n482_), .ZN(new_n2399_));
  NAND4_X1   g02335(.A1(new_n2397_), .A2(new_n2394_), .A3(new_n2398_), .A4(new_n2399_), .ZN(new_n2400_));
  NOR2_X1    g02336(.A1(new_n945_), .A2(new_n1355_), .ZN(new_n2401_));
  NAND3_X1   g02337(.A1(new_n2401_), .A2(new_n854_), .A3(new_n880_), .ZN(new_n2402_));
  NAND4_X1   g02338(.A1(new_n293_), .A2(new_n361_), .A3(new_n808_), .A4(new_n207_), .ZN(new_n2403_));
  NOR2_X1    g02339(.A1(new_n988_), .A2(new_n935_), .ZN(new_n2404_));
  NAND3_X1   g02340(.A1(new_n2402_), .A2(new_n2404_), .A3(new_n2403_), .ZN(new_n2405_));
  NOR2_X1    g02341(.A1(new_n2400_), .A2(new_n2405_), .ZN(new_n2406_));
  NAND4_X1   g02342(.A1(new_n1219_), .A2(new_n2406_), .A3(new_n1201_), .A4(new_n2393_), .ZN(new_n2407_));
  NOR2_X1    g02343(.A1(new_n2407_), .A2(new_n2388_), .ZN(new_n2408_));
  NOR2_X1    g02344(.A1(new_n2367_), .A2(new_n2408_), .ZN(new_n2409_));
  INV_X1     g02345(.I(new_n2409_), .ZN(new_n2410_));
  NAND3_X1   g02346(.A1(new_n2364_), .A2(new_n2366_), .A3(new_n2410_), .ZN(new_n2411_));
  INV_X1     g02347(.I(new_n2408_), .ZN(new_n2412_));
  NOR2_X1    g02348(.A1(new_n1241_), .A2(new_n2412_), .ZN(new_n2413_));
  INV_X1     g02349(.I(new_n2413_), .ZN(new_n2414_));
  NOR2_X1    g02350(.A1(new_n505_), .A2(new_n1236_), .ZN(new_n2415_));
  NOR3_X1    g02351(.A1(new_n565_), .A2(new_n490_), .A3(new_n531_), .ZN(new_n2416_));
  NAND4_X1   g02352(.A1(new_n2416_), .A2(new_n667_), .A3(new_n1227_), .A4(new_n2415_), .ZN(new_n2417_));
  INV_X1     g02353(.I(new_n2417_), .ZN(new_n2418_));
  NOR3_X1    g02354(.A1(new_n495_), .A2(new_n117_), .A3(new_n744_), .ZN(new_n2419_));
  INV_X1     g02355(.I(new_n2419_), .ZN(new_n2420_));
  NOR4_X1    g02356(.A1(new_n251_), .A2(new_n491_), .A3(new_n1138_), .A4(new_n90_), .ZN(new_n2421_));
  NAND2_X1   g02357(.A1(new_n295_), .A2(new_n360_), .ZN(new_n2422_));
  NOR4_X1    g02358(.A1(new_n2420_), .A2(new_n1755_), .A3(new_n2421_), .A4(new_n2422_), .ZN(new_n2423_));
  NOR4_X1    g02359(.A1(new_n958_), .A2(new_n891_), .A3(new_n1043_), .A4(new_n1875_), .ZN(new_n2424_));
  NOR4_X1    g02360(.A1(new_n647_), .A2(new_n936_), .A3(new_n316_), .A4(new_n1858_), .ZN(new_n2425_));
  NAND4_X1   g02361(.A1(new_n2418_), .A2(new_n2423_), .A3(new_n2424_), .A4(new_n2425_), .ZN(new_n2426_));
  NOR4_X1    g02362(.A1(new_n788_), .A2(new_n335_), .A3(new_n652_), .A4(new_n236_), .ZN(new_n2427_));
  NOR2_X1    g02363(.A1(new_n553_), .A2(new_n388_), .ZN(new_n2428_));
  INV_X1     g02364(.I(new_n2428_), .ZN(new_n2429_));
  NOR3_X1    g02365(.A1(new_n2427_), .A2(new_n2429_), .A3(new_n558_), .ZN(new_n2430_));
  INV_X1     g02366(.I(new_n2430_), .ZN(new_n2431_));
  NOR2_X1    g02367(.A1(new_n119_), .A2(new_n397_), .ZN(new_n2432_));
  NAND4_X1   g02368(.A1(new_n987_), .A2(new_n2245_), .A3(new_n2432_), .A4(new_n978_), .ZN(new_n2433_));
  NAND2_X1   g02369(.A1(new_n1472_), .A2(new_n126_), .ZN(new_n2434_));
  NOR4_X1    g02370(.A1(new_n2431_), .A2(new_n1730_), .A3(new_n2433_), .A4(new_n2434_), .ZN(new_n2435_));
  NOR4_X1    g02371(.A1(new_n326_), .A2(new_n648_), .A3(new_n770_), .A4(new_n482_), .ZN(new_n2436_));
  NOR2_X1    g02372(.A1(new_n602_), .A2(new_n955_), .ZN(new_n2437_));
  INV_X1     g02373(.I(new_n2437_), .ZN(new_n2438_));
  INV_X1     g02374(.I(new_n598_), .ZN(new_n2439_));
  NOR2_X1    g02375(.A1(new_n2439_), .A2(new_n751_), .ZN(new_n2440_));
  INV_X1     g02376(.I(new_n2440_), .ZN(new_n2441_));
  NOR3_X1    g02377(.A1(new_n2441_), .A2(new_n261_), .A3(new_n468_), .ZN(new_n2442_));
  NOR3_X1    g02378(.A1(new_n2442_), .A2(new_n2436_), .A3(new_n2438_), .ZN(new_n2443_));
  NOR2_X1    g02379(.A1(new_n486_), .A2(new_n654_), .ZN(new_n2444_));
  INV_X1     g02380(.I(new_n2444_), .ZN(new_n2445_));
  NOR2_X1    g02381(.A1(new_n2445_), .A2(new_n297_), .ZN(new_n2446_));
  INV_X1     g02382(.I(new_n2446_), .ZN(new_n2447_));
  NOR4_X1    g02383(.A1(new_n239_), .A2(new_n260_), .A3(new_n384_), .A4(new_n1167_), .ZN(new_n2448_));
  NOR3_X1    g02384(.A1(new_n2447_), .A2(new_n571_), .A3(new_n2448_), .ZN(new_n2449_));
  NAND4_X1   g02385(.A1(new_n1544_), .A2(new_n2435_), .A3(new_n2443_), .A4(new_n2449_), .ZN(new_n2450_));
  NOR2_X1    g02386(.A1(new_n2450_), .A2(new_n2426_), .ZN(new_n2451_));
  NOR2_X1    g02387(.A1(new_n2451_), .A2(new_n2408_), .ZN(new_n2452_));
  AOI21_X1   g02388(.A1(new_n2411_), .A2(new_n2414_), .B(new_n2452_), .ZN(new_n2453_));
  INV_X1     g02389(.I(new_n2451_), .ZN(new_n2454_));
  NOR2_X1    g02390(.A1(new_n2454_), .A2(new_n2412_), .ZN(new_n2455_));
  NOR2_X1    g02391(.A1(new_n593_), .A2(new_n359_), .ZN(new_n2456_));
  INV_X1     g02392(.I(new_n2456_), .ZN(new_n2457_));
  INV_X1     g02393(.I(new_n1730_), .ZN(new_n2458_));
  NAND2_X1   g02394(.A1(new_n2458_), .A2(new_n1958_), .ZN(new_n2459_));
  NAND4_X1   g02395(.A1(new_n987_), .A2(new_n1358_), .A3(new_n1002_), .A4(new_n819_), .ZN(new_n2460_));
  NOR4_X1    g02396(.A1(new_n2459_), .A2(new_n2457_), .A3(new_n2460_), .A4(new_n1094_), .ZN(new_n2461_));
  NAND3_X1   g02397(.A1(new_n1311_), .A2(new_n1216_), .A3(new_n311_), .ZN(new_n2462_));
  NOR3_X1    g02398(.A1(new_n1652_), .A2(new_n420_), .A3(new_n689_), .ZN(new_n2463_));
  NAND2_X1   g02399(.A1(new_n1628_), .A2(new_n1494_), .ZN(new_n2464_));
  NOR4_X1    g02400(.A1(new_n2463_), .A2(new_n804_), .A3(new_n2462_), .A4(new_n2464_), .ZN(new_n2465_));
  NOR4_X1    g02401(.A1(new_n343_), .A2(new_n866_), .A3(new_n2439_), .A4(new_n136_), .ZN(new_n2466_));
  NAND4_X1   g02402(.A1(new_n628_), .A2(new_n1403_), .A3(new_n1444_), .A4(new_n843_), .ZN(new_n2467_));
  NOR4_X1    g02403(.A1(new_n950_), .A2(new_n1750_), .A3(new_n2466_), .A4(new_n2467_), .ZN(new_n2468_));
  NAND3_X1   g02404(.A1(new_n2468_), .A2(new_n2461_), .A3(new_n2465_), .ZN(new_n2469_));
  INV_X1     g02405(.I(new_n1201_), .ZN(new_n2470_));
  NAND4_X1   g02406(.A1(new_n1506_), .A2(new_n1796_), .A3(new_n832_), .A4(new_n669_), .ZN(new_n2471_));
  NOR4_X1    g02407(.A1(new_n1175_), .A2(new_n460_), .A3(new_n670_), .A4(new_n413_), .ZN(new_n2472_));
  NOR4_X1    g02408(.A1(new_n267_), .A2(new_n217_), .A3(new_n510_), .A4(new_n587_), .ZN(new_n2473_));
  NOR2_X1    g02409(.A1(new_n2473_), .A2(new_n2472_), .ZN(new_n2474_));
  NAND4_X1   g02410(.A1(new_n2474_), .A2(new_n492_), .A3(new_n2154_), .A4(new_n2471_), .ZN(new_n2475_));
  NOR4_X1    g02411(.A1(new_n740_), .A2(new_n590_), .A3(new_n1146_), .A4(new_n1167_), .ZN(new_n2476_));
  NOR4_X1    g02412(.A1(new_n1498_), .A2(new_n261_), .A3(new_n304_), .A4(new_n2476_), .ZN(new_n2477_));
  NOR4_X1    g02413(.A1(new_n618_), .A2(new_n70_), .A3(new_n335_), .A4(new_n695_), .ZN(new_n2478_));
  NOR2_X1    g02414(.A1(new_n783_), .A2(new_n192_), .ZN(new_n2479_));
  INV_X1     g02415(.I(new_n2479_), .ZN(new_n2480_));
  NOR2_X1    g02416(.A1(new_n637_), .A2(new_n496_), .ZN(new_n2481_));
  INV_X1     g02417(.I(new_n2481_), .ZN(new_n2482_));
  NOR4_X1    g02418(.A1(new_n2482_), .A2(new_n2480_), .A3(new_n365_), .A4(new_n772_), .ZN(new_n2483_));
  NAND3_X1   g02419(.A1(new_n2477_), .A2(new_n2483_), .A3(new_n2478_), .ZN(new_n2484_));
  NOR3_X1    g02420(.A1(new_n939_), .A2(new_n135_), .A3(new_n264_), .ZN(new_n2485_));
  NOR2_X1    g02421(.A1(new_n1461_), .A2(new_n533_), .ZN(new_n2486_));
  NAND4_X1   g02422(.A1(new_n1960_), .A2(new_n221_), .A3(new_n250_), .A4(new_n824_), .ZN(new_n2487_));
  NOR4_X1    g02423(.A1(new_n255_), .A2(new_n553_), .A3(new_n430_), .A4(new_n329_), .ZN(new_n2488_));
  INV_X1     g02424(.I(new_n2488_), .ZN(new_n2489_));
  NAND4_X1   g02425(.A1(new_n2485_), .A2(new_n2486_), .A3(new_n2487_), .A4(new_n2489_), .ZN(new_n2490_));
  OR4_X2     g02426(.A1(new_n2470_), .A2(new_n2484_), .A3(new_n2475_), .A4(new_n2490_), .Z(new_n2491_));
  NOR2_X1    g02427(.A1(new_n2491_), .A2(new_n2469_), .ZN(new_n2492_));
  NOR2_X1    g02428(.A1(new_n2492_), .A2(new_n2451_), .ZN(new_n2493_));
  INV_X1     g02429(.I(new_n2493_), .ZN(new_n2494_));
  OAI21_X1   g02430(.A1(new_n2453_), .A2(new_n2455_), .B(new_n2494_), .ZN(new_n2495_));
  INV_X1     g02431(.I(new_n2492_), .ZN(new_n2496_));
  NOR2_X1    g02432(.A1(new_n2496_), .A2(new_n2454_), .ZN(new_n2497_));
  INV_X1     g02433(.I(new_n2497_), .ZN(new_n2498_));
  NOR2_X1    g02434(.A1(new_n1121_), .A2(new_n2492_), .ZN(new_n2499_));
  AOI21_X1   g02435(.A1(new_n2495_), .A2(new_n2498_), .B(new_n2499_), .ZN(new_n2500_));
  NOR2_X1    g02436(.A1(new_n1122_), .A2(new_n2496_), .ZN(new_n2501_));
  NOR3_X1    g02437(.A1(new_n2500_), .A2(new_n1008_), .A3(new_n2501_), .ZN(new_n2502_));
  OAI21_X1   g02438(.A1(new_n2502_), .A2(new_n1181_), .B(new_n1122_), .ZN(new_n2503_));
  INV_X1     g02439(.I(new_n1008_), .ZN(new_n2504_));
  NOR2_X1    g02440(.A1(new_n2500_), .A2(new_n2501_), .ZN(new_n2505_));
  OAI21_X1   g02441(.A1(new_n2505_), .A2(new_n2504_), .B(new_n1181_), .ZN(new_n2506_));
  AOI21_X1   g02442(.A1(new_n2503_), .A2(new_n2506_), .B(new_n1008_), .ZN(new_n2507_));
  OAI21_X1   g02443(.A1(new_n2507_), .A2(new_n897_), .B(new_n814_), .ZN(new_n2508_));
  NAND2_X1   g02444(.A1(new_n2503_), .A2(new_n2506_), .ZN(new_n2509_));
  OAI21_X1   g02445(.A1(new_n2509_), .A2(new_n2504_), .B(new_n897_), .ZN(new_n2510_));
  INV_X1     g02446(.I(new_n2013_), .ZN(new_n2511_));
  NOR2_X1    g02447(.A1(new_n2482_), .A2(new_n2511_), .ZN(new_n2512_));
  NOR4_X1    g02448(.A1(new_n117_), .A2(new_n192_), .A3(new_n804_), .A4(new_n574_), .ZN(new_n2513_));
  NAND3_X1   g02449(.A1(new_n457_), .A2(new_n628_), .A3(new_n934_), .ZN(new_n2514_));
  NOR4_X1    g02450(.A1(new_n2514_), .A2(new_n879_), .A3(new_n2137_), .A4(new_n2513_), .ZN(new_n2515_));
  NAND4_X1   g02451(.A1(new_n2515_), .A2(new_n1246_), .A3(new_n1256_), .A4(new_n2512_), .ZN(new_n2516_));
  NOR3_X1    g02452(.A1(new_n219_), .A2(new_n403_), .A3(new_n560_), .ZN(new_n2517_));
  NOR3_X1    g02453(.A1(new_n687_), .A2(new_n366_), .A3(new_n329_), .ZN(new_n2518_));
  NAND4_X1   g02454(.A1(new_n2518_), .A2(new_n780_), .A3(new_n1001_), .A4(new_n2517_), .ZN(new_n2519_));
  NOR3_X1    g02455(.A1(new_n2516_), .A2(new_n1171_), .A3(new_n2519_), .ZN(new_n2520_));
  NOR2_X1    g02456(.A1(new_n225_), .A2(new_n347_), .ZN(new_n2521_));
  NAND4_X1   g02457(.A1(new_n1575_), .A2(new_n2432_), .A3(new_n2521_), .A4(new_n655_), .ZN(new_n2522_));
  NAND3_X1   g02458(.A1(new_n1530_), .A2(new_n675_), .A3(new_n222_), .ZN(new_n2523_));
  NAND3_X1   g02459(.A1(new_n2437_), .A2(new_n1605_), .A3(new_n677_), .ZN(new_n2524_));
  NOR3_X1    g02460(.A1(new_n2522_), .A2(new_n2524_), .A3(new_n2523_), .ZN(new_n2525_));
  NAND2_X1   g02461(.A1(new_n2520_), .A2(new_n2525_), .ZN(new_n2526_));
  NOR2_X1    g02462(.A1(new_n413_), .A2(new_n718_), .ZN(new_n2527_));
  INV_X1     g02463(.I(new_n2527_), .ZN(new_n2528_));
  NOR4_X1    g02464(.A1(new_n1160_), .A2(new_n1145_), .A3(new_n2193_), .A4(new_n2445_), .ZN(new_n2529_));
  NOR2_X1    g02465(.A1(new_n238_), .A2(new_n453_), .ZN(new_n2530_));
  NOR4_X1    g02466(.A1(new_n424_), .A2(new_n90_), .A3(new_n305_), .A4(new_n841_), .ZN(new_n2531_));
  NAND4_X1   g02467(.A1(new_n2529_), .A2(new_n266_), .A3(new_n2530_), .A4(new_n2531_), .ZN(new_n2532_));
  NOR4_X1    g02468(.A1(new_n2532_), .A2(new_n988_), .A3(new_n1511_), .A4(new_n2528_), .ZN(new_n2533_));
  INV_X1     g02469(.I(new_n2533_), .ZN(new_n2534_));
  NOR4_X1    g02470(.A1(new_n1116_), .A2(new_n1664_), .A3(new_n125_), .A4(new_n1236_), .ZN(new_n2535_));
  NAND4_X1   g02471(.A1(new_n2535_), .A2(new_n627_), .A3(new_n1063_), .A4(new_n442_), .ZN(new_n2536_));
  INV_X1     g02472(.I(new_n2536_), .ZN(new_n2537_));
  NOR4_X1    g02473(.A1(new_n465_), .A2(new_n235_), .A3(new_n763_), .A4(new_n320_), .ZN(new_n2538_));
  INV_X1     g02474(.I(new_n2538_), .ZN(new_n2539_));
  NOR3_X1    g02475(.A1(new_n936_), .A2(new_n365_), .A3(new_n447_), .ZN(new_n2540_));
  NAND4_X1   g02476(.A1(new_n2537_), .A2(new_n1047_), .A3(new_n2539_), .A4(new_n2540_), .ZN(new_n2541_));
  NOR2_X1    g02477(.A1(new_n2534_), .A2(new_n2541_), .ZN(new_n2542_));
  INV_X1     g02478(.I(new_n1534_), .ZN(new_n2543_));
  NOR2_X1    g02479(.A1(new_n960_), .A2(new_n1243_), .ZN(new_n2544_));
  INV_X1     g02480(.I(new_n2544_), .ZN(new_n2545_));
  NAND3_X1   g02481(.A1(new_n360_), .A2(new_n1454_), .A3(new_n669_), .ZN(new_n2546_));
  NOR3_X1    g02482(.A1(new_n774_), .A2(new_n1944_), .A3(new_n1146_), .ZN(new_n2547_));
  INV_X1     g02483(.I(new_n2547_), .ZN(new_n2548_));
  NOR4_X1    g02484(.A1(new_n2543_), .A2(new_n2545_), .A3(new_n2546_), .A4(new_n2548_), .ZN(new_n2549_));
  NAND3_X1   g02485(.A1(new_n1311_), .A2(new_n188_), .A3(new_n356_), .ZN(new_n2550_));
  NAND2_X1   g02486(.A1(new_n319_), .A2(new_n880_), .ZN(new_n2551_));
  NOR4_X1    g02487(.A1(new_n2550_), .A2(new_n213_), .A3(new_n2551_), .A4(new_n553_), .ZN(new_n2552_));
  INV_X1     g02488(.I(new_n1161_), .ZN(new_n2553_));
  NOR2_X1    g02489(.A1(new_n714_), .A2(new_n603_), .ZN(new_n2554_));
  NAND4_X1   g02490(.A1(new_n2553_), .A2(new_n539_), .A3(new_n2191_), .A4(new_n2554_), .ZN(new_n2555_));
  NAND3_X1   g02491(.A1(new_n276_), .A2(new_n808_), .A3(new_n1638_), .ZN(new_n2556_));
  NOR3_X1    g02492(.A1(new_n2555_), .A2(new_n917_), .A3(new_n2556_), .ZN(new_n2557_));
  NAND4_X1   g02493(.A1(new_n2542_), .A2(new_n2549_), .A3(new_n2552_), .A4(new_n2557_), .ZN(new_n2558_));
  NOR2_X1    g02494(.A1(new_n2558_), .A2(new_n2526_), .ZN(new_n2559_));
  NOR2_X1    g02495(.A1(new_n2559_), .A2(new_n813_), .ZN(new_n2560_));
  INV_X1     g02496(.I(new_n2560_), .ZN(new_n2561_));
  NAND3_X1   g02497(.A1(new_n2508_), .A2(new_n2510_), .A3(new_n2561_), .ZN(new_n2562_));
  INV_X1     g02498(.I(new_n2559_), .ZN(new_n2563_));
  NOR2_X1    g02499(.A1(new_n2563_), .A2(new_n814_), .ZN(new_n2564_));
  INV_X1     g02500(.I(new_n2564_), .ZN(new_n2565_));
  NAND2_X1   g02501(.A1(new_n2562_), .A2(new_n2565_), .ZN(new_n2566_));
  INV_X1     g02502(.I(new_n529_), .ZN(new_n2567_));
  NAND2_X1   g02503(.A1(new_n2563_), .A2(new_n2567_), .ZN(new_n2568_));
  NAND2_X1   g02504(.A1(new_n2566_), .A2(new_n2568_), .ZN(new_n2569_));
  NOR2_X1    g02505(.A1(new_n2563_), .A2(new_n2567_), .ZN(new_n2570_));
  INV_X1     g02506(.I(new_n2570_), .ZN(new_n2571_));
  NOR3_X1    g02507(.A1(new_n106_), .A2(new_n170_), .A3(new_n152_), .ZN(new_n2572_));
  NAND4_X1   g02508(.A1(new_n2465_), .A2(new_n1489_), .A3(new_n1095_), .A4(new_n2572_), .ZN(new_n2573_));
  NAND4_X1   g02509(.A1(new_n1404_), .A2(new_n1829_), .A3(new_n572_), .A4(new_n1605_), .ZN(new_n2574_));
  NOR3_X1    g02510(.A1(new_n491_), .A2(new_n584_), .A3(new_n535_), .ZN(new_n2575_));
  NAND4_X1   g02511(.A1(new_n2574_), .A2(new_n1968_), .A3(new_n2575_), .A4(new_n2527_), .ZN(new_n2576_));
  NOR4_X1    g02512(.A1(new_n495_), .A2(new_n485_), .A3(new_n1035_), .A4(new_n376_), .ZN(new_n2577_));
  NOR4_X1    g02513(.A1(new_n2577_), .A2(new_n387_), .A3(new_n906_), .A4(new_n510_), .ZN(new_n2578_));
  INV_X1     g02514(.I(new_n2578_), .ZN(new_n2579_));
  NOR4_X1    g02515(.A1(new_n132_), .A2(new_n262_), .A3(new_n732_), .A4(new_n1092_), .ZN(new_n2580_));
  NOR4_X1    g02516(.A1(new_n2580_), .A2(new_n70_), .A3(new_n459_), .A4(new_n1627_), .ZN(new_n2581_));
  INV_X1     g02517(.I(new_n1399_), .ZN(new_n2582_));
  NOR2_X1    g02518(.A1(new_n2582_), .A2(new_n544_), .ZN(new_n2583_));
  NAND4_X1   g02519(.A1(new_n2581_), .A2(new_n2583_), .A3(new_n641_), .A4(new_n1001_), .ZN(new_n2584_));
  NOR4_X1    g02520(.A1(new_n2573_), .A2(new_n2576_), .A3(new_n2584_), .A4(new_n2579_), .ZN(new_n2585_));
  INV_X1     g02521(.I(new_n1740_), .ZN(new_n2586_));
  NOR2_X1    g02522(.A1(new_n2438_), .A2(new_n487_), .ZN(new_n2587_));
  NOR2_X1    g02523(.A1(new_n531_), .A2(new_n719_), .ZN(new_n2588_));
  NAND4_X1   g02524(.A1(new_n2587_), .A2(new_n775_), .A3(new_n1375_), .A4(new_n2588_), .ZN(new_n2589_));
  NOR4_X1    g02525(.A1(new_n740_), .A2(new_n236_), .A3(new_n1262_), .A4(new_n577_), .ZN(new_n2590_));
  NOR2_X1    g02526(.A1(new_n211_), .A2(new_n1167_), .ZN(new_n2591_));
  NAND3_X1   g02527(.A1(new_n2591_), .A2(new_n187_), .A3(new_n342_), .ZN(new_n2592_));
  NAND4_X1   g02528(.A1(new_n2590_), .A2(new_n2489_), .A3(new_n2592_), .A4(new_n2148_), .ZN(new_n2593_));
  NAND4_X1   g02529(.A1(new_n790_), .A2(new_n274_), .A3(new_n391_), .A4(new_n1538_), .ZN(new_n2594_));
  NOR4_X1    g02530(.A1(new_n2589_), .A2(new_n2586_), .A3(new_n2593_), .A4(new_n2594_), .ZN(new_n2595_));
  NAND2_X1   g02531(.A1(new_n2585_), .A2(new_n2595_), .ZN(new_n2596_));
  NOR2_X1    g02532(.A1(new_n763_), .A2(new_n714_), .ZN(new_n2597_));
  INV_X1     g02533(.I(new_n2597_), .ZN(new_n2598_));
  NOR3_X1    g02534(.A1(new_n2598_), .A2(new_n618_), .A3(new_n630_), .ZN(new_n2599_));
  NOR3_X1    g02535(.A1(new_n899_), .A2(new_n330_), .A3(new_n506_), .ZN(new_n2600_));
  INV_X1     g02536(.I(new_n2600_), .ZN(new_n2601_));
  NOR4_X1    g02537(.A1(new_n352_), .A2(new_n1531_), .A3(new_n684_), .A4(new_n741_), .ZN(new_n2602_));
  NOR4_X1    g02538(.A1(new_n948_), .A2(new_n1589_), .A3(new_n2601_), .A4(new_n2602_), .ZN(new_n2603_));
  NOR4_X1    g02539(.A1(new_n415_), .A2(new_n625_), .A3(new_n212_), .A4(new_n247_), .ZN(new_n2604_));
  NAND2_X1   g02540(.A1(new_n351_), .A2(new_n1325_), .ZN(new_n2605_));
  NAND2_X1   g02541(.A1(new_n1446_), .A2(new_n809_), .ZN(new_n2606_));
  NAND2_X1   g02542(.A1(new_n543_), .A2(new_n2606_), .ZN(new_n2607_));
  NOR4_X1    g02543(.A1(new_n2607_), .A2(new_n81_), .A3(new_n2604_), .A4(new_n2605_), .ZN(new_n2608_));
  NOR4_X1    g02544(.A1(new_n137_), .A2(new_n837_), .A3(new_n488_), .A4(new_n1146_), .ZN(new_n2609_));
  INV_X1     g02545(.I(new_n1656_), .ZN(new_n2610_));
  NAND4_X1   g02546(.A1(new_n2610_), .A2(new_n197_), .A3(new_n1590_), .A4(new_n707_), .ZN(new_n2611_));
  NOR2_X1    g02547(.A1(new_n2611_), .A2(new_n2609_), .ZN(new_n2612_));
  NAND4_X1   g02548(.A1(new_n2612_), .A2(new_n2603_), .A3(new_n2608_), .A4(new_n2599_), .ZN(new_n2613_));
  NOR2_X1    g02549(.A1(new_n2596_), .A2(new_n2613_), .ZN(new_n2614_));
  INV_X1     g02550(.I(new_n2614_), .ZN(new_n2615_));
  NAND3_X1   g02551(.A1(new_n2569_), .A2(new_n2571_), .A3(new_n2615_), .ZN(new_n2616_));
  AOI21_X1   g02552(.A1(new_n2616_), .A2(new_n694_), .B(new_n529_), .ZN(new_n2617_));
  NAND2_X1   g02553(.A1(new_n2569_), .A2(new_n2571_), .ZN(new_n2618_));
  AOI21_X1   g02554(.A1(new_n2618_), .A2(new_n2614_), .B(new_n694_), .ZN(new_n2619_));
  NOR2_X1    g02555(.A1(new_n232_), .A2(new_n741_), .ZN(new_n2620_));
  NAND3_X1   g02556(.A1(new_n2219_), .A2(new_n2620_), .A3(new_n1765_), .ZN(new_n2621_));
  NOR2_X1    g02557(.A1(new_n740_), .A2(new_n474_), .ZN(new_n2622_));
  NOR2_X1    g02558(.A1(new_n135_), .A2(new_n1152_), .ZN(new_n2623_));
  NOR2_X1    g02559(.A1(new_n817_), .A2(new_n1031_), .ZN(new_n2624_));
  NAND4_X1   g02560(.A1(new_n253_), .A2(new_n2622_), .A3(new_n2623_), .A4(new_n2624_), .ZN(new_n2625_));
  NOR4_X1    g02561(.A1(new_n837_), .A2(new_n944_), .A3(new_n397_), .A4(new_n329_), .ZN(new_n2626_));
  NOR4_X1    g02562(.A1(new_n225_), .A2(new_n297_), .A3(new_n305_), .A4(new_n682_), .ZN(new_n2627_));
  NOR4_X1    g02563(.A1(new_n2625_), .A2(new_n2621_), .A3(new_n2626_), .A4(new_n2627_), .ZN(new_n2628_));
  INV_X1     g02564(.I(new_n2628_), .ZN(new_n2629_));
  NOR2_X1    g02565(.A1(new_n2289_), .A2(new_n2282_), .ZN(new_n2630_));
  NAND2_X1   g02566(.A1(new_n1025_), .A2(new_n471_), .ZN(new_n2631_));
  NOR4_X1    g02567(.A1(new_n2631_), .A2(new_n149_), .A3(new_n2439_), .A4(new_n388_), .ZN(new_n2632_));
  NOR4_X1    g02568(.A1(new_n637_), .A2(new_n603_), .A3(new_n173_), .A4(new_n376_), .ZN(new_n2633_));
  NOR2_X1    g02569(.A1(new_n647_), .A2(new_n1011_), .ZN(new_n2634_));
  NAND4_X1   g02570(.A1(new_n2630_), .A2(new_n2632_), .A3(new_n2633_), .A4(new_n2634_), .ZN(new_n2635_));
  NOR4_X1    g02571(.A1(new_n130_), .A2(new_n304_), .A3(new_n447_), .A4(new_n324_), .ZN(new_n2636_));
  NOR4_X1    g02572(.A1(new_n2636_), .A2(new_n428_), .A3(new_n381_), .A4(new_n556_), .ZN(new_n2637_));
  NAND3_X1   g02573(.A1(new_n2637_), .A2(new_n1853_), .A3(new_n1689_), .ZN(new_n2638_));
  NAND4_X1   g02574(.A1(new_n1628_), .A2(new_n1091_), .A3(new_n1605_), .A4(new_n274_), .ZN(new_n2639_));
  NAND3_X1   g02575(.A1(new_n1021_), .A2(new_n662_), .A3(new_n1315_), .ZN(new_n2640_));
  NAND4_X1   g02576(.A1(new_n2640_), .A2(new_n1436_), .A3(new_n1968_), .A4(new_n2639_), .ZN(new_n2641_));
  NOR4_X1    g02577(.A1(new_n2629_), .A2(new_n2635_), .A3(new_n2638_), .A4(new_n2641_), .ZN(new_n2642_));
  NAND3_X1   g02578(.A1(new_n967_), .A2(new_n1767_), .A3(new_n631_), .ZN(new_n2643_));
  NOR2_X1    g02579(.A1(new_n582_), .A2(new_n359_), .ZN(new_n2644_));
  NAND4_X1   g02580(.A1(new_n545_), .A2(new_n2444_), .A3(new_n2644_), .A4(new_n1699_), .ZN(new_n2645_));
  NOR2_X1    g02581(.A1(new_n791_), .A2(new_n764_), .ZN(new_n2646_));
  INV_X1     g02582(.I(new_n2646_), .ZN(new_n2647_));
  NOR3_X1    g02583(.A1(new_n2647_), .A2(new_n226_), .A3(new_n1236_), .ZN(new_n2648_));
  NOR3_X1    g02584(.A1(new_n244_), .A2(new_n594_), .A3(new_n930_), .ZN(new_n2649_));
  INV_X1     g02585(.I(new_n2649_), .ZN(new_n2650_));
  NOR4_X1    g02586(.A1(new_n2650_), .A2(new_n2643_), .A3(new_n2645_), .A4(new_n2648_), .ZN(new_n2651_));
  NOR4_X1    g02587(.A1(new_n906_), .A2(new_n288_), .A3(new_n584_), .A4(new_n487_), .ZN(new_n2652_));
  NAND3_X1   g02588(.A1(new_n2652_), .A2(new_n554_), .A3(new_n1319_), .ZN(new_n2653_));
  NOR2_X1    g02589(.A1(new_n387_), .A2(new_n510_), .ZN(new_n2654_));
  NAND4_X1   g02590(.A1(new_n1349_), .A2(new_n187_), .A3(new_n2654_), .A4(new_n436_), .ZN(new_n2655_));
  NOR2_X1    g02591(.A1(new_n2653_), .A2(new_n2655_), .ZN(new_n2656_));
  INV_X1     g02592(.I(new_n1782_), .ZN(new_n2657_));
  NOR3_X1    g02593(.A1(new_n577_), .A2(new_n1035_), .A3(new_n731_), .ZN(new_n2658_));
  NOR3_X1    g02594(.A1(new_n1962_), .A2(new_n782_), .A3(new_n841_), .ZN(new_n2659_));
  NAND4_X1   g02595(.A1(new_n469_), .A2(new_n1088_), .A3(new_n655_), .A4(new_n394_), .ZN(new_n2660_));
  NAND4_X1   g02596(.A1(new_n2660_), .A2(new_n2657_), .A3(new_n2659_), .A4(new_n2658_), .ZN(new_n2661_));
  INV_X1     g02597(.I(new_n2661_), .ZN(new_n2662_));
  AND3_X2    g02598(.A1(new_n2651_), .A2(new_n2656_), .A3(new_n2662_), .Z(new_n2663_));
  NAND2_X1   g02599(.A1(new_n2663_), .A2(new_n2642_), .ZN(new_n2664_));
  INV_X1     g02600(.I(new_n2664_), .ZN(new_n2665_));
  NOR2_X1    g02601(.A1(new_n2614_), .A2(new_n2665_), .ZN(new_n2666_));
  NOR3_X1    g02602(.A1(new_n2617_), .A2(new_n2619_), .A3(new_n2666_), .ZN(new_n2667_));
  NOR2_X1    g02603(.A1(new_n2615_), .A2(new_n2664_), .ZN(new_n2668_));
  NOR2_X1    g02604(.A1(new_n2667_), .A2(new_n2668_), .ZN(new_n2669_));
  NOR3_X1    g02605(.A1(new_n337_), .A2(new_n227_), .A3(new_n384_), .ZN(new_n2670_));
  NOR2_X1    g02606(.A1(new_n1365_), .A2(new_n1954_), .ZN(new_n2671_));
  NAND4_X1   g02607(.A1(new_n2670_), .A2(new_n2671_), .A3(new_n1766_), .A4(new_n1781_), .ZN(new_n2672_));
  NOR4_X1    g02608(.A1(new_n495_), .A2(new_n190_), .A3(new_n420_), .A4(new_n475_), .ZN(new_n2673_));
  NOR4_X1    g02609(.A1(new_n1531_), .A2(new_n183_), .A3(new_n517_), .A4(new_n132_), .ZN(new_n2674_));
  NOR3_X1    g02610(.A1(new_n2673_), .A2(new_n1487_), .A3(new_n2674_), .ZN(new_n2675_));
  NOR2_X1    g02611(.A1(new_n236_), .A2(new_n419_), .ZN(new_n2676_));
  INV_X1     g02612(.I(new_n2676_), .ZN(new_n2677_));
  NOR4_X1    g02613(.A1(new_n406_), .A2(new_n163_), .A3(new_n255_), .A4(new_n286_), .ZN(new_n2678_));
  NOR4_X1    g02614(.A1(new_n2678_), .A2(new_n496_), .A3(new_n2677_), .A4(new_n541_), .ZN(new_n2679_));
  NAND3_X1   g02615(.A1(new_n792_), .A2(new_n913_), .A3(new_n797_), .ZN(new_n2680_));
  NAND4_X1   g02616(.A1(new_n2679_), .A2(new_n2675_), .A3(new_n947_), .A4(new_n2680_), .ZN(new_n2681_));
  NOR4_X1    g02617(.A1(new_n607_), .A2(new_n491_), .A3(new_n561_), .A4(new_n611_), .ZN(new_n2682_));
  INV_X1     g02618(.I(new_n2682_), .ZN(new_n2683_));
  NOR2_X1    g02619(.A1(new_n2149_), .A2(new_n763_), .ZN(new_n2684_));
  NAND4_X1   g02620(.A1(new_n2684_), .A2(new_n452_), .A3(new_n532_), .A4(new_n2683_), .ZN(new_n2685_));
  NOR3_X1    g02621(.A1(new_n2681_), .A2(new_n2685_), .A3(new_n2672_), .ZN(new_n2686_));
  NOR4_X1    g02622(.A1(new_n251_), .A2(new_n1084_), .A3(new_n670_), .A4(new_n352_), .ZN(new_n2687_));
  NOR3_X1    g02623(.A1(new_n2687_), .A2(new_n1152_), .A3(new_n779_), .ZN(new_n2688_));
  NOR4_X1    g02624(.A1(new_n226_), .A2(new_n388_), .A3(new_n817_), .A4(new_n1073_), .ZN(new_n2689_));
  INV_X1     g02625(.I(new_n2689_), .ZN(new_n2690_));
  NOR2_X1    g02626(.A1(new_n121_), .A2(new_n397_), .ZN(new_n2691_));
  NAND4_X1   g02627(.A1(new_n2688_), .A2(new_n2659_), .A3(new_n2690_), .A4(new_n2691_), .ZN(new_n2692_));
  NOR4_X1    g02628(.A1(new_n2692_), .A2(new_n2638_), .A3(new_n2653_), .A4(new_n2655_), .ZN(new_n2693_));
  NAND3_X1   g02629(.A1(new_n301_), .A2(new_n1662_), .A3(new_n222_), .ZN(new_n2694_));
  NOR4_X1    g02630(.A1(new_n2284_), .A2(new_n788_), .A3(new_n736_), .A4(new_n2694_), .ZN(new_n2695_));
  NAND2_X1   g02631(.A1(new_n2695_), .A2(new_n269_), .ZN(new_n2696_));
  INV_X1     g02632(.I(new_n2696_), .ZN(new_n2697_));
  NOR2_X1    g02633(.A1(new_n744_), .A2(new_n749_), .ZN(new_n2698_));
  NAND4_X1   g02634(.A1(new_n2693_), .A2(new_n2686_), .A3(new_n2697_), .A4(new_n2698_), .ZN(new_n2699_));
  NAND4_X1   g02635(.A1(new_n819_), .A2(new_n1930_), .A3(new_n319_), .A4(new_n432_), .ZN(new_n2700_));
  NOR2_X1    g02636(.A1(new_n2061_), .A2(new_n2700_), .ZN(new_n2701_));
  NOR2_X1    g02637(.A1(new_n2445_), .A2(new_n460_), .ZN(new_n2702_));
  INV_X1     g02638(.I(new_n1165_), .ZN(new_n2703_));
  INV_X1     g02639(.I(new_n1237_), .ZN(new_n2704_));
  NOR3_X1    g02640(.A1(new_n2703_), .A2(new_n2704_), .A3(new_n935_), .ZN(new_n2705_));
  AND4_X2    g02641(.A1(new_n2608_), .A2(new_n2701_), .A3(new_n2702_), .A4(new_n2705_), .Z(new_n2706_));
  NOR4_X1    g02642(.A1(new_n945_), .A2(new_n136_), .A3(new_n548_), .A4(new_n347_), .ZN(new_n2707_));
  NOR3_X1    g02643(.A1(new_n366_), .A2(new_n604_), .A3(new_n698_), .ZN(new_n2708_));
  INV_X1     g02644(.I(new_n2708_), .ZN(new_n2709_));
  NOR4_X1    g02645(.A1(new_n2709_), .A2(new_n2707_), .A3(new_n1157_), .A4(new_n1754_), .ZN(new_n2710_));
  INV_X1     g02646(.I(new_n2710_), .ZN(new_n2711_));
  NOR2_X1    g02647(.A1(new_n252_), .A2(new_n149_), .ZN(new_n2712_));
  NAND4_X1   g02648(.A1(new_n2712_), .A2(new_n992_), .A3(new_n1605_), .A4(new_n383_), .ZN(new_n2713_));
  NOR4_X1    g02649(.A1(new_n2711_), .A2(new_n1175_), .A3(new_n576_), .A4(new_n2713_), .ZN(new_n2714_));
  NAND2_X1   g02650(.A1(new_n2706_), .A2(new_n2714_), .ZN(new_n2715_));
  NOR2_X1    g02651(.A1(new_n2715_), .A2(new_n2699_), .ZN(new_n2716_));
  XOR2_X1    g02652(.A1(new_n2716_), .A2(new_n2664_), .Z(new_n2717_));
  INV_X1     g02653(.I(new_n694_), .ZN(new_n2718_));
  AOI22_X1   g02654(.A1(new_n2562_), .A2(new_n2565_), .B1(new_n2567_), .B2(new_n2563_), .ZN(new_n2719_));
  NOR3_X1    g02655(.A1(new_n2719_), .A2(new_n2570_), .A3(new_n2614_), .ZN(new_n2720_));
  OAI21_X1   g02656(.A1(new_n2720_), .A2(new_n2718_), .B(new_n2567_), .ZN(new_n2721_));
  NOR2_X1    g02657(.A1(new_n2719_), .A2(new_n2570_), .ZN(new_n2722_));
  OAI21_X1   g02658(.A1(new_n2722_), .A2(new_n2615_), .B(new_n2718_), .ZN(new_n2723_));
  INV_X1     g02659(.I(new_n2666_), .ZN(new_n2724_));
  NAND3_X1   g02660(.A1(new_n2721_), .A2(new_n2723_), .A3(new_n2724_), .ZN(new_n2725_));
  INV_X1     g02661(.I(new_n2668_), .ZN(new_n2726_));
  NOR2_X1    g02662(.A1(new_n2716_), .A2(new_n2665_), .ZN(new_n2727_));
  INV_X1     g02663(.I(new_n2716_), .ZN(new_n2728_));
  NOR2_X1    g02664(.A1(new_n2728_), .A2(new_n2664_), .ZN(new_n2729_));
  NOR2_X1    g02665(.A1(new_n2729_), .A2(new_n2727_), .ZN(new_n2730_));
  INV_X1     g02666(.I(new_n2730_), .ZN(new_n2731_));
  NAND3_X1   g02667(.A1(new_n2725_), .A2(new_n2726_), .A3(new_n2731_), .ZN(new_n2732_));
  OAI21_X1   g02668(.A1(new_n2669_), .A2(new_n2717_), .B(new_n2732_), .ZN(new_n2733_));
  XNOR2_X1   g02669(.A1(\a[26] ), .A2(\a[27] ), .ZN(new_n2734_));
  XNOR2_X1   g02670(.A1(\a[28] ), .A2(\a[29] ), .ZN(new_n2735_));
  NOR2_X1    g02671(.A1(new_n2735_), .A2(new_n2734_), .ZN(new_n2736_));
  INV_X1     g02672(.I(new_n2736_), .ZN(new_n2737_));
  NOR2_X1    g02673(.A1(new_n82_), .A2(\a[28] ), .ZN(new_n2738_));
  NAND2_X1   g02674(.A1(new_n2738_), .A2(\a[26] ), .ZN(new_n2739_));
  NOR2_X1    g02675(.A1(new_n67_), .A2(\a[27] ), .ZN(new_n2740_));
  NAND2_X1   g02676(.A1(new_n2740_), .A2(new_n72_), .ZN(new_n2741_));
  AND2_X2    g02677(.A1(new_n2739_), .A2(new_n2741_), .Z(new_n2742_));
  XNOR2_X1   g02678(.A1(\a[26] ), .A2(\a[28] ), .ZN(new_n2743_));
  NAND2_X1   g02679(.A1(new_n2734_), .A2(new_n2743_), .ZN(new_n2744_));
  XNOR2_X1   g02680(.A1(\a[26] ), .A2(\a[29] ), .ZN(new_n2745_));
  AND2_X2    g02681(.A1(new_n2744_), .A2(new_n2745_), .Z(new_n2746_));
  INV_X1     g02682(.I(new_n2746_), .ZN(new_n2747_));
  OAI22_X1   g02683(.A1(new_n2614_), .A2(new_n2747_), .B1(new_n2665_), .B2(new_n2742_), .ZN(new_n2748_));
  INV_X1     g02684(.I(new_n2734_), .ZN(new_n2749_));
  NOR2_X1    g02685(.A1(new_n2749_), .A2(new_n2735_), .ZN(new_n2750_));
  NAND2_X1   g02686(.A1(new_n2728_), .A2(new_n2750_), .ZN(new_n2751_));
  AOI21_X1   g02687(.A1(new_n2751_), .A2(new_n2748_), .B(new_n2737_), .ZN(new_n2752_));
  NAND2_X1   g02688(.A1(new_n2733_), .A2(new_n2752_), .ZN(new_n2753_));
  XOR2_X1    g02689(.A1(new_n2753_), .A2(\a[29] ), .Z(new_n2754_));
  XOR2_X1    g02690(.A1(new_n694_), .A2(new_n2567_), .Z(new_n2755_));
  XOR2_X1    g02691(.A1(new_n694_), .A2(new_n529_), .Z(new_n2756_));
  NOR3_X1    g02692(.A1(new_n2719_), .A2(new_n2570_), .A3(new_n2756_), .ZN(new_n2757_));
  INV_X1     g02693(.I(new_n2757_), .ZN(new_n2758_));
  OAI21_X1   g02694(.A1(new_n2722_), .A2(new_n2755_), .B(new_n2758_), .ZN(new_n2759_));
  NAND2_X1   g02695(.A1(new_n74_), .A2(\a[30] ), .ZN(new_n2760_));
  NAND2_X1   g02696(.A1(new_n68_), .A2(\a[29] ), .ZN(new_n2761_));
  NAND2_X1   g02697(.A1(new_n2760_), .A2(new_n2761_), .ZN(new_n2762_));
  NAND2_X1   g02698(.A1(new_n2762_), .A2(\a[31] ), .ZN(new_n2763_));
  INV_X1     g02699(.I(new_n2763_), .ZN(new_n2764_));
  NAND2_X1   g02700(.A1(\a[29] ), .A2(\a[30] ), .ZN(new_n2765_));
  NOR2_X1    g02701(.A1(new_n2765_), .A2(\a[31] ), .ZN(new_n2766_));
  AOI21_X1   g02702(.A1(\a[31] ), .A2(new_n354_), .B(new_n2766_), .ZN(new_n2767_));
  OAI21_X1   g02703(.A1(new_n529_), .A2(new_n2767_), .B(new_n2764_), .ZN(new_n2768_));
  INV_X1     g02704(.I(\a[31] ), .ZN(new_n2769_));
  NOR2_X1    g02705(.A1(new_n2765_), .A2(new_n2769_), .ZN(new_n2770_));
  INV_X1     g02706(.I(new_n2770_), .ZN(new_n2771_));
  NAND2_X1   g02707(.A1(new_n2762_), .A2(new_n2769_), .ZN(new_n2772_));
  OAI22_X1   g02708(.A1(new_n2559_), .A2(new_n2771_), .B1(new_n694_), .B2(new_n2772_), .ZN(new_n2773_));
  NOR2_X1    g02709(.A1(new_n2773_), .A2(new_n2768_), .ZN(new_n2774_));
  NAND2_X1   g02710(.A1(new_n2759_), .A2(new_n2774_), .ZN(new_n2775_));
  NOR3_X1    g02711(.A1(new_n2338_), .A2(new_n695_), .A3(new_n776_), .ZN(new_n2776_));
  INV_X1     g02712(.I(new_n2776_), .ZN(new_n2777_));
  NAND2_X1   g02713(.A1(new_n1403_), .A2(new_n221_), .ZN(new_n2778_));
  NOR4_X1    g02714(.A1(new_n81_), .A2(new_n782_), .A3(new_n487_), .A4(new_n715_), .ZN(new_n2779_));
  INV_X1     g02715(.I(new_n2779_), .ZN(new_n2780_));
  NOR3_X1    g02716(.A1(new_n898_), .A2(new_n232_), .A3(new_n418_), .ZN(new_n2781_));
  NAND2_X1   g02717(.A1(new_n2780_), .A2(new_n2781_), .ZN(new_n2782_));
  NOR4_X1    g02718(.A1(new_n2782_), .A2(new_n347_), .A3(new_n2777_), .A4(new_n2778_), .ZN(new_n2783_));
  NOR4_X1    g02719(.A1(new_n384_), .A2(new_n899_), .A3(new_n474_), .A4(new_n561_), .ZN(new_n2784_));
  NAND4_X1   g02720(.A1(new_n511_), .A2(new_n1666_), .A3(new_n302_), .A4(new_n1935_), .ZN(new_n2785_));
  NAND3_X1   g02721(.A1(new_n875_), .A2(new_n271_), .A3(new_n501_), .ZN(new_n2786_));
  NOR4_X1    g02722(.A1(new_n607_), .A2(new_n324_), .A3(new_n584_), .A4(new_n867_), .ZN(new_n2787_));
  NOR4_X1    g02723(.A1(new_n2787_), .A2(new_n172_), .A3(new_n573_), .A4(new_n604_), .ZN(new_n2788_));
  NAND4_X1   g02724(.A1(new_n2788_), .A2(new_n827_), .A3(new_n1329_), .A4(new_n1942_), .ZN(new_n2789_));
  NOR4_X1    g02725(.A1(new_n2789_), .A2(new_n2784_), .A3(new_n2785_), .A4(new_n2786_), .ZN(new_n2790_));
  NAND2_X1   g02726(.A1(new_n2790_), .A2(new_n2783_), .ZN(new_n2791_));
  NAND4_X1   g02727(.A1(new_n292_), .A2(new_n322_), .A3(new_n512_), .A4(new_n1070_), .ZN(new_n2792_));
  NAND4_X1   g02728(.A1(new_n248_), .A2(new_n442_), .A3(new_n1025_), .A4(new_n1436_), .ZN(new_n2793_));
  NAND2_X1   g02729(.A1(new_n2793_), .A2(new_n2792_), .ZN(new_n2794_));
  NOR2_X1    g02730(.A1(new_n76_), .A2(new_n286_), .ZN(new_n2795_));
  NOR4_X1    g02731(.A1(new_n563_), .A2(new_n1985_), .A3(new_n663_), .A4(new_n177_), .ZN(new_n2796_));
  NAND4_X1   g02732(.A1(new_n2796_), .A2(new_n852_), .A3(new_n1516_), .A4(new_n2795_), .ZN(new_n2797_));
  NOR4_X1    g02733(.A1(new_n611_), .A2(new_n783_), .A3(new_n610_), .A4(new_n163_), .ZN(new_n2798_));
  NOR2_X1    g02734(.A1(new_n929_), .A2(new_n2798_), .ZN(new_n2799_));
  NOR4_X1    g02735(.A1(new_n1355_), .A2(new_n191_), .A3(new_n268_), .A4(new_n282_), .ZN(new_n2800_));
  NOR2_X1    g02736(.A1(new_n505_), .A2(new_n260_), .ZN(new_n2801_));
  AOI21_X1   g02737(.A1(new_n2332_), .A2(new_n2801_), .B(new_n2800_), .ZN(new_n2802_));
  NAND4_X1   g02738(.A1(new_n438_), .A2(new_n672_), .A3(new_n984_), .A4(new_n222_), .ZN(new_n2803_));
  NAND4_X1   g02739(.A1(new_n612_), .A2(new_n2375_), .A3(new_n110_), .A4(new_n246_), .ZN(new_n2804_));
  NOR4_X1    g02740(.A1(new_n2804_), .A2(new_n2803_), .A3(new_n299_), .A4(new_n825_), .ZN(new_n2805_));
  NAND3_X1   g02741(.A1(new_n2805_), .A2(new_n2802_), .A3(new_n2799_), .ZN(new_n2806_));
  NOR4_X1    g02742(.A1(new_n2791_), .A2(new_n2794_), .A3(new_n2797_), .A4(new_n2806_), .ZN(new_n2807_));
  NAND2_X1   g02743(.A1(new_n2807_), .A2(new_n1428_), .ZN(new_n2808_));
  INV_X1     g02744(.I(new_n2808_), .ZN(new_n2809_));
  NOR2_X1    g02745(.A1(new_n475_), .A2(new_n490_), .ZN(new_n2810_));
  INV_X1     g02746(.I(new_n2810_), .ZN(new_n2811_));
  NAND2_X1   g02747(.A1(new_n160_), .A2(new_n378_), .ZN(new_n2812_));
  NOR3_X1    g02748(.A1(new_n946_), .A2(new_n326_), .A3(new_n264_), .ZN(new_n2813_));
  NOR4_X1    g02749(.A1(new_n119_), .A2(new_n130_), .A3(new_n396_), .A4(new_n437_), .ZN(new_n2814_));
  INV_X1     g02750(.I(new_n2814_), .ZN(new_n2815_));
  NAND4_X1   g02751(.A1(new_n2539_), .A2(new_n2815_), .A3(new_n1387_), .A4(new_n2813_), .ZN(new_n2816_));
  NOR4_X1    g02752(.A1(new_n2816_), .A2(new_n1391_), .A3(new_n2811_), .A4(new_n2812_), .ZN(new_n2817_));
  INV_X1     g02753(.I(new_n2817_), .ZN(new_n2818_));
  NOR4_X1    g02754(.A1(new_n324_), .A2(new_n753_), .A3(new_n359_), .A4(new_n937_), .ZN(new_n2819_));
  NOR4_X1    g02755(.A1(new_n136_), .A2(new_n242_), .A3(new_n260_), .A4(new_n330_), .ZN(new_n2820_));
  INV_X1     g02756(.I(new_n2820_), .ZN(new_n2821_));
  NOR4_X1    g02757(.A1(new_n2821_), .A2(new_n2819_), .A3(new_n687_), .A4(new_n873_), .ZN(new_n2822_));
  NOR4_X1    g02758(.A1(new_n286_), .A2(new_n584_), .A3(new_n1355_), .A4(new_n660_), .ZN(new_n2823_));
  NOR4_X1    g02759(.A1(new_n495_), .A2(new_n656_), .A3(new_n955_), .A4(new_n779_), .ZN(new_n2824_));
  NOR2_X1    g02760(.A1(new_n267_), .A2(new_n453_), .ZN(new_n2825_));
  INV_X1     g02761(.I(new_n2825_), .ZN(new_n2826_));
  NOR3_X1    g02762(.A1(new_n2826_), .A2(new_n2823_), .A3(new_n2824_), .ZN(new_n2827_));
  NOR2_X1    g02763(.A1(new_n212_), .A2(new_n297_), .ZN(new_n2828_));
  INV_X1     g02764(.I(new_n2828_), .ZN(new_n2829_));
  NOR4_X1    g02765(.A1(new_n2829_), .A2(new_n1157_), .A3(new_n124_), .A4(new_n463_), .ZN(new_n2830_));
  NAND4_X1   g02766(.A1(new_n2830_), .A2(new_n313_), .A3(new_n983_), .A4(new_n980_), .ZN(new_n2831_));
  INV_X1     g02767(.I(new_n2831_), .ZN(new_n2832_));
  NAND4_X1   g02768(.A1(new_n2832_), .A2(new_n1928_), .A3(new_n2822_), .A4(new_n2827_), .ZN(new_n2833_));
  NOR2_X1    g02769(.A1(new_n2833_), .A2(new_n2818_), .ZN(new_n2834_));
  INV_X1     g02770(.I(new_n1499_), .ZN(new_n2835_));
  NOR4_X1    g02771(.A1(new_n866_), .A2(new_n549_), .A3(new_n587_), .A4(new_n1984_), .ZN(new_n2836_));
  NOR4_X1    g02772(.A1(new_n2836_), .A2(new_n216_), .A3(new_n268_), .A4(new_n607_), .ZN(new_n2837_));
  NOR2_X1    g02773(.A1(new_n367_), .A2(new_n734_), .ZN(new_n2838_));
  INV_X1     g02774(.I(new_n2838_), .ZN(new_n2839_));
  NOR4_X1    g02775(.A1(new_n2839_), .A2(new_n615_), .A3(new_n306_), .A4(new_n774_), .ZN(new_n2840_));
  NOR2_X1    g02776(.A1(new_n1039_), .A2(new_n1381_), .ZN(new_n2841_));
  NAND4_X1   g02777(.A1(new_n2837_), .A2(new_n2840_), .A3(new_n2835_), .A4(new_n2841_), .ZN(new_n2842_));
  NOR3_X1    g02778(.A1(new_n2445_), .A2(new_n397_), .A3(new_n531_), .ZN(new_n2843_));
  NOR3_X1    g02779(.A1(new_n200_), .A2(new_n213_), .A3(new_n752_), .ZN(new_n2844_));
  NAND4_X1   g02780(.A1(new_n322_), .A2(new_n522_), .A3(new_n1892_), .A4(new_n501_), .ZN(new_n2845_));
  NAND4_X1   g02781(.A1(new_n2843_), .A2(new_n2844_), .A3(new_n1554_), .A4(new_n2845_), .ZN(new_n2846_));
  NOR3_X1    g02782(.A1(new_n2842_), .A2(new_n2846_), .A3(new_n1297_), .ZN(new_n2847_));
  NAND2_X1   g02783(.A1(new_n2834_), .A2(new_n2847_), .ZN(new_n2848_));
  NOR4_X1    g02784(.A1(new_n717_), .A2(new_n1994_), .A3(new_n170_), .A4(new_n817_), .ZN(new_n2849_));
  NOR4_X1    g02785(.A1(new_n2096_), .A2(new_n286_), .A3(new_n374_), .A4(new_n1146_), .ZN(new_n2850_));
  NAND3_X1   g02786(.A1(new_n1825_), .A2(new_n1829_), .A3(new_n572_), .ZN(new_n2851_));
  NOR4_X1    g02787(.A1(new_n2851_), .A2(new_n119_), .A3(new_n297_), .A4(new_n561_), .ZN(new_n2852_));
  NAND3_X1   g02788(.A1(new_n2850_), .A2(new_n2849_), .A3(new_n2852_), .ZN(new_n2853_));
  NOR4_X1    g02789(.A1(new_n172_), .A2(new_n214_), .A3(new_n596_), .A4(new_n577_), .ZN(new_n2854_));
  NOR2_X1    g02790(.A1(new_n1984_), .A2(new_n163_), .ZN(new_n2855_));
  NAND4_X1   g02791(.A1(new_n2855_), .A2(new_n1441_), .A3(new_n1530_), .A4(new_n1190_), .ZN(new_n2856_));
  NOR2_X1    g02792(.A1(new_n2856_), .A2(new_n2854_), .ZN(new_n2857_));
  NAND3_X1   g02793(.A1(new_n690_), .A2(new_n808_), .A3(new_n378_), .ZN(new_n2858_));
  NOR4_X1    g02794(.A1(new_n281_), .A2(new_n304_), .A3(new_n413_), .A4(new_n518_), .ZN(new_n2859_));
  NOR4_X1    g02795(.A1(new_n446_), .A2(new_n154_), .A3(new_n463_), .A4(new_n437_), .ZN(new_n2860_));
  NOR4_X1    g02796(.A1(new_n2860_), .A2(new_n1034_), .A3(new_n2858_), .A4(new_n2859_), .ZN(new_n2861_));
  NOR2_X1    g02797(.A1(new_n260_), .A2(new_n487_), .ZN(new_n2862_));
  NAND4_X1   g02798(.A1(new_n218_), .A2(new_n2862_), .A3(new_n382_), .A4(new_n1018_), .ZN(new_n2863_));
  NOR2_X1    g02799(.A1(new_n2863_), .A2(new_n2385_), .ZN(new_n2864_));
  NAND3_X1   g02800(.A1(new_n2861_), .A2(new_n2864_), .A3(new_n2857_), .ZN(new_n2865_));
  NOR2_X1    g02801(.A1(new_n2853_), .A2(new_n2865_), .ZN(new_n2866_));
  INV_X1     g02802(.I(new_n240_), .ZN(new_n2867_));
  NOR4_X1    g02803(.A1(new_n1245_), .A2(new_n1054_), .A3(new_n1730_), .A4(new_n1976_), .ZN(new_n2868_));
  NOR4_X1    g02804(.A1(new_n1620_), .A2(new_n419_), .A3(new_n734_), .A4(new_n764_), .ZN(new_n2869_));
  INV_X1     g02805(.I(new_n2399_), .ZN(new_n2870_));
  NOR4_X1    g02806(.A1(new_n541_), .A2(new_n496_), .A3(new_n670_), .A4(new_n776_), .ZN(new_n2871_));
  NOR3_X1    g02807(.A1(new_n2871_), .A2(new_n2870_), .A3(new_n697_), .ZN(new_n2872_));
  NAND4_X1   g02808(.A1(new_n711_), .A2(new_n2868_), .A3(new_n2872_), .A4(new_n2869_), .ZN(new_n2873_));
  NOR4_X1    g02809(.A1(new_n534_), .A2(new_n724_), .A3(new_n397_), .A4(new_n955_), .ZN(new_n2874_));
  NAND2_X1   g02810(.A1(new_n187_), .A2(new_n824_), .ZN(new_n2875_));
  NOR4_X1    g02811(.A1(new_n2342_), .A2(new_n604_), .A3(new_n2306_), .A4(new_n2875_), .ZN(new_n2876_));
  INV_X1     g02812(.I(new_n2876_), .ZN(new_n2877_));
  NOR4_X1    g02813(.A1(new_n2873_), .A2(new_n2867_), .A3(new_n2874_), .A4(new_n2877_), .ZN(new_n2878_));
  NOR3_X1    g02814(.A1(new_n763_), .A2(new_n124_), .A3(new_n930_), .ZN(new_n2879_));
  INV_X1     g02815(.I(new_n2879_), .ZN(new_n2880_));
  NOR4_X1    g02816(.A1(new_n774_), .A2(new_n430_), .A3(new_n488_), .A4(new_n770_), .ZN(new_n2881_));
  NAND3_X1   g02817(.A1(new_n2390_), .A2(new_n598_), .A3(new_n643_), .ZN(new_n2882_));
  NOR3_X1    g02818(.A1(new_n2881_), .A2(new_n2880_), .A3(new_n2882_), .ZN(new_n2883_));
  INV_X1     g02819(.I(new_n2219_), .ZN(new_n2884_));
  NOR4_X1    g02820(.A1(new_n2884_), .A2(new_n929_), .A3(new_n533_), .A4(new_n1103_), .ZN(new_n2885_));
  NOR2_X1    g02821(.A1(new_n1084_), .A2(new_n634_), .ZN(new_n2886_));
  NAND4_X1   g02822(.A1(new_n2079_), .A2(new_n1963_), .A3(new_n2591_), .A4(new_n2886_), .ZN(new_n2887_));
  INV_X1     g02823(.I(new_n2887_), .ZN(new_n2888_));
  NAND4_X1   g02824(.A1(new_n2888_), .A2(new_n461_), .A3(new_n2883_), .A4(new_n2885_), .ZN(new_n2889_));
  INV_X1     g02825(.I(new_n2889_), .ZN(new_n2890_));
  AND2_X2    g02826(.A1(new_n2878_), .A2(new_n2890_), .Z(new_n2891_));
  NAND2_X1   g02827(.A1(new_n2891_), .A2(new_n2866_), .ZN(new_n2892_));
  INV_X1     g02828(.I(new_n2892_), .ZN(new_n2893_));
  NOR2_X1    g02829(.A1(new_n2893_), .A2(\a[23] ), .ZN(new_n2894_));
  NOR2_X1    g02830(.A1(new_n2894_), .A2(new_n2848_), .ZN(new_n2895_));
  NOR2_X1    g02831(.A1(new_n2892_), .A2(new_n84_), .ZN(new_n2896_));
  NOR2_X1    g02832(.A1(new_n2895_), .A2(new_n2896_), .ZN(new_n2897_));
  NOR2_X1    g02833(.A1(new_n2897_), .A2(new_n2809_), .ZN(new_n2898_));
  INV_X1     g02834(.I(new_n2898_), .ZN(new_n2899_));
  NAND2_X1   g02835(.A1(new_n2897_), .A2(new_n2809_), .ZN(new_n2900_));
  AOI21_X1   g02836(.A1(new_n2899_), .A2(new_n2900_), .B(new_n2775_), .ZN(new_n2901_));
  INV_X1     g02837(.I(new_n2775_), .ZN(new_n2902_));
  XOR2_X1    g02838(.A1(new_n2897_), .A2(new_n2808_), .Z(new_n2903_));
  NOR2_X1    g02839(.A1(new_n2902_), .A2(new_n2903_), .ZN(new_n2904_));
  NOR2_X1    g02840(.A1(new_n2904_), .A2(new_n2901_), .ZN(new_n2905_));
  INV_X1     g02841(.I(new_n2905_), .ZN(new_n2906_));
  AOI21_X1   g02842(.A1(new_n2503_), .A2(new_n2506_), .B(new_n897_), .ZN(new_n2907_));
  INV_X1     g02843(.I(new_n2907_), .ZN(new_n2908_));
  NAND3_X1   g02844(.A1(new_n2503_), .A2(new_n2506_), .A3(new_n897_), .ZN(new_n2909_));
  NAND2_X1   g02845(.A1(new_n2908_), .A2(new_n2909_), .ZN(new_n2910_));
  XOR2_X1    g02846(.A1(new_n1008_), .A2(new_n897_), .Z(new_n2911_));
  INV_X1     g02847(.I(new_n2911_), .ZN(new_n2912_));
  NAND3_X1   g02848(.A1(new_n2910_), .A2(new_n814_), .A3(new_n2912_), .ZN(new_n2913_));
  INV_X1     g02849(.I(new_n2909_), .ZN(new_n2914_));
  OAI21_X1   g02850(.A1(new_n2914_), .A2(new_n2907_), .B(new_n2912_), .ZN(new_n2915_));
  NAND2_X1   g02851(.A1(new_n2915_), .A2(new_n813_), .ZN(new_n2916_));
  NAND2_X1   g02852(.A1(new_n2913_), .A2(new_n2916_), .ZN(new_n2917_));
  OAI21_X1   g02853(.A1(new_n896_), .A2(new_n2767_), .B(new_n2764_), .ZN(new_n2918_));
  OAI22_X1   g02854(.A1(new_n813_), .A2(new_n2772_), .B1(new_n1008_), .B2(new_n2771_), .ZN(new_n2919_));
  NOR2_X1    g02855(.A1(new_n2919_), .A2(new_n2918_), .ZN(new_n2920_));
  NAND2_X1   g02856(.A1(new_n2917_), .A2(new_n2920_), .ZN(new_n2921_));
  INV_X1     g02857(.I(new_n2921_), .ZN(new_n2922_));
  NOR3_X1    g02858(.A1(new_n147_), .A2(new_n615_), .A3(new_n262_), .ZN(new_n2923_));
  INV_X1     g02859(.I(new_n2923_), .ZN(new_n2924_));
  NOR4_X1    g02860(.A1(new_n488_), .A2(new_n498_), .A3(new_n556_), .A4(new_n376_), .ZN(new_n2925_));
  NOR4_X1    g02861(.A1(new_n2924_), .A2(new_n751_), .A3(new_n213_), .A4(new_n2925_), .ZN(new_n2926_));
  NAND4_X1   g02862(.A1(new_n436_), .A2(new_n871_), .A3(new_n1725_), .A4(new_n665_), .ZN(new_n2927_));
  NAND3_X1   g02863(.A1(new_n1961_), .A2(new_n313_), .A3(new_n592_), .ZN(new_n2928_));
  NOR4_X1    g02864(.A1(new_n2928_), .A2(new_n988_), .A3(new_n154_), .A4(new_n2927_), .ZN(new_n2929_));
  INV_X1     g02865(.I(new_n2624_), .ZN(new_n2930_));
  NOR4_X1    g02866(.A1(new_n2930_), .A2(new_n98_), .A3(new_n280_), .A4(new_n298_), .ZN(new_n2931_));
  INV_X1     g02867(.I(new_n1356_), .ZN(new_n2932_));
  NAND2_X1   g02868(.A1(new_n829_), .A2(new_n1952_), .ZN(new_n2933_));
  NOR3_X1    g02869(.A1(new_n2932_), .A2(new_n2933_), .A3(new_n1944_), .ZN(new_n2934_));
  NAND4_X1   g02870(.A1(new_n2934_), .A2(new_n2926_), .A3(new_n2929_), .A4(new_n2931_), .ZN(new_n2935_));
  NOR2_X1    g02871(.A1(new_n2935_), .A2(new_n2475_), .ZN(new_n2936_));
  NOR2_X1    g02872(.A1(new_n102_), .A2(new_n117_), .ZN(new_n2937_));
  NOR4_X1    g02873(.A1(new_n2937_), .A2(new_n211_), .A3(new_n406_), .A4(new_n531_), .ZN(new_n2938_));
  NAND3_X1   g02874(.A1(new_n2122_), .A2(new_n965_), .A3(new_n797_), .ZN(new_n2939_));
  NOR2_X1    g02875(.A1(new_n648_), .A2(new_n801_), .ZN(new_n2940_));
  NAND4_X1   g02876(.A1(new_n2938_), .A2(new_n606_), .A3(new_n2939_), .A4(new_n2940_), .ZN(new_n2941_));
  NOR2_X1    g02877(.A1(new_n772_), .A2(new_n660_), .ZN(new_n2942_));
  NAND4_X1   g02878(.A1(new_n2597_), .A2(new_n888_), .A3(new_n2942_), .A4(new_n2233_), .ZN(new_n2943_));
  NOR2_X1    g02879(.A1(new_n1152_), .A2(new_n719_), .ZN(new_n2944_));
  NAND4_X1   g02880(.A1(new_n2622_), .A2(new_n2944_), .A3(new_n641_), .A4(new_n2244_), .ZN(new_n2945_));
  NOR3_X1    g02881(.A1(new_n465_), .A2(new_n163_), .A3(new_n506_), .ZN(new_n2946_));
  NAND4_X1   g02882(.A1(new_n2946_), .A2(new_n351_), .A3(new_n1129_), .A4(new_n1068_), .ZN(new_n2947_));
  OR4_X2     g02883(.A1(new_n2941_), .A2(new_n2943_), .A3(new_n2945_), .A4(new_n2947_), .Z(new_n2948_));
  NOR3_X1    g02884(.A1(new_n2948_), .A2(new_n1661_), .A3(new_n1675_), .ZN(new_n2949_));
  NAND2_X1   g02885(.A1(new_n2949_), .A2(new_n2936_), .ZN(new_n2950_));
  INV_X1     g02886(.I(new_n2950_), .ZN(new_n2951_));
  INV_X1     g02887(.I(new_n1443_), .ZN(new_n2952_));
  NOR4_X1    g02888(.A1(new_n1045_), .A2(new_n1379_), .A3(new_n713_), .A4(new_n1247_), .ZN(new_n2953_));
  NOR2_X1    g02889(.A1(new_n956_), .A2(new_n226_), .ZN(new_n2954_));
  INV_X1     g02890(.I(new_n2954_), .ZN(new_n2955_));
  NOR4_X1    g02891(.A1(new_n320_), .A2(new_n518_), .A3(new_n736_), .A4(new_n749_), .ZN(new_n2956_));
  NOR3_X1    g02892(.A1(new_n102_), .A2(new_n751_), .A3(new_n841_), .ZN(new_n2957_));
  INV_X1     g02893(.I(new_n2957_), .ZN(new_n2958_));
  NOR3_X1    g02894(.A1(new_n2955_), .A2(new_n2956_), .A3(new_n2958_), .ZN(new_n2959_));
  NOR3_X1    g02895(.A1(new_n1014_), .A2(new_n625_), .A3(new_n637_), .ZN(new_n2960_));
  NOR4_X1    g02896(.A1(new_n640_), .A2(new_n297_), .A3(new_n366_), .A4(new_n776_), .ZN(new_n2961_));
  NOR4_X1    g02897(.A1(new_n2961_), .A2(new_n173_), .A3(new_n388_), .A4(new_n946_), .ZN(new_n2962_));
  NAND4_X1   g02898(.A1(new_n2960_), .A2(new_n957_), .A3(new_n2962_), .A4(new_n1001_), .ZN(new_n2963_));
  INV_X1     g02899(.I(new_n2963_), .ZN(new_n2964_));
  NAND4_X1   g02900(.A1(new_n2964_), .A2(new_n2952_), .A3(new_n2953_), .A4(new_n2959_), .ZN(new_n2965_));
  INV_X1     g02901(.I(new_n2965_), .ZN(new_n2966_));
  NOR4_X1    g02902(.A1(new_n324_), .A2(new_n611_), .A3(new_n721_), .A4(new_n660_), .ZN(new_n2967_));
  NAND2_X1   g02903(.A1(new_n1205_), .A2(new_n2624_), .ZN(new_n2968_));
  NAND3_X1   g02904(.A1(new_n2862_), .A2(new_n197_), .A3(new_n773_), .ZN(new_n2969_));
  NOR3_X1    g02905(.A1(new_n1011_), .A2(new_n548_), .A3(new_n213_), .ZN(new_n2970_));
  INV_X1     g02906(.I(new_n2970_), .ZN(new_n2971_));
  NOR4_X1    g02907(.A1(new_n2968_), .A2(new_n2971_), .A3(new_n2969_), .A4(new_n2967_), .ZN(new_n2972_));
  NAND3_X1   g02908(.A1(new_n184_), .A2(new_n551_), .A3(new_n999_), .ZN(new_n2973_));
  NOR4_X1    g02909(.A1(new_n2973_), .A2(new_n261_), .A3(new_n304_), .A4(new_n1996_), .ZN(new_n2974_));
  NOR2_X1    g02910(.A1(new_n740_), .A2(new_n535_), .ZN(new_n2975_));
  INV_X1     g02911(.I(new_n2975_), .ZN(new_n2976_));
  NAND4_X1   g02912(.A1(new_n1336_), .A2(new_n1126_), .A3(new_n624_), .A4(new_n1952_), .ZN(new_n2977_));
  NOR4_X1    g02913(.A1(new_n2976_), .A2(new_n2977_), .A3(new_n1615_), .A4(new_n2083_), .ZN(new_n2978_));
  NAND3_X1   g02914(.A1(new_n2978_), .A2(new_n2972_), .A3(new_n2974_), .ZN(new_n2979_));
  INV_X1     g02915(.I(new_n2979_), .ZN(new_n2980_));
  INV_X1     g02916(.I(new_n692_), .ZN(new_n2981_));
  INV_X1     g02917(.I(new_n138_), .ZN(new_n2982_));
  NOR2_X1    g02918(.A1(new_n2826_), .A2(new_n2982_), .ZN(new_n2983_));
  NOR4_X1    g02919(.A1(new_n465_), .A2(new_n515_), .A3(new_n241_), .A4(new_n944_), .ZN(new_n2984_));
  NOR2_X1    g02920(.A1(new_n2984_), .A2(new_n1643_), .ZN(new_n2985_));
  NAND4_X1   g02921(.A1(new_n2983_), .A2(new_n473_), .A3(new_n852_), .A4(new_n2985_), .ZN(new_n2986_));
  NOR3_X1    g02922(.A1(new_n333_), .A2(new_n359_), .A3(new_n610_), .ZN(new_n2987_));
  NOR4_X1    g02923(.A1(new_n788_), .A2(new_n198_), .A3(new_n192_), .A4(new_n262_), .ZN(new_n2988_));
  NAND2_X1   g02924(.A1(new_n2988_), .A2(new_n2987_), .ZN(new_n2989_));
  NOR4_X1    g02925(.A1(new_n486_), .A2(new_n772_), .A3(new_n744_), .A4(new_n468_), .ZN(new_n2990_));
  NOR4_X1    g02926(.A1(new_n117_), .A2(new_n698_), .A3(new_n428_), .A4(new_n92_), .ZN(new_n2991_));
  NOR3_X1    g02927(.A1(new_n2989_), .A2(new_n2990_), .A3(new_n2991_), .ZN(new_n2992_));
  INV_X1     g02928(.I(new_n2992_), .ZN(new_n2993_));
  INV_X1     g02929(.I(new_n819_), .ZN(new_n2994_));
  NOR3_X1    g02930(.A1(new_n2994_), .A2(new_n573_), .A3(new_n217_), .ZN(new_n2995_));
  NOR3_X1    g02931(.A1(new_n770_), .A2(new_n449_), .A3(new_n352_), .ZN(new_n2996_));
  NOR3_X1    g02932(.A1(new_n149_), .A2(new_n638_), .A3(new_n330_), .ZN(new_n2997_));
  NAND4_X1   g02933(.A1(new_n2995_), .A2(new_n2996_), .A3(new_n2997_), .A4(new_n1751_), .ZN(new_n2998_));
  NOR4_X1    g02934(.A1(new_n2981_), .A2(new_n2986_), .A3(new_n2993_), .A4(new_n2998_), .ZN(new_n2999_));
  NAND3_X1   g02935(.A1(new_n2966_), .A2(new_n2999_), .A3(new_n2980_), .ZN(new_n3000_));
  INV_X1     g02936(.I(new_n3000_), .ZN(new_n3001_));
  NAND4_X1   g02937(.A1(new_n382_), .A2(new_n2240_), .A3(new_n880_), .A4(new_n1601_), .ZN(new_n3002_));
  NAND4_X1   g02938(.A1(new_n2691_), .A2(new_n542_), .A3(new_n2113_), .A4(new_n3002_), .ZN(new_n3003_));
  NAND2_X1   g02939(.A1(new_n2164_), .A2(new_n2082_), .ZN(new_n3004_));
  NAND4_X1   g02940(.A1(new_n1329_), .A2(new_n911_), .A3(new_n953_), .A4(new_n1153_), .ZN(new_n3005_));
  NOR4_X1    g02941(.A1(new_n3003_), .A2(new_n2457_), .A3(new_n3004_), .A4(new_n3005_), .ZN(new_n3006_));
  AND3_X2    g02942(.A1(new_n3006_), .A2(new_n224_), .A3(new_n2378_), .Z(new_n3007_));
  INV_X1     g02943(.I(new_n1794_), .ZN(new_n3008_));
  NOR3_X1    g02944(.A1(new_n1620_), .A2(new_n124_), .A3(new_n607_), .ZN(new_n3009_));
  NAND4_X1   g02945(.A1(new_n2587_), .A2(new_n1284_), .A3(new_n3008_), .A4(new_n3009_), .ZN(new_n3010_));
  NAND3_X1   g02946(.A1(new_n353_), .A2(new_n568_), .A3(new_n809_), .ZN(new_n3011_));
  NOR4_X1    g02947(.A1(new_n2047_), .A2(new_n3011_), .A3(new_n490_), .A4(new_n465_), .ZN(new_n3012_));
  NOR2_X1    g02948(.A1(new_n232_), .A2(new_n506_), .ZN(new_n3013_));
  NAND4_X1   g02949(.A1(new_n336_), .A2(new_n1380_), .A3(new_n3013_), .A4(new_n113_), .ZN(new_n3014_));
  NOR4_X1    g02950(.A1(new_n3014_), .A2(new_n2146_), .A3(new_n1493_), .A4(new_n2234_), .ZN(new_n3015_));
  NAND2_X1   g02951(.A1(new_n3015_), .A2(new_n3012_), .ZN(new_n3016_));
  NOR2_X1    g02952(.A1(new_n3010_), .A2(new_n3016_), .ZN(new_n3017_));
  NOR4_X1    g02953(.A1(new_n994_), .A2(new_n332_), .A3(new_n177_), .A4(new_n1782_), .ZN(new_n3018_));
  NAND4_X1   g02954(.A1(new_n481_), .A2(new_n1448_), .A3(new_n686_), .A4(new_n1662_), .ZN(new_n3019_));
  NAND4_X1   g02955(.A1(new_n1489_), .A2(new_n807_), .A3(new_n1468_), .A4(new_n1059_), .ZN(new_n3020_));
  NAND4_X1   g02956(.A1(new_n3018_), .A2(new_n2923_), .A3(new_n3019_), .A4(new_n3020_), .ZN(new_n3021_));
  INV_X1     g02957(.I(new_n347_), .ZN(new_n3022_));
  NAND3_X1   g02958(.A1(new_n3022_), .A2(new_n1105_), .A3(new_n832_), .ZN(new_n3023_));
  NOR3_X1    g02959(.A1(new_n86_), .A2(new_n776_), .A3(new_n468_), .ZN(new_n3024_));
  NAND4_X1   g02960(.A1(new_n1816_), .A2(new_n1088_), .A3(new_n441_), .A4(new_n395_), .ZN(new_n3025_));
  NAND2_X1   g02961(.A1(new_n3025_), .A2(new_n3024_), .ZN(new_n3026_));
  NOR4_X1    g02962(.A1(new_n3026_), .A2(new_n1039_), .A3(new_n1160_), .A4(new_n3023_), .ZN(new_n3027_));
  INV_X1     g02963(.I(new_n3027_), .ZN(new_n3028_));
  NOR3_X1    g02964(.A1(new_n3028_), .A2(new_n3021_), .A3(new_n1517_), .ZN(new_n3029_));
  AND2_X2    g02965(.A1(new_n3029_), .A2(new_n3017_), .Z(new_n3030_));
  NAND2_X1   g02966(.A1(new_n3030_), .A2(new_n3007_), .ZN(new_n3031_));
  INV_X1     g02967(.I(new_n3031_), .ZN(new_n3032_));
  NOR2_X1    g02968(.A1(new_n3032_), .A2(\a[20] ), .ZN(new_n3033_));
  INV_X1     g02969(.I(new_n3033_), .ZN(new_n3034_));
  INV_X1     g02970(.I(\a[20] ), .ZN(new_n3035_));
  NOR2_X1    g02971(.A1(new_n3031_), .A2(new_n3035_), .ZN(new_n3036_));
  AOI21_X1   g02972(.A1(new_n3034_), .A2(new_n3001_), .B(new_n3036_), .ZN(new_n3037_));
  NAND2_X1   g02973(.A1(new_n3037_), .A2(new_n2951_), .ZN(new_n3038_));
  NAND2_X1   g02974(.A1(new_n2922_), .A2(new_n3038_), .ZN(new_n3039_));
  OR2_X2     g02975(.A1(new_n3037_), .A2(new_n2951_), .Z(new_n3040_));
  NAND2_X1   g02976(.A1(new_n3039_), .A2(new_n3040_), .ZN(new_n3041_));
  INV_X1     g02977(.I(new_n3041_), .ZN(new_n3042_));
  NOR2_X1    g02978(.A1(new_n2951_), .A2(new_n2848_), .ZN(new_n3043_));
  INV_X1     g02979(.I(new_n2848_), .ZN(new_n3044_));
  NOR2_X1    g02980(.A1(new_n3044_), .A2(new_n2950_), .ZN(new_n3045_));
  INV_X1     g02981(.I(new_n3045_), .ZN(new_n3046_));
  OAI21_X1   g02982(.A1(new_n3042_), .A2(new_n3043_), .B(new_n3046_), .ZN(new_n3047_));
  XOR2_X1    g02983(.A1(new_n2559_), .A2(new_n529_), .Z(new_n3048_));
  NAND2_X1   g02984(.A1(new_n2566_), .A2(new_n3048_), .ZN(new_n3049_));
  AND2_X2    g02985(.A1(new_n2571_), .A2(new_n2568_), .Z(new_n3050_));
  OAI21_X1   g02986(.A1(new_n2566_), .A2(new_n3050_), .B(new_n3049_), .ZN(new_n3051_));
  OAI21_X1   g02987(.A1(new_n813_), .A2(new_n2771_), .B(new_n2764_), .ZN(new_n3052_));
  OAI22_X1   g02988(.A1(new_n2559_), .A2(new_n2767_), .B1(new_n529_), .B2(new_n2772_), .ZN(new_n3053_));
  NOR2_X1    g02989(.A1(new_n3053_), .A2(new_n3052_), .ZN(new_n3054_));
  NAND2_X1   g02990(.A1(new_n3051_), .A2(new_n3054_), .ZN(new_n3055_));
  OAI21_X1   g02991(.A1(new_n2894_), .A2(new_n2896_), .B(new_n3044_), .ZN(new_n3056_));
  XOR2_X1    g02992(.A1(new_n2892_), .A2(\a[23] ), .Z(new_n3057_));
  OAI21_X1   g02993(.A1(new_n3044_), .A2(new_n3057_), .B(new_n3056_), .ZN(new_n3058_));
  INV_X1     g02994(.I(new_n3058_), .ZN(new_n3059_));
  NAND2_X1   g02995(.A1(new_n3055_), .A2(new_n3059_), .ZN(new_n3060_));
  NOR2_X1    g02996(.A1(new_n3055_), .A2(new_n3059_), .ZN(new_n3061_));
  AOI21_X1   g02997(.A1(new_n3047_), .A2(new_n3060_), .B(new_n3061_), .ZN(new_n3062_));
  INV_X1     g02998(.I(new_n3062_), .ZN(new_n3063_));
  NOR2_X1    g02999(.A1(new_n2906_), .A2(new_n3063_), .ZN(new_n3064_));
  NOR2_X1    g03000(.A1(new_n2754_), .A2(new_n3064_), .ZN(new_n3065_));
  NOR2_X1    g03001(.A1(new_n2905_), .A2(new_n3062_), .ZN(new_n3066_));
  NOR2_X1    g03002(.A1(new_n3065_), .A2(new_n3066_), .ZN(new_n3067_));
  INV_X1     g03003(.I(new_n3067_), .ZN(new_n3068_));
  INV_X1     g03004(.I(new_n2755_), .ZN(new_n3069_));
  NOR3_X1    g03005(.A1(new_n2719_), .A2(new_n2718_), .A3(new_n2570_), .ZN(new_n3070_));
  OAI21_X1   g03006(.A1(new_n2719_), .A2(new_n2570_), .B(new_n2718_), .ZN(new_n3071_));
  INV_X1     g03007(.I(new_n3071_), .ZN(new_n3072_));
  OAI21_X1   g03008(.A1(new_n3072_), .A2(new_n3070_), .B(new_n3069_), .ZN(new_n3073_));
  XOR2_X1    g03009(.A1(new_n3073_), .A2(new_n2615_), .Z(new_n3074_));
  NOR2_X1    g03010(.A1(new_n2614_), .A2(new_n2772_), .ZN(new_n3075_));
  NOR2_X1    g03011(.A1(new_n529_), .A2(new_n2771_), .ZN(new_n3076_));
  NOR2_X1    g03012(.A1(new_n694_), .A2(new_n2767_), .ZN(new_n3077_));
  NOR4_X1    g03013(.A1(new_n3077_), .A2(new_n2763_), .A3(new_n3075_), .A4(new_n3076_), .ZN(new_n3078_));
  NAND2_X1   g03014(.A1(new_n3074_), .A2(new_n3078_), .ZN(new_n3079_));
  NOR3_X1    g03015(.A1(new_n1266_), .A2(new_n569_), .A3(new_n1434_), .ZN(new_n3080_));
  NAND2_X1   g03016(.A1(new_n2437_), .A2(new_n2328_), .ZN(new_n3081_));
  NOR4_X1    g03017(.A1(new_n3081_), .A2(new_n774_), .A3(new_n841_), .A4(new_n1865_), .ZN(new_n3082_));
  NAND4_X1   g03018(.A1(new_n414_), .A2(new_n435_), .A3(new_n522_), .A4(new_n1325_), .ZN(new_n3083_));
  NAND4_X1   g03019(.A1(new_n3082_), .A2(new_n3080_), .A3(new_n986_), .A4(new_n3083_), .ZN(new_n3084_));
  NOR4_X1    g03020(.A1(new_n1355_), .A2(new_n1084_), .A3(new_n352_), .A4(new_n1138_), .ZN(new_n3085_));
  NOR3_X1    g03021(.A1(new_n3085_), .A2(new_n459_), .A3(new_n604_), .ZN(new_n3086_));
  NOR2_X1    g03022(.A1(new_n638_), .A2(new_n783_), .ZN(new_n3087_));
  NOR2_X1    g03023(.A1(new_n1157_), .A2(new_n577_), .ZN(new_n3088_));
  NAND4_X1   g03024(.A1(new_n3086_), .A2(new_n1426_), .A3(new_n3087_), .A4(new_n3088_), .ZN(new_n3089_));
  NOR3_X1    g03025(.A1(new_n591_), .A2(new_n584_), .A3(new_n430_), .ZN(new_n3090_));
  NOR3_X1    g03026(.A1(new_n488_), .A2(new_n510_), .A3(new_n556_), .ZN(new_n3091_));
  NOR2_X1    g03027(.A1(new_n381_), .A2(new_n453_), .ZN(new_n3092_));
  NAND4_X1   g03028(.A1(new_n3090_), .A2(new_n3091_), .A3(new_n2038_), .A4(new_n3092_), .ZN(new_n3093_));
  NAND4_X1   g03029(.A1(new_n690_), .A2(new_n508_), .A3(new_n1454_), .A4(new_n999_), .ZN(new_n3094_));
  NOR3_X1    g03030(.A1(new_n541_), .A2(new_n384_), .A3(new_n1168_), .ZN(new_n3095_));
  NAND4_X1   g03031(.A1(new_n423_), .A2(new_n872_), .A3(new_n1796_), .A4(new_n1662_), .ZN(new_n3096_));
  NAND3_X1   g03032(.A1(new_n3095_), .A2(new_n3094_), .A3(new_n3096_), .ZN(new_n3097_));
  NOR4_X1    g03033(.A1(new_n3084_), .A2(new_n3089_), .A3(new_n3093_), .A4(new_n3097_), .ZN(new_n3098_));
  NOR2_X1    g03034(.A1(new_n714_), .A2(new_n910_), .ZN(new_n3099_));
  INV_X1     g03035(.I(new_n3099_), .ZN(new_n3100_));
  NOR2_X1    g03036(.A1(new_n267_), .A2(new_n637_), .ZN(new_n3101_));
  INV_X1     g03037(.I(new_n3101_), .ZN(new_n3102_));
  NOR4_X1    g03038(.A1(new_n3102_), .A2(new_n254_), .A3(new_n1632_), .A4(new_n3100_), .ZN(new_n3103_));
  NOR3_X1    g03039(.A1(new_n216_), .A2(new_n238_), .A3(new_n449_), .ZN(new_n3104_));
  NAND4_X1   g03040(.A1(new_n220_), .A2(new_n197_), .A3(new_n1305_), .A4(new_n1892_), .ZN(new_n3105_));
  NAND4_X1   g03041(.A1(new_n3103_), .A2(new_n2404_), .A3(new_n3104_), .A4(new_n3105_), .ZN(new_n3106_));
  NOR2_X1    g03042(.A1(new_n195_), .A2(new_n3106_), .ZN(new_n3107_));
  AOI21_X1   g03043(.A1(new_n3098_), .A2(new_n3107_), .B(new_n2808_), .ZN(new_n3108_));
  NAND2_X1   g03044(.A1(new_n3107_), .A2(new_n3098_), .ZN(new_n3109_));
  NOR2_X1    g03045(.A1(new_n2809_), .A2(new_n3109_), .ZN(new_n3110_));
  NOR2_X1    g03046(.A1(new_n3110_), .A2(new_n3108_), .ZN(new_n3111_));
  NOR2_X1    g03047(.A1(new_n3079_), .A2(new_n3111_), .ZN(new_n3112_));
  INV_X1     g03048(.I(new_n3079_), .ZN(new_n3113_));
  XOR2_X1    g03049(.A1(new_n2808_), .A2(new_n3109_), .Z(new_n3114_));
  NOR2_X1    g03050(.A1(new_n3113_), .A2(new_n3114_), .ZN(new_n3115_));
  NOR2_X1    g03051(.A1(new_n3115_), .A2(new_n3112_), .ZN(new_n3116_));
  AOI21_X1   g03052(.A1(new_n2902_), .A2(new_n2900_), .B(new_n2898_), .ZN(new_n3117_));
  NAND2_X1   g03053(.A1(new_n3116_), .A2(new_n3117_), .ZN(new_n3118_));
  NOR2_X1    g03054(.A1(new_n3116_), .A2(new_n3117_), .ZN(new_n3119_));
  AOI21_X1   g03055(.A1(new_n3068_), .A2(new_n3118_), .B(new_n3119_), .ZN(new_n3120_));
  NOR2_X1    g03056(.A1(new_n1984_), .A2(new_n297_), .ZN(new_n3121_));
  NAND2_X1   g03057(.A1(new_n543_), .A2(new_n3121_), .ZN(new_n3122_));
  NOR4_X1    g03058(.A1(new_n239_), .A2(new_n591_), .A3(new_n899_), .A4(new_n490_), .ZN(new_n3123_));
  NAND3_X1   g03059(.A1(new_n1712_), .A2(new_n1025_), .A3(new_n564_), .ZN(new_n3124_));
  NOR4_X1    g03060(.A1(new_n3122_), .A2(new_n3124_), .A3(new_n2703_), .A4(new_n3123_), .ZN(new_n3125_));
  NOR4_X1    g03061(.A1(new_n289_), .A2(new_n482_), .A3(new_n1146_), .A4(new_n652_), .ZN(new_n3126_));
  NAND2_X1   g03062(.A1(new_n1921_), .A2(new_n1065_), .ZN(new_n3127_));
  NOR3_X1    g03063(.A1(new_n3126_), .A2(new_n783_), .A3(new_n3127_), .ZN(new_n3128_));
  NOR2_X1    g03064(.A1(new_n753_), .A2(new_n1175_), .ZN(new_n3129_));
  NAND4_X1   g03065(.A1(new_n816_), .A2(new_n2444_), .A3(new_n3129_), .A4(new_n1315_), .ZN(new_n3130_));
  NOR4_X1    g03066(.A1(new_n3130_), .A2(new_n2582_), .A3(new_n1589_), .A4(new_n1620_), .ZN(new_n3131_));
  NAND3_X1   g03067(.A1(new_n3125_), .A2(new_n3131_), .A3(new_n3128_), .ZN(new_n3132_));
  INV_X1     g03068(.I(new_n3132_), .ZN(new_n3133_));
  NOR2_X1    g03069(.A1(new_n2713_), .A2(new_n202_), .ZN(new_n3134_));
  NAND3_X1   g03070(.A1(new_n3133_), .A2(new_n1572_), .A3(new_n3134_), .ZN(new_n3135_));
  NOR4_X1    g03071(.A1(new_n3100_), .A2(new_n937_), .A3(new_n468_), .A4(new_n656_), .ZN(new_n3136_));
  INV_X1     g03072(.I(new_n1126_), .ZN(new_n3137_));
  NOR3_X1    g03073(.A1(new_n1197_), .A2(new_n1014_), .A3(new_n3137_), .ZN(new_n3138_));
  NAND4_X1   g03074(.A1(new_n3022_), .A2(new_n551_), .A3(new_n1393_), .A4(new_n1106_), .ZN(new_n3139_));
  NOR2_X1    g03075(.A1(new_n950_), .A2(new_n3139_), .ZN(new_n3140_));
  NAND4_X1   g03076(.A1(new_n3140_), .A2(new_n635_), .A3(new_n3136_), .A4(new_n3138_), .ZN(new_n3141_));
  NOR2_X1    g03077(.A1(new_n3135_), .A2(new_n3141_), .ZN(new_n3142_));
  NAND4_X1   g03078(.A1(new_n2725_), .A2(new_n2664_), .A3(new_n2726_), .A4(new_n2716_), .ZN(new_n3143_));
  NAND2_X1   g03079(.A1(new_n2725_), .A2(new_n2726_), .ZN(new_n3144_));
  NAND3_X1   g03080(.A1(new_n3144_), .A2(new_n2665_), .A3(new_n2728_), .ZN(new_n3145_));
  INV_X1     g03081(.I(new_n2037_), .ZN(new_n3146_));
  NOR3_X1    g03082(.A1(new_n576_), .A2(new_n1087_), .A3(new_n1076_), .ZN(new_n3147_));
  INV_X1     g03083(.I(new_n3147_), .ZN(new_n3148_));
  NOR4_X1    g03084(.A1(new_n216_), .A2(new_n603_), .A3(new_n698_), .A4(new_n741_), .ZN(new_n3149_));
  NOR3_X1    g03085(.A1(new_n1420_), .A2(new_n247_), .A3(new_n474_), .ZN(new_n3150_));
  INV_X1     g03086(.I(new_n3150_), .ZN(new_n3151_));
  NOR3_X1    g03087(.A1(new_n3151_), .A2(new_n3148_), .A3(new_n3149_), .ZN(new_n3152_));
  NAND4_X1   g03088(.A1(new_n3152_), .A2(new_n2701_), .A3(new_n80_), .A4(new_n274_), .ZN(new_n3153_));
  NOR2_X1    g03089(.A1(new_n3153_), .A2(new_n3146_), .ZN(new_n3154_));
  INV_X1     g03090(.I(new_n3154_), .ZN(new_n3155_));
  INV_X1     g03091(.I(new_n344_), .ZN(new_n3156_));
  NAND3_X1   g03092(.A1(new_n103_), .A2(new_n1242_), .A3(new_n1770_), .ZN(new_n3157_));
  NAND3_X1   g03093(.A1(new_n922_), .A2(new_n220_), .A3(new_n983_), .ZN(new_n3158_));
  NOR2_X1    g03094(.A1(new_n198_), .A2(new_n192_), .ZN(new_n3159_));
  NAND2_X1   g03095(.A1(new_n2125_), .A2(new_n3159_), .ZN(new_n3160_));
  NOR4_X1    g03096(.A1(new_n3160_), .A2(new_n696_), .A3(new_n3157_), .A4(new_n3158_), .ZN(new_n3161_));
  NOR4_X1    g03097(.A1(new_n1149_), .A2(new_n1346_), .A3(new_n413_), .A4(new_n640_), .ZN(new_n3162_));
  NAND2_X1   g03098(.A1(new_n3161_), .A2(new_n3162_), .ZN(new_n3163_));
  NOR4_X1    g03099(.A1(new_n3163_), .A2(new_n244_), .A3(new_n3156_), .A4(new_n3081_), .ZN(new_n3164_));
  INV_X1     g03100(.I(new_n3164_), .ZN(new_n3165_));
  NOR2_X1    g03101(.A1(new_n3155_), .A2(new_n3165_), .ZN(new_n3166_));
  NOR3_X1    g03102(.A1(new_n3141_), .A2(new_n202_), .A3(new_n2338_), .ZN(new_n3167_));
  NAND2_X1   g03103(.A1(new_n3166_), .A2(new_n3167_), .ZN(new_n3168_));
  XOR2_X1    g03104(.A1(new_n3168_), .A2(new_n2716_), .Z(new_n3169_));
  INV_X1     g03105(.I(new_n3169_), .ZN(new_n3170_));
  NAND3_X1   g03106(.A1(new_n3145_), .A2(new_n3143_), .A3(new_n3170_), .ZN(new_n3171_));
  NOR2_X1    g03107(.A1(new_n3171_), .A2(new_n3142_), .ZN(new_n3172_));
  AND2_X2    g03108(.A1(new_n3171_), .A2(new_n3142_), .Z(new_n3173_));
  OR2_X2     g03109(.A1(new_n3173_), .A2(new_n3172_), .Z(new_n3174_));
  INV_X1     g03110(.I(new_n2750_), .ZN(new_n3175_));
  INV_X1     g03111(.I(new_n3168_), .ZN(new_n3176_));
  OAI22_X1   g03112(.A1(new_n3176_), .A2(new_n2742_), .B1(new_n3175_), .B2(new_n3142_), .ZN(new_n3177_));
  NAND2_X1   g03113(.A1(new_n2728_), .A2(new_n2746_), .ZN(new_n3178_));
  AOI21_X1   g03114(.A1(new_n3177_), .A2(new_n3178_), .B(new_n2737_), .ZN(new_n3179_));
  NAND2_X1   g03115(.A1(new_n3174_), .A2(new_n3179_), .ZN(new_n3180_));
  XOR2_X1    g03116(.A1(new_n3180_), .A2(\a[29] ), .Z(new_n3181_));
  NOR2_X1    g03117(.A1(new_n3079_), .A2(new_n3108_), .ZN(new_n3182_));
  NOR2_X1    g03118(.A1(new_n3182_), .A2(new_n3110_), .ZN(new_n3183_));
  INV_X1     g03119(.I(new_n3183_), .ZN(new_n3184_));
  NAND2_X1   g03120(.A1(new_n2721_), .A2(new_n2723_), .ZN(new_n3185_));
  XOR2_X1    g03121(.A1(new_n2614_), .A2(new_n2664_), .Z(new_n3186_));
  OAI22_X1   g03122(.A1(new_n2617_), .A2(new_n2619_), .B1(new_n2666_), .B2(new_n2668_), .ZN(new_n3187_));
  OAI21_X1   g03123(.A1(new_n3185_), .A2(new_n3186_), .B(new_n3187_), .ZN(new_n3188_));
  INV_X1     g03124(.I(new_n2767_), .ZN(new_n3189_));
  NAND2_X1   g03125(.A1(new_n2615_), .A2(new_n3189_), .ZN(new_n3190_));
  NAND2_X1   g03126(.A1(new_n2718_), .A2(new_n2770_), .ZN(new_n3191_));
  AOI21_X1   g03127(.A1(new_n2760_), .A2(new_n2761_), .B(new_n2769_), .ZN(new_n3192_));
  NAND4_X1   g03128(.A1(new_n3188_), .A2(new_n3190_), .A3(new_n3191_), .A4(new_n3192_), .ZN(new_n3193_));
  NOR4_X1    g03129(.A1(new_n147_), .A2(new_n190_), .A3(new_n460_), .A4(new_n718_), .ZN(new_n3194_));
  NAND2_X1   g03130(.A1(new_n790_), .A2(new_n508_), .ZN(new_n3195_));
  NOR4_X1    g03131(.A1(new_n2342_), .A2(new_n3194_), .A3(new_n1343_), .A4(new_n3195_), .ZN(new_n3196_));
  NOR4_X1    g03132(.A1(new_n1262_), .A2(new_n428_), .A3(new_n505_), .A4(new_n654_), .ZN(new_n3197_));
  INV_X1     g03133(.I(new_n517_), .ZN(new_n3198_));
  NAND3_X1   g03134(.A1(new_n233_), .A2(new_n3198_), .A3(new_n464_), .ZN(new_n3199_));
  NOR4_X1    g03135(.A1(new_n381_), .A2(new_n703_), .A3(new_n715_), .A4(new_n376_), .ZN(new_n3200_));
  NOR3_X1    g03136(.A1(new_n3197_), .A2(new_n3200_), .A3(new_n3199_), .ZN(new_n3201_));
  NOR3_X1    g03137(.A1(new_n3102_), .A2(new_n1264_), .A3(new_n1151_), .ZN(new_n3202_));
  INV_X1     g03138(.I(new_n454_), .ZN(new_n3203_));
  INV_X1     g03139(.I(new_n1319_), .ZN(new_n3204_));
  NOR4_X1    g03140(.A1(new_n3203_), .A2(new_n3204_), .A3(new_n1381_), .A4(new_n713_), .ZN(new_n3205_));
  NAND4_X1   g03141(.A1(new_n3202_), .A2(new_n3196_), .A3(new_n3205_), .A4(new_n3201_), .ZN(new_n3206_));
  NOR4_X1    g03142(.A1(new_n740_), .A2(new_n335_), .A3(new_n899_), .A4(new_n930_), .ZN(new_n3207_));
  INV_X1     g03143(.I(new_n3207_), .ZN(new_n3208_));
  NOR4_X1    g03144(.A1(new_n607_), .A2(new_n241_), .A3(new_n347_), .A4(new_n1146_), .ZN(new_n3209_));
  INV_X1     g03145(.I(new_n3209_), .ZN(new_n3210_));
  NOR3_X1    g03146(.A1(new_n936_), .A2(new_n170_), .A3(new_n306_), .ZN(new_n3211_));
  NAND4_X1   g03147(.A1(new_n3210_), .A2(new_n3208_), .A3(new_n2869_), .A4(new_n3211_), .ZN(new_n3212_));
  INV_X1     g03148(.I(new_n889_), .ZN(new_n3213_));
  NOR4_X1    g03149(.A1(new_n525_), .A2(new_n3213_), .A3(new_n400_), .A4(new_n730_), .ZN(new_n3214_));
  NOR4_X1    g03150(.A1(new_n289_), .A2(new_n482_), .A3(new_n437_), .A4(new_n736_), .ZN(new_n3215_));
  INV_X1     g03151(.I(new_n3215_), .ZN(new_n3216_));
  NOR2_X1    g03152(.A1(new_n788_), .A2(new_n684_), .ZN(new_n3217_));
  INV_X1     g03153(.I(new_n3217_), .ZN(new_n3218_));
  NOR3_X1    g03154(.A1(new_n3218_), .A2(new_n388_), .A3(new_n644_), .ZN(new_n3219_));
  INV_X1     g03155(.I(new_n1608_), .ZN(new_n3220_));
  NOR4_X1    g03156(.A1(new_n1149_), .A2(new_n343_), .A3(new_n574_), .A4(new_n1138_), .ZN(new_n3221_));
  INV_X1     g03157(.I(new_n3221_), .ZN(new_n3222_));
  NOR4_X1    g03158(.A1(new_n3222_), .A2(new_n1433_), .A3(new_n3220_), .A4(new_n2829_), .ZN(new_n3223_));
  NAND4_X1   g03159(.A1(new_n3223_), .A2(new_n3214_), .A3(new_n3216_), .A4(new_n3219_), .ZN(new_n3224_));
  OR3_X2     g03160(.A1(new_n3224_), .A2(new_n1966_), .A3(new_n3212_), .Z(new_n3225_));
  NOR2_X1    g03161(.A1(new_n3225_), .A2(new_n3206_), .ZN(new_n3226_));
  NOR2_X1    g03162(.A1(new_n3226_), .A2(\a[26] ), .ZN(new_n3227_));
  INV_X1     g03163(.I(new_n3226_), .ZN(new_n3228_));
  NOR2_X1    g03164(.A1(new_n3228_), .A2(new_n72_), .ZN(new_n3229_));
  NOR2_X1    g03165(.A1(new_n3229_), .A2(new_n3227_), .ZN(new_n3230_));
  NOR2_X1    g03166(.A1(new_n3230_), .A2(new_n2808_), .ZN(new_n3231_));
  XOR2_X1    g03167(.A1(new_n3226_), .A2(\a[26] ), .Z(new_n3232_));
  AOI21_X1   g03168(.A1(new_n2808_), .A2(new_n3232_), .B(new_n3231_), .ZN(new_n3233_));
  NAND2_X1   g03169(.A1(new_n3193_), .A2(new_n3233_), .ZN(new_n3234_));
  INV_X1     g03170(.I(new_n3234_), .ZN(new_n3235_));
  NOR2_X1    g03171(.A1(new_n3193_), .A2(new_n3233_), .ZN(new_n3236_));
  OAI21_X1   g03172(.A1(new_n3235_), .A2(new_n3236_), .B(new_n3184_), .ZN(new_n3237_));
  XNOR2_X1   g03173(.A1(new_n3193_), .A2(new_n3233_), .ZN(new_n3238_));
  OAI21_X1   g03174(.A1(new_n3184_), .A2(new_n3238_), .B(new_n3237_), .ZN(new_n3239_));
  INV_X1     g03175(.I(new_n3239_), .ZN(new_n3240_));
  NAND2_X1   g03176(.A1(new_n3181_), .A2(new_n3240_), .ZN(new_n3241_));
  NOR2_X1    g03177(.A1(new_n3181_), .A2(new_n3240_), .ZN(new_n3242_));
  INV_X1     g03178(.I(new_n3242_), .ZN(new_n3243_));
  AOI21_X1   g03179(.A1(new_n3243_), .A2(new_n3241_), .B(new_n3120_), .ZN(new_n3244_));
  XOR2_X1    g03180(.A1(new_n3181_), .A2(new_n3240_), .Z(new_n3245_));
  AOI21_X1   g03181(.A1(new_n3120_), .A2(new_n3245_), .B(new_n3244_), .ZN(new_n3246_));
  INV_X1     g03182(.I(new_n3142_), .ZN(new_n3247_));
  INV_X1     g03183(.I(new_n2729_), .ZN(new_n3248_));
  AOI21_X1   g03184(.A1(new_n2725_), .A2(new_n2726_), .B(new_n2727_), .ZN(new_n3249_));
  INV_X1     g03185(.I(new_n3249_), .ZN(new_n3250_));
  NAND2_X1   g03186(.A1(new_n3250_), .A2(new_n3248_), .ZN(new_n3251_));
  OAI21_X1   g03187(.A1(new_n3251_), .A2(new_n2716_), .B(new_n3176_), .ZN(new_n3252_));
  NAND2_X1   g03188(.A1(new_n3252_), .A2(new_n3247_), .ZN(new_n3253_));
  INV_X1     g03189(.I(new_n3253_), .ZN(new_n3254_));
  NOR2_X1    g03190(.A1(new_n71_), .A2(\a[23] ), .ZN(new_n3255_));
  NOR2_X1    g03191(.A1(new_n84_), .A2(\a[24] ), .ZN(new_n3256_));
  NOR2_X1    g03192(.A1(new_n3255_), .A2(new_n3256_), .ZN(new_n3257_));
  NOR2_X1    g03193(.A1(new_n470_), .A2(new_n99_), .ZN(new_n3258_));
  NOR2_X1    g03194(.A1(new_n3257_), .A2(new_n3258_), .ZN(new_n3259_));
  INV_X1     g03195(.I(new_n3259_), .ZN(new_n3260_));
  NOR2_X1    g03196(.A1(new_n84_), .A2(\a[26] ), .ZN(new_n3261_));
  NOR2_X1    g03197(.A1(new_n72_), .A2(\a[23] ), .ZN(new_n3262_));
  NOR2_X1    g03198(.A1(new_n84_), .A2(\a[25] ), .ZN(new_n3263_));
  NOR2_X1    g03199(.A1(new_n78_), .A2(\a[23] ), .ZN(new_n3264_));
  INV_X1     g03200(.I(new_n3257_), .ZN(new_n3265_));
  NOR3_X1    g03201(.A1(new_n3265_), .A2(new_n3263_), .A3(new_n3264_), .ZN(new_n3266_));
  NOR3_X1    g03202(.A1(new_n3266_), .A2(new_n3261_), .A3(new_n3262_), .ZN(new_n3267_));
  INV_X1     g03203(.I(new_n3267_), .ZN(new_n3268_));
  OAI22_X1   g03204(.A1(new_n3254_), .A2(new_n3260_), .B1(new_n3142_), .B2(new_n3268_), .ZN(new_n3269_));
  XOR2_X1    g03205(.A1(new_n3269_), .A2(new_n72_), .Z(new_n3270_));
  OAI21_X1   g03206(.A1(new_n3249_), .A2(new_n2729_), .B(new_n3170_), .ZN(new_n3271_));
  XOR2_X1    g03207(.A1(new_n3168_), .A2(new_n2728_), .Z(new_n3272_));
  OAI21_X1   g03208(.A1(new_n3251_), .A2(new_n3272_), .B(new_n3271_), .ZN(new_n3273_));
  OAI22_X1   g03209(.A1(new_n3176_), .A2(new_n3175_), .B1(new_n2665_), .B2(new_n2747_), .ZN(new_n3274_));
  INV_X1     g03210(.I(new_n2742_), .ZN(new_n3275_));
  NAND2_X1   g03211(.A1(new_n2728_), .A2(new_n3275_), .ZN(new_n3276_));
  AOI21_X1   g03212(.A1(new_n3274_), .A2(new_n3276_), .B(new_n2737_), .ZN(new_n3277_));
  NAND2_X1   g03213(.A1(new_n3273_), .A2(new_n3277_), .ZN(new_n3278_));
  XOR2_X1    g03214(.A1(new_n3278_), .A2(\a[29] ), .Z(new_n3279_));
  INV_X1     g03215(.I(new_n3279_), .ZN(new_n3280_));
  XOR2_X1    g03216(.A1(new_n3270_), .A2(new_n3280_), .Z(new_n3281_));
  INV_X1     g03217(.I(new_n3281_), .ZN(new_n3282_));
  XOR2_X1    g03218(.A1(new_n3116_), .A2(new_n3117_), .Z(new_n3283_));
  INV_X1     g03219(.I(new_n3119_), .ZN(new_n3284_));
  AOI21_X1   g03220(.A1(new_n3118_), .A2(new_n3284_), .B(new_n3068_), .ZN(new_n3285_));
  AOI21_X1   g03221(.A1(new_n3068_), .A2(new_n3283_), .B(new_n3285_), .ZN(new_n3286_));
  OAI21_X1   g03222(.A1(new_n3270_), .A2(new_n3286_), .B(new_n3282_), .ZN(new_n3287_));
  NAND2_X1   g03223(.A1(new_n3246_), .A2(new_n3287_), .ZN(new_n3288_));
  INV_X1     g03224(.I(new_n3288_), .ZN(new_n3289_));
  NOR2_X1    g03225(.A1(new_n3246_), .A2(new_n3287_), .ZN(new_n3290_));
  NOR2_X1    g03226(.A1(new_n3289_), .A2(new_n3290_), .ZN(new_n3291_));
  INV_X1     g03227(.I(new_n3291_), .ZN(new_n3292_));
  XOR2_X1    g03228(.A1(new_n3286_), .A2(new_n3269_), .Z(new_n3293_));
  XOR2_X1    g03229(.A1(new_n3293_), .A2(\a[26] ), .Z(new_n3294_));
  XOR2_X1    g03230(.A1(new_n3294_), .A2(new_n3280_), .Z(new_n3295_));
  INV_X1     g03231(.I(\a[21] ), .ZN(new_n3296_));
  NOR2_X1    g03232(.A1(new_n3296_), .A2(\a[20] ), .ZN(new_n3297_));
  NOR2_X1    g03233(.A1(new_n3035_), .A2(\a[21] ), .ZN(new_n3298_));
  NOR2_X1    g03234(.A1(new_n3297_), .A2(new_n3298_), .ZN(new_n3299_));
  XNOR2_X1   g03235(.A1(\a[22] ), .A2(\a[23] ), .ZN(new_n3300_));
  NOR2_X1    g03236(.A1(new_n3299_), .A2(new_n3300_), .ZN(new_n3301_));
  INV_X1     g03237(.I(new_n3301_), .ZN(new_n3302_));
  NOR2_X1    g03238(.A1(new_n3035_), .A2(\a[22] ), .ZN(new_n3303_));
  INV_X1     g03239(.I(\a[22] ), .ZN(new_n3304_));
  NOR3_X1    g03240(.A1(new_n3304_), .A2(\a[20] ), .A3(\a[21] ), .ZN(new_n3305_));
  AOI21_X1   g03241(.A1(\a[21] ), .A2(new_n3303_), .B(new_n3305_), .ZN(new_n3306_));
  INV_X1     g03242(.I(new_n3299_), .ZN(new_n3307_));
  XOR2_X1    g03243(.A1(\a[20] ), .A2(\a[22] ), .Z(new_n3308_));
  XNOR2_X1   g03244(.A1(\a[20] ), .A2(\a[23] ), .ZN(new_n3309_));
  OAI21_X1   g03245(.A1(new_n3307_), .A2(new_n3308_), .B(new_n3309_), .ZN(new_n3310_));
  OAI22_X1   g03246(.A1(new_n2614_), .A2(new_n3310_), .B1(new_n2665_), .B2(new_n3306_), .ZN(new_n3311_));
  NOR2_X1    g03247(.A1(new_n3307_), .A2(new_n3300_), .ZN(new_n3312_));
  NAND2_X1   g03248(.A1(new_n2728_), .A2(new_n3312_), .ZN(new_n3313_));
  AOI21_X1   g03249(.A1(new_n3313_), .A2(new_n3311_), .B(new_n3302_), .ZN(new_n3314_));
  NAND2_X1   g03250(.A1(new_n2733_), .A2(new_n3314_), .ZN(new_n3315_));
  XOR2_X1    g03251(.A1(new_n3315_), .A2(\a[23] ), .Z(new_n3316_));
  NOR2_X1    g03252(.A1(new_n3265_), .A2(new_n3258_), .ZN(new_n3317_));
  INV_X1     g03253(.I(new_n3317_), .ZN(new_n3318_));
  OAI22_X1   g03254(.A1(new_n2559_), .A2(new_n3268_), .B1(new_n694_), .B2(new_n3318_), .ZN(new_n3319_));
  NOR2_X1    g03255(.A1(new_n78_), .A2(\a[24] ), .ZN(new_n3320_));
  NOR2_X1    g03256(.A1(new_n84_), .A2(new_n71_), .ZN(new_n3321_));
  AOI22_X1   g03257(.A1(new_n3321_), .A2(new_n78_), .B1(new_n3320_), .B2(new_n84_), .ZN(new_n3322_));
  INV_X1     g03258(.I(new_n3322_), .ZN(new_n3323_));
  NAND2_X1   g03259(.A1(new_n2567_), .A2(new_n3323_), .ZN(new_n3324_));
  AOI21_X1   g03260(.A1(new_n3319_), .A2(new_n3324_), .B(new_n3260_), .ZN(new_n3325_));
  NAND2_X1   g03261(.A1(new_n2759_), .A2(new_n3325_), .ZN(new_n3326_));
  XOR2_X1    g03262(.A1(new_n3326_), .A2(\a[26] ), .Z(new_n3327_));
  XOR2_X1    g03263(.A1(new_n1121_), .A2(new_n1180_), .Z(new_n3328_));
  XNOR2_X1   g03264(.A1(new_n1121_), .A2(new_n1180_), .ZN(new_n3329_));
  MUX2_X1    g03265(.I0(new_n3328_), .I1(new_n3329_), .S(new_n2505_), .Z(new_n3330_));
  NAND2_X1   g03266(.A1(new_n1122_), .A2(new_n3189_), .ZN(new_n3331_));
  INV_X1     g03267(.I(new_n2772_), .ZN(new_n3332_));
  AOI22_X1   g03268(.A1(new_n2496_), .A2(new_n2770_), .B1(new_n1181_), .B2(new_n3332_), .ZN(new_n3333_));
  NAND4_X1   g03269(.A1(new_n3330_), .A2(new_n2764_), .A3(new_n3331_), .A4(new_n3333_), .ZN(new_n3334_));
  NOR4_X1    g03270(.A1(new_n415_), .A2(new_n333_), .A3(new_n420_), .A4(new_n817_), .ZN(new_n3335_));
  NOR4_X1    g03271(.A1(new_n294_), .A2(new_n498_), .A3(new_n719_), .A4(new_n449_), .ZN(new_n3336_));
  NOR3_X1    g03272(.A1(new_n617_), .A2(new_n268_), .A3(new_n1531_), .ZN(new_n3337_));
  INV_X1     g03273(.I(new_n3337_), .ZN(new_n3338_));
  NOR4_X1    g03274(.A1(new_n3338_), .A2(new_n571_), .A3(new_n3335_), .A4(new_n3336_), .ZN(new_n3339_));
  NAND2_X1   g03275(.A1(new_n641_), .A2(new_n649_), .ZN(new_n3340_));
  NOR4_X1    g03276(.A1(new_n1278_), .A2(new_n1055_), .A3(new_n3340_), .A4(new_n2270_), .ZN(new_n3341_));
  NOR4_X1    g03277(.A1(new_n1206_), .A2(new_n2234_), .A3(new_n782_), .A4(new_n280_), .ZN(new_n3342_));
  INV_X1     g03278(.I(new_n2398_), .ZN(new_n3343_));
  NOR4_X1    g03279(.A1(new_n172_), .A2(new_n591_), .A3(new_n482_), .A4(new_n1236_), .ZN(new_n3344_));
  NOR4_X1    g03280(.A1(new_n3343_), .A2(new_n3344_), .A3(new_n81_), .A4(new_n267_), .ZN(new_n3345_));
  NAND4_X1   g03281(.A1(new_n3341_), .A2(new_n3339_), .A3(new_n3342_), .A4(new_n3345_), .ZN(new_n3346_));
  NOR4_X1    g03282(.A1(new_n541_), .A2(new_n203_), .A3(new_n910_), .A4(new_n736_), .ZN(new_n3347_));
  NOR4_X1    g03283(.A1(new_n1984_), .A2(new_n398_), .A3(new_n487_), .A4(new_n772_), .ZN(new_n3348_));
  NOR4_X1    g03284(.A1(new_n1262_), .A2(new_n556_), .A3(new_n902_), .A4(new_n310_), .ZN(new_n3349_));
  NOR3_X1    g03285(.A1(new_n3213_), .A2(new_n1175_), .A3(new_n211_), .ZN(new_n3350_));
  INV_X1     g03286(.I(new_n3350_), .ZN(new_n3351_));
  NOR4_X1    g03287(.A1(new_n3351_), .A2(new_n3347_), .A3(new_n3348_), .A4(new_n3349_), .ZN(new_n3352_));
  INV_X1     g03288(.I(new_n2245_), .ZN(new_n3353_));
  NAND3_X1   g03289(.A1(new_n765_), .A2(new_n1424_), .A3(new_n1923_), .ZN(new_n3354_));
  NOR4_X1    g03290(.A1(new_n3354_), .A2(new_n1198_), .A3(new_n2092_), .A4(new_n3353_), .ZN(new_n3355_));
  NAND3_X1   g03291(.A1(new_n3352_), .A2(new_n532_), .A3(new_n3355_), .ZN(new_n3356_));
  NOR3_X1    g03292(.A1(new_n3346_), .A2(new_n2526_), .A3(new_n3356_), .ZN(new_n3357_));
  INV_X1     g03293(.I(new_n750_), .ZN(new_n3358_));
  NAND2_X1   g03294(.A1(new_n438_), .A2(new_n1395_), .ZN(new_n3359_));
  NOR4_X1    g03295(.A1(new_n865_), .A2(new_n1116_), .A3(new_n3359_), .A4(new_n956_), .ZN(new_n3360_));
  NOR4_X1    g03296(.A1(new_n415_), .A2(new_n714_), .A3(new_n736_), .A4(new_n796_), .ZN(new_n3361_));
  NOR4_X1    g03297(.A1(new_n203_), .A2(new_n226_), .A3(new_n491_), .A4(new_n286_), .ZN(new_n3362_));
  NOR2_X1    g03298(.A1(new_n3361_), .A2(new_n3362_), .ZN(new_n3363_));
  NAND2_X1   g03299(.A1(new_n3360_), .A2(new_n3363_), .ZN(new_n3364_));
  NOR2_X1    g03300(.A1(new_n267_), .A2(new_n420_), .ZN(new_n3365_));
  NAND4_X1   g03301(.A1(new_n3365_), .A2(new_n1497_), .A3(new_n1700_), .A4(new_n2040_), .ZN(new_n3366_));
  NOR4_X1    g03302(.A1(new_n3364_), .A2(new_n2068_), .A3(new_n3358_), .A4(new_n3366_), .ZN(new_n3367_));
  NOR2_X1    g03303(.A1(new_n2629_), .A2(new_n1737_), .ZN(new_n3368_));
  NAND3_X1   g03304(.A1(new_n623_), .A2(new_n3367_), .A3(new_n3368_), .ZN(new_n3369_));
  INV_X1     g03305(.I(new_n3369_), .ZN(new_n3370_));
  OAI21_X1   g03306(.A1(new_n3370_), .A2(\a[17] ), .B(new_n3357_), .ZN(new_n3371_));
  INV_X1     g03307(.I(\a[17] ), .ZN(new_n3372_));
  NOR2_X1    g03308(.A1(new_n3369_), .A2(new_n3372_), .ZN(new_n3373_));
  INV_X1     g03309(.I(new_n3373_), .ZN(new_n3374_));
  AOI21_X1   g03310(.A1(new_n3371_), .A2(new_n3374_), .B(new_n3032_), .ZN(new_n3375_));
  NAND2_X1   g03311(.A1(new_n3371_), .A2(new_n3374_), .ZN(new_n3376_));
  NOR2_X1    g03312(.A1(new_n3376_), .A2(new_n3031_), .ZN(new_n3377_));
  NOR2_X1    g03313(.A1(new_n3377_), .A2(new_n3375_), .ZN(new_n3378_));
  NOR2_X1    g03314(.A1(new_n3334_), .A2(new_n3378_), .ZN(new_n3379_));
  XOR2_X1    g03315(.A1(new_n3376_), .A2(new_n3032_), .Z(new_n3380_));
  INV_X1     g03316(.I(new_n3380_), .ZN(new_n3381_));
  AOI21_X1   g03317(.A1(new_n3334_), .A2(new_n3381_), .B(new_n3379_), .ZN(new_n3382_));
  OAI22_X1   g03318(.A1(new_n813_), .A2(new_n3175_), .B1(new_n1008_), .B2(new_n2747_), .ZN(new_n3383_));
  NAND2_X1   g03319(.A1(new_n897_), .A2(new_n3275_), .ZN(new_n3384_));
  AOI21_X1   g03320(.A1(new_n3383_), .A2(new_n3384_), .B(new_n2737_), .ZN(new_n3385_));
  NAND2_X1   g03321(.A1(new_n2917_), .A2(new_n3385_), .ZN(new_n3386_));
  XOR2_X1    g03322(.A1(new_n3386_), .A2(\a[29] ), .Z(new_n3387_));
  XNOR2_X1   g03323(.A1(new_n1121_), .A2(new_n2492_), .ZN(new_n3388_));
  AOI21_X1   g03324(.A1(new_n2495_), .A2(new_n2498_), .B(new_n3388_), .ZN(new_n3389_));
  NAND2_X1   g03325(.A1(new_n2495_), .A2(new_n2498_), .ZN(new_n3390_));
  NOR2_X1    g03326(.A1(new_n2501_), .A2(new_n2499_), .ZN(new_n3391_));
  NOR2_X1    g03327(.A1(new_n3390_), .A2(new_n3391_), .ZN(new_n3392_));
  OR2_X2     g03328(.A1(new_n3392_), .A2(new_n3389_), .Z(new_n3393_));
  OAI21_X1   g03329(.A1(new_n2451_), .A2(new_n2771_), .B(new_n2764_), .ZN(new_n3394_));
  OAI22_X1   g03330(.A1(new_n1121_), .A2(new_n2772_), .B1(new_n2492_), .B2(new_n2767_), .ZN(new_n3395_));
  NOR2_X1    g03331(.A1(new_n3394_), .A2(new_n3395_), .ZN(new_n3396_));
  AND2_X2    g03332(.A1(new_n3393_), .A2(new_n3396_), .Z(new_n3397_));
  NAND2_X1   g03333(.A1(new_n2411_), .A2(new_n2414_), .ZN(new_n3398_));
  XNOR2_X1   g03334(.A1(new_n2451_), .A2(new_n2408_), .ZN(new_n3399_));
  INV_X1     g03335(.I(new_n3399_), .ZN(new_n3400_));
  NAND2_X1   g03336(.A1(new_n3398_), .A2(new_n3400_), .ZN(new_n3401_));
  NOR2_X1    g03337(.A1(new_n2455_), .A2(new_n2452_), .ZN(new_n3402_));
  OAI21_X1   g03338(.A1(new_n3398_), .A2(new_n3402_), .B(new_n3401_), .ZN(new_n3403_));
  OAI21_X1   g03339(.A1(new_n2408_), .A2(new_n2767_), .B(new_n2764_), .ZN(new_n3404_));
  OAI22_X1   g03340(.A1(new_n2367_), .A2(new_n2771_), .B1(new_n2451_), .B2(new_n2772_), .ZN(new_n3405_));
  NOR2_X1    g03341(.A1(new_n3405_), .A2(new_n3404_), .ZN(new_n3406_));
  NAND2_X1   g03342(.A1(new_n3403_), .A2(new_n3406_), .ZN(new_n3407_));
  NOR3_X1    g03343(.A1(new_n1262_), .A2(new_n548_), .A3(new_n459_), .ZN(new_n3408_));
  NOR3_X1    g03344(.A1(new_n1043_), .A2(new_n324_), .A3(new_n510_), .ZN(new_n3409_));
  NOR3_X1    g03345(.A1(new_n590_), .A2(new_n428_), .A3(new_n474_), .ZN(new_n3410_));
  NAND4_X1   g03346(.A1(new_n3409_), .A2(new_n3024_), .A3(new_n3408_), .A4(new_n3410_), .ZN(new_n3411_));
  NAND2_X1   g03347(.A1(new_n405_), .A2(new_n383_), .ZN(new_n3412_));
  NOR4_X1    g03348(.A1(new_n2232_), .A2(new_n1730_), .A3(new_n3412_), .A4(new_n1079_), .ZN(new_n3413_));
  NAND3_X1   g03349(.A1(new_n1660_), .A2(new_n2124_), .A3(new_n3413_), .ZN(new_n3414_));
  NOR3_X1    g03350(.A1(new_n3414_), .A2(new_n2049_), .A3(new_n3411_), .ZN(new_n3415_));
  NAND2_X1   g03351(.A1(new_n1601_), .A2(new_n1059_), .ZN(new_n3416_));
  NOR4_X1    g03352(.A1(new_n2023_), .A2(new_n2234_), .A3(new_n3416_), .A4(new_n299_), .ZN(new_n3417_));
  NOR2_X1    g03353(.A1(new_n1808_), .A2(new_n491_), .ZN(new_n3418_));
  INV_X1     g03354(.I(new_n3418_), .ZN(new_n3419_));
  NOR4_X1    g03355(.A1(new_n593_), .A2(new_n703_), .A3(new_n191_), .A4(new_n310_), .ZN(new_n3420_));
  NOR4_X1    g03356(.A1(new_n267_), .A2(new_n398_), .A3(new_n731_), .A4(new_n430_), .ZN(new_n3421_));
  NOR4_X1    g03357(.A1(new_n1777_), .A2(new_n3419_), .A3(new_n3420_), .A4(new_n3421_), .ZN(new_n3422_));
  NAND4_X1   g03358(.A1(new_n951_), .A2(new_n1651_), .A3(new_n3417_), .A4(new_n3422_), .ZN(new_n3423_));
  NOR3_X1    g03359(.A1(new_n573_), .A2(new_n396_), .A3(new_n930_), .ZN(new_n3424_));
  NOR2_X1    g03360(.A1(new_n1614_), .A2(new_n730_), .ZN(new_n3425_));
  NAND4_X1   g03361(.A1(new_n3425_), .A2(new_n1472_), .A3(new_n1738_), .A4(new_n3424_), .ZN(new_n3426_));
  NOR4_X1    g03362(.A1(new_n2439_), .A2(new_n252_), .A3(new_n294_), .A4(new_n574_), .ZN(new_n3427_));
  INV_X1     g03363(.I(new_n3427_), .ZN(new_n3428_));
  NAND4_X1   g03364(.A1(new_n1335_), .A2(new_n293_), .A3(new_n564_), .A4(new_n1095_), .ZN(new_n3429_));
  NAND4_X1   g03365(.A1(new_n313_), .A2(new_n1605_), .A3(new_n1066_), .A4(new_n1393_), .ZN(new_n3430_));
  NAND4_X1   g03366(.A1(new_n631_), .A2(new_n3099_), .A3(new_n524_), .A4(new_n1690_), .ZN(new_n3431_));
  NOR2_X1    g03367(.A1(new_n2180_), .A2(new_n3431_), .ZN(new_n3432_));
  NAND4_X1   g03368(.A1(new_n3432_), .A2(new_n3428_), .A3(new_n3429_), .A4(new_n3430_), .ZN(new_n3433_));
  NOR3_X1    g03369(.A1(new_n3423_), .A2(new_n3426_), .A3(new_n3433_), .ZN(new_n3434_));
  NAND2_X1   g03370(.A1(new_n3434_), .A2(new_n3415_), .ZN(new_n3435_));
  NOR4_X1    g03371(.A1(new_n3218_), .A2(new_n238_), .A3(new_n485_), .A4(new_n1152_), .ZN(new_n3436_));
  NOR4_X1    g03372(.A1(new_n226_), .A2(new_n304_), .A3(new_n837_), .A4(new_n261_), .ZN(new_n3437_));
  NOR3_X1    g03373(.A1(new_n1988_), .A2(new_n496_), .A3(new_n505_), .ZN(new_n3438_));
  NOR3_X1    g03374(.A1(new_n3351_), .A2(new_n3437_), .A3(new_n3438_), .ZN(new_n3439_));
  AND2_X2    g03375(.A1(new_n3439_), .A2(new_n3436_), .Z(new_n3440_));
  NOR4_X1    g03376(.A1(new_n912_), .A2(new_n2042_), .A3(new_n164_), .A4(new_n320_), .ZN(new_n3441_));
  NOR4_X1    g03377(.A1(new_n593_), .A2(new_n202_), .A3(new_n577_), .A4(new_n902_), .ZN(new_n3442_));
  NOR4_X1    g03378(.A1(new_n241_), .A2(new_n610_), .A3(new_n1236_), .A4(new_n517_), .ZN(new_n3443_));
  NOR3_X1    g03379(.A1(new_n3442_), .A2(new_n3427_), .A3(new_n3443_), .ZN(new_n3444_));
  NAND4_X1   g03380(.A1(new_n3440_), .A2(new_n679_), .A3(new_n3441_), .A4(new_n3444_), .ZN(new_n3445_));
  INV_X1     g03381(.I(new_n3445_), .ZN(new_n3446_));
  NOR2_X1    g03382(.A1(new_n359_), .A2(new_n459_), .ZN(new_n3447_));
  NAND4_X1   g03383(.A1(new_n775_), .A2(new_n1354_), .A3(new_n1159_), .A4(new_n3447_), .ZN(new_n3448_));
  NOR4_X1    g03384(.A1(new_n147_), .A2(new_n403_), .A3(new_n420_), .A4(new_n1168_), .ZN(new_n3449_));
  NOR2_X1    g03385(.A1(new_n584_), .A2(new_n227_), .ZN(new_n3450_));
  NOR2_X1    g03386(.A1(new_n644_), .A2(new_n102_), .ZN(new_n3451_));
  AOI21_X1   g03387(.A1(new_n3450_), .A2(new_n3451_), .B(new_n3449_), .ZN(new_n3452_));
  INV_X1     g03388(.I(new_n3452_), .ZN(new_n3453_));
  NOR4_X1    g03389(.A1(new_n1048_), .A2(new_n906_), .A3(new_n770_), .A4(new_n172_), .ZN(new_n3454_));
  NOR4_X1    g03390(.A1(new_n3454_), .A2(new_n347_), .A3(new_n518_), .A4(new_n544_), .ZN(new_n3455_));
  INV_X1     g03391(.I(new_n3455_), .ZN(new_n3456_));
  NAND4_X1   g03392(.A1(new_n1657_), .A2(new_n399_), .A3(new_n646_), .A4(new_n1111_), .ZN(new_n3457_));
  NOR4_X1    g03393(.A1(new_n3457_), .A2(new_n3456_), .A3(new_n3448_), .A4(new_n3453_), .ZN(new_n3458_));
  NOR2_X1    g03394(.A1(new_n381_), .A2(new_n681_), .ZN(new_n3459_));
  INV_X1     g03395(.I(new_n3459_), .ZN(new_n3460_));
  NOR4_X1    g03396(.A1(new_n3460_), .A2(new_n3353_), .A3(new_n594_), .A4(new_n718_), .ZN(new_n3461_));
  INV_X1     g03397(.I(new_n3461_), .ZN(new_n3462_));
  NOR4_X1    g03398(.A1(new_n256_), .A2(new_n437_), .A3(new_n721_), .A4(new_n776_), .ZN(new_n3463_));
  NOR4_X1    g03399(.A1(new_n3462_), .A2(new_n1203_), .A3(new_n1648_), .A4(new_n3463_), .ZN(new_n3464_));
  NAND2_X1   g03400(.A1(new_n1816_), .A2(new_n1058_), .ZN(new_n3465_));
  NAND2_X1   g03401(.A1(new_n1601_), .A2(new_n572_), .ZN(new_n3466_));
  NOR4_X1    g03402(.A1(new_n2261_), .A2(new_n596_), .A3(new_n3465_), .A4(new_n3466_), .ZN(new_n3467_));
  NAND3_X1   g03403(.A1(new_n483_), .A2(new_n871_), .A3(new_n809_), .ZN(new_n3468_));
  INV_X1     g03404(.I(new_n3468_), .ZN(new_n3469_));
  INV_X1     g03405(.I(new_n1318_), .ZN(new_n3470_));
  NOR2_X1    g03406(.A1(new_n3470_), .A2(new_n1264_), .ZN(new_n3471_));
  NOR3_X1    g03407(.A1(new_n76_), .A2(new_n648_), .A3(new_n556_), .ZN(new_n3472_));
  NOR3_X1    g03408(.A1(new_n2306_), .A2(new_n282_), .A3(new_n428_), .ZN(new_n3473_));
  NAND4_X1   g03409(.A1(new_n3471_), .A2(new_n2657_), .A3(new_n3472_), .A4(new_n3473_), .ZN(new_n3474_));
  NOR4_X1    g03410(.A1(new_n3474_), .A2(new_n567_), .A3(new_n2420_), .A4(new_n3469_), .ZN(new_n3475_));
  AND3_X2    g03411(.A1(new_n3475_), .A2(new_n3464_), .A3(new_n3467_), .Z(new_n3476_));
  NAND3_X1   g03412(.A1(new_n3446_), .A2(new_n3458_), .A3(new_n3476_), .ZN(new_n3477_));
  INV_X1     g03413(.I(new_n3477_), .ZN(new_n3478_));
  INV_X1     g03414(.I(new_n1772_), .ZN(new_n3479_));
  NOR3_X1    g03415(.A1(new_n172_), .A2(new_n307_), .A3(new_n190_), .ZN(new_n3480_));
  NAND4_X1   g03416(.A1(new_n1222_), .A2(new_n3198_), .A3(new_n110_), .A4(new_n808_), .ZN(new_n3481_));
  NAND4_X1   g03417(.A1(new_n3479_), .A2(new_n3481_), .A3(new_n1474_), .A4(new_n3480_), .ZN(new_n3482_));
  NOR4_X1    g03418(.A1(new_n343_), .A2(new_n898_), .A3(new_n262_), .A4(new_n1531_), .ZN(new_n3483_));
  NOR2_X1    g03419(.A1(new_n106_), .A2(new_n255_), .ZN(new_n3484_));
  INV_X1     g03420(.I(new_n3484_), .ZN(new_n3485_));
  NOR3_X1    g03421(.A1(new_n3483_), .A2(new_n3485_), .A3(new_n865_), .ZN(new_n3486_));
  INV_X1     g03422(.I(new_n3486_), .ZN(new_n3487_));
  NOR4_X1    g03423(.A1(new_n541_), .A2(new_n534_), .A3(new_n225_), .A4(new_n804_), .ZN(new_n3488_));
  NOR2_X1    g03424(.A1(new_n2441_), .A2(new_n3488_), .ZN(new_n3489_));
  NAND4_X1   g03425(.A1(new_n3489_), .A2(new_n629_), .A3(new_n2091_), .A4(new_n1329_), .ZN(new_n3490_));
  NOR4_X1    g03426(.A1(new_n3490_), .A2(new_n3487_), .A3(new_n3426_), .A4(new_n3482_), .ZN(new_n3491_));
  NOR4_X1    g03427(.A1(new_n495_), .A2(new_n281_), .A3(new_n817_), .A4(new_n306_), .ZN(new_n3492_));
  NOR3_X1    g03428(.A1(new_n666_), .A2(new_n264_), .A3(new_n359_), .ZN(new_n3493_));
  NAND2_X1   g03429(.A1(new_n3493_), .A2(new_n3410_), .ZN(new_n3494_));
  NOR2_X1    g03430(.A1(new_n3494_), .A2(new_n3492_), .ZN(new_n3495_));
  NAND3_X1   g03431(.A1(new_n795_), .A2(new_n985_), .A3(new_n1935_), .ZN(new_n3496_));
  NOR4_X1    g03432(.A1(new_n214_), .A2(new_n239_), .A3(new_n841_), .A4(new_n749_), .ZN(new_n3497_));
  NOR4_X1    g03433(.A1(new_n2447_), .A2(new_n1962_), .A3(new_n3496_), .A4(new_n3497_), .ZN(new_n3498_));
  NAND4_X1   g03434(.A1(new_n3498_), .A2(new_n1809_), .A3(new_n2552_), .A4(new_n3495_), .ZN(new_n3499_));
  NOR4_X1    g03435(.A1(new_n2482_), .A2(new_n406_), .A3(new_n561_), .A4(new_n1915_), .ZN(new_n3500_));
  NOR2_X1    g03436(.A1(new_n2647_), .A2(new_n98_), .ZN(new_n3501_));
  INV_X1     g03437(.I(new_n420_), .ZN(new_n3502_));
  NAND4_X1   g03438(.A1(new_n3502_), .A2(new_n469_), .A3(new_n373_), .A4(new_n551_), .ZN(new_n3503_));
  NAND4_X1   g03439(.A1(new_n612_), .A2(new_n311_), .A3(new_n1100_), .A4(new_n1605_), .ZN(new_n3504_));
  NAND4_X1   g03440(.A1(new_n3500_), .A2(new_n3501_), .A3(new_n3503_), .A4(new_n3504_), .ZN(new_n3505_));
  NOR3_X1    g03441(.A1(new_n288_), .A2(new_n753_), .A3(new_n413_), .ZN(new_n3506_));
  NOR3_X1    g03442(.A1(new_n247_), .A2(new_n584_), .A3(new_n660_), .ZN(new_n3507_));
  NAND4_X1   g03443(.A1(new_n2079_), .A2(new_n1923_), .A3(new_n3506_), .A4(new_n3507_), .ZN(new_n3508_));
  NAND4_X1   g03444(.A1(new_n295_), .A2(new_n1396_), .A3(new_n984_), .A4(new_n80_), .ZN(new_n3509_));
  NOR3_X1    g03445(.A1(new_n505_), .A2(new_n779_), .A3(new_n837_), .ZN(new_n3510_));
  NOR2_X1    g03446(.A1(new_n1048_), .A2(new_n453_), .ZN(new_n3511_));
  INV_X1     g03447(.I(new_n3511_), .ZN(new_n3512_));
  NAND4_X1   g03448(.A1(new_n1668_), .A2(new_n631_), .A3(new_n509_), .A4(new_n1468_), .ZN(new_n3513_));
  NOR4_X1    g03449(.A1(new_n3513_), .A2(new_n3512_), .A3(new_n1183_), .A4(new_n650_), .ZN(new_n3514_));
  NAND4_X1   g03450(.A1(new_n3514_), .A2(new_n3009_), .A3(new_n3509_), .A4(new_n3510_), .ZN(new_n3515_));
  NOR4_X1    g03451(.A1(new_n3499_), .A2(new_n3505_), .A3(new_n3508_), .A4(new_n3515_), .ZN(new_n3516_));
  NAND2_X1   g03452(.A1(new_n3516_), .A2(new_n3491_), .ZN(new_n3517_));
  INV_X1     g03453(.I(new_n3517_), .ZN(new_n3518_));
  NOR2_X1    g03454(.A1(new_n3518_), .A2(\a[14] ), .ZN(new_n3519_));
  INV_X1     g03455(.I(new_n3519_), .ZN(new_n3520_));
  INV_X1     g03456(.I(\a[14] ), .ZN(new_n3521_));
  NOR2_X1    g03457(.A1(new_n3517_), .A2(new_n3521_), .ZN(new_n3522_));
  AOI21_X1   g03458(.A1(new_n3520_), .A2(new_n3478_), .B(new_n3522_), .ZN(new_n3523_));
  INV_X1     g03459(.I(new_n3523_), .ZN(new_n3524_));
  NOR2_X1    g03460(.A1(new_n3524_), .A2(new_n3435_), .ZN(new_n3525_));
  NAND2_X1   g03461(.A1(new_n3524_), .A2(new_n3435_), .ZN(new_n3526_));
  OAI21_X1   g03462(.A1(new_n3407_), .A2(new_n3525_), .B(new_n3526_), .ZN(new_n3527_));
  INV_X1     g03463(.I(new_n3435_), .ZN(new_n3528_));
  NOR2_X1    g03464(.A1(new_n3528_), .A2(new_n3369_), .ZN(new_n3529_));
  INV_X1     g03465(.I(new_n3529_), .ZN(new_n3530_));
  NOR2_X1    g03466(.A1(new_n3370_), .A2(new_n3435_), .ZN(new_n3531_));
  AOI21_X1   g03467(.A1(new_n3527_), .A2(new_n3530_), .B(new_n3531_), .ZN(new_n3532_));
  INV_X1     g03468(.I(new_n3532_), .ZN(new_n3533_));
  NOR2_X1    g03469(.A1(new_n3370_), .A2(\a[17] ), .ZN(new_n3534_));
  NOR2_X1    g03470(.A1(new_n3534_), .A2(new_n3373_), .ZN(new_n3535_));
  INV_X1     g03471(.I(new_n3535_), .ZN(new_n3536_));
  XOR2_X1    g03472(.A1(new_n3369_), .A2(\a[17] ), .Z(new_n3537_));
  NOR2_X1    g03473(.A1(new_n3537_), .A2(new_n3357_), .ZN(new_n3538_));
  AOI21_X1   g03474(.A1(new_n3357_), .A2(new_n3536_), .B(new_n3538_), .ZN(new_n3539_));
  INV_X1     g03475(.I(new_n3539_), .ZN(new_n3540_));
  NOR2_X1    g03476(.A1(new_n3533_), .A2(new_n3540_), .ZN(new_n3541_));
  INV_X1     g03477(.I(new_n3541_), .ZN(new_n3542_));
  NOR2_X1    g03478(.A1(new_n3532_), .A2(new_n3539_), .ZN(new_n3543_));
  AOI21_X1   g03479(.A1(new_n3542_), .A2(new_n3397_), .B(new_n3543_), .ZN(new_n3544_));
  INV_X1     g03480(.I(new_n3544_), .ZN(new_n3545_));
  XOR2_X1    g03481(.A1(new_n3387_), .A2(new_n3545_), .Z(new_n3546_));
  NOR2_X1    g03482(.A1(new_n3546_), .A2(new_n3382_), .ZN(new_n3547_));
  INV_X1     g03483(.I(new_n3382_), .ZN(new_n3548_));
  AND2_X2    g03484(.A1(new_n3387_), .A2(new_n3544_), .Z(new_n3549_));
  NOR2_X1    g03485(.A1(new_n3387_), .A2(new_n3544_), .ZN(new_n3550_));
  NOR2_X1    g03486(.A1(new_n3549_), .A2(new_n3550_), .ZN(new_n3551_));
  NOR2_X1    g03487(.A1(new_n3551_), .A2(new_n3548_), .ZN(new_n3552_));
  NOR2_X1    g03488(.A1(new_n3552_), .A2(new_n3547_), .ZN(new_n3553_));
  NOR3_X1    g03489(.A1(new_n2500_), .A2(new_n1181_), .A3(new_n2501_), .ZN(new_n3554_));
  INV_X1     g03490(.I(new_n3554_), .ZN(new_n3555_));
  OAI21_X1   g03491(.A1(new_n2500_), .A2(new_n2501_), .B(new_n1181_), .ZN(new_n3556_));
  NAND2_X1   g03492(.A1(new_n3555_), .A2(new_n3556_), .ZN(new_n3557_));
  NAND3_X1   g03493(.A1(new_n3557_), .A2(new_n2504_), .A3(new_n3328_), .ZN(new_n3558_));
  INV_X1     g03494(.I(new_n3556_), .ZN(new_n3559_));
  OAI21_X1   g03495(.A1(new_n3559_), .A2(new_n3554_), .B(new_n3328_), .ZN(new_n3560_));
  NAND2_X1   g03496(.A1(new_n3560_), .A2(new_n1008_), .ZN(new_n3561_));
  NAND2_X1   g03497(.A1(new_n3561_), .A2(new_n3558_), .ZN(new_n3562_));
  OAI22_X1   g03498(.A1(new_n1008_), .A2(new_n3175_), .B1(new_n1121_), .B2(new_n2747_), .ZN(new_n3563_));
  NAND2_X1   g03499(.A1(new_n1181_), .A2(new_n3275_), .ZN(new_n3564_));
  AOI21_X1   g03500(.A1(new_n3563_), .A2(new_n3564_), .B(new_n2737_), .ZN(new_n3565_));
  NAND2_X1   g03501(.A1(new_n3562_), .A2(new_n3565_), .ZN(new_n3566_));
  XOR2_X1    g03502(.A1(new_n3566_), .A2(\a[29] ), .Z(new_n3567_));
  INV_X1     g03503(.I(new_n3567_), .ZN(new_n3568_));
  OAI21_X1   g03504(.A1(new_n3529_), .A2(new_n3531_), .B(new_n3527_), .ZN(new_n3569_));
  XOR2_X1    g03505(.A1(new_n3435_), .A2(new_n3369_), .Z(new_n3570_));
  OAI21_X1   g03506(.A1(new_n3527_), .A2(new_n3570_), .B(new_n3569_), .ZN(new_n3571_));
  NOR2_X1    g03507(.A1(new_n2453_), .A2(new_n2455_), .ZN(new_n3572_));
  XNOR2_X1   g03508(.A1(new_n2492_), .A2(new_n2451_), .ZN(new_n3573_));
  NOR2_X1    g03509(.A1(new_n3572_), .A2(new_n3573_), .ZN(new_n3574_));
  NOR2_X1    g03510(.A1(new_n2497_), .A2(new_n2493_), .ZN(new_n3575_));
  NOR3_X1    g03511(.A1(new_n2453_), .A2(new_n2455_), .A3(new_n3575_), .ZN(new_n3576_));
  OR2_X2     g03512(.A1(new_n3574_), .A2(new_n3576_), .Z(new_n3577_));
  NOR2_X1    g03513(.A1(new_n2408_), .A2(new_n2771_), .ZN(new_n3578_));
  INV_X1     g03514(.I(new_n3578_), .ZN(new_n3579_));
  AOI22_X1   g03515(.A1(new_n2496_), .A2(new_n3332_), .B1(new_n2454_), .B2(new_n3189_), .ZN(new_n3580_));
  NAND4_X1   g03516(.A1(new_n3577_), .A2(new_n2764_), .A3(new_n3579_), .A4(new_n3580_), .ZN(new_n3581_));
  INV_X1     g03517(.I(new_n3581_), .ZN(new_n3582_));
  NOR2_X1    g03518(.A1(new_n3571_), .A2(new_n3582_), .ZN(new_n3583_));
  INV_X1     g03519(.I(new_n3583_), .ZN(new_n3584_));
  NAND2_X1   g03520(.A1(new_n3568_), .A2(new_n3584_), .ZN(new_n3585_));
  NAND2_X1   g03521(.A1(new_n3571_), .A2(new_n3582_), .ZN(new_n3586_));
  NAND2_X1   g03522(.A1(new_n3585_), .A2(new_n3586_), .ZN(new_n3587_));
  INV_X1     g03523(.I(new_n3587_), .ZN(new_n3588_));
  INV_X1     g03524(.I(new_n3397_), .ZN(new_n3589_));
  XOR2_X1    g03525(.A1(new_n3532_), .A2(new_n3540_), .Z(new_n3590_));
  OAI21_X1   g03526(.A1(new_n3541_), .A2(new_n3543_), .B(new_n3589_), .ZN(new_n3591_));
  OAI21_X1   g03527(.A1(new_n3589_), .A2(new_n3590_), .B(new_n3591_), .ZN(new_n3592_));
  XOR2_X1    g03528(.A1(new_n1008_), .A2(new_n896_), .Z(new_n3593_));
  INV_X1     g03529(.I(new_n3593_), .ZN(new_n3594_));
  NAND2_X1   g03530(.A1(new_n2509_), .A2(new_n3594_), .ZN(new_n3595_));
  OAI21_X1   g03531(.A1(new_n2509_), .A2(new_n2911_), .B(new_n3595_), .ZN(new_n3596_));
  OAI22_X1   g03532(.A1(new_n896_), .A2(new_n3175_), .B1(new_n1180_), .B2(new_n2747_), .ZN(new_n3597_));
  NAND2_X1   g03533(.A1(new_n2504_), .A2(new_n3275_), .ZN(new_n3598_));
  AOI21_X1   g03534(.A1(new_n3598_), .A2(new_n3597_), .B(new_n2737_), .ZN(new_n3599_));
  NAND2_X1   g03535(.A1(new_n3596_), .A2(new_n3599_), .ZN(new_n3600_));
  XOR2_X1    g03536(.A1(new_n3600_), .A2(\a[29] ), .Z(new_n3601_));
  AND2_X2    g03537(.A1(new_n3601_), .A2(new_n3592_), .Z(new_n3602_));
  NOR2_X1    g03538(.A1(new_n3588_), .A2(new_n3602_), .ZN(new_n3603_));
  NOR2_X1    g03539(.A1(new_n3601_), .A2(new_n3592_), .ZN(new_n3604_));
  NOR3_X1    g03540(.A1(new_n3553_), .A2(new_n3603_), .A3(new_n3604_), .ZN(new_n3605_));
  INV_X1     g03541(.I(new_n3553_), .ZN(new_n3606_));
  NOR2_X1    g03542(.A1(new_n3603_), .A2(new_n3604_), .ZN(new_n3607_));
  NOR2_X1    g03543(.A1(new_n3606_), .A2(new_n3607_), .ZN(new_n3608_));
  NOR2_X1    g03544(.A1(new_n3608_), .A2(new_n3605_), .ZN(new_n3609_));
  NOR2_X1    g03545(.A1(new_n3609_), .A2(new_n3327_), .ZN(new_n3610_));
  INV_X1     g03546(.I(new_n3327_), .ZN(new_n3611_));
  XOR2_X1    g03547(.A1(new_n3553_), .A2(new_n3607_), .Z(new_n3612_));
  NOR2_X1    g03548(.A1(new_n3612_), .A2(new_n3611_), .ZN(new_n3613_));
  OAI22_X1   g03549(.A1(new_n813_), .A2(new_n3268_), .B1(new_n529_), .B2(new_n3318_), .ZN(new_n3614_));
  NAND2_X1   g03550(.A1(new_n2563_), .A2(new_n3323_), .ZN(new_n3615_));
  AOI21_X1   g03551(.A1(new_n3615_), .A2(new_n3614_), .B(new_n3260_), .ZN(new_n3616_));
  NAND2_X1   g03552(.A1(new_n3051_), .A2(new_n3616_), .ZN(new_n3617_));
  XOR2_X1    g03553(.A1(new_n3617_), .A2(\a[26] ), .Z(new_n3618_));
  INV_X1     g03554(.I(new_n3618_), .ZN(new_n3619_));
  NAND2_X1   g03555(.A1(new_n2508_), .A2(new_n2510_), .ZN(new_n3620_));
  XNOR2_X1   g03556(.A1(new_n2559_), .A2(new_n813_), .ZN(new_n3621_));
  NOR2_X1    g03557(.A1(new_n3620_), .A2(new_n3621_), .ZN(new_n3622_));
  AOI22_X1   g03558(.A1(new_n2508_), .A2(new_n2510_), .B1(new_n2561_), .B2(new_n2565_), .ZN(new_n3623_));
  OR2_X2     g03559(.A1(new_n3622_), .A2(new_n3623_), .Z(new_n3624_));
  OAI22_X1   g03560(.A1(new_n2559_), .A2(new_n3318_), .B1(new_n896_), .B2(new_n3268_), .ZN(new_n3625_));
  NAND2_X1   g03561(.A1(new_n814_), .A2(new_n3323_), .ZN(new_n3626_));
  AOI21_X1   g03562(.A1(new_n3625_), .A2(new_n3626_), .B(new_n3260_), .ZN(new_n3627_));
  NAND2_X1   g03563(.A1(new_n3624_), .A2(new_n3627_), .ZN(new_n3628_));
  XOR2_X1    g03564(.A1(new_n3628_), .A2(\a[26] ), .Z(new_n3629_));
  INV_X1     g03565(.I(new_n3629_), .ZN(new_n3630_));
  AOI21_X1   g03566(.A1(new_n3584_), .A2(new_n3586_), .B(new_n3567_), .ZN(new_n3631_));
  XOR2_X1    g03567(.A1(new_n3571_), .A2(new_n3581_), .Z(new_n3632_));
  NOR2_X1    g03568(.A1(new_n3568_), .A2(new_n3632_), .ZN(new_n3633_));
  NOR2_X1    g03569(.A1(new_n3633_), .A2(new_n3631_), .ZN(new_n3634_));
  INV_X1     g03570(.I(new_n3634_), .ZN(new_n3635_));
  OAI22_X1   g03571(.A1(new_n1180_), .A2(new_n3175_), .B1(new_n2492_), .B2(new_n2747_), .ZN(new_n3636_));
  NAND2_X1   g03572(.A1(new_n1122_), .A2(new_n3275_), .ZN(new_n3637_));
  AOI21_X1   g03573(.A1(new_n3637_), .A2(new_n3636_), .B(new_n2737_), .ZN(new_n3638_));
  NAND2_X1   g03574(.A1(new_n3330_), .A2(new_n3638_), .ZN(new_n3639_));
  XOR2_X1    g03575(.A1(new_n3639_), .A2(new_n74_), .Z(new_n3640_));
  INV_X1     g03576(.I(new_n3525_), .ZN(new_n3641_));
  AOI21_X1   g03577(.A1(new_n3641_), .A2(new_n3526_), .B(new_n3407_), .ZN(new_n3642_));
  XOR2_X1    g03578(.A1(new_n3523_), .A2(new_n3528_), .Z(new_n3643_));
  AOI21_X1   g03579(.A1(new_n3407_), .A2(new_n3643_), .B(new_n3642_), .ZN(new_n3644_));
  NAND3_X1   g03580(.A1(new_n2362_), .A2(new_n1408_), .A3(new_n1453_), .ZN(new_n3645_));
  NAND4_X1   g03581(.A1(new_n2358_), .A2(new_n1409_), .A3(new_n2359_), .A4(new_n2361_), .ZN(new_n3646_));
  XOR2_X1    g03582(.A1(new_n1408_), .A2(new_n1333_), .Z(new_n3647_));
  INV_X1     g03583(.I(new_n3647_), .ZN(new_n3648_));
  NAND2_X1   g03584(.A1(new_n3646_), .A2(new_n3648_), .ZN(new_n3649_));
  INV_X1     g03585(.I(new_n3649_), .ZN(new_n3650_));
  NAND3_X1   g03586(.A1(new_n3650_), .A2(new_n1241_), .A3(new_n3645_), .ZN(new_n3651_));
  INV_X1     g03587(.I(new_n3645_), .ZN(new_n3652_));
  OAI21_X1   g03588(.A1(new_n3652_), .A2(new_n3649_), .B(new_n2367_), .ZN(new_n3653_));
  NAND2_X1   g03589(.A1(new_n3651_), .A2(new_n3653_), .ZN(new_n3654_));
  NOR2_X1    g03590(.A1(new_n1333_), .A2(new_n2767_), .ZN(new_n3655_));
  NOR2_X1    g03591(.A1(new_n1409_), .A2(new_n2771_), .ZN(new_n3656_));
  NOR2_X1    g03592(.A1(new_n2367_), .A2(new_n2772_), .ZN(new_n3657_));
  NOR4_X1    g03593(.A1(new_n3656_), .A2(new_n3657_), .A3(new_n2763_), .A4(new_n3655_), .ZN(new_n3658_));
  NAND2_X1   g03594(.A1(new_n3654_), .A2(new_n3658_), .ZN(new_n3659_));
  INV_X1     g03595(.I(new_n3659_), .ZN(new_n3660_));
  NAND2_X1   g03596(.A1(new_n1222_), .A2(new_n479_), .ZN(new_n3661_));
  NOR4_X1    g03597(.A1(new_n3661_), .A2(new_n456_), .A3(new_n682_), .A4(new_n1092_), .ZN(new_n3662_));
  NOR2_X1    g03598(.A1(new_n988_), .A2(new_n2284_), .ZN(new_n3663_));
  NOR4_X1    g03599(.A1(new_n226_), .A2(new_n654_), .A3(new_n1031_), .A4(new_n419_), .ZN(new_n3664_));
  NOR2_X1    g03600(.A1(new_n3664_), .A2(new_n1797_), .ZN(new_n3665_));
  NAND4_X1   g03601(.A1(new_n3662_), .A2(new_n3663_), .A3(new_n1825_), .A4(new_n3665_), .ZN(new_n3666_));
  NOR4_X1    g03602(.A1(new_n366_), .A2(new_n582_), .A3(new_n459_), .A4(new_n724_), .ZN(new_n3667_));
  NAND4_X1   g03603(.A1(new_n439_), .A2(new_n880_), .A3(new_n980_), .A4(new_n1465_), .ZN(new_n3668_));
  NAND4_X1   g03604(.A1(new_n612_), .A2(new_n1091_), .A3(new_n686_), .A4(new_n832_), .ZN(new_n3669_));
  NAND4_X1   g03605(.A1(new_n3669_), .A2(new_n144_), .A3(new_n1025_), .A4(new_n2944_), .ZN(new_n3670_));
  NOR2_X1    g03606(.A1(new_n252_), .A2(new_n236_), .ZN(new_n3671_));
  NAND4_X1   g03607(.A1(new_n1751_), .A2(new_n3671_), .A3(new_n938_), .A4(new_n2192_), .ZN(new_n3672_));
  OR3_X2     g03608(.A1(new_n3670_), .A2(new_n1496_), .A3(new_n3672_), .Z(new_n3673_));
  NOR4_X1    g03609(.A1(new_n3673_), .A2(new_n3666_), .A3(new_n3667_), .A4(new_n3668_), .ZN(new_n3674_));
  NOR4_X1    g03610(.A1(new_n2438_), .A2(new_n332_), .A3(new_n617_), .A4(new_n1461_), .ZN(new_n3675_));
  INV_X1     g03611(.I(new_n714_), .ZN(new_n3676_));
  NAND4_X1   g03612(.A1(new_n3676_), .A2(new_n207_), .A3(new_n1646_), .A4(new_n322_), .ZN(new_n3677_));
  NAND4_X1   g03613(.A1(new_n1628_), .A2(new_n628_), .A3(new_n934_), .A4(new_n1590_), .ZN(new_n3678_));
  NOR3_X1    g03614(.A1(new_n1365_), .A2(new_n844_), .A3(new_n930_), .ZN(new_n3679_));
  INV_X1     g03615(.I(new_n3679_), .ZN(new_n3680_));
  NAND4_X1   g03616(.A1(new_n664_), .A2(new_n3365_), .A3(new_n1767_), .A4(new_n2810_), .ZN(new_n3681_));
  NOR3_X1    g03617(.A1(new_n3680_), .A2(new_n821_), .A3(new_n3681_), .ZN(new_n3682_));
  NAND4_X1   g03618(.A1(new_n3682_), .A2(new_n3675_), .A3(new_n3677_), .A4(new_n3678_), .ZN(new_n3683_));
  NOR3_X1    g03619(.A1(new_n3218_), .A2(new_n1048_), .A3(new_n1589_), .ZN(new_n3684_));
  INV_X1     g03620(.I(new_n2795_), .ZN(new_n3685_));
  NOR3_X1    g03621(.A1(new_n2083_), .A2(new_n3685_), .A3(new_n1200_), .ZN(new_n3686_));
  INV_X1     g03622(.I(new_n887_), .ZN(new_n3687_));
  NOR3_X1    g03623(.A1(new_n746_), .A2(new_n3687_), .A3(new_n912_), .ZN(new_n3688_));
  NOR4_X1    g03624(.A1(new_n106_), .A2(new_n268_), .A3(new_n732_), .A4(new_n506_), .ZN(new_n3689_));
  NOR4_X1    g03625(.A1(new_n751_), .A2(new_n447_), .A3(new_n1167_), .A4(new_n468_), .ZN(new_n3690_));
  NOR4_X1    g03626(.A1(new_n3093_), .A2(new_n3209_), .A3(new_n3689_), .A4(new_n3690_), .ZN(new_n3691_));
  NAND4_X1   g03627(.A1(new_n3691_), .A2(new_n3684_), .A3(new_n3686_), .A4(new_n3688_), .ZN(new_n3692_));
  NOR2_X1    g03628(.A1(new_n3683_), .A2(new_n3692_), .ZN(new_n3693_));
  NAND2_X1   g03629(.A1(new_n3693_), .A2(new_n3674_), .ZN(new_n3694_));
  INV_X1     g03630(.I(new_n3694_), .ZN(new_n3695_));
  NOR2_X1    g03631(.A1(new_n3695_), .A2(new_n3517_), .ZN(new_n3696_));
  INV_X1     g03632(.I(new_n3696_), .ZN(new_n3697_));
  NOR2_X1    g03633(.A1(new_n3518_), .A2(new_n3694_), .ZN(new_n3698_));
  AOI21_X1   g03634(.A1(new_n3660_), .A2(new_n3697_), .B(new_n3698_), .ZN(new_n3699_));
  INV_X1     g03635(.I(new_n3699_), .ZN(new_n3700_));
  INV_X1     g03636(.I(new_n2364_), .ZN(new_n3701_));
  INV_X1     g03637(.I(new_n2366_), .ZN(new_n3702_));
  NOR2_X1    g03638(.A1(new_n3701_), .A2(new_n3702_), .ZN(new_n3703_));
  XOR2_X1    g03639(.A1(new_n1241_), .A2(new_n2408_), .Z(new_n3704_));
  NOR3_X1    g03640(.A1(new_n3701_), .A2(new_n3702_), .A3(new_n3704_), .ZN(new_n3705_));
  INV_X1     g03641(.I(new_n3705_), .ZN(new_n3706_));
  NOR2_X1    g03642(.A1(new_n2409_), .A2(new_n2413_), .ZN(new_n3707_));
  OAI21_X1   g03643(.A1(new_n3703_), .A2(new_n3707_), .B(new_n3706_), .ZN(new_n3708_));
  NOR2_X1    g03644(.A1(new_n1333_), .A2(new_n2771_), .ZN(new_n3709_));
  NOR2_X1    g03645(.A1(new_n2408_), .A2(new_n2772_), .ZN(new_n3710_));
  NOR2_X1    g03646(.A1(new_n2367_), .A2(new_n2767_), .ZN(new_n3711_));
  NOR4_X1    g03647(.A1(new_n3711_), .A2(new_n3709_), .A3(new_n3710_), .A4(new_n2763_), .ZN(new_n3712_));
  NOR2_X1    g03648(.A1(new_n3519_), .A2(new_n3522_), .ZN(new_n3713_));
  NOR2_X1    g03649(.A1(new_n3713_), .A2(new_n3477_), .ZN(new_n3714_));
  XOR2_X1    g03650(.A1(new_n3517_), .A2(\a[14] ), .Z(new_n3715_));
  INV_X1     g03651(.I(new_n3715_), .ZN(new_n3716_));
  AOI21_X1   g03652(.A1(new_n3477_), .A2(new_n3716_), .B(new_n3714_), .ZN(new_n3717_));
  INV_X1     g03653(.I(new_n3717_), .ZN(new_n3718_));
  AOI21_X1   g03654(.A1(new_n3708_), .A2(new_n3712_), .B(new_n3718_), .ZN(new_n3719_));
  INV_X1     g03655(.I(new_n3719_), .ZN(new_n3720_));
  NAND2_X1   g03656(.A1(new_n3720_), .A2(new_n3700_), .ZN(new_n3721_));
  NAND2_X1   g03657(.A1(new_n3708_), .A2(new_n3712_), .ZN(new_n3722_));
  NOR2_X1    g03658(.A1(new_n3722_), .A2(new_n3717_), .ZN(new_n3723_));
  INV_X1     g03659(.I(new_n3723_), .ZN(new_n3724_));
  NAND2_X1   g03660(.A1(new_n3721_), .A2(new_n3724_), .ZN(new_n3725_));
  INV_X1     g03661(.I(new_n3725_), .ZN(new_n3726_));
  NAND2_X1   g03662(.A1(new_n3726_), .A2(new_n3644_), .ZN(new_n3727_));
  NOR2_X1    g03663(.A1(new_n3726_), .A2(new_n3644_), .ZN(new_n3728_));
  AOI21_X1   g03664(.A1(new_n3640_), .A2(new_n3727_), .B(new_n3728_), .ZN(new_n3729_));
  INV_X1     g03665(.I(new_n3729_), .ZN(new_n3730_));
  NOR2_X1    g03666(.A1(new_n3635_), .A2(new_n3730_), .ZN(new_n3731_));
  INV_X1     g03667(.I(new_n3731_), .ZN(new_n3732_));
  NOR2_X1    g03668(.A1(new_n3634_), .A2(new_n3729_), .ZN(new_n3733_));
  AOI21_X1   g03669(.A1(new_n3732_), .A2(new_n3630_), .B(new_n3733_), .ZN(new_n3734_));
  INV_X1     g03670(.I(new_n3734_), .ZN(new_n3735_));
  OAI21_X1   g03671(.A1(new_n3602_), .A2(new_n3604_), .B(new_n3587_), .ZN(new_n3736_));
  XNOR2_X1   g03672(.A1(new_n3601_), .A2(new_n3592_), .ZN(new_n3737_));
  OAI21_X1   g03673(.A1(new_n3587_), .A2(new_n3737_), .B(new_n3736_), .ZN(new_n3738_));
  NOR2_X1    g03674(.A1(new_n3735_), .A2(new_n3738_), .ZN(new_n3739_));
  INV_X1     g03675(.I(new_n3739_), .ZN(new_n3740_));
  NAND2_X1   g03676(.A1(new_n3735_), .A2(new_n3738_), .ZN(new_n3741_));
  INV_X1     g03677(.I(new_n3741_), .ZN(new_n3742_));
  AOI21_X1   g03678(.A1(new_n3619_), .A2(new_n3740_), .B(new_n3742_), .ZN(new_n3743_));
  INV_X1     g03679(.I(new_n3743_), .ZN(new_n3744_));
  NOR3_X1    g03680(.A1(new_n3744_), .A2(new_n3610_), .A3(new_n3613_), .ZN(new_n3745_));
  NOR2_X1    g03681(.A1(new_n3610_), .A2(new_n3613_), .ZN(new_n3746_));
  NOR2_X1    g03682(.A1(new_n3746_), .A2(new_n3743_), .ZN(new_n3747_));
  NOR2_X1    g03683(.A1(new_n3747_), .A2(new_n3745_), .ZN(new_n3748_));
  NOR2_X1    g03684(.A1(new_n3748_), .A2(new_n3316_), .ZN(new_n3749_));
  INV_X1     g03685(.I(new_n3316_), .ZN(new_n3750_));
  XOR2_X1    g03686(.A1(new_n3746_), .A2(new_n3744_), .Z(new_n3751_));
  NOR2_X1    g03687(.A1(new_n3751_), .A2(new_n3750_), .ZN(new_n3752_));
  NOR2_X1    g03688(.A1(new_n3752_), .A2(new_n3749_), .ZN(new_n3753_));
  XOR2_X1    g03689(.A1(new_n3168_), .A2(new_n3142_), .Z(new_n3754_));
  INV_X1     g03690(.I(new_n3754_), .ZN(new_n3755_));
  XOR2_X1    g03691(.A1(new_n2716_), .A2(new_n3247_), .Z(new_n3756_));
  NAND3_X1   g03692(.A1(new_n3145_), .A2(new_n3143_), .A3(new_n3756_), .ZN(new_n3757_));
  AND2_X2    g03693(.A1(new_n3757_), .A2(new_n3755_), .Z(new_n3758_));
  INV_X1     g03694(.I(\a[18] ), .ZN(new_n3759_));
  NOR2_X1    g03695(.A1(new_n3759_), .A2(\a[17] ), .ZN(new_n3760_));
  NOR2_X1    g03696(.A1(new_n3372_), .A2(\a[18] ), .ZN(new_n3761_));
  NOR2_X1    g03697(.A1(new_n3760_), .A2(new_n3761_), .ZN(new_n3762_));
  INV_X1     g03698(.I(new_n3762_), .ZN(new_n3763_));
  INV_X1     g03699(.I(\a[19] ), .ZN(new_n3764_));
  NOR2_X1    g03700(.A1(new_n3764_), .A2(\a[17] ), .ZN(new_n3765_));
  NOR2_X1    g03701(.A1(new_n3372_), .A2(\a[19] ), .ZN(new_n3766_));
  OR2_X2     g03702(.A1(new_n3765_), .A2(new_n3766_), .Z(new_n3767_));
  XNOR2_X1   g03703(.A1(\a[17] ), .A2(\a[20] ), .ZN(new_n3768_));
  OAI21_X1   g03704(.A1(new_n3763_), .A2(new_n3767_), .B(new_n3768_), .ZN(new_n3769_));
  INV_X1     g03705(.I(new_n3769_), .ZN(new_n3770_));
  NAND2_X1   g03706(.A1(new_n3168_), .A2(new_n3770_), .ZN(new_n3771_));
  XNOR2_X1   g03707(.A1(\a[19] ), .A2(\a[20] ), .ZN(new_n3772_));
  NOR2_X1    g03708(.A1(new_n3762_), .A2(new_n3772_), .ZN(new_n3773_));
  NOR3_X1    g03709(.A1(new_n3764_), .A2(\a[17] ), .A3(\a[18] ), .ZN(new_n3774_));
  AOI21_X1   g03710(.A1(\a[18] ), .A2(new_n3766_), .B(new_n3774_), .ZN(new_n3775_));
  INV_X1     g03711(.I(new_n3775_), .ZN(new_n3776_));
  NAND2_X1   g03712(.A1(new_n3247_), .A2(new_n3776_), .ZN(new_n3777_));
  NAND4_X1   g03713(.A1(new_n3758_), .A2(new_n3771_), .A3(new_n3773_), .A4(new_n3777_), .ZN(new_n3778_));
  XOR2_X1    g03714(.A1(new_n3778_), .A2(\a[20] ), .Z(new_n3779_));
  INV_X1     g03715(.I(new_n3312_), .ZN(new_n3780_));
  OAI22_X1   g03716(.A1(new_n694_), .A2(new_n3310_), .B1(new_n2665_), .B2(new_n3780_), .ZN(new_n3781_));
  INV_X1     g03717(.I(new_n3306_), .ZN(new_n3782_));
  NAND2_X1   g03718(.A1(new_n2615_), .A2(new_n3782_), .ZN(new_n3783_));
  AOI21_X1   g03719(.A1(new_n3781_), .A2(new_n3783_), .B(new_n3302_), .ZN(new_n3784_));
  NAND2_X1   g03720(.A1(new_n3188_), .A2(new_n3784_), .ZN(new_n3785_));
  XOR2_X1    g03721(.A1(new_n3785_), .A2(\a[23] ), .Z(new_n3786_));
  INV_X1     g03722(.I(new_n3786_), .ZN(new_n3787_));
  XOR2_X1    g03723(.A1(new_n3734_), .A2(new_n3738_), .Z(new_n3788_));
  NOR2_X1    g03724(.A1(new_n3788_), .A2(new_n3618_), .ZN(new_n3789_));
  AOI21_X1   g03725(.A1(new_n3740_), .A2(new_n3741_), .B(new_n3619_), .ZN(new_n3790_));
  NOR2_X1    g03726(.A1(new_n3790_), .A2(new_n3789_), .ZN(new_n3791_));
  OAI22_X1   g03727(.A1(new_n2614_), .A2(new_n3780_), .B1(new_n529_), .B2(new_n3310_), .ZN(new_n3792_));
  NAND2_X1   g03728(.A1(new_n2718_), .A2(new_n3782_), .ZN(new_n3793_));
  AOI21_X1   g03729(.A1(new_n3793_), .A2(new_n3792_), .B(new_n3302_), .ZN(new_n3794_));
  NAND2_X1   g03730(.A1(new_n3074_), .A2(new_n3794_), .ZN(new_n3795_));
  XOR2_X1    g03731(.A1(new_n3795_), .A2(\a[23] ), .Z(new_n3796_));
  INV_X1     g03732(.I(new_n3796_), .ZN(new_n3797_));
  OAI21_X1   g03733(.A1(new_n3731_), .A2(new_n3733_), .B(new_n3630_), .ZN(new_n3798_));
  XOR2_X1    g03734(.A1(new_n3634_), .A2(new_n3730_), .Z(new_n3799_));
  OAI21_X1   g03735(.A1(new_n3630_), .A2(new_n3799_), .B(new_n3798_), .ZN(new_n3800_));
  OAI22_X1   g03736(.A1(new_n813_), .A2(new_n3318_), .B1(new_n1008_), .B2(new_n3268_), .ZN(new_n3801_));
  NAND2_X1   g03737(.A1(new_n897_), .A2(new_n3323_), .ZN(new_n3802_));
  AOI21_X1   g03738(.A1(new_n3801_), .A2(new_n3802_), .B(new_n3260_), .ZN(new_n3803_));
  NAND2_X1   g03739(.A1(new_n2917_), .A2(new_n3803_), .ZN(new_n3804_));
  XOR2_X1    g03740(.A1(new_n3804_), .A2(\a[26] ), .Z(new_n3805_));
  OAI22_X1   g03741(.A1(new_n1121_), .A2(new_n3175_), .B1(new_n2451_), .B2(new_n2747_), .ZN(new_n3806_));
  NAND2_X1   g03742(.A1(new_n2496_), .A2(new_n3275_), .ZN(new_n3807_));
  AOI21_X1   g03743(.A1(new_n3806_), .A2(new_n3807_), .B(new_n2737_), .ZN(new_n3808_));
  NAND2_X1   g03744(.A1(new_n3393_), .A2(new_n3808_), .ZN(new_n3809_));
  XOR2_X1    g03745(.A1(new_n3809_), .A2(\a[29] ), .Z(new_n3810_));
  INV_X1     g03746(.I(new_n3810_), .ZN(new_n3811_));
  OAI22_X1   g03747(.A1(new_n2367_), .A2(new_n2747_), .B1(new_n2451_), .B2(new_n3175_), .ZN(new_n3812_));
  NAND2_X1   g03748(.A1(new_n2412_), .A2(new_n3275_), .ZN(new_n3813_));
  AOI21_X1   g03749(.A1(new_n3812_), .A2(new_n3813_), .B(new_n2737_), .ZN(new_n3814_));
  NAND2_X1   g03750(.A1(new_n3403_), .A2(new_n3814_), .ZN(new_n3815_));
  XOR2_X1    g03751(.A1(new_n3815_), .A2(\a[29] ), .Z(new_n3816_));
  INV_X1     g03752(.I(new_n3816_), .ZN(new_n3817_));
  NOR2_X1    g03753(.A1(new_n1409_), .A2(new_n1453_), .ZN(new_n3818_));
  INV_X1     g03754(.I(new_n3818_), .ZN(new_n3819_));
  NAND2_X1   g03755(.A1(new_n2362_), .A2(new_n3819_), .ZN(new_n3820_));
  NOR2_X1    g03756(.A1(new_n2359_), .A2(new_n1408_), .ZN(new_n3821_));
  INV_X1     g03757(.I(new_n3821_), .ZN(new_n3822_));
  AOI21_X1   g03758(.A1(new_n3820_), .A2(new_n3822_), .B(new_n3647_), .ZN(new_n3823_));
  INV_X1     g03759(.I(new_n3823_), .ZN(new_n3824_));
  XNOR2_X1   g03760(.A1(new_n1408_), .A2(new_n1333_), .ZN(new_n3825_));
  INV_X1     g03761(.I(new_n3825_), .ZN(new_n3826_));
  NAND3_X1   g03762(.A1(new_n3820_), .A2(new_n3822_), .A3(new_n3826_), .ZN(new_n3827_));
  NAND2_X1   g03763(.A1(new_n3824_), .A2(new_n3827_), .ZN(new_n3828_));
  NOR2_X1    g03764(.A1(new_n1333_), .A2(new_n2772_), .ZN(new_n3829_));
  NOR2_X1    g03765(.A1(new_n1453_), .A2(new_n2771_), .ZN(new_n3830_));
  NOR2_X1    g03766(.A1(new_n1409_), .A2(new_n2767_), .ZN(new_n3831_));
  NOR4_X1    g03767(.A1(new_n3831_), .A2(new_n2763_), .A3(new_n3829_), .A4(new_n3830_), .ZN(new_n3832_));
  NAND2_X1   g03768(.A1(new_n3828_), .A2(new_n3832_), .ZN(new_n3833_));
  INV_X1     g03769(.I(new_n2320_), .ZN(new_n3834_));
  NOR3_X1    g03770(.A1(new_n3220_), .A2(new_n549_), .A3(new_n1858_), .ZN(new_n3835_));
  INV_X1     g03771(.I(new_n3835_), .ZN(new_n3836_));
  NOR3_X1    g03772(.A1(new_n666_), .A2(new_n130_), .A3(new_n791_), .ZN(new_n3837_));
  NOR2_X1    g03773(.A1(new_n3412_), .A2(new_n1055_), .ZN(new_n3838_));
  NAND4_X1   g03774(.A1(new_n442_), .A2(new_n2375_), .A3(new_n434_), .A4(new_n1058_), .ZN(new_n3839_));
  NOR3_X1    g03775(.A1(new_n217_), .A2(new_n261_), .A3(new_n430_), .ZN(new_n3840_));
  NAND4_X1   g03776(.A1(new_n3838_), .A2(new_n3839_), .A3(new_n3837_), .A4(new_n3840_), .ZN(new_n3841_));
  NOR4_X1    g03777(.A1(new_n3834_), .A2(new_n3508_), .A3(new_n3836_), .A4(new_n3841_), .ZN(new_n3842_));
  INV_X1     g03778(.I(new_n3842_), .ZN(new_n3843_));
  NOR4_X1    g03779(.A1(new_n164_), .A2(new_n170_), .A3(new_n294_), .A4(new_n419_), .ZN(new_n3844_));
  INV_X1     g03780(.I(new_n3844_), .ZN(new_n3845_));
  NOR3_X1    g03781(.A1(new_n225_), .A2(new_n638_), .A3(new_n744_), .ZN(new_n3846_));
  NAND4_X1   g03782(.A1(new_n1221_), .A2(new_n436_), .A3(new_n999_), .A4(new_n441_), .ZN(new_n3847_));
  NAND4_X1   g03783(.A1(new_n1281_), .A2(new_n3845_), .A3(new_n3846_), .A4(new_n3847_), .ZN(new_n3848_));
  NOR4_X1    g03784(.A1(new_n740_), .A2(new_n515_), .A3(new_n460_), .A4(new_n561_), .ZN(new_n3849_));
  NOR4_X1    g03785(.A1(new_n3849_), .A2(new_n937_), .A3(new_n418_), .A4(new_n1995_), .ZN(new_n3850_));
  INV_X1     g03786(.I(new_n3850_), .ZN(new_n3851_));
  NAND2_X1   g03787(.A1(new_n2862_), .A2(new_n1679_), .ZN(new_n3852_));
  NOR4_X1    g03788(.A1(new_n3851_), .A2(new_n3848_), .A3(new_n2248_), .A4(new_n3852_), .ZN(new_n3853_));
  INV_X1     g03789(.I(new_n3853_), .ZN(new_n3854_));
  INV_X1     g03790(.I(new_n2620_), .ZN(new_n3855_));
  NAND2_X1   g03791(.A1(new_n677_), .A2(new_n1025_), .ZN(new_n3856_));
  NOR3_X1    g03792(.A1(new_n3460_), .A2(new_n2439_), .A3(new_n424_), .ZN(new_n3857_));
  NOR4_X1    g03793(.A1(new_n1714_), .A2(new_n190_), .A3(new_n1175_), .A4(new_n345_), .ZN(new_n3858_));
  NAND4_X1   g03794(.A1(new_n3857_), .A2(new_n452_), .A3(new_n3858_), .A4(new_n653_), .ZN(new_n3859_));
  NOR4_X1    g03795(.A1(new_n3859_), .A2(new_n1328_), .A3(new_n3855_), .A4(new_n3856_), .ZN(new_n3860_));
  INV_X1     g03796(.I(new_n3860_), .ZN(new_n3861_));
  NOR4_X1    g03797(.A1(new_n3843_), .A2(new_n728_), .A3(new_n3861_), .A4(new_n3854_), .ZN(new_n3862_));
  NAND4_X1   g03798(.A1(new_n138_), .A2(new_n1358_), .A3(new_n2944_), .A4(new_n1840_), .ZN(new_n3863_));
  NOR4_X1    g03799(.A1(new_n251_), .A2(new_n584_), .A3(new_n791_), .A4(new_n280_), .ZN(new_n3864_));
  NAND2_X1   g03800(.A1(new_n540_), .A2(new_n502_), .ZN(new_n3865_));
  NOR4_X1    g03801(.A1(new_n3863_), .A2(new_n268_), .A3(new_n3864_), .A4(new_n3865_), .ZN(new_n3866_));
  NOR3_X1    g03802(.A1(new_n906_), .A2(new_n1531_), .A3(new_n397_), .ZN(new_n3867_));
  NOR2_X1    g03803(.A1(new_n634_), .A2(new_n625_), .ZN(new_n3868_));
  NOR4_X1    g03804(.A1(new_n1984_), .A2(new_n591_), .A3(new_n76_), .A4(new_n485_), .ZN(new_n3869_));
  NOR4_X1    g03805(.A1(new_n117_), .A2(new_n198_), .A3(new_n515_), .A4(new_n535_), .ZN(new_n3870_));
  NOR2_X1    g03806(.A1(new_n3869_), .A2(new_n3870_), .ZN(new_n3871_));
  AND4_X2    g03807(.A1(new_n1599_), .A2(new_n3871_), .A3(new_n3867_), .A4(new_n3868_), .Z(new_n3872_));
  NOR4_X1    g03808(.A1(new_n1276_), .A2(new_n825_), .A3(new_n3353_), .A4(new_n2098_), .ZN(new_n3873_));
  NAND4_X1   g03809(.A1(new_n3872_), .A2(new_n1135_), .A3(new_n3866_), .A4(new_n3873_), .ZN(new_n3874_));
  NOR4_X1    g03810(.A1(new_n602_), .A2(new_n644_), .A3(new_n714_), .A4(new_n307_), .ZN(new_n3875_));
  NOR4_X1    g03811(.A1(new_n945_), .A2(new_n752_), .A3(new_n460_), .A4(new_n744_), .ZN(new_n3876_));
  INV_X1     g03812(.I(new_n3876_), .ZN(new_n3877_));
  NAND4_X1   g03813(.A1(new_n385_), .A2(new_n3502_), .A3(new_n690_), .A4(new_n361_), .ZN(new_n3878_));
  NAND4_X1   g03814(.A1(new_n2370_), .A2(new_n3875_), .A3(new_n3877_), .A4(new_n3878_), .ZN(new_n3879_));
  NAND4_X1   g03815(.A1(new_n766_), .A2(new_n1679_), .A3(new_n1712_), .A4(new_n1883_), .ZN(new_n3880_));
  NOR2_X1    g03816(.A1(new_n534_), .A2(new_n172_), .ZN(new_n3881_));
  NAND4_X1   g03817(.A1(new_n3881_), .A2(new_n1495_), .A3(new_n389_), .A4(new_n1526_), .ZN(new_n3882_));
  NOR4_X1    g03818(.A1(new_n3028_), .A2(new_n3882_), .A3(new_n3879_), .A4(new_n3880_), .ZN(new_n3883_));
  INV_X1     g03819(.I(new_n3883_), .ZN(new_n3884_));
  NOR4_X1    g03820(.A1(new_n3884_), .A2(new_n2818_), .A3(new_n3861_), .A4(new_n3874_), .ZN(new_n3885_));
  NOR2_X1    g03821(.A1(new_n3885_), .A2(\a[11] ), .ZN(new_n3886_));
  INV_X1     g03822(.I(new_n3886_), .ZN(new_n3887_));
  NAND2_X1   g03823(.A1(new_n3885_), .A2(\a[11] ), .ZN(new_n3888_));
  INV_X1     g03824(.I(new_n3888_), .ZN(new_n3889_));
  AOI21_X1   g03825(.A1(new_n3862_), .A2(new_n3887_), .B(new_n3889_), .ZN(new_n3890_));
  NOR2_X1    g03826(.A1(new_n3890_), .A2(new_n3518_), .ZN(new_n3891_));
  INV_X1     g03827(.I(new_n3891_), .ZN(new_n3892_));
  NAND2_X1   g03828(.A1(new_n3890_), .A2(new_n3518_), .ZN(new_n3893_));
  AOI21_X1   g03829(.A1(new_n3892_), .A2(new_n3893_), .B(new_n3833_), .ZN(new_n3894_));
  INV_X1     g03830(.I(new_n3833_), .ZN(new_n3895_));
  XOR2_X1    g03831(.A1(new_n3890_), .A2(new_n3517_), .Z(new_n3896_));
  NOR2_X1    g03832(.A1(new_n3895_), .A2(new_n3896_), .ZN(new_n3897_));
  NOR2_X1    g03833(.A1(new_n3897_), .A2(new_n3894_), .ZN(new_n3898_));
  INV_X1     g03834(.I(new_n3898_), .ZN(new_n3899_));
  XOR2_X1    g03835(.A1(new_n1453_), .A2(new_n1408_), .Z(new_n3900_));
  AOI21_X1   g03836(.A1(new_n2358_), .A2(new_n2361_), .B(new_n3900_), .ZN(new_n3901_));
  INV_X1     g03837(.I(new_n3901_), .ZN(new_n3902_));
  NOR2_X1    g03838(.A1(new_n3821_), .A2(new_n3818_), .ZN(new_n3903_));
  OAI21_X1   g03839(.A1(new_n2362_), .A2(new_n3903_), .B(new_n3902_), .ZN(new_n3904_));
  AOI21_X1   g03840(.A1(new_n2354_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n3905_));
  OAI21_X1   g03841(.A1(new_n1409_), .A2(new_n2772_), .B(new_n3905_), .ZN(new_n3906_));
  AOI21_X1   g03842(.A1(new_n2359_), .A2(new_n3189_), .B(new_n3906_), .ZN(new_n3907_));
  AND2_X2    g03843(.A1(new_n3904_), .A2(new_n3907_), .Z(new_n3908_));
  NAND2_X1   g03844(.A1(new_n2314_), .A2(new_n2316_), .ZN(new_n3909_));
  XOR2_X1    g03845(.A1(new_n2310_), .A2(new_n2351_), .Z(new_n3910_));
  AOI21_X1   g03846(.A1(new_n2314_), .A2(new_n2316_), .B(new_n3910_), .ZN(new_n3911_));
  INV_X1     g03847(.I(new_n3911_), .ZN(new_n3912_));
  NOR2_X1    g03848(.A1(new_n2352_), .A2(new_n2355_), .ZN(new_n3913_));
  OAI21_X1   g03849(.A1(new_n3909_), .A2(new_n3913_), .B(new_n3912_), .ZN(new_n3914_));
  NOR2_X1    g03850(.A1(new_n2311_), .A2(new_n2767_), .ZN(new_n3915_));
  NOR2_X1    g03851(.A1(new_n2351_), .A2(new_n2772_), .ZN(new_n3916_));
  NOR2_X1    g03852(.A1(new_n2251_), .A2(new_n2771_), .ZN(new_n3917_));
  NOR4_X1    g03853(.A1(new_n3915_), .A2(new_n2763_), .A3(new_n3916_), .A4(new_n3917_), .ZN(new_n3918_));
  NAND2_X1   g03854(.A1(new_n3914_), .A2(new_n3918_), .ZN(new_n3919_));
  INV_X1     g03855(.I(new_n3919_), .ZN(new_n3920_));
  NAND4_X1   g03856(.A1(new_n1217_), .A2(new_n627_), .A3(new_n184_), .A4(new_n414_), .ZN(new_n3921_));
  NOR4_X1    g03857(.A1(new_n137_), .A2(new_n463_), .A3(new_n486_), .A4(new_n388_), .ZN(new_n3922_));
  INV_X1     g03858(.I(new_n3922_), .ZN(new_n3923_));
  NAND2_X1   g03859(.A1(new_n3501_), .A2(new_n3923_), .ZN(new_n3924_));
  NOR4_X1    g03860(.A1(new_n365_), .A2(new_n490_), .A3(new_n611_), .A4(new_n517_), .ZN(new_n3925_));
  NAND3_X1   g03861(.A1(new_n1540_), .A2(new_n1144_), .A3(new_n3925_), .ZN(new_n3926_));
  NOR4_X1    g03862(.A1(new_n251_), .A2(new_n106_), .A3(new_n783_), .A4(new_n242_), .ZN(new_n3927_));
  NOR4_X1    g03863(.A1(new_n866_), .A2(new_n910_), .A3(new_n428_), .A4(new_n594_), .ZN(new_n3928_));
  NOR3_X1    g03864(.A1(new_n2880_), .A2(new_n3928_), .A3(new_n3927_), .ZN(new_n3929_));
  NOR4_X1    g03865(.A1(new_n644_), .A2(new_n310_), .A3(new_n347_), .A4(new_n574_), .ZN(new_n3930_));
  NOR4_X1    g03866(.A1(new_n3930_), .A2(new_n2020_), .A3(new_n398_), .A4(new_n681_), .ZN(new_n3931_));
  NAND2_X1   g03867(.A1(new_n3929_), .A2(new_n3931_), .ZN(new_n3932_));
  NOR4_X1    g03868(.A1(new_n3932_), .A2(new_n3921_), .A3(new_n3924_), .A4(new_n3926_), .ZN(new_n3933_));
  NAND4_X1   g03869(.A1(new_n1222_), .A2(new_n1335_), .A3(new_n1446_), .A4(new_n405_), .ZN(new_n3934_));
  NOR3_X1    g03870(.A1(new_n1211_), .A2(new_n715_), .A3(new_n2338_), .ZN(new_n3935_));
  NAND4_X1   g03871(.A1(new_n982_), .A2(new_n628_), .A3(new_n231_), .A4(new_n709_), .ZN(new_n3936_));
  AND3_X2    g03872(.A1(new_n3935_), .A2(new_n3934_), .A3(new_n3936_), .Z(new_n3937_));
  INV_X1     g03873(.I(new_n2862_), .ZN(new_n3938_));
  NOR3_X1    g03874(.A1(new_n2457_), .A2(new_n1139_), .A3(new_n3938_), .ZN(new_n3939_));
  NOR4_X1    g03875(.A1(new_n954_), .A2(new_n825_), .A3(new_n1994_), .A4(new_n2052_), .ZN(new_n3940_));
  NAND4_X1   g03876(.A1(new_n3937_), .A2(new_n3467_), .A3(new_n3939_), .A4(new_n3940_), .ZN(new_n3941_));
  NAND4_X1   g03877(.A1(new_n309_), .A2(new_n686_), .A3(new_n999_), .A4(new_n409_), .ZN(new_n3942_));
  NOR2_X1    g03878(.A1(new_n465_), .A2(new_n333_), .ZN(new_n3943_));
  INV_X1     g03879(.I(new_n3943_), .ZN(new_n3944_));
  NOR4_X1    g03880(.A1(new_n3944_), .A2(new_n3942_), .A3(new_n1167_), .A4(new_n902_), .ZN(new_n3945_));
  NOR4_X1    g03881(.A1(new_n602_), .A2(new_n666_), .A3(new_n289_), .A4(new_n689_), .ZN(new_n3946_));
  NOR2_X1    g03882(.A1(new_n166_), .A2(new_n3946_), .ZN(new_n3947_));
  NOR3_X1    g03883(.A1(new_n714_), .A2(new_n485_), .A3(new_n352_), .ZN(new_n3948_));
  NAND4_X1   g03884(.A1(new_n1562_), .A2(new_n358_), .A3(new_n840_), .A4(new_n3948_), .ZN(new_n3949_));
  INV_X1     g03885(.I(new_n3949_), .ZN(new_n3950_));
  NAND4_X1   g03886(.A1(new_n3950_), .A2(new_n2231_), .A3(new_n3945_), .A4(new_n3947_), .ZN(new_n3951_));
  NOR4_X1    g03887(.A1(new_n945_), .A2(new_n86_), .A3(new_n548_), .A4(new_n460_), .ZN(new_n3952_));
  NOR4_X1    g03888(.A1(new_n3952_), .A2(new_n955_), .A3(new_n2582_), .A4(new_n841_), .ZN(new_n3953_));
  NAND4_X1   g03889(.A1(new_n3953_), .A2(new_n708_), .A3(new_n1699_), .A4(new_n2145_), .ZN(new_n3954_));
  NOR3_X1    g03890(.A1(new_n326_), .A2(new_n437_), .A3(new_n721_), .ZN(new_n3955_));
  NOR2_X1    g03891(.A1(new_n515_), .A2(new_n719_), .ZN(new_n3956_));
  NAND4_X1   g03892(.A1(new_n3955_), .A2(new_n1766_), .A3(new_n2290_), .A4(new_n3956_), .ZN(new_n3957_));
  NOR4_X1    g03893(.A1(new_n3941_), .A2(new_n3951_), .A3(new_n3954_), .A4(new_n3957_), .ZN(new_n3958_));
  NAND2_X1   g03894(.A1(new_n3958_), .A2(new_n3933_), .ZN(new_n3959_));
  NOR4_X1    g03895(.A1(new_n607_), .A2(new_n241_), .A3(new_n772_), .A4(new_n652_), .ZN(new_n3960_));
  NOR3_X1    g03896(.A1(new_n3960_), .A2(new_n161_), .A3(new_n618_), .ZN(new_n3961_));
  NOR3_X1    g03897(.A1(new_n1211_), .A2(new_n1337_), .A3(new_n625_), .ZN(new_n3962_));
  INV_X1     g03898(.I(new_n3962_), .ZN(new_n3963_));
  NAND2_X1   g03899(.A1(new_n2339_), .A2(new_n1814_), .ZN(new_n3964_));
  NOR4_X1    g03900(.A1(new_n3963_), .A2(new_n3964_), .A3(new_n2982_), .A4(new_n1620_), .ZN(new_n3965_));
  NAND2_X1   g03901(.A1(new_n1565_), .A2(new_n723_), .ZN(new_n3966_));
  NOR4_X1    g03902(.A1(new_n415_), .A2(new_n387_), .A3(new_n403_), .A4(new_n418_), .ZN(new_n3967_));
  NOR4_X1    g03903(.A1(new_n102_), .A2(new_n236_), .A3(new_n930_), .A4(new_n506_), .ZN(new_n3968_));
  NOR4_X1    g03904(.A1(new_n3966_), .A2(new_n2598_), .A3(new_n3967_), .A4(new_n3968_), .ZN(new_n3969_));
  NOR3_X1    g03905(.A1(new_n1157_), .A2(new_n261_), .A3(new_n343_), .ZN(new_n3970_));
  NAND4_X1   g03906(.A1(new_n3970_), .A2(new_n934_), .A3(new_n564_), .A4(new_n1144_), .ZN(new_n3971_));
  NOR4_X1    g03907(.A1(new_n219_), .A2(new_n260_), .A3(new_n381_), .A4(new_n638_), .ZN(new_n3972_));
  NOR3_X1    g03908(.A1(new_n3971_), .A2(new_n2488_), .A3(new_n3972_), .ZN(new_n3973_));
  NAND4_X1   g03909(.A1(new_n3973_), .A2(new_n3965_), .A3(new_n3961_), .A4(new_n3969_), .ZN(new_n3974_));
  INV_X1     g03910(.I(new_n3974_), .ZN(new_n3975_));
  NOR4_X1    g03911(.A1(new_n326_), .A2(new_n732_), .A3(new_n640_), .A4(new_n152_), .ZN(new_n3976_));
  NOR3_X1    g03912(.A1(new_n449_), .A2(new_n719_), .A3(new_n535_), .ZN(new_n3977_));
  INV_X1     g03913(.I(new_n3977_), .ZN(new_n3978_));
  NOR4_X1    g03914(.A1(new_n3978_), .A2(new_n3976_), .A3(new_n125_), .A4(new_n298_), .ZN(new_n3979_));
  INV_X1     g03915(.I(new_n3979_), .ZN(new_n3980_));
  NAND2_X1   g03916(.A1(new_n1891_), .A2(new_n672_), .ZN(new_n3981_));
  NOR4_X1    g03917(.A1(new_n939_), .A2(new_n3981_), .A3(new_n170_), .A4(new_n2994_), .ZN(new_n3982_));
  NOR3_X1    g03918(.A1(new_n267_), .A2(new_n648_), .A3(new_n764_), .ZN(new_n3983_));
  NAND3_X1   g03919(.A1(new_n3982_), .A2(new_n2547_), .A3(new_n3983_), .ZN(new_n3984_));
  NAND4_X1   g03920(.A1(new_n1414_), .A2(new_n253_), .A3(new_n1958_), .A4(new_n1044_), .ZN(new_n3985_));
  NOR4_X1    g03921(.A1(new_n3980_), .A2(new_n3984_), .A3(new_n3456_), .A4(new_n3985_), .ZN(new_n3986_));
  NAND4_X1   g03922(.A1(new_n690_), .A2(new_n834_), .A3(new_n1063_), .A4(new_n1638_), .ZN(new_n3987_));
  NOR4_X1    g03923(.A1(new_n1160_), .A2(new_n744_), .A3(new_n1922_), .A4(new_n1531_), .ZN(new_n3988_));
  NOR4_X1    g03924(.A1(new_n950_), .A2(new_n192_), .A3(new_n203_), .A4(new_n703_), .ZN(new_n3989_));
  INV_X1     g03925(.I(new_n657_), .ZN(new_n3990_));
  INV_X1     g03926(.I(new_n827_), .ZN(new_n3991_));
  NOR4_X1    g03927(.A1(new_n3990_), .A2(new_n3991_), .A3(new_n1243_), .A4(new_n1985_), .ZN(new_n3992_));
  NAND4_X1   g03928(.A1(new_n3989_), .A2(new_n3987_), .A3(new_n3988_), .A4(new_n3992_), .ZN(new_n3993_));
  NAND4_X1   g03929(.A1(new_n612_), .A2(new_n188_), .A3(new_n1590_), .A4(new_n1395_), .ZN(new_n3994_));
  NAND3_X1   g03930(.A1(new_n3447_), .A2(new_n207_), .A3(new_n395_), .ZN(new_n3995_));
  NAND3_X1   g03931(.A1(new_n3995_), .A2(new_n3994_), .A3(new_n336_), .ZN(new_n3996_));
  NOR3_X1    g03932(.A1(new_n190_), .A2(new_n227_), .A3(new_n741_), .ZN(new_n3997_));
  INV_X1     g03933(.I(new_n3997_), .ZN(new_n3998_));
  NAND2_X1   g03934(.A1(new_n1263_), .A2(new_n1126_), .ZN(new_n3999_));
  NOR4_X1    g03935(.A1(new_n644_), .A2(new_n226_), .A3(new_n306_), .A4(new_n610_), .ZN(new_n4000_));
  NOR4_X1    g03936(.A1(new_n591_), .A2(new_n817_), .A3(new_n715_), .A4(new_n376_), .ZN(new_n4001_));
  NOR4_X1    g03937(.A1(new_n3999_), .A2(new_n3998_), .A3(new_n4000_), .A4(new_n4001_), .ZN(new_n4002_));
  INV_X1     g03938(.I(new_n4002_), .ZN(new_n4003_));
  NOR3_X1    g03939(.A1(new_n3993_), .A2(new_n3996_), .A3(new_n4003_), .ZN(new_n4004_));
  NAND3_X1   g03940(.A1(new_n4004_), .A2(new_n3975_), .A3(new_n3986_), .ZN(new_n4005_));
  INV_X1     g03941(.I(new_n4005_), .ZN(new_n4006_));
  NOR2_X1    g03942(.A1(new_n4006_), .A2(\a[8] ), .ZN(new_n4007_));
  NOR2_X1    g03943(.A1(new_n4007_), .A2(new_n3959_), .ZN(new_n4008_));
  INV_X1     g03944(.I(\a[8] ), .ZN(new_n4009_));
  NOR2_X1    g03945(.A1(new_n4005_), .A2(new_n4009_), .ZN(new_n4010_));
  NOR2_X1    g03946(.A1(new_n4008_), .A2(new_n4010_), .ZN(new_n4011_));
  NAND2_X1   g03947(.A1(new_n4011_), .A2(new_n3862_), .ZN(new_n4012_));
  NAND2_X1   g03948(.A1(new_n3920_), .A2(new_n4012_), .ZN(new_n4013_));
  INV_X1     g03949(.I(new_n3862_), .ZN(new_n4014_));
  OAI21_X1   g03950(.A1(new_n4008_), .A2(new_n4010_), .B(new_n4014_), .ZN(new_n4015_));
  NAND2_X1   g03951(.A1(new_n4013_), .A2(new_n4015_), .ZN(new_n4016_));
  NOR4_X1    g03952(.A1(new_n681_), .A2(new_n456_), .A3(new_n320_), .A4(new_n744_), .ZN(new_n4017_));
  NOR3_X1    g03953(.A1(new_n1415_), .A2(new_n640_), .A3(new_n343_), .ZN(new_n4018_));
  INV_X1     g03954(.I(new_n4018_), .ZN(new_n4019_));
  NAND3_X1   g03955(.A1(new_n399_), .A2(new_n1646_), .A3(new_n1832_), .ZN(new_n4020_));
  NOR4_X1    g03956(.A1(new_n4019_), .A2(new_n4020_), .A3(new_n2472_), .A4(new_n4017_), .ZN(new_n4021_));
  INV_X1     g03957(.I(new_n1745_), .ZN(new_n4022_));
  NAND4_X1   g03958(.A1(new_n599_), .A2(new_n293_), .A3(new_n521_), .A4(new_n1590_), .ZN(new_n4023_));
  NAND2_X1   g03959(.A1(new_n4023_), .A2(new_n1700_), .ZN(new_n4024_));
  NAND3_X1   g03960(.A1(new_n1105_), .A2(new_n1853_), .A3(new_n739_), .ZN(new_n4025_));
  NOR4_X1    g03961(.A1(new_n4024_), .A2(new_n1499_), .A3(new_n4025_), .A4(new_n4022_), .ZN(new_n4026_));
  NAND2_X1   g03962(.A1(new_n4021_), .A2(new_n4026_), .ZN(new_n4027_));
  NOR4_X1    g03963(.A1(new_n4027_), .A2(new_n2187_), .A3(new_n2335_), .A4(new_n2831_), .ZN(new_n4028_));
  NAND2_X1   g03964(.A1(new_n4028_), .A2(new_n1051_), .ZN(new_n4029_));
  NAND2_X1   g03965(.A1(new_n4029_), .A2(new_n3862_), .ZN(new_n4030_));
  NOR2_X1    g03966(.A1(new_n4029_), .A2(new_n3862_), .ZN(new_n4031_));
  AOI21_X1   g03967(.A1(new_n4016_), .A2(new_n4030_), .B(new_n4031_), .ZN(new_n4032_));
  AOI21_X1   g03968(.A1(new_n3887_), .A2(new_n3888_), .B(new_n4014_), .ZN(new_n4033_));
  INV_X1     g03969(.I(\a[11] ), .ZN(new_n4034_));
  XOR2_X1    g03970(.A1(new_n3885_), .A2(new_n4034_), .Z(new_n4035_));
  NOR2_X1    g03971(.A1(new_n4035_), .A2(new_n3862_), .ZN(new_n4036_));
  NOR2_X1    g03972(.A1(new_n4036_), .A2(new_n4033_), .ZN(new_n4037_));
  NAND2_X1   g03973(.A1(new_n4032_), .A2(new_n4037_), .ZN(new_n4038_));
  NAND2_X1   g03974(.A1(new_n4038_), .A2(new_n3908_), .ZN(new_n4039_));
  NOR2_X1    g03975(.A1(new_n4032_), .A2(new_n4037_), .ZN(new_n4040_));
  INV_X1     g03976(.I(new_n4040_), .ZN(new_n4041_));
  NAND2_X1   g03977(.A1(new_n4039_), .A2(new_n4041_), .ZN(new_n4042_));
  NOR2_X1    g03978(.A1(new_n3899_), .A2(new_n4042_), .ZN(new_n4043_));
  INV_X1     g03979(.I(new_n4043_), .ZN(new_n4044_));
  NAND2_X1   g03980(.A1(new_n3899_), .A2(new_n4042_), .ZN(new_n4045_));
  INV_X1     g03981(.I(new_n4045_), .ZN(new_n4046_));
  AOI21_X1   g03982(.A1(new_n3817_), .A2(new_n4044_), .B(new_n4046_), .ZN(new_n4047_));
  INV_X1     g03983(.I(new_n4047_), .ZN(new_n4048_));
  OAI21_X1   g03984(.A1(new_n3696_), .A2(new_n3698_), .B(new_n3660_), .ZN(new_n4049_));
  XOR2_X1    g03985(.A1(new_n3517_), .A2(new_n3694_), .Z(new_n4050_));
  OAI21_X1   g03986(.A1(new_n3660_), .A2(new_n4050_), .B(new_n4049_), .ZN(new_n4051_));
  AOI21_X1   g03987(.A1(new_n3895_), .A2(new_n3893_), .B(new_n3891_), .ZN(new_n4052_));
  INV_X1     g03988(.I(new_n4052_), .ZN(new_n4053_));
  NOR2_X1    g03989(.A1(new_n4051_), .A2(new_n4053_), .ZN(new_n4054_));
  INV_X1     g03990(.I(new_n4054_), .ZN(new_n4055_));
  AND2_X2    g03991(.A1(new_n4051_), .A2(new_n4053_), .Z(new_n4056_));
  AOI21_X1   g03992(.A1(new_n4048_), .A2(new_n4055_), .B(new_n4056_), .ZN(new_n4057_));
  INV_X1     g03993(.I(new_n4057_), .ZN(new_n4058_));
  AOI21_X1   g03994(.A1(new_n3724_), .A2(new_n3720_), .B(new_n3699_), .ZN(new_n4059_));
  XOR2_X1    g03995(.A1(new_n3722_), .A2(new_n3718_), .Z(new_n4060_));
  NOR2_X1    g03996(.A1(new_n4060_), .A2(new_n3700_), .ZN(new_n4061_));
  NOR2_X1    g03997(.A1(new_n4061_), .A2(new_n4059_), .ZN(new_n4062_));
  INV_X1     g03998(.I(new_n4062_), .ZN(new_n4063_));
  NOR2_X1    g03999(.A1(new_n4058_), .A2(new_n4063_), .ZN(new_n4064_));
  INV_X1     g04000(.I(new_n4064_), .ZN(new_n4065_));
  NOR2_X1    g04001(.A1(new_n4057_), .A2(new_n4062_), .ZN(new_n4066_));
  AOI21_X1   g04002(.A1(new_n4065_), .A2(new_n3811_), .B(new_n4066_), .ZN(new_n4067_));
  NOR2_X1    g04003(.A1(new_n3805_), .A2(new_n4067_), .ZN(new_n4068_));
  XOR2_X1    g04004(.A1(new_n3644_), .A2(new_n3725_), .Z(new_n4069_));
  INV_X1     g04005(.I(new_n4069_), .ZN(new_n4070_));
  INV_X1     g04006(.I(new_n3728_), .ZN(new_n4071_));
  AOI21_X1   g04007(.A1(new_n4071_), .A2(new_n3727_), .B(new_n3640_), .ZN(new_n4072_));
  AOI21_X1   g04008(.A1(new_n3640_), .A2(new_n4070_), .B(new_n4072_), .ZN(new_n4073_));
  INV_X1     g04009(.I(new_n3805_), .ZN(new_n4074_));
  INV_X1     g04010(.I(new_n4067_), .ZN(new_n4075_));
  NOR2_X1    g04011(.A1(new_n4074_), .A2(new_n4075_), .ZN(new_n4076_));
  INV_X1     g04012(.I(new_n4076_), .ZN(new_n4077_));
  AOI21_X1   g04013(.A1(new_n4077_), .A2(new_n4073_), .B(new_n4068_), .ZN(new_n4078_));
  INV_X1     g04014(.I(new_n4078_), .ZN(new_n4079_));
  NOR2_X1    g04015(.A1(new_n3800_), .A2(new_n4079_), .ZN(new_n4080_));
  INV_X1     g04016(.I(new_n4080_), .ZN(new_n4081_));
  AND2_X2    g04017(.A1(new_n3800_), .A2(new_n4079_), .Z(new_n4082_));
  AOI21_X1   g04018(.A1(new_n3797_), .A2(new_n4081_), .B(new_n4082_), .ZN(new_n4083_));
  INV_X1     g04019(.I(new_n4083_), .ZN(new_n4084_));
  NOR2_X1    g04020(.A1(new_n3791_), .A2(new_n4084_), .ZN(new_n4085_));
  INV_X1     g04021(.I(new_n4085_), .ZN(new_n4086_));
  NOR3_X1    g04022(.A1(new_n4083_), .A2(new_n3790_), .A3(new_n3789_), .ZN(new_n4087_));
  AOI21_X1   g04023(.A1(new_n4086_), .A2(new_n3787_), .B(new_n4087_), .ZN(new_n4088_));
  AND2_X2    g04024(.A1(new_n4088_), .A2(new_n3779_), .Z(new_n4089_));
  NOR2_X1    g04025(.A1(new_n4088_), .A2(new_n3779_), .ZN(new_n4090_));
  NOR2_X1    g04026(.A1(new_n4089_), .A2(new_n4090_), .ZN(new_n4091_));
  XOR2_X1    g04027(.A1(new_n4088_), .A2(new_n3779_), .Z(new_n4092_));
  NAND2_X1   g04028(.A1(new_n4092_), .A2(new_n3753_), .ZN(new_n4093_));
  OAI21_X1   g04029(.A1(new_n3753_), .A2(new_n4091_), .B(new_n4093_), .ZN(new_n4094_));
  INV_X1     g04030(.I(new_n3773_), .ZN(new_n4095_));
  NOR2_X1    g04031(.A1(new_n3763_), .A2(new_n3772_), .ZN(new_n4096_));
  INV_X1     g04032(.I(new_n4096_), .ZN(new_n4097_));
  OAI22_X1   g04033(.A1(new_n3176_), .A2(new_n4097_), .B1(new_n2665_), .B2(new_n3769_), .ZN(new_n4098_));
  NAND2_X1   g04034(.A1(new_n2728_), .A2(new_n3776_), .ZN(new_n4099_));
  AOI21_X1   g04035(.A1(new_n4098_), .A2(new_n4099_), .B(new_n4095_), .ZN(new_n4100_));
  NAND2_X1   g04036(.A1(new_n3273_), .A2(new_n4100_), .ZN(new_n4101_));
  XOR2_X1    g04037(.A1(new_n4101_), .A2(\a[20] ), .Z(new_n4102_));
  INV_X1     g04038(.I(new_n4102_), .ZN(new_n4103_));
  OAI21_X1   g04039(.A1(new_n4082_), .A2(new_n4080_), .B(new_n3797_), .ZN(new_n4104_));
  XOR2_X1    g04040(.A1(new_n3800_), .A2(new_n4078_), .Z(new_n4105_));
  OAI21_X1   g04041(.A1(new_n3797_), .A2(new_n4105_), .B(new_n4104_), .ZN(new_n4106_));
  OAI22_X1   g04042(.A1(new_n2559_), .A2(new_n3310_), .B1(new_n694_), .B2(new_n3780_), .ZN(new_n4107_));
  NAND2_X1   g04043(.A1(new_n2567_), .A2(new_n3782_), .ZN(new_n4108_));
  AOI21_X1   g04044(.A1(new_n4107_), .A2(new_n4108_), .B(new_n3302_), .ZN(new_n4109_));
  NAND2_X1   g04045(.A1(new_n2759_), .A2(new_n4109_), .ZN(new_n4110_));
  XOR2_X1    g04046(.A1(new_n4110_), .A2(\a[23] ), .Z(new_n4111_));
  INV_X1     g04047(.I(new_n4111_), .ZN(new_n4112_));
  XNOR2_X1   g04048(.A1(new_n3805_), .A2(new_n4067_), .ZN(new_n4113_));
  OAI21_X1   g04049(.A1(new_n4076_), .A2(new_n4068_), .B(new_n4073_), .ZN(new_n4114_));
  OAI21_X1   g04050(.A1(new_n4073_), .A2(new_n4113_), .B(new_n4114_), .ZN(new_n4115_));
  OAI22_X1   g04051(.A1(new_n896_), .A2(new_n3318_), .B1(new_n1180_), .B2(new_n3268_), .ZN(new_n4116_));
  NAND2_X1   g04052(.A1(new_n2504_), .A2(new_n3323_), .ZN(new_n4117_));
  AOI21_X1   g04053(.A1(new_n4117_), .A2(new_n4116_), .B(new_n3260_), .ZN(new_n4118_));
  NAND2_X1   g04054(.A1(new_n3596_), .A2(new_n4118_), .ZN(new_n4119_));
  XOR2_X1    g04055(.A1(new_n4119_), .A2(\a[26] ), .Z(new_n4120_));
  INV_X1     g04056(.I(new_n4120_), .ZN(new_n4121_));
  XOR2_X1    g04057(.A1(new_n4057_), .A2(new_n4063_), .Z(new_n4122_));
  OAI21_X1   g04058(.A1(new_n4064_), .A2(new_n4066_), .B(new_n3810_), .ZN(new_n4123_));
  OAI21_X1   g04059(.A1(new_n4122_), .A2(new_n3810_), .B(new_n4123_), .ZN(new_n4124_));
  INV_X1     g04060(.I(new_n4124_), .ZN(new_n4125_));
  OAI22_X1   g04061(.A1(new_n1008_), .A2(new_n3318_), .B1(new_n1121_), .B2(new_n3268_), .ZN(new_n4126_));
  NAND2_X1   g04062(.A1(new_n1181_), .A2(new_n3323_), .ZN(new_n4127_));
  AOI21_X1   g04063(.A1(new_n4126_), .A2(new_n4127_), .B(new_n3260_), .ZN(new_n4128_));
  NAND2_X1   g04064(.A1(new_n3562_), .A2(new_n4128_), .ZN(new_n4129_));
  XOR2_X1    g04065(.A1(new_n4129_), .A2(\a[26] ), .Z(new_n4130_));
  INV_X1     g04066(.I(new_n4130_), .ZN(new_n4131_));
  XOR2_X1    g04067(.A1(new_n4051_), .A2(new_n4052_), .Z(new_n4132_));
  OAI21_X1   g04068(.A1(new_n4054_), .A2(new_n4056_), .B(new_n4047_), .ZN(new_n4133_));
  OAI21_X1   g04069(.A1(new_n4047_), .A2(new_n4132_), .B(new_n4133_), .ZN(new_n4134_));
  OAI22_X1   g04070(.A1(new_n2492_), .A2(new_n3175_), .B1(new_n2408_), .B2(new_n2747_), .ZN(new_n4135_));
  NAND2_X1   g04071(.A1(new_n2454_), .A2(new_n3275_), .ZN(new_n4136_));
  AOI21_X1   g04072(.A1(new_n4136_), .A2(new_n4135_), .B(new_n2737_), .ZN(new_n4137_));
  NAND2_X1   g04073(.A1(new_n3577_), .A2(new_n4137_), .ZN(new_n4138_));
  XOR2_X1    g04074(.A1(new_n4138_), .A2(\a[29] ), .Z(new_n4139_));
  NAND2_X1   g04075(.A1(new_n4134_), .A2(new_n4139_), .ZN(new_n4140_));
  NOR2_X1    g04076(.A1(new_n4134_), .A2(new_n4139_), .ZN(new_n4141_));
  AOI21_X1   g04077(.A1(new_n4131_), .A2(new_n4140_), .B(new_n4141_), .ZN(new_n4142_));
  INV_X1     g04078(.I(new_n4142_), .ZN(new_n4143_));
  NOR2_X1    g04079(.A1(new_n4125_), .A2(new_n4143_), .ZN(new_n4144_));
  INV_X1     g04080(.I(new_n4144_), .ZN(new_n4145_));
  NOR2_X1    g04081(.A1(new_n4124_), .A2(new_n4142_), .ZN(new_n4146_));
  AOI21_X1   g04082(.A1(new_n4145_), .A2(new_n4121_), .B(new_n4146_), .ZN(new_n4147_));
  INV_X1     g04083(.I(new_n4147_), .ZN(new_n4148_));
  NOR2_X1    g04084(.A1(new_n4148_), .A2(new_n4115_), .ZN(new_n4149_));
  INV_X1     g04085(.I(new_n4149_), .ZN(new_n4150_));
  NAND2_X1   g04086(.A1(new_n4148_), .A2(new_n4115_), .ZN(new_n4151_));
  INV_X1     g04087(.I(new_n4151_), .ZN(new_n4152_));
  AOI21_X1   g04088(.A1(new_n4112_), .A2(new_n4150_), .B(new_n4152_), .ZN(new_n4153_));
  INV_X1     g04089(.I(new_n4153_), .ZN(new_n4154_));
  NOR2_X1    g04090(.A1(new_n4106_), .A2(new_n4154_), .ZN(new_n4155_));
  INV_X1     g04091(.I(new_n4155_), .ZN(new_n4156_));
  AND2_X2    g04092(.A1(new_n4106_), .A2(new_n4154_), .Z(new_n4157_));
  AOI21_X1   g04093(.A1(new_n4156_), .A2(new_n4103_), .B(new_n4157_), .ZN(new_n4158_));
  XOR2_X1    g04094(.A1(new_n3791_), .A2(new_n4083_), .Z(new_n4159_));
  OAI21_X1   g04095(.A1(new_n4085_), .A2(new_n4087_), .B(new_n3786_), .ZN(new_n4160_));
  OAI21_X1   g04096(.A1(new_n4159_), .A2(new_n3786_), .B(new_n4160_), .ZN(new_n4161_));
  INV_X1     g04097(.I(new_n4161_), .ZN(new_n4162_));
  OAI22_X1   g04098(.A1(new_n3176_), .A2(new_n3775_), .B1(new_n3142_), .B2(new_n4097_), .ZN(new_n4163_));
  NAND2_X1   g04099(.A1(new_n2728_), .A2(new_n3770_), .ZN(new_n4164_));
  AOI21_X1   g04100(.A1(new_n4163_), .A2(new_n4164_), .B(new_n4095_), .ZN(new_n4165_));
  NAND2_X1   g04101(.A1(new_n3174_), .A2(new_n4165_), .ZN(new_n4166_));
  XOR2_X1    g04102(.A1(new_n4166_), .A2(\a[20] ), .Z(new_n4167_));
  INV_X1     g04103(.I(new_n4167_), .ZN(new_n4168_));
  NOR2_X1    g04104(.A1(new_n4162_), .A2(new_n4168_), .ZN(new_n4169_));
  NOR2_X1    g04105(.A1(new_n4169_), .A2(new_n4158_), .ZN(new_n4170_));
  NOR2_X1    g04106(.A1(new_n4161_), .A2(new_n4167_), .ZN(new_n4171_));
  NOR2_X1    g04107(.A1(new_n4170_), .A2(new_n4171_), .ZN(new_n4172_));
  NOR2_X1    g04108(.A1(new_n4094_), .A2(new_n4172_), .ZN(new_n4173_));
  INV_X1     g04109(.I(new_n4173_), .ZN(new_n4174_));
  OAI22_X1   g04110(.A1(new_n2614_), .A2(new_n3769_), .B1(new_n2665_), .B2(new_n3775_), .ZN(new_n4175_));
  NAND2_X1   g04111(.A1(new_n2728_), .A2(new_n4096_), .ZN(new_n4176_));
  AOI21_X1   g04112(.A1(new_n4176_), .A2(new_n4175_), .B(new_n4095_), .ZN(new_n4177_));
  NAND2_X1   g04113(.A1(new_n2733_), .A2(new_n4177_), .ZN(new_n4178_));
  XOR2_X1    g04114(.A1(new_n4178_), .A2(\a[20] ), .Z(new_n4179_));
  AOI21_X1   g04115(.A1(new_n4150_), .A2(new_n4151_), .B(new_n4111_), .ZN(new_n4180_));
  XOR2_X1    g04116(.A1(new_n4115_), .A2(new_n4147_), .Z(new_n4181_));
  NOR2_X1    g04117(.A1(new_n4181_), .A2(new_n4112_), .ZN(new_n4182_));
  NOR2_X1    g04118(.A1(new_n4180_), .A2(new_n4182_), .ZN(new_n4183_));
  OAI22_X1   g04119(.A1(new_n813_), .A2(new_n3310_), .B1(new_n529_), .B2(new_n3780_), .ZN(new_n4184_));
  NAND2_X1   g04120(.A1(new_n2563_), .A2(new_n3782_), .ZN(new_n4185_));
  AOI21_X1   g04121(.A1(new_n4185_), .A2(new_n4184_), .B(new_n3302_), .ZN(new_n4186_));
  NAND2_X1   g04122(.A1(new_n3051_), .A2(new_n4186_), .ZN(new_n4187_));
  XOR2_X1    g04123(.A1(new_n4187_), .A2(\a[23] ), .Z(new_n4188_));
  INV_X1     g04124(.I(new_n4188_), .ZN(new_n4189_));
  XOR2_X1    g04125(.A1(new_n4124_), .A2(new_n4143_), .Z(new_n4190_));
  OAI21_X1   g04126(.A1(new_n4144_), .A2(new_n4146_), .B(new_n4120_), .ZN(new_n4191_));
  OAI21_X1   g04127(.A1(new_n4120_), .A2(new_n4190_), .B(new_n4191_), .ZN(new_n4192_));
  INV_X1     g04128(.I(new_n4192_), .ZN(new_n4193_));
  OAI22_X1   g04129(.A1(new_n2559_), .A2(new_n3780_), .B1(new_n896_), .B2(new_n3310_), .ZN(new_n4194_));
  NAND2_X1   g04130(.A1(new_n814_), .A2(new_n3782_), .ZN(new_n4195_));
  AOI21_X1   g04131(.A1(new_n4194_), .A2(new_n4195_), .B(new_n3302_), .ZN(new_n4196_));
  NAND2_X1   g04132(.A1(new_n3624_), .A2(new_n4196_), .ZN(new_n4197_));
  XOR2_X1    g04133(.A1(new_n4197_), .A2(\a[23] ), .Z(new_n4198_));
  INV_X1     g04134(.I(new_n4198_), .ZN(new_n4199_));
  INV_X1     g04135(.I(new_n4140_), .ZN(new_n4200_));
  OAI21_X1   g04136(.A1(new_n4200_), .A2(new_n4141_), .B(new_n4131_), .ZN(new_n4201_));
  XOR2_X1    g04137(.A1(new_n4134_), .A2(new_n4139_), .Z(new_n4202_));
  NAND2_X1   g04138(.A1(new_n4202_), .A2(new_n4130_), .ZN(new_n4203_));
  NAND2_X1   g04139(.A1(new_n4203_), .A2(new_n4201_), .ZN(new_n4204_));
  OAI22_X1   g04140(.A1(new_n1180_), .A2(new_n3318_), .B1(new_n2492_), .B2(new_n3268_), .ZN(new_n4205_));
  NAND2_X1   g04141(.A1(new_n1122_), .A2(new_n3323_), .ZN(new_n4206_));
  AOI21_X1   g04142(.A1(new_n4206_), .A2(new_n4205_), .B(new_n3260_), .ZN(new_n4207_));
  NAND2_X1   g04143(.A1(new_n3330_), .A2(new_n4207_), .ZN(new_n4208_));
  XOR2_X1    g04144(.A1(new_n4208_), .A2(\a[26] ), .Z(new_n4209_));
  INV_X1     g04145(.I(new_n4209_), .ZN(new_n4210_));
  XOR2_X1    g04146(.A1(new_n4042_), .A2(new_n3898_), .Z(new_n4211_));
  NOR2_X1    g04147(.A1(new_n4211_), .A2(new_n3816_), .ZN(new_n4212_));
  AOI21_X1   g04148(.A1(new_n4044_), .A2(new_n4045_), .B(new_n3817_), .ZN(new_n4213_));
  NOR2_X1    g04149(.A1(new_n4213_), .A2(new_n4212_), .ZN(new_n4214_));
  OAI22_X1   g04150(.A1(new_n1409_), .A2(new_n2747_), .B1(new_n2367_), .B2(new_n3175_), .ZN(new_n4215_));
  NAND2_X1   g04151(.A1(new_n1334_), .A2(new_n3275_), .ZN(new_n4216_));
  AOI21_X1   g04152(.A1(new_n4215_), .A2(new_n4216_), .B(new_n2737_), .ZN(new_n4217_));
  NAND2_X1   g04153(.A1(new_n3654_), .A2(new_n4217_), .ZN(new_n4218_));
  XOR2_X1    g04154(.A1(new_n4218_), .A2(new_n74_), .Z(new_n4219_));
  INV_X1     g04155(.I(new_n4031_), .ZN(new_n4220_));
  AOI22_X1   g04156(.A1(new_n4013_), .A2(new_n4015_), .B1(new_n4030_), .B2(new_n4220_), .ZN(new_n4221_));
  XOR2_X1    g04157(.A1(new_n4029_), .A2(new_n4014_), .Z(new_n4222_));
  NOR2_X1    g04158(.A1(new_n4016_), .A2(new_n4222_), .ZN(new_n4223_));
  NOR2_X1    g04159(.A1(new_n4223_), .A2(new_n4221_), .ZN(new_n4224_));
  XNOR2_X1   g04160(.A1(new_n1453_), .A2(new_n2351_), .ZN(new_n4225_));
  INV_X1     g04161(.I(new_n4225_), .ZN(new_n4226_));
  OAI21_X1   g04162(.A1(new_n2353_), .A2(new_n2355_), .B(new_n4226_), .ZN(new_n4227_));
  NOR2_X1    g04163(.A1(new_n2360_), .A2(new_n2356_), .ZN(new_n4228_));
  NOR3_X1    g04164(.A1(new_n2353_), .A2(new_n2355_), .A3(new_n4228_), .ZN(new_n4229_));
  INV_X1     g04165(.I(new_n4229_), .ZN(new_n4230_));
  NAND2_X1   g04166(.A1(new_n4230_), .A2(new_n4227_), .ZN(new_n4231_));
  AOI21_X1   g04167(.A1(new_n2354_), .A2(new_n3189_), .B(new_n2763_), .ZN(new_n4232_));
  OAI21_X1   g04168(.A1(new_n2311_), .A2(new_n2771_), .B(new_n4232_), .ZN(new_n4233_));
  AOI21_X1   g04169(.A1(new_n2359_), .A2(new_n3332_), .B(new_n4233_), .ZN(new_n4234_));
  AND2_X2    g04170(.A1(new_n4231_), .A2(new_n4234_), .Z(new_n4235_));
  INV_X1     g04171(.I(new_n4235_), .ZN(new_n4236_));
  NAND2_X1   g04172(.A1(new_n4224_), .A2(new_n4236_), .ZN(new_n4237_));
  NAND2_X1   g04173(.A1(new_n4219_), .A2(new_n4237_), .ZN(new_n4238_));
  OAI21_X1   g04174(.A1(new_n4223_), .A2(new_n4221_), .B(new_n4235_), .ZN(new_n4239_));
  AND2_X2    g04175(.A1(new_n4238_), .A2(new_n4239_), .Z(new_n4240_));
  INV_X1     g04176(.I(new_n4240_), .ZN(new_n4241_));
  XNOR2_X1   g04177(.A1(new_n4032_), .A2(new_n4037_), .ZN(new_n4242_));
  INV_X1     g04178(.I(new_n4242_), .ZN(new_n4243_));
  AOI21_X1   g04179(.A1(new_n4041_), .A2(new_n4038_), .B(new_n3908_), .ZN(new_n4244_));
  AOI21_X1   g04180(.A1(new_n4243_), .A2(new_n3908_), .B(new_n4244_), .ZN(new_n4245_));
  OAI22_X1   g04181(.A1(new_n2367_), .A2(new_n2742_), .B1(new_n2408_), .B2(new_n3175_), .ZN(new_n4246_));
  NAND2_X1   g04182(.A1(new_n1334_), .A2(new_n2746_), .ZN(new_n4247_));
  AOI21_X1   g04183(.A1(new_n4246_), .A2(new_n4247_), .B(new_n2737_), .ZN(new_n4248_));
  NAND2_X1   g04184(.A1(new_n3708_), .A2(new_n4248_), .ZN(new_n4249_));
  XOR2_X1    g04185(.A1(new_n4249_), .A2(new_n74_), .Z(new_n4250_));
  NOR2_X1    g04186(.A1(new_n4250_), .A2(new_n4245_), .ZN(new_n4251_));
  INV_X1     g04187(.I(new_n4251_), .ZN(new_n4252_));
  INV_X1     g04188(.I(new_n4245_), .ZN(new_n4253_));
  XOR2_X1    g04189(.A1(new_n4249_), .A2(\a[29] ), .Z(new_n4254_));
  NOR2_X1    g04190(.A1(new_n4253_), .A2(new_n4254_), .ZN(new_n4255_));
  AOI21_X1   g04191(.A1(new_n4252_), .A2(new_n4241_), .B(new_n4255_), .ZN(new_n4256_));
  INV_X1     g04192(.I(new_n4256_), .ZN(new_n4257_));
  NOR2_X1    g04193(.A1(new_n4257_), .A2(new_n4214_), .ZN(new_n4258_));
  INV_X1     g04194(.I(new_n4258_), .ZN(new_n4259_));
  NOR3_X1    g04195(.A1(new_n4256_), .A2(new_n4212_), .A3(new_n4213_), .ZN(new_n4260_));
  AOI21_X1   g04196(.A1(new_n4259_), .A2(new_n4210_), .B(new_n4260_), .ZN(new_n4261_));
  INV_X1     g04197(.I(new_n4261_), .ZN(new_n4262_));
  NOR2_X1    g04198(.A1(new_n4204_), .A2(new_n4262_), .ZN(new_n4263_));
  INV_X1     g04199(.I(new_n4263_), .ZN(new_n4264_));
  NAND2_X1   g04200(.A1(new_n4204_), .A2(new_n4262_), .ZN(new_n4265_));
  INV_X1     g04201(.I(new_n4265_), .ZN(new_n4266_));
  AOI21_X1   g04202(.A1(new_n4199_), .A2(new_n4264_), .B(new_n4266_), .ZN(new_n4267_));
  INV_X1     g04203(.I(new_n4267_), .ZN(new_n4268_));
  NOR2_X1    g04204(.A1(new_n4193_), .A2(new_n4268_), .ZN(new_n4269_));
  INV_X1     g04205(.I(new_n4269_), .ZN(new_n4270_));
  NOR2_X1    g04206(.A1(new_n4192_), .A2(new_n4267_), .ZN(new_n4271_));
  AOI21_X1   g04207(.A1(new_n4270_), .A2(new_n4189_), .B(new_n4271_), .ZN(new_n4272_));
  AND2_X2    g04208(.A1(new_n4183_), .A2(new_n4272_), .Z(new_n4273_));
  NOR2_X1    g04209(.A1(new_n4183_), .A2(new_n4272_), .ZN(new_n4274_));
  NOR2_X1    g04210(.A1(new_n4273_), .A2(new_n4274_), .ZN(new_n4275_));
  NOR2_X1    g04211(.A1(new_n4275_), .A2(new_n4179_), .ZN(new_n4276_));
  INV_X1     g04212(.I(new_n4179_), .ZN(new_n4277_));
  XNOR2_X1   g04213(.A1(new_n4183_), .A2(new_n4272_), .ZN(new_n4278_));
  NOR2_X1    g04214(.A1(new_n4278_), .A2(new_n4277_), .ZN(new_n4279_));
  NOR2_X1    g04215(.A1(new_n4276_), .A2(new_n4279_), .ZN(new_n4280_));
  INV_X1     g04216(.I(\a[15] ), .ZN(new_n4281_));
  NOR2_X1    g04217(.A1(new_n4281_), .A2(\a[14] ), .ZN(new_n4282_));
  NOR2_X1    g04218(.A1(new_n3521_), .A2(\a[15] ), .ZN(new_n4283_));
  NOR2_X1    g04219(.A1(new_n4282_), .A2(new_n4283_), .ZN(new_n4284_));
  INV_X1     g04220(.I(new_n4284_), .ZN(new_n4285_));
  INV_X1     g04221(.I(\a[16] ), .ZN(new_n4286_));
  NOR2_X1    g04222(.A1(new_n4286_), .A2(\a[14] ), .ZN(new_n4287_));
  NOR2_X1    g04223(.A1(new_n3521_), .A2(\a[16] ), .ZN(new_n4288_));
  OR2_X2     g04224(.A1(new_n4287_), .A2(new_n4288_), .Z(new_n4289_));
  XNOR2_X1   g04225(.A1(\a[14] ), .A2(\a[17] ), .ZN(new_n4290_));
  OAI21_X1   g04226(.A1(new_n4285_), .A2(new_n4289_), .B(new_n4290_), .ZN(new_n4291_));
  INV_X1     g04227(.I(new_n4291_), .ZN(new_n4292_));
  NAND2_X1   g04228(.A1(new_n3168_), .A2(new_n4292_), .ZN(new_n4293_));
  XNOR2_X1   g04229(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n4294_));
  NOR2_X1    g04230(.A1(new_n4284_), .A2(new_n4294_), .ZN(new_n4295_));
  NOR3_X1    g04231(.A1(new_n4286_), .A2(\a[14] ), .A3(\a[15] ), .ZN(new_n4296_));
  AOI21_X1   g04232(.A1(\a[15] ), .A2(new_n4288_), .B(new_n4296_), .ZN(new_n4297_));
  INV_X1     g04233(.I(new_n4297_), .ZN(new_n4298_));
  NAND2_X1   g04234(.A1(new_n3247_), .A2(new_n4298_), .ZN(new_n4299_));
  NAND4_X1   g04235(.A1(new_n3758_), .A2(new_n4293_), .A3(new_n4295_), .A4(new_n4299_), .ZN(new_n4300_));
  XOR2_X1    g04236(.A1(new_n4300_), .A2(\a[17] ), .Z(new_n4301_));
  INV_X1     g04237(.I(new_n4301_), .ZN(new_n4302_));
  OAI22_X1   g04238(.A1(new_n694_), .A2(new_n3769_), .B1(new_n2665_), .B2(new_n4097_), .ZN(new_n4303_));
  NAND2_X1   g04239(.A1(new_n2615_), .A2(new_n3776_), .ZN(new_n4304_));
  AOI21_X1   g04240(.A1(new_n4303_), .A2(new_n4304_), .B(new_n4095_), .ZN(new_n4305_));
  NAND2_X1   g04241(.A1(new_n3188_), .A2(new_n4305_), .ZN(new_n4306_));
  XOR2_X1    g04242(.A1(new_n4306_), .A2(\a[20] ), .Z(new_n4307_));
  XNOR2_X1   g04243(.A1(new_n4192_), .A2(new_n4267_), .ZN(new_n4308_));
  OAI21_X1   g04244(.A1(new_n4269_), .A2(new_n4271_), .B(new_n4188_), .ZN(new_n4309_));
  OAI21_X1   g04245(.A1(new_n4308_), .A2(new_n4188_), .B(new_n4309_), .ZN(new_n4310_));
  INV_X1     g04246(.I(new_n4310_), .ZN(new_n4311_));
  OAI22_X1   g04247(.A1(new_n2614_), .A2(new_n4097_), .B1(new_n529_), .B2(new_n3769_), .ZN(new_n4312_));
  NAND2_X1   g04248(.A1(new_n2718_), .A2(new_n3776_), .ZN(new_n4313_));
  AOI21_X1   g04249(.A1(new_n4313_), .A2(new_n4312_), .B(new_n4095_), .ZN(new_n4314_));
  NAND2_X1   g04250(.A1(new_n3074_), .A2(new_n4314_), .ZN(new_n4315_));
  XOR2_X1    g04251(.A1(new_n4315_), .A2(\a[20] ), .Z(new_n4316_));
  INV_X1     g04252(.I(new_n4316_), .ZN(new_n4317_));
  AOI21_X1   g04253(.A1(new_n4264_), .A2(new_n4265_), .B(new_n4198_), .ZN(new_n4318_));
  XOR2_X1    g04254(.A1(new_n4204_), .A2(new_n4261_), .Z(new_n4319_));
  NOR2_X1    g04255(.A1(new_n4319_), .A2(new_n4199_), .ZN(new_n4320_));
  NOR2_X1    g04256(.A1(new_n4320_), .A2(new_n4318_), .ZN(new_n4321_));
  OAI21_X1   g04257(.A1(new_n4258_), .A2(new_n4260_), .B(new_n4210_), .ZN(new_n4322_));
  XOR2_X1    g04258(.A1(new_n4214_), .A2(new_n4256_), .Z(new_n4323_));
  OAI21_X1   g04259(.A1(new_n4323_), .A2(new_n4210_), .B(new_n4322_), .ZN(new_n4324_));
  OAI22_X1   g04260(.A1(new_n813_), .A2(new_n3780_), .B1(new_n1008_), .B2(new_n3310_), .ZN(new_n4325_));
  NAND2_X1   g04261(.A1(new_n897_), .A2(new_n3782_), .ZN(new_n4326_));
  AOI21_X1   g04262(.A1(new_n4325_), .A2(new_n4326_), .B(new_n3302_), .ZN(new_n4327_));
  NAND2_X1   g04263(.A1(new_n2917_), .A2(new_n4327_), .ZN(new_n4328_));
  XOR2_X1    g04264(.A1(new_n4328_), .A2(\a[23] ), .Z(new_n4329_));
  INV_X1     g04265(.I(new_n4329_), .ZN(new_n4330_));
  OAI22_X1   g04266(.A1(new_n1121_), .A2(new_n3318_), .B1(new_n2451_), .B2(new_n3268_), .ZN(new_n4331_));
  NAND2_X1   g04267(.A1(new_n2496_), .A2(new_n3323_), .ZN(new_n4332_));
  AOI21_X1   g04268(.A1(new_n4331_), .A2(new_n4332_), .B(new_n3260_), .ZN(new_n4333_));
  NAND2_X1   g04269(.A1(new_n3393_), .A2(new_n4333_), .ZN(new_n4334_));
  XOR2_X1    g04270(.A1(new_n4334_), .A2(\a[26] ), .Z(new_n4335_));
  INV_X1     g04271(.I(new_n4335_), .ZN(new_n4336_));
  OAI22_X1   g04272(.A1(new_n2492_), .A2(new_n3318_), .B1(new_n2408_), .B2(new_n3268_), .ZN(new_n4337_));
  NAND2_X1   g04273(.A1(new_n2454_), .A2(new_n3323_), .ZN(new_n4338_));
  AOI21_X1   g04274(.A1(new_n4338_), .A2(new_n4337_), .B(new_n3260_), .ZN(new_n4339_));
  NAND2_X1   g04275(.A1(new_n3577_), .A2(new_n4339_), .ZN(new_n4340_));
  XOR2_X1    g04276(.A1(new_n4340_), .A2(\a[26] ), .Z(new_n4341_));
  INV_X1     g04277(.I(new_n4341_), .ZN(new_n4342_));
  NAND2_X1   g04278(.A1(new_n4237_), .A2(new_n4239_), .ZN(new_n4343_));
  XOR2_X1    g04279(.A1(new_n4224_), .A2(new_n4235_), .Z(new_n4344_));
  NOR2_X1    g04280(.A1(new_n4344_), .A2(new_n4219_), .ZN(new_n4345_));
  AOI21_X1   g04281(.A1(new_n4219_), .A2(new_n4343_), .B(new_n4345_), .ZN(new_n4346_));
  OAI22_X1   g04282(.A1(new_n1409_), .A2(new_n2742_), .B1(new_n1333_), .B2(new_n3175_), .ZN(new_n4347_));
  NAND2_X1   g04283(.A1(new_n2359_), .A2(new_n2746_), .ZN(new_n4348_));
  AOI21_X1   g04284(.A1(new_n4347_), .A2(new_n4348_), .B(new_n2737_), .ZN(new_n4349_));
  NAND2_X1   g04285(.A1(new_n3828_), .A2(new_n4349_), .ZN(new_n4350_));
  XOR2_X1    g04286(.A1(new_n4350_), .A2(\a[29] ), .Z(new_n4351_));
  INV_X1     g04287(.I(new_n4351_), .ZN(new_n4352_));
  AOI21_X1   g04288(.A1(new_n4012_), .A2(new_n4015_), .B(new_n3919_), .ZN(new_n4353_));
  XOR2_X1    g04289(.A1(new_n4011_), .A2(new_n4014_), .Z(new_n4354_));
  NOR2_X1    g04290(.A1(new_n3920_), .A2(new_n4354_), .ZN(new_n4355_));
  NOR2_X1    g04291(.A1(new_n4355_), .A2(new_n4353_), .ZN(new_n4356_));
  XOR2_X1    g04292(.A1(new_n1547_), .A2(new_n1503_), .Z(new_n4357_));
  INV_X1     g04293(.I(new_n4357_), .ZN(new_n4358_));
  OAI21_X1   g04294(.A1(new_n2206_), .A2(new_n2207_), .B(new_n4358_), .ZN(new_n4359_));
  XNOR2_X1   g04295(.A1(new_n1547_), .A2(new_n1503_), .ZN(new_n4360_));
  INV_X1     g04296(.I(new_n4360_), .ZN(new_n4361_));
  NAND2_X1   g04297(.A1(new_n2254_), .A2(new_n4361_), .ZN(new_n4362_));
  NAND2_X1   g04298(.A1(new_n4362_), .A2(new_n4359_), .ZN(new_n4363_));
  NOR2_X1    g04299(.A1(new_n1503_), .A2(new_n2767_), .ZN(new_n4364_));
  INV_X1     g04300(.I(new_n1547_), .ZN(new_n4365_));
  NOR2_X1    g04301(.A1(new_n4365_), .A2(new_n2772_), .ZN(new_n4366_));
  NOR2_X1    g04302(.A1(new_n2198_), .A2(new_n2771_), .ZN(new_n4367_));
  NOR4_X1    g04303(.A1(new_n4366_), .A2(new_n2763_), .A3(new_n4364_), .A4(new_n4367_), .ZN(new_n4368_));
  NAND2_X1   g04304(.A1(new_n4363_), .A2(new_n4368_), .ZN(new_n4369_));
  INV_X1     g04305(.I(new_n4369_), .ZN(new_n4370_));
  INV_X1     g04306(.I(new_n3959_), .ZN(new_n4371_));
  NOR4_X1    g04307(.A1(new_n465_), .A2(new_n119_), .A3(new_n183_), .A4(new_n955_), .ZN(new_n4372_));
  NOR2_X1    g04308(.A1(new_n930_), .A2(new_n170_), .ZN(new_n4373_));
  NAND4_X1   g04309(.A1(new_n1173_), .A2(new_n309_), .A3(new_n1322_), .A4(new_n4373_), .ZN(new_n4374_));
  NOR4_X1    g04310(.A1(new_n774_), .A2(new_n70_), .A3(new_n235_), .A4(new_n841_), .ZN(new_n4375_));
  NAND4_X1   g04311(.A1(new_n771_), .A2(new_n967_), .A3(new_n1856_), .A4(new_n4375_), .ZN(new_n4376_));
  INV_X1     g04312(.I(new_n2554_), .ZN(new_n4377_));
  NOR4_X1    g04313(.A1(new_n4377_), .A2(new_n258_), .A3(new_n306_), .A4(new_n428_), .ZN(new_n4378_));
  NAND4_X1   g04314(.A1(new_n4378_), .A2(new_n1585_), .A3(new_n521_), .A4(new_n686_), .ZN(new_n4379_));
  INV_X1     g04315(.I(new_n4379_), .ZN(new_n4380_));
  NAND2_X1   g04316(.A1(new_n4380_), .A2(new_n738_), .ZN(new_n4381_));
  NOR4_X1    g04317(.A1(new_n4381_), .A2(new_n4372_), .A3(new_n4374_), .A4(new_n4376_), .ZN(new_n4382_));
  NAND4_X1   g04318(.A1(new_n3446_), .A2(new_n2783_), .A3(new_n2790_), .A4(new_n4382_), .ZN(new_n4383_));
  INV_X1     g04319(.I(new_n4383_), .ZN(new_n4384_));
  NOR2_X1    g04320(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n4385_));
  INV_X1     g04321(.I(new_n4385_), .ZN(new_n4386_));
  INV_X1     g04322(.I(\a[2] ), .ZN(new_n4387_));
  NOR2_X1    g04323(.A1(new_n4387_), .A2(new_n65_), .ZN(new_n4388_));
  AOI21_X1   g04324(.A1(new_n4384_), .A2(new_n4386_), .B(new_n4388_), .ZN(new_n4389_));
  NAND2_X1   g04325(.A1(new_n4389_), .A2(new_n4371_), .ZN(new_n4390_));
  NAND2_X1   g04326(.A1(new_n4370_), .A2(new_n4390_), .ZN(new_n4391_));
  OR2_X2     g04327(.A1(new_n4389_), .A2(new_n4371_), .Z(new_n4392_));
  NAND2_X1   g04328(.A1(new_n4391_), .A2(new_n4392_), .ZN(new_n4393_));
  INV_X1     g04329(.I(new_n3957_), .ZN(new_n4394_));
  NAND4_X1   g04330(.A1(new_n351_), .A2(new_n378_), .A3(new_n1448_), .A4(new_n1465_), .ZN(new_n4395_));
  NAND4_X1   g04331(.A1(new_n272_), .A2(new_n293_), .A3(new_n1572_), .A4(new_n823_), .ZN(new_n4396_));
  NOR3_X1    g04332(.A1(new_n596_), .A2(new_n418_), .A3(new_n715_), .ZN(new_n4397_));
  AND3_X2    g04333(.A1(new_n4395_), .A2(new_n4396_), .A3(new_n4397_), .Z(new_n4398_));
  NOR4_X1    g04334(.A1(new_n2135_), .A2(new_n988_), .A3(new_n2930_), .A4(new_n1134_), .ZN(new_n4399_));
  NAND4_X1   g04335(.A1(new_n4394_), .A2(new_n4399_), .A3(new_n3961_), .A4(new_n4398_), .ZN(new_n4400_));
  NOR4_X1    g04336(.A1(new_n1339_), .A2(new_n407_), .A3(new_n447_), .A4(new_n1984_), .ZN(new_n4401_));
  NAND3_X1   g04337(.A1(new_n1194_), .A2(new_n1585_), .A3(new_n2328_), .ZN(new_n4402_));
  NAND3_X1   g04338(.A1(new_n4401_), .A2(new_n2844_), .A3(new_n4402_), .ZN(new_n4403_));
  NOR3_X1    g04339(.A1(new_n1161_), .A2(new_n202_), .A3(new_n697_), .ZN(new_n4404_));
  NAND4_X1   g04340(.A1(new_n4404_), .A2(new_n1472_), .A3(new_n2339_), .A4(new_n2975_), .ZN(new_n4405_));
  NOR2_X1    g04341(.A1(new_n4403_), .A2(new_n4405_), .ZN(new_n4406_));
  NAND2_X1   g04342(.A1(new_n4406_), .A2(new_n1682_), .ZN(new_n4407_));
  NOR3_X1    g04343(.A1(new_n4407_), .A2(new_n2965_), .A3(new_n4400_), .ZN(new_n4408_));
  NOR2_X1    g04344(.A1(new_n3959_), .A2(new_n4408_), .ZN(new_n4409_));
  INV_X1     g04345(.I(new_n4409_), .ZN(new_n4410_));
  INV_X1     g04346(.I(new_n4408_), .ZN(new_n4411_));
  NOR2_X1    g04347(.A1(new_n4371_), .A2(new_n4411_), .ZN(new_n4412_));
  AOI21_X1   g04348(.A1(new_n4393_), .A2(new_n4410_), .B(new_n4412_), .ZN(new_n4413_));
  INV_X1     g04349(.I(new_n4413_), .ZN(new_n4414_));
  NAND2_X1   g04350(.A1(new_n2253_), .A2(new_n2256_), .ZN(new_n4415_));
  XOR2_X1    g04351(.A1(new_n2310_), .A2(new_n2251_), .Z(new_n4416_));
  NAND2_X1   g04352(.A1(new_n2313_), .A2(new_n2316_), .ZN(new_n4417_));
  NAND2_X1   g04353(.A1(new_n4415_), .A2(new_n4417_), .ZN(new_n4418_));
  OAI21_X1   g04354(.A1(new_n4415_), .A2(new_n4416_), .B(new_n4418_), .ZN(new_n4419_));
  NOR2_X1    g04355(.A1(new_n2311_), .A2(new_n2772_), .ZN(new_n4420_));
  NOR2_X1    g04356(.A1(new_n4365_), .A2(new_n2771_), .ZN(new_n4421_));
  NOR2_X1    g04357(.A1(new_n2251_), .A2(new_n2767_), .ZN(new_n4422_));
  NOR4_X1    g04358(.A1(new_n4420_), .A2(new_n2763_), .A3(new_n4421_), .A4(new_n4422_), .ZN(new_n4423_));
  NAND2_X1   g04359(.A1(new_n4419_), .A2(new_n4423_), .ZN(new_n4424_));
  OAI21_X1   g04360(.A1(new_n4007_), .A2(new_n4010_), .B(new_n4371_), .ZN(new_n4425_));
  XOR2_X1    g04361(.A1(new_n4005_), .A2(\a[8] ), .Z(new_n4426_));
  OAI21_X1   g04362(.A1(new_n4371_), .A2(new_n4426_), .B(new_n4425_), .ZN(new_n4427_));
  INV_X1     g04363(.I(new_n4427_), .ZN(new_n4428_));
  NAND2_X1   g04364(.A1(new_n4424_), .A2(new_n4428_), .ZN(new_n4429_));
  NAND2_X1   g04365(.A1(new_n4414_), .A2(new_n4429_), .ZN(new_n4430_));
  NAND3_X1   g04366(.A1(new_n4419_), .A2(new_n4423_), .A3(new_n4427_), .ZN(new_n4431_));
  NAND2_X1   g04367(.A1(new_n4430_), .A2(new_n4431_), .ZN(new_n4432_));
  INV_X1     g04368(.I(new_n4432_), .ZN(new_n4433_));
  NAND2_X1   g04369(.A1(new_n4433_), .A2(new_n4356_), .ZN(new_n4434_));
  NOR2_X1    g04370(.A1(new_n4433_), .A2(new_n4356_), .ZN(new_n4435_));
  AOI21_X1   g04371(.A1(new_n4352_), .A2(new_n4434_), .B(new_n4435_), .ZN(new_n4436_));
  NAND2_X1   g04372(.A1(new_n4346_), .A2(new_n4436_), .ZN(new_n4437_));
  NOR2_X1    g04373(.A1(new_n4346_), .A2(new_n4436_), .ZN(new_n4438_));
  AOI21_X1   g04374(.A1(new_n4342_), .A2(new_n4437_), .B(new_n4438_), .ZN(new_n4439_));
  NOR2_X1    g04375(.A1(new_n4255_), .A2(new_n4251_), .ZN(new_n4440_));
  NOR2_X1    g04376(.A1(new_n4440_), .A2(new_n4240_), .ZN(new_n4441_));
  XOR2_X1    g04377(.A1(new_n4254_), .A2(new_n4245_), .Z(new_n4442_));
  NOR2_X1    g04378(.A1(new_n4442_), .A2(new_n4241_), .ZN(new_n4443_));
  NOR2_X1    g04379(.A1(new_n4443_), .A2(new_n4441_), .ZN(new_n4444_));
  NAND2_X1   g04380(.A1(new_n4444_), .A2(new_n4439_), .ZN(new_n4445_));
  NOR2_X1    g04381(.A1(new_n4444_), .A2(new_n4439_), .ZN(new_n4446_));
  AOI21_X1   g04382(.A1(new_n4336_), .A2(new_n4445_), .B(new_n4446_), .ZN(new_n4447_));
  INV_X1     g04383(.I(new_n4447_), .ZN(new_n4448_));
  NOR2_X1    g04384(.A1(new_n4330_), .A2(new_n4448_), .ZN(new_n4449_));
  INV_X1     g04385(.I(new_n4449_), .ZN(new_n4450_));
  NOR2_X1    g04386(.A1(new_n4329_), .A2(new_n4447_), .ZN(new_n4451_));
  AOI21_X1   g04387(.A1(new_n4450_), .A2(new_n4324_), .B(new_n4451_), .ZN(new_n4452_));
  NAND2_X1   g04388(.A1(new_n4321_), .A2(new_n4452_), .ZN(new_n4453_));
  NOR2_X1    g04389(.A1(new_n4321_), .A2(new_n4452_), .ZN(new_n4454_));
  AOI21_X1   g04390(.A1(new_n4317_), .A2(new_n4453_), .B(new_n4454_), .ZN(new_n4455_));
  INV_X1     g04391(.I(new_n4455_), .ZN(new_n4456_));
  NOR2_X1    g04392(.A1(new_n4311_), .A2(new_n4456_), .ZN(new_n4457_));
  NOR2_X1    g04393(.A1(new_n4310_), .A2(new_n4455_), .ZN(new_n4458_));
  INV_X1     g04394(.I(new_n4458_), .ZN(new_n4459_));
  OAI21_X1   g04395(.A1(new_n4307_), .A2(new_n4457_), .B(new_n4459_), .ZN(new_n4460_));
  NOR2_X1    g04396(.A1(new_n4460_), .A2(new_n4302_), .ZN(new_n4461_));
  NAND2_X1   g04397(.A1(new_n4460_), .A2(new_n4302_), .ZN(new_n4462_));
  INV_X1     g04398(.I(new_n4462_), .ZN(new_n4463_));
  NOR2_X1    g04399(.A1(new_n4463_), .A2(new_n4461_), .ZN(new_n4464_));
  XOR2_X1    g04400(.A1(new_n4460_), .A2(new_n4302_), .Z(new_n4465_));
  NAND2_X1   g04401(.A1(new_n4465_), .A2(new_n4280_), .ZN(new_n4466_));
  OAI21_X1   g04402(.A1(new_n4280_), .A2(new_n4464_), .B(new_n4466_), .ZN(new_n4467_));
  INV_X1     g04403(.I(new_n4295_), .ZN(new_n4468_));
  NOR2_X1    g04404(.A1(new_n4285_), .A2(new_n4294_), .ZN(new_n4469_));
  INV_X1     g04405(.I(new_n4469_), .ZN(new_n4470_));
  OAI22_X1   g04406(.A1(new_n3176_), .A2(new_n4470_), .B1(new_n2665_), .B2(new_n4291_), .ZN(new_n4471_));
  NAND2_X1   g04407(.A1(new_n2728_), .A2(new_n4298_), .ZN(new_n4472_));
  AOI21_X1   g04408(.A1(new_n4471_), .A2(new_n4472_), .B(new_n4468_), .ZN(new_n4473_));
  NAND2_X1   g04409(.A1(new_n3273_), .A2(new_n4473_), .ZN(new_n4474_));
  XOR2_X1    g04410(.A1(new_n4474_), .A2(\a[17] ), .Z(new_n4475_));
  INV_X1     g04411(.I(new_n4475_), .ZN(new_n4476_));
  INV_X1     g04412(.I(new_n4454_), .ZN(new_n4477_));
  AOI21_X1   g04413(.A1(new_n4477_), .A2(new_n4453_), .B(new_n4316_), .ZN(new_n4478_));
  XNOR2_X1   g04414(.A1(new_n4321_), .A2(new_n4452_), .ZN(new_n4479_));
  NOR2_X1    g04415(.A1(new_n4479_), .A2(new_n4317_), .ZN(new_n4480_));
  NOR2_X1    g04416(.A1(new_n4480_), .A2(new_n4478_), .ZN(new_n4481_));
  INV_X1     g04417(.I(new_n4481_), .ZN(new_n4482_));
  OAI22_X1   g04418(.A1(new_n2559_), .A2(new_n3769_), .B1(new_n694_), .B2(new_n4097_), .ZN(new_n4483_));
  NAND2_X1   g04419(.A1(new_n2567_), .A2(new_n3776_), .ZN(new_n4484_));
  AOI21_X1   g04420(.A1(new_n4483_), .A2(new_n4484_), .B(new_n4095_), .ZN(new_n4485_));
  NAND2_X1   g04421(.A1(new_n2759_), .A2(new_n4485_), .ZN(new_n4486_));
  XOR2_X1    g04422(.A1(new_n4486_), .A2(\a[20] ), .Z(new_n4487_));
  INV_X1     g04423(.I(new_n4487_), .ZN(new_n4488_));
  OAI21_X1   g04424(.A1(new_n4449_), .A2(new_n4451_), .B(new_n4324_), .ZN(new_n4489_));
  XOR2_X1    g04425(.A1(new_n4329_), .A2(new_n4448_), .Z(new_n4490_));
  OAI21_X1   g04426(.A1(new_n4324_), .A2(new_n4490_), .B(new_n4489_), .ZN(new_n4491_));
  OAI22_X1   g04427(.A1(new_n896_), .A2(new_n3780_), .B1(new_n1180_), .B2(new_n3310_), .ZN(new_n4492_));
  NAND2_X1   g04428(.A1(new_n2504_), .A2(new_n3782_), .ZN(new_n4493_));
  AOI21_X1   g04429(.A1(new_n4493_), .A2(new_n4492_), .B(new_n3302_), .ZN(new_n4494_));
  NAND2_X1   g04430(.A1(new_n3596_), .A2(new_n4494_), .ZN(new_n4495_));
  XOR2_X1    g04431(.A1(new_n4495_), .A2(\a[23] ), .Z(new_n4496_));
  INV_X1     g04432(.I(new_n4496_), .ZN(new_n4497_));
  XOR2_X1    g04433(.A1(new_n4444_), .A2(new_n4439_), .Z(new_n4498_));
  NAND2_X1   g04434(.A1(new_n4498_), .A2(new_n4336_), .ZN(new_n4499_));
  INV_X1     g04435(.I(new_n4446_), .ZN(new_n4500_));
  NAND2_X1   g04436(.A1(new_n4500_), .A2(new_n4445_), .ZN(new_n4501_));
  NAND2_X1   g04437(.A1(new_n4501_), .A2(new_n4335_), .ZN(new_n4502_));
  NAND2_X1   g04438(.A1(new_n4502_), .A2(new_n4499_), .ZN(new_n4503_));
  OAI22_X1   g04439(.A1(new_n1008_), .A2(new_n3780_), .B1(new_n1121_), .B2(new_n3310_), .ZN(new_n4504_));
  NAND2_X1   g04440(.A1(new_n1181_), .A2(new_n3782_), .ZN(new_n4505_));
  AOI21_X1   g04441(.A1(new_n4504_), .A2(new_n4505_), .B(new_n3302_), .ZN(new_n4506_));
  NAND2_X1   g04442(.A1(new_n3562_), .A2(new_n4506_), .ZN(new_n4507_));
  XOR2_X1    g04443(.A1(new_n4507_), .A2(\a[23] ), .Z(new_n4508_));
  INV_X1     g04444(.I(new_n4508_), .ZN(new_n4509_));
  INV_X1     g04445(.I(new_n4438_), .ZN(new_n4510_));
  AOI21_X1   g04446(.A1(new_n4510_), .A2(new_n4437_), .B(new_n4341_), .ZN(new_n4511_));
  XNOR2_X1   g04447(.A1(new_n4346_), .A2(new_n4436_), .ZN(new_n4512_));
  NOR2_X1    g04448(.A1(new_n4512_), .A2(new_n4342_), .ZN(new_n4513_));
  NOR2_X1    g04449(.A1(new_n4513_), .A2(new_n4511_), .ZN(new_n4514_));
  OAI22_X1   g04450(.A1(new_n2367_), .A2(new_n3268_), .B1(new_n2451_), .B2(new_n3318_), .ZN(new_n4515_));
  NAND2_X1   g04451(.A1(new_n2412_), .A2(new_n3323_), .ZN(new_n4516_));
  AOI21_X1   g04452(.A1(new_n4515_), .A2(new_n4516_), .B(new_n3260_), .ZN(new_n4517_));
  NAND2_X1   g04453(.A1(new_n3403_), .A2(new_n4517_), .ZN(new_n4518_));
  XOR2_X1    g04454(.A1(new_n4518_), .A2(new_n72_), .Z(new_n4519_));
  INV_X1     g04455(.I(new_n4519_), .ZN(new_n4520_));
  XOR2_X1    g04456(.A1(new_n4356_), .A2(new_n4432_), .Z(new_n4521_));
  NOR2_X1    g04457(.A1(new_n4351_), .A2(new_n4521_), .ZN(new_n4522_));
  INV_X1     g04458(.I(new_n4435_), .ZN(new_n4523_));
  NAND2_X1   g04459(.A1(new_n4523_), .A2(new_n4434_), .ZN(new_n4524_));
  AOI21_X1   g04460(.A1(new_n4351_), .A2(new_n4524_), .B(new_n4522_), .ZN(new_n4525_));
  OAI22_X1   g04461(.A1(new_n1409_), .A2(new_n3175_), .B1(new_n2351_), .B2(new_n2747_), .ZN(new_n4526_));
  NAND2_X1   g04462(.A1(new_n2359_), .A2(new_n3275_), .ZN(new_n4527_));
  AOI21_X1   g04463(.A1(new_n4526_), .A2(new_n4527_), .B(new_n2737_), .ZN(new_n4528_));
  NAND2_X1   g04464(.A1(new_n3904_), .A2(new_n4528_), .ZN(new_n4529_));
  XOR2_X1    g04465(.A1(new_n4529_), .A2(\a[29] ), .Z(new_n4530_));
  INV_X1     g04466(.I(new_n4530_), .ZN(new_n4531_));
  OAI22_X1   g04467(.A1(new_n2251_), .A2(new_n2747_), .B1(new_n2351_), .B2(new_n3175_), .ZN(new_n4532_));
  NAND2_X1   g04468(.A1(new_n2310_), .A2(new_n3275_), .ZN(new_n4533_));
  AOI21_X1   g04469(.A1(new_n4533_), .A2(new_n4532_), .B(new_n2737_), .ZN(new_n4534_));
  NAND2_X1   g04470(.A1(new_n3914_), .A2(new_n4534_), .ZN(new_n4535_));
  XOR2_X1    g04471(.A1(new_n4535_), .A2(\a[29] ), .Z(new_n4536_));
  AOI21_X1   g04472(.A1(new_n4390_), .A2(new_n4392_), .B(new_n4369_), .ZN(new_n4537_));
  XOR2_X1    g04473(.A1(new_n4389_), .A2(new_n3959_), .Z(new_n4538_));
  NOR2_X1    g04474(.A1(new_n4370_), .A2(new_n4538_), .ZN(new_n4539_));
  NOR2_X1    g04475(.A1(new_n4539_), .A2(new_n4537_), .ZN(new_n4540_));
  AOI22_X1   g04476(.A1(new_n2072_), .A2(new_n1613_), .B1(new_n2075_), .B2(new_n2074_), .ZN(new_n4541_));
  XOR2_X1    g04477(.A1(new_n2102_), .A2(new_n2107_), .Z(new_n4542_));
  NAND2_X1   g04478(.A1(new_n4541_), .A2(new_n4542_), .ZN(new_n4543_));
  NOR2_X1    g04479(.A1(new_n2104_), .A2(new_n2108_), .ZN(new_n4544_));
  OAI21_X1   g04480(.A1(new_n4541_), .A2(new_n4544_), .B(new_n4543_), .ZN(new_n4545_));
  NOR2_X1    g04481(.A1(new_n2071_), .A2(new_n2767_), .ZN(new_n4546_));
  NOR2_X1    g04482(.A1(new_n2103_), .A2(new_n2772_), .ZN(new_n4547_));
  NOR2_X1    g04483(.A1(new_n1678_), .A2(new_n2771_), .ZN(new_n4548_));
  NOR4_X1    g04484(.A1(new_n4547_), .A2(new_n2763_), .A3(new_n4546_), .A4(new_n4548_), .ZN(new_n4549_));
  NAND2_X1   g04485(.A1(new_n4545_), .A2(new_n4549_), .ZN(new_n4550_));
  NOR3_X1    g04486(.A1(new_n4019_), .A2(new_n2543_), .A3(new_n1822_), .ZN(new_n4551_));
  NAND2_X1   g04487(.A1(new_n765_), .A2(new_n1770_), .ZN(new_n4552_));
  NAND2_X1   g04488(.A1(new_n1356_), .A2(new_n3101_), .ZN(new_n4553_));
  NOR2_X1    g04489(.A1(new_n604_), .A2(new_n192_), .ZN(new_n4554_));
  NOR2_X1    g04490(.A1(new_n262_), .A2(new_n475_), .ZN(new_n4555_));
  NAND4_X1   g04491(.A1(new_n1510_), .A2(new_n4554_), .A3(new_n4555_), .A4(new_n606_), .ZN(new_n4556_));
  NOR4_X1    g04492(.A1(new_n3949_), .A2(new_n4552_), .A3(new_n4553_), .A4(new_n4556_), .ZN(new_n4557_));
  NAND2_X1   g04493(.A1(new_n4551_), .A2(new_n4557_), .ZN(new_n4558_));
  INV_X1     g04494(.I(new_n4558_), .ZN(new_n4559_));
  NAND4_X1   g04495(.A1(new_n1628_), .A2(new_n2375_), .A3(new_n1590_), .A4(new_n432_), .ZN(new_n4560_));
  NOR2_X1    g04496(.A1(new_n2023_), .A2(new_n1988_), .ZN(new_n4561_));
  NAND3_X1   g04497(.A1(new_n3219_), .A2(new_n4560_), .A3(new_n4561_), .ZN(new_n4562_));
  NOR3_X1    g04498(.A1(new_n365_), .A2(new_n294_), .A3(new_n560_), .ZN(new_n4563_));
  NAND4_X1   g04499(.A1(new_n775_), .A2(new_n4563_), .A3(new_n1921_), .A4(new_n1853_), .ZN(new_n4564_));
  NAND2_X1   g04500(.A1(new_n845_), .A2(new_n2795_), .ZN(new_n4565_));
  NOR4_X1    g04501(.A1(new_n4562_), .A2(new_n3485_), .A3(new_n4564_), .A4(new_n4565_), .ZN(new_n4566_));
  NAND4_X1   g04502(.A1(new_n4559_), .A2(new_n1957_), .A3(new_n3196_), .A4(new_n4566_), .ZN(new_n4567_));
  NOR2_X1    g04503(.A1(new_n4567_), .A2(new_n1280_), .ZN(new_n4568_));
  NOR2_X1    g04504(.A1(new_n4568_), .A2(new_n4387_), .ZN(new_n4569_));
  NAND2_X1   g04505(.A1(new_n4568_), .A2(new_n4387_), .ZN(new_n4570_));
  OAI21_X1   g04506(.A1(new_n4550_), .A2(new_n4569_), .B(new_n4570_), .ZN(new_n4571_));
  NAND2_X1   g04507(.A1(new_n1842_), .A2(new_n1823_), .ZN(new_n4572_));
  INV_X1     g04508(.I(new_n4572_), .ZN(new_n4573_));
  INV_X1     g04509(.I(new_n894_), .ZN(new_n4574_));
  NOR4_X1    g04510(.A1(new_n710_), .A2(new_n1197_), .A3(new_n1045_), .A4(new_n1431_), .ZN(new_n4575_));
  NOR3_X1    g04511(.A1(new_n121_), .A2(new_n1154_), .A3(new_n2811_), .ZN(new_n4576_));
  NAND2_X1   g04512(.A1(new_n2802_), .A2(new_n2799_), .ZN(new_n4577_));
  NOR2_X1    g04513(.A1(new_n398_), .A2(new_n468_), .ZN(new_n4578_));
  NAND4_X1   g04514(.A1(new_n1165_), .A2(new_n938_), .A3(new_n3671_), .A4(new_n4578_), .ZN(new_n4579_));
  NOR4_X1    g04515(.A1(new_n495_), .A2(new_n654_), .A3(new_n698_), .A4(new_n930_), .ZN(new_n4580_));
  NOR4_X1    g04516(.A1(new_n4577_), .A2(new_n500_), .A3(new_n4579_), .A4(new_n4580_), .ZN(new_n4581_));
  NAND4_X1   g04517(.A1(new_n4581_), .A2(new_n3486_), .A3(new_n4575_), .A4(new_n4576_), .ZN(new_n4582_));
  NOR2_X1    g04518(.A1(new_n4582_), .A2(new_n4574_), .ZN(new_n4583_));
  AOI21_X1   g04519(.A1(new_n4583_), .A2(new_n4573_), .B(new_n4387_), .ZN(new_n4584_));
  INV_X1     g04520(.I(new_n4584_), .ZN(new_n4585_));
  NAND2_X1   g04521(.A1(new_n4571_), .A2(new_n4585_), .ZN(new_n4586_));
  NAND2_X1   g04522(.A1(new_n4583_), .A2(new_n4573_), .ZN(new_n4587_));
  NOR2_X1    g04523(.A1(new_n4587_), .A2(\a[2] ), .ZN(new_n4588_));
  INV_X1     g04524(.I(new_n4588_), .ZN(new_n4589_));
  NAND2_X1   g04525(.A1(new_n4586_), .A2(new_n4589_), .ZN(new_n4590_));
  NOR3_X1    g04526(.A1(new_n1595_), .A2(new_n137_), .A3(new_n211_), .ZN(new_n4591_));
  NAND4_X1   g04527(.A1(new_n4591_), .A2(new_n1831_), .A3(new_n922_), .A4(new_n643_), .ZN(new_n4592_));
  NAND2_X1   g04528(.A1(new_n3087_), .A2(new_n2795_), .ZN(new_n4593_));
  NOR4_X1    g04529(.A1(new_n4592_), .A2(new_n2391_), .A3(new_n3512_), .A4(new_n4593_), .ZN(new_n4594_));
  NOR3_X1    g04530(.A1(new_n1787_), .A2(new_n640_), .A3(new_n841_), .ZN(new_n4595_));
  INV_X1     g04531(.I(new_n4595_), .ZN(new_n4596_));
  NAND2_X1   g04532(.A1(new_n2527_), .A2(new_n285_), .ZN(new_n4597_));
  NOR4_X1    g04533(.A1(new_n4596_), .A2(new_n415_), .A3(new_n4597_), .A4(new_n3127_), .ZN(new_n4598_));
  NAND3_X1   g04534(.A1(new_n120_), .A2(new_n233_), .A3(new_n856_), .ZN(new_n4599_));
  NOR4_X1    g04535(.A1(new_n2543_), .A2(new_n3864_), .A3(new_n4020_), .A4(new_n4599_), .ZN(new_n4600_));
  NAND4_X1   g04536(.A1(new_n4600_), .A2(new_n380_), .A3(new_n4594_), .A4(new_n4598_), .ZN(new_n4601_));
  NAND2_X1   g04537(.A1(new_n2141_), .A2(new_n1567_), .ZN(new_n4602_));
  NOR2_X1    g04538(.A1(new_n4602_), .A2(new_n4601_), .ZN(new_n4603_));
  NOR2_X1    g04539(.A1(new_n4603_), .A2(new_n4387_), .ZN(new_n4604_));
  INV_X1     g04540(.I(new_n4604_), .ZN(new_n4605_));
  NAND2_X1   g04541(.A1(new_n4590_), .A2(new_n4605_), .ZN(new_n4606_));
  NAND2_X1   g04542(.A1(new_n4603_), .A2(new_n4387_), .ZN(new_n4607_));
  NAND2_X1   g04543(.A1(new_n4606_), .A2(new_n4607_), .ZN(new_n4608_));
  XNOR2_X1   g04544(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n4609_));
  INV_X1     g04545(.I(new_n4609_), .ZN(new_n4610_));
  NOR2_X1    g04546(.A1(new_n4388_), .A2(new_n4385_), .ZN(new_n4611_));
  NOR2_X1    g04547(.A1(new_n4384_), .A2(new_n4611_), .ZN(new_n4612_));
  AOI21_X1   g04548(.A1(new_n4384_), .A2(new_n4610_), .B(new_n4612_), .ZN(new_n4613_));
  INV_X1     g04549(.I(new_n4613_), .ZN(new_n4614_));
  NAND2_X1   g04550(.A1(new_n2201_), .A2(new_n2204_), .ZN(new_n4615_));
  XOR2_X1    g04551(.A1(new_n1503_), .A2(new_n2198_), .Z(new_n4616_));
  NAND2_X1   g04552(.A1(new_n4615_), .A2(new_n4616_), .ZN(new_n4617_));
  OR2_X2     g04553(.A1(new_n2207_), .A2(new_n2205_), .Z(new_n4618_));
  NAND3_X1   g04554(.A1(new_n2201_), .A2(new_n2204_), .A3(new_n4618_), .ZN(new_n4619_));
  NAND2_X1   g04555(.A1(new_n4617_), .A2(new_n4619_), .ZN(new_n4620_));
  NOR2_X1    g04556(.A1(new_n1503_), .A2(new_n2772_), .ZN(new_n4621_));
  NOR2_X1    g04557(.A1(new_n2198_), .A2(new_n2767_), .ZN(new_n4622_));
  NOR2_X1    g04558(.A1(new_n2158_), .A2(new_n2771_), .ZN(new_n4623_));
  NOR4_X1    g04559(.A1(new_n4623_), .A2(new_n4621_), .A3(new_n2763_), .A4(new_n4622_), .ZN(new_n4624_));
  NAND2_X1   g04560(.A1(new_n4620_), .A2(new_n4624_), .ZN(new_n4625_));
  NAND2_X1   g04561(.A1(new_n4625_), .A2(new_n4614_), .ZN(new_n4626_));
  NAND2_X1   g04562(.A1(new_n4608_), .A2(new_n4626_), .ZN(new_n4627_));
  NOR2_X1    g04563(.A1(new_n4625_), .A2(new_n4614_), .ZN(new_n4628_));
  INV_X1     g04564(.I(new_n4628_), .ZN(new_n4629_));
  NAND2_X1   g04565(.A1(new_n4627_), .A2(new_n4629_), .ZN(new_n4630_));
  INV_X1     g04566(.I(new_n4630_), .ZN(new_n4631_));
  NAND2_X1   g04567(.A1(new_n4631_), .A2(new_n4540_), .ZN(new_n4632_));
  INV_X1     g04568(.I(new_n4632_), .ZN(new_n4633_));
  NOR2_X1    g04569(.A1(new_n4631_), .A2(new_n4540_), .ZN(new_n4634_));
  INV_X1     g04570(.I(new_n4634_), .ZN(new_n4635_));
  OAI21_X1   g04571(.A1(new_n4536_), .A2(new_n4633_), .B(new_n4635_), .ZN(new_n4636_));
  INV_X1     g04572(.I(new_n4412_), .ZN(new_n4637_));
  NAND2_X1   g04573(.A1(new_n4637_), .A2(new_n4410_), .ZN(new_n4638_));
  XNOR2_X1   g04574(.A1(new_n3959_), .A2(new_n4408_), .ZN(new_n4639_));
  NOR2_X1    g04575(.A1(new_n4393_), .A2(new_n4639_), .ZN(new_n4640_));
  AOI21_X1   g04576(.A1(new_n4393_), .A2(new_n4638_), .B(new_n4640_), .ZN(new_n4641_));
  NOR3_X1    g04577(.A1(new_n2206_), .A2(new_n1547_), .A3(new_n2207_), .ZN(new_n4642_));
  INV_X1     g04578(.I(new_n4642_), .ZN(new_n4643_));
  OAI21_X1   g04579(.A1(new_n2206_), .A2(new_n2207_), .B(new_n1547_), .ZN(new_n4644_));
  NAND2_X1   g04580(.A1(new_n4643_), .A2(new_n4644_), .ZN(new_n4645_));
  NAND3_X1   g04581(.A1(new_n4645_), .A2(new_n2255_), .A3(new_n4358_), .ZN(new_n4646_));
  INV_X1     g04582(.I(new_n4644_), .ZN(new_n4647_));
  OAI21_X1   g04583(.A1(new_n4647_), .A2(new_n4642_), .B(new_n4358_), .ZN(new_n4648_));
  NAND2_X1   g04584(.A1(new_n4648_), .A2(new_n2251_), .ZN(new_n4649_));
  NAND2_X1   g04585(.A1(new_n4649_), .A2(new_n4646_), .ZN(new_n4650_));
  NOR2_X1    g04586(.A1(new_n1503_), .A2(new_n2771_), .ZN(new_n4651_));
  NOR2_X1    g04587(.A1(new_n2251_), .A2(new_n2772_), .ZN(new_n4652_));
  NOR2_X1    g04588(.A1(new_n4365_), .A2(new_n2767_), .ZN(new_n4653_));
  NOR4_X1    g04589(.A1(new_n4652_), .A2(new_n2763_), .A3(new_n4651_), .A4(new_n4653_), .ZN(new_n4654_));
  AND2_X2    g04590(.A1(new_n4650_), .A2(new_n4654_), .Z(new_n4655_));
  INV_X1     g04591(.I(new_n4655_), .ZN(new_n4656_));
  NAND2_X1   g04592(.A1(new_n4641_), .A2(new_n4656_), .ZN(new_n4657_));
  NOR2_X1    g04593(.A1(new_n4641_), .A2(new_n4656_), .ZN(new_n4658_));
  AOI21_X1   g04594(.A1(new_n4636_), .A2(new_n4657_), .B(new_n4658_), .ZN(new_n4659_));
  AOI21_X1   g04595(.A1(new_n4429_), .A2(new_n4431_), .B(new_n4413_), .ZN(new_n4660_));
  XOR2_X1    g04596(.A1(new_n4424_), .A2(new_n4428_), .Z(new_n4661_));
  AOI21_X1   g04597(.A1(new_n4661_), .A2(new_n4413_), .B(new_n4660_), .ZN(new_n4662_));
  NAND2_X1   g04598(.A1(new_n4659_), .A2(new_n4662_), .ZN(new_n4663_));
  NAND2_X1   g04599(.A1(new_n4663_), .A2(new_n4531_), .ZN(new_n4664_));
  OR2_X2     g04600(.A1(new_n4659_), .A2(new_n4662_), .Z(new_n4665_));
  NAND2_X1   g04601(.A1(new_n4664_), .A2(new_n4665_), .ZN(new_n4666_));
  NOR2_X1    g04602(.A1(new_n4525_), .A2(new_n4666_), .ZN(new_n4667_));
  NOR2_X1    g04603(.A1(new_n4520_), .A2(new_n4667_), .ZN(new_n4668_));
  AND2_X2    g04604(.A1(new_n4525_), .A2(new_n4666_), .Z(new_n4669_));
  NOR2_X1    g04605(.A1(new_n4668_), .A2(new_n4669_), .ZN(new_n4670_));
  NAND2_X1   g04606(.A1(new_n4514_), .A2(new_n4670_), .ZN(new_n4671_));
  NOR2_X1    g04607(.A1(new_n4514_), .A2(new_n4670_), .ZN(new_n4672_));
  AOI21_X1   g04608(.A1(new_n4509_), .A2(new_n4671_), .B(new_n4672_), .ZN(new_n4673_));
  NAND2_X1   g04609(.A1(new_n4503_), .A2(new_n4673_), .ZN(new_n4674_));
  NOR2_X1    g04610(.A1(new_n4503_), .A2(new_n4673_), .ZN(new_n4675_));
  AOI21_X1   g04611(.A1(new_n4497_), .A2(new_n4674_), .B(new_n4675_), .ZN(new_n4676_));
  INV_X1     g04612(.I(new_n4676_), .ZN(new_n4677_));
  NOR2_X1    g04613(.A1(new_n4491_), .A2(new_n4677_), .ZN(new_n4678_));
  INV_X1     g04614(.I(new_n4678_), .ZN(new_n4679_));
  NAND2_X1   g04615(.A1(new_n4491_), .A2(new_n4677_), .ZN(new_n4680_));
  INV_X1     g04616(.I(new_n4680_), .ZN(new_n4681_));
  AOI21_X1   g04617(.A1(new_n4488_), .A2(new_n4679_), .B(new_n4681_), .ZN(new_n4682_));
  INV_X1     g04618(.I(new_n4682_), .ZN(new_n4683_));
  NOR2_X1    g04619(.A1(new_n4482_), .A2(new_n4683_), .ZN(new_n4684_));
  INV_X1     g04620(.I(new_n4684_), .ZN(new_n4685_));
  NOR2_X1    g04621(.A1(new_n4481_), .A2(new_n4682_), .ZN(new_n4686_));
  AOI21_X1   g04622(.A1(new_n4685_), .A2(new_n4476_), .B(new_n4686_), .ZN(new_n4687_));
  INV_X1     g04623(.I(new_n4687_), .ZN(new_n4688_));
  XOR2_X1    g04624(.A1(new_n4310_), .A2(new_n4456_), .Z(new_n4689_));
  OAI21_X1   g04625(.A1(new_n4457_), .A2(new_n4458_), .B(new_n4307_), .ZN(new_n4690_));
  OAI21_X1   g04626(.A1(new_n4307_), .A2(new_n4689_), .B(new_n4690_), .ZN(new_n4691_));
  OAI22_X1   g04627(.A1(new_n3176_), .A2(new_n4297_), .B1(new_n3142_), .B2(new_n4470_), .ZN(new_n4692_));
  NAND2_X1   g04628(.A1(new_n2728_), .A2(new_n4292_), .ZN(new_n4693_));
  AOI21_X1   g04629(.A1(new_n4692_), .A2(new_n4693_), .B(new_n4468_), .ZN(new_n4694_));
  NAND2_X1   g04630(.A1(new_n3174_), .A2(new_n4694_), .ZN(new_n4695_));
  XOR2_X1    g04631(.A1(new_n4695_), .A2(\a[17] ), .Z(new_n4696_));
  NAND2_X1   g04632(.A1(new_n4691_), .A2(new_n4696_), .ZN(new_n4697_));
  NOR2_X1    g04633(.A1(new_n4691_), .A2(new_n4696_), .ZN(new_n4698_));
  AOI21_X1   g04634(.A1(new_n4688_), .A2(new_n4697_), .B(new_n4698_), .ZN(new_n4699_));
  NOR2_X1    g04635(.A1(new_n4467_), .A2(new_n4699_), .ZN(new_n4700_));
  INV_X1     g04636(.I(\a[9] ), .ZN(new_n4701_));
  NOR2_X1    g04637(.A1(new_n4701_), .A2(\a[8] ), .ZN(new_n4702_));
  NOR2_X1    g04638(.A1(new_n4009_), .A2(\a[9] ), .ZN(new_n4703_));
  NOR2_X1    g04639(.A1(new_n4702_), .A2(new_n4703_), .ZN(new_n4704_));
  XNOR2_X1   g04640(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n4705_));
  NOR2_X1    g04641(.A1(new_n4704_), .A2(new_n4705_), .ZN(new_n4706_));
  INV_X1     g04642(.I(new_n4706_), .ZN(new_n4707_));
  INV_X1     g04643(.I(new_n4704_), .ZN(new_n4708_));
  NOR2_X1    g04644(.A1(new_n4708_), .A2(new_n4705_), .ZN(new_n4709_));
  INV_X1     g04645(.I(new_n4709_), .ZN(new_n4710_));
  INV_X1     g04646(.I(\a[10] ), .ZN(new_n4711_));
  NOR2_X1    g04647(.A1(new_n4711_), .A2(\a[8] ), .ZN(new_n4712_));
  NOR2_X1    g04648(.A1(new_n4009_), .A2(\a[10] ), .ZN(new_n4713_));
  OR2_X2     g04649(.A1(new_n4712_), .A2(new_n4713_), .Z(new_n4714_));
  XNOR2_X1   g04650(.A1(\a[8] ), .A2(\a[11] ), .ZN(new_n4715_));
  OAI21_X1   g04651(.A1(new_n4708_), .A2(new_n4714_), .B(new_n4715_), .ZN(new_n4716_));
  OAI22_X1   g04652(.A1(new_n2559_), .A2(new_n4710_), .B1(new_n896_), .B2(new_n4716_), .ZN(new_n4717_));
  NOR3_X1    g04653(.A1(new_n4711_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n4718_));
  AOI21_X1   g04654(.A1(\a[9] ), .A2(new_n4713_), .B(new_n4718_), .ZN(new_n4719_));
  INV_X1     g04655(.I(new_n4719_), .ZN(new_n4720_));
  NAND2_X1   g04656(.A1(new_n814_), .A2(new_n4720_), .ZN(new_n4721_));
  AOI21_X1   g04657(.A1(new_n4717_), .A2(new_n4721_), .B(new_n4707_), .ZN(new_n4722_));
  NAND2_X1   g04658(.A1(new_n3624_), .A2(new_n4722_), .ZN(new_n4723_));
  XOR2_X1    g04659(.A1(new_n4723_), .A2(\a[11] ), .Z(new_n4724_));
  OAI22_X1   g04660(.A1(new_n2367_), .A2(new_n4297_), .B1(new_n2408_), .B2(new_n4470_), .ZN(new_n4725_));
  NAND2_X1   g04661(.A1(new_n1334_), .A2(new_n4292_), .ZN(new_n4726_));
  AOI21_X1   g04662(.A1(new_n4725_), .A2(new_n4726_), .B(new_n4468_), .ZN(new_n4727_));
  AND3_X2    g04663(.A1(new_n3708_), .A2(new_n3372_), .A3(new_n4727_), .Z(new_n4728_));
  AOI21_X1   g04664(.A1(new_n3708_), .A2(new_n4727_), .B(new_n3372_), .ZN(new_n4729_));
  NOR2_X1    g04665(.A1(new_n4728_), .A2(new_n4729_), .ZN(new_n4730_));
  INV_X1     g04666(.I(new_n4730_), .ZN(new_n4731_));
  OAI22_X1   g04667(.A1(new_n4365_), .A2(new_n3318_), .B1(new_n2198_), .B2(new_n3268_), .ZN(new_n4732_));
  NAND2_X1   g04668(.A1(new_n1504_), .A2(new_n3323_), .ZN(new_n4733_));
  AOI21_X1   g04669(.A1(new_n4732_), .A2(new_n4733_), .B(new_n3260_), .ZN(new_n4734_));
  NAND2_X1   g04670(.A1(new_n4363_), .A2(new_n4734_), .ZN(new_n4735_));
  XOR2_X1    g04671(.A1(new_n4735_), .A2(\a[26] ), .Z(new_n4736_));
  INV_X1     g04672(.I(new_n4736_), .ZN(new_n4737_));
  OAI21_X1   g04673(.A1(new_n1941_), .A2(new_n2000_), .B(new_n1763_), .ZN(new_n4738_));
  NOR4_X1    g04674(.A1(new_n505_), .A2(new_n90_), .A3(new_n119_), .A4(new_n1035_), .ZN(new_n4739_));
  NOR4_X1    g04675(.A1(new_n4739_), .A2(new_n268_), .A3(new_n1640_), .A4(new_n796_), .ZN(new_n4740_));
  NAND2_X1   g04676(.A1(new_n2055_), .A2(new_n677_), .ZN(new_n4741_));
  NOR4_X1    g04677(.A1(new_n4741_), .A2(new_n1914_), .A3(new_n1591_), .A4(new_n1183_), .ZN(new_n4742_));
  NOR4_X1    g04678(.A1(new_n1373_), .A2(new_n1771_), .A3(new_n1772_), .A4(new_n1769_), .ZN(new_n4743_));
  NAND4_X1   g04679(.A1(new_n4743_), .A2(new_n4740_), .A3(new_n4742_), .A4(new_n1776_), .ZN(new_n4744_));
  NOR4_X1    g04680(.A1(new_n4744_), .A2(new_n1900_), .A3(new_n1786_), .A4(new_n1799_), .ZN(new_n4745_));
  NOR2_X1    g04681(.A1(new_n1939_), .A2(new_n1882_), .ZN(new_n4746_));
  NOR2_X1    g04682(.A1(new_n1862_), .A2(new_n1729_), .ZN(new_n4747_));
  OAI21_X1   g04683(.A1(new_n4747_), .A2(new_n4746_), .B(new_n4745_), .ZN(new_n4748_));
  NOR2_X1    g04684(.A1(new_n548_), .A2(new_n304_), .ZN(new_n4749_));
  NOR4_X1    g04685(.A1(new_n4749_), .A2(new_n247_), .A3(new_n260_), .A4(new_n468_), .ZN(new_n4750_));
  NAND4_X1   g04686(.A1(new_n2938_), .A2(new_n4750_), .A3(new_n1945_), .A4(new_n1946_), .ZN(new_n4751_));
  NOR2_X1    g04687(.A1(new_n638_), .A2(new_n1073_), .ZN(new_n4752_));
  NOR2_X1    g04688(.A1(new_n956_), .A2(new_n4752_), .ZN(new_n4753_));
  NOR2_X1    g04689(.A1(new_n305_), .A2(new_n1035_), .ZN(new_n4754_));
  NOR4_X1    g04690(.A1(new_n995_), .A2(new_n4754_), .A3(new_n163_), .A4(new_n1962_), .ZN(new_n4755_));
  NAND4_X1   g04691(.A1(new_n4755_), .A2(new_n1244_), .A3(new_n4753_), .A4(new_n1326_), .ZN(new_n4756_));
  NOR4_X1    g04692(.A1(new_n4751_), .A2(new_n4756_), .A3(new_n1951_), .A4(new_n1956_), .ZN(new_n4757_));
  INV_X1     g04693(.I(new_n500_), .ZN(new_n4758_));
  NOR2_X1    g04694(.A1(new_n565_), .A2(new_n656_), .ZN(new_n4759_));
  NOR2_X1    g04695(.A1(new_n936_), .A2(new_n135_), .ZN(new_n4760_));
  NAND4_X1   g04696(.A1(new_n1921_), .A2(new_n1491_), .A3(new_n672_), .A4(new_n432_), .ZN(new_n4761_));
  NAND4_X1   g04697(.A1(new_n4759_), .A2(new_n4760_), .A3(new_n4758_), .A4(new_n4761_), .ZN(new_n4762_));
  NAND2_X1   g04698(.A1(new_n1977_), .A2(new_n1975_), .ZN(new_n4763_));
  NOR3_X1    g04699(.A1(new_n4763_), .A2(new_n291_), .A3(new_n4762_), .ZN(new_n4764_));
  NOR2_X1    g04700(.A1(new_n1998_), .A2(new_n1983_), .ZN(new_n4765_));
  NAND3_X1   g04701(.A1(new_n4757_), .A2(new_n4765_), .A3(new_n4764_), .ZN(new_n4766_));
  NAND3_X1   g04702(.A1(new_n4766_), .A2(new_n1729_), .A3(new_n1862_), .ZN(new_n4767_));
  NAND3_X1   g04703(.A1(new_n4748_), .A2(new_n1764_), .A3(new_n4767_), .ZN(new_n4768_));
  NAND2_X1   g04704(.A1(new_n4738_), .A2(new_n4768_), .ZN(new_n4769_));
  NAND2_X1   g04705(.A1(new_n1763_), .A2(new_n1729_), .ZN(new_n4770_));
  NAND4_X1   g04706(.A1(new_n1749_), .A2(new_n1882_), .A3(new_n1762_), .A4(new_n1567_), .ZN(new_n4771_));
  NAND2_X1   g04707(.A1(new_n4770_), .A2(new_n4771_), .ZN(new_n4772_));
  NAND3_X1   g04708(.A1(new_n4769_), .A2(new_n1613_), .A3(new_n4772_), .ZN(new_n4773_));
  AOI21_X1   g04709(.A1(new_n4748_), .A2(new_n4767_), .B(new_n1764_), .ZN(new_n4774_));
  NOR3_X1    g04710(.A1(new_n1941_), .A2(new_n1763_), .A3(new_n2000_), .ZN(new_n4775_));
  OAI21_X1   g04711(.A1(new_n4774_), .A2(new_n4775_), .B(new_n4772_), .ZN(new_n4776_));
  NAND2_X1   g04712(.A1(new_n4776_), .A2(new_n1612_), .ZN(new_n4777_));
  NAND2_X1   g04713(.A1(new_n4777_), .A2(new_n4773_), .ZN(new_n4778_));
  NOR2_X1    g04714(.A1(new_n1612_), .A2(new_n2772_), .ZN(new_n4779_));
  NOR2_X1    g04715(.A1(new_n1764_), .A2(new_n2767_), .ZN(new_n4780_));
  NOR2_X1    g04716(.A1(new_n1729_), .A2(new_n2771_), .ZN(new_n4781_));
  NOR4_X1    g04717(.A1(new_n4780_), .A2(new_n4779_), .A3(new_n2763_), .A4(new_n4781_), .ZN(new_n4782_));
  NAND2_X1   g04718(.A1(new_n4778_), .A2(new_n4782_), .ZN(new_n4783_));
  NOR4_X1    g04719(.A1(new_n1669_), .A2(new_n666_), .A3(new_n736_), .A4(new_n1092_), .ZN(new_n4784_));
  NAND4_X1   g04720(.A1(new_n313_), .A2(new_n287_), .A3(new_n707_), .A4(new_n1305_), .ZN(new_n4785_));
  NAND4_X1   g04721(.A1(new_n480_), .A2(new_n481_), .A3(new_n1444_), .A4(new_n182_), .ZN(new_n4786_));
  NAND4_X1   g04722(.A1(new_n4784_), .A2(new_n257_), .A3(new_n4785_), .A4(new_n4786_), .ZN(new_n4787_));
  NOR3_X1    g04723(.A1(new_n3213_), .A2(new_n535_), .A3(new_n654_), .ZN(new_n4788_));
  NOR2_X1    g04724(.A1(new_n2047_), .A2(new_n3991_), .ZN(new_n4789_));
  NOR3_X1    g04725(.A1(new_n330_), .A2(new_n596_), .A3(new_n682_), .ZN(new_n4790_));
  NAND4_X1   g04726(.A1(new_n4788_), .A2(new_n4789_), .A3(new_n2154_), .A4(new_n4790_), .ZN(new_n4791_));
  NOR4_X1    g04727(.A1(new_n2589_), .A2(new_n4787_), .A3(new_n1626_), .A4(new_n4791_), .ZN(new_n4792_));
  NAND3_X1   g04728(.A1(new_n1515_), .A2(new_n978_), .A3(new_n1100_), .ZN(new_n4793_));
  NOR2_X1    g04729(.A1(new_n946_), .A2(new_n172_), .ZN(new_n4794_));
  NAND4_X1   g04730(.A1(new_n4793_), .A2(new_n1446_), .A3(new_n2188_), .A4(new_n4794_), .ZN(new_n4795_));
  NOR2_X1    g04731(.A1(new_n203_), .A2(new_n268_), .ZN(new_n4796_));
  NAND4_X1   g04732(.A1(new_n162_), .A2(new_n545_), .A3(new_n4796_), .A4(new_n1338_), .ZN(new_n4797_));
  NOR4_X1    g04733(.A1(new_n2884_), .A2(new_n262_), .A3(new_n648_), .A4(new_n634_), .ZN(new_n4798_));
  NOR4_X1    g04734(.A1(new_n565_), .A2(new_n2338_), .A3(new_n406_), .A4(new_n345_), .ZN(new_n4799_));
  NAND2_X1   g04735(.A1(new_n4798_), .A2(new_n4799_), .ZN(new_n4800_));
  NOR4_X1    g04736(.A1(new_n4800_), .A2(new_n4024_), .A3(new_n4795_), .A4(new_n4797_), .ZN(new_n4801_));
  NAND3_X1   g04737(.A1(new_n4792_), .A2(new_n3933_), .A3(new_n4801_), .ZN(new_n4802_));
  OR2_X2     g04738(.A1(new_n4783_), .A2(new_n4802_), .Z(new_n4803_));
  NOR3_X1    g04739(.A1(new_n1813_), .A2(new_n1862_), .A3(new_n1729_), .ZN(new_n4804_));
  NOR3_X1    g04740(.A1(new_n1941_), .A2(new_n1882_), .A3(new_n2000_), .ZN(new_n4805_));
  OAI21_X1   g04741(.A1(new_n4805_), .A2(new_n4804_), .B(new_n1764_), .ZN(new_n4806_));
  AOI21_X1   g04742(.A1(new_n4745_), .A2(new_n1939_), .B(new_n1729_), .ZN(new_n4807_));
  AOI21_X1   g04743(.A1(new_n4748_), .A2(new_n4767_), .B(new_n1882_), .ZN(new_n4808_));
  OAI21_X1   g04744(.A1(new_n4808_), .A2(new_n4807_), .B(new_n1763_), .ZN(new_n4809_));
  NAND2_X1   g04745(.A1(new_n4806_), .A2(new_n4809_), .ZN(new_n4810_));
  NOR2_X1    g04746(.A1(new_n1939_), .A2(new_n2771_), .ZN(new_n4811_));
  NOR2_X1    g04747(.A1(new_n1764_), .A2(new_n2772_), .ZN(new_n4812_));
  NOR2_X1    g04748(.A1(new_n1729_), .A2(new_n2767_), .ZN(new_n4813_));
  NOR4_X1    g04749(.A1(new_n4812_), .A2(new_n2763_), .A3(new_n4811_), .A4(new_n4813_), .ZN(new_n4814_));
  NAND2_X1   g04750(.A1(new_n4810_), .A2(new_n4814_), .ZN(new_n4815_));
  NAND2_X1   g04751(.A1(new_n554_), .A2(new_n476_), .ZN(new_n4816_));
  NOR4_X1    g04752(.A1(new_n198_), .A2(new_n837_), .A3(new_n1531_), .A4(new_n817_), .ZN(new_n4817_));
  NOR4_X1    g04753(.A1(new_n2338_), .A2(new_n898_), .A3(new_n556_), .A4(new_n910_), .ZN(new_n4818_));
  NAND4_X1   g04754(.A1(new_n4818_), .A2(new_n913_), .A3(new_n592_), .A4(new_n1419_), .ZN(new_n4819_));
  NOR4_X1    g04755(.A1(new_n4819_), .A2(new_n1415_), .A3(new_n4816_), .A4(new_n4817_), .ZN(new_n4820_));
  NOR4_X1    g04756(.A1(new_n326_), .A2(new_n90_), .A3(new_n312_), .A4(new_n376_), .ZN(new_n4821_));
  NOR4_X1    g04757(.A1(new_n2703_), .A2(new_n2881_), .A3(new_n603_), .A4(new_n4821_), .ZN(new_n4822_));
  NAND2_X1   g04758(.A1(new_n641_), .A2(new_n646_), .ZN(new_n4823_));
  NAND4_X1   g04759(.A1(new_n1804_), .A2(new_n627_), .A3(new_n390_), .A4(new_n409_), .ZN(new_n4824_));
  NOR4_X1    g04760(.A1(new_n4824_), .A2(new_n177_), .A3(new_n687_), .A4(new_n4823_), .ZN(new_n4825_));
  NOR3_X1    g04761(.A1(new_n343_), .A2(new_n944_), .A3(new_n1073_), .ZN(new_n4826_));
  NAND4_X1   g04762(.A1(new_n4826_), .A2(new_n221_), .A3(new_n564_), .A4(new_n1354_), .ZN(new_n4827_));
  NOR4_X1    g04763(.A1(new_n4827_), .A2(new_n1079_), .A3(new_n2381_), .A4(new_n3485_), .ZN(new_n4828_));
  NAND4_X1   g04764(.A1(new_n4820_), .A2(new_n4828_), .A3(new_n4822_), .A4(new_n4825_), .ZN(new_n4829_));
  NOR2_X1    g04765(.A1(new_n2030_), .A2(new_n4829_), .ZN(new_n4830_));
  INV_X1     g04766(.I(new_n4830_), .ZN(new_n4831_));
  NOR2_X1    g04767(.A1(new_n4815_), .A2(new_n4831_), .ZN(new_n4832_));
  NAND4_X1   g04768(.A1(new_n1939_), .A2(new_n4757_), .A3(new_n4764_), .A4(new_n4765_), .ZN(new_n4833_));
  NAND2_X1   g04769(.A1(new_n1862_), .A2(new_n4745_), .ZN(new_n4834_));
  NAND2_X1   g04770(.A1(new_n1813_), .A2(new_n1939_), .ZN(new_n4835_));
  NAND2_X1   g04771(.A1(new_n4835_), .A2(new_n4834_), .ZN(new_n4836_));
  NAND3_X1   g04772(.A1(new_n4836_), .A2(new_n1882_), .A3(new_n4833_), .ZN(new_n4837_));
  NOR2_X1    g04773(.A1(new_n1813_), .A2(new_n1939_), .ZN(new_n4838_));
  NOR2_X1    g04774(.A1(new_n1862_), .A2(new_n4745_), .ZN(new_n4839_));
  OAI21_X1   g04775(.A1(new_n4838_), .A2(new_n4839_), .B(new_n4833_), .ZN(new_n4840_));
  NAND2_X1   g04776(.A1(new_n4840_), .A2(new_n1729_), .ZN(new_n4841_));
  NAND2_X1   g04777(.A1(new_n4841_), .A2(new_n4837_), .ZN(new_n4842_));
  NOR3_X1    g04778(.A1(new_n1730_), .A2(new_n453_), .A3(new_n899_), .ZN(new_n4843_));
  NOR3_X1    g04779(.A1(new_n289_), .A2(new_n582_), .A3(new_n90_), .ZN(new_n4844_));
  NOR4_X1    g04780(.A1(new_n604_), .A2(new_n235_), .A3(new_n242_), .A4(new_n280_), .ZN(new_n4845_));
  INV_X1     g04781(.I(new_n4845_), .ZN(new_n4846_));
  AND3_X2    g04782(.A1(new_n4846_), .A2(new_n4843_), .A3(new_n4844_), .Z(new_n4847_));
  INV_X1     g04783(.I(new_n4847_), .ZN(new_n4848_));
  NOR4_X1    g04784(.A1(new_n1262_), .A2(new_n945_), .A3(new_n326_), .A4(new_n304_), .ZN(new_n4849_));
  NOR4_X1    g04785(.A1(new_n4849_), .A2(new_n310_), .A3(new_n715_), .A4(new_n776_), .ZN(new_n4850_));
  INV_X1     g04786(.I(new_n4850_), .ZN(new_n4851_));
  NOR2_X1    g04787(.A1(new_n2333_), .A2(new_n2331_), .ZN(new_n4852_));
  NOR2_X1    g04788(.A1(new_n415_), .A2(new_n367_), .ZN(new_n4853_));
  NAND4_X1   g04789(.A1(new_n4852_), .A2(new_n723_), .A3(new_n1223_), .A4(new_n4853_), .ZN(new_n4854_));
  NOR4_X1    g04790(.A1(new_n4848_), .A2(new_n1846_), .A3(new_n4851_), .A4(new_n4854_), .ZN(new_n4855_));
  NOR4_X1    g04791(.A1(new_n1048_), .A2(new_n413_), .A3(new_n574_), .A4(new_n594_), .ZN(new_n4856_));
  OR3_X2     g04792(.A1(new_n4856_), .A2(new_n682_), .A3(new_n2930_), .Z(new_n4857_));
  NOR4_X1    g04793(.A1(new_n4857_), .A2(new_n1410_), .A3(new_n2323_), .A4(new_n3855_), .ZN(new_n4858_));
  NOR4_X1    g04794(.A1(new_n212_), .A2(new_n288_), .A3(new_n403_), .A4(new_n902_), .ZN(new_n4859_));
  NOR3_X1    g04795(.A1(new_n1213_), .A2(new_n418_), .A3(new_n732_), .ZN(new_n4860_));
  INV_X1     g04796(.I(new_n4860_), .ZN(new_n4861_));
  NOR4_X1    g04797(.A1(new_n365_), .A2(new_n505_), .A3(new_n172_), .A4(new_n1073_), .ZN(new_n4862_));
  NOR3_X1    g04798(.A1(new_n4861_), .A2(new_n4859_), .A3(new_n4862_), .ZN(new_n4863_));
  NAND2_X1   g04799(.A1(new_n1562_), .A2(new_n2456_), .ZN(new_n4864_));
  NOR2_X1    g04800(.A1(new_n86_), .A2(new_n333_), .ZN(new_n4865_));
  NAND4_X1   g04801(.A1(new_n688_), .A2(new_n875_), .A3(new_n4865_), .A4(new_n1126_), .ZN(new_n4866_));
  NOR4_X1    g04802(.A1(new_n4866_), .A2(new_n4864_), .A3(new_n1323_), .A4(new_n1434_), .ZN(new_n4867_));
  AND3_X2    g04803(.A1(new_n4858_), .A2(new_n4863_), .A3(new_n4867_), .Z(new_n4868_));
  NAND3_X1   g04804(.A1(new_n4868_), .A2(new_n1362_), .A3(new_n4855_), .ZN(new_n4869_));
  INV_X1     g04805(.I(new_n4869_), .ZN(new_n4870_));
  NOR2_X1    g04806(.A1(new_n1939_), .A2(new_n2767_), .ZN(new_n4871_));
  NOR2_X1    g04807(.A1(new_n1729_), .A2(new_n2772_), .ZN(new_n4872_));
  NOR2_X1    g04808(.A1(new_n4745_), .A2(new_n2771_), .ZN(new_n4873_));
  NOR4_X1    g04809(.A1(new_n4871_), .A2(new_n4872_), .A3(new_n4873_), .A4(new_n2763_), .ZN(new_n4874_));
  NAND3_X1   g04810(.A1(new_n4842_), .A2(new_n4870_), .A3(new_n4874_), .ZN(new_n4875_));
  NOR2_X1    g04811(.A1(new_n4766_), .A2(new_n1862_), .ZN(new_n4876_));
  NAND2_X1   g04812(.A1(new_n1999_), .A2(new_n1813_), .ZN(new_n4877_));
  AOI22_X1   g04813(.A1(new_n4877_), .A2(new_n1862_), .B1(new_n4876_), .B2(new_n1813_), .ZN(new_n4878_));
  NOR2_X1    g04814(.A1(new_n1939_), .A2(new_n2772_), .ZN(new_n4879_));
  NOR2_X1    g04815(.A1(new_n4745_), .A2(new_n2767_), .ZN(new_n4880_));
  OAI21_X1   g04816(.A1(new_n1999_), .A2(new_n2771_), .B(new_n2764_), .ZN(new_n4881_));
  NOR4_X1    g04817(.A1(new_n4878_), .A2(new_n4879_), .A3(new_n4880_), .A4(new_n4881_), .ZN(new_n4882_));
  NOR3_X1    g04818(.A1(new_n552_), .A2(new_n264_), .A3(new_n388_), .ZN(new_n4883_));
  NOR4_X1    g04819(.A1(new_n235_), .A2(new_n282_), .A3(new_n381_), .A4(new_n370_), .ZN(new_n4884_));
  NOR3_X1    g04820(.A1(new_n4883_), .A2(new_n1788_), .A3(new_n4884_), .ZN(new_n4885_));
  INV_X1     g04821(.I(new_n722_), .ZN(new_n4886_));
  NOR4_X1    g04822(.A1(new_n717_), .A2(new_n4886_), .A3(new_n2098_), .A4(new_n1053_), .ZN(new_n4887_));
  NOR2_X1    g04823(.A1(new_n584_), .A2(new_n286_), .ZN(new_n4888_));
  NOR4_X1    g04824(.A1(new_n553_), .A2(new_n654_), .A3(new_n428_), .A4(new_n329_), .ZN(new_n4889_));
  NOR2_X1    g04825(.A1(new_n596_), .A2(new_n776_), .ZN(new_n4890_));
  AOI21_X1   g04826(.A1(new_n4888_), .A2(new_n4890_), .B(new_n4889_), .ZN(new_n4891_));
  NOR4_X1    g04827(.A1(new_n687_), .A2(new_n136_), .A3(new_n413_), .A4(new_n474_), .ZN(new_n4892_));
  INV_X1     g04828(.I(new_n2191_), .ZN(new_n4893_));
  NOR4_X1    g04829(.A1(new_n958_), .A2(new_n2480_), .A3(new_n4893_), .A4(new_n1019_), .ZN(new_n4894_));
  NAND2_X1   g04830(.A1(new_n4894_), .A2(new_n4892_), .ZN(new_n4895_));
  INV_X1     g04831(.I(new_n4895_), .ZN(new_n4896_));
  AND3_X2    g04832(.A1(new_n4896_), .A2(new_n4887_), .A3(new_n4891_), .Z(new_n4897_));
  NOR2_X1    g04833(.A1(new_n3346_), .A2(new_n2889_), .ZN(new_n4898_));
  NAND4_X1   g04834(.A1(new_n4898_), .A2(new_n2116_), .A3(new_n4885_), .A4(new_n4897_), .ZN(new_n4899_));
  INV_X1     g04835(.I(new_n4899_), .ZN(new_n4900_));
  OR2_X2     g04836(.A1(new_n4882_), .A2(new_n4900_), .Z(new_n4901_));
  NAND2_X1   g04837(.A1(new_n4842_), .A2(new_n4874_), .ZN(new_n4902_));
  NAND2_X1   g04838(.A1(new_n4902_), .A2(new_n4869_), .ZN(new_n4903_));
  NAND2_X1   g04839(.A1(new_n4903_), .A2(new_n4901_), .ZN(new_n4904_));
  AOI22_X1   g04840(.A1(new_n4904_), .A2(new_n4875_), .B1(new_n4815_), .B2(new_n4831_), .ZN(new_n4905_));
  NOR2_X1    g04841(.A1(new_n4905_), .A2(new_n4832_), .ZN(new_n4906_));
  INV_X1     g04842(.I(new_n4906_), .ZN(new_n4907_));
  NAND2_X1   g04843(.A1(new_n4783_), .A2(new_n4802_), .ZN(new_n4908_));
  NAND2_X1   g04844(.A1(new_n4907_), .A2(new_n4908_), .ZN(new_n4909_));
  NAND2_X1   g04845(.A1(new_n4909_), .A2(new_n4803_), .ZN(new_n4910_));
  NAND2_X1   g04846(.A1(new_n4748_), .A2(new_n4767_), .ZN(new_n4911_));
  OAI21_X1   g04847(.A1(new_n4911_), .A2(new_n1612_), .B(new_n1764_), .ZN(new_n4912_));
  NAND2_X1   g04848(.A1(new_n4912_), .A2(new_n1882_), .ZN(new_n4913_));
  XOR2_X1    g04849(.A1(new_n1678_), .A2(new_n1612_), .Z(new_n4914_));
  NAND3_X1   g04850(.A1(new_n4913_), .A2(new_n2004_), .A3(new_n4914_), .ZN(new_n4915_));
  XOR2_X1    g04851(.A1(new_n1678_), .A2(new_n1612_), .Z(new_n4916_));
  OAI21_X1   g04852(.A1(new_n2006_), .A2(new_n4916_), .B(new_n4915_), .ZN(new_n4917_));
  NOR2_X1    g04853(.A1(new_n1612_), .A2(new_n2767_), .ZN(new_n4918_));
  NOR2_X1    g04854(.A1(new_n1678_), .A2(new_n2772_), .ZN(new_n4919_));
  NOR2_X1    g04855(.A1(new_n1764_), .A2(new_n2771_), .ZN(new_n4920_));
  NOR4_X1    g04856(.A1(new_n4919_), .A2(new_n2763_), .A3(new_n4920_), .A4(new_n4918_), .ZN(new_n4921_));
  NAND2_X1   g04857(.A1(new_n4917_), .A2(new_n4921_), .ZN(new_n4922_));
  INV_X1     g04858(.I(new_n878_), .ZN(new_n4923_));
  NOR2_X1    g04859(.A1(new_n236_), .A2(new_n125_), .ZN(new_n4924_));
  AOI21_X1   g04860(.A1(new_n2401_), .A2(new_n4924_), .B(new_n939_), .ZN(new_n4925_));
  NOR2_X1    g04861(.A1(new_n2270_), .A2(new_n2511_), .ZN(new_n4926_));
  NOR4_X1    g04862(.A1(new_n1498_), .A2(new_n932_), .A3(new_n1589_), .A4(new_n1995_), .ZN(new_n4927_));
  NAND4_X1   g04863(.A1(new_n4927_), .A2(new_n2294_), .A3(new_n4925_), .A4(new_n4926_), .ZN(new_n4928_));
  NOR4_X1    g04864(.A1(new_n567_), .A2(new_n490_), .A3(new_n607_), .A4(new_n3218_), .ZN(new_n4929_));
  NOR3_X1    g04865(.A1(new_n1211_), .A2(new_n183_), .A3(new_n219_), .ZN(new_n4930_));
  NAND2_X1   g04866(.A1(new_n1222_), .A2(new_n501_), .ZN(new_n4931_));
  NOR3_X1    g04867(.A1(new_n4931_), .A2(new_n752_), .A3(new_n670_), .ZN(new_n4932_));
  INV_X1     g04868(.I(new_n4932_), .ZN(new_n4933_));
  NAND4_X1   g04869(.A1(new_n4929_), .A2(new_n3866_), .A3(new_n4930_), .A4(new_n4933_), .ZN(new_n4934_));
  NAND4_X1   g04870(.A1(new_n3846_), .A2(new_n599_), .A3(new_n1590_), .A4(new_n1100_), .ZN(new_n4935_));
  NOR3_X1    g04871(.A1(new_n406_), .A2(new_n86_), .A3(new_n307_), .ZN(new_n4936_));
  INV_X1     g04872(.I(new_n4936_), .ZN(new_n4937_));
  NOR4_X1    g04873(.A1(new_n615_), .A2(new_n955_), .A3(new_n510_), .A4(new_n459_), .ZN(new_n4938_));
  NOR3_X1    g04874(.A1(new_n4937_), .A2(new_n4935_), .A3(new_n4938_), .ZN(new_n4939_));
  INV_X1     g04875(.I(new_n3345_), .ZN(new_n4940_));
  NAND4_X1   g04876(.A1(new_n827_), .A2(new_n1767_), .A3(new_n3121_), .A4(new_n2191_), .ZN(new_n4941_));
  NOR2_X1    g04877(.A1(new_n4940_), .A2(new_n4941_), .ZN(new_n4942_));
  AND2_X2    g04878(.A1(new_n4942_), .A2(new_n4939_), .Z(new_n4943_));
  INV_X1     g04879(.I(new_n4943_), .ZN(new_n4944_));
  NOR4_X1    g04880(.A1(new_n4944_), .A2(new_n4923_), .A3(new_n4928_), .A4(new_n4934_), .ZN(new_n4945_));
  INV_X1     g04881(.I(new_n4945_), .ZN(new_n4946_));
  NAND2_X1   g04882(.A1(new_n4922_), .A2(new_n4946_), .ZN(new_n4947_));
  NOR2_X1    g04883(.A1(new_n4922_), .A2(new_n4946_), .ZN(new_n4948_));
  INV_X1     g04884(.I(new_n4948_), .ZN(new_n4949_));
  NAND2_X1   g04885(.A1(new_n4949_), .A2(new_n4947_), .ZN(new_n4950_));
  NAND2_X1   g04886(.A1(new_n4910_), .A2(new_n4950_), .ZN(new_n4951_));
  XOR2_X1    g04887(.A1(new_n4922_), .A2(new_n4945_), .Z(new_n4952_));
  OAI21_X1   g04888(.A1(new_n4910_), .A2(new_n4952_), .B(new_n4951_), .ZN(new_n4953_));
  AOI21_X1   g04889(.A1(new_n4541_), .A2(new_n2105_), .B(new_n2108_), .ZN(new_n4954_));
  XOR2_X1    g04890(.A1(new_n2102_), .A2(new_n2158_), .Z(new_n4955_));
  NOR2_X1    g04891(.A1(new_n2159_), .A2(new_n2162_), .ZN(new_n4956_));
  INV_X1     g04892(.I(new_n4956_), .ZN(new_n4957_));
  NAND3_X1   g04893(.A1(new_n2106_), .A2(new_n2109_), .A3(new_n4957_), .ZN(new_n4958_));
  OAI21_X1   g04894(.A1(new_n4954_), .A2(new_n4955_), .B(new_n4958_), .ZN(new_n4959_));
  OAI22_X1   g04895(.A1(new_n2103_), .A2(new_n2742_), .B1(new_n2158_), .B2(new_n3175_), .ZN(new_n4960_));
  NAND2_X1   g04896(.A1(new_n2107_), .A2(new_n2746_), .ZN(new_n4961_));
  AOI21_X1   g04897(.A1(new_n4960_), .A2(new_n4961_), .B(new_n2737_), .ZN(new_n4962_));
  NAND2_X1   g04898(.A1(new_n4959_), .A2(new_n4962_), .ZN(new_n4963_));
  XOR2_X1    g04899(.A1(new_n4963_), .A2(new_n74_), .Z(new_n4964_));
  XOR2_X1    g04900(.A1(new_n4964_), .A2(new_n4953_), .Z(new_n4965_));
  INV_X1     g04901(.I(new_n4965_), .ZN(new_n4966_));
  NOR2_X1    g04902(.A1(new_n1999_), .A2(new_n2734_), .ZN(new_n4967_));
  INV_X1     g04903(.I(new_n4967_), .ZN(new_n4968_));
  OAI22_X1   g04904(.A1(new_n1729_), .A2(new_n3318_), .B1(new_n4745_), .B2(new_n3268_), .ZN(new_n4969_));
  NAND2_X1   g04905(.A1(new_n1862_), .A2(new_n3323_), .ZN(new_n4970_));
  AOI21_X1   g04906(.A1(new_n4969_), .A2(new_n4970_), .B(new_n3260_), .ZN(new_n4971_));
  NAND2_X1   g04907(.A1(new_n4842_), .A2(new_n4971_), .ZN(new_n4972_));
  XOR2_X1    g04908(.A1(new_n4972_), .A2(new_n72_), .Z(new_n4973_));
  NAND2_X1   g04909(.A1(new_n4973_), .A2(new_n4968_), .ZN(new_n4974_));
  AOI22_X1   g04910(.A1(new_n4766_), .A2(new_n3267_), .B1(new_n1813_), .B2(new_n3323_), .ZN(new_n4975_));
  AOI21_X1   g04911(.A1(new_n1862_), .A2(new_n3317_), .B(new_n4975_), .ZN(new_n4976_));
  NOR3_X1    g04912(.A1(new_n4976_), .A2(new_n4878_), .A3(new_n3260_), .ZN(new_n4977_));
  XOR2_X1    g04913(.A1(new_n4977_), .A2(new_n72_), .Z(new_n4978_));
  NOR2_X1    g04914(.A1(new_n1999_), .A2(new_n4745_), .ZN(new_n4979_));
  NOR2_X1    g04915(.A1(new_n4766_), .A2(new_n1813_), .ZN(new_n4980_));
  NOR2_X1    g04916(.A1(new_n4979_), .A2(new_n4980_), .ZN(new_n4981_));
  NAND2_X1   g04917(.A1(new_n1813_), .A2(new_n3317_), .ZN(new_n4982_));
  NAND2_X1   g04918(.A1(new_n4766_), .A2(new_n3323_), .ZN(new_n4983_));
  NAND4_X1   g04919(.A1(new_n4981_), .A2(new_n3259_), .A3(new_n4982_), .A4(new_n4983_), .ZN(new_n4984_));
  XOR2_X1    g04920(.A1(new_n4984_), .A2(\a[26] ), .Z(new_n4985_));
  NOR2_X1    g04921(.A1(new_n1999_), .A2(new_n3257_), .ZN(new_n4986_));
  NOR2_X1    g04922(.A1(new_n4986_), .A2(new_n72_), .ZN(new_n4987_));
  NAND3_X1   g04923(.A1(new_n4978_), .A2(new_n4985_), .A3(new_n4987_), .ZN(new_n4988_));
  INV_X1     g04924(.I(new_n4988_), .ZN(new_n4989_));
  NOR2_X1    g04925(.A1(new_n4973_), .A2(new_n4968_), .ZN(new_n4990_));
  OAI21_X1   g04926(.A1(new_n4989_), .A2(new_n4990_), .B(new_n4974_), .ZN(new_n4991_));
  NAND2_X1   g04927(.A1(new_n1813_), .A2(new_n2750_), .ZN(new_n4992_));
  NAND2_X1   g04928(.A1(new_n4766_), .A2(new_n3275_), .ZN(new_n4993_));
  NAND4_X1   g04929(.A1(new_n4981_), .A2(new_n2736_), .A3(new_n4992_), .A4(new_n4993_), .ZN(new_n4994_));
  XOR2_X1    g04930(.A1(new_n4994_), .A2(new_n74_), .Z(new_n4995_));
  NOR2_X1    g04931(.A1(new_n4967_), .A2(new_n74_), .ZN(new_n4996_));
  XNOR2_X1   g04932(.A1(new_n4995_), .A2(new_n4996_), .ZN(new_n4997_));
  OAI22_X1   g04933(.A1(new_n1764_), .A2(new_n3318_), .B1(new_n1729_), .B2(new_n3322_), .ZN(new_n4998_));
  NAND2_X1   g04934(.A1(new_n1862_), .A2(new_n3267_), .ZN(new_n4999_));
  AOI21_X1   g04935(.A1(new_n4998_), .A2(new_n4999_), .B(new_n3260_), .ZN(new_n5000_));
  NAND2_X1   g04936(.A1(new_n4810_), .A2(new_n5000_), .ZN(new_n5001_));
  XOR2_X1    g04937(.A1(new_n5001_), .A2(\a[26] ), .Z(new_n5002_));
  NAND2_X1   g04938(.A1(new_n5002_), .A2(new_n4997_), .ZN(new_n5003_));
  NOR2_X1    g04939(.A1(new_n5002_), .A2(new_n4997_), .ZN(new_n5004_));
  AOI21_X1   g04940(.A1(new_n4991_), .A2(new_n5003_), .B(new_n5004_), .ZN(new_n5005_));
  AOI22_X1   g04941(.A1(new_n4766_), .A2(new_n2746_), .B1(new_n1813_), .B2(new_n3275_), .ZN(new_n5006_));
  AOI21_X1   g04942(.A1(new_n1862_), .A2(new_n2750_), .B(new_n5006_), .ZN(new_n5007_));
  NOR3_X1    g04943(.A1(new_n5007_), .A2(new_n4878_), .A3(new_n2737_), .ZN(new_n5008_));
  XOR2_X1    g04944(.A1(new_n5008_), .A2(\a[29] ), .Z(new_n5009_));
  NOR3_X1    g04945(.A1(new_n4994_), .A2(new_n74_), .A3(new_n4967_), .ZN(new_n5010_));
  XOR2_X1    g04946(.A1(new_n5009_), .A2(new_n5010_), .Z(new_n5011_));
  OAI22_X1   g04947(.A1(new_n1764_), .A2(new_n3322_), .B1(new_n1729_), .B2(new_n3268_), .ZN(new_n5012_));
  NAND2_X1   g04948(.A1(new_n1613_), .A2(new_n3317_), .ZN(new_n5013_));
  AOI21_X1   g04949(.A1(new_n5013_), .A2(new_n5012_), .B(new_n3260_), .ZN(new_n5014_));
  NAND2_X1   g04950(.A1(new_n4778_), .A2(new_n5014_), .ZN(new_n5015_));
  XOR2_X1    g04951(.A1(new_n5015_), .A2(new_n72_), .Z(new_n5016_));
  NOR2_X1    g04952(.A1(new_n5016_), .A2(new_n5011_), .ZN(new_n5017_));
  NAND2_X1   g04953(.A1(new_n5016_), .A2(new_n5011_), .ZN(new_n5018_));
  OAI21_X1   g04954(.A1(new_n5005_), .A2(new_n5017_), .B(new_n5018_), .ZN(new_n5019_));
  NOR4_X1    g04955(.A1(new_n5009_), .A2(new_n74_), .A3(new_n4967_), .A4(new_n4995_), .ZN(new_n5020_));
  NOR2_X1    g04956(.A1(new_n2764_), .A2(new_n3332_), .ZN(new_n5021_));
  NOR2_X1    g04957(.A1(new_n1999_), .A2(new_n5021_), .ZN(new_n5022_));
  OAI22_X1   g04958(.A1(new_n1729_), .A2(new_n3175_), .B1(new_n4745_), .B2(new_n2747_), .ZN(new_n5023_));
  NAND2_X1   g04959(.A1(new_n1862_), .A2(new_n3275_), .ZN(new_n5024_));
  AOI21_X1   g04960(.A1(new_n5023_), .A2(new_n5024_), .B(new_n2737_), .ZN(new_n5025_));
  NAND2_X1   g04961(.A1(new_n4842_), .A2(new_n5025_), .ZN(new_n5026_));
  XOR2_X1    g04962(.A1(new_n5026_), .A2(\a[29] ), .Z(new_n5027_));
  NOR2_X1    g04963(.A1(new_n5027_), .A2(new_n5022_), .ZN(new_n5028_));
  INV_X1     g04964(.I(new_n5022_), .ZN(new_n5029_));
  XOR2_X1    g04965(.A1(new_n5026_), .A2(new_n74_), .Z(new_n5030_));
  NOR2_X1    g04966(.A1(new_n5030_), .A2(new_n5029_), .ZN(new_n5031_));
  OAI21_X1   g04967(.A1(new_n5028_), .A2(new_n5031_), .B(new_n5020_), .ZN(new_n5032_));
  INV_X1     g04968(.I(new_n5009_), .ZN(new_n5033_));
  NAND2_X1   g04969(.A1(new_n5033_), .A2(new_n5010_), .ZN(new_n5034_));
  NOR2_X1    g04970(.A1(new_n5030_), .A2(new_n5022_), .ZN(new_n5035_));
  NOR2_X1    g04971(.A1(new_n5027_), .A2(new_n5029_), .ZN(new_n5036_));
  OAI21_X1   g04972(.A1(new_n5035_), .A2(new_n5036_), .B(new_n5034_), .ZN(new_n5037_));
  NAND2_X1   g04973(.A1(new_n5032_), .A2(new_n5037_), .ZN(new_n5038_));
  OAI22_X1   g04974(.A1(new_n1678_), .A2(new_n3318_), .B1(new_n1764_), .B2(new_n3268_), .ZN(new_n5039_));
  NAND2_X1   g04975(.A1(new_n1613_), .A2(new_n3323_), .ZN(new_n5040_));
  AOI21_X1   g04976(.A1(new_n5039_), .A2(new_n5040_), .B(new_n3260_), .ZN(new_n5041_));
  NAND2_X1   g04977(.A1(new_n4917_), .A2(new_n5041_), .ZN(new_n5042_));
  XOR2_X1    g04978(.A1(new_n5042_), .A2(\a[26] ), .Z(new_n5043_));
  NAND2_X1   g04979(.A1(new_n5038_), .A2(new_n5043_), .ZN(new_n5044_));
  NOR2_X1    g04980(.A1(new_n5038_), .A2(new_n5043_), .ZN(new_n5045_));
  AOI21_X1   g04981(.A1(new_n5019_), .A2(new_n5044_), .B(new_n5045_), .ZN(new_n5046_));
  NAND2_X1   g04982(.A1(new_n5030_), .A2(new_n5029_), .ZN(new_n5047_));
  OAI21_X1   g04983(.A1(new_n5020_), .A2(new_n5031_), .B(new_n5047_), .ZN(new_n5048_));
  OAI22_X1   g04984(.A1(new_n1764_), .A2(new_n3175_), .B1(new_n1729_), .B2(new_n2742_), .ZN(new_n5049_));
  NAND2_X1   g04985(.A1(new_n1862_), .A2(new_n2746_), .ZN(new_n5050_));
  AOI21_X1   g04986(.A1(new_n5049_), .A2(new_n5050_), .B(new_n2737_), .ZN(new_n5051_));
  NAND2_X1   g04987(.A1(new_n4810_), .A2(new_n5051_), .ZN(new_n5052_));
  XOR2_X1    g04988(.A1(new_n5052_), .A2(new_n74_), .Z(new_n5053_));
  AOI22_X1   g04989(.A1(new_n4766_), .A2(new_n3189_), .B1(new_n1813_), .B2(new_n3332_), .ZN(new_n5054_));
  AOI21_X1   g04990(.A1(new_n4981_), .A2(new_n2764_), .B(new_n5054_), .ZN(new_n5055_));
  NOR2_X1    g04991(.A1(new_n5053_), .A2(new_n5055_), .ZN(new_n5056_));
  XOR2_X1    g04992(.A1(new_n5052_), .A2(\a[29] ), .Z(new_n5057_));
  INV_X1     g04993(.I(new_n5055_), .ZN(new_n5058_));
  NOR2_X1    g04994(.A1(new_n5057_), .A2(new_n5058_), .ZN(new_n5059_));
  OAI21_X1   g04995(.A1(new_n5056_), .A2(new_n5059_), .B(new_n5048_), .ZN(new_n5060_));
  NAND2_X1   g04996(.A1(new_n5027_), .A2(new_n5022_), .ZN(new_n5061_));
  AOI21_X1   g04997(.A1(new_n5034_), .A2(new_n5061_), .B(new_n5028_), .ZN(new_n5062_));
  NOR2_X1    g04998(.A1(new_n5057_), .A2(new_n5055_), .ZN(new_n5063_));
  NOR2_X1    g04999(.A1(new_n5053_), .A2(new_n5058_), .ZN(new_n5064_));
  OAI21_X1   g05000(.A1(new_n5063_), .A2(new_n5064_), .B(new_n5062_), .ZN(new_n5065_));
  NAND2_X1   g05001(.A1(new_n5065_), .A2(new_n5060_), .ZN(new_n5066_));
  AOI21_X1   g05002(.A1(new_n4913_), .A2(new_n2004_), .B(new_n2074_), .ZN(new_n5067_));
  NOR3_X1    g05003(.A1(new_n2003_), .A2(new_n2005_), .A3(new_n1678_), .ZN(new_n5068_));
  OAI21_X1   g05004(.A1(new_n5068_), .A2(new_n5067_), .B(new_n4914_), .ZN(new_n5069_));
  XOR2_X1    g05005(.A1(new_n5069_), .A2(new_n2107_), .Z(new_n5070_));
  OAI22_X1   g05006(.A1(new_n1678_), .A2(new_n3322_), .B1(new_n2071_), .B2(new_n3318_), .ZN(new_n5071_));
  NAND2_X1   g05007(.A1(new_n1613_), .A2(new_n3267_), .ZN(new_n5072_));
  AOI21_X1   g05008(.A1(new_n5071_), .A2(new_n5072_), .B(new_n3260_), .ZN(new_n5073_));
  NAND3_X1   g05009(.A1(new_n5070_), .A2(new_n72_), .A3(new_n5073_), .ZN(new_n5074_));
  AOI21_X1   g05010(.A1(new_n5070_), .A2(new_n5073_), .B(new_n72_), .ZN(new_n5075_));
  INV_X1     g05011(.I(new_n5075_), .ZN(new_n5076_));
  NAND2_X1   g05012(.A1(new_n5076_), .A2(new_n5074_), .ZN(new_n5077_));
  NOR2_X1    g05013(.A1(new_n5077_), .A2(new_n5066_), .ZN(new_n5078_));
  NAND2_X1   g05014(.A1(new_n5077_), .A2(new_n5066_), .ZN(new_n5079_));
  OAI21_X1   g05015(.A1(new_n5046_), .A2(new_n5078_), .B(new_n5079_), .ZN(new_n5080_));
  NAND2_X1   g05016(.A1(new_n5053_), .A2(new_n5055_), .ZN(new_n5081_));
  OAI21_X1   g05017(.A1(new_n5062_), .A2(new_n5056_), .B(new_n5081_), .ZN(new_n5082_));
  OAI22_X1   g05018(.A1(new_n1764_), .A2(new_n2742_), .B1(new_n1729_), .B2(new_n2747_), .ZN(new_n5083_));
  NAND2_X1   g05019(.A1(new_n1613_), .A2(new_n2750_), .ZN(new_n5084_));
  AOI21_X1   g05020(.A1(new_n5084_), .A2(new_n5083_), .B(new_n2737_), .ZN(new_n5085_));
  NAND2_X1   g05021(.A1(new_n4778_), .A2(new_n5085_), .ZN(new_n5086_));
  XOR2_X1    g05022(.A1(new_n5086_), .A2(\a[29] ), .Z(new_n5087_));
  NAND2_X1   g05023(.A1(new_n4882_), .A2(new_n4900_), .ZN(new_n5088_));
  AND2_X2    g05024(.A1(new_n4901_), .A2(new_n5088_), .Z(new_n5089_));
  INV_X1     g05025(.I(new_n5089_), .ZN(new_n5090_));
  NOR2_X1    g05026(.A1(new_n5087_), .A2(new_n5090_), .ZN(new_n5091_));
  XOR2_X1    g05027(.A1(new_n5086_), .A2(new_n74_), .Z(new_n5092_));
  NOR2_X1    g05028(.A1(new_n5092_), .A2(new_n5089_), .ZN(new_n5093_));
  OAI21_X1   g05029(.A1(new_n5091_), .A2(new_n5093_), .B(new_n5082_), .ZN(new_n5094_));
  NAND2_X1   g05030(.A1(new_n5087_), .A2(new_n5089_), .ZN(new_n5095_));
  NAND2_X1   g05031(.A1(new_n5092_), .A2(new_n5090_), .ZN(new_n5096_));
  AOI21_X1   g05032(.A1(new_n5095_), .A2(new_n5096_), .B(new_n5082_), .ZN(new_n5097_));
  INV_X1     g05033(.I(new_n5097_), .ZN(new_n5098_));
  OAI22_X1   g05034(.A1(new_n2103_), .A2(new_n3318_), .B1(new_n1678_), .B2(new_n3268_), .ZN(new_n5099_));
  NAND2_X1   g05035(.A1(new_n2107_), .A2(new_n3323_), .ZN(new_n5100_));
  AOI21_X1   g05036(.A1(new_n5099_), .A2(new_n5100_), .B(new_n3260_), .ZN(new_n5101_));
  NAND3_X1   g05037(.A1(new_n4545_), .A2(new_n72_), .A3(new_n5101_), .ZN(new_n5102_));
  AND3_X2    g05038(.A1(new_n2073_), .A2(new_n2076_), .A3(new_n4542_), .Z(new_n5103_));
  NOR2_X1    g05039(.A1(new_n4541_), .A2(new_n4544_), .ZN(new_n5104_));
  OAI21_X1   g05040(.A1(new_n5103_), .A2(new_n5104_), .B(new_n5101_), .ZN(new_n5105_));
  NAND2_X1   g05041(.A1(new_n5105_), .A2(\a[26] ), .ZN(new_n5106_));
  NAND2_X1   g05042(.A1(new_n5102_), .A2(new_n5106_), .ZN(new_n5107_));
  AOI21_X1   g05043(.A1(new_n5098_), .A2(new_n5094_), .B(new_n5107_), .ZN(new_n5108_));
  INV_X1     g05044(.I(new_n5108_), .ZN(new_n5109_));
  INV_X1     g05045(.I(new_n5094_), .ZN(new_n5110_));
  INV_X1     g05046(.I(new_n5107_), .ZN(new_n5111_));
  NOR3_X1    g05047(.A1(new_n5111_), .A2(new_n5110_), .A3(new_n5097_), .ZN(new_n5112_));
  AOI21_X1   g05048(.A1(new_n5109_), .A2(new_n5080_), .B(new_n5112_), .ZN(new_n5113_));
  NOR2_X1    g05049(.A1(new_n5087_), .A2(new_n5089_), .ZN(new_n5114_));
  AOI21_X1   g05050(.A1(new_n5082_), .A2(new_n5095_), .B(new_n5114_), .ZN(new_n5115_));
  OAI22_X1   g05051(.A1(new_n1678_), .A2(new_n3175_), .B1(new_n1764_), .B2(new_n2747_), .ZN(new_n5116_));
  NAND2_X1   g05052(.A1(new_n1613_), .A2(new_n3275_), .ZN(new_n5117_));
  AOI21_X1   g05053(.A1(new_n5116_), .A2(new_n5117_), .B(new_n2737_), .ZN(new_n5118_));
  NAND3_X1   g05054(.A1(new_n4917_), .A2(new_n74_), .A3(new_n5118_), .ZN(new_n5119_));
  NAND2_X1   g05055(.A1(new_n4917_), .A2(new_n5118_), .ZN(new_n5120_));
  NAND2_X1   g05056(.A1(new_n5120_), .A2(\a[29] ), .ZN(new_n5121_));
  NAND2_X1   g05057(.A1(new_n5121_), .A2(new_n5119_), .ZN(new_n5122_));
  XOR2_X1    g05058(.A1(new_n4902_), .A2(new_n4870_), .Z(new_n5123_));
  NOR2_X1    g05059(.A1(new_n5123_), .A2(new_n4901_), .ZN(new_n5124_));
  NAND2_X1   g05060(.A1(new_n4903_), .A2(new_n4875_), .ZN(new_n5125_));
  AOI21_X1   g05061(.A1(new_n4901_), .A2(new_n5125_), .B(new_n5124_), .ZN(new_n5126_));
  NAND2_X1   g05062(.A1(new_n5122_), .A2(new_n5126_), .ZN(new_n5127_));
  INV_X1     g05063(.I(new_n5122_), .ZN(new_n5128_));
  INV_X1     g05064(.I(new_n5126_), .ZN(new_n5129_));
  NAND2_X1   g05065(.A1(new_n5128_), .A2(new_n5129_), .ZN(new_n5130_));
  AOI21_X1   g05066(.A1(new_n5127_), .A2(new_n5130_), .B(new_n5115_), .ZN(new_n5131_));
  INV_X1     g05067(.I(new_n5115_), .ZN(new_n5132_));
  NOR2_X1    g05068(.A1(new_n5129_), .A2(new_n5122_), .ZN(new_n5133_));
  NOR2_X1    g05069(.A1(new_n5128_), .A2(new_n5126_), .ZN(new_n5134_));
  NOR2_X1    g05070(.A1(new_n5134_), .A2(new_n5133_), .ZN(new_n5135_));
  NOR2_X1    g05071(.A1(new_n5132_), .A2(new_n5135_), .ZN(new_n5136_));
  NOR2_X1    g05072(.A1(new_n5136_), .A2(new_n5131_), .ZN(new_n5137_));
  OAI22_X1   g05073(.A1(new_n2103_), .A2(new_n3322_), .B1(new_n2158_), .B2(new_n3318_), .ZN(new_n5138_));
  NAND2_X1   g05074(.A1(new_n2107_), .A2(new_n3267_), .ZN(new_n5139_));
  AOI21_X1   g05075(.A1(new_n5138_), .A2(new_n5139_), .B(new_n3260_), .ZN(new_n5140_));
  NAND3_X1   g05076(.A1(new_n4959_), .A2(new_n72_), .A3(new_n5140_), .ZN(new_n5141_));
  AOI21_X1   g05077(.A1(new_n4959_), .A2(new_n5140_), .B(new_n72_), .ZN(new_n5142_));
  INV_X1     g05078(.I(new_n5142_), .ZN(new_n5143_));
  NAND2_X1   g05079(.A1(new_n5143_), .A2(new_n5141_), .ZN(new_n5144_));
  NOR2_X1    g05080(.A1(new_n5137_), .A2(new_n5144_), .ZN(new_n5145_));
  NAND2_X1   g05081(.A1(new_n5137_), .A2(new_n5144_), .ZN(new_n5146_));
  OAI21_X1   g05082(.A1(new_n5113_), .A2(new_n5145_), .B(new_n5146_), .ZN(new_n5147_));
  NAND2_X1   g05083(.A1(new_n5129_), .A2(new_n5122_), .ZN(new_n5148_));
  OAI21_X1   g05084(.A1(new_n5115_), .A2(new_n5133_), .B(new_n5148_), .ZN(new_n5149_));
  OAI22_X1   g05085(.A1(new_n1678_), .A2(new_n2742_), .B1(new_n2071_), .B2(new_n3175_), .ZN(new_n5150_));
  NAND2_X1   g05086(.A1(new_n1613_), .A2(new_n2746_), .ZN(new_n5151_));
  AOI21_X1   g05087(.A1(new_n5150_), .A2(new_n5151_), .B(new_n2737_), .ZN(new_n5152_));
  NAND3_X1   g05088(.A1(new_n5070_), .A2(new_n74_), .A3(new_n5152_), .ZN(new_n5153_));
  INV_X1     g05089(.I(new_n5153_), .ZN(new_n5154_));
  AOI21_X1   g05090(.A1(new_n5070_), .A2(new_n5152_), .B(new_n74_), .ZN(new_n5155_));
  NOR2_X1    g05091(.A1(new_n5154_), .A2(new_n5155_), .ZN(new_n5156_));
  NAND2_X1   g05092(.A1(new_n4904_), .A2(new_n4875_), .ZN(new_n5157_));
  XOR2_X1    g05093(.A1(new_n4815_), .A2(new_n4830_), .Z(new_n5158_));
  XOR2_X1    g05094(.A1(new_n4815_), .A2(new_n4830_), .Z(new_n5159_));
  NOR2_X1    g05095(.A1(new_n5159_), .A2(new_n5157_), .ZN(new_n5160_));
  AOI21_X1   g05096(.A1(new_n5157_), .A2(new_n5158_), .B(new_n5160_), .ZN(new_n5161_));
  INV_X1     g05097(.I(new_n5161_), .ZN(new_n5162_));
  NOR2_X1    g05098(.A1(new_n5156_), .A2(new_n5162_), .ZN(new_n5163_));
  INV_X1     g05099(.I(new_n5155_), .ZN(new_n5164_));
  NAND2_X1   g05100(.A1(new_n5164_), .A2(new_n5153_), .ZN(new_n5165_));
  NOR2_X1    g05101(.A1(new_n5165_), .A2(new_n5161_), .ZN(new_n5166_));
  OAI21_X1   g05102(.A1(new_n5166_), .A2(new_n5163_), .B(new_n5149_), .ZN(new_n5167_));
  INV_X1     g05103(.I(new_n5149_), .ZN(new_n5168_));
  NOR2_X1    g05104(.A1(new_n5165_), .A2(new_n5162_), .ZN(new_n5169_));
  NOR2_X1    g05105(.A1(new_n5156_), .A2(new_n5161_), .ZN(new_n5170_));
  OAI21_X1   g05106(.A1(new_n5169_), .A2(new_n5170_), .B(new_n5168_), .ZN(new_n5171_));
  NAND2_X1   g05107(.A1(new_n5171_), .A2(new_n5167_), .ZN(new_n5172_));
  XNOR2_X1   g05108(.A1(new_n2158_), .A2(new_n2198_), .ZN(new_n5173_));
  INV_X1     g05109(.I(new_n5173_), .ZN(new_n5174_));
  OAI21_X1   g05110(.A1(new_n2160_), .A2(new_n2162_), .B(new_n5174_), .ZN(new_n5175_));
  INV_X1     g05111(.I(new_n5175_), .ZN(new_n5176_));
  NOR2_X1    g05112(.A1(new_n2203_), .A2(new_n2199_), .ZN(new_n5177_));
  NOR3_X1    g05113(.A1(new_n2160_), .A2(new_n2162_), .A3(new_n5177_), .ZN(new_n5178_));
  OAI22_X1   g05114(.A1(new_n2103_), .A2(new_n3268_), .B1(new_n2198_), .B2(new_n3318_), .ZN(new_n5179_));
  NAND2_X1   g05115(.A1(new_n2161_), .A2(new_n3323_), .ZN(new_n5180_));
  AOI21_X1   g05116(.A1(new_n5179_), .A2(new_n5180_), .B(new_n3260_), .ZN(new_n5181_));
  OAI21_X1   g05117(.A1(new_n5176_), .A2(new_n5178_), .B(new_n5181_), .ZN(new_n5182_));
  XOR2_X1    g05118(.A1(new_n5182_), .A2(\a[26] ), .Z(new_n5183_));
  NAND2_X1   g05119(.A1(new_n5172_), .A2(new_n5183_), .ZN(new_n5184_));
  INV_X1     g05120(.I(new_n5167_), .ZN(new_n5185_));
  NAND2_X1   g05121(.A1(new_n5156_), .A2(new_n5161_), .ZN(new_n5186_));
  NAND2_X1   g05122(.A1(new_n5165_), .A2(new_n5162_), .ZN(new_n5187_));
  AOI21_X1   g05123(.A1(new_n5187_), .A2(new_n5186_), .B(new_n5149_), .ZN(new_n5188_));
  NOR3_X1    g05124(.A1(new_n5183_), .A2(new_n5185_), .A3(new_n5188_), .ZN(new_n5189_));
  AOI21_X1   g05125(.A1(new_n5147_), .A2(new_n5184_), .B(new_n5189_), .ZN(new_n5190_));
  AOI21_X1   g05126(.A1(new_n5186_), .A2(new_n5149_), .B(new_n5170_), .ZN(new_n5191_));
  OAI22_X1   g05127(.A1(new_n2103_), .A2(new_n3175_), .B1(new_n1678_), .B2(new_n2747_), .ZN(new_n5192_));
  NAND2_X1   g05128(.A1(new_n2107_), .A2(new_n3275_), .ZN(new_n5193_));
  AOI21_X1   g05129(.A1(new_n5192_), .A2(new_n5193_), .B(new_n2737_), .ZN(new_n5194_));
  NAND3_X1   g05130(.A1(new_n4545_), .A2(new_n74_), .A3(new_n5194_), .ZN(new_n5195_));
  AOI21_X1   g05131(.A1(new_n4545_), .A2(new_n5194_), .B(new_n74_), .ZN(new_n5196_));
  INV_X1     g05132(.I(new_n5196_), .ZN(new_n5197_));
  AOI21_X1   g05133(.A1(new_n4908_), .A2(new_n4803_), .B(new_n4906_), .ZN(new_n5198_));
  XNOR2_X1   g05134(.A1(new_n4783_), .A2(new_n4802_), .ZN(new_n5199_));
  NOR2_X1    g05135(.A1(new_n4907_), .A2(new_n5199_), .ZN(new_n5200_));
  NOR2_X1    g05136(.A1(new_n5200_), .A2(new_n5198_), .ZN(new_n5201_));
  INV_X1     g05137(.I(new_n5201_), .ZN(new_n5202_));
  AOI21_X1   g05138(.A1(new_n5197_), .A2(new_n5195_), .B(new_n5202_), .ZN(new_n5203_));
  INV_X1     g05139(.I(new_n5195_), .ZN(new_n5204_));
  NOR3_X1    g05140(.A1(new_n5204_), .A2(new_n5201_), .A3(new_n5196_), .ZN(new_n5205_));
  NOR2_X1    g05141(.A1(new_n5203_), .A2(new_n5205_), .ZN(new_n5206_));
  NOR2_X1    g05142(.A1(new_n5206_), .A2(new_n5191_), .ZN(new_n5207_));
  NAND3_X1   g05143(.A1(new_n5197_), .A2(new_n5201_), .A3(new_n5195_), .ZN(new_n5208_));
  OAI21_X1   g05144(.A1(new_n5204_), .A2(new_n5196_), .B(new_n5202_), .ZN(new_n5209_));
  NAND2_X1   g05145(.A1(new_n5209_), .A2(new_n5208_), .ZN(new_n5210_));
  AOI21_X1   g05146(.A1(new_n5191_), .A2(new_n5210_), .B(new_n5207_), .ZN(new_n5211_));
  OAI22_X1   g05147(.A1(new_n2158_), .A2(new_n3268_), .B1(new_n2198_), .B2(new_n3322_), .ZN(new_n5212_));
  NAND2_X1   g05148(.A1(new_n1504_), .A2(new_n3317_), .ZN(new_n5213_));
  AOI21_X1   g05149(.A1(new_n5213_), .A2(new_n5212_), .B(new_n3260_), .ZN(new_n5214_));
  NAND3_X1   g05150(.A1(new_n4620_), .A2(new_n72_), .A3(new_n5214_), .ZN(new_n5215_));
  AOI21_X1   g05151(.A1(new_n4620_), .A2(new_n5214_), .B(new_n72_), .ZN(new_n5216_));
  INV_X1     g05152(.I(new_n5216_), .ZN(new_n5217_));
  NAND2_X1   g05153(.A1(new_n5217_), .A2(new_n5215_), .ZN(new_n5218_));
  NOR2_X1    g05154(.A1(new_n5211_), .A2(new_n5218_), .ZN(new_n5219_));
  NAND2_X1   g05155(.A1(new_n5211_), .A2(new_n5218_), .ZN(new_n5220_));
  OAI21_X1   g05156(.A1(new_n5190_), .A2(new_n5219_), .B(new_n5220_), .ZN(new_n5221_));
  NOR3_X1    g05157(.A1(new_n5202_), .A2(new_n5204_), .A3(new_n5196_), .ZN(new_n5222_));
  OAI21_X1   g05158(.A1(new_n5191_), .A2(new_n5222_), .B(new_n5209_), .ZN(new_n5223_));
  INV_X1     g05159(.I(new_n5223_), .ZN(new_n5224_));
  NOR2_X1    g05160(.A1(new_n5221_), .A2(new_n5224_), .ZN(new_n5225_));
  XOR2_X1    g05161(.A1(new_n4972_), .A2(\a[26] ), .Z(new_n5226_));
  NOR2_X1    g05162(.A1(new_n5226_), .A2(new_n4967_), .ZN(new_n5227_));
  NAND2_X1   g05163(.A1(new_n5226_), .A2(new_n4967_), .ZN(new_n5228_));
  AOI21_X1   g05164(.A1(new_n4988_), .A2(new_n5228_), .B(new_n5227_), .ZN(new_n5229_));
  XOR2_X1    g05165(.A1(new_n4995_), .A2(new_n4996_), .Z(new_n5230_));
  XOR2_X1    g05166(.A1(new_n5001_), .A2(new_n72_), .Z(new_n5231_));
  NOR2_X1    g05167(.A1(new_n5231_), .A2(new_n5230_), .ZN(new_n5232_));
  NAND2_X1   g05168(.A1(new_n5231_), .A2(new_n5230_), .ZN(new_n5233_));
  OAI21_X1   g05169(.A1(new_n5229_), .A2(new_n5232_), .B(new_n5233_), .ZN(new_n5234_));
  INV_X1     g05170(.I(new_n5011_), .ZN(new_n5235_));
  XOR2_X1    g05171(.A1(new_n5015_), .A2(\a[26] ), .Z(new_n5236_));
  NAND2_X1   g05172(.A1(new_n5236_), .A2(new_n5235_), .ZN(new_n5237_));
  NOR2_X1    g05173(.A1(new_n5236_), .A2(new_n5235_), .ZN(new_n5238_));
  AOI21_X1   g05174(.A1(new_n5234_), .A2(new_n5237_), .B(new_n5238_), .ZN(new_n5239_));
  AND2_X2    g05175(.A1(new_n5032_), .A2(new_n5037_), .Z(new_n5240_));
  XOR2_X1    g05176(.A1(new_n5042_), .A2(new_n72_), .Z(new_n5241_));
  NOR2_X1    g05177(.A1(new_n5240_), .A2(new_n5241_), .ZN(new_n5242_));
  NAND2_X1   g05178(.A1(new_n5240_), .A2(new_n5241_), .ZN(new_n5243_));
  OAI21_X1   g05179(.A1(new_n5239_), .A2(new_n5242_), .B(new_n5243_), .ZN(new_n5244_));
  NOR2_X1    g05180(.A1(new_n5056_), .A2(new_n5059_), .ZN(new_n5245_));
  NOR2_X1    g05181(.A1(new_n5063_), .A2(new_n5064_), .ZN(new_n5246_));
  MUX2_X1    g05182(.I0(new_n5246_), .I1(new_n5245_), .S(new_n5048_), .Z(new_n5247_));
  INV_X1     g05183(.I(new_n5074_), .ZN(new_n5248_));
  NOR2_X1    g05184(.A1(new_n5248_), .A2(new_n5075_), .ZN(new_n5249_));
  NAND2_X1   g05185(.A1(new_n5247_), .A2(new_n5249_), .ZN(new_n5250_));
  NOR2_X1    g05186(.A1(new_n5247_), .A2(new_n5249_), .ZN(new_n5251_));
  AOI21_X1   g05187(.A1(new_n5244_), .A2(new_n5250_), .B(new_n5251_), .ZN(new_n5252_));
  NAND3_X1   g05188(.A1(new_n5098_), .A2(new_n5107_), .A3(new_n5094_), .ZN(new_n5253_));
  OAI21_X1   g05189(.A1(new_n5252_), .A2(new_n5108_), .B(new_n5253_), .ZN(new_n5254_));
  NAND2_X1   g05190(.A1(new_n5130_), .A2(new_n5127_), .ZN(new_n5255_));
  NAND2_X1   g05191(.A1(new_n5132_), .A2(new_n5255_), .ZN(new_n5256_));
  OAI21_X1   g05192(.A1(new_n5133_), .A2(new_n5134_), .B(new_n5115_), .ZN(new_n5257_));
  NAND2_X1   g05193(.A1(new_n5256_), .A2(new_n5257_), .ZN(new_n5258_));
  AOI21_X1   g05194(.A1(new_n2106_), .A2(new_n2109_), .B(new_n4955_), .ZN(new_n5259_));
  INV_X1     g05195(.I(new_n4958_), .ZN(new_n5260_));
  OAI21_X1   g05196(.A1(new_n5260_), .A2(new_n5259_), .B(new_n5140_), .ZN(new_n5261_));
  NOR2_X1    g05197(.A1(new_n5261_), .A2(\a[26] ), .ZN(new_n5262_));
  NOR2_X1    g05198(.A1(new_n5262_), .A2(new_n5142_), .ZN(new_n5263_));
  NAND2_X1   g05199(.A1(new_n5258_), .A2(new_n5263_), .ZN(new_n5264_));
  NOR2_X1    g05200(.A1(new_n5258_), .A2(new_n5263_), .ZN(new_n5265_));
  AOI21_X1   g05201(.A1(new_n5254_), .A2(new_n5264_), .B(new_n5265_), .ZN(new_n5266_));
  XOR2_X1    g05202(.A1(new_n5182_), .A2(new_n72_), .Z(new_n5267_));
  AOI21_X1   g05203(.A1(new_n5167_), .A2(new_n5171_), .B(new_n5267_), .ZN(new_n5268_));
  NAND3_X1   g05204(.A1(new_n5267_), .A2(new_n5171_), .A3(new_n5167_), .ZN(new_n5269_));
  OAI21_X1   g05205(.A1(new_n5266_), .A2(new_n5268_), .B(new_n5269_), .ZN(new_n5270_));
  NOR2_X1    g05206(.A1(new_n5168_), .A2(new_n5169_), .ZN(new_n5271_));
  OAI22_X1   g05207(.A1(new_n5271_), .A2(new_n5170_), .B1(new_n5203_), .B2(new_n5205_), .ZN(new_n5272_));
  AOI21_X1   g05208(.A1(new_n5197_), .A2(new_n5195_), .B(new_n5201_), .ZN(new_n5273_));
  OAI21_X1   g05209(.A1(new_n5222_), .A2(new_n5273_), .B(new_n5191_), .ZN(new_n5274_));
  NAND2_X1   g05210(.A1(new_n5272_), .A2(new_n5274_), .ZN(new_n5275_));
  INV_X1     g05211(.I(new_n5215_), .ZN(new_n5276_));
  NOR2_X1    g05212(.A1(new_n5276_), .A2(new_n5216_), .ZN(new_n5277_));
  NAND2_X1   g05213(.A1(new_n5275_), .A2(new_n5277_), .ZN(new_n5278_));
  NAND2_X1   g05214(.A1(new_n5270_), .A2(new_n5278_), .ZN(new_n5279_));
  AOI21_X1   g05215(.A1(new_n5279_), .A2(new_n5220_), .B(new_n5223_), .ZN(new_n5280_));
  OAI21_X1   g05216(.A1(new_n5225_), .A2(new_n5280_), .B(new_n4966_), .ZN(new_n5281_));
  NAND3_X1   g05217(.A1(new_n5279_), .A2(new_n5220_), .A3(new_n5223_), .ZN(new_n5282_));
  NAND2_X1   g05218(.A1(new_n5221_), .A2(new_n5224_), .ZN(new_n5283_));
  NAND3_X1   g05219(.A1(new_n5283_), .A2(new_n5282_), .A3(new_n4965_), .ZN(new_n5284_));
  AOI21_X1   g05220(.A1(new_n5281_), .A2(new_n5284_), .B(new_n4737_), .ZN(new_n5285_));
  AOI21_X1   g05221(.A1(new_n5283_), .A2(new_n5282_), .B(new_n4965_), .ZN(new_n5286_));
  NOR3_X1    g05222(.A1(new_n5225_), .A2(new_n5280_), .A3(new_n4966_), .ZN(new_n5287_));
  NOR3_X1    g05223(.A1(new_n5287_), .A2(new_n5286_), .A3(new_n4736_), .ZN(new_n5288_));
  NAND2_X1   g05224(.A1(new_n2310_), .A2(new_n3782_), .ZN(new_n5289_));
  NAND2_X1   g05225(.A1(new_n2354_), .A2(new_n3312_), .ZN(new_n5290_));
  INV_X1     g05226(.I(new_n3310_), .ZN(new_n5291_));
  AOI21_X1   g05227(.A1(new_n2255_), .A2(new_n5291_), .B(new_n3302_), .ZN(new_n5292_));
  NAND4_X1   g05228(.A1(new_n3914_), .A2(new_n5289_), .A3(new_n5290_), .A4(new_n5292_), .ZN(new_n5293_));
  XOR2_X1    g05229(.A1(new_n5293_), .A2(new_n84_), .Z(new_n5294_));
  NOR3_X1    g05230(.A1(new_n5288_), .A2(new_n5285_), .A3(new_n5294_), .ZN(new_n5295_));
  OAI21_X1   g05231(.A1(new_n5287_), .A2(new_n5286_), .B(new_n4736_), .ZN(new_n5296_));
  NAND3_X1   g05232(.A1(new_n5281_), .A2(new_n5284_), .A3(new_n4737_), .ZN(new_n5297_));
  XOR2_X1    g05233(.A1(new_n5293_), .A2(\a[23] ), .Z(new_n5298_));
  AOI21_X1   g05234(.A1(new_n5296_), .A2(new_n5297_), .B(new_n5298_), .ZN(new_n5299_));
  OAI22_X1   g05235(.A1(new_n2251_), .A2(new_n3780_), .B1(new_n4365_), .B2(new_n3306_), .ZN(new_n5300_));
  NAND2_X1   g05236(.A1(new_n1504_), .A2(new_n5291_), .ZN(new_n5301_));
  AOI21_X1   g05237(.A1(new_n5300_), .A2(new_n5301_), .B(new_n3302_), .ZN(new_n5302_));
  NAND3_X1   g05238(.A1(new_n4650_), .A2(new_n84_), .A3(new_n5302_), .ZN(new_n5303_));
  AOI21_X1   g05239(.A1(new_n4650_), .A2(new_n5302_), .B(new_n84_), .ZN(new_n5304_));
  INV_X1     g05240(.I(new_n5304_), .ZN(new_n5305_));
  NAND2_X1   g05241(.A1(new_n5305_), .A2(new_n5303_), .ZN(new_n5306_));
  AOI21_X1   g05242(.A1(new_n5184_), .A2(new_n5269_), .B(new_n5266_), .ZN(new_n5307_));
  NAND3_X1   g05243(.A1(new_n5183_), .A2(new_n5171_), .A3(new_n5167_), .ZN(new_n5308_));
  NAND2_X1   g05244(.A1(new_n5172_), .A2(new_n5267_), .ZN(new_n5309_));
  AOI21_X1   g05245(.A1(new_n5308_), .A2(new_n5309_), .B(new_n5147_), .ZN(new_n5310_));
  NOR2_X1    g05246(.A1(new_n5310_), .A2(new_n5307_), .ZN(new_n5311_));
  NAND2_X1   g05247(.A1(new_n5306_), .A2(new_n5311_), .ZN(new_n5312_));
  INV_X1     g05248(.I(new_n5303_), .ZN(new_n5313_));
  NOR2_X1    g05249(.A1(new_n5313_), .A2(new_n5304_), .ZN(new_n5314_));
  OAI21_X1   g05250(.A1(new_n5268_), .A2(new_n5189_), .B(new_n5147_), .ZN(new_n5315_));
  NAND2_X1   g05251(.A1(new_n5309_), .A2(new_n5308_), .ZN(new_n5316_));
  NAND2_X1   g05252(.A1(new_n5316_), .A2(new_n5266_), .ZN(new_n5317_));
  NAND2_X1   g05253(.A1(new_n5317_), .A2(new_n5315_), .ZN(new_n5318_));
  NAND2_X1   g05254(.A1(new_n5314_), .A2(new_n5318_), .ZN(new_n5319_));
  OAI21_X1   g05255(.A1(new_n5145_), .A2(new_n5265_), .B(new_n5254_), .ZN(new_n5320_));
  NOR3_X1    g05256(.A1(new_n5144_), .A2(new_n5136_), .A3(new_n5131_), .ZN(new_n5321_));
  AOI21_X1   g05257(.A1(new_n5256_), .A2(new_n5257_), .B(new_n5263_), .ZN(new_n5322_));
  OAI21_X1   g05258(.A1(new_n5321_), .A2(new_n5322_), .B(new_n5113_), .ZN(new_n5323_));
  OAI22_X1   g05259(.A1(new_n4365_), .A2(new_n3780_), .B1(new_n2198_), .B2(new_n3310_), .ZN(new_n5324_));
  NAND2_X1   g05260(.A1(new_n1504_), .A2(new_n3782_), .ZN(new_n5325_));
  AOI21_X1   g05261(.A1(new_n5324_), .A2(new_n5325_), .B(new_n3302_), .ZN(new_n5326_));
  NAND3_X1   g05262(.A1(new_n4363_), .A2(new_n84_), .A3(new_n5326_), .ZN(new_n5327_));
  AOI21_X1   g05263(.A1(new_n4363_), .A2(new_n5326_), .B(new_n84_), .ZN(new_n5328_));
  INV_X1     g05264(.I(new_n5328_), .ZN(new_n5329_));
  NAND4_X1   g05265(.A1(new_n5323_), .A2(new_n5320_), .A3(new_n5327_), .A4(new_n5329_), .ZN(new_n5330_));
  AOI21_X1   g05266(.A1(new_n5264_), .A2(new_n5146_), .B(new_n5113_), .ZN(new_n5331_));
  NOR2_X1    g05267(.A1(new_n5321_), .A2(new_n5322_), .ZN(new_n5332_));
  NOR2_X1    g05268(.A1(new_n5332_), .A2(new_n5254_), .ZN(new_n5333_));
  INV_X1     g05269(.I(new_n5327_), .ZN(new_n5334_));
  NOR4_X1    g05270(.A1(new_n5331_), .A2(new_n5333_), .A3(new_n5334_), .A4(new_n5328_), .ZN(new_n5335_));
  AOI22_X1   g05271(.A1(new_n5323_), .A2(new_n5320_), .B1(new_n5327_), .B2(new_n5329_), .ZN(new_n5336_));
  NOR2_X1    g05272(.A1(new_n5336_), .A2(new_n5335_), .ZN(new_n5337_));
  AOI21_X1   g05273(.A1(new_n5109_), .A2(new_n5253_), .B(new_n5252_), .ZN(new_n5338_));
  NAND3_X1   g05274(.A1(new_n5111_), .A2(new_n5094_), .A3(new_n5098_), .ZN(new_n5339_));
  OAI21_X1   g05275(.A1(new_n5110_), .A2(new_n5097_), .B(new_n5107_), .ZN(new_n5340_));
  AOI21_X1   g05276(.A1(new_n5339_), .A2(new_n5340_), .B(new_n5080_), .ZN(new_n5341_));
  OAI22_X1   g05277(.A1(new_n2158_), .A2(new_n3310_), .B1(new_n2198_), .B2(new_n3306_), .ZN(new_n5342_));
  NAND2_X1   g05278(.A1(new_n1504_), .A2(new_n3312_), .ZN(new_n5343_));
  AOI21_X1   g05279(.A1(new_n5343_), .A2(new_n5342_), .B(new_n3302_), .ZN(new_n5344_));
  NAND3_X1   g05280(.A1(new_n4620_), .A2(new_n84_), .A3(new_n5344_), .ZN(new_n5345_));
  INV_X1     g05281(.I(new_n5345_), .ZN(new_n5346_));
  AOI21_X1   g05282(.A1(new_n4620_), .A2(new_n5344_), .B(new_n84_), .ZN(new_n5347_));
  NOR4_X1    g05283(.A1(new_n5338_), .A2(new_n5341_), .A3(new_n5346_), .A4(new_n5347_), .ZN(new_n5348_));
  INV_X1     g05284(.I(new_n5348_), .ZN(new_n5349_));
  OR3_X2     g05285(.A1(new_n2160_), .A2(new_n2162_), .A3(new_n5177_), .Z(new_n5350_));
  NAND2_X1   g05286(.A1(new_n5350_), .A2(new_n5175_), .ZN(new_n5351_));
  OAI22_X1   g05287(.A1(new_n2103_), .A2(new_n3310_), .B1(new_n2198_), .B2(new_n3780_), .ZN(new_n5352_));
  NAND2_X1   g05288(.A1(new_n2161_), .A2(new_n3782_), .ZN(new_n5353_));
  AOI21_X1   g05289(.A1(new_n5352_), .A2(new_n5353_), .B(new_n3302_), .ZN(new_n5354_));
  NAND3_X1   g05290(.A1(new_n5351_), .A2(new_n84_), .A3(new_n5354_), .ZN(new_n5355_));
  OAI21_X1   g05291(.A1(new_n5176_), .A2(new_n5178_), .B(new_n5354_), .ZN(new_n5356_));
  NAND2_X1   g05292(.A1(new_n5356_), .A2(\a[23] ), .ZN(new_n5357_));
  AND2_X2    g05293(.A1(new_n5357_), .A2(new_n5355_), .Z(new_n5358_));
  OAI21_X1   g05294(.A1(new_n5078_), .A2(new_n5251_), .B(new_n5244_), .ZN(new_n5359_));
  NOR2_X1    g05295(.A1(new_n5247_), .A2(new_n5077_), .ZN(new_n5360_));
  NOR2_X1    g05296(.A1(new_n5249_), .A2(new_n5066_), .ZN(new_n5361_));
  OAI21_X1   g05297(.A1(new_n5360_), .A2(new_n5361_), .B(new_n5046_), .ZN(new_n5362_));
  NAND2_X1   g05298(.A1(new_n5359_), .A2(new_n5362_), .ZN(new_n5363_));
  NAND2_X1   g05299(.A1(new_n5363_), .A2(new_n5358_), .ZN(new_n5364_));
  INV_X1     g05300(.I(new_n4986_), .ZN(new_n5365_));
  OAI22_X1   g05301(.A1(new_n1729_), .A2(new_n3780_), .B1(new_n4745_), .B2(new_n3310_), .ZN(new_n5366_));
  NAND2_X1   g05302(.A1(new_n1862_), .A2(new_n3782_), .ZN(new_n5367_));
  AOI21_X1   g05303(.A1(new_n5366_), .A2(new_n5367_), .B(new_n3302_), .ZN(new_n5368_));
  NAND2_X1   g05304(.A1(new_n4842_), .A2(new_n5368_), .ZN(new_n5369_));
  XOR2_X1    g05305(.A1(new_n5369_), .A2(new_n84_), .Z(new_n5370_));
  NAND2_X1   g05306(.A1(new_n5370_), .A2(new_n5365_), .ZN(new_n5371_));
  AOI22_X1   g05307(.A1(new_n4766_), .A2(new_n5291_), .B1(new_n1813_), .B2(new_n3782_), .ZN(new_n5372_));
  AOI21_X1   g05308(.A1(new_n1862_), .A2(new_n3312_), .B(new_n5372_), .ZN(new_n5373_));
  NOR3_X1    g05309(.A1(new_n5373_), .A2(new_n4878_), .A3(new_n3302_), .ZN(new_n5374_));
  XOR2_X1    g05310(.A1(new_n5374_), .A2(new_n84_), .Z(new_n5375_));
  NAND2_X1   g05311(.A1(new_n1813_), .A2(new_n3312_), .ZN(new_n5376_));
  NAND2_X1   g05312(.A1(new_n4766_), .A2(new_n3782_), .ZN(new_n5377_));
  NAND4_X1   g05313(.A1(new_n4981_), .A2(new_n3301_), .A3(new_n5376_), .A4(new_n5377_), .ZN(new_n5378_));
  XOR2_X1    g05314(.A1(new_n5378_), .A2(\a[23] ), .Z(new_n5379_));
  NOR2_X1    g05315(.A1(new_n1999_), .A2(new_n3299_), .ZN(new_n5380_));
  NOR2_X1    g05316(.A1(new_n5380_), .A2(new_n84_), .ZN(new_n5381_));
  NAND3_X1   g05317(.A1(new_n5375_), .A2(new_n5379_), .A3(new_n5381_), .ZN(new_n5382_));
  INV_X1     g05318(.I(new_n5382_), .ZN(new_n5383_));
  NOR2_X1    g05319(.A1(new_n5370_), .A2(new_n5365_), .ZN(new_n5384_));
  OAI21_X1   g05320(.A1(new_n5383_), .A2(new_n5384_), .B(new_n5371_), .ZN(new_n5385_));
  XOR2_X1    g05321(.A1(new_n4985_), .A2(new_n4987_), .Z(new_n5386_));
  OAI22_X1   g05322(.A1(new_n1764_), .A2(new_n3780_), .B1(new_n1729_), .B2(new_n3306_), .ZN(new_n5387_));
  NAND2_X1   g05323(.A1(new_n1862_), .A2(new_n5291_), .ZN(new_n5388_));
  AOI21_X1   g05324(.A1(new_n5387_), .A2(new_n5388_), .B(new_n3302_), .ZN(new_n5389_));
  NAND2_X1   g05325(.A1(new_n4810_), .A2(new_n5389_), .ZN(new_n5390_));
  XOR2_X1    g05326(.A1(new_n5390_), .A2(\a[23] ), .Z(new_n5391_));
  NAND2_X1   g05327(.A1(new_n5391_), .A2(new_n5386_), .ZN(new_n5392_));
  NOR2_X1    g05328(.A1(new_n5391_), .A2(new_n5386_), .ZN(new_n5393_));
  AOI21_X1   g05329(.A1(new_n5385_), .A2(new_n5392_), .B(new_n5393_), .ZN(new_n5394_));
  NAND2_X1   g05330(.A1(new_n4985_), .A2(new_n4987_), .ZN(new_n5395_));
  XOR2_X1    g05331(.A1(new_n5395_), .A2(new_n4978_), .Z(new_n5396_));
  OAI22_X1   g05332(.A1(new_n1764_), .A2(new_n3306_), .B1(new_n1729_), .B2(new_n3310_), .ZN(new_n5397_));
  NAND2_X1   g05333(.A1(new_n1613_), .A2(new_n3312_), .ZN(new_n5398_));
  AOI21_X1   g05334(.A1(new_n5398_), .A2(new_n5397_), .B(new_n3302_), .ZN(new_n5399_));
  NAND2_X1   g05335(.A1(new_n4778_), .A2(new_n5399_), .ZN(new_n5400_));
  XOR2_X1    g05336(.A1(new_n5400_), .A2(new_n84_), .Z(new_n5401_));
  NOR2_X1    g05337(.A1(new_n5401_), .A2(new_n5396_), .ZN(new_n5402_));
  NAND2_X1   g05338(.A1(new_n5401_), .A2(new_n5396_), .ZN(new_n5403_));
  OAI21_X1   g05339(.A1(new_n5394_), .A2(new_n5402_), .B(new_n5403_), .ZN(new_n5404_));
  NOR2_X1    g05340(.A1(new_n4973_), .A2(new_n4967_), .ZN(new_n5405_));
  NOR2_X1    g05341(.A1(new_n5226_), .A2(new_n4968_), .ZN(new_n5406_));
  OAI21_X1   g05342(.A1(new_n5405_), .A2(new_n5406_), .B(new_n4989_), .ZN(new_n5407_));
  OAI21_X1   g05343(.A1(new_n5227_), .A2(new_n4990_), .B(new_n4988_), .ZN(new_n5408_));
  NAND2_X1   g05344(.A1(new_n5407_), .A2(new_n5408_), .ZN(new_n5409_));
  OAI22_X1   g05345(.A1(new_n1678_), .A2(new_n3780_), .B1(new_n1764_), .B2(new_n3310_), .ZN(new_n5410_));
  NAND2_X1   g05346(.A1(new_n1613_), .A2(new_n3782_), .ZN(new_n5411_));
  AOI21_X1   g05347(.A1(new_n5410_), .A2(new_n5411_), .B(new_n3302_), .ZN(new_n5412_));
  NAND2_X1   g05348(.A1(new_n4917_), .A2(new_n5412_), .ZN(new_n5413_));
  XOR2_X1    g05349(.A1(new_n5413_), .A2(new_n84_), .Z(new_n5414_));
  OAI21_X1   g05350(.A1(new_n5409_), .A2(new_n5414_), .B(new_n5404_), .ZN(new_n5415_));
  NAND2_X1   g05351(.A1(new_n5409_), .A2(new_n5414_), .ZN(new_n5416_));
  NAND2_X1   g05352(.A1(new_n5415_), .A2(new_n5416_), .ZN(new_n5417_));
  NAND2_X1   g05353(.A1(new_n5002_), .A2(new_n5230_), .ZN(new_n5418_));
  NAND2_X1   g05354(.A1(new_n5231_), .A2(new_n4997_), .ZN(new_n5419_));
  NAND2_X1   g05355(.A1(new_n5419_), .A2(new_n5418_), .ZN(new_n5420_));
  NAND2_X1   g05356(.A1(new_n5420_), .A2(new_n4991_), .ZN(new_n5421_));
  OAI21_X1   g05357(.A1(new_n5232_), .A2(new_n5004_), .B(new_n5229_), .ZN(new_n5422_));
  NAND2_X1   g05358(.A1(new_n5421_), .A2(new_n5422_), .ZN(new_n5423_));
  OAI22_X1   g05359(.A1(new_n1678_), .A2(new_n3306_), .B1(new_n2071_), .B2(new_n3780_), .ZN(new_n5424_));
  NAND2_X1   g05360(.A1(new_n1613_), .A2(new_n5291_), .ZN(new_n5425_));
  AOI21_X1   g05361(.A1(new_n5424_), .A2(new_n5425_), .B(new_n3302_), .ZN(new_n5426_));
  NAND2_X1   g05362(.A1(new_n5070_), .A2(new_n5426_), .ZN(new_n5427_));
  XOR2_X1    g05363(.A1(new_n5427_), .A2(\a[23] ), .Z(new_n5428_));
  NAND2_X1   g05364(.A1(new_n5428_), .A2(new_n5423_), .ZN(new_n5429_));
  NOR2_X1    g05365(.A1(new_n5428_), .A2(new_n5423_), .ZN(new_n5430_));
  AOI21_X1   g05366(.A1(new_n5417_), .A2(new_n5429_), .B(new_n5430_), .ZN(new_n5431_));
  XOR2_X1    g05367(.A1(new_n5236_), .A2(new_n5011_), .Z(new_n5432_));
  OAI21_X1   g05368(.A1(new_n5017_), .A2(new_n5238_), .B(new_n5005_), .ZN(new_n5433_));
  OAI21_X1   g05369(.A1(new_n5005_), .A2(new_n5432_), .B(new_n5433_), .ZN(new_n5434_));
  OAI22_X1   g05370(.A1(new_n2103_), .A2(new_n3780_), .B1(new_n1678_), .B2(new_n3310_), .ZN(new_n5435_));
  NAND2_X1   g05371(.A1(new_n2107_), .A2(new_n3782_), .ZN(new_n5436_));
  AOI21_X1   g05372(.A1(new_n5435_), .A2(new_n5436_), .B(new_n3302_), .ZN(new_n5437_));
  NAND2_X1   g05373(.A1(new_n4545_), .A2(new_n5437_), .ZN(new_n5438_));
  NOR2_X1    g05374(.A1(new_n5438_), .A2(\a[23] ), .ZN(new_n5439_));
  AOI21_X1   g05375(.A1(new_n4545_), .A2(new_n5437_), .B(new_n84_), .ZN(new_n5440_));
  NOR2_X1    g05376(.A1(new_n5439_), .A2(new_n5440_), .ZN(new_n5441_));
  NAND2_X1   g05377(.A1(new_n5434_), .A2(new_n5441_), .ZN(new_n5442_));
  INV_X1     g05378(.I(new_n5442_), .ZN(new_n5443_));
  NOR2_X1    g05379(.A1(new_n5432_), .A2(new_n5005_), .ZN(new_n5444_));
  INV_X1     g05380(.I(new_n5433_), .ZN(new_n5445_));
  NOR2_X1    g05381(.A1(new_n5445_), .A2(new_n5444_), .ZN(new_n5446_));
  INV_X1     g05382(.I(new_n5441_), .ZN(new_n5447_));
  NAND2_X1   g05383(.A1(new_n5447_), .A2(new_n5446_), .ZN(new_n5448_));
  OAI21_X1   g05384(.A1(new_n5431_), .A2(new_n5443_), .B(new_n5448_), .ZN(new_n5449_));
  OAI22_X1   g05385(.A1(new_n2103_), .A2(new_n3306_), .B1(new_n2158_), .B2(new_n3780_), .ZN(new_n5450_));
  NAND2_X1   g05386(.A1(new_n2107_), .A2(new_n5291_), .ZN(new_n5451_));
  AOI21_X1   g05387(.A1(new_n5450_), .A2(new_n5451_), .B(new_n3302_), .ZN(new_n5452_));
  NAND3_X1   g05388(.A1(new_n4959_), .A2(new_n84_), .A3(new_n5452_), .ZN(new_n5453_));
  INV_X1     g05389(.I(new_n5453_), .ZN(new_n5454_));
  AOI21_X1   g05390(.A1(new_n4959_), .A2(new_n5452_), .B(new_n84_), .ZN(new_n5455_));
  NOR2_X1    g05391(.A1(new_n5038_), .A2(new_n5241_), .ZN(new_n5456_));
  INV_X1     g05392(.I(new_n5456_), .ZN(new_n5457_));
  NAND2_X1   g05393(.A1(new_n5038_), .A2(new_n5241_), .ZN(new_n5458_));
  AOI21_X1   g05394(.A1(new_n5457_), .A2(new_n5458_), .B(new_n5239_), .ZN(new_n5459_));
  AOI21_X1   g05395(.A1(new_n5243_), .A2(new_n5044_), .B(new_n5019_), .ZN(new_n5460_));
  NOR4_X1    g05396(.A1(new_n5459_), .A2(new_n5460_), .A3(new_n5454_), .A4(new_n5455_), .ZN(new_n5461_));
  INV_X1     g05397(.I(new_n5455_), .ZN(new_n5462_));
  INV_X1     g05398(.I(new_n5458_), .ZN(new_n5463_));
  OAI21_X1   g05399(.A1(new_n5463_), .A2(new_n5456_), .B(new_n5019_), .ZN(new_n5464_));
  OAI21_X1   g05400(.A1(new_n5242_), .A2(new_n5045_), .B(new_n5239_), .ZN(new_n5465_));
  AOI22_X1   g05401(.A1(new_n5464_), .A2(new_n5465_), .B1(new_n5462_), .B2(new_n5453_), .ZN(new_n5466_));
  NOR2_X1    g05402(.A1(new_n5466_), .A2(new_n5461_), .ZN(new_n5467_));
  NOR2_X1    g05403(.A1(new_n5449_), .A2(new_n5467_), .ZN(new_n5468_));
  AOI21_X1   g05404(.A1(new_n5250_), .A2(new_n5079_), .B(new_n5046_), .ZN(new_n5469_));
  NAND2_X1   g05405(.A1(new_n5249_), .A2(new_n5066_), .ZN(new_n5470_));
  NAND2_X1   g05406(.A1(new_n5247_), .A2(new_n5077_), .ZN(new_n5471_));
  AOI21_X1   g05407(.A1(new_n5470_), .A2(new_n5471_), .B(new_n5244_), .ZN(new_n5472_));
  NOR3_X1    g05408(.A1(new_n5358_), .A2(new_n5469_), .A3(new_n5472_), .ZN(new_n5473_));
  NAND2_X1   g05409(.A1(new_n5357_), .A2(new_n5355_), .ZN(new_n5474_));
  AOI21_X1   g05410(.A1(new_n5359_), .A2(new_n5362_), .B(new_n5474_), .ZN(new_n5475_));
  NAND2_X1   g05411(.A1(new_n5462_), .A2(new_n5453_), .ZN(new_n5476_));
  NOR2_X1    g05412(.A1(new_n5459_), .A2(new_n5460_), .ZN(new_n5477_));
  NOR2_X1    g05413(.A1(new_n5477_), .A2(new_n5476_), .ZN(new_n5478_));
  INV_X1     g05414(.I(new_n5478_), .ZN(new_n5479_));
  OAI21_X1   g05415(.A1(new_n5473_), .A2(new_n5475_), .B(new_n5479_), .ZN(new_n5480_));
  OAI21_X1   g05416(.A1(new_n5480_), .A2(new_n5468_), .B(new_n5364_), .ZN(new_n5481_));
  OAI21_X1   g05417(.A1(new_n5108_), .A2(new_n5112_), .B(new_n5080_), .ZN(new_n5482_));
  NAND2_X1   g05418(.A1(new_n5339_), .A2(new_n5340_), .ZN(new_n5483_));
  NAND2_X1   g05419(.A1(new_n5483_), .A2(new_n5252_), .ZN(new_n5484_));
  INV_X1     g05420(.I(new_n5347_), .ZN(new_n5485_));
  AOI22_X1   g05421(.A1(new_n5484_), .A2(new_n5482_), .B1(new_n5345_), .B2(new_n5485_), .ZN(new_n5486_));
  OAI21_X1   g05422(.A1(new_n5481_), .A2(new_n5486_), .B(new_n5349_), .ZN(new_n5487_));
  NAND3_X1   g05423(.A1(new_n5487_), .A2(new_n5337_), .A3(new_n5330_), .ZN(new_n5488_));
  AOI22_X1   g05424(.A1(new_n5488_), .A2(new_n5306_), .B1(new_n5312_), .B2(new_n5319_), .ZN(new_n5489_));
  NAND2_X1   g05425(.A1(new_n5220_), .A2(new_n5278_), .ZN(new_n5490_));
  NAND2_X1   g05426(.A1(new_n5490_), .A2(new_n5270_), .ZN(new_n5491_));
  NOR2_X1    g05427(.A1(new_n5275_), .A2(new_n5218_), .ZN(new_n5492_));
  NOR2_X1    g05428(.A1(new_n5211_), .A2(new_n5277_), .ZN(new_n5493_));
  OAI21_X1   g05429(.A1(new_n5492_), .A2(new_n5493_), .B(new_n5190_), .ZN(new_n5494_));
  OAI22_X1   g05430(.A1(new_n2311_), .A2(new_n3780_), .B1(new_n4365_), .B2(new_n3310_), .ZN(new_n5495_));
  NAND2_X1   g05431(.A1(new_n2255_), .A2(new_n3782_), .ZN(new_n5496_));
  AOI21_X1   g05432(.A1(new_n5495_), .A2(new_n5496_), .B(new_n3302_), .ZN(new_n5497_));
  NAND3_X1   g05433(.A1(new_n4419_), .A2(new_n84_), .A3(new_n5497_), .ZN(new_n5498_));
  INV_X1     g05434(.I(new_n5498_), .ZN(new_n5499_));
  AOI21_X1   g05435(.A1(new_n4419_), .A2(new_n5497_), .B(new_n84_), .ZN(new_n5500_));
  NOR2_X1    g05436(.A1(new_n5499_), .A2(new_n5500_), .ZN(new_n5501_));
  NAND3_X1   g05437(.A1(new_n5501_), .A2(new_n5491_), .A3(new_n5494_), .ZN(new_n5502_));
  AOI21_X1   g05438(.A1(new_n5491_), .A2(new_n5494_), .B(new_n5501_), .ZN(new_n5503_));
  AOI21_X1   g05439(.A1(new_n5489_), .A2(new_n5502_), .B(new_n5503_), .ZN(new_n5504_));
  NOR3_X1    g05440(.A1(new_n5295_), .A2(new_n5299_), .A3(new_n5504_), .ZN(new_n5505_));
  XOR2_X1    g05441(.A1(new_n5293_), .A2(\a[23] ), .Z(new_n5506_));
  NAND3_X1   g05442(.A1(new_n5296_), .A2(new_n5297_), .A3(new_n5506_), .ZN(new_n5507_));
  XOR2_X1    g05443(.A1(new_n5293_), .A2(new_n84_), .Z(new_n5508_));
  OAI21_X1   g05444(.A1(new_n5288_), .A2(new_n5285_), .B(new_n5508_), .ZN(new_n5509_));
  NOR2_X1    g05445(.A1(new_n5314_), .A2(new_n5318_), .ZN(new_n5510_));
  NOR2_X1    g05446(.A1(new_n5306_), .A2(new_n5311_), .ZN(new_n5511_));
  OAI22_X1   g05447(.A1(new_n5331_), .A2(new_n5333_), .B1(new_n5334_), .B2(new_n5328_), .ZN(new_n5512_));
  NAND2_X1   g05448(.A1(new_n5330_), .A2(new_n5512_), .ZN(new_n5513_));
  INV_X1     g05449(.I(new_n5364_), .ZN(new_n5514_));
  AOI22_X1   g05450(.A1(new_n5415_), .A2(new_n5416_), .B1(new_n5423_), .B2(new_n5428_), .ZN(new_n5515_));
  OAI21_X1   g05451(.A1(new_n5515_), .A2(new_n5430_), .B(new_n5442_), .ZN(new_n5516_));
  NAND4_X1   g05452(.A1(new_n5464_), .A2(new_n5465_), .A3(new_n5462_), .A4(new_n5453_), .ZN(new_n5517_));
  OAI22_X1   g05453(.A1(new_n5459_), .A2(new_n5460_), .B1(new_n5454_), .B2(new_n5455_), .ZN(new_n5518_));
  NAND2_X1   g05454(.A1(new_n5518_), .A2(new_n5517_), .ZN(new_n5519_));
  NAND3_X1   g05455(.A1(new_n5519_), .A2(new_n5516_), .A3(new_n5448_), .ZN(new_n5520_));
  NAND3_X1   g05456(.A1(new_n5474_), .A2(new_n5359_), .A3(new_n5362_), .ZN(new_n5521_));
  NAND2_X1   g05457(.A1(new_n5363_), .A2(new_n5358_), .ZN(new_n5522_));
  AOI21_X1   g05458(.A1(new_n5522_), .A2(new_n5521_), .B(new_n5478_), .ZN(new_n5523_));
  AOI21_X1   g05459(.A1(new_n5523_), .A2(new_n5520_), .B(new_n5514_), .ZN(new_n5524_));
  NOR2_X1    g05460(.A1(new_n5486_), .A2(new_n5348_), .ZN(new_n5525_));
  AOI21_X1   g05461(.A1(new_n5524_), .A2(new_n5525_), .B(new_n5348_), .ZN(new_n5526_));
  NOR3_X1    g05462(.A1(new_n5526_), .A2(new_n5335_), .A3(new_n5513_), .ZN(new_n5527_));
  OAI22_X1   g05463(.A1(new_n5527_), .A2(new_n5314_), .B1(new_n5511_), .B2(new_n5510_), .ZN(new_n5528_));
  INV_X1     g05464(.I(new_n5502_), .ZN(new_n5529_));
  NAND2_X1   g05465(.A1(new_n5491_), .A2(new_n5494_), .ZN(new_n5530_));
  INV_X1     g05466(.I(new_n5500_), .ZN(new_n5531_));
  NAND2_X1   g05467(.A1(new_n5531_), .A2(new_n5498_), .ZN(new_n5532_));
  NAND2_X1   g05468(.A1(new_n5530_), .A2(new_n5532_), .ZN(new_n5533_));
  OAI21_X1   g05469(.A1(new_n5528_), .A2(new_n5529_), .B(new_n5533_), .ZN(new_n5534_));
  AOI21_X1   g05470(.A1(new_n5509_), .A2(new_n5507_), .B(new_n5534_), .ZN(new_n5535_));
  INV_X1     g05471(.I(new_n3827_), .ZN(new_n5536_));
  OAI22_X1   g05472(.A1(new_n1409_), .A2(new_n3775_), .B1(new_n1333_), .B2(new_n4097_), .ZN(new_n5537_));
  NAND2_X1   g05473(.A1(new_n2359_), .A2(new_n3770_), .ZN(new_n5538_));
  AOI21_X1   g05474(.A1(new_n5537_), .A2(new_n5538_), .B(new_n4095_), .ZN(new_n5539_));
  OAI21_X1   g05475(.A1(new_n5536_), .A2(new_n3823_), .B(new_n5539_), .ZN(new_n5540_));
  XOR2_X1    g05476(.A1(new_n5540_), .A2(\a[20] ), .Z(new_n5541_));
  OAI21_X1   g05477(.A1(new_n5505_), .A2(new_n5535_), .B(new_n5541_), .ZN(new_n5542_));
  NOR2_X1    g05478(.A1(new_n5481_), .A2(new_n5525_), .ZN(new_n5543_));
  NOR3_X1    g05479(.A1(new_n5524_), .A2(new_n5348_), .A3(new_n5486_), .ZN(new_n5544_));
  OAI22_X1   g05480(.A1(new_n2311_), .A2(new_n4097_), .B1(new_n4365_), .B2(new_n3769_), .ZN(new_n5545_));
  NAND2_X1   g05481(.A1(new_n2255_), .A2(new_n3776_), .ZN(new_n5546_));
  AOI21_X1   g05482(.A1(new_n5545_), .A2(new_n5546_), .B(new_n4095_), .ZN(new_n5547_));
  NAND3_X1   g05483(.A1(new_n4419_), .A2(new_n3035_), .A3(new_n5547_), .ZN(new_n5548_));
  INV_X1     g05484(.I(new_n5548_), .ZN(new_n5549_));
  AOI21_X1   g05485(.A1(new_n4419_), .A2(new_n5547_), .B(new_n3035_), .ZN(new_n5550_));
  NOR2_X1    g05486(.A1(new_n5549_), .A2(new_n5550_), .ZN(new_n5551_));
  NOR3_X1    g05487(.A1(new_n5551_), .A2(new_n5543_), .A3(new_n5544_), .ZN(new_n5552_));
  NOR2_X1    g05488(.A1(new_n5487_), .A2(new_n5513_), .ZN(new_n5553_));
  NOR2_X1    g05489(.A1(new_n5526_), .A2(new_n5337_), .ZN(new_n5554_));
  NOR2_X1    g05490(.A1(new_n3909_), .A2(new_n3913_), .ZN(new_n5555_));
  OAI22_X1   g05491(.A1(new_n2251_), .A2(new_n3769_), .B1(new_n2351_), .B2(new_n4097_), .ZN(new_n5556_));
  NAND2_X1   g05492(.A1(new_n2310_), .A2(new_n3776_), .ZN(new_n5557_));
  AOI21_X1   g05493(.A1(new_n5557_), .A2(new_n5556_), .B(new_n4095_), .ZN(new_n5558_));
  OAI21_X1   g05494(.A1(new_n5555_), .A2(new_n3911_), .B(new_n5558_), .ZN(new_n5559_));
  NOR2_X1    g05495(.A1(new_n5559_), .A2(\a[20] ), .ZN(new_n5560_));
  AOI21_X1   g05496(.A1(new_n3914_), .A2(new_n5558_), .B(new_n3035_), .ZN(new_n5561_));
  NOR2_X1    g05497(.A1(new_n5561_), .A2(new_n5560_), .ZN(new_n5562_));
  OAI21_X1   g05498(.A1(new_n5554_), .A2(new_n5553_), .B(new_n5562_), .ZN(new_n5563_));
  NOR3_X1    g05499(.A1(new_n5554_), .A2(new_n5553_), .A3(new_n5562_), .ZN(new_n5564_));
  AOI21_X1   g05500(.A1(new_n5563_), .A2(new_n5552_), .B(new_n5564_), .ZN(new_n5565_));
  NOR2_X1    g05501(.A1(new_n5527_), .A2(new_n5306_), .ZN(new_n5566_));
  NOR2_X1    g05502(.A1(new_n5488_), .A2(new_n5314_), .ZN(new_n5567_));
  OAI21_X1   g05503(.A1(new_n5566_), .A2(new_n5567_), .B(new_n5311_), .ZN(new_n5568_));
  NAND2_X1   g05504(.A1(new_n5488_), .A2(new_n5314_), .ZN(new_n5569_));
  NAND4_X1   g05505(.A1(new_n5487_), .A2(new_n5306_), .A3(new_n5337_), .A4(new_n5330_), .ZN(new_n5570_));
  NAND3_X1   g05506(.A1(new_n5569_), .A2(new_n5318_), .A3(new_n5570_), .ZN(new_n5571_));
  OAI22_X1   g05507(.A1(new_n1453_), .A2(new_n4097_), .B1(new_n2351_), .B2(new_n3775_), .ZN(new_n5572_));
  NAND2_X1   g05508(.A1(new_n2310_), .A2(new_n3770_), .ZN(new_n5573_));
  AOI21_X1   g05509(.A1(new_n5573_), .A2(new_n5572_), .B(new_n4095_), .ZN(new_n5574_));
  NAND2_X1   g05510(.A1(new_n4231_), .A2(new_n5574_), .ZN(new_n5575_));
  XOR2_X1    g05511(.A1(new_n5575_), .A2(new_n3035_), .Z(new_n5576_));
  AOI21_X1   g05512(.A1(new_n5568_), .A2(new_n5571_), .B(new_n5576_), .ZN(new_n5577_));
  NOR2_X1    g05513(.A1(new_n5577_), .A2(new_n5565_), .ZN(new_n5578_));
  AOI21_X1   g05514(.A1(new_n5569_), .A2(new_n5570_), .B(new_n5318_), .ZN(new_n5579_));
  NOR3_X1    g05515(.A1(new_n5566_), .A2(new_n5567_), .A3(new_n5311_), .ZN(new_n5580_));
  XOR2_X1    g05516(.A1(new_n5575_), .A2(\a[20] ), .Z(new_n5581_));
  NOR3_X1    g05517(.A1(new_n5580_), .A2(new_n5579_), .A3(new_n5581_), .ZN(new_n5582_));
  NAND2_X1   g05518(.A1(new_n5530_), .A2(new_n5501_), .ZN(new_n5583_));
  NAND3_X1   g05519(.A1(new_n5532_), .A2(new_n5491_), .A3(new_n5494_), .ZN(new_n5584_));
  AOI21_X1   g05520(.A1(new_n5583_), .A2(new_n5584_), .B(new_n5528_), .ZN(new_n5585_));
  AOI21_X1   g05521(.A1(new_n5502_), .A2(new_n5533_), .B(new_n5489_), .ZN(new_n5586_));
  NOR2_X1    g05522(.A1(new_n5585_), .A2(new_n5586_), .ZN(new_n5587_));
  OAI22_X1   g05523(.A1(new_n1409_), .A2(new_n4097_), .B1(new_n2351_), .B2(new_n3769_), .ZN(new_n5588_));
  NAND2_X1   g05524(.A1(new_n2359_), .A2(new_n3776_), .ZN(new_n5589_));
  AOI21_X1   g05525(.A1(new_n5588_), .A2(new_n5589_), .B(new_n4095_), .ZN(new_n5590_));
  NAND3_X1   g05526(.A1(new_n3904_), .A2(new_n3035_), .A3(new_n5590_), .ZN(new_n5591_));
  NAND2_X1   g05527(.A1(new_n3904_), .A2(new_n5590_), .ZN(new_n5592_));
  NAND2_X1   g05528(.A1(new_n5592_), .A2(\a[20] ), .ZN(new_n5593_));
  NAND2_X1   g05529(.A1(new_n5593_), .A2(new_n5591_), .ZN(new_n5594_));
  OAI22_X1   g05530(.A1(new_n5578_), .A2(new_n5582_), .B1(new_n5587_), .B2(new_n5594_), .ZN(new_n5595_));
  NAND2_X1   g05531(.A1(new_n5587_), .A2(new_n5594_), .ZN(new_n5596_));
  NAND3_X1   g05532(.A1(new_n5509_), .A2(new_n5507_), .A3(new_n5534_), .ZN(new_n5597_));
  OAI21_X1   g05533(.A1(new_n5295_), .A2(new_n5299_), .B(new_n5504_), .ZN(new_n5598_));
  XOR2_X1    g05534(.A1(new_n5540_), .A2(new_n3035_), .Z(new_n5599_));
  NAND3_X1   g05535(.A1(new_n5598_), .A2(new_n5597_), .A3(new_n5599_), .ZN(new_n5600_));
  NAND4_X1   g05536(.A1(new_n5595_), .A2(new_n5542_), .A3(new_n5600_), .A4(new_n5596_), .ZN(new_n5601_));
  AOI21_X1   g05537(.A1(new_n5598_), .A2(new_n5597_), .B(new_n5599_), .ZN(new_n5602_));
  NOR2_X1    g05538(.A1(new_n5544_), .A2(new_n5543_), .ZN(new_n5603_));
  INV_X1     g05539(.I(new_n5550_), .ZN(new_n5604_));
  NAND2_X1   g05540(.A1(new_n5604_), .A2(new_n5548_), .ZN(new_n5605_));
  NAND2_X1   g05541(.A1(new_n5603_), .A2(new_n5605_), .ZN(new_n5606_));
  INV_X1     g05542(.I(new_n5563_), .ZN(new_n5607_));
  NOR2_X1    g05543(.A1(new_n5554_), .A2(new_n5553_), .ZN(new_n5608_));
  INV_X1     g05544(.I(new_n5562_), .ZN(new_n5609_));
  NAND2_X1   g05545(.A1(new_n5608_), .A2(new_n5609_), .ZN(new_n5610_));
  OAI21_X1   g05546(.A1(new_n5606_), .A2(new_n5607_), .B(new_n5610_), .ZN(new_n5611_));
  OAI21_X1   g05547(.A1(new_n5580_), .A2(new_n5579_), .B(new_n5581_), .ZN(new_n5612_));
  NAND2_X1   g05548(.A1(new_n5612_), .A2(new_n5611_), .ZN(new_n5613_));
  NAND3_X1   g05549(.A1(new_n5568_), .A2(new_n5571_), .A3(new_n5576_), .ZN(new_n5614_));
  NAND2_X1   g05550(.A1(new_n5583_), .A2(new_n5584_), .ZN(new_n5615_));
  NAND2_X1   g05551(.A1(new_n5615_), .A2(new_n5489_), .ZN(new_n5616_));
  OAI21_X1   g05552(.A1(new_n5529_), .A2(new_n5503_), .B(new_n5528_), .ZN(new_n5617_));
  AOI21_X1   g05553(.A1(new_n5617_), .A2(new_n5616_), .B(new_n5594_), .ZN(new_n5618_));
  AOI21_X1   g05554(.A1(new_n5613_), .A2(new_n5614_), .B(new_n5618_), .ZN(new_n5619_));
  NAND2_X1   g05555(.A1(new_n5617_), .A2(new_n5616_), .ZN(new_n5620_));
  INV_X1     g05556(.I(new_n5594_), .ZN(new_n5621_));
  NOR2_X1    g05557(.A1(new_n5620_), .A2(new_n5621_), .ZN(new_n5622_));
  NOR3_X1    g05558(.A1(new_n5505_), .A2(new_n5535_), .A3(new_n5541_), .ZN(new_n5623_));
  OAI22_X1   g05559(.A1(new_n5619_), .A2(new_n5622_), .B1(new_n5623_), .B2(new_n5602_), .ZN(new_n5624_));
  AOI21_X1   g05560(.A1(new_n2411_), .A2(new_n2414_), .B(new_n3399_), .ZN(new_n5625_));
  NOR2_X1    g05561(.A1(new_n3398_), .A2(new_n3402_), .ZN(new_n5626_));
  OAI21_X1   g05562(.A1(new_n2408_), .A2(new_n4297_), .B(new_n4295_), .ZN(new_n5627_));
  OAI22_X1   g05563(.A1(new_n2367_), .A2(new_n4291_), .B1(new_n2451_), .B2(new_n4470_), .ZN(new_n5628_));
  NOR2_X1    g05564(.A1(new_n5628_), .A2(new_n5627_), .ZN(new_n5629_));
  OAI21_X1   g05565(.A1(new_n5626_), .A2(new_n5625_), .B(new_n5629_), .ZN(new_n5630_));
  XOR2_X1    g05566(.A1(new_n5630_), .A2(\a[17] ), .Z(new_n5631_));
  NAND3_X1   g05567(.A1(new_n5624_), .A2(new_n5601_), .A3(new_n5631_), .ZN(new_n5632_));
  NOR3_X1    g05568(.A1(new_n3652_), .A2(new_n2367_), .A3(new_n3649_), .ZN(new_n5633_));
  AOI21_X1   g05569(.A1(new_n3650_), .A2(new_n3645_), .B(new_n1241_), .ZN(new_n5634_));
  OAI22_X1   g05570(.A1(new_n1409_), .A2(new_n4291_), .B1(new_n2367_), .B2(new_n4470_), .ZN(new_n5635_));
  NAND2_X1   g05571(.A1(new_n1334_), .A2(new_n4298_), .ZN(new_n5636_));
  AOI21_X1   g05572(.A1(new_n5635_), .A2(new_n5636_), .B(new_n4468_), .ZN(new_n5637_));
  OAI21_X1   g05573(.A1(new_n5634_), .A2(new_n5633_), .B(new_n5637_), .ZN(new_n5638_));
  NOR2_X1    g05574(.A1(new_n5638_), .A2(\a[17] ), .ZN(new_n5639_));
  AOI21_X1   g05575(.A1(new_n3654_), .A2(new_n5637_), .B(new_n3372_), .ZN(new_n5640_));
  NOR2_X1    g05576(.A1(new_n5639_), .A2(new_n5640_), .ZN(new_n5641_));
  AOI21_X1   g05577(.A1(new_n5612_), .A2(new_n5614_), .B(new_n5565_), .ZN(new_n5642_));
  NAND3_X1   g05578(.A1(new_n5568_), .A2(new_n5571_), .A3(new_n5581_), .ZN(new_n5643_));
  OAI21_X1   g05579(.A1(new_n5580_), .A2(new_n5579_), .B(new_n5576_), .ZN(new_n5644_));
  AOI21_X1   g05580(.A1(new_n5644_), .A2(new_n5643_), .B(new_n5611_), .ZN(new_n5645_));
  NOR3_X1    g05581(.A1(new_n5645_), .A2(new_n5642_), .A3(new_n5641_), .ZN(new_n5646_));
  INV_X1     g05582(.I(new_n5641_), .ZN(new_n5647_));
  OAI21_X1   g05583(.A1(new_n5577_), .A2(new_n5582_), .B(new_n5611_), .ZN(new_n5648_));
  NOR3_X1    g05584(.A1(new_n5580_), .A2(new_n5579_), .A3(new_n5576_), .ZN(new_n5649_));
  AOI21_X1   g05585(.A1(new_n5568_), .A2(new_n5571_), .B(new_n5581_), .ZN(new_n5650_));
  OAI21_X1   g05586(.A1(new_n5650_), .A2(new_n5649_), .B(new_n5565_), .ZN(new_n5651_));
  AOI21_X1   g05587(.A1(new_n5648_), .A2(new_n5651_), .B(new_n5647_), .ZN(new_n5652_));
  NOR2_X1    g05588(.A1(new_n5652_), .A2(new_n5646_), .ZN(new_n5653_));
  NAND2_X1   g05589(.A1(new_n5648_), .A2(new_n5651_), .ZN(new_n5654_));
  NAND2_X1   g05590(.A1(new_n5654_), .A2(new_n5641_), .ZN(new_n5655_));
  OAI21_X1   g05591(.A1(new_n5607_), .A2(new_n5564_), .B(new_n5552_), .ZN(new_n5656_));
  NOR3_X1    g05592(.A1(new_n5609_), .A2(new_n5554_), .A3(new_n5553_), .ZN(new_n5657_));
  NOR2_X1    g05593(.A1(new_n5608_), .A2(new_n5562_), .ZN(new_n5658_));
  OAI21_X1   g05594(.A1(new_n5658_), .A2(new_n5657_), .B(new_n5606_), .ZN(new_n5659_));
  OAI22_X1   g05595(.A1(new_n1409_), .A2(new_n4297_), .B1(new_n1333_), .B2(new_n4470_), .ZN(new_n5660_));
  NAND2_X1   g05596(.A1(new_n2359_), .A2(new_n4292_), .ZN(new_n5661_));
  AOI21_X1   g05597(.A1(new_n5660_), .A2(new_n5661_), .B(new_n4468_), .ZN(new_n5662_));
  NAND3_X1   g05598(.A1(new_n3828_), .A2(new_n3372_), .A3(new_n5662_), .ZN(new_n5663_));
  OAI21_X1   g05599(.A1(new_n5536_), .A2(new_n3823_), .B(new_n5662_), .ZN(new_n5664_));
  NAND2_X1   g05600(.A1(new_n5664_), .A2(\a[17] ), .ZN(new_n5665_));
  NAND4_X1   g05601(.A1(new_n5659_), .A2(new_n5656_), .A3(new_n5663_), .A4(new_n5665_), .ZN(new_n5666_));
  AOI21_X1   g05602(.A1(new_n5610_), .A2(new_n5563_), .B(new_n5606_), .ZN(new_n5667_));
  NAND2_X1   g05603(.A1(new_n5608_), .A2(new_n5562_), .ZN(new_n5668_));
  OAI21_X1   g05604(.A1(new_n5553_), .A2(new_n5554_), .B(new_n5609_), .ZN(new_n5669_));
  AOI21_X1   g05605(.A1(new_n5668_), .A2(new_n5669_), .B(new_n5552_), .ZN(new_n5670_));
  INV_X1     g05606(.I(new_n5663_), .ZN(new_n5671_));
  AOI21_X1   g05607(.A1(new_n3828_), .A2(new_n5662_), .B(new_n3372_), .ZN(new_n5672_));
  NOR4_X1    g05608(.A1(new_n5670_), .A2(new_n5671_), .A3(new_n5667_), .A4(new_n5672_), .ZN(new_n5673_));
  AOI22_X1   g05609(.A1(new_n5659_), .A2(new_n5656_), .B1(new_n5663_), .B2(new_n5665_), .ZN(new_n5674_));
  NOR2_X1    g05610(.A1(new_n5673_), .A2(new_n5674_), .ZN(new_n5675_));
  OAI21_X1   g05611(.A1(new_n5543_), .A2(new_n5544_), .B(new_n5551_), .ZN(new_n5676_));
  NOR2_X1    g05612(.A1(new_n1453_), .A2(new_n4297_), .ZN(new_n5677_));
  NOR2_X1    g05613(.A1(new_n1409_), .A2(new_n4470_), .ZN(new_n5678_));
  NOR2_X1    g05614(.A1(new_n2351_), .A2(new_n4291_), .ZN(new_n5679_));
  NOR4_X1    g05615(.A1(new_n5678_), .A2(new_n4468_), .A3(new_n5677_), .A4(new_n5679_), .ZN(new_n5680_));
  NAND2_X1   g05616(.A1(new_n3904_), .A2(new_n5680_), .ZN(new_n5681_));
  XOR2_X1    g05617(.A1(new_n5681_), .A2(new_n3372_), .Z(new_n5682_));
  NAND3_X1   g05618(.A1(new_n5682_), .A2(new_n5606_), .A3(new_n5676_), .ZN(new_n5683_));
  INV_X1     g05619(.I(new_n4227_), .ZN(new_n5684_));
  OAI22_X1   g05620(.A1(new_n1453_), .A2(new_n4470_), .B1(new_n2351_), .B2(new_n4297_), .ZN(new_n5685_));
  NAND2_X1   g05621(.A1(new_n2310_), .A2(new_n4292_), .ZN(new_n5686_));
  AOI21_X1   g05622(.A1(new_n5686_), .A2(new_n5685_), .B(new_n4468_), .ZN(new_n5687_));
  OAI21_X1   g05623(.A1(new_n5684_), .A2(new_n4229_), .B(new_n5687_), .ZN(new_n5688_));
  XOR2_X1    g05624(.A1(new_n5688_), .A2(\a[17] ), .Z(new_n5689_));
  INV_X1     g05625(.I(new_n5363_), .ZN(new_n5690_));
  AOI21_X1   g05626(.A1(new_n5520_), .A2(new_n5479_), .B(new_n5474_), .ZN(new_n5691_));
  OAI21_X1   g05627(.A1(new_n5449_), .A2(new_n5467_), .B(new_n5479_), .ZN(new_n5692_));
  NOR2_X1    g05628(.A1(new_n5692_), .A2(new_n5358_), .ZN(new_n5693_));
  OAI21_X1   g05629(.A1(new_n5693_), .A2(new_n5691_), .B(new_n5690_), .ZN(new_n5694_));
  NAND2_X1   g05630(.A1(new_n5692_), .A2(new_n5358_), .ZN(new_n5695_));
  NAND3_X1   g05631(.A1(new_n5520_), .A2(new_n5474_), .A3(new_n5479_), .ZN(new_n5696_));
  NAND3_X1   g05632(.A1(new_n5695_), .A2(new_n5696_), .A3(new_n5363_), .ZN(new_n5697_));
  NAND2_X1   g05633(.A1(new_n5694_), .A2(new_n5697_), .ZN(new_n5698_));
  NOR2_X1    g05634(.A1(new_n5449_), .A2(new_n5519_), .ZN(new_n5699_));
  AOI21_X1   g05635(.A1(new_n5516_), .A2(new_n5448_), .B(new_n5467_), .ZN(new_n5700_));
  INV_X1     g05636(.I(new_n4359_), .ZN(new_n5701_));
  NOR3_X1    g05637(.A1(new_n2206_), .A2(new_n2207_), .A3(new_n4360_), .ZN(new_n5702_));
  OAI22_X1   g05638(.A1(new_n4365_), .A2(new_n4097_), .B1(new_n2198_), .B2(new_n3769_), .ZN(new_n5703_));
  NAND2_X1   g05639(.A1(new_n1504_), .A2(new_n3776_), .ZN(new_n5704_));
  AOI21_X1   g05640(.A1(new_n5703_), .A2(new_n5704_), .B(new_n4095_), .ZN(new_n5705_));
  OAI21_X1   g05641(.A1(new_n5701_), .A2(new_n5702_), .B(new_n5705_), .ZN(new_n5706_));
  XOR2_X1    g05642(.A1(new_n5706_), .A2(\a[20] ), .Z(new_n5707_));
  OAI21_X1   g05643(.A1(new_n5699_), .A2(new_n5700_), .B(new_n5707_), .ZN(new_n5708_));
  NAND3_X1   g05644(.A1(new_n5467_), .A2(new_n5516_), .A3(new_n5448_), .ZN(new_n5709_));
  NAND2_X1   g05645(.A1(new_n5449_), .A2(new_n5519_), .ZN(new_n5710_));
  NAND3_X1   g05646(.A1(new_n4363_), .A2(new_n3035_), .A3(new_n5705_), .ZN(new_n5711_));
  NAND2_X1   g05647(.A1(new_n5706_), .A2(\a[20] ), .ZN(new_n5712_));
  NAND2_X1   g05648(.A1(new_n5712_), .A2(new_n5711_), .ZN(new_n5713_));
  NAND3_X1   g05649(.A1(new_n5710_), .A2(new_n5713_), .A3(new_n5709_), .ZN(new_n5714_));
  AOI21_X1   g05650(.A1(new_n5442_), .A2(new_n5448_), .B(new_n5431_), .ZN(new_n5715_));
  NOR2_X1    g05651(.A1(new_n5447_), .A2(new_n5434_), .ZN(new_n5716_));
  NOR2_X1    g05652(.A1(new_n5446_), .A2(new_n5441_), .ZN(new_n5717_));
  OAI21_X1   g05653(.A1(new_n5716_), .A2(new_n5717_), .B(new_n5431_), .ZN(new_n5718_));
  INV_X1     g05654(.I(new_n5718_), .ZN(new_n5719_));
  OAI22_X1   g05655(.A1(new_n2158_), .A2(new_n3769_), .B1(new_n2198_), .B2(new_n3775_), .ZN(new_n5720_));
  NAND2_X1   g05656(.A1(new_n1504_), .A2(new_n4096_), .ZN(new_n5721_));
  AOI21_X1   g05657(.A1(new_n5721_), .A2(new_n5720_), .B(new_n4095_), .ZN(new_n5722_));
  NAND3_X1   g05658(.A1(new_n4620_), .A2(new_n3035_), .A3(new_n5722_), .ZN(new_n5723_));
  INV_X1     g05659(.I(new_n5723_), .ZN(new_n5724_));
  AOI21_X1   g05660(.A1(new_n4620_), .A2(new_n5722_), .B(new_n3035_), .ZN(new_n5725_));
  NOR2_X1    g05661(.A1(new_n5724_), .A2(new_n5725_), .ZN(new_n5726_));
  INV_X1     g05662(.I(new_n5726_), .ZN(new_n5727_));
  OAI21_X1   g05663(.A1(new_n5719_), .A2(new_n5715_), .B(new_n5727_), .ZN(new_n5728_));
  NAND3_X1   g05664(.A1(new_n5708_), .A2(new_n5728_), .A3(new_n5714_), .ZN(new_n5729_));
  NOR2_X1    g05665(.A1(new_n4648_), .A2(new_n2251_), .ZN(new_n5730_));
  AOI21_X1   g05666(.A1(new_n4645_), .A2(new_n4358_), .B(new_n2255_), .ZN(new_n5731_));
  OAI22_X1   g05667(.A1(new_n2251_), .A2(new_n4097_), .B1(new_n4365_), .B2(new_n3775_), .ZN(new_n5732_));
  NAND2_X1   g05668(.A1(new_n1504_), .A2(new_n3770_), .ZN(new_n5733_));
  AOI21_X1   g05669(.A1(new_n5732_), .A2(new_n5733_), .B(new_n4095_), .ZN(new_n5734_));
  OAI21_X1   g05670(.A1(new_n5730_), .A2(new_n5731_), .B(new_n5734_), .ZN(new_n5735_));
  XOR2_X1    g05671(.A1(new_n5735_), .A2(\a[20] ), .Z(new_n5736_));
  NAND2_X1   g05672(.A1(new_n5729_), .A2(new_n5736_), .ZN(new_n5737_));
  AOI21_X1   g05673(.A1(new_n5710_), .A2(new_n5709_), .B(new_n5713_), .ZN(new_n5738_));
  NOR3_X1    g05674(.A1(new_n5707_), .A2(new_n5699_), .A3(new_n5700_), .ZN(new_n5739_));
  INV_X1     g05675(.I(new_n5715_), .ZN(new_n5740_));
  AOI21_X1   g05676(.A1(new_n5740_), .A2(new_n5718_), .B(new_n5726_), .ZN(new_n5741_));
  NOR3_X1    g05677(.A1(new_n5739_), .A2(new_n5738_), .A3(new_n5741_), .ZN(new_n5742_));
  XOR2_X1    g05678(.A1(new_n5735_), .A2(new_n3035_), .Z(new_n5743_));
  NAND2_X1   g05679(.A1(new_n5742_), .A2(new_n5743_), .ZN(new_n5744_));
  AOI21_X1   g05680(.A1(new_n5737_), .A2(new_n5744_), .B(new_n5698_), .ZN(new_n5745_));
  AOI21_X1   g05681(.A1(new_n5695_), .A2(new_n5696_), .B(new_n5363_), .ZN(new_n5746_));
  NOR3_X1    g05682(.A1(new_n5693_), .A2(new_n5691_), .A3(new_n5690_), .ZN(new_n5747_));
  NOR2_X1    g05683(.A1(new_n5747_), .A2(new_n5746_), .ZN(new_n5748_));
  NOR2_X1    g05684(.A1(new_n5742_), .A2(new_n5743_), .ZN(new_n5749_));
  NOR2_X1    g05685(.A1(new_n5729_), .A2(new_n5736_), .ZN(new_n5750_));
  NOR3_X1    g05686(.A1(new_n5750_), .A2(new_n5749_), .A3(new_n5748_), .ZN(new_n5751_));
  OAI21_X1   g05687(.A1(new_n5745_), .A2(new_n5751_), .B(new_n5689_), .ZN(new_n5752_));
  OAI22_X1   g05688(.A1(new_n2251_), .A2(new_n4291_), .B1(new_n2351_), .B2(new_n4470_), .ZN(new_n5753_));
  NAND2_X1   g05689(.A1(new_n2310_), .A2(new_n4298_), .ZN(new_n5754_));
  AOI21_X1   g05690(.A1(new_n5754_), .A2(new_n5753_), .B(new_n4468_), .ZN(new_n5755_));
  NAND3_X1   g05691(.A1(new_n3914_), .A2(new_n3372_), .A3(new_n5755_), .ZN(new_n5756_));
  OAI21_X1   g05692(.A1(new_n5555_), .A2(new_n3911_), .B(new_n5755_), .ZN(new_n5757_));
  NAND2_X1   g05693(.A1(new_n5757_), .A2(\a[17] ), .ZN(new_n5758_));
  NAND2_X1   g05694(.A1(new_n5756_), .A2(new_n5758_), .ZN(new_n5759_));
  NOR3_X1    g05695(.A1(new_n5728_), .A2(new_n5739_), .A3(new_n5738_), .ZN(new_n5760_));
  AOI21_X1   g05696(.A1(new_n5708_), .A2(new_n5714_), .B(new_n5741_), .ZN(new_n5761_));
  NOR3_X1    g05697(.A1(new_n5759_), .A2(new_n5760_), .A3(new_n5761_), .ZN(new_n5762_));
  XOR2_X1    g05698(.A1(new_n5757_), .A2(\a[17] ), .Z(new_n5763_));
  INV_X1     g05699(.I(new_n5760_), .ZN(new_n5764_));
  INV_X1     g05700(.I(new_n5761_), .ZN(new_n5765_));
  AOI21_X1   g05701(.A1(new_n5764_), .A2(new_n5765_), .B(new_n5763_), .ZN(new_n5766_));
  INV_X1     g05702(.I(new_n5380_), .ZN(new_n5767_));
  OAI22_X1   g05703(.A1(new_n1729_), .A2(new_n4097_), .B1(new_n4745_), .B2(new_n3769_), .ZN(new_n5768_));
  NAND2_X1   g05704(.A1(new_n1862_), .A2(new_n3776_), .ZN(new_n5769_));
  AOI21_X1   g05705(.A1(new_n5768_), .A2(new_n5769_), .B(new_n4095_), .ZN(new_n5770_));
  NAND2_X1   g05706(.A1(new_n4842_), .A2(new_n5770_), .ZN(new_n5771_));
  XOR2_X1    g05707(.A1(new_n5771_), .A2(new_n3035_), .Z(new_n5772_));
  NAND2_X1   g05708(.A1(new_n5772_), .A2(new_n5767_), .ZN(new_n5773_));
  AOI22_X1   g05709(.A1(new_n4766_), .A2(new_n3770_), .B1(new_n1813_), .B2(new_n3776_), .ZN(new_n5774_));
  AOI21_X1   g05710(.A1(new_n1862_), .A2(new_n4096_), .B(new_n5774_), .ZN(new_n5775_));
  NOR3_X1    g05711(.A1(new_n5775_), .A2(new_n4878_), .A3(new_n4095_), .ZN(new_n5776_));
  XOR2_X1    g05712(.A1(new_n5776_), .A2(new_n3035_), .Z(new_n5777_));
  NAND2_X1   g05713(.A1(new_n1813_), .A2(new_n4096_), .ZN(new_n5778_));
  NAND2_X1   g05714(.A1(new_n4766_), .A2(new_n3776_), .ZN(new_n5779_));
  NAND4_X1   g05715(.A1(new_n4981_), .A2(new_n3773_), .A3(new_n5778_), .A4(new_n5779_), .ZN(new_n5780_));
  XOR2_X1    g05716(.A1(new_n5780_), .A2(\a[20] ), .Z(new_n5781_));
  NOR2_X1    g05717(.A1(new_n1999_), .A2(new_n3762_), .ZN(new_n5782_));
  NOR2_X1    g05718(.A1(new_n5782_), .A2(new_n3035_), .ZN(new_n5783_));
  NAND3_X1   g05719(.A1(new_n5777_), .A2(new_n5781_), .A3(new_n5783_), .ZN(new_n5784_));
  XOR2_X1    g05720(.A1(new_n5771_), .A2(\a[20] ), .Z(new_n5785_));
  NAND2_X1   g05721(.A1(new_n5785_), .A2(new_n5380_), .ZN(new_n5786_));
  NAND2_X1   g05722(.A1(new_n5786_), .A2(new_n5784_), .ZN(new_n5787_));
  NAND2_X1   g05723(.A1(new_n5787_), .A2(new_n5773_), .ZN(new_n5788_));
  XOR2_X1    g05724(.A1(new_n5379_), .A2(new_n5381_), .Z(new_n5789_));
  OAI22_X1   g05725(.A1(new_n1764_), .A2(new_n4097_), .B1(new_n1729_), .B2(new_n3775_), .ZN(new_n5790_));
  NAND2_X1   g05726(.A1(new_n1862_), .A2(new_n3770_), .ZN(new_n5791_));
  AOI21_X1   g05727(.A1(new_n5790_), .A2(new_n5791_), .B(new_n4095_), .ZN(new_n5792_));
  NAND2_X1   g05728(.A1(new_n4810_), .A2(new_n5792_), .ZN(new_n5793_));
  XOR2_X1    g05729(.A1(new_n5793_), .A2(\a[20] ), .Z(new_n5794_));
  NAND2_X1   g05730(.A1(new_n5794_), .A2(new_n5789_), .ZN(new_n5795_));
  NOR2_X1    g05731(.A1(new_n5794_), .A2(new_n5789_), .ZN(new_n5796_));
  AOI21_X1   g05732(.A1(new_n5788_), .A2(new_n5795_), .B(new_n5796_), .ZN(new_n5797_));
  NAND2_X1   g05733(.A1(new_n5379_), .A2(new_n5381_), .ZN(new_n5798_));
  XOR2_X1    g05734(.A1(new_n5798_), .A2(new_n5375_), .Z(new_n5799_));
  OAI22_X1   g05735(.A1(new_n1764_), .A2(new_n3775_), .B1(new_n1729_), .B2(new_n3769_), .ZN(new_n5800_));
  NAND2_X1   g05736(.A1(new_n1613_), .A2(new_n4096_), .ZN(new_n5801_));
  AOI21_X1   g05737(.A1(new_n5801_), .A2(new_n5800_), .B(new_n4095_), .ZN(new_n5802_));
  NAND2_X1   g05738(.A1(new_n4778_), .A2(new_n5802_), .ZN(new_n5803_));
  XOR2_X1    g05739(.A1(new_n5803_), .A2(new_n3035_), .Z(new_n5804_));
  NOR2_X1    g05740(.A1(new_n5804_), .A2(new_n5799_), .ZN(new_n5805_));
  NAND2_X1   g05741(.A1(new_n5804_), .A2(new_n5799_), .ZN(new_n5806_));
  OAI21_X1   g05742(.A1(new_n5797_), .A2(new_n5805_), .B(new_n5806_), .ZN(new_n5807_));
  XOR2_X1    g05743(.A1(new_n5369_), .A2(\a[23] ), .Z(new_n5808_));
  XOR2_X1    g05744(.A1(new_n5808_), .A2(new_n4986_), .Z(new_n5809_));
  NAND2_X1   g05745(.A1(new_n5809_), .A2(new_n5383_), .ZN(new_n5810_));
  NAND2_X1   g05746(.A1(new_n5808_), .A2(new_n4986_), .ZN(new_n5811_));
  AOI21_X1   g05747(.A1(new_n5371_), .A2(new_n5811_), .B(new_n5383_), .ZN(new_n5812_));
  INV_X1     g05748(.I(new_n5812_), .ZN(new_n5813_));
  OAI22_X1   g05749(.A1(new_n1678_), .A2(new_n4097_), .B1(new_n1764_), .B2(new_n3769_), .ZN(new_n5814_));
  NAND2_X1   g05750(.A1(new_n1613_), .A2(new_n3776_), .ZN(new_n5815_));
  AOI21_X1   g05751(.A1(new_n5814_), .A2(new_n5815_), .B(new_n4095_), .ZN(new_n5816_));
  NAND2_X1   g05752(.A1(new_n4917_), .A2(new_n5816_), .ZN(new_n5817_));
  XOR2_X1    g05753(.A1(new_n5817_), .A2(\a[20] ), .Z(new_n5818_));
  NAND3_X1   g05754(.A1(new_n5810_), .A2(new_n5818_), .A3(new_n5813_), .ZN(new_n5819_));
  AOI21_X1   g05755(.A1(new_n5810_), .A2(new_n5813_), .B(new_n5818_), .ZN(new_n5820_));
  AOI21_X1   g05756(.A1(new_n5807_), .A2(new_n5819_), .B(new_n5820_), .ZN(new_n5821_));
  NOR2_X1    g05757(.A1(new_n5808_), .A2(new_n4986_), .ZN(new_n5822_));
  AOI21_X1   g05758(.A1(new_n5382_), .A2(new_n5811_), .B(new_n5822_), .ZN(new_n5823_));
  XNOR2_X1   g05759(.A1(new_n4985_), .A2(new_n4987_), .ZN(new_n5824_));
  NAND2_X1   g05760(.A1(new_n5391_), .A2(new_n5824_), .ZN(new_n5825_));
  XOR2_X1    g05761(.A1(new_n5390_), .A2(new_n84_), .Z(new_n5826_));
  NAND2_X1   g05762(.A1(new_n5826_), .A2(new_n5386_), .ZN(new_n5827_));
  AOI21_X1   g05763(.A1(new_n5825_), .A2(new_n5827_), .B(new_n5823_), .ZN(new_n5828_));
  NAND2_X1   g05764(.A1(new_n5826_), .A2(new_n5824_), .ZN(new_n5829_));
  AOI21_X1   g05765(.A1(new_n5392_), .A2(new_n5829_), .B(new_n5385_), .ZN(new_n5830_));
  NOR2_X1    g05766(.A1(new_n5828_), .A2(new_n5830_), .ZN(new_n5831_));
  OAI22_X1   g05767(.A1(new_n1678_), .A2(new_n3775_), .B1(new_n2071_), .B2(new_n4097_), .ZN(new_n5832_));
  NAND2_X1   g05768(.A1(new_n1613_), .A2(new_n3770_), .ZN(new_n5833_));
  AOI21_X1   g05769(.A1(new_n5832_), .A2(new_n5833_), .B(new_n4095_), .ZN(new_n5834_));
  NAND3_X1   g05770(.A1(new_n5070_), .A2(new_n3035_), .A3(new_n5834_), .ZN(new_n5835_));
  AOI21_X1   g05771(.A1(new_n5070_), .A2(new_n5834_), .B(new_n3035_), .ZN(new_n5836_));
  INV_X1     g05772(.I(new_n5836_), .ZN(new_n5837_));
  NAND2_X1   g05773(.A1(new_n5837_), .A2(new_n5835_), .ZN(new_n5838_));
  NOR2_X1    g05774(.A1(new_n5838_), .A2(new_n5831_), .ZN(new_n5839_));
  NOR2_X1    g05775(.A1(new_n5821_), .A2(new_n5839_), .ZN(new_n5840_));
  NAND2_X1   g05776(.A1(new_n5825_), .A2(new_n5827_), .ZN(new_n5841_));
  NAND2_X1   g05777(.A1(new_n5829_), .A2(new_n5392_), .ZN(new_n5842_));
  MUX2_X1    g05778(.I0(new_n5842_), .I1(new_n5841_), .S(new_n5385_), .Z(new_n5843_));
  INV_X1     g05779(.I(new_n5835_), .ZN(new_n5844_));
  NOR2_X1    g05780(.A1(new_n5844_), .A2(new_n5836_), .ZN(new_n5845_));
  NOR2_X1    g05781(.A1(new_n5843_), .A2(new_n5845_), .ZN(new_n5846_));
  NOR2_X1    g05782(.A1(new_n5840_), .A2(new_n5846_), .ZN(new_n5847_));
  NOR2_X1    g05783(.A1(new_n5826_), .A2(new_n5824_), .ZN(new_n5848_));
  OAI21_X1   g05784(.A1(new_n5823_), .A2(new_n5848_), .B(new_n5829_), .ZN(new_n5849_));
  XNOR2_X1   g05785(.A1(new_n5395_), .A2(new_n4978_), .ZN(new_n5850_));
  XOR2_X1    g05786(.A1(new_n5400_), .A2(\a[23] ), .Z(new_n5851_));
  XOR2_X1    g05787(.A1(new_n5851_), .A2(new_n5850_), .Z(new_n5852_));
  NAND2_X1   g05788(.A1(new_n5852_), .A2(new_n5849_), .ZN(new_n5853_));
  NAND2_X1   g05789(.A1(new_n5851_), .A2(new_n5850_), .ZN(new_n5854_));
  AOI21_X1   g05790(.A1(new_n5854_), .A2(new_n5403_), .B(new_n5849_), .ZN(new_n5855_));
  INV_X1     g05791(.I(new_n5855_), .ZN(new_n5856_));
  OAI22_X1   g05792(.A1(new_n2103_), .A2(new_n4097_), .B1(new_n1678_), .B2(new_n3769_), .ZN(new_n5857_));
  NAND2_X1   g05793(.A1(new_n2107_), .A2(new_n3776_), .ZN(new_n5858_));
  AOI21_X1   g05794(.A1(new_n5857_), .A2(new_n5858_), .B(new_n4095_), .ZN(new_n5859_));
  NAND3_X1   g05795(.A1(new_n4545_), .A2(new_n3035_), .A3(new_n5859_), .ZN(new_n5860_));
  OAI21_X1   g05796(.A1(new_n5103_), .A2(new_n5104_), .B(new_n5859_), .ZN(new_n5861_));
  NAND2_X1   g05797(.A1(new_n5861_), .A2(\a[20] ), .ZN(new_n5862_));
  NAND2_X1   g05798(.A1(new_n5860_), .A2(new_n5862_), .ZN(new_n5863_));
  AOI21_X1   g05799(.A1(new_n5856_), .A2(new_n5853_), .B(new_n5863_), .ZN(new_n5864_));
  NAND2_X1   g05800(.A1(new_n5856_), .A2(new_n5853_), .ZN(new_n5865_));
  INV_X1     g05801(.I(new_n5863_), .ZN(new_n5866_));
  NOR2_X1    g05802(.A1(new_n5865_), .A2(new_n5866_), .ZN(new_n5867_));
  NOR2_X1    g05803(.A1(new_n5867_), .A2(new_n5864_), .ZN(new_n5868_));
  NOR2_X1    g05804(.A1(new_n5868_), .A2(new_n5847_), .ZN(new_n5869_));
  INV_X1     g05805(.I(new_n5869_), .ZN(new_n5870_));
  AOI21_X1   g05806(.A1(new_n5849_), .A2(new_n5852_), .B(new_n5855_), .ZN(new_n5871_));
  XOR2_X1    g05807(.A1(new_n5871_), .A2(new_n5863_), .Z(new_n5872_));
  NAND2_X1   g05808(.A1(new_n5872_), .A2(new_n5847_), .ZN(new_n5873_));
  OAI22_X1   g05809(.A1(new_n2158_), .A2(new_n4291_), .B1(new_n2198_), .B2(new_n4297_), .ZN(new_n5874_));
  NAND2_X1   g05810(.A1(new_n1504_), .A2(new_n4469_), .ZN(new_n5875_));
  AOI21_X1   g05811(.A1(new_n5875_), .A2(new_n5874_), .B(new_n4468_), .ZN(new_n5876_));
  NAND2_X1   g05812(.A1(new_n4620_), .A2(new_n5876_), .ZN(new_n5877_));
  XOR2_X1    g05813(.A1(new_n5877_), .A2(\a[17] ), .Z(new_n5878_));
  AOI21_X1   g05814(.A1(new_n5870_), .A2(new_n5873_), .B(new_n5878_), .ZN(new_n5879_));
  INV_X1     g05815(.I(new_n5867_), .ZN(new_n5880_));
  OAI22_X1   g05816(.A1(new_n5840_), .A2(new_n5846_), .B1(new_n5871_), .B2(new_n5863_), .ZN(new_n5881_));
  AOI21_X1   g05817(.A1(new_n5407_), .A2(new_n5408_), .B(new_n5414_), .ZN(new_n5882_));
  XOR2_X1    g05818(.A1(new_n5413_), .A2(\a[23] ), .Z(new_n5883_));
  NOR2_X1    g05819(.A1(new_n5409_), .A2(new_n5883_), .ZN(new_n5884_));
  OAI21_X1   g05820(.A1(new_n5882_), .A2(new_n5884_), .B(new_n5404_), .ZN(new_n5885_));
  NOR2_X1    g05821(.A1(new_n5851_), .A2(new_n5850_), .ZN(new_n5886_));
  AOI21_X1   g05822(.A1(new_n5849_), .A2(new_n5854_), .B(new_n5886_), .ZN(new_n5887_));
  NOR2_X1    g05823(.A1(new_n5409_), .A2(new_n5414_), .ZN(new_n5888_));
  INV_X1     g05824(.I(new_n5416_), .ZN(new_n5889_));
  OAI21_X1   g05825(.A1(new_n5889_), .A2(new_n5888_), .B(new_n5887_), .ZN(new_n5890_));
  OAI22_X1   g05826(.A1(new_n2103_), .A2(new_n3775_), .B1(new_n2158_), .B2(new_n4097_), .ZN(new_n5891_));
  NAND2_X1   g05827(.A1(new_n2107_), .A2(new_n3770_), .ZN(new_n5892_));
  AOI21_X1   g05828(.A1(new_n5891_), .A2(new_n5892_), .B(new_n4095_), .ZN(new_n5893_));
  NAND3_X1   g05829(.A1(new_n4959_), .A2(new_n3035_), .A3(new_n5893_), .ZN(new_n5894_));
  OAI21_X1   g05830(.A1(new_n5260_), .A2(new_n5259_), .B(new_n5893_), .ZN(new_n5895_));
  NAND2_X1   g05831(.A1(new_n5895_), .A2(\a[20] ), .ZN(new_n5896_));
  NAND2_X1   g05832(.A1(new_n5896_), .A2(new_n5894_), .ZN(new_n5897_));
  NAND3_X1   g05833(.A1(new_n5897_), .A2(new_n5890_), .A3(new_n5885_), .ZN(new_n5898_));
  NAND2_X1   g05834(.A1(new_n5890_), .A2(new_n5885_), .ZN(new_n5899_));
  NAND3_X1   g05835(.A1(new_n5899_), .A2(new_n5894_), .A3(new_n5896_), .ZN(new_n5900_));
  NAND4_X1   g05836(.A1(new_n5881_), .A2(new_n5880_), .A3(new_n5900_), .A4(new_n5898_), .ZN(new_n5901_));
  NOR2_X1    g05837(.A1(new_n5785_), .A2(new_n5380_), .ZN(new_n5902_));
  AOI21_X1   g05838(.A1(new_n5784_), .A2(new_n5786_), .B(new_n5902_), .ZN(new_n5903_));
  XNOR2_X1   g05839(.A1(new_n5379_), .A2(new_n5381_), .ZN(new_n5904_));
  XOR2_X1    g05840(.A1(new_n5793_), .A2(new_n3035_), .Z(new_n5905_));
  NOR2_X1    g05841(.A1(new_n5905_), .A2(new_n5904_), .ZN(new_n5906_));
  NAND2_X1   g05842(.A1(new_n5905_), .A2(new_n5904_), .ZN(new_n5907_));
  OAI21_X1   g05843(.A1(new_n5903_), .A2(new_n5906_), .B(new_n5907_), .ZN(new_n5908_));
  INV_X1     g05844(.I(new_n5799_), .ZN(new_n5909_));
  XOR2_X1    g05845(.A1(new_n5803_), .A2(\a[20] ), .Z(new_n5910_));
  NAND2_X1   g05846(.A1(new_n5909_), .A2(new_n5910_), .ZN(new_n5911_));
  NOR2_X1    g05847(.A1(new_n5909_), .A2(new_n5910_), .ZN(new_n5912_));
  AOI21_X1   g05848(.A1(new_n5908_), .A2(new_n5911_), .B(new_n5912_), .ZN(new_n5913_));
  INV_X1     g05849(.I(new_n5819_), .ZN(new_n5914_));
  XOR2_X1    g05850(.A1(new_n5370_), .A2(new_n4986_), .Z(new_n5915_));
  NOR2_X1    g05851(.A1(new_n5915_), .A2(new_n5382_), .ZN(new_n5916_));
  XOR2_X1    g05852(.A1(new_n5817_), .A2(new_n3035_), .Z(new_n5917_));
  OAI21_X1   g05853(.A1(new_n5916_), .A2(new_n5812_), .B(new_n5917_), .ZN(new_n5918_));
  OAI21_X1   g05854(.A1(new_n5914_), .A2(new_n5913_), .B(new_n5918_), .ZN(new_n5919_));
  NAND2_X1   g05855(.A1(new_n5843_), .A2(new_n5845_), .ZN(new_n5920_));
  NAND2_X1   g05856(.A1(new_n5919_), .A2(new_n5920_), .ZN(new_n5921_));
  INV_X1     g05857(.I(new_n5846_), .ZN(new_n5922_));
  AOI21_X1   g05858(.A1(new_n5921_), .A2(new_n5922_), .B(new_n5864_), .ZN(new_n5923_));
  INV_X1     g05859(.I(new_n5898_), .ZN(new_n5924_));
  AOI21_X1   g05860(.A1(new_n5885_), .A2(new_n5890_), .B(new_n5897_), .ZN(new_n5925_));
  OAI22_X1   g05861(.A1(new_n5923_), .A2(new_n5867_), .B1(new_n5924_), .B2(new_n5925_), .ZN(new_n5926_));
  OAI22_X1   g05862(.A1(new_n4365_), .A2(new_n4470_), .B1(new_n2198_), .B2(new_n4291_), .ZN(new_n5927_));
  NAND2_X1   g05863(.A1(new_n1504_), .A2(new_n4298_), .ZN(new_n5928_));
  AOI21_X1   g05864(.A1(new_n5927_), .A2(new_n5928_), .B(new_n4468_), .ZN(new_n5929_));
  NAND3_X1   g05865(.A1(new_n4363_), .A2(new_n3372_), .A3(new_n5929_), .ZN(new_n5930_));
  AOI21_X1   g05866(.A1(new_n4363_), .A2(new_n5929_), .B(new_n3372_), .ZN(new_n5931_));
  INV_X1     g05867(.I(new_n5931_), .ZN(new_n5932_));
  NAND4_X1   g05868(.A1(new_n5926_), .A2(new_n5901_), .A3(new_n5932_), .A4(new_n5930_), .ZN(new_n5933_));
  AOI22_X1   g05869(.A1(new_n5926_), .A2(new_n5901_), .B1(new_n5932_), .B2(new_n5930_), .ZN(new_n5934_));
  AOI21_X1   g05870(.A1(new_n5879_), .A2(new_n5933_), .B(new_n5934_), .ZN(new_n5935_));
  XOR2_X1    g05871(.A1(new_n5428_), .A2(new_n5423_), .Z(new_n5936_));
  INV_X1     g05872(.I(new_n5430_), .ZN(new_n5937_));
  AOI21_X1   g05873(.A1(new_n5937_), .A2(new_n5429_), .B(new_n5417_), .ZN(new_n5938_));
  AOI21_X1   g05874(.A1(new_n5936_), .A2(new_n5417_), .B(new_n5938_), .ZN(new_n5939_));
  OAI22_X1   g05875(.A1(new_n2103_), .A2(new_n3769_), .B1(new_n2198_), .B2(new_n4097_), .ZN(new_n5940_));
  NAND2_X1   g05876(.A1(new_n2161_), .A2(new_n3776_), .ZN(new_n5941_));
  AOI21_X1   g05877(.A1(new_n5940_), .A2(new_n5941_), .B(new_n4095_), .ZN(new_n5942_));
  NAND2_X1   g05878(.A1(new_n5351_), .A2(new_n5942_), .ZN(new_n5943_));
  XOR2_X1    g05879(.A1(new_n5943_), .A2(new_n3035_), .Z(new_n5944_));
  AOI21_X1   g05880(.A1(new_n5901_), .A2(new_n5900_), .B(new_n5944_), .ZN(new_n5945_));
  NOR4_X1    g05881(.A1(new_n5923_), .A2(new_n5924_), .A3(new_n5925_), .A4(new_n5867_), .ZN(new_n5946_));
  INV_X1     g05882(.I(new_n5944_), .ZN(new_n5947_));
  NOR3_X1    g05883(.A1(new_n5946_), .A2(new_n5947_), .A3(new_n5925_), .ZN(new_n5948_));
  OAI21_X1   g05884(.A1(new_n5945_), .A2(new_n5948_), .B(new_n5939_), .ZN(new_n5949_));
  INV_X1     g05885(.I(new_n5939_), .ZN(new_n5950_));
  OAI21_X1   g05886(.A1(new_n5946_), .A2(new_n5925_), .B(new_n5947_), .ZN(new_n5951_));
  NAND3_X1   g05887(.A1(new_n5901_), .A2(new_n5900_), .A3(new_n5944_), .ZN(new_n5952_));
  NAND3_X1   g05888(.A1(new_n5951_), .A2(new_n5952_), .A3(new_n5950_), .ZN(new_n5953_));
  NAND2_X1   g05889(.A1(new_n5949_), .A2(new_n5953_), .ZN(new_n5954_));
  OAI22_X1   g05890(.A1(new_n2251_), .A2(new_n4470_), .B1(new_n4365_), .B2(new_n4297_), .ZN(new_n5955_));
  NAND2_X1   g05891(.A1(new_n1504_), .A2(new_n4292_), .ZN(new_n5956_));
  AOI21_X1   g05892(.A1(new_n5955_), .A2(new_n5956_), .B(new_n4468_), .ZN(new_n5957_));
  NAND3_X1   g05893(.A1(new_n4650_), .A2(new_n3372_), .A3(new_n5957_), .ZN(new_n5958_));
  OAI21_X1   g05894(.A1(new_n5730_), .A2(new_n5731_), .B(new_n5957_), .ZN(new_n5959_));
  NAND2_X1   g05895(.A1(new_n5959_), .A2(\a[17] ), .ZN(new_n5960_));
  NAND2_X1   g05896(.A1(new_n5960_), .A2(new_n5958_), .ZN(new_n5961_));
  INV_X1     g05897(.I(new_n5961_), .ZN(new_n5962_));
  AOI21_X1   g05898(.A1(new_n5954_), .A2(new_n5962_), .B(new_n5935_), .ZN(new_n5963_));
  NOR2_X1    g05899(.A1(new_n5954_), .A2(new_n5962_), .ZN(new_n5964_));
  NOR2_X1    g05900(.A1(new_n5963_), .A2(new_n5964_), .ZN(new_n5965_));
  OAI22_X1   g05901(.A1(new_n2311_), .A2(new_n4470_), .B1(new_n4365_), .B2(new_n4291_), .ZN(new_n5966_));
  NAND2_X1   g05902(.A1(new_n2255_), .A2(new_n4298_), .ZN(new_n5967_));
  AOI21_X1   g05903(.A1(new_n5966_), .A2(new_n5967_), .B(new_n4468_), .ZN(new_n5968_));
  NAND3_X1   g05904(.A1(new_n4419_), .A2(new_n3372_), .A3(new_n5968_), .ZN(new_n5969_));
  INV_X1     g05905(.I(new_n5969_), .ZN(new_n5970_));
  AOI21_X1   g05906(.A1(new_n4419_), .A2(new_n5968_), .B(new_n3372_), .ZN(new_n5971_));
  NOR2_X1    g05907(.A1(new_n5970_), .A2(new_n5971_), .ZN(new_n5972_));
  NOR4_X1    g05908(.A1(new_n5965_), .A2(new_n5766_), .A3(new_n5762_), .A4(new_n5972_), .ZN(new_n5973_));
  NOR3_X1    g05909(.A1(new_n5719_), .A2(new_n5727_), .A3(new_n5715_), .ZN(new_n5974_));
  AOI21_X1   g05910(.A1(new_n5740_), .A2(new_n5718_), .B(new_n5726_), .ZN(new_n5975_));
  NOR2_X1    g05911(.A1(new_n5974_), .A2(new_n5975_), .ZN(new_n5976_));
  NOR3_X1    g05912(.A1(new_n5963_), .A2(new_n5964_), .A3(new_n5972_), .ZN(new_n5977_));
  XOR2_X1    g05913(.A1(new_n5871_), .A2(new_n5866_), .Z(new_n5978_));
  NOR3_X1    g05914(.A1(new_n5978_), .A2(new_n5840_), .A3(new_n5846_), .ZN(new_n5979_));
  XOR2_X1    g05915(.A1(new_n5877_), .A2(new_n3372_), .Z(new_n5980_));
  OAI21_X1   g05916(.A1(new_n5869_), .A2(new_n5979_), .B(new_n5980_), .ZN(new_n5981_));
  INV_X1     g05917(.I(new_n5933_), .ZN(new_n5982_));
  NAND2_X1   g05918(.A1(new_n5926_), .A2(new_n5901_), .ZN(new_n5983_));
  NAND2_X1   g05919(.A1(new_n5932_), .A2(new_n5930_), .ZN(new_n5984_));
  NAND2_X1   g05920(.A1(new_n5983_), .A2(new_n5984_), .ZN(new_n5985_));
  OAI21_X1   g05921(.A1(new_n5982_), .A2(new_n5981_), .B(new_n5985_), .ZN(new_n5986_));
  AOI21_X1   g05922(.A1(new_n5951_), .A2(new_n5952_), .B(new_n5950_), .ZN(new_n5987_));
  NOR3_X1    g05923(.A1(new_n5945_), .A2(new_n5948_), .A3(new_n5939_), .ZN(new_n5988_));
  NOR2_X1    g05924(.A1(new_n5988_), .A2(new_n5987_), .ZN(new_n5989_));
  OAI21_X1   g05925(.A1(new_n5989_), .A2(new_n5961_), .B(new_n5986_), .ZN(new_n5990_));
  NAND3_X1   g05926(.A1(new_n5961_), .A2(new_n5949_), .A3(new_n5953_), .ZN(new_n5991_));
  INV_X1     g05927(.I(new_n5972_), .ZN(new_n5992_));
  AOI21_X1   g05928(.A1(new_n5990_), .A2(new_n5991_), .B(new_n5992_), .ZN(new_n5993_));
  OAI21_X1   g05929(.A1(new_n5993_), .A2(new_n5977_), .B(new_n5976_), .ZN(new_n5994_));
  NOR2_X1    g05930(.A1(new_n5994_), .A2(new_n5973_), .ZN(new_n5995_));
  NOR3_X1    g05931(.A1(new_n5745_), .A2(new_n5751_), .A3(new_n5689_), .ZN(new_n5996_));
  XOR2_X1    g05932(.A1(new_n5688_), .A2(new_n3372_), .Z(new_n5997_));
  OAI21_X1   g05933(.A1(new_n5750_), .A2(new_n5749_), .B(new_n5748_), .ZN(new_n5998_));
  NAND3_X1   g05934(.A1(new_n5737_), .A2(new_n5744_), .A3(new_n5698_), .ZN(new_n5999_));
  AOI21_X1   g05935(.A1(new_n5998_), .A2(new_n5999_), .B(new_n5997_), .ZN(new_n6000_));
  AOI21_X1   g05936(.A1(new_n5764_), .A2(new_n5765_), .B(new_n5759_), .ZN(new_n6001_));
  INV_X1     g05937(.I(new_n6001_), .ZN(new_n6002_));
  OAI21_X1   g05938(.A1(new_n5996_), .A2(new_n6000_), .B(new_n6002_), .ZN(new_n6003_));
  OAI21_X1   g05939(.A1(new_n5995_), .A2(new_n6003_), .B(new_n5752_), .ZN(new_n6004_));
  AOI21_X1   g05940(.A1(new_n5606_), .A2(new_n5676_), .B(\a[17] ), .ZN(new_n6005_));
  NOR2_X1    g05941(.A1(new_n5603_), .A2(new_n5605_), .ZN(new_n6006_));
  NOR3_X1    g05942(.A1(new_n6006_), .A2(new_n5552_), .A3(new_n3372_), .ZN(new_n6007_));
  OAI21_X1   g05943(.A1(new_n6007_), .A2(new_n6005_), .B(new_n5681_), .ZN(new_n6008_));
  INV_X1     g05944(.I(new_n5681_), .ZN(new_n6009_));
  OAI21_X1   g05945(.A1(new_n6006_), .A2(new_n5552_), .B(new_n3372_), .ZN(new_n6010_));
  NAND3_X1   g05946(.A1(new_n5606_), .A2(new_n5676_), .A3(\a[17] ), .ZN(new_n6011_));
  NAND3_X1   g05947(.A1(new_n6010_), .A2(new_n6011_), .A3(new_n6009_), .ZN(new_n6012_));
  NAND2_X1   g05948(.A1(new_n6008_), .A2(new_n6012_), .ZN(new_n6013_));
  OAI21_X1   g05949(.A1(new_n6004_), .A2(new_n6013_), .B(new_n5683_), .ZN(new_n6014_));
  NAND3_X1   g05950(.A1(new_n6014_), .A2(new_n5666_), .A3(new_n5675_), .ZN(new_n6015_));
  OAI21_X1   g05951(.A1(new_n6015_), .A2(new_n5653_), .B(new_n5655_), .ZN(new_n6016_));
  NAND2_X1   g05952(.A1(new_n5613_), .A2(new_n5614_), .ZN(new_n6017_));
  OAI21_X1   g05953(.A1(new_n5618_), .A2(new_n5622_), .B(new_n6017_), .ZN(new_n6018_));
  NOR2_X1    g05954(.A1(new_n5578_), .A2(new_n5582_), .ZN(new_n6019_));
  NOR2_X1    g05955(.A1(new_n5620_), .A2(new_n5594_), .ZN(new_n6020_));
  NOR2_X1    g05956(.A1(new_n5587_), .A2(new_n5621_), .ZN(new_n6021_));
  OAI21_X1   g05957(.A1(new_n6020_), .A2(new_n6021_), .B(new_n6019_), .ZN(new_n6022_));
  NAND2_X1   g05958(.A1(new_n6018_), .A2(new_n6022_), .ZN(new_n6023_));
  NOR4_X1    g05959(.A1(new_n5619_), .A2(new_n5623_), .A3(new_n5602_), .A4(new_n5622_), .ZN(new_n6024_));
  AOI22_X1   g05960(.A1(new_n5595_), .A2(new_n5596_), .B1(new_n5542_), .B2(new_n5600_), .ZN(new_n6025_));
  XOR2_X1    g05961(.A1(new_n5630_), .A2(new_n3372_), .Z(new_n6026_));
  OAI21_X1   g05962(.A1(new_n6025_), .A2(new_n6024_), .B(new_n6026_), .ZN(new_n6027_));
  NAND4_X1   g05963(.A1(new_n6016_), .A2(new_n6027_), .A3(new_n5632_), .A4(new_n6023_), .ZN(new_n6028_));
  XOR2_X1    g05964(.A1(new_n5630_), .A2(new_n3372_), .Z(new_n6029_));
  NOR3_X1    g05965(.A1(new_n6025_), .A2(new_n6024_), .A3(new_n6029_), .ZN(new_n6030_));
  NAND3_X1   g05966(.A1(new_n5647_), .A2(new_n5648_), .A3(new_n5651_), .ZN(new_n6031_));
  OAI21_X1   g05967(.A1(new_n5645_), .A2(new_n5642_), .B(new_n5641_), .ZN(new_n6032_));
  NAND2_X1   g05968(.A1(new_n6031_), .A2(new_n6032_), .ZN(new_n6033_));
  OAI22_X1   g05969(.A1(new_n5670_), .A2(new_n5667_), .B1(new_n5671_), .B2(new_n5672_), .ZN(new_n6034_));
  NAND2_X1   g05970(.A1(new_n6034_), .A2(new_n5666_), .ZN(new_n6035_));
  XOR2_X1    g05971(.A1(new_n5681_), .A2(\a[17] ), .Z(new_n6036_));
  NOR3_X1    g05972(.A1(new_n6036_), .A2(new_n5552_), .A3(new_n6006_), .ZN(new_n6037_));
  INV_X1     g05973(.I(new_n5752_), .ZN(new_n6038_));
  NAND3_X1   g05974(.A1(new_n5763_), .A2(new_n5765_), .A3(new_n5764_), .ZN(new_n6039_));
  OAI21_X1   g05975(.A1(new_n5760_), .A2(new_n5761_), .B(new_n5759_), .ZN(new_n6040_));
  AOI21_X1   g05976(.A1(new_n5949_), .A2(new_n5953_), .B(new_n5961_), .ZN(new_n6041_));
  OAI21_X1   g05977(.A1(new_n6041_), .A2(new_n5935_), .B(new_n5991_), .ZN(new_n6042_));
  NAND4_X1   g05978(.A1(new_n6040_), .A2(new_n6039_), .A3(new_n6042_), .A4(new_n5992_), .ZN(new_n6043_));
  NAND3_X1   g05979(.A1(new_n5990_), .A2(new_n5991_), .A3(new_n5992_), .ZN(new_n6044_));
  OAI21_X1   g05980(.A1(new_n5963_), .A2(new_n5964_), .B(new_n5972_), .ZN(new_n6045_));
  NAND2_X1   g05981(.A1(new_n6044_), .A2(new_n6045_), .ZN(new_n6046_));
  NAND3_X1   g05982(.A1(new_n6046_), .A2(new_n6043_), .A3(new_n5976_), .ZN(new_n6047_));
  NAND3_X1   g05983(.A1(new_n5998_), .A2(new_n5999_), .A3(new_n5997_), .ZN(new_n6048_));
  OAI21_X1   g05984(.A1(new_n5745_), .A2(new_n5751_), .B(new_n5689_), .ZN(new_n6049_));
  AOI21_X1   g05985(.A1(new_n6049_), .A2(new_n6048_), .B(new_n6001_), .ZN(new_n6050_));
  AOI21_X1   g05986(.A1(new_n6047_), .A2(new_n6050_), .B(new_n6038_), .ZN(new_n6051_));
  AOI21_X1   g05987(.A1(new_n6010_), .A2(new_n6011_), .B(new_n6009_), .ZN(new_n6052_));
  NOR3_X1    g05988(.A1(new_n6007_), .A2(new_n6005_), .A3(new_n5681_), .ZN(new_n6053_));
  NOR2_X1    g05989(.A1(new_n6053_), .A2(new_n6052_), .ZN(new_n6054_));
  AOI21_X1   g05990(.A1(new_n6051_), .A2(new_n6054_), .B(new_n6037_), .ZN(new_n6055_));
  NOR3_X1    g05991(.A1(new_n6055_), .A2(new_n5673_), .A3(new_n6035_), .ZN(new_n6056_));
  OAI21_X1   g05992(.A1(new_n6056_), .A2(new_n5641_), .B(new_n6033_), .ZN(new_n6057_));
  NOR2_X1    g05993(.A1(new_n5622_), .A2(new_n5618_), .ZN(new_n6058_));
  NOR2_X1    g05994(.A1(new_n6058_), .A2(new_n6019_), .ZN(new_n6059_));
  NOR2_X1    g05995(.A1(new_n6021_), .A2(new_n6020_), .ZN(new_n6060_));
  NOR2_X1    g05996(.A1(new_n6060_), .A2(new_n6017_), .ZN(new_n6061_));
  NOR2_X1    g05997(.A1(new_n6061_), .A2(new_n6059_), .ZN(new_n6062_));
  XOR2_X1    g05998(.A1(new_n5630_), .A2(\a[17] ), .Z(new_n6063_));
  AOI21_X1   g05999(.A1(new_n5624_), .A2(new_n5601_), .B(new_n6063_), .ZN(new_n6064_));
  OAI22_X1   g06000(.A1(new_n6057_), .A2(new_n6062_), .B1(new_n6064_), .B2(new_n6030_), .ZN(new_n6065_));
  NAND2_X1   g06001(.A1(new_n6056_), .A2(new_n6033_), .ZN(new_n6066_));
  NAND3_X1   g06002(.A1(new_n6066_), .A2(new_n5655_), .A3(new_n6023_), .ZN(new_n6067_));
  NAND2_X1   g06003(.A1(new_n6016_), .A2(new_n6062_), .ZN(new_n6068_));
  NAND2_X1   g06004(.A1(new_n6068_), .A2(new_n6067_), .ZN(new_n6069_));
  NAND4_X1   g06005(.A1(new_n6069_), .A2(new_n4731_), .A3(new_n6028_), .A4(new_n6065_), .ZN(new_n6070_));
  NAND2_X1   g06006(.A1(new_n6065_), .A2(new_n6028_), .ZN(new_n6071_));
  NOR2_X1    g06007(.A1(new_n6016_), .A2(new_n6062_), .ZN(new_n6072_));
  NOR2_X1    g06008(.A1(new_n6057_), .A2(new_n6023_), .ZN(new_n6073_));
  OAI21_X1   g06009(.A1(new_n6073_), .A2(new_n6072_), .B(new_n4731_), .ZN(new_n6074_));
  NAND2_X1   g06010(.A1(new_n6071_), .A2(new_n6074_), .ZN(new_n6075_));
  INV_X1     g06011(.I(\a[12] ), .ZN(new_n6076_));
  NOR2_X1    g06012(.A1(new_n6076_), .A2(\a[11] ), .ZN(new_n6077_));
  NOR2_X1    g06013(.A1(new_n4034_), .A2(\a[12] ), .ZN(new_n6078_));
  NOR2_X1    g06014(.A1(new_n6077_), .A2(new_n6078_), .ZN(new_n6079_));
  XNOR2_X1   g06015(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n6080_));
  NOR2_X1    g06016(.A1(new_n6079_), .A2(new_n6080_), .ZN(new_n6081_));
  INV_X1     g06017(.I(new_n6081_), .ZN(new_n6082_));
  INV_X1     g06018(.I(new_n6079_), .ZN(new_n6083_));
  INV_X1     g06019(.I(\a[13] ), .ZN(new_n6084_));
  NOR2_X1    g06020(.A1(new_n6084_), .A2(\a[11] ), .ZN(new_n6085_));
  NOR2_X1    g06021(.A1(new_n4034_), .A2(\a[13] ), .ZN(new_n6086_));
  OR2_X2     g06022(.A1(new_n6085_), .A2(new_n6086_), .Z(new_n6087_));
  XNOR2_X1   g06023(.A1(\a[11] ), .A2(\a[14] ), .ZN(new_n6088_));
  OAI21_X1   g06024(.A1(new_n6083_), .A2(new_n6087_), .B(new_n6088_), .ZN(new_n6089_));
  NOR2_X1    g06025(.A1(new_n6083_), .A2(new_n6080_), .ZN(new_n6090_));
  INV_X1     g06026(.I(new_n6090_), .ZN(new_n6091_));
  OAI22_X1   g06027(.A1(new_n1180_), .A2(new_n6091_), .B1(new_n2492_), .B2(new_n6089_), .ZN(new_n6092_));
  NOR3_X1    g06028(.A1(new_n6084_), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n6093_));
  AOI21_X1   g06029(.A1(\a[12] ), .A2(new_n6086_), .B(new_n6093_), .ZN(new_n6094_));
  INV_X1     g06030(.I(new_n6094_), .ZN(new_n6095_));
  NAND2_X1   g06031(.A1(new_n1122_), .A2(new_n6095_), .ZN(new_n6096_));
  AOI21_X1   g06032(.A1(new_n6096_), .A2(new_n6092_), .B(new_n6082_), .ZN(new_n6097_));
  NAND2_X1   g06033(.A1(new_n3330_), .A2(new_n6097_), .ZN(new_n6098_));
  XOR2_X1    g06034(.A1(new_n6098_), .A2(new_n3521_), .Z(new_n6099_));
  AOI21_X1   g06035(.A1(new_n6075_), .A2(new_n6070_), .B(new_n6099_), .ZN(new_n6100_));
  NOR2_X1    g06036(.A1(new_n6062_), .A2(new_n4731_), .ZN(new_n6101_));
  NOR2_X1    g06037(.A1(new_n6023_), .A2(new_n4730_), .ZN(new_n6102_));
  OAI21_X1   g06038(.A1(new_n6101_), .A2(new_n6102_), .B(new_n6016_), .ZN(new_n6103_));
  NOR2_X1    g06039(.A1(new_n6023_), .A2(new_n4731_), .ZN(new_n6104_));
  NOR2_X1    g06040(.A1(new_n6062_), .A2(new_n4730_), .ZN(new_n6105_));
  OAI21_X1   g06041(.A1(new_n6105_), .A2(new_n6104_), .B(new_n6057_), .ZN(new_n6106_));
  OAI22_X1   g06042(.A1(new_n1121_), .A2(new_n6091_), .B1(new_n2451_), .B2(new_n6089_), .ZN(new_n6107_));
  NAND2_X1   g06043(.A1(new_n2496_), .A2(new_n6095_), .ZN(new_n6108_));
  AOI21_X1   g06044(.A1(new_n6107_), .A2(new_n6108_), .B(new_n6082_), .ZN(new_n6109_));
  NAND3_X1   g06045(.A1(new_n3393_), .A2(new_n3521_), .A3(new_n6109_), .ZN(new_n6110_));
  NAND2_X1   g06046(.A1(new_n3393_), .A2(new_n6109_), .ZN(new_n6111_));
  NAND2_X1   g06047(.A1(new_n6111_), .A2(\a[14] ), .ZN(new_n6112_));
  NAND2_X1   g06048(.A1(new_n6112_), .A2(new_n6110_), .ZN(new_n6113_));
  NAND3_X1   g06049(.A1(new_n6103_), .A2(new_n6106_), .A3(new_n6113_), .ZN(new_n6114_));
  INV_X1     g06050(.I(new_n6114_), .ZN(new_n6115_));
  NOR2_X1    g06051(.A1(new_n6071_), .A2(new_n6074_), .ZN(new_n6116_));
  AOI22_X1   g06052(.A1(new_n6069_), .A2(new_n4731_), .B1(new_n6028_), .B2(new_n6065_), .ZN(new_n6117_));
  XOR2_X1    g06053(.A1(new_n6098_), .A2(\a[14] ), .Z(new_n6118_));
  NOR3_X1    g06054(.A1(new_n6116_), .A2(new_n6117_), .A3(new_n6118_), .ZN(new_n6119_));
  NOR3_X1    g06055(.A1(new_n6119_), .A2(new_n6100_), .A3(new_n6115_), .ZN(new_n6120_));
  OAI21_X1   g06056(.A1(new_n6116_), .A2(new_n6117_), .B(new_n6118_), .ZN(new_n6121_));
  NAND3_X1   g06057(.A1(new_n6075_), .A2(new_n6070_), .A3(new_n6099_), .ZN(new_n6122_));
  AOI21_X1   g06058(.A1(new_n6121_), .A2(new_n6122_), .B(new_n6114_), .ZN(new_n6123_));
  NOR2_X1    g06059(.A1(new_n2915_), .A2(new_n813_), .ZN(new_n6124_));
  AOI21_X1   g06060(.A1(new_n2910_), .A2(new_n2912_), .B(new_n814_), .ZN(new_n6125_));
  OAI21_X1   g06061(.A1(new_n896_), .A2(new_n4719_), .B(new_n4706_), .ZN(new_n6126_));
  OAI22_X1   g06062(.A1(new_n813_), .A2(new_n4710_), .B1(new_n1008_), .B2(new_n4716_), .ZN(new_n6127_));
  NOR2_X1    g06063(.A1(new_n6127_), .A2(new_n6126_), .ZN(new_n6128_));
  OAI21_X1   g06064(.A1(new_n6125_), .A2(new_n6124_), .B(new_n6128_), .ZN(new_n6129_));
  XOR2_X1    g06065(.A1(new_n6129_), .A2(new_n4034_), .Z(new_n6130_));
  NOR3_X1    g06066(.A1(new_n6120_), .A2(new_n6130_), .A3(new_n6123_), .ZN(new_n6131_));
  NAND3_X1   g06067(.A1(new_n6121_), .A2(new_n6122_), .A3(new_n6114_), .ZN(new_n6132_));
  OAI21_X1   g06068(.A1(new_n6119_), .A2(new_n6100_), .B(new_n6115_), .ZN(new_n6133_));
  XOR2_X1    g06069(.A1(new_n6129_), .A2(\a[11] ), .Z(new_n6134_));
  NAND3_X1   g06070(.A1(new_n6133_), .A2(new_n6134_), .A3(new_n6132_), .ZN(new_n6135_));
  NAND3_X1   g06071(.A1(new_n2917_), .A2(new_n4034_), .A3(new_n6128_), .ZN(new_n6136_));
  NAND2_X1   g06072(.A1(new_n6129_), .A2(\a[11] ), .ZN(new_n6137_));
  NAND2_X1   g06073(.A1(new_n6137_), .A2(new_n6136_), .ZN(new_n6138_));
  OAI21_X1   g06074(.A1(new_n6120_), .A2(new_n6123_), .B(new_n6138_), .ZN(new_n6139_));
  NAND2_X1   g06075(.A1(new_n6135_), .A2(new_n6139_), .ZN(new_n6140_));
  OAI22_X1   g06076(.A1(new_n896_), .A2(new_n4710_), .B1(new_n1180_), .B2(new_n4716_), .ZN(new_n6141_));
  NAND2_X1   g06077(.A1(new_n2504_), .A2(new_n4720_), .ZN(new_n6142_));
  AOI21_X1   g06078(.A1(new_n6142_), .A2(new_n6141_), .B(new_n4707_), .ZN(new_n6143_));
  AND3_X2    g06079(.A1(new_n3596_), .A2(new_n4034_), .A3(new_n6143_), .Z(new_n6144_));
  AOI21_X1   g06080(.A1(new_n3596_), .A2(new_n6143_), .B(new_n4034_), .ZN(new_n6145_));
  NOR2_X1    g06081(.A1(new_n6144_), .A2(new_n6145_), .ZN(new_n6146_));
  INV_X1     g06082(.I(new_n6146_), .ZN(new_n6147_));
  AOI21_X1   g06083(.A1(new_n6103_), .A2(new_n6106_), .B(new_n6113_), .ZN(new_n6148_));
  NOR2_X1    g06084(.A1(new_n6115_), .A2(new_n6148_), .ZN(new_n6149_));
  NOR2_X1    g06085(.A1(new_n6147_), .A2(new_n6149_), .ZN(new_n6150_));
  NOR2_X1    g06086(.A1(new_n3560_), .A2(new_n1008_), .ZN(new_n6151_));
  AOI21_X1   g06087(.A1(new_n3557_), .A2(new_n3328_), .B(new_n2504_), .ZN(new_n6152_));
  OAI22_X1   g06088(.A1(new_n1008_), .A2(new_n4710_), .B1(new_n1121_), .B2(new_n4716_), .ZN(new_n6153_));
  NAND2_X1   g06089(.A1(new_n1181_), .A2(new_n4720_), .ZN(new_n6154_));
  AOI21_X1   g06090(.A1(new_n6153_), .A2(new_n6154_), .B(new_n4707_), .ZN(new_n6155_));
  OAI21_X1   g06091(.A1(new_n6151_), .A2(new_n6152_), .B(new_n6155_), .ZN(new_n6156_));
  XOR2_X1    g06092(.A1(new_n6156_), .A2(\a[11] ), .Z(new_n6157_));
  XOR2_X1    g06093(.A1(new_n6156_), .A2(new_n4034_), .Z(new_n6158_));
  NAND2_X1   g06094(.A1(new_n6015_), .A2(new_n5641_), .ZN(new_n6159_));
  NOR4_X1    g06095(.A1(new_n6055_), .A2(new_n5641_), .A3(new_n6035_), .A4(new_n5673_), .ZN(new_n6160_));
  INV_X1     g06096(.I(new_n6160_), .ZN(new_n6161_));
  AOI21_X1   g06097(.A1(new_n6161_), .A2(new_n6159_), .B(new_n5654_), .ZN(new_n6162_));
  INV_X1     g06098(.I(new_n5654_), .ZN(new_n6163_));
  NOR2_X1    g06099(.A1(new_n6056_), .A2(new_n5647_), .ZN(new_n6164_));
  NOR3_X1    g06100(.A1(new_n6164_), .A2(new_n6163_), .A3(new_n6160_), .ZN(new_n6165_));
  NOR2_X1    g06101(.A1(new_n6162_), .A2(new_n6165_), .ZN(new_n6166_));
  NAND2_X1   g06102(.A1(new_n6055_), .A2(new_n5675_), .ZN(new_n6167_));
  NAND2_X1   g06103(.A1(new_n6014_), .A2(new_n6035_), .ZN(new_n6168_));
  OAI22_X1   g06104(.A1(new_n2367_), .A2(new_n6089_), .B1(new_n2451_), .B2(new_n6091_), .ZN(new_n6169_));
  NAND2_X1   g06105(.A1(new_n2412_), .A2(new_n6095_), .ZN(new_n6170_));
  AOI21_X1   g06106(.A1(new_n6169_), .A2(new_n6170_), .B(new_n6082_), .ZN(new_n6171_));
  OAI21_X1   g06107(.A1(new_n5626_), .A2(new_n5625_), .B(new_n6171_), .ZN(new_n6172_));
  XOR2_X1    g06108(.A1(new_n6172_), .A2(new_n3521_), .Z(new_n6173_));
  AOI21_X1   g06109(.A1(new_n6168_), .A2(new_n6167_), .B(new_n6173_), .ZN(new_n6174_));
  NOR2_X1    g06110(.A1(new_n6014_), .A2(new_n6035_), .ZN(new_n6175_));
  NOR2_X1    g06111(.A1(new_n6055_), .A2(new_n5675_), .ZN(new_n6176_));
  XOR2_X1    g06112(.A1(new_n6172_), .A2(\a[14] ), .Z(new_n6177_));
  NOR3_X1    g06113(.A1(new_n6175_), .A2(new_n6176_), .A3(new_n6177_), .ZN(new_n6178_));
  OAI22_X1   g06114(.A1(new_n2367_), .A2(new_n6094_), .B1(new_n2408_), .B2(new_n6091_), .ZN(new_n6179_));
  INV_X1     g06115(.I(new_n6089_), .ZN(new_n6180_));
  NAND2_X1   g06116(.A1(new_n1334_), .A2(new_n6180_), .ZN(new_n6181_));
  AOI21_X1   g06117(.A1(new_n6179_), .A2(new_n6181_), .B(new_n6082_), .ZN(new_n6182_));
  NAND3_X1   g06118(.A1(new_n3708_), .A2(new_n3521_), .A3(new_n6182_), .ZN(new_n6183_));
  AOI21_X1   g06119(.A1(new_n3708_), .A2(new_n6182_), .B(new_n3521_), .ZN(new_n6184_));
  INV_X1     g06120(.I(new_n6184_), .ZN(new_n6185_));
  NAND2_X1   g06121(.A1(new_n6185_), .A2(new_n6183_), .ZN(new_n6186_));
  NOR2_X1    g06122(.A1(new_n6004_), .A2(new_n6054_), .ZN(new_n6187_));
  NOR2_X1    g06123(.A1(new_n6051_), .A2(new_n6013_), .ZN(new_n6188_));
  NOR2_X1    g06124(.A1(new_n6187_), .A2(new_n6188_), .ZN(new_n6189_));
  NOR2_X1    g06125(.A1(new_n6189_), .A2(new_n6186_), .ZN(new_n6190_));
  NOR3_X1    g06126(.A1(new_n6174_), .A2(new_n6178_), .A3(new_n6190_), .ZN(new_n6191_));
  OAI22_X1   g06127(.A1(new_n2492_), .A2(new_n6091_), .B1(new_n2408_), .B2(new_n6089_), .ZN(new_n6192_));
  NAND2_X1   g06128(.A1(new_n2454_), .A2(new_n6095_), .ZN(new_n6193_));
  AOI21_X1   g06129(.A1(new_n6193_), .A2(new_n6192_), .B(new_n6082_), .ZN(new_n6194_));
  NAND2_X1   g06130(.A1(new_n3577_), .A2(new_n6194_), .ZN(new_n6195_));
  XOR2_X1    g06131(.A1(new_n6195_), .A2(new_n3521_), .Z(new_n6196_));
  NOR2_X1    g06132(.A1(new_n6191_), .A2(new_n6196_), .ZN(new_n6197_));
  OAI21_X1   g06133(.A1(new_n6175_), .A2(new_n6176_), .B(new_n6177_), .ZN(new_n6198_));
  NAND3_X1   g06134(.A1(new_n6168_), .A2(new_n6167_), .A3(new_n6173_), .ZN(new_n6199_));
  INV_X1     g06135(.I(new_n6183_), .ZN(new_n6200_));
  NOR2_X1    g06136(.A1(new_n6200_), .A2(new_n6184_), .ZN(new_n6201_));
  XOR2_X1    g06137(.A1(new_n6051_), .A2(new_n6054_), .Z(new_n6202_));
  NAND2_X1   g06138(.A1(new_n6202_), .A2(new_n6201_), .ZN(new_n6203_));
  NAND3_X1   g06139(.A1(new_n6198_), .A2(new_n6203_), .A3(new_n6199_), .ZN(new_n6204_));
  XOR2_X1    g06140(.A1(new_n6195_), .A2(\a[14] ), .Z(new_n6205_));
  NOR2_X1    g06141(.A1(new_n6204_), .A2(new_n6205_), .ZN(new_n6206_));
  OAI21_X1   g06142(.A1(new_n6206_), .A2(new_n6197_), .B(new_n6166_), .ZN(new_n6207_));
  OAI21_X1   g06143(.A1(new_n6164_), .A2(new_n6160_), .B(new_n6163_), .ZN(new_n6208_));
  NAND3_X1   g06144(.A1(new_n6161_), .A2(new_n6159_), .A3(new_n5654_), .ZN(new_n6209_));
  NAND2_X1   g06145(.A1(new_n6209_), .A2(new_n6208_), .ZN(new_n6210_));
  NAND2_X1   g06146(.A1(new_n6204_), .A2(new_n6205_), .ZN(new_n6211_));
  NAND2_X1   g06147(.A1(new_n6191_), .A2(new_n6196_), .ZN(new_n6212_));
  NAND3_X1   g06148(.A1(new_n6211_), .A2(new_n6212_), .A3(new_n6210_), .ZN(new_n6213_));
  NAND3_X1   g06149(.A1(new_n6158_), .A2(new_n6207_), .A3(new_n6213_), .ZN(new_n6214_));
  AOI21_X1   g06150(.A1(new_n6211_), .A2(new_n6212_), .B(new_n6210_), .ZN(new_n6215_));
  NOR3_X1    g06151(.A1(new_n6206_), .A2(new_n6197_), .A3(new_n6166_), .ZN(new_n6216_));
  OAI21_X1   g06152(.A1(new_n6215_), .A2(new_n6216_), .B(new_n6157_), .ZN(new_n6217_));
  NAND2_X1   g06153(.A1(new_n6217_), .A2(new_n6214_), .ZN(new_n6218_));
  OAI22_X1   g06154(.A1(new_n1180_), .A2(new_n4710_), .B1(new_n2492_), .B2(new_n4716_), .ZN(new_n6219_));
  NAND2_X1   g06155(.A1(new_n1122_), .A2(new_n4720_), .ZN(new_n6220_));
  AOI21_X1   g06156(.A1(new_n6220_), .A2(new_n6219_), .B(new_n4707_), .ZN(new_n6221_));
  NAND2_X1   g06157(.A1(new_n3330_), .A2(new_n6221_), .ZN(new_n6222_));
  NOR2_X1    g06158(.A1(new_n6222_), .A2(\a[11] ), .ZN(new_n6223_));
  INV_X1     g06159(.I(new_n6223_), .ZN(new_n6224_));
  NAND2_X1   g06160(.A1(new_n6222_), .A2(\a[11] ), .ZN(new_n6225_));
  NOR2_X1    g06161(.A1(new_n6202_), .A2(new_n6201_), .ZN(new_n6226_));
  NAND3_X1   g06162(.A1(new_n6198_), .A2(new_n6226_), .A3(new_n6199_), .ZN(new_n6227_));
  AOI21_X1   g06163(.A1(new_n6198_), .A2(new_n6199_), .B(new_n6226_), .ZN(new_n6228_));
  INV_X1     g06164(.I(new_n6228_), .ZN(new_n6229_));
  NAND4_X1   g06165(.A1(new_n6229_), .A2(new_n6224_), .A3(new_n6225_), .A4(new_n6227_), .ZN(new_n6230_));
  INV_X1     g06166(.I(new_n6230_), .ZN(new_n6231_));
  INV_X1     g06167(.I(new_n6225_), .ZN(new_n6232_));
  INV_X1     g06168(.I(new_n6227_), .ZN(new_n6233_));
  OAI22_X1   g06169(.A1(new_n6233_), .A2(new_n6228_), .B1(new_n6232_), .B2(new_n6223_), .ZN(new_n6234_));
  NAND2_X1   g06170(.A1(new_n6234_), .A2(new_n6230_), .ZN(new_n6235_));
  OAI21_X1   g06171(.A1(new_n2492_), .A2(new_n4719_), .B(new_n4706_), .ZN(new_n6236_));
  OAI22_X1   g06172(.A1(new_n1121_), .A2(new_n4710_), .B1(new_n2451_), .B2(new_n4716_), .ZN(new_n6237_));
  NOR2_X1    g06173(.A1(new_n6237_), .A2(new_n6236_), .ZN(new_n6238_));
  NAND2_X1   g06174(.A1(new_n3393_), .A2(new_n6238_), .ZN(new_n6239_));
  XOR2_X1    g06175(.A1(new_n6239_), .A2(\a[11] ), .Z(new_n6240_));
  NOR3_X1    g06176(.A1(new_n6240_), .A2(new_n6190_), .A3(new_n6226_), .ZN(new_n6241_));
  OAI22_X1   g06177(.A1(new_n2492_), .A2(new_n4710_), .B1(new_n2408_), .B2(new_n4716_), .ZN(new_n6242_));
  NAND2_X1   g06178(.A1(new_n2454_), .A2(new_n4720_), .ZN(new_n6243_));
  AOI21_X1   g06179(.A1(new_n6243_), .A2(new_n6242_), .B(new_n4707_), .ZN(new_n6244_));
  NAND2_X1   g06180(.A1(new_n3577_), .A2(new_n6244_), .ZN(new_n6245_));
  XOR2_X1    g06181(.A1(new_n6245_), .A2(\a[11] ), .Z(new_n6246_));
  NOR2_X1    g06182(.A1(new_n5745_), .A2(new_n5751_), .ZN(new_n6247_));
  NOR2_X1    g06183(.A1(new_n5995_), .A2(new_n6001_), .ZN(new_n6248_));
  NOR2_X1    g06184(.A1(new_n6248_), .A2(new_n5997_), .ZN(new_n6249_));
  NAND2_X1   g06185(.A1(new_n6047_), .A2(new_n6002_), .ZN(new_n6250_));
  NOR2_X1    g06186(.A1(new_n6250_), .A2(new_n5689_), .ZN(new_n6251_));
  OAI21_X1   g06187(.A1(new_n6249_), .A2(new_n6251_), .B(new_n6247_), .ZN(new_n6252_));
  INV_X1     g06188(.I(new_n6247_), .ZN(new_n6253_));
  NAND2_X1   g06189(.A1(new_n6250_), .A2(new_n5689_), .ZN(new_n6254_));
  NAND2_X1   g06190(.A1(new_n6248_), .A2(new_n5997_), .ZN(new_n6255_));
  NAND3_X1   g06191(.A1(new_n6255_), .A2(new_n6254_), .A3(new_n6253_), .ZN(new_n6256_));
  NAND2_X1   g06192(.A1(new_n6252_), .A2(new_n6256_), .ZN(new_n6257_));
  OAI22_X1   g06193(.A1(new_n1409_), .A2(new_n6094_), .B1(new_n1333_), .B2(new_n6091_), .ZN(new_n6258_));
  NAND2_X1   g06194(.A1(new_n2359_), .A2(new_n6180_), .ZN(new_n6259_));
  AOI21_X1   g06195(.A1(new_n6258_), .A2(new_n6259_), .B(new_n6082_), .ZN(new_n6260_));
  NAND2_X1   g06196(.A1(new_n3828_), .A2(new_n6260_), .ZN(new_n6261_));
  XOR2_X1    g06197(.A1(new_n6261_), .A2(\a[14] ), .Z(new_n6262_));
  NOR2_X1    g06198(.A1(new_n5965_), .A2(new_n5972_), .ZN(new_n6263_));
  INV_X1     g06199(.I(new_n6263_), .ZN(new_n6264_));
  NAND2_X1   g06200(.A1(new_n6040_), .A2(new_n6039_), .ZN(new_n6265_));
  NOR2_X1    g06201(.A1(new_n5994_), .A2(new_n6265_), .ZN(new_n6266_));
  NOR2_X1    g06202(.A1(new_n5766_), .A2(new_n5762_), .ZN(new_n6267_));
  AOI21_X1   g06203(.A1(new_n6046_), .A2(new_n5976_), .B(new_n6267_), .ZN(new_n6268_));
  NOR3_X1    g06204(.A1(new_n6266_), .A2(new_n6268_), .A3(new_n6264_), .ZN(new_n6269_));
  NAND3_X1   g06205(.A1(new_n6046_), .A2(new_n5976_), .A3(new_n6267_), .ZN(new_n6270_));
  NAND2_X1   g06206(.A1(new_n5994_), .A2(new_n6265_), .ZN(new_n6271_));
  AOI21_X1   g06207(.A1(new_n6271_), .A2(new_n6270_), .B(new_n6263_), .ZN(new_n6272_));
  OAI21_X1   g06208(.A1(new_n6269_), .A2(new_n6272_), .B(new_n6262_), .ZN(new_n6273_));
  XOR2_X1    g06209(.A1(new_n6261_), .A2(new_n3521_), .Z(new_n6274_));
  NAND3_X1   g06210(.A1(new_n6271_), .A2(new_n6270_), .A3(new_n6263_), .ZN(new_n6275_));
  OAI21_X1   g06211(.A1(new_n6266_), .A2(new_n6268_), .B(new_n6264_), .ZN(new_n6276_));
  NAND3_X1   g06212(.A1(new_n6276_), .A2(new_n6275_), .A3(new_n6274_), .ZN(new_n6277_));
  NOR2_X1    g06213(.A1(new_n1453_), .A2(new_n6094_), .ZN(new_n6278_));
  NOR2_X1    g06214(.A1(new_n1409_), .A2(new_n6091_), .ZN(new_n6279_));
  NOR2_X1    g06215(.A1(new_n2351_), .A2(new_n6089_), .ZN(new_n6280_));
  NOR4_X1    g06216(.A1(new_n6279_), .A2(new_n6082_), .A3(new_n6278_), .A4(new_n6280_), .ZN(new_n6281_));
  NAND2_X1   g06217(.A1(new_n3904_), .A2(new_n6281_), .ZN(new_n6282_));
  NAND2_X1   g06218(.A1(new_n6282_), .A2(\a[14] ), .ZN(new_n6283_));
  NAND3_X1   g06219(.A1(new_n3904_), .A2(new_n3521_), .A3(new_n6281_), .ZN(new_n6284_));
  NOR3_X1    g06220(.A1(new_n5976_), .A2(new_n5970_), .A3(new_n5971_), .ZN(new_n6285_));
  INV_X1     g06221(.I(new_n5976_), .ZN(new_n6286_));
  NOR2_X1    g06222(.A1(new_n5972_), .A2(new_n6286_), .ZN(new_n6287_));
  OAI21_X1   g06223(.A1(new_n6285_), .A2(new_n6287_), .B(new_n6042_), .ZN(new_n6288_));
  NAND2_X1   g06224(.A1(new_n5972_), .A2(new_n5976_), .ZN(new_n6289_));
  OAI21_X1   g06225(.A1(new_n5970_), .A2(new_n5971_), .B(new_n6286_), .ZN(new_n6290_));
  NAND2_X1   g06226(.A1(new_n6290_), .A2(new_n6289_), .ZN(new_n6291_));
  NAND2_X1   g06227(.A1(new_n6291_), .A2(new_n5965_), .ZN(new_n6292_));
  NAND4_X1   g06228(.A1(new_n6292_), .A2(new_n6283_), .A3(new_n6288_), .A4(new_n6284_), .ZN(new_n6293_));
  XOR2_X1    g06229(.A1(new_n5910_), .A2(new_n5799_), .Z(new_n6294_));
  NOR2_X1    g06230(.A1(new_n6294_), .A2(new_n5797_), .ZN(new_n6295_));
  AOI21_X1   g06231(.A1(new_n5911_), .A2(new_n5806_), .B(new_n5908_), .ZN(new_n6296_));
  NOR2_X1    g06232(.A1(new_n6295_), .A2(new_n6296_), .ZN(new_n6297_));
  OAI22_X1   g06233(.A1(new_n2103_), .A2(new_n4470_), .B1(new_n1678_), .B2(new_n4291_), .ZN(new_n6298_));
  NAND2_X1   g06234(.A1(new_n2107_), .A2(new_n4298_), .ZN(new_n6299_));
  AOI21_X1   g06235(.A1(new_n6298_), .A2(new_n6299_), .B(new_n4468_), .ZN(new_n6300_));
  NAND2_X1   g06236(.A1(new_n4545_), .A2(new_n6300_), .ZN(new_n6301_));
  XOR2_X1    g06237(.A1(new_n6301_), .A2(\a[17] ), .Z(new_n6302_));
  XOR2_X1    g06238(.A1(new_n6302_), .A2(new_n6297_), .Z(new_n6303_));
  OAI22_X1   g06239(.A1(new_n2158_), .A2(new_n6089_), .B1(new_n2198_), .B2(new_n6094_), .ZN(new_n6304_));
  OAI21_X1   g06240(.A1(new_n1503_), .A2(new_n6091_), .B(new_n6304_), .ZN(new_n6305_));
  AOI21_X1   g06241(.A1(new_n4620_), .A2(new_n6081_), .B(new_n6305_), .ZN(new_n6306_));
  XOR2_X1    g06242(.A1(new_n6306_), .A2(new_n3521_), .Z(new_n6307_));
  NOR2_X1    g06243(.A1(new_n6307_), .A2(new_n6303_), .ZN(new_n6308_));
  OAI22_X1   g06244(.A1(new_n4365_), .A2(new_n6091_), .B1(new_n2198_), .B2(new_n6089_), .ZN(new_n6309_));
  NAND2_X1   g06245(.A1(new_n1504_), .A2(new_n6095_), .ZN(new_n6310_));
  AOI21_X1   g06246(.A1(new_n6309_), .A2(new_n6310_), .B(new_n6082_), .ZN(new_n6311_));
  NAND3_X1   g06247(.A1(new_n4363_), .A2(new_n3521_), .A3(new_n6311_), .ZN(new_n6312_));
  INV_X1     g06248(.I(new_n6312_), .ZN(new_n6313_));
  AOI21_X1   g06249(.A1(new_n4363_), .A2(new_n6311_), .B(new_n3521_), .ZN(new_n6314_));
  NOR2_X1    g06250(.A1(new_n6313_), .A2(new_n6314_), .ZN(new_n6315_));
  INV_X1     g06251(.I(new_n6302_), .ZN(new_n6316_));
  NAND2_X1   g06252(.A1(new_n6316_), .A2(new_n6297_), .ZN(new_n6317_));
  AOI21_X1   g06253(.A1(new_n5810_), .A2(new_n5813_), .B(new_n5917_), .ZN(new_n6318_));
  NOR3_X1    g06254(.A1(new_n5916_), .A2(new_n5818_), .A3(new_n5812_), .ZN(new_n6319_));
  OAI21_X1   g06255(.A1(new_n6319_), .A2(new_n6318_), .B(new_n5807_), .ZN(new_n6320_));
  OAI21_X1   g06256(.A1(new_n5914_), .A2(new_n5820_), .B(new_n5913_), .ZN(new_n6321_));
  OAI22_X1   g06257(.A1(new_n2103_), .A2(new_n4297_), .B1(new_n2158_), .B2(new_n4470_), .ZN(new_n6322_));
  NAND2_X1   g06258(.A1(new_n2107_), .A2(new_n4292_), .ZN(new_n6323_));
  AOI21_X1   g06259(.A1(new_n6322_), .A2(new_n6323_), .B(new_n4468_), .ZN(new_n6324_));
  NAND3_X1   g06260(.A1(new_n4959_), .A2(new_n3372_), .A3(new_n6324_), .ZN(new_n6325_));
  AOI21_X1   g06261(.A1(new_n4959_), .A2(new_n6324_), .B(new_n3372_), .ZN(new_n6326_));
  INV_X1     g06262(.I(new_n6326_), .ZN(new_n6327_));
  NAND2_X1   g06263(.A1(new_n6327_), .A2(new_n6325_), .ZN(new_n6328_));
  NAND3_X1   g06264(.A1(new_n6328_), .A2(new_n6320_), .A3(new_n6321_), .ZN(new_n6329_));
  NAND2_X1   g06265(.A1(new_n6320_), .A2(new_n6321_), .ZN(new_n6330_));
  INV_X1     g06266(.I(new_n6325_), .ZN(new_n6331_));
  NOR2_X1    g06267(.A1(new_n6331_), .A2(new_n6326_), .ZN(new_n6332_));
  NAND2_X1   g06268(.A1(new_n6330_), .A2(new_n6332_), .ZN(new_n6333_));
  NAND3_X1   g06269(.A1(new_n6333_), .A2(new_n6317_), .A3(new_n6329_), .ZN(new_n6334_));
  NOR3_X1    g06270(.A1(new_n6302_), .A2(new_n6295_), .A3(new_n6296_), .ZN(new_n6335_));
  NOR2_X1    g06271(.A1(new_n6330_), .A2(new_n6332_), .ZN(new_n6336_));
  AOI21_X1   g06272(.A1(new_n6320_), .A2(new_n6321_), .B(new_n6328_), .ZN(new_n6337_));
  OAI21_X1   g06273(.A1(new_n6336_), .A2(new_n6337_), .B(new_n6335_), .ZN(new_n6338_));
  NAND3_X1   g06274(.A1(new_n6315_), .A2(new_n6334_), .A3(new_n6338_), .ZN(new_n6339_));
  INV_X1     g06275(.I(new_n6314_), .ZN(new_n6340_));
  AOI22_X1   g06276(.A1(new_n6312_), .A2(new_n6340_), .B1(new_n6338_), .B2(new_n6334_), .ZN(new_n6341_));
  AOI21_X1   g06277(.A1(new_n6339_), .A2(new_n6308_), .B(new_n6341_), .ZN(new_n6342_));
  XOR2_X1    g06278(.A1(new_n5845_), .A2(new_n5831_), .Z(new_n6343_));
  NOR2_X1    g06279(.A1(new_n6343_), .A2(new_n5821_), .ZN(new_n6344_));
  NAND2_X1   g06280(.A1(new_n5922_), .A2(new_n5920_), .ZN(new_n6345_));
  AOI21_X1   g06281(.A1(new_n5821_), .A2(new_n6345_), .B(new_n6344_), .ZN(new_n6346_));
  OAI22_X1   g06282(.A1(new_n2103_), .A2(new_n4291_), .B1(new_n2198_), .B2(new_n4470_), .ZN(new_n6347_));
  NAND2_X1   g06283(.A1(new_n2161_), .A2(new_n4298_), .ZN(new_n6348_));
  AOI21_X1   g06284(.A1(new_n6347_), .A2(new_n6348_), .B(new_n4468_), .ZN(new_n6349_));
  NAND2_X1   g06285(.A1(new_n5351_), .A2(new_n6349_), .ZN(new_n6350_));
  XOR2_X1    g06286(.A1(new_n6350_), .A2(new_n3372_), .Z(new_n6351_));
  AOI21_X1   g06287(.A1(new_n6334_), .A2(new_n6333_), .B(new_n6351_), .ZN(new_n6352_));
  NOR3_X1    g06288(.A1(new_n6336_), .A2(new_n6337_), .A3(new_n6335_), .ZN(new_n6353_));
  INV_X1     g06289(.I(new_n6351_), .ZN(new_n6354_));
  NOR3_X1    g06290(.A1(new_n6353_), .A2(new_n6354_), .A3(new_n6337_), .ZN(new_n6355_));
  OAI21_X1   g06291(.A1(new_n6355_), .A2(new_n6352_), .B(new_n6346_), .ZN(new_n6356_));
  INV_X1     g06292(.I(new_n6346_), .ZN(new_n6357_));
  OAI21_X1   g06293(.A1(new_n6353_), .A2(new_n6337_), .B(new_n6354_), .ZN(new_n6358_));
  NAND3_X1   g06294(.A1(new_n6334_), .A2(new_n6333_), .A3(new_n6351_), .ZN(new_n6359_));
  NAND3_X1   g06295(.A1(new_n6358_), .A2(new_n6359_), .A3(new_n6357_), .ZN(new_n6360_));
  NAND2_X1   g06296(.A1(new_n6360_), .A2(new_n6356_), .ZN(new_n6361_));
  OAI22_X1   g06297(.A1(new_n2251_), .A2(new_n6091_), .B1(new_n4365_), .B2(new_n6094_), .ZN(new_n6362_));
  NAND2_X1   g06298(.A1(new_n1504_), .A2(new_n6180_), .ZN(new_n6363_));
  AOI21_X1   g06299(.A1(new_n6362_), .A2(new_n6363_), .B(new_n6082_), .ZN(new_n6364_));
  NAND2_X1   g06300(.A1(new_n4650_), .A2(new_n6364_), .ZN(new_n6365_));
  NOR2_X1    g06301(.A1(new_n6365_), .A2(\a[14] ), .ZN(new_n6366_));
  AOI21_X1   g06302(.A1(new_n4650_), .A2(new_n6364_), .B(new_n3521_), .ZN(new_n6367_));
  NOR2_X1    g06303(.A1(new_n6366_), .A2(new_n6367_), .ZN(new_n6368_));
  AOI21_X1   g06304(.A1(new_n6361_), .A2(new_n6368_), .B(new_n6342_), .ZN(new_n6369_));
  NOR2_X1    g06305(.A1(new_n6361_), .A2(new_n6368_), .ZN(new_n6370_));
  NAND3_X1   g06306(.A1(new_n5870_), .A2(new_n5878_), .A3(new_n5873_), .ZN(new_n6371_));
  NAND2_X1   g06307(.A1(new_n5981_), .A2(new_n6371_), .ZN(new_n6372_));
  OAI22_X1   g06308(.A1(new_n2311_), .A2(new_n6091_), .B1(new_n4365_), .B2(new_n6089_), .ZN(new_n6373_));
  NAND2_X1   g06309(.A1(new_n2255_), .A2(new_n6095_), .ZN(new_n6374_));
  AOI21_X1   g06310(.A1(new_n6373_), .A2(new_n6374_), .B(new_n6082_), .ZN(new_n6375_));
  NAND3_X1   g06311(.A1(new_n4419_), .A2(new_n3521_), .A3(new_n6375_), .ZN(new_n6376_));
  AOI21_X1   g06312(.A1(new_n4419_), .A2(new_n6375_), .B(new_n3521_), .ZN(new_n6377_));
  INV_X1     g06313(.I(new_n6377_), .ZN(new_n6378_));
  NAND3_X1   g06314(.A1(new_n6372_), .A2(new_n6378_), .A3(new_n6376_), .ZN(new_n6379_));
  OAI21_X1   g06315(.A1(new_n6369_), .A2(new_n6370_), .B(new_n6379_), .ZN(new_n6380_));
  NOR3_X1    g06316(.A1(new_n5980_), .A2(new_n5979_), .A3(new_n5869_), .ZN(new_n6381_));
  NOR2_X1    g06317(.A1(new_n5879_), .A2(new_n6381_), .ZN(new_n6382_));
  INV_X1     g06318(.I(new_n6376_), .ZN(new_n6383_));
  OAI21_X1   g06319(.A1(new_n6383_), .A2(new_n6377_), .B(new_n6382_), .ZN(new_n6384_));
  NAND2_X1   g06320(.A1(new_n6380_), .A2(new_n6384_), .ZN(new_n6385_));
  AOI21_X1   g06321(.A1(new_n5901_), .A2(new_n5926_), .B(new_n5984_), .ZN(new_n6386_));
  AOI21_X1   g06322(.A1(new_n5930_), .A2(new_n5932_), .B(new_n5983_), .ZN(new_n6387_));
  OAI21_X1   g06323(.A1(new_n6386_), .A2(new_n6387_), .B(new_n5879_), .ZN(new_n6388_));
  OAI21_X1   g06324(.A1(new_n5982_), .A2(new_n5934_), .B(new_n5981_), .ZN(new_n6389_));
  NAND2_X1   g06325(.A1(new_n6388_), .A2(new_n6389_), .ZN(new_n6390_));
  OAI22_X1   g06326(.A1(new_n2251_), .A2(new_n6089_), .B1(new_n2351_), .B2(new_n6091_), .ZN(new_n6391_));
  NAND2_X1   g06327(.A1(new_n2310_), .A2(new_n6095_), .ZN(new_n6392_));
  AOI21_X1   g06328(.A1(new_n6392_), .A2(new_n6391_), .B(new_n6082_), .ZN(new_n6393_));
  NAND3_X1   g06329(.A1(new_n3914_), .A2(new_n3521_), .A3(new_n6393_), .ZN(new_n6394_));
  INV_X1     g06330(.I(new_n6394_), .ZN(new_n6395_));
  AOI21_X1   g06331(.A1(new_n3914_), .A2(new_n6393_), .B(new_n3521_), .ZN(new_n6396_));
  NOR2_X1    g06332(.A1(new_n6395_), .A2(new_n6396_), .ZN(new_n6397_));
  NAND2_X1   g06333(.A1(new_n6390_), .A2(new_n6397_), .ZN(new_n6398_));
  NOR2_X1    g06334(.A1(new_n6390_), .A2(new_n6397_), .ZN(new_n6399_));
  AOI21_X1   g06335(.A1(new_n6385_), .A2(new_n6398_), .B(new_n6399_), .ZN(new_n6400_));
  NAND2_X1   g06336(.A1(new_n5989_), .A2(new_n5962_), .ZN(new_n6401_));
  NAND2_X1   g06337(.A1(new_n5954_), .A2(new_n5961_), .ZN(new_n6402_));
  AOI21_X1   g06338(.A1(new_n6401_), .A2(new_n6402_), .B(new_n5935_), .ZN(new_n6403_));
  NAND2_X1   g06339(.A1(new_n5954_), .A2(new_n5962_), .ZN(new_n6404_));
  AOI21_X1   g06340(.A1(new_n6404_), .A2(new_n5991_), .B(new_n5986_), .ZN(new_n6405_));
  NOR2_X1    g06341(.A1(new_n6403_), .A2(new_n6405_), .ZN(new_n6406_));
  OAI22_X1   g06342(.A1(new_n1453_), .A2(new_n6091_), .B1(new_n2351_), .B2(new_n6094_), .ZN(new_n6407_));
  NAND2_X1   g06343(.A1(new_n2310_), .A2(new_n6180_), .ZN(new_n6408_));
  AOI21_X1   g06344(.A1(new_n6408_), .A2(new_n6407_), .B(new_n6082_), .ZN(new_n6409_));
  NAND2_X1   g06345(.A1(new_n4231_), .A2(new_n6409_), .ZN(new_n6410_));
  XOR2_X1    g06346(.A1(new_n6410_), .A2(\a[14] ), .Z(new_n6411_));
  INV_X1     g06347(.I(new_n6411_), .ZN(new_n6412_));
  NOR2_X1    g06348(.A1(new_n6406_), .A2(new_n6412_), .ZN(new_n6413_));
  NAND2_X1   g06349(.A1(new_n6406_), .A2(new_n6412_), .ZN(new_n6414_));
  OAI21_X1   g06350(.A1(new_n6400_), .A2(new_n6413_), .B(new_n6414_), .ZN(new_n6415_));
  AOI22_X1   g06351(.A1(new_n6292_), .A2(new_n6288_), .B1(new_n6283_), .B2(new_n6284_), .ZN(new_n6416_));
  OAI21_X1   g06352(.A1(new_n6415_), .A2(new_n6416_), .B(new_n6293_), .ZN(new_n6417_));
  NAND3_X1   g06353(.A1(new_n6273_), .A2(new_n6277_), .A3(new_n6417_), .ZN(new_n6418_));
  OAI22_X1   g06354(.A1(new_n1409_), .A2(new_n6089_), .B1(new_n2367_), .B2(new_n6091_), .ZN(new_n6419_));
  NAND2_X1   g06355(.A1(new_n1334_), .A2(new_n6095_), .ZN(new_n6420_));
  AOI21_X1   g06356(.A1(new_n6419_), .A2(new_n6420_), .B(new_n6082_), .ZN(new_n6421_));
  NAND2_X1   g06357(.A1(new_n3654_), .A2(new_n6421_), .ZN(new_n6422_));
  XOR2_X1    g06358(.A1(new_n6422_), .A2(\a[14] ), .Z(new_n6423_));
  NAND2_X1   g06359(.A1(new_n6418_), .A2(new_n6423_), .ZN(new_n6424_));
  INV_X1     g06360(.I(new_n6423_), .ZN(new_n6425_));
  NAND4_X1   g06361(.A1(new_n6273_), .A2(new_n6277_), .A3(new_n6417_), .A4(new_n6425_), .ZN(new_n6426_));
  AOI21_X1   g06362(.A1(new_n6424_), .A2(new_n6426_), .B(new_n6257_), .ZN(new_n6427_));
  AOI21_X1   g06363(.A1(new_n6255_), .A2(new_n6254_), .B(new_n6253_), .ZN(new_n6428_));
  NOR3_X1    g06364(.A1(new_n6249_), .A2(new_n6251_), .A3(new_n6247_), .ZN(new_n6429_));
  NOR2_X1    g06365(.A1(new_n6428_), .A2(new_n6429_), .ZN(new_n6430_));
  AOI21_X1   g06366(.A1(new_n6276_), .A2(new_n6275_), .B(new_n6274_), .ZN(new_n6431_));
  NOR3_X1    g06367(.A1(new_n6269_), .A2(new_n6272_), .A3(new_n6262_), .ZN(new_n6432_));
  INV_X1     g06368(.I(new_n6293_), .ZN(new_n6433_));
  INV_X1     g06369(.I(new_n6308_), .ZN(new_n6434_));
  NAND2_X1   g06370(.A1(new_n6340_), .A2(new_n6312_), .ZN(new_n6435_));
  NAND2_X1   g06371(.A1(new_n6338_), .A2(new_n6334_), .ZN(new_n6436_));
  NOR2_X1    g06372(.A1(new_n6435_), .A2(new_n6436_), .ZN(new_n6437_));
  NAND2_X1   g06373(.A1(new_n6435_), .A2(new_n6436_), .ZN(new_n6438_));
  OAI21_X1   g06374(.A1(new_n6434_), .A2(new_n6437_), .B(new_n6438_), .ZN(new_n6439_));
  AOI21_X1   g06375(.A1(new_n6358_), .A2(new_n6359_), .B(new_n6357_), .ZN(new_n6440_));
  NOR3_X1    g06376(.A1(new_n6355_), .A2(new_n6352_), .A3(new_n6346_), .ZN(new_n6441_));
  NOR2_X1    g06377(.A1(new_n6440_), .A2(new_n6441_), .ZN(new_n6442_));
  XOR2_X1    g06378(.A1(new_n6365_), .A2(new_n3521_), .Z(new_n6443_));
  OAI21_X1   g06379(.A1(new_n6443_), .A2(new_n6442_), .B(new_n6439_), .ZN(new_n6444_));
  NAND2_X1   g06380(.A1(new_n6443_), .A2(new_n6442_), .ZN(new_n6445_));
  NAND2_X1   g06381(.A1(new_n6444_), .A2(new_n6445_), .ZN(new_n6446_));
  INV_X1     g06382(.I(new_n6384_), .ZN(new_n6447_));
  AOI21_X1   g06383(.A1(new_n6446_), .A2(new_n6379_), .B(new_n6447_), .ZN(new_n6448_));
  INV_X1     g06384(.I(new_n6396_), .ZN(new_n6449_));
  NAND2_X1   g06385(.A1(new_n6449_), .A2(new_n6394_), .ZN(new_n6450_));
  AOI21_X1   g06386(.A1(new_n6388_), .A2(new_n6389_), .B(new_n6450_), .ZN(new_n6451_));
  NAND3_X1   g06387(.A1(new_n6450_), .A2(new_n6388_), .A3(new_n6389_), .ZN(new_n6452_));
  OAI21_X1   g06388(.A1(new_n6448_), .A2(new_n6451_), .B(new_n6452_), .ZN(new_n6453_));
  OAI21_X1   g06389(.A1(new_n6403_), .A2(new_n6405_), .B(new_n6411_), .ZN(new_n6454_));
  NOR3_X1    g06390(.A1(new_n6411_), .A2(new_n6403_), .A3(new_n6405_), .ZN(new_n6455_));
  AOI21_X1   g06391(.A1(new_n6453_), .A2(new_n6454_), .B(new_n6455_), .ZN(new_n6456_));
  NAND2_X1   g06392(.A1(new_n6283_), .A2(new_n6284_), .ZN(new_n6457_));
  INV_X1     g06393(.I(new_n6288_), .ZN(new_n6458_));
  AOI21_X1   g06394(.A1(new_n6289_), .A2(new_n6290_), .B(new_n6042_), .ZN(new_n6459_));
  OAI21_X1   g06395(.A1(new_n6458_), .A2(new_n6459_), .B(new_n6457_), .ZN(new_n6460_));
  AOI21_X1   g06396(.A1(new_n6456_), .A2(new_n6460_), .B(new_n6433_), .ZN(new_n6461_));
  NOR3_X1    g06397(.A1(new_n6432_), .A2(new_n6431_), .A3(new_n6461_), .ZN(new_n6462_));
  NOR2_X1    g06398(.A1(new_n6462_), .A2(new_n6425_), .ZN(new_n6463_));
  INV_X1     g06399(.I(new_n6426_), .ZN(new_n6464_));
  NOR3_X1    g06400(.A1(new_n6463_), .A2(new_n6464_), .A3(new_n6430_), .ZN(new_n6465_));
  NOR3_X1    g06401(.A1(new_n6465_), .A2(new_n6427_), .A3(new_n6246_), .ZN(new_n6466_));
  XOR2_X1    g06402(.A1(new_n6245_), .A2(new_n4034_), .Z(new_n6467_));
  OAI21_X1   g06403(.A1(new_n6463_), .A2(new_n6464_), .B(new_n6430_), .ZN(new_n6468_));
  NAND3_X1   g06404(.A1(new_n6424_), .A2(new_n6257_), .A3(new_n6426_), .ZN(new_n6469_));
  AOI21_X1   g06405(.A1(new_n6468_), .A2(new_n6469_), .B(new_n6467_), .ZN(new_n6470_));
  OAI22_X1   g06406(.A1(new_n2367_), .A2(new_n4716_), .B1(new_n2451_), .B2(new_n4710_), .ZN(new_n6471_));
  NAND2_X1   g06407(.A1(new_n2412_), .A2(new_n4720_), .ZN(new_n6472_));
  AOI21_X1   g06408(.A1(new_n6471_), .A2(new_n6472_), .B(new_n4707_), .ZN(new_n6473_));
  NAND2_X1   g06409(.A1(new_n3403_), .A2(new_n6473_), .ZN(new_n6474_));
  XOR2_X1    g06410(.A1(new_n6474_), .A2(\a[11] ), .Z(new_n6475_));
  NAND3_X1   g06411(.A1(new_n6273_), .A2(new_n6277_), .A3(new_n6461_), .ZN(new_n6476_));
  OAI21_X1   g06412(.A1(new_n6432_), .A2(new_n6431_), .B(new_n6417_), .ZN(new_n6477_));
  NAND2_X1   g06413(.A1(new_n6477_), .A2(new_n6476_), .ZN(new_n6478_));
  OAI22_X1   g06414(.A1(new_n2367_), .A2(new_n4719_), .B1(new_n2408_), .B2(new_n4710_), .ZN(new_n6479_));
  INV_X1     g06415(.I(new_n4716_), .ZN(new_n6480_));
  NAND2_X1   g06416(.A1(new_n1334_), .A2(new_n6480_), .ZN(new_n6481_));
  AOI21_X1   g06417(.A1(new_n6479_), .A2(new_n6481_), .B(new_n4707_), .ZN(new_n6482_));
  AND3_X2    g06418(.A1(new_n3708_), .A2(new_n4034_), .A3(new_n6482_), .Z(new_n6483_));
  AOI21_X1   g06419(.A1(new_n3708_), .A2(new_n6482_), .B(new_n4034_), .ZN(new_n6484_));
  NOR2_X1    g06420(.A1(new_n6483_), .A2(new_n6484_), .ZN(new_n6485_));
  NAND2_X1   g06421(.A1(new_n6460_), .A2(new_n6293_), .ZN(new_n6486_));
  XOR2_X1    g06422(.A1(new_n6486_), .A2(new_n6415_), .Z(new_n6487_));
  NOR2_X1    g06423(.A1(new_n6487_), .A2(new_n6485_), .ZN(new_n6488_));
  AOI21_X1   g06424(.A1(new_n6478_), .A2(new_n6475_), .B(new_n6488_), .ZN(new_n6489_));
  OAI22_X1   g06425(.A1(new_n6470_), .A2(new_n6466_), .B1(new_n6246_), .B2(new_n6489_), .ZN(new_n6490_));
  NOR2_X1    g06426(.A1(new_n6226_), .A2(new_n6190_), .ZN(new_n6491_));
  XOR2_X1    g06427(.A1(new_n6239_), .A2(new_n4034_), .Z(new_n6492_));
  NOR2_X1    g06428(.A1(new_n6492_), .A2(new_n6491_), .ZN(new_n6493_));
  NOR2_X1    g06429(.A1(new_n6241_), .A2(new_n6493_), .ZN(new_n6494_));
  AOI21_X1   g06430(.A1(new_n6490_), .A2(new_n6494_), .B(new_n6241_), .ZN(new_n6495_));
  NOR3_X1    g06431(.A1(new_n6495_), .A2(new_n6231_), .A3(new_n6235_), .ZN(new_n6496_));
  OAI21_X1   g06432(.A1(new_n6496_), .A2(new_n6157_), .B(new_n6218_), .ZN(new_n6497_));
  INV_X1     g06433(.I(new_n6148_), .ZN(new_n6498_));
  NAND2_X1   g06434(.A1(new_n6498_), .A2(new_n6114_), .ZN(new_n6499_));
  NOR2_X1    g06435(.A1(new_n6499_), .A2(new_n6146_), .ZN(new_n6500_));
  NOR2_X1    g06436(.A1(new_n6150_), .A2(new_n6500_), .ZN(new_n6501_));
  AOI21_X1   g06437(.A1(new_n6497_), .A2(new_n6501_), .B(new_n6150_), .ZN(new_n6502_));
  NOR3_X1    g06438(.A1(new_n6502_), .A2(new_n6140_), .A3(new_n6131_), .ZN(new_n6503_));
  NAND2_X1   g06439(.A1(new_n5221_), .A2(new_n4737_), .ZN(new_n6504_));
  XOR2_X1    g06440(.A1(new_n4965_), .A2(new_n5223_), .Z(new_n6505_));
  OAI21_X1   g06441(.A1(new_n5221_), .A2(new_n4737_), .B(new_n6505_), .ZN(new_n6506_));
  NAND2_X1   g06442(.A1(new_n6506_), .A2(new_n6504_), .ZN(new_n6507_));
  INV_X1     g06443(.I(new_n6507_), .ZN(new_n6508_));
  INV_X1     g06444(.I(new_n4953_), .ZN(new_n6509_));
  INV_X1     g06445(.I(new_n4964_), .ZN(new_n6510_));
  NAND2_X1   g06446(.A1(new_n6510_), .A2(new_n6509_), .ZN(new_n6511_));
  NOR2_X1    g06447(.A1(new_n6510_), .A2(new_n6509_), .ZN(new_n6512_));
  AOI21_X1   g06448(.A1(new_n5223_), .A2(new_n6511_), .B(new_n6512_), .ZN(new_n6513_));
  NAND2_X1   g06449(.A1(new_n4910_), .A2(new_n4947_), .ZN(new_n6514_));
  NAND2_X1   g06450(.A1(new_n6514_), .A2(new_n4949_), .ZN(new_n6515_));
  NOR2_X1    g06451(.A1(new_n2071_), .A2(new_n2772_), .ZN(new_n6516_));
  NOR2_X1    g06452(.A1(new_n1612_), .A2(new_n2771_), .ZN(new_n6517_));
  NOR2_X1    g06453(.A1(new_n1678_), .A2(new_n2767_), .ZN(new_n6518_));
  NOR4_X1    g06454(.A1(new_n6518_), .A2(new_n6517_), .A3(new_n6516_), .A4(new_n2763_), .ZN(new_n6519_));
  NAND2_X1   g06455(.A1(new_n5070_), .A2(new_n6519_), .ZN(new_n6520_));
  INV_X1     g06456(.I(new_n3440_), .ZN(new_n6521_));
  NOR4_X1    g06457(.A1(new_n239_), .A2(new_n640_), .A3(new_n817_), .A4(new_n1073_), .ZN(new_n6522_));
  INV_X1     g06458(.I(new_n6522_), .ZN(new_n6523_));
  NAND3_X1   g06459(.A1(new_n6523_), .A2(new_n269_), .A3(new_n2781_), .ZN(new_n6524_));
  NOR4_X1    g06460(.A1(new_n3944_), .A2(new_n124_), .A3(new_n242_), .A4(new_n560_), .ZN(new_n6525_));
  INV_X1     g06461(.I(new_n6525_), .ZN(new_n6526_));
  NOR4_X1    g06462(.A1(new_n1151_), .A2(new_n4377_), .A3(new_n1045_), .A4(new_n1995_), .ZN(new_n6527_));
  NOR3_X1    g06463(.A1(new_n945_), .A2(new_n92_), .A3(new_n173_), .ZN(new_n6528_));
  NAND4_X1   g06464(.A1(new_n6528_), .A2(new_n707_), .A3(new_n807_), .A4(new_n765_), .ZN(new_n6529_));
  INV_X1     g06465(.I(new_n6529_), .ZN(new_n6530_));
  NAND2_X1   g06466(.A1(new_n6530_), .A2(new_n6527_), .ZN(new_n6531_));
  NOR4_X1    g06467(.A1(new_n6521_), .A2(new_n6524_), .A3(new_n6526_), .A4(new_n6531_), .ZN(new_n6532_));
  NAND4_X1   g06468(.A1(new_n1091_), .A2(new_n1403_), .A3(new_n1506_), .A4(new_n1448_), .ZN(new_n6533_));
  NAND2_X1   g06469(.A1(new_n1205_), .A2(new_n1319_), .ZN(new_n6534_));
  NAND3_X1   g06470(.A1(new_n1840_), .A2(new_n469_), .A3(new_n1067_), .ZN(new_n6535_));
  NAND4_X1   g06471(.A1(new_n6535_), .A2(new_n1311_), .A3(new_n1454_), .A4(new_n676_), .ZN(new_n6536_));
  NAND4_X1   g06472(.A1(new_n3489_), .A2(new_n389_), .A3(new_n1460_), .A4(new_n3459_), .ZN(new_n6537_));
  NOR4_X1    g06473(.A1(new_n6537_), .A2(new_n6533_), .A3(new_n6534_), .A4(new_n6536_), .ZN(new_n6538_));
  AND2_X2    g06474(.A1(new_n6538_), .A2(new_n2242_), .Z(new_n6539_));
  NAND3_X1   g06475(.A1(new_n6532_), .A2(new_n3458_), .A3(new_n6539_), .ZN(new_n6540_));
  AND2_X2    g06476(.A1(new_n6520_), .A2(new_n6540_), .Z(new_n6541_));
  NOR2_X1    g06477(.A1(new_n6520_), .A2(new_n6540_), .ZN(new_n6542_));
  OAI21_X1   g06478(.A1(new_n6541_), .A2(new_n6542_), .B(new_n6515_), .ZN(new_n6543_));
  XOR2_X1    g06479(.A1(new_n6520_), .A2(new_n6540_), .Z(new_n6544_));
  NAND3_X1   g06480(.A1(new_n6544_), .A2(new_n6514_), .A3(new_n4949_), .ZN(new_n6545_));
  NAND2_X1   g06481(.A1(new_n6543_), .A2(new_n6545_), .ZN(new_n6546_));
  OAI22_X1   g06482(.A1(new_n2103_), .A2(new_n2747_), .B1(new_n2198_), .B2(new_n3175_), .ZN(new_n6547_));
  NAND2_X1   g06483(.A1(new_n2161_), .A2(new_n3275_), .ZN(new_n6548_));
  AOI21_X1   g06484(.A1(new_n6547_), .A2(new_n6548_), .B(new_n2737_), .ZN(new_n6549_));
  NAND2_X1   g06485(.A1(new_n5351_), .A2(new_n6549_), .ZN(new_n6550_));
  XOR2_X1    g06486(.A1(new_n6550_), .A2(\a[29] ), .Z(new_n6551_));
  XOR2_X1    g06487(.A1(new_n6551_), .A2(new_n6546_), .Z(new_n6552_));
  OR2_X2     g06488(.A1(new_n6552_), .A2(new_n6513_), .Z(new_n6553_));
  INV_X1     g06489(.I(new_n6551_), .ZN(new_n6554_));
  NOR2_X1    g06490(.A1(new_n6554_), .A2(new_n6546_), .ZN(new_n6555_));
  NAND2_X1   g06491(.A1(new_n6554_), .A2(new_n6546_), .ZN(new_n6556_));
  INV_X1     g06492(.I(new_n6556_), .ZN(new_n6557_));
  OAI21_X1   g06493(.A1(new_n6557_), .A2(new_n6555_), .B(new_n6513_), .ZN(new_n6558_));
  NAND2_X1   g06494(.A1(new_n6553_), .A2(new_n6558_), .ZN(new_n6559_));
  OAI22_X1   g06495(.A1(new_n2251_), .A2(new_n3318_), .B1(new_n4365_), .B2(new_n3322_), .ZN(new_n6560_));
  NAND2_X1   g06496(.A1(new_n1504_), .A2(new_n3267_), .ZN(new_n6561_));
  AOI21_X1   g06497(.A1(new_n6560_), .A2(new_n6561_), .B(new_n3260_), .ZN(new_n6562_));
  NAND2_X1   g06498(.A1(new_n4650_), .A2(new_n6562_), .ZN(new_n6563_));
  XOR2_X1    g06499(.A1(new_n6563_), .A2(\a[26] ), .Z(new_n6564_));
  NAND2_X1   g06500(.A1(new_n6559_), .A2(new_n6564_), .ZN(new_n6565_));
  INV_X1     g06501(.I(new_n6559_), .ZN(new_n6566_));
  INV_X1     g06502(.I(new_n6564_), .ZN(new_n6567_));
  NAND2_X1   g06503(.A1(new_n6566_), .A2(new_n6567_), .ZN(new_n6568_));
  AOI21_X1   g06504(.A1(new_n6568_), .A2(new_n6565_), .B(new_n6508_), .ZN(new_n6569_));
  NAND2_X1   g06505(.A1(new_n6566_), .A2(new_n6564_), .ZN(new_n6570_));
  NAND2_X1   g06506(.A1(new_n6567_), .A2(new_n6559_), .ZN(new_n6571_));
  AOI21_X1   g06507(.A1(new_n6570_), .A2(new_n6571_), .B(new_n6507_), .ZN(new_n6572_));
  NOR2_X1    g06508(.A1(new_n6569_), .A2(new_n6572_), .ZN(new_n6573_));
  INV_X1     g06509(.I(new_n6573_), .ZN(new_n6574_));
  OAI22_X1   g06510(.A1(new_n1453_), .A2(new_n3780_), .B1(new_n2351_), .B2(new_n3306_), .ZN(new_n6575_));
  NAND2_X1   g06511(.A1(new_n2310_), .A2(new_n5291_), .ZN(new_n6576_));
  AOI21_X1   g06512(.A1(new_n6576_), .A2(new_n6575_), .B(new_n3302_), .ZN(new_n6577_));
  NAND2_X1   g06513(.A1(new_n4231_), .A2(new_n6577_), .ZN(new_n6578_));
  XOR2_X1    g06514(.A1(new_n6578_), .A2(\a[23] ), .Z(new_n6579_));
  INV_X1     g06515(.I(new_n6579_), .ZN(new_n6580_));
  NAND3_X1   g06516(.A1(new_n5509_), .A2(new_n5507_), .A3(new_n5504_), .ZN(new_n6581_));
  AOI21_X1   g06517(.A1(new_n6581_), .A2(new_n5507_), .B(new_n6580_), .ZN(new_n6582_));
  INV_X1     g06518(.I(new_n6582_), .ZN(new_n6583_));
  NAND3_X1   g06519(.A1(new_n6581_), .A2(new_n6580_), .A3(new_n5507_), .ZN(new_n6584_));
  AOI21_X1   g06520(.A1(new_n6583_), .A2(new_n6584_), .B(new_n6574_), .ZN(new_n6585_));
  INV_X1     g06521(.I(new_n6584_), .ZN(new_n6586_));
  NOR3_X1    g06522(.A1(new_n6586_), .A2(new_n6573_), .A3(new_n6582_), .ZN(new_n6587_));
  NOR2_X1    g06523(.A1(new_n6585_), .A2(new_n6587_), .ZN(new_n6588_));
  INV_X1     g06524(.I(new_n6588_), .ZN(new_n6589_));
  NAND2_X1   g06525(.A1(new_n5601_), .A2(new_n5542_), .ZN(new_n6590_));
  OAI22_X1   g06526(.A1(new_n1409_), .A2(new_n3769_), .B1(new_n2367_), .B2(new_n4097_), .ZN(new_n6591_));
  NAND2_X1   g06527(.A1(new_n1334_), .A2(new_n3776_), .ZN(new_n6592_));
  AOI21_X1   g06528(.A1(new_n6591_), .A2(new_n6592_), .B(new_n4095_), .ZN(new_n6593_));
  NAND2_X1   g06529(.A1(new_n3654_), .A2(new_n6593_), .ZN(new_n6594_));
  XOR2_X1    g06530(.A1(new_n6594_), .A2(\a[20] ), .Z(new_n6595_));
  NAND2_X1   g06531(.A1(new_n6590_), .A2(new_n6595_), .ZN(new_n6596_));
  NOR2_X1    g06532(.A1(new_n6024_), .A2(new_n5602_), .ZN(new_n6597_));
  INV_X1     g06533(.I(new_n6595_), .ZN(new_n6598_));
  NAND2_X1   g06534(.A1(new_n6597_), .A2(new_n6598_), .ZN(new_n6599_));
  AOI21_X1   g06535(.A1(new_n6596_), .A2(new_n6599_), .B(new_n6589_), .ZN(new_n6600_));
  NOR2_X1    g06536(.A1(new_n6597_), .A2(new_n6598_), .ZN(new_n6601_));
  NOR2_X1    g06537(.A1(new_n6590_), .A2(new_n6595_), .ZN(new_n6602_));
  NOR3_X1    g06538(.A1(new_n6601_), .A2(new_n6602_), .A3(new_n6588_), .ZN(new_n6603_));
  NOR2_X1    g06539(.A1(new_n6600_), .A2(new_n6603_), .ZN(new_n6604_));
  OAI22_X1   g06540(.A1(new_n2492_), .A2(new_n4470_), .B1(new_n2408_), .B2(new_n4291_), .ZN(new_n6605_));
  NAND2_X1   g06541(.A1(new_n2454_), .A2(new_n4298_), .ZN(new_n6606_));
  AOI21_X1   g06542(.A1(new_n6606_), .A2(new_n6605_), .B(new_n4468_), .ZN(new_n6607_));
  NAND2_X1   g06543(.A1(new_n3577_), .A2(new_n6607_), .ZN(new_n6608_));
  XOR2_X1    g06544(.A1(new_n6608_), .A2(\a[17] ), .Z(new_n6609_));
  INV_X1     g06545(.I(new_n6609_), .ZN(new_n6610_));
  NOR2_X1    g06546(.A1(new_n6104_), .A2(new_n6057_), .ZN(new_n6611_));
  NOR4_X1    g06547(.A1(new_n6611_), .A2(new_n6030_), .A3(new_n6064_), .A4(new_n6105_), .ZN(new_n6612_));
  XOR2_X1    g06548(.A1(new_n6612_), .A2(new_n6610_), .Z(new_n6613_));
  XOR2_X1    g06549(.A1(new_n6613_), .A2(new_n6604_), .Z(new_n6614_));
  OAI22_X1   g06550(.A1(new_n1008_), .A2(new_n6091_), .B1(new_n1121_), .B2(new_n6089_), .ZN(new_n6615_));
  NAND2_X1   g06551(.A1(new_n1181_), .A2(new_n6095_), .ZN(new_n6616_));
  AOI21_X1   g06552(.A1(new_n6615_), .A2(new_n6616_), .B(new_n6082_), .ZN(new_n6617_));
  NAND2_X1   g06553(.A1(new_n3562_), .A2(new_n6617_), .ZN(new_n6618_));
  XOR2_X1    g06554(.A1(new_n6618_), .A2(\a[14] ), .Z(new_n6619_));
  INV_X1     g06555(.I(new_n6619_), .ZN(new_n6620_));
  AOI21_X1   g06556(.A1(new_n6132_), .A2(new_n6121_), .B(new_n6620_), .ZN(new_n6621_));
  INV_X1     g06557(.I(new_n6621_), .ZN(new_n6622_));
  NAND3_X1   g06558(.A1(new_n6132_), .A2(new_n6620_), .A3(new_n6121_), .ZN(new_n6623_));
  AOI21_X1   g06559(.A1(new_n6622_), .A2(new_n6623_), .B(new_n6614_), .ZN(new_n6624_));
  XNOR2_X1   g06560(.A1(new_n6613_), .A2(new_n6604_), .ZN(new_n6625_));
  NOR3_X1    g06561(.A1(new_n6120_), .A2(new_n6619_), .A3(new_n6100_), .ZN(new_n6626_));
  NOR3_X1    g06562(.A1(new_n6625_), .A2(new_n6621_), .A3(new_n6626_), .ZN(new_n6627_));
  NOR3_X1    g06563(.A1(new_n6624_), .A2(new_n6627_), .A3(new_n4724_), .ZN(new_n6628_));
  OAI21_X1   g06564(.A1(new_n6621_), .A2(new_n6626_), .B(new_n6625_), .ZN(new_n6629_));
  NAND3_X1   g06565(.A1(new_n6622_), .A2(new_n6614_), .A3(new_n6623_), .ZN(new_n6630_));
  INV_X1     g06566(.I(new_n4724_), .ZN(new_n6631_));
  AOI21_X1   g06567(.A1(new_n6629_), .A2(new_n6630_), .B(new_n6631_), .ZN(new_n6632_));
  OAI22_X1   g06568(.A1(new_n6632_), .A2(new_n6628_), .B1(new_n6503_), .B2(new_n4724_), .ZN(new_n6633_));
  NOR2_X1    g06569(.A1(new_n2559_), .A2(new_n4719_), .ZN(new_n6634_));
  OAI22_X1   g06570(.A1(new_n813_), .A2(new_n4716_), .B1(new_n529_), .B2(new_n4710_), .ZN(new_n6635_));
  NOR3_X1    g06571(.A1(new_n6634_), .A2(new_n4707_), .A3(new_n6635_), .ZN(new_n6636_));
  NAND2_X1   g06572(.A1(new_n3051_), .A2(new_n6636_), .ZN(new_n6637_));
  INV_X1     g06573(.I(new_n6637_), .ZN(new_n6638_));
  NOR3_X1    g06574(.A1(new_n6600_), .A2(new_n6603_), .A3(new_n6609_), .ZN(new_n6639_));
  OAI21_X1   g06575(.A1(new_n6601_), .A2(new_n6602_), .B(new_n6588_), .ZN(new_n6640_));
  NAND3_X1   g06576(.A1(new_n6589_), .A2(new_n6599_), .A3(new_n6596_), .ZN(new_n6641_));
  AOI21_X1   g06577(.A1(new_n6641_), .A2(new_n6640_), .B(new_n6610_), .ZN(new_n6642_));
  OAI22_X1   g06578(.A1(new_n6639_), .A2(new_n6642_), .B1(new_n6609_), .B2(new_n6612_), .ZN(new_n6643_));
  INV_X1     g06579(.I(new_n6581_), .ZN(new_n6644_));
  NOR3_X1    g06580(.A1(new_n6569_), .A2(new_n6572_), .A3(new_n6579_), .ZN(new_n6645_));
  NOR2_X1    g06581(.A1(new_n6573_), .A2(new_n6580_), .ZN(new_n6646_));
  OAI21_X1   g06582(.A1(new_n6646_), .A2(new_n6645_), .B(new_n5507_), .ZN(new_n6647_));
  OAI22_X1   g06583(.A1(new_n6647_), .A2(new_n6644_), .B1(new_n6573_), .B2(new_n6580_), .ZN(new_n6648_));
  INV_X1     g06584(.I(new_n6648_), .ZN(new_n6649_));
  NAND2_X1   g06585(.A1(new_n6565_), .A2(new_n6507_), .ZN(new_n6650_));
  NAND2_X1   g06586(.A1(new_n6650_), .A2(new_n6568_), .ZN(new_n6651_));
  OAI21_X1   g06587(.A1(new_n6513_), .A2(new_n6555_), .B(new_n6556_), .ZN(new_n6652_));
  INV_X1     g06588(.I(new_n6652_), .ZN(new_n6653_));
  OAI22_X1   g06589(.A1(new_n2158_), .A2(new_n2747_), .B1(new_n2198_), .B2(new_n2742_), .ZN(new_n6654_));
  NAND2_X1   g06590(.A1(new_n1504_), .A2(new_n2750_), .ZN(new_n6655_));
  AOI21_X1   g06591(.A1(new_n6655_), .A2(new_n6654_), .B(new_n2737_), .ZN(new_n6656_));
  NAND3_X1   g06592(.A1(new_n4620_), .A2(new_n74_), .A3(new_n6656_), .ZN(new_n6657_));
  AOI21_X1   g06593(.A1(new_n4620_), .A2(new_n6656_), .B(new_n74_), .ZN(new_n6658_));
  INV_X1     g06594(.I(new_n6658_), .ZN(new_n6659_));
  NAND2_X1   g06595(.A1(new_n6659_), .A2(new_n6657_), .ZN(new_n6660_));
  AOI21_X1   g06596(.A1(new_n6514_), .A2(new_n4949_), .B(new_n6541_), .ZN(new_n6661_));
  NOR2_X1    g06597(.A1(new_n6661_), .A2(new_n6542_), .ZN(new_n6662_));
  INV_X1     g06598(.I(new_n4569_), .ZN(new_n6663_));
  NAND2_X1   g06599(.A1(new_n6663_), .A2(new_n4570_), .ZN(new_n6664_));
  NAND3_X1   g06600(.A1(new_n4545_), .A2(new_n4549_), .A3(new_n6664_), .ZN(new_n6665_));
  XOR2_X1    g06601(.A1(new_n4568_), .A2(new_n4387_), .Z(new_n6666_));
  NAND2_X1   g06602(.A1(new_n4550_), .A2(new_n6666_), .ZN(new_n6667_));
  NAND2_X1   g06603(.A1(new_n6667_), .A2(new_n6665_), .ZN(new_n6668_));
  INV_X1     g06604(.I(new_n6668_), .ZN(new_n6669_));
  XOR2_X1    g06605(.A1(new_n6662_), .A2(new_n6669_), .Z(new_n6670_));
  NOR3_X1    g06606(.A1(new_n6661_), .A2(new_n6542_), .A3(new_n6668_), .ZN(new_n6671_));
  NOR2_X1    g06607(.A1(new_n6662_), .A2(new_n6669_), .ZN(new_n6672_));
  NOR2_X1    g06608(.A1(new_n6672_), .A2(new_n6671_), .ZN(new_n6673_));
  NOR2_X1    g06609(.A1(new_n6660_), .A2(new_n6673_), .ZN(new_n6674_));
  AOI21_X1   g06610(.A1(new_n6660_), .A2(new_n6670_), .B(new_n6674_), .ZN(new_n6675_));
  OAI22_X1   g06611(.A1(new_n2311_), .A2(new_n3318_), .B1(new_n4365_), .B2(new_n3268_), .ZN(new_n6676_));
  NAND2_X1   g06612(.A1(new_n2255_), .A2(new_n3323_), .ZN(new_n6677_));
  AOI21_X1   g06613(.A1(new_n6676_), .A2(new_n6677_), .B(new_n3260_), .ZN(new_n6678_));
  NAND3_X1   g06614(.A1(new_n4419_), .A2(new_n72_), .A3(new_n6678_), .ZN(new_n6679_));
  AOI21_X1   g06615(.A1(new_n4419_), .A2(new_n6678_), .B(new_n72_), .ZN(new_n6680_));
  INV_X1     g06616(.I(new_n6680_), .ZN(new_n6681_));
  NAND3_X1   g06617(.A1(new_n6681_), .A2(new_n6675_), .A3(new_n6679_), .ZN(new_n6682_));
  NAND2_X1   g06618(.A1(new_n6670_), .A2(new_n6660_), .ZN(new_n6683_));
  OAI21_X1   g06619(.A1(new_n6660_), .A2(new_n6673_), .B(new_n6683_), .ZN(new_n6684_));
  INV_X1     g06620(.I(new_n6679_), .ZN(new_n6685_));
  OAI21_X1   g06621(.A1(new_n6685_), .A2(new_n6680_), .B(new_n6684_), .ZN(new_n6686_));
  AOI21_X1   g06622(.A1(new_n6686_), .A2(new_n6682_), .B(new_n6653_), .ZN(new_n6687_));
  NAND3_X1   g06623(.A1(new_n6681_), .A2(new_n6684_), .A3(new_n6679_), .ZN(new_n6688_));
  OAI21_X1   g06624(.A1(new_n6685_), .A2(new_n6680_), .B(new_n6675_), .ZN(new_n6689_));
  AOI21_X1   g06625(.A1(new_n6688_), .A2(new_n6689_), .B(new_n6652_), .ZN(new_n6690_));
  NOR2_X1    g06626(.A1(new_n6687_), .A2(new_n6690_), .ZN(new_n6691_));
  INV_X1     g06627(.I(new_n6691_), .ZN(new_n6692_));
  OAI22_X1   g06628(.A1(new_n1409_), .A2(new_n3780_), .B1(new_n2351_), .B2(new_n3310_), .ZN(new_n6693_));
  NAND2_X1   g06629(.A1(new_n2359_), .A2(new_n3782_), .ZN(new_n6694_));
  AOI21_X1   g06630(.A1(new_n6693_), .A2(new_n6694_), .B(new_n3302_), .ZN(new_n6695_));
  NAND2_X1   g06631(.A1(new_n3904_), .A2(new_n6695_), .ZN(new_n6696_));
  NOR2_X1    g06632(.A1(new_n6696_), .A2(\a[23] ), .ZN(new_n6697_));
  NAND2_X1   g06633(.A1(new_n6696_), .A2(\a[23] ), .ZN(new_n6698_));
  INV_X1     g06634(.I(new_n6698_), .ZN(new_n6699_));
  NOR3_X1    g06635(.A1(new_n6692_), .A2(new_n6699_), .A3(new_n6697_), .ZN(new_n6700_));
  INV_X1     g06636(.I(new_n6697_), .ZN(new_n6701_));
  AOI21_X1   g06637(.A1(new_n6701_), .A2(new_n6698_), .B(new_n6691_), .ZN(new_n6702_));
  OAI21_X1   g06638(.A1(new_n6700_), .A2(new_n6702_), .B(new_n6651_), .ZN(new_n6703_));
  INV_X1     g06639(.I(new_n6703_), .ZN(new_n6704_));
  NAND3_X1   g06640(.A1(new_n6692_), .A2(new_n6701_), .A3(new_n6698_), .ZN(new_n6705_));
  OAI21_X1   g06641(.A1(new_n6699_), .A2(new_n6697_), .B(new_n6691_), .ZN(new_n6706_));
  AOI21_X1   g06642(.A1(new_n6705_), .A2(new_n6706_), .B(new_n6651_), .ZN(new_n6707_));
  NOR2_X1    g06643(.A1(new_n6704_), .A2(new_n6707_), .ZN(new_n6708_));
  OAI22_X1   g06644(.A1(new_n2367_), .A2(new_n3775_), .B1(new_n2408_), .B2(new_n4097_), .ZN(new_n6709_));
  NAND2_X1   g06645(.A1(new_n1334_), .A2(new_n3770_), .ZN(new_n6710_));
  AOI21_X1   g06646(.A1(new_n6709_), .A2(new_n6710_), .B(new_n4095_), .ZN(new_n6711_));
  NAND3_X1   g06647(.A1(new_n3708_), .A2(new_n3035_), .A3(new_n6711_), .ZN(new_n6712_));
  AOI21_X1   g06648(.A1(new_n3708_), .A2(new_n6711_), .B(new_n3035_), .ZN(new_n6713_));
  INV_X1     g06649(.I(new_n6713_), .ZN(new_n6714_));
  NAND3_X1   g06650(.A1(new_n6708_), .A2(new_n6712_), .A3(new_n6714_), .ZN(new_n6715_));
  INV_X1     g06651(.I(new_n6707_), .ZN(new_n6716_));
  AOI22_X1   g06652(.A1(new_n6712_), .A2(new_n6714_), .B1(new_n6716_), .B2(new_n6703_), .ZN(new_n6717_));
  INV_X1     g06653(.I(new_n6717_), .ZN(new_n6718_));
  AOI21_X1   g06654(.A1(new_n6718_), .A2(new_n6715_), .B(new_n6649_), .ZN(new_n6719_));
  NAND2_X1   g06655(.A1(new_n6716_), .A2(new_n6703_), .ZN(new_n6720_));
  NAND3_X1   g06656(.A1(new_n6720_), .A2(new_n6712_), .A3(new_n6714_), .ZN(new_n6721_));
  INV_X1     g06657(.I(new_n6712_), .ZN(new_n6722_));
  OAI21_X1   g06658(.A1(new_n6722_), .A2(new_n6713_), .B(new_n6708_), .ZN(new_n6723_));
  AOI21_X1   g06659(.A1(new_n6723_), .A2(new_n6721_), .B(new_n6648_), .ZN(new_n6724_));
  NOR2_X1    g06660(.A1(new_n6719_), .A2(new_n6724_), .ZN(new_n6725_));
  AOI21_X1   g06661(.A1(new_n2496_), .A2(new_n4298_), .B(new_n4468_), .ZN(new_n6726_));
  AOI22_X1   g06662(.A1(new_n1122_), .A2(new_n4469_), .B1(new_n2454_), .B2(new_n4292_), .ZN(new_n6727_));
  NAND3_X1   g06663(.A1(new_n3393_), .A2(new_n6726_), .A3(new_n6727_), .ZN(new_n6728_));
  XOR2_X1    g06664(.A1(new_n6728_), .A2(new_n3372_), .Z(new_n6729_));
  NOR2_X1    g06665(.A1(new_n6725_), .A2(new_n6729_), .ZN(new_n6730_));
  NOR3_X1    g06666(.A1(new_n6720_), .A2(new_n6722_), .A3(new_n6713_), .ZN(new_n6731_));
  OAI21_X1   g06667(.A1(new_n6731_), .A2(new_n6717_), .B(new_n6648_), .ZN(new_n6732_));
  NOR3_X1    g06668(.A1(new_n6708_), .A2(new_n6722_), .A3(new_n6713_), .ZN(new_n6733_));
  AOI21_X1   g06669(.A1(new_n6712_), .A2(new_n6714_), .B(new_n6720_), .ZN(new_n6734_));
  OAI21_X1   g06670(.A1(new_n6734_), .A2(new_n6733_), .B(new_n6649_), .ZN(new_n6735_));
  NAND2_X1   g06671(.A1(new_n6735_), .A2(new_n6732_), .ZN(new_n6736_));
  XOR2_X1    g06672(.A1(new_n6728_), .A2(\a[17] ), .Z(new_n6737_));
  NOR2_X1    g06673(.A1(new_n6737_), .A2(new_n6736_), .ZN(new_n6738_));
  NOR2_X1    g06674(.A1(new_n6730_), .A2(new_n6738_), .ZN(new_n6739_));
  OAI22_X1   g06675(.A1(new_n896_), .A2(new_n6091_), .B1(new_n1180_), .B2(new_n6089_), .ZN(new_n6740_));
  NAND2_X1   g06676(.A1(new_n2504_), .A2(new_n6095_), .ZN(new_n6741_));
  AOI21_X1   g06677(.A1(new_n6741_), .A2(new_n6740_), .B(new_n6082_), .ZN(new_n6742_));
  NAND3_X1   g06678(.A1(new_n3596_), .A2(new_n3521_), .A3(new_n6742_), .ZN(new_n6743_));
  AOI21_X1   g06679(.A1(new_n3596_), .A2(new_n6742_), .B(new_n3521_), .ZN(new_n6744_));
  INV_X1     g06680(.I(new_n6744_), .ZN(new_n6745_));
  NAND3_X1   g06681(.A1(new_n6739_), .A2(new_n6745_), .A3(new_n6743_), .ZN(new_n6746_));
  NAND2_X1   g06682(.A1(new_n6737_), .A2(new_n6736_), .ZN(new_n6747_));
  NAND2_X1   g06683(.A1(new_n6725_), .A2(new_n6729_), .ZN(new_n6748_));
  NAND2_X1   g06684(.A1(new_n6748_), .A2(new_n6747_), .ZN(new_n6749_));
  INV_X1     g06685(.I(new_n6743_), .ZN(new_n6750_));
  OAI21_X1   g06686(.A1(new_n6750_), .A2(new_n6744_), .B(new_n6749_), .ZN(new_n6751_));
  AOI21_X1   g06687(.A1(new_n6751_), .A2(new_n6746_), .B(new_n6643_), .ZN(new_n6752_));
  INV_X1     g06688(.I(new_n6643_), .ZN(new_n6753_));
  NAND3_X1   g06689(.A1(new_n6749_), .A2(new_n6745_), .A3(new_n6743_), .ZN(new_n6754_));
  OAI21_X1   g06690(.A1(new_n6750_), .A2(new_n6744_), .B(new_n6739_), .ZN(new_n6755_));
  AOI21_X1   g06691(.A1(new_n6755_), .A2(new_n6754_), .B(new_n6753_), .ZN(new_n6756_));
  OAI21_X1   g06692(.A1(new_n6756_), .A2(new_n6752_), .B(new_n4034_), .ZN(new_n6757_));
  NOR3_X1    g06693(.A1(new_n6749_), .A2(new_n6744_), .A3(new_n6750_), .ZN(new_n6758_));
  AOI21_X1   g06694(.A1(new_n6743_), .A2(new_n6745_), .B(new_n6739_), .ZN(new_n6759_));
  OAI21_X1   g06695(.A1(new_n6759_), .A2(new_n6758_), .B(new_n6753_), .ZN(new_n6760_));
  NOR3_X1    g06696(.A1(new_n6739_), .A2(new_n6744_), .A3(new_n6750_), .ZN(new_n6761_));
  AOI21_X1   g06697(.A1(new_n6743_), .A2(new_n6745_), .B(new_n6749_), .ZN(new_n6762_));
  OAI21_X1   g06698(.A1(new_n6762_), .A2(new_n6761_), .B(new_n6643_), .ZN(new_n6763_));
  NAND3_X1   g06699(.A1(new_n6760_), .A2(new_n6763_), .A3(\a[11] ), .ZN(new_n6764_));
  AOI21_X1   g06700(.A1(new_n6757_), .A2(new_n6764_), .B(new_n6638_), .ZN(new_n6765_));
  AOI21_X1   g06701(.A1(new_n6760_), .A2(new_n6763_), .B(\a[11] ), .ZN(new_n6766_));
  NOR3_X1    g06702(.A1(new_n6756_), .A2(new_n6752_), .A3(new_n4034_), .ZN(new_n6767_));
  NOR3_X1    g06703(.A1(new_n6766_), .A2(new_n6767_), .A3(new_n6637_), .ZN(new_n6768_));
  NOR2_X1    g06704(.A1(new_n6768_), .A2(new_n6765_), .ZN(new_n6769_));
  INV_X1     g06705(.I(\a[6] ), .ZN(new_n6770_));
  NOR2_X1    g06706(.A1(new_n6770_), .A2(\a[5] ), .ZN(new_n6771_));
  NOR2_X1    g06707(.A1(new_n65_), .A2(\a[6] ), .ZN(new_n6772_));
  NOR2_X1    g06708(.A1(new_n6771_), .A2(new_n6772_), .ZN(new_n6773_));
  XNOR2_X1   g06709(.A1(\a[7] ), .A2(\a[8] ), .ZN(new_n6774_));
  NOR2_X1    g06710(.A1(new_n6773_), .A2(new_n6774_), .ZN(new_n6775_));
  INV_X1     g06711(.I(new_n6775_), .ZN(new_n6776_));
  INV_X1     g06712(.I(new_n6773_), .ZN(new_n6777_));
  INV_X1     g06713(.I(\a[7] ), .ZN(new_n6778_));
  NOR2_X1    g06714(.A1(new_n6778_), .A2(\a[5] ), .ZN(new_n6779_));
  NOR2_X1    g06715(.A1(new_n65_), .A2(\a[7] ), .ZN(new_n6780_));
  OR2_X2     g06716(.A1(new_n6779_), .A2(new_n6780_), .Z(new_n6781_));
  XNOR2_X1   g06717(.A1(\a[5] ), .A2(\a[8] ), .ZN(new_n6782_));
  OAI21_X1   g06718(.A1(new_n6777_), .A2(new_n6781_), .B(new_n6782_), .ZN(new_n6783_));
  NOR2_X1    g06719(.A1(new_n6777_), .A2(new_n6774_), .ZN(new_n6784_));
  INV_X1     g06720(.I(new_n6784_), .ZN(new_n6785_));
  OAI22_X1   g06721(.A1(new_n694_), .A2(new_n6783_), .B1(new_n2665_), .B2(new_n6785_), .ZN(new_n6786_));
  NOR3_X1    g06722(.A1(new_n6778_), .A2(\a[5] ), .A3(\a[6] ), .ZN(new_n6787_));
  AOI21_X1   g06723(.A1(\a[6] ), .A2(new_n6780_), .B(new_n6787_), .ZN(new_n6788_));
  INV_X1     g06724(.I(new_n6788_), .ZN(new_n6789_));
  NAND2_X1   g06725(.A1(new_n2615_), .A2(new_n6789_), .ZN(new_n6790_));
  AOI21_X1   g06726(.A1(new_n6786_), .A2(new_n6790_), .B(new_n6776_), .ZN(new_n6791_));
  NAND3_X1   g06727(.A1(new_n3188_), .A2(new_n4009_), .A3(new_n6791_), .ZN(new_n6792_));
  AOI21_X1   g06728(.A1(new_n3188_), .A2(new_n6791_), .B(new_n4009_), .ZN(new_n6793_));
  INV_X1     g06729(.I(new_n6793_), .ZN(new_n6794_));
  NAND3_X1   g06730(.A1(new_n6794_), .A2(new_n6769_), .A3(new_n6792_), .ZN(new_n6795_));
  OAI21_X1   g06731(.A1(new_n6766_), .A2(new_n6767_), .B(new_n6637_), .ZN(new_n6796_));
  NAND3_X1   g06732(.A1(new_n6757_), .A2(new_n6764_), .A3(new_n6638_), .ZN(new_n6797_));
  NAND2_X1   g06733(.A1(new_n6796_), .A2(new_n6797_), .ZN(new_n6798_));
  INV_X1     g06734(.I(new_n6792_), .ZN(new_n6799_));
  OAI21_X1   g06735(.A1(new_n6799_), .A2(new_n6793_), .B(new_n6798_), .ZN(new_n6800_));
  AOI21_X1   g06736(.A1(new_n6800_), .A2(new_n6795_), .B(new_n6633_), .ZN(new_n6801_));
  NAND2_X1   g06737(.A1(new_n6499_), .A2(new_n6146_), .ZN(new_n6802_));
  NOR3_X1    g06738(.A1(new_n6157_), .A2(new_n6216_), .A3(new_n6215_), .ZN(new_n6803_));
  AOI21_X1   g06739(.A1(new_n6207_), .A2(new_n6213_), .B(new_n6158_), .ZN(new_n6804_));
  NOR2_X1    g06740(.A1(new_n6804_), .A2(new_n6803_), .ZN(new_n6805_));
  OAI21_X1   g06741(.A1(new_n6215_), .A2(new_n6216_), .B(new_n6157_), .ZN(new_n6806_));
  INV_X1     g06742(.I(new_n6241_), .ZN(new_n6807_));
  NAND3_X1   g06743(.A1(new_n6468_), .A2(new_n6469_), .A3(new_n6467_), .ZN(new_n6808_));
  OAI21_X1   g06744(.A1(new_n6465_), .A2(new_n6427_), .B(new_n6246_), .ZN(new_n6809_));
  NAND2_X1   g06745(.A1(new_n6478_), .A2(new_n6475_), .ZN(new_n6810_));
  INV_X1     g06746(.I(new_n6485_), .ZN(new_n6811_));
  XOR2_X1    g06747(.A1(new_n6486_), .A2(new_n6456_), .Z(new_n6812_));
  NAND2_X1   g06748(.A1(new_n6812_), .A2(new_n6811_), .ZN(new_n6813_));
  NAND2_X1   g06749(.A1(new_n6810_), .A2(new_n6813_), .ZN(new_n6814_));
  AOI22_X1   g06750(.A1(new_n6809_), .A2(new_n6808_), .B1(new_n6467_), .B2(new_n6814_), .ZN(new_n6815_));
  OAI21_X1   g06751(.A1(new_n6815_), .A2(new_n6493_), .B(new_n6807_), .ZN(new_n6816_));
  NAND3_X1   g06752(.A1(new_n6816_), .A2(new_n6230_), .A3(new_n6234_), .ZN(new_n6817_));
  OAI21_X1   g06753(.A1(new_n6817_), .A2(new_n6805_), .B(new_n6806_), .ZN(new_n6818_));
  NAND2_X1   g06754(.A1(new_n6147_), .A2(new_n6149_), .ZN(new_n6819_));
  NAND2_X1   g06755(.A1(new_n6819_), .A2(new_n6802_), .ZN(new_n6820_));
  OAI21_X1   g06756(.A1(new_n6818_), .A2(new_n6820_), .B(new_n6802_), .ZN(new_n6821_));
  NAND3_X1   g06757(.A1(new_n6821_), .A2(new_n6135_), .A3(new_n6139_), .ZN(new_n6822_));
  NAND3_X1   g06758(.A1(new_n6629_), .A2(new_n6630_), .A3(new_n6631_), .ZN(new_n6823_));
  OAI21_X1   g06759(.A1(new_n6624_), .A2(new_n6627_), .B(new_n4724_), .ZN(new_n6824_));
  AOI22_X1   g06760(.A1(new_n6823_), .A2(new_n6824_), .B1(new_n6631_), .B2(new_n6822_), .ZN(new_n6825_));
  NAND3_X1   g06761(.A1(new_n6794_), .A2(new_n6798_), .A3(new_n6792_), .ZN(new_n6826_));
  OAI21_X1   g06762(.A1(new_n6799_), .A2(new_n6793_), .B(new_n6769_), .ZN(new_n6827_));
  AOI21_X1   g06763(.A1(new_n6827_), .A2(new_n6826_), .B(new_n6825_), .ZN(new_n6828_));
  NOR2_X1    g06764(.A1(new_n6828_), .A2(new_n6801_), .ZN(new_n6829_));
  INV_X1     g06765(.I(\a[3] ), .ZN(new_n6830_));
  NOR2_X1    g06766(.A1(new_n6830_), .A2(\a[2] ), .ZN(new_n6831_));
  NOR2_X1    g06767(.A1(new_n4387_), .A2(\a[3] ), .ZN(new_n6832_));
  NOR2_X1    g06768(.A1(new_n6831_), .A2(new_n6832_), .ZN(new_n6833_));
  XNOR2_X1   g06769(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n6834_));
  NOR2_X1    g06770(.A1(new_n6833_), .A2(new_n6834_), .ZN(new_n6835_));
  INV_X1     g06771(.I(new_n6835_), .ZN(new_n6836_));
  INV_X1     g06772(.I(new_n6833_), .ZN(new_n6837_));
  NOR2_X1    g06773(.A1(new_n6837_), .A2(new_n6834_), .ZN(new_n6838_));
  INV_X1     g06774(.I(new_n6838_), .ZN(new_n6839_));
  NOR3_X1    g06775(.A1(new_n4387_), .A2(new_n6830_), .A3(\a[4] ), .ZN(new_n6840_));
  NAND3_X1   g06776(.A1(new_n4387_), .A2(new_n6830_), .A3(\a[4] ), .ZN(new_n6841_));
  INV_X1     g06777(.I(new_n6841_), .ZN(new_n6842_));
  NOR2_X1    g06778(.A1(new_n6842_), .A2(new_n6840_), .ZN(new_n6843_));
  OAI22_X1   g06779(.A1(new_n3176_), .A2(new_n6843_), .B1(new_n3142_), .B2(new_n6839_), .ZN(new_n6844_));
  XNOR2_X1   g06780(.A1(\a[2] ), .A2(\a[4] ), .ZN(new_n6845_));
  AOI21_X1   g06781(.A1(new_n6833_), .A2(new_n6845_), .B(new_n4610_), .ZN(new_n6846_));
  NAND2_X1   g06782(.A1(new_n2728_), .A2(new_n6846_), .ZN(new_n6847_));
  AOI21_X1   g06783(.A1(new_n6844_), .A2(new_n6847_), .B(new_n6836_), .ZN(new_n6848_));
  OAI21_X1   g06784(.A1(new_n3173_), .A2(new_n3172_), .B(new_n6848_), .ZN(new_n6849_));
  NOR2_X1    g06785(.A1(new_n6849_), .A2(\a[5] ), .ZN(new_n6850_));
  NAND2_X1   g06786(.A1(new_n6849_), .A2(\a[5] ), .ZN(new_n6851_));
  INV_X1     g06787(.I(new_n6851_), .ZN(new_n6852_));
  OAI21_X1   g06788(.A1(new_n6850_), .A2(new_n6852_), .B(new_n6829_), .ZN(new_n6853_));
  NAND2_X1   g06789(.A1(new_n6629_), .A2(new_n6630_), .ZN(new_n6854_));
  NAND2_X1   g06790(.A1(new_n6822_), .A2(new_n4724_), .ZN(new_n6855_));
  NAND4_X1   g06791(.A1(new_n6821_), .A2(new_n6631_), .A3(new_n6135_), .A4(new_n6139_), .ZN(new_n6856_));
  AOI21_X1   g06792(.A1(new_n6855_), .A2(new_n6856_), .B(new_n6854_), .ZN(new_n6857_));
  NOR2_X1    g06793(.A1(new_n6624_), .A2(new_n6627_), .ZN(new_n6858_));
  NOR2_X1    g06794(.A1(new_n6503_), .A2(new_n6631_), .ZN(new_n6859_));
  NOR4_X1    g06795(.A1(new_n6502_), .A2(new_n6140_), .A3(new_n4724_), .A4(new_n6131_), .ZN(new_n6860_));
  NOR3_X1    g06796(.A1(new_n6859_), .A2(new_n6858_), .A3(new_n6860_), .ZN(new_n6861_));
  NOR2_X1    g06797(.A1(new_n6861_), .A2(new_n6857_), .ZN(new_n6862_));
  OAI22_X1   g06798(.A1(new_n2614_), .A2(new_n6785_), .B1(new_n529_), .B2(new_n6783_), .ZN(new_n6863_));
  NAND2_X1   g06799(.A1(new_n2718_), .A2(new_n6789_), .ZN(new_n6864_));
  AOI21_X1   g06800(.A1(new_n6864_), .A2(new_n6863_), .B(new_n6776_), .ZN(new_n6865_));
  NAND3_X1   g06801(.A1(new_n3074_), .A2(new_n4009_), .A3(new_n6865_), .ZN(new_n6866_));
  AOI21_X1   g06802(.A1(new_n3074_), .A2(new_n6865_), .B(new_n4009_), .ZN(new_n6867_));
  INV_X1     g06803(.I(new_n6867_), .ZN(new_n6868_));
  NAND2_X1   g06804(.A1(new_n6868_), .A2(new_n6866_), .ZN(new_n6869_));
  AOI22_X1   g06805(.A1(new_n6133_), .A2(new_n6132_), .B1(new_n6136_), .B2(new_n6137_), .ZN(new_n6870_));
  NOR2_X1    g06806(.A1(new_n6870_), .A2(new_n6131_), .ZN(new_n6871_));
  NAND2_X1   g06807(.A1(new_n6502_), .A2(new_n6871_), .ZN(new_n6872_));
  NAND2_X1   g06808(.A1(new_n6821_), .A2(new_n6140_), .ZN(new_n6873_));
  OAI22_X1   g06809(.A1(new_n2559_), .A2(new_n6783_), .B1(new_n694_), .B2(new_n6785_), .ZN(new_n6874_));
  NAND2_X1   g06810(.A1(new_n2567_), .A2(new_n6789_), .ZN(new_n6875_));
  AOI21_X1   g06811(.A1(new_n6874_), .A2(new_n6875_), .B(new_n6776_), .ZN(new_n6876_));
  NAND3_X1   g06812(.A1(new_n2759_), .A2(new_n4009_), .A3(new_n6876_), .ZN(new_n6877_));
  AOI21_X1   g06813(.A1(new_n2759_), .A2(new_n6876_), .B(new_n4009_), .ZN(new_n6878_));
  INV_X1     g06814(.I(new_n6878_), .ZN(new_n6879_));
  NAND2_X1   g06815(.A1(new_n6879_), .A2(new_n6877_), .ZN(new_n6880_));
  AOI21_X1   g06816(.A1(new_n6872_), .A2(new_n6873_), .B(new_n6880_), .ZN(new_n6881_));
  NOR2_X1    g06817(.A1(new_n6821_), .A2(new_n6140_), .ZN(new_n6882_));
  NOR2_X1    g06818(.A1(new_n6502_), .A2(new_n6871_), .ZN(new_n6883_));
  INV_X1     g06819(.I(new_n6877_), .ZN(new_n6884_));
  NOR2_X1    g06820(.A1(new_n6884_), .A2(new_n6878_), .ZN(new_n6885_));
  NOR3_X1    g06821(.A1(new_n6883_), .A2(new_n6882_), .A3(new_n6885_), .ZN(new_n6886_));
  OAI22_X1   g06822(.A1(new_n813_), .A2(new_n6783_), .B1(new_n529_), .B2(new_n6785_), .ZN(new_n6887_));
  NAND2_X1   g06823(.A1(new_n2563_), .A2(new_n6789_), .ZN(new_n6888_));
  AOI21_X1   g06824(.A1(new_n6888_), .A2(new_n6887_), .B(new_n6776_), .ZN(new_n6889_));
  NAND2_X1   g06825(.A1(new_n3051_), .A2(new_n6889_), .ZN(new_n6890_));
  XOR2_X1    g06826(.A1(new_n6890_), .A2(\a[8] ), .Z(new_n6891_));
  NOR2_X1    g06827(.A1(new_n6818_), .A2(new_n6501_), .ZN(new_n6892_));
  NOR2_X1    g06828(.A1(new_n6497_), .A2(new_n6820_), .ZN(new_n6893_));
  OAI21_X1   g06829(.A1(new_n6893_), .A2(new_n6892_), .B(new_n6891_), .ZN(new_n6894_));
  INV_X1     g06830(.I(new_n6894_), .ZN(new_n6895_));
  NOR3_X1    g06831(.A1(new_n6881_), .A2(new_n6886_), .A3(new_n6895_), .ZN(new_n6896_));
  NOR2_X1    g06832(.A1(new_n6896_), .A2(new_n6869_), .ZN(new_n6897_));
  INV_X1     g06833(.I(new_n6866_), .ZN(new_n6898_));
  NOR2_X1    g06834(.A1(new_n6898_), .A2(new_n6867_), .ZN(new_n6899_));
  NOR4_X1    g06835(.A1(new_n6899_), .A2(new_n6881_), .A3(new_n6886_), .A4(new_n6895_), .ZN(new_n6900_));
  OAI21_X1   g06836(.A1(new_n6897_), .A2(new_n6900_), .B(new_n6862_), .ZN(new_n6901_));
  OAI21_X1   g06837(.A1(new_n6859_), .A2(new_n6860_), .B(new_n6858_), .ZN(new_n6902_));
  NAND3_X1   g06838(.A1(new_n6855_), .A2(new_n6854_), .A3(new_n6856_), .ZN(new_n6903_));
  NAND2_X1   g06839(.A1(new_n6902_), .A2(new_n6903_), .ZN(new_n6904_));
  OAI21_X1   g06840(.A1(new_n6883_), .A2(new_n6882_), .B(new_n6885_), .ZN(new_n6905_));
  NAND3_X1   g06841(.A1(new_n6872_), .A2(new_n6873_), .A3(new_n6880_), .ZN(new_n6906_));
  NAND3_X1   g06842(.A1(new_n6905_), .A2(new_n6906_), .A3(new_n6894_), .ZN(new_n6907_));
  NAND2_X1   g06843(.A1(new_n6907_), .A2(new_n6899_), .ZN(new_n6908_));
  NAND4_X1   g06844(.A1(new_n6869_), .A2(new_n6905_), .A3(new_n6906_), .A4(new_n6894_), .ZN(new_n6909_));
  NAND3_X1   g06845(.A1(new_n6908_), .A2(new_n6904_), .A3(new_n6909_), .ZN(new_n6910_));
  NOR2_X1    g06846(.A1(new_n3176_), .A2(new_n6839_), .ZN(new_n6911_));
  NOR2_X1    g06847(.A1(new_n2716_), .A2(new_n6843_), .ZN(new_n6912_));
  INV_X1     g06848(.I(new_n6846_), .ZN(new_n6913_));
  NOR2_X1    g06849(.A1(new_n2665_), .A2(new_n6913_), .ZN(new_n6914_));
  NOR4_X1    g06850(.A1(new_n6911_), .A2(new_n6912_), .A3(new_n6914_), .A4(new_n6836_), .ZN(new_n6915_));
  NAND2_X1   g06851(.A1(new_n3273_), .A2(new_n6915_), .ZN(new_n6916_));
  XOR2_X1    g06852(.A1(new_n6916_), .A2(\a[5] ), .Z(new_n6917_));
  AOI21_X1   g06853(.A1(new_n6901_), .A2(new_n6910_), .B(new_n6917_), .ZN(new_n6918_));
  NAND3_X1   g06854(.A1(new_n6901_), .A2(new_n6910_), .A3(new_n6917_), .ZN(new_n6919_));
  INV_X1     g06855(.I(\a[0] ), .ZN(new_n6920_));
  XNOR2_X1   g06856(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n6921_));
  NOR2_X1    g06857(.A1(new_n6921_), .A2(new_n6920_), .ZN(new_n6922_));
  NOR2_X1    g06858(.A1(\a[0] ), .A2(\a[1] ), .ZN(new_n6923_));
  INV_X1     g06859(.I(new_n6923_), .ZN(new_n6924_));
  NOR2_X1    g06860(.A1(new_n6924_), .A2(new_n4387_), .ZN(new_n6925_));
  AOI22_X1   g06861(.A1(new_n3253_), .A2(new_n6922_), .B1(new_n3247_), .B2(new_n6925_), .ZN(new_n6926_));
  XOR2_X1    g06862(.A1(new_n6926_), .A2(new_n4387_), .Z(new_n6927_));
  AOI21_X1   g06863(.A1(new_n6919_), .A2(new_n6927_), .B(new_n6918_), .ZN(new_n6928_));
  NOR3_X1    g06864(.A1(new_n6799_), .A2(new_n6798_), .A3(new_n6793_), .ZN(new_n6929_));
  AOI21_X1   g06865(.A1(new_n6794_), .A2(new_n6792_), .B(new_n6769_), .ZN(new_n6930_));
  OAI21_X1   g06866(.A1(new_n6930_), .A2(new_n6929_), .B(new_n6825_), .ZN(new_n6931_));
  NOR3_X1    g06867(.A1(new_n6769_), .A2(new_n6799_), .A3(new_n6793_), .ZN(new_n6932_));
  AOI21_X1   g06868(.A1(new_n6794_), .A2(new_n6792_), .B(new_n6798_), .ZN(new_n6933_));
  OAI21_X1   g06869(.A1(new_n6933_), .A2(new_n6932_), .B(new_n6633_), .ZN(new_n6934_));
  NAND2_X1   g06870(.A1(new_n6931_), .A2(new_n6934_), .ZN(new_n6935_));
  INV_X1     g06871(.I(new_n6850_), .ZN(new_n6936_));
  NAND3_X1   g06872(.A1(new_n6935_), .A2(new_n6936_), .A3(new_n6851_), .ZN(new_n6937_));
  NAND2_X1   g06873(.A1(new_n6853_), .A2(new_n6937_), .ZN(new_n6938_));
  NAND2_X1   g06874(.A1(new_n6928_), .A2(new_n6938_), .ZN(new_n6939_));
  AOI21_X1   g06875(.A1(new_n6908_), .A2(new_n6909_), .B(new_n6904_), .ZN(new_n6940_));
  NOR3_X1    g06876(.A1(new_n6897_), .A2(new_n6862_), .A3(new_n6900_), .ZN(new_n6941_));
  XOR2_X1    g06877(.A1(new_n6916_), .A2(new_n65_), .Z(new_n6942_));
  OAI21_X1   g06878(.A1(new_n6940_), .A2(new_n6941_), .B(new_n6942_), .ZN(new_n6943_));
  NOR3_X1    g06879(.A1(new_n6940_), .A2(new_n6941_), .A3(new_n6942_), .ZN(new_n6944_));
  XOR2_X1    g06880(.A1(new_n6926_), .A2(\a[2] ), .Z(new_n6945_));
  OAI21_X1   g06881(.A1(new_n6944_), .A2(new_n6945_), .B(new_n6943_), .ZN(new_n6946_));
  NOR3_X1    g06882(.A1(new_n6829_), .A2(new_n6852_), .A3(new_n6850_), .ZN(new_n6947_));
  AOI21_X1   g06883(.A1(new_n6936_), .A2(new_n6851_), .B(new_n6935_), .ZN(new_n6948_));
  NOR2_X1    g06884(.A1(new_n6948_), .A2(new_n6947_), .ZN(new_n6949_));
  AOI21_X1   g06885(.A1(new_n6825_), .A2(new_n6826_), .B(new_n6933_), .ZN(new_n6950_));
  INV_X1     g06886(.I(new_n6950_), .ZN(new_n6951_));
  OAI21_X1   g06887(.A1(new_n3142_), .A2(new_n6843_), .B(new_n6835_), .ZN(new_n6952_));
  AOI21_X1   g06888(.A1(new_n3168_), .A2(new_n6846_), .B(new_n6952_), .ZN(new_n6953_));
  NAND4_X1   g06889(.A1(new_n3757_), .A2(new_n65_), .A3(new_n3755_), .A4(new_n6953_), .ZN(new_n6954_));
  NAND3_X1   g06890(.A1(new_n3757_), .A2(new_n3755_), .A3(new_n6953_), .ZN(new_n6955_));
  NAND2_X1   g06891(.A1(new_n6955_), .A2(\a[5] ), .ZN(new_n6956_));
  NAND2_X1   g06892(.A1(new_n6956_), .A2(new_n6954_), .ZN(new_n6957_));
  INV_X1     g06893(.I(new_n6957_), .ZN(new_n6958_));
  AOI21_X1   g06894(.A1(new_n2725_), .A2(new_n2726_), .B(new_n2717_), .ZN(new_n6959_));
  INV_X1     g06895(.I(new_n2732_), .ZN(new_n6960_));
  OAI22_X1   g06896(.A1(new_n2614_), .A2(new_n6783_), .B1(new_n2665_), .B2(new_n6788_), .ZN(new_n6961_));
  NAND2_X1   g06897(.A1(new_n2728_), .A2(new_n6784_), .ZN(new_n6962_));
  AOI21_X1   g06898(.A1(new_n6962_), .A2(new_n6961_), .B(new_n6776_), .ZN(new_n6963_));
  OAI21_X1   g06899(.A1(new_n6960_), .A2(new_n6959_), .B(new_n6963_), .ZN(new_n6964_));
  NOR2_X1    g06900(.A1(new_n6964_), .A2(\a[8] ), .ZN(new_n6965_));
  AOI21_X1   g06901(.A1(new_n2733_), .A2(new_n6963_), .B(new_n4009_), .ZN(new_n6966_));
  NOR2_X1    g06902(.A1(new_n6965_), .A2(new_n6966_), .ZN(new_n6967_));
  NOR2_X1    g06903(.A1(new_n2722_), .A2(new_n2755_), .ZN(new_n6968_));
  OAI22_X1   g06904(.A1(new_n2559_), .A2(new_n4716_), .B1(new_n694_), .B2(new_n4710_), .ZN(new_n6969_));
  NAND2_X1   g06905(.A1(new_n2567_), .A2(new_n4720_), .ZN(new_n6970_));
  AOI21_X1   g06906(.A1(new_n6969_), .A2(new_n6970_), .B(new_n4707_), .ZN(new_n6971_));
  OAI21_X1   g06907(.A1(new_n6968_), .A2(new_n2757_), .B(new_n6971_), .ZN(new_n6972_));
  XOR2_X1    g06908(.A1(new_n6972_), .A2(new_n4034_), .Z(new_n6973_));
  OAI21_X1   g06909(.A1(new_n6643_), .A2(new_n6761_), .B(new_n6755_), .ZN(new_n6974_));
  OAI22_X1   g06910(.A1(new_n1180_), .A2(new_n4470_), .B1(new_n2492_), .B2(new_n4291_), .ZN(new_n6975_));
  NAND2_X1   g06911(.A1(new_n1122_), .A2(new_n4298_), .ZN(new_n6976_));
  AOI21_X1   g06912(.A1(new_n6976_), .A2(new_n6975_), .B(new_n4468_), .ZN(new_n6977_));
  NAND2_X1   g06913(.A1(new_n3330_), .A2(new_n6977_), .ZN(new_n6978_));
  XOR2_X1    g06914(.A1(new_n6978_), .A2(\a[17] ), .Z(new_n6979_));
  OAI22_X1   g06915(.A1(new_n2367_), .A2(new_n3769_), .B1(new_n2451_), .B2(new_n4097_), .ZN(new_n6980_));
  NAND2_X1   g06916(.A1(new_n2412_), .A2(new_n3776_), .ZN(new_n6981_));
  AOI21_X1   g06917(.A1(new_n6980_), .A2(new_n6981_), .B(new_n4095_), .ZN(new_n6982_));
  NAND3_X1   g06918(.A1(new_n3403_), .A2(new_n3035_), .A3(new_n6982_), .ZN(new_n6983_));
  INV_X1     g06919(.I(new_n6983_), .ZN(new_n6984_));
  AOI21_X1   g06920(.A1(new_n3403_), .A2(new_n6982_), .B(new_n3035_), .ZN(new_n6985_));
  NOR2_X1    g06921(.A1(new_n6984_), .A2(new_n6985_), .ZN(new_n6986_));
  INV_X1     g06922(.I(new_n6689_), .ZN(new_n6987_));
  AOI21_X1   g06923(.A1(new_n6652_), .A2(new_n6688_), .B(new_n6987_), .ZN(new_n6988_));
  OAI22_X1   g06924(.A1(new_n2251_), .A2(new_n3268_), .B1(new_n2351_), .B2(new_n3318_), .ZN(new_n6989_));
  NAND2_X1   g06925(.A1(new_n2310_), .A2(new_n3323_), .ZN(new_n6990_));
  AOI21_X1   g06926(.A1(new_n6990_), .A2(new_n6989_), .B(new_n3260_), .ZN(new_n6991_));
  NAND3_X1   g06927(.A1(new_n3914_), .A2(new_n72_), .A3(new_n6991_), .ZN(new_n6992_));
  OAI21_X1   g06928(.A1(new_n5555_), .A2(new_n3911_), .B(new_n6991_), .ZN(new_n6993_));
  NAND2_X1   g06929(.A1(new_n6993_), .A2(\a[26] ), .ZN(new_n6994_));
  NAND2_X1   g06930(.A1(new_n6992_), .A2(new_n6994_), .ZN(new_n6995_));
  INV_X1     g06931(.I(new_n6672_), .ZN(new_n6996_));
  INV_X1     g06932(.I(new_n6657_), .ZN(new_n6997_));
  INV_X1     g06933(.I(new_n6671_), .ZN(new_n6998_));
  OAI21_X1   g06934(.A1(new_n6997_), .A2(new_n6658_), .B(new_n6998_), .ZN(new_n6999_));
  NAND2_X1   g06935(.A1(new_n4589_), .A2(new_n4585_), .ZN(new_n7000_));
  NAND2_X1   g06936(.A1(new_n4571_), .A2(new_n7000_), .ZN(new_n7001_));
  XOR2_X1    g06937(.A1(new_n4587_), .A2(new_n4387_), .Z(new_n7002_));
  OAI21_X1   g06938(.A1(new_n4571_), .A2(new_n7002_), .B(new_n7001_), .ZN(new_n7003_));
  AOI21_X1   g06939(.A1(new_n2760_), .A2(new_n2761_), .B(new_n2769_), .ZN(new_n7004_));
  OAI21_X1   g06940(.A1(new_n2103_), .A2(new_n2767_), .B(new_n7004_), .ZN(new_n7005_));
  AOI21_X1   g06941(.A1(new_n2107_), .A2(new_n2770_), .B(new_n7005_), .ZN(new_n7006_));
  NAND2_X1   g06942(.A1(new_n4959_), .A2(new_n7006_), .ZN(new_n7007_));
  INV_X1     g06943(.I(new_n7007_), .ZN(new_n7008_));
  NOR2_X1    g06944(.A1(new_n7003_), .A2(new_n7008_), .ZN(new_n7009_));
  INV_X1     g06945(.I(new_n7009_), .ZN(new_n7010_));
  NAND2_X1   g06946(.A1(new_n7003_), .A2(new_n7008_), .ZN(new_n7011_));
  AOI22_X1   g06947(.A1(new_n6999_), .A2(new_n6996_), .B1(new_n7010_), .B2(new_n7011_), .ZN(new_n7012_));
  AOI21_X1   g06948(.A1(new_n6659_), .A2(new_n6657_), .B(new_n6671_), .ZN(new_n7013_));
  XOR2_X1    g06949(.A1(new_n7003_), .A2(new_n7007_), .Z(new_n7014_));
  NOR3_X1    g06950(.A1(new_n7014_), .A2(new_n6672_), .A3(new_n7013_), .ZN(new_n7015_));
  NOR2_X1    g06951(.A1(new_n7015_), .A2(new_n7012_), .ZN(new_n7016_));
  OAI22_X1   g06952(.A1(new_n4365_), .A2(new_n3175_), .B1(new_n2198_), .B2(new_n2747_), .ZN(new_n7017_));
  NAND2_X1   g06953(.A1(new_n1504_), .A2(new_n3275_), .ZN(new_n7018_));
  AOI21_X1   g06954(.A1(new_n7017_), .A2(new_n7018_), .B(new_n2737_), .ZN(new_n7019_));
  NAND2_X1   g06955(.A1(new_n4363_), .A2(new_n7019_), .ZN(new_n7020_));
  XOR2_X1    g06956(.A1(new_n7020_), .A2(\a[29] ), .Z(new_n7021_));
  NAND2_X1   g06957(.A1(new_n7016_), .A2(new_n7021_), .ZN(new_n7022_));
  XOR2_X1    g06958(.A1(new_n7020_), .A2(new_n74_), .Z(new_n7023_));
  OAI21_X1   g06959(.A1(new_n7012_), .A2(new_n7015_), .B(new_n7023_), .ZN(new_n7024_));
  NAND2_X1   g06960(.A1(new_n7022_), .A2(new_n7024_), .ZN(new_n7025_));
  OAI21_X1   g06961(.A1(new_n7012_), .A2(new_n7015_), .B(new_n7021_), .ZN(new_n7026_));
  INV_X1     g06962(.I(new_n7011_), .ZN(new_n7027_));
  OAI22_X1   g06963(.A1(new_n7013_), .A2(new_n6672_), .B1(new_n7027_), .B2(new_n7009_), .ZN(new_n7028_));
  XOR2_X1    g06964(.A1(new_n7003_), .A2(new_n7008_), .Z(new_n7029_));
  NAND3_X1   g06965(.A1(new_n7029_), .A2(new_n6999_), .A3(new_n6996_), .ZN(new_n7030_));
  NAND3_X1   g06966(.A1(new_n7030_), .A2(new_n7023_), .A3(new_n7028_), .ZN(new_n7031_));
  NAND2_X1   g06967(.A1(new_n7026_), .A2(new_n7031_), .ZN(new_n7032_));
  MUX2_X1    g06968(.I0(new_n7032_), .I1(new_n7025_), .S(new_n6995_), .Z(new_n7033_));
  AOI21_X1   g06969(.A1(new_n3824_), .A2(new_n3827_), .B(new_n3302_), .ZN(new_n7034_));
  NOR2_X1    g06970(.A1(new_n1333_), .A2(new_n3780_), .ZN(new_n7035_));
  NOR2_X1    g06971(.A1(new_n1409_), .A2(new_n3306_), .ZN(new_n7036_));
  OAI22_X1   g06972(.A1(new_n7036_), .A2(new_n7035_), .B1(new_n1453_), .B2(new_n3310_), .ZN(new_n7037_));
  OAI21_X1   g06973(.A1(new_n7034_), .A2(new_n7037_), .B(new_n7033_), .ZN(new_n7038_));
  INV_X1     g06974(.I(new_n6995_), .ZN(new_n7039_));
  AOI22_X1   g06975(.A1(new_n7022_), .A2(new_n7024_), .B1(new_n6994_), .B2(new_n6992_), .ZN(new_n7040_));
  AOI21_X1   g06976(.A1(new_n7039_), .A2(new_n7032_), .B(new_n7040_), .ZN(new_n7041_));
  OAI21_X1   g06977(.A1(new_n5536_), .A2(new_n3823_), .B(new_n3301_), .ZN(new_n7042_));
  INV_X1     g06978(.I(new_n7037_), .ZN(new_n7043_));
  NAND3_X1   g06979(.A1(new_n7041_), .A2(new_n7042_), .A3(new_n7043_), .ZN(new_n7044_));
  AOI21_X1   g06980(.A1(new_n7038_), .A2(new_n7044_), .B(\a[23] ), .ZN(new_n7045_));
  AOI21_X1   g06981(.A1(new_n7042_), .A2(new_n7043_), .B(new_n7041_), .ZN(new_n7046_));
  NOR3_X1    g06982(.A1(new_n7033_), .A2(new_n7034_), .A3(new_n7037_), .ZN(new_n7047_));
  NOR3_X1    g06983(.A1(new_n7046_), .A2(new_n7047_), .A3(new_n84_), .ZN(new_n7048_));
  OAI21_X1   g06984(.A1(new_n7045_), .A2(new_n7048_), .B(new_n6988_), .ZN(new_n7049_));
  INV_X1     g06985(.I(new_n6988_), .ZN(new_n7050_));
  OAI21_X1   g06986(.A1(new_n7046_), .A2(new_n7047_), .B(new_n84_), .ZN(new_n7051_));
  NAND3_X1   g06987(.A1(new_n7038_), .A2(new_n7044_), .A3(\a[23] ), .ZN(new_n7052_));
  NAND3_X1   g06988(.A1(new_n7052_), .A2(new_n7051_), .A3(new_n7050_), .ZN(new_n7053_));
  AOI21_X1   g06989(.A1(new_n6701_), .A2(new_n6698_), .B(new_n6692_), .ZN(new_n7054_));
  AOI21_X1   g06990(.A1(new_n6651_), .A2(new_n6705_), .B(new_n7054_), .ZN(new_n7055_));
  NAND3_X1   g06991(.A1(new_n7049_), .A2(new_n7053_), .A3(new_n7055_), .ZN(new_n7056_));
  AOI21_X1   g06992(.A1(new_n7052_), .A2(new_n7051_), .B(new_n7050_), .ZN(new_n7057_));
  NOR3_X1    g06993(.A1(new_n7045_), .A2(new_n7048_), .A3(new_n6988_), .ZN(new_n7058_));
  NAND2_X1   g06994(.A1(new_n6705_), .A2(new_n6651_), .ZN(new_n7059_));
  NAND2_X1   g06995(.A1(new_n7059_), .A2(new_n6706_), .ZN(new_n7060_));
  OAI21_X1   g06996(.A1(new_n7057_), .A2(new_n7058_), .B(new_n7060_), .ZN(new_n7061_));
  AOI21_X1   g06997(.A1(new_n7061_), .A2(new_n7056_), .B(new_n6986_), .ZN(new_n7062_));
  INV_X1     g06998(.I(new_n6985_), .ZN(new_n7063_));
  NAND2_X1   g06999(.A1(new_n7063_), .A2(new_n6983_), .ZN(new_n7064_));
  OAI21_X1   g07000(.A1(new_n7057_), .A2(new_n7058_), .B(new_n7055_), .ZN(new_n7065_));
  NAND3_X1   g07001(.A1(new_n7049_), .A2(new_n7053_), .A3(new_n7060_), .ZN(new_n7066_));
  AOI21_X1   g07002(.A1(new_n7066_), .A2(new_n7065_), .B(new_n7064_), .ZN(new_n7067_));
  OAI21_X1   g07003(.A1(new_n6649_), .A2(new_n6733_), .B(new_n6723_), .ZN(new_n7068_));
  NOR3_X1    g07004(.A1(new_n7068_), .A2(new_n7062_), .A3(new_n7067_), .ZN(new_n7069_));
  INV_X1     g07005(.I(new_n7069_), .ZN(new_n7070_));
  OAI21_X1   g07006(.A1(new_n7062_), .A2(new_n7067_), .B(new_n7068_), .ZN(new_n7071_));
  AOI21_X1   g07007(.A1(new_n7070_), .A2(new_n7071_), .B(new_n6979_), .ZN(new_n7072_));
  INV_X1     g07008(.I(new_n6979_), .ZN(new_n7073_));
  NOR2_X1    g07009(.A1(new_n7067_), .A2(new_n7062_), .ZN(new_n7074_));
  XOR2_X1    g07010(.A1(new_n7074_), .A2(new_n7068_), .Z(new_n7075_));
  NOR2_X1    g07011(.A1(new_n7075_), .A2(new_n7073_), .ZN(new_n7076_));
  NOR2_X1    g07012(.A1(new_n7076_), .A2(new_n7072_), .ZN(new_n7077_));
  OAI22_X1   g07013(.A1(new_n813_), .A2(new_n6091_), .B1(new_n1008_), .B2(new_n6089_), .ZN(new_n7078_));
  NAND2_X1   g07014(.A1(new_n897_), .A2(new_n6095_), .ZN(new_n7079_));
  AOI21_X1   g07015(.A1(new_n7078_), .A2(new_n7079_), .B(new_n6082_), .ZN(new_n7080_));
  NAND3_X1   g07016(.A1(new_n2917_), .A2(new_n3521_), .A3(new_n7080_), .ZN(new_n7081_));
  OAI21_X1   g07017(.A1(new_n6125_), .A2(new_n6124_), .B(new_n7080_), .ZN(new_n7082_));
  NAND2_X1   g07018(.A1(new_n7082_), .A2(\a[14] ), .ZN(new_n7083_));
  NAND3_X1   g07019(.A1(new_n7083_), .A2(new_n7081_), .A3(new_n6748_), .ZN(new_n7084_));
  NOR2_X1    g07020(.A1(new_n7082_), .A2(\a[14] ), .ZN(new_n7085_));
  AOI21_X1   g07021(.A1(new_n2917_), .A2(new_n7080_), .B(new_n3521_), .ZN(new_n7086_));
  OAI21_X1   g07022(.A1(new_n7085_), .A2(new_n7086_), .B(new_n6738_), .ZN(new_n7087_));
  AOI21_X1   g07023(.A1(new_n7087_), .A2(new_n7084_), .B(new_n7077_), .ZN(new_n7088_));
  INV_X1     g07024(.I(new_n7071_), .ZN(new_n7089_));
  OAI21_X1   g07025(.A1(new_n7069_), .A2(new_n7089_), .B(new_n7073_), .ZN(new_n7090_));
  OAI21_X1   g07026(.A1(new_n7073_), .A2(new_n7075_), .B(new_n7090_), .ZN(new_n7091_));
  NAND3_X1   g07027(.A1(new_n7083_), .A2(new_n7081_), .A3(new_n6738_), .ZN(new_n7092_));
  AOI21_X1   g07028(.A1(new_n7083_), .A2(new_n7081_), .B(new_n6738_), .ZN(new_n7093_));
  INV_X1     g07029(.I(new_n7093_), .ZN(new_n7094_));
  AOI21_X1   g07030(.A1(new_n7094_), .A2(new_n7092_), .B(new_n7091_), .ZN(new_n7095_));
  NOR3_X1    g07031(.A1(new_n7095_), .A2(new_n7088_), .A3(new_n6974_), .ZN(new_n7096_));
  AOI21_X1   g07032(.A1(new_n6753_), .A2(new_n6754_), .B(new_n6762_), .ZN(new_n7097_));
  INV_X1     g07033(.I(new_n7088_), .ZN(new_n7098_));
  INV_X1     g07034(.I(new_n7092_), .ZN(new_n7099_));
  OAI21_X1   g07035(.A1(new_n7099_), .A2(new_n7093_), .B(new_n7077_), .ZN(new_n7100_));
  AOI21_X1   g07036(.A1(new_n7098_), .A2(new_n7100_), .B(new_n7097_), .ZN(new_n7101_));
  OAI21_X1   g07037(.A1(new_n7101_), .A2(new_n7096_), .B(new_n6973_), .ZN(new_n7102_));
  XOR2_X1    g07038(.A1(new_n6972_), .A2(\a[11] ), .Z(new_n7103_));
  NOR3_X1    g07039(.A1(new_n7095_), .A2(new_n7088_), .A3(new_n7097_), .ZN(new_n7104_));
  AOI21_X1   g07040(.A1(new_n7098_), .A2(new_n7100_), .B(new_n6974_), .ZN(new_n7105_));
  OAI21_X1   g07041(.A1(new_n7105_), .A2(new_n7104_), .B(new_n7103_), .ZN(new_n7106_));
  NOR2_X1    g07042(.A1(new_n6756_), .A2(new_n6752_), .ZN(new_n7107_));
  NOR2_X1    g07043(.A1(new_n6638_), .A2(new_n4034_), .ZN(new_n7108_));
  NOR2_X1    g07044(.A1(new_n6637_), .A2(\a[11] ), .ZN(new_n7109_));
  OAI21_X1   g07045(.A1(new_n7108_), .A2(new_n7109_), .B(new_n7107_), .ZN(new_n7110_));
  NAND3_X1   g07046(.A1(new_n7106_), .A2(new_n7102_), .A3(new_n7110_), .ZN(new_n7111_));
  NAND3_X1   g07047(.A1(new_n7098_), .A2(new_n7100_), .A3(new_n7097_), .ZN(new_n7112_));
  OAI21_X1   g07048(.A1(new_n7095_), .A2(new_n7088_), .B(new_n6974_), .ZN(new_n7113_));
  AOI21_X1   g07049(.A1(new_n7112_), .A2(new_n7113_), .B(new_n7103_), .ZN(new_n7114_));
  NAND3_X1   g07050(.A1(new_n7098_), .A2(new_n7100_), .A3(new_n6974_), .ZN(new_n7115_));
  OAI21_X1   g07051(.A1(new_n7095_), .A2(new_n7088_), .B(new_n7097_), .ZN(new_n7116_));
  AOI21_X1   g07052(.A1(new_n7115_), .A2(new_n7116_), .B(new_n6973_), .ZN(new_n7117_));
  INV_X1     g07053(.I(new_n7110_), .ZN(new_n7118_));
  OAI21_X1   g07054(.A1(new_n7114_), .A2(new_n7117_), .B(new_n7118_), .ZN(new_n7119_));
  AOI21_X1   g07055(.A1(new_n7111_), .A2(new_n7119_), .B(new_n6967_), .ZN(new_n7120_));
  NAND3_X1   g07056(.A1(new_n2733_), .A2(new_n4009_), .A3(new_n6963_), .ZN(new_n7121_));
  NAND2_X1   g07057(.A1(new_n6964_), .A2(\a[8] ), .ZN(new_n7122_));
  NAND2_X1   g07058(.A1(new_n7122_), .A2(new_n7121_), .ZN(new_n7123_));
  OAI21_X1   g07059(.A1(new_n7114_), .A2(new_n7117_), .B(new_n7110_), .ZN(new_n7124_));
  NAND3_X1   g07060(.A1(new_n7106_), .A2(new_n7102_), .A3(new_n7118_), .ZN(new_n7125_));
  AOI21_X1   g07061(.A1(new_n7124_), .A2(new_n7125_), .B(new_n7123_), .ZN(new_n7126_));
  NOR3_X1    g07062(.A1(new_n6958_), .A2(new_n7120_), .A3(new_n7126_), .ZN(new_n7127_));
  NOR3_X1    g07063(.A1(new_n7114_), .A2(new_n7117_), .A3(new_n7118_), .ZN(new_n7128_));
  AOI21_X1   g07064(.A1(new_n7106_), .A2(new_n7102_), .B(new_n7110_), .ZN(new_n7129_));
  OAI21_X1   g07065(.A1(new_n7129_), .A2(new_n7128_), .B(new_n7123_), .ZN(new_n7130_));
  AOI21_X1   g07066(.A1(new_n7106_), .A2(new_n7102_), .B(new_n7118_), .ZN(new_n7131_));
  NOR3_X1    g07067(.A1(new_n7114_), .A2(new_n7117_), .A3(new_n7110_), .ZN(new_n7132_));
  OAI21_X1   g07068(.A1(new_n7131_), .A2(new_n7132_), .B(new_n6967_), .ZN(new_n7133_));
  AOI21_X1   g07069(.A1(new_n7133_), .A2(new_n7130_), .B(new_n6957_), .ZN(new_n7134_));
  OAI21_X1   g07070(.A1(new_n7127_), .A2(new_n7134_), .B(new_n6951_), .ZN(new_n7135_));
  NOR3_X1    g07071(.A1(new_n7120_), .A2(new_n7126_), .A3(new_n6957_), .ZN(new_n7136_));
  AOI22_X1   g07072(.A1(new_n7133_), .A2(new_n7130_), .B1(new_n6954_), .B2(new_n6956_), .ZN(new_n7137_));
  OAI21_X1   g07073(.A1(new_n7137_), .A2(new_n7136_), .B(new_n6950_), .ZN(new_n7138_));
  NAND2_X1   g07074(.A1(new_n7135_), .A2(new_n7138_), .ZN(new_n7139_));
  NOR3_X1    g07075(.A1(new_n6946_), .A2(new_n7139_), .A3(new_n6949_), .ZN(new_n7140_));
  AOI22_X1   g07076(.A1(new_n6928_), .A2(new_n6938_), .B1(new_n7135_), .B2(new_n7138_), .ZN(new_n7141_));
  OAI22_X1   g07077(.A1(new_n7141_), .A2(new_n7140_), .B1(new_n6853_), .B2(new_n6939_), .ZN(new_n7142_));
  OAI22_X1   g07078(.A1(new_n3254_), .A2(new_n6836_), .B1(new_n3142_), .B2(new_n6913_), .ZN(new_n7143_));
  INV_X1     g07079(.I(new_n3271_), .ZN(new_n7144_));
  NOR3_X1    g07080(.A1(new_n3249_), .A2(new_n2729_), .A3(new_n3272_), .ZN(new_n7145_));
  OAI22_X1   g07081(.A1(new_n3176_), .A2(new_n6785_), .B1(new_n2665_), .B2(new_n6783_), .ZN(new_n7146_));
  NAND2_X1   g07082(.A1(new_n2728_), .A2(new_n6789_), .ZN(new_n7147_));
  AOI21_X1   g07083(.A1(new_n7146_), .A2(new_n7147_), .B(new_n6776_), .ZN(new_n7148_));
  OAI21_X1   g07084(.A1(new_n7144_), .A2(new_n7145_), .B(new_n7148_), .ZN(new_n7149_));
  NOR2_X1    g07085(.A1(new_n7149_), .A2(\a[8] ), .ZN(new_n7150_));
  AOI21_X1   g07086(.A1(new_n3273_), .A2(new_n7148_), .B(new_n4009_), .ZN(new_n7151_));
  NOR2_X1    g07087(.A1(new_n7150_), .A2(new_n7151_), .ZN(new_n7152_));
  NOR2_X1    g07088(.A1(new_n3073_), .A2(new_n2614_), .ZN(new_n7153_));
  INV_X1     g07089(.I(new_n3070_), .ZN(new_n7154_));
  NAND2_X1   g07090(.A1(new_n7154_), .A2(new_n3071_), .ZN(new_n7155_));
  AOI21_X1   g07091(.A1(new_n7155_), .A2(new_n3069_), .B(new_n2615_), .ZN(new_n7156_));
  OAI22_X1   g07092(.A1(new_n2614_), .A2(new_n4710_), .B1(new_n529_), .B2(new_n4716_), .ZN(new_n7157_));
  NAND2_X1   g07093(.A1(new_n2718_), .A2(new_n4720_), .ZN(new_n7158_));
  AOI21_X1   g07094(.A1(new_n7158_), .A2(new_n7157_), .B(new_n4707_), .ZN(new_n7159_));
  OAI21_X1   g07095(.A1(new_n7153_), .A2(new_n7156_), .B(new_n7159_), .ZN(new_n7160_));
  NOR2_X1    g07096(.A1(new_n7160_), .A2(\a[11] ), .ZN(new_n7161_));
  AOI21_X1   g07097(.A1(new_n3074_), .A2(new_n7159_), .B(new_n4034_), .ZN(new_n7162_));
  AOI21_X1   g07098(.A1(new_n7073_), .A2(new_n7070_), .B(new_n7089_), .ZN(new_n7163_));
  OAI22_X1   g07099(.A1(new_n1008_), .A2(new_n4470_), .B1(new_n1121_), .B2(new_n4291_), .ZN(new_n7164_));
  NAND2_X1   g07100(.A1(new_n1181_), .A2(new_n4298_), .ZN(new_n7165_));
  AOI21_X1   g07101(.A1(new_n7164_), .A2(new_n7165_), .B(new_n4468_), .ZN(new_n7166_));
  NAND3_X1   g07102(.A1(new_n3562_), .A2(new_n3372_), .A3(new_n7166_), .ZN(new_n7167_));
  OAI21_X1   g07103(.A1(new_n6151_), .A2(new_n6152_), .B(new_n7166_), .ZN(new_n7168_));
  NAND2_X1   g07104(.A1(new_n7168_), .A2(\a[17] ), .ZN(new_n7169_));
  OAI22_X1   g07105(.A1(new_n2492_), .A2(new_n4097_), .B1(new_n2408_), .B2(new_n3769_), .ZN(new_n7170_));
  NAND2_X1   g07106(.A1(new_n2454_), .A2(new_n3776_), .ZN(new_n7171_));
  AOI21_X1   g07107(.A1(new_n7171_), .A2(new_n7170_), .B(new_n4095_), .ZN(new_n7172_));
  OAI21_X1   g07108(.A1(new_n3574_), .A2(new_n3576_), .B(new_n7172_), .ZN(new_n7173_));
  NOR2_X1    g07109(.A1(new_n7173_), .A2(\a[20] ), .ZN(new_n7174_));
  INV_X1     g07110(.I(new_n7174_), .ZN(new_n7175_));
  NAND2_X1   g07111(.A1(new_n7173_), .A2(\a[20] ), .ZN(new_n7176_));
  OAI22_X1   g07112(.A1(new_n1409_), .A2(new_n3310_), .B1(new_n2367_), .B2(new_n3780_), .ZN(new_n7177_));
  NAND2_X1   g07113(.A1(new_n1334_), .A2(new_n3782_), .ZN(new_n7178_));
  AOI21_X1   g07114(.A1(new_n7177_), .A2(new_n7178_), .B(new_n3302_), .ZN(new_n7179_));
  OAI21_X1   g07115(.A1(new_n5634_), .A2(new_n5633_), .B(new_n7179_), .ZN(new_n7180_));
  NOR2_X1    g07116(.A1(new_n7180_), .A2(\a[23] ), .ZN(new_n7181_));
  NAND2_X1   g07117(.A1(new_n7180_), .A2(\a[23] ), .ZN(new_n7182_));
  INV_X1     g07118(.I(new_n7182_), .ZN(new_n7183_));
  OAI22_X1   g07119(.A1(new_n1453_), .A2(new_n3318_), .B1(new_n2351_), .B2(new_n3322_), .ZN(new_n7184_));
  NAND2_X1   g07120(.A1(new_n2310_), .A2(new_n3267_), .ZN(new_n7185_));
  AOI21_X1   g07121(.A1(new_n7185_), .A2(new_n7184_), .B(new_n3260_), .ZN(new_n7186_));
  NAND3_X1   g07122(.A1(new_n4231_), .A2(new_n72_), .A3(new_n7186_), .ZN(new_n7187_));
  OAI21_X1   g07123(.A1(new_n5684_), .A2(new_n4229_), .B(new_n7186_), .ZN(new_n7188_));
  NAND2_X1   g07124(.A1(new_n7188_), .A2(\a[26] ), .ZN(new_n7189_));
  NAND2_X1   g07125(.A1(new_n7189_), .A2(new_n7187_), .ZN(new_n7190_));
  AOI21_X1   g07126(.A1(new_n6999_), .A2(new_n6996_), .B(new_n7009_), .ZN(new_n7191_));
  NOR2_X1    g07127(.A1(new_n7191_), .A2(new_n7027_), .ZN(new_n7192_));
  AOI22_X1   g07128(.A1(new_n4586_), .A2(new_n4589_), .B1(new_n4605_), .B2(new_n4607_), .ZN(new_n7193_));
  INV_X1     g07129(.I(new_n7193_), .ZN(new_n7194_));
  XOR2_X1    g07130(.A1(new_n4603_), .A2(\a[2] ), .Z(new_n7195_));
  INV_X1     g07131(.I(new_n7195_), .ZN(new_n7196_));
  NAND3_X1   g07132(.A1(new_n4586_), .A2(new_n4589_), .A3(new_n7196_), .ZN(new_n7197_));
  NOR2_X1    g07133(.A1(new_n2103_), .A2(new_n2771_), .ZN(new_n7198_));
  INV_X1     g07134(.I(new_n7198_), .ZN(new_n7199_));
  AOI22_X1   g07135(.A1(new_n2161_), .A2(new_n3189_), .B1(new_n2202_), .B2(new_n3332_), .ZN(new_n7200_));
  NAND4_X1   g07136(.A1(new_n5351_), .A2(new_n2764_), .A3(new_n7199_), .A4(new_n7200_), .ZN(new_n7201_));
  NAND3_X1   g07137(.A1(new_n7194_), .A2(new_n7197_), .A3(new_n7201_), .ZN(new_n7202_));
  INV_X1     g07138(.I(new_n7202_), .ZN(new_n7203_));
  INV_X1     g07139(.I(new_n7197_), .ZN(new_n7204_));
  INV_X1     g07140(.I(new_n7201_), .ZN(new_n7205_));
  OAI21_X1   g07141(.A1(new_n7204_), .A2(new_n7193_), .B(new_n7205_), .ZN(new_n7206_));
  INV_X1     g07142(.I(new_n7206_), .ZN(new_n7207_));
  NOR2_X1    g07143(.A1(new_n7203_), .A2(new_n7207_), .ZN(new_n7208_));
  OAI21_X1   g07144(.A1(new_n7013_), .A2(new_n6672_), .B(new_n7010_), .ZN(new_n7209_));
  OAI21_X1   g07145(.A1(new_n7204_), .A2(new_n7193_), .B(new_n7201_), .ZN(new_n7210_));
  NAND3_X1   g07146(.A1(new_n7194_), .A2(new_n7197_), .A3(new_n7205_), .ZN(new_n7211_));
  NAND2_X1   g07147(.A1(new_n7211_), .A2(new_n7210_), .ZN(new_n7212_));
  NAND3_X1   g07148(.A1(new_n7209_), .A2(new_n7011_), .A3(new_n7212_), .ZN(new_n7213_));
  OAI21_X1   g07149(.A1(new_n7192_), .A2(new_n7208_), .B(new_n7213_), .ZN(new_n7214_));
  OAI22_X1   g07150(.A1(new_n2251_), .A2(new_n3175_), .B1(new_n4365_), .B2(new_n2742_), .ZN(new_n7215_));
  NAND2_X1   g07151(.A1(new_n1504_), .A2(new_n2746_), .ZN(new_n7216_));
  AOI21_X1   g07152(.A1(new_n7215_), .A2(new_n7216_), .B(new_n2737_), .ZN(new_n7217_));
  NAND3_X1   g07153(.A1(new_n4650_), .A2(new_n74_), .A3(new_n7217_), .ZN(new_n7218_));
  AOI21_X1   g07154(.A1(new_n4650_), .A2(new_n7217_), .B(new_n74_), .ZN(new_n7219_));
  INV_X1     g07155(.I(new_n7219_), .ZN(new_n7220_));
  NAND2_X1   g07156(.A1(new_n7220_), .A2(new_n7218_), .ZN(new_n7221_));
  NOR2_X1    g07157(.A1(new_n7214_), .A2(new_n7221_), .ZN(new_n7222_));
  AOI22_X1   g07158(.A1(new_n7209_), .A2(new_n7011_), .B1(new_n7202_), .B2(new_n7206_), .ZN(new_n7223_));
  INV_X1     g07159(.I(new_n7212_), .ZN(new_n7224_));
  NOR3_X1    g07160(.A1(new_n7224_), .A2(new_n7191_), .A3(new_n7027_), .ZN(new_n7225_));
  NOR2_X1    g07161(.A1(new_n7225_), .A2(new_n7223_), .ZN(new_n7226_));
  INV_X1     g07162(.I(new_n7218_), .ZN(new_n7227_));
  NOR2_X1    g07163(.A1(new_n7227_), .A2(new_n7219_), .ZN(new_n7228_));
  NOR2_X1    g07164(.A1(new_n7226_), .A2(new_n7228_), .ZN(new_n7229_));
  OAI21_X1   g07165(.A1(new_n7222_), .A2(new_n7229_), .B(new_n7190_), .ZN(new_n7230_));
  NOR2_X1    g07166(.A1(new_n7188_), .A2(\a[26] ), .ZN(new_n7231_));
  AOI21_X1   g07167(.A1(new_n4231_), .A2(new_n7186_), .B(new_n72_), .ZN(new_n7232_));
  NOR2_X1    g07168(.A1(new_n7231_), .A2(new_n7232_), .ZN(new_n7233_));
  NOR2_X1    g07169(.A1(new_n7226_), .A2(new_n7221_), .ZN(new_n7234_));
  NOR2_X1    g07170(.A1(new_n7214_), .A2(new_n7228_), .ZN(new_n7235_));
  OAI21_X1   g07171(.A1(new_n7234_), .A2(new_n7235_), .B(new_n7233_), .ZN(new_n7236_));
  INV_X1     g07172(.I(new_n7024_), .ZN(new_n7237_));
  AOI21_X1   g07173(.A1(new_n6995_), .A2(new_n7022_), .B(new_n7237_), .ZN(new_n7238_));
  NAND3_X1   g07174(.A1(new_n7236_), .A2(new_n7230_), .A3(new_n7238_), .ZN(new_n7239_));
  INV_X1     g07175(.I(new_n7239_), .ZN(new_n7240_));
  AOI21_X1   g07176(.A1(new_n7236_), .A2(new_n7230_), .B(new_n7238_), .ZN(new_n7241_));
  OAI22_X1   g07177(.A1(new_n7240_), .A2(new_n7241_), .B1(new_n7183_), .B2(new_n7181_), .ZN(new_n7242_));
  INV_X1     g07178(.I(new_n7181_), .ZN(new_n7243_));
  INV_X1     g07179(.I(new_n7222_), .ZN(new_n7244_));
  NAND2_X1   g07180(.A1(new_n7214_), .A2(new_n7221_), .ZN(new_n7245_));
  AOI21_X1   g07181(.A1(new_n7244_), .A2(new_n7245_), .B(new_n7233_), .ZN(new_n7246_));
  NOR2_X1    g07182(.A1(new_n7234_), .A2(new_n7235_), .ZN(new_n7247_));
  NOR2_X1    g07183(.A1(new_n7247_), .A2(new_n7190_), .ZN(new_n7248_));
  OAI21_X1   g07184(.A1(new_n7248_), .A2(new_n7246_), .B(new_n7238_), .ZN(new_n7249_));
  INV_X1     g07185(.I(new_n7238_), .ZN(new_n7250_));
  NAND3_X1   g07186(.A1(new_n7236_), .A2(new_n7230_), .A3(new_n7250_), .ZN(new_n7251_));
  NAND2_X1   g07187(.A1(new_n7249_), .A2(new_n7251_), .ZN(new_n7252_));
  NAND3_X1   g07188(.A1(new_n7252_), .A2(new_n7243_), .A3(new_n7182_), .ZN(new_n7253_));
  NOR2_X1    g07189(.A1(new_n7041_), .A2(new_n6988_), .ZN(new_n7254_));
  NAND2_X1   g07190(.A1(new_n7041_), .A2(new_n6988_), .ZN(new_n7255_));
  OAI21_X1   g07191(.A1(new_n7034_), .A2(new_n7037_), .B(\a[23] ), .ZN(new_n7256_));
  NAND3_X1   g07192(.A1(new_n7042_), .A2(new_n84_), .A3(new_n7043_), .ZN(new_n7257_));
  NAND2_X1   g07193(.A1(new_n7256_), .A2(new_n7257_), .ZN(new_n7258_));
  AOI21_X1   g07194(.A1(new_n7258_), .A2(new_n7255_), .B(new_n7254_), .ZN(new_n7259_));
  NAND3_X1   g07195(.A1(new_n7253_), .A2(new_n7242_), .A3(new_n7259_), .ZN(new_n7260_));
  INV_X1     g07196(.I(new_n7241_), .ZN(new_n7261_));
  AOI22_X1   g07197(.A1(new_n7261_), .A2(new_n7239_), .B1(new_n7243_), .B2(new_n7182_), .ZN(new_n7262_));
  NAND2_X1   g07198(.A1(new_n7243_), .A2(new_n7182_), .ZN(new_n7263_));
  AOI21_X1   g07199(.A1(new_n7236_), .A2(new_n7230_), .B(new_n7250_), .ZN(new_n7264_));
  NOR3_X1    g07200(.A1(new_n7248_), .A2(new_n7246_), .A3(new_n7238_), .ZN(new_n7265_));
  NOR2_X1    g07201(.A1(new_n7265_), .A2(new_n7264_), .ZN(new_n7266_));
  NOR2_X1    g07202(.A1(new_n7263_), .A2(new_n7266_), .ZN(new_n7267_));
  INV_X1     g07203(.I(new_n7254_), .ZN(new_n7268_));
  AOI21_X1   g07204(.A1(new_n7042_), .A2(new_n7043_), .B(new_n84_), .ZN(new_n7269_));
  NOR3_X1    g07205(.A1(new_n7034_), .A2(\a[23] ), .A3(new_n7037_), .ZN(new_n7270_));
  OAI21_X1   g07206(.A1(new_n7269_), .A2(new_n7270_), .B(new_n7255_), .ZN(new_n7271_));
  NAND2_X1   g07207(.A1(new_n7271_), .A2(new_n7268_), .ZN(new_n7272_));
  OAI21_X1   g07208(.A1(new_n7267_), .A2(new_n7262_), .B(new_n7272_), .ZN(new_n7273_));
  AOI22_X1   g07209(.A1(new_n7175_), .A2(new_n7176_), .B1(new_n7273_), .B2(new_n7260_), .ZN(new_n7274_));
  NAND2_X1   g07210(.A1(new_n7175_), .A2(new_n7176_), .ZN(new_n7275_));
  AOI21_X1   g07211(.A1(new_n7253_), .A2(new_n7242_), .B(new_n7272_), .ZN(new_n7276_));
  NOR3_X1    g07212(.A1(new_n7267_), .A2(new_n7262_), .A3(new_n7259_), .ZN(new_n7277_));
  NOR2_X1    g07213(.A1(new_n7277_), .A2(new_n7276_), .ZN(new_n7278_));
  NOR2_X1    g07214(.A1(new_n7275_), .A2(new_n7278_), .ZN(new_n7279_));
  NOR3_X1    g07215(.A1(new_n7057_), .A2(new_n7058_), .A3(new_n7060_), .ZN(new_n7280_));
  OAI21_X1   g07216(.A1(new_n6986_), .A2(new_n7280_), .B(new_n7061_), .ZN(new_n7281_));
  NOR3_X1    g07217(.A1(new_n7279_), .A2(new_n7274_), .A3(new_n7281_), .ZN(new_n7282_));
  INV_X1     g07218(.I(new_n7176_), .ZN(new_n7283_));
  NOR3_X1    g07219(.A1(new_n7267_), .A2(new_n7262_), .A3(new_n7272_), .ZN(new_n7284_));
  AOI21_X1   g07220(.A1(new_n7253_), .A2(new_n7242_), .B(new_n7259_), .ZN(new_n7285_));
  OAI22_X1   g07221(.A1(new_n7174_), .A2(new_n7283_), .B1(new_n7284_), .B2(new_n7285_), .ZN(new_n7286_));
  OAI21_X1   g07222(.A1(new_n7267_), .A2(new_n7262_), .B(new_n7259_), .ZN(new_n7287_));
  NAND3_X1   g07223(.A1(new_n7253_), .A2(new_n7242_), .A3(new_n7272_), .ZN(new_n7288_));
  NAND2_X1   g07224(.A1(new_n7287_), .A2(new_n7288_), .ZN(new_n7289_));
  NAND3_X1   g07225(.A1(new_n7289_), .A2(new_n7175_), .A3(new_n7176_), .ZN(new_n7290_));
  AOI21_X1   g07226(.A1(new_n7049_), .A2(new_n7053_), .B(new_n7055_), .ZN(new_n7291_));
  AOI21_X1   g07227(.A1(new_n7064_), .A2(new_n7056_), .B(new_n7291_), .ZN(new_n7292_));
  AOI21_X1   g07228(.A1(new_n7290_), .A2(new_n7286_), .B(new_n7292_), .ZN(new_n7293_));
  NOR2_X1    g07229(.A1(new_n7282_), .A2(new_n7293_), .ZN(new_n7294_));
  AOI21_X1   g07230(.A1(new_n7167_), .A2(new_n7169_), .B(new_n7294_), .ZN(new_n7295_));
  NOR2_X1    g07231(.A1(new_n7168_), .A2(\a[17] ), .ZN(new_n7296_));
  AOI21_X1   g07232(.A1(new_n3562_), .A2(new_n7166_), .B(new_n3372_), .ZN(new_n7297_));
  AOI21_X1   g07233(.A1(new_n7290_), .A2(new_n7286_), .B(new_n7281_), .ZN(new_n7298_));
  NOR3_X1    g07234(.A1(new_n7279_), .A2(new_n7274_), .A3(new_n7292_), .ZN(new_n7299_));
  NOR2_X1    g07235(.A1(new_n7299_), .A2(new_n7298_), .ZN(new_n7300_));
  NOR3_X1    g07236(.A1(new_n7300_), .A2(new_n7296_), .A3(new_n7297_), .ZN(new_n7301_));
  OAI21_X1   g07237(.A1(new_n813_), .A2(new_n6094_), .B(new_n6081_), .ZN(new_n7302_));
  OAI22_X1   g07238(.A1(new_n2559_), .A2(new_n6091_), .B1(new_n896_), .B2(new_n6089_), .ZN(new_n7303_));
  NOR2_X1    g07239(.A1(new_n7303_), .A2(new_n7302_), .ZN(new_n7304_));
  OAI21_X1   g07240(.A1(new_n3622_), .A2(new_n3623_), .B(new_n7304_), .ZN(new_n7305_));
  OAI21_X1   g07241(.A1(new_n7295_), .A2(new_n7301_), .B(new_n7305_), .ZN(new_n7306_));
  OAI22_X1   g07242(.A1(new_n7296_), .A2(new_n7297_), .B1(new_n7282_), .B2(new_n7293_), .ZN(new_n7307_));
  OAI21_X1   g07243(.A1(new_n7279_), .A2(new_n7274_), .B(new_n7292_), .ZN(new_n7308_));
  NAND3_X1   g07244(.A1(new_n7290_), .A2(new_n7281_), .A3(new_n7286_), .ZN(new_n7309_));
  NAND2_X1   g07245(.A1(new_n7308_), .A2(new_n7309_), .ZN(new_n7310_));
  NAND3_X1   g07246(.A1(new_n7310_), .A2(new_n7169_), .A3(new_n7167_), .ZN(new_n7311_));
  NAND4_X1   g07247(.A1(new_n3624_), .A2(new_n7307_), .A3(new_n7311_), .A4(new_n7304_), .ZN(new_n7312_));
  AOI21_X1   g07248(.A1(new_n7312_), .A2(new_n7306_), .B(\a[14] ), .ZN(new_n7313_));
  AOI22_X1   g07249(.A1(new_n3624_), .A2(new_n7304_), .B1(new_n7311_), .B2(new_n7307_), .ZN(new_n7314_));
  NOR3_X1    g07250(.A1(new_n7295_), .A2(new_n7301_), .A3(new_n7305_), .ZN(new_n7315_));
  NOR3_X1    g07251(.A1(new_n7314_), .A2(new_n7315_), .A3(new_n3521_), .ZN(new_n7316_));
  OAI21_X1   g07252(.A1(new_n7316_), .A2(new_n7313_), .B(new_n7163_), .ZN(new_n7317_));
  INV_X1     g07253(.I(new_n7163_), .ZN(new_n7318_));
  OAI21_X1   g07254(.A1(new_n7314_), .A2(new_n7315_), .B(new_n3521_), .ZN(new_n7319_));
  NAND3_X1   g07255(.A1(new_n7312_), .A2(new_n7306_), .A3(\a[14] ), .ZN(new_n7320_));
  NAND3_X1   g07256(.A1(new_n7319_), .A2(new_n7320_), .A3(new_n7318_), .ZN(new_n7321_));
  AOI21_X1   g07257(.A1(new_n7083_), .A2(new_n7081_), .B(new_n6748_), .ZN(new_n7322_));
  AOI21_X1   g07258(.A1(new_n7091_), .A2(new_n7084_), .B(new_n7322_), .ZN(new_n7323_));
  NAND3_X1   g07259(.A1(new_n7317_), .A2(new_n7321_), .A3(new_n7323_), .ZN(new_n7324_));
  AOI21_X1   g07260(.A1(new_n7319_), .A2(new_n7320_), .B(new_n7318_), .ZN(new_n7325_));
  NOR3_X1    g07261(.A1(new_n7316_), .A2(new_n7313_), .A3(new_n7163_), .ZN(new_n7326_));
  NOR3_X1    g07262(.A1(new_n7085_), .A2(new_n7086_), .A3(new_n6738_), .ZN(new_n7327_));
  OAI21_X1   g07263(.A1(new_n7077_), .A2(new_n7327_), .B(new_n7087_), .ZN(new_n7328_));
  OAI21_X1   g07264(.A1(new_n7326_), .A2(new_n7325_), .B(new_n7328_), .ZN(new_n7329_));
  NAND2_X1   g07265(.A1(new_n7329_), .A2(new_n7324_), .ZN(new_n7330_));
  OAI21_X1   g07266(.A1(new_n7161_), .A2(new_n7162_), .B(new_n7330_), .ZN(new_n7331_));
  NAND3_X1   g07267(.A1(new_n3074_), .A2(new_n4034_), .A3(new_n7159_), .ZN(new_n7332_));
  NAND2_X1   g07268(.A1(new_n7160_), .A2(\a[11] ), .ZN(new_n7333_));
  OAI21_X1   g07269(.A1(new_n7326_), .A2(new_n7325_), .B(new_n7323_), .ZN(new_n7334_));
  NAND3_X1   g07270(.A1(new_n7317_), .A2(new_n7321_), .A3(new_n7328_), .ZN(new_n7335_));
  NAND2_X1   g07271(.A1(new_n7334_), .A2(new_n7335_), .ZN(new_n7336_));
  NAND3_X1   g07272(.A1(new_n7336_), .A2(new_n7332_), .A3(new_n7333_), .ZN(new_n7337_));
  AOI21_X1   g07273(.A1(new_n6973_), .A2(new_n7112_), .B(new_n7101_), .ZN(new_n7338_));
  NAND3_X1   g07274(.A1(new_n7331_), .A2(new_n7337_), .A3(new_n7338_), .ZN(new_n7339_));
  AOI22_X1   g07275(.A1(new_n7332_), .A2(new_n7333_), .B1(new_n7324_), .B2(new_n7329_), .ZN(new_n7340_));
  AOI21_X1   g07276(.A1(new_n7317_), .A2(new_n7321_), .B(new_n7328_), .ZN(new_n7341_));
  NOR3_X1    g07277(.A1(new_n7326_), .A2(new_n7325_), .A3(new_n7323_), .ZN(new_n7342_));
  NOR2_X1    g07278(.A1(new_n7342_), .A2(new_n7341_), .ZN(new_n7343_));
  NOR3_X1    g07279(.A1(new_n7343_), .A2(new_n7161_), .A3(new_n7162_), .ZN(new_n7344_));
  INV_X1     g07280(.I(new_n7338_), .ZN(new_n7345_));
  OAI21_X1   g07281(.A1(new_n7344_), .A2(new_n7340_), .B(new_n7345_), .ZN(new_n7346_));
  AOI21_X1   g07282(.A1(new_n7339_), .A2(new_n7346_), .B(new_n7152_), .ZN(new_n7347_));
  NAND3_X1   g07283(.A1(new_n3273_), .A2(new_n4009_), .A3(new_n7148_), .ZN(new_n7348_));
  NAND2_X1   g07284(.A1(new_n7149_), .A2(\a[8] ), .ZN(new_n7349_));
  NAND2_X1   g07285(.A1(new_n7349_), .A2(new_n7348_), .ZN(new_n7350_));
  OAI21_X1   g07286(.A1(new_n7344_), .A2(new_n7340_), .B(new_n7338_), .ZN(new_n7351_));
  NAND3_X1   g07287(.A1(new_n7331_), .A2(new_n7337_), .A3(new_n7345_), .ZN(new_n7352_));
  AOI21_X1   g07288(.A1(new_n7351_), .A2(new_n7352_), .B(new_n7350_), .ZN(new_n7353_));
  AOI21_X1   g07289(.A1(new_n7123_), .A2(new_n7111_), .B(new_n7129_), .ZN(new_n7354_));
  NOR3_X1    g07290(.A1(new_n7347_), .A2(new_n7353_), .A3(new_n7354_), .ZN(new_n7355_));
  NOR3_X1    g07291(.A1(new_n7344_), .A2(new_n7345_), .A3(new_n7340_), .ZN(new_n7356_));
  AOI21_X1   g07292(.A1(new_n7331_), .A2(new_n7337_), .B(new_n7338_), .ZN(new_n7357_));
  OAI21_X1   g07293(.A1(new_n7356_), .A2(new_n7357_), .B(new_n7350_), .ZN(new_n7358_));
  INV_X1     g07294(.I(new_n7351_), .ZN(new_n7359_));
  NOR3_X1    g07295(.A1(new_n7344_), .A2(new_n7340_), .A3(new_n7338_), .ZN(new_n7360_));
  OAI21_X1   g07296(.A1(new_n7359_), .A2(new_n7360_), .B(new_n7152_), .ZN(new_n7361_));
  INV_X1     g07297(.I(new_n7354_), .ZN(new_n7362_));
  AOI21_X1   g07298(.A1(new_n7361_), .A2(new_n7358_), .B(new_n7362_), .ZN(new_n7363_));
  OAI21_X1   g07299(.A1(new_n7363_), .A2(new_n7355_), .B(new_n65_), .ZN(new_n7364_));
  NAND3_X1   g07300(.A1(new_n7361_), .A2(new_n7358_), .A3(new_n7362_), .ZN(new_n7365_));
  OAI21_X1   g07301(.A1(new_n7347_), .A2(new_n7353_), .B(new_n7354_), .ZN(new_n7366_));
  NAND3_X1   g07302(.A1(new_n7365_), .A2(new_n7366_), .A3(\a[5] ), .ZN(new_n7367_));
  AOI21_X1   g07303(.A1(new_n7364_), .A2(new_n7367_), .B(new_n7143_), .ZN(new_n7368_));
  INV_X1     g07304(.I(new_n7143_), .ZN(new_n7369_));
  AOI21_X1   g07305(.A1(new_n7365_), .A2(new_n7366_), .B(\a[5] ), .ZN(new_n7370_));
  NOR3_X1    g07306(.A1(new_n7363_), .A2(new_n7355_), .A3(new_n65_), .ZN(new_n7371_));
  NOR3_X1    g07307(.A1(new_n7371_), .A2(new_n7370_), .A3(new_n7369_), .ZN(new_n7372_));
  NOR2_X1    g07308(.A1(new_n7136_), .A2(new_n6950_), .ZN(new_n7373_));
  NOR2_X1    g07309(.A1(new_n7373_), .A2(new_n7137_), .ZN(new_n7374_));
  INV_X1     g07310(.I(new_n7374_), .ZN(new_n7375_));
  NOR3_X1    g07311(.A1(new_n7372_), .A2(new_n7368_), .A3(new_n7375_), .ZN(new_n7376_));
  OAI21_X1   g07312(.A1(new_n7372_), .A2(new_n7368_), .B(new_n7375_), .ZN(new_n7377_));
  OAI21_X1   g07313(.A1(new_n7142_), .A2(new_n7376_), .B(new_n7377_), .ZN(new_n7378_));
  INV_X1     g07314(.I(new_n7329_), .ZN(new_n7379_));
  NOR2_X1    g07315(.A1(new_n7326_), .A2(new_n7325_), .ZN(new_n7380_));
  AOI22_X1   g07316(.A1(new_n7332_), .A2(new_n7333_), .B1(new_n7380_), .B2(new_n7323_), .ZN(new_n7381_));
  NOR2_X1    g07317(.A1(new_n7381_), .A2(new_n7379_), .ZN(new_n7382_));
  INV_X1     g07318(.I(new_n7382_), .ZN(new_n7383_));
  OAI22_X1   g07319(.A1(new_n813_), .A2(new_n6089_), .B1(new_n529_), .B2(new_n6091_), .ZN(new_n7384_));
  NAND2_X1   g07320(.A1(new_n2563_), .A2(new_n6095_), .ZN(new_n7385_));
  AOI21_X1   g07321(.A1(new_n7385_), .A2(new_n7384_), .B(new_n6082_), .ZN(new_n7386_));
  NAND2_X1   g07322(.A1(new_n3051_), .A2(new_n7386_), .ZN(new_n7387_));
  XOR2_X1    g07323(.A1(new_n7387_), .A2(\a[14] ), .Z(new_n7388_));
  INV_X1     g07324(.I(new_n7388_), .ZN(new_n7389_));
  OAI22_X1   g07325(.A1(new_n896_), .A2(new_n4470_), .B1(new_n1180_), .B2(new_n4291_), .ZN(new_n7390_));
  NAND2_X1   g07326(.A1(new_n2504_), .A2(new_n4298_), .ZN(new_n7391_));
  AOI21_X1   g07327(.A1(new_n7391_), .A2(new_n7390_), .B(new_n4468_), .ZN(new_n7392_));
  NAND2_X1   g07328(.A1(new_n3596_), .A2(new_n7392_), .ZN(new_n7393_));
  XOR2_X1    g07329(.A1(new_n7393_), .A2(\a[17] ), .Z(new_n7394_));
  INV_X1     g07330(.I(new_n7293_), .ZN(new_n7395_));
  OAI22_X1   g07331(.A1(new_n1121_), .A2(new_n4097_), .B1(new_n2451_), .B2(new_n3769_), .ZN(new_n7396_));
  NAND2_X1   g07332(.A1(new_n2496_), .A2(new_n3776_), .ZN(new_n7397_));
  AOI21_X1   g07333(.A1(new_n7396_), .A2(new_n7397_), .B(new_n4095_), .ZN(new_n7398_));
  NAND2_X1   g07334(.A1(new_n3393_), .A2(new_n7398_), .ZN(new_n7399_));
  XOR2_X1    g07335(.A1(new_n7399_), .A2(\a[20] ), .Z(new_n7400_));
  OAI22_X1   g07336(.A1(new_n2367_), .A2(new_n3306_), .B1(new_n2408_), .B2(new_n3780_), .ZN(new_n7401_));
  NAND2_X1   g07337(.A1(new_n1334_), .A2(new_n5291_), .ZN(new_n7402_));
  AOI21_X1   g07338(.A1(new_n7401_), .A2(new_n7402_), .B(new_n3302_), .ZN(new_n7403_));
  NAND2_X1   g07339(.A1(new_n3708_), .A2(new_n7403_), .ZN(new_n7404_));
  XOR2_X1    g07340(.A1(new_n7404_), .A2(\a[23] ), .Z(new_n7405_));
  OAI22_X1   g07341(.A1(new_n1409_), .A2(new_n3318_), .B1(new_n2351_), .B2(new_n3268_), .ZN(new_n7406_));
  NAND2_X1   g07342(.A1(new_n2359_), .A2(new_n3323_), .ZN(new_n7407_));
  AOI21_X1   g07343(.A1(new_n7406_), .A2(new_n7407_), .B(new_n3260_), .ZN(new_n7408_));
  NAND2_X1   g07344(.A1(new_n3904_), .A2(new_n7408_), .ZN(new_n7409_));
  XOR2_X1    g07345(.A1(new_n7409_), .A2(new_n72_), .Z(new_n7410_));
  OAI21_X1   g07346(.A1(new_n7233_), .A2(new_n7222_), .B(new_n7245_), .ZN(new_n7411_));
  INV_X1     g07347(.I(new_n7411_), .ZN(new_n7412_));
  OAI21_X1   g07348(.A1(new_n7192_), .A2(new_n7203_), .B(new_n7206_), .ZN(new_n7413_));
  INV_X1     g07349(.I(new_n7413_), .ZN(new_n7414_));
  OAI22_X1   g07350(.A1(new_n2311_), .A2(new_n3175_), .B1(new_n4365_), .B2(new_n2747_), .ZN(new_n7415_));
  NAND2_X1   g07351(.A1(new_n2255_), .A2(new_n3275_), .ZN(new_n7416_));
  AOI21_X1   g07352(.A1(new_n7415_), .A2(new_n7416_), .B(new_n2737_), .ZN(new_n7417_));
  NAND2_X1   g07353(.A1(new_n4419_), .A2(new_n7417_), .ZN(new_n7418_));
  XOR2_X1    g07354(.A1(new_n7418_), .A2(new_n74_), .Z(new_n7419_));
  NAND2_X1   g07355(.A1(new_n4629_), .A2(new_n4626_), .ZN(new_n7420_));
  XOR2_X1    g07356(.A1(new_n4625_), .A2(new_n4613_), .Z(new_n7421_));
  NOR2_X1    g07357(.A1(new_n7421_), .A2(new_n4608_), .ZN(new_n7422_));
  AOI21_X1   g07358(.A1(new_n4608_), .A2(new_n7420_), .B(new_n7422_), .ZN(new_n7423_));
  INV_X1     g07359(.I(new_n7423_), .ZN(new_n7424_));
  OR2_X2     g07360(.A1(new_n7419_), .A2(new_n7424_), .Z(new_n7425_));
  NAND2_X1   g07361(.A1(new_n7419_), .A2(new_n7424_), .ZN(new_n7426_));
  AOI21_X1   g07362(.A1(new_n7425_), .A2(new_n7426_), .B(new_n7414_), .ZN(new_n7427_));
  XOR2_X1    g07363(.A1(new_n7419_), .A2(new_n7423_), .Z(new_n7428_));
  NOR2_X1    g07364(.A1(new_n7428_), .A2(new_n7413_), .ZN(new_n7429_));
  NOR2_X1    g07365(.A1(new_n7429_), .A2(new_n7427_), .ZN(new_n7430_));
  XOR2_X1    g07366(.A1(new_n7430_), .A2(new_n7412_), .Z(new_n7431_));
  NAND2_X1   g07367(.A1(new_n7430_), .A2(new_n7412_), .ZN(new_n7432_));
  OAI21_X1   g07368(.A1(new_n7429_), .A2(new_n7427_), .B(new_n7411_), .ZN(new_n7433_));
  AOI21_X1   g07369(.A1(new_n7432_), .A2(new_n7433_), .B(new_n7410_), .ZN(new_n7434_));
  AOI21_X1   g07370(.A1(new_n7431_), .A2(new_n7410_), .B(new_n7434_), .ZN(new_n7435_));
  AOI21_X1   g07371(.A1(new_n7263_), .A2(new_n7239_), .B(new_n7241_), .ZN(new_n7436_));
  NAND2_X1   g07372(.A1(new_n7435_), .A2(new_n7436_), .ZN(new_n7437_));
  NOR2_X1    g07373(.A1(new_n7435_), .A2(new_n7436_), .ZN(new_n7438_));
  INV_X1     g07374(.I(new_n7438_), .ZN(new_n7439_));
  AOI21_X1   g07375(.A1(new_n7439_), .A2(new_n7437_), .B(new_n7405_), .ZN(new_n7440_));
  INV_X1     g07376(.I(new_n7405_), .ZN(new_n7441_));
  INV_X1     g07377(.I(new_n7436_), .ZN(new_n7442_));
  NOR2_X1    g07378(.A1(new_n7435_), .A2(new_n7442_), .ZN(new_n7443_));
  INV_X1     g07379(.I(new_n7443_), .ZN(new_n7444_));
  NAND2_X1   g07380(.A1(new_n7435_), .A2(new_n7442_), .ZN(new_n7445_));
  AOI21_X1   g07381(.A1(new_n7444_), .A2(new_n7445_), .B(new_n7441_), .ZN(new_n7446_));
  NOR2_X1    g07382(.A1(new_n7440_), .A2(new_n7446_), .ZN(new_n7447_));
  AOI21_X1   g07383(.A1(new_n7275_), .A2(new_n7260_), .B(new_n7285_), .ZN(new_n7448_));
  NAND2_X1   g07384(.A1(new_n7447_), .A2(new_n7448_), .ZN(new_n7449_));
  NOR2_X1    g07385(.A1(new_n7447_), .A2(new_n7448_), .ZN(new_n7450_));
  INV_X1     g07386(.I(new_n7450_), .ZN(new_n7451_));
  AOI21_X1   g07387(.A1(new_n7451_), .A2(new_n7449_), .B(new_n7400_), .ZN(new_n7452_));
  INV_X1     g07388(.I(new_n7400_), .ZN(new_n7453_));
  OR2_X2     g07389(.A1(new_n7440_), .A2(new_n7446_), .Z(new_n7454_));
  NAND2_X1   g07390(.A1(new_n7454_), .A2(new_n7448_), .ZN(new_n7455_));
  INV_X1     g07391(.I(new_n7448_), .ZN(new_n7456_));
  NAND2_X1   g07392(.A1(new_n7447_), .A2(new_n7456_), .ZN(new_n7457_));
  AOI21_X1   g07393(.A1(new_n7455_), .A2(new_n7457_), .B(new_n7453_), .ZN(new_n7458_));
  NOR2_X1    g07394(.A1(new_n7452_), .A2(new_n7458_), .ZN(new_n7459_));
  NAND2_X1   g07395(.A1(new_n7290_), .A2(new_n7286_), .ZN(new_n7460_));
  OAI22_X1   g07396(.A1(new_n7296_), .A2(new_n7297_), .B1(new_n7460_), .B2(new_n7281_), .ZN(new_n7461_));
  NAND3_X1   g07397(.A1(new_n7459_), .A2(new_n7395_), .A3(new_n7461_), .ZN(new_n7462_));
  INV_X1     g07398(.I(new_n7449_), .ZN(new_n7463_));
  OAI21_X1   g07399(.A1(new_n7463_), .A2(new_n7450_), .B(new_n7453_), .ZN(new_n7464_));
  NOR2_X1    g07400(.A1(new_n7447_), .A2(new_n7456_), .ZN(new_n7465_));
  NOR2_X1    g07401(.A1(new_n7454_), .A2(new_n7448_), .ZN(new_n7466_));
  OAI21_X1   g07402(.A1(new_n7466_), .A2(new_n7465_), .B(new_n7400_), .ZN(new_n7467_));
  NAND2_X1   g07403(.A1(new_n7464_), .A2(new_n7467_), .ZN(new_n7468_));
  NAND2_X1   g07404(.A1(new_n7461_), .A2(new_n7395_), .ZN(new_n7469_));
  NAND2_X1   g07405(.A1(new_n7468_), .A2(new_n7469_), .ZN(new_n7470_));
  AOI21_X1   g07406(.A1(new_n7462_), .A2(new_n7470_), .B(new_n7394_), .ZN(new_n7471_));
  INV_X1     g07407(.I(new_n7394_), .ZN(new_n7472_));
  NAND3_X1   g07408(.A1(new_n7468_), .A2(new_n7395_), .A3(new_n7461_), .ZN(new_n7473_));
  NAND2_X1   g07409(.A1(new_n7459_), .A2(new_n7469_), .ZN(new_n7474_));
  AOI21_X1   g07410(.A1(new_n7473_), .A2(new_n7474_), .B(new_n7472_), .ZN(new_n7475_));
  AOI21_X1   g07411(.A1(new_n7307_), .A2(new_n7311_), .B(new_n7163_), .ZN(new_n7476_));
  NOR2_X1    g07412(.A1(new_n7295_), .A2(new_n7301_), .ZN(new_n7477_));
  XOR2_X1    g07413(.A1(new_n7305_), .A2(\a[14] ), .Z(new_n7478_));
  AOI21_X1   g07414(.A1(new_n7163_), .A2(new_n7477_), .B(new_n7478_), .ZN(new_n7479_));
  NOR2_X1    g07415(.A1(new_n7479_), .A2(new_n7476_), .ZN(new_n7480_));
  INV_X1     g07416(.I(new_n7480_), .ZN(new_n7481_));
  NOR3_X1    g07417(.A1(new_n7475_), .A2(new_n7471_), .A3(new_n7481_), .ZN(new_n7482_));
  NOR2_X1    g07418(.A1(new_n7475_), .A2(new_n7471_), .ZN(new_n7483_));
  NOR2_X1    g07419(.A1(new_n7483_), .A2(new_n7480_), .ZN(new_n7484_));
  OAI21_X1   g07420(.A1(new_n7484_), .A2(new_n7482_), .B(new_n7389_), .ZN(new_n7485_));
  NOR2_X1    g07421(.A1(new_n7483_), .A2(new_n7481_), .ZN(new_n7486_));
  NOR3_X1    g07422(.A1(new_n7475_), .A2(new_n7471_), .A3(new_n7480_), .ZN(new_n7487_));
  OAI21_X1   g07423(.A1(new_n7486_), .A2(new_n7487_), .B(new_n7388_), .ZN(new_n7488_));
  OAI22_X1   g07424(.A1(new_n694_), .A2(new_n4716_), .B1(new_n2665_), .B2(new_n4710_), .ZN(new_n7489_));
  NAND2_X1   g07425(.A1(new_n2615_), .A2(new_n4720_), .ZN(new_n7490_));
  AOI21_X1   g07426(.A1(new_n7489_), .A2(new_n7490_), .B(new_n4707_), .ZN(new_n7491_));
  NAND2_X1   g07427(.A1(new_n3188_), .A2(new_n7491_), .ZN(new_n7492_));
  XOR2_X1    g07428(.A1(new_n7492_), .A2(\a[11] ), .Z(new_n7493_));
  NAND3_X1   g07429(.A1(new_n7485_), .A2(new_n7488_), .A3(new_n7493_), .ZN(new_n7494_));
  INV_X1     g07430(.I(new_n7494_), .ZN(new_n7495_));
  AOI21_X1   g07431(.A1(new_n7485_), .A2(new_n7488_), .B(new_n7493_), .ZN(new_n7496_));
  OAI21_X1   g07432(.A1(new_n7495_), .A2(new_n7496_), .B(new_n7383_), .ZN(new_n7497_));
  NAND2_X1   g07433(.A1(new_n7485_), .A2(new_n7488_), .ZN(new_n7498_));
  NAND2_X1   g07434(.A1(new_n7498_), .A2(new_n7493_), .ZN(new_n7499_));
  INV_X1     g07435(.I(new_n7499_), .ZN(new_n7500_));
  NOR2_X1    g07436(.A1(new_n7498_), .A2(new_n7493_), .ZN(new_n7501_));
  NOR2_X1    g07437(.A1(new_n7500_), .A2(new_n7501_), .ZN(new_n7502_));
  OAI21_X1   g07438(.A1(new_n7502_), .A2(new_n7383_), .B(new_n7497_), .ZN(new_n7503_));
  OAI21_X1   g07439(.A1(new_n7152_), .A2(new_n7356_), .B(new_n7346_), .ZN(new_n7504_));
  NOR2_X1    g07440(.A1(new_n3142_), .A2(new_n6785_), .ZN(new_n7505_));
  NOR2_X1    g07441(.A1(new_n3176_), .A2(new_n6788_), .ZN(new_n7506_));
  OAI22_X1   g07442(.A1(new_n7506_), .A2(new_n7505_), .B1(new_n2716_), .B2(new_n6783_), .ZN(new_n7507_));
  AOI21_X1   g07443(.A1(new_n3174_), .A2(new_n6775_), .B(new_n7507_), .ZN(new_n7508_));
  NOR2_X1    g07444(.A1(new_n7508_), .A2(new_n7504_), .ZN(new_n7509_));
  AND2_X2    g07445(.A1(new_n7508_), .A2(new_n7504_), .Z(new_n7510_));
  OAI21_X1   g07446(.A1(new_n7510_), .A2(new_n7509_), .B(new_n4009_), .ZN(new_n7511_));
  NOR3_X1    g07447(.A1(new_n7510_), .A2(new_n7509_), .A3(new_n4009_), .ZN(new_n7512_));
  INV_X1     g07448(.I(new_n7512_), .ZN(new_n7513_));
  AOI21_X1   g07449(.A1(new_n7513_), .A2(new_n7511_), .B(new_n7503_), .ZN(new_n7514_));
  INV_X1     g07450(.I(new_n7496_), .ZN(new_n7515_));
  AOI21_X1   g07451(.A1(new_n7515_), .A2(new_n7494_), .B(new_n7382_), .ZN(new_n7516_));
  INV_X1     g07452(.I(new_n7501_), .ZN(new_n7517_));
  NAND2_X1   g07453(.A1(new_n7517_), .A2(new_n7499_), .ZN(new_n7518_));
  AOI21_X1   g07454(.A1(new_n7518_), .A2(new_n7382_), .B(new_n7516_), .ZN(new_n7519_));
  INV_X1     g07455(.I(new_n7511_), .ZN(new_n7520_));
  NOR3_X1    g07456(.A1(new_n7520_), .A2(new_n7519_), .A3(new_n7512_), .ZN(new_n7521_));
  NOR2_X1    g07457(.A1(new_n7347_), .A2(new_n7353_), .ZN(new_n7522_));
  NOR2_X1    g07458(.A1(new_n7522_), .A2(new_n7354_), .ZN(new_n7523_));
  XOR2_X1    g07459(.A1(new_n7143_), .A2(new_n65_), .Z(new_n7524_));
  NOR4_X1    g07460(.A1(new_n7524_), .A2(new_n7347_), .A3(new_n7353_), .A4(new_n7362_), .ZN(new_n7525_));
  NOR2_X1    g07461(.A1(new_n7525_), .A2(new_n7523_), .ZN(new_n7526_));
  OAI21_X1   g07462(.A1(new_n7514_), .A2(new_n7521_), .B(new_n7526_), .ZN(new_n7527_));
  NOR3_X1    g07463(.A1(new_n7514_), .A2(new_n7521_), .A3(new_n7526_), .ZN(new_n7528_));
  AOI21_X1   g07464(.A1(new_n7378_), .A2(new_n7527_), .B(new_n7528_), .ZN(new_n7529_));
  INV_X1     g07465(.I(new_n6783_), .ZN(new_n7530_));
  NAND2_X1   g07466(.A1(new_n3168_), .A2(new_n7530_), .ZN(new_n7531_));
  NAND2_X1   g07467(.A1(new_n3247_), .A2(new_n6789_), .ZN(new_n7532_));
  NAND4_X1   g07468(.A1(new_n3758_), .A2(new_n6775_), .A3(new_n7531_), .A4(new_n7532_), .ZN(new_n7533_));
  XOR2_X1    g07469(.A1(new_n7533_), .A2(\a[8] ), .Z(new_n7534_));
  OAI22_X1   g07470(.A1(new_n2614_), .A2(new_n4716_), .B1(new_n2665_), .B2(new_n4719_), .ZN(new_n7535_));
  NAND2_X1   g07471(.A1(new_n2728_), .A2(new_n4709_), .ZN(new_n7536_));
  AOI21_X1   g07472(.A1(new_n7536_), .A2(new_n7535_), .B(new_n4707_), .ZN(new_n7537_));
  NAND2_X1   g07473(.A1(new_n2733_), .A2(new_n7537_), .ZN(new_n7538_));
  XOR2_X1    g07474(.A1(new_n7538_), .A2(\a[11] ), .Z(new_n7539_));
  OAI22_X1   g07475(.A1(new_n2559_), .A2(new_n6089_), .B1(new_n694_), .B2(new_n6091_), .ZN(new_n7540_));
  NAND2_X1   g07476(.A1(new_n2567_), .A2(new_n6095_), .ZN(new_n7541_));
  AOI21_X1   g07477(.A1(new_n7540_), .A2(new_n7541_), .B(new_n6082_), .ZN(new_n7542_));
  NAND2_X1   g07478(.A1(new_n2759_), .A2(new_n7542_), .ZN(new_n7543_));
  XOR2_X1    g07479(.A1(new_n7543_), .A2(new_n3521_), .Z(new_n7544_));
  INV_X1     g07480(.I(new_n7544_), .ZN(new_n7545_));
  OAI22_X1   g07481(.A1(new_n1180_), .A2(new_n4097_), .B1(new_n2492_), .B2(new_n3769_), .ZN(new_n7546_));
  NAND2_X1   g07482(.A1(new_n1122_), .A2(new_n3776_), .ZN(new_n7547_));
  AOI21_X1   g07483(.A1(new_n7547_), .A2(new_n7546_), .B(new_n4095_), .ZN(new_n7548_));
  NAND2_X1   g07484(.A1(new_n3330_), .A2(new_n7548_), .ZN(new_n7549_));
  XOR2_X1    g07485(.A1(new_n7549_), .A2(new_n3035_), .Z(new_n7550_));
  OAI22_X1   g07486(.A1(new_n2367_), .A2(new_n3310_), .B1(new_n2451_), .B2(new_n3780_), .ZN(new_n7551_));
  NAND2_X1   g07487(.A1(new_n2412_), .A2(new_n3782_), .ZN(new_n7552_));
  AOI21_X1   g07488(.A1(new_n7551_), .A2(new_n7552_), .B(new_n3302_), .ZN(new_n7553_));
  NAND2_X1   g07489(.A1(new_n3403_), .A2(new_n7553_), .ZN(new_n7554_));
  XOR2_X1    g07490(.A1(new_n7554_), .A2(\a[23] ), .Z(new_n7555_));
  OAI22_X1   g07491(.A1(new_n1409_), .A2(new_n3322_), .B1(new_n1333_), .B2(new_n3318_), .ZN(new_n7556_));
  NAND2_X1   g07492(.A1(new_n2359_), .A2(new_n3267_), .ZN(new_n7557_));
  AOI21_X1   g07493(.A1(new_n7556_), .A2(new_n7557_), .B(new_n3260_), .ZN(new_n7558_));
  NAND2_X1   g07494(.A1(new_n3828_), .A2(new_n7558_), .ZN(new_n7559_));
  XOR2_X1    g07495(.A1(new_n7559_), .A2(\a[26] ), .Z(new_n7560_));
  XOR2_X1    g07496(.A1(new_n4540_), .A2(new_n4630_), .Z(new_n7561_));
  OR2_X2     g07497(.A1(new_n4536_), .A2(new_n7561_), .Z(new_n7562_));
  OAI21_X1   g07498(.A1(new_n4633_), .A2(new_n4634_), .B(new_n4536_), .ZN(new_n7563_));
  NAND2_X1   g07499(.A1(new_n7562_), .A2(new_n7563_), .ZN(new_n7564_));
  NAND2_X1   g07500(.A1(new_n7425_), .A2(new_n7413_), .ZN(new_n7565_));
  NAND3_X1   g07501(.A1(new_n7564_), .A2(new_n7426_), .A3(new_n7565_), .ZN(new_n7566_));
  NAND2_X1   g07502(.A1(new_n7565_), .A2(new_n7426_), .ZN(new_n7567_));
  NAND3_X1   g07503(.A1(new_n7567_), .A2(new_n7562_), .A3(new_n7563_), .ZN(new_n7568_));
  AOI21_X1   g07504(.A1(new_n7568_), .A2(new_n7566_), .B(new_n7560_), .ZN(new_n7569_));
  INV_X1     g07505(.I(new_n7560_), .ZN(new_n7570_));
  XOR2_X1    g07506(.A1(new_n7564_), .A2(new_n7567_), .Z(new_n7571_));
  NOR2_X1    g07507(.A1(new_n7571_), .A2(new_n7570_), .ZN(new_n7572_));
  NOR2_X1    g07508(.A1(new_n7572_), .A2(new_n7569_), .ZN(new_n7573_));
  NAND2_X1   g07509(.A1(new_n7432_), .A2(new_n7410_), .ZN(new_n7574_));
  NAND3_X1   g07510(.A1(new_n7573_), .A2(new_n7433_), .A3(new_n7574_), .ZN(new_n7575_));
  NAND2_X1   g07511(.A1(new_n7574_), .A2(new_n7433_), .ZN(new_n7576_));
  OAI21_X1   g07512(.A1(new_n7569_), .A2(new_n7572_), .B(new_n7576_), .ZN(new_n7577_));
  AOI21_X1   g07513(.A1(new_n7575_), .A2(new_n7577_), .B(new_n7555_), .ZN(new_n7578_));
  INV_X1     g07514(.I(new_n7555_), .ZN(new_n7579_));
  XOR2_X1    g07515(.A1(new_n7573_), .A2(new_n7576_), .Z(new_n7580_));
  NOR2_X1    g07516(.A1(new_n7580_), .A2(new_n7579_), .ZN(new_n7581_));
  NOR2_X1    g07517(.A1(new_n7581_), .A2(new_n7578_), .ZN(new_n7582_));
  OAI21_X1   g07518(.A1(new_n7405_), .A2(new_n7443_), .B(new_n7445_), .ZN(new_n7583_));
  INV_X1     g07519(.I(new_n7583_), .ZN(new_n7584_));
  NAND2_X1   g07520(.A1(new_n7582_), .A2(new_n7584_), .ZN(new_n7585_));
  INV_X1     g07521(.I(new_n7585_), .ZN(new_n7586_));
  NOR2_X1    g07522(.A1(new_n7582_), .A2(new_n7584_), .ZN(new_n7587_));
  OAI21_X1   g07523(.A1(new_n7586_), .A2(new_n7587_), .B(new_n7550_), .ZN(new_n7588_));
  XOR2_X1    g07524(.A1(new_n7582_), .A2(new_n7583_), .Z(new_n7589_));
  OAI21_X1   g07525(.A1(new_n7550_), .A2(new_n7589_), .B(new_n7588_), .ZN(new_n7590_));
  OAI22_X1   g07526(.A1(new_n813_), .A2(new_n4470_), .B1(new_n1008_), .B2(new_n4291_), .ZN(new_n7591_));
  NAND2_X1   g07527(.A1(new_n897_), .A2(new_n4298_), .ZN(new_n7592_));
  AOI21_X1   g07528(.A1(new_n7591_), .A2(new_n7592_), .B(new_n4468_), .ZN(new_n7593_));
  NAND2_X1   g07529(.A1(new_n2917_), .A2(new_n7593_), .ZN(new_n7594_));
  XOR2_X1    g07530(.A1(new_n7594_), .A2(\a[17] ), .Z(new_n7595_));
  OAI21_X1   g07531(.A1(new_n7400_), .A2(new_n7465_), .B(new_n7457_), .ZN(new_n7596_));
  INV_X1     g07532(.I(new_n7596_), .ZN(new_n7597_));
  NAND2_X1   g07533(.A1(new_n7595_), .A2(new_n7597_), .ZN(new_n7598_));
  XOR2_X1    g07534(.A1(new_n7594_), .A2(new_n3372_), .Z(new_n7599_));
  NAND2_X1   g07535(.A1(new_n7599_), .A2(new_n7596_), .ZN(new_n7600_));
  NAND2_X1   g07536(.A1(new_n7598_), .A2(new_n7600_), .ZN(new_n7601_));
  NAND2_X1   g07537(.A1(new_n7601_), .A2(new_n7590_), .ZN(new_n7602_));
  INV_X1     g07538(.I(new_n7602_), .ZN(new_n7603_));
  XOR2_X1    g07539(.A1(new_n7595_), .A2(new_n7596_), .Z(new_n7604_));
  NOR2_X1    g07540(.A1(new_n7604_), .A2(new_n7590_), .ZN(new_n7605_));
  NOR2_X1    g07541(.A1(new_n7603_), .A2(new_n7605_), .ZN(new_n7606_));
  NOR2_X1    g07542(.A1(new_n7459_), .A2(new_n7469_), .ZN(new_n7607_));
  OAI21_X1   g07543(.A1(new_n7394_), .A2(new_n7607_), .B(new_n7474_), .ZN(new_n7608_));
  INV_X1     g07544(.I(new_n7608_), .ZN(new_n7609_));
  NAND2_X1   g07545(.A1(new_n7606_), .A2(new_n7609_), .ZN(new_n7610_));
  OAI21_X1   g07546(.A1(new_n7590_), .A2(new_n7604_), .B(new_n7602_), .ZN(new_n7611_));
  NAND2_X1   g07547(.A1(new_n7611_), .A2(new_n7608_), .ZN(new_n7612_));
  AOI21_X1   g07548(.A1(new_n7610_), .A2(new_n7612_), .B(new_n7545_), .ZN(new_n7613_));
  NAND2_X1   g07549(.A1(new_n7611_), .A2(new_n7609_), .ZN(new_n7614_));
  NAND2_X1   g07550(.A1(new_n7606_), .A2(new_n7608_), .ZN(new_n7615_));
  AOI21_X1   g07551(.A1(new_n7615_), .A2(new_n7614_), .B(new_n7544_), .ZN(new_n7616_));
  INV_X1     g07552(.I(new_n7487_), .ZN(new_n7617_));
  OAI21_X1   g07553(.A1(new_n7483_), .A2(new_n7481_), .B(new_n7389_), .ZN(new_n7618_));
  NAND2_X1   g07554(.A1(new_n7618_), .A2(new_n7617_), .ZN(new_n7619_));
  NOR3_X1    g07555(.A1(new_n7613_), .A2(new_n7616_), .A3(new_n7619_), .ZN(new_n7620_));
  INV_X1     g07556(.I(new_n7620_), .ZN(new_n7621_));
  OAI21_X1   g07557(.A1(new_n7613_), .A2(new_n7616_), .B(new_n7619_), .ZN(new_n7622_));
  AOI21_X1   g07558(.A1(new_n7621_), .A2(new_n7622_), .B(new_n7539_), .ZN(new_n7623_));
  INV_X1     g07559(.I(new_n7539_), .ZN(new_n7624_));
  INV_X1     g07560(.I(new_n7619_), .ZN(new_n7625_));
  OAI21_X1   g07561(.A1(new_n7613_), .A2(new_n7616_), .B(new_n7625_), .ZN(new_n7626_));
  NOR2_X1    g07562(.A1(new_n7611_), .A2(new_n7608_), .ZN(new_n7627_));
  INV_X1     g07563(.I(new_n7612_), .ZN(new_n7628_));
  OAI21_X1   g07564(.A1(new_n7628_), .A2(new_n7627_), .B(new_n7544_), .ZN(new_n7629_));
  INV_X1     g07565(.I(new_n7616_), .ZN(new_n7630_));
  NAND3_X1   g07566(.A1(new_n7630_), .A2(new_n7629_), .A3(new_n7619_), .ZN(new_n7631_));
  AOI21_X1   g07567(.A1(new_n7631_), .A2(new_n7626_), .B(new_n7624_), .ZN(new_n7632_));
  AOI21_X1   g07568(.A1(new_n7383_), .A2(new_n7499_), .B(new_n7501_), .ZN(new_n7633_));
  OAI21_X1   g07569(.A1(new_n7623_), .A2(new_n7632_), .B(new_n7633_), .ZN(new_n7634_));
  INV_X1     g07570(.I(new_n7622_), .ZN(new_n7635_));
  OAI21_X1   g07571(.A1(new_n7635_), .A2(new_n7620_), .B(new_n7624_), .ZN(new_n7636_));
  AOI21_X1   g07572(.A1(new_n7630_), .A2(new_n7629_), .B(new_n7619_), .ZN(new_n7637_));
  NOR3_X1    g07573(.A1(new_n7613_), .A2(new_n7616_), .A3(new_n7625_), .ZN(new_n7638_));
  OAI21_X1   g07574(.A1(new_n7637_), .A2(new_n7638_), .B(new_n7539_), .ZN(new_n7639_));
  INV_X1     g07575(.I(new_n7633_), .ZN(new_n7640_));
  NAND3_X1   g07576(.A1(new_n7640_), .A2(new_n7636_), .A3(new_n7639_), .ZN(new_n7641_));
  AOI21_X1   g07577(.A1(new_n7641_), .A2(new_n7634_), .B(new_n7534_), .ZN(new_n7642_));
  INV_X1     g07578(.I(new_n7534_), .ZN(new_n7643_));
  NAND3_X1   g07579(.A1(new_n7636_), .A2(new_n7639_), .A3(new_n7633_), .ZN(new_n7644_));
  OAI21_X1   g07580(.A1(new_n7623_), .A2(new_n7632_), .B(new_n7640_), .ZN(new_n7645_));
  AOI21_X1   g07581(.A1(new_n7645_), .A2(new_n7644_), .B(new_n7643_), .ZN(new_n7646_));
  NOR2_X1    g07582(.A1(new_n7646_), .A2(new_n7642_), .ZN(new_n7647_));
  XOR2_X1    g07583(.A1(new_n7508_), .A2(\a[8] ), .Z(new_n7648_));
  INV_X1     g07584(.I(new_n7648_), .ZN(new_n7649_));
  NAND2_X1   g07585(.A1(new_n7519_), .A2(new_n7649_), .ZN(new_n7650_));
  NAND2_X1   g07586(.A1(new_n7503_), .A2(new_n7648_), .ZN(new_n7651_));
  AOI22_X1   g07587(.A1(new_n7650_), .A2(new_n7651_), .B1(new_n7504_), .B2(new_n7649_), .ZN(new_n7652_));
  NOR2_X1    g07588(.A1(new_n7647_), .A2(new_n7652_), .ZN(new_n7653_));
  NAND2_X1   g07589(.A1(new_n7647_), .A2(new_n7652_), .ZN(new_n7654_));
  OAI21_X1   g07590(.A1(new_n7529_), .A2(new_n7653_), .B(new_n7654_), .ZN(new_n7655_));
  OAI22_X1   g07591(.A1(new_n3254_), .A2(new_n6776_), .B1(new_n3142_), .B2(new_n6783_), .ZN(new_n7656_));
  OAI22_X1   g07592(.A1(new_n3176_), .A2(new_n4710_), .B1(new_n2665_), .B2(new_n4716_), .ZN(new_n7657_));
  NAND2_X1   g07593(.A1(new_n2728_), .A2(new_n4720_), .ZN(new_n7658_));
  AOI21_X1   g07594(.A1(new_n7657_), .A2(new_n7658_), .B(new_n4707_), .ZN(new_n7659_));
  NAND2_X1   g07595(.A1(new_n3273_), .A2(new_n7659_), .ZN(new_n7660_));
  XOR2_X1    g07596(.A1(new_n7660_), .A2(\a[11] ), .Z(new_n7661_));
  OAI22_X1   g07597(.A1(new_n2614_), .A2(new_n6091_), .B1(new_n529_), .B2(new_n6089_), .ZN(new_n7662_));
  NAND2_X1   g07598(.A1(new_n2718_), .A2(new_n6095_), .ZN(new_n7663_));
  AOI21_X1   g07599(.A1(new_n7663_), .A2(new_n7662_), .B(new_n6082_), .ZN(new_n7664_));
  NAND2_X1   g07600(.A1(new_n3074_), .A2(new_n7664_), .ZN(new_n7665_));
  XOR2_X1    g07601(.A1(new_n7665_), .A2(\a[14] ), .Z(new_n7666_));
  OAI22_X1   g07602(.A1(new_n2559_), .A2(new_n4470_), .B1(new_n896_), .B2(new_n4291_), .ZN(new_n7667_));
  NAND2_X1   g07603(.A1(new_n814_), .A2(new_n4298_), .ZN(new_n7668_));
  AOI21_X1   g07604(.A1(new_n7667_), .A2(new_n7668_), .B(new_n4468_), .ZN(new_n7669_));
  NAND2_X1   g07605(.A1(new_n3624_), .A2(new_n7669_), .ZN(new_n7670_));
  XOR2_X1    g07606(.A1(new_n7670_), .A2(\a[17] ), .Z(new_n7671_));
  OAI22_X1   g07607(.A1(new_n1008_), .A2(new_n4097_), .B1(new_n1121_), .B2(new_n3769_), .ZN(new_n7672_));
  NAND2_X1   g07608(.A1(new_n1181_), .A2(new_n3776_), .ZN(new_n7673_));
  AOI21_X1   g07609(.A1(new_n7672_), .A2(new_n7673_), .B(new_n4095_), .ZN(new_n7674_));
  NAND2_X1   g07610(.A1(new_n3562_), .A2(new_n7674_), .ZN(new_n7675_));
  XOR2_X1    g07611(.A1(new_n7675_), .A2(new_n3035_), .Z(new_n7676_));
  OAI22_X1   g07612(.A1(new_n2492_), .A2(new_n3780_), .B1(new_n2408_), .B2(new_n3310_), .ZN(new_n7677_));
  NAND2_X1   g07613(.A1(new_n2454_), .A2(new_n3782_), .ZN(new_n7678_));
  AOI21_X1   g07614(.A1(new_n7678_), .A2(new_n7677_), .B(new_n3302_), .ZN(new_n7679_));
  NAND2_X1   g07615(.A1(new_n3577_), .A2(new_n7679_), .ZN(new_n7680_));
  XOR2_X1    g07616(.A1(new_n7680_), .A2(new_n84_), .Z(new_n7681_));
  OAI22_X1   g07617(.A1(new_n1409_), .A2(new_n3268_), .B1(new_n2367_), .B2(new_n3318_), .ZN(new_n7682_));
  NAND2_X1   g07618(.A1(new_n1334_), .A2(new_n3323_), .ZN(new_n7683_));
  AOI21_X1   g07619(.A1(new_n7682_), .A2(new_n7683_), .B(new_n3260_), .ZN(new_n7684_));
  NAND2_X1   g07620(.A1(new_n3654_), .A2(new_n7684_), .ZN(new_n7685_));
  XOR2_X1    g07621(.A1(new_n7685_), .A2(new_n72_), .Z(new_n7686_));
  INV_X1     g07622(.I(new_n7686_), .ZN(new_n7687_));
  XOR2_X1    g07623(.A1(new_n4535_), .A2(new_n74_), .Z(new_n7688_));
  NAND2_X1   g07624(.A1(new_n7688_), .A2(new_n4632_), .ZN(new_n7689_));
  INV_X1     g07625(.I(new_n4658_), .ZN(new_n7690_));
  AOI22_X1   g07626(.A1(new_n7689_), .A2(new_n4635_), .B1(new_n4657_), .B2(new_n7690_), .ZN(new_n7691_));
  XOR2_X1    g07627(.A1(new_n4641_), .A2(new_n4655_), .Z(new_n7692_));
  NOR2_X1    g07628(.A1(new_n4636_), .A2(new_n7692_), .ZN(new_n7693_));
  NOR2_X1    g07629(.A1(new_n7691_), .A2(new_n7693_), .ZN(new_n7694_));
  OAI22_X1   g07630(.A1(new_n1453_), .A2(new_n3175_), .B1(new_n2351_), .B2(new_n2742_), .ZN(new_n7695_));
  NAND2_X1   g07631(.A1(new_n2310_), .A2(new_n2746_), .ZN(new_n7696_));
  AOI21_X1   g07632(.A1(new_n7696_), .A2(new_n7695_), .B(new_n2737_), .ZN(new_n7697_));
  NAND2_X1   g07633(.A1(new_n4231_), .A2(new_n7697_), .ZN(new_n7698_));
  XOR2_X1    g07634(.A1(new_n7698_), .A2(\a[29] ), .Z(new_n7699_));
  NAND2_X1   g07635(.A1(new_n7694_), .A2(new_n7699_), .ZN(new_n7700_));
  OR2_X2     g07636(.A1(new_n7691_), .A2(new_n7693_), .Z(new_n7701_));
  INV_X1     g07637(.I(new_n7699_), .ZN(new_n7702_));
  NAND2_X1   g07638(.A1(new_n7701_), .A2(new_n7702_), .ZN(new_n7703_));
  AOI21_X1   g07639(.A1(new_n7703_), .A2(new_n7700_), .B(new_n7687_), .ZN(new_n7704_));
  NAND2_X1   g07640(.A1(new_n7701_), .A2(new_n7699_), .ZN(new_n7705_));
  NAND2_X1   g07641(.A1(new_n7694_), .A2(new_n7702_), .ZN(new_n7706_));
  AOI21_X1   g07642(.A1(new_n7705_), .A2(new_n7706_), .B(new_n7686_), .ZN(new_n7707_));
  OR2_X2     g07643(.A1(new_n7704_), .A2(new_n7707_), .Z(new_n7708_));
  NAND2_X1   g07644(.A1(new_n7570_), .A2(new_n7566_), .ZN(new_n7709_));
  NAND2_X1   g07645(.A1(new_n7709_), .A2(new_n7568_), .ZN(new_n7710_));
  NOR2_X1    g07646(.A1(new_n7708_), .A2(new_n7710_), .ZN(new_n7711_));
  NOR2_X1    g07647(.A1(new_n7704_), .A2(new_n7707_), .ZN(new_n7712_));
  INV_X1     g07648(.I(new_n7710_), .ZN(new_n7713_));
  NOR2_X1    g07649(.A1(new_n7712_), .A2(new_n7713_), .ZN(new_n7714_));
  OAI21_X1   g07650(.A1(new_n7711_), .A2(new_n7714_), .B(new_n7681_), .ZN(new_n7715_));
  XOR2_X1    g07651(.A1(new_n7680_), .A2(\a[23] ), .Z(new_n7716_));
  NOR2_X1    g07652(.A1(new_n7712_), .A2(new_n7710_), .ZN(new_n7717_));
  NOR2_X1    g07653(.A1(new_n7708_), .A2(new_n7713_), .ZN(new_n7718_));
  OAI21_X1   g07654(.A1(new_n7718_), .A2(new_n7717_), .B(new_n7716_), .ZN(new_n7719_));
  NAND2_X1   g07655(.A1(new_n7715_), .A2(new_n7719_), .ZN(new_n7720_));
  NAND2_X1   g07656(.A1(new_n7575_), .A2(new_n7579_), .ZN(new_n7721_));
  NAND2_X1   g07657(.A1(new_n7721_), .A2(new_n7577_), .ZN(new_n7722_));
  NOR2_X1    g07658(.A1(new_n7720_), .A2(new_n7722_), .ZN(new_n7723_));
  INV_X1     g07659(.I(new_n7722_), .ZN(new_n7724_));
  AOI21_X1   g07660(.A1(new_n7715_), .A2(new_n7719_), .B(new_n7724_), .ZN(new_n7725_));
  OAI21_X1   g07661(.A1(new_n7725_), .A2(new_n7723_), .B(new_n7676_), .ZN(new_n7726_));
  INV_X1     g07662(.I(new_n7676_), .ZN(new_n7727_));
  NAND2_X1   g07663(.A1(new_n7720_), .A2(new_n7724_), .ZN(new_n7728_));
  NAND3_X1   g07664(.A1(new_n7715_), .A2(new_n7719_), .A3(new_n7722_), .ZN(new_n7729_));
  NAND2_X1   g07665(.A1(new_n7728_), .A2(new_n7729_), .ZN(new_n7730_));
  NAND2_X1   g07666(.A1(new_n7730_), .A2(new_n7727_), .ZN(new_n7731_));
  NAND2_X1   g07667(.A1(new_n7731_), .A2(new_n7726_), .ZN(new_n7732_));
  AOI21_X1   g07668(.A1(new_n7550_), .A2(new_n7585_), .B(new_n7587_), .ZN(new_n7733_));
  INV_X1     g07669(.I(new_n7733_), .ZN(new_n7734_));
  NOR2_X1    g07670(.A1(new_n7732_), .A2(new_n7734_), .ZN(new_n7735_));
  INV_X1     g07671(.I(new_n7735_), .ZN(new_n7736_));
  NAND2_X1   g07672(.A1(new_n7732_), .A2(new_n7734_), .ZN(new_n7737_));
  AOI21_X1   g07673(.A1(new_n7736_), .A2(new_n7737_), .B(new_n7671_), .ZN(new_n7738_));
  INV_X1     g07674(.I(new_n7671_), .ZN(new_n7739_));
  NAND2_X1   g07675(.A1(new_n7732_), .A2(new_n7733_), .ZN(new_n7740_));
  NAND3_X1   g07676(.A1(new_n7734_), .A2(new_n7726_), .A3(new_n7731_), .ZN(new_n7741_));
  AOI21_X1   g07677(.A1(new_n7740_), .A2(new_n7741_), .B(new_n7739_), .ZN(new_n7742_));
  NAND2_X1   g07678(.A1(new_n7590_), .A2(new_n7598_), .ZN(new_n7743_));
  NAND2_X1   g07679(.A1(new_n7743_), .A2(new_n7600_), .ZN(new_n7744_));
  NOR3_X1    g07680(.A1(new_n7738_), .A2(new_n7744_), .A3(new_n7742_), .ZN(new_n7745_));
  INV_X1     g07681(.I(new_n7745_), .ZN(new_n7746_));
  OAI21_X1   g07682(.A1(new_n7738_), .A2(new_n7742_), .B(new_n7744_), .ZN(new_n7747_));
  AOI21_X1   g07683(.A1(new_n7746_), .A2(new_n7747_), .B(new_n7666_), .ZN(new_n7748_));
  XOR2_X1    g07684(.A1(new_n7665_), .A2(new_n3521_), .Z(new_n7749_));
  INV_X1     g07685(.I(new_n7737_), .ZN(new_n7750_));
  OAI21_X1   g07686(.A1(new_n7750_), .A2(new_n7735_), .B(new_n7739_), .ZN(new_n7751_));
  INV_X1     g07687(.I(new_n7742_), .ZN(new_n7752_));
  AOI21_X1   g07688(.A1(new_n7752_), .A2(new_n7751_), .B(new_n7744_), .ZN(new_n7753_));
  INV_X1     g07689(.I(new_n7753_), .ZN(new_n7754_));
  NAND3_X1   g07690(.A1(new_n7752_), .A2(new_n7751_), .A3(new_n7744_), .ZN(new_n7755_));
  AOI21_X1   g07691(.A1(new_n7754_), .A2(new_n7755_), .B(new_n7749_), .ZN(new_n7756_));
  NOR2_X1    g07692(.A1(new_n7756_), .A2(new_n7748_), .ZN(new_n7757_));
  OAI21_X1   g07693(.A1(new_n7545_), .A2(new_n7627_), .B(new_n7612_), .ZN(new_n7758_));
  INV_X1     g07694(.I(new_n7758_), .ZN(new_n7759_));
  NAND2_X1   g07695(.A1(new_n7757_), .A2(new_n7759_), .ZN(new_n7760_));
  INV_X1     g07696(.I(new_n7747_), .ZN(new_n7761_));
  OAI21_X1   g07697(.A1(new_n7761_), .A2(new_n7745_), .B(new_n7749_), .ZN(new_n7762_));
  INV_X1     g07698(.I(new_n7744_), .ZN(new_n7763_));
  NOR3_X1    g07699(.A1(new_n7763_), .A2(new_n7738_), .A3(new_n7742_), .ZN(new_n7764_));
  OAI21_X1   g07700(.A1(new_n7753_), .A2(new_n7764_), .B(new_n7666_), .ZN(new_n7765_));
  NAND2_X1   g07701(.A1(new_n7762_), .A2(new_n7765_), .ZN(new_n7766_));
  NAND2_X1   g07702(.A1(new_n7766_), .A2(new_n7758_), .ZN(new_n7767_));
  AOI21_X1   g07703(.A1(new_n7760_), .A2(new_n7767_), .B(new_n7661_), .ZN(new_n7768_));
  INV_X1     g07704(.I(new_n7661_), .ZN(new_n7769_));
  NAND2_X1   g07705(.A1(new_n7766_), .A2(new_n7759_), .ZN(new_n7770_));
  NAND2_X1   g07706(.A1(new_n7757_), .A2(new_n7758_), .ZN(new_n7771_));
  AOI21_X1   g07707(.A1(new_n7771_), .A2(new_n7770_), .B(new_n7769_), .ZN(new_n7772_));
  OAI21_X1   g07708(.A1(new_n7539_), .A2(new_n7620_), .B(new_n7622_), .ZN(new_n7773_));
  INV_X1     g07709(.I(new_n7773_), .ZN(new_n7774_));
  NOR3_X1    g07710(.A1(new_n7774_), .A2(new_n7768_), .A3(new_n7772_), .ZN(new_n7775_));
  NOR2_X1    g07711(.A1(new_n7766_), .A2(new_n7758_), .ZN(new_n7776_));
  NOR2_X1    g07712(.A1(new_n7757_), .A2(new_n7759_), .ZN(new_n7777_));
  OAI21_X1   g07713(.A1(new_n7777_), .A2(new_n7776_), .B(new_n7769_), .ZN(new_n7778_));
  INV_X1     g07714(.I(new_n7772_), .ZN(new_n7779_));
  AOI21_X1   g07715(.A1(new_n7779_), .A2(new_n7778_), .B(new_n7773_), .ZN(new_n7780_));
  OAI21_X1   g07716(.A1(new_n7780_), .A2(new_n7775_), .B(new_n4009_), .ZN(new_n7781_));
  NAND3_X1   g07717(.A1(new_n7779_), .A2(new_n7778_), .A3(new_n7773_), .ZN(new_n7782_));
  OAI21_X1   g07718(.A1(new_n7768_), .A2(new_n7772_), .B(new_n7774_), .ZN(new_n7783_));
  NAND3_X1   g07719(.A1(new_n7782_), .A2(new_n7783_), .A3(\a[8] ), .ZN(new_n7784_));
  AOI21_X1   g07720(.A1(new_n7781_), .A2(new_n7784_), .B(new_n7656_), .ZN(new_n7785_));
  INV_X1     g07721(.I(new_n7656_), .ZN(new_n7786_));
  AOI21_X1   g07722(.A1(new_n7782_), .A2(new_n7783_), .B(\a[8] ), .ZN(new_n7787_));
  NOR3_X1    g07723(.A1(new_n7780_), .A2(new_n4009_), .A3(new_n7775_), .ZN(new_n7788_));
  NOR3_X1    g07724(.A1(new_n7787_), .A2(new_n7788_), .A3(new_n7786_), .ZN(new_n7789_));
  NOR2_X1    g07725(.A1(new_n7789_), .A2(new_n7785_), .ZN(new_n7790_));
  INV_X1     g07726(.I(new_n7790_), .ZN(new_n7791_));
  OAI22_X1   g07727(.A1(new_n694_), .A2(new_n6089_), .B1(new_n2665_), .B2(new_n6091_), .ZN(new_n7792_));
  NAND2_X1   g07728(.A1(new_n2615_), .A2(new_n6095_), .ZN(new_n7793_));
  AOI21_X1   g07729(.A1(new_n7792_), .A2(new_n7793_), .B(new_n6082_), .ZN(new_n7794_));
  NAND2_X1   g07730(.A1(new_n3188_), .A2(new_n7794_), .ZN(new_n7795_));
  XOR2_X1    g07731(.A1(new_n7795_), .A2(\a[14] ), .Z(new_n7796_));
  INV_X1     g07732(.I(new_n7796_), .ZN(new_n7797_));
  OAI22_X1   g07733(.A1(new_n813_), .A2(new_n4291_), .B1(new_n529_), .B2(new_n4470_), .ZN(new_n7798_));
  NAND2_X1   g07734(.A1(new_n2563_), .A2(new_n4298_), .ZN(new_n7799_));
  AOI21_X1   g07735(.A1(new_n7799_), .A2(new_n7798_), .B(new_n4468_), .ZN(new_n7800_));
  NAND2_X1   g07736(.A1(new_n3051_), .A2(new_n7800_), .ZN(new_n7801_));
  XOR2_X1    g07737(.A1(new_n7801_), .A2(\a[17] ), .Z(new_n7802_));
  OAI22_X1   g07738(.A1(new_n896_), .A2(new_n4097_), .B1(new_n1180_), .B2(new_n3769_), .ZN(new_n7803_));
  NAND2_X1   g07739(.A1(new_n2504_), .A2(new_n3776_), .ZN(new_n7804_));
  AOI21_X1   g07740(.A1(new_n7804_), .A2(new_n7803_), .B(new_n4095_), .ZN(new_n7805_));
  NAND2_X1   g07741(.A1(new_n3596_), .A2(new_n7805_), .ZN(new_n7806_));
  XOR2_X1    g07742(.A1(new_n7806_), .A2(\a[20] ), .Z(new_n7807_));
  OAI22_X1   g07743(.A1(new_n1121_), .A2(new_n3780_), .B1(new_n2451_), .B2(new_n3310_), .ZN(new_n7808_));
  NAND2_X1   g07744(.A1(new_n2496_), .A2(new_n3782_), .ZN(new_n7809_));
  AOI21_X1   g07745(.A1(new_n7808_), .A2(new_n7809_), .B(new_n3302_), .ZN(new_n7810_));
  NAND2_X1   g07746(.A1(new_n3393_), .A2(new_n7810_), .ZN(new_n7811_));
  XOR2_X1    g07747(.A1(new_n7811_), .A2(\a[23] ), .Z(new_n7812_));
  OAI22_X1   g07748(.A1(new_n2367_), .A2(new_n3322_), .B1(new_n2408_), .B2(new_n3318_), .ZN(new_n7813_));
  NAND2_X1   g07749(.A1(new_n1334_), .A2(new_n3267_), .ZN(new_n7814_));
  AOI21_X1   g07750(.A1(new_n7813_), .A2(new_n7814_), .B(new_n3260_), .ZN(new_n7815_));
  NAND2_X1   g07751(.A1(new_n3708_), .A2(new_n7815_), .ZN(new_n7816_));
  XOR2_X1    g07752(.A1(new_n7816_), .A2(\a[26] ), .Z(new_n7817_));
  XNOR2_X1   g07753(.A1(new_n4659_), .A2(new_n4662_), .ZN(new_n7818_));
  NOR2_X1    g07754(.A1(new_n7818_), .A2(new_n4530_), .ZN(new_n7819_));
  AOI21_X1   g07755(.A1(new_n4665_), .A2(new_n4663_), .B(new_n4531_), .ZN(new_n7820_));
  NOR2_X1    g07756(.A1(new_n7819_), .A2(new_n7820_), .ZN(new_n7821_));
  NAND2_X1   g07757(.A1(new_n7700_), .A2(new_n7686_), .ZN(new_n7822_));
  NAND2_X1   g07758(.A1(new_n7822_), .A2(new_n7703_), .ZN(new_n7823_));
  INV_X1     g07759(.I(new_n7823_), .ZN(new_n7824_));
  NAND2_X1   g07760(.A1(new_n7824_), .A2(new_n7821_), .ZN(new_n7825_));
  INV_X1     g07761(.I(new_n7821_), .ZN(new_n7826_));
  NAND2_X1   g07762(.A1(new_n7826_), .A2(new_n7823_), .ZN(new_n7827_));
  AOI21_X1   g07763(.A1(new_n7827_), .A2(new_n7825_), .B(new_n7817_), .ZN(new_n7828_));
  INV_X1     g07764(.I(new_n7817_), .ZN(new_n7829_));
  NOR2_X1    g07765(.A1(new_n7821_), .A2(new_n7823_), .ZN(new_n7830_));
  NOR2_X1    g07766(.A1(new_n7826_), .A2(new_n7824_), .ZN(new_n7831_));
  NOR2_X1    g07767(.A1(new_n7831_), .A2(new_n7830_), .ZN(new_n7832_));
  NOR2_X1    g07768(.A1(new_n7832_), .A2(new_n7829_), .ZN(new_n7833_));
  NOR2_X1    g07769(.A1(new_n7833_), .A2(new_n7828_), .ZN(new_n7834_));
  NOR2_X1    g07770(.A1(new_n7711_), .A2(new_n7716_), .ZN(new_n7835_));
  NOR2_X1    g07771(.A1(new_n7835_), .A2(new_n7714_), .ZN(new_n7836_));
  NAND2_X1   g07772(.A1(new_n7834_), .A2(new_n7836_), .ZN(new_n7837_));
  INV_X1     g07773(.I(new_n7834_), .ZN(new_n7838_));
  INV_X1     g07774(.I(new_n7836_), .ZN(new_n7839_));
  NAND2_X1   g07775(.A1(new_n7838_), .A2(new_n7839_), .ZN(new_n7840_));
  AOI21_X1   g07776(.A1(new_n7840_), .A2(new_n7837_), .B(new_n7812_), .ZN(new_n7841_));
  INV_X1     g07777(.I(new_n7812_), .ZN(new_n7842_));
  NAND2_X1   g07778(.A1(new_n7838_), .A2(new_n7836_), .ZN(new_n7843_));
  NAND2_X1   g07779(.A1(new_n7839_), .A2(new_n7834_), .ZN(new_n7844_));
  AOI21_X1   g07780(.A1(new_n7843_), .A2(new_n7844_), .B(new_n7842_), .ZN(new_n7845_));
  NOR2_X1    g07781(.A1(new_n7841_), .A2(new_n7845_), .ZN(new_n7846_));
  INV_X1     g07782(.I(new_n7725_), .ZN(new_n7847_));
  OAI21_X1   g07783(.A1(new_n7720_), .A2(new_n7722_), .B(new_n7676_), .ZN(new_n7848_));
  NAND2_X1   g07784(.A1(new_n7848_), .A2(new_n7847_), .ZN(new_n7849_));
  INV_X1     g07785(.I(new_n7849_), .ZN(new_n7850_));
  NAND2_X1   g07786(.A1(new_n7846_), .A2(new_n7850_), .ZN(new_n7851_));
  OR2_X2     g07787(.A1(new_n7841_), .A2(new_n7845_), .Z(new_n7852_));
  NAND2_X1   g07788(.A1(new_n7852_), .A2(new_n7849_), .ZN(new_n7853_));
  AOI21_X1   g07789(.A1(new_n7853_), .A2(new_n7851_), .B(new_n7807_), .ZN(new_n7854_));
  INV_X1     g07790(.I(new_n7807_), .ZN(new_n7855_));
  NAND2_X1   g07791(.A1(new_n7852_), .A2(new_n7850_), .ZN(new_n7856_));
  NAND2_X1   g07792(.A1(new_n7846_), .A2(new_n7849_), .ZN(new_n7857_));
  AOI21_X1   g07793(.A1(new_n7856_), .A2(new_n7857_), .B(new_n7855_), .ZN(new_n7858_));
  OAI21_X1   g07794(.A1(new_n7671_), .A2(new_n7735_), .B(new_n7737_), .ZN(new_n7859_));
  NOR3_X1    g07795(.A1(new_n7854_), .A2(new_n7858_), .A3(new_n7859_), .ZN(new_n7860_));
  INV_X1     g07796(.I(new_n7860_), .ZN(new_n7861_));
  OAI21_X1   g07797(.A1(new_n7854_), .A2(new_n7858_), .B(new_n7859_), .ZN(new_n7862_));
  AOI21_X1   g07798(.A1(new_n7861_), .A2(new_n7862_), .B(new_n7802_), .ZN(new_n7863_));
  INV_X1     g07799(.I(new_n7802_), .ZN(new_n7864_));
  INV_X1     g07800(.I(new_n7859_), .ZN(new_n7865_));
  OAI21_X1   g07801(.A1(new_n7854_), .A2(new_n7858_), .B(new_n7865_), .ZN(new_n7866_));
  NOR3_X1    g07802(.A1(new_n7854_), .A2(new_n7858_), .A3(new_n7865_), .ZN(new_n7867_));
  INV_X1     g07803(.I(new_n7867_), .ZN(new_n7868_));
  AOI21_X1   g07804(.A1(new_n7868_), .A2(new_n7866_), .B(new_n7864_), .ZN(new_n7869_));
  NOR2_X1    g07805(.A1(new_n7869_), .A2(new_n7863_), .ZN(new_n7870_));
  AOI21_X1   g07806(.A1(new_n7749_), .A2(new_n7746_), .B(new_n7761_), .ZN(new_n7871_));
  INV_X1     g07807(.I(new_n7871_), .ZN(new_n7872_));
  NOR2_X1    g07808(.A1(new_n7870_), .A2(new_n7872_), .ZN(new_n7873_));
  INV_X1     g07809(.I(new_n7862_), .ZN(new_n7874_));
  OAI21_X1   g07810(.A1(new_n7874_), .A2(new_n7860_), .B(new_n7864_), .ZN(new_n7875_));
  INV_X1     g07811(.I(new_n7866_), .ZN(new_n7876_));
  OAI21_X1   g07812(.A1(new_n7876_), .A2(new_n7867_), .B(new_n7802_), .ZN(new_n7877_));
  NAND2_X1   g07813(.A1(new_n7877_), .A2(new_n7875_), .ZN(new_n7878_));
  NOR2_X1    g07814(.A1(new_n7878_), .A2(new_n7871_), .ZN(new_n7879_));
  OAI21_X1   g07815(.A1(new_n7873_), .A2(new_n7879_), .B(new_n7797_), .ZN(new_n7880_));
  NOR2_X1    g07816(.A1(new_n7878_), .A2(new_n7872_), .ZN(new_n7881_));
  NOR2_X1    g07817(.A1(new_n7870_), .A2(new_n7871_), .ZN(new_n7882_));
  OAI21_X1   g07818(.A1(new_n7882_), .A2(new_n7881_), .B(new_n7796_), .ZN(new_n7883_));
  AND2_X2    g07819(.A1(new_n7880_), .A2(new_n7883_), .Z(new_n7884_));
  NAND2_X1   g07820(.A1(new_n7760_), .A2(new_n7769_), .ZN(new_n7885_));
  NOR2_X1    g07821(.A1(new_n3142_), .A2(new_n4710_), .ZN(new_n7886_));
  NOR2_X1    g07822(.A1(new_n3176_), .A2(new_n4719_), .ZN(new_n7887_));
  OAI22_X1   g07823(.A1(new_n7887_), .A2(new_n7886_), .B1(new_n2716_), .B2(new_n4716_), .ZN(new_n7888_));
  AOI21_X1   g07824(.A1(new_n3174_), .A2(new_n4706_), .B(new_n7888_), .ZN(new_n7889_));
  INV_X1     g07825(.I(new_n7889_), .ZN(new_n7890_));
  NAND3_X1   g07826(.A1(new_n7885_), .A2(new_n7767_), .A3(new_n7890_), .ZN(new_n7891_));
  NOR2_X1    g07827(.A1(new_n7776_), .A2(new_n7661_), .ZN(new_n7892_));
  OAI21_X1   g07828(.A1(new_n7892_), .A2(new_n7777_), .B(new_n7889_), .ZN(new_n7893_));
  AOI21_X1   g07829(.A1(new_n7891_), .A2(new_n7893_), .B(\a[11] ), .ZN(new_n7894_));
  NOR3_X1    g07830(.A1(new_n7892_), .A2(new_n7777_), .A3(new_n7889_), .ZN(new_n7895_));
  AOI21_X1   g07831(.A1(new_n7769_), .A2(new_n7760_), .B(new_n7777_), .ZN(new_n7896_));
  NOR2_X1    g07832(.A1(new_n7896_), .A2(new_n7890_), .ZN(new_n7897_));
  NOR3_X1    g07833(.A1(new_n7897_), .A2(new_n7895_), .A3(new_n4034_), .ZN(new_n7898_));
  OAI21_X1   g07834(.A1(new_n7898_), .A2(new_n7894_), .B(new_n7884_), .ZN(new_n7899_));
  NAND2_X1   g07835(.A1(new_n7880_), .A2(new_n7883_), .ZN(new_n7900_));
  OAI21_X1   g07836(.A1(new_n7897_), .A2(new_n7895_), .B(new_n4034_), .ZN(new_n7901_));
  NAND3_X1   g07837(.A1(new_n7891_), .A2(new_n7893_), .A3(\a[11] ), .ZN(new_n7902_));
  NAND3_X1   g07838(.A1(new_n7901_), .A2(new_n7902_), .A3(new_n7900_), .ZN(new_n7903_));
  AOI21_X1   g07839(.A1(new_n7779_), .A2(new_n7778_), .B(new_n7774_), .ZN(new_n7904_));
  XOR2_X1    g07840(.A1(new_n7656_), .A2(new_n4009_), .Z(new_n7905_));
  NOR4_X1    g07841(.A1(new_n7768_), .A2(new_n7772_), .A3(new_n7773_), .A4(new_n7905_), .ZN(new_n7906_));
  NOR2_X1    g07842(.A1(new_n7904_), .A2(new_n7906_), .ZN(new_n7907_));
  INV_X1     g07843(.I(new_n7907_), .ZN(new_n7908_));
  NAND3_X1   g07844(.A1(new_n7899_), .A2(new_n7908_), .A3(new_n7903_), .ZN(new_n7909_));
  AOI21_X1   g07845(.A1(new_n7901_), .A2(new_n7902_), .B(new_n7900_), .ZN(new_n7910_));
  NOR3_X1    g07846(.A1(new_n7898_), .A2(new_n7884_), .A3(new_n7894_), .ZN(new_n7911_));
  OAI21_X1   g07847(.A1(new_n7911_), .A2(new_n7910_), .B(new_n7907_), .ZN(new_n7912_));
  AOI21_X1   g07848(.A1(new_n7636_), .A2(new_n7639_), .B(new_n7633_), .ZN(new_n7913_));
  AOI21_X1   g07849(.A1(new_n7643_), .A2(new_n7644_), .B(new_n7913_), .ZN(new_n7914_));
  INV_X1     g07850(.I(new_n7914_), .ZN(new_n7915_));
  NAND3_X1   g07851(.A1(new_n7909_), .A2(new_n7912_), .A3(new_n7915_), .ZN(new_n7916_));
  NAND3_X1   g07852(.A1(new_n7655_), .A2(new_n7791_), .A3(new_n7916_), .ZN(new_n7917_));
  NOR3_X1    g07853(.A1(new_n7908_), .A2(new_n7911_), .A3(new_n7910_), .ZN(new_n7918_));
  INV_X1     g07854(.I(new_n7918_), .ZN(new_n7919_));
  NAND2_X1   g07855(.A1(new_n7917_), .A2(new_n7919_), .ZN(new_n7920_));
  NOR2_X1    g07856(.A1(new_n6946_), .A2(new_n6949_), .ZN(new_n7921_));
  NAND4_X1   g07857(.A1(new_n6928_), .A2(new_n6938_), .A3(new_n7135_), .A4(new_n7138_), .ZN(new_n7922_));
  OAI21_X1   g07858(.A1(new_n6946_), .A2(new_n6949_), .B(new_n7139_), .ZN(new_n7923_));
  AOI22_X1   g07859(.A1(new_n7922_), .A2(new_n7923_), .B1(new_n7921_), .B2(new_n6948_), .ZN(new_n7924_));
  OAI21_X1   g07860(.A1(new_n7371_), .A2(new_n7370_), .B(new_n7369_), .ZN(new_n7925_));
  NAND3_X1   g07861(.A1(new_n7364_), .A2(new_n7367_), .A3(new_n7143_), .ZN(new_n7926_));
  NAND3_X1   g07862(.A1(new_n7925_), .A2(new_n7926_), .A3(new_n7374_), .ZN(new_n7927_));
  AOI21_X1   g07863(.A1(new_n7925_), .A2(new_n7926_), .B(new_n7374_), .ZN(new_n7928_));
  AOI21_X1   g07864(.A1(new_n7924_), .A2(new_n7927_), .B(new_n7928_), .ZN(new_n7929_));
  OAI21_X1   g07865(.A1(new_n7520_), .A2(new_n7512_), .B(new_n7519_), .ZN(new_n7930_));
  NAND3_X1   g07866(.A1(new_n7513_), .A2(new_n7503_), .A3(new_n7511_), .ZN(new_n7931_));
  INV_X1     g07867(.I(new_n7526_), .ZN(new_n7932_));
  AOI21_X1   g07868(.A1(new_n7930_), .A2(new_n7931_), .B(new_n7932_), .ZN(new_n7933_));
  NAND3_X1   g07869(.A1(new_n7930_), .A2(new_n7932_), .A3(new_n7931_), .ZN(new_n7934_));
  OAI21_X1   g07870(.A1(new_n7929_), .A2(new_n7933_), .B(new_n7934_), .ZN(new_n7935_));
  AOI21_X1   g07871(.A1(new_n7636_), .A2(new_n7639_), .B(new_n7640_), .ZN(new_n7936_));
  NOR3_X1    g07872(.A1(new_n7623_), .A2(new_n7632_), .A3(new_n7633_), .ZN(new_n7937_));
  OAI21_X1   g07873(.A1(new_n7936_), .A2(new_n7937_), .B(new_n7643_), .ZN(new_n7938_));
  NOR3_X1    g07874(.A1(new_n7640_), .A2(new_n7623_), .A3(new_n7632_), .ZN(new_n7939_));
  OAI21_X1   g07875(.A1(new_n7939_), .A2(new_n7913_), .B(new_n7534_), .ZN(new_n7940_));
  NAND2_X1   g07876(.A1(new_n7938_), .A2(new_n7940_), .ZN(new_n7941_));
  INV_X1     g07877(.I(new_n7504_), .ZN(new_n7942_));
  NOR2_X1    g07878(.A1(new_n7503_), .A2(new_n7648_), .ZN(new_n7943_));
  NOR2_X1    g07879(.A1(new_n7519_), .A2(new_n7649_), .ZN(new_n7944_));
  OAI22_X1   g07880(.A1(new_n7944_), .A2(new_n7943_), .B1(new_n7942_), .B2(new_n7648_), .ZN(new_n7945_));
  NAND2_X1   g07881(.A1(new_n7941_), .A2(new_n7945_), .ZN(new_n7946_));
  NOR2_X1    g07882(.A1(new_n7941_), .A2(new_n7945_), .ZN(new_n7947_));
  AOI21_X1   g07883(.A1(new_n7935_), .A2(new_n7946_), .B(new_n7947_), .ZN(new_n7948_));
  NOR3_X1    g07884(.A1(new_n7911_), .A2(new_n7910_), .A3(new_n7907_), .ZN(new_n7949_));
  AOI21_X1   g07885(.A1(new_n7899_), .A2(new_n7903_), .B(new_n7908_), .ZN(new_n7950_));
  NOR3_X1    g07886(.A1(new_n7950_), .A2(new_n7949_), .A3(new_n7914_), .ZN(new_n7951_));
  NOR3_X1    g07887(.A1(new_n7948_), .A2(new_n7951_), .A3(new_n7790_), .ZN(new_n7952_));
  NAND2_X1   g07888(.A1(new_n3168_), .A2(new_n6480_), .ZN(new_n7953_));
  NAND2_X1   g07889(.A1(new_n3247_), .A2(new_n4720_), .ZN(new_n7954_));
  NAND4_X1   g07890(.A1(new_n3758_), .A2(new_n4706_), .A3(new_n7953_), .A4(new_n7954_), .ZN(new_n7955_));
  XOR2_X1    g07891(.A1(new_n7955_), .A2(\a[11] ), .Z(new_n7956_));
  INV_X1     g07892(.I(new_n7956_), .ZN(new_n7957_));
  OAI22_X1   g07893(.A1(new_n2614_), .A2(new_n6089_), .B1(new_n2665_), .B2(new_n6094_), .ZN(new_n7958_));
  NAND2_X1   g07894(.A1(new_n2728_), .A2(new_n6090_), .ZN(new_n7959_));
  AOI21_X1   g07895(.A1(new_n7959_), .A2(new_n7958_), .B(new_n6082_), .ZN(new_n7960_));
  NAND2_X1   g07896(.A1(new_n2733_), .A2(new_n7960_), .ZN(new_n7961_));
  XOR2_X1    g07897(.A1(new_n7961_), .A2(\a[14] ), .Z(new_n7962_));
  INV_X1     g07898(.I(new_n7962_), .ZN(new_n7963_));
  OAI22_X1   g07899(.A1(new_n2559_), .A2(new_n4291_), .B1(new_n694_), .B2(new_n4470_), .ZN(new_n7964_));
  NAND2_X1   g07900(.A1(new_n2567_), .A2(new_n4298_), .ZN(new_n7965_));
  AOI21_X1   g07901(.A1(new_n7964_), .A2(new_n7965_), .B(new_n4468_), .ZN(new_n7966_));
  NAND2_X1   g07902(.A1(new_n2759_), .A2(new_n7966_), .ZN(new_n7967_));
  XOR2_X1    g07903(.A1(new_n7967_), .A2(\a[17] ), .Z(new_n7968_));
  INV_X1     g07904(.I(new_n7968_), .ZN(new_n7969_));
  OAI22_X1   g07905(.A1(new_n1180_), .A2(new_n3780_), .B1(new_n2492_), .B2(new_n3310_), .ZN(new_n7970_));
  NAND2_X1   g07906(.A1(new_n1122_), .A2(new_n3782_), .ZN(new_n7971_));
  AOI21_X1   g07907(.A1(new_n7971_), .A2(new_n7970_), .B(new_n3302_), .ZN(new_n7972_));
  NAND2_X1   g07908(.A1(new_n3330_), .A2(new_n7972_), .ZN(new_n7973_));
  XOR2_X1    g07909(.A1(new_n7973_), .A2(\a[23] ), .Z(new_n7974_));
  INV_X1     g07910(.I(new_n7974_), .ZN(new_n7975_));
  OAI21_X1   g07911(.A1(new_n4669_), .A2(new_n4667_), .B(new_n4519_), .ZN(new_n7976_));
  XOR2_X1    g07912(.A1(new_n4525_), .A2(new_n4666_), .Z(new_n7977_));
  NAND2_X1   g07913(.A1(new_n7977_), .A2(new_n4520_), .ZN(new_n7978_));
  NOR2_X1    g07914(.A1(new_n7830_), .A2(new_n7817_), .ZN(new_n7979_));
  NOR2_X1    g07915(.A1(new_n7979_), .A2(new_n7831_), .ZN(new_n7980_));
  NAND3_X1   g07916(.A1(new_n7980_), .A2(new_n7978_), .A3(new_n7976_), .ZN(new_n7981_));
  NAND2_X1   g07917(.A1(new_n7978_), .A2(new_n7976_), .ZN(new_n7982_));
  OAI21_X1   g07918(.A1(new_n7831_), .A2(new_n7979_), .B(new_n7982_), .ZN(new_n7983_));
  NAND2_X1   g07919(.A1(new_n7983_), .A2(new_n7981_), .ZN(new_n7984_));
  NAND2_X1   g07920(.A1(new_n7984_), .A2(new_n7975_), .ZN(new_n7985_));
  XNOR2_X1   g07921(.A1(new_n7982_), .A2(new_n7980_), .ZN(new_n7986_));
  NAND2_X1   g07922(.A1(new_n7986_), .A2(new_n7974_), .ZN(new_n7987_));
  OAI22_X1   g07923(.A1(new_n813_), .A2(new_n4097_), .B1(new_n1008_), .B2(new_n3769_), .ZN(new_n7988_));
  NAND2_X1   g07924(.A1(new_n897_), .A2(new_n3776_), .ZN(new_n7989_));
  AOI21_X1   g07925(.A1(new_n7988_), .A2(new_n7989_), .B(new_n4095_), .ZN(new_n7990_));
  NAND2_X1   g07926(.A1(new_n2917_), .A2(new_n7990_), .ZN(new_n7991_));
  XOR2_X1    g07927(.A1(new_n7991_), .A2(new_n3035_), .Z(new_n7992_));
  INV_X1     g07928(.I(new_n7992_), .ZN(new_n7993_));
  INV_X1     g07929(.I(new_n7844_), .ZN(new_n7994_));
  AOI21_X1   g07930(.A1(new_n7842_), .A2(new_n7843_), .B(new_n7994_), .ZN(new_n7995_));
  NAND2_X1   g07931(.A1(new_n7993_), .A2(new_n7995_), .ZN(new_n7996_));
  INV_X1     g07932(.I(new_n7995_), .ZN(new_n7997_));
  NAND2_X1   g07933(.A1(new_n7997_), .A2(new_n7992_), .ZN(new_n7998_));
  AOI22_X1   g07934(.A1(new_n7998_), .A2(new_n7996_), .B1(new_n7985_), .B2(new_n7987_), .ZN(new_n7999_));
  NAND2_X1   g07935(.A1(new_n7987_), .A2(new_n7985_), .ZN(new_n8000_));
  XOR2_X1    g07936(.A1(new_n7995_), .A2(new_n7992_), .Z(new_n8001_));
  NOR2_X1    g07937(.A1(new_n8001_), .A2(new_n8000_), .ZN(new_n8002_));
  NOR2_X1    g07938(.A1(new_n8002_), .A2(new_n7999_), .ZN(new_n8003_));
  INV_X1     g07939(.I(new_n8003_), .ZN(new_n8004_));
  NAND2_X1   g07940(.A1(new_n7856_), .A2(new_n7855_), .ZN(new_n8005_));
  NAND2_X1   g07941(.A1(new_n8005_), .A2(new_n7857_), .ZN(new_n8006_));
  NOR2_X1    g07942(.A1(new_n8004_), .A2(new_n8006_), .ZN(new_n8007_));
  INV_X1     g07943(.I(new_n8006_), .ZN(new_n8008_));
  NOR2_X1    g07944(.A1(new_n8008_), .A2(new_n8003_), .ZN(new_n8009_));
  OAI21_X1   g07945(.A1(new_n8007_), .A2(new_n8009_), .B(new_n7969_), .ZN(new_n8010_));
  XOR2_X1    g07946(.A1(new_n8003_), .A2(new_n8006_), .Z(new_n8011_));
  OAI21_X1   g07947(.A1(new_n7969_), .A2(new_n8011_), .B(new_n8010_), .ZN(new_n8012_));
  AOI21_X1   g07948(.A1(new_n7864_), .A2(new_n7866_), .B(new_n7867_), .ZN(new_n8013_));
  INV_X1     g07949(.I(new_n8013_), .ZN(new_n8014_));
  NOR2_X1    g07950(.A1(new_n8012_), .A2(new_n8014_), .ZN(new_n8015_));
  OR2_X2     g07951(.A1(new_n8011_), .A2(new_n7969_), .Z(new_n8016_));
  AOI21_X1   g07952(.A1(new_n8016_), .A2(new_n8010_), .B(new_n8013_), .ZN(new_n8017_));
  OAI21_X1   g07953(.A1(new_n8017_), .A2(new_n8015_), .B(new_n7963_), .ZN(new_n8018_));
  XOR2_X1    g07954(.A1(new_n8012_), .A2(new_n8013_), .Z(new_n8019_));
  OAI21_X1   g07955(.A1(new_n8019_), .A2(new_n7963_), .B(new_n8018_), .ZN(new_n8020_));
  INV_X1     g07956(.I(new_n7879_), .ZN(new_n8021_));
  OAI21_X1   g07957(.A1(new_n7870_), .A2(new_n7872_), .B(new_n7797_), .ZN(new_n8022_));
  NAND2_X1   g07958(.A1(new_n8021_), .A2(new_n8022_), .ZN(new_n8023_));
  XOR2_X1    g07959(.A1(new_n8020_), .A2(new_n8023_), .Z(new_n8024_));
  NOR2_X1    g07960(.A1(new_n8020_), .A2(new_n8023_), .ZN(new_n8025_));
  INV_X1     g07961(.I(new_n8025_), .ZN(new_n8026_));
  NAND2_X1   g07962(.A1(new_n8020_), .A2(new_n8023_), .ZN(new_n8027_));
  AOI21_X1   g07963(.A1(new_n8026_), .A2(new_n8027_), .B(new_n7957_), .ZN(new_n8028_));
  AOI21_X1   g07964(.A1(new_n8024_), .A2(new_n7957_), .B(new_n8028_), .ZN(new_n8029_));
  OAI21_X1   g07965(.A1(new_n7952_), .A2(new_n7918_), .B(new_n8029_), .ZN(new_n8030_));
  NAND2_X1   g07966(.A1(new_n8024_), .A2(new_n7957_), .ZN(new_n8031_));
  INV_X1     g07967(.I(new_n8027_), .ZN(new_n8032_));
  OAI21_X1   g07968(.A1(new_n8032_), .A2(new_n8025_), .B(new_n7956_), .ZN(new_n8033_));
  NAND2_X1   g07969(.A1(new_n8031_), .A2(new_n8033_), .ZN(new_n8034_));
  NAND3_X1   g07970(.A1(new_n7917_), .A2(new_n7919_), .A3(new_n8034_), .ZN(new_n8035_));
  NOR2_X1    g07971(.A1(new_n7884_), .A2(new_n7896_), .ZN(new_n8036_));
  XOR2_X1    g07972(.A1(new_n7889_), .A2(\a[11] ), .Z(new_n8037_));
  NOR4_X1    g07973(.A1(new_n7900_), .A2(new_n7777_), .A3(new_n7892_), .A4(new_n8037_), .ZN(new_n8038_));
  NOR2_X1    g07974(.A1(new_n8036_), .A2(new_n8038_), .ZN(new_n8039_));
  INV_X1     g07975(.I(new_n8039_), .ZN(new_n8040_));
  AOI22_X1   g07976(.A1(new_n8030_), .A2(new_n8035_), .B1(new_n7920_), .B2(new_n8040_), .ZN(new_n8041_));
  AOI22_X1   g07977(.A1(new_n3253_), .A2(new_n4706_), .B1(new_n3247_), .B2(new_n6480_), .ZN(new_n8042_));
  INV_X1     g07978(.I(new_n8042_), .ZN(new_n8043_));
  OAI22_X1   g07979(.A1(new_n3176_), .A2(new_n6091_), .B1(new_n2665_), .B2(new_n6089_), .ZN(new_n8044_));
  NAND2_X1   g07980(.A1(new_n2728_), .A2(new_n6095_), .ZN(new_n8045_));
  AOI21_X1   g07981(.A1(new_n8044_), .A2(new_n8045_), .B(new_n6082_), .ZN(new_n8046_));
  NAND2_X1   g07982(.A1(new_n3273_), .A2(new_n8046_), .ZN(new_n8047_));
  XOR2_X1    g07983(.A1(new_n8047_), .A2(\a[14] ), .Z(new_n8048_));
  OAI22_X1   g07984(.A1(new_n2614_), .A2(new_n4470_), .B1(new_n529_), .B2(new_n4291_), .ZN(new_n8049_));
  NAND2_X1   g07985(.A1(new_n2718_), .A2(new_n4298_), .ZN(new_n8050_));
  AOI21_X1   g07986(.A1(new_n8050_), .A2(new_n8049_), .B(new_n4468_), .ZN(new_n8051_));
  NAND2_X1   g07987(.A1(new_n3074_), .A2(new_n8051_), .ZN(new_n8052_));
  XOR2_X1    g07988(.A1(new_n8052_), .A2(new_n3372_), .Z(new_n8053_));
  INV_X1     g07989(.I(new_n8053_), .ZN(new_n8054_));
  OAI22_X1   g07990(.A1(new_n2559_), .A2(new_n4097_), .B1(new_n896_), .B2(new_n3769_), .ZN(new_n8055_));
  NAND2_X1   g07991(.A1(new_n814_), .A2(new_n3776_), .ZN(new_n8056_));
  AOI21_X1   g07992(.A1(new_n8055_), .A2(new_n8056_), .B(new_n4095_), .ZN(new_n8057_));
  NAND2_X1   g07993(.A1(new_n3624_), .A2(new_n8057_), .ZN(new_n8058_));
  XOR2_X1    g07994(.A1(new_n8058_), .A2(\a[20] ), .Z(new_n8059_));
  INV_X1     g07995(.I(new_n4672_), .ZN(new_n8060_));
  AOI21_X1   g07996(.A1(new_n8060_), .A2(new_n4671_), .B(new_n4508_), .ZN(new_n8061_));
  INV_X1     g07997(.I(new_n4670_), .ZN(new_n8062_));
  XOR2_X1    g07998(.A1(new_n4514_), .A2(new_n8062_), .Z(new_n8063_));
  NOR2_X1    g07999(.A1(new_n8063_), .A2(new_n4509_), .ZN(new_n8064_));
  NOR2_X1    g08000(.A1(new_n8064_), .A2(new_n8061_), .ZN(new_n8065_));
  NAND2_X1   g08001(.A1(new_n7975_), .A2(new_n7981_), .ZN(new_n8066_));
  NAND2_X1   g08002(.A1(new_n8066_), .A2(new_n7983_), .ZN(new_n8067_));
  INV_X1     g08003(.I(new_n8067_), .ZN(new_n8068_));
  NAND2_X1   g08004(.A1(new_n8065_), .A2(new_n8068_), .ZN(new_n8069_));
  NOR2_X1    g08005(.A1(new_n8065_), .A2(new_n8068_), .ZN(new_n8070_));
  INV_X1     g08006(.I(new_n8070_), .ZN(new_n8071_));
  AOI21_X1   g08007(.A1(new_n8071_), .A2(new_n8069_), .B(new_n8059_), .ZN(new_n8072_));
  INV_X1     g08008(.I(new_n8059_), .ZN(new_n8073_));
  XOR2_X1    g08009(.A1(new_n8065_), .A2(new_n8067_), .Z(new_n8074_));
  NOR2_X1    g08010(.A1(new_n8074_), .A2(new_n8073_), .ZN(new_n8075_));
  NOR2_X1    g08011(.A1(new_n8075_), .A2(new_n8072_), .ZN(new_n8076_));
  NAND2_X1   g08012(.A1(new_n7996_), .A2(new_n8000_), .ZN(new_n8077_));
  NAND2_X1   g08013(.A1(new_n8077_), .A2(new_n7998_), .ZN(new_n8078_));
  INV_X1     g08014(.I(new_n8078_), .ZN(new_n8079_));
  NAND2_X1   g08015(.A1(new_n8076_), .A2(new_n8079_), .ZN(new_n8080_));
  OAI21_X1   g08016(.A1(new_n8075_), .A2(new_n8072_), .B(new_n8078_), .ZN(new_n8081_));
  AOI21_X1   g08017(.A1(new_n8080_), .A2(new_n8081_), .B(new_n8054_), .ZN(new_n8082_));
  XOR2_X1    g08018(.A1(new_n8076_), .A2(new_n8078_), .Z(new_n8083_));
  NOR2_X1    g08019(.A1(new_n8083_), .A2(new_n8053_), .ZN(new_n8084_));
  NOR2_X1    g08020(.A1(new_n8084_), .A2(new_n8082_), .ZN(new_n8085_));
  NAND2_X1   g08021(.A1(new_n8008_), .A2(new_n8003_), .ZN(new_n8086_));
  AOI21_X1   g08022(.A1(new_n7969_), .A2(new_n8086_), .B(new_n8009_), .ZN(new_n8087_));
  NAND2_X1   g08023(.A1(new_n8085_), .A2(new_n8087_), .ZN(new_n8088_));
  NOR2_X1    g08024(.A1(new_n8085_), .A2(new_n8087_), .ZN(new_n8089_));
  INV_X1     g08025(.I(new_n8089_), .ZN(new_n8090_));
  AOI21_X1   g08026(.A1(new_n8090_), .A2(new_n8088_), .B(new_n8048_), .ZN(new_n8091_));
  INV_X1     g08027(.I(new_n8048_), .ZN(new_n8092_));
  INV_X1     g08028(.I(new_n8087_), .ZN(new_n8093_));
  XOR2_X1    g08029(.A1(new_n8085_), .A2(new_n8093_), .Z(new_n8094_));
  NOR2_X1    g08030(.A1(new_n8094_), .A2(new_n8092_), .ZN(new_n8095_));
  INV_X1     g08031(.I(new_n8015_), .ZN(new_n8096_));
  AOI21_X1   g08032(.A1(new_n8096_), .A2(new_n7963_), .B(new_n8017_), .ZN(new_n8097_));
  NOR3_X1    g08033(.A1(new_n8095_), .A2(new_n8091_), .A3(new_n8097_), .ZN(new_n8098_));
  OAI21_X1   g08034(.A1(new_n8095_), .A2(new_n8091_), .B(new_n8097_), .ZN(new_n8099_));
  INV_X1     g08035(.I(new_n8099_), .ZN(new_n8100_));
  OAI21_X1   g08036(.A1(new_n8100_), .A2(new_n8098_), .B(new_n4034_), .ZN(new_n8101_));
  INV_X1     g08037(.I(new_n8098_), .ZN(new_n8102_));
  NAND3_X1   g08038(.A1(new_n8102_), .A2(new_n8099_), .A3(\a[11] ), .ZN(new_n8103_));
  AOI21_X1   g08039(.A1(new_n8101_), .A2(new_n8103_), .B(new_n8043_), .ZN(new_n8104_));
  AOI21_X1   g08040(.A1(new_n8102_), .A2(new_n8099_), .B(\a[11] ), .ZN(new_n8105_));
  NOR3_X1    g08041(.A1(new_n8100_), .A2(new_n8098_), .A3(new_n4034_), .ZN(new_n8106_));
  NOR3_X1    g08042(.A1(new_n8105_), .A2(new_n8106_), .A3(new_n8042_), .ZN(new_n8107_));
  NOR2_X1    g08043(.A1(new_n8107_), .A2(new_n8104_), .ZN(new_n8108_));
  INV_X1     g08044(.I(new_n8108_), .ZN(new_n8109_));
  NOR2_X1    g08045(.A1(new_n8095_), .A2(new_n8091_), .ZN(new_n8110_));
  NOR2_X1    g08046(.A1(new_n8110_), .A2(new_n8097_), .ZN(new_n8111_));
  INV_X1     g08047(.I(new_n8097_), .ZN(new_n8112_));
  XOR2_X1    g08048(.A1(new_n8042_), .A2(\a[11] ), .Z(new_n8113_));
  NOR4_X1    g08049(.A1(new_n8095_), .A2(new_n8091_), .A3(new_n8112_), .A4(new_n8113_), .ZN(new_n8114_));
  NOR2_X1    g08050(.A1(new_n8111_), .A2(new_n8114_), .ZN(new_n8115_));
  AOI21_X1   g08051(.A1(new_n8092_), .A2(new_n8088_), .B(new_n8089_), .ZN(new_n8116_));
  INV_X1     g08052(.I(new_n8116_), .ZN(new_n8117_));
  OAI22_X1   g08053(.A1(new_n3176_), .A2(new_n6094_), .B1(new_n3142_), .B2(new_n6091_), .ZN(new_n8118_));
  NAND2_X1   g08054(.A1(new_n2728_), .A2(new_n6180_), .ZN(new_n8119_));
  AOI21_X1   g08055(.A1(new_n8118_), .A2(new_n8119_), .B(new_n6082_), .ZN(new_n8120_));
  NAND2_X1   g08056(.A1(new_n3174_), .A2(new_n8120_), .ZN(new_n8121_));
  XOR2_X1    g08057(.A1(new_n8121_), .A2(\a[14] ), .Z(new_n8122_));
  INV_X1     g08058(.I(new_n8122_), .ZN(new_n8123_));
  OAI22_X1   g08059(.A1(new_n694_), .A2(new_n4291_), .B1(new_n2665_), .B2(new_n4470_), .ZN(new_n8124_));
  NAND2_X1   g08060(.A1(new_n2615_), .A2(new_n4298_), .ZN(new_n8125_));
  AOI21_X1   g08061(.A1(new_n8124_), .A2(new_n8125_), .B(new_n4468_), .ZN(new_n8126_));
  NAND2_X1   g08062(.A1(new_n3188_), .A2(new_n8126_), .ZN(new_n8127_));
  XOR2_X1    g08063(.A1(new_n8127_), .A2(\a[17] ), .Z(new_n8128_));
  OAI22_X1   g08064(.A1(new_n813_), .A2(new_n3769_), .B1(new_n529_), .B2(new_n4097_), .ZN(new_n8129_));
  NAND2_X1   g08065(.A1(new_n2563_), .A2(new_n3776_), .ZN(new_n8130_));
  AOI21_X1   g08066(.A1(new_n8130_), .A2(new_n8129_), .B(new_n4095_), .ZN(new_n8131_));
  NAND2_X1   g08067(.A1(new_n3051_), .A2(new_n8131_), .ZN(new_n8132_));
  XOR2_X1    g08068(.A1(new_n8132_), .A2(\a[20] ), .Z(new_n8133_));
  INV_X1     g08069(.I(new_n8133_), .ZN(new_n8134_));
  XNOR2_X1   g08070(.A1(new_n4503_), .A2(new_n4673_), .ZN(new_n8135_));
  NOR2_X1    g08071(.A1(new_n8135_), .A2(new_n4496_), .ZN(new_n8136_));
  INV_X1     g08072(.I(new_n4675_), .ZN(new_n8137_));
  AOI21_X1   g08073(.A1(new_n8137_), .A2(new_n4674_), .B(new_n4497_), .ZN(new_n8138_));
  NOR2_X1    g08074(.A1(new_n8136_), .A2(new_n8138_), .ZN(new_n8139_));
  AOI21_X1   g08075(.A1(new_n8065_), .A2(new_n8068_), .B(new_n8059_), .ZN(new_n8140_));
  NOR2_X1    g08076(.A1(new_n8140_), .A2(new_n8070_), .ZN(new_n8141_));
  INV_X1     g08077(.I(new_n8141_), .ZN(new_n8142_));
  XOR2_X1    g08078(.A1(new_n8139_), .A2(new_n8142_), .Z(new_n8143_));
  NAND2_X1   g08079(.A1(new_n8143_), .A2(new_n8134_), .ZN(new_n8144_));
  NOR2_X1    g08080(.A1(new_n8139_), .A2(new_n8142_), .ZN(new_n8145_));
  NOR3_X1    g08081(.A1(new_n8136_), .A2(new_n8138_), .A3(new_n8141_), .ZN(new_n8146_));
  OAI21_X1   g08082(.A1(new_n8145_), .A2(new_n8146_), .B(new_n8133_), .ZN(new_n8147_));
  NAND2_X1   g08083(.A1(new_n8144_), .A2(new_n8147_), .ZN(new_n8148_));
  INV_X1     g08084(.I(new_n8081_), .ZN(new_n8149_));
  AOI21_X1   g08085(.A1(new_n8076_), .A2(new_n8079_), .B(new_n8054_), .ZN(new_n8150_));
  NOR2_X1    g08086(.A1(new_n8150_), .A2(new_n8149_), .ZN(new_n8151_));
  INV_X1     g08087(.I(new_n8151_), .ZN(new_n8152_));
  XOR2_X1    g08088(.A1(new_n8148_), .A2(new_n8152_), .Z(new_n8153_));
  NAND2_X1   g08089(.A1(new_n8148_), .A2(new_n8151_), .ZN(new_n8154_));
  NAND3_X1   g08090(.A1(new_n8152_), .A2(new_n8144_), .A3(new_n8147_), .ZN(new_n8155_));
  NAND2_X1   g08091(.A1(new_n8154_), .A2(new_n8155_), .ZN(new_n8156_));
  NAND2_X1   g08092(.A1(new_n8156_), .A2(new_n8128_), .ZN(new_n8157_));
  OAI21_X1   g08093(.A1(new_n8128_), .A2(new_n8153_), .B(new_n8157_), .ZN(new_n8158_));
  NOR2_X1    g08094(.A1(new_n8158_), .A2(new_n8123_), .ZN(new_n8159_));
  NAND2_X1   g08095(.A1(new_n8158_), .A2(new_n8123_), .ZN(new_n8160_));
  INV_X1     g08096(.I(new_n8160_), .ZN(new_n8161_));
  OAI21_X1   g08097(.A1(new_n8161_), .A2(new_n8159_), .B(new_n8117_), .ZN(new_n8162_));
  NOR2_X1    g08098(.A1(new_n8158_), .A2(new_n8122_), .ZN(new_n8163_));
  NAND2_X1   g08099(.A1(new_n8158_), .A2(new_n8122_), .ZN(new_n8164_));
  INV_X1     g08100(.I(new_n8164_), .ZN(new_n8165_));
  OAI21_X1   g08101(.A1(new_n8165_), .A2(new_n8163_), .B(new_n8116_), .ZN(new_n8166_));
  NAND3_X1   g08102(.A1(new_n8162_), .A2(new_n8166_), .A3(new_n8115_), .ZN(new_n8167_));
  OR2_X2     g08103(.A1(new_n8111_), .A2(new_n8114_), .Z(new_n8168_));
  INV_X1     g08104(.I(new_n8159_), .ZN(new_n8169_));
  AOI21_X1   g08105(.A1(new_n8169_), .A2(new_n8160_), .B(new_n8116_), .ZN(new_n8170_));
  INV_X1     g08106(.I(new_n8163_), .ZN(new_n8171_));
  AOI21_X1   g08107(.A1(new_n8171_), .A2(new_n8164_), .B(new_n8117_), .ZN(new_n8172_));
  OAI21_X1   g08108(.A1(new_n8170_), .A2(new_n8172_), .B(new_n8168_), .ZN(new_n8173_));
  OAI21_X1   g08109(.A1(new_n7956_), .A2(new_n8025_), .B(new_n8027_), .ZN(new_n8174_));
  NAND3_X1   g08110(.A1(new_n8173_), .A2(new_n8167_), .A3(new_n8174_), .ZN(new_n8175_));
  NAND3_X1   g08111(.A1(new_n8041_), .A2(new_n8109_), .A3(new_n8175_), .ZN(new_n8176_));
  AOI21_X1   g08112(.A1(new_n8162_), .A2(new_n8166_), .B(new_n8168_), .ZN(new_n8177_));
  INV_X1     g08113(.I(new_n8177_), .ZN(new_n8178_));
  NAND2_X1   g08114(.A1(new_n8176_), .A2(new_n8178_), .ZN(new_n8179_));
  NOR2_X1    g08115(.A1(new_n7952_), .A2(new_n7918_), .ZN(new_n8180_));
  AOI21_X1   g08116(.A1(new_n7917_), .A2(new_n7919_), .B(new_n8034_), .ZN(new_n8181_));
  NOR3_X1    g08117(.A1(new_n7952_), .A2(new_n7918_), .A3(new_n8029_), .ZN(new_n8182_));
  OAI22_X1   g08118(.A1(new_n8182_), .A2(new_n8181_), .B1(new_n8180_), .B2(new_n8039_), .ZN(new_n8183_));
  NOR3_X1    g08119(.A1(new_n8168_), .A2(new_n8172_), .A3(new_n8170_), .ZN(new_n8184_));
  AOI21_X1   g08120(.A1(new_n8162_), .A2(new_n8166_), .B(new_n8115_), .ZN(new_n8185_));
  INV_X1     g08121(.I(new_n8174_), .ZN(new_n8186_));
  NOR3_X1    g08122(.A1(new_n8184_), .A2(new_n8185_), .A3(new_n8186_), .ZN(new_n8187_));
  NOR3_X1    g08123(.A1(new_n8183_), .A2(new_n8108_), .A3(new_n8187_), .ZN(new_n8188_));
  NAND2_X1   g08124(.A1(new_n3168_), .A2(new_n6180_), .ZN(new_n8189_));
  NAND2_X1   g08125(.A1(new_n3247_), .A2(new_n6095_), .ZN(new_n8190_));
  NAND4_X1   g08126(.A1(new_n3758_), .A2(new_n6081_), .A3(new_n8189_), .A4(new_n8190_), .ZN(new_n8191_));
  XOR2_X1    g08127(.A1(new_n8191_), .A2(\a[14] ), .Z(new_n8192_));
  OAI22_X1   g08128(.A1(new_n2614_), .A2(new_n4291_), .B1(new_n2665_), .B2(new_n4297_), .ZN(new_n8193_));
  NAND2_X1   g08129(.A1(new_n2728_), .A2(new_n4469_), .ZN(new_n8194_));
  AOI21_X1   g08130(.A1(new_n8194_), .A2(new_n8193_), .B(new_n4468_), .ZN(new_n8195_));
  NAND2_X1   g08131(.A1(new_n2733_), .A2(new_n8195_), .ZN(new_n8196_));
  XOR2_X1    g08132(.A1(new_n8196_), .A2(\a[17] ), .Z(new_n8197_));
  AOI21_X1   g08133(.A1(new_n4679_), .A2(new_n4680_), .B(new_n4487_), .ZN(new_n8198_));
  XOR2_X1    g08134(.A1(new_n4491_), .A2(new_n4676_), .Z(new_n8199_));
  NOR2_X1    g08135(.A1(new_n8199_), .A2(new_n4488_), .ZN(new_n8200_));
  NOR2_X1    g08136(.A1(new_n8145_), .A2(new_n8133_), .ZN(new_n8201_));
  NOR4_X1    g08137(.A1(new_n8200_), .A2(new_n8198_), .A3(new_n8201_), .A4(new_n8146_), .ZN(new_n8202_));
  NOR2_X1    g08138(.A1(new_n8200_), .A2(new_n8198_), .ZN(new_n8203_));
  NOR2_X1    g08139(.A1(new_n8201_), .A2(new_n8146_), .ZN(new_n8204_));
  NOR2_X1    g08140(.A1(new_n8203_), .A2(new_n8204_), .ZN(new_n8205_));
  NOR2_X1    g08141(.A1(new_n8205_), .A2(new_n8202_), .ZN(new_n8206_));
  NOR2_X1    g08142(.A1(new_n8206_), .A2(new_n8197_), .ZN(new_n8207_));
  INV_X1     g08143(.I(new_n8197_), .ZN(new_n8208_));
  XNOR2_X1   g08144(.A1(new_n8203_), .A2(new_n8204_), .ZN(new_n8209_));
  NOR2_X1    g08145(.A1(new_n8209_), .A2(new_n8208_), .ZN(new_n8210_));
  NOR2_X1    g08146(.A1(new_n8210_), .A2(new_n8207_), .ZN(new_n8211_));
  INV_X1     g08147(.I(new_n8128_), .ZN(new_n8212_));
  NAND2_X1   g08148(.A1(new_n8154_), .A2(new_n8212_), .ZN(new_n8213_));
  NAND2_X1   g08149(.A1(new_n8213_), .A2(new_n8155_), .ZN(new_n8214_));
  XOR2_X1    g08150(.A1(new_n8211_), .A2(new_n8214_), .Z(new_n8215_));
  NOR2_X1    g08151(.A1(new_n8215_), .A2(new_n8192_), .ZN(new_n8216_));
  INV_X1     g08152(.I(new_n8192_), .ZN(new_n8217_));
  INV_X1     g08153(.I(new_n8211_), .ZN(new_n8218_));
  NOR2_X1    g08154(.A1(new_n8218_), .A2(new_n8214_), .ZN(new_n8219_));
  INV_X1     g08155(.I(new_n8219_), .ZN(new_n8220_));
  NAND2_X1   g08156(.A1(new_n8218_), .A2(new_n8214_), .ZN(new_n8221_));
  AOI21_X1   g08157(.A1(new_n8220_), .A2(new_n8221_), .B(new_n8217_), .ZN(new_n8222_));
  NOR2_X1    g08158(.A1(new_n8222_), .A2(new_n8216_), .ZN(new_n8223_));
  OAI21_X1   g08159(.A1(new_n8188_), .A2(new_n8177_), .B(new_n8223_), .ZN(new_n8224_));
  INV_X1     g08160(.I(new_n8223_), .ZN(new_n8225_));
  NAND3_X1   g08161(.A1(new_n8176_), .A2(new_n8178_), .A3(new_n8225_), .ZN(new_n8226_));
  AOI21_X1   g08162(.A1(new_n8117_), .A2(new_n8164_), .B(new_n8163_), .ZN(new_n8227_));
  INV_X1     g08163(.I(new_n8227_), .ZN(new_n8228_));
  AOI22_X1   g08164(.A1(new_n8224_), .A2(new_n8226_), .B1(new_n8179_), .B2(new_n8228_), .ZN(new_n8229_));
  AOI22_X1   g08165(.A1(new_n3253_), .A2(new_n6081_), .B1(new_n3247_), .B2(new_n6180_), .ZN(new_n8230_));
  INV_X1     g08166(.I(new_n8230_), .ZN(new_n8231_));
  OAI21_X1   g08167(.A1(new_n4684_), .A2(new_n4686_), .B(new_n4476_), .ZN(new_n8232_));
  XOR2_X1    g08168(.A1(new_n4481_), .A2(new_n4683_), .Z(new_n8233_));
  OAI21_X1   g08169(.A1(new_n4476_), .A2(new_n8233_), .B(new_n8232_), .ZN(new_n8234_));
  INV_X1     g08170(.I(new_n8202_), .ZN(new_n8235_));
  AOI21_X1   g08171(.A1(new_n8235_), .A2(new_n8208_), .B(new_n8205_), .ZN(new_n8236_));
  XOR2_X1    g08172(.A1(new_n8234_), .A2(new_n8236_), .Z(new_n8237_));
  XOR2_X1    g08173(.A1(new_n8237_), .A2(\a[14] ), .Z(new_n8238_));
  NOR2_X1    g08174(.A1(new_n8238_), .A2(new_n8231_), .ZN(new_n8239_));
  AND2_X2    g08175(.A1(new_n8238_), .A2(new_n8231_), .Z(new_n8240_));
  NOR2_X1    g08176(.A1(new_n8240_), .A2(new_n8239_), .ZN(new_n8241_));
  INV_X1     g08177(.I(new_n8241_), .ZN(new_n8242_));
  INV_X1     g08178(.I(new_n8236_), .ZN(new_n8243_));
  XOR2_X1    g08179(.A1(new_n8230_), .A2(\a[14] ), .Z(new_n8244_));
  NOR3_X1    g08180(.A1(new_n8234_), .A2(new_n8243_), .A3(new_n8244_), .ZN(new_n8245_));
  AOI21_X1   g08181(.A1(new_n8234_), .A2(new_n8243_), .B(new_n8245_), .ZN(new_n8246_));
  XNOR2_X1   g08182(.A1(new_n4691_), .A2(new_n4696_), .ZN(new_n8247_));
  INV_X1     g08183(.I(new_n4697_), .ZN(new_n8248_));
  OAI21_X1   g08184(.A1(new_n8248_), .A2(new_n4698_), .B(new_n4687_), .ZN(new_n8249_));
  OAI21_X1   g08185(.A1(new_n4687_), .A2(new_n8247_), .B(new_n8249_), .ZN(new_n8250_));
  XOR2_X1    g08186(.A1(new_n8250_), .A2(new_n8246_), .Z(new_n8251_));
  OAI21_X1   g08187(.A1(new_n8192_), .A2(new_n8219_), .B(new_n8221_), .ZN(new_n8252_));
  INV_X1     g08188(.I(new_n8252_), .ZN(new_n8253_));
  NOR2_X1    g08189(.A1(new_n8251_), .A2(new_n8253_), .ZN(new_n8254_));
  INV_X1     g08190(.I(new_n8254_), .ZN(new_n8255_));
  NAND3_X1   g08191(.A1(new_n8229_), .A2(new_n8242_), .A3(new_n8255_), .ZN(new_n8256_));
  XOR2_X1    g08192(.A1(new_n4467_), .A2(new_n4699_), .Z(new_n8257_));
  NAND2_X1   g08193(.A1(new_n8250_), .A2(new_n8246_), .ZN(new_n8258_));
  INV_X1     g08194(.I(new_n8258_), .ZN(new_n8259_));
  NOR2_X1    g08195(.A1(new_n8257_), .A2(new_n8259_), .ZN(new_n8260_));
  AOI21_X1   g08196(.A1(new_n8256_), .A2(new_n8260_), .B(new_n4700_), .ZN(new_n8261_));
  AOI22_X1   g08197(.A1(new_n3253_), .A2(new_n4295_), .B1(new_n3247_), .B2(new_n4292_), .ZN(new_n8262_));
  INV_X1     g08198(.I(new_n8262_), .ZN(new_n8263_));
  OAI21_X1   g08199(.A1(new_n4157_), .A2(new_n4155_), .B(new_n4103_), .ZN(new_n8264_));
  XOR2_X1    g08200(.A1(new_n4106_), .A2(new_n4153_), .Z(new_n8265_));
  OAI21_X1   g08201(.A1(new_n4103_), .A2(new_n8265_), .B(new_n8264_), .ZN(new_n8266_));
  INV_X1     g08202(.I(new_n4273_), .ZN(new_n8267_));
  AOI21_X1   g08203(.A1(new_n8267_), .A2(new_n4277_), .B(new_n4274_), .ZN(new_n8268_));
  XOR2_X1    g08204(.A1(new_n8266_), .A2(new_n8268_), .Z(new_n8269_));
  XOR2_X1    g08205(.A1(new_n8269_), .A2(\a[17] ), .Z(new_n8270_));
  NOR2_X1    g08206(.A1(new_n8270_), .A2(new_n8263_), .ZN(new_n8271_));
  NAND2_X1   g08207(.A1(new_n8270_), .A2(new_n8263_), .ZN(new_n8272_));
  INV_X1     g08208(.I(new_n8272_), .ZN(new_n8273_));
  NOR2_X1    g08209(.A1(new_n8273_), .A2(new_n8271_), .ZN(new_n8274_));
  INV_X1     g08210(.I(new_n8268_), .ZN(new_n8275_));
  XOR2_X1    g08211(.A1(new_n8262_), .A2(\a[17] ), .Z(new_n8276_));
  NOR3_X1    g08212(.A1(new_n8275_), .A2(new_n8266_), .A3(new_n8276_), .ZN(new_n8277_));
  AOI21_X1   g08213(.A1(new_n8266_), .A2(new_n8275_), .B(new_n8277_), .ZN(new_n8278_));
  XOR2_X1    g08214(.A1(new_n4161_), .A2(new_n4168_), .Z(new_n8279_));
  OAI21_X1   g08215(.A1(new_n4169_), .A2(new_n4171_), .B(new_n4158_), .ZN(new_n8280_));
  OAI21_X1   g08216(.A1(new_n4158_), .A2(new_n8279_), .B(new_n8280_), .ZN(new_n8281_));
  XNOR2_X1   g08217(.A1(new_n8281_), .A2(new_n8278_), .ZN(new_n8282_));
  OAI21_X1   g08218(.A1(new_n4280_), .A2(new_n4461_), .B(new_n4462_), .ZN(new_n8283_));
  NAND2_X1   g08219(.A1(new_n8282_), .A2(new_n8283_), .ZN(new_n8284_));
  INV_X1     g08220(.I(new_n8284_), .ZN(new_n8285_));
  NOR3_X1    g08221(.A1(new_n8261_), .A2(new_n8274_), .A3(new_n8285_), .ZN(new_n8286_));
  XOR2_X1    g08222(.A1(new_n4094_), .A2(new_n4172_), .Z(new_n8287_));
  NAND2_X1   g08223(.A1(new_n8281_), .A2(new_n8278_), .ZN(new_n8288_));
  INV_X1     g08224(.I(new_n8288_), .ZN(new_n8289_));
  NOR2_X1    g08225(.A1(new_n8287_), .A2(new_n8289_), .ZN(new_n8290_));
  INV_X1     g08226(.I(new_n8290_), .ZN(new_n8291_));
  OAI21_X1   g08227(.A1(new_n8286_), .A2(new_n8291_), .B(new_n4174_), .ZN(new_n8292_));
  AOI22_X1   g08228(.A1(new_n3253_), .A2(new_n3773_), .B1(new_n3247_), .B2(new_n3770_), .ZN(new_n8293_));
  INV_X1     g08229(.I(new_n8293_), .ZN(new_n8294_));
  OAI22_X1   g08230(.A1(new_n3176_), .A2(new_n3780_), .B1(new_n2665_), .B2(new_n3310_), .ZN(new_n8295_));
  NAND2_X1   g08231(.A1(new_n2728_), .A2(new_n3782_), .ZN(new_n8296_));
  AOI21_X1   g08232(.A1(new_n8295_), .A2(new_n8296_), .B(new_n3302_), .ZN(new_n8297_));
  NAND2_X1   g08233(.A1(new_n3273_), .A2(new_n8297_), .ZN(new_n8298_));
  XOR2_X1    g08234(.A1(new_n8298_), .A2(\a[23] ), .Z(new_n8299_));
  OAI22_X1   g08235(.A1(new_n2614_), .A2(new_n3318_), .B1(new_n529_), .B2(new_n3268_), .ZN(new_n8300_));
  NAND2_X1   g08236(.A1(new_n2718_), .A2(new_n3323_), .ZN(new_n8301_));
  AOI21_X1   g08237(.A1(new_n8301_), .A2(new_n8300_), .B(new_n3260_), .ZN(new_n8302_));
  NAND2_X1   g08238(.A1(new_n3074_), .A2(new_n8302_), .ZN(new_n8303_));
  XOR2_X1    g08239(.A1(new_n8303_), .A2(\a[26] ), .Z(new_n8304_));
  INV_X1     g08240(.I(new_n3549_), .ZN(new_n8305_));
  AOI21_X1   g08241(.A1(new_n8305_), .A2(new_n3548_), .B(new_n3550_), .ZN(new_n8306_));
  OAI21_X1   g08242(.A1(new_n1180_), .A2(new_n2767_), .B(new_n2764_), .ZN(new_n8307_));
  OAI22_X1   g08243(.A1(new_n1008_), .A2(new_n2772_), .B1(new_n1121_), .B2(new_n2771_), .ZN(new_n8308_));
  NOR2_X1    g08244(.A1(new_n8308_), .A2(new_n8307_), .ZN(new_n8309_));
  NAND2_X1   g08245(.A1(new_n3562_), .A2(new_n8309_), .ZN(new_n8310_));
  INV_X1     g08246(.I(new_n970_), .ZN(new_n8311_));
  NOR2_X1    g08247(.A1(new_n413_), .A2(new_n772_), .ZN(new_n8312_));
  NAND4_X1   g08248(.A1(new_n597_), .A2(new_n2091_), .A3(new_n8312_), .A4(new_n1526_), .ZN(new_n8313_));
  INV_X1     g08249(.I(new_n1367_), .ZN(new_n8314_));
  NOR3_X1    g08250(.A1(new_n8314_), .A2(new_n173_), .A3(new_n721_), .ZN(new_n8315_));
  NAND2_X1   g08251(.A1(new_n3989_), .A2(new_n8315_), .ZN(new_n8316_));
  NOR3_X1    g08252(.A1(new_n8316_), .A2(new_n3963_), .A3(new_n8313_), .ZN(new_n8317_));
  NOR4_X1    g08253(.A1(new_n147_), .A2(new_n505_), .A3(new_n130_), .A4(new_n468_), .ZN(new_n8318_));
  NAND2_X1   g08254(.A1(new_n612_), .A2(new_n1018_), .ZN(new_n8319_));
  NOR4_X1    g08255(.A1(new_n8318_), .A2(new_n8319_), .A3(new_n695_), .A4(new_n1787_), .ZN(new_n8320_));
  NOR4_X1    g08256(.A1(new_n615_), .A2(new_n282_), .A3(new_n312_), .A4(new_n335_), .ZN(new_n8321_));
  NOR3_X1    g08257(.A1(new_n579_), .A2(new_n737_), .A3(new_n8321_), .ZN(new_n8322_));
  NAND3_X1   g08258(.A1(new_n8317_), .A2(new_n8320_), .A3(new_n8322_), .ZN(new_n8323_));
  NAND4_X1   g08259(.A1(new_n3502_), .A2(new_n221_), .A3(new_n1327_), .A4(new_n1838_), .ZN(new_n8324_));
  NOR4_X1    g08260(.A1(new_n8324_), .A2(new_n2870_), .A3(new_n238_), .A4(new_n453_), .ZN(new_n8325_));
  NOR3_X1    g08261(.A1(new_n988_), .A2(new_n2811_), .A3(new_n1078_), .ZN(new_n8326_));
  NAND4_X1   g08262(.A1(new_n8325_), .A2(new_n8326_), .A3(new_n1458_), .A4(new_n2489_), .ZN(new_n8327_));
  NOR4_X1    g08263(.A1(new_n8323_), .A2(new_n8311_), .A3(new_n2017_), .A4(new_n8327_), .ZN(new_n8328_));
  NAND2_X1   g08264(.A1(new_n8328_), .A2(new_n3986_), .ZN(new_n8329_));
  NAND2_X1   g08265(.A1(new_n8329_), .A2(new_n3032_), .ZN(new_n8330_));
  NOR2_X1    g08266(.A1(new_n8329_), .A2(new_n3032_), .ZN(new_n8331_));
  INV_X1     g08267(.I(new_n8331_), .ZN(new_n8332_));
  AOI21_X1   g08268(.A1(new_n8330_), .A2(new_n8332_), .B(new_n8310_), .ZN(new_n8333_));
  INV_X1     g08269(.I(new_n8310_), .ZN(new_n8334_));
  XOR2_X1    g08270(.A1(new_n8329_), .A2(new_n3031_), .Z(new_n8335_));
  NOR2_X1    g08271(.A1(new_n8334_), .A2(new_n8335_), .ZN(new_n8336_));
  NOR2_X1    g08272(.A1(new_n8336_), .A2(new_n8333_), .ZN(new_n8337_));
  NOR2_X1    g08273(.A1(new_n3334_), .A2(new_n3377_), .ZN(new_n8338_));
  NOR2_X1    g08274(.A1(new_n8338_), .A2(new_n3375_), .ZN(new_n8339_));
  INV_X1     g08275(.I(new_n8339_), .ZN(new_n8340_));
  XOR2_X1    g08276(.A1(new_n8337_), .A2(new_n8340_), .Z(new_n8341_));
  NOR2_X1    g08277(.A1(new_n8306_), .A2(new_n8341_), .ZN(new_n8342_));
  INV_X1     g08278(.I(new_n8306_), .ZN(new_n8343_));
  NOR3_X1    g08279(.A1(new_n8336_), .A2(new_n8333_), .A3(new_n8340_), .ZN(new_n8344_));
  NOR2_X1    g08280(.A1(new_n8337_), .A2(new_n8339_), .ZN(new_n8345_));
  NOR2_X1    g08281(.A1(new_n8345_), .A2(new_n8344_), .ZN(new_n8346_));
  NOR2_X1    g08282(.A1(new_n8343_), .A2(new_n8346_), .ZN(new_n8347_));
  NOR2_X1    g08283(.A1(new_n8347_), .A2(new_n8342_), .ZN(new_n8348_));
  OAI22_X1   g08284(.A1(new_n2559_), .A2(new_n3175_), .B1(new_n896_), .B2(new_n2747_), .ZN(new_n8349_));
  NAND2_X1   g08285(.A1(new_n814_), .A2(new_n3275_), .ZN(new_n8350_));
  AOI21_X1   g08286(.A1(new_n8349_), .A2(new_n8350_), .B(new_n2737_), .ZN(new_n8351_));
  NAND2_X1   g08287(.A1(new_n3624_), .A2(new_n8351_), .ZN(new_n8352_));
  XOR2_X1    g08288(.A1(new_n8352_), .A2(\a[29] ), .Z(new_n8353_));
  INV_X1     g08289(.I(new_n8353_), .ZN(new_n8354_));
  NOR2_X1    g08290(.A1(new_n8348_), .A2(new_n8354_), .ZN(new_n8355_));
  INV_X1     g08291(.I(new_n8348_), .ZN(new_n8356_));
  NOR2_X1    g08292(.A1(new_n8356_), .A2(new_n8353_), .ZN(new_n8357_));
  NOR2_X1    g08293(.A1(new_n8357_), .A2(new_n8355_), .ZN(new_n8358_));
  NOR2_X1    g08294(.A1(new_n8358_), .A2(new_n8304_), .ZN(new_n8359_));
  INV_X1     g08295(.I(new_n8304_), .ZN(new_n8360_));
  XOR2_X1    g08296(.A1(new_n8348_), .A2(new_n8353_), .Z(new_n8361_));
  NOR2_X1    g08297(.A1(new_n8361_), .A2(new_n8360_), .ZN(new_n8362_));
  INV_X1     g08298(.I(new_n3605_), .ZN(new_n8363_));
  AOI21_X1   g08299(.A1(new_n8363_), .A2(new_n3611_), .B(new_n3608_), .ZN(new_n8364_));
  INV_X1     g08300(.I(new_n8364_), .ZN(new_n8365_));
  NOR3_X1    g08301(.A1(new_n8359_), .A2(new_n8362_), .A3(new_n8365_), .ZN(new_n8366_));
  NOR2_X1    g08302(.A1(new_n8359_), .A2(new_n8362_), .ZN(new_n8367_));
  NOR2_X1    g08303(.A1(new_n8367_), .A2(new_n8364_), .ZN(new_n8368_));
  NOR2_X1    g08304(.A1(new_n8368_), .A2(new_n8366_), .ZN(new_n8369_));
  NOR2_X1    g08305(.A1(new_n8369_), .A2(new_n8299_), .ZN(new_n8370_));
  INV_X1     g08306(.I(new_n8299_), .ZN(new_n8371_));
  XOR2_X1    g08307(.A1(new_n8367_), .A2(new_n8365_), .Z(new_n8372_));
  NOR2_X1    g08308(.A1(new_n8372_), .A2(new_n8371_), .ZN(new_n8373_));
  NOR2_X1    g08309(.A1(new_n8373_), .A2(new_n8370_), .ZN(new_n8374_));
  INV_X1     g08310(.I(new_n3745_), .ZN(new_n8375_));
  AOI21_X1   g08311(.A1(new_n8375_), .A2(new_n3750_), .B(new_n3747_), .ZN(new_n8376_));
  XOR2_X1    g08312(.A1(new_n8374_), .A2(new_n8376_), .Z(new_n8377_));
  XOR2_X1    g08313(.A1(new_n8377_), .A2(new_n3035_), .Z(new_n8378_));
  NOR2_X1    g08314(.A1(new_n8378_), .A2(new_n8294_), .ZN(new_n8379_));
  NAND2_X1   g08315(.A1(new_n8378_), .A2(new_n8294_), .ZN(new_n8380_));
  INV_X1     g08316(.I(new_n8380_), .ZN(new_n8381_));
  NOR2_X1    g08317(.A1(new_n8381_), .A2(new_n8379_), .ZN(new_n8382_));
  INV_X1     g08318(.I(new_n8382_), .ZN(new_n8383_));
  INV_X1     g08319(.I(new_n8366_), .ZN(new_n8384_));
  AOI21_X1   g08320(.A1(new_n8384_), .A2(new_n8371_), .B(new_n8368_), .ZN(new_n8385_));
  OAI22_X1   g08321(.A1(new_n3176_), .A2(new_n3306_), .B1(new_n3142_), .B2(new_n3780_), .ZN(new_n8386_));
  NAND2_X1   g08322(.A1(new_n2728_), .A2(new_n5291_), .ZN(new_n8387_));
  AOI21_X1   g08323(.A1(new_n8386_), .A2(new_n8387_), .B(new_n3302_), .ZN(new_n8388_));
  NAND2_X1   g08324(.A1(new_n3174_), .A2(new_n8388_), .ZN(new_n8389_));
  XOR2_X1    g08325(.A1(new_n8389_), .A2(\a[23] ), .Z(new_n8390_));
  INV_X1     g08326(.I(new_n8390_), .ZN(new_n8391_));
  OAI22_X1   g08327(.A1(new_n694_), .A2(new_n3268_), .B1(new_n2665_), .B2(new_n3318_), .ZN(new_n8392_));
  NAND2_X1   g08328(.A1(new_n2615_), .A2(new_n3323_), .ZN(new_n8393_));
  AOI21_X1   g08329(.A1(new_n8392_), .A2(new_n8393_), .B(new_n3260_), .ZN(new_n8394_));
  NAND2_X1   g08330(.A1(new_n3188_), .A2(new_n8394_), .ZN(new_n8395_));
  XOR2_X1    g08331(.A1(new_n8395_), .A2(\a[26] ), .Z(new_n8396_));
  OAI22_X1   g08332(.A1(new_n813_), .A2(new_n2747_), .B1(new_n529_), .B2(new_n3175_), .ZN(new_n8397_));
  NAND2_X1   g08333(.A1(new_n2563_), .A2(new_n3275_), .ZN(new_n8398_));
  AOI21_X1   g08334(.A1(new_n8398_), .A2(new_n8397_), .B(new_n2737_), .ZN(new_n8399_));
  NAND2_X1   g08335(.A1(new_n3051_), .A2(new_n8399_), .ZN(new_n8400_));
  XOR2_X1    g08336(.A1(new_n8400_), .A2(\a[29] ), .Z(new_n8401_));
  INV_X1     g08337(.I(new_n8401_), .ZN(new_n8402_));
  INV_X1     g08338(.I(new_n8344_), .ZN(new_n8403_));
  AOI21_X1   g08339(.A1(new_n8343_), .A2(new_n8403_), .B(new_n8345_), .ZN(new_n8404_));
  AOI21_X1   g08340(.A1(new_n8334_), .A2(new_n8330_), .B(new_n8331_), .ZN(new_n8405_));
  OAI21_X1   g08341(.A1(new_n1008_), .A2(new_n2767_), .B(new_n2764_), .ZN(new_n8406_));
  OAI22_X1   g08342(.A1(new_n896_), .A2(new_n2772_), .B1(new_n1180_), .B2(new_n2771_), .ZN(new_n8407_));
  NOR2_X1    g08343(.A1(new_n8406_), .A2(new_n8407_), .ZN(new_n8408_));
  NOR2_X1    g08344(.A1(new_n3033_), .A2(new_n3036_), .ZN(new_n8409_));
  NOR2_X1    g08345(.A1(new_n8409_), .A2(new_n3000_), .ZN(new_n8410_));
  XOR2_X1    g08346(.A1(new_n3031_), .A2(\a[20] ), .Z(new_n8411_));
  INV_X1     g08347(.I(new_n8411_), .ZN(new_n8412_));
  AOI21_X1   g08348(.A1(new_n3000_), .A2(new_n8412_), .B(new_n8410_), .ZN(new_n8413_));
  INV_X1     g08349(.I(new_n8413_), .ZN(new_n8414_));
  AOI21_X1   g08350(.A1(new_n3596_), .A2(new_n8408_), .B(new_n8414_), .ZN(new_n8415_));
  NAND2_X1   g08351(.A1(new_n3596_), .A2(new_n8408_), .ZN(new_n8416_));
  NOR2_X1    g08352(.A1(new_n8416_), .A2(new_n8413_), .ZN(new_n8417_));
  NOR2_X1    g08353(.A1(new_n8417_), .A2(new_n8415_), .ZN(new_n8418_));
  NOR2_X1    g08354(.A1(new_n8418_), .A2(new_n8405_), .ZN(new_n8419_));
  INV_X1     g08355(.I(new_n8405_), .ZN(new_n8420_));
  XOR2_X1    g08356(.A1(new_n8416_), .A2(new_n8414_), .Z(new_n8421_));
  NOR2_X1    g08357(.A1(new_n8421_), .A2(new_n8420_), .ZN(new_n8422_));
  NOR2_X1    g08358(.A1(new_n8422_), .A2(new_n8419_), .ZN(new_n8423_));
  XOR2_X1    g08359(.A1(new_n8404_), .A2(new_n8423_), .Z(new_n8424_));
  NAND2_X1   g08360(.A1(new_n8424_), .A2(new_n8402_), .ZN(new_n8425_));
  AND2_X2    g08361(.A1(new_n8404_), .A2(new_n8423_), .Z(new_n8426_));
  NOR2_X1    g08362(.A1(new_n8404_), .A2(new_n8423_), .ZN(new_n8427_));
  OAI21_X1   g08363(.A1(new_n8426_), .A2(new_n8427_), .B(new_n8401_), .ZN(new_n8428_));
  NAND2_X1   g08364(.A1(new_n8425_), .A2(new_n8428_), .ZN(new_n8429_));
  INV_X1     g08365(.I(new_n8355_), .ZN(new_n8430_));
  AOI21_X1   g08366(.A1(new_n8360_), .A2(new_n8430_), .B(new_n8357_), .ZN(new_n8431_));
  AND2_X2    g08367(.A1(new_n8429_), .A2(new_n8431_), .Z(new_n8432_));
  INV_X1     g08368(.I(new_n8432_), .ZN(new_n8433_));
  NOR2_X1    g08369(.A1(new_n8429_), .A2(new_n8431_), .ZN(new_n8434_));
  INV_X1     g08370(.I(new_n8434_), .ZN(new_n8435_));
  AOI21_X1   g08371(.A1(new_n8433_), .A2(new_n8435_), .B(new_n8396_), .ZN(new_n8436_));
  INV_X1     g08372(.I(new_n8396_), .ZN(new_n8437_));
  XNOR2_X1   g08373(.A1(new_n8429_), .A2(new_n8431_), .ZN(new_n8438_));
  NOR2_X1    g08374(.A1(new_n8438_), .A2(new_n8437_), .ZN(new_n8439_));
  NOR3_X1    g08375(.A1(new_n8436_), .A2(new_n8439_), .A3(new_n8391_), .ZN(new_n8440_));
  NOR2_X1    g08376(.A1(new_n8436_), .A2(new_n8439_), .ZN(new_n8441_));
  NOR2_X1    g08377(.A1(new_n8441_), .A2(new_n8390_), .ZN(new_n8442_));
  NOR2_X1    g08378(.A1(new_n8442_), .A2(new_n8440_), .ZN(new_n8443_));
  NOR2_X1    g08379(.A1(new_n8443_), .A2(new_n8385_), .ZN(new_n8444_));
  INV_X1     g08380(.I(new_n8385_), .ZN(new_n8445_));
  XOR2_X1    g08381(.A1(new_n8441_), .A2(new_n8391_), .Z(new_n8446_));
  NOR2_X1    g08382(.A1(new_n8446_), .A2(new_n8445_), .ZN(new_n8447_));
  NOR2_X1    g08383(.A1(new_n8447_), .A2(new_n8444_), .ZN(new_n8448_));
  INV_X1     g08384(.I(new_n8374_), .ZN(new_n8449_));
  INV_X1     g08385(.I(new_n8376_), .ZN(new_n8450_));
  XOR2_X1    g08386(.A1(new_n8293_), .A2(\a[20] ), .Z(new_n8451_));
  NOR3_X1    g08387(.A1(new_n8449_), .A2(new_n8450_), .A3(new_n8451_), .ZN(new_n8452_));
  AOI21_X1   g08388(.A1(new_n8449_), .A2(new_n8450_), .B(new_n8452_), .ZN(new_n8453_));
  XNOR2_X1   g08389(.A1(new_n8448_), .A2(new_n8453_), .ZN(new_n8454_));
  NOR2_X1    g08390(.A1(new_n3753_), .A2(new_n4089_), .ZN(new_n8455_));
  NOR2_X1    g08391(.A1(new_n8455_), .A2(new_n4090_), .ZN(new_n8456_));
  INV_X1     g08392(.I(new_n8456_), .ZN(new_n8457_));
  NAND2_X1   g08393(.A1(new_n8454_), .A2(new_n8457_), .ZN(new_n8458_));
  NAND3_X1   g08394(.A1(new_n8292_), .A2(new_n8383_), .A3(new_n8458_), .ZN(new_n8459_));
  NAND2_X1   g08395(.A1(new_n8448_), .A2(new_n8453_), .ZN(new_n8460_));
  NAND2_X1   g08396(.A1(new_n8459_), .A2(new_n8460_), .ZN(new_n8461_));
  INV_X1     g08397(.I(new_n4700_), .ZN(new_n8462_));
  NOR2_X1    g08398(.A1(new_n8188_), .A2(new_n8177_), .ZN(new_n8463_));
  AOI21_X1   g08399(.A1(new_n8176_), .A2(new_n8178_), .B(new_n8225_), .ZN(new_n8464_));
  NOR3_X1    g08400(.A1(new_n8188_), .A2(new_n8177_), .A3(new_n8223_), .ZN(new_n8465_));
  OAI22_X1   g08401(.A1(new_n8465_), .A2(new_n8464_), .B1(new_n8463_), .B2(new_n8227_), .ZN(new_n8466_));
  NOR3_X1    g08402(.A1(new_n8466_), .A2(new_n8241_), .A3(new_n8254_), .ZN(new_n8467_));
  INV_X1     g08403(.I(new_n8260_), .ZN(new_n8468_));
  OAI21_X1   g08404(.A1(new_n8467_), .A2(new_n8468_), .B(new_n8462_), .ZN(new_n8469_));
  INV_X1     g08405(.I(new_n8274_), .ZN(new_n8470_));
  NAND3_X1   g08406(.A1(new_n8469_), .A2(new_n8470_), .A3(new_n8284_), .ZN(new_n8471_));
  AOI21_X1   g08407(.A1(new_n8471_), .A2(new_n8290_), .B(new_n4173_), .ZN(new_n8472_));
  INV_X1     g08408(.I(new_n8458_), .ZN(new_n8473_));
  NOR3_X1    g08409(.A1(new_n8472_), .A2(new_n8382_), .A3(new_n8473_), .ZN(new_n8474_));
  INV_X1     g08410(.I(new_n8460_), .ZN(new_n8475_));
  OAI22_X1   g08411(.A1(new_n2614_), .A2(new_n3268_), .B1(new_n2665_), .B2(new_n3322_), .ZN(new_n8476_));
  NAND2_X1   g08412(.A1(new_n2728_), .A2(new_n3317_), .ZN(new_n8477_));
  AOI21_X1   g08413(.A1(new_n8477_), .A2(new_n8476_), .B(new_n3260_), .ZN(new_n8478_));
  NAND2_X1   g08414(.A1(new_n2733_), .A2(new_n8478_), .ZN(new_n8479_));
  XOR2_X1    g08415(.A1(new_n8479_), .A2(\a[26] ), .Z(new_n8480_));
  OAI22_X1   g08416(.A1(new_n2559_), .A2(new_n2747_), .B1(new_n694_), .B2(new_n3175_), .ZN(new_n8481_));
  NAND2_X1   g08417(.A1(new_n2567_), .A2(new_n3275_), .ZN(new_n8482_));
  AOI21_X1   g08418(.A1(new_n8481_), .A2(new_n8482_), .B(new_n2737_), .ZN(new_n8483_));
  NAND2_X1   g08419(.A1(new_n2759_), .A2(new_n8483_), .ZN(new_n8484_));
  XOR2_X1    g08420(.A1(new_n8484_), .A2(\a[29] ), .Z(new_n8485_));
  INV_X1     g08421(.I(new_n8485_), .ZN(new_n8486_));
  AOI21_X1   g08422(.A1(new_n3038_), .A2(new_n3040_), .B(new_n2921_), .ZN(new_n8487_));
  XOR2_X1    g08423(.A1(new_n3037_), .A2(new_n2950_), .Z(new_n8488_));
  NOR2_X1    g08424(.A1(new_n2922_), .A2(new_n8488_), .ZN(new_n8489_));
  NOR2_X1    g08425(.A1(new_n8489_), .A2(new_n8487_), .ZN(new_n8490_));
  INV_X1     g08426(.I(new_n8415_), .ZN(new_n8491_));
  AOI21_X1   g08427(.A1(new_n8420_), .A2(new_n8491_), .B(new_n8417_), .ZN(new_n8492_));
  XOR2_X1    g08428(.A1(new_n8490_), .A2(new_n8492_), .Z(new_n8493_));
  INV_X1     g08429(.I(new_n8492_), .ZN(new_n8494_));
  NOR3_X1    g08430(.A1(new_n8494_), .A2(new_n8487_), .A3(new_n8489_), .ZN(new_n8495_));
  INV_X1     g08431(.I(new_n8495_), .ZN(new_n8496_));
  NOR2_X1    g08432(.A1(new_n8490_), .A2(new_n8492_), .ZN(new_n8497_));
  INV_X1     g08433(.I(new_n8497_), .ZN(new_n8498_));
  AOI21_X1   g08434(.A1(new_n8496_), .A2(new_n8498_), .B(new_n8486_), .ZN(new_n8499_));
  AOI21_X1   g08435(.A1(new_n8486_), .A2(new_n8493_), .B(new_n8499_), .ZN(new_n8500_));
  NOR2_X1    g08436(.A1(new_n8426_), .A2(new_n8401_), .ZN(new_n8501_));
  NOR2_X1    g08437(.A1(new_n8501_), .A2(new_n8427_), .ZN(new_n8502_));
  XOR2_X1    g08438(.A1(new_n8502_), .A2(new_n8500_), .Z(new_n8503_));
  NOR2_X1    g08439(.A1(new_n8503_), .A2(new_n8480_), .ZN(new_n8504_));
  INV_X1     g08440(.I(new_n8480_), .ZN(new_n8505_));
  INV_X1     g08441(.I(new_n8502_), .ZN(new_n8506_));
  NOR2_X1    g08442(.A1(new_n8506_), .A2(new_n8500_), .ZN(new_n8507_));
  INV_X1     g08443(.I(new_n8507_), .ZN(new_n8508_));
  NAND2_X1   g08444(.A1(new_n8506_), .A2(new_n8500_), .ZN(new_n8509_));
  AOI21_X1   g08445(.A1(new_n8508_), .A2(new_n8509_), .B(new_n8505_), .ZN(new_n8510_));
  NOR2_X1    g08446(.A1(new_n8510_), .A2(new_n8504_), .ZN(new_n8511_));
  NAND2_X1   g08447(.A1(new_n3168_), .A2(new_n5291_), .ZN(new_n8512_));
  NAND2_X1   g08448(.A1(new_n3247_), .A2(new_n3782_), .ZN(new_n8513_));
  NAND4_X1   g08449(.A1(new_n3758_), .A2(new_n3301_), .A3(new_n8512_), .A4(new_n8513_), .ZN(new_n8514_));
  XOR2_X1    g08450(.A1(new_n8514_), .A2(\a[23] ), .Z(new_n8515_));
  NAND2_X1   g08451(.A1(new_n8433_), .A2(new_n8437_), .ZN(new_n8516_));
  AOI21_X1   g08452(.A1(new_n8516_), .A2(new_n8435_), .B(new_n8515_), .ZN(new_n8517_));
  INV_X1     g08453(.I(new_n8515_), .ZN(new_n8518_));
  NAND2_X1   g08454(.A1(new_n8516_), .A2(new_n8435_), .ZN(new_n8519_));
  NOR2_X1    g08455(.A1(new_n8519_), .A2(new_n8518_), .ZN(new_n8520_));
  NOR2_X1    g08456(.A1(new_n8520_), .A2(new_n8517_), .ZN(new_n8521_));
  NOR2_X1    g08457(.A1(new_n8521_), .A2(new_n8511_), .ZN(new_n8522_));
  XOR2_X1    g08458(.A1(new_n8519_), .A2(new_n8515_), .Z(new_n8523_));
  INV_X1     g08459(.I(new_n8523_), .ZN(new_n8524_));
  AOI21_X1   g08460(.A1(new_n8524_), .A2(new_n8511_), .B(new_n8522_), .ZN(new_n8525_));
  OAI21_X1   g08461(.A1(new_n8474_), .A2(new_n8475_), .B(new_n8525_), .ZN(new_n8526_));
  INV_X1     g08462(.I(new_n8525_), .ZN(new_n8527_));
  NAND3_X1   g08463(.A1(new_n8459_), .A2(new_n8460_), .A3(new_n8527_), .ZN(new_n8528_));
  INV_X1     g08464(.I(new_n8440_), .ZN(new_n8529_));
  AOI21_X1   g08465(.A1(new_n8529_), .A2(new_n8445_), .B(new_n8442_), .ZN(new_n8530_));
  INV_X1     g08466(.I(new_n8530_), .ZN(new_n8531_));
  AOI22_X1   g08467(.A1(new_n8526_), .A2(new_n8528_), .B1(new_n8461_), .B2(new_n8531_), .ZN(new_n8532_));
  AOI22_X1   g08468(.A1(new_n3253_), .A2(new_n3301_), .B1(new_n3247_), .B2(new_n5291_), .ZN(new_n8533_));
  INV_X1     g08469(.I(new_n8533_), .ZN(new_n8534_));
  OAI22_X1   g08470(.A1(new_n3176_), .A2(new_n3318_), .B1(new_n2665_), .B2(new_n3268_), .ZN(new_n8535_));
  NAND2_X1   g08471(.A1(new_n2728_), .A2(new_n3323_), .ZN(new_n8536_));
  AOI21_X1   g08472(.A1(new_n8535_), .A2(new_n8536_), .B(new_n3260_), .ZN(new_n8537_));
  NAND2_X1   g08473(.A1(new_n3273_), .A2(new_n8537_), .ZN(new_n8538_));
  XOR2_X1    g08474(.A1(new_n8538_), .A2(\a[26] ), .Z(new_n8539_));
  AOI21_X1   g08475(.A1(new_n8486_), .A2(new_n8496_), .B(new_n8497_), .ZN(new_n8540_));
  INV_X1     g08476(.I(new_n8540_), .ZN(new_n8541_));
  OAI21_X1   g08477(.A1(new_n3043_), .A2(new_n3045_), .B(new_n3041_), .ZN(new_n8542_));
  XOR2_X1    g08478(.A1(new_n2950_), .A2(new_n2848_), .Z(new_n8543_));
  OAI21_X1   g08479(.A1(new_n3041_), .A2(new_n8543_), .B(new_n8542_), .ZN(new_n8544_));
  INV_X1     g08480(.I(new_n8544_), .ZN(new_n8545_));
  NOR2_X1    g08481(.A1(new_n896_), .A2(new_n2771_), .ZN(new_n8546_));
  INV_X1     g08482(.I(new_n8546_), .ZN(new_n8547_));
  AOI22_X1   g08483(.A1(new_n2563_), .A2(new_n3332_), .B1(new_n814_), .B2(new_n3189_), .ZN(new_n8548_));
  NAND4_X1   g08484(.A1(new_n3624_), .A2(new_n2764_), .A3(new_n8547_), .A4(new_n8548_), .ZN(new_n8549_));
  NOR2_X1    g08485(.A1(new_n8545_), .A2(new_n8549_), .ZN(new_n8550_));
  INV_X1     g08486(.I(new_n8550_), .ZN(new_n8551_));
  NAND2_X1   g08487(.A1(new_n8545_), .A2(new_n8549_), .ZN(new_n8552_));
  NAND2_X1   g08488(.A1(new_n8551_), .A2(new_n8552_), .ZN(new_n8553_));
  NAND2_X1   g08489(.A1(new_n8553_), .A2(new_n8541_), .ZN(new_n8554_));
  XOR2_X1    g08490(.A1(new_n8544_), .A2(new_n8549_), .Z(new_n8555_));
  OAI21_X1   g08491(.A1(new_n8541_), .A2(new_n8555_), .B(new_n8554_), .ZN(new_n8556_));
  OAI22_X1   g08492(.A1(new_n2614_), .A2(new_n3175_), .B1(new_n529_), .B2(new_n2747_), .ZN(new_n8557_));
  NAND2_X1   g08493(.A1(new_n2718_), .A2(new_n3275_), .ZN(new_n8558_));
  AOI21_X1   g08494(.A1(new_n8558_), .A2(new_n8557_), .B(new_n2737_), .ZN(new_n8559_));
  NAND2_X1   g08495(.A1(new_n3074_), .A2(new_n8559_), .ZN(new_n8560_));
  XOR2_X1    g08496(.A1(new_n8560_), .A2(\a[29] ), .Z(new_n8561_));
  INV_X1     g08497(.I(new_n8561_), .ZN(new_n8562_));
  NOR2_X1    g08498(.A1(new_n8556_), .A2(new_n8562_), .ZN(new_n8563_));
  INV_X1     g08499(.I(new_n8563_), .ZN(new_n8564_));
  NAND2_X1   g08500(.A1(new_n8556_), .A2(new_n8562_), .ZN(new_n8565_));
  AOI21_X1   g08501(.A1(new_n8564_), .A2(new_n8565_), .B(new_n8539_), .ZN(new_n8566_));
  INV_X1     g08502(.I(new_n8539_), .ZN(new_n8567_));
  XOR2_X1    g08503(.A1(new_n8556_), .A2(new_n8561_), .Z(new_n8568_));
  NOR2_X1    g08504(.A1(new_n8568_), .A2(new_n8567_), .ZN(new_n8569_));
  NOR2_X1    g08505(.A1(new_n8569_), .A2(new_n8566_), .ZN(new_n8570_));
  OAI21_X1   g08506(.A1(new_n8480_), .A2(new_n8507_), .B(new_n8509_), .ZN(new_n8571_));
  INV_X1     g08507(.I(new_n8571_), .ZN(new_n8572_));
  XOR2_X1    g08508(.A1(new_n8570_), .A2(new_n8572_), .Z(new_n8573_));
  XOR2_X1    g08509(.A1(new_n8573_), .A2(new_n84_), .Z(new_n8574_));
  NOR2_X1    g08510(.A1(new_n8574_), .A2(new_n8534_), .ZN(new_n8575_));
  NAND2_X1   g08511(.A1(new_n8574_), .A2(new_n8534_), .ZN(new_n8576_));
  INV_X1     g08512(.I(new_n8576_), .ZN(new_n8577_));
  NOR2_X1    g08513(.A1(new_n8577_), .A2(new_n8575_), .ZN(new_n8578_));
  INV_X1     g08514(.I(new_n8578_), .ZN(new_n8579_));
  NOR2_X1    g08515(.A1(new_n8570_), .A2(new_n8572_), .ZN(new_n8580_));
  XOR2_X1    g08516(.A1(new_n8533_), .A2(\a[23] ), .Z(new_n8581_));
  NOR4_X1    g08517(.A1(new_n8571_), .A2(new_n8566_), .A3(new_n8569_), .A4(new_n8581_), .ZN(new_n8582_));
  NOR2_X1    g08518(.A1(new_n8580_), .A2(new_n8582_), .ZN(new_n8583_));
  OAI21_X1   g08519(.A1(new_n8539_), .A2(new_n8563_), .B(new_n8565_), .ZN(new_n8584_));
  AOI21_X1   g08520(.A1(new_n8541_), .A2(new_n8552_), .B(new_n8550_), .ZN(new_n8585_));
  OAI22_X1   g08521(.A1(new_n694_), .A2(new_n2747_), .B1(new_n2665_), .B2(new_n3175_), .ZN(new_n8586_));
  NAND2_X1   g08522(.A1(new_n2615_), .A2(new_n3275_), .ZN(new_n8587_));
  AOI21_X1   g08523(.A1(new_n8586_), .A2(new_n8587_), .B(new_n2737_), .ZN(new_n8588_));
  NAND2_X1   g08524(.A1(new_n3188_), .A2(new_n8588_), .ZN(new_n8589_));
  XOR2_X1    g08525(.A1(new_n8589_), .A2(\a[29] ), .Z(new_n8590_));
  XOR2_X1    g08526(.A1(new_n3055_), .A2(new_n3059_), .Z(new_n8591_));
  AND2_X2    g08527(.A1(new_n3047_), .A2(new_n8591_), .Z(new_n8592_));
  INV_X1     g08528(.I(new_n3061_), .ZN(new_n8593_));
  AOI21_X1   g08529(.A1(new_n3060_), .A2(new_n8593_), .B(new_n3047_), .ZN(new_n8594_));
  NOR3_X1    g08530(.A1(new_n8590_), .A2(new_n8592_), .A3(new_n8594_), .ZN(new_n8595_));
  INV_X1     g08531(.I(new_n8595_), .ZN(new_n8596_));
  INV_X1     g08532(.I(new_n8590_), .ZN(new_n8597_));
  NOR2_X1    g08533(.A1(new_n8592_), .A2(new_n8594_), .ZN(new_n8598_));
  NOR2_X1    g08534(.A1(new_n8597_), .A2(new_n8598_), .ZN(new_n8599_));
  INV_X1     g08535(.I(new_n8599_), .ZN(new_n8600_));
  AOI21_X1   g08536(.A1(new_n8600_), .A2(new_n8596_), .B(new_n8585_), .ZN(new_n8601_));
  INV_X1     g08537(.I(new_n8585_), .ZN(new_n8602_));
  XOR2_X1    g08538(.A1(new_n8590_), .A2(new_n8598_), .Z(new_n8603_));
  NOR2_X1    g08539(.A1(new_n8603_), .A2(new_n8602_), .ZN(new_n8604_));
  NOR2_X1    g08540(.A1(new_n8601_), .A2(new_n8604_), .ZN(new_n8605_));
  OAI22_X1   g08541(.A1(new_n3176_), .A2(new_n3322_), .B1(new_n3142_), .B2(new_n3318_), .ZN(new_n8606_));
  NAND2_X1   g08542(.A1(new_n2728_), .A2(new_n3267_), .ZN(new_n8607_));
  AOI21_X1   g08543(.A1(new_n8606_), .A2(new_n8607_), .B(new_n3260_), .ZN(new_n8608_));
  NAND2_X1   g08544(.A1(new_n3174_), .A2(new_n8608_), .ZN(new_n8609_));
  XOR2_X1    g08545(.A1(new_n8609_), .A2(\a[26] ), .Z(new_n8610_));
  XNOR2_X1   g08546(.A1(new_n8605_), .A2(new_n8610_), .ZN(new_n8611_));
  AND2_X2    g08547(.A1(new_n8605_), .A2(new_n8610_), .Z(new_n8612_));
  NOR2_X1    g08548(.A1(new_n8605_), .A2(new_n8610_), .ZN(new_n8613_));
  NOR2_X1    g08549(.A1(new_n8612_), .A2(new_n8613_), .ZN(new_n8614_));
  MUX2_X1    g08550(.I0(new_n8614_), .I1(new_n8611_), .S(new_n8584_), .Z(new_n8615_));
  XOR2_X1    g08551(.A1(new_n8583_), .A2(new_n8615_), .Z(new_n8616_));
  INV_X1     g08552(.I(new_n8520_), .ZN(new_n8617_));
  AOI21_X1   g08553(.A1(new_n8617_), .A2(new_n8511_), .B(new_n8517_), .ZN(new_n8618_));
  INV_X1     g08554(.I(new_n8618_), .ZN(new_n8619_));
  NAND2_X1   g08555(.A1(new_n8619_), .A2(new_n8616_), .ZN(new_n8620_));
  NAND3_X1   g08556(.A1(new_n8532_), .A2(new_n8579_), .A3(new_n8620_), .ZN(new_n8621_));
  NOR3_X1    g08557(.A1(new_n8615_), .A2(new_n8580_), .A3(new_n8582_), .ZN(new_n8622_));
  INV_X1     g08558(.I(new_n8622_), .ZN(new_n8623_));
  NAND2_X1   g08559(.A1(new_n8621_), .A2(new_n8623_), .ZN(new_n8624_));
  NOR2_X1    g08560(.A1(new_n8474_), .A2(new_n8475_), .ZN(new_n8625_));
  AOI21_X1   g08561(.A1(new_n8459_), .A2(new_n8460_), .B(new_n8527_), .ZN(new_n8626_));
  NOR3_X1    g08562(.A1(new_n8474_), .A2(new_n8475_), .A3(new_n8525_), .ZN(new_n8627_));
  OAI22_X1   g08563(.A1(new_n8627_), .A2(new_n8626_), .B1(new_n8625_), .B2(new_n8530_), .ZN(new_n8628_));
  INV_X1     g08564(.I(new_n8620_), .ZN(new_n8629_));
  NOR3_X1    g08565(.A1(new_n8628_), .A2(new_n8578_), .A3(new_n8629_), .ZN(new_n8630_));
  NAND2_X1   g08566(.A1(new_n3168_), .A2(new_n3267_), .ZN(new_n8631_));
  NAND2_X1   g08567(.A1(new_n3247_), .A2(new_n3323_), .ZN(new_n8632_));
  NAND4_X1   g08568(.A1(new_n3758_), .A2(new_n3259_), .A3(new_n8631_), .A4(new_n8632_), .ZN(new_n8633_));
  XOR2_X1    g08569(.A1(new_n8633_), .A2(\a[26] ), .Z(new_n8634_));
  NAND2_X1   g08570(.A1(new_n8600_), .A2(new_n8602_), .ZN(new_n8635_));
  NAND2_X1   g08571(.A1(new_n8635_), .A2(new_n8596_), .ZN(new_n8636_));
  XNOR2_X1   g08572(.A1(new_n2905_), .A2(new_n3062_), .ZN(new_n8637_));
  OAI21_X1   g08573(.A1(new_n3064_), .A2(new_n3066_), .B(new_n2754_), .ZN(new_n8638_));
  OAI21_X1   g08574(.A1(new_n2754_), .A2(new_n8637_), .B(new_n8638_), .ZN(new_n8639_));
  XOR2_X1    g08575(.A1(new_n8636_), .A2(new_n8639_), .Z(new_n8640_));
  NOR2_X1    g08576(.A1(new_n8640_), .A2(new_n8634_), .ZN(new_n8641_));
  INV_X1     g08577(.I(new_n8634_), .ZN(new_n8642_));
  INV_X1     g08578(.I(new_n8636_), .ZN(new_n8643_));
  NOR2_X1    g08579(.A1(new_n8643_), .A2(new_n8639_), .ZN(new_n8644_));
  INV_X1     g08580(.I(new_n8644_), .ZN(new_n8645_));
  NAND2_X1   g08581(.A1(new_n8643_), .A2(new_n8639_), .ZN(new_n8646_));
  AOI21_X1   g08582(.A1(new_n8645_), .A2(new_n8646_), .B(new_n8642_), .ZN(new_n8647_));
  NOR2_X1    g08583(.A1(new_n8647_), .A2(new_n8641_), .ZN(new_n8648_));
  OAI21_X1   g08584(.A1(new_n8630_), .A2(new_n8622_), .B(new_n8648_), .ZN(new_n8649_));
  INV_X1     g08585(.I(new_n8648_), .ZN(new_n8650_));
  NAND3_X1   g08586(.A1(new_n8621_), .A2(new_n8623_), .A3(new_n8650_), .ZN(new_n8651_));
  INV_X1     g08587(.I(new_n8612_), .ZN(new_n8652_));
  AOI21_X1   g08588(.A1(new_n8652_), .A2(new_n8584_), .B(new_n8613_), .ZN(new_n8653_));
  INV_X1     g08589(.I(new_n8653_), .ZN(new_n8654_));
  AOI22_X1   g08590(.A1(new_n8649_), .A2(new_n8651_), .B1(new_n8624_), .B2(new_n8654_), .ZN(new_n8655_));
  AOI21_X1   g08591(.A1(new_n8642_), .A2(new_n8646_), .B(new_n8644_), .ZN(new_n8656_));
  INV_X1     g08592(.I(new_n8656_), .ZN(new_n8657_));
  OAI21_X1   g08593(.A1(new_n8655_), .A2(new_n3295_), .B(new_n8657_), .ZN(new_n8658_));
  NOR2_X1    g08594(.A1(new_n8658_), .A2(new_n3292_), .ZN(new_n8659_));
  AND2_X2    g08595(.A1(new_n8658_), .A2(new_n3292_), .Z(new_n8660_));
  NOR2_X1    g08596(.A1(new_n8660_), .A2(new_n8659_), .ZN(new_n8661_));
  INV_X1     g08597(.I(new_n8661_), .ZN(new_n8662_));
  NOR2_X1    g08598(.A1(new_n8630_), .A2(new_n8622_), .ZN(new_n8663_));
  AOI21_X1   g08599(.A1(new_n8621_), .A2(new_n8623_), .B(new_n8650_), .ZN(new_n8664_));
  NOR3_X1    g08600(.A1(new_n8630_), .A2(new_n8622_), .A3(new_n8648_), .ZN(new_n8665_));
  OAI22_X1   g08601(.A1(new_n8665_), .A2(new_n8664_), .B1(new_n8663_), .B2(new_n8653_), .ZN(new_n8666_));
  XOR2_X1    g08602(.A1(new_n3295_), .A2(new_n8656_), .Z(new_n8667_));
  NOR2_X1    g08603(.A1(new_n8666_), .A2(new_n8667_), .ZN(new_n8668_));
  NOR2_X1    g08604(.A1(new_n3295_), .A2(new_n8657_), .ZN(new_n8669_));
  INV_X1     g08605(.I(new_n8669_), .ZN(new_n8670_));
  NAND2_X1   g08606(.A1(new_n3295_), .A2(new_n8657_), .ZN(new_n8671_));
  AOI21_X1   g08607(.A1(new_n8670_), .A2(new_n8671_), .B(new_n8655_), .ZN(new_n8672_));
  NOR2_X1    g08608(.A1(new_n8672_), .A2(new_n8668_), .ZN(new_n8673_));
  INV_X1     g08609(.I(new_n8673_), .ZN(new_n8674_));
  NAND2_X1   g08610(.A1(new_n8532_), .A2(new_n8579_), .ZN(new_n8675_));
  XOR2_X1    g08611(.A1(new_n8675_), .A2(new_n8616_), .Z(new_n8676_));
  XOR2_X1    g08612(.A1(new_n8532_), .A2(new_n8579_), .Z(new_n8677_));
  NAND2_X1   g08613(.A1(new_n8677_), .A2(new_n8619_), .ZN(new_n8678_));
  NOR2_X1    g08614(.A1(new_n8676_), .A2(new_n8678_), .ZN(new_n8679_));
  AND2_X2    g08615(.A1(new_n8676_), .A2(new_n8678_), .Z(new_n8680_));
  NOR2_X1    g08616(.A1(new_n8680_), .A2(new_n8679_), .ZN(new_n8681_));
  INV_X1     g08617(.I(new_n8681_), .ZN(new_n8682_));
  NAND2_X1   g08618(.A1(new_n8649_), .A2(new_n8651_), .ZN(new_n8683_));
  NAND2_X1   g08619(.A1(new_n8683_), .A2(new_n8653_), .ZN(new_n8684_));
  INV_X1     g08620(.I(new_n8684_), .ZN(new_n8685_));
  NOR2_X1    g08621(.A1(new_n8683_), .A2(new_n8653_), .ZN(new_n8686_));
  NOR2_X1    g08622(.A1(new_n8685_), .A2(new_n8686_), .ZN(new_n8687_));
  INV_X1     g08623(.I(new_n8687_), .ZN(new_n8688_));
  NOR2_X1    g08624(.A1(new_n8682_), .A2(new_n8688_), .ZN(new_n8689_));
  XOR2_X1    g08625(.A1(new_n8578_), .A2(new_n8619_), .Z(new_n8690_));
  NOR2_X1    g08626(.A1(new_n8628_), .A2(new_n8690_), .ZN(new_n8691_));
  XOR2_X1    g08627(.A1(new_n8578_), .A2(new_n8618_), .Z(new_n8692_));
  NOR2_X1    g08628(.A1(new_n8532_), .A2(new_n8692_), .ZN(new_n8693_));
  NOR2_X1    g08629(.A1(new_n8691_), .A2(new_n8693_), .ZN(new_n8694_));
  NAND2_X1   g08630(.A1(new_n8681_), .A2(new_n8694_), .ZN(new_n8695_));
  INV_X1     g08631(.I(new_n8694_), .ZN(new_n8696_));
  NOR2_X1    g08632(.A1(new_n8627_), .A2(new_n8626_), .ZN(new_n8697_));
  NOR2_X1    g08633(.A1(new_n8697_), .A2(new_n8531_), .ZN(new_n8698_));
  NAND2_X1   g08634(.A1(new_n8697_), .A2(new_n8531_), .ZN(new_n8699_));
  INV_X1     g08635(.I(new_n8699_), .ZN(new_n8700_));
  NOR2_X1    g08636(.A1(new_n8700_), .A2(new_n8698_), .ZN(new_n8701_));
  INV_X1     g08637(.I(new_n8701_), .ZN(new_n8702_));
  NOR2_X1    g08638(.A1(new_n8702_), .A2(new_n8696_), .ZN(new_n8703_));
  NAND2_X1   g08639(.A1(new_n8292_), .A2(new_n8383_), .ZN(new_n8704_));
  XOR2_X1    g08640(.A1(new_n8704_), .A2(new_n8454_), .Z(new_n8705_));
  XOR2_X1    g08641(.A1(new_n8292_), .A2(new_n8383_), .Z(new_n8706_));
  NAND2_X1   g08642(.A1(new_n8706_), .A2(new_n8457_), .ZN(new_n8707_));
  NOR2_X1    g08643(.A1(new_n8705_), .A2(new_n8707_), .ZN(new_n8708_));
  AND2_X2    g08644(.A1(new_n8705_), .A2(new_n8707_), .Z(new_n8709_));
  NOR2_X1    g08645(.A1(new_n8709_), .A2(new_n8708_), .ZN(new_n8710_));
  INV_X1     g08646(.I(new_n8710_), .ZN(new_n8711_));
  NOR2_X1    g08647(.A1(new_n8702_), .A2(new_n8711_), .ZN(new_n8712_));
  INV_X1     g08648(.I(new_n8712_), .ZN(new_n8713_));
  XOR2_X1    g08649(.A1(new_n8382_), .A2(new_n8457_), .Z(new_n8714_));
  NOR2_X1    g08650(.A1(new_n8472_), .A2(new_n8714_), .ZN(new_n8715_));
  XOR2_X1    g08651(.A1(new_n8382_), .A2(new_n8456_), .Z(new_n8716_));
  NOR2_X1    g08652(.A1(new_n8292_), .A2(new_n8716_), .ZN(new_n8717_));
  NOR2_X1    g08653(.A1(new_n8715_), .A2(new_n8717_), .ZN(new_n8718_));
  INV_X1     g08654(.I(new_n8718_), .ZN(new_n8719_));
  NOR2_X1    g08655(.A1(new_n8711_), .A2(new_n8719_), .ZN(new_n8720_));
  NAND2_X1   g08656(.A1(new_n8471_), .A2(new_n8288_), .ZN(new_n8721_));
  XOR2_X1    g08657(.A1(new_n8721_), .A2(new_n4094_), .Z(new_n8722_));
  AND2_X2    g08658(.A1(new_n8722_), .A2(new_n4172_), .Z(new_n8723_));
  NOR2_X1    g08659(.A1(new_n8722_), .A2(new_n4172_), .ZN(new_n8724_));
  NOR2_X1    g08660(.A1(new_n8723_), .A2(new_n8724_), .ZN(new_n8725_));
  INV_X1     g08661(.I(new_n8725_), .ZN(new_n8726_));
  NOR2_X1    g08662(.A1(new_n8726_), .A2(new_n8719_), .ZN(new_n8727_));
  INV_X1     g08663(.I(new_n8727_), .ZN(new_n8728_));
  NAND2_X1   g08664(.A1(new_n8469_), .A2(new_n8470_), .ZN(new_n8729_));
  XOR2_X1    g08665(.A1(new_n8729_), .A2(new_n8282_), .Z(new_n8730_));
  XOR2_X1    g08666(.A1(new_n8261_), .A2(new_n8274_), .Z(new_n8731_));
  NAND2_X1   g08667(.A1(new_n8731_), .A2(new_n8283_), .ZN(new_n8732_));
  NOR2_X1    g08668(.A1(new_n8730_), .A2(new_n8732_), .ZN(new_n8733_));
  AND2_X2    g08669(.A1(new_n8730_), .A2(new_n8732_), .Z(new_n8734_));
  NOR2_X1    g08670(.A1(new_n8734_), .A2(new_n8733_), .ZN(new_n8735_));
  INV_X1     g08671(.I(new_n8735_), .ZN(new_n8736_));
  NOR2_X1    g08672(.A1(new_n8726_), .A2(new_n8736_), .ZN(new_n8737_));
  NOR2_X1    g08673(.A1(new_n8466_), .A2(new_n8241_), .ZN(new_n8738_));
  XOR2_X1    g08674(.A1(new_n8738_), .A2(new_n8251_), .Z(new_n8739_));
  XOR2_X1    g08675(.A1(new_n8229_), .A2(new_n8242_), .Z(new_n8740_));
  NAND2_X1   g08676(.A1(new_n8740_), .A2(new_n8252_), .ZN(new_n8741_));
  NOR2_X1    g08677(.A1(new_n8739_), .A2(new_n8741_), .ZN(new_n8742_));
  NAND2_X1   g08678(.A1(new_n8739_), .A2(new_n8741_), .ZN(new_n8743_));
  INV_X1     g08679(.I(new_n8743_), .ZN(new_n8744_));
  NOR2_X1    g08680(.A1(new_n8744_), .A2(new_n8742_), .ZN(new_n8745_));
  INV_X1     g08681(.I(new_n8745_), .ZN(new_n8746_));
  NAND2_X1   g08682(.A1(new_n8256_), .A2(new_n8258_), .ZN(new_n8747_));
  XOR2_X1    g08683(.A1(new_n8747_), .A2(new_n4467_), .Z(new_n8748_));
  AND2_X2    g08684(.A1(new_n8748_), .A2(new_n4699_), .Z(new_n8749_));
  NOR2_X1    g08685(.A1(new_n8748_), .A2(new_n4699_), .ZN(new_n8750_));
  NOR2_X1    g08686(.A1(new_n8749_), .A2(new_n8750_), .ZN(new_n8751_));
  INV_X1     g08687(.I(new_n8751_), .ZN(new_n8752_));
  NOR2_X1    g08688(.A1(new_n8752_), .A2(new_n8746_), .ZN(new_n8753_));
  XOR2_X1    g08689(.A1(new_n8241_), .A2(new_n8252_), .Z(new_n8754_));
  NOR2_X1    g08690(.A1(new_n8754_), .A2(new_n8466_), .ZN(new_n8755_));
  XOR2_X1    g08691(.A1(new_n8241_), .A2(new_n8253_), .Z(new_n8756_));
  NOR2_X1    g08692(.A1(new_n8756_), .A2(new_n8229_), .ZN(new_n8757_));
  NOR2_X1    g08693(.A1(new_n8755_), .A2(new_n8757_), .ZN(new_n8758_));
  NAND2_X1   g08694(.A1(new_n8745_), .A2(new_n8758_), .ZN(new_n8759_));
  INV_X1     g08695(.I(new_n8759_), .ZN(new_n8760_));
  INV_X1     g08696(.I(new_n8758_), .ZN(new_n8761_));
  NAND2_X1   g08697(.A1(new_n8224_), .A2(new_n8226_), .ZN(new_n8762_));
  NAND2_X1   g08698(.A1(new_n8762_), .A2(new_n8227_), .ZN(new_n8763_));
  INV_X1     g08699(.I(new_n8763_), .ZN(new_n8764_));
  NOR2_X1    g08700(.A1(new_n8762_), .A2(new_n8227_), .ZN(new_n8765_));
  NOR2_X1    g08701(.A1(new_n8764_), .A2(new_n8765_), .ZN(new_n8766_));
  NOR2_X1    g08702(.A1(new_n8184_), .A2(new_n8185_), .ZN(new_n8767_));
  NAND2_X1   g08703(.A1(new_n8041_), .A2(new_n8109_), .ZN(new_n8768_));
  XOR2_X1    g08704(.A1(new_n8768_), .A2(new_n8767_), .Z(new_n8769_));
  XOR2_X1    g08705(.A1(new_n8041_), .A2(new_n8109_), .Z(new_n8770_));
  NAND2_X1   g08706(.A1(new_n8770_), .A2(new_n8174_), .ZN(new_n8771_));
  NOR2_X1    g08707(.A1(new_n8769_), .A2(new_n8771_), .ZN(new_n8772_));
  AND2_X2    g08708(.A1(new_n8769_), .A2(new_n8771_), .Z(new_n8773_));
  NOR2_X1    g08709(.A1(new_n8773_), .A2(new_n8772_), .ZN(new_n8774_));
  XOR2_X1    g08710(.A1(new_n7941_), .A2(new_n7652_), .Z(new_n8775_));
  NOR2_X1    g08711(.A1(new_n8775_), .A2(new_n7529_), .ZN(new_n8776_));
  AOI21_X1   g08712(.A1(new_n7946_), .A2(new_n7654_), .B(new_n7935_), .ZN(new_n8777_));
  NOR2_X1    g08713(.A1(new_n8776_), .A2(new_n8777_), .ZN(new_n8778_));
  INV_X1     g08714(.I(new_n8778_), .ZN(new_n8779_));
  NAND3_X1   g08715(.A1(new_n7930_), .A2(new_n7931_), .A3(new_n7526_), .ZN(new_n8780_));
  OAI21_X1   g08716(.A1(new_n7514_), .A2(new_n7521_), .B(new_n7932_), .ZN(new_n8781_));
  AOI21_X1   g08717(.A1(new_n8780_), .A2(new_n8781_), .B(new_n7929_), .ZN(new_n8782_));
  AOI21_X1   g08718(.A1(new_n7527_), .A2(new_n7934_), .B(new_n7378_), .ZN(new_n8783_));
  NOR2_X1    g08719(.A1(new_n8782_), .A2(new_n8783_), .ZN(new_n8784_));
  INV_X1     g08720(.I(new_n8784_), .ZN(new_n8785_));
  XOR2_X1    g08721(.A1(new_n6928_), .A2(new_n6949_), .Z(new_n8786_));
  NAND3_X1   g08722(.A1(new_n6901_), .A2(new_n6910_), .A3(new_n6942_), .ZN(new_n8787_));
  INV_X1     g08723(.I(new_n8787_), .ZN(new_n8788_));
  AOI21_X1   g08724(.A1(new_n6901_), .A2(new_n6910_), .B(new_n6942_), .ZN(new_n8789_));
  OAI21_X1   g08725(.A1(new_n8788_), .A2(new_n8789_), .B(new_n4387_), .ZN(new_n8790_));
  OAI21_X1   g08726(.A1(new_n6940_), .A2(new_n6941_), .B(new_n6917_), .ZN(new_n8791_));
  NAND3_X1   g08727(.A1(new_n8791_), .A2(new_n8787_), .A3(\a[2] ), .ZN(new_n8792_));
  NAND2_X1   g08728(.A1(new_n8790_), .A2(new_n8792_), .ZN(new_n8793_));
  NAND2_X1   g08729(.A1(new_n8793_), .A2(new_n6926_), .ZN(new_n8794_));
  INV_X1     g08730(.I(new_n6926_), .ZN(new_n8795_));
  NAND3_X1   g08731(.A1(new_n8790_), .A2(new_n8792_), .A3(new_n8795_), .ZN(new_n8796_));
  NAND2_X1   g08732(.A1(new_n8794_), .A2(new_n8796_), .ZN(new_n8797_));
  OAI22_X1   g08733(.A1(new_n2614_), .A2(new_n6839_), .B1(new_n529_), .B2(new_n6913_), .ZN(new_n8798_));
  INV_X1     g08734(.I(new_n6843_), .ZN(new_n8799_));
  NAND2_X1   g08735(.A1(new_n2718_), .A2(new_n8799_), .ZN(new_n8800_));
  AOI21_X1   g08736(.A1(new_n8800_), .A2(new_n8798_), .B(new_n6836_), .ZN(new_n8801_));
  NAND2_X1   g08737(.A1(new_n3074_), .A2(new_n8801_), .ZN(new_n8802_));
  XOR2_X1    g08738(.A1(new_n8802_), .A2(new_n65_), .Z(new_n8803_));
  NOR2_X1    g08739(.A1(new_n6216_), .A2(new_n6215_), .ZN(new_n8804_));
  INV_X1     g08740(.I(new_n8804_), .ZN(new_n8805_));
  XOR2_X1    g08741(.A1(new_n6817_), .A2(new_n6157_), .Z(new_n8806_));
  NOR2_X1    g08742(.A1(new_n8806_), .A2(new_n8805_), .ZN(new_n8807_));
  XOR2_X1    g08743(.A1(new_n6817_), .A2(new_n6158_), .Z(new_n8808_));
  NOR2_X1    g08744(.A1(new_n8808_), .A2(new_n8804_), .ZN(new_n8809_));
  NOR2_X1    g08745(.A1(new_n8809_), .A2(new_n8807_), .ZN(new_n8810_));
  XOR2_X1    g08746(.A1(new_n6816_), .A2(new_n6235_), .Z(new_n8811_));
  OAI22_X1   g08747(.A1(new_n813_), .A2(new_n6785_), .B1(new_n1008_), .B2(new_n6783_), .ZN(new_n8812_));
  NAND2_X1   g08748(.A1(new_n897_), .A2(new_n6789_), .ZN(new_n8813_));
  AOI21_X1   g08749(.A1(new_n8812_), .A2(new_n8813_), .B(new_n6776_), .ZN(new_n8814_));
  NAND2_X1   g08750(.A1(new_n2917_), .A2(new_n8814_), .ZN(new_n8815_));
  XOR2_X1    g08751(.A1(new_n8815_), .A2(\a[8] ), .Z(new_n8816_));
  INV_X1     g08752(.I(new_n8816_), .ZN(new_n8817_));
  NOR2_X1    g08753(.A1(new_n8811_), .A2(new_n8817_), .ZN(new_n8818_));
  XOR2_X1    g08754(.A1(new_n6495_), .A2(new_n6235_), .Z(new_n8819_));
  NOR2_X1    g08755(.A1(new_n8819_), .A2(new_n8816_), .ZN(new_n8820_));
  OAI22_X1   g08756(.A1(new_n896_), .A2(new_n6785_), .B1(new_n1180_), .B2(new_n6783_), .ZN(new_n8821_));
  NAND2_X1   g08757(.A1(new_n2504_), .A2(new_n6789_), .ZN(new_n8822_));
  AOI21_X1   g08758(.A1(new_n8822_), .A2(new_n8821_), .B(new_n6776_), .ZN(new_n8823_));
  NAND2_X1   g08759(.A1(new_n3596_), .A2(new_n8823_), .ZN(new_n8824_));
  XOR2_X1    g08760(.A1(new_n8824_), .A2(\a[8] ), .Z(new_n8825_));
  XOR2_X1    g08761(.A1(new_n6490_), .A2(new_n6494_), .Z(new_n8826_));
  NAND2_X1   g08762(.A1(new_n8826_), .A2(new_n8825_), .ZN(new_n8827_));
  INV_X1     g08763(.I(new_n8827_), .ZN(new_n8828_));
  NOR3_X1    g08764(.A1(new_n8818_), .A2(new_n8820_), .A3(new_n8828_), .ZN(new_n8829_));
  OAI22_X1   g08765(.A1(new_n2559_), .A2(new_n6785_), .B1(new_n896_), .B2(new_n6783_), .ZN(new_n8830_));
  NAND2_X1   g08766(.A1(new_n814_), .A2(new_n6789_), .ZN(new_n8831_));
  AOI21_X1   g08767(.A1(new_n8830_), .A2(new_n8831_), .B(new_n6776_), .ZN(new_n8832_));
  NAND2_X1   g08768(.A1(new_n3624_), .A2(new_n8832_), .ZN(new_n8833_));
  XOR2_X1    g08769(.A1(new_n8833_), .A2(\a[8] ), .Z(new_n8834_));
  INV_X1     g08770(.I(new_n8834_), .ZN(new_n8835_));
  NOR2_X1    g08771(.A1(new_n8829_), .A2(new_n8835_), .ZN(new_n8836_));
  NAND2_X1   g08772(.A1(new_n8819_), .A2(new_n8816_), .ZN(new_n8837_));
  NAND2_X1   g08773(.A1(new_n8811_), .A2(new_n8817_), .ZN(new_n8838_));
  NAND4_X1   g08774(.A1(new_n8838_), .A2(new_n8837_), .A3(new_n8827_), .A4(new_n8835_), .ZN(new_n8839_));
  INV_X1     g08775(.I(new_n8839_), .ZN(new_n8840_));
  OAI21_X1   g08776(.A1(new_n8836_), .A2(new_n8840_), .B(new_n8810_), .ZN(new_n8841_));
  XOR2_X1    g08777(.A1(new_n8808_), .A2(new_n8805_), .Z(new_n8842_));
  NAND3_X1   g08778(.A1(new_n8838_), .A2(new_n8837_), .A3(new_n8827_), .ZN(new_n8843_));
  NAND2_X1   g08779(.A1(new_n8843_), .A2(new_n8834_), .ZN(new_n8844_));
  NAND3_X1   g08780(.A1(new_n8842_), .A2(new_n8844_), .A3(new_n8839_), .ZN(new_n8845_));
  NAND3_X1   g08781(.A1(new_n8845_), .A2(new_n8841_), .A3(new_n8803_), .ZN(new_n8846_));
  XOR2_X1    g08782(.A1(new_n8802_), .A2(\a[5] ), .Z(new_n8847_));
  AOI21_X1   g08783(.A1(new_n8844_), .A2(new_n8839_), .B(new_n8842_), .ZN(new_n8848_));
  NOR3_X1    g08784(.A1(new_n8810_), .A2(new_n8836_), .A3(new_n8840_), .ZN(new_n8849_));
  OAI21_X1   g08785(.A1(new_n8848_), .A2(new_n8849_), .B(new_n8847_), .ZN(new_n8850_));
  INV_X1     g08786(.I(new_n8825_), .ZN(new_n8851_));
  XOR2_X1    g08787(.A1(new_n6815_), .A2(new_n6494_), .Z(new_n8852_));
  NAND2_X1   g08788(.A1(new_n8852_), .A2(new_n8851_), .ZN(new_n8853_));
  INV_X1     g08789(.I(new_n8853_), .ZN(new_n8854_));
  NAND3_X1   g08790(.A1(new_n8838_), .A2(new_n8837_), .A3(new_n8854_), .ZN(new_n8855_));
  OAI21_X1   g08791(.A1(new_n8818_), .A2(new_n8820_), .B(new_n8853_), .ZN(new_n8856_));
  OAI22_X1   g08792(.A1(new_n2559_), .A2(new_n6913_), .B1(new_n694_), .B2(new_n6839_), .ZN(new_n8857_));
  NAND2_X1   g08793(.A1(new_n2567_), .A2(new_n8799_), .ZN(new_n8858_));
  AOI21_X1   g08794(.A1(new_n8857_), .A2(new_n8858_), .B(new_n6836_), .ZN(new_n8859_));
  NAND2_X1   g08795(.A1(new_n2759_), .A2(new_n8859_), .ZN(new_n8860_));
  XOR2_X1    g08796(.A1(new_n8860_), .A2(\a[5] ), .Z(new_n8861_));
  NAND3_X1   g08797(.A1(new_n8856_), .A2(new_n8855_), .A3(new_n8861_), .ZN(new_n8862_));
  NOR3_X1    g08798(.A1(new_n8818_), .A2(new_n8820_), .A3(new_n8853_), .ZN(new_n8863_));
  AOI21_X1   g08799(.A1(new_n8838_), .A2(new_n8837_), .B(new_n8854_), .ZN(new_n8864_));
  XOR2_X1    g08800(.A1(new_n8860_), .A2(new_n65_), .Z(new_n8865_));
  OAI21_X1   g08801(.A1(new_n8864_), .A2(new_n8863_), .B(new_n8865_), .ZN(new_n8866_));
  NAND2_X1   g08802(.A1(new_n8827_), .A2(new_n8853_), .ZN(new_n8867_));
  OAI21_X1   g08803(.A1(new_n2559_), .A2(new_n6843_), .B(new_n6835_), .ZN(new_n8868_));
  OAI22_X1   g08804(.A1(new_n813_), .A2(new_n6913_), .B1(new_n529_), .B2(new_n6839_), .ZN(new_n8869_));
  NOR2_X1    g08805(.A1(new_n8868_), .A2(new_n8869_), .ZN(new_n8870_));
  NAND2_X1   g08806(.A1(new_n3051_), .A2(new_n8870_), .ZN(new_n8871_));
  XOR2_X1    g08807(.A1(new_n8871_), .A2(\a[5] ), .Z(new_n8872_));
  NOR2_X1    g08808(.A1(new_n8867_), .A2(new_n8872_), .ZN(new_n8873_));
  INV_X1     g08809(.I(new_n8873_), .ZN(new_n8874_));
  OAI22_X1   g08810(.A1(new_n2559_), .A2(new_n6839_), .B1(new_n896_), .B2(new_n6913_), .ZN(new_n8875_));
  NAND2_X1   g08811(.A1(new_n814_), .A2(new_n8799_), .ZN(new_n8876_));
  AOI21_X1   g08812(.A1(new_n8875_), .A2(new_n8876_), .B(new_n6836_), .ZN(new_n8877_));
  AND3_X2    g08813(.A1(new_n3624_), .A2(new_n65_), .A3(new_n8877_), .Z(new_n8878_));
  AOI21_X1   g08814(.A1(new_n3624_), .A2(new_n8877_), .B(new_n65_), .ZN(new_n8879_));
  NOR2_X1    g08815(.A1(new_n8878_), .A2(new_n8879_), .ZN(new_n8880_));
  INV_X1     g08816(.I(new_n8880_), .ZN(new_n8881_));
  NAND2_X1   g08817(.A1(new_n6468_), .A2(new_n6469_), .ZN(new_n8882_));
  XOR2_X1    g08818(.A1(new_n6489_), .A2(new_n6246_), .Z(new_n8883_));
  XOR2_X1    g08819(.A1(new_n8883_), .A2(new_n8882_), .Z(new_n8884_));
  NAND3_X1   g08820(.A1(new_n6475_), .A2(new_n6477_), .A3(new_n6476_), .ZN(new_n8885_));
  INV_X1     g08821(.I(new_n8885_), .ZN(new_n8886_));
  AOI21_X1   g08822(.A1(new_n6476_), .A2(new_n6477_), .B(new_n6475_), .ZN(new_n8887_));
  NOR3_X1    g08823(.A1(new_n8886_), .A2(new_n6813_), .A3(new_n8887_), .ZN(new_n8888_));
  INV_X1     g08824(.I(new_n8887_), .ZN(new_n8889_));
  AOI21_X1   g08825(.A1(new_n8889_), .A2(new_n8885_), .B(new_n6488_), .ZN(new_n8890_));
  OAI22_X1   g08826(.A1(new_n1180_), .A2(new_n6785_), .B1(new_n2492_), .B2(new_n6783_), .ZN(new_n8891_));
  NAND2_X1   g08827(.A1(new_n1122_), .A2(new_n6789_), .ZN(new_n8892_));
  AOI21_X1   g08828(.A1(new_n8892_), .A2(new_n8891_), .B(new_n6776_), .ZN(new_n8893_));
  AND3_X2    g08829(.A1(new_n3330_), .A2(new_n4009_), .A3(new_n8893_), .Z(new_n8894_));
  AOI21_X1   g08830(.A1(new_n3330_), .A2(new_n8893_), .B(new_n4009_), .ZN(new_n8895_));
  NOR2_X1    g08831(.A1(new_n8894_), .A2(new_n8895_), .ZN(new_n8896_));
  OAI21_X1   g08832(.A1(new_n8890_), .A2(new_n8888_), .B(new_n8896_), .ZN(new_n8897_));
  NOR3_X1    g08833(.A1(new_n8890_), .A2(new_n8888_), .A3(new_n8896_), .ZN(new_n8898_));
  INV_X1     g08834(.I(new_n8898_), .ZN(new_n8899_));
  NAND2_X1   g08835(.A1(new_n6487_), .A2(new_n6485_), .ZN(new_n8900_));
  NAND2_X1   g08836(.A1(new_n6813_), .A2(new_n8900_), .ZN(new_n8901_));
  OAI21_X1   g08837(.A1(new_n2492_), .A2(new_n6788_), .B(new_n6775_), .ZN(new_n8902_));
  OAI22_X1   g08838(.A1(new_n1121_), .A2(new_n6785_), .B1(new_n2451_), .B2(new_n6783_), .ZN(new_n8903_));
  NOR2_X1    g08839(.A1(new_n8903_), .A2(new_n8902_), .ZN(new_n8904_));
  NAND2_X1   g08840(.A1(new_n3393_), .A2(new_n8904_), .ZN(new_n8905_));
  INV_X1     g08841(.I(new_n8905_), .ZN(new_n8906_));
  NOR2_X1    g08842(.A1(new_n8906_), .A2(new_n4009_), .ZN(new_n8907_));
  NOR2_X1    g08843(.A1(new_n8905_), .A2(\a[8] ), .ZN(new_n8908_));
  NOR2_X1    g08844(.A1(new_n8907_), .A2(new_n8908_), .ZN(new_n8909_));
  NOR2_X1    g08845(.A1(new_n6812_), .A2(new_n6811_), .ZN(new_n8910_));
  OAI21_X1   g08846(.A1(new_n8910_), .A2(new_n6488_), .B(new_n4009_), .ZN(new_n8911_));
  NAND3_X1   g08847(.A1(new_n6813_), .A2(new_n8900_), .A3(\a[8] ), .ZN(new_n8912_));
  AOI21_X1   g08848(.A1(new_n8911_), .A2(new_n8912_), .B(new_n8906_), .ZN(new_n8913_));
  AOI21_X1   g08849(.A1(new_n6813_), .A2(new_n8900_), .B(\a[8] ), .ZN(new_n8914_));
  NOR3_X1    g08850(.A1(new_n8910_), .A2(new_n6488_), .A3(new_n4009_), .ZN(new_n8915_));
  NOR3_X1    g08851(.A1(new_n8914_), .A2(new_n8915_), .A3(new_n8905_), .ZN(new_n8916_));
  OAI22_X1   g08852(.A1(new_n8916_), .A2(new_n8913_), .B1(new_n8901_), .B2(new_n8909_), .ZN(new_n8917_));
  NAND3_X1   g08853(.A1(new_n8899_), .A2(new_n8917_), .A3(new_n8897_), .ZN(new_n8918_));
  OAI22_X1   g08854(.A1(new_n1008_), .A2(new_n6785_), .B1(new_n1121_), .B2(new_n6783_), .ZN(new_n8919_));
  NAND2_X1   g08855(.A1(new_n1181_), .A2(new_n6789_), .ZN(new_n8920_));
  AOI21_X1   g08856(.A1(new_n8919_), .A2(new_n8920_), .B(new_n6776_), .ZN(new_n8921_));
  NAND2_X1   g08857(.A1(new_n3562_), .A2(new_n8921_), .ZN(new_n8922_));
  XOR2_X1    g08858(.A1(new_n8922_), .A2(\a[8] ), .Z(new_n8923_));
  NAND2_X1   g08859(.A1(new_n8918_), .A2(new_n8923_), .ZN(new_n8924_));
  INV_X1     g08860(.I(new_n8923_), .ZN(new_n8925_));
  NAND4_X1   g08861(.A1(new_n8925_), .A2(new_n8899_), .A3(new_n8917_), .A4(new_n8897_), .ZN(new_n8926_));
  AOI21_X1   g08862(.A1(new_n8924_), .A2(new_n8926_), .B(new_n8884_), .ZN(new_n8927_));
  XNOR2_X1   g08863(.A1(new_n8883_), .A2(new_n8882_), .ZN(new_n8928_));
  INV_X1     g08864(.I(new_n8897_), .ZN(new_n8929_));
  NOR2_X1    g08865(.A1(new_n8909_), .A2(new_n8901_), .ZN(new_n8930_));
  INV_X1     g08866(.I(new_n8913_), .ZN(new_n8931_));
  NAND3_X1   g08867(.A1(new_n8911_), .A2(new_n8912_), .A3(new_n8906_), .ZN(new_n8932_));
  AOI21_X1   g08868(.A1(new_n8931_), .A2(new_n8932_), .B(new_n8930_), .ZN(new_n8933_));
  NOR3_X1    g08869(.A1(new_n8933_), .A2(new_n8929_), .A3(new_n8898_), .ZN(new_n8934_));
  NOR2_X1    g08870(.A1(new_n8934_), .A2(new_n8925_), .ZN(new_n8935_));
  NOR2_X1    g08871(.A1(new_n8918_), .A2(new_n8923_), .ZN(new_n8936_));
  NOR3_X1    g08872(.A1(new_n8935_), .A2(new_n8936_), .A3(new_n8928_), .ZN(new_n8937_));
  NOR2_X1    g08873(.A1(new_n8937_), .A2(new_n8927_), .ZN(new_n8938_));
  NOR2_X1    g08874(.A1(new_n8938_), .A2(new_n8881_), .ZN(new_n8939_));
  INV_X1     g08875(.I(new_n8939_), .ZN(new_n8940_));
  OAI22_X1   g08876(.A1(new_n813_), .A2(new_n6839_), .B1(new_n1008_), .B2(new_n6913_), .ZN(new_n8941_));
  NAND2_X1   g08877(.A1(new_n897_), .A2(new_n8799_), .ZN(new_n8942_));
  AOI21_X1   g08878(.A1(new_n8941_), .A2(new_n8942_), .B(new_n6836_), .ZN(new_n8943_));
  AND3_X2    g08879(.A1(new_n2917_), .A2(new_n65_), .A3(new_n8943_), .Z(new_n8944_));
  AOI21_X1   g08880(.A1(new_n2917_), .A2(new_n8943_), .B(new_n65_), .ZN(new_n8945_));
  NOR2_X1    g08881(.A1(new_n8944_), .A2(new_n8945_), .ZN(new_n8946_));
  INV_X1     g08882(.I(new_n8946_), .ZN(new_n8947_));
  NAND3_X1   g08883(.A1(new_n8933_), .A2(new_n8899_), .A3(new_n8897_), .ZN(new_n8948_));
  OAI21_X1   g08884(.A1(new_n8929_), .A2(new_n8898_), .B(new_n8917_), .ZN(new_n8949_));
  NAND2_X1   g08885(.A1(new_n8948_), .A2(new_n8949_), .ZN(new_n8950_));
  NOR2_X1    g08886(.A1(new_n8947_), .A2(new_n8950_), .ZN(new_n8951_));
  NOR3_X1    g08887(.A1(new_n8929_), .A2(new_n8898_), .A3(new_n8917_), .ZN(new_n8952_));
  AOI21_X1   g08888(.A1(new_n8899_), .A2(new_n8897_), .B(new_n8933_), .ZN(new_n8953_));
  NOR2_X1    g08889(.A1(new_n8953_), .A2(new_n8952_), .ZN(new_n8954_));
  NOR2_X1    g08890(.A1(new_n8954_), .A2(new_n8946_), .ZN(new_n8955_));
  INV_X1     g08891(.I(new_n5782_), .ZN(new_n8956_));
  OAI22_X1   g08892(.A1(new_n1729_), .A2(new_n4470_), .B1(new_n4745_), .B2(new_n4291_), .ZN(new_n8957_));
  NAND2_X1   g08893(.A1(new_n1862_), .A2(new_n4298_), .ZN(new_n8958_));
  AOI21_X1   g08894(.A1(new_n8957_), .A2(new_n8958_), .B(new_n4468_), .ZN(new_n8959_));
  NAND2_X1   g08895(.A1(new_n4842_), .A2(new_n8959_), .ZN(new_n8960_));
  XOR2_X1    g08896(.A1(new_n8960_), .A2(new_n3372_), .Z(new_n8961_));
  NAND2_X1   g08897(.A1(new_n8961_), .A2(new_n8956_), .ZN(new_n8962_));
  AOI22_X1   g08898(.A1(new_n4766_), .A2(new_n4292_), .B1(new_n1813_), .B2(new_n4298_), .ZN(new_n8963_));
  AOI21_X1   g08899(.A1(new_n1862_), .A2(new_n4469_), .B(new_n8963_), .ZN(new_n8964_));
  NOR3_X1    g08900(.A1(new_n8964_), .A2(new_n4878_), .A3(new_n4468_), .ZN(new_n8965_));
  XOR2_X1    g08901(.A1(new_n8965_), .A2(\a[17] ), .Z(new_n8966_));
  NAND2_X1   g08902(.A1(new_n1813_), .A2(new_n4469_), .ZN(new_n8967_));
  NAND2_X1   g08903(.A1(new_n4766_), .A2(new_n4298_), .ZN(new_n8968_));
  NAND4_X1   g08904(.A1(new_n4981_), .A2(new_n4295_), .A3(new_n8967_), .A4(new_n8968_), .ZN(new_n8969_));
  XOR2_X1    g08905(.A1(new_n8969_), .A2(\a[17] ), .Z(new_n8970_));
  NOR2_X1    g08906(.A1(new_n1999_), .A2(new_n4284_), .ZN(new_n8971_));
  NOR2_X1    g08907(.A1(new_n8971_), .A2(new_n3372_), .ZN(new_n8972_));
  NAND2_X1   g08908(.A1(new_n8970_), .A2(new_n8972_), .ZN(new_n8973_));
  NOR2_X1    g08909(.A1(new_n8973_), .A2(new_n8966_), .ZN(new_n8974_));
  NOR2_X1    g08910(.A1(new_n8961_), .A2(new_n8956_), .ZN(new_n8975_));
  OAI21_X1   g08911(.A1(new_n8974_), .A2(new_n8975_), .B(new_n8962_), .ZN(new_n8976_));
  XOR2_X1    g08912(.A1(new_n5781_), .A2(new_n5783_), .Z(new_n8977_));
  OAI22_X1   g08913(.A1(new_n1764_), .A2(new_n4470_), .B1(new_n1729_), .B2(new_n4297_), .ZN(new_n8978_));
  NAND2_X1   g08914(.A1(new_n1862_), .A2(new_n4292_), .ZN(new_n8979_));
  AOI21_X1   g08915(.A1(new_n8978_), .A2(new_n8979_), .B(new_n4468_), .ZN(new_n8980_));
  NAND2_X1   g08916(.A1(new_n4810_), .A2(new_n8980_), .ZN(new_n8981_));
  XOR2_X1    g08917(.A1(new_n8981_), .A2(\a[17] ), .Z(new_n8982_));
  NAND2_X1   g08918(.A1(new_n8982_), .A2(new_n8977_), .ZN(new_n8983_));
  NAND2_X1   g08919(.A1(new_n8976_), .A2(new_n8983_), .ZN(new_n8984_));
  OR2_X2     g08920(.A1(new_n8982_), .A2(new_n8977_), .Z(new_n8985_));
  NAND2_X1   g08921(.A1(new_n8984_), .A2(new_n8985_), .ZN(new_n8986_));
  OAI22_X1   g08922(.A1(new_n1764_), .A2(new_n4297_), .B1(new_n1729_), .B2(new_n4291_), .ZN(new_n8987_));
  NAND2_X1   g08923(.A1(new_n1613_), .A2(new_n4469_), .ZN(new_n8988_));
  AOI21_X1   g08924(.A1(new_n8988_), .A2(new_n8987_), .B(new_n4468_), .ZN(new_n8989_));
  NAND2_X1   g08925(.A1(new_n4778_), .A2(new_n8989_), .ZN(new_n8990_));
  XOR2_X1    g08926(.A1(new_n8990_), .A2(new_n3372_), .Z(new_n8991_));
  NAND2_X1   g08927(.A1(new_n5781_), .A2(new_n5783_), .ZN(new_n8992_));
  XOR2_X1    g08928(.A1(new_n8992_), .A2(new_n5777_), .Z(new_n8993_));
  NOR2_X1    g08929(.A1(new_n8991_), .A2(new_n8993_), .ZN(new_n8994_));
  XOR2_X1    g08930(.A1(new_n8990_), .A2(\a[17] ), .Z(new_n8995_));
  INV_X1     g08931(.I(new_n8993_), .ZN(new_n8996_));
  NOR2_X1    g08932(.A1(new_n8996_), .A2(new_n8995_), .ZN(new_n8997_));
  NOR2_X1    g08933(.A1(new_n8997_), .A2(new_n8994_), .ZN(new_n8998_));
  XOR2_X1    g08934(.A1(new_n8998_), .A2(new_n8986_), .Z(new_n8999_));
  OAI22_X1   g08935(.A1(new_n2103_), .A2(new_n6091_), .B1(new_n1678_), .B2(new_n6089_), .ZN(new_n9000_));
  NAND2_X1   g08936(.A1(new_n2107_), .A2(new_n6095_), .ZN(new_n9001_));
  AOI21_X1   g08937(.A1(new_n9000_), .A2(new_n9001_), .B(new_n6082_), .ZN(new_n9002_));
  NAND2_X1   g08938(.A1(new_n4545_), .A2(new_n9002_), .ZN(new_n9003_));
  XOR2_X1    g08939(.A1(new_n9003_), .A2(new_n3521_), .Z(new_n9004_));
  XNOR2_X1   g08940(.A1(new_n8999_), .A2(new_n9004_), .ZN(new_n9005_));
  OAI22_X1   g08941(.A1(new_n2158_), .A2(new_n4716_), .B1(new_n2198_), .B2(new_n4719_), .ZN(new_n9006_));
  OAI21_X1   g08942(.A1(new_n1503_), .A2(new_n4710_), .B(new_n9006_), .ZN(new_n9007_));
  AOI21_X1   g08943(.A1(new_n4620_), .A2(new_n4706_), .B(new_n9007_), .ZN(new_n9008_));
  XOR2_X1    g08944(.A1(new_n9008_), .A2(new_n4034_), .Z(new_n9009_));
  OAI22_X1   g08945(.A1(new_n4365_), .A2(new_n4710_), .B1(new_n2198_), .B2(new_n4716_), .ZN(new_n9010_));
  NAND2_X1   g08946(.A1(new_n1504_), .A2(new_n4720_), .ZN(new_n9011_));
  AOI21_X1   g08947(.A1(new_n9010_), .A2(new_n9011_), .B(new_n4707_), .ZN(new_n9012_));
  NAND3_X1   g08948(.A1(new_n4363_), .A2(new_n4034_), .A3(new_n9012_), .ZN(new_n9013_));
  NAND2_X1   g08949(.A1(new_n4363_), .A2(new_n9012_), .ZN(new_n9014_));
  NAND2_X1   g08950(.A1(new_n9014_), .A2(\a[11] ), .ZN(new_n9015_));
  NAND2_X1   g08951(.A1(new_n9015_), .A2(new_n9013_), .ZN(new_n9016_));
  NAND2_X1   g08952(.A1(new_n8999_), .A2(new_n9004_), .ZN(new_n9017_));
  XOR2_X1    g08953(.A1(new_n5785_), .A2(new_n5767_), .Z(new_n9018_));
  NOR2_X1    g08954(.A1(new_n5772_), .A2(new_n5767_), .ZN(new_n9019_));
  OAI21_X1   g08955(.A1(new_n5902_), .A2(new_n9019_), .B(new_n5784_), .ZN(new_n9020_));
  OAI21_X1   g08956(.A1(new_n9018_), .A2(new_n5784_), .B(new_n9020_), .ZN(new_n9021_));
  OAI22_X1   g08957(.A1(new_n1678_), .A2(new_n4470_), .B1(new_n1764_), .B2(new_n4291_), .ZN(new_n9022_));
  NAND2_X1   g08958(.A1(new_n1613_), .A2(new_n4298_), .ZN(new_n9023_));
  AOI21_X1   g08959(.A1(new_n9022_), .A2(new_n9023_), .B(new_n4468_), .ZN(new_n9024_));
  NAND2_X1   g08960(.A1(new_n4917_), .A2(new_n9024_), .ZN(new_n9025_));
  XOR2_X1    g08961(.A1(new_n9025_), .A2(new_n3372_), .Z(new_n9026_));
  XNOR2_X1   g08962(.A1(new_n9021_), .A2(new_n9026_), .ZN(new_n9027_));
  INV_X1     g08963(.I(new_n8994_), .ZN(new_n9028_));
  OAI21_X1   g08964(.A1(new_n8986_), .A2(new_n8997_), .B(new_n9028_), .ZN(new_n9029_));
  INV_X1     g08965(.I(new_n9029_), .ZN(new_n9030_));
  NAND2_X1   g08966(.A1(new_n9027_), .A2(new_n9030_), .ZN(new_n9031_));
  XOR2_X1    g08967(.A1(new_n9021_), .A2(new_n9026_), .Z(new_n9032_));
  NAND2_X1   g08968(.A1(new_n9032_), .A2(new_n9029_), .ZN(new_n9033_));
  OAI22_X1   g08969(.A1(new_n2103_), .A2(new_n6094_), .B1(new_n2158_), .B2(new_n6091_), .ZN(new_n9034_));
  NAND2_X1   g08970(.A1(new_n2107_), .A2(new_n6180_), .ZN(new_n9035_));
  AOI21_X1   g08971(.A1(new_n9034_), .A2(new_n9035_), .B(new_n6082_), .ZN(new_n9036_));
  NAND2_X1   g08972(.A1(new_n4959_), .A2(new_n9036_), .ZN(new_n9037_));
  XOR2_X1    g08973(.A1(new_n9037_), .A2(new_n3521_), .Z(new_n9038_));
  NAND3_X1   g08974(.A1(new_n9038_), .A2(new_n9031_), .A3(new_n9033_), .ZN(new_n9039_));
  NOR2_X1    g08975(.A1(new_n9032_), .A2(new_n9029_), .ZN(new_n9040_));
  NOR2_X1    g08976(.A1(new_n9027_), .A2(new_n9030_), .ZN(new_n9041_));
  XOR2_X1    g08977(.A1(new_n9037_), .A2(\a[14] ), .Z(new_n9042_));
  OAI21_X1   g08978(.A1(new_n9040_), .A2(new_n9041_), .B(new_n9042_), .ZN(new_n9043_));
  NAND3_X1   g08979(.A1(new_n9043_), .A2(new_n9039_), .A3(new_n9017_), .ZN(new_n9044_));
  INV_X1     g08980(.I(new_n9017_), .ZN(new_n9045_));
  NOR3_X1    g08981(.A1(new_n9042_), .A2(new_n9041_), .A3(new_n9040_), .ZN(new_n9046_));
  AOI21_X1   g08982(.A1(new_n9031_), .A2(new_n9033_), .B(new_n9038_), .ZN(new_n9047_));
  OAI21_X1   g08983(.A1(new_n9047_), .A2(new_n9046_), .B(new_n9045_), .ZN(new_n9048_));
  NAND2_X1   g08984(.A1(new_n9048_), .A2(new_n9044_), .ZN(new_n9049_));
  NOR2_X1    g08985(.A1(new_n9049_), .A2(new_n9016_), .ZN(new_n9050_));
  NOR3_X1    g08986(.A1(new_n9050_), .A2(new_n9005_), .A3(new_n9009_), .ZN(new_n9051_));
  AOI22_X1   g08987(.A1(new_n9048_), .A2(new_n9044_), .B1(new_n9015_), .B2(new_n9013_), .ZN(new_n9052_));
  XOR2_X1    g08988(.A1(new_n5794_), .A2(new_n5904_), .Z(new_n9053_));
  NOR2_X1    g08989(.A1(new_n9053_), .A2(new_n5903_), .ZN(new_n9054_));
  AOI21_X1   g08990(.A1(new_n5795_), .A2(new_n5907_), .B(new_n5788_), .ZN(new_n9055_));
  NOR2_X1    g08991(.A1(new_n9054_), .A2(new_n9055_), .ZN(new_n9056_));
  INV_X1     g08992(.I(new_n9056_), .ZN(new_n9057_));
  NOR2_X1    g08993(.A1(new_n9021_), .A2(new_n9026_), .ZN(new_n9058_));
  OAI22_X1   g08994(.A1(new_n1678_), .A2(new_n4297_), .B1(new_n2071_), .B2(new_n4470_), .ZN(new_n9059_));
  NAND2_X1   g08995(.A1(new_n1613_), .A2(new_n4292_), .ZN(new_n9060_));
  AOI21_X1   g08996(.A1(new_n9059_), .A2(new_n9060_), .B(new_n4468_), .ZN(new_n9061_));
  NAND2_X1   g08997(.A1(new_n5070_), .A2(new_n9061_), .ZN(new_n9062_));
  XOR2_X1    g08998(.A1(new_n9062_), .A2(\a[17] ), .Z(new_n9063_));
  OAI21_X1   g08999(.A1(new_n9040_), .A2(new_n9058_), .B(new_n9063_), .ZN(new_n9064_));
  INV_X1     g09000(.I(new_n9058_), .ZN(new_n9065_));
  INV_X1     g09001(.I(new_n9063_), .ZN(new_n9066_));
  NAND3_X1   g09002(.A1(new_n9031_), .A2(new_n9065_), .A3(new_n9066_), .ZN(new_n9067_));
  AOI21_X1   g09003(.A1(new_n9067_), .A2(new_n9064_), .B(new_n9057_), .ZN(new_n9068_));
  AOI21_X1   g09004(.A1(new_n9031_), .A2(new_n9065_), .B(new_n9066_), .ZN(new_n9069_));
  NOR3_X1    g09005(.A1(new_n9040_), .A2(new_n9058_), .A3(new_n9063_), .ZN(new_n9070_));
  NOR3_X1    g09006(.A1(new_n9069_), .A2(new_n9070_), .A3(new_n9056_), .ZN(new_n9071_));
  OR2_X2     g09007(.A1(new_n9071_), .A2(new_n9068_), .Z(new_n9072_));
  NOR3_X1    g09008(.A1(new_n9047_), .A2(new_n9046_), .A3(new_n9045_), .ZN(new_n9073_));
  OAI22_X1   g09009(.A1(new_n2103_), .A2(new_n6089_), .B1(new_n2198_), .B2(new_n6091_), .ZN(new_n9074_));
  NAND2_X1   g09010(.A1(new_n2161_), .A2(new_n6095_), .ZN(new_n9075_));
  AOI21_X1   g09011(.A1(new_n9074_), .A2(new_n9075_), .B(new_n6082_), .ZN(new_n9076_));
  NAND2_X1   g09012(.A1(new_n5351_), .A2(new_n9076_), .ZN(new_n9077_));
  XOR2_X1    g09013(.A1(new_n9077_), .A2(\a[14] ), .Z(new_n9078_));
  OAI21_X1   g09014(.A1(new_n9073_), .A2(new_n9047_), .B(new_n9078_), .ZN(new_n9079_));
  INV_X1     g09015(.I(new_n9078_), .ZN(new_n9080_));
  NAND3_X1   g09016(.A1(new_n9044_), .A2(new_n9043_), .A3(new_n9080_), .ZN(new_n9081_));
  AOI21_X1   g09017(.A1(new_n9079_), .A2(new_n9081_), .B(new_n9072_), .ZN(new_n9082_));
  NOR2_X1    g09018(.A1(new_n9071_), .A2(new_n9068_), .ZN(new_n9083_));
  AOI21_X1   g09019(.A1(new_n9044_), .A2(new_n9043_), .B(new_n9080_), .ZN(new_n9084_));
  NOR3_X1    g09020(.A1(new_n9073_), .A2(new_n9047_), .A3(new_n9078_), .ZN(new_n9085_));
  NOR3_X1    g09021(.A1(new_n9085_), .A2(new_n9084_), .A3(new_n9083_), .ZN(new_n9086_));
  NOR2_X1    g09022(.A1(new_n9082_), .A2(new_n9086_), .ZN(new_n9087_));
  OAI22_X1   g09023(.A1(new_n2251_), .A2(new_n4710_), .B1(new_n4365_), .B2(new_n4719_), .ZN(new_n9088_));
  NAND2_X1   g09024(.A1(new_n1504_), .A2(new_n6480_), .ZN(new_n9089_));
  AOI21_X1   g09025(.A1(new_n9088_), .A2(new_n9089_), .B(new_n4707_), .ZN(new_n9090_));
  NAND2_X1   g09026(.A1(new_n4650_), .A2(new_n9090_), .ZN(new_n9091_));
  XOR2_X1    g09027(.A1(new_n9091_), .A2(new_n4034_), .Z(new_n9092_));
  OAI22_X1   g09028(.A1(new_n9087_), .A2(new_n9092_), .B1(new_n9051_), .B2(new_n9052_), .ZN(new_n9093_));
  NAND2_X1   g09029(.A1(new_n9087_), .A2(new_n9092_), .ZN(new_n9094_));
  XNOR2_X1   g09030(.A1(new_n6307_), .A2(new_n6303_), .ZN(new_n9095_));
  INV_X1     g09031(.I(new_n9095_), .ZN(new_n9096_));
  OAI22_X1   g09032(.A1(new_n2311_), .A2(new_n4710_), .B1(new_n4365_), .B2(new_n4716_), .ZN(new_n9097_));
  NAND2_X1   g09033(.A1(new_n2255_), .A2(new_n4720_), .ZN(new_n9098_));
  AOI21_X1   g09034(.A1(new_n9097_), .A2(new_n9098_), .B(new_n4707_), .ZN(new_n9099_));
  NAND3_X1   g09035(.A1(new_n4419_), .A2(new_n4034_), .A3(new_n9099_), .ZN(new_n9100_));
  INV_X1     g09036(.I(new_n9100_), .ZN(new_n9101_));
  AOI21_X1   g09037(.A1(new_n4419_), .A2(new_n9099_), .B(new_n4034_), .ZN(new_n9102_));
  NOR2_X1    g09038(.A1(new_n9101_), .A2(new_n9102_), .ZN(new_n9103_));
  NAND2_X1   g09039(.A1(new_n9096_), .A2(new_n9103_), .ZN(new_n9104_));
  INV_X1     g09040(.I(new_n9102_), .ZN(new_n9105_));
  NAND2_X1   g09041(.A1(new_n9105_), .A2(new_n9100_), .ZN(new_n9106_));
  NAND2_X1   g09042(.A1(new_n9106_), .A2(new_n9095_), .ZN(new_n9107_));
  AOI22_X1   g09043(.A1(new_n9093_), .A2(new_n9094_), .B1(new_n9104_), .B2(new_n9107_), .ZN(new_n9108_));
  NOR2_X1    g09044(.A1(new_n9009_), .A2(new_n9005_), .ZN(new_n9109_));
  XOR2_X1    g09045(.A1(new_n9014_), .A2(\a[11] ), .Z(new_n9110_));
  NAND3_X1   g09046(.A1(new_n9110_), .A2(new_n9044_), .A3(new_n9048_), .ZN(new_n9111_));
  AOI21_X1   g09047(.A1(new_n9111_), .A2(new_n9109_), .B(new_n9052_), .ZN(new_n9112_));
  OAI21_X1   g09048(.A1(new_n9085_), .A2(new_n9084_), .B(new_n9083_), .ZN(new_n9113_));
  NAND3_X1   g09049(.A1(new_n9072_), .A2(new_n9079_), .A3(new_n9081_), .ZN(new_n9114_));
  NAND2_X1   g09050(.A1(new_n9114_), .A2(new_n9113_), .ZN(new_n9115_));
  XOR2_X1    g09051(.A1(new_n9091_), .A2(\a[11] ), .Z(new_n9116_));
  AOI21_X1   g09052(.A1(new_n9115_), .A2(new_n9116_), .B(new_n9112_), .ZN(new_n9117_));
  NOR2_X1    g09053(.A1(new_n9115_), .A2(new_n9116_), .ZN(new_n9118_));
  XOR2_X1    g09054(.A1(new_n9103_), .A2(new_n9095_), .Z(new_n9119_));
  NOR3_X1    g09055(.A1(new_n9119_), .A2(new_n9117_), .A3(new_n9118_), .ZN(new_n9120_));
  NOR2_X1    g09056(.A1(new_n9120_), .A2(new_n9108_), .ZN(new_n9121_));
  NAND2_X1   g09057(.A1(new_n2359_), .A2(new_n6789_), .ZN(new_n9122_));
  NAND2_X1   g09058(.A1(new_n1408_), .A2(new_n6784_), .ZN(new_n9123_));
  AOI21_X1   g09059(.A1(new_n2354_), .A2(new_n7530_), .B(new_n6776_), .ZN(new_n9124_));
  NAND4_X1   g09060(.A1(new_n3904_), .A2(new_n9122_), .A3(new_n9123_), .A4(new_n9124_), .ZN(new_n9125_));
  XOR2_X1    g09061(.A1(new_n9125_), .A2(new_n4009_), .Z(new_n9126_));
  INV_X1     g09062(.I(new_n9126_), .ZN(new_n9127_));
  NOR2_X1    g09063(.A1(new_n9127_), .A2(new_n9121_), .ZN(new_n9128_));
  INV_X1     g09064(.I(new_n9107_), .ZN(new_n9129_));
  AOI22_X1   g09065(.A1(new_n9093_), .A2(new_n9094_), .B1(new_n9096_), .B2(new_n9103_), .ZN(new_n9130_));
  NAND3_X1   g09066(.A1(new_n6435_), .A2(new_n6334_), .A3(new_n6338_), .ZN(new_n9131_));
  NAND2_X1   g09067(.A1(new_n6436_), .A2(new_n6315_), .ZN(new_n9132_));
  AOI21_X1   g09068(.A1(new_n9131_), .A2(new_n9132_), .B(new_n6434_), .ZN(new_n9133_));
  AOI21_X1   g09069(.A1(new_n6438_), .A2(new_n6339_), .B(new_n6308_), .ZN(new_n9134_));
  NOR2_X1    g09070(.A1(new_n9133_), .A2(new_n9134_), .ZN(new_n9135_));
  OAI22_X1   g09071(.A1(new_n2251_), .A2(new_n4716_), .B1(new_n2351_), .B2(new_n4710_), .ZN(new_n9136_));
  NAND2_X1   g09072(.A1(new_n2310_), .A2(new_n4720_), .ZN(new_n9137_));
  AOI21_X1   g09073(.A1(new_n9137_), .A2(new_n9136_), .B(new_n4707_), .ZN(new_n9138_));
  NAND3_X1   g09074(.A1(new_n3914_), .A2(new_n4034_), .A3(new_n9138_), .ZN(new_n9139_));
  AOI21_X1   g09075(.A1(new_n3914_), .A2(new_n9138_), .B(new_n4034_), .ZN(new_n9140_));
  INV_X1     g09076(.I(new_n9140_), .ZN(new_n9141_));
  NAND2_X1   g09077(.A1(new_n9141_), .A2(new_n9139_), .ZN(new_n9142_));
  NOR2_X1    g09078(.A1(new_n9142_), .A2(new_n9135_), .ZN(new_n9143_));
  NAND2_X1   g09079(.A1(new_n9131_), .A2(new_n9132_), .ZN(new_n9144_));
  NAND2_X1   g09080(.A1(new_n9144_), .A2(new_n6308_), .ZN(new_n9145_));
  OAI21_X1   g09081(.A1(new_n6437_), .A2(new_n6341_), .B(new_n6434_), .ZN(new_n9146_));
  NAND2_X1   g09082(.A1(new_n9145_), .A2(new_n9146_), .ZN(new_n9147_));
  INV_X1     g09083(.I(new_n9139_), .ZN(new_n9148_));
  NOR2_X1    g09084(.A1(new_n9148_), .A2(new_n9140_), .ZN(new_n9149_));
  NOR2_X1    g09085(.A1(new_n9147_), .A2(new_n9149_), .ZN(new_n9150_));
  OAI22_X1   g09086(.A1(new_n9130_), .A2(new_n9129_), .B1(new_n9143_), .B2(new_n9150_), .ZN(new_n9151_));
  OAI21_X1   g09087(.A1(new_n9117_), .A2(new_n9118_), .B(new_n9104_), .ZN(new_n9152_));
  NAND2_X1   g09088(.A1(new_n9149_), .A2(new_n9135_), .ZN(new_n9153_));
  NAND2_X1   g09089(.A1(new_n9147_), .A2(new_n9142_), .ZN(new_n9154_));
  NAND2_X1   g09090(.A1(new_n9154_), .A2(new_n9153_), .ZN(new_n9155_));
  NAND3_X1   g09091(.A1(new_n9155_), .A2(new_n9107_), .A3(new_n9152_), .ZN(new_n9156_));
  OAI22_X1   g09092(.A1(new_n1409_), .A2(new_n6788_), .B1(new_n1333_), .B2(new_n6785_), .ZN(new_n9157_));
  NAND2_X1   g09093(.A1(new_n2359_), .A2(new_n7530_), .ZN(new_n9158_));
  AOI21_X1   g09094(.A1(new_n9157_), .A2(new_n9158_), .B(new_n6776_), .ZN(new_n9159_));
  NAND3_X1   g09095(.A1(new_n3828_), .A2(new_n4009_), .A3(new_n9159_), .ZN(new_n9160_));
  INV_X1     g09096(.I(new_n9160_), .ZN(new_n9161_));
  AOI21_X1   g09097(.A1(new_n3828_), .A2(new_n9159_), .B(new_n4009_), .ZN(new_n9162_));
  NOR2_X1    g09098(.A1(new_n9161_), .A2(new_n9162_), .ZN(new_n9163_));
  NAND3_X1   g09099(.A1(new_n9163_), .A2(new_n9151_), .A3(new_n9156_), .ZN(new_n9164_));
  INV_X1     g09100(.I(new_n9162_), .ZN(new_n9165_));
  AOI22_X1   g09101(.A1(new_n9156_), .A2(new_n9151_), .B1(new_n9160_), .B2(new_n9165_), .ZN(new_n9166_));
  AOI21_X1   g09102(.A1(new_n9128_), .A2(new_n9164_), .B(new_n9166_), .ZN(new_n9167_));
  AOI21_X1   g09103(.A1(new_n9152_), .A2(new_n9107_), .B(new_n9143_), .ZN(new_n9168_));
  NAND2_X1   g09104(.A1(new_n6442_), .A2(new_n6368_), .ZN(new_n9169_));
  NAND2_X1   g09105(.A1(new_n6443_), .A2(new_n6361_), .ZN(new_n9170_));
  AOI21_X1   g09106(.A1(new_n9170_), .A2(new_n9169_), .B(new_n6342_), .ZN(new_n9171_));
  NAND2_X1   g09107(.A1(new_n6361_), .A2(new_n6368_), .ZN(new_n9172_));
  AOI21_X1   g09108(.A1(new_n6445_), .A2(new_n9172_), .B(new_n6439_), .ZN(new_n9173_));
  OAI22_X1   g09109(.A1(new_n1453_), .A2(new_n4710_), .B1(new_n2351_), .B2(new_n4719_), .ZN(new_n9174_));
  NAND2_X1   g09110(.A1(new_n2310_), .A2(new_n6480_), .ZN(new_n9175_));
  AOI21_X1   g09111(.A1(new_n9175_), .A2(new_n9174_), .B(new_n4707_), .ZN(new_n9176_));
  NAND2_X1   g09112(.A1(new_n4231_), .A2(new_n9176_), .ZN(new_n9177_));
  XOR2_X1    g09113(.A1(new_n9177_), .A2(new_n4034_), .Z(new_n9178_));
  NOR3_X1    g09114(.A1(new_n9178_), .A2(new_n9171_), .A3(new_n9173_), .ZN(new_n9179_));
  OAI21_X1   g09115(.A1(new_n9171_), .A2(new_n9173_), .B(new_n9178_), .ZN(new_n9180_));
  INV_X1     g09116(.I(new_n9180_), .ZN(new_n9181_));
  OAI22_X1   g09117(.A1(new_n9181_), .A2(new_n9179_), .B1(new_n9150_), .B2(new_n9168_), .ZN(new_n9182_));
  NOR2_X1    g09118(.A1(new_n9168_), .A2(new_n9150_), .ZN(new_n9183_));
  INV_X1     g09119(.I(new_n9171_), .ZN(new_n9184_));
  INV_X1     g09120(.I(new_n9172_), .ZN(new_n9185_));
  OAI21_X1   g09121(.A1(new_n9185_), .A2(new_n6370_), .B(new_n6342_), .ZN(new_n9186_));
  AOI21_X1   g09122(.A1(new_n9184_), .A2(new_n9186_), .B(new_n9178_), .ZN(new_n9187_));
  XOR2_X1    g09123(.A1(new_n9177_), .A2(\a[11] ), .Z(new_n9188_));
  NOR3_X1    g09124(.A1(new_n9188_), .A2(new_n9171_), .A3(new_n9173_), .ZN(new_n9189_));
  OAI21_X1   g09125(.A1(new_n9187_), .A2(new_n9189_), .B(new_n9183_), .ZN(new_n9190_));
  OAI22_X1   g09126(.A1(new_n1409_), .A2(new_n6783_), .B1(new_n2367_), .B2(new_n6785_), .ZN(new_n9191_));
  NAND2_X1   g09127(.A1(new_n1334_), .A2(new_n6789_), .ZN(new_n9192_));
  AOI21_X1   g09128(.A1(new_n9191_), .A2(new_n9192_), .B(new_n6776_), .ZN(new_n9193_));
  NAND2_X1   g09129(.A1(new_n3654_), .A2(new_n9193_), .ZN(new_n9194_));
  XOR2_X1    g09130(.A1(new_n9194_), .A2(new_n4009_), .Z(new_n9195_));
  AOI21_X1   g09131(.A1(new_n9190_), .A2(new_n9182_), .B(new_n9195_), .ZN(new_n9196_));
  NAND3_X1   g09132(.A1(new_n9190_), .A2(new_n9182_), .A3(new_n9195_), .ZN(new_n9197_));
  OAI21_X1   g09133(.A1(new_n9196_), .A2(new_n9167_), .B(new_n9197_), .ZN(new_n9198_));
  OAI22_X1   g09134(.A1(new_n2367_), .A2(new_n6788_), .B1(new_n2408_), .B2(new_n6785_), .ZN(new_n9199_));
  NAND2_X1   g09135(.A1(new_n1334_), .A2(new_n7530_), .ZN(new_n9200_));
  AOI21_X1   g09136(.A1(new_n9199_), .A2(new_n9200_), .B(new_n6776_), .ZN(new_n9201_));
  NAND3_X1   g09137(.A1(new_n3708_), .A2(new_n4009_), .A3(new_n9201_), .ZN(new_n9202_));
  NOR2_X1    g09138(.A1(new_n3703_), .A2(new_n3707_), .ZN(new_n9203_));
  OAI21_X1   g09139(.A1(new_n9203_), .A2(new_n3705_), .B(new_n9201_), .ZN(new_n9204_));
  NAND2_X1   g09140(.A1(new_n9204_), .A2(\a[8] ), .ZN(new_n9205_));
  NAND2_X1   g09141(.A1(new_n9202_), .A2(new_n9205_), .ZN(new_n9206_));
  NAND2_X1   g09142(.A1(new_n9142_), .A2(new_n9135_), .ZN(new_n9207_));
  NAND2_X1   g09143(.A1(new_n9147_), .A2(new_n9149_), .ZN(new_n9208_));
  OAI21_X1   g09144(.A1(new_n9130_), .A2(new_n9129_), .B(new_n9208_), .ZN(new_n9209_));
  AOI21_X1   g09145(.A1(new_n9209_), .A2(new_n9207_), .B(new_n9187_), .ZN(new_n9210_));
  NOR2_X1    g09146(.A1(new_n9210_), .A2(new_n9189_), .ZN(new_n9211_));
  NOR2_X1    g09147(.A1(new_n1453_), .A2(new_n4719_), .ZN(new_n9212_));
  NOR2_X1    g09148(.A1(new_n1409_), .A2(new_n4710_), .ZN(new_n9213_));
  NOR2_X1    g09149(.A1(new_n2351_), .A2(new_n4716_), .ZN(new_n9214_));
  NOR4_X1    g09150(.A1(new_n9213_), .A2(new_n4707_), .A3(new_n9212_), .A4(new_n9214_), .ZN(new_n9215_));
  AOI21_X1   g09151(.A1(new_n3904_), .A2(new_n9215_), .B(new_n4034_), .ZN(new_n9216_));
  INV_X1     g09152(.I(new_n9216_), .ZN(new_n9217_));
  NAND3_X1   g09153(.A1(new_n3904_), .A2(new_n4034_), .A3(new_n9215_), .ZN(new_n9218_));
  NAND2_X1   g09154(.A1(new_n6384_), .A2(new_n6379_), .ZN(new_n9219_));
  NAND2_X1   g09155(.A1(new_n6446_), .A2(new_n9219_), .ZN(new_n9220_));
  NAND3_X1   g09156(.A1(new_n6378_), .A2(new_n6382_), .A3(new_n6376_), .ZN(new_n9221_));
  OAI21_X1   g09157(.A1(new_n6383_), .A2(new_n6377_), .B(new_n6372_), .ZN(new_n9222_));
  NAND2_X1   g09158(.A1(new_n9222_), .A2(new_n9221_), .ZN(new_n9223_));
  NAND3_X1   g09159(.A1(new_n9223_), .A2(new_n6444_), .A3(new_n6445_), .ZN(new_n9224_));
  NAND4_X1   g09160(.A1(new_n9220_), .A2(new_n9217_), .A3(new_n9218_), .A4(new_n9224_), .ZN(new_n9225_));
  INV_X1     g09161(.I(new_n9218_), .ZN(new_n9226_));
  AOI22_X1   g09162(.A1(new_n6444_), .A2(new_n6445_), .B1(new_n6379_), .B2(new_n6384_), .ZN(new_n9227_));
  NOR3_X1    g09163(.A1(new_n6372_), .A2(new_n6383_), .A3(new_n6377_), .ZN(new_n9228_));
  AOI21_X1   g09164(.A1(new_n6378_), .A2(new_n6376_), .B(new_n6382_), .ZN(new_n9229_));
  NOR2_X1    g09165(.A1(new_n9229_), .A2(new_n9228_), .ZN(new_n9230_));
  NOR3_X1    g09166(.A1(new_n9230_), .A2(new_n6369_), .A3(new_n6370_), .ZN(new_n9231_));
  OAI22_X1   g09167(.A1(new_n9231_), .A2(new_n9227_), .B1(new_n9226_), .B2(new_n9216_), .ZN(new_n9232_));
  NAND2_X1   g09168(.A1(new_n9225_), .A2(new_n9232_), .ZN(new_n9233_));
  NAND2_X1   g09169(.A1(new_n9211_), .A2(new_n9233_), .ZN(new_n9234_));
  INV_X1     g09170(.I(new_n9189_), .ZN(new_n9235_));
  NOR2_X1    g09171(.A1(new_n9173_), .A2(new_n9171_), .ZN(new_n9236_));
  OAI22_X1   g09172(.A1(new_n9168_), .A2(new_n9150_), .B1(new_n9236_), .B2(new_n9178_), .ZN(new_n9237_));
  NAND2_X1   g09173(.A1(new_n9237_), .A2(new_n9235_), .ZN(new_n9238_));
  NOR4_X1    g09174(.A1(new_n9231_), .A2(new_n9227_), .A3(new_n9226_), .A4(new_n9216_), .ZN(new_n9239_));
  AOI22_X1   g09175(.A1(new_n9220_), .A2(new_n9224_), .B1(new_n9217_), .B2(new_n9218_), .ZN(new_n9240_));
  NOR2_X1    g09176(.A1(new_n9240_), .A2(new_n9239_), .ZN(new_n9241_));
  NAND2_X1   g09177(.A1(new_n9238_), .A2(new_n9241_), .ZN(new_n9242_));
  AOI21_X1   g09178(.A1(new_n9234_), .A2(new_n9242_), .B(new_n9206_), .ZN(new_n9243_));
  INV_X1     g09179(.I(new_n9206_), .ZN(new_n9244_));
  NAND2_X1   g09180(.A1(new_n9234_), .A2(new_n9242_), .ZN(new_n9245_));
  NOR2_X1    g09181(.A1(new_n9245_), .A2(new_n9244_), .ZN(new_n9246_));
  OAI21_X1   g09182(.A1(new_n9246_), .A2(new_n9243_), .B(new_n9198_), .ZN(new_n9247_));
  INV_X1     g09183(.I(new_n9198_), .ZN(new_n9248_));
  XOR2_X1    g09184(.A1(new_n9245_), .A2(new_n9244_), .Z(new_n9249_));
  NAND2_X1   g09185(.A1(new_n9249_), .A2(new_n9248_), .ZN(new_n9250_));
  NAND2_X1   g09186(.A1(new_n2496_), .A2(new_n8799_), .ZN(new_n9251_));
  AOI22_X1   g09187(.A1(new_n1122_), .A2(new_n6838_), .B1(new_n2454_), .B2(new_n6846_), .ZN(new_n9252_));
  NAND4_X1   g09188(.A1(new_n3393_), .A2(new_n6835_), .A3(new_n9251_), .A4(new_n9252_), .ZN(new_n9253_));
  XOR2_X1    g09189(.A1(new_n9253_), .A2(\a[5] ), .Z(new_n9254_));
  AOI21_X1   g09190(.A1(new_n9250_), .A2(new_n9247_), .B(new_n9254_), .ZN(new_n9255_));
  INV_X1     g09191(.I(new_n9255_), .ZN(new_n9256_));
  OAI21_X1   g09192(.A1(new_n6451_), .A2(new_n6399_), .B(new_n6385_), .ZN(new_n9257_));
  NAND3_X1   g09193(.A1(new_n6397_), .A2(new_n6388_), .A3(new_n6389_), .ZN(new_n9258_));
  NAND2_X1   g09194(.A1(new_n6390_), .A2(new_n6450_), .ZN(new_n9259_));
  NAND2_X1   g09195(.A1(new_n9259_), .A2(new_n9258_), .ZN(new_n9260_));
  NAND2_X1   g09196(.A1(new_n9260_), .A2(new_n6448_), .ZN(new_n9261_));
  OAI22_X1   g09197(.A1(new_n1409_), .A2(new_n4719_), .B1(new_n1333_), .B2(new_n4710_), .ZN(new_n9262_));
  NAND2_X1   g09198(.A1(new_n2359_), .A2(new_n6480_), .ZN(new_n9263_));
  AOI21_X1   g09199(.A1(new_n9262_), .A2(new_n9263_), .B(new_n4707_), .ZN(new_n9264_));
  NAND3_X1   g09200(.A1(new_n3828_), .A2(new_n4034_), .A3(new_n9264_), .ZN(new_n9265_));
  AOI21_X1   g09201(.A1(new_n3828_), .A2(new_n9264_), .B(new_n4034_), .ZN(new_n9266_));
  INV_X1     g09202(.I(new_n9266_), .ZN(new_n9267_));
  NAND4_X1   g09203(.A1(new_n9257_), .A2(new_n9261_), .A3(new_n9265_), .A4(new_n9267_), .ZN(new_n9268_));
  AOI22_X1   g09204(.A1(new_n6398_), .A2(new_n6452_), .B1(new_n6380_), .B2(new_n6384_), .ZN(new_n9269_));
  AOI21_X1   g09205(.A1(new_n9258_), .A2(new_n9259_), .B(new_n6385_), .ZN(new_n9270_));
  INV_X1     g09206(.I(new_n9265_), .ZN(new_n9271_));
  OAI22_X1   g09207(.A1(new_n9270_), .A2(new_n9269_), .B1(new_n9271_), .B2(new_n9266_), .ZN(new_n9272_));
  NAND3_X1   g09208(.A1(new_n9241_), .A2(new_n9237_), .A3(new_n9235_), .ZN(new_n9273_));
  NAND4_X1   g09209(.A1(new_n9273_), .A2(new_n9225_), .A3(new_n9268_), .A4(new_n9272_), .ZN(new_n9274_));
  NAND2_X1   g09210(.A1(new_n9272_), .A2(new_n9268_), .ZN(new_n9275_));
  NAND2_X1   g09211(.A1(new_n9273_), .A2(new_n9225_), .ZN(new_n9276_));
  NAND2_X1   g09212(.A1(new_n9276_), .A2(new_n9275_), .ZN(new_n9277_));
  OAI22_X1   g09213(.A1(new_n2367_), .A2(new_n6783_), .B1(new_n2451_), .B2(new_n6785_), .ZN(new_n9278_));
  NAND2_X1   g09214(.A1(new_n2412_), .A2(new_n6789_), .ZN(new_n9279_));
  AOI21_X1   g09215(.A1(new_n9278_), .A2(new_n9279_), .B(new_n6776_), .ZN(new_n9280_));
  NAND3_X1   g09216(.A1(new_n3403_), .A2(new_n4009_), .A3(new_n9280_), .ZN(new_n9281_));
  NAND2_X1   g09217(.A1(new_n3403_), .A2(new_n9280_), .ZN(new_n9282_));
  NAND2_X1   g09218(.A1(new_n9282_), .A2(\a[8] ), .ZN(new_n9283_));
  NAND2_X1   g09219(.A1(new_n9283_), .A2(new_n9281_), .ZN(new_n9284_));
  NAND3_X1   g09220(.A1(new_n9277_), .A2(new_n9284_), .A3(new_n9274_), .ZN(new_n9285_));
  NOR3_X1    g09221(.A1(new_n9210_), .A2(new_n9233_), .A3(new_n9189_), .ZN(new_n9286_));
  NOR3_X1    g09222(.A1(new_n9275_), .A2(new_n9286_), .A3(new_n9239_), .ZN(new_n9287_));
  AOI22_X1   g09223(.A1(new_n9273_), .A2(new_n9225_), .B1(new_n9268_), .B2(new_n9272_), .ZN(new_n9288_));
  XOR2_X1    g09224(.A1(new_n9282_), .A2(\a[8] ), .Z(new_n9289_));
  OAI21_X1   g09225(.A1(new_n9287_), .A2(new_n9288_), .B(new_n9289_), .ZN(new_n9290_));
  NAND2_X1   g09226(.A1(new_n9290_), .A2(new_n9285_), .ZN(new_n9291_));
  INV_X1     g09227(.I(new_n9245_), .ZN(new_n9292_));
  NOR2_X1    g09228(.A1(new_n9198_), .A2(new_n9244_), .ZN(new_n9293_));
  OAI21_X1   g09229(.A1(new_n9108_), .A2(new_n9120_), .B(new_n9126_), .ZN(new_n9294_));
  AOI22_X1   g09230(.A1(new_n9152_), .A2(new_n9107_), .B1(new_n9208_), .B2(new_n9207_), .ZN(new_n9295_));
  NOR4_X1    g09231(.A1(new_n9148_), .A2(new_n9133_), .A3(new_n9134_), .A4(new_n9140_), .ZN(new_n9296_));
  NOR2_X1    g09232(.A1(new_n9149_), .A2(new_n9135_), .ZN(new_n9297_));
  NOR2_X1    g09233(.A1(new_n9297_), .A2(new_n9296_), .ZN(new_n9298_));
  NOR3_X1    g09234(.A1(new_n9298_), .A2(new_n9130_), .A3(new_n9129_), .ZN(new_n9299_));
  NOR4_X1    g09235(.A1(new_n9299_), .A2(new_n9295_), .A3(new_n9161_), .A4(new_n9162_), .ZN(new_n9300_));
  OAI22_X1   g09236(.A1(new_n9299_), .A2(new_n9295_), .B1(new_n9161_), .B2(new_n9162_), .ZN(new_n9301_));
  OAI21_X1   g09237(.A1(new_n9294_), .A2(new_n9300_), .B(new_n9301_), .ZN(new_n9302_));
  INV_X1     g09238(.I(new_n9179_), .ZN(new_n9303_));
  AOI22_X1   g09239(.A1(new_n9303_), .A2(new_n9180_), .B1(new_n9209_), .B2(new_n9207_), .ZN(new_n9304_));
  NOR2_X1    g09240(.A1(new_n9187_), .A2(new_n9189_), .ZN(new_n9305_));
  NOR3_X1    g09241(.A1(new_n9305_), .A2(new_n9150_), .A3(new_n9168_), .ZN(new_n9306_));
  XOR2_X1    g09242(.A1(new_n9194_), .A2(\a[8] ), .Z(new_n9307_));
  OAI21_X1   g09243(.A1(new_n9306_), .A2(new_n9304_), .B(new_n9307_), .ZN(new_n9308_));
  NAND2_X1   g09244(.A1(new_n9308_), .A2(new_n9302_), .ZN(new_n9309_));
  AOI21_X1   g09245(.A1(new_n9309_), .A2(new_n9197_), .B(new_n9206_), .ZN(new_n9310_));
  OAI21_X1   g09246(.A1(new_n9293_), .A2(new_n9310_), .B(new_n9292_), .ZN(new_n9311_));
  NOR2_X1    g09247(.A1(new_n9311_), .A2(new_n9291_), .ZN(new_n9312_));
  NOR3_X1    g09248(.A1(new_n9289_), .A2(new_n9287_), .A3(new_n9288_), .ZN(new_n9313_));
  AOI21_X1   g09249(.A1(new_n9277_), .A2(new_n9274_), .B(new_n9284_), .ZN(new_n9314_));
  NOR2_X1    g09250(.A1(new_n9314_), .A2(new_n9313_), .ZN(new_n9315_));
  NAND3_X1   g09251(.A1(new_n9309_), .A2(new_n9197_), .A3(new_n9206_), .ZN(new_n9316_));
  NAND2_X1   g09252(.A1(new_n9198_), .A2(new_n9244_), .ZN(new_n9317_));
  AOI21_X1   g09253(.A1(new_n9317_), .A2(new_n9316_), .B(new_n9245_), .ZN(new_n9318_));
  NOR2_X1    g09254(.A1(new_n9318_), .A2(new_n9315_), .ZN(new_n9319_));
  NOR2_X1    g09255(.A1(new_n9248_), .A2(new_n9244_), .ZN(new_n9320_));
  INV_X1     g09256(.I(new_n9320_), .ZN(new_n9321_));
  NOR3_X1    g09257(.A1(new_n9312_), .A2(new_n9319_), .A3(new_n9321_), .ZN(new_n9322_));
  NAND2_X1   g09258(.A1(new_n9318_), .A2(new_n9315_), .ZN(new_n9323_));
  NAND2_X1   g09259(.A1(new_n9311_), .A2(new_n9291_), .ZN(new_n9324_));
  AOI21_X1   g09260(.A1(new_n9324_), .A2(new_n9323_), .B(new_n9320_), .ZN(new_n9325_));
  OAI22_X1   g09261(.A1(new_n1180_), .A2(new_n6839_), .B1(new_n2492_), .B2(new_n6913_), .ZN(new_n9326_));
  NAND2_X1   g09262(.A1(new_n1122_), .A2(new_n8799_), .ZN(new_n9327_));
  AOI21_X1   g09263(.A1(new_n9327_), .A2(new_n9326_), .B(new_n6836_), .ZN(new_n9328_));
  NAND2_X1   g09264(.A1(new_n3330_), .A2(new_n9328_), .ZN(new_n9329_));
  XOR2_X1    g09265(.A1(new_n9329_), .A2(\a[5] ), .Z(new_n9330_));
  INV_X1     g09266(.I(new_n9330_), .ZN(new_n9331_));
  NOR3_X1    g09267(.A1(new_n9325_), .A2(new_n9322_), .A3(new_n9331_), .ZN(new_n9332_));
  OAI21_X1   g09268(.A1(new_n9325_), .A2(new_n9322_), .B(new_n9331_), .ZN(new_n9333_));
  OAI21_X1   g09269(.A1(new_n9256_), .A2(new_n9332_), .B(new_n9333_), .ZN(new_n9334_));
  XOR2_X1    g09270(.A1(new_n6406_), .A2(new_n6412_), .Z(new_n9335_));
  NAND2_X1   g09271(.A1(new_n9335_), .A2(new_n6453_), .ZN(new_n9336_));
  OAI21_X1   g09272(.A1(new_n6413_), .A2(new_n6455_), .B(new_n6400_), .ZN(new_n9337_));
  NAND2_X1   g09273(.A1(new_n9336_), .A2(new_n9337_), .ZN(new_n9338_));
  NOR2_X1    g09274(.A1(new_n9286_), .A2(new_n9239_), .ZN(new_n9339_));
  NAND2_X1   g09275(.A1(new_n9272_), .A2(new_n9268_), .ZN(new_n9340_));
  OAI22_X1   g09276(.A1(new_n1409_), .A2(new_n4716_), .B1(new_n2367_), .B2(new_n4710_), .ZN(new_n9341_));
  NAND2_X1   g09277(.A1(new_n1334_), .A2(new_n4720_), .ZN(new_n9342_));
  AOI21_X1   g09278(.A1(new_n9341_), .A2(new_n9342_), .B(new_n4707_), .ZN(new_n9343_));
  NAND2_X1   g09279(.A1(new_n3654_), .A2(new_n9343_), .ZN(new_n9344_));
  XOR2_X1    g09280(.A1(new_n9344_), .A2(\a[11] ), .Z(new_n9345_));
  OAI21_X1   g09281(.A1(new_n9339_), .A2(new_n9340_), .B(new_n9345_), .ZN(new_n9346_));
  INV_X1     g09282(.I(new_n9340_), .ZN(new_n9347_));
  INV_X1     g09283(.I(new_n9345_), .ZN(new_n9348_));
  NAND3_X1   g09284(.A1(new_n9347_), .A2(new_n9276_), .A3(new_n9348_), .ZN(new_n9349_));
  AOI21_X1   g09285(.A1(new_n9349_), .A2(new_n9346_), .B(new_n9338_), .ZN(new_n9350_));
  INV_X1     g09286(.I(new_n9338_), .ZN(new_n9351_));
  AOI21_X1   g09287(.A1(new_n9347_), .A2(new_n9276_), .B(new_n9348_), .ZN(new_n9352_));
  NOR3_X1    g09288(.A1(new_n9339_), .A2(new_n9340_), .A3(new_n9345_), .ZN(new_n9353_));
  NOR3_X1    g09289(.A1(new_n9352_), .A2(new_n9353_), .A3(new_n9351_), .ZN(new_n9354_));
  NOR2_X1    g09290(.A1(new_n9350_), .A2(new_n9354_), .ZN(new_n9355_));
  NOR2_X1    g09291(.A1(new_n9238_), .A2(new_n9241_), .ZN(new_n9356_));
  NOR2_X1    g09292(.A1(new_n9211_), .A2(new_n9233_), .ZN(new_n9357_));
  OAI21_X1   g09293(.A1(new_n9356_), .A2(new_n9357_), .B(new_n9244_), .ZN(new_n9358_));
  NOR2_X1    g09294(.A1(new_n9358_), .A2(new_n9198_), .ZN(new_n9359_));
  NOR3_X1    g09295(.A1(new_n9359_), .A2(new_n9314_), .A3(new_n9243_), .ZN(new_n9360_));
  OAI22_X1   g09296(.A1(new_n2492_), .A2(new_n6785_), .B1(new_n2408_), .B2(new_n6783_), .ZN(new_n9361_));
  NAND2_X1   g09297(.A1(new_n2454_), .A2(new_n6789_), .ZN(new_n9362_));
  AOI21_X1   g09298(.A1(new_n9362_), .A2(new_n9361_), .B(new_n6776_), .ZN(new_n9363_));
  NAND2_X1   g09299(.A1(new_n3577_), .A2(new_n9363_), .ZN(new_n9364_));
  XOR2_X1    g09300(.A1(new_n9364_), .A2(\a[8] ), .Z(new_n9365_));
  INV_X1     g09301(.I(new_n9365_), .ZN(new_n9366_));
  AOI21_X1   g09302(.A1(new_n9360_), .A2(new_n9315_), .B(new_n9366_), .ZN(new_n9367_));
  NAND3_X1   g09303(.A1(new_n9243_), .A2(new_n9309_), .A3(new_n9197_), .ZN(new_n9368_));
  NAND4_X1   g09304(.A1(new_n9290_), .A2(new_n9368_), .A3(new_n9285_), .A4(new_n9358_), .ZN(new_n9369_));
  NOR2_X1    g09305(.A1(new_n9369_), .A2(new_n9365_), .ZN(new_n9370_));
  OAI21_X1   g09306(.A1(new_n9367_), .A2(new_n9370_), .B(new_n9355_), .ZN(new_n9371_));
  INV_X1     g09307(.I(new_n9355_), .ZN(new_n9372_));
  NAND2_X1   g09308(.A1(new_n9369_), .A2(new_n9365_), .ZN(new_n9373_));
  NAND3_X1   g09309(.A1(new_n9360_), .A2(new_n9315_), .A3(new_n9366_), .ZN(new_n9374_));
  NAND3_X1   g09310(.A1(new_n9374_), .A2(new_n9373_), .A3(new_n9372_), .ZN(new_n9375_));
  NAND2_X1   g09311(.A1(new_n9375_), .A2(new_n9371_), .ZN(new_n9376_));
  OAI22_X1   g09312(.A1(new_n1008_), .A2(new_n6839_), .B1(new_n1121_), .B2(new_n6913_), .ZN(new_n9377_));
  NAND2_X1   g09313(.A1(new_n1181_), .A2(new_n8799_), .ZN(new_n9378_));
  AOI21_X1   g09314(.A1(new_n9377_), .A2(new_n9378_), .B(new_n6836_), .ZN(new_n9379_));
  NAND2_X1   g09315(.A1(new_n3562_), .A2(new_n9379_), .ZN(new_n9380_));
  XOR2_X1    g09316(.A1(new_n9380_), .A2(new_n65_), .Z(new_n9381_));
  INV_X1     g09317(.I(new_n9381_), .ZN(new_n9382_));
  NAND2_X1   g09318(.A1(new_n9376_), .A2(new_n9382_), .ZN(new_n9383_));
  NAND3_X1   g09319(.A1(new_n9381_), .A2(new_n9375_), .A3(new_n9371_), .ZN(new_n9384_));
  INV_X1     g09320(.I(new_n9384_), .ZN(new_n9385_));
  AOI21_X1   g09321(.A1(new_n9334_), .A2(new_n9383_), .B(new_n9385_), .ZN(new_n9386_));
  OAI22_X1   g09322(.A1(new_n896_), .A2(new_n6839_), .B1(new_n1180_), .B2(new_n6913_), .ZN(new_n9387_));
  NAND2_X1   g09323(.A1(new_n2504_), .A2(new_n8799_), .ZN(new_n9388_));
  AOI21_X1   g09324(.A1(new_n9388_), .A2(new_n9387_), .B(new_n6836_), .ZN(new_n9389_));
  NAND2_X1   g09325(.A1(new_n3596_), .A2(new_n9389_), .ZN(new_n9390_));
  XOR2_X1    g09326(.A1(new_n9390_), .A2(\a[5] ), .Z(new_n9391_));
  NOR4_X1    g09327(.A1(new_n8955_), .A2(new_n8951_), .A3(new_n9386_), .A4(new_n9391_), .ZN(new_n9392_));
  NOR2_X1    g09328(.A1(new_n8916_), .A2(new_n8913_), .ZN(new_n9393_));
  NAND3_X1   g09329(.A1(new_n9324_), .A2(new_n9323_), .A3(new_n9320_), .ZN(new_n9394_));
  OAI21_X1   g09330(.A1(new_n9312_), .A2(new_n9319_), .B(new_n9321_), .ZN(new_n9395_));
  NAND3_X1   g09331(.A1(new_n9395_), .A2(new_n9394_), .A3(new_n9330_), .ZN(new_n9396_));
  AOI21_X1   g09332(.A1(new_n9395_), .A2(new_n9394_), .B(new_n9330_), .ZN(new_n9397_));
  AOI21_X1   g09333(.A1(new_n9255_), .A2(new_n9396_), .B(new_n9397_), .ZN(new_n9398_));
  AOI21_X1   g09334(.A1(new_n9371_), .A2(new_n9375_), .B(new_n9381_), .ZN(new_n9399_));
  OAI21_X1   g09335(.A1(new_n9398_), .A2(new_n9399_), .B(new_n9384_), .ZN(new_n9400_));
  NOR2_X1    g09336(.A1(new_n9400_), .A2(new_n9391_), .ZN(new_n9401_));
  INV_X1     g09337(.I(new_n9391_), .ZN(new_n9402_));
  NOR2_X1    g09338(.A1(new_n9386_), .A2(new_n9402_), .ZN(new_n9403_));
  OAI21_X1   g09339(.A1(new_n9403_), .A2(new_n9401_), .B(new_n9393_), .ZN(new_n9404_));
  NOR2_X1    g09340(.A1(new_n9404_), .A2(new_n9392_), .ZN(new_n9405_));
  NOR3_X1    g09341(.A1(new_n8937_), .A2(new_n8927_), .A3(new_n8880_), .ZN(new_n9406_));
  OAI21_X1   g09342(.A1(new_n8935_), .A2(new_n8936_), .B(new_n8928_), .ZN(new_n9407_));
  NAND3_X1   g09343(.A1(new_n8924_), .A2(new_n8926_), .A3(new_n8884_), .ZN(new_n9408_));
  AOI21_X1   g09344(.A1(new_n9407_), .A2(new_n9408_), .B(new_n8881_), .ZN(new_n9409_));
  NOR2_X1    g09345(.A1(new_n8954_), .A2(new_n8947_), .ZN(new_n9410_));
  INV_X1     g09346(.I(new_n9410_), .ZN(new_n9411_));
  OAI21_X1   g09347(.A1(new_n9409_), .A2(new_n9406_), .B(new_n9411_), .ZN(new_n9412_));
  OAI21_X1   g09348(.A1(new_n9405_), .A2(new_n9412_), .B(new_n8940_), .ZN(new_n9413_));
  AOI21_X1   g09349(.A1(new_n8827_), .A2(new_n8853_), .B(\a[5] ), .ZN(new_n9414_));
  NAND3_X1   g09350(.A1(new_n8827_), .A2(new_n8853_), .A3(\a[5] ), .ZN(new_n9415_));
  INV_X1     g09351(.I(new_n9415_), .ZN(new_n9416_));
  OAI21_X1   g09352(.A1(new_n9416_), .A2(new_n9414_), .B(new_n8871_), .ZN(new_n9417_));
  INV_X1     g09353(.I(new_n8871_), .ZN(new_n9418_));
  INV_X1     g09354(.I(new_n9414_), .ZN(new_n9419_));
  NAND3_X1   g09355(.A1(new_n9419_), .A2(new_n9415_), .A3(new_n9418_), .ZN(new_n9420_));
  NAND2_X1   g09356(.A1(new_n9420_), .A2(new_n9417_), .ZN(new_n9421_));
  OAI21_X1   g09357(.A1(new_n9413_), .A2(new_n9421_), .B(new_n8874_), .ZN(new_n9422_));
  NAND3_X1   g09358(.A1(new_n9422_), .A2(new_n8862_), .A3(new_n8866_), .ZN(new_n9423_));
  AOI22_X1   g09359(.A1(new_n9423_), .A2(new_n8803_), .B1(new_n8846_), .B2(new_n8850_), .ZN(new_n9424_));
  OAI22_X1   g09360(.A1(new_n694_), .A2(new_n6913_), .B1(new_n2665_), .B2(new_n6839_), .ZN(new_n9425_));
  NAND2_X1   g09361(.A1(new_n2615_), .A2(new_n8799_), .ZN(new_n9426_));
  AOI21_X1   g09362(.A1(new_n9425_), .A2(new_n9426_), .B(new_n6836_), .ZN(new_n9427_));
  AND3_X2    g09363(.A1(new_n3188_), .A2(new_n65_), .A3(new_n9427_), .Z(new_n9428_));
  AOI21_X1   g09364(.A1(new_n3188_), .A2(new_n9427_), .B(new_n65_), .ZN(new_n9429_));
  NOR2_X1    g09365(.A1(new_n9428_), .A2(new_n9429_), .ZN(new_n9430_));
  INV_X1     g09366(.I(new_n9430_), .ZN(new_n9431_));
  NAND2_X1   g09367(.A1(new_n9424_), .A2(new_n9431_), .ZN(new_n9432_));
  NAND2_X1   g09368(.A1(new_n8850_), .A2(new_n8846_), .ZN(new_n9433_));
  INV_X1     g09369(.I(new_n8862_), .ZN(new_n9434_));
  NAND2_X1   g09370(.A1(new_n8866_), .A2(new_n8862_), .ZN(new_n9435_));
  NAND2_X1   g09371(.A1(new_n8954_), .A2(new_n8946_), .ZN(new_n9436_));
  NAND2_X1   g09372(.A1(new_n8947_), .A2(new_n8950_), .ZN(new_n9437_));
  NAND4_X1   g09373(.A1(new_n9436_), .A2(new_n9437_), .A3(new_n9400_), .A4(new_n9402_), .ZN(new_n9438_));
  INV_X1     g09374(.I(new_n9393_), .ZN(new_n9439_));
  NAND2_X1   g09375(.A1(new_n9386_), .A2(new_n9402_), .ZN(new_n9440_));
  NAND2_X1   g09376(.A1(new_n9396_), .A2(new_n9255_), .ZN(new_n9441_));
  AOI21_X1   g09377(.A1(new_n9441_), .A2(new_n9333_), .B(new_n9399_), .ZN(new_n9442_));
  OAI21_X1   g09378(.A1(new_n9442_), .A2(new_n9385_), .B(new_n9391_), .ZN(new_n9443_));
  AOI21_X1   g09379(.A1(new_n9440_), .A2(new_n9443_), .B(new_n9439_), .ZN(new_n9444_));
  NAND2_X1   g09380(.A1(new_n9444_), .A2(new_n9438_), .ZN(new_n9445_));
  NAND3_X1   g09381(.A1(new_n9407_), .A2(new_n9408_), .A3(new_n8881_), .ZN(new_n9446_));
  OAI21_X1   g09382(.A1(new_n8937_), .A2(new_n8927_), .B(new_n8880_), .ZN(new_n9447_));
  AOI21_X1   g09383(.A1(new_n9446_), .A2(new_n9447_), .B(new_n9410_), .ZN(new_n9448_));
  AOI21_X1   g09384(.A1(new_n9445_), .A2(new_n9448_), .B(new_n8939_), .ZN(new_n9449_));
  AOI21_X1   g09385(.A1(new_n9419_), .A2(new_n9415_), .B(new_n9418_), .ZN(new_n9450_));
  NOR3_X1    g09386(.A1(new_n9416_), .A2(new_n9414_), .A3(new_n8871_), .ZN(new_n9451_));
  NOR2_X1    g09387(.A1(new_n9450_), .A2(new_n9451_), .ZN(new_n9452_));
  AOI21_X1   g09388(.A1(new_n9449_), .A2(new_n9452_), .B(new_n8873_), .ZN(new_n9453_));
  NOR3_X1    g09389(.A1(new_n9453_), .A2(new_n9434_), .A3(new_n9435_), .ZN(new_n9454_));
  OAI21_X1   g09390(.A1(new_n8847_), .A2(new_n9454_), .B(new_n9433_), .ZN(new_n9455_));
  INV_X1     g09391(.I(new_n6891_), .ZN(new_n9456_));
  NOR2_X1    g09392(.A1(new_n6893_), .A2(new_n6892_), .ZN(new_n9457_));
  NAND2_X1   g09393(.A1(new_n9457_), .A2(new_n9456_), .ZN(new_n9458_));
  NAND2_X1   g09394(.A1(new_n9458_), .A2(new_n6894_), .ZN(new_n9459_));
  NAND2_X1   g09395(.A1(new_n9459_), .A2(new_n9430_), .ZN(new_n9460_));
  INV_X1     g09396(.I(new_n9460_), .ZN(new_n9461_));
  NAND2_X1   g09397(.A1(new_n9455_), .A2(new_n9461_), .ZN(new_n9462_));
  NAND2_X1   g09398(.A1(new_n9462_), .A2(new_n9432_), .ZN(new_n9463_));
  NAND2_X1   g09399(.A1(new_n6905_), .A2(new_n6906_), .ZN(new_n9464_));
  XOR2_X1    g09400(.A1(new_n9464_), .A2(new_n9458_), .Z(new_n9465_));
  INV_X1     g09401(.I(new_n9465_), .ZN(new_n9466_));
  NAND2_X1   g09402(.A1(new_n9463_), .A2(new_n9466_), .ZN(new_n9467_));
  AND2_X2    g09403(.A1(new_n2733_), .A2(new_n6835_), .Z(new_n9468_));
  OAI22_X1   g09404(.A1(new_n2665_), .A2(new_n6843_), .B1(new_n2614_), .B2(new_n6913_), .ZN(new_n9469_));
  OAI21_X1   g09405(.A1(new_n2716_), .A2(new_n6839_), .B(new_n9469_), .ZN(new_n9470_));
  NOR2_X1    g09406(.A1(new_n9468_), .A2(new_n9470_), .ZN(new_n9471_));
  XOR2_X1    g09407(.A1(new_n9471_), .A2(\a[5] ), .Z(new_n9472_));
  OAI21_X1   g09408(.A1(new_n9463_), .A2(new_n9466_), .B(new_n9472_), .ZN(new_n9473_));
  NAND2_X1   g09409(.A1(new_n9473_), .A2(new_n9467_), .ZN(new_n9474_));
  AND3_X2    g09410(.A1(new_n9474_), .A2(new_n8786_), .A3(new_n8797_), .Z(new_n9475_));
  AOI22_X1   g09411(.A1(new_n8794_), .A2(new_n8796_), .B1(new_n9473_), .B2(new_n9467_), .ZN(new_n9476_));
  NOR2_X1    g09412(.A1(new_n9476_), .A2(new_n8786_), .ZN(new_n9477_));
  NOR2_X1    g09413(.A1(new_n9475_), .A2(new_n9477_), .ZN(new_n9478_));
  INV_X1     g09414(.I(new_n9478_), .ZN(new_n9479_));
  XNOR2_X1   g09415(.A1(new_n9459_), .A2(new_n9430_), .ZN(new_n9480_));
  INV_X1     g09416(.I(new_n9480_), .ZN(new_n9481_));
  INV_X1     g09417(.I(new_n6922_), .ZN(new_n9482_));
  NAND2_X1   g09418(.A1(new_n6920_), .A2(\a[1] ), .ZN(new_n9483_));
  NOR2_X1    g09419(.A1(new_n3176_), .A2(new_n9483_), .ZN(new_n9484_));
  INV_X1     g09420(.I(new_n6925_), .ZN(new_n9485_));
  NOR2_X1    g09421(.A1(new_n2716_), .A2(new_n9485_), .ZN(new_n9486_));
  XOR2_X1    g09422(.A1(\a[1] ), .A2(\a[2] ), .Z(new_n9487_));
  NOR2_X1    g09423(.A1(new_n9487_), .A2(new_n6920_), .ZN(new_n9488_));
  INV_X1     g09424(.I(new_n9488_), .ZN(new_n9489_));
  NOR2_X1    g09425(.A1(new_n3142_), .A2(new_n9489_), .ZN(new_n9490_));
  NOR4_X1    g09426(.A1(new_n9484_), .A2(new_n9482_), .A3(new_n9486_), .A4(new_n9490_), .ZN(new_n9491_));
  AOI21_X1   g09427(.A1(new_n3174_), .A2(new_n9491_), .B(\a[2] ), .ZN(new_n9492_));
  NAND3_X1   g09428(.A1(new_n3174_), .A2(\a[2] ), .A3(new_n9491_), .ZN(new_n9493_));
  INV_X1     g09429(.I(new_n9493_), .ZN(new_n9494_));
  NOR3_X1    g09430(.A1(new_n9494_), .A2(new_n9481_), .A3(new_n9492_), .ZN(new_n9495_));
  INV_X1     g09431(.I(new_n9492_), .ZN(new_n9496_));
  AOI21_X1   g09432(.A1(new_n9496_), .A2(new_n9493_), .B(new_n9480_), .ZN(new_n9497_));
  OAI21_X1   g09433(.A1(new_n9495_), .A2(new_n9497_), .B(new_n9424_), .ZN(new_n9498_));
  NOR3_X1    g09434(.A1(new_n9494_), .A2(new_n9480_), .A3(new_n9492_), .ZN(new_n9499_));
  AOI21_X1   g09435(.A1(new_n9496_), .A2(new_n9493_), .B(new_n9481_), .ZN(new_n9500_));
  OAI21_X1   g09436(.A1(new_n9500_), .A2(new_n9499_), .B(new_n9455_), .ZN(new_n9501_));
  OAI22_X1   g09437(.A1(new_n3176_), .A2(new_n9489_), .B1(new_n2665_), .B2(new_n9485_), .ZN(new_n9502_));
  INV_X1     g09438(.I(new_n9483_), .ZN(new_n9503_));
  NAND2_X1   g09439(.A1(new_n2728_), .A2(new_n9503_), .ZN(new_n9504_));
  AOI21_X1   g09440(.A1(new_n9502_), .A2(new_n9504_), .B(new_n9482_), .ZN(new_n9505_));
  NAND2_X1   g09441(.A1(new_n3273_), .A2(new_n9505_), .ZN(new_n9506_));
  XOR2_X1    g09442(.A1(new_n9506_), .A2(\a[2] ), .Z(new_n9507_));
  NOR2_X1    g09443(.A1(new_n8848_), .A2(new_n8849_), .ZN(new_n9508_));
  INV_X1     g09444(.I(new_n9508_), .ZN(new_n9509_));
  NAND2_X1   g09445(.A1(new_n9423_), .A2(new_n8847_), .ZN(new_n9510_));
  NOR4_X1    g09446(.A1(new_n9453_), .A2(new_n8847_), .A3(new_n9434_), .A4(new_n9435_), .ZN(new_n9511_));
  INV_X1     g09447(.I(new_n9511_), .ZN(new_n9512_));
  AOI21_X1   g09448(.A1(new_n9510_), .A2(new_n9512_), .B(new_n9509_), .ZN(new_n9513_));
  NOR2_X1    g09449(.A1(new_n9454_), .A2(new_n8803_), .ZN(new_n9514_));
  NOR3_X1    g09450(.A1(new_n9514_), .A2(new_n9508_), .A3(new_n9511_), .ZN(new_n9515_));
  NOR3_X1    g09451(.A1(new_n9513_), .A2(new_n9515_), .A3(new_n9507_), .ZN(new_n9516_));
  NAND3_X1   g09452(.A1(new_n9516_), .A2(new_n9501_), .A3(new_n9498_), .ZN(new_n9517_));
  NAND3_X1   g09453(.A1(new_n9496_), .A2(new_n9480_), .A3(new_n9493_), .ZN(new_n9518_));
  OAI21_X1   g09454(.A1(new_n9494_), .A2(new_n9492_), .B(new_n9481_), .ZN(new_n9519_));
  AOI21_X1   g09455(.A1(new_n9519_), .A2(new_n9518_), .B(new_n9455_), .ZN(new_n9520_));
  NAND3_X1   g09456(.A1(new_n9496_), .A2(new_n9481_), .A3(new_n9493_), .ZN(new_n9521_));
  OAI21_X1   g09457(.A1(new_n9494_), .A2(new_n9492_), .B(new_n9480_), .ZN(new_n9522_));
  AOI21_X1   g09458(.A1(new_n9521_), .A2(new_n9522_), .B(new_n9424_), .ZN(new_n9523_));
  INV_X1     g09459(.I(new_n9507_), .ZN(new_n9524_));
  OAI21_X1   g09460(.A1(new_n9514_), .A2(new_n9511_), .B(new_n9508_), .ZN(new_n9525_));
  NAND3_X1   g09461(.A1(new_n9510_), .A2(new_n9512_), .A3(new_n9509_), .ZN(new_n9526_));
  NAND3_X1   g09462(.A1(new_n9526_), .A2(new_n9525_), .A3(new_n9524_), .ZN(new_n9527_));
  OAI21_X1   g09463(.A1(new_n9520_), .A2(new_n9523_), .B(new_n9527_), .ZN(new_n9528_));
  NAND2_X1   g09464(.A1(new_n9528_), .A2(new_n9517_), .ZN(new_n9529_));
  XNOR2_X1   g09465(.A1(new_n9453_), .A2(new_n9435_), .ZN(new_n9530_));
  INV_X1     g09466(.I(new_n9530_), .ZN(new_n9531_));
  OAI22_X1   g09467(.A1(new_n2614_), .A2(new_n9489_), .B1(new_n529_), .B2(new_n9485_), .ZN(new_n9532_));
  NAND2_X1   g09468(.A1(new_n2718_), .A2(new_n9503_), .ZN(new_n9533_));
  AOI21_X1   g09469(.A1(new_n9533_), .A2(new_n9532_), .B(new_n9482_), .ZN(new_n9534_));
  NAND2_X1   g09470(.A1(new_n3074_), .A2(new_n9534_), .ZN(new_n9535_));
  XOR2_X1    g09471(.A1(new_n9535_), .A2(\a[2] ), .Z(new_n9536_));
  INV_X1     g09472(.I(new_n9536_), .ZN(new_n9537_));
  AOI21_X1   g09473(.A1(new_n9445_), .A2(new_n9411_), .B(new_n8881_), .ZN(new_n9538_));
  NOR3_X1    g09474(.A1(new_n9405_), .A2(new_n8880_), .A3(new_n9410_), .ZN(new_n9539_));
  OAI21_X1   g09475(.A1(new_n9539_), .A2(new_n9538_), .B(new_n8938_), .ZN(new_n9540_));
  NOR3_X1    g09476(.A1(new_n9539_), .A2(new_n9538_), .A3(new_n8938_), .ZN(new_n9541_));
  INV_X1     g09477(.I(new_n9541_), .ZN(new_n9542_));
  AOI21_X1   g09478(.A1(new_n9542_), .A2(new_n9540_), .B(new_n9537_), .ZN(new_n9543_));
  INV_X1     g09479(.I(new_n9543_), .ZN(new_n9544_));
  NOR2_X1    g09480(.A1(new_n1333_), .A2(new_n9485_), .ZN(new_n9545_));
  NOR2_X1    g09481(.A1(new_n2408_), .A2(new_n9489_), .ZN(new_n9546_));
  NOR2_X1    g09482(.A1(new_n2367_), .A2(new_n9483_), .ZN(new_n9547_));
  NOR4_X1    g09483(.A1(new_n9547_), .A2(new_n9545_), .A3(new_n9546_), .A4(new_n9482_), .ZN(new_n9548_));
  NAND2_X1   g09484(.A1(new_n3708_), .A2(new_n9548_), .ZN(new_n9549_));
  XOR2_X1    g09485(.A1(new_n9549_), .A2(new_n4387_), .Z(new_n9550_));
  XNOR2_X1   g09486(.A1(new_n9009_), .A2(new_n9005_), .ZN(new_n9551_));
  OAI22_X1   g09487(.A1(new_n2311_), .A2(new_n6785_), .B1(new_n4365_), .B2(new_n6783_), .ZN(new_n9552_));
  NAND2_X1   g09488(.A1(new_n2255_), .A2(new_n6789_), .ZN(new_n9553_));
  AOI21_X1   g09489(.A1(new_n9552_), .A2(new_n9553_), .B(new_n6776_), .ZN(new_n9554_));
  NAND2_X1   g09490(.A1(new_n4419_), .A2(new_n9554_), .ZN(new_n9555_));
  XOR2_X1    g09491(.A1(new_n9555_), .A2(\a[8] ), .Z(new_n9556_));
  XOR2_X1    g09492(.A1(new_n9556_), .A2(new_n9551_), .Z(new_n9557_));
  NAND2_X1   g09493(.A1(new_n2359_), .A2(new_n8799_), .ZN(new_n9558_));
  NAND2_X1   g09494(.A1(new_n1408_), .A2(new_n6838_), .ZN(new_n9559_));
  AOI21_X1   g09495(.A1(new_n2354_), .A2(new_n6846_), .B(new_n6836_), .ZN(new_n9560_));
  NAND4_X1   g09496(.A1(new_n3904_), .A2(new_n9558_), .A3(new_n9559_), .A4(new_n9560_), .ZN(new_n9561_));
  XOR2_X1    g09497(.A1(new_n9561_), .A2(\a[5] ), .Z(new_n9562_));
  NOR2_X1    g09498(.A1(new_n9562_), .A2(new_n9557_), .ZN(new_n9563_));
  INV_X1     g09499(.I(new_n9563_), .ZN(new_n9564_));
  NAND2_X1   g09500(.A1(new_n9562_), .A2(new_n9557_), .ZN(new_n9565_));
  NAND2_X1   g09501(.A1(new_n9564_), .A2(new_n9565_), .ZN(new_n9566_));
  INV_X1     g09502(.I(new_n9566_), .ZN(new_n9567_));
  NOR2_X1    g09503(.A1(new_n9550_), .A2(new_n9567_), .ZN(new_n9568_));
  NAND2_X1   g09504(.A1(new_n1334_), .A2(new_n9488_), .ZN(new_n9569_));
  NAND2_X1   g09505(.A1(new_n2359_), .A2(new_n6925_), .ZN(new_n9570_));
  AOI21_X1   g09506(.A1(new_n1408_), .A2(new_n9503_), .B(new_n9482_), .ZN(new_n9571_));
  NAND4_X1   g09507(.A1(new_n3828_), .A2(new_n9569_), .A3(new_n9570_), .A4(new_n9571_), .ZN(new_n9572_));
  XOR2_X1    g09508(.A1(new_n9572_), .A2(\a[2] ), .Z(new_n9573_));
  INV_X1     g09509(.I(new_n9573_), .ZN(new_n9574_));
  NAND2_X1   g09510(.A1(new_n1504_), .A2(new_n6925_), .ZN(new_n9575_));
  NAND2_X1   g09511(.A1(new_n2255_), .A2(new_n9488_), .ZN(new_n9576_));
  AOI21_X1   g09512(.A1(new_n1547_), .A2(new_n9503_), .B(new_n9482_), .ZN(new_n9577_));
  NAND4_X1   g09513(.A1(new_n4650_), .A2(new_n9575_), .A3(new_n9576_), .A4(new_n9577_), .ZN(new_n9578_));
  XOR2_X1    g09514(.A1(new_n9578_), .A2(\a[2] ), .Z(new_n9579_));
  NOR2_X1    g09515(.A1(new_n1503_), .A2(new_n9489_), .ZN(new_n9580_));
  NOR2_X1    g09516(.A1(new_n2198_), .A2(new_n9483_), .ZN(new_n9581_));
  NOR2_X1    g09517(.A1(new_n2158_), .A2(new_n9485_), .ZN(new_n9582_));
  NOR4_X1    g09518(.A1(new_n9582_), .A2(new_n9580_), .A3(new_n9482_), .A4(new_n9581_), .ZN(new_n9583_));
  NAND2_X1   g09519(.A1(new_n4620_), .A2(new_n9583_), .ZN(new_n9584_));
  XOR2_X1    g09520(.A1(new_n9584_), .A2(\a[2] ), .Z(new_n9585_));
  NOR2_X1    g09521(.A1(new_n5069_), .A2(new_n2071_), .ZN(new_n9586_));
  OAI21_X1   g09522(.A1(new_n2003_), .A2(new_n2005_), .B(new_n1678_), .ZN(new_n9587_));
  NAND3_X1   g09523(.A1(new_n4913_), .A2(new_n2074_), .A3(new_n2004_), .ZN(new_n9588_));
  NAND2_X1   g09524(.A1(new_n9587_), .A2(new_n9588_), .ZN(new_n9589_));
  AOI21_X1   g09525(.A1(new_n9589_), .A2(new_n4914_), .B(new_n2107_), .ZN(new_n9590_));
  NOR2_X1    g09526(.A1(new_n2071_), .A2(new_n9489_), .ZN(new_n9591_));
  NOR2_X1    g09527(.A1(new_n1612_), .A2(new_n9485_), .ZN(new_n9592_));
  NOR2_X1    g09528(.A1(new_n1678_), .A2(new_n9483_), .ZN(new_n9593_));
  NOR4_X1    g09529(.A1(new_n9593_), .A2(new_n9592_), .A3(new_n9591_), .A4(new_n9482_), .ZN(new_n9594_));
  OAI21_X1   g09530(.A1(new_n9586_), .A2(new_n9590_), .B(new_n9594_), .ZN(new_n9595_));
  XOR2_X1    g09531(.A1(new_n9595_), .A2(\a[2] ), .Z(new_n9596_));
  NOR2_X1    g09532(.A1(new_n1612_), .A2(new_n9489_), .ZN(new_n9597_));
  NOR2_X1    g09533(.A1(new_n1764_), .A2(new_n9483_), .ZN(new_n9598_));
  NOR2_X1    g09534(.A1(new_n1729_), .A2(new_n9485_), .ZN(new_n9599_));
  NOR4_X1    g09535(.A1(new_n9598_), .A2(new_n9597_), .A3(new_n9482_), .A4(new_n9599_), .ZN(new_n9600_));
  AOI21_X1   g09536(.A1(new_n4778_), .A2(new_n9600_), .B(new_n4387_), .ZN(new_n9601_));
  NOR2_X1    g09537(.A1(new_n4776_), .A2(new_n1612_), .ZN(new_n9602_));
  AOI21_X1   g09538(.A1(new_n4769_), .A2(new_n4772_), .B(new_n1613_), .ZN(new_n9603_));
  OAI21_X1   g09539(.A1(new_n9602_), .A2(new_n9603_), .B(new_n9600_), .ZN(new_n9604_));
  NOR2_X1    g09540(.A1(new_n9604_), .A2(\a[2] ), .ZN(new_n9605_));
  NOR2_X1    g09541(.A1(new_n9605_), .A2(new_n9601_), .ZN(new_n9606_));
  NOR2_X1    g09542(.A1(new_n1999_), .A2(new_n6833_), .ZN(new_n9607_));
  NOR2_X1    g09543(.A1(new_n1999_), .A2(new_n9485_), .ZN(new_n9608_));
  NAND4_X1   g09544(.A1(new_n4573_), .A2(new_n1812_), .A3(new_n1861_), .A4(new_n9489_), .ZN(new_n9609_));
  NAND4_X1   g09545(.A1(new_n1800_), .A2(new_n1778_), .A3(new_n1812_), .A4(new_n9483_), .ZN(new_n9610_));
  NAND2_X1   g09546(.A1(new_n9609_), .A2(new_n9610_), .ZN(new_n9611_));
  OAI21_X1   g09547(.A1(new_n9611_), .A2(new_n9608_), .B(\a[2] ), .ZN(new_n9612_));
  NOR2_X1    g09548(.A1(new_n9482_), .A2(new_n4387_), .ZN(new_n9613_));
  NAND3_X1   g09549(.A1(new_n1999_), .A2(new_n1813_), .A3(new_n1862_), .ZN(new_n9614_));
  OAI21_X1   g09550(.A1(new_n4766_), .A2(new_n4745_), .B(new_n1939_), .ZN(new_n9615_));
  AOI21_X1   g09551(.A1(new_n9614_), .A2(new_n9615_), .B(new_n9613_), .ZN(new_n9616_));
  INV_X1     g09552(.I(new_n9613_), .ZN(new_n9617_));
  NAND2_X1   g09553(.A1(new_n4766_), .A2(new_n4745_), .ZN(new_n9618_));
  AOI21_X1   g09554(.A1(new_n4877_), .A2(new_n9618_), .B(new_n9617_), .ZN(new_n9619_));
  NOR2_X1    g09555(.A1(new_n6922_), .A2(new_n9488_), .ZN(new_n9620_));
  OAI21_X1   g09556(.A1(new_n1999_), .A2(new_n9620_), .B(\a[2] ), .ZN(new_n9621_));
  NAND3_X1   g09557(.A1(new_n4766_), .A2(\a[2] ), .A3(new_n9503_), .ZN(new_n9622_));
  NAND2_X1   g09558(.A1(new_n9488_), .A2(\a[2] ), .ZN(new_n9623_));
  NAND4_X1   g09559(.A1(new_n9621_), .A2(new_n9622_), .A3(new_n4745_), .A4(new_n9623_), .ZN(new_n9624_));
  NOR3_X1    g09560(.A1(new_n9624_), .A2(new_n9616_), .A3(new_n9619_), .ZN(new_n9625_));
  NAND3_X1   g09561(.A1(new_n9625_), .A2(new_n9607_), .A3(new_n9612_), .ZN(new_n9626_));
  INV_X1     g09562(.I(new_n9626_), .ZN(new_n9627_));
  NOR2_X1    g09563(.A1(new_n4840_), .A2(new_n1729_), .ZN(new_n9628_));
  AOI21_X1   g09564(.A1(new_n4836_), .A2(new_n4833_), .B(new_n1882_), .ZN(new_n9629_));
  NOR2_X1    g09565(.A1(new_n1939_), .A2(new_n9483_), .ZN(new_n9630_));
  NOR2_X1    g09566(.A1(new_n1729_), .A2(new_n9489_), .ZN(new_n9631_));
  NOR2_X1    g09567(.A1(new_n4745_), .A2(new_n9485_), .ZN(new_n9632_));
  NOR4_X1    g09568(.A1(new_n9630_), .A2(new_n9631_), .A3(new_n9632_), .A4(new_n9482_), .ZN(new_n9633_));
  OAI21_X1   g09569(.A1(new_n9628_), .A2(new_n9629_), .B(new_n9633_), .ZN(new_n9634_));
  NAND2_X1   g09570(.A1(new_n9634_), .A2(\a[2] ), .ZN(new_n9635_));
  NAND3_X1   g09571(.A1(new_n4842_), .A2(new_n4387_), .A3(new_n9633_), .ZN(new_n9636_));
  NAND2_X1   g09572(.A1(new_n9635_), .A2(new_n9636_), .ZN(new_n9637_));
  AOI21_X1   g09573(.A1(new_n9625_), .A2(new_n9612_), .B(new_n9607_), .ZN(new_n9638_));
  AOI21_X1   g09574(.A1(new_n9637_), .A2(new_n9638_), .B(new_n9627_), .ZN(new_n9639_));
  AOI22_X1   g09575(.A1(new_n4766_), .A2(new_n8799_), .B1(new_n1813_), .B2(new_n6838_), .ZN(new_n9640_));
  AOI21_X1   g09576(.A1(new_n4981_), .A2(new_n6835_), .B(new_n9640_), .ZN(new_n9641_));
  NAND2_X1   g09577(.A1(new_n9607_), .A2(\a[5] ), .ZN(new_n9642_));
  XOR2_X1    g09578(.A1(new_n9641_), .A2(new_n9642_), .Z(new_n9643_));
  INV_X1     g09579(.I(new_n4804_), .ZN(new_n9644_));
  NAND3_X1   g09580(.A1(new_n4748_), .A2(new_n1729_), .A3(new_n4767_), .ZN(new_n9645_));
  AOI21_X1   g09581(.A1(new_n9645_), .A2(new_n9644_), .B(new_n1763_), .ZN(new_n9646_));
  INV_X1     g09582(.I(new_n4807_), .ZN(new_n9647_));
  OAI21_X1   g09583(.A1(new_n1941_), .A2(new_n2000_), .B(new_n1729_), .ZN(new_n9648_));
  AOI21_X1   g09584(.A1(new_n9648_), .A2(new_n9647_), .B(new_n1764_), .ZN(new_n9649_));
  NOR2_X1    g09585(.A1(new_n1939_), .A2(new_n9485_), .ZN(new_n9650_));
  NOR2_X1    g09586(.A1(new_n1763_), .A2(new_n9488_), .ZN(new_n9651_));
  NOR2_X1    g09587(.A1(new_n1729_), .A2(new_n9483_), .ZN(new_n9652_));
  NOR4_X1    g09588(.A1(new_n9651_), .A2(new_n9482_), .A3(new_n9650_), .A4(new_n9652_), .ZN(new_n9653_));
  OAI21_X1   g09589(.A1(new_n9649_), .A2(new_n9646_), .B(new_n9653_), .ZN(new_n9654_));
  NOR2_X1    g09590(.A1(new_n9654_), .A2(\a[2] ), .ZN(new_n9655_));
  AOI21_X1   g09591(.A1(new_n4810_), .A2(new_n9653_), .B(new_n4387_), .ZN(new_n9656_));
  NOR3_X1    g09592(.A1(new_n9656_), .A2(new_n9655_), .A3(new_n9643_), .ZN(new_n9657_));
  NOR2_X1    g09593(.A1(new_n9657_), .A2(new_n9639_), .ZN(new_n9658_));
  OAI21_X1   g09594(.A1(new_n9656_), .A2(new_n9655_), .B(new_n9643_), .ZN(new_n9659_));
  INV_X1     g09595(.I(new_n9659_), .ZN(new_n9660_));
  NOR3_X1    g09596(.A1(new_n9658_), .A2(new_n9606_), .A3(new_n9660_), .ZN(new_n9661_));
  NAND2_X1   g09597(.A1(new_n9604_), .A2(\a[2] ), .ZN(new_n9662_));
  NAND3_X1   g09598(.A1(new_n4778_), .A2(new_n4387_), .A3(new_n9600_), .ZN(new_n9663_));
  NAND2_X1   g09599(.A1(new_n9662_), .A2(new_n9663_), .ZN(new_n9664_));
  AOI21_X1   g09600(.A1(new_n4842_), .A2(new_n9633_), .B(new_n4387_), .ZN(new_n9665_));
  NOR2_X1    g09601(.A1(new_n9634_), .A2(\a[2] ), .ZN(new_n9666_));
  OAI21_X1   g09602(.A1(new_n9666_), .A2(new_n9665_), .B(new_n9638_), .ZN(new_n9667_));
  NAND2_X1   g09603(.A1(new_n9667_), .A2(new_n9626_), .ZN(new_n9668_));
  XNOR2_X1   g09604(.A1(new_n9641_), .A2(new_n9642_), .ZN(new_n9669_));
  NAND3_X1   g09605(.A1(new_n4810_), .A2(new_n4387_), .A3(new_n9653_), .ZN(new_n9670_));
  NAND2_X1   g09606(.A1(new_n9654_), .A2(\a[2] ), .ZN(new_n9671_));
  NAND3_X1   g09607(.A1(new_n9670_), .A2(new_n9671_), .A3(new_n9669_), .ZN(new_n9672_));
  NAND2_X1   g09608(.A1(new_n9672_), .A2(new_n9668_), .ZN(new_n9673_));
  AOI21_X1   g09609(.A1(new_n9673_), .A2(new_n9659_), .B(new_n9664_), .ZN(new_n9674_));
  INV_X1     g09610(.I(new_n9641_), .ZN(new_n9675_));
  NOR3_X1    g09611(.A1(new_n9675_), .A2(new_n65_), .A3(new_n9607_), .ZN(new_n9676_));
  AOI22_X1   g09612(.A1(new_n4766_), .A2(new_n6846_), .B1(new_n1813_), .B2(new_n8799_), .ZN(new_n9677_));
  AOI21_X1   g09613(.A1(new_n1862_), .A2(new_n6838_), .B(new_n9677_), .ZN(new_n9678_));
  NOR3_X1    g09614(.A1(new_n9678_), .A2(new_n4878_), .A3(new_n6836_), .ZN(new_n9679_));
  XOR2_X1    g09615(.A1(new_n9679_), .A2(\a[5] ), .Z(new_n9680_));
  XOR2_X1    g09616(.A1(new_n9680_), .A2(new_n9676_), .Z(new_n9681_));
  OAI22_X1   g09617(.A1(new_n9674_), .A2(new_n9661_), .B1(new_n9606_), .B2(new_n9681_), .ZN(new_n9682_));
  XOR2_X1    g09618(.A1(new_n9679_), .A2(new_n65_), .Z(new_n9683_));
  NOR2_X1    g09619(.A1(new_n1999_), .A2(new_n6773_), .ZN(new_n9684_));
  OAI22_X1   g09620(.A1(new_n1729_), .A2(new_n6839_), .B1(new_n4745_), .B2(new_n6913_), .ZN(new_n9685_));
  NAND2_X1   g09621(.A1(new_n1862_), .A2(new_n8799_), .ZN(new_n9686_));
  AOI21_X1   g09622(.A1(new_n9685_), .A2(new_n9686_), .B(new_n6836_), .ZN(new_n9687_));
  NAND3_X1   g09623(.A1(new_n4842_), .A2(new_n65_), .A3(new_n9687_), .ZN(new_n9688_));
  AOI21_X1   g09624(.A1(new_n4842_), .A2(new_n9687_), .B(new_n65_), .ZN(new_n9689_));
  INV_X1     g09625(.I(new_n9689_), .ZN(new_n9690_));
  NAND3_X1   g09626(.A1(new_n9690_), .A2(new_n9684_), .A3(new_n9688_), .ZN(new_n9691_));
  INV_X1     g09627(.I(new_n9684_), .ZN(new_n9692_));
  INV_X1     g09628(.I(new_n9688_), .ZN(new_n9693_));
  OAI21_X1   g09629(.A1(new_n9693_), .A2(new_n9689_), .B(new_n9692_), .ZN(new_n9694_));
  AOI22_X1   g09630(.A1(new_n9691_), .A2(new_n9694_), .B1(new_n9676_), .B2(new_n9683_), .ZN(new_n9695_));
  NOR3_X1    g09631(.A1(new_n9693_), .A2(new_n9692_), .A3(new_n9689_), .ZN(new_n9696_));
  AOI21_X1   g09632(.A1(new_n9690_), .A2(new_n9688_), .B(new_n9684_), .ZN(new_n9697_));
  NAND2_X1   g09633(.A1(new_n9683_), .A2(new_n9676_), .ZN(new_n9698_));
  NOR3_X1    g09634(.A1(new_n9698_), .A2(new_n9697_), .A3(new_n9696_), .ZN(new_n9699_));
  NOR2_X1    g09635(.A1(new_n9695_), .A2(new_n9699_), .ZN(new_n9700_));
  OAI22_X1   g09636(.A1(new_n1678_), .A2(new_n9489_), .B1(new_n1764_), .B2(new_n9485_), .ZN(new_n9701_));
  NAND2_X1   g09637(.A1(new_n1613_), .A2(new_n9503_), .ZN(new_n9702_));
  AOI21_X1   g09638(.A1(new_n9701_), .A2(new_n9702_), .B(new_n9482_), .ZN(new_n9703_));
  NAND3_X1   g09639(.A1(new_n4917_), .A2(new_n4387_), .A3(new_n9703_), .ZN(new_n9704_));
  NAND2_X1   g09640(.A1(new_n4917_), .A2(new_n9703_), .ZN(new_n9705_));
  NAND2_X1   g09641(.A1(new_n9705_), .A2(\a[2] ), .ZN(new_n9706_));
  NAND2_X1   g09642(.A1(new_n9706_), .A2(new_n9704_), .ZN(new_n9707_));
  NOR2_X1    g09643(.A1(new_n9707_), .A2(new_n9700_), .ZN(new_n9708_));
  NAND2_X1   g09644(.A1(new_n9707_), .A2(new_n9700_), .ZN(new_n9709_));
  OAI21_X1   g09645(.A1(new_n9682_), .A2(new_n9708_), .B(new_n9709_), .ZN(new_n9710_));
  NAND2_X1   g09646(.A1(new_n9710_), .A2(new_n9596_), .ZN(new_n9711_));
  NOR2_X1    g09647(.A1(new_n9710_), .A2(new_n9596_), .ZN(new_n9712_));
  XOR2_X1    g09648(.A1(new_n9595_), .A2(new_n4387_), .Z(new_n9713_));
  AOI21_X1   g09649(.A1(new_n9673_), .A2(new_n9659_), .B(new_n9664_), .ZN(new_n9714_));
  NAND3_X1   g09650(.A1(new_n9673_), .A2(new_n9664_), .A3(new_n9659_), .ZN(new_n9715_));
  OAI21_X1   g09651(.A1(new_n9658_), .A2(new_n9660_), .B(new_n9606_), .ZN(new_n9716_));
  INV_X1     g09652(.I(new_n9681_), .ZN(new_n9717_));
  AOI21_X1   g09653(.A1(new_n9716_), .A2(new_n9715_), .B(new_n9717_), .ZN(new_n9718_));
  OAI21_X1   g09654(.A1(new_n9696_), .A2(new_n9697_), .B(new_n9698_), .ZN(new_n9719_));
  NAND4_X1   g09655(.A1(new_n9691_), .A2(new_n9694_), .A3(new_n9676_), .A4(new_n9683_), .ZN(new_n9720_));
  NAND2_X1   g09656(.A1(new_n9719_), .A2(new_n9720_), .ZN(new_n9721_));
  NAND3_X1   g09657(.A1(new_n9721_), .A2(new_n9704_), .A3(new_n9706_), .ZN(new_n9722_));
  OAI21_X1   g09658(.A1(new_n9718_), .A2(new_n9714_), .B(new_n9722_), .ZN(new_n9723_));
  AOI21_X1   g09659(.A1(new_n9723_), .A2(new_n9709_), .B(new_n9713_), .ZN(new_n9724_));
  OAI22_X1   g09660(.A1(new_n1764_), .A2(new_n6839_), .B1(new_n1729_), .B2(new_n6843_), .ZN(new_n9725_));
  NAND2_X1   g09661(.A1(new_n1862_), .A2(new_n6846_), .ZN(new_n9726_));
  AOI21_X1   g09662(.A1(new_n9725_), .A2(new_n9726_), .B(new_n6836_), .ZN(new_n9727_));
  NAND2_X1   g09663(.A1(new_n4810_), .A2(new_n9727_), .ZN(new_n9728_));
  XOR2_X1    g09664(.A1(new_n9728_), .A2(\a[5] ), .Z(new_n9729_));
  NAND2_X1   g09665(.A1(new_n1813_), .A2(new_n6784_), .ZN(new_n9730_));
  NAND2_X1   g09666(.A1(new_n4766_), .A2(new_n6789_), .ZN(new_n9731_));
  NAND4_X1   g09667(.A1(new_n4981_), .A2(new_n6775_), .A3(new_n9730_), .A4(new_n9731_), .ZN(new_n9732_));
  XOR2_X1    g09668(.A1(new_n9732_), .A2(\a[8] ), .Z(new_n9733_));
  NAND2_X1   g09669(.A1(new_n9692_), .A2(\a[8] ), .ZN(new_n9734_));
  XOR2_X1    g09670(.A1(new_n9733_), .A2(new_n9734_), .Z(new_n9735_));
  NOR3_X1    g09671(.A1(new_n9697_), .A2(new_n9696_), .A3(new_n9680_), .ZN(new_n9736_));
  NOR3_X1    g09672(.A1(new_n9693_), .A2(new_n9692_), .A3(new_n9689_), .ZN(new_n9737_));
  OAI21_X1   g09673(.A1(new_n9736_), .A2(new_n9676_), .B(new_n9737_), .ZN(new_n9738_));
  INV_X1     g09674(.I(new_n9676_), .ZN(new_n9739_));
  NAND3_X1   g09675(.A1(new_n9691_), .A2(new_n9694_), .A3(new_n9683_), .ZN(new_n9740_));
  INV_X1     g09676(.I(new_n9737_), .ZN(new_n9741_));
  NAND3_X1   g09677(.A1(new_n9740_), .A2(new_n9739_), .A3(new_n9741_), .ZN(new_n9742_));
  NAND3_X1   g09678(.A1(new_n9738_), .A2(new_n9742_), .A3(new_n9735_), .ZN(new_n9743_));
  INV_X1     g09679(.I(new_n9735_), .ZN(new_n9744_));
  AOI21_X1   g09680(.A1(new_n9740_), .A2(new_n9739_), .B(new_n9741_), .ZN(new_n9745_));
  NOR3_X1    g09681(.A1(new_n9736_), .A2(new_n9676_), .A3(new_n9737_), .ZN(new_n9746_));
  OAI21_X1   g09682(.A1(new_n9746_), .A2(new_n9745_), .B(new_n9744_), .ZN(new_n9747_));
  AOI21_X1   g09683(.A1(new_n9747_), .A2(new_n9743_), .B(new_n9729_), .ZN(new_n9748_));
  INV_X1     g09684(.I(new_n9729_), .ZN(new_n9749_));
  NAND3_X1   g09685(.A1(new_n9738_), .A2(new_n9742_), .A3(new_n9744_), .ZN(new_n9750_));
  OAI21_X1   g09686(.A1(new_n9746_), .A2(new_n9745_), .B(new_n9735_), .ZN(new_n9751_));
  AOI21_X1   g09687(.A1(new_n9751_), .A2(new_n9750_), .B(new_n9749_), .ZN(new_n9752_));
  NOR2_X1    g09688(.A1(new_n9748_), .A2(new_n9752_), .ZN(new_n9753_));
  OAI21_X1   g09689(.A1(new_n9712_), .A2(new_n9724_), .B(new_n9753_), .ZN(new_n9754_));
  OAI22_X1   g09690(.A1(new_n2103_), .A2(new_n9489_), .B1(new_n1678_), .B2(new_n9485_), .ZN(new_n9755_));
  NAND2_X1   g09691(.A1(new_n2107_), .A2(new_n9503_), .ZN(new_n9756_));
  AOI21_X1   g09692(.A1(new_n9755_), .A2(new_n9756_), .B(new_n9482_), .ZN(new_n9757_));
  NAND3_X1   g09693(.A1(new_n4545_), .A2(new_n4387_), .A3(new_n9757_), .ZN(new_n9758_));
  OAI21_X1   g09694(.A1(new_n5103_), .A2(new_n5104_), .B(new_n9757_), .ZN(new_n9759_));
  NAND2_X1   g09695(.A1(new_n9759_), .A2(\a[2] ), .ZN(new_n9760_));
  AND2_X2    g09696(.A1(new_n9758_), .A2(new_n9760_), .Z(new_n9761_));
  AOI21_X1   g09697(.A1(new_n9754_), .A2(new_n9711_), .B(new_n9761_), .ZN(new_n9762_));
  NAND3_X1   g09698(.A1(new_n9723_), .A2(new_n9713_), .A3(new_n9709_), .ZN(new_n9763_));
  NAND2_X1   g09699(.A1(new_n9710_), .A2(new_n9596_), .ZN(new_n9764_));
  NOR3_X1    g09700(.A1(new_n9746_), .A2(new_n9745_), .A3(new_n9744_), .ZN(new_n9765_));
  AOI21_X1   g09701(.A1(new_n9738_), .A2(new_n9742_), .B(new_n9735_), .ZN(new_n9766_));
  OAI21_X1   g09702(.A1(new_n9765_), .A2(new_n9766_), .B(new_n9749_), .ZN(new_n9767_));
  NOR3_X1    g09703(.A1(new_n9746_), .A2(new_n9745_), .A3(new_n9735_), .ZN(new_n9768_));
  AOI21_X1   g09704(.A1(new_n9738_), .A2(new_n9742_), .B(new_n9744_), .ZN(new_n9769_));
  OAI21_X1   g09705(.A1(new_n9768_), .A2(new_n9769_), .B(new_n9729_), .ZN(new_n9770_));
  NAND2_X1   g09706(.A1(new_n9767_), .A2(new_n9770_), .ZN(new_n9771_));
  AOI22_X1   g09707(.A1(new_n9764_), .A2(new_n9763_), .B1(new_n9771_), .B2(new_n9713_), .ZN(new_n9772_));
  NAND2_X1   g09708(.A1(new_n9750_), .A2(new_n9749_), .ZN(new_n9773_));
  NAND2_X1   g09709(.A1(new_n4766_), .A2(new_n7530_), .ZN(new_n9774_));
  NAND2_X1   g09710(.A1(new_n1813_), .A2(new_n6789_), .ZN(new_n9775_));
  AOI22_X1   g09711(.A1(new_n9774_), .A2(new_n9775_), .B1(new_n1862_), .B2(new_n6784_), .ZN(new_n9776_));
  NOR3_X1    g09712(.A1(new_n4878_), .A2(new_n9776_), .A3(new_n6776_), .ZN(new_n9777_));
  XOR2_X1    g09713(.A1(new_n9777_), .A2(\a[8] ), .Z(new_n9778_));
  NOR3_X1    g09714(.A1(new_n9732_), .A2(new_n4009_), .A3(new_n9684_), .ZN(new_n9779_));
  XOR2_X1    g09715(.A1(new_n9778_), .A2(new_n9779_), .Z(new_n9780_));
  INV_X1     g09716(.I(new_n9780_), .ZN(new_n9781_));
  OAI22_X1   g09717(.A1(new_n1764_), .A2(new_n6843_), .B1(new_n1729_), .B2(new_n6913_), .ZN(new_n9782_));
  NAND2_X1   g09718(.A1(new_n1613_), .A2(new_n6838_), .ZN(new_n9783_));
  AOI21_X1   g09719(.A1(new_n9783_), .A2(new_n9782_), .B(new_n6836_), .ZN(new_n9784_));
  NAND2_X1   g09720(.A1(new_n4778_), .A2(new_n9784_), .ZN(new_n9785_));
  XOR2_X1    g09721(.A1(new_n9785_), .A2(\a[5] ), .Z(new_n9786_));
  NAND2_X1   g09722(.A1(new_n9786_), .A2(new_n9781_), .ZN(new_n9787_));
  XOR2_X1    g09723(.A1(new_n9785_), .A2(new_n65_), .Z(new_n9788_));
  NAND2_X1   g09724(.A1(new_n9788_), .A2(new_n9780_), .ZN(new_n9789_));
  NAND2_X1   g09725(.A1(new_n9787_), .A2(new_n9789_), .ZN(new_n9790_));
  AOI21_X1   g09726(.A1(new_n9751_), .A2(new_n9773_), .B(new_n9790_), .ZN(new_n9791_));
  NAND2_X1   g09727(.A1(new_n9773_), .A2(new_n9751_), .ZN(new_n9792_));
  NOR2_X1    g09728(.A1(new_n9788_), .A2(new_n9780_), .ZN(new_n9793_));
  NOR2_X1    g09729(.A1(new_n9786_), .A2(new_n9781_), .ZN(new_n9794_));
  NOR2_X1    g09730(.A1(new_n9793_), .A2(new_n9794_), .ZN(new_n9795_));
  NOR2_X1    g09731(.A1(new_n9792_), .A2(new_n9795_), .ZN(new_n9796_));
  OAI21_X1   g09732(.A1(new_n9791_), .A2(new_n9796_), .B(new_n9761_), .ZN(new_n9797_));
  NOR2_X1    g09733(.A1(new_n9797_), .A2(new_n9772_), .ZN(new_n9798_));
  OAI22_X1   g09734(.A1(new_n2103_), .A2(new_n9483_), .B1(new_n2158_), .B2(new_n9489_), .ZN(new_n9799_));
  NAND2_X1   g09735(.A1(new_n2107_), .A2(new_n6925_), .ZN(new_n9800_));
  AOI21_X1   g09736(.A1(new_n9799_), .A2(new_n9800_), .B(new_n9482_), .ZN(new_n9801_));
  NAND2_X1   g09737(.A1(new_n4959_), .A2(new_n9801_), .ZN(new_n9802_));
  XOR2_X1    g09738(.A1(new_n9802_), .A2(\a[2] ), .Z(new_n9803_));
  INV_X1     g09739(.I(new_n9803_), .ZN(new_n9804_));
  OAI21_X1   g09740(.A1(new_n9798_), .A2(new_n9762_), .B(new_n9804_), .ZN(new_n9805_));
  NAND2_X1   g09741(.A1(new_n9758_), .A2(new_n9760_), .ZN(new_n9806_));
  NAND2_X1   g09742(.A1(new_n9772_), .A2(new_n9806_), .ZN(new_n9807_));
  NOR2_X1    g09743(.A1(new_n9768_), .A2(new_n9729_), .ZN(new_n9808_));
  OAI21_X1   g09744(.A1(new_n9769_), .A2(new_n9808_), .B(new_n9795_), .ZN(new_n9809_));
  NAND3_X1   g09745(.A1(new_n9790_), .A2(new_n9773_), .A3(new_n9751_), .ZN(new_n9810_));
  AOI21_X1   g09746(.A1(new_n9809_), .A2(new_n9810_), .B(new_n9806_), .ZN(new_n9811_));
  NAND3_X1   g09747(.A1(new_n9754_), .A2(new_n9711_), .A3(new_n9811_), .ZN(new_n9812_));
  NAND3_X1   g09748(.A1(new_n9807_), .A2(new_n9812_), .A3(new_n9803_), .ZN(new_n9813_));
  NAND2_X1   g09749(.A1(new_n9792_), .A2(new_n9787_), .ZN(new_n9814_));
  NAND2_X1   g09750(.A1(new_n9814_), .A2(new_n9789_), .ZN(new_n9815_));
  OAI22_X1   g09751(.A1(new_n1678_), .A2(new_n6839_), .B1(new_n1764_), .B2(new_n6913_), .ZN(new_n9816_));
  NAND2_X1   g09752(.A1(new_n1613_), .A2(new_n8799_), .ZN(new_n9817_));
  AOI21_X1   g09753(.A1(new_n9816_), .A2(new_n9817_), .B(new_n6836_), .ZN(new_n9818_));
  NAND2_X1   g09754(.A1(new_n4917_), .A2(new_n9818_), .ZN(new_n9819_));
  XOR2_X1    g09755(.A1(new_n9819_), .A2(\a[5] ), .Z(new_n9820_));
  INV_X1     g09756(.I(new_n9820_), .ZN(new_n9821_));
  INV_X1     g09757(.I(new_n9777_), .ZN(new_n9822_));
  NOR4_X1    g09758(.A1(new_n9822_), .A2(new_n4009_), .A3(new_n9684_), .A4(new_n9732_), .ZN(new_n9823_));
  INV_X1     g09759(.I(new_n9823_), .ZN(new_n9824_));
  NOR2_X1    g09760(.A1(new_n1999_), .A2(new_n4704_), .ZN(new_n9825_));
  INV_X1     g09761(.I(new_n9825_), .ZN(new_n9826_));
  OAI22_X1   g09762(.A1(new_n1729_), .A2(new_n6785_), .B1(new_n4745_), .B2(new_n6783_), .ZN(new_n9827_));
  NAND2_X1   g09763(.A1(new_n1862_), .A2(new_n6789_), .ZN(new_n9828_));
  AOI21_X1   g09764(.A1(new_n9827_), .A2(new_n9828_), .B(new_n6776_), .ZN(new_n9829_));
  NAND2_X1   g09765(.A1(new_n4842_), .A2(new_n9829_), .ZN(new_n9830_));
  XOR2_X1    g09766(.A1(new_n9830_), .A2(\a[8] ), .Z(new_n9831_));
  XOR2_X1    g09767(.A1(new_n9831_), .A2(new_n9826_), .Z(new_n9832_));
  NAND2_X1   g09768(.A1(new_n9832_), .A2(new_n9824_), .ZN(new_n9833_));
  XOR2_X1    g09769(.A1(new_n9831_), .A2(new_n9825_), .Z(new_n9834_));
  NAND2_X1   g09770(.A1(new_n9834_), .A2(new_n9823_), .ZN(new_n9835_));
  NAND2_X1   g09771(.A1(new_n9835_), .A2(new_n9833_), .ZN(new_n9836_));
  XOR2_X1    g09772(.A1(new_n9836_), .A2(new_n9821_), .Z(new_n9837_));
  XOR2_X1    g09773(.A1(new_n9815_), .A2(new_n9837_), .Z(new_n9838_));
  NAND2_X1   g09774(.A1(new_n9813_), .A2(new_n9838_), .ZN(new_n9839_));
  NOR2_X1    g09775(.A1(new_n9836_), .A2(new_n9821_), .ZN(new_n9840_));
  AOI21_X1   g09776(.A1(new_n9814_), .A2(new_n9789_), .B(new_n9840_), .ZN(new_n9841_));
  AOI21_X1   g09777(.A1(new_n9833_), .A2(new_n9835_), .B(new_n9820_), .ZN(new_n9842_));
  XOR2_X1    g09778(.A1(new_n9823_), .A2(new_n9825_), .Z(new_n9843_));
  NAND2_X1   g09779(.A1(new_n9843_), .A2(new_n9831_), .ZN(new_n9844_));
  NAND2_X1   g09780(.A1(new_n9823_), .A2(new_n9825_), .ZN(new_n9845_));
  NAND2_X1   g09781(.A1(new_n1813_), .A2(new_n4709_), .ZN(new_n9846_));
  NAND2_X1   g09782(.A1(new_n4766_), .A2(new_n4720_), .ZN(new_n9847_));
  NAND4_X1   g09783(.A1(new_n4981_), .A2(new_n4706_), .A3(new_n9846_), .A4(new_n9847_), .ZN(new_n9848_));
  XOR2_X1    g09784(.A1(new_n9848_), .A2(new_n4034_), .Z(new_n9849_));
  NOR2_X1    g09785(.A1(new_n9825_), .A2(new_n4034_), .ZN(new_n9850_));
  XOR2_X1    g09786(.A1(new_n9849_), .A2(new_n9850_), .Z(new_n9851_));
  INV_X1     g09787(.I(new_n9851_), .ZN(new_n9852_));
  AOI21_X1   g09788(.A1(new_n9844_), .A2(new_n9845_), .B(new_n9852_), .ZN(new_n9853_));
  INV_X1     g09789(.I(new_n9831_), .ZN(new_n9854_));
  XOR2_X1    g09790(.A1(new_n9823_), .A2(new_n9826_), .Z(new_n9855_));
  OAI21_X1   g09791(.A1(new_n9855_), .A2(new_n9854_), .B(new_n9845_), .ZN(new_n9856_));
  NOR2_X1    g09792(.A1(new_n9856_), .A2(new_n9851_), .ZN(new_n9857_));
  OAI22_X1   g09793(.A1(new_n1764_), .A2(new_n6785_), .B1(new_n1729_), .B2(new_n6788_), .ZN(new_n9858_));
  NAND2_X1   g09794(.A1(new_n1862_), .A2(new_n7530_), .ZN(new_n9859_));
  AOI21_X1   g09795(.A1(new_n9858_), .A2(new_n9859_), .B(new_n6776_), .ZN(new_n9860_));
  NAND2_X1   g09796(.A1(new_n4810_), .A2(new_n9860_), .ZN(new_n9861_));
  XOR2_X1    g09797(.A1(new_n9861_), .A2(\a[8] ), .Z(new_n9862_));
  OAI21_X1   g09798(.A1(new_n9857_), .A2(new_n9853_), .B(new_n9862_), .ZN(new_n9863_));
  NAND2_X1   g09799(.A1(new_n9856_), .A2(new_n9851_), .ZN(new_n9864_));
  NAND3_X1   g09800(.A1(new_n9844_), .A2(new_n9852_), .A3(new_n9845_), .ZN(new_n9865_));
  INV_X1     g09801(.I(new_n9862_), .ZN(new_n9866_));
  NAND3_X1   g09802(.A1(new_n9864_), .A2(new_n9865_), .A3(new_n9866_), .ZN(new_n9867_));
  NAND2_X1   g09803(.A1(new_n9863_), .A2(new_n9867_), .ZN(new_n9868_));
  OAI22_X1   g09804(.A1(new_n1678_), .A2(new_n6843_), .B1(new_n2071_), .B2(new_n6839_), .ZN(new_n9869_));
  NAND2_X1   g09805(.A1(new_n1613_), .A2(new_n6846_), .ZN(new_n9870_));
  AOI21_X1   g09806(.A1(new_n9869_), .A2(new_n9870_), .B(new_n6836_), .ZN(new_n9871_));
  NAND2_X1   g09807(.A1(new_n5070_), .A2(new_n9871_), .ZN(new_n9872_));
  XOR2_X1    g09808(.A1(new_n9872_), .A2(new_n65_), .Z(new_n9873_));
  NOR2_X1    g09809(.A1(new_n9873_), .A2(new_n9868_), .ZN(new_n9874_));
  AOI21_X1   g09810(.A1(new_n9864_), .A2(new_n9865_), .B(new_n9866_), .ZN(new_n9875_));
  NOR3_X1    g09811(.A1(new_n9857_), .A2(new_n9853_), .A3(new_n9862_), .ZN(new_n9876_));
  NOR2_X1    g09812(.A1(new_n9876_), .A2(new_n9875_), .ZN(new_n9877_));
  XOR2_X1    g09813(.A1(new_n9872_), .A2(\a[5] ), .Z(new_n9878_));
  NOR2_X1    g09814(.A1(new_n9878_), .A2(new_n9877_), .ZN(new_n9879_));
  OAI22_X1   g09815(.A1(new_n9841_), .A2(new_n9842_), .B1(new_n9874_), .B2(new_n9879_), .ZN(new_n9880_));
  NOR2_X1    g09816(.A1(new_n9841_), .A2(new_n9842_), .ZN(new_n9881_));
  NAND2_X1   g09817(.A1(new_n9878_), .A2(new_n9868_), .ZN(new_n9882_));
  NAND2_X1   g09818(.A1(new_n9873_), .A2(new_n9877_), .ZN(new_n9883_));
  NAND2_X1   g09819(.A1(new_n9882_), .A2(new_n9883_), .ZN(new_n9884_));
  NAND2_X1   g09820(.A1(new_n9881_), .A2(new_n9884_), .ZN(new_n9885_));
  OAI22_X1   g09821(.A1(new_n2103_), .A2(new_n9485_), .B1(new_n2198_), .B2(new_n9489_), .ZN(new_n9886_));
  NAND2_X1   g09822(.A1(new_n2161_), .A2(new_n9503_), .ZN(new_n9887_));
  AOI21_X1   g09823(.A1(new_n9886_), .A2(new_n9887_), .B(new_n9482_), .ZN(new_n9888_));
  NAND3_X1   g09824(.A1(new_n5351_), .A2(new_n4387_), .A3(new_n9888_), .ZN(new_n9889_));
  NAND2_X1   g09825(.A1(new_n5351_), .A2(new_n9888_), .ZN(new_n9890_));
  NAND2_X1   g09826(.A1(new_n9890_), .A2(\a[2] ), .ZN(new_n9891_));
  NAND2_X1   g09827(.A1(new_n9891_), .A2(new_n9889_), .ZN(new_n9892_));
  AOI21_X1   g09828(.A1(new_n9885_), .A2(new_n9880_), .B(new_n9892_), .ZN(new_n9893_));
  AOI21_X1   g09829(.A1(new_n9839_), .A2(new_n9805_), .B(new_n9893_), .ZN(new_n9894_));
  INV_X1     g09830(.I(new_n9880_), .ZN(new_n9895_));
  NOR2_X1    g09831(.A1(new_n9873_), .A2(new_n9877_), .ZN(new_n9896_));
  NOR2_X1    g09832(.A1(new_n9878_), .A2(new_n9868_), .ZN(new_n9897_));
  NOR2_X1    g09833(.A1(new_n9896_), .A2(new_n9897_), .ZN(new_n9898_));
  NOR3_X1    g09834(.A1(new_n9898_), .A2(new_n9841_), .A3(new_n9842_), .ZN(new_n9899_));
  INV_X1     g09835(.I(new_n9892_), .ZN(new_n9900_));
  NOR3_X1    g09836(.A1(new_n9895_), .A2(new_n9900_), .A3(new_n9899_), .ZN(new_n9901_));
  NOR3_X1    g09837(.A1(new_n9894_), .A2(new_n9585_), .A3(new_n9901_), .ZN(new_n9902_));
  INV_X1     g09838(.I(new_n9585_), .ZN(new_n9903_));
  INV_X1     g09839(.I(new_n9805_), .ZN(new_n9904_));
  NOR3_X1    g09840(.A1(new_n9798_), .A2(new_n9762_), .A3(new_n9804_), .ZN(new_n9905_));
  XNOR2_X1   g09841(.A1(new_n9815_), .A2(new_n9837_), .ZN(new_n9906_));
  NOR2_X1    g09842(.A1(new_n9905_), .A2(new_n9906_), .ZN(new_n9907_));
  OAI21_X1   g09843(.A1(new_n9895_), .A2(new_n9899_), .B(new_n9900_), .ZN(new_n9908_));
  OAI21_X1   g09844(.A1(new_n9907_), .A2(new_n9904_), .B(new_n9908_), .ZN(new_n9909_));
  INV_X1     g09845(.I(new_n9901_), .ZN(new_n9910_));
  AOI21_X1   g09846(.A1(new_n9909_), .A2(new_n9910_), .B(new_n9903_), .ZN(new_n9911_));
  OAI21_X1   g09847(.A1(new_n9841_), .A2(new_n9842_), .B(new_n9882_), .ZN(new_n9912_));
  NAND2_X1   g09848(.A1(new_n9912_), .A2(new_n9883_), .ZN(new_n9913_));
  OAI22_X1   g09849(.A1(new_n2103_), .A2(new_n6839_), .B1(new_n1678_), .B2(new_n6913_), .ZN(new_n9914_));
  NAND2_X1   g09850(.A1(new_n2107_), .A2(new_n8799_), .ZN(new_n9915_));
  AOI21_X1   g09851(.A1(new_n9914_), .A2(new_n9915_), .B(new_n6836_), .ZN(new_n9916_));
  NAND2_X1   g09852(.A1(new_n4545_), .A2(new_n9916_), .ZN(new_n9917_));
  XOR2_X1    g09853(.A1(new_n9917_), .A2(\a[5] ), .Z(new_n9918_));
  INV_X1     g09854(.I(new_n9918_), .ZN(new_n9919_));
  NOR2_X1    g09855(.A1(new_n9856_), .A2(new_n9851_), .ZN(new_n9920_));
  NOR2_X1    g09856(.A1(new_n9875_), .A2(new_n9920_), .ZN(new_n9921_));
  AOI22_X1   g09857(.A1(new_n4766_), .A2(new_n6480_), .B1(new_n1813_), .B2(new_n4720_), .ZN(new_n9922_));
  AOI21_X1   g09858(.A1(new_n1862_), .A2(new_n4709_), .B(new_n9922_), .ZN(new_n9923_));
  NOR3_X1    g09859(.A1(new_n9923_), .A2(new_n4878_), .A3(new_n4707_), .ZN(new_n9924_));
  XOR2_X1    g09860(.A1(new_n9924_), .A2(\a[11] ), .Z(new_n9925_));
  NOR3_X1    g09861(.A1(new_n9848_), .A2(new_n4034_), .A3(new_n9825_), .ZN(new_n9926_));
  XOR2_X1    g09862(.A1(new_n9925_), .A2(new_n9926_), .Z(new_n9927_));
  OAI22_X1   g09863(.A1(new_n1764_), .A2(new_n6788_), .B1(new_n1729_), .B2(new_n6783_), .ZN(new_n9928_));
  NAND2_X1   g09864(.A1(new_n1613_), .A2(new_n6784_), .ZN(new_n9929_));
  AOI21_X1   g09865(.A1(new_n9929_), .A2(new_n9928_), .B(new_n6776_), .ZN(new_n9930_));
  NAND2_X1   g09866(.A1(new_n4778_), .A2(new_n9930_), .ZN(new_n9931_));
  XOR2_X1    g09867(.A1(new_n9931_), .A2(\a[8] ), .Z(new_n9932_));
  XOR2_X1    g09868(.A1(new_n9932_), .A2(new_n9927_), .Z(new_n9933_));
  NOR2_X1    g09869(.A1(new_n9921_), .A2(new_n9933_), .ZN(new_n9934_));
  INV_X1     g09870(.I(new_n9927_), .ZN(new_n9935_));
  NAND2_X1   g09871(.A1(new_n9932_), .A2(new_n9935_), .ZN(new_n9936_));
  NOR2_X1    g09872(.A1(new_n9932_), .A2(new_n9935_), .ZN(new_n9937_));
  INV_X1     g09873(.I(new_n9937_), .ZN(new_n9938_));
  NAND2_X1   g09874(.A1(new_n9938_), .A2(new_n9936_), .ZN(new_n9939_));
  AOI21_X1   g09875(.A1(new_n9921_), .A2(new_n9939_), .B(new_n9934_), .ZN(new_n9940_));
  XOR2_X1    g09876(.A1(new_n9940_), .A2(new_n9919_), .Z(new_n9941_));
  NOR2_X1    g09877(.A1(new_n9940_), .A2(new_n9919_), .ZN(new_n9942_));
  INV_X1     g09878(.I(new_n9940_), .ZN(new_n9943_));
  NOR2_X1    g09879(.A1(new_n9943_), .A2(new_n9918_), .ZN(new_n9944_));
  NOR2_X1    g09880(.A1(new_n9944_), .A2(new_n9942_), .ZN(new_n9945_));
  NOR2_X1    g09881(.A1(new_n9945_), .A2(new_n9913_), .ZN(new_n9946_));
  AOI21_X1   g09882(.A1(new_n9913_), .A2(new_n9941_), .B(new_n9946_), .ZN(new_n9947_));
  OAI22_X1   g09883(.A1(new_n9911_), .A2(new_n9902_), .B1(new_n9947_), .B2(new_n9585_), .ZN(new_n9948_));
  NOR2_X1    g09884(.A1(new_n1999_), .A2(new_n6079_), .ZN(new_n9949_));
  INV_X1     g09885(.I(new_n9949_), .ZN(new_n9950_));
  XOR2_X1    g09886(.A1(new_n9924_), .A2(new_n4034_), .Z(new_n9951_));
  NAND2_X1   g09887(.A1(new_n9951_), .A2(new_n9926_), .ZN(new_n9952_));
  NAND2_X1   g09888(.A1(new_n9952_), .A2(new_n9950_), .ZN(new_n9953_));
  NAND3_X1   g09889(.A1(new_n9951_), .A2(new_n9926_), .A3(new_n9949_), .ZN(new_n9954_));
  OAI22_X1   g09890(.A1(new_n1729_), .A2(new_n4710_), .B1(new_n4745_), .B2(new_n4716_), .ZN(new_n9955_));
  NAND2_X1   g09891(.A1(new_n1862_), .A2(new_n4720_), .ZN(new_n9956_));
  AOI21_X1   g09892(.A1(new_n9955_), .A2(new_n9956_), .B(new_n4707_), .ZN(new_n9957_));
  NAND2_X1   g09893(.A1(new_n4842_), .A2(new_n9957_), .ZN(new_n9958_));
  XOR2_X1    g09894(.A1(new_n9958_), .A2(\a[11] ), .Z(new_n9959_));
  NAND3_X1   g09895(.A1(new_n9953_), .A2(new_n9954_), .A3(new_n9959_), .ZN(new_n9960_));
  NAND2_X1   g09896(.A1(new_n9953_), .A2(new_n9954_), .ZN(new_n9961_));
  INV_X1     g09897(.I(new_n9959_), .ZN(new_n9962_));
  NAND2_X1   g09898(.A1(new_n9961_), .A2(new_n9962_), .ZN(new_n9963_));
  NAND2_X1   g09899(.A1(new_n9963_), .A2(new_n9960_), .ZN(new_n9964_));
  OAI22_X1   g09900(.A1(new_n1678_), .A2(new_n6785_), .B1(new_n1764_), .B2(new_n6783_), .ZN(new_n9965_));
  NAND2_X1   g09901(.A1(new_n1613_), .A2(new_n6789_), .ZN(new_n9966_));
  AOI21_X1   g09902(.A1(new_n9965_), .A2(new_n9966_), .B(new_n6776_), .ZN(new_n9967_));
  NAND2_X1   g09903(.A1(new_n4917_), .A2(new_n9967_), .ZN(new_n9968_));
  XOR2_X1    g09904(.A1(new_n9968_), .A2(\a[8] ), .Z(new_n9969_));
  XOR2_X1    g09905(.A1(new_n9964_), .A2(new_n9969_), .Z(new_n9970_));
  OAI21_X1   g09906(.A1(new_n9856_), .A2(new_n9851_), .B(new_n9863_), .ZN(new_n9971_));
  AOI21_X1   g09907(.A1(new_n9971_), .A2(new_n9936_), .B(new_n9937_), .ZN(new_n9972_));
  OAI22_X1   g09908(.A1(new_n2103_), .A2(new_n6843_), .B1(new_n2158_), .B2(new_n6839_), .ZN(new_n9973_));
  NAND2_X1   g09909(.A1(new_n2107_), .A2(new_n6846_), .ZN(new_n9974_));
  AOI21_X1   g09910(.A1(new_n9973_), .A2(new_n9974_), .B(new_n6836_), .ZN(new_n9975_));
  NAND2_X1   g09911(.A1(new_n4959_), .A2(new_n9975_), .ZN(new_n9976_));
  XOR2_X1    g09912(.A1(new_n9976_), .A2(new_n65_), .Z(new_n9977_));
  NAND2_X1   g09913(.A1(new_n9977_), .A2(new_n9972_), .ZN(new_n9978_));
  INV_X1     g09914(.I(new_n9972_), .ZN(new_n9979_));
  XOR2_X1    g09915(.A1(new_n9976_), .A2(\a[5] ), .Z(new_n9980_));
  NAND2_X1   g09916(.A1(new_n9979_), .A2(new_n9980_), .ZN(new_n9981_));
  AOI21_X1   g09917(.A1(new_n9981_), .A2(new_n9978_), .B(new_n9970_), .ZN(new_n9982_));
  XOR2_X1    g09918(.A1(new_n9977_), .A2(new_n9972_), .Z(new_n9983_));
  AOI21_X1   g09919(.A1(new_n9983_), .A2(new_n9970_), .B(new_n9982_), .ZN(new_n9984_));
  NOR2_X1    g09920(.A1(new_n9913_), .A2(new_n9940_), .ZN(new_n9985_));
  INV_X1     g09921(.I(new_n9985_), .ZN(new_n9986_));
  NAND3_X1   g09922(.A1(new_n9984_), .A2(new_n9986_), .A3(new_n9919_), .ZN(new_n9987_));
  INV_X1     g09923(.I(new_n9970_), .ZN(new_n9988_));
  INV_X1     g09924(.I(new_n9978_), .ZN(new_n9989_));
  NOR2_X1    g09925(.A1(new_n9977_), .A2(new_n9972_), .ZN(new_n9990_));
  OAI21_X1   g09926(.A1(new_n9989_), .A2(new_n9990_), .B(new_n9988_), .ZN(new_n9991_));
  XOR2_X1    g09927(.A1(new_n9980_), .A2(new_n9972_), .Z(new_n9992_));
  OAI21_X1   g09928(.A1(new_n9992_), .A2(new_n9988_), .B(new_n9991_), .ZN(new_n9993_));
  OAI21_X1   g09929(.A1(new_n9918_), .A2(new_n9985_), .B(new_n9993_), .ZN(new_n9994_));
  OAI22_X1   g09930(.A1(new_n4365_), .A2(new_n9489_), .B1(new_n2198_), .B2(new_n9485_), .ZN(new_n9995_));
  NAND2_X1   g09931(.A1(new_n1504_), .A2(new_n9503_), .ZN(new_n9996_));
  AOI21_X1   g09932(.A1(new_n9995_), .A2(new_n9996_), .B(new_n9482_), .ZN(new_n9997_));
  NAND2_X1   g09933(.A1(new_n4363_), .A2(new_n9997_), .ZN(new_n9998_));
  XOR2_X1    g09934(.A1(new_n9998_), .A2(\a[2] ), .Z(new_n9999_));
  INV_X1     g09935(.I(new_n9999_), .ZN(new_n10000_));
  AOI21_X1   g09936(.A1(new_n9994_), .A2(new_n9987_), .B(new_n10000_), .ZN(new_n10001_));
  NAND3_X1   g09937(.A1(new_n9994_), .A2(new_n9987_), .A3(new_n10000_), .ZN(new_n10002_));
  OAI21_X1   g09938(.A1(new_n9948_), .A2(new_n10001_), .B(new_n10002_), .ZN(new_n10003_));
  NOR2_X1    g09939(.A1(new_n10003_), .A2(new_n9579_), .ZN(new_n10004_));
  INV_X1     g09940(.I(new_n9579_), .ZN(new_n10005_));
  NAND3_X1   g09941(.A1(new_n9909_), .A2(new_n9903_), .A3(new_n9910_), .ZN(new_n10006_));
  OAI21_X1   g09942(.A1(new_n9894_), .A2(new_n9901_), .B(new_n9585_), .ZN(new_n10007_));
  NAND2_X1   g09943(.A1(new_n9941_), .A2(new_n9913_), .ZN(new_n10008_));
  OAI21_X1   g09944(.A1(new_n9913_), .A2(new_n9945_), .B(new_n10008_), .ZN(new_n10009_));
  AOI22_X1   g09945(.A1(new_n10006_), .A2(new_n10007_), .B1(new_n9903_), .B2(new_n10009_), .ZN(new_n10010_));
  NOR3_X1    g09946(.A1(new_n9993_), .A2(new_n9918_), .A3(new_n9985_), .ZN(new_n10011_));
  AOI21_X1   g09947(.A1(new_n9986_), .A2(new_n9919_), .B(new_n9984_), .ZN(new_n10012_));
  OAI21_X1   g09948(.A1(new_n10011_), .A2(new_n10012_), .B(new_n9999_), .ZN(new_n10013_));
  NAND2_X1   g09949(.A1(new_n10010_), .A2(new_n10013_), .ZN(new_n10014_));
  AOI21_X1   g09950(.A1(new_n10014_), .A2(new_n10002_), .B(new_n10005_), .ZN(new_n10015_));
  NAND2_X1   g09951(.A1(new_n9960_), .A2(new_n9954_), .ZN(new_n10016_));
  NAND2_X1   g09952(.A1(new_n1813_), .A2(new_n6090_), .ZN(new_n10017_));
  NAND2_X1   g09953(.A1(new_n4766_), .A2(new_n6095_), .ZN(new_n10018_));
  NAND4_X1   g09954(.A1(new_n4981_), .A2(new_n6081_), .A3(new_n10017_), .A4(new_n10018_), .ZN(new_n10019_));
  XOR2_X1    g09955(.A1(new_n10019_), .A2(\a[14] ), .Z(new_n10020_));
  NOR2_X1    g09956(.A1(new_n9949_), .A2(new_n3521_), .ZN(new_n10021_));
  INV_X1     g09957(.I(new_n10021_), .ZN(new_n10022_));
  XOR2_X1    g09958(.A1(new_n10020_), .A2(new_n10022_), .Z(new_n10023_));
  NAND2_X1   g09959(.A1(new_n10016_), .A2(new_n10023_), .ZN(new_n10024_));
  INV_X1     g09960(.I(new_n10023_), .ZN(new_n10025_));
  NAND3_X1   g09961(.A1(new_n9960_), .A2(new_n9954_), .A3(new_n10025_), .ZN(new_n10026_));
  OAI22_X1   g09962(.A1(new_n1764_), .A2(new_n4710_), .B1(new_n1729_), .B2(new_n4719_), .ZN(new_n10027_));
  NAND2_X1   g09963(.A1(new_n1862_), .A2(new_n6480_), .ZN(new_n10028_));
  AOI21_X1   g09964(.A1(new_n10027_), .A2(new_n10028_), .B(new_n4707_), .ZN(new_n10029_));
  NAND2_X1   g09965(.A1(new_n4810_), .A2(new_n10029_), .ZN(new_n10030_));
  XOR2_X1    g09966(.A1(new_n10030_), .A2(\a[11] ), .Z(new_n10031_));
  INV_X1     g09967(.I(new_n10031_), .ZN(new_n10032_));
  AOI21_X1   g09968(.A1(new_n10024_), .A2(new_n10026_), .B(new_n10032_), .ZN(new_n10033_));
  AND3_X2    g09969(.A1(new_n10024_), .A2(new_n10026_), .A3(new_n10032_), .Z(new_n10034_));
  NOR2_X1    g09970(.A1(new_n10034_), .A2(new_n10033_), .ZN(new_n10035_));
  NAND3_X1   g09971(.A1(new_n9969_), .A2(new_n9963_), .A3(new_n9960_), .ZN(new_n10036_));
  OAI21_X1   g09972(.A1(new_n9979_), .A2(new_n9970_), .B(new_n10036_), .ZN(new_n10037_));
  OAI22_X1   g09973(.A1(new_n1678_), .A2(new_n6788_), .B1(new_n2071_), .B2(new_n6785_), .ZN(new_n10038_));
  NAND2_X1   g09974(.A1(new_n1613_), .A2(new_n7530_), .ZN(new_n10039_));
  AOI21_X1   g09975(.A1(new_n10038_), .A2(new_n10039_), .B(new_n6776_), .ZN(new_n10040_));
  NAND2_X1   g09976(.A1(new_n5070_), .A2(new_n10040_), .ZN(new_n10041_));
  XOR2_X1    g09977(.A1(new_n10041_), .A2(\a[8] ), .Z(new_n10042_));
  XOR2_X1    g09978(.A1(new_n10037_), .A2(new_n10042_), .Z(new_n10043_));
  XOR2_X1    g09979(.A1(new_n10043_), .A2(new_n10035_), .Z(new_n10044_));
  INV_X1     g09980(.I(new_n9942_), .ZN(new_n10045_));
  NOR2_X1    g09981(.A1(new_n9913_), .A2(new_n10045_), .ZN(new_n10046_));
  NOR2_X1    g09982(.A1(new_n9992_), .A2(new_n9988_), .ZN(new_n10047_));
  XOR2_X1    g09983(.A1(new_n9972_), .A2(new_n9970_), .Z(new_n10048_));
  OAI21_X1   g09984(.A1(new_n10048_), .A2(new_n9977_), .B(new_n10045_), .ZN(new_n10049_));
  OR3_X2     g09985(.A1(new_n10047_), .A2(new_n10049_), .A3(new_n9982_), .Z(new_n10050_));
  OAI22_X1   g09986(.A1(new_n2103_), .A2(new_n6913_), .B1(new_n2198_), .B2(new_n6839_), .ZN(new_n10051_));
  NAND2_X1   g09987(.A1(new_n2161_), .A2(new_n8799_), .ZN(new_n10052_));
  AOI21_X1   g09988(.A1(new_n10051_), .A2(new_n10052_), .B(new_n6836_), .ZN(new_n10053_));
  NAND2_X1   g09989(.A1(new_n5351_), .A2(new_n10053_), .ZN(new_n10054_));
  XOR2_X1    g09990(.A1(new_n10054_), .A2(\a[5] ), .Z(new_n10055_));
  OAI21_X1   g09991(.A1(new_n10050_), .A2(new_n10046_), .B(new_n10055_), .ZN(new_n10056_));
  INV_X1     g09992(.I(new_n10046_), .ZN(new_n10057_));
  NOR2_X1    g09993(.A1(new_n9993_), .A2(new_n10049_), .ZN(new_n10058_));
  INV_X1     g09994(.I(new_n10055_), .ZN(new_n10059_));
  NAND3_X1   g09995(.A1(new_n10058_), .A2(new_n10057_), .A3(new_n10059_), .ZN(new_n10060_));
  AOI21_X1   g09996(.A1(new_n10056_), .A2(new_n10060_), .B(new_n10044_), .ZN(new_n10061_));
  XNOR2_X1   g09997(.A1(new_n10043_), .A2(new_n10035_), .ZN(new_n10062_));
  AOI21_X1   g09998(.A1(new_n10058_), .A2(new_n10057_), .B(new_n10059_), .ZN(new_n10063_));
  NOR3_X1    g09999(.A1(new_n10050_), .A2(new_n10046_), .A3(new_n10055_), .ZN(new_n10064_));
  NOR3_X1    g10000(.A1(new_n10063_), .A2(new_n10064_), .A3(new_n10062_), .ZN(new_n10065_));
  NOR2_X1    g10001(.A1(new_n10065_), .A2(new_n10061_), .ZN(new_n10066_));
  OAI22_X1   g10002(.A1(new_n10004_), .A2(new_n10015_), .B1(new_n9579_), .B2(new_n10066_), .ZN(new_n10067_));
  OAI22_X1   g10003(.A1(new_n2158_), .A2(new_n6913_), .B1(new_n2198_), .B2(new_n6843_), .ZN(new_n10068_));
  OAI21_X1   g10004(.A1(new_n1503_), .A2(new_n6839_), .B(new_n10068_), .ZN(new_n10069_));
  AOI21_X1   g10005(.A1(new_n4620_), .A2(new_n6835_), .B(new_n10069_), .ZN(new_n10070_));
  AOI22_X1   g10006(.A1(new_n10024_), .A2(new_n10026_), .B1(new_n10016_), .B2(new_n10032_), .ZN(new_n10071_));
  OAI22_X1   g10007(.A1(new_n1764_), .A2(new_n4719_), .B1(new_n1729_), .B2(new_n4716_), .ZN(new_n10072_));
  NAND2_X1   g10008(.A1(new_n1613_), .A2(new_n4709_), .ZN(new_n10073_));
  AOI21_X1   g10009(.A1(new_n10073_), .A2(new_n10072_), .B(new_n4707_), .ZN(new_n10074_));
  NAND2_X1   g10010(.A1(new_n4778_), .A2(new_n10074_), .ZN(new_n10075_));
  XOR2_X1    g10011(.A1(new_n10075_), .A2(\a[11] ), .Z(new_n10076_));
  AOI22_X1   g10012(.A1(new_n4766_), .A2(new_n6180_), .B1(new_n1813_), .B2(new_n6095_), .ZN(new_n10077_));
  AOI21_X1   g10013(.A1(new_n1862_), .A2(new_n6090_), .B(new_n10077_), .ZN(new_n10078_));
  NOR3_X1    g10014(.A1(new_n10078_), .A2(new_n4878_), .A3(new_n6082_), .ZN(new_n10079_));
  XOR2_X1    g10015(.A1(new_n10079_), .A2(new_n3521_), .Z(new_n10080_));
  NOR3_X1    g10016(.A1(new_n10019_), .A2(new_n3521_), .A3(new_n9949_), .ZN(new_n10081_));
  XNOR2_X1   g10017(.A1(new_n10080_), .A2(new_n10081_), .ZN(new_n10082_));
  INV_X1     g10018(.I(new_n10082_), .ZN(new_n10083_));
  NAND2_X1   g10019(.A1(new_n10083_), .A2(new_n10076_), .ZN(new_n10084_));
  INV_X1     g10020(.I(new_n10084_), .ZN(new_n10085_));
  NOR2_X1    g10021(.A1(new_n10083_), .A2(new_n10076_), .ZN(new_n10086_));
  NOR2_X1    g10022(.A1(new_n10085_), .A2(new_n10086_), .ZN(new_n10087_));
  NOR2_X1    g10023(.A1(new_n10071_), .A2(new_n10087_), .ZN(new_n10088_));
  NAND2_X1   g10024(.A1(new_n10071_), .A2(new_n10087_), .ZN(new_n10089_));
  INV_X1     g10025(.I(new_n10089_), .ZN(new_n10090_));
  NOR2_X1    g10026(.A1(new_n10090_), .A2(new_n10088_), .ZN(new_n10091_));
  OAI22_X1   g10027(.A1(new_n2103_), .A2(new_n6785_), .B1(new_n1678_), .B2(new_n6783_), .ZN(new_n10092_));
  NAND2_X1   g10028(.A1(new_n2107_), .A2(new_n6789_), .ZN(new_n10093_));
  AOI21_X1   g10029(.A1(new_n10092_), .A2(new_n10093_), .B(new_n6776_), .ZN(new_n10094_));
  NAND2_X1   g10030(.A1(new_n4545_), .A2(new_n10094_), .ZN(new_n10095_));
  XOR2_X1    g10031(.A1(new_n10095_), .A2(\a[8] ), .Z(new_n10096_));
  XOR2_X1    g10032(.A1(new_n10091_), .A2(new_n10096_), .Z(new_n10097_));
  XOR2_X1    g10033(.A1(new_n10097_), .A2(\a[5] ), .Z(new_n10098_));
  XOR2_X1    g10034(.A1(new_n10098_), .A2(new_n10070_), .Z(new_n10099_));
  OAI22_X1   g10035(.A1(new_n2311_), .A2(new_n9489_), .B1(new_n4365_), .B2(new_n9485_), .ZN(new_n10100_));
  NAND2_X1   g10036(.A1(new_n2255_), .A2(new_n9503_), .ZN(new_n10101_));
  AOI21_X1   g10037(.A1(new_n10100_), .A2(new_n10101_), .B(new_n9482_), .ZN(new_n10102_));
  NAND2_X1   g10038(.A1(new_n4419_), .A2(new_n10102_), .ZN(new_n10103_));
  XOR2_X1    g10039(.A1(new_n10103_), .A2(new_n4387_), .Z(new_n10104_));
  NOR2_X1    g10040(.A1(new_n10099_), .A2(new_n10104_), .ZN(new_n10105_));
  NAND2_X1   g10041(.A1(new_n10099_), .A2(new_n10104_), .ZN(new_n10106_));
  OAI21_X1   g10042(.A1(new_n10067_), .A2(new_n10105_), .B(new_n10106_), .ZN(new_n10107_));
  OAI22_X1   g10043(.A1(new_n2251_), .A2(new_n9485_), .B1(new_n2351_), .B2(new_n9489_), .ZN(new_n10108_));
  NAND2_X1   g10044(.A1(new_n2310_), .A2(new_n9503_), .ZN(new_n10109_));
  AOI21_X1   g10045(.A1(new_n10109_), .A2(new_n10108_), .B(new_n9482_), .ZN(new_n10110_));
  NAND2_X1   g10046(.A1(new_n3914_), .A2(new_n10110_), .ZN(new_n10111_));
  XOR2_X1    g10047(.A1(new_n10111_), .A2(\a[2] ), .Z(new_n10112_));
  INV_X1     g10048(.I(new_n10112_), .ZN(new_n10113_));
  NAND2_X1   g10049(.A1(new_n10107_), .A2(new_n10113_), .ZN(new_n10114_));
  NAND3_X1   g10050(.A1(new_n10014_), .A2(new_n10005_), .A3(new_n10002_), .ZN(new_n10115_));
  NAND2_X1   g10051(.A1(new_n10003_), .A2(new_n9579_), .ZN(new_n10116_));
  OAI21_X1   g10052(.A1(new_n10064_), .A2(new_n10063_), .B(new_n10062_), .ZN(new_n10117_));
  NAND3_X1   g10053(.A1(new_n10056_), .A2(new_n10060_), .A3(new_n10044_), .ZN(new_n10118_));
  NAND2_X1   g10054(.A1(new_n10117_), .A2(new_n10118_), .ZN(new_n10119_));
  AOI22_X1   g10055(.A1(new_n10116_), .A2(new_n10115_), .B1(new_n10005_), .B2(new_n10119_), .ZN(new_n10120_));
  INV_X1     g10056(.I(new_n10105_), .ZN(new_n10121_));
  NAND2_X1   g10057(.A1(new_n10120_), .A2(new_n10121_), .ZN(new_n10122_));
  XOR2_X1    g10058(.A1(new_n10070_), .A2(new_n65_), .Z(new_n10123_));
  OR2_X2     g10059(.A1(new_n10097_), .A2(new_n10123_), .Z(new_n10124_));
  NOR3_X1    g10060(.A1(new_n10090_), .A2(new_n10088_), .A3(new_n10096_), .ZN(new_n10125_));
  INV_X1     g10061(.I(new_n10125_), .ZN(new_n10126_));
  NAND2_X1   g10062(.A1(new_n10080_), .A2(new_n10081_), .ZN(new_n10127_));
  INV_X1     g10063(.I(new_n8971_), .ZN(new_n10128_));
  OAI22_X1   g10064(.A1(new_n1729_), .A2(new_n6091_), .B1(new_n4745_), .B2(new_n6089_), .ZN(new_n10129_));
  NAND2_X1   g10065(.A1(new_n1862_), .A2(new_n6095_), .ZN(new_n10130_));
  AOI21_X1   g10066(.A1(new_n10129_), .A2(new_n10130_), .B(new_n6082_), .ZN(new_n10131_));
  NAND2_X1   g10067(.A1(new_n4842_), .A2(new_n10131_), .ZN(new_n10132_));
  XOR2_X1    g10068(.A1(new_n10132_), .A2(\a[14] ), .Z(new_n10133_));
  XOR2_X1    g10069(.A1(new_n10133_), .A2(new_n10128_), .Z(new_n10134_));
  NOR2_X1    g10070(.A1(new_n10133_), .A2(new_n8971_), .ZN(new_n10135_));
  XOR2_X1    g10071(.A1(new_n10132_), .A2(new_n3521_), .Z(new_n10136_));
  NOR2_X1    g10072(.A1(new_n10136_), .A2(new_n10128_), .ZN(new_n10137_));
  OAI21_X1   g10073(.A1(new_n10135_), .A2(new_n10137_), .B(new_n10127_), .ZN(new_n10138_));
  OAI21_X1   g10074(.A1(new_n10134_), .A2(new_n10127_), .B(new_n10138_), .ZN(new_n10139_));
  OAI22_X1   g10075(.A1(new_n1678_), .A2(new_n4710_), .B1(new_n1764_), .B2(new_n4716_), .ZN(new_n10140_));
  NAND2_X1   g10076(.A1(new_n1613_), .A2(new_n4720_), .ZN(new_n10141_));
  AOI21_X1   g10077(.A1(new_n10140_), .A2(new_n10141_), .B(new_n4707_), .ZN(new_n10142_));
  NAND2_X1   g10078(.A1(new_n4917_), .A2(new_n10142_), .ZN(new_n10143_));
  XOR2_X1    g10079(.A1(new_n10143_), .A2(new_n4034_), .Z(new_n10144_));
  XOR2_X1    g10080(.A1(new_n10139_), .A2(new_n10144_), .Z(new_n10145_));
  OAI21_X1   g10081(.A1(new_n10071_), .A2(new_n10086_), .B(new_n10084_), .ZN(new_n10146_));
  NOR2_X1    g10082(.A1(new_n10146_), .A2(new_n10145_), .ZN(new_n10147_));
  INV_X1     g10083(.I(new_n10147_), .ZN(new_n10148_));
  NAND2_X1   g10084(.A1(new_n10146_), .A2(new_n10145_), .ZN(new_n10149_));
  OAI22_X1   g10085(.A1(new_n2103_), .A2(new_n6788_), .B1(new_n2158_), .B2(new_n6785_), .ZN(new_n10150_));
  NAND2_X1   g10086(.A1(new_n2107_), .A2(new_n7530_), .ZN(new_n10151_));
  AOI21_X1   g10087(.A1(new_n10150_), .A2(new_n10151_), .B(new_n6776_), .ZN(new_n10152_));
  NAND2_X1   g10088(.A1(new_n4959_), .A2(new_n10152_), .ZN(new_n10153_));
  XOR2_X1    g10089(.A1(new_n10153_), .A2(\a[8] ), .Z(new_n10154_));
  INV_X1     g10090(.I(new_n10154_), .ZN(new_n10155_));
  NAND3_X1   g10091(.A1(new_n10155_), .A2(new_n10148_), .A3(new_n10149_), .ZN(new_n10156_));
  INV_X1     g10092(.I(new_n10149_), .ZN(new_n10157_));
  OAI21_X1   g10093(.A1(new_n10157_), .A2(new_n10147_), .B(new_n10154_), .ZN(new_n10158_));
  NAND3_X1   g10094(.A1(new_n10156_), .A2(new_n10158_), .A3(new_n10126_), .ZN(new_n10159_));
  INV_X1     g10095(.I(new_n10159_), .ZN(new_n10160_));
  AOI21_X1   g10096(.A1(new_n10156_), .A2(new_n10158_), .B(new_n10126_), .ZN(new_n10161_));
  NOR2_X1    g10097(.A1(new_n10160_), .A2(new_n10161_), .ZN(new_n10162_));
  OAI22_X1   g10098(.A1(new_n4365_), .A2(new_n6839_), .B1(new_n2198_), .B2(new_n6913_), .ZN(new_n10163_));
  NAND2_X1   g10099(.A1(new_n1504_), .A2(new_n8799_), .ZN(new_n10164_));
  AOI21_X1   g10100(.A1(new_n10163_), .A2(new_n10164_), .B(new_n6836_), .ZN(new_n10165_));
  NAND2_X1   g10101(.A1(new_n4363_), .A2(new_n10165_), .ZN(new_n10166_));
  XOR2_X1    g10102(.A1(new_n10166_), .A2(\a[5] ), .Z(new_n10167_));
  XNOR2_X1   g10103(.A1(new_n10162_), .A2(new_n10167_), .ZN(new_n10168_));
  OR2_X2     g10104(.A1(new_n10168_), .A2(new_n10124_), .Z(new_n10169_));
  NAND2_X1   g10105(.A1(new_n10168_), .A2(new_n10124_), .ZN(new_n10170_));
  AOI21_X1   g10106(.A1(new_n10169_), .A2(new_n10170_), .B(new_n10113_), .ZN(new_n10171_));
  NAND3_X1   g10107(.A1(new_n10122_), .A2(new_n10106_), .A3(new_n10171_), .ZN(new_n10172_));
  OAI22_X1   g10108(.A1(new_n1453_), .A2(new_n9489_), .B1(new_n2351_), .B2(new_n9483_), .ZN(new_n10173_));
  NAND2_X1   g10109(.A1(new_n2310_), .A2(new_n6925_), .ZN(new_n10174_));
  AOI21_X1   g10110(.A1(new_n10174_), .A2(new_n10173_), .B(new_n9482_), .ZN(new_n10175_));
  NAND2_X1   g10111(.A1(new_n4231_), .A2(new_n10175_), .ZN(new_n10176_));
  XOR2_X1    g10112(.A1(new_n10176_), .A2(\a[2] ), .Z(new_n10177_));
  AOI21_X1   g10113(.A1(new_n10114_), .A2(new_n10172_), .B(new_n10177_), .ZN(new_n10178_));
  AOI21_X1   g10114(.A1(new_n10122_), .A2(new_n10106_), .B(new_n10112_), .ZN(new_n10179_));
  INV_X1     g10115(.I(new_n10171_), .ZN(new_n10180_));
  NOR2_X1    g10116(.A1(new_n10107_), .A2(new_n10180_), .ZN(new_n10181_));
  INV_X1     g10117(.I(new_n10177_), .ZN(new_n10182_));
  AOI21_X1   g10118(.A1(new_n10124_), .A2(new_n10167_), .B(new_n10162_), .ZN(new_n10183_));
  NOR2_X1    g10119(.A1(new_n10124_), .A2(new_n10167_), .ZN(new_n10184_));
  NOR2_X1    g10120(.A1(new_n10183_), .A2(new_n10184_), .ZN(new_n10185_));
  INV_X1     g10121(.I(new_n10185_), .ZN(new_n10186_));
  INV_X1     g10122(.I(new_n10137_), .ZN(new_n10187_));
  AOI21_X1   g10123(.A1(new_n10187_), .A2(new_n10127_), .B(new_n10135_), .ZN(new_n10188_));
  XNOR2_X1   g10124(.A1(new_n8970_), .A2(new_n8972_), .ZN(new_n10189_));
  OAI22_X1   g10125(.A1(new_n1764_), .A2(new_n6091_), .B1(new_n1729_), .B2(new_n6094_), .ZN(new_n10190_));
  NAND2_X1   g10126(.A1(new_n1862_), .A2(new_n6180_), .ZN(new_n10191_));
  AOI21_X1   g10127(.A1(new_n10190_), .A2(new_n10191_), .B(new_n6082_), .ZN(new_n10192_));
  NAND2_X1   g10128(.A1(new_n4810_), .A2(new_n10192_), .ZN(new_n10193_));
  XOR2_X1    g10129(.A1(new_n10193_), .A2(new_n3521_), .Z(new_n10194_));
  XNOR2_X1   g10130(.A1(new_n10194_), .A2(new_n10189_), .ZN(new_n10195_));
  NOR2_X1    g10131(.A1(new_n10195_), .A2(new_n10188_), .ZN(new_n10196_));
  INV_X1     g10132(.I(new_n10188_), .ZN(new_n10197_));
  NOR2_X1    g10133(.A1(new_n10194_), .A2(new_n10189_), .ZN(new_n10198_));
  INV_X1     g10134(.I(new_n10198_), .ZN(new_n10199_));
  NAND2_X1   g10135(.A1(new_n10194_), .A2(new_n10189_), .ZN(new_n10200_));
  AOI21_X1   g10136(.A1(new_n10199_), .A2(new_n10200_), .B(new_n10197_), .ZN(new_n10201_));
  NOR2_X1    g10137(.A1(new_n10201_), .A2(new_n10196_), .ZN(new_n10202_));
  INV_X1     g10138(.I(new_n10202_), .ZN(new_n10203_));
  NOR2_X1    g10139(.A1(new_n10139_), .A2(new_n10144_), .ZN(new_n10204_));
  OAI22_X1   g10140(.A1(new_n1678_), .A2(new_n4719_), .B1(new_n2071_), .B2(new_n4710_), .ZN(new_n10205_));
  NAND2_X1   g10141(.A1(new_n1613_), .A2(new_n6480_), .ZN(new_n10206_));
  AOI21_X1   g10142(.A1(new_n10205_), .A2(new_n10206_), .B(new_n4707_), .ZN(new_n10207_));
  NAND2_X1   g10143(.A1(new_n5070_), .A2(new_n10207_), .ZN(new_n10208_));
  XOR2_X1    g10144(.A1(new_n10208_), .A2(\a[11] ), .Z(new_n10209_));
  OAI21_X1   g10145(.A1(new_n10147_), .A2(new_n10204_), .B(new_n10209_), .ZN(new_n10210_));
  NOR3_X1    g10146(.A1(new_n10147_), .A2(new_n10204_), .A3(new_n10209_), .ZN(new_n10211_));
  INV_X1     g10147(.I(new_n10211_), .ZN(new_n10212_));
  AOI21_X1   g10148(.A1(new_n10212_), .A2(new_n10210_), .B(new_n10203_), .ZN(new_n10213_));
  INV_X1     g10149(.I(new_n10210_), .ZN(new_n10214_));
  NOR3_X1    g10150(.A1(new_n10214_), .A2(new_n10202_), .A3(new_n10211_), .ZN(new_n10215_));
  NOR2_X1    g10151(.A1(new_n10213_), .A2(new_n10215_), .ZN(new_n10216_));
  INV_X1     g10152(.I(new_n10216_), .ZN(new_n10217_));
  OAI22_X1   g10153(.A1(new_n2103_), .A2(new_n6783_), .B1(new_n2198_), .B2(new_n6785_), .ZN(new_n10218_));
  NAND2_X1   g10154(.A1(new_n2161_), .A2(new_n6789_), .ZN(new_n10219_));
  AOI21_X1   g10155(.A1(new_n10218_), .A2(new_n10219_), .B(new_n6776_), .ZN(new_n10220_));
  NAND2_X1   g10156(.A1(new_n5351_), .A2(new_n10220_), .ZN(new_n10221_));
  XOR2_X1    g10157(.A1(new_n10221_), .A2(\a[8] ), .Z(new_n10222_));
  INV_X1     g10158(.I(new_n10222_), .ZN(new_n10223_));
  AOI21_X1   g10159(.A1(new_n10159_), .A2(new_n10158_), .B(new_n10223_), .ZN(new_n10224_));
  INV_X1     g10160(.I(new_n10224_), .ZN(new_n10225_));
  NAND3_X1   g10161(.A1(new_n10159_), .A2(new_n10158_), .A3(new_n10223_), .ZN(new_n10226_));
  AOI21_X1   g10162(.A1(new_n10225_), .A2(new_n10226_), .B(new_n10217_), .ZN(new_n10227_));
  INV_X1     g10163(.I(new_n10226_), .ZN(new_n10228_));
  NOR3_X1    g10164(.A1(new_n10228_), .A2(new_n10216_), .A3(new_n10224_), .ZN(new_n10229_));
  NOR2_X1    g10165(.A1(new_n10227_), .A2(new_n10229_), .ZN(new_n10230_));
  OAI22_X1   g10166(.A1(new_n2251_), .A2(new_n6839_), .B1(new_n4365_), .B2(new_n6843_), .ZN(new_n10231_));
  NAND2_X1   g10167(.A1(new_n1504_), .A2(new_n6846_), .ZN(new_n10232_));
  AOI21_X1   g10168(.A1(new_n10231_), .A2(new_n10232_), .B(new_n6836_), .ZN(new_n10233_));
  NAND2_X1   g10169(.A1(new_n4650_), .A2(new_n10233_), .ZN(new_n10234_));
  XOR2_X1    g10170(.A1(new_n10234_), .A2(\a[5] ), .Z(new_n10235_));
  INV_X1     g10171(.I(new_n10235_), .ZN(new_n10236_));
  NAND2_X1   g10172(.A1(new_n10230_), .A2(new_n10236_), .ZN(new_n10237_));
  NOR2_X1    g10173(.A1(new_n10230_), .A2(new_n10236_), .ZN(new_n10238_));
  INV_X1     g10174(.I(new_n10238_), .ZN(new_n10239_));
  NAND3_X1   g10175(.A1(new_n10239_), .A2(new_n10186_), .A3(new_n10237_), .ZN(new_n10240_));
  INV_X1     g10176(.I(new_n10237_), .ZN(new_n10241_));
  OAI21_X1   g10177(.A1(new_n10241_), .A2(new_n10238_), .B(new_n10185_), .ZN(new_n10242_));
  AOI21_X1   g10178(.A1(new_n10242_), .A2(new_n10240_), .B(new_n10182_), .ZN(new_n10243_));
  INV_X1     g10179(.I(new_n10243_), .ZN(new_n10244_));
  NOR3_X1    g10180(.A1(new_n10181_), .A2(new_n10179_), .A3(new_n10244_), .ZN(new_n10245_));
  NAND2_X1   g10181(.A1(new_n4620_), .A2(new_n6775_), .ZN(new_n10246_));
  AOI22_X1   g10182(.A1(new_n2161_), .A2(new_n7530_), .B1(new_n2202_), .B2(new_n6789_), .ZN(new_n10247_));
  AOI21_X1   g10183(.A1(new_n1504_), .A2(new_n6784_), .B(new_n10247_), .ZN(new_n10248_));
  NAND2_X1   g10184(.A1(new_n10246_), .A2(new_n10248_), .ZN(new_n10249_));
  OAI21_X1   g10185(.A1(new_n10188_), .A2(new_n10198_), .B(new_n10200_), .ZN(new_n10250_));
  OAI22_X1   g10186(.A1(new_n1764_), .A2(new_n6094_), .B1(new_n1729_), .B2(new_n6089_), .ZN(new_n10251_));
  NAND2_X1   g10187(.A1(new_n1613_), .A2(new_n6090_), .ZN(new_n10252_));
  AOI21_X1   g10188(.A1(new_n10252_), .A2(new_n10251_), .B(new_n6082_), .ZN(new_n10253_));
  NAND2_X1   g10189(.A1(new_n4778_), .A2(new_n10253_), .ZN(new_n10254_));
  XOR2_X1    g10190(.A1(new_n10254_), .A2(\a[14] ), .Z(new_n10255_));
  XOR2_X1    g10191(.A1(new_n8973_), .A2(new_n8966_), .Z(new_n10256_));
  NAND2_X1   g10192(.A1(new_n10255_), .A2(new_n10256_), .ZN(new_n10257_));
  INV_X1     g10193(.I(new_n10257_), .ZN(new_n10258_));
  NOR2_X1    g10194(.A1(new_n10255_), .A2(new_n10256_), .ZN(new_n10259_));
  NOR2_X1    g10195(.A1(new_n10258_), .A2(new_n10259_), .ZN(new_n10260_));
  XOR2_X1    g10196(.A1(new_n10260_), .A2(new_n10250_), .Z(new_n10261_));
  OAI22_X1   g10197(.A1(new_n2103_), .A2(new_n4710_), .B1(new_n1678_), .B2(new_n4716_), .ZN(new_n10262_));
  NAND2_X1   g10198(.A1(new_n2107_), .A2(new_n4720_), .ZN(new_n10263_));
  AOI21_X1   g10199(.A1(new_n10262_), .A2(new_n10263_), .B(new_n4707_), .ZN(new_n10264_));
  NAND2_X1   g10200(.A1(new_n4545_), .A2(new_n10264_), .ZN(new_n10265_));
  XOR2_X1    g10201(.A1(new_n10265_), .A2(\a[11] ), .Z(new_n10266_));
  XOR2_X1    g10202(.A1(new_n10261_), .A2(new_n10266_), .Z(new_n10267_));
  XOR2_X1    g10203(.A1(new_n10267_), .A2(new_n4009_), .Z(new_n10268_));
  XOR2_X1    g10204(.A1(new_n10268_), .A2(new_n10249_), .Z(new_n10269_));
  INV_X1     g10205(.I(new_n10269_), .ZN(new_n10270_));
  NOR2_X1    g10206(.A1(new_n10185_), .A2(new_n10235_), .ZN(new_n10271_));
  INV_X1     g10207(.I(new_n10230_), .ZN(new_n10272_));
  AOI21_X1   g10208(.A1(new_n10185_), .A2(new_n10235_), .B(new_n10272_), .ZN(new_n10273_));
  OAI22_X1   g10209(.A1(new_n2311_), .A2(new_n6839_), .B1(new_n4365_), .B2(new_n6913_), .ZN(new_n10274_));
  NAND2_X1   g10210(.A1(new_n2255_), .A2(new_n8799_), .ZN(new_n10275_));
  AOI21_X1   g10211(.A1(new_n10274_), .A2(new_n10275_), .B(new_n6836_), .ZN(new_n10276_));
  NAND2_X1   g10212(.A1(new_n4419_), .A2(new_n10276_), .ZN(new_n10277_));
  XOR2_X1    g10213(.A1(new_n10277_), .A2(\a[5] ), .Z(new_n10278_));
  INV_X1     g10214(.I(new_n10278_), .ZN(new_n10279_));
  NOR3_X1    g10215(.A1(new_n10273_), .A2(new_n10271_), .A3(new_n10279_), .ZN(new_n10280_));
  INV_X1     g10216(.I(new_n10271_), .ZN(new_n10281_));
  OAI21_X1   g10217(.A1(new_n10186_), .A2(new_n10236_), .B(new_n10230_), .ZN(new_n10282_));
  AOI21_X1   g10218(.A1(new_n10282_), .A2(new_n10281_), .B(new_n10278_), .ZN(new_n10283_));
  OAI21_X1   g10219(.A1(new_n10280_), .A2(new_n10283_), .B(new_n10270_), .ZN(new_n10284_));
  INV_X1     g10220(.I(new_n10284_), .ZN(new_n10285_));
  AOI21_X1   g10221(.A1(new_n10282_), .A2(new_n10281_), .B(new_n10279_), .ZN(new_n10286_));
  INV_X1     g10222(.I(new_n10286_), .ZN(new_n10287_));
  NAND3_X1   g10223(.A1(new_n10282_), .A2(new_n10281_), .A3(new_n10279_), .ZN(new_n10288_));
  AOI21_X1   g10224(.A1(new_n10287_), .A2(new_n10288_), .B(new_n10270_), .ZN(new_n10289_));
  OAI22_X1   g10225(.A1(new_n1409_), .A2(new_n9489_), .B1(new_n2351_), .B2(new_n9485_), .ZN(new_n10290_));
  NAND2_X1   g10226(.A1(new_n2359_), .A2(new_n9503_), .ZN(new_n10291_));
  AOI21_X1   g10227(.A1(new_n10290_), .A2(new_n10291_), .B(new_n9482_), .ZN(new_n10292_));
  NAND2_X1   g10228(.A1(new_n3904_), .A2(new_n10292_), .ZN(new_n10293_));
  XOR2_X1    g10229(.A1(new_n10293_), .A2(\a[2] ), .Z(new_n10294_));
  OAI21_X1   g10230(.A1(new_n10285_), .A2(new_n10289_), .B(new_n10294_), .ZN(new_n10295_));
  OAI21_X1   g10231(.A1(new_n10245_), .A2(new_n10178_), .B(new_n10295_), .ZN(new_n10296_));
  NOR3_X1    g10232(.A1(new_n10285_), .A2(new_n10289_), .A3(new_n10294_), .ZN(new_n10297_));
  INV_X1     g10233(.I(new_n10297_), .ZN(new_n10298_));
  NAND3_X1   g10234(.A1(new_n10296_), .A2(new_n9574_), .A3(new_n10298_), .ZN(new_n10299_));
  OAI21_X1   g10235(.A1(new_n10181_), .A2(new_n10179_), .B(new_n10182_), .ZN(new_n10300_));
  NAND3_X1   g10236(.A1(new_n10114_), .A2(new_n10172_), .A3(new_n10243_), .ZN(new_n10301_));
  INV_X1     g10237(.I(new_n10288_), .ZN(new_n10302_));
  OAI21_X1   g10238(.A1(new_n10302_), .A2(new_n10286_), .B(new_n10269_), .ZN(new_n10303_));
  INV_X1     g10239(.I(new_n10294_), .ZN(new_n10304_));
  AOI21_X1   g10240(.A1(new_n10303_), .A2(new_n10284_), .B(new_n10304_), .ZN(new_n10305_));
  AOI21_X1   g10241(.A1(new_n10300_), .A2(new_n10301_), .B(new_n10305_), .ZN(new_n10306_));
  OAI21_X1   g10242(.A1(new_n10306_), .A2(new_n10297_), .B(new_n9573_), .ZN(new_n10307_));
  XOR2_X1    g10243(.A1(new_n10249_), .A2(\a[8] ), .Z(new_n10308_));
  NOR2_X1    g10244(.A1(new_n10308_), .A2(new_n10267_), .ZN(new_n10309_));
  INV_X1     g10245(.I(new_n10266_), .ZN(new_n10310_));
  NAND2_X1   g10246(.A1(new_n10310_), .A2(new_n10261_), .ZN(new_n10311_));
  XOR2_X1    g10247(.A1(new_n8961_), .A2(new_n8956_), .Z(new_n10312_));
  NAND2_X1   g10248(.A1(new_n10312_), .A2(new_n8974_), .ZN(new_n10313_));
  INV_X1     g10249(.I(new_n8962_), .ZN(new_n10314_));
  OAI22_X1   g10250(.A1(new_n10314_), .A2(new_n8975_), .B1(new_n8966_), .B2(new_n8973_), .ZN(new_n10315_));
  NAND2_X1   g10251(.A1(new_n10313_), .A2(new_n10315_), .ZN(new_n10316_));
  OAI22_X1   g10252(.A1(new_n1678_), .A2(new_n6091_), .B1(new_n1764_), .B2(new_n6089_), .ZN(new_n10317_));
  NAND2_X1   g10253(.A1(new_n1613_), .A2(new_n6095_), .ZN(new_n10318_));
  AOI21_X1   g10254(.A1(new_n10317_), .A2(new_n10318_), .B(new_n6082_), .ZN(new_n10319_));
  NAND2_X1   g10255(.A1(new_n4917_), .A2(new_n10319_), .ZN(new_n10320_));
  XOR2_X1    g10256(.A1(new_n10320_), .A2(new_n3521_), .Z(new_n10321_));
  XOR2_X1    g10257(.A1(new_n10316_), .A2(new_n10321_), .Z(new_n10322_));
  OAI21_X1   g10258(.A1(new_n10250_), .A2(new_n10259_), .B(new_n10257_), .ZN(new_n10323_));
  XOR2_X1    g10259(.A1(new_n10322_), .A2(new_n10323_), .Z(new_n10324_));
  OAI22_X1   g10260(.A1(new_n2103_), .A2(new_n4719_), .B1(new_n2158_), .B2(new_n4710_), .ZN(new_n10325_));
  NAND2_X1   g10261(.A1(new_n2107_), .A2(new_n6480_), .ZN(new_n10326_));
  AOI21_X1   g10262(.A1(new_n10325_), .A2(new_n10326_), .B(new_n4707_), .ZN(new_n10327_));
  NAND2_X1   g10263(.A1(new_n4959_), .A2(new_n10327_), .ZN(new_n10328_));
  XOR2_X1    g10264(.A1(new_n10328_), .A2(new_n4034_), .Z(new_n10329_));
  XOR2_X1    g10265(.A1(new_n10324_), .A2(new_n10329_), .Z(new_n10330_));
  XOR2_X1    g10266(.A1(new_n10330_), .A2(new_n10311_), .Z(new_n10331_));
  OAI22_X1   g10267(.A1(new_n4365_), .A2(new_n6785_), .B1(new_n2198_), .B2(new_n6783_), .ZN(new_n10332_));
  NAND2_X1   g10268(.A1(new_n1504_), .A2(new_n6789_), .ZN(new_n10333_));
  AOI21_X1   g10269(.A1(new_n10332_), .A2(new_n10333_), .B(new_n6776_), .ZN(new_n10334_));
  NAND2_X1   g10270(.A1(new_n4363_), .A2(new_n10334_), .ZN(new_n10335_));
  XOR2_X1    g10271(.A1(new_n10335_), .A2(\a[8] ), .Z(new_n10336_));
  NAND2_X1   g10272(.A1(new_n10331_), .A2(new_n10336_), .ZN(new_n10337_));
  XNOR2_X1   g10273(.A1(new_n10330_), .A2(new_n10311_), .ZN(new_n10338_));
  INV_X1     g10274(.I(new_n10336_), .ZN(new_n10339_));
  NAND2_X1   g10275(.A1(new_n10338_), .A2(new_n10339_), .ZN(new_n10340_));
  NAND2_X1   g10276(.A1(new_n10340_), .A2(new_n10337_), .ZN(new_n10341_));
  OAI22_X1   g10277(.A1(new_n2251_), .A2(new_n6913_), .B1(new_n2351_), .B2(new_n6839_), .ZN(new_n10342_));
  NAND2_X1   g10278(.A1(new_n2310_), .A2(new_n8799_), .ZN(new_n10343_));
  AOI21_X1   g10279(.A1(new_n10343_), .A2(new_n10342_), .B(new_n6836_), .ZN(new_n10344_));
  NAND2_X1   g10280(.A1(new_n3914_), .A2(new_n10344_), .ZN(new_n10345_));
  XOR2_X1    g10281(.A1(new_n10345_), .A2(\a[5] ), .Z(new_n10346_));
  INV_X1     g10282(.I(new_n10346_), .ZN(new_n10347_));
  NOR2_X1    g10283(.A1(new_n10341_), .A2(new_n10347_), .ZN(new_n10348_));
  NAND2_X1   g10284(.A1(new_n10341_), .A2(new_n10347_), .ZN(new_n10349_));
  INV_X1     g10285(.I(new_n10349_), .ZN(new_n10350_));
  OAI21_X1   g10286(.A1(new_n10350_), .A2(new_n10348_), .B(new_n10309_), .ZN(new_n10351_));
  INV_X1     g10287(.I(new_n10309_), .ZN(new_n10352_));
  NOR2_X1    g10288(.A1(new_n10338_), .A2(new_n10339_), .ZN(new_n10353_));
  NOR2_X1    g10289(.A1(new_n10331_), .A2(new_n10336_), .ZN(new_n10354_));
  NOR2_X1    g10290(.A1(new_n10353_), .A2(new_n10354_), .ZN(new_n10355_));
  NOR2_X1    g10291(.A1(new_n10355_), .A2(new_n10347_), .ZN(new_n10356_));
  NOR2_X1    g10292(.A1(new_n10341_), .A2(new_n10346_), .ZN(new_n10357_));
  OAI21_X1   g10293(.A1(new_n10356_), .A2(new_n10357_), .B(new_n10352_), .ZN(new_n10358_));
  NAND2_X1   g10294(.A1(new_n10351_), .A2(new_n10358_), .ZN(new_n10359_));
  OAI21_X1   g10295(.A1(new_n10273_), .A2(new_n10271_), .B(new_n10269_), .ZN(new_n10360_));
  NOR2_X1    g10296(.A1(new_n10359_), .A2(new_n10360_), .ZN(new_n10361_));
  NAND2_X1   g10297(.A1(new_n10355_), .A2(new_n10346_), .ZN(new_n10362_));
  AOI21_X1   g10298(.A1(new_n10349_), .A2(new_n10362_), .B(new_n10352_), .ZN(new_n10363_));
  NAND2_X1   g10299(.A1(new_n10341_), .A2(new_n10346_), .ZN(new_n10364_));
  NAND2_X1   g10300(.A1(new_n10355_), .A2(new_n10347_), .ZN(new_n10365_));
  AOI21_X1   g10301(.A1(new_n10365_), .A2(new_n10364_), .B(new_n10309_), .ZN(new_n10366_));
  NOR2_X1    g10302(.A1(new_n10363_), .A2(new_n10366_), .ZN(new_n10367_));
  INV_X1     g10303(.I(new_n10360_), .ZN(new_n10368_));
  NOR2_X1    g10304(.A1(new_n10367_), .A2(new_n10368_), .ZN(new_n10369_));
  NAND3_X1   g10305(.A1(new_n10282_), .A2(new_n10270_), .A3(new_n10281_), .ZN(new_n10370_));
  AND3_X2    g10306(.A1(new_n10360_), .A2(new_n10278_), .A3(new_n10370_), .Z(new_n10371_));
  NOR3_X1    g10307(.A1(new_n10361_), .A2(new_n10369_), .A3(new_n10371_), .ZN(new_n10372_));
  AND4_X2    g10308(.A1(new_n10278_), .A2(new_n10359_), .A3(new_n10360_), .A4(new_n10370_), .Z(new_n10373_));
  OR2_X2     g10309(.A1(new_n10372_), .A2(new_n10373_), .Z(new_n10374_));
  AOI22_X1   g10310(.A1(new_n10299_), .A2(new_n10307_), .B1(new_n10374_), .B2(new_n9574_), .ZN(new_n10375_));
  XOR2_X1    g10311(.A1(new_n8982_), .A2(new_n8977_), .Z(new_n10376_));
  AOI21_X1   g10312(.A1(new_n8985_), .A2(new_n8983_), .B(new_n8976_), .ZN(new_n10377_));
  AOI21_X1   g10313(.A1(new_n8976_), .A2(new_n10376_), .B(new_n10377_), .ZN(new_n10378_));
  NOR2_X1    g10314(.A1(new_n10322_), .A2(new_n10323_), .ZN(new_n10379_));
  NOR2_X1    g10315(.A1(new_n10316_), .A2(new_n10321_), .ZN(new_n10380_));
  NOR2_X1    g10316(.A1(new_n10379_), .A2(new_n10380_), .ZN(new_n10381_));
  OAI22_X1   g10317(.A1(new_n1678_), .A2(new_n6094_), .B1(new_n2071_), .B2(new_n6091_), .ZN(new_n10382_));
  NAND2_X1   g10318(.A1(new_n1613_), .A2(new_n6180_), .ZN(new_n10383_));
  AOI21_X1   g10319(.A1(new_n10382_), .A2(new_n10383_), .B(new_n6082_), .ZN(new_n10384_));
  NAND2_X1   g10320(.A1(new_n5070_), .A2(new_n10384_), .ZN(new_n10385_));
  XOR2_X1    g10321(.A1(new_n10385_), .A2(\a[14] ), .Z(new_n10386_));
  XOR2_X1    g10322(.A1(new_n10381_), .A2(new_n10386_), .Z(new_n10387_));
  XNOR2_X1   g10323(.A1(new_n10387_), .A2(new_n10378_), .ZN(new_n10388_));
  NOR2_X1    g10324(.A1(new_n10324_), .A2(new_n10329_), .ZN(new_n10389_));
  AOI21_X1   g10325(.A1(new_n10330_), .A2(new_n10311_), .B(new_n10389_), .ZN(new_n10390_));
  OAI22_X1   g10326(.A1(new_n2103_), .A2(new_n4716_), .B1(new_n2198_), .B2(new_n4710_), .ZN(new_n10391_));
  NAND2_X1   g10327(.A1(new_n2161_), .A2(new_n4720_), .ZN(new_n10392_));
  AOI21_X1   g10328(.A1(new_n10391_), .A2(new_n10392_), .B(new_n4707_), .ZN(new_n10393_));
  NAND2_X1   g10329(.A1(new_n5351_), .A2(new_n10393_), .ZN(new_n10394_));
  XOR2_X1    g10330(.A1(new_n10394_), .A2(new_n4034_), .Z(new_n10395_));
  XOR2_X1    g10331(.A1(new_n10390_), .A2(new_n10395_), .Z(new_n10396_));
  XNOR2_X1   g10332(.A1(new_n10396_), .A2(new_n10388_), .ZN(new_n10397_));
  OAI21_X1   g10333(.A1(new_n10309_), .A2(new_n10354_), .B(new_n10337_), .ZN(new_n10398_));
  OAI22_X1   g10334(.A1(new_n2251_), .A2(new_n6785_), .B1(new_n4365_), .B2(new_n6788_), .ZN(new_n10399_));
  NAND2_X1   g10335(.A1(new_n1504_), .A2(new_n7530_), .ZN(new_n10400_));
  AOI21_X1   g10336(.A1(new_n10399_), .A2(new_n10400_), .B(new_n6776_), .ZN(new_n10401_));
  NAND2_X1   g10337(.A1(new_n4650_), .A2(new_n10401_), .ZN(new_n10402_));
  XOR2_X1    g10338(.A1(new_n10402_), .A2(\a[8] ), .Z(new_n10403_));
  NAND2_X1   g10339(.A1(new_n10398_), .A2(new_n10403_), .ZN(new_n10404_));
  NOR2_X1    g10340(.A1(new_n10398_), .A2(new_n10403_), .ZN(new_n10405_));
  INV_X1     g10341(.I(new_n10405_), .ZN(new_n10406_));
  AOI21_X1   g10342(.A1(new_n10406_), .A2(new_n10404_), .B(new_n10397_), .ZN(new_n10407_));
  XOR2_X1    g10343(.A1(new_n10396_), .A2(new_n10388_), .Z(new_n10408_));
  INV_X1     g10344(.I(new_n10404_), .ZN(new_n10409_));
  NOR3_X1    g10345(.A1(new_n10409_), .A2(new_n10408_), .A3(new_n10405_), .ZN(new_n10410_));
  NOR2_X1    g10346(.A1(new_n10407_), .A2(new_n10410_), .ZN(new_n10411_));
  NAND2_X1   g10347(.A1(new_n10355_), .A2(new_n10309_), .ZN(new_n10412_));
  NAND2_X1   g10348(.A1(new_n10341_), .A2(new_n10352_), .ZN(new_n10413_));
  NAND2_X1   g10349(.A1(new_n10412_), .A2(new_n10413_), .ZN(new_n10414_));
  AOI22_X1   g10350(.A1(new_n10360_), .A2(new_n10279_), .B1(new_n10414_), .B2(new_n10346_), .ZN(new_n10415_));
  OAI22_X1   g10351(.A1(new_n1453_), .A2(new_n6839_), .B1(new_n2351_), .B2(new_n6843_), .ZN(new_n10416_));
  NAND2_X1   g10352(.A1(new_n2310_), .A2(new_n6846_), .ZN(new_n10417_));
  AOI21_X1   g10353(.A1(new_n10417_), .A2(new_n10416_), .B(new_n6836_), .ZN(new_n10418_));
  NAND2_X1   g10354(.A1(new_n4231_), .A2(new_n10418_), .ZN(new_n10419_));
  XOR2_X1    g10355(.A1(new_n10419_), .A2(\a[5] ), .Z(new_n10420_));
  INV_X1     g10356(.I(new_n10420_), .ZN(new_n10421_));
  AOI21_X1   g10357(.A1(new_n10415_), .A2(new_n10367_), .B(new_n10421_), .ZN(new_n10422_));
  NAND2_X1   g10358(.A1(new_n10360_), .A2(new_n10279_), .ZN(new_n10423_));
  NAND2_X1   g10359(.A1(new_n10414_), .A2(new_n10346_), .ZN(new_n10424_));
  NAND2_X1   g10360(.A1(new_n10423_), .A2(new_n10424_), .ZN(new_n10425_));
  NOR3_X1    g10361(.A1(new_n10425_), .A2(new_n10359_), .A3(new_n10420_), .ZN(new_n10426_));
  OAI21_X1   g10362(.A1(new_n10426_), .A2(new_n10422_), .B(new_n10411_), .ZN(new_n10427_));
  INV_X1     g10363(.I(new_n10411_), .ZN(new_n10428_));
  OAI21_X1   g10364(.A1(new_n10425_), .A2(new_n10359_), .B(new_n10420_), .ZN(new_n10429_));
  NAND3_X1   g10365(.A1(new_n10415_), .A2(new_n10367_), .A3(new_n10421_), .ZN(new_n10430_));
  NAND3_X1   g10366(.A1(new_n10429_), .A2(new_n10428_), .A3(new_n10430_), .ZN(new_n10431_));
  NAND2_X1   g10367(.A1(new_n10427_), .A2(new_n10431_), .ZN(new_n10432_));
  OAI22_X1   g10368(.A1(new_n1409_), .A2(new_n9485_), .B1(new_n2367_), .B2(new_n9489_), .ZN(new_n10433_));
  NAND2_X1   g10369(.A1(new_n1334_), .A2(new_n9503_), .ZN(new_n10434_));
  AOI21_X1   g10370(.A1(new_n10433_), .A2(new_n10434_), .B(new_n9482_), .ZN(new_n10435_));
  NAND2_X1   g10371(.A1(new_n3654_), .A2(new_n10435_), .ZN(new_n10436_));
  XOR2_X1    g10372(.A1(new_n10436_), .A2(\a[2] ), .Z(new_n10437_));
  NAND2_X1   g10373(.A1(new_n10432_), .A2(new_n10437_), .ZN(new_n10438_));
  NAND2_X1   g10374(.A1(new_n9550_), .A2(new_n9567_), .ZN(new_n10439_));
  XOR2_X1    g10375(.A1(new_n9549_), .A2(\a[2] ), .Z(new_n10440_));
  NAND2_X1   g10376(.A1(new_n10440_), .A2(new_n9566_), .ZN(new_n10441_));
  NAND2_X1   g10377(.A1(new_n10439_), .A2(new_n10441_), .ZN(new_n10442_));
  OAI21_X1   g10378(.A1(new_n10432_), .A2(new_n10437_), .B(new_n10442_), .ZN(new_n10443_));
  AOI21_X1   g10379(.A1(new_n10375_), .A2(new_n10438_), .B(new_n10443_), .ZN(new_n10444_));
  OAI22_X1   g10380(.A1(new_n2367_), .A2(new_n9485_), .B1(new_n2451_), .B2(new_n9489_), .ZN(new_n10445_));
  NAND2_X1   g10381(.A1(new_n2412_), .A2(new_n9503_), .ZN(new_n10446_));
  AOI21_X1   g10382(.A1(new_n10445_), .A2(new_n10446_), .B(new_n9482_), .ZN(new_n10447_));
  NAND2_X1   g10383(.A1(new_n3403_), .A2(new_n10447_), .ZN(new_n10448_));
  XOR2_X1    g10384(.A1(new_n10448_), .A2(new_n4387_), .Z(new_n10449_));
  OAI21_X1   g10385(.A1(new_n10444_), .A2(new_n9568_), .B(new_n10449_), .ZN(new_n10450_));
  INV_X1     g10386(.I(new_n9568_), .ZN(new_n10451_));
  NOR3_X1    g10387(.A1(new_n10306_), .A2(new_n9573_), .A3(new_n10297_), .ZN(new_n10452_));
  AOI21_X1   g10388(.A1(new_n10296_), .A2(new_n10298_), .B(new_n9574_), .ZN(new_n10453_));
  NOR2_X1    g10389(.A1(new_n10372_), .A2(new_n10373_), .ZN(new_n10454_));
  OAI22_X1   g10390(.A1(new_n10453_), .A2(new_n10452_), .B1(new_n9573_), .B2(new_n10454_), .ZN(new_n10455_));
  AOI21_X1   g10391(.A1(new_n10429_), .A2(new_n10430_), .B(new_n10428_), .ZN(new_n10456_));
  NOR3_X1    g10392(.A1(new_n10426_), .A2(new_n10422_), .A3(new_n10411_), .ZN(new_n10457_));
  NOR2_X1    g10393(.A1(new_n10456_), .A2(new_n10457_), .ZN(new_n10458_));
  INV_X1     g10394(.I(new_n10437_), .ZN(new_n10459_));
  NOR2_X1    g10395(.A1(new_n10458_), .A2(new_n10459_), .ZN(new_n10460_));
  AOI22_X1   g10396(.A1(new_n10458_), .A2(new_n10459_), .B1(new_n10439_), .B2(new_n10441_), .ZN(new_n10461_));
  OAI21_X1   g10397(.A1(new_n10455_), .A2(new_n10460_), .B(new_n10461_), .ZN(new_n10462_));
  INV_X1     g10398(.I(new_n9551_), .ZN(new_n10463_));
  NOR2_X1    g10399(.A1(new_n9556_), .A2(new_n10463_), .ZN(new_n10464_));
  XOR2_X1    g10400(.A1(new_n9049_), .A2(new_n9016_), .Z(new_n10465_));
  NOR2_X1    g10401(.A1(new_n9050_), .A2(new_n9052_), .ZN(new_n10466_));
  NOR2_X1    g10402(.A1(new_n10466_), .A2(new_n9109_), .ZN(new_n10467_));
  AOI21_X1   g10403(.A1(new_n10465_), .A2(new_n9109_), .B(new_n10467_), .ZN(new_n10468_));
  INV_X1     g10404(.I(new_n10468_), .ZN(new_n10469_));
  OAI22_X1   g10405(.A1(new_n2251_), .A2(new_n6783_), .B1(new_n2351_), .B2(new_n6785_), .ZN(new_n10470_));
  NAND2_X1   g10406(.A1(new_n2310_), .A2(new_n6789_), .ZN(new_n10471_));
  AOI21_X1   g10407(.A1(new_n10471_), .A2(new_n10470_), .B(new_n6776_), .ZN(new_n10472_));
  NAND2_X1   g10408(.A1(new_n3914_), .A2(new_n10472_), .ZN(new_n10473_));
  XOR2_X1    g10409(.A1(new_n10473_), .A2(\a[8] ), .Z(new_n10474_));
  NOR2_X1    g10410(.A1(new_n10469_), .A2(new_n10474_), .ZN(new_n10475_));
  INV_X1     g10411(.I(new_n10474_), .ZN(new_n10476_));
  NOR2_X1    g10412(.A1(new_n10476_), .A2(new_n10468_), .ZN(new_n10477_));
  NOR3_X1    g10413(.A1(new_n10475_), .A2(new_n10477_), .A3(new_n10464_), .ZN(new_n10478_));
  INV_X1     g10414(.I(new_n10464_), .ZN(new_n10479_));
  NAND2_X1   g10415(.A1(new_n10476_), .A2(new_n10468_), .ZN(new_n10480_));
  NAND2_X1   g10416(.A1(new_n10469_), .A2(new_n10474_), .ZN(new_n10481_));
  AOI21_X1   g10417(.A1(new_n10481_), .A2(new_n10480_), .B(new_n10479_), .ZN(new_n10482_));
  NOR2_X1    g10418(.A1(new_n10478_), .A2(new_n10482_), .ZN(new_n10483_));
  OAI22_X1   g10419(.A1(new_n1409_), .A2(new_n6843_), .B1(new_n1333_), .B2(new_n6839_), .ZN(new_n10484_));
  NAND2_X1   g10420(.A1(new_n2359_), .A2(new_n6846_), .ZN(new_n10485_));
  AOI21_X1   g10421(.A1(new_n10484_), .A2(new_n10485_), .B(new_n6836_), .ZN(new_n10486_));
  NAND2_X1   g10422(.A1(new_n3828_), .A2(new_n10486_), .ZN(new_n10487_));
  XOR2_X1    g10423(.A1(new_n10487_), .A2(\a[5] ), .Z(new_n10488_));
  NAND2_X1   g10424(.A1(new_n10483_), .A2(new_n10488_), .ZN(new_n10489_));
  INV_X1     g10425(.I(new_n10483_), .ZN(new_n10490_));
  INV_X1     g10426(.I(new_n10488_), .ZN(new_n10491_));
  NAND2_X1   g10427(.A1(new_n10490_), .A2(new_n10491_), .ZN(new_n10492_));
  NAND2_X1   g10428(.A1(new_n10492_), .A2(new_n10489_), .ZN(new_n10493_));
  NAND2_X1   g10429(.A1(new_n10493_), .A2(new_n9564_), .ZN(new_n10494_));
  NAND3_X1   g10430(.A1(new_n10492_), .A2(new_n9563_), .A3(new_n10489_), .ZN(new_n10495_));
  AND2_X2    g10431(.A1(new_n10494_), .A2(new_n10495_), .Z(new_n10496_));
  NOR2_X1    g10432(.A1(new_n10496_), .A2(new_n10449_), .ZN(new_n10497_));
  NAND3_X1   g10433(.A1(new_n10462_), .A2(new_n10451_), .A3(new_n10497_), .ZN(new_n10498_));
  OAI22_X1   g10434(.A1(new_n2492_), .A2(new_n9489_), .B1(new_n2408_), .B2(new_n9485_), .ZN(new_n10499_));
  NAND2_X1   g10435(.A1(new_n2454_), .A2(new_n9503_), .ZN(new_n10500_));
  AOI21_X1   g10436(.A1(new_n10500_), .A2(new_n10499_), .B(new_n9482_), .ZN(new_n10501_));
  NAND2_X1   g10437(.A1(new_n3577_), .A2(new_n10501_), .ZN(new_n10502_));
  XOR2_X1    g10438(.A1(new_n10502_), .A2(new_n4387_), .Z(new_n10503_));
  INV_X1     g10439(.I(new_n10503_), .ZN(new_n10504_));
  AOI21_X1   g10440(.A1(new_n10450_), .A2(new_n10498_), .B(new_n10504_), .ZN(new_n10505_));
  INV_X1     g10441(.I(new_n10449_), .ZN(new_n10506_));
  AOI21_X1   g10442(.A1(new_n10462_), .A2(new_n10451_), .B(new_n10506_), .ZN(new_n10507_));
  NOR4_X1    g10443(.A1(new_n10444_), .A2(new_n9568_), .A3(new_n10449_), .A4(new_n10496_), .ZN(new_n10508_));
  AOI21_X1   g10444(.A1(new_n9564_), .A2(new_n10488_), .B(new_n10483_), .ZN(new_n10509_));
  NOR2_X1    g10445(.A1(new_n9564_), .A2(new_n10488_), .ZN(new_n10510_));
  NOR2_X1    g10446(.A1(new_n10509_), .A2(new_n10510_), .ZN(new_n10511_));
  XOR2_X1    g10447(.A1(new_n9115_), .A2(new_n9116_), .Z(new_n10512_));
  OAI21_X1   g10448(.A1(new_n9051_), .A2(new_n9052_), .B(new_n10512_), .ZN(new_n10513_));
  NOR2_X1    g10449(.A1(new_n9087_), .A2(new_n9092_), .ZN(new_n10514_));
  OAI21_X1   g10450(.A1(new_n10514_), .A2(new_n9118_), .B(new_n9112_), .ZN(new_n10515_));
  OAI22_X1   g10451(.A1(new_n1453_), .A2(new_n6785_), .B1(new_n2351_), .B2(new_n6788_), .ZN(new_n10516_));
  NAND2_X1   g10452(.A1(new_n2310_), .A2(new_n7530_), .ZN(new_n10517_));
  AOI21_X1   g10453(.A1(new_n10517_), .A2(new_n10516_), .B(new_n6776_), .ZN(new_n10518_));
  NAND2_X1   g10454(.A1(new_n4231_), .A2(new_n10518_), .ZN(new_n10519_));
  XOR2_X1    g10455(.A1(new_n10519_), .A2(\a[8] ), .Z(new_n10520_));
  OAI21_X1   g10456(.A1(new_n10478_), .A2(new_n10477_), .B(new_n10520_), .ZN(new_n10521_));
  OR3_X2     g10457(.A1(new_n10478_), .A2(new_n10477_), .A3(new_n10520_), .Z(new_n10522_));
  NAND2_X1   g10458(.A1(new_n10522_), .A2(new_n10521_), .ZN(new_n10523_));
  NAND3_X1   g10459(.A1(new_n10523_), .A2(new_n10513_), .A3(new_n10515_), .ZN(new_n10524_));
  NAND2_X1   g10460(.A1(new_n10513_), .A2(new_n10515_), .ZN(new_n10525_));
  NAND3_X1   g10461(.A1(new_n10522_), .A2(new_n10525_), .A3(new_n10521_), .ZN(new_n10526_));
  OAI22_X1   g10462(.A1(new_n1409_), .A2(new_n6913_), .B1(new_n2367_), .B2(new_n6839_), .ZN(new_n10527_));
  NAND2_X1   g10463(.A1(new_n1334_), .A2(new_n8799_), .ZN(new_n10528_));
  AOI21_X1   g10464(.A1(new_n10527_), .A2(new_n10528_), .B(new_n6836_), .ZN(new_n10529_));
  NAND2_X1   g10465(.A1(new_n3654_), .A2(new_n10529_), .ZN(new_n10530_));
  XOR2_X1    g10466(.A1(new_n10530_), .A2(\a[5] ), .Z(new_n10531_));
  INV_X1     g10467(.I(new_n10531_), .ZN(new_n10532_));
  NAND3_X1   g10468(.A1(new_n10524_), .A2(new_n10526_), .A3(new_n10532_), .ZN(new_n10533_));
  INV_X1     g10469(.I(new_n10533_), .ZN(new_n10534_));
  AOI21_X1   g10470(.A1(new_n10524_), .A2(new_n10526_), .B(new_n10532_), .ZN(new_n10535_));
  OAI21_X1   g10471(.A1(new_n10534_), .A2(new_n10535_), .B(new_n10511_), .ZN(new_n10536_));
  INV_X1     g10472(.I(new_n10511_), .ZN(new_n10537_));
  INV_X1     g10473(.I(new_n10535_), .ZN(new_n10538_));
  NAND3_X1   g10474(.A1(new_n10538_), .A2(new_n10537_), .A3(new_n10533_), .ZN(new_n10539_));
  AOI21_X1   g10475(.A1(new_n10539_), .A2(new_n10536_), .B(new_n10503_), .ZN(new_n10540_));
  INV_X1     g10476(.I(new_n10540_), .ZN(new_n10541_));
  NOR3_X1    g10477(.A1(new_n10508_), .A2(new_n10507_), .A3(new_n10541_), .ZN(new_n10542_));
  NAND2_X1   g10478(.A1(new_n9127_), .A2(new_n9121_), .ZN(new_n10543_));
  AND2_X2    g10479(.A1(new_n10543_), .A2(new_n9294_), .Z(new_n10544_));
  NAND2_X1   g10480(.A1(new_n10524_), .A2(new_n10526_), .ZN(new_n10545_));
  OAI21_X1   g10481(.A1(new_n10509_), .A2(new_n10510_), .B(new_n10532_), .ZN(new_n10546_));
  NAND2_X1   g10482(.A1(new_n10511_), .A2(new_n10531_), .ZN(new_n10547_));
  INV_X1     g10483(.I(new_n10547_), .ZN(new_n10548_));
  OAI21_X1   g10484(.A1(new_n10548_), .A2(new_n10545_), .B(new_n10546_), .ZN(new_n10549_));
  OAI22_X1   g10485(.A1(new_n2367_), .A2(new_n6843_), .B1(new_n2408_), .B2(new_n6839_), .ZN(new_n10550_));
  NAND2_X1   g10486(.A1(new_n1334_), .A2(new_n6846_), .ZN(new_n10551_));
  AOI21_X1   g10487(.A1(new_n10550_), .A2(new_n10551_), .B(new_n6836_), .ZN(new_n10552_));
  NAND2_X1   g10488(.A1(new_n3708_), .A2(new_n10552_), .ZN(new_n10553_));
  XOR2_X1    g10489(.A1(new_n10553_), .A2(\a[5] ), .Z(new_n10554_));
  INV_X1     g10490(.I(new_n10554_), .ZN(new_n10555_));
  NOR2_X1    g10491(.A1(new_n10549_), .A2(new_n10555_), .ZN(new_n10556_));
  INV_X1     g10492(.I(new_n10556_), .ZN(new_n10557_));
  NAND2_X1   g10493(.A1(new_n10549_), .A2(new_n10555_), .ZN(new_n10558_));
  AOI21_X1   g10494(.A1(new_n10557_), .A2(new_n10558_), .B(new_n10544_), .ZN(new_n10559_));
  INV_X1     g10495(.I(new_n10544_), .ZN(new_n10560_));
  NAND2_X1   g10496(.A1(new_n10549_), .A2(new_n10554_), .ZN(new_n10561_));
  NOR2_X1    g10497(.A1(new_n10549_), .A2(new_n10554_), .ZN(new_n10562_));
  INV_X1     g10498(.I(new_n10562_), .ZN(new_n10563_));
  AOI21_X1   g10499(.A1(new_n10563_), .A2(new_n10561_), .B(new_n10560_), .ZN(new_n10564_));
  OAI22_X1   g10500(.A1(new_n1121_), .A2(new_n9489_), .B1(new_n2451_), .B2(new_n9485_), .ZN(new_n10565_));
  NAND2_X1   g10501(.A1(new_n2496_), .A2(new_n9503_), .ZN(new_n10566_));
  AOI21_X1   g10502(.A1(new_n10565_), .A2(new_n10566_), .B(new_n9482_), .ZN(new_n10567_));
  NAND2_X1   g10503(.A1(new_n3393_), .A2(new_n10567_), .ZN(new_n10568_));
  XOR2_X1    g10504(.A1(new_n10568_), .A2(\a[2] ), .Z(new_n10569_));
  OAI21_X1   g10505(.A1(new_n10559_), .A2(new_n10564_), .B(new_n10569_), .ZN(new_n10570_));
  OAI21_X1   g10506(.A1(new_n10542_), .A2(new_n10505_), .B(new_n10570_), .ZN(new_n10571_));
  NOR3_X1    g10507(.A1(new_n10559_), .A2(new_n10564_), .A3(new_n10569_), .ZN(new_n10572_));
  INV_X1     g10508(.I(new_n10572_), .ZN(new_n10573_));
  NOR2_X1    g10509(.A1(new_n9299_), .A2(new_n9295_), .ZN(new_n10574_));
  XNOR2_X1   g10510(.A1(new_n10574_), .A2(new_n9163_), .ZN(new_n10575_));
  NOR2_X1    g10511(.A1(new_n10575_), .A2(new_n9294_), .ZN(new_n10576_));
  AOI21_X1   g10512(.A1(new_n9164_), .A2(new_n9301_), .B(new_n9128_), .ZN(new_n10577_));
  OAI22_X1   g10513(.A1(new_n2367_), .A2(new_n6913_), .B1(new_n2451_), .B2(new_n6839_), .ZN(new_n10578_));
  NAND2_X1   g10514(.A1(new_n2412_), .A2(new_n8799_), .ZN(new_n10579_));
  AOI21_X1   g10515(.A1(new_n10578_), .A2(new_n10579_), .B(new_n6836_), .ZN(new_n10580_));
  NAND2_X1   g10516(.A1(new_n3403_), .A2(new_n10580_), .ZN(new_n10581_));
  XOR2_X1    g10517(.A1(new_n10581_), .A2(\a[5] ), .Z(new_n10582_));
  OR3_X2     g10518(.A1(new_n10576_), .A2(new_n10577_), .A3(new_n10582_), .Z(new_n10583_));
  OAI21_X1   g10519(.A1(new_n10576_), .A2(new_n10577_), .B(new_n10582_), .ZN(new_n10584_));
  NAND2_X1   g10520(.A1(new_n10583_), .A2(new_n10584_), .ZN(new_n10585_));
  NAND2_X1   g10521(.A1(new_n10549_), .A2(new_n10544_), .ZN(new_n10586_));
  NOR2_X1    g10522(.A1(new_n10586_), .A2(new_n10585_), .ZN(new_n10587_));
  INV_X1     g10523(.I(new_n10587_), .ZN(new_n10588_));
  NAND2_X1   g10524(.A1(new_n10586_), .A2(new_n10585_), .ZN(new_n10589_));
  NOR2_X1    g10525(.A1(new_n10549_), .A2(new_n10544_), .ZN(new_n10590_));
  INV_X1     g10526(.I(new_n10590_), .ZN(new_n10591_));
  NAND3_X1   g10527(.A1(new_n10591_), .A2(new_n10586_), .A3(new_n10554_), .ZN(new_n10592_));
  NAND3_X1   g10528(.A1(new_n10592_), .A2(new_n10588_), .A3(new_n10589_), .ZN(new_n10593_));
  NAND4_X1   g10529(.A1(new_n10591_), .A2(new_n10586_), .A3(new_n10585_), .A4(new_n10554_), .ZN(new_n10594_));
  OAI22_X1   g10530(.A1(new_n1180_), .A2(new_n9489_), .B1(new_n2492_), .B2(new_n9485_), .ZN(new_n10595_));
  NAND2_X1   g10531(.A1(new_n1122_), .A2(new_n9503_), .ZN(new_n10596_));
  AOI21_X1   g10532(.A1(new_n10596_), .A2(new_n10595_), .B(new_n9482_), .ZN(new_n10597_));
  NAND2_X1   g10533(.A1(new_n3330_), .A2(new_n10597_), .ZN(new_n10598_));
  XOR2_X1    g10534(.A1(new_n10598_), .A2(\a[2] ), .Z(new_n10599_));
  INV_X1     g10535(.I(new_n10599_), .ZN(new_n10600_));
  AOI21_X1   g10536(.A1(new_n10593_), .A2(new_n10594_), .B(new_n10600_), .ZN(new_n10601_));
  AOI21_X1   g10537(.A1(new_n10571_), .A2(new_n10573_), .B(new_n10601_), .ZN(new_n10602_));
  INV_X1     g10538(.I(new_n10589_), .ZN(new_n10603_));
  INV_X1     g10539(.I(new_n10586_), .ZN(new_n10604_));
  NOR3_X1    g10540(.A1(new_n10604_), .A2(new_n10590_), .A3(new_n10555_), .ZN(new_n10605_));
  NOR3_X1    g10541(.A1(new_n10605_), .A2(new_n10603_), .A3(new_n10587_), .ZN(new_n10606_));
  INV_X1     g10542(.I(new_n10594_), .ZN(new_n10607_));
  NOR3_X1    g10543(.A1(new_n10606_), .A2(new_n10607_), .A3(new_n10599_), .ZN(new_n10608_));
  NAND2_X1   g10544(.A1(new_n9190_), .A2(new_n9182_), .ZN(new_n10609_));
  XOR2_X1    g10545(.A1(new_n10609_), .A2(new_n9195_), .Z(new_n10610_));
  NAND2_X1   g10546(.A1(new_n9308_), .A2(new_n9197_), .ZN(new_n10611_));
  NAND2_X1   g10547(.A1(new_n10611_), .A2(new_n9167_), .ZN(new_n10612_));
  OAI21_X1   g10548(.A1(new_n10610_), .A2(new_n9167_), .B(new_n10612_), .ZN(new_n10613_));
  INV_X1     g10549(.I(new_n10613_), .ZN(new_n10614_));
  AOI21_X1   g10550(.A1(new_n10549_), .A2(new_n10544_), .B(new_n10554_), .ZN(new_n10615_));
  NAND2_X1   g10551(.A1(new_n10583_), .A2(new_n10584_), .ZN(new_n10616_));
  OAI22_X1   g10552(.A1(new_n2492_), .A2(new_n6839_), .B1(new_n2408_), .B2(new_n6913_), .ZN(new_n10617_));
  NAND2_X1   g10553(.A1(new_n2454_), .A2(new_n8799_), .ZN(new_n10618_));
  AOI21_X1   g10554(.A1(new_n10618_), .A2(new_n10617_), .B(new_n6836_), .ZN(new_n10619_));
  NAND2_X1   g10555(.A1(new_n3577_), .A2(new_n10619_), .ZN(new_n10620_));
  XOR2_X1    g10556(.A1(new_n10620_), .A2(\a[5] ), .Z(new_n10621_));
  OAI21_X1   g10557(.A1(new_n10615_), .A2(new_n10616_), .B(new_n10621_), .ZN(new_n10622_));
  INV_X1     g10558(.I(new_n10622_), .ZN(new_n10623_));
  NOR3_X1    g10559(.A1(new_n10615_), .A2(new_n10616_), .A3(new_n10621_), .ZN(new_n10624_));
  OAI21_X1   g10560(.A1(new_n10623_), .A2(new_n10624_), .B(new_n10614_), .ZN(new_n10625_));
  INV_X1     g10561(.I(new_n10624_), .ZN(new_n10626_));
  NAND3_X1   g10562(.A1(new_n10626_), .A2(new_n10622_), .A3(new_n10613_), .ZN(new_n10627_));
  NAND2_X1   g10563(.A1(new_n10625_), .A2(new_n10627_), .ZN(new_n10628_));
  OAI22_X1   g10564(.A1(new_n1008_), .A2(new_n9489_), .B1(new_n1121_), .B2(new_n9485_), .ZN(new_n10629_));
  NAND2_X1   g10565(.A1(new_n1181_), .A2(new_n9503_), .ZN(new_n10630_));
  AOI21_X1   g10566(.A1(new_n10629_), .A2(new_n10630_), .B(new_n9482_), .ZN(new_n10631_));
  NAND2_X1   g10567(.A1(new_n3562_), .A2(new_n10631_), .ZN(new_n10632_));
  XOR2_X1    g10568(.A1(new_n10632_), .A2(new_n4387_), .Z(new_n10633_));
  INV_X1     g10569(.I(new_n10633_), .ZN(new_n10634_));
  NAND2_X1   g10570(.A1(new_n10628_), .A2(new_n10634_), .ZN(new_n10635_));
  OAI21_X1   g10571(.A1(new_n10602_), .A2(new_n10608_), .B(new_n10635_), .ZN(new_n10636_));
  NOR2_X1    g10572(.A1(new_n10628_), .A2(new_n10634_), .ZN(new_n10637_));
  INV_X1     g10573(.I(new_n10637_), .ZN(new_n10638_));
  OAI22_X1   g10574(.A1(new_n896_), .A2(new_n9489_), .B1(new_n1180_), .B2(new_n9485_), .ZN(new_n10639_));
  NAND2_X1   g10575(.A1(new_n2504_), .A2(new_n9503_), .ZN(new_n10640_));
  AOI21_X1   g10576(.A1(new_n10640_), .A2(new_n10639_), .B(new_n9482_), .ZN(new_n10641_));
  NAND2_X1   g10577(.A1(new_n3596_), .A2(new_n10641_), .ZN(new_n10642_));
  XOR2_X1    g10578(.A1(new_n10642_), .A2(\a[2] ), .Z(new_n10643_));
  AOI21_X1   g10579(.A1(new_n10636_), .A2(new_n10638_), .B(new_n10643_), .ZN(new_n10644_));
  OAI21_X1   g10580(.A1(new_n10508_), .A2(new_n10507_), .B(new_n10503_), .ZN(new_n10645_));
  NAND3_X1   g10581(.A1(new_n10450_), .A2(new_n10498_), .A3(new_n10540_), .ZN(new_n10646_));
  INV_X1     g10582(.I(new_n10558_), .ZN(new_n10647_));
  OAI21_X1   g10583(.A1(new_n10647_), .A2(new_n10556_), .B(new_n10560_), .ZN(new_n10648_));
  INV_X1     g10584(.I(new_n10545_), .ZN(new_n10649_));
  INV_X1     g10585(.I(new_n10546_), .ZN(new_n10650_));
  AOI21_X1   g10586(.A1(new_n10649_), .A2(new_n10547_), .B(new_n10650_), .ZN(new_n10651_));
  NOR2_X1    g10587(.A1(new_n10651_), .A2(new_n10555_), .ZN(new_n10652_));
  OAI21_X1   g10588(.A1(new_n10652_), .A2(new_n10562_), .B(new_n10544_), .ZN(new_n10653_));
  INV_X1     g10589(.I(new_n10569_), .ZN(new_n10654_));
  AOI21_X1   g10590(.A1(new_n10648_), .A2(new_n10653_), .B(new_n10654_), .ZN(new_n10655_));
  AOI21_X1   g10591(.A1(new_n10645_), .A2(new_n10646_), .B(new_n10655_), .ZN(new_n10656_));
  OAI21_X1   g10592(.A1(new_n10606_), .A2(new_n10607_), .B(new_n10599_), .ZN(new_n10657_));
  OAI21_X1   g10593(.A1(new_n10656_), .A2(new_n10572_), .B(new_n10657_), .ZN(new_n10658_));
  INV_X1     g10594(.I(new_n10608_), .ZN(new_n10659_));
  AOI21_X1   g10595(.A1(new_n10626_), .A2(new_n10622_), .B(new_n10613_), .ZN(new_n10660_));
  NOR3_X1    g10596(.A1(new_n10623_), .A2(new_n10614_), .A3(new_n10624_), .ZN(new_n10661_));
  NOR2_X1    g10597(.A1(new_n10660_), .A2(new_n10661_), .ZN(new_n10662_));
  NOR2_X1    g10598(.A1(new_n10662_), .A2(new_n10633_), .ZN(new_n10663_));
  AOI21_X1   g10599(.A1(new_n10658_), .A2(new_n10659_), .B(new_n10663_), .ZN(new_n10664_));
  NAND2_X1   g10600(.A1(new_n9250_), .A2(new_n9247_), .ZN(new_n10665_));
  XOR2_X1    g10601(.A1(new_n9253_), .A2(new_n65_), .Z(new_n10666_));
  NOR2_X1    g10602(.A1(new_n10665_), .A2(new_n10666_), .ZN(new_n10667_));
  OAI21_X1   g10603(.A1(new_n9255_), .A2(new_n10667_), .B(new_n10643_), .ZN(new_n10668_));
  NOR3_X1    g10604(.A1(new_n10664_), .A2(new_n10637_), .A3(new_n10668_), .ZN(new_n10669_));
  OAI22_X1   g10605(.A1(new_n813_), .A2(new_n9489_), .B1(new_n1008_), .B2(new_n9485_), .ZN(new_n10670_));
  NAND2_X1   g10606(.A1(new_n897_), .A2(new_n9503_), .ZN(new_n10671_));
  AOI21_X1   g10607(.A1(new_n10670_), .A2(new_n10671_), .B(new_n9482_), .ZN(new_n10672_));
  NAND2_X1   g10608(.A1(new_n2917_), .A2(new_n10672_), .ZN(new_n10673_));
  XOR2_X1    g10609(.A1(new_n10673_), .A2(\a[2] ), .Z(new_n10674_));
  INV_X1     g10610(.I(new_n10674_), .ZN(new_n10675_));
  OAI21_X1   g10611(.A1(new_n10644_), .A2(new_n10669_), .B(new_n10675_), .ZN(new_n10676_));
  INV_X1     g10612(.I(new_n10643_), .ZN(new_n10677_));
  OAI21_X1   g10613(.A1(new_n10664_), .A2(new_n10637_), .B(new_n10677_), .ZN(new_n10678_));
  INV_X1     g10614(.I(new_n10668_), .ZN(new_n10679_));
  NAND3_X1   g10615(.A1(new_n10636_), .A2(new_n10638_), .A3(new_n10679_), .ZN(new_n10680_));
  NOR3_X1    g10616(.A1(new_n9332_), .A2(new_n9397_), .A3(new_n9256_), .ZN(new_n10681_));
  AOI21_X1   g10617(.A1(new_n9333_), .A2(new_n9396_), .B(new_n9255_), .ZN(new_n10682_));
  OAI21_X1   g10618(.A1(new_n10681_), .A2(new_n10682_), .B(new_n10674_), .ZN(new_n10683_));
  INV_X1     g10619(.I(new_n10683_), .ZN(new_n10684_));
  NAND3_X1   g10620(.A1(new_n10680_), .A2(new_n10678_), .A3(new_n10684_), .ZN(new_n10685_));
  OAI22_X1   g10621(.A1(new_n2559_), .A2(new_n9489_), .B1(new_n896_), .B2(new_n9485_), .ZN(new_n10686_));
  NAND2_X1   g10622(.A1(new_n814_), .A2(new_n9503_), .ZN(new_n10687_));
  AOI21_X1   g10623(.A1(new_n10686_), .A2(new_n10687_), .B(new_n9482_), .ZN(new_n10688_));
  NAND2_X1   g10624(.A1(new_n3624_), .A2(new_n10688_), .ZN(new_n10689_));
  XOR2_X1    g10625(.A1(new_n10689_), .A2(\a[2] ), .Z(new_n10690_));
  AOI21_X1   g10626(.A1(new_n10676_), .A2(new_n10685_), .B(new_n10690_), .ZN(new_n10691_));
  AOI21_X1   g10627(.A1(new_n10680_), .A2(new_n10678_), .B(new_n10674_), .ZN(new_n10692_));
  NOR3_X1    g10628(.A1(new_n10644_), .A2(new_n10669_), .A3(new_n10683_), .ZN(new_n10693_));
  INV_X1     g10629(.I(new_n10690_), .ZN(new_n10694_));
  NAND2_X1   g10630(.A1(new_n9383_), .A2(new_n9384_), .ZN(new_n10695_));
  XOR2_X1    g10631(.A1(new_n10695_), .A2(new_n9398_), .Z(new_n10696_));
  NOR4_X1    g10632(.A1(new_n10692_), .A2(new_n10693_), .A3(new_n10694_), .A4(new_n10696_), .ZN(new_n10697_));
  XOR2_X1    g10633(.A1(new_n9391_), .A2(new_n9393_), .Z(new_n10698_));
  INV_X1     g10634(.I(new_n10698_), .ZN(new_n10699_));
  XOR2_X1    g10635(.A1(new_n9391_), .A2(new_n9439_), .Z(new_n10700_));
  NOR2_X1    g10636(.A1(new_n9400_), .A2(new_n10700_), .ZN(new_n10701_));
  AOI21_X1   g10637(.A1(new_n9400_), .A2(new_n10699_), .B(new_n10701_), .ZN(new_n10702_));
  INV_X1     g10638(.I(new_n10702_), .ZN(new_n10703_));
  OAI22_X1   g10639(.A1(new_n813_), .A2(new_n9485_), .B1(new_n529_), .B2(new_n9489_), .ZN(new_n10704_));
  NAND2_X1   g10640(.A1(new_n2563_), .A2(new_n9503_), .ZN(new_n10705_));
  AOI21_X1   g10641(.A1(new_n10705_), .A2(new_n10704_), .B(new_n9482_), .ZN(new_n10706_));
  NAND2_X1   g10642(.A1(new_n3051_), .A2(new_n10706_), .ZN(new_n10707_));
  XOR2_X1    g10643(.A1(new_n10707_), .A2(\a[2] ), .Z(new_n10708_));
  NAND2_X1   g10644(.A1(new_n10703_), .A2(new_n10708_), .ZN(new_n10709_));
  OAI21_X1   g10645(.A1(new_n10697_), .A2(new_n10691_), .B(new_n10709_), .ZN(new_n10710_));
  NOR2_X1    g10646(.A1(new_n10703_), .A2(new_n10708_), .ZN(new_n10711_));
  INV_X1     g10647(.I(new_n10711_), .ZN(new_n10712_));
  NOR2_X1    g10648(.A1(new_n9386_), .A2(new_n9391_), .ZN(new_n10713_));
  NAND2_X1   g10649(.A1(new_n9436_), .A2(new_n9437_), .ZN(new_n10714_));
  XOR2_X1    g10650(.A1(new_n9404_), .A2(new_n10714_), .Z(new_n10715_));
  NAND2_X1   g10651(.A1(new_n10715_), .A2(new_n10713_), .ZN(new_n10716_));
  INV_X1     g10652(.I(new_n10713_), .ZN(new_n10717_));
  XOR2_X1    g10653(.A1(new_n9444_), .A2(new_n10714_), .Z(new_n10718_));
  NAND2_X1   g10654(.A1(new_n10718_), .A2(new_n10717_), .ZN(new_n10719_));
  OAI22_X1   g10655(.A1(new_n2559_), .A2(new_n9485_), .B1(new_n694_), .B2(new_n9489_), .ZN(new_n10720_));
  NAND2_X1   g10656(.A1(new_n2567_), .A2(new_n9503_), .ZN(new_n10721_));
  AOI21_X1   g10657(.A1(new_n10720_), .A2(new_n10721_), .B(new_n9482_), .ZN(new_n10722_));
  NAND2_X1   g10658(.A1(new_n2759_), .A2(new_n10722_), .ZN(new_n10723_));
  XOR2_X1    g10659(.A1(new_n10723_), .A2(\a[2] ), .Z(new_n10724_));
  INV_X1     g10660(.I(new_n10724_), .ZN(new_n10725_));
  AOI21_X1   g10661(.A1(new_n10716_), .A2(new_n10719_), .B(new_n10725_), .ZN(new_n10726_));
  AOI21_X1   g10662(.A1(new_n10710_), .A2(new_n10712_), .B(new_n10726_), .ZN(new_n10727_));
  NOR2_X1    g10663(.A1(new_n10718_), .A2(new_n10717_), .ZN(new_n10728_));
  NOR2_X1    g10664(.A1(new_n10715_), .A2(new_n10713_), .ZN(new_n10729_));
  NOR3_X1    g10665(.A1(new_n10729_), .A2(new_n10728_), .A3(new_n10724_), .ZN(new_n10730_));
  NOR3_X1    g10666(.A1(new_n10727_), .A2(new_n9544_), .A3(new_n10730_), .ZN(new_n10731_));
  OAI22_X1   g10667(.A1(new_n694_), .A2(new_n9485_), .B1(new_n2665_), .B2(new_n9489_), .ZN(new_n10732_));
  NAND2_X1   g10668(.A1(new_n2615_), .A2(new_n9503_), .ZN(new_n10733_));
  AOI21_X1   g10669(.A1(new_n10732_), .A2(new_n10733_), .B(new_n9482_), .ZN(new_n10734_));
  NAND2_X1   g10670(.A1(new_n3188_), .A2(new_n10734_), .ZN(new_n10735_));
  XOR2_X1    g10671(.A1(new_n10735_), .A2(new_n4387_), .Z(new_n10736_));
  NOR2_X1    g10672(.A1(new_n10736_), .A2(new_n9421_), .ZN(new_n10737_));
  XOR2_X1    g10673(.A1(new_n10735_), .A2(\a[2] ), .Z(new_n10738_));
  NOR2_X1    g10674(.A1(new_n10738_), .A2(new_n9452_), .ZN(new_n10739_));
  OR2_X2     g10675(.A1(new_n10737_), .A2(new_n10739_), .Z(new_n10740_));
  NAND2_X1   g10676(.A1(new_n10738_), .A2(new_n9421_), .ZN(new_n10741_));
  NAND2_X1   g10677(.A1(new_n10736_), .A2(new_n9452_), .ZN(new_n10742_));
  AOI21_X1   g10678(.A1(new_n10741_), .A2(new_n10742_), .B(new_n9413_), .ZN(new_n10743_));
  AOI21_X1   g10679(.A1(new_n10740_), .A2(new_n9413_), .B(new_n10743_), .ZN(new_n10744_));
  XOR2_X1    g10680(.A1(new_n9449_), .A2(new_n9452_), .Z(new_n10745_));
  NAND2_X1   g10681(.A1(new_n10745_), .A2(new_n10738_), .ZN(new_n10746_));
  NAND3_X1   g10682(.A1(new_n9544_), .A2(new_n10744_), .A3(new_n10746_), .ZN(new_n10747_));
  NAND2_X1   g10683(.A1(new_n2615_), .A2(new_n6925_), .ZN(new_n10748_));
  NAND2_X1   g10684(.A1(new_n2728_), .A2(new_n9488_), .ZN(new_n10749_));
  AOI21_X1   g10685(.A1(new_n2664_), .A2(new_n9503_), .B(new_n9482_), .ZN(new_n10750_));
  NAND4_X1   g10686(.A1(new_n2733_), .A2(new_n10748_), .A3(new_n10749_), .A4(new_n10750_), .ZN(new_n10751_));
  XOR2_X1    g10687(.A1(new_n10751_), .A2(new_n4387_), .Z(new_n10752_));
  OAI21_X1   g10688(.A1(new_n10731_), .A2(new_n10747_), .B(new_n10752_), .ZN(new_n10753_));
  OAI21_X1   g10689(.A1(new_n10692_), .A2(new_n10693_), .B(new_n10694_), .ZN(new_n10754_));
  NOR2_X1    g10690(.A1(new_n10696_), .A2(new_n10694_), .ZN(new_n10755_));
  NAND3_X1   g10691(.A1(new_n10676_), .A2(new_n10685_), .A3(new_n10755_), .ZN(new_n10756_));
  INV_X1     g10692(.I(new_n10709_), .ZN(new_n10757_));
  AOI21_X1   g10693(.A1(new_n10754_), .A2(new_n10756_), .B(new_n10757_), .ZN(new_n10758_));
  OAI21_X1   g10694(.A1(new_n10729_), .A2(new_n10728_), .B(new_n10724_), .ZN(new_n10759_));
  OAI21_X1   g10695(.A1(new_n10758_), .A2(new_n10711_), .B(new_n10759_), .ZN(new_n10760_));
  INV_X1     g10696(.I(new_n10730_), .ZN(new_n10761_));
  NAND3_X1   g10697(.A1(new_n10760_), .A2(new_n9543_), .A3(new_n10761_), .ZN(new_n10762_));
  OAI21_X1   g10698(.A1(new_n10737_), .A2(new_n10739_), .B(new_n9413_), .ZN(new_n10763_));
  AND2_X2    g10699(.A1(new_n10741_), .A2(new_n10742_), .Z(new_n10764_));
  OAI21_X1   g10700(.A1(new_n10764_), .A2(new_n9413_), .B(new_n10763_), .ZN(new_n10765_));
  XOR2_X1    g10701(.A1(new_n9449_), .A2(new_n9421_), .Z(new_n10766_));
  NOR2_X1    g10702(.A1(new_n10766_), .A2(new_n10736_), .ZN(new_n10767_));
  NOR3_X1    g10703(.A1(new_n10765_), .A2(new_n9543_), .A3(new_n10767_), .ZN(new_n10768_));
  INV_X1     g10704(.I(new_n10752_), .ZN(new_n10769_));
  NAND3_X1   g10705(.A1(new_n10762_), .A2(new_n10768_), .A3(new_n10769_), .ZN(new_n10770_));
  AOI21_X1   g10706(.A1(new_n10753_), .A2(new_n10770_), .B(new_n9531_), .ZN(new_n10771_));
  AOI21_X1   g10707(.A1(new_n10762_), .A2(new_n10768_), .B(new_n10769_), .ZN(new_n10772_));
  NOR3_X1    g10708(.A1(new_n10731_), .A2(new_n10747_), .A3(new_n10752_), .ZN(new_n10773_));
  NOR3_X1    g10709(.A1(new_n10773_), .A2(new_n10772_), .A3(new_n9530_), .ZN(new_n10774_));
  NOR2_X1    g10710(.A1(new_n10774_), .A2(new_n10771_), .ZN(new_n10775_));
  AOI21_X1   g10711(.A1(new_n9526_), .A2(new_n9525_), .B(new_n9524_), .ZN(new_n10776_));
  NOR2_X1    g10712(.A1(new_n9516_), .A2(new_n10776_), .ZN(new_n10777_));
  INV_X1     g10713(.I(new_n9540_), .ZN(new_n10778_));
  NOR2_X1    g10714(.A1(new_n10778_), .A2(new_n9541_), .ZN(new_n10779_));
  NOR3_X1    g10715(.A1(new_n10727_), .A2(new_n9536_), .A3(new_n10730_), .ZN(new_n10780_));
  AOI21_X1   g10716(.A1(new_n10760_), .A2(new_n10761_), .B(new_n9537_), .ZN(new_n10781_));
  OAI21_X1   g10717(.A1(new_n10780_), .A2(new_n10781_), .B(new_n10779_), .ZN(new_n10782_));
  NOR2_X1    g10718(.A1(new_n10782_), .A2(new_n10765_), .ZN(new_n10783_));
  NAND3_X1   g10719(.A1(new_n10760_), .A2(new_n9537_), .A3(new_n10761_), .ZN(new_n10784_));
  OAI21_X1   g10720(.A1(new_n10727_), .A2(new_n10730_), .B(new_n9536_), .ZN(new_n10785_));
  NAND2_X1   g10721(.A1(new_n10785_), .A2(new_n10784_), .ZN(new_n10786_));
  AOI21_X1   g10722(.A1(new_n10786_), .A2(new_n10779_), .B(new_n10744_), .ZN(new_n10787_));
  AOI21_X1   g10723(.A1(new_n10760_), .A2(new_n10761_), .B(new_n9536_), .ZN(new_n10788_));
  INV_X1     g10724(.I(new_n10788_), .ZN(new_n10789_));
  NOR3_X1    g10725(.A1(new_n10783_), .A2(new_n10787_), .A3(new_n10789_), .ZN(new_n10790_));
  NAND3_X1   g10726(.A1(new_n10786_), .A2(new_n10779_), .A3(new_n10744_), .ZN(new_n10791_));
  NAND2_X1   g10727(.A1(new_n10782_), .A2(new_n10765_), .ZN(new_n10792_));
  AOI21_X1   g10728(.A1(new_n10792_), .A2(new_n10791_), .B(new_n10788_), .ZN(new_n10793_));
  NOR2_X1    g10729(.A1(new_n10790_), .A2(new_n10793_), .ZN(new_n10794_));
  NOR3_X1    g10730(.A1(new_n10775_), .A2(new_n9529_), .A3(new_n10777_), .ZN(new_n10795_));
  NOR3_X1    g10731(.A1(new_n9527_), .A2(new_n9520_), .A3(new_n9523_), .ZN(new_n10796_));
  AOI21_X1   g10732(.A1(new_n9498_), .A2(new_n9501_), .B(new_n9516_), .ZN(new_n10797_));
  NOR2_X1    g10733(.A1(new_n10797_), .A2(new_n10796_), .ZN(new_n10798_));
  NAND2_X1   g10734(.A1(new_n10775_), .A2(new_n10798_), .ZN(new_n10799_));
  INV_X1     g10735(.I(new_n10777_), .ZN(new_n10800_));
  NOR4_X1    g10736(.A1(new_n10775_), .A2(new_n10790_), .A3(new_n10793_), .A4(new_n10798_), .ZN(new_n10801_));
  OAI21_X1   g10737(.A1(new_n10801_), .A2(new_n10800_), .B(new_n10799_), .ZN(new_n10802_));
  INV_X1     g10738(.I(new_n9471_), .ZN(new_n10803_));
  NAND3_X1   g10739(.A1(new_n9462_), .A2(new_n9432_), .A3(new_n9466_), .ZN(new_n10804_));
  NOR2_X1    g10740(.A1(new_n9455_), .A2(new_n9430_), .ZN(new_n10805_));
  NOR2_X1    g10741(.A1(new_n9424_), .A2(new_n9460_), .ZN(new_n10806_));
  OAI21_X1   g10742(.A1(new_n10805_), .A2(new_n10806_), .B(new_n9465_), .ZN(new_n10807_));
  AOI21_X1   g10743(.A1(new_n10807_), .A2(new_n10804_), .B(\a[5] ), .ZN(new_n10808_));
  NOR3_X1    g10744(.A1(new_n10805_), .A2(new_n10806_), .A3(new_n9465_), .ZN(new_n10809_));
  AOI21_X1   g10745(.A1(new_n9462_), .A2(new_n9432_), .B(new_n9466_), .ZN(new_n10810_));
  NOR3_X1    g10746(.A1(new_n10809_), .A2(new_n10810_), .A3(new_n65_), .ZN(new_n10811_));
  OAI21_X1   g10747(.A1(new_n10811_), .A2(new_n10808_), .B(new_n10803_), .ZN(new_n10812_));
  OAI21_X1   g10748(.A1(new_n10809_), .A2(new_n10810_), .B(new_n65_), .ZN(new_n10813_));
  NAND3_X1   g10749(.A1(new_n10807_), .A2(new_n10804_), .A3(\a[5] ), .ZN(new_n10814_));
  NAND3_X1   g10750(.A1(new_n10813_), .A2(new_n10814_), .A3(new_n9471_), .ZN(new_n10815_));
  NOR2_X1    g10751(.A1(new_n9494_), .A2(new_n9492_), .ZN(new_n10816_));
  INV_X1     g10752(.I(new_n10816_), .ZN(new_n10817_));
  NAND2_X1   g10753(.A1(new_n9424_), .A2(new_n9481_), .ZN(new_n10818_));
  NAND2_X1   g10754(.A1(new_n9455_), .A2(new_n9480_), .ZN(new_n10819_));
  AOI21_X1   g10755(.A1(new_n10819_), .A2(new_n10818_), .B(new_n10817_), .ZN(new_n10820_));
  NAND2_X1   g10756(.A1(new_n3168_), .A2(new_n6925_), .ZN(new_n10821_));
  NAND2_X1   g10757(.A1(new_n3247_), .A2(new_n9503_), .ZN(new_n10822_));
  NAND4_X1   g10758(.A1(new_n3758_), .A2(new_n6922_), .A3(new_n10821_), .A4(new_n10822_), .ZN(new_n10823_));
  XOR2_X1    g10759(.A1(new_n10823_), .A2(\a[2] ), .Z(new_n10824_));
  OAI21_X1   g10760(.A1(new_n10820_), .A2(new_n9516_), .B(new_n10824_), .ZN(new_n10825_));
  NOR2_X1    g10761(.A1(new_n9455_), .A2(new_n9480_), .ZN(new_n10826_));
  NOR2_X1    g10762(.A1(new_n9424_), .A2(new_n9481_), .ZN(new_n10827_));
  OAI21_X1   g10763(.A1(new_n10826_), .A2(new_n10827_), .B(new_n10816_), .ZN(new_n10828_));
  INV_X1     g10764(.I(new_n10824_), .ZN(new_n10829_));
  NAND3_X1   g10765(.A1(new_n10828_), .A2(new_n9527_), .A3(new_n10829_), .ZN(new_n10830_));
  NAND2_X1   g10766(.A1(new_n10825_), .A2(new_n10830_), .ZN(new_n10831_));
  NAND3_X1   g10767(.A1(new_n10812_), .A2(new_n10815_), .A3(new_n10831_), .ZN(new_n10832_));
  AOI21_X1   g10768(.A1(new_n10813_), .A2(new_n10814_), .B(new_n9471_), .ZN(new_n10833_));
  NOR3_X1    g10769(.A1(new_n10811_), .A2(new_n10808_), .A3(new_n10803_), .ZN(new_n10834_));
  AOI21_X1   g10770(.A1(new_n10828_), .A2(new_n9527_), .B(new_n10829_), .ZN(new_n10835_));
  NOR3_X1    g10771(.A1(new_n10820_), .A2(new_n9516_), .A3(new_n10824_), .ZN(new_n10836_));
  NOR2_X1    g10772(.A1(new_n10835_), .A2(new_n10836_), .ZN(new_n10837_));
  OAI21_X1   g10773(.A1(new_n10834_), .A2(new_n10833_), .B(new_n10837_), .ZN(new_n10838_));
  NAND2_X1   g10774(.A1(new_n10838_), .A2(new_n10832_), .ZN(new_n10839_));
  AOI21_X1   g10775(.A1(new_n10802_), .A2(new_n9529_), .B(new_n10839_), .ZN(new_n10840_));
  NOR2_X1    g10776(.A1(new_n10840_), .A2(new_n10795_), .ZN(new_n10841_));
  NOR3_X1    g10777(.A1(new_n10834_), .A2(new_n10833_), .A3(new_n10837_), .ZN(new_n10842_));
  AOI21_X1   g10778(.A1(new_n10812_), .A2(new_n10815_), .B(new_n10831_), .ZN(new_n10843_));
  NOR2_X1    g10779(.A1(new_n10842_), .A2(new_n10843_), .ZN(new_n10844_));
  NOR2_X1    g10780(.A1(new_n8797_), .A2(new_n9474_), .ZN(new_n10845_));
  NOR2_X1    g10781(.A1(new_n10845_), .A2(new_n9476_), .ZN(new_n10846_));
  OAI21_X1   g10782(.A1(new_n9478_), .A2(new_n10844_), .B(new_n10846_), .ZN(new_n10847_));
  AOI21_X1   g10783(.A1(new_n9478_), .A2(new_n10844_), .B(new_n10846_), .ZN(new_n10848_));
  AOI21_X1   g10784(.A1(new_n10841_), .A2(new_n10847_), .B(new_n10848_), .ZN(new_n10849_));
  NOR2_X1    g10785(.A1(new_n10849_), .A2(new_n9479_), .ZN(new_n10850_));
  AOI21_X1   g10786(.A1(new_n7922_), .A2(new_n7923_), .B(new_n6948_), .ZN(new_n10851_));
  NOR3_X1    g10787(.A1(new_n7141_), .A2(new_n7140_), .A3(new_n6853_), .ZN(new_n10852_));
  NOR2_X1    g10788(.A1(new_n10851_), .A2(new_n10852_), .ZN(new_n10853_));
  INV_X1     g10789(.I(new_n10853_), .ZN(new_n10854_));
  AOI21_X1   g10790(.A1(new_n10849_), .A2(new_n9479_), .B(new_n10854_), .ZN(new_n10855_));
  NOR2_X1    g10791(.A1(new_n10855_), .A2(new_n10850_), .ZN(new_n10856_));
  OAI21_X1   g10792(.A1(new_n7372_), .A2(new_n7368_), .B(new_n7374_), .ZN(new_n10857_));
  NAND3_X1   g10793(.A1(new_n7925_), .A2(new_n7926_), .A3(new_n7375_), .ZN(new_n10858_));
  AOI21_X1   g10794(.A1(new_n10857_), .A2(new_n10858_), .B(new_n7142_), .ZN(new_n10859_));
  AOI21_X1   g10795(.A1(new_n7927_), .A2(new_n7377_), .B(new_n7924_), .ZN(new_n10860_));
  NOR2_X1    g10796(.A1(new_n10860_), .A2(new_n10859_), .ZN(new_n10861_));
  INV_X1     g10797(.I(new_n10861_), .ZN(new_n10862_));
  OAI21_X1   g10798(.A1(new_n8784_), .A2(new_n10853_), .B(new_n10861_), .ZN(new_n10863_));
  NAND2_X1   g10799(.A1(new_n8784_), .A2(new_n10853_), .ZN(new_n10864_));
  AOI22_X1   g10800(.A1(new_n10856_), .A2(new_n10863_), .B1(new_n10862_), .B2(new_n10864_), .ZN(new_n10865_));
  AOI21_X1   g10801(.A1(new_n10865_), .A2(new_n8785_), .B(new_n8779_), .ZN(new_n10866_));
  XOR2_X1    g10802(.A1(new_n7790_), .A2(new_n7915_), .Z(new_n10867_));
  NOR2_X1    g10803(.A1(new_n10867_), .A2(new_n7948_), .ZN(new_n10868_));
  XOR2_X1    g10804(.A1(new_n7790_), .A2(new_n7914_), .Z(new_n10869_));
  NOR2_X1    g10805(.A1(new_n10869_), .A2(new_n7655_), .ZN(new_n10870_));
  NOR2_X1    g10806(.A1(new_n10868_), .A2(new_n10870_), .ZN(new_n10871_));
  INV_X1     g10807(.I(new_n10871_), .ZN(new_n10872_));
  NAND2_X1   g10808(.A1(new_n10856_), .A2(new_n10863_), .ZN(new_n10873_));
  NAND2_X1   g10809(.A1(new_n10864_), .A2(new_n10862_), .ZN(new_n10874_));
  NAND2_X1   g10810(.A1(new_n10873_), .A2(new_n10874_), .ZN(new_n10875_));
  AOI21_X1   g10811(.A1(new_n10875_), .A2(new_n8784_), .B(new_n8778_), .ZN(new_n10876_));
  NOR2_X1    g10812(.A1(new_n10876_), .A2(new_n10872_), .ZN(new_n10877_));
  NOR2_X1    g10813(.A1(new_n7950_), .A2(new_n7949_), .ZN(new_n10878_));
  NAND2_X1   g10814(.A1(new_n7655_), .A2(new_n7791_), .ZN(new_n10879_));
  XOR2_X1    g10815(.A1(new_n10879_), .A2(new_n10878_), .Z(new_n10880_));
  XOR2_X1    g10816(.A1(new_n7655_), .A2(new_n7791_), .Z(new_n10881_));
  NAND2_X1   g10817(.A1(new_n10881_), .A2(new_n7915_), .ZN(new_n10882_));
  NOR2_X1    g10818(.A1(new_n10880_), .A2(new_n10882_), .ZN(new_n10883_));
  AND2_X2    g10819(.A1(new_n10880_), .A2(new_n10882_), .Z(new_n10884_));
  NOR2_X1    g10820(.A1(new_n10884_), .A2(new_n10883_), .ZN(new_n10885_));
  INV_X1     g10821(.I(new_n10885_), .ZN(new_n10886_));
  OAI21_X1   g10822(.A1(new_n8182_), .A2(new_n8181_), .B(new_n8039_), .ZN(new_n10887_));
  NAND3_X1   g10823(.A1(new_n8030_), .A2(new_n8035_), .A3(new_n8040_), .ZN(new_n10888_));
  NAND2_X1   g10824(.A1(new_n10887_), .A2(new_n10888_), .ZN(new_n10889_));
  AOI21_X1   g10825(.A1(new_n10872_), .A2(new_n10889_), .B(new_n10886_), .ZN(new_n10890_));
  OR3_X2     g10826(.A1(new_n10877_), .A2(new_n10866_), .A3(new_n10890_), .Z(new_n10891_));
  INV_X1     g10827(.I(new_n10889_), .ZN(new_n10892_));
  AOI21_X1   g10828(.A1(new_n10892_), .A2(new_n10871_), .B(new_n10885_), .ZN(new_n10893_));
  INV_X1     g10829(.I(new_n10893_), .ZN(new_n10894_));
  XOR2_X1    g10830(.A1(new_n8108_), .A2(new_n8174_), .Z(new_n10895_));
  NOR2_X1    g10831(.A1(new_n10895_), .A2(new_n8183_), .ZN(new_n10896_));
  XOR2_X1    g10832(.A1(new_n8108_), .A2(new_n8186_), .Z(new_n10897_));
  NOR2_X1    g10833(.A1(new_n10897_), .A2(new_n8041_), .ZN(new_n10898_));
  NOR2_X1    g10834(.A1(new_n10898_), .A2(new_n10896_), .ZN(new_n10899_));
  OAI21_X1   g10835(.A1(new_n8774_), .A2(new_n10892_), .B(new_n10899_), .ZN(new_n10900_));
  NAND3_X1   g10836(.A1(new_n10891_), .A2(new_n10894_), .A3(new_n10900_), .ZN(new_n10901_));
  AOI21_X1   g10837(.A1(new_n8774_), .A2(new_n10892_), .B(new_n10899_), .ZN(new_n10902_));
  INV_X1     g10838(.I(new_n10902_), .ZN(new_n10903_));
  NAND2_X1   g10839(.A1(new_n10901_), .A2(new_n10903_), .ZN(new_n10904_));
  OAI21_X1   g10840(.A1(new_n10904_), .A2(new_n8774_), .B(new_n8766_), .ZN(new_n10905_));
  INV_X1     g10841(.I(new_n8774_), .ZN(new_n10906_));
  AOI21_X1   g10842(.A1(new_n10901_), .A2(new_n10903_), .B(new_n10906_), .ZN(new_n10907_));
  OAI21_X1   g10843(.A1(new_n10875_), .A2(new_n8784_), .B(new_n8778_), .ZN(new_n10908_));
  OAI21_X1   g10844(.A1(new_n10872_), .A2(new_n10876_), .B(new_n10908_), .ZN(new_n10909_));
  NOR2_X1    g10845(.A1(new_n10909_), .A2(new_n10890_), .ZN(new_n10910_));
  INV_X1     g10846(.I(new_n10900_), .ZN(new_n10911_));
  NOR3_X1    g10847(.A1(new_n10911_), .A2(new_n10910_), .A3(new_n10893_), .ZN(new_n10912_));
  NOR3_X1    g10848(.A1(new_n10912_), .A2(new_n8774_), .A3(new_n10902_), .ZN(new_n10913_));
  OAI21_X1   g10849(.A1(new_n10907_), .A2(new_n8766_), .B(new_n8758_), .ZN(new_n10914_));
  AOI22_X1   g10850(.A1(new_n10914_), .A2(new_n10905_), .B1(new_n8746_), .B2(new_n8761_), .ZN(new_n10915_));
  NOR2_X1    g10851(.A1(new_n10915_), .A2(new_n8760_), .ZN(new_n10916_));
  NOR2_X1    g10852(.A1(new_n8751_), .A2(new_n8745_), .ZN(new_n10917_));
  NOR2_X1    g10853(.A1(new_n10916_), .A2(new_n10917_), .ZN(new_n10918_));
  NOR2_X1    g10854(.A1(new_n10918_), .A2(new_n8753_), .ZN(new_n10919_));
  XOR2_X1    g10855(.A1(new_n8274_), .A2(new_n8283_), .Z(new_n10920_));
  NOR2_X1    g10856(.A1(new_n8261_), .A2(new_n10920_), .ZN(new_n10921_));
  XNOR2_X1   g10857(.A1(new_n8274_), .A2(new_n8283_), .ZN(new_n10922_));
  NOR2_X1    g10858(.A1(new_n8469_), .A2(new_n10922_), .ZN(new_n10923_));
  NOR2_X1    g10859(.A1(new_n10923_), .A2(new_n10921_), .ZN(new_n10924_));
  OAI21_X1   g10860(.A1(new_n8735_), .A2(new_n8751_), .B(new_n10924_), .ZN(new_n10925_));
  NAND2_X1   g10861(.A1(new_n10919_), .A2(new_n10925_), .ZN(new_n10926_));
  INV_X1     g10862(.I(new_n10924_), .ZN(new_n10927_));
  OAI21_X1   g10863(.A1(new_n8736_), .A2(new_n8752_), .B(new_n10927_), .ZN(new_n10928_));
  NOR2_X1    g10864(.A1(new_n8725_), .A2(new_n8735_), .ZN(new_n10929_));
  AOI21_X1   g10865(.A1(new_n10926_), .A2(new_n10928_), .B(new_n10929_), .ZN(new_n10930_));
  NOR2_X1    g10866(.A1(new_n8725_), .A2(new_n8718_), .ZN(new_n10931_));
  INV_X1     g10867(.I(new_n10931_), .ZN(new_n10932_));
  OAI21_X1   g10868(.A1(new_n10930_), .A2(new_n8737_), .B(new_n10932_), .ZN(new_n10933_));
  NAND2_X1   g10869(.A1(new_n10933_), .A2(new_n8728_), .ZN(new_n10934_));
  NAND2_X1   g10870(.A1(new_n8711_), .A2(new_n8719_), .ZN(new_n10935_));
  AOI21_X1   g10871(.A1(new_n10934_), .A2(new_n10935_), .B(new_n8720_), .ZN(new_n10936_));
  NOR2_X1    g10872(.A1(new_n8701_), .A2(new_n8710_), .ZN(new_n10937_));
  OAI21_X1   g10873(.A1(new_n10936_), .A2(new_n10937_), .B(new_n8713_), .ZN(new_n10938_));
  NOR2_X1    g10874(.A1(new_n8701_), .A2(new_n8694_), .ZN(new_n10939_));
  INV_X1     g10875(.I(new_n10939_), .ZN(new_n10940_));
  AOI21_X1   g10876(.A1(new_n10938_), .A2(new_n10940_), .B(new_n8703_), .ZN(new_n10941_));
  NOR2_X1    g10877(.A1(new_n8681_), .A2(new_n8694_), .ZN(new_n10942_));
  OAI21_X1   g10878(.A1(new_n10941_), .A2(new_n10942_), .B(new_n8695_), .ZN(new_n10943_));
  NOR2_X1    g10879(.A1(new_n8681_), .A2(new_n8687_), .ZN(new_n10944_));
  INV_X1     g10880(.I(new_n10944_), .ZN(new_n10945_));
  AOI21_X1   g10881(.A1(new_n10943_), .A2(new_n10945_), .B(new_n8689_), .ZN(new_n10946_));
  NOR2_X1    g10882(.A1(new_n10946_), .A2(new_n8674_), .ZN(new_n10947_));
  AOI22_X1   g10883(.A1(new_n10933_), .A2(new_n8728_), .B1(new_n8711_), .B2(new_n8719_), .ZN(new_n10948_));
  INV_X1     g10884(.I(new_n10937_), .ZN(new_n10949_));
  OAI21_X1   g10885(.A1(new_n10948_), .A2(new_n8720_), .B(new_n10949_), .ZN(new_n10950_));
  AOI21_X1   g10886(.A1(new_n10950_), .A2(new_n8713_), .B(new_n10939_), .ZN(new_n10951_));
  INV_X1     g10887(.I(new_n10942_), .ZN(new_n10952_));
  OAI21_X1   g10888(.A1(new_n10951_), .A2(new_n8703_), .B(new_n10952_), .ZN(new_n10953_));
  AOI21_X1   g10889(.A1(new_n10953_), .A2(new_n8695_), .B(new_n10944_), .ZN(new_n10954_));
  NOR3_X1    g10890(.A1(new_n10954_), .A2(new_n8673_), .A3(new_n8689_), .ZN(new_n10955_));
  XNOR2_X1   g10891(.A1(new_n8673_), .A2(new_n8687_), .ZN(new_n10956_));
  NOR4_X1    g10892(.A1(new_n10947_), .A2(new_n8662_), .A3(new_n10955_), .A4(new_n10956_), .ZN(new_n10957_));
  INV_X1     g10893(.I(new_n10947_), .ZN(new_n10958_));
  NOR2_X1    g10894(.A1(new_n10955_), .A2(new_n10956_), .ZN(new_n10959_));
  AOI21_X1   g10895(.A1(new_n10958_), .A2(new_n10959_), .B(new_n8661_), .ZN(new_n10960_));
  AOI21_X1   g10896(.A1(new_n8688_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n10961_));
  OAI21_X1   g10897(.A1(new_n2767_), .A2(new_n8673_), .B(new_n10961_), .ZN(new_n10962_));
  AOI21_X1   g10898(.A1(new_n8662_), .A2(new_n3332_), .B(new_n10962_), .ZN(new_n10963_));
  OAI21_X1   g10899(.A1(new_n10960_), .A2(new_n10957_), .B(new_n10963_), .ZN(new_n10964_));
  NOR2_X1    g10900(.A1(new_n10964_), .A2(new_n341_), .ZN(new_n10965_));
  INV_X1     g10901(.I(new_n10965_), .ZN(new_n10966_));
  NOR4_X1    g10902(.A1(new_n1976_), .A2(new_n1784_), .A3(new_n81_), .A4(new_n267_), .ZN(new_n10967_));
  NAND4_X1   g10903(.A1(new_n1404_), .A2(new_n113_), .A3(new_n1190_), .A4(new_n840_), .ZN(new_n10968_));
  NAND3_X1   g10904(.A1(new_n10967_), .A2(new_n6523_), .A3(new_n10968_), .ZN(new_n10969_));
  NOR2_X1    g10905(.A1(new_n4749_), .A2(new_n468_), .ZN(new_n10970_));
  NOR3_X1    g10906(.A1(new_n944_), .A2(new_n149_), .A3(new_n152_), .ZN(new_n10971_));
  NAND4_X1   g10907(.A1(new_n10970_), .A2(new_n807_), .A3(new_n1628_), .A4(new_n10971_), .ZN(new_n10972_));
  NAND4_X1   g10908(.A1(new_n685_), .A2(new_n385_), .A3(new_n1647_), .A4(new_n665_), .ZN(new_n10973_));
  NAND4_X1   g10909(.A1(new_n10973_), .A2(new_n872_), .A3(new_n1444_), .A4(new_n1572_), .ZN(new_n10974_));
  OR4_X2     g10910(.A1(new_n3836_), .A2(new_n10969_), .A3(new_n10972_), .A4(new_n10974_), .Z(new_n10975_));
  NAND4_X1   g10911(.A1(new_n797_), .A2(new_n842_), .A3(new_n301_), .A4(new_n1067_), .ZN(new_n10976_));
  NOR4_X1    g10912(.A1(new_n147_), .A2(new_n154_), .A3(new_n294_), .A4(new_n574_), .ZN(new_n10977_));
  NAND4_X1   g10913(.A1(new_n442_), .A2(new_n1129_), .A3(new_n508_), .A4(new_n187_), .ZN(new_n10978_));
  NAND4_X1   g10914(.A1(new_n1026_), .A2(new_n349_), .A3(new_n391_), .A4(new_n405_), .ZN(new_n10979_));
  NAND2_X1   g10915(.A1(new_n10979_), .A2(new_n10978_), .ZN(new_n10980_));
  NOR4_X1    g10916(.A1(new_n10980_), .A2(new_n712_), .A3(new_n1213_), .A4(new_n1276_), .ZN(new_n10981_));
  NAND4_X1   g10917(.A1(new_n10981_), .A2(new_n3493_), .A3(new_n10976_), .A4(new_n10977_), .ZN(new_n10982_));
  NAND3_X1   g10918(.A1(new_n2332_), .A2(new_n362_), .A3(new_n509_), .ZN(new_n10983_));
  NOR2_X1    g10919(.A1(new_n869_), .A2(new_n2839_), .ZN(new_n10984_));
  NAND4_X1   g10920(.A1(new_n2119_), .A2(new_n598_), .A3(new_n414_), .A4(new_n999_), .ZN(new_n10985_));
  NAND4_X1   g10921(.A1(new_n10984_), .A2(new_n3506_), .A3(new_n10983_), .A4(new_n10985_), .ZN(new_n10986_));
  NOR3_X1    g10922(.A1(new_n119_), .A2(new_n403_), .A3(new_n226_), .ZN(new_n10987_));
  NAND4_X1   g10923(.A1(new_n1329_), .A2(new_n1590_), .A3(new_n829_), .A4(new_n10987_), .ZN(new_n10988_));
  NOR4_X1    g10924(.A1(new_n10982_), .A2(new_n10975_), .A3(new_n10986_), .A4(new_n10988_), .ZN(new_n10989_));
  NAND2_X1   g10925(.A1(new_n10989_), .A2(new_n4573_), .ZN(new_n10990_));
  NOR4_X1    g10926(.A1(new_n1247_), .A2(new_n3856_), .A3(new_n906_), .A4(new_n459_), .ZN(new_n10991_));
  NAND2_X1   g10927(.A1(new_n220_), .A2(new_n188_), .ZN(new_n10992_));
  NAND2_X1   g10928(.A1(new_n438_), .A2(new_n1058_), .ZN(new_n10993_));
  NOR4_X1    g10929(.A1(new_n891_), .A2(new_n10993_), .A3(new_n835_), .A4(new_n873_), .ZN(new_n10994_));
  INV_X1     g10930(.I(new_n10994_), .ZN(new_n10995_));
  NOR4_X1    g10931(.A1(new_n10995_), .A2(new_n866_), .A3(new_n1313_), .A4(new_n10992_), .ZN(new_n10996_));
  NAND4_X1   g10932(.A1(new_n10996_), .A2(new_n645_), .A3(new_n1901_), .A4(new_n10991_), .ZN(new_n10997_));
  NOR2_X1    g10933(.A1(new_n932_), .A2(new_n1079_), .ZN(new_n10998_));
  NOR2_X1    g10934(.A1(new_n289_), .A2(new_n553_), .ZN(new_n10999_));
  NAND2_X1   g10935(.A1(new_n10999_), .A2(new_n410_), .ZN(new_n11000_));
  NOR4_X1    g10936(.A1(new_n11000_), .A2(new_n2982_), .A3(new_n463_), .A4(new_n732_), .ZN(new_n11001_));
  NOR4_X1    g10937(.A1(new_n2439_), .A2(new_n590_), .A3(new_n721_), .A4(new_n216_), .ZN(new_n11002_));
  NOR2_X1    g10938(.A1(new_n2955_), .A2(new_n11002_), .ZN(new_n11003_));
  NAND4_X1   g10939(.A1(new_n11003_), .A2(new_n2479_), .A3(new_n11001_), .A4(new_n10998_), .ZN(new_n11004_));
  NOR4_X1    g10940(.A1(new_n10997_), .A2(new_n1983_), .A3(new_n2417_), .A4(new_n11004_), .ZN(new_n11005_));
  NAND2_X1   g10941(.A1(new_n11005_), .A2(new_n2273_), .ZN(new_n11006_));
  NOR2_X1    g10942(.A1(new_n11006_), .A2(new_n10990_), .ZN(new_n11007_));
  AOI22_X1   g10943(.A1(new_n3253_), .A2(new_n2764_), .B1(new_n2770_), .B2(new_n3247_), .ZN(new_n11008_));
  INV_X1     g10944(.I(new_n3152_), .ZN(new_n11009_));
  NOR4_X1    g10945(.A1(new_n2034_), .A2(new_n782_), .A3(new_n1073_), .A4(new_n1962_), .ZN(new_n11010_));
  NAND4_X1   g10946(.A1(new_n3125_), .A2(new_n11010_), .A3(new_n1767_), .A4(new_n2634_), .ZN(new_n11011_));
  NOR2_X1    g10947(.A1(new_n1175_), .A2(new_n930_), .ZN(new_n11012_));
  AOI21_X1   g10948(.A1(new_n1246_), .A2(new_n11012_), .B(new_n2234_), .ZN(new_n11013_));
  NAND3_X1   g10949(.A1(new_n380_), .A2(new_n2697_), .A3(new_n11013_), .ZN(new_n11014_));
  NOR4_X1    g10950(.A1(new_n11009_), .A2(new_n11014_), .A3(new_n3954_), .A4(new_n11011_), .ZN(new_n11015_));
  NAND2_X1   g10951(.A1(new_n11015_), .A2(new_n2686_), .ZN(new_n11016_));
  NOR4_X1    g10952(.A1(new_n2438_), .A2(new_n347_), .A3(new_n945_), .A4(new_n763_), .ZN(new_n11017_));
  NAND3_X1   g10953(.A1(new_n11017_), .A2(new_n344_), .A3(new_n949_), .ZN(new_n11018_));
  INV_X1     g10954(.I(new_n11018_), .ZN(new_n11019_));
  NOR3_X1    g10955(.A1(new_n681_), .A2(new_n1168_), .A3(new_n749_), .ZN(new_n11020_));
  INV_X1     g10956(.I(new_n11020_), .ZN(new_n11021_));
  NOR4_X1    g10957(.A1(new_n2650_), .A2(new_n3137_), .A3(new_n1589_), .A4(new_n11021_), .ZN(new_n11022_));
  NAND4_X1   g10958(.A1(new_n3154_), .A2(new_n3128_), .A3(new_n11019_), .A4(new_n11022_), .ZN(new_n11023_));
  INV_X1     g10959(.I(new_n11023_), .ZN(new_n11024_));
  NOR2_X1    g10960(.A1(new_n11024_), .A2(new_n11016_), .ZN(new_n11025_));
  INV_X1     g10961(.I(new_n11016_), .ZN(new_n11026_));
  NOR2_X1    g10962(.A1(new_n11026_), .A2(new_n11023_), .ZN(new_n11027_));
  INV_X1     g10963(.I(new_n11027_), .ZN(new_n11028_));
  OAI21_X1   g10964(.A1(new_n11008_), .A2(new_n11025_), .B(new_n11028_), .ZN(new_n11029_));
  NOR3_X1    g10965(.A1(new_n379_), .A2(new_n647_), .A3(new_n1011_), .ZN(new_n11030_));
  INV_X1     g10966(.I(new_n11030_), .ZN(new_n11031_));
  NOR2_X1    g10967(.A1(new_n582_), .A2(new_n1035_), .ZN(new_n11032_));
  NAND4_X1   g10968(.A1(new_n11032_), .A2(new_n3022_), .A3(new_n551_), .A4(new_n832_), .ZN(new_n11033_));
  NOR4_X1    g10969(.A1(new_n2699_), .A2(new_n3163_), .A3(new_n11031_), .A4(new_n11033_), .ZN(new_n11034_));
  XOR2_X1    g10970(.A1(new_n11034_), .A2(new_n11016_), .Z(new_n11035_));
  INV_X1     g10971(.I(new_n11035_), .ZN(new_n11036_));
  NOR2_X1    g10972(.A1(new_n11029_), .A2(new_n11036_), .ZN(new_n11037_));
  INV_X1     g10973(.I(new_n11037_), .ZN(new_n11038_));
  AOI22_X1   g10974(.A1(new_n3168_), .A2(new_n2770_), .B1(new_n3189_), .B2(new_n3247_), .ZN(new_n11039_));
  AOI21_X1   g10975(.A1(new_n3758_), .A2(new_n2764_), .B(new_n11039_), .ZN(new_n11040_));
  NAND4_X1   g10976(.A1(new_n2642_), .A2(new_n502_), .A3(new_n2458_), .A4(new_n3868_), .ZN(new_n11041_));
  INV_X1     g10977(.I(new_n11041_), .ZN(new_n11042_));
  NAND2_X1   g10978(.A1(new_n2697_), .A2(new_n11013_), .ZN(new_n11043_));
  NOR2_X1    g10979(.A1(new_n684_), .A2(new_n125_), .ZN(new_n11044_));
  INV_X1     g10980(.I(new_n2294_), .ZN(new_n11045_));
  NOR4_X1    g10981(.A1(new_n11045_), .A2(new_n1276_), .A3(new_n1341_), .A4(new_n2445_), .ZN(new_n11046_));
  NAND4_X1   g10982(.A1(new_n11046_), .A2(new_n2656_), .A3(new_n665_), .A4(new_n11044_), .ZN(new_n11047_));
  NOR4_X1    g10983(.A1(new_n11043_), .A2(new_n2672_), .A3(new_n11047_), .A4(new_n11018_), .ZN(new_n11048_));
  NAND2_X1   g10984(.A1(new_n11042_), .A2(new_n11048_), .ZN(new_n11049_));
  NOR4_X1    g10985(.A1(new_n4886_), .A2(new_n647_), .A3(new_n1247_), .A4(new_n1864_), .ZN(new_n11050_));
  NOR3_X1    g10986(.A1(new_n3419_), .A2(new_n191_), .A3(new_n1381_), .ZN(new_n11051_));
  AND3_X2    g10987(.A1(new_n2292_), .A2(new_n11051_), .A3(new_n11050_), .Z(new_n11052_));
  NAND3_X1   g10988(.A1(new_n720_), .A2(new_n540_), .A3(new_n685_), .ZN(new_n11053_));
  NOR4_X1    g10989(.A1(new_n11053_), .A2(new_n163_), .A3(new_n1984_), .A4(new_n3412_), .ZN(new_n11054_));
  NAND4_X1   g10990(.A1(new_n408_), .A2(new_n966_), .A3(new_n1322_), .A4(new_n1096_), .ZN(new_n11055_));
  NOR3_X1    g10991(.A1(new_n241_), .A2(new_n381_), .A3(new_n791_), .ZN(new_n11056_));
  NAND3_X1   g10992(.A1(new_n11054_), .A2(new_n11055_), .A3(new_n11056_), .ZN(new_n11057_));
  NAND4_X1   g10993(.A1(new_n220_), .A2(new_n287_), .A3(new_n1396_), .A4(new_n1095_), .ZN(new_n11058_));
  NAND4_X1   g10994(.A1(new_n965_), .A2(new_n797_), .A3(new_n1759_), .A4(new_n309_), .ZN(new_n11059_));
  NAND4_X1   g10995(.A1(new_n3877_), .A2(new_n2382_), .A3(new_n11058_), .A4(new_n11059_), .ZN(new_n11060_));
  NOR3_X1    g10996(.A1(new_n11057_), .A2(new_n11060_), .A3(new_n1041_), .ZN(new_n11061_));
  NOR4_X1    g10997(.A1(new_n960_), .A2(new_n70_), .A3(new_n81_), .A4(new_n630_), .ZN(new_n11062_));
  INV_X1     g10998(.I(new_n11062_), .ZN(new_n11063_));
  NOR4_X1    g10999(.A1(new_n252_), .A2(new_n437_), .A3(new_n596_), .A4(new_n475_), .ZN(new_n11064_));
  NOR4_X1    g11000(.A1(new_n495_), .A2(new_n239_), .A3(new_n376_), .A4(new_n731_), .ZN(new_n11065_));
  NOR4_X1    g11001(.A1(new_n11063_), .A2(new_n3156_), .A3(new_n11064_), .A4(new_n11065_), .ZN(new_n11066_));
  NAND4_X1   g11002(.A1(new_n11066_), .A2(new_n221_), .A3(new_n2178_), .A4(new_n1647_), .ZN(new_n11067_));
  NOR2_X1    g11003(.A1(new_n11067_), .A2(new_n1709_), .ZN(new_n11068_));
  NAND3_X1   g11004(.A1(new_n11068_), .A2(new_n11052_), .A3(new_n11061_), .ZN(new_n11069_));
  INV_X1     g11005(.I(new_n11069_), .ZN(new_n11070_));
  NOR2_X1    g11006(.A1(new_n11070_), .A2(\a[29] ), .ZN(new_n11071_));
  NOR2_X1    g11007(.A1(new_n11069_), .A2(new_n74_), .ZN(new_n11072_));
  INV_X1     g11008(.I(new_n11072_), .ZN(new_n11073_));
  OAI21_X1   g11009(.A1(new_n11049_), .A2(new_n11071_), .B(new_n11073_), .ZN(new_n11074_));
  NOR2_X1    g11010(.A1(new_n11074_), .A2(new_n11016_), .ZN(new_n11075_));
  INV_X1     g11011(.I(new_n11075_), .ZN(new_n11076_));
  NAND2_X1   g11012(.A1(new_n11074_), .A2(new_n11016_), .ZN(new_n11077_));
  NAND2_X1   g11013(.A1(new_n11076_), .A2(new_n11077_), .ZN(new_n11078_));
  XOR2_X1    g11014(.A1(new_n11074_), .A2(new_n11026_), .Z(new_n11079_));
  NOR2_X1    g11015(.A1(new_n11040_), .A2(new_n11079_), .ZN(new_n11080_));
  AOI21_X1   g11016(.A1(new_n11040_), .A2(new_n11078_), .B(new_n11080_), .ZN(new_n11081_));
  INV_X1     g11017(.I(new_n11081_), .ZN(new_n11082_));
  NOR2_X1    g11018(.A1(new_n2614_), .A2(new_n2771_), .ZN(new_n11083_));
  NOR2_X1    g11019(.A1(new_n2716_), .A2(new_n2772_), .ZN(new_n11084_));
  NOR2_X1    g11020(.A1(new_n2665_), .A2(new_n2767_), .ZN(new_n11085_));
  NOR4_X1    g11021(.A1(new_n11084_), .A2(new_n2763_), .A3(new_n11083_), .A4(new_n11085_), .ZN(new_n11086_));
  INV_X1     g11022(.I(new_n800_), .ZN(new_n11087_));
  INV_X1     g11023(.I(new_n3983_), .ZN(new_n11088_));
  NOR4_X1    g11024(.A1(new_n203_), .A2(new_n1531_), .A3(new_n396_), .A4(new_n149_), .ZN(new_n11089_));
  NOR4_X1    g11025(.A1(new_n262_), .A2(new_n603_), .A3(new_n330_), .A4(new_n347_), .ZN(new_n11090_));
  NOR3_X1    g11026(.A1(new_n11088_), .A2(new_n11089_), .A3(new_n11090_), .ZN(new_n11091_));
  NAND3_X1   g11027(.A1(new_n716_), .A2(new_n2283_), .A3(new_n1689_), .ZN(new_n11092_));
  NOR4_X1    g11028(.A1(new_n11092_), .A2(new_n1202_), .A3(new_n576_), .A4(new_n3353_), .ZN(new_n11093_));
  NAND2_X1   g11029(.A1(new_n11091_), .A2(new_n11093_), .ZN(new_n11094_));
  NAND4_X1   g11030(.A1(new_n1026_), .A2(new_n992_), .A3(new_n394_), .A4(new_n390_), .ZN(new_n11095_));
  NOR4_X1    g11031(.A1(new_n172_), .A2(new_n225_), .A3(new_n604_), .A4(new_n192_), .ZN(new_n11096_));
  NAND4_X1   g11032(.A1(new_n11096_), .A2(new_n572_), .A3(new_n222_), .A4(new_n1961_), .ZN(new_n11097_));
  NOR4_X1    g11033(.A1(new_n11097_), .A2(new_n104_), .A3(new_n687_), .A4(new_n1243_), .ZN(new_n11098_));
  NAND4_X1   g11034(.A1(new_n11098_), .A2(new_n2587_), .A3(new_n4844_), .A4(new_n11095_), .ZN(new_n11099_));
  NOR4_X1    g11035(.A1(new_n2982_), .A2(new_n4931_), .A3(new_n1323_), .A4(new_n2551_), .ZN(new_n11100_));
  NAND4_X1   g11036(.A1(new_n287_), .A2(new_n1706_), .A3(new_n464_), .A4(new_n1494_), .ZN(new_n11101_));
  NOR2_X1    g11037(.A1(new_n212_), .A2(new_n724_), .ZN(new_n11102_));
  NAND4_X1   g11038(.A1(new_n11100_), .A2(new_n832_), .A3(new_n11101_), .A4(new_n11102_), .ZN(new_n11103_));
  NOR4_X1    g11039(.A1(new_n11099_), .A2(new_n11087_), .A3(new_n11094_), .A4(new_n11103_), .ZN(new_n11104_));
  NAND2_X1   g11040(.A1(new_n11104_), .A2(new_n3415_), .ZN(new_n11105_));
  INV_X1     g11041(.I(new_n11105_), .ZN(new_n11106_));
  NOR2_X1    g11042(.A1(new_n3227_), .A2(new_n2808_), .ZN(new_n11107_));
  NOR2_X1    g11043(.A1(new_n11107_), .A2(new_n3229_), .ZN(new_n11108_));
  NAND2_X1   g11044(.A1(new_n11108_), .A2(new_n11106_), .ZN(new_n11109_));
  NAND3_X1   g11045(.A1(new_n2733_), .A2(new_n11086_), .A3(new_n11109_), .ZN(new_n11110_));
  OAI21_X1   g11046(.A1(new_n11107_), .A2(new_n3229_), .B(new_n11105_), .ZN(new_n11111_));
  NAND2_X1   g11047(.A1(new_n11110_), .A2(new_n11111_), .ZN(new_n11112_));
  NOR2_X1    g11048(.A1(new_n11106_), .A2(new_n11069_), .ZN(new_n11113_));
  INV_X1     g11049(.I(new_n11113_), .ZN(new_n11114_));
  NOR2_X1    g11050(.A1(new_n11070_), .A2(new_n11105_), .ZN(new_n11115_));
  AOI21_X1   g11051(.A1(new_n11112_), .A2(new_n11114_), .B(new_n11115_), .ZN(new_n11116_));
  INV_X1     g11052(.I(new_n11116_), .ZN(new_n11117_));
  NOR2_X1    g11053(.A1(new_n3176_), .A2(new_n2767_), .ZN(new_n11118_));
  NOR2_X1    g11054(.A1(new_n2716_), .A2(new_n2771_), .ZN(new_n11119_));
  NAND2_X1   g11055(.A1(new_n2762_), .A2(\a[31] ), .ZN(new_n11120_));
  NOR3_X1    g11056(.A1(new_n11118_), .A2(new_n11119_), .A3(new_n11120_), .ZN(new_n11121_));
  NAND2_X1   g11057(.A1(new_n3174_), .A2(new_n11121_), .ZN(new_n11122_));
  INV_X1     g11058(.I(new_n11122_), .ZN(new_n11123_));
  NOR2_X1    g11059(.A1(new_n11071_), .A2(new_n11072_), .ZN(new_n11124_));
  NOR2_X1    g11060(.A1(new_n11124_), .A2(new_n11049_), .ZN(new_n11125_));
  XOR2_X1    g11061(.A1(new_n11069_), .A2(\a[29] ), .Z(new_n11126_));
  INV_X1     g11062(.I(new_n11126_), .ZN(new_n11127_));
  AOI21_X1   g11063(.A1(new_n11049_), .A2(new_n11127_), .B(new_n11125_), .ZN(new_n11128_));
  INV_X1     g11064(.I(new_n11128_), .ZN(new_n11129_));
  NOR2_X1    g11065(.A1(new_n11123_), .A2(new_n11129_), .ZN(new_n11130_));
  INV_X1     g11066(.I(new_n11130_), .ZN(new_n11131_));
  NOR2_X1    g11067(.A1(new_n11122_), .A2(new_n11128_), .ZN(new_n11132_));
  AOI21_X1   g11068(.A1(new_n11131_), .A2(new_n11117_), .B(new_n11132_), .ZN(new_n11133_));
  NOR2_X1    g11069(.A1(new_n11133_), .A2(new_n11082_), .ZN(new_n11134_));
  OAI21_X1   g11070(.A1(new_n11113_), .A2(new_n11115_), .B(new_n11112_), .ZN(new_n11135_));
  XOR2_X1    g11071(.A1(new_n11069_), .A2(new_n11105_), .Z(new_n11136_));
  OAI21_X1   g11072(.A1(new_n11112_), .A2(new_n11136_), .B(new_n11135_), .ZN(new_n11137_));
  AOI21_X1   g11073(.A1(new_n2664_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n11138_));
  OAI21_X1   g11074(.A1(new_n2716_), .A2(new_n2767_), .B(new_n11138_), .ZN(new_n11139_));
  AOI21_X1   g11075(.A1(new_n3332_), .A2(new_n3168_), .B(new_n11139_), .ZN(new_n11140_));
  AND2_X2    g11076(.A1(new_n3273_), .A2(new_n11140_), .Z(new_n11141_));
  NOR2_X1    g11077(.A1(new_n11137_), .A2(new_n11141_), .ZN(new_n11142_));
  OAI22_X1   g11078(.A1(new_n3254_), .A2(new_n2737_), .B1(new_n2747_), .B2(new_n3142_), .ZN(new_n11143_));
  XOR2_X1    g11079(.A1(new_n11143_), .A2(new_n74_), .Z(new_n11144_));
  NOR2_X1    g11080(.A1(new_n11144_), .A2(new_n11142_), .ZN(new_n11145_));
  AOI21_X1   g11081(.A1(new_n11137_), .A2(new_n11141_), .B(new_n11145_), .ZN(new_n11146_));
  XOR2_X1    g11082(.A1(new_n11122_), .A2(new_n11129_), .Z(new_n11147_));
  OAI21_X1   g11083(.A1(new_n11130_), .A2(new_n11132_), .B(new_n11116_), .ZN(new_n11148_));
  OAI21_X1   g11084(.A1(new_n11116_), .A2(new_n11147_), .B(new_n11148_), .ZN(new_n11149_));
  XNOR2_X1   g11085(.A1(new_n11146_), .A2(new_n11149_), .ZN(new_n11150_));
  INV_X1     g11086(.I(new_n11150_), .ZN(new_n11151_));
  XOR2_X1    g11087(.A1(new_n11137_), .A2(new_n11143_), .Z(new_n11152_));
  XOR2_X1    g11088(.A1(new_n11152_), .A2(new_n74_), .Z(new_n11153_));
  XOR2_X1    g11089(.A1(new_n11153_), .A2(new_n11141_), .Z(new_n11154_));
  NAND2_X1   g11090(.A1(new_n2733_), .A2(new_n11086_), .ZN(new_n11155_));
  AOI21_X1   g11091(.A1(new_n11109_), .A2(new_n11111_), .B(new_n11155_), .ZN(new_n11156_));
  XOR2_X1    g11092(.A1(new_n11108_), .A2(new_n11105_), .Z(new_n11157_));
  AOI21_X1   g11093(.A1(new_n2733_), .A2(new_n11086_), .B(new_n11157_), .ZN(new_n11158_));
  NOR2_X1    g11094(.A1(new_n11156_), .A2(new_n11158_), .ZN(new_n11159_));
  NAND2_X1   g11095(.A1(new_n3168_), .A2(new_n2746_), .ZN(new_n11160_));
  NAND2_X1   g11096(.A1(new_n3247_), .A2(new_n3275_), .ZN(new_n11161_));
  NAND4_X1   g11097(.A1(new_n3758_), .A2(new_n2736_), .A3(new_n11160_), .A4(new_n11161_), .ZN(new_n11162_));
  XOR2_X1    g11098(.A1(new_n11162_), .A2(\a[29] ), .Z(new_n11163_));
  INV_X1     g11099(.I(new_n11163_), .ZN(new_n11164_));
  AOI21_X1   g11100(.A1(new_n3184_), .A2(new_n3234_), .B(new_n3236_), .ZN(new_n11165_));
  INV_X1     g11101(.I(new_n11165_), .ZN(new_n11166_));
  NOR2_X1    g11102(.A1(new_n11164_), .A2(new_n11166_), .ZN(new_n11167_));
  NOR2_X1    g11103(.A1(new_n11167_), .A2(new_n11159_), .ZN(new_n11168_));
  NOR2_X1    g11104(.A1(new_n11163_), .A2(new_n11165_), .ZN(new_n11169_));
  NOR2_X1    g11105(.A1(new_n11168_), .A2(new_n11169_), .ZN(new_n11170_));
  NAND2_X1   g11106(.A1(new_n11154_), .A2(new_n11170_), .ZN(new_n11171_));
  NOR2_X1    g11107(.A1(new_n11167_), .A2(new_n11169_), .ZN(new_n11172_));
  NOR2_X1    g11108(.A1(new_n11172_), .A2(new_n11159_), .ZN(new_n11173_));
  XOR2_X1    g11109(.A1(new_n11163_), .A2(new_n11166_), .Z(new_n11174_));
  INV_X1     g11110(.I(new_n11174_), .ZN(new_n11175_));
  AOI21_X1   g11111(.A1(new_n11159_), .A2(new_n11175_), .B(new_n11173_), .ZN(new_n11176_));
  INV_X1     g11112(.I(new_n11176_), .ZN(new_n11177_));
  INV_X1     g11113(.I(new_n3120_), .ZN(new_n11178_));
  AOI21_X1   g11114(.A1(new_n11178_), .A2(new_n3241_), .B(new_n3242_), .ZN(new_n11179_));
  NOR2_X1    g11115(.A1(new_n11177_), .A2(new_n11179_), .ZN(new_n11180_));
  INV_X1     g11116(.I(new_n11180_), .ZN(new_n11181_));
  NOR2_X1    g11117(.A1(new_n8669_), .A2(new_n3292_), .ZN(new_n11182_));
  OAI21_X1   g11118(.A1(new_n8655_), .A2(new_n8670_), .B(new_n11182_), .ZN(new_n11183_));
  XNOR2_X1   g11119(.A1(new_n11176_), .A2(new_n11179_), .ZN(new_n11184_));
  NOR2_X1    g11120(.A1(new_n11184_), .A2(new_n3289_), .ZN(new_n11185_));
  INV_X1     g11121(.I(new_n11185_), .ZN(new_n11186_));
  OAI21_X1   g11122(.A1(new_n11183_), .A2(new_n11186_), .B(new_n11181_), .ZN(new_n11187_));
  XNOR2_X1   g11123(.A1(new_n11154_), .A2(new_n11170_), .ZN(new_n11188_));
  OAI21_X1   g11124(.A1(new_n11187_), .A2(new_n11188_), .B(new_n11171_), .ZN(new_n11189_));
  XOR2_X1    g11125(.A1(new_n11133_), .A2(new_n11082_), .Z(new_n11190_));
  NAND2_X1   g11126(.A1(new_n11146_), .A2(new_n11149_), .ZN(new_n11191_));
  INV_X1     g11127(.I(new_n11191_), .ZN(new_n11192_));
  NOR2_X1    g11128(.A1(new_n11192_), .A2(new_n11190_), .ZN(new_n11193_));
  INV_X1     g11129(.I(new_n11193_), .ZN(new_n11194_));
  AOI21_X1   g11130(.A1(new_n11189_), .A2(new_n11151_), .B(new_n11194_), .ZN(new_n11195_));
  NOR2_X1    g11131(.A1(new_n11025_), .A2(new_n11027_), .ZN(new_n11196_));
  XNOR2_X1   g11132(.A1(new_n11023_), .A2(new_n11016_), .ZN(new_n11197_));
  NAND2_X1   g11133(.A1(new_n11008_), .A2(new_n11197_), .ZN(new_n11198_));
  OAI21_X1   g11134(.A1(new_n11008_), .A2(new_n11196_), .B(new_n11198_), .ZN(new_n11199_));
  NAND2_X1   g11135(.A1(new_n11040_), .A2(new_n11076_), .ZN(new_n11200_));
  NAND2_X1   g11136(.A1(new_n11200_), .A2(new_n11077_), .ZN(new_n11201_));
  NOR2_X1    g11137(.A1(new_n11199_), .A2(new_n11201_), .ZN(new_n11202_));
  INV_X1     g11138(.I(new_n11202_), .ZN(new_n11203_));
  OAI21_X1   g11139(.A1(new_n11195_), .A2(new_n11134_), .B(new_n11203_), .ZN(new_n11204_));
  XOR2_X1    g11140(.A1(new_n11029_), .A2(new_n11036_), .Z(new_n11205_));
  NAND2_X1   g11141(.A1(new_n11199_), .A2(new_n11201_), .ZN(new_n11206_));
  NAND2_X1   g11142(.A1(new_n11205_), .A2(new_n11206_), .ZN(new_n11207_));
  INV_X1     g11143(.I(new_n11207_), .ZN(new_n11208_));
  NAND2_X1   g11144(.A1(new_n11026_), .A2(new_n11034_), .ZN(new_n11209_));
  NOR4_X1    g11145(.A1(new_n420_), .A2(new_n611_), .A3(new_n684_), .A4(new_n660_), .ZN(new_n11210_));
  NAND2_X1   g11146(.A1(new_n2178_), .A2(new_n1935_), .ZN(new_n11211_));
  NOR4_X1    g11147(.A1(new_n3348_), .A2(new_n11211_), .A3(new_n11210_), .A4(new_n682_), .ZN(new_n11212_));
  AND4_X2    g11148(.A1(new_n747_), .A2(new_n11212_), .A3(new_n2553_), .A4(new_n2456_), .Z(new_n11213_));
  NOR3_X1    g11149(.A1(new_n2083_), .A2(new_n879_), .A3(new_n1323_), .ZN(new_n11214_));
  NOR3_X1    g11150(.A1(new_n1145_), .A2(new_n1262_), .A3(new_n474_), .ZN(new_n11215_));
  NOR2_X1    g11151(.A1(new_n1206_), .A2(new_n1365_), .ZN(new_n11216_));
  NAND4_X1   g11152(.A1(new_n11214_), .A2(new_n11215_), .A3(new_n11216_), .A4(new_n4799_), .ZN(new_n11217_));
  NOR2_X1    g11153(.A1(new_n2543_), .A2(new_n2171_), .ZN(new_n11218_));
  NAND2_X1   g11154(.A1(new_n11218_), .A2(new_n4826_), .ZN(new_n11219_));
  NOR3_X1    g11155(.A1(new_n11219_), .A2(new_n1450_), .A3(new_n11217_), .ZN(new_n11220_));
  NAND4_X1   g11156(.A1(new_n341_), .A2(new_n3098_), .A3(new_n11213_), .A4(new_n11220_), .ZN(new_n11221_));
  INV_X1     g11157(.I(new_n11221_), .ZN(new_n11222_));
  NOR2_X1    g11158(.A1(new_n1014_), .A2(new_n764_), .ZN(new_n11223_));
  NAND4_X1   g11159(.A1(new_n11222_), .A2(new_n635_), .A3(new_n3136_), .A4(new_n11223_), .ZN(new_n11224_));
  NAND2_X1   g11160(.A1(new_n11224_), .A2(new_n11209_), .ZN(new_n11225_));
  NAND4_X1   g11161(.A1(new_n11204_), .A2(new_n11038_), .A3(new_n11208_), .A4(new_n11225_), .ZN(new_n11226_));
  NAND2_X1   g11162(.A1(new_n4097_), .A2(new_n3775_), .ZN(new_n11227_));
  NOR3_X1    g11163(.A1(new_n11227_), .A2(new_n3770_), .A3(new_n3773_), .ZN(new_n11228_));
  NOR2_X1    g11164(.A1(new_n11228_), .A2(new_n3035_), .ZN(new_n11229_));
  INV_X1     g11165(.I(new_n11228_), .ZN(new_n11230_));
  NAND2_X1   g11166(.A1(new_n11226_), .A2(new_n11230_), .ZN(new_n11231_));
  AOI22_X1   g11167(.A1(new_n11231_), .A2(new_n3035_), .B1(new_n11226_), .B2(new_n11229_), .ZN(new_n11232_));
  NAND2_X1   g11168(.A1(new_n11006_), .A2(new_n10990_), .ZN(new_n11233_));
  AOI21_X1   g11169(.A1(new_n11232_), .A2(new_n11233_), .B(new_n11007_), .ZN(new_n11234_));
  NAND2_X1   g11170(.A1(new_n10964_), .A2(new_n341_), .ZN(new_n11235_));
  INV_X1     g11171(.I(new_n11235_), .ZN(new_n11236_));
  OAI21_X1   g11172(.A1(new_n11234_), .A2(new_n11236_), .B(new_n10966_), .ZN(new_n11237_));
  INV_X1     g11173(.I(new_n341_), .ZN(new_n11238_));
  NOR3_X1    g11174(.A1(new_n1264_), .A2(new_n1875_), .A3(new_n1630_), .ZN(new_n11239_));
  NOR4_X1    g11175(.A1(new_n2601_), .A2(new_n3203_), .A3(new_n130_), .A4(new_n136_), .ZN(new_n11240_));
  NOR4_X1    g11176(.A1(new_n1355_), .A2(new_n214_), .A3(new_n577_), .A4(new_n1138_), .ZN(new_n11241_));
  INV_X1     g11177(.I(new_n11241_), .ZN(new_n11242_));
  NAND4_X1   g11178(.A1(new_n11240_), .A2(new_n3090_), .A3(new_n11239_), .A4(new_n11242_), .ZN(new_n11243_));
  INV_X1     g11179(.I(new_n476_), .ZN(new_n11244_));
  NOR3_X1    g11180(.A1(new_n946_), .A2(new_n397_), .A3(new_n714_), .ZN(new_n11245_));
  NAND4_X1   g11181(.A1(new_n11245_), .A2(new_n1358_), .A3(new_n1314_), .A4(new_n351_), .ZN(new_n11246_));
  NOR4_X1    g11182(.A1(new_n11246_), .A2(new_n11244_), .A3(new_n2137_), .A4(new_n3855_), .ZN(new_n11247_));
  NAND4_X1   g11183(.A1(new_n11247_), .A2(new_n614_), .A3(new_n2850_), .A4(new_n4404_), .ZN(new_n11248_));
  NOR3_X1    g11184(.A1(new_n11248_), .A2(new_n10975_), .A3(new_n11243_), .ZN(new_n11249_));
  NAND2_X1   g11185(.A1(new_n11249_), .A2(new_n3491_), .ZN(new_n11250_));
  INV_X1     g11186(.I(new_n11250_), .ZN(new_n11251_));
  NOR2_X1    g11187(.A1(new_n11238_), .A2(new_n11251_), .ZN(new_n11252_));
  NOR2_X1    g11188(.A1(new_n341_), .A2(new_n11250_), .ZN(new_n11253_));
  NOR2_X1    g11189(.A1(new_n11252_), .A2(new_n11253_), .ZN(new_n11254_));
  INV_X1     g11190(.I(new_n11254_), .ZN(new_n11255_));
  XNOR2_X1   g11191(.A1(new_n341_), .A2(new_n11250_), .ZN(new_n11256_));
  NOR2_X1    g11192(.A1(new_n11237_), .A2(new_n11256_), .ZN(new_n11257_));
  AOI21_X1   g11193(.A1(new_n11237_), .A2(new_n11255_), .B(new_n11257_), .ZN(new_n11258_));
  INV_X1     g11194(.I(new_n11133_), .ZN(new_n11259_));
  AOI21_X1   g11195(.A1(new_n11189_), .A2(new_n11151_), .B(new_n11192_), .ZN(new_n11260_));
  XOR2_X1    g11196(.A1(new_n11260_), .A2(new_n11082_), .Z(new_n11261_));
  NOR2_X1    g11197(.A1(new_n11261_), .A2(new_n11259_), .ZN(new_n11262_));
  AND2_X2    g11198(.A1(new_n11261_), .A2(new_n11259_), .Z(new_n11263_));
  NOR2_X1    g11199(.A1(new_n11263_), .A2(new_n11262_), .ZN(new_n11264_));
  INV_X1     g11200(.I(new_n11188_), .ZN(new_n11265_));
  NOR2_X1    g11201(.A1(new_n11187_), .A2(new_n11265_), .ZN(new_n11266_));
  INV_X1     g11202(.I(new_n11182_), .ZN(new_n11267_));
  AOI21_X1   g11203(.A1(new_n8666_), .A2(new_n8669_), .B(new_n11267_), .ZN(new_n11268_));
  AOI21_X1   g11204(.A1(new_n11268_), .A2(new_n11185_), .B(new_n11180_), .ZN(new_n11269_));
  NOR2_X1    g11205(.A1(new_n11269_), .A2(new_n11188_), .ZN(new_n11270_));
  NOR2_X1    g11206(.A1(new_n11270_), .A2(new_n11266_), .ZN(new_n11271_));
  INV_X1     g11207(.I(new_n11271_), .ZN(new_n11272_));
  INV_X1     g11208(.I(new_n11171_), .ZN(new_n11273_));
  AOI21_X1   g11209(.A1(new_n11269_), .A2(new_n11265_), .B(new_n11273_), .ZN(new_n11274_));
  NOR2_X1    g11210(.A1(new_n11274_), .A2(new_n11151_), .ZN(new_n11275_));
  NOR2_X1    g11211(.A1(new_n11189_), .A2(new_n11150_), .ZN(new_n11276_));
  NOR2_X1    g11212(.A1(new_n11275_), .A2(new_n11276_), .ZN(new_n11277_));
  XOR2_X1    g11213(.A1(new_n11277_), .A2(new_n11272_), .Z(new_n11278_));
  INV_X1     g11214(.I(new_n11278_), .ZN(new_n11279_));
  NAND2_X1   g11215(.A1(new_n11268_), .A2(new_n3288_), .ZN(new_n11280_));
  XOR2_X1    g11216(.A1(new_n11280_), .A2(new_n11177_), .Z(new_n11281_));
  AND2_X2    g11217(.A1(new_n11281_), .A2(new_n11179_), .Z(new_n11282_));
  NOR2_X1    g11218(.A1(new_n11281_), .A2(new_n11179_), .ZN(new_n11283_));
  NOR2_X1    g11219(.A1(new_n11282_), .A2(new_n11283_), .ZN(new_n11284_));
  INV_X1     g11220(.I(new_n11284_), .ZN(new_n11285_));
  NOR2_X1    g11221(.A1(new_n11285_), .A2(new_n11272_), .ZN(new_n11286_));
  NOR2_X1    g11222(.A1(new_n11285_), .A2(new_n8662_), .ZN(new_n11287_));
  INV_X1     g11223(.I(new_n11287_), .ZN(new_n11288_));
  INV_X1     g11224(.I(new_n8689_), .ZN(new_n11289_));
  INV_X1     g11225(.I(new_n10943_), .ZN(new_n11290_));
  OAI21_X1   g11226(.A1(new_n11290_), .A2(new_n10944_), .B(new_n11289_), .ZN(new_n11291_));
  AOI21_X1   g11227(.A1(new_n8662_), .A2(new_n8688_), .B(new_n8674_), .ZN(new_n11292_));
  AOI21_X1   g11228(.A1(new_n8661_), .A2(new_n8687_), .B(new_n8673_), .ZN(new_n11293_));
  INV_X1     g11229(.I(new_n11293_), .ZN(new_n11294_));
  OAI21_X1   g11230(.A1(new_n11291_), .A2(new_n11292_), .B(new_n11294_), .ZN(new_n11295_));
  NOR2_X1    g11231(.A1(new_n11284_), .A2(new_n8661_), .ZN(new_n11296_));
  INV_X1     g11232(.I(new_n11296_), .ZN(new_n11297_));
  NAND2_X1   g11233(.A1(new_n11295_), .A2(new_n11297_), .ZN(new_n11298_));
  NOR2_X1    g11234(.A1(new_n11284_), .A2(new_n11271_), .ZN(new_n11299_));
  AOI21_X1   g11235(.A1(new_n11298_), .A2(new_n11288_), .B(new_n11299_), .ZN(new_n11300_));
  NOR2_X1    g11236(.A1(new_n11300_), .A2(new_n11286_), .ZN(new_n11301_));
  XOR2_X1    g11237(.A1(new_n11301_), .A2(new_n11271_), .Z(new_n11302_));
  NAND3_X1   g11238(.A1(new_n11302_), .A2(new_n11264_), .A3(new_n11279_), .ZN(new_n11303_));
  INV_X1     g11239(.I(new_n11264_), .ZN(new_n11304_));
  NAND2_X1   g11240(.A1(new_n11298_), .A2(new_n11288_), .ZN(new_n11305_));
  AOI21_X1   g11241(.A1(new_n11305_), .A2(new_n11284_), .B(new_n11271_), .ZN(new_n11306_));
  NOR2_X1    g11242(.A1(new_n11301_), .A2(new_n11272_), .ZN(new_n11307_));
  OAI21_X1   g11243(.A1(new_n11307_), .A2(new_n11306_), .B(new_n11279_), .ZN(new_n11308_));
  NAND2_X1   g11244(.A1(new_n11308_), .A2(new_n11304_), .ZN(new_n11309_));
  NAND2_X1   g11245(.A1(new_n11303_), .A2(new_n11309_), .ZN(new_n11310_));
  INV_X1     g11246(.I(new_n11277_), .ZN(new_n11311_));
  AOI22_X1   g11247(.A1(new_n11311_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n11272_), .ZN(new_n11312_));
  NOR2_X1    g11248(.A1(new_n11264_), .A2(new_n3175_), .ZN(new_n11313_));
  OAI21_X1   g11249(.A1(new_n11313_), .A2(new_n11312_), .B(new_n2736_), .ZN(new_n11314_));
  NOR3_X1    g11250(.A1(new_n11310_), .A2(\a[29] ), .A3(new_n11314_), .ZN(new_n11315_));
  NOR2_X1    g11251(.A1(new_n11310_), .A2(new_n11314_), .ZN(new_n11316_));
  NOR2_X1    g11252(.A1(new_n11316_), .A2(new_n74_), .ZN(new_n11317_));
  NOR2_X1    g11253(.A1(new_n11317_), .A2(new_n11315_), .ZN(new_n11318_));
  INV_X1     g11254(.I(new_n11295_), .ZN(new_n11319_));
  XOR2_X1    g11255(.A1(new_n11284_), .A2(new_n8662_), .Z(new_n11320_));
  NOR2_X1    g11256(.A1(new_n11319_), .A2(new_n11320_), .ZN(new_n11321_));
  AOI21_X1   g11257(.A1(new_n11288_), .A2(new_n11297_), .B(new_n11295_), .ZN(new_n11322_));
  OR2_X2     g11258(.A1(new_n11321_), .A2(new_n11322_), .Z(new_n11323_));
  AOI21_X1   g11259(.A1(new_n8674_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n11324_));
  OAI21_X1   g11260(.A1(new_n8661_), .A2(new_n2767_), .B(new_n11324_), .ZN(new_n11325_));
  AOI21_X1   g11261(.A1(new_n11285_), .A2(new_n3332_), .B(new_n11325_), .ZN(new_n11326_));
  AND2_X2    g11262(.A1(new_n11323_), .A2(new_n11326_), .Z(new_n11327_));
  XOR2_X1    g11263(.A1(new_n11318_), .A2(new_n11327_), .Z(new_n11328_));
  NOR2_X1    g11264(.A1(new_n11328_), .A2(new_n11258_), .ZN(new_n11329_));
  INV_X1     g11265(.I(new_n11258_), .ZN(new_n11330_));
  INV_X1     g11266(.I(new_n11318_), .ZN(new_n11331_));
  NOR2_X1    g11267(.A1(new_n11331_), .A2(new_n11327_), .ZN(new_n11332_));
  INV_X1     g11268(.I(new_n11332_), .ZN(new_n11333_));
  NAND2_X1   g11269(.A1(new_n11331_), .A2(new_n11327_), .ZN(new_n11334_));
  AOI21_X1   g11270(.A1(new_n11333_), .A2(new_n11334_), .B(new_n11330_), .ZN(new_n11335_));
  NOR2_X1    g11271(.A1(new_n11335_), .A2(new_n11329_), .ZN(new_n11336_));
  OAI21_X1   g11272(.A1(new_n11264_), .A2(new_n11271_), .B(new_n11277_), .ZN(new_n11337_));
  AOI21_X1   g11273(.A1(new_n11264_), .A2(new_n11271_), .B(new_n11277_), .ZN(new_n11338_));
  AOI21_X1   g11274(.A1(new_n11301_), .A2(new_n11337_), .B(new_n11338_), .ZN(new_n11339_));
  NOR2_X1    g11275(.A1(new_n11195_), .A2(new_n11134_), .ZN(new_n11340_));
  XNOR2_X1   g11276(.A1(new_n11199_), .A2(new_n11201_), .ZN(new_n11341_));
  NOR2_X1    g11277(.A1(new_n11340_), .A2(new_n11341_), .ZN(new_n11342_));
  INV_X1     g11278(.I(new_n11340_), .ZN(new_n11343_));
  AOI21_X1   g11279(.A1(new_n11203_), .A2(new_n11206_), .B(new_n11343_), .ZN(new_n11344_));
  NOR2_X1    g11280(.A1(new_n11344_), .A2(new_n11342_), .ZN(new_n11345_));
  INV_X1     g11281(.I(new_n11345_), .ZN(new_n11346_));
  NAND2_X1   g11282(.A1(new_n11343_), .A2(new_n11199_), .ZN(new_n11347_));
  XOR2_X1    g11283(.A1(new_n11347_), .A2(new_n11205_), .Z(new_n11348_));
  XNOR2_X1   g11284(.A1(new_n11340_), .A2(new_n11199_), .ZN(new_n11349_));
  NAND2_X1   g11285(.A1(new_n11349_), .A2(new_n11201_), .ZN(new_n11350_));
  NOR2_X1    g11286(.A1(new_n11348_), .A2(new_n11350_), .ZN(new_n11351_));
  AND2_X2    g11287(.A1(new_n11348_), .A2(new_n11350_), .Z(new_n11352_));
  NOR2_X1    g11288(.A1(new_n11352_), .A2(new_n11351_), .ZN(new_n11353_));
  INV_X1     g11289(.I(new_n11353_), .ZN(new_n11354_));
  AOI21_X1   g11290(.A1(new_n11354_), .A2(new_n11304_), .B(new_n11346_), .ZN(new_n11355_));
  INV_X1     g11291(.I(new_n11355_), .ZN(new_n11356_));
  AND2_X2    g11292(.A1(new_n11339_), .A2(new_n11356_), .Z(new_n11357_));
  AOI21_X1   g11293(.A1(new_n11353_), .A2(new_n11264_), .B(new_n11345_), .ZN(new_n11358_));
  NOR2_X1    g11294(.A1(new_n11357_), .A2(new_n11358_), .ZN(new_n11359_));
  INV_X1     g11295(.I(new_n11209_), .ZN(new_n11360_));
  INV_X1     g11296(.I(new_n11134_), .ZN(new_n11361_));
  OAI21_X1   g11297(.A1(new_n11274_), .A2(new_n11150_), .B(new_n11193_), .ZN(new_n11362_));
  AOI21_X1   g11298(.A1(new_n11362_), .A2(new_n11361_), .B(new_n11202_), .ZN(new_n11363_));
  NOR2_X1    g11299(.A1(new_n11363_), .A2(new_n11207_), .ZN(new_n11364_));
  NAND2_X1   g11300(.A1(new_n11364_), .A2(new_n11038_), .ZN(new_n11365_));
  XOR2_X1    g11301(.A1(new_n11365_), .A2(new_n11224_), .Z(new_n11366_));
  OR2_X2     g11302(.A1(new_n11366_), .A2(new_n11360_), .Z(new_n11367_));
  NAND2_X1   g11303(.A1(new_n11366_), .A2(new_n11360_), .ZN(new_n11368_));
  NAND2_X1   g11304(.A1(new_n11367_), .A2(new_n11368_), .ZN(new_n11369_));
  INV_X1     g11305(.I(new_n11369_), .ZN(new_n11370_));
  NOR2_X1    g11306(.A1(new_n11370_), .A2(new_n11354_), .ZN(new_n11371_));
  INV_X1     g11307(.I(new_n11371_), .ZN(new_n11372_));
  NOR2_X1    g11308(.A1(new_n11369_), .A2(new_n11353_), .ZN(new_n11373_));
  INV_X1     g11309(.I(new_n11373_), .ZN(new_n11374_));
  AOI21_X1   g11310(.A1(new_n11372_), .A2(new_n11374_), .B(new_n11359_), .ZN(new_n11375_));
  OR2_X2     g11311(.A1(new_n11357_), .A2(new_n11358_), .Z(new_n11376_));
  XNOR2_X1   g11312(.A1(new_n11369_), .A2(new_n11353_), .ZN(new_n11377_));
  NOR2_X1    g11313(.A1(new_n11376_), .A2(new_n11377_), .ZN(new_n11378_));
  NOR2_X1    g11314(.A1(new_n11378_), .A2(new_n11375_), .ZN(new_n11379_));
  OAI22_X1   g11315(.A1(new_n11353_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n11345_), .ZN(new_n11380_));
  NAND2_X1   g11316(.A1(new_n11370_), .A2(new_n3317_), .ZN(new_n11381_));
  AOI21_X1   g11317(.A1(new_n11381_), .A2(new_n11380_), .B(new_n3260_), .ZN(new_n11382_));
  NAND2_X1   g11318(.A1(new_n11379_), .A2(new_n11382_), .ZN(new_n11383_));
  XOR2_X1    g11319(.A1(new_n11383_), .A2(\a[26] ), .Z(new_n11384_));
  XOR2_X1    g11320(.A1(new_n10964_), .A2(new_n11238_), .Z(new_n11385_));
  OAI21_X1   g11321(.A1(new_n11236_), .A2(new_n10965_), .B(new_n11234_), .ZN(new_n11386_));
  OAI21_X1   g11322(.A1(new_n11234_), .A2(new_n11385_), .B(new_n11386_), .ZN(new_n11387_));
  NOR2_X1    g11323(.A1(new_n11301_), .A2(new_n11278_), .ZN(new_n11388_));
  XOR2_X1    g11324(.A1(new_n11277_), .A2(new_n11271_), .Z(new_n11389_));
  NOR3_X1    g11325(.A1(new_n11300_), .A2(new_n11286_), .A3(new_n11389_), .ZN(new_n11390_));
  OR2_X2     g11326(.A1(new_n11388_), .A2(new_n11390_), .Z(new_n11391_));
  OAI22_X1   g11327(.A1(new_n11284_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n11271_), .ZN(new_n11392_));
  NAND2_X1   g11328(.A1(new_n11311_), .A2(new_n2750_), .ZN(new_n11393_));
  AOI21_X1   g11329(.A1(new_n11392_), .A2(new_n11393_), .B(new_n2737_), .ZN(new_n11394_));
  NAND2_X1   g11330(.A1(new_n11391_), .A2(new_n11394_), .ZN(new_n11395_));
  XOR2_X1    g11331(.A1(new_n11395_), .A2(\a[29] ), .Z(new_n11396_));
  OR2_X2     g11332(.A1(new_n11396_), .A2(new_n11387_), .Z(new_n11397_));
  NOR3_X1    g11333(.A1(new_n289_), .A2(new_n591_), .A3(new_n654_), .ZN(new_n11398_));
  NOR3_X1    g11334(.A1(new_n2930_), .A2(new_n90_), .A3(new_n374_), .ZN(new_n11399_));
  NOR4_X1    g11335(.A1(new_n281_), .A2(new_n366_), .A3(new_n403_), .A4(new_n782_), .ZN(new_n11400_));
  INV_X1     g11336(.I(new_n11400_), .ZN(new_n11401_));
  NAND4_X1   g11337(.A1(new_n11399_), .A2(new_n3510_), .A3(new_n11398_), .A4(new_n11401_), .ZN(new_n11402_));
  NOR4_X1    g11338(.A1(new_n1457_), .A2(new_n170_), .A3(new_n510_), .A4(new_n695_), .ZN(new_n11403_));
  NOR4_X1    g11339(.A1(new_n1415_), .A2(new_n713_), .A3(new_n1247_), .A4(new_n2677_), .ZN(new_n11404_));
  NAND3_X1   g11340(.A1(new_n11404_), .A2(new_n1231_), .A3(new_n11403_), .ZN(new_n11405_));
  NOR3_X1    g11341(.A1(new_n11405_), .A2(new_n1480_), .A3(new_n11402_), .ZN(new_n11406_));
  INV_X1     g11342(.I(new_n1485_), .ZN(new_n11407_));
  NAND4_X1   g11343(.A1(new_n653_), .A2(new_n2275_), .A3(new_n331_), .A4(new_n1883_), .ZN(new_n11408_));
  NAND4_X1   g11344(.A1(new_n373_), .A2(new_n467_), .A3(new_n709_), .A4(new_n1216_), .ZN(new_n11409_));
  NAND4_X1   g11345(.A1(new_n2119_), .A2(new_n182_), .A3(new_n1025_), .A4(new_n309_), .ZN(new_n11410_));
  NAND4_X1   g11346(.A1(new_n2544_), .A2(new_n3479_), .A3(new_n11409_), .A4(new_n11410_), .ZN(new_n11411_));
  NOR3_X1    g11347(.A1(new_n11407_), .A2(new_n11411_), .A3(new_n11408_), .ZN(new_n11412_));
  NAND3_X1   g11348(.A1(new_n11406_), .A2(new_n3933_), .A3(new_n11412_), .ZN(new_n11413_));
  INV_X1     g11349(.I(new_n11413_), .ZN(new_n11414_));
  NAND2_X1   g11350(.A1(new_n10990_), .A2(new_n11414_), .ZN(new_n11415_));
  XNOR2_X1   g11351(.A1(new_n8681_), .A2(new_n8687_), .ZN(new_n11416_));
  INV_X1     g11352(.I(new_n11416_), .ZN(new_n11417_));
  NAND2_X1   g11353(.A1(new_n10943_), .A2(new_n11417_), .ZN(new_n11418_));
  NOR2_X1    g11354(.A1(new_n8689_), .A2(new_n10944_), .ZN(new_n11419_));
  OAI21_X1   g11355(.A1(new_n10943_), .A2(new_n11419_), .B(new_n11418_), .ZN(new_n11420_));
  NOR2_X1    g11356(.A1(new_n8687_), .A2(new_n2772_), .ZN(new_n11421_));
  NOR2_X1    g11357(.A1(new_n8681_), .A2(new_n2767_), .ZN(new_n11422_));
  NOR2_X1    g11358(.A1(new_n8694_), .A2(new_n2771_), .ZN(new_n11423_));
  NOR4_X1    g11359(.A1(new_n11422_), .A2(new_n11421_), .A3(new_n2763_), .A4(new_n11423_), .ZN(new_n11424_));
  INV_X1     g11360(.I(new_n10990_), .ZN(new_n11425_));
  NAND2_X1   g11361(.A1(new_n11425_), .A2(new_n11413_), .ZN(new_n11426_));
  NAND3_X1   g11362(.A1(new_n11420_), .A2(new_n11424_), .A3(new_n11426_), .ZN(new_n11427_));
  XOR2_X1    g11363(.A1(new_n8673_), .A2(new_n8687_), .Z(new_n11428_));
  INV_X1     g11364(.I(new_n11428_), .ZN(new_n11429_));
  NAND2_X1   g11365(.A1(new_n10946_), .A2(new_n11429_), .ZN(new_n11430_));
  OAI21_X1   g11366(.A1(new_n10946_), .A2(new_n10956_), .B(new_n11430_), .ZN(new_n11431_));
  NOR2_X1    g11367(.A1(new_n8673_), .A2(new_n2772_), .ZN(new_n11432_));
  NOR2_X1    g11368(.A1(new_n8687_), .A2(new_n2767_), .ZN(new_n11433_));
  NOR2_X1    g11369(.A1(new_n8681_), .A2(new_n2771_), .ZN(new_n11434_));
  NOR4_X1    g11370(.A1(new_n11432_), .A2(new_n11434_), .A3(new_n11433_), .A4(new_n2763_), .ZN(new_n11435_));
  NAND2_X1   g11371(.A1(new_n11431_), .A2(new_n11435_), .ZN(new_n11436_));
  AOI21_X1   g11372(.A1(new_n11415_), .A2(new_n11427_), .B(new_n11436_), .ZN(new_n11437_));
  INV_X1     g11373(.I(new_n11007_), .ZN(new_n11438_));
  AOI21_X1   g11374(.A1(new_n11438_), .A2(new_n11233_), .B(new_n11232_), .ZN(new_n11439_));
  XNOR2_X1   g11375(.A1(new_n11006_), .A2(new_n10990_), .ZN(new_n11440_));
  INV_X1     g11376(.I(new_n11440_), .ZN(new_n11441_));
  AOI21_X1   g11377(.A1(new_n11232_), .A2(new_n11441_), .B(new_n11439_), .ZN(new_n11442_));
  NAND2_X1   g11378(.A1(new_n11427_), .A2(new_n11415_), .ZN(new_n11443_));
  INV_X1     g11379(.I(new_n11436_), .ZN(new_n11444_));
  NOR2_X1    g11380(.A1(new_n11444_), .A2(new_n11443_), .ZN(new_n11445_));
  INV_X1     g11381(.I(new_n11445_), .ZN(new_n11446_));
  AOI21_X1   g11382(.A1(new_n11446_), .A2(new_n11442_), .B(new_n11437_), .ZN(new_n11447_));
  INV_X1     g11383(.I(new_n11447_), .ZN(new_n11448_));
  NAND2_X1   g11384(.A1(new_n11396_), .A2(new_n11387_), .ZN(new_n11449_));
  NAND2_X1   g11385(.A1(new_n11449_), .A2(new_n11448_), .ZN(new_n11450_));
  NAND2_X1   g11386(.A1(new_n11450_), .A2(new_n11397_), .ZN(new_n11451_));
  XOR2_X1    g11387(.A1(new_n11384_), .A2(new_n11451_), .Z(new_n11452_));
  NOR2_X1    g11388(.A1(new_n11452_), .A2(new_n11336_), .ZN(new_n11453_));
  INV_X1     g11389(.I(new_n11384_), .ZN(new_n11454_));
  NOR2_X1    g11390(.A1(new_n11454_), .A2(new_n11451_), .ZN(new_n11455_));
  INV_X1     g11391(.I(new_n11455_), .ZN(new_n11456_));
  NAND2_X1   g11392(.A1(new_n11454_), .A2(new_n11451_), .ZN(new_n11457_));
  NAND2_X1   g11393(.A1(new_n11456_), .A2(new_n11457_), .ZN(new_n11458_));
  AOI21_X1   g11394(.A1(new_n11336_), .A2(new_n11458_), .B(new_n11453_), .ZN(new_n11459_));
  INV_X1     g11395(.I(new_n11225_), .ZN(new_n11460_));
  NOR4_X1    g11396(.A1(new_n11363_), .A2(new_n11037_), .A3(new_n11207_), .A4(new_n11460_), .ZN(new_n11461_));
  NOR3_X1    g11397(.A1(new_n11037_), .A2(new_n11209_), .A3(new_n11224_), .ZN(new_n11462_));
  NAND2_X1   g11398(.A1(new_n11364_), .A2(new_n11462_), .ZN(new_n11463_));
  AOI21_X1   g11399(.A1(new_n11376_), .A2(new_n11353_), .B(new_n11369_), .ZN(new_n11464_));
  NOR3_X1    g11400(.A1(new_n11464_), .A2(new_n11461_), .A3(new_n11463_), .ZN(new_n11465_));
  INV_X1     g11401(.I(new_n11463_), .ZN(new_n11466_));
  AOI21_X1   g11402(.A1(new_n11464_), .A2(new_n11466_), .B(new_n11226_), .ZN(new_n11467_));
  OR2_X2     g11403(.A1(new_n11465_), .A2(new_n11467_), .Z(new_n11468_));
  NAND2_X1   g11404(.A1(new_n3780_), .A2(new_n3306_), .ZN(new_n11469_));
  AND3_X2    g11405(.A1(new_n11463_), .A2(new_n5291_), .A3(new_n11469_), .Z(new_n11470_));
  NOR4_X1    g11406(.A1(new_n11468_), .A2(new_n3302_), .A3(new_n11461_), .A4(new_n11470_), .ZN(new_n11471_));
  XOR2_X1    g11407(.A1(new_n11471_), .A2(new_n84_), .Z(new_n11472_));
  NOR2_X1    g11408(.A1(new_n11459_), .A2(new_n11472_), .ZN(new_n11473_));
  NOR3_X1    g11409(.A1(new_n3874_), .A2(new_n236_), .A3(new_n324_), .ZN(new_n11474_));
  NAND2_X1   g11410(.A1(new_n1790_), .A2(new_n1793_), .ZN(new_n11475_));
  INV_X1     g11411(.I(new_n2542_), .ZN(new_n11476_));
  NAND4_X1   g11412(.A1(new_n3198_), .A2(new_n271_), .A3(new_n1590_), .A4(new_n1096_), .ZN(new_n11477_));
  INV_X1     g11413(.I(new_n2622_), .ZN(new_n11478_));
  NOR2_X1    g11414(.A1(new_n11478_), .A2(new_n3218_), .ZN(new_n11479_));
  NAND4_X1   g11415(.A1(new_n311_), .A2(new_n701_), .A3(new_n435_), .A4(new_n1216_), .ZN(new_n11480_));
  NAND4_X1   g11416(.A1(new_n11479_), .A2(new_n3970_), .A3(new_n11477_), .A4(new_n11480_), .ZN(new_n11481_));
  NOR4_X1    g11417(.A1(new_n11476_), .A2(new_n11475_), .A3(new_n2400_), .A4(new_n11481_), .ZN(new_n11482_));
  NAND2_X1   g11418(.A1(new_n11482_), .A2(new_n11474_), .ZN(new_n11483_));
  NOR4_X1    g11419(.A1(new_n774_), .A2(new_n456_), .A3(new_n1084_), .A4(new_n591_), .ZN(new_n11484_));
  NOR3_X1    g11420(.A1(new_n11484_), .A2(new_n939_), .A3(new_n1381_), .ZN(new_n11485_));
  NOR4_X1    g11421(.A1(new_n3470_), .A2(new_n234_), .A3(new_n437_), .A4(new_n2306_), .ZN(new_n11486_));
  NAND4_X1   g11422(.A1(new_n903_), .A2(new_n2931_), .A3(new_n11485_), .A4(new_n11486_), .ZN(new_n11487_));
  INV_X1     g11423(.I(new_n3497_), .ZN(new_n11488_));
  NOR2_X1    g11424(.A1(new_n1410_), .A2(new_n2092_), .ZN(new_n11489_));
  NAND4_X1   g11425(.A1(new_n1216_), .A2(new_n423_), .A3(new_n551_), .A4(new_n1059_), .ZN(new_n11490_));
  NAND3_X1   g11426(.A1(new_n11489_), .A2(new_n11488_), .A3(new_n11490_), .ZN(new_n11491_));
  NOR4_X1    g11427(.A1(new_n11487_), .A2(new_n2212_), .A3(new_n2228_), .A4(new_n11491_), .ZN(new_n11492_));
  NAND2_X1   g11428(.A1(new_n6539_), .A2(new_n11492_), .ZN(new_n11493_));
  NOR2_X1    g11429(.A1(new_n11483_), .A2(new_n11493_), .ZN(new_n11494_));
  INV_X1     g11430(.I(new_n11494_), .ZN(new_n11495_));
  NAND2_X1   g11431(.A1(new_n6091_), .A2(new_n6094_), .ZN(new_n11496_));
  NOR3_X1    g11432(.A1(new_n11496_), .A2(new_n6081_), .A3(new_n6180_), .ZN(new_n11497_));
  NOR2_X1    g11433(.A1(new_n11497_), .A2(new_n3521_), .ZN(new_n11498_));
  INV_X1     g11434(.I(new_n11498_), .ZN(new_n11499_));
  NOR2_X1    g11435(.A1(new_n11461_), .A2(new_n11499_), .ZN(new_n11500_));
  NOR2_X1    g11436(.A1(new_n11461_), .A2(new_n11497_), .ZN(new_n11501_));
  NOR2_X1    g11437(.A1(new_n11501_), .A2(\a[14] ), .ZN(new_n11502_));
  NOR2_X1    g11438(.A1(new_n11502_), .A2(new_n11500_), .ZN(new_n11503_));
  NAND2_X1   g11439(.A1(new_n11483_), .A2(new_n11493_), .ZN(new_n11504_));
  NAND2_X1   g11440(.A1(new_n11503_), .A2(new_n11504_), .ZN(new_n11505_));
  NAND2_X1   g11441(.A1(new_n11505_), .A2(new_n11495_), .ZN(new_n11506_));
  NOR2_X1    g11442(.A1(new_n460_), .A2(new_n899_), .ZN(new_n11507_));
  NOR2_X1    g11443(.A1(new_n2976_), .A2(new_n1381_), .ZN(new_n11508_));
  NAND4_X1   g11444(.A1(new_n913_), .A2(new_n1129_), .A3(new_n301_), .A4(new_n1446_), .ZN(new_n11509_));
  NAND4_X1   g11445(.A1(new_n1628_), .A2(new_n438_), .A3(new_n1753_), .A4(new_n675_), .ZN(new_n11510_));
  NAND4_X1   g11446(.A1(new_n11508_), .A2(new_n11507_), .A3(new_n11509_), .A4(new_n11510_), .ZN(new_n11511_));
  NOR4_X1    g11447(.A1(new_n714_), .A2(new_n117_), .A3(new_n381_), .A4(new_n262_), .ZN(new_n11512_));
  NOR3_X1    g11448(.A1(new_n11512_), .A2(new_n86_), .A3(new_n1167_), .ZN(new_n11513_));
  INV_X1     g11449(.I(new_n11513_), .ZN(new_n11514_));
  NOR4_X1    g11450(.A1(new_n11511_), .A2(new_n3505_), .A3(new_n4592_), .A4(new_n11514_), .ZN(new_n11515_));
  NAND4_X1   g11451(.A1(new_n11515_), .A2(new_n1832_), .A3(new_n1662_), .A4(new_n773_), .ZN(new_n11516_));
  INV_X1     g11452(.I(new_n11516_), .ZN(new_n11517_));
  NOR4_X1    g11453(.A1(new_n1245_), .A2(new_n316_), .A3(new_n730_), .A4(new_n1954_), .ZN(new_n11518_));
  INV_X1     g11454(.I(new_n11518_), .ZN(new_n11519_));
  NOR4_X1    g11455(.A1(new_n81_), .A2(new_n76_), .A3(new_n247_), .A4(new_n718_), .ZN(new_n11520_));
  NOR4_X1    g11456(.A1(new_n11519_), .A2(new_n183_), .A3(new_n908_), .A4(new_n11520_), .ZN(new_n11521_));
  INV_X1     g11457(.I(new_n11521_), .ZN(new_n11522_));
  INV_X1     g11458(.I(new_n2339_), .ZN(new_n11523_));
  NOR2_X1    g11459(.A1(new_n11523_), .A2(new_n4022_), .ZN(new_n11524_));
  NAND4_X1   g11460(.A1(new_n1335_), .A2(new_n208_), .A3(new_n665_), .A4(new_n188_), .ZN(new_n11525_));
  NAND4_X1   g11461(.A1(new_n11524_), .A2(new_n1291_), .A3(new_n1467_), .A4(new_n11525_), .ZN(new_n11526_));
  NOR3_X1    g11462(.A1(new_n198_), .A2(new_n312_), .A3(new_n430_), .ZN(new_n11527_));
  NAND4_X1   g11463(.A1(new_n2788_), .A2(new_n516_), .A3(new_n2275_), .A4(new_n11527_), .ZN(new_n11528_));
  NOR4_X1    g11464(.A1(new_n11522_), .A2(new_n1978_), .A3(new_n11526_), .A4(new_n11528_), .ZN(new_n11529_));
  NAND2_X1   g11465(.A1(new_n11517_), .A2(new_n11529_), .ZN(new_n11530_));
  XOR2_X1    g11466(.A1(new_n8710_), .A2(new_n8719_), .Z(new_n11531_));
  AOI21_X1   g11467(.A1(new_n10933_), .A2(new_n8728_), .B(new_n11531_), .ZN(new_n11532_));
  INV_X1     g11468(.I(new_n11532_), .ZN(new_n11533_));
  INV_X1     g11469(.I(new_n8720_), .ZN(new_n11534_));
  AND2_X2    g11470(.A1(new_n11534_), .A2(new_n10935_), .Z(new_n11535_));
  OAI21_X1   g11471(.A1(new_n10934_), .A2(new_n11535_), .B(new_n11533_), .ZN(new_n11536_));
  AOI21_X1   g11472(.A1(new_n8719_), .A2(new_n3189_), .B(new_n2763_), .ZN(new_n11537_));
  OAI21_X1   g11473(.A1(new_n8725_), .A2(new_n2771_), .B(new_n11537_), .ZN(new_n11538_));
  AOI21_X1   g11474(.A1(new_n8711_), .A2(new_n3332_), .B(new_n11538_), .ZN(new_n11539_));
  AOI21_X1   g11475(.A1(new_n11536_), .A2(new_n11539_), .B(new_n11530_), .ZN(new_n11540_));
  INV_X1     g11476(.I(new_n11540_), .ZN(new_n11541_));
  NAND2_X1   g11477(.A1(new_n11506_), .A2(new_n11541_), .ZN(new_n11542_));
  INV_X1     g11478(.I(new_n11530_), .ZN(new_n11543_));
  NAND2_X1   g11479(.A1(new_n11536_), .A2(new_n11539_), .ZN(new_n11544_));
  NOR2_X1    g11480(.A1(new_n11544_), .A2(new_n11543_), .ZN(new_n11545_));
  INV_X1     g11481(.I(new_n11545_), .ZN(new_n11546_));
  NAND2_X1   g11482(.A1(new_n11542_), .A2(new_n11546_), .ZN(new_n11547_));
  NOR4_X1    g11483(.A1(new_n1146_), .A2(new_n549_), .A3(new_n611_), .A4(new_n732_), .ZN(new_n11548_));
  NOR4_X1    g11484(.A1(new_n11548_), .A2(new_n397_), .A3(new_n633_), .A4(new_n1991_), .ZN(new_n11549_));
  INV_X1     g11485(.I(new_n11549_), .ZN(new_n11550_));
  NOR2_X1    g11486(.A1(new_n335_), .A2(new_n841_), .ZN(new_n11551_));
  NAND4_X1   g11487(.A1(new_n2013_), .A2(new_n2219_), .A3(new_n2795_), .A4(new_n11551_), .ZN(new_n11552_));
  NAND3_X1   g11488(.A1(new_n1086_), .A2(new_n80_), .A3(new_n992_), .ZN(new_n11553_));
  NAND2_X1   g11489(.A1(new_n1767_), .A2(new_n722_), .ZN(new_n11554_));
  NOR4_X1    g11490(.A1(new_n11550_), .A2(new_n11552_), .A3(new_n11553_), .A4(new_n11554_), .ZN(new_n11555_));
  INV_X1     g11491(.I(new_n1351_), .ZN(new_n11556_));
  NOR4_X1    g11492(.A1(new_n214_), .A2(new_n510_), .A3(new_n660_), .A4(new_n902_), .ZN(new_n11557_));
  NOR3_X1    g11493(.A1(new_n11556_), .A2(new_n1735_), .A3(new_n11557_), .ZN(new_n11558_));
  AND2_X2    g11494(.A1(new_n3969_), .A2(new_n11558_), .Z(new_n11559_));
  NAND4_X1   g11495(.A1(new_n11559_), .A2(new_n1655_), .A3(new_n3029_), .A4(new_n11555_), .ZN(new_n11560_));
  NOR2_X1    g11496(.A1(new_n11543_), .A2(new_n11560_), .ZN(new_n11561_));
  INV_X1     g11497(.I(new_n11561_), .ZN(new_n11562_));
  NAND2_X1   g11498(.A1(new_n11543_), .A2(new_n11560_), .ZN(new_n11563_));
  INV_X1     g11499(.I(new_n11563_), .ZN(new_n11564_));
  AOI21_X1   g11500(.A1(new_n11547_), .A2(new_n11562_), .B(new_n11564_), .ZN(new_n11565_));
  INV_X1     g11501(.I(new_n11565_), .ZN(new_n11566_));
  NAND2_X1   g11502(.A1(new_n4470_), .A2(new_n4297_), .ZN(new_n11567_));
  NOR3_X1    g11503(.A1(new_n11567_), .A2(new_n4292_), .A3(new_n4295_), .ZN(new_n11568_));
  NOR2_X1    g11504(.A1(new_n11568_), .A2(new_n3372_), .ZN(new_n11569_));
  INV_X1     g11505(.I(new_n11569_), .ZN(new_n11570_));
  NOR2_X1    g11506(.A1(new_n11461_), .A2(new_n11570_), .ZN(new_n11571_));
  NOR2_X1    g11507(.A1(new_n11461_), .A2(new_n11568_), .ZN(new_n11572_));
  NOR2_X1    g11508(.A1(new_n11572_), .A2(\a[17] ), .ZN(new_n11573_));
  NOR2_X1    g11509(.A1(new_n11573_), .A2(new_n11571_), .ZN(new_n11574_));
  NOR3_X1    g11510(.A1(new_n805_), .A2(new_n152_), .A3(new_n698_), .ZN(new_n11575_));
  NAND4_X1   g11511(.A1(new_n1018_), .A2(new_n1506_), .A3(new_n669_), .A4(new_n432_), .ZN(new_n11576_));
  NAND4_X1   g11512(.A1(new_n246_), .A2(new_n807_), .A3(new_n840_), .A4(new_n672_), .ZN(new_n11577_));
  NOR2_X1    g11513(.A1(new_n4752_), .A2(new_n163_), .ZN(new_n11578_));
  NAND4_X1   g11514(.A1(new_n11575_), .A2(new_n11578_), .A3(new_n11576_), .A4(new_n11577_), .ZN(new_n11579_));
  NOR4_X1    g11515(.A1(new_n2703_), .A2(new_n906_), .A3(new_n603_), .A4(new_n1157_), .ZN(new_n11580_));
  NAND4_X1   g11516(.A1(new_n11580_), .A2(new_n201_), .A3(new_n1608_), .A4(new_n2339_), .ZN(new_n11581_));
  NOR4_X1    g11517(.A1(new_n11581_), .A2(new_n1906_), .A3(new_n10986_), .A4(new_n11579_), .ZN(new_n11582_));
  NOR2_X1    g11518(.A1(new_n11067_), .A2(new_n3692_), .ZN(new_n11583_));
  NAND2_X1   g11519(.A1(new_n11583_), .A2(new_n11582_), .ZN(new_n11584_));
  NAND2_X1   g11520(.A1(new_n11584_), .A2(new_n11560_), .ZN(new_n11585_));
  NOR2_X1    g11521(.A1(new_n11584_), .A2(new_n11560_), .ZN(new_n11586_));
  INV_X1     g11522(.I(new_n11586_), .ZN(new_n11587_));
  AOI21_X1   g11523(.A1(new_n11585_), .A2(new_n11587_), .B(new_n11574_), .ZN(new_n11588_));
  XNOR2_X1   g11524(.A1(new_n11584_), .A2(new_n11560_), .ZN(new_n11589_));
  INV_X1     g11525(.I(new_n11589_), .ZN(new_n11590_));
  AOI21_X1   g11526(.A1(new_n11574_), .A2(new_n11590_), .B(new_n11588_), .ZN(new_n11591_));
  OAI21_X1   g11527(.A1(new_n8703_), .A2(new_n10939_), .B(new_n10938_), .ZN(new_n11592_));
  XOR2_X1    g11528(.A1(new_n8701_), .A2(new_n8694_), .Z(new_n11593_));
  NAND3_X1   g11529(.A1(new_n10950_), .A2(new_n8713_), .A3(new_n11593_), .ZN(new_n11594_));
  AND2_X2    g11530(.A1(new_n11592_), .A2(new_n11594_), .Z(new_n11595_));
  NOR2_X1    g11531(.A1(new_n8694_), .A2(new_n2772_), .ZN(new_n11596_));
  NOR2_X1    g11532(.A1(new_n8701_), .A2(new_n2767_), .ZN(new_n11597_));
  OAI21_X1   g11533(.A1(new_n8710_), .A2(new_n2771_), .B(new_n2763_), .ZN(new_n11598_));
  NOR4_X1    g11534(.A1(new_n11595_), .A2(new_n11596_), .A3(new_n11597_), .A4(new_n11598_), .ZN(new_n11599_));
  NOR2_X1    g11535(.A1(new_n11591_), .A2(new_n11599_), .ZN(new_n11600_));
  INV_X1     g11536(.I(new_n11600_), .ZN(new_n11601_));
  NAND2_X1   g11537(.A1(new_n11591_), .A2(new_n11599_), .ZN(new_n11602_));
  INV_X1     g11538(.I(new_n11602_), .ZN(new_n11603_));
  AOI21_X1   g11539(.A1(new_n11566_), .A2(new_n11601_), .B(new_n11603_), .ZN(new_n11604_));
  NAND2_X1   g11540(.A1(new_n11574_), .A2(new_n11585_), .ZN(new_n11605_));
  NAND2_X1   g11541(.A1(new_n11605_), .A2(new_n11587_), .ZN(new_n11606_));
  INV_X1     g11542(.I(new_n8695_), .ZN(new_n11607_));
  OAI22_X1   g11543(.A1(new_n10951_), .A2(new_n8703_), .B1(new_n11607_), .B2(new_n10942_), .ZN(new_n11608_));
  XOR2_X1    g11544(.A1(new_n8681_), .A2(new_n8696_), .Z(new_n11609_));
  INV_X1     g11545(.I(new_n11609_), .ZN(new_n11610_));
  NAND2_X1   g11546(.A1(new_n10941_), .A2(new_n11610_), .ZN(new_n11611_));
  NAND2_X1   g11547(.A1(new_n11611_), .A2(new_n11608_), .ZN(new_n11612_));
  NAND2_X1   g11548(.A1(new_n8682_), .A2(new_n3332_), .ZN(new_n11613_));
  NAND2_X1   g11549(.A1(new_n8696_), .A2(new_n3189_), .ZN(new_n11614_));
  AOI21_X1   g11550(.A1(new_n8702_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n11615_));
  NAND4_X1   g11551(.A1(new_n11612_), .A2(new_n11613_), .A3(new_n11614_), .A4(new_n11615_), .ZN(new_n11616_));
  XOR2_X1    g11552(.A1(new_n11616_), .A2(new_n10990_), .Z(new_n11617_));
  INV_X1     g11553(.I(new_n11617_), .ZN(new_n11618_));
  NOR2_X1    g11554(.A1(new_n11616_), .A2(new_n11425_), .ZN(new_n11619_));
  INV_X1     g11555(.I(new_n11619_), .ZN(new_n11620_));
  NAND2_X1   g11556(.A1(new_n11616_), .A2(new_n11425_), .ZN(new_n11621_));
  AOI21_X1   g11557(.A1(new_n11620_), .A2(new_n11621_), .B(new_n11606_), .ZN(new_n11622_));
  AOI21_X1   g11558(.A1(new_n11618_), .A2(new_n11606_), .B(new_n11622_), .ZN(new_n11623_));
  NOR2_X1    g11559(.A1(new_n10960_), .A2(new_n10957_), .ZN(new_n11624_));
  OAI22_X1   g11560(.A1(new_n8673_), .A2(new_n2742_), .B1(new_n8687_), .B2(new_n2747_), .ZN(new_n11625_));
  NAND2_X1   g11561(.A1(new_n8662_), .A2(new_n2750_), .ZN(new_n11626_));
  AOI21_X1   g11562(.A1(new_n11626_), .A2(new_n11625_), .B(new_n2737_), .ZN(new_n11627_));
  NAND2_X1   g11563(.A1(new_n11624_), .A2(new_n11627_), .ZN(new_n11628_));
  XOR2_X1    g11564(.A1(new_n11628_), .A2(\a[29] ), .Z(new_n11629_));
  INV_X1     g11565(.I(new_n11629_), .ZN(new_n11630_));
  NOR2_X1    g11566(.A1(new_n11630_), .A2(new_n11623_), .ZN(new_n11631_));
  NOR2_X1    g11567(.A1(new_n11631_), .A2(new_n11604_), .ZN(new_n11632_));
  INV_X1     g11568(.I(new_n11623_), .ZN(new_n11633_));
  NOR2_X1    g11569(.A1(new_n11629_), .A2(new_n11633_), .ZN(new_n11634_));
  NOR2_X1    g11570(.A1(new_n11632_), .A2(new_n11634_), .ZN(new_n11635_));
  AOI21_X1   g11571(.A1(new_n11606_), .A2(new_n11621_), .B(new_n11619_), .ZN(new_n11636_));
  INV_X1     g11572(.I(new_n11636_), .ZN(new_n11637_));
  NAND2_X1   g11573(.A1(new_n11420_), .A2(new_n11424_), .ZN(new_n11638_));
  AOI21_X1   g11574(.A1(new_n11415_), .A2(new_n11426_), .B(new_n11638_), .ZN(new_n11639_));
  XOR2_X1    g11575(.A1(new_n10990_), .A2(new_n11413_), .Z(new_n11640_));
  AOI21_X1   g11576(.A1(new_n11420_), .A2(new_n11424_), .B(new_n11640_), .ZN(new_n11641_));
  NOR3_X1    g11577(.A1(new_n11637_), .A2(new_n11639_), .A3(new_n11641_), .ZN(new_n11642_));
  NOR2_X1    g11578(.A1(new_n11635_), .A2(new_n11642_), .ZN(new_n11643_));
  NOR2_X1    g11579(.A1(new_n11639_), .A2(new_n11641_), .ZN(new_n11644_));
  NOR2_X1    g11580(.A1(new_n11644_), .A2(new_n11636_), .ZN(new_n11645_));
  NOR2_X1    g11581(.A1(new_n11643_), .A2(new_n11645_), .ZN(new_n11646_));
  INV_X1     g11582(.I(new_n11646_), .ZN(new_n11647_));
  XOR2_X1    g11583(.A1(new_n11436_), .A2(new_n11443_), .Z(new_n11648_));
  OAI21_X1   g11584(.A1(new_n11445_), .A2(new_n11437_), .B(new_n11442_), .ZN(new_n11649_));
  OAI21_X1   g11585(.A1(new_n11442_), .A2(new_n11648_), .B(new_n11649_), .ZN(new_n11650_));
  OAI21_X1   g11586(.A1(new_n11286_), .A2(new_n11299_), .B(new_n11305_), .ZN(new_n11651_));
  XOR2_X1    g11587(.A1(new_n11284_), .A2(new_n11272_), .Z(new_n11652_));
  INV_X1     g11588(.I(new_n11652_), .ZN(new_n11653_));
  NAND3_X1   g11589(.A1(new_n11298_), .A2(new_n11288_), .A3(new_n11653_), .ZN(new_n11654_));
  AND2_X2    g11590(.A1(new_n11651_), .A2(new_n11654_), .Z(new_n11655_));
  OAI22_X1   g11591(.A1(new_n11284_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8661_), .ZN(new_n11656_));
  NAND2_X1   g11592(.A1(new_n11272_), .A2(new_n2750_), .ZN(new_n11657_));
  AOI21_X1   g11593(.A1(new_n11656_), .A2(new_n11657_), .B(new_n2737_), .ZN(new_n11658_));
  NAND2_X1   g11594(.A1(new_n11655_), .A2(new_n11658_), .ZN(new_n11659_));
  XOR2_X1    g11595(.A1(new_n11659_), .A2(\a[29] ), .Z(new_n11660_));
  INV_X1     g11596(.I(new_n11660_), .ZN(new_n11661_));
  NOR2_X1    g11597(.A1(new_n11661_), .A2(new_n11650_), .ZN(new_n11662_));
  INV_X1     g11598(.I(new_n11662_), .ZN(new_n11663_));
  INV_X1     g11599(.I(new_n11650_), .ZN(new_n11664_));
  NOR2_X1    g11600(.A1(new_n11660_), .A2(new_n11664_), .ZN(new_n11665_));
  AOI21_X1   g11601(.A1(new_n11647_), .A2(new_n11663_), .B(new_n11665_), .ZN(new_n11666_));
  INV_X1     g11602(.I(new_n11666_), .ZN(new_n11667_));
  XNOR2_X1   g11603(.A1(new_n11396_), .A2(new_n11387_), .ZN(new_n11668_));
  NAND2_X1   g11604(.A1(new_n11397_), .A2(new_n11449_), .ZN(new_n11669_));
  NAND2_X1   g11605(.A1(new_n11669_), .A2(new_n11447_), .ZN(new_n11670_));
  OAI21_X1   g11606(.A1(new_n11447_), .A2(new_n11668_), .B(new_n11670_), .ZN(new_n11671_));
  XOR2_X1    g11607(.A1(new_n11339_), .A2(new_n11304_), .Z(new_n11672_));
  XOR2_X1    g11608(.A1(new_n11339_), .A2(new_n11346_), .Z(new_n11673_));
  INV_X1     g11609(.I(new_n11673_), .ZN(new_n11674_));
  NOR3_X1    g11610(.A1(new_n11674_), .A2(new_n11672_), .A3(new_n11354_), .ZN(new_n11675_));
  INV_X1     g11611(.I(new_n11672_), .ZN(new_n11676_));
  AOI21_X1   g11612(.A1(new_n11676_), .A2(new_n11673_), .B(new_n11353_), .ZN(new_n11677_));
  OR2_X2     g11613(.A1(new_n11675_), .A2(new_n11677_), .Z(new_n11678_));
  OAI22_X1   g11614(.A1(new_n11264_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n11345_), .ZN(new_n11679_));
  NAND2_X1   g11615(.A1(new_n11354_), .A2(new_n3317_), .ZN(new_n11680_));
  AOI21_X1   g11616(.A1(new_n11680_), .A2(new_n11679_), .B(new_n3260_), .ZN(new_n11681_));
  NAND2_X1   g11617(.A1(new_n11678_), .A2(new_n11681_), .ZN(new_n11682_));
  XOR2_X1    g11618(.A1(new_n11682_), .A2(\a[26] ), .Z(new_n11683_));
  NAND2_X1   g11619(.A1(new_n11671_), .A2(new_n11683_), .ZN(new_n11684_));
  NOR2_X1    g11620(.A1(new_n11671_), .A2(new_n11683_), .ZN(new_n11685_));
  AOI21_X1   g11621(.A1(new_n11667_), .A2(new_n11684_), .B(new_n11685_), .ZN(new_n11686_));
  INV_X1     g11622(.I(new_n11686_), .ZN(new_n11687_));
  NAND2_X1   g11623(.A1(new_n11459_), .A2(new_n11472_), .ZN(new_n11688_));
  AOI21_X1   g11624(.A1(new_n11687_), .A2(new_n11688_), .B(new_n11473_), .ZN(new_n11689_));
  INV_X1     g11625(.I(new_n11336_), .ZN(new_n11690_));
  OAI21_X1   g11626(.A1(new_n11690_), .A2(new_n11455_), .B(new_n11457_), .ZN(new_n11691_));
  OAI21_X1   g11627(.A1(new_n11359_), .A2(new_n11373_), .B(new_n11372_), .ZN(new_n11692_));
  INV_X1     g11628(.I(new_n11692_), .ZN(new_n11693_));
  NOR2_X1    g11629(.A1(new_n11466_), .A2(new_n11461_), .ZN(new_n11694_));
  XOR2_X1    g11630(.A1(new_n11369_), .A2(new_n11694_), .Z(new_n11695_));
  NOR2_X1    g11631(.A1(new_n11693_), .A2(new_n11695_), .ZN(new_n11696_));
  INV_X1     g11632(.I(new_n11694_), .ZN(new_n11697_));
  XOR2_X1    g11633(.A1(new_n11369_), .A2(new_n11697_), .Z(new_n11698_));
  NOR2_X1    g11634(.A1(new_n11692_), .A2(new_n11698_), .ZN(new_n11699_));
  OR2_X2     g11635(.A1(new_n11696_), .A2(new_n11699_), .Z(new_n11700_));
  OAI22_X1   g11636(.A1(new_n11353_), .A2(new_n3268_), .B1(new_n3318_), .B2(new_n11697_), .ZN(new_n11701_));
  NAND2_X1   g11637(.A1(new_n11370_), .A2(new_n3323_), .ZN(new_n11702_));
  AOI21_X1   g11638(.A1(new_n11702_), .A2(new_n11701_), .B(new_n3260_), .ZN(new_n11703_));
  NAND2_X1   g11639(.A1(new_n11700_), .A2(new_n11703_), .ZN(new_n11704_));
  XOR2_X1    g11640(.A1(new_n11704_), .A2(\a[26] ), .Z(new_n11705_));
  INV_X1     g11641(.I(new_n11252_), .ZN(new_n11706_));
  OAI21_X1   g11642(.A1(new_n341_), .A2(new_n11250_), .B(new_n11237_), .ZN(new_n11707_));
  INV_X1     g11643(.I(new_n11655_), .ZN(new_n11708_));
  NOR3_X1    g11644(.A1(new_n11469_), .A2(new_n3301_), .A3(new_n5291_), .ZN(new_n11709_));
  NOR2_X1    g11645(.A1(new_n11709_), .A2(new_n84_), .ZN(new_n11710_));
  INV_X1     g11646(.I(new_n11709_), .ZN(new_n11711_));
  NAND2_X1   g11647(.A1(new_n11226_), .A2(new_n11711_), .ZN(new_n11712_));
  AOI22_X1   g11648(.A1(new_n11712_), .A2(new_n84_), .B1(new_n11226_), .B2(new_n11710_), .ZN(new_n11713_));
  NOR4_X1    g11649(.A1(new_n640_), .A2(new_n286_), .A3(new_n475_), .A4(new_n397_), .ZN(new_n11714_));
  NAND4_X1   g11650(.A1(new_n4930_), .A2(new_n221_), .A3(new_n2307_), .A4(new_n564_), .ZN(new_n11715_));
  OR2_X2     g11651(.A1(new_n11715_), .A2(new_n11714_), .Z(new_n11716_));
  NAND4_X1   g11652(.A1(new_n1256_), .A2(new_n425_), .A3(new_n575_), .A4(new_n2942_), .ZN(new_n11717_));
  NOR4_X1    g11653(.A1(new_n3666_), .A2(new_n11716_), .A3(new_n2579_), .A4(new_n11717_), .ZN(new_n11718_));
  NOR4_X1    g11654(.A1(new_n555_), .A2(new_n2396_), .A3(new_n294_), .A4(new_n681_), .ZN(new_n11719_));
  NOR4_X1    g11655(.A1(new_n1355_), .A2(new_n365_), .A3(new_n235_), .A4(new_n256_), .ZN(new_n11720_));
  INV_X1     g11656(.I(new_n11720_), .ZN(new_n11721_));
  NAND4_X1   g11657(.A1(new_n11719_), .A2(new_n839_), .A3(new_n11721_), .A4(new_n11575_), .ZN(new_n11722_));
  INV_X1     g11658(.I(new_n11722_), .ZN(new_n11723_));
  NAND4_X1   g11659(.A1(new_n1263_), .A2(new_n1497_), .A3(new_n1044_), .A4(new_n1390_), .ZN(new_n11724_));
  NOR3_X1    g11660(.A1(new_n898_), .A2(new_n388_), .A3(new_n689_), .ZN(new_n11725_));
  NAND4_X1   g11661(.A1(new_n11725_), .A2(new_n243_), .A3(new_n685_), .A4(new_n840_), .ZN(new_n11726_));
  NOR3_X1    g11662(.A1(new_n465_), .A2(new_n106_), .A3(new_n1175_), .ZN(new_n11727_));
  INV_X1     g11663(.I(new_n11727_), .ZN(new_n11728_));
  NOR4_X1    g11664(.A1(new_n11726_), .A2(new_n11724_), .A3(new_n1683_), .A4(new_n11728_), .ZN(new_n11729_));
  NAND4_X1   g11665(.A1(new_n11718_), .A2(new_n11515_), .A3(new_n11723_), .A4(new_n11729_), .ZN(new_n11730_));
  NAND2_X1   g11666(.A1(new_n11730_), .A2(new_n11250_), .ZN(new_n11731_));
  NOR2_X1    g11667(.A1(new_n11730_), .A2(new_n11250_), .ZN(new_n11732_));
  INV_X1     g11668(.I(new_n11732_), .ZN(new_n11733_));
  AOI21_X1   g11669(.A1(new_n11731_), .A2(new_n11733_), .B(new_n11713_), .ZN(new_n11734_));
  XNOR2_X1   g11670(.A1(new_n11730_), .A2(new_n11250_), .ZN(new_n11735_));
  INV_X1     g11671(.I(new_n11735_), .ZN(new_n11736_));
  AOI21_X1   g11672(.A1(new_n11713_), .A2(new_n11736_), .B(new_n11734_), .ZN(new_n11737_));
  NOR2_X1    g11673(.A1(new_n11284_), .A2(new_n2767_), .ZN(new_n11738_));
  NOR2_X1    g11674(.A1(new_n11271_), .A2(new_n2772_), .ZN(new_n11739_));
  NOR2_X1    g11675(.A1(new_n8661_), .A2(new_n2771_), .ZN(new_n11740_));
  NOR4_X1    g11676(.A1(new_n11738_), .A2(new_n2764_), .A3(new_n11739_), .A4(new_n11740_), .ZN(new_n11741_));
  AOI21_X1   g11677(.A1(new_n11708_), .A2(new_n11741_), .B(new_n11737_), .ZN(new_n11742_));
  INV_X1     g11678(.I(new_n11742_), .ZN(new_n11743_));
  INV_X1     g11679(.I(new_n11737_), .ZN(new_n11744_));
  NAND2_X1   g11680(.A1(new_n11708_), .A2(new_n11741_), .ZN(new_n11745_));
  NOR2_X1    g11681(.A1(new_n11745_), .A2(new_n11744_), .ZN(new_n11746_));
  INV_X1     g11682(.I(new_n11746_), .ZN(new_n11747_));
  AOI22_X1   g11683(.A1(new_n11743_), .A2(new_n11747_), .B1(new_n11706_), .B2(new_n11707_), .ZN(new_n11748_));
  NAND2_X1   g11684(.A1(new_n11707_), .A2(new_n11706_), .ZN(new_n11749_));
  XOR2_X1    g11685(.A1(new_n11745_), .A2(new_n11737_), .Z(new_n11750_));
  NOR2_X1    g11686(.A1(new_n11750_), .A2(new_n11749_), .ZN(new_n11751_));
  NOR2_X1    g11687(.A1(new_n11751_), .A2(new_n11748_), .ZN(new_n11752_));
  OAI21_X1   g11688(.A1(new_n11258_), .A2(new_n11332_), .B(new_n11334_), .ZN(new_n11753_));
  XOR2_X1    g11689(.A1(new_n11264_), .A2(new_n11346_), .Z(new_n11754_));
  XOR2_X1    g11690(.A1(new_n11264_), .A2(new_n11346_), .Z(new_n11755_));
  NAND2_X1   g11691(.A1(new_n11339_), .A2(new_n11755_), .ZN(new_n11756_));
  OAI21_X1   g11692(.A1(new_n11339_), .A2(new_n11754_), .B(new_n11756_), .ZN(new_n11757_));
  OAI22_X1   g11693(.A1(new_n11264_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n11277_), .ZN(new_n11758_));
  NAND2_X1   g11694(.A1(new_n11346_), .A2(new_n2750_), .ZN(new_n11759_));
  AOI21_X1   g11695(.A1(new_n11758_), .A2(new_n11759_), .B(new_n2737_), .ZN(new_n11760_));
  NAND2_X1   g11696(.A1(new_n11757_), .A2(new_n11760_), .ZN(new_n11761_));
  XOR2_X1    g11697(.A1(new_n11761_), .A2(\a[29] ), .Z(new_n11762_));
  INV_X1     g11698(.I(new_n11762_), .ZN(new_n11763_));
  NOR2_X1    g11699(.A1(new_n11753_), .A2(new_n11763_), .ZN(new_n11764_));
  INV_X1     g11700(.I(new_n11764_), .ZN(new_n11765_));
  NAND2_X1   g11701(.A1(new_n11753_), .A2(new_n11763_), .ZN(new_n11766_));
  AOI21_X1   g11702(.A1(new_n11765_), .A2(new_n11766_), .B(new_n11752_), .ZN(new_n11767_));
  XOR2_X1    g11703(.A1(new_n11753_), .A2(new_n11762_), .Z(new_n11768_));
  NOR3_X1    g11704(.A1(new_n11768_), .A2(new_n11748_), .A3(new_n11751_), .ZN(new_n11769_));
  NOR2_X1    g11705(.A1(new_n11769_), .A2(new_n11767_), .ZN(new_n11770_));
  AND2_X2    g11706(.A1(new_n11770_), .A2(new_n11705_), .Z(new_n11771_));
  NOR2_X1    g11707(.A1(new_n11770_), .A2(new_n11705_), .ZN(new_n11772_));
  OAI21_X1   g11708(.A1(new_n11771_), .A2(new_n11772_), .B(new_n11691_), .ZN(new_n11773_));
  INV_X1     g11709(.I(new_n11691_), .ZN(new_n11774_));
  XOR2_X1    g11710(.A1(new_n11770_), .A2(new_n11705_), .Z(new_n11775_));
  NAND2_X1   g11711(.A1(new_n11775_), .A2(new_n11774_), .ZN(new_n11776_));
  NAND2_X1   g11712(.A1(new_n11776_), .A2(new_n11773_), .ZN(new_n11777_));
  NOR2_X1    g11713(.A1(new_n6924_), .A2(\a[2] ), .ZN(new_n11778_));
  NOR2_X1    g11714(.A1(new_n11778_), .A2(new_n4387_), .ZN(new_n11779_));
  NAND2_X1   g11715(.A1(new_n11226_), .A2(new_n11779_), .ZN(new_n11780_));
  OAI21_X1   g11716(.A1(new_n11461_), .A2(new_n6923_), .B(new_n4387_), .ZN(new_n11781_));
  NAND2_X1   g11717(.A1(new_n11781_), .A2(new_n11780_), .ZN(new_n11782_));
  INV_X1     g11718(.I(new_n11779_), .ZN(new_n11783_));
  NOR2_X1    g11719(.A1(new_n11461_), .A2(new_n11783_), .ZN(new_n11784_));
  AOI21_X1   g11720(.A1(new_n11226_), .A2(new_n6924_), .B(\a[2] ), .ZN(new_n11785_));
  NAND3_X1   g11721(.A1(new_n10865_), .A2(new_n8778_), .A3(new_n8785_), .ZN(new_n11786_));
  INV_X1     g11722(.I(new_n11786_), .ZN(new_n11787_));
  NAND2_X1   g11723(.A1(new_n10875_), .A2(new_n8784_), .ZN(new_n11788_));
  NAND2_X1   g11724(.A1(new_n10865_), .A2(new_n8785_), .ZN(new_n11789_));
  INV_X1     g11725(.I(new_n11789_), .ZN(new_n11790_));
  NOR2_X1    g11726(.A1(new_n11788_), .A2(new_n8778_), .ZN(new_n11791_));
  OAI21_X1   g11727(.A1(new_n11791_), .A2(new_n11787_), .B(new_n10872_), .ZN(new_n11792_));
  OAI21_X1   g11728(.A1(new_n10876_), .A2(new_n10866_), .B(new_n10871_), .ZN(new_n11793_));
  NAND2_X1   g11729(.A1(new_n11792_), .A2(new_n11793_), .ZN(new_n11794_));
  NAND2_X1   g11730(.A1(new_n10872_), .A2(new_n3332_), .ZN(new_n11795_));
  NAND2_X1   g11731(.A1(new_n8779_), .A2(new_n3189_), .ZN(new_n11796_));
  AOI21_X1   g11732(.A1(new_n8785_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n11797_));
  NAND4_X1   g11733(.A1(new_n11794_), .A2(new_n11795_), .A3(new_n11796_), .A4(new_n11797_), .ZN(new_n11798_));
  INV_X1     g11734(.I(new_n2299_), .ZN(new_n11799_));
  NOR3_X1    g11735(.A1(new_n1289_), .A2(new_n850_), .A3(new_n1620_), .ZN(new_n11800_));
  NOR3_X1    g11736(.A1(new_n607_), .A2(new_n1084_), .A3(new_n910_), .ZN(new_n11801_));
  INV_X1     g11737(.I(new_n11801_), .ZN(new_n11802_));
  NOR4_X1    g11738(.A1(new_n1984_), .A2(new_n294_), .A3(new_n574_), .A4(new_n70_), .ZN(new_n11803_));
  NOR4_X1    g11739(.A1(new_n3876_), .A2(new_n11802_), .A3(new_n2859_), .A4(new_n11803_), .ZN(new_n11804_));
  NOR4_X1    g11740(.A1(new_n1433_), .A2(new_n2065_), .A3(new_n238_), .A4(new_n463_), .ZN(new_n11805_));
  NAND4_X1   g11741(.A1(new_n11805_), .A2(new_n207_), .A3(new_n1395_), .A4(new_n451_), .ZN(new_n11806_));
  INV_X1     g11742(.I(new_n11806_), .ZN(new_n11807_));
  NAND4_X1   g11743(.A1(new_n11807_), .A2(new_n11799_), .A3(new_n11800_), .A4(new_n11804_), .ZN(new_n11808_));
  NOR2_X1    g11744(.A1(new_n415_), .A2(new_n487_), .ZN(new_n11809_));
  NAND4_X1   g11745(.A1(new_n11809_), .A2(new_n662_), .A3(new_n204_), .A4(new_n2269_), .ZN(new_n11810_));
  NOR2_X1    g11746(.A1(new_n11808_), .A2(new_n11810_), .ZN(new_n11811_));
  NAND4_X1   g11747(.A1(new_n978_), .A2(new_n1725_), .A3(new_n655_), .A4(new_n250_), .ZN(new_n11812_));
  NOR2_X1    g11748(.A1(new_n381_), .A2(new_n172_), .ZN(new_n11813_));
  NAND4_X1   g11749(.A1(new_n583_), .A2(new_n438_), .A3(new_n11812_), .A4(new_n11813_), .ZN(new_n11814_));
  NOR2_X1    g11750(.A1(new_n714_), .A2(new_n227_), .ZN(new_n11815_));
  INV_X1     g11751(.I(new_n11815_), .ZN(new_n11816_));
  NOR2_X1    g11752(.A1(new_n11816_), .A2(new_n106_), .ZN(new_n11817_));
  NOR4_X1    g11753(.A1(new_n217_), .A2(new_n640_), .A3(new_n333_), .A4(new_n1168_), .ZN(new_n11818_));
  INV_X1     g11754(.I(new_n11818_), .ZN(new_n11819_));
  NAND4_X1   g11755(.A1(new_n628_), .A2(new_n1190_), .A3(new_n1468_), .A4(new_n1557_), .ZN(new_n11820_));
  NAND4_X1   g11756(.A1(new_n1411_), .A2(new_n11817_), .A3(new_n11819_), .A4(new_n11820_), .ZN(new_n11821_));
  INV_X1     g11757(.I(new_n1991_), .ZN(new_n11822_));
  NAND3_X1   g11758(.A1(new_n1329_), .A2(new_n927_), .A3(new_n11822_), .ZN(new_n11823_));
  NOR4_X1    g11759(.A1(new_n11821_), .A2(new_n2305_), .A3(new_n11814_), .A4(new_n11823_), .ZN(new_n11824_));
  NAND3_X1   g11760(.A1(new_n11811_), .A2(new_n11412_), .A3(new_n11824_), .ZN(new_n11825_));
  NAND2_X1   g11761(.A1(new_n11798_), .A2(new_n11825_), .ZN(new_n11826_));
  OAI21_X1   g11762(.A1(new_n11785_), .A2(new_n11784_), .B(new_n11826_), .ZN(new_n11827_));
  NOR2_X1    g11763(.A1(new_n11798_), .A2(new_n11825_), .ZN(new_n11828_));
  INV_X1     g11764(.I(new_n11828_), .ZN(new_n11829_));
  NOR4_X1    g11765(.A1(new_n213_), .A2(new_n1531_), .A3(new_n648_), .A4(new_n487_), .ZN(new_n11830_));
  NAND4_X1   g11766(.A1(new_n766_), .A2(new_n2395_), .A3(new_n2521_), .A4(new_n410_), .ZN(new_n11831_));
  NAND3_X1   g11767(.A1(new_n1810_), .A2(new_n2828_), .A3(new_n911_), .ZN(new_n11832_));
  NOR4_X1    g11768(.A1(new_n11831_), .A2(new_n472_), .A3(new_n11830_), .A4(new_n11832_), .ZN(new_n11833_));
  NOR4_X1    g11769(.A1(new_n11818_), .A2(new_n866_), .A3(new_n304_), .A4(new_n1944_), .ZN(new_n11834_));
  NOR3_X1    g11770(.A1(new_n891_), .A2(new_n2234_), .A3(new_n611_), .ZN(new_n11835_));
  AND3_X2    g11771(.A1(new_n3086_), .A2(new_n11834_), .A3(new_n11835_), .Z(new_n11836_));
  NAND2_X1   g11772(.A1(new_n2024_), .A2(new_n2957_), .ZN(new_n11837_));
  NOR4_X1    g11773(.A1(new_n11837_), .A2(new_n1410_), .A3(new_n855_), .A4(new_n2092_), .ZN(new_n11838_));
  NAND4_X1   g11774(.A1(new_n11838_), .A2(new_n11836_), .A3(new_n1909_), .A4(new_n11833_), .ZN(new_n11839_));
  NAND3_X1   g11775(.A1(new_n162_), .A2(new_n11507_), .A3(new_n832_), .ZN(new_n11840_));
  NAND4_X1   g11776(.A1(new_n2835_), .A2(new_n2274_), .A3(new_n3365_), .A4(new_n1700_), .ZN(new_n11841_));
  NOR4_X1    g11777(.A1(new_n2149_), .A2(new_n1264_), .A3(new_n954_), .A4(new_n1157_), .ZN(new_n11842_));
  NOR4_X1    g11778(.A1(new_n602_), .A2(new_n2439_), .A3(new_n398_), .A4(new_n763_), .ZN(new_n11843_));
  INV_X1     g11779(.I(new_n11843_), .ZN(new_n11844_));
  NAND4_X1   g11780(.A1(new_n11842_), .A2(new_n1638_), .A3(new_n1282_), .A4(new_n11844_), .ZN(new_n11845_));
  OR3_X2     g11781(.A1(new_n11845_), .A2(new_n997_), .A3(new_n1041_), .Z(new_n11846_));
  NOR4_X1    g11782(.A1(new_n11846_), .A2(new_n323_), .A3(new_n11840_), .A4(new_n11841_), .ZN(new_n11847_));
  INV_X1     g11783(.I(new_n11847_), .ZN(new_n11848_));
  NOR2_X1    g11784(.A1(new_n11848_), .A2(new_n11839_), .ZN(new_n11849_));
  NOR3_X1    g11785(.A1(new_n11785_), .A2(new_n11784_), .A3(new_n11849_), .ZN(new_n11850_));
  AOI21_X1   g11786(.A1(new_n11827_), .A2(new_n11829_), .B(new_n11850_), .ZN(new_n11851_));
  INV_X1     g11787(.I(new_n11849_), .ZN(new_n11852_));
  AOI21_X1   g11788(.A1(new_n11781_), .A2(new_n11780_), .B(new_n11852_), .ZN(new_n11853_));
  INV_X1     g11789(.I(new_n2834_), .ZN(new_n11854_));
  NAND3_X1   g11790(.A1(new_n757_), .A2(new_n442_), .A3(new_n1212_), .ZN(new_n11855_));
  NOR2_X1    g11791(.A1(new_n906_), .A2(new_n459_), .ZN(new_n11856_));
  NAND2_X1   g11792(.A1(new_n1817_), .A2(new_n11856_), .ZN(new_n11857_));
  NOR4_X1    g11793(.A1(new_n415_), .A2(new_n261_), .A3(new_n125_), .A4(new_n594_), .ZN(new_n11858_));
  NOR4_X1    g11794(.A1(new_n945_), .A2(new_n637_), .A3(new_n239_), .A4(new_n698_), .ZN(new_n11859_));
  NOR4_X1    g11795(.A1(new_n11857_), .A2(new_n11859_), .A3(new_n11855_), .A4(new_n11858_), .ZN(new_n11860_));
  NAND4_X1   g11796(.A1(new_n2783_), .A2(new_n1182_), .A3(new_n11860_), .A4(new_n1975_), .ZN(new_n11861_));
  NOR3_X1    g11797(.A1(new_n11854_), .A2(new_n2573_), .A3(new_n11861_), .ZN(new_n11862_));
  OAI22_X1   g11798(.A1(new_n11851_), .A2(new_n11853_), .B1(new_n11782_), .B2(new_n11862_), .ZN(new_n11863_));
  INV_X1     g11799(.I(new_n11862_), .ZN(new_n11864_));
  AOI21_X1   g11800(.A1(new_n11781_), .A2(new_n11780_), .B(new_n11864_), .ZN(new_n11865_));
  INV_X1     g11801(.I(new_n11865_), .ZN(new_n11866_));
  NAND2_X1   g11802(.A1(new_n11863_), .A2(new_n11866_), .ZN(new_n11867_));
  NOR2_X1    g11803(.A1(new_n6838_), .A2(new_n8799_), .ZN(new_n11868_));
  INV_X1     g11804(.I(new_n11868_), .ZN(new_n11869_));
  NOR3_X1    g11805(.A1(new_n11869_), .A2(new_n6846_), .A3(new_n6835_), .ZN(new_n11870_));
  NOR2_X1    g11806(.A1(new_n11870_), .A2(new_n65_), .ZN(new_n11871_));
  NAND2_X1   g11807(.A1(new_n11226_), .A2(new_n11871_), .ZN(new_n11872_));
  OAI21_X1   g11808(.A1(new_n11461_), .A2(new_n11870_), .B(new_n65_), .ZN(new_n11873_));
  NAND2_X1   g11809(.A1(new_n11873_), .A2(new_n11872_), .ZN(new_n11874_));
  NOR3_X1    g11810(.A1(new_n1915_), .A2(new_n1782_), .A3(new_n198_), .ZN(new_n11875_));
  INV_X1     g11811(.I(new_n11875_), .ZN(new_n11876_));
  NOR4_X1    g11812(.A1(new_n424_), .A2(new_n261_), .A3(new_n594_), .A4(new_n817_), .ZN(new_n11877_));
  NOR4_X1    g11813(.A1(new_n732_), .A2(new_n154_), .A3(new_n376_), .A4(new_n506_), .ZN(new_n11878_));
  NOR4_X1    g11814(.A1(new_n1259_), .A2(new_n11876_), .A3(new_n11877_), .A4(new_n11878_), .ZN(new_n11879_));
  NAND4_X1   g11815(.A1(new_n1414_), .A2(new_n657_), .A3(new_n820_), .A4(new_n2810_), .ZN(new_n11880_));
  NOR4_X1    g11816(.A1(new_n86_), .A2(new_n137_), .A3(new_n531_), .A4(new_n335_), .ZN(new_n11881_));
  NOR3_X1    g11817(.A1(new_n11880_), .A2(new_n2955_), .A3(new_n11881_), .ZN(new_n11882_));
  NOR2_X1    g11818(.A1(new_n4827_), .A2(new_n4564_), .ZN(new_n11883_));
  NAND4_X1   g11819(.A1(new_n11879_), .A2(new_n2857_), .A3(new_n11882_), .A4(new_n11883_), .ZN(new_n11884_));
  NOR2_X1    g11820(.A1(new_n11884_), .A2(new_n11839_), .ZN(new_n11885_));
  NOR2_X1    g11821(.A1(new_n11874_), .A2(new_n11885_), .ZN(new_n11886_));
  INV_X1     g11822(.I(new_n11871_), .ZN(new_n11887_));
  NOR2_X1    g11823(.A1(new_n11461_), .A2(new_n11887_), .ZN(new_n11888_));
  INV_X1     g11824(.I(new_n11870_), .ZN(new_n11889_));
  AOI21_X1   g11825(.A1(new_n11226_), .A2(new_n11889_), .B(\a[5] ), .ZN(new_n11890_));
  NOR2_X1    g11826(.A1(new_n11890_), .A2(new_n11888_), .ZN(new_n11891_));
  INV_X1     g11827(.I(new_n11885_), .ZN(new_n11892_));
  NOR2_X1    g11828(.A1(new_n11891_), .A2(new_n11892_), .ZN(new_n11893_));
  OAI21_X1   g11829(.A1(new_n11893_), .A2(new_n11886_), .B(new_n11782_), .ZN(new_n11894_));
  INV_X1     g11830(.I(new_n11782_), .ZN(new_n11895_));
  NOR2_X1    g11831(.A1(new_n11891_), .A2(new_n11885_), .ZN(new_n11896_));
  NOR3_X1    g11832(.A1(new_n11890_), .A2(new_n11888_), .A3(new_n11892_), .ZN(new_n11897_));
  OAI21_X1   g11833(.A1(new_n11896_), .A2(new_n11897_), .B(new_n11895_), .ZN(new_n11898_));
  INV_X1     g11834(.I(new_n10899_), .ZN(new_n11899_));
  NAND3_X1   g11835(.A1(new_n10891_), .A2(new_n10892_), .A3(new_n10894_), .ZN(new_n11900_));
  INV_X1     g11836(.I(new_n11900_), .ZN(new_n11901_));
  AOI21_X1   g11837(.A1(new_n10891_), .A2(new_n10894_), .B(new_n10892_), .ZN(new_n11902_));
  OAI21_X1   g11838(.A1(new_n11901_), .A2(new_n11902_), .B(new_n11899_), .ZN(new_n11903_));
  OAI21_X1   g11839(.A1(new_n10910_), .A2(new_n10893_), .B(new_n10892_), .ZN(new_n11904_));
  NAND3_X1   g11840(.A1(new_n10891_), .A2(new_n10889_), .A3(new_n10894_), .ZN(new_n11905_));
  NAND2_X1   g11841(.A1(new_n11905_), .A2(new_n11904_), .ZN(new_n11906_));
  NAND2_X1   g11842(.A1(new_n11906_), .A2(new_n10899_), .ZN(new_n11907_));
  NAND2_X1   g11843(.A1(new_n11903_), .A2(new_n11907_), .ZN(new_n11908_));
  NOR2_X1    g11844(.A1(new_n10899_), .A2(new_n2772_), .ZN(new_n11909_));
  NOR2_X1    g11845(.A1(new_n10892_), .A2(new_n2767_), .ZN(new_n11910_));
  NOR2_X1    g11846(.A1(new_n10885_), .A2(new_n2771_), .ZN(new_n11911_));
  NOR4_X1    g11847(.A1(new_n11909_), .A2(new_n2764_), .A3(new_n11910_), .A4(new_n11911_), .ZN(new_n11912_));
  NAND2_X1   g11848(.A1(new_n11908_), .A2(new_n11912_), .ZN(new_n11913_));
  NAND3_X1   g11849(.A1(new_n11894_), .A2(new_n11898_), .A3(new_n11913_), .ZN(new_n11914_));
  AOI21_X1   g11850(.A1(new_n11894_), .A2(new_n11898_), .B(new_n11913_), .ZN(new_n11915_));
  AOI21_X1   g11851(.A1(new_n11867_), .A2(new_n11914_), .B(new_n11915_), .ZN(new_n11916_));
  NAND2_X1   g11852(.A1(new_n11874_), .A2(new_n11892_), .ZN(new_n11917_));
  AOI21_X1   g11853(.A1(new_n11917_), .A2(new_n11895_), .B(new_n11897_), .ZN(new_n11918_));
  NOR3_X1    g11854(.A1(new_n670_), .A2(new_n910_), .A3(new_n449_), .ZN(new_n11919_));
  NAND4_X1   g11855(.A1(new_n2125_), .A2(new_n773_), .A3(new_n1096_), .A4(new_n11919_), .ZN(new_n11920_));
  NOR4_X1    g11856(.A1(new_n11920_), .A2(new_n544_), .A3(new_n756_), .A4(new_n2930_), .ZN(new_n11921_));
  NAND2_X1   g11857(.A1(new_n246_), .A2(new_n349_), .ZN(new_n11922_));
  NOR3_X1    g11858(.A1(new_n1197_), .A2(new_n482_), .A3(new_n531_), .ZN(new_n11923_));
  NAND4_X1   g11859(.A1(new_n11923_), .A2(new_n628_), .A3(new_n790_), .A4(new_n3502_), .ZN(new_n11924_));
  NOR4_X1    g11860(.A1(new_n11924_), .A2(new_n1614_), .A3(new_n2193_), .A4(new_n11922_), .ZN(new_n11925_));
  INV_X1     g11861(.I(new_n10970_), .ZN(new_n11926_));
  NOR3_X1    g11862(.A1(new_n11926_), .A2(new_n802_), .A3(new_n2523_), .ZN(new_n11927_));
  NAND4_X1   g11863(.A1(new_n11925_), .A2(new_n3012_), .A3(new_n11921_), .A4(new_n11927_), .ZN(new_n11928_));
  NAND2_X1   g11864(.A1(new_n1601_), .A2(new_n1070_), .ZN(new_n11929_));
  NAND3_X1   g11865(.A1(new_n875_), .A2(new_n913_), .A3(new_n1805_), .ZN(new_n11930_));
  NAND2_X1   g11866(.A1(new_n3337_), .A2(new_n1296_), .ZN(new_n11931_));
  NOR4_X1    g11867(.A1(new_n11931_), .A2(new_n734_), .A3(new_n11929_), .A4(new_n11930_), .ZN(new_n11932_));
  NAND4_X1   g11868(.A1(new_n11932_), .A2(new_n931_), .A3(new_n993_), .A4(new_n2040_), .ZN(new_n11933_));
  NOR3_X1    g11869(.A1(new_n11928_), .A2(new_n11722_), .A3(new_n11933_), .ZN(new_n11934_));
  NAND2_X1   g11870(.A1(new_n11934_), .A2(new_n1676_), .ZN(new_n11935_));
  AOI21_X1   g11871(.A1(new_n10891_), .A2(new_n10894_), .B(new_n10889_), .ZN(new_n11936_));
  NOR3_X1    g11872(.A1(new_n10910_), .A2(new_n10892_), .A3(new_n10893_), .ZN(new_n11937_));
  NOR2_X1    g11873(.A1(new_n11936_), .A2(new_n11937_), .ZN(new_n11938_));
  OAI21_X1   g11874(.A1(new_n10910_), .A2(new_n10893_), .B(new_n10899_), .ZN(new_n11939_));
  NAND3_X1   g11875(.A1(new_n10891_), .A2(new_n10894_), .A3(new_n11899_), .ZN(new_n11940_));
  NAND2_X1   g11876(.A1(new_n11940_), .A2(new_n11939_), .ZN(new_n11941_));
  NOR3_X1    g11877(.A1(new_n11938_), .A2(new_n11941_), .A3(new_n10906_), .ZN(new_n11942_));
  INV_X1     g11878(.I(new_n11942_), .ZN(new_n11943_));
  OAI21_X1   g11879(.A1(new_n11938_), .A2(new_n11941_), .B(new_n10906_), .ZN(new_n11944_));
  NAND2_X1   g11880(.A1(new_n11943_), .A2(new_n11944_), .ZN(new_n11945_));
  NAND2_X1   g11881(.A1(new_n10906_), .A2(new_n3332_), .ZN(new_n11946_));
  NAND2_X1   g11882(.A1(new_n11899_), .A2(new_n3189_), .ZN(new_n11947_));
  AOI21_X1   g11883(.A1(new_n10889_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n11948_));
  NAND4_X1   g11884(.A1(new_n11945_), .A2(new_n11946_), .A3(new_n11947_), .A4(new_n11948_), .ZN(new_n11949_));
  XOR2_X1    g11885(.A1(new_n11949_), .A2(new_n11935_), .Z(new_n11950_));
  NOR2_X1    g11886(.A1(new_n11918_), .A2(new_n11950_), .ZN(new_n11951_));
  NAND3_X1   g11887(.A1(new_n11873_), .A2(new_n11872_), .A3(new_n11885_), .ZN(new_n11952_));
  OAI21_X1   g11888(.A1(new_n11896_), .A2(new_n11782_), .B(new_n11952_), .ZN(new_n11953_));
  INV_X1     g11889(.I(new_n11935_), .ZN(new_n11954_));
  NOR2_X1    g11890(.A1(new_n11949_), .A2(new_n11954_), .ZN(new_n11955_));
  INV_X1     g11891(.I(new_n11955_), .ZN(new_n11956_));
  NAND2_X1   g11892(.A1(new_n11949_), .A2(new_n11954_), .ZN(new_n11957_));
  AOI21_X1   g11893(.A1(new_n11956_), .A2(new_n11957_), .B(new_n11953_), .ZN(new_n11958_));
  AND2_X2    g11894(.A1(new_n10914_), .A2(new_n10905_), .Z(new_n11959_));
  XOR2_X1    g11895(.A1(new_n8746_), .A2(new_n8758_), .Z(new_n11960_));
  NAND2_X1   g11896(.A1(new_n8746_), .A2(new_n8761_), .ZN(new_n11961_));
  NAND2_X1   g11897(.A1(new_n11961_), .A2(new_n8759_), .ZN(new_n11962_));
  NAND2_X1   g11898(.A1(new_n11959_), .A2(new_n11962_), .ZN(new_n11963_));
  OAI21_X1   g11899(.A1(new_n11959_), .A2(new_n11960_), .B(new_n11963_), .ZN(new_n11964_));
  OAI22_X1   g11900(.A1(new_n8758_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8766_), .ZN(new_n11965_));
  NAND2_X1   g11901(.A1(new_n8746_), .A2(new_n2750_), .ZN(new_n11966_));
  AOI21_X1   g11902(.A1(new_n11966_), .A2(new_n11965_), .B(new_n2737_), .ZN(new_n11967_));
  NAND2_X1   g11903(.A1(new_n11964_), .A2(new_n11967_), .ZN(new_n11968_));
  XOR2_X1    g11904(.A1(new_n11968_), .A2(\a[29] ), .Z(new_n11969_));
  OAI21_X1   g11905(.A1(new_n11958_), .A2(new_n11951_), .B(new_n11969_), .ZN(new_n11970_));
  INV_X1     g11906(.I(new_n11970_), .ZN(new_n11971_));
  INV_X1     g11907(.I(new_n11950_), .ZN(new_n11972_));
  NAND2_X1   g11908(.A1(new_n11953_), .A2(new_n11972_), .ZN(new_n11973_));
  INV_X1     g11909(.I(new_n11957_), .ZN(new_n11974_));
  OAI21_X1   g11910(.A1(new_n11955_), .A2(new_n11974_), .B(new_n11918_), .ZN(new_n11975_));
  INV_X1     g11911(.I(new_n11969_), .ZN(new_n11976_));
  NAND3_X1   g11912(.A1(new_n11975_), .A2(new_n11973_), .A3(new_n11976_), .ZN(new_n11977_));
  OAI21_X1   g11913(.A1(new_n11971_), .A2(new_n11916_), .B(new_n11977_), .ZN(new_n11978_));
  AOI21_X1   g11914(.A1(new_n11953_), .A2(new_n11957_), .B(new_n11955_), .ZN(new_n11979_));
  NAND4_X1   g11915(.A1(new_n3935_), .A2(new_n1805_), .A3(new_n983_), .A4(new_n1712_), .ZN(new_n11980_));
  NAND4_X1   g11916(.A1(new_n922_), .A2(new_n2375_), .A3(new_n568_), .A4(new_n592_), .ZN(new_n11981_));
  NOR3_X1    g11917(.A1(new_n1206_), .A2(new_n398_), .A3(new_n459_), .ZN(new_n11982_));
  NAND2_X1   g11918(.A1(new_n11982_), .A2(new_n11981_), .ZN(new_n11983_));
  NAND4_X1   g11919(.A1(new_n575_), .A2(new_n870_), .A3(new_n1963_), .A4(new_n2012_), .ZN(new_n11984_));
  NOR4_X1    g11920(.A1(new_n11980_), .A2(new_n392_), .A3(new_n11983_), .A4(new_n11984_), .ZN(new_n11985_));
  NAND4_X1   g11921(.A1(new_n2221_), .A2(new_n1476_), .A3(new_n494_), .A4(new_n11985_), .ZN(new_n11986_));
  NAND2_X1   g11922(.A1(new_n11954_), .A2(new_n11986_), .ZN(new_n11987_));
  NOR2_X1    g11923(.A1(new_n11954_), .A2(new_n11986_), .ZN(new_n11988_));
  INV_X1     g11924(.I(new_n11988_), .ZN(new_n11989_));
  AOI21_X1   g11925(.A1(new_n11987_), .A2(new_n11989_), .B(new_n11979_), .ZN(new_n11990_));
  XOR2_X1    g11926(.A1(new_n11935_), .A2(new_n11986_), .Z(new_n11991_));
  INV_X1     g11927(.I(new_n11991_), .ZN(new_n11992_));
  NAND2_X1   g11928(.A1(new_n11979_), .A2(new_n11992_), .ZN(new_n11993_));
  INV_X1     g11929(.I(new_n11993_), .ZN(new_n11994_));
  NOR2_X1    g11930(.A1(new_n11994_), .A2(new_n11990_), .ZN(new_n11995_));
  INV_X1     g11931(.I(new_n8766_), .ZN(new_n11996_));
  OAI21_X1   g11932(.A1(new_n10913_), .A2(new_n10907_), .B(new_n11996_), .ZN(new_n11997_));
  NOR3_X1    g11933(.A1(new_n10912_), .A2(new_n10906_), .A3(new_n10902_), .ZN(new_n11998_));
  AOI21_X1   g11934(.A1(new_n10901_), .A2(new_n10903_), .B(new_n8774_), .ZN(new_n11999_));
  OAI21_X1   g11935(.A1(new_n11998_), .A2(new_n11999_), .B(new_n8766_), .ZN(new_n12000_));
  NAND2_X1   g11936(.A1(new_n11997_), .A2(new_n12000_), .ZN(new_n12001_));
  INV_X1     g11937(.I(new_n12001_), .ZN(new_n12002_));
  NOR2_X1    g11938(.A1(new_n8766_), .A2(new_n2772_), .ZN(new_n12003_));
  NOR2_X1    g11939(.A1(new_n8774_), .A2(new_n2767_), .ZN(new_n12004_));
  OAI21_X1   g11940(.A1(new_n10899_), .A2(new_n2771_), .B(new_n2764_), .ZN(new_n12005_));
  NOR4_X1    g11941(.A1(new_n12002_), .A2(new_n12003_), .A3(new_n12004_), .A4(new_n12005_), .ZN(new_n12006_));
  INV_X1     g11942(.I(new_n12006_), .ZN(new_n12007_));
  NAND2_X1   g11943(.A1(new_n11995_), .A2(new_n12007_), .ZN(new_n12008_));
  OAI21_X1   g11944(.A1(new_n11994_), .A2(new_n11990_), .B(new_n12006_), .ZN(new_n12009_));
  INV_X1     g11945(.I(new_n12009_), .ZN(new_n12010_));
  AOI21_X1   g11946(.A1(new_n11978_), .A2(new_n12008_), .B(new_n12010_), .ZN(new_n12011_));
  INV_X1     g11947(.I(new_n12011_), .ZN(new_n12012_));
  NAND2_X1   g11948(.A1(new_n11953_), .A2(new_n11957_), .ZN(new_n12013_));
  NAND2_X1   g11949(.A1(new_n12013_), .A2(new_n11956_), .ZN(new_n12014_));
  NAND2_X1   g11950(.A1(new_n12014_), .A2(new_n11987_), .ZN(new_n12015_));
  NAND2_X1   g11951(.A1(new_n6785_), .A2(new_n6788_), .ZN(new_n12016_));
  NOR3_X1    g11952(.A1(new_n12016_), .A2(new_n6775_), .A3(new_n7530_), .ZN(new_n12017_));
  NOR2_X1    g11953(.A1(new_n12017_), .A2(new_n4009_), .ZN(new_n12018_));
  INV_X1     g11954(.I(new_n12018_), .ZN(new_n12019_));
  NOR2_X1    g11955(.A1(new_n11461_), .A2(new_n12019_), .ZN(new_n12020_));
  INV_X1     g11956(.I(new_n12017_), .ZN(new_n12021_));
  AOI21_X1   g11957(.A1(new_n11226_), .A2(new_n12021_), .B(\a[8] ), .ZN(new_n12022_));
  NOR2_X1    g11958(.A1(new_n12022_), .A2(new_n12020_), .ZN(new_n12023_));
  NAND2_X1   g11959(.A1(new_n2406_), .A2(new_n2393_), .ZN(new_n12024_));
  NAND4_X1   g11960(.A1(new_n3676_), .A2(new_n1311_), .A3(new_n1446_), .A4(new_n501_), .ZN(new_n12025_));
  NOR2_X1    g11961(.A1(new_n1915_), .A2(new_n1053_), .ZN(new_n12026_));
  NAND4_X1   g11962(.A1(new_n2265_), .A2(new_n2181_), .A3(new_n12025_), .A4(new_n12026_), .ZN(new_n12027_));
  INV_X1     g11963(.I(new_n3840_), .ZN(new_n12028_));
  NAND4_X1   g11964(.A1(new_n1164_), .A2(new_n1489_), .A3(new_n1327_), .A4(new_n1174_), .ZN(new_n12029_));
  NOR4_X1    g11965(.A1(new_n593_), .A2(new_n225_), .A3(new_n752_), .A4(new_n560_), .ZN(new_n12030_));
  NOR3_X1    g11966(.A1(new_n12029_), .A2(new_n12028_), .A3(new_n12030_), .ZN(new_n12031_));
  NAND3_X1   g11967(.A1(new_n3502_), .A2(new_n843_), .A3(new_n1009_), .ZN(new_n12032_));
  NOR4_X1    g11968(.A1(new_n298_), .A2(new_n596_), .A3(new_n719_), .A4(new_n902_), .ZN(new_n12033_));
  NOR2_X1    g11969(.A1(new_n12032_), .A2(new_n12033_), .ZN(new_n12034_));
  INV_X1     g11970(.I(new_n852_), .ZN(new_n12035_));
  NOR3_X1    g11971(.A1(new_n12035_), .A2(new_n1656_), .A3(new_n2270_), .ZN(new_n12036_));
  NAND4_X1   g11972(.A1(new_n12031_), .A2(new_n1505_), .A3(new_n12034_), .A4(new_n12036_), .ZN(new_n12037_));
  OR4_X2     g11973(.A1(new_n12024_), .A2(new_n3206_), .A3(new_n12027_), .A4(new_n12037_), .Z(new_n12038_));
  NOR2_X1    g11974(.A1(new_n11935_), .A2(new_n12038_), .ZN(new_n12039_));
  INV_X1     g11975(.I(new_n12039_), .ZN(new_n12040_));
  NAND2_X1   g11976(.A1(new_n11935_), .A2(new_n12038_), .ZN(new_n12041_));
  AOI21_X1   g11977(.A1(new_n12040_), .A2(new_n12041_), .B(new_n12023_), .ZN(new_n12042_));
  XNOR2_X1   g11978(.A1(new_n11935_), .A2(new_n12038_), .ZN(new_n12043_));
  INV_X1     g11979(.I(new_n12043_), .ZN(new_n12044_));
  AOI21_X1   g11980(.A1(new_n12023_), .A2(new_n12044_), .B(new_n12042_), .ZN(new_n12045_));
  NOR3_X1    g11981(.A1(new_n10904_), .A2(new_n11996_), .A3(new_n8774_), .ZN(new_n12046_));
  OAI21_X1   g11982(.A1(new_n10912_), .A2(new_n10902_), .B(new_n8774_), .ZN(new_n12047_));
  NOR2_X1    g11983(.A1(new_n12047_), .A2(new_n8766_), .ZN(new_n12048_));
  OAI21_X1   g11984(.A1(new_n12048_), .A2(new_n12046_), .B(new_n8761_), .ZN(new_n12049_));
  INV_X1     g11985(.I(new_n10905_), .ZN(new_n12050_));
  NOR2_X1    g11986(.A1(new_n10907_), .A2(new_n8766_), .ZN(new_n12051_));
  OAI21_X1   g11987(.A1(new_n12050_), .A2(new_n12051_), .B(new_n8758_), .ZN(new_n12052_));
  NAND2_X1   g11988(.A1(new_n12052_), .A2(new_n12049_), .ZN(new_n12053_));
  NOR2_X1    g11989(.A1(new_n8758_), .A2(new_n2772_), .ZN(new_n12054_));
  NOR2_X1    g11990(.A1(new_n8766_), .A2(new_n2767_), .ZN(new_n12055_));
  NOR2_X1    g11991(.A1(new_n8774_), .A2(new_n2771_), .ZN(new_n12056_));
  NOR4_X1    g11992(.A1(new_n12054_), .A2(new_n2764_), .A3(new_n12056_), .A4(new_n12055_), .ZN(new_n12057_));
  NAND2_X1   g11993(.A1(new_n12053_), .A2(new_n12057_), .ZN(new_n12058_));
  INV_X1     g11994(.I(new_n12058_), .ZN(new_n12059_));
  NOR2_X1    g11995(.A1(new_n12045_), .A2(new_n12059_), .ZN(new_n12060_));
  INV_X1     g11996(.I(new_n12060_), .ZN(new_n12061_));
  NAND2_X1   g11997(.A1(new_n12045_), .A2(new_n12059_), .ZN(new_n12062_));
  AOI22_X1   g11998(.A1(new_n12015_), .A2(new_n11989_), .B1(new_n12061_), .B2(new_n12062_), .ZN(new_n12063_));
  INV_X1     g11999(.I(new_n11987_), .ZN(new_n12064_));
  OAI21_X1   g12000(.A1(new_n11979_), .A2(new_n12064_), .B(new_n11989_), .ZN(new_n12065_));
  XOR2_X1    g12001(.A1(new_n12045_), .A2(new_n12058_), .Z(new_n12066_));
  NOR2_X1    g12002(.A1(new_n12066_), .A2(new_n12065_), .ZN(new_n12067_));
  NOR2_X1    g12003(.A1(new_n12063_), .A2(new_n12067_), .ZN(new_n12068_));
  XOR2_X1    g12004(.A1(new_n8751_), .A2(new_n10927_), .Z(new_n12069_));
  XOR2_X1    g12005(.A1(new_n8751_), .A2(new_n10927_), .Z(new_n12070_));
  NAND2_X1   g12006(.A1(new_n10919_), .A2(new_n12070_), .ZN(new_n12071_));
  OAI21_X1   g12007(.A1(new_n10919_), .A2(new_n12069_), .B(new_n12071_), .ZN(new_n12072_));
  OAI22_X1   g12008(.A1(new_n8751_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8745_), .ZN(new_n12073_));
  NAND2_X1   g12009(.A1(new_n10927_), .A2(new_n2750_), .ZN(new_n12074_));
  AOI21_X1   g12010(.A1(new_n12073_), .A2(new_n12074_), .B(new_n2737_), .ZN(new_n12075_));
  NAND2_X1   g12011(.A1(new_n12072_), .A2(new_n12075_), .ZN(new_n12076_));
  XOR2_X1    g12012(.A1(new_n12076_), .A2(\a[29] ), .Z(new_n12077_));
  NAND2_X1   g12013(.A1(new_n12068_), .A2(new_n12077_), .ZN(new_n12078_));
  NOR2_X1    g12014(.A1(new_n12068_), .A2(new_n12077_), .ZN(new_n12079_));
  AOI21_X1   g12015(.A1(new_n12012_), .A2(new_n12078_), .B(new_n12079_), .ZN(new_n12080_));
  INV_X1     g12016(.I(new_n12080_), .ZN(new_n12081_));
  NAND2_X1   g12017(.A1(new_n12061_), .A2(new_n12065_), .ZN(new_n12082_));
  NAND2_X1   g12018(.A1(new_n12082_), .A2(new_n12062_), .ZN(new_n12083_));
  NAND2_X1   g12019(.A1(new_n12023_), .A2(new_n12041_), .ZN(new_n12084_));
  NAND2_X1   g12020(.A1(new_n12084_), .A2(new_n12040_), .ZN(new_n12085_));
  INV_X1     g12021(.I(new_n11879_), .ZN(new_n12086_));
  NAND4_X1   g12022(.A1(new_n667_), .A2(new_n1221_), .A3(new_n1446_), .A4(new_n808_), .ZN(new_n12087_));
  NAND4_X1   g12023(.A1(new_n451_), .A2(new_n568_), .A3(new_n1396_), .A4(new_n672_), .ZN(new_n12088_));
  NAND4_X1   g12024(.A1(new_n12087_), .A2(new_n2167_), .A3(new_n11056_), .A4(new_n12088_), .ZN(new_n12089_));
  NOR2_X1    g12025(.A1(new_n541_), .A2(new_n574_), .ZN(new_n12090_));
  NAND4_X1   g12026(.A1(new_n12090_), .A2(new_n3868_), .A3(new_n93_), .A4(new_n1395_), .ZN(new_n12091_));
  NOR2_X1    g12027(.A1(new_n2582_), .A2(new_n1365_), .ZN(new_n12092_));
  NAND4_X1   g12028(.A1(new_n3342_), .A2(new_n1575_), .A3(new_n12092_), .A4(new_n1767_), .ZN(new_n12093_));
  NOR4_X1    g12029(.A1(new_n12086_), .A2(new_n12089_), .A3(new_n12091_), .A4(new_n12093_), .ZN(new_n12094_));
  NOR2_X1    g12030(.A1(new_n4558_), .A2(new_n1966_), .ZN(new_n12095_));
  NAND2_X1   g12031(.A1(new_n12094_), .A2(new_n12095_), .ZN(new_n12096_));
  NAND2_X1   g12032(.A1(new_n8746_), .A2(new_n3332_), .ZN(new_n12097_));
  NAND2_X1   g12033(.A1(new_n8761_), .A2(new_n3189_), .ZN(new_n12098_));
  AOI21_X1   g12034(.A1(new_n11996_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n12099_));
  NAND4_X1   g12035(.A1(new_n11964_), .A2(new_n12097_), .A3(new_n12098_), .A4(new_n12099_), .ZN(new_n12100_));
  XOR2_X1    g12036(.A1(new_n12100_), .A2(new_n12096_), .Z(new_n12101_));
  INV_X1     g12037(.I(new_n12101_), .ZN(new_n12102_));
  INV_X1     g12038(.I(new_n12096_), .ZN(new_n12103_));
  NAND2_X1   g12039(.A1(new_n12100_), .A2(new_n12103_), .ZN(new_n12104_));
  NOR2_X1    g12040(.A1(new_n12100_), .A2(new_n12103_), .ZN(new_n12105_));
  INV_X1     g12041(.I(new_n12105_), .ZN(new_n12106_));
  AOI21_X1   g12042(.A1(new_n12104_), .A2(new_n12106_), .B(new_n12085_), .ZN(new_n12107_));
  AOI21_X1   g12043(.A1(new_n12085_), .A2(new_n12102_), .B(new_n12107_), .ZN(new_n12108_));
  INV_X1     g12044(.I(new_n8753_), .ZN(new_n12109_));
  OAI22_X1   g12045(.A1(new_n10915_), .A2(new_n8760_), .B1(new_n8745_), .B2(new_n8751_), .ZN(new_n12110_));
  AOI21_X1   g12046(.A1(new_n12110_), .A2(new_n12109_), .B(new_n10927_), .ZN(new_n12111_));
  INV_X1     g12047(.I(new_n12069_), .ZN(new_n12112_));
  NAND3_X1   g12048(.A1(new_n12110_), .A2(new_n12109_), .A3(new_n10927_), .ZN(new_n12113_));
  NAND2_X1   g12049(.A1(new_n12113_), .A2(new_n12112_), .ZN(new_n12114_));
  NOR3_X1    g12050(.A1(new_n12114_), .A2(new_n8736_), .A3(new_n12111_), .ZN(new_n12115_));
  OAI21_X1   g12051(.A1(new_n12114_), .A2(new_n12111_), .B(new_n8736_), .ZN(new_n12116_));
  INV_X1     g12052(.I(new_n12116_), .ZN(new_n12117_));
  NOR2_X1    g12053(.A1(new_n12117_), .A2(new_n12115_), .ZN(new_n12118_));
  OAI22_X1   g12054(.A1(new_n8751_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n10924_), .ZN(new_n12119_));
  NAND2_X1   g12055(.A1(new_n8736_), .A2(new_n2750_), .ZN(new_n12120_));
  AOI21_X1   g12056(.A1(new_n12120_), .A2(new_n12119_), .B(new_n2737_), .ZN(new_n12121_));
  NAND2_X1   g12057(.A1(new_n12118_), .A2(new_n12121_), .ZN(new_n12122_));
  XOR2_X1    g12058(.A1(new_n12122_), .A2(\a[29] ), .Z(new_n12123_));
  XOR2_X1    g12059(.A1(new_n12108_), .A2(new_n12123_), .Z(new_n12124_));
  INV_X1     g12060(.I(new_n12124_), .ZN(new_n12125_));
  INV_X1     g12061(.I(new_n12108_), .ZN(new_n12126_));
  NAND2_X1   g12062(.A1(new_n12126_), .A2(new_n12123_), .ZN(new_n12127_));
  NOR2_X1    g12063(.A1(new_n12126_), .A2(new_n12123_), .ZN(new_n12128_));
  INV_X1     g12064(.I(new_n12128_), .ZN(new_n12129_));
  AOI21_X1   g12065(.A1(new_n12129_), .A2(new_n12127_), .B(new_n12083_), .ZN(new_n12130_));
  AOI21_X1   g12066(.A1(new_n12083_), .A2(new_n12125_), .B(new_n12130_), .ZN(new_n12131_));
  OAI22_X1   g12067(.A1(new_n8725_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n8718_), .ZN(new_n12132_));
  NAND2_X1   g12068(.A1(new_n8711_), .A2(new_n3317_), .ZN(new_n12133_));
  AOI21_X1   g12069(.A1(new_n12133_), .A2(new_n12132_), .B(new_n3260_), .ZN(new_n12134_));
  NAND2_X1   g12070(.A1(new_n11536_), .A2(new_n12134_), .ZN(new_n12135_));
  XOR2_X1    g12071(.A1(new_n12135_), .A2(\a[26] ), .Z(new_n12136_));
  INV_X1     g12072(.I(new_n12136_), .ZN(new_n12137_));
  NOR2_X1    g12073(.A1(new_n12131_), .A2(new_n12137_), .ZN(new_n12138_));
  INV_X1     g12074(.I(new_n12138_), .ZN(new_n12139_));
  NAND2_X1   g12075(.A1(new_n12131_), .A2(new_n12137_), .ZN(new_n12140_));
  INV_X1     g12076(.I(new_n12140_), .ZN(new_n12141_));
  AOI21_X1   g12077(.A1(new_n12081_), .A2(new_n12139_), .B(new_n12141_), .ZN(new_n12142_));
  INV_X1     g12078(.I(new_n12142_), .ZN(new_n12143_));
  NAND2_X1   g12079(.A1(new_n12083_), .A2(new_n12127_), .ZN(new_n12144_));
  AOI21_X1   g12080(.A1(new_n12085_), .A2(new_n12104_), .B(new_n12105_), .ZN(new_n12145_));
  NAND3_X1   g12081(.A1(new_n1319_), .A2(new_n1816_), .A3(new_n1096_), .ZN(new_n12146_));
  NAND2_X1   g12082(.A1(new_n1354_), .A2(new_n476_), .ZN(new_n12147_));
  NAND3_X1   g12083(.A1(new_n1395_), .A2(new_n1327_), .A3(new_n761_), .ZN(new_n12148_));
  NOR4_X1    g12084(.A1(new_n12147_), .A2(new_n12146_), .A3(new_n11818_), .A4(new_n12148_), .ZN(new_n12149_));
  NAND2_X1   g12085(.A1(new_n1256_), .A2(new_n399_), .ZN(new_n12150_));
  NOR4_X1    g12086(.A1(new_n514_), .A2(new_n12150_), .A3(new_n200_), .A4(new_n1341_), .ZN(new_n12151_));
  NOR4_X1    g12087(.A1(new_n958_), .A2(new_n534_), .A3(new_n256_), .A4(new_n633_), .ZN(new_n12152_));
  INV_X1     g12088(.I(new_n12152_), .ZN(new_n12153_));
  NOR2_X1    g12089(.A1(new_n12153_), .A2(new_n1936_), .ZN(new_n12154_));
  NAND3_X1   g12090(.A1(new_n12154_), .A2(new_n12149_), .A3(new_n12151_), .ZN(new_n12155_));
  NOR2_X1    g12091(.A1(new_n12155_), .A2(new_n1464_), .ZN(new_n12156_));
  NAND3_X1   g12092(.A1(new_n2038_), .A2(new_n1237_), .A3(new_n1126_), .ZN(new_n12157_));
  NOR3_X1    g12093(.A1(new_n1382_), .A2(new_n264_), .A3(new_n459_), .ZN(new_n12158_));
  NOR3_X1    g12094(.A1(new_n117_), .A2(new_n485_), .A3(new_n376_), .ZN(new_n12159_));
  INV_X1     g12095(.I(new_n12159_), .ZN(new_n12160_));
  NOR3_X1    g12096(.A1(new_n12157_), .A2(new_n12158_), .A3(new_n12160_), .ZN(new_n12161_));
  INV_X1     g12097(.I(new_n12161_), .ZN(new_n12162_));
  NOR4_X1    g12098(.A1(new_n1137_), .A2(new_n523_), .A3(new_n935_), .A4(new_n1954_), .ZN(new_n12163_));
  INV_X1     g12099(.I(new_n2346_), .ZN(new_n12164_));
  NOR4_X1    g12100(.A1(new_n12164_), .A2(new_n137_), .A3(new_n866_), .A4(new_n2677_), .ZN(new_n12165_));
  NOR2_X1    g12101(.A1(new_n127_), .A2(new_n825_), .ZN(new_n12166_));
  NAND4_X1   g12102(.A1(new_n675_), .A2(new_n1805_), .A3(new_n319_), .A4(new_n1491_), .ZN(new_n12167_));
  NAND4_X1   g12103(.A1(new_n12165_), .A2(new_n12163_), .A3(new_n12166_), .A4(new_n12167_), .ZN(new_n12168_));
  NOR3_X1    g12104(.A1(new_n12168_), .A2(new_n3433_), .A3(new_n12162_), .ZN(new_n12169_));
  AOI21_X1   g12105(.A1(new_n12156_), .A2(new_n12169_), .B(new_n12096_), .ZN(new_n12170_));
  NAND2_X1   g12106(.A1(new_n12169_), .A2(new_n12156_), .ZN(new_n12171_));
  NOR2_X1    g12107(.A1(new_n12103_), .A2(new_n12171_), .ZN(new_n12172_));
  NOR2_X1    g12108(.A1(new_n12172_), .A2(new_n12170_), .ZN(new_n12173_));
  XNOR2_X1   g12109(.A1(new_n12096_), .A2(new_n12171_), .ZN(new_n12174_));
  NAND2_X1   g12110(.A1(new_n12145_), .A2(new_n12174_), .ZN(new_n12175_));
  OAI21_X1   g12111(.A1(new_n12145_), .A2(new_n12173_), .B(new_n12175_), .ZN(new_n12176_));
  NAND2_X1   g12112(.A1(new_n10926_), .A2(new_n10928_), .ZN(new_n12177_));
  OAI21_X1   g12113(.A1(new_n8737_), .A2(new_n10929_), .B(new_n12177_), .ZN(new_n12178_));
  XOR2_X1    g12114(.A1(new_n8725_), .A2(new_n8735_), .Z(new_n12179_));
  NAND3_X1   g12115(.A1(new_n10926_), .A2(new_n10928_), .A3(new_n12179_), .ZN(new_n12180_));
  AND2_X2    g12116(.A1(new_n12178_), .A2(new_n12180_), .Z(new_n12181_));
  OAI22_X1   g12117(.A1(new_n8735_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n10924_), .ZN(new_n12182_));
  NAND2_X1   g12118(.A1(new_n8726_), .A2(new_n2750_), .ZN(new_n12183_));
  AOI21_X1   g12119(.A1(new_n12183_), .A2(new_n12182_), .B(new_n2737_), .ZN(new_n12184_));
  NAND2_X1   g12120(.A1(new_n12181_), .A2(new_n12184_), .ZN(new_n12185_));
  XOR2_X1    g12121(.A1(new_n12185_), .A2(\a[29] ), .Z(new_n12186_));
  XOR2_X1    g12122(.A1(new_n8751_), .A2(new_n8746_), .Z(new_n12187_));
  OAI21_X1   g12123(.A1(new_n8753_), .A2(new_n10917_), .B(new_n10916_), .ZN(new_n12188_));
  OAI21_X1   g12124(.A1(new_n10916_), .A2(new_n12187_), .B(new_n12188_), .ZN(new_n12189_));
  AOI21_X1   g12125(.A1(new_n8761_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n12190_));
  OAI21_X1   g12126(.A1(new_n8745_), .A2(new_n2767_), .B(new_n12190_), .ZN(new_n12191_));
  AOI21_X1   g12127(.A1(new_n3332_), .A2(new_n8752_), .B(new_n12191_), .ZN(new_n12192_));
  AND2_X2    g12128(.A1(new_n12189_), .A2(new_n12192_), .Z(new_n12193_));
  INV_X1     g12129(.I(new_n12193_), .ZN(new_n12194_));
  XOR2_X1    g12130(.A1(new_n12186_), .A2(new_n12194_), .Z(new_n12195_));
  AND2_X2    g12131(.A1(new_n12176_), .A2(new_n12195_), .Z(new_n12196_));
  AND2_X2    g12132(.A1(new_n12186_), .A2(new_n12194_), .Z(new_n12197_));
  INV_X1     g12133(.I(new_n12197_), .ZN(new_n12198_));
  NOR2_X1    g12134(.A1(new_n12186_), .A2(new_n12194_), .ZN(new_n12199_));
  INV_X1     g12135(.I(new_n12199_), .ZN(new_n12200_));
  AOI21_X1   g12136(.A1(new_n12198_), .A2(new_n12200_), .B(new_n12176_), .ZN(new_n12201_));
  AOI21_X1   g12137(.A1(new_n8713_), .A2(new_n10949_), .B(new_n10936_), .ZN(new_n12202_));
  XNOR2_X1   g12138(.A1(new_n8701_), .A2(new_n8710_), .ZN(new_n12203_));
  NOR3_X1    g12139(.A1(new_n10948_), .A2(new_n8720_), .A3(new_n12203_), .ZN(new_n12204_));
  NOR2_X1    g12140(.A1(new_n12202_), .A2(new_n12204_), .ZN(new_n12205_));
  OAI22_X1   g12141(.A1(new_n8710_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8718_), .ZN(new_n12206_));
  NAND2_X1   g12142(.A1(new_n8702_), .A2(new_n3317_), .ZN(new_n12207_));
  AOI21_X1   g12143(.A1(new_n12207_), .A2(new_n12206_), .B(new_n3260_), .ZN(new_n12208_));
  NAND2_X1   g12144(.A1(new_n12205_), .A2(new_n12208_), .ZN(new_n12209_));
  XOR2_X1    g12145(.A1(new_n12209_), .A2(\a[26] ), .Z(new_n12210_));
  OAI21_X1   g12146(.A1(new_n12196_), .A2(new_n12201_), .B(new_n12210_), .ZN(new_n12211_));
  NOR2_X1    g12147(.A1(new_n12196_), .A2(new_n12201_), .ZN(new_n12212_));
  INV_X1     g12148(.I(new_n12210_), .ZN(new_n12213_));
  NAND2_X1   g12149(.A1(new_n12212_), .A2(new_n12213_), .ZN(new_n12214_));
  AOI22_X1   g12150(.A1(new_n12214_), .A2(new_n12211_), .B1(new_n12129_), .B2(new_n12144_), .ZN(new_n12215_));
  NAND2_X1   g12151(.A1(new_n12144_), .A2(new_n12129_), .ZN(new_n12216_));
  XOR2_X1    g12152(.A1(new_n12212_), .A2(new_n12210_), .Z(new_n12217_));
  NOR2_X1    g12153(.A1(new_n12217_), .A2(new_n12216_), .ZN(new_n12218_));
  NOR2_X1    g12154(.A1(new_n12218_), .A2(new_n12215_), .ZN(new_n12219_));
  INV_X1     g12155(.I(new_n12219_), .ZN(new_n12220_));
  OAI22_X1   g12156(.A1(new_n8681_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8694_), .ZN(new_n12221_));
  NAND2_X1   g12157(.A1(new_n8688_), .A2(new_n3312_), .ZN(new_n12222_));
  AOI21_X1   g12158(.A1(new_n12222_), .A2(new_n12221_), .B(new_n3302_), .ZN(new_n12223_));
  NAND2_X1   g12159(.A1(new_n11420_), .A2(new_n12223_), .ZN(new_n12224_));
  XOR2_X1    g12160(.A1(new_n12224_), .A2(\a[23] ), .Z(new_n12225_));
  INV_X1     g12161(.I(new_n12225_), .ZN(new_n12226_));
  NOR2_X1    g12162(.A1(new_n12220_), .A2(new_n12226_), .ZN(new_n12227_));
  INV_X1     g12163(.I(new_n12227_), .ZN(new_n12228_));
  NOR2_X1    g12164(.A1(new_n12219_), .A2(new_n12225_), .ZN(new_n12229_));
  AOI21_X1   g12165(.A1(new_n12228_), .A2(new_n12143_), .B(new_n12229_), .ZN(new_n12230_));
  INV_X1     g12166(.I(new_n12230_), .ZN(new_n12231_));
  OAI22_X1   g12167(.A1(new_n3322_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n3268_), .ZN(new_n12232_));
  NAND2_X1   g12168(.A1(new_n8696_), .A2(new_n3317_), .ZN(new_n12233_));
  AOI21_X1   g12169(.A1(new_n12232_), .A2(new_n12233_), .B(new_n3260_), .ZN(new_n12234_));
  NAND2_X1   g12170(.A1(new_n11595_), .A2(new_n12234_), .ZN(new_n12235_));
  XOR2_X1    g12171(.A1(new_n12235_), .A2(\a[26] ), .Z(new_n12236_));
  NOR2_X1    g12172(.A1(new_n10930_), .A2(new_n8737_), .ZN(new_n12237_));
  XOR2_X1    g12173(.A1(new_n8725_), .A2(new_n8719_), .Z(new_n12238_));
  NOR2_X1    g12174(.A1(new_n12237_), .A2(new_n12238_), .ZN(new_n12239_));
  NOR2_X1    g12175(.A1(new_n8727_), .A2(new_n10931_), .ZN(new_n12240_));
  NOR3_X1    g12176(.A1(new_n10930_), .A2(new_n8737_), .A3(new_n12240_), .ZN(new_n12241_));
  OR2_X2     g12177(.A1(new_n12239_), .A2(new_n12241_), .Z(new_n12242_));
  OAI22_X1   g12178(.A1(new_n8725_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8735_), .ZN(new_n12243_));
  NAND2_X1   g12179(.A1(new_n8719_), .A2(new_n2750_), .ZN(new_n12244_));
  AOI21_X1   g12180(.A1(new_n12243_), .A2(new_n12244_), .B(new_n2737_), .ZN(new_n12245_));
  NAND2_X1   g12181(.A1(new_n12242_), .A2(new_n12245_), .ZN(new_n12246_));
  XOR2_X1    g12182(.A1(new_n12246_), .A2(\a[29] ), .Z(new_n12247_));
  INV_X1     g12183(.I(new_n12247_), .ZN(new_n12248_));
  NAND2_X1   g12184(.A1(new_n12216_), .A2(new_n12211_), .ZN(new_n12249_));
  NAND2_X1   g12185(.A1(new_n12249_), .A2(new_n12214_), .ZN(new_n12250_));
  NAND2_X1   g12186(.A1(new_n12176_), .A2(new_n12198_), .ZN(new_n12251_));
  NAND2_X1   g12187(.A1(new_n12251_), .A2(new_n12200_), .ZN(new_n12252_));
  NOR2_X1    g12188(.A1(new_n12145_), .A2(new_n12170_), .ZN(new_n12253_));
  NOR2_X1    g12189(.A1(new_n12253_), .A2(new_n12172_), .ZN(new_n12254_));
  NAND2_X1   g12190(.A1(new_n4710_), .A2(new_n4719_), .ZN(new_n12255_));
  NOR3_X1    g12191(.A1(new_n12255_), .A2(new_n4706_), .A3(new_n6480_), .ZN(new_n12256_));
  NOR2_X1    g12192(.A1(new_n12256_), .A2(new_n4034_), .ZN(new_n12257_));
  INV_X1     g12193(.I(new_n12257_), .ZN(new_n12258_));
  NOR2_X1    g12194(.A1(new_n11461_), .A2(new_n12258_), .ZN(new_n12259_));
  NOR2_X1    g12195(.A1(new_n11461_), .A2(new_n12256_), .ZN(new_n12260_));
  NOR2_X1    g12196(.A1(new_n12260_), .A2(\a[11] ), .ZN(new_n12261_));
  NOR2_X1    g12197(.A1(new_n12261_), .A2(new_n12259_), .ZN(new_n12262_));
  INV_X1     g12198(.I(new_n1207_), .ZN(new_n12263_));
  NAND3_X1   g12199(.A1(new_n1404_), .A2(new_n1638_), .A3(new_n1096_), .ZN(new_n12264_));
  NOR4_X1    g12200(.A1(new_n12263_), .A2(new_n136_), .A3(new_n239_), .A4(new_n12264_), .ZN(new_n12265_));
  INV_X1     g12201(.I(new_n3493_), .ZN(new_n12266_));
  NOR4_X1    g12202(.A1(new_n289_), .A2(new_n487_), .A3(new_n560_), .A4(new_n163_), .ZN(new_n12267_));
  NOR3_X1    g12203(.A1(new_n12266_), .A2(new_n12267_), .A3(new_n2462_), .ZN(new_n12268_));
  NOR3_X1    g12204(.A1(new_n2389_), .A2(new_n1200_), .A3(new_n1864_), .ZN(new_n12269_));
  INV_X1     g12205(.I(new_n1623_), .ZN(new_n12270_));
  NOR2_X1    g12206(.A1(new_n2538_), .A2(new_n12270_), .ZN(new_n12271_));
  NAND4_X1   g12207(.A1(new_n12265_), .A2(new_n12268_), .A3(new_n12269_), .A4(new_n12271_), .ZN(new_n12272_));
  NOR2_X1    g12208(.A1(new_n622_), .A2(new_n12272_), .ZN(new_n12273_));
  NAND4_X1   g12209(.A1(new_n12273_), .A2(new_n878_), .A3(new_n2374_), .A4(new_n4406_), .ZN(new_n12274_));
  NAND2_X1   g12210(.A1(new_n12096_), .A2(new_n12274_), .ZN(new_n12275_));
  NOR2_X1    g12211(.A1(new_n12096_), .A2(new_n12274_), .ZN(new_n12276_));
  INV_X1     g12212(.I(new_n12276_), .ZN(new_n12277_));
  AOI21_X1   g12213(.A1(new_n12275_), .A2(new_n12277_), .B(new_n12262_), .ZN(new_n12278_));
  XNOR2_X1   g12214(.A1(new_n12096_), .A2(new_n12274_), .ZN(new_n12279_));
  INV_X1     g12215(.I(new_n12279_), .ZN(new_n12280_));
  AOI21_X1   g12216(.A1(new_n12262_), .A2(new_n12280_), .B(new_n12278_), .ZN(new_n12281_));
  NOR2_X1    g12217(.A1(new_n8751_), .A2(new_n2767_), .ZN(new_n12282_));
  NOR2_X1    g12218(.A1(new_n10924_), .A2(new_n2772_), .ZN(new_n12283_));
  NOR2_X1    g12219(.A1(new_n8745_), .A2(new_n2771_), .ZN(new_n12284_));
  NOR4_X1    g12220(.A1(new_n12282_), .A2(new_n2763_), .A3(new_n12283_), .A4(new_n12284_), .ZN(new_n12285_));
  NAND2_X1   g12221(.A1(new_n12072_), .A2(new_n12285_), .ZN(new_n12286_));
  INV_X1     g12222(.I(new_n12286_), .ZN(new_n12287_));
  NOR2_X1    g12223(.A1(new_n12281_), .A2(new_n12287_), .ZN(new_n12288_));
  NAND2_X1   g12224(.A1(new_n12281_), .A2(new_n12287_), .ZN(new_n12289_));
  INV_X1     g12225(.I(new_n12289_), .ZN(new_n12290_));
  NOR2_X1    g12226(.A1(new_n12290_), .A2(new_n12288_), .ZN(new_n12291_));
  XOR2_X1    g12227(.A1(new_n12281_), .A2(new_n12287_), .Z(new_n12292_));
  NAND2_X1   g12228(.A1(new_n12292_), .A2(new_n12254_), .ZN(new_n12293_));
  OAI21_X1   g12229(.A1(new_n12254_), .A2(new_n12291_), .B(new_n12293_), .ZN(new_n12294_));
  XOR2_X1    g12230(.A1(new_n12294_), .A2(new_n12252_), .Z(new_n12295_));
  XOR2_X1    g12231(.A1(new_n12295_), .A2(new_n12250_), .Z(new_n12296_));
  XOR2_X1    g12232(.A1(new_n12296_), .A2(new_n12248_), .Z(new_n12297_));
  XOR2_X1    g12233(.A1(new_n12297_), .A2(new_n12236_), .Z(new_n12298_));
  OAI22_X1   g12234(.A1(new_n3310_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n3306_), .ZN(new_n12299_));
  NAND2_X1   g12235(.A1(new_n8674_), .A2(new_n3312_), .ZN(new_n12300_));
  AOI21_X1   g12236(.A1(new_n12300_), .A2(new_n12299_), .B(new_n3302_), .ZN(new_n12301_));
  NAND2_X1   g12237(.A1(new_n11431_), .A2(new_n12301_), .ZN(new_n12302_));
  XOR2_X1    g12238(.A1(new_n12302_), .A2(\a[23] ), .Z(new_n12303_));
  NAND2_X1   g12239(.A1(new_n12298_), .A2(new_n12303_), .ZN(new_n12304_));
  NAND2_X1   g12240(.A1(new_n12304_), .A2(new_n12231_), .ZN(new_n12305_));
  OR2_X2     g12241(.A1(new_n12298_), .A2(new_n12303_), .Z(new_n12306_));
  NAND2_X1   g12242(.A1(new_n12305_), .A2(new_n12306_), .ZN(new_n12307_));
  INV_X1     g12243(.I(new_n12236_), .ZN(new_n12308_));
  XOR2_X1    g12244(.A1(new_n12295_), .A2(new_n12248_), .Z(new_n12309_));
  NOR3_X1    g12245(.A1(new_n12309_), .A2(new_n12308_), .A3(new_n12250_), .ZN(new_n12310_));
  AOI21_X1   g12246(.A1(new_n12308_), .A2(new_n12250_), .B(new_n12310_), .ZN(new_n12311_));
  OAI21_X1   g12247(.A1(new_n12248_), .A2(new_n12294_), .B(new_n12252_), .ZN(new_n12312_));
  NAND2_X1   g12248(.A1(new_n12294_), .A2(new_n12248_), .ZN(new_n12313_));
  AND2_X2    g12249(.A1(new_n12312_), .A2(new_n12313_), .Z(new_n12314_));
  OAI21_X1   g12250(.A1(new_n12254_), .A2(new_n12288_), .B(new_n12289_), .ZN(new_n12315_));
  INV_X1     g12251(.I(new_n12315_), .ZN(new_n12316_));
  NAND2_X1   g12252(.A1(new_n12262_), .A2(new_n12275_), .ZN(new_n12317_));
  NAND2_X1   g12253(.A1(new_n12317_), .A2(new_n12277_), .ZN(new_n12318_));
  INV_X1     g12254(.I(new_n12111_), .ZN(new_n12319_));
  AOI21_X1   g12255(.A1(new_n10919_), .A2(new_n10927_), .B(new_n12069_), .ZN(new_n12320_));
  NAND3_X1   g12256(.A1(new_n12320_), .A2(new_n8735_), .A3(new_n12319_), .ZN(new_n12321_));
  NAND2_X1   g12257(.A1(new_n12321_), .A2(new_n12116_), .ZN(new_n12322_));
  NAND2_X1   g12258(.A1(new_n8736_), .A2(new_n3332_), .ZN(new_n12323_));
  NAND2_X1   g12259(.A1(new_n8752_), .A2(new_n2770_), .ZN(new_n12324_));
  AOI21_X1   g12260(.A1(new_n10927_), .A2(new_n3189_), .B(new_n2764_), .ZN(new_n12325_));
  NAND4_X1   g12261(.A1(new_n12322_), .A2(new_n12323_), .A3(new_n12324_), .A4(new_n12325_), .ZN(new_n12326_));
  XOR2_X1    g12262(.A1(new_n12326_), .A2(new_n11483_), .Z(new_n12327_));
  INV_X1     g12263(.I(new_n12327_), .ZN(new_n12328_));
  INV_X1     g12264(.I(new_n11483_), .ZN(new_n12329_));
  NOR2_X1    g12265(.A1(new_n12326_), .A2(new_n12329_), .ZN(new_n12330_));
  INV_X1     g12266(.I(new_n12330_), .ZN(new_n12331_));
  NAND2_X1   g12267(.A1(new_n12326_), .A2(new_n12329_), .ZN(new_n12332_));
  AOI21_X1   g12268(.A1(new_n12331_), .A2(new_n12332_), .B(new_n12318_), .ZN(new_n12333_));
  AOI21_X1   g12269(.A1(new_n12318_), .A2(new_n12328_), .B(new_n12333_), .ZN(new_n12334_));
  OAI22_X1   g12270(.A1(new_n8725_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n8718_), .ZN(new_n12335_));
  NAND2_X1   g12271(.A1(new_n8711_), .A2(new_n2750_), .ZN(new_n12336_));
  AOI21_X1   g12272(.A1(new_n12336_), .A2(new_n12335_), .B(new_n2737_), .ZN(new_n12337_));
  NAND2_X1   g12273(.A1(new_n11536_), .A2(new_n12337_), .ZN(new_n12338_));
  XOR2_X1    g12274(.A1(new_n12338_), .A2(\a[29] ), .Z(new_n12339_));
  XOR2_X1    g12275(.A1(new_n12334_), .A2(new_n12339_), .Z(new_n12340_));
  NOR2_X1    g12276(.A1(new_n12340_), .A2(new_n12316_), .ZN(new_n12341_));
  INV_X1     g12277(.I(new_n12339_), .ZN(new_n12342_));
  NOR2_X1    g12278(.A1(new_n12334_), .A2(new_n12342_), .ZN(new_n12343_));
  INV_X1     g12279(.I(new_n12343_), .ZN(new_n12344_));
  NAND2_X1   g12280(.A1(new_n12334_), .A2(new_n12342_), .ZN(new_n12345_));
  AOI21_X1   g12281(.A1(new_n12344_), .A2(new_n12345_), .B(new_n12315_), .ZN(new_n12346_));
  INV_X1     g12282(.I(new_n11612_), .ZN(new_n12347_));
  OAI22_X1   g12283(.A1(new_n8701_), .A2(new_n3268_), .B1(new_n8694_), .B2(new_n3322_), .ZN(new_n12348_));
  NAND2_X1   g12284(.A1(new_n8682_), .A2(new_n3317_), .ZN(new_n12349_));
  AOI21_X1   g12285(.A1(new_n12349_), .A2(new_n12348_), .B(new_n3260_), .ZN(new_n12350_));
  NAND2_X1   g12286(.A1(new_n12347_), .A2(new_n12350_), .ZN(new_n12351_));
  XOR2_X1    g12287(.A1(new_n12351_), .A2(\a[26] ), .Z(new_n12352_));
  OAI21_X1   g12288(.A1(new_n12341_), .A2(new_n12346_), .B(new_n12352_), .ZN(new_n12353_));
  NOR2_X1    g12289(.A1(new_n12341_), .A2(new_n12346_), .ZN(new_n12354_));
  INV_X1     g12290(.I(new_n12352_), .ZN(new_n12355_));
  NAND2_X1   g12291(.A1(new_n12354_), .A2(new_n12355_), .ZN(new_n12356_));
  AOI21_X1   g12292(.A1(new_n12353_), .A2(new_n12356_), .B(new_n12314_), .ZN(new_n12357_));
  INV_X1     g12293(.I(new_n12314_), .ZN(new_n12358_));
  XOR2_X1    g12294(.A1(new_n12354_), .A2(new_n12352_), .Z(new_n12359_));
  NOR2_X1    g12295(.A1(new_n12359_), .A2(new_n12358_), .ZN(new_n12360_));
  OAI22_X1   g12296(.A1(new_n8673_), .A2(new_n3306_), .B1(new_n8687_), .B2(new_n3310_), .ZN(new_n12361_));
  NAND2_X1   g12297(.A1(new_n8662_), .A2(new_n3312_), .ZN(new_n12362_));
  AOI21_X1   g12298(.A1(new_n12362_), .A2(new_n12361_), .B(new_n3302_), .ZN(new_n12363_));
  NAND2_X1   g12299(.A1(new_n11624_), .A2(new_n12363_), .ZN(new_n12364_));
  XOR2_X1    g12300(.A1(new_n12364_), .A2(\a[23] ), .Z(new_n12365_));
  INV_X1     g12301(.I(new_n12365_), .ZN(new_n12366_));
  NOR3_X1    g12302(.A1(new_n12360_), .A2(new_n12357_), .A3(new_n12366_), .ZN(new_n12367_));
  NOR2_X1    g12303(.A1(new_n12360_), .A2(new_n12357_), .ZN(new_n12368_));
  NOR2_X1    g12304(.A1(new_n12368_), .A2(new_n12365_), .ZN(new_n12369_));
  NOR2_X1    g12305(.A1(new_n12369_), .A2(new_n12367_), .ZN(new_n12370_));
  NOR2_X1    g12306(.A1(new_n12370_), .A2(new_n12311_), .ZN(new_n12371_));
  INV_X1     g12307(.I(new_n12311_), .ZN(new_n12372_));
  XOR2_X1    g12308(.A1(new_n12368_), .A2(new_n12366_), .Z(new_n12373_));
  NOR2_X1    g12309(.A1(new_n12373_), .A2(new_n12372_), .ZN(new_n12374_));
  NOR2_X1    g12310(.A1(new_n12374_), .A2(new_n12371_), .ZN(new_n12375_));
  INV_X1     g12311(.I(new_n12375_), .ZN(new_n12376_));
  OAI22_X1   g12312(.A1(new_n11284_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n11271_), .ZN(new_n12377_));
  NAND2_X1   g12313(.A1(new_n11311_), .A2(new_n4096_), .ZN(new_n12378_));
  AOI21_X1   g12314(.A1(new_n12377_), .A2(new_n12378_), .B(new_n4095_), .ZN(new_n12379_));
  NAND2_X1   g12315(.A1(new_n11391_), .A2(new_n12379_), .ZN(new_n12380_));
  XOR2_X1    g12316(.A1(new_n12380_), .A2(\a[20] ), .Z(new_n12381_));
  INV_X1     g12317(.I(new_n12381_), .ZN(new_n12382_));
  NOR2_X1    g12318(.A1(new_n12376_), .A2(new_n12382_), .ZN(new_n12383_));
  NOR2_X1    g12319(.A1(new_n12375_), .A2(new_n12381_), .ZN(new_n12384_));
  OAI21_X1   g12320(.A1(new_n12383_), .A2(new_n12384_), .B(new_n12307_), .ZN(new_n12385_));
  XOR2_X1    g12321(.A1(new_n12375_), .A2(new_n12382_), .Z(new_n12386_));
  OAI21_X1   g12322(.A1(new_n12307_), .A2(new_n12386_), .B(new_n12385_), .ZN(new_n12387_));
  NOR2_X1    g12323(.A1(new_n12227_), .A2(new_n12229_), .ZN(new_n12388_));
  NOR2_X1    g12324(.A1(new_n12388_), .A2(new_n12142_), .ZN(new_n12389_));
  XOR2_X1    g12325(.A1(new_n12219_), .A2(new_n12226_), .Z(new_n12390_));
  INV_X1     g12326(.I(new_n12390_), .ZN(new_n12391_));
  AOI21_X1   g12327(.A1(new_n12142_), .A2(new_n12391_), .B(new_n12389_), .ZN(new_n12392_));
  INV_X1     g12328(.I(new_n12392_), .ZN(new_n12393_));
  NOR2_X1    g12329(.A1(new_n12141_), .A2(new_n12138_), .ZN(new_n12394_));
  NOR2_X1    g12330(.A1(new_n12394_), .A2(new_n12080_), .ZN(new_n12395_));
  XOR2_X1    g12331(.A1(new_n12131_), .A2(new_n12137_), .Z(new_n12396_));
  AOI21_X1   g12332(.A1(new_n12080_), .A2(new_n12396_), .B(new_n12395_), .ZN(new_n12397_));
  INV_X1     g12333(.I(new_n12397_), .ZN(new_n12398_));
  OAI22_X1   g12334(.A1(new_n8735_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n10924_), .ZN(new_n12399_));
  NAND2_X1   g12335(.A1(new_n8726_), .A2(new_n3317_), .ZN(new_n12400_));
  AOI21_X1   g12336(.A1(new_n12400_), .A2(new_n12399_), .B(new_n3260_), .ZN(new_n12401_));
  NAND2_X1   g12337(.A1(new_n12181_), .A2(new_n12401_), .ZN(new_n12402_));
  XOR2_X1    g12338(.A1(new_n12402_), .A2(\a[26] ), .Z(new_n12403_));
  OAI22_X1   g12339(.A1(new_n8745_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8758_), .ZN(new_n12404_));
  NAND2_X1   g12340(.A1(new_n8752_), .A2(new_n2750_), .ZN(new_n12405_));
  AOI21_X1   g12341(.A1(new_n12405_), .A2(new_n12404_), .B(new_n2737_), .ZN(new_n12406_));
  NAND2_X1   g12342(.A1(new_n12189_), .A2(new_n12406_), .ZN(new_n12407_));
  XOR2_X1    g12343(.A1(new_n12407_), .A2(\a[29] ), .Z(new_n12408_));
  NOR2_X1    g12344(.A1(new_n12403_), .A2(new_n12408_), .ZN(new_n12409_));
  INV_X1     g12345(.I(new_n11826_), .ZN(new_n12410_));
  AOI21_X1   g12346(.A1(new_n11781_), .A2(new_n11780_), .B(new_n12410_), .ZN(new_n12411_));
  NAND3_X1   g12347(.A1(new_n11781_), .A2(new_n11780_), .A3(new_n11852_), .ZN(new_n12412_));
  OAI21_X1   g12348(.A1(new_n12411_), .A2(new_n11828_), .B(new_n12412_), .ZN(new_n12413_));
  OAI21_X1   g12349(.A1(new_n11785_), .A2(new_n11784_), .B(new_n11849_), .ZN(new_n12414_));
  NOR3_X1    g12350(.A1(new_n11785_), .A2(new_n11784_), .A3(new_n11862_), .ZN(new_n12415_));
  AOI21_X1   g12351(.A1(new_n12413_), .A2(new_n12414_), .B(new_n12415_), .ZN(new_n12416_));
  NOR2_X1    g12352(.A1(new_n12416_), .A2(new_n11865_), .ZN(new_n12417_));
  NAND2_X1   g12353(.A1(new_n11891_), .A2(new_n11892_), .ZN(new_n12418_));
  NAND2_X1   g12354(.A1(new_n11874_), .A2(new_n11885_), .ZN(new_n12419_));
  AOI21_X1   g12355(.A1(new_n12418_), .A2(new_n12419_), .B(new_n11895_), .ZN(new_n12420_));
  AOI21_X1   g12356(.A1(new_n11917_), .A2(new_n11952_), .B(new_n11782_), .ZN(new_n12421_));
  INV_X1     g12357(.I(new_n11913_), .ZN(new_n12422_));
  NOR3_X1    g12358(.A1(new_n12420_), .A2(new_n12421_), .A3(new_n12422_), .ZN(new_n12423_));
  OAI21_X1   g12359(.A1(new_n12420_), .A2(new_n12421_), .B(new_n12422_), .ZN(new_n12424_));
  OAI21_X1   g12360(.A1(new_n12417_), .A2(new_n12423_), .B(new_n12424_), .ZN(new_n12425_));
  INV_X1     g12361(.I(new_n11977_), .ZN(new_n12426_));
  AOI21_X1   g12362(.A1(new_n12425_), .A2(new_n11970_), .B(new_n12426_), .ZN(new_n12427_));
  INV_X1     g12363(.I(new_n11990_), .ZN(new_n12428_));
  NAND2_X1   g12364(.A1(new_n12428_), .A2(new_n11993_), .ZN(new_n12429_));
  NAND2_X1   g12365(.A1(new_n12429_), .A2(new_n12007_), .ZN(new_n12430_));
  NOR3_X1    g12366(.A1(new_n11994_), .A2(new_n11990_), .A3(new_n12007_), .ZN(new_n12431_));
  INV_X1     g12367(.I(new_n12431_), .ZN(new_n12432_));
  AOI21_X1   g12368(.A1(new_n12430_), .A2(new_n12432_), .B(new_n12427_), .ZN(new_n12433_));
  AOI21_X1   g12369(.A1(new_n12008_), .A2(new_n12009_), .B(new_n11978_), .ZN(new_n12434_));
  NOR2_X1    g12370(.A1(new_n12433_), .A2(new_n12434_), .ZN(new_n12435_));
  NAND2_X1   g12371(.A1(new_n12403_), .A2(new_n12408_), .ZN(new_n12436_));
  AOI21_X1   g12372(.A1(new_n12435_), .A2(new_n12436_), .B(new_n12409_), .ZN(new_n12437_));
  INV_X1     g12373(.I(new_n12437_), .ZN(new_n12438_));
  OAI22_X1   g12374(.A1(new_n8725_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8735_), .ZN(new_n12439_));
  NAND2_X1   g12375(.A1(new_n8719_), .A2(new_n3317_), .ZN(new_n12440_));
  AOI21_X1   g12376(.A1(new_n12439_), .A2(new_n12440_), .B(new_n3260_), .ZN(new_n12441_));
  NAND2_X1   g12377(.A1(new_n12242_), .A2(new_n12441_), .ZN(new_n12442_));
  XOR2_X1    g12378(.A1(new_n12442_), .A2(\a[26] ), .Z(new_n12443_));
  INV_X1     g12379(.I(new_n12443_), .ZN(new_n12444_));
  NAND2_X1   g12380(.A1(new_n12438_), .A2(new_n12444_), .ZN(new_n12445_));
  XNOR2_X1   g12381(.A1(new_n12068_), .A2(new_n12077_), .ZN(new_n12446_));
  NOR2_X1    g12382(.A1(new_n12446_), .A2(new_n12011_), .ZN(new_n12447_));
  INV_X1     g12383(.I(new_n12079_), .ZN(new_n12448_));
  AOI21_X1   g12384(.A1(new_n12448_), .A2(new_n12078_), .B(new_n12012_), .ZN(new_n12449_));
  NOR2_X1    g12385(.A1(new_n12447_), .A2(new_n12449_), .ZN(new_n12450_));
  OAI21_X1   g12386(.A1(new_n12438_), .A2(new_n12444_), .B(new_n12450_), .ZN(new_n12451_));
  NAND2_X1   g12387(.A1(new_n12451_), .A2(new_n12445_), .ZN(new_n12452_));
  INV_X1     g12388(.I(new_n12452_), .ZN(new_n12453_));
  OAI22_X1   g12389(.A1(new_n8701_), .A2(new_n3310_), .B1(new_n8694_), .B2(new_n3306_), .ZN(new_n12454_));
  NAND2_X1   g12390(.A1(new_n8682_), .A2(new_n3312_), .ZN(new_n12455_));
  AOI21_X1   g12391(.A1(new_n12455_), .A2(new_n12454_), .B(new_n3302_), .ZN(new_n12456_));
  NAND2_X1   g12392(.A1(new_n12347_), .A2(new_n12456_), .ZN(new_n12457_));
  XOR2_X1    g12393(.A1(new_n12457_), .A2(\a[23] ), .Z(new_n12458_));
  NAND2_X1   g12394(.A1(new_n12453_), .A2(new_n12458_), .ZN(new_n12459_));
  INV_X1     g12395(.I(new_n12458_), .ZN(new_n12460_));
  NAND2_X1   g12396(.A1(new_n12452_), .A2(new_n12460_), .ZN(new_n12461_));
  INV_X1     g12397(.I(new_n12461_), .ZN(new_n12462_));
  AOI21_X1   g12398(.A1(new_n12398_), .A2(new_n12459_), .B(new_n12462_), .ZN(new_n12463_));
  OAI22_X1   g12399(.A1(new_n8661_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n8673_), .ZN(new_n12464_));
  NAND2_X1   g12400(.A1(new_n11285_), .A2(new_n4096_), .ZN(new_n12465_));
  AOI21_X1   g12401(.A1(new_n12465_), .A2(new_n12464_), .B(new_n4095_), .ZN(new_n12466_));
  NAND2_X1   g12402(.A1(new_n11323_), .A2(new_n12466_), .ZN(new_n12467_));
  XOR2_X1    g12403(.A1(new_n12467_), .A2(\a[20] ), .Z(new_n12468_));
  NAND2_X1   g12404(.A1(new_n12463_), .A2(new_n12468_), .ZN(new_n12469_));
  NOR2_X1    g12405(.A1(new_n12463_), .A2(new_n12468_), .ZN(new_n12470_));
  AOI21_X1   g12406(.A1(new_n12393_), .A2(new_n12469_), .B(new_n12470_), .ZN(new_n12471_));
  OAI22_X1   g12407(.A1(new_n11284_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n8661_), .ZN(new_n12472_));
  NAND2_X1   g12408(.A1(new_n11272_), .A2(new_n4096_), .ZN(new_n12473_));
  AOI21_X1   g12409(.A1(new_n12472_), .A2(new_n12473_), .B(new_n4095_), .ZN(new_n12474_));
  NAND2_X1   g12410(.A1(new_n11655_), .A2(new_n12474_), .ZN(new_n12475_));
  XOR2_X1    g12411(.A1(new_n12475_), .A2(\a[20] ), .Z(new_n12476_));
  NOR2_X1    g12412(.A1(new_n12471_), .A2(new_n12476_), .ZN(new_n12477_));
  XNOR2_X1   g12413(.A1(new_n12298_), .A2(new_n12303_), .ZN(new_n12478_));
  NOR2_X1    g12414(.A1(new_n12478_), .A2(new_n12230_), .ZN(new_n12479_));
  AOI21_X1   g12415(.A1(new_n12306_), .A2(new_n12304_), .B(new_n12231_), .ZN(new_n12480_));
  NOR2_X1    g12416(.A1(new_n12479_), .A2(new_n12480_), .ZN(new_n12481_));
  NAND2_X1   g12417(.A1(new_n12471_), .A2(new_n12476_), .ZN(new_n12482_));
  AOI21_X1   g12418(.A1(new_n12481_), .A2(new_n12482_), .B(new_n12477_), .ZN(new_n12483_));
  OAI22_X1   g12419(.A1(new_n11264_), .A2(new_n4291_), .B1(new_n4297_), .B2(new_n11345_), .ZN(new_n12484_));
  NAND2_X1   g12420(.A1(new_n11354_), .A2(new_n4469_), .ZN(new_n12485_));
  AOI21_X1   g12421(.A1(new_n12485_), .A2(new_n12484_), .B(new_n4468_), .ZN(new_n12486_));
  NAND2_X1   g12422(.A1(new_n11678_), .A2(new_n12486_), .ZN(new_n12487_));
  XOR2_X1    g12423(.A1(new_n12487_), .A2(\a[17] ), .Z(new_n12488_));
  NAND2_X1   g12424(.A1(new_n12483_), .A2(new_n12488_), .ZN(new_n12489_));
  NAND2_X1   g12425(.A1(new_n12489_), .A2(new_n12387_), .ZN(new_n12490_));
  NOR2_X1    g12426(.A1(new_n12483_), .A2(new_n12488_), .ZN(new_n12491_));
  INV_X1     g12427(.I(new_n12491_), .ZN(new_n12492_));
  NAND2_X1   g12428(.A1(new_n12490_), .A2(new_n12492_), .ZN(new_n12493_));
  INV_X1     g12429(.I(new_n12383_), .ZN(new_n12494_));
  AOI21_X1   g12430(.A1(new_n12494_), .A2(new_n12307_), .B(new_n12384_), .ZN(new_n12495_));
  OAI21_X1   g12431(.A1(new_n12316_), .A2(new_n12343_), .B(new_n12345_), .ZN(new_n12496_));
  INV_X1     g12432(.I(new_n12496_), .ZN(new_n12497_));
  NAND2_X1   g12433(.A1(new_n12318_), .A2(new_n12332_), .ZN(new_n12498_));
  NAND2_X1   g12434(.A1(new_n12498_), .A2(new_n12331_), .ZN(new_n12499_));
  INV_X1     g12435(.I(new_n12181_), .ZN(new_n12500_));
  NOR2_X1    g12436(.A1(new_n8725_), .A2(new_n2772_), .ZN(new_n12501_));
  NOR2_X1    g12437(.A1(new_n8735_), .A2(new_n2767_), .ZN(new_n12502_));
  NOR2_X1    g12438(.A1(new_n10924_), .A2(new_n2771_), .ZN(new_n12503_));
  NOR4_X1    g12439(.A1(new_n12501_), .A2(new_n2764_), .A3(new_n12502_), .A4(new_n12503_), .ZN(new_n12504_));
  NAND2_X1   g12440(.A1(new_n12500_), .A2(new_n12504_), .ZN(new_n12505_));
  INV_X1     g12441(.I(new_n2156_), .ZN(new_n12506_));
  NOR2_X1    g12442(.A1(new_n2777_), .A2(new_n2546_), .ZN(new_n12507_));
  NAND4_X1   g12443(.A1(new_n382_), .A2(new_n1706_), .A3(new_n1436_), .A4(new_n540_), .ZN(new_n12508_));
  NAND4_X1   g12444(.A1(new_n385_), .A2(new_n1719_), .A3(new_n467_), .A4(new_n643_), .ZN(new_n12509_));
  NAND3_X1   g12445(.A1(new_n12509_), .A2(new_n391_), .A3(new_n1088_), .ZN(new_n12510_));
  NAND3_X1   g12446(.A1(new_n2307_), .A2(new_n1575_), .A3(new_n1460_), .ZN(new_n12511_));
  NAND2_X1   g12447(.A1(new_n2368_), .A2(new_n188_), .ZN(new_n12512_));
  NOR4_X1    g12448(.A1(new_n12510_), .A2(new_n12511_), .A3(new_n2488_), .A4(new_n12512_), .ZN(new_n12513_));
  NAND4_X1   g12449(.A1(new_n12513_), .A2(new_n12166_), .A3(new_n12507_), .A4(new_n12508_), .ZN(new_n12514_));
  NOR2_X1    g12450(.A1(new_n932_), .A2(new_n1417_), .ZN(new_n12515_));
  NAND4_X1   g12451(.A1(new_n2837_), .A2(new_n12515_), .A3(new_n1657_), .A4(new_n3365_), .ZN(new_n12516_));
  NOR3_X1    g12452(.A1(new_n1784_), .A2(new_n135_), .A3(new_n615_), .ZN(new_n12517_));
  INV_X1     g12453(.I(new_n12517_), .ZN(new_n12518_));
  NAND2_X1   g12454(.A1(new_n1471_), .A2(new_n1765_), .ZN(new_n12519_));
  NOR4_X1    g12455(.A1(new_n212_), .A2(new_n235_), .A3(new_n226_), .A4(new_n397_), .ZN(new_n12520_));
  NOR4_X1    g12456(.A1(new_n12518_), .A2(new_n2969_), .A3(new_n12519_), .A4(new_n12520_), .ZN(new_n12521_));
  AND3_X2    g12457(.A1(new_n1321_), .A2(new_n971_), .A3(new_n2444_), .Z(new_n12522_));
  NAND4_X1   g12458(.A1(new_n2375_), .A2(new_n221_), .A3(new_n383_), .A4(new_n677_), .ZN(new_n12523_));
  NAND4_X1   g12459(.A1(new_n248_), .A2(new_n807_), .A3(new_n423_), .A4(new_n1638_), .ZN(new_n12524_));
  NAND4_X1   g12460(.A1(new_n12521_), .A2(new_n12522_), .A3(new_n12523_), .A4(new_n12524_), .ZN(new_n12525_));
  NOR4_X1    g12461(.A1(new_n12506_), .A2(new_n12514_), .A3(new_n12516_), .A4(new_n12525_), .ZN(new_n12526_));
  OR2_X2     g12462(.A1(new_n11483_), .A2(new_n12526_), .Z(new_n12527_));
  NAND2_X1   g12463(.A1(new_n11483_), .A2(new_n12526_), .ZN(new_n12528_));
  AOI21_X1   g12464(.A1(new_n12527_), .A2(new_n12528_), .B(new_n12505_), .ZN(new_n12529_));
  XNOR2_X1   g12465(.A1(new_n11483_), .A2(new_n12526_), .ZN(new_n12530_));
  AOI21_X1   g12466(.A1(new_n12500_), .A2(new_n12504_), .B(new_n12530_), .ZN(new_n12531_));
  NOR2_X1    g12467(.A1(new_n12529_), .A2(new_n12531_), .ZN(new_n12532_));
  XOR2_X1    g12468(.A1(new_n12499_), .A2(new_n12532_), .Z(new_n12533_));
  NOR2_X1    g12469(.A1(new_n12497_), .A2(new_n12533_), .ZN(new_n12534_));
  INV_X1     g12470(.I(new_n12532_), .ZN(new_n12535_));
  NOR2_X1    g12471(.A1(new_n12499_), .A2(new_n12535_), .ZN(new_n12536_));
  INV_X1     g12472(.I(new_n12536_), .ZN(new_n12537_));
  NAND2_X1   g12473(.A1(new_n12499_), .A2(new_n12535_), .ZN(new_n12538_));
  AOI21_X1   g12474(.A1(new_n12537_), .A2(new_n12538_), .B(new_n12496_), .ZN(new_n12539_));
  NOR2_X1    g12475(.A1(new_n12534_), .A2(new_n12539_), .ZN(new_n12540_));
  OAI22_X1   g12476(.A1(new_n8681_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8694_), .ZN(new_n12541_));
  NAND2_X1   g12477(.A1(new_n8688_), .A2(new_n3317_), .ZN(new_n12542_));
  AOI21_X1   g12478(.A1(new_n12542_), .A2(new_n12541_), .B(new_n3260_), .ZN(new_n12543_));
  NAND2_X1   g12479(.A1(new_n11420_), .A2(new_n12543_), .ZN(new_n12544_));
  XOR2_X1    g12480(.A1(new_n12544_), .A2(\a[26] ), .Z(new_n12545_));
  OAI22_X1   g12481(.A1(new_n8710_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8718_), .ZN(new_n12546_));
  NAND2_X1   g12482(.A1(new_n8702_), .A2(new_n2750_), .ZN(new_n12547_));
  AOI21_X1   g12483(.A1(new_n12547_), .A2(new_n12546_), .B(new_n2737_), .ZN(new_n12548_));
  NAND2_X1   g12484(.A1(new_n12205_), .A2(new_n12548_), .ZN(new_n12549_));
  XOR2_X1    g12485(.A1(new_n12549_), .A2(\a[29] ), .Z(new_n12550_));
  XNOR2_X1   g12486(.A1(new_n12545_), .A2(new_n12550_), .ZN(new_n12551_));
  NOR2_X1    g12487(.A1(new_n12540_), .A2(new_n12551_), .ZN(new_n12552_));
  NOR2_X1    g12488(.A1(new_n12545_), .A2(new_n12550_), .ZN(new_n12553_));
  NAND2_X1   g12489(.A1(new_n12545_), .A2(new_n12550_), .ZN(new_n12554_));
  INV_X1     g12490(.I(new_n12554_), .ZN(new_n12555_));
  NOR2_X1    g12491(.A1(new_n12555_), .A2(new_n12553_), .ZN(new_n12556_));
  INV_X1     g12492(.I(new_n12556_), .ZN(new_n12557_));
  AOI21_X1   g12493(.A1(new_n12540_), .A2(new_n12557_), .B(new_n12552_), .ZN(new_n12558_));
  INV_X1     g12494(.I(new_n12558_), .ZN(new_n12559_));
  NAND2_X1   g12495(.A1(new_n12358_), .A2(new_n12353_), .ZN(new_n12560_));
  NAND2_X1   g12496(.A1(new_n12560_), .A2(new_n12356_), .ZN(new_n12561_));
  OAI22_X1   g12497(.A1(new_n8661_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8673_), .ZN(new_n12562_));
  NAND2_X1   g12498(.A1(new_n11285_), .A2(new_n3312_), .ZN(new_n12563_));
  AOI21_X1   g12499(.A1(new_n12563_), .A2(new_n12562_), .B(new_n3302_), .ZN(new_n12564_));
  NAND2_X1   g12500(.A1(new_n11323_), .A2(new_n12564_), .ZN(new_n12565_));
  XOR2_X1    g12501(.A1(new_n12565_), .A2(\a[23] ), .Z(new_n12566_));
  INV_X1     g12502(.I(new_n12566_), .ZN(new_n12567_));
  NOR2_X1    g12503(.A1(new_n12561_), .A2(new_n12567_), .ZN(new_n12568_));
  NAND2_X1   g12504(.A1(new_n12561_), .A2(new_n12567_), .ZN(new_n12569_));
  INV_X1     g12505(.I(new_n12569_), .ZN(new_n12570_));
  OAI21_X1   g12506(.A1(new_n12570_), .A2(new_n12568_), .B(new_n12559_), .ZN(new_n12571_));
  XOR2_X1    g12507(.A1(new_n12561_), .A2(new_n12566_), .Z(new_n12572_));
  OAI21_X1   g12508(.A1(new_n12559_), .A2(new_n12572_), .B(new_n12571_), .ZN(new_n12573_));
  INV_X1     g12509(.I(new_n12573_), .ZN(new_n12574_));
  INV_X1     g12510(.I(new_n12367_), .ZN(new_n12575_));
  AOI21_X1   g12511(.A1(new_n12372_), .A2(new_n12575_), .B(new_n12369_), .ZN(new_n12576_));
  AOI22_X1   g12512(.A1(new_n11311_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n11272_), .ZN(new_n12577_));
  NOR2_X1    g12513(.A1(new_n11264_), .A2(new_n4097_), .ZN(new_n12578_));
  OAI21_X1   g12514(.A1(new_n12578_), .A2(new_n12577_), .B(new_n3773_), .ZN(new_n12579_));
  NOR2_X1    g12515(.A1(new_n11310_), .A2(new_n12579_), .ZN(new_n12580_));
  XOR2_X1    g12516(.A1(new_n12580_), .A2(new_n3035_), .Z(new_n12581_));
  AND2_X2    g12517(.A1(new_n12576_), .A2(new_n12581_), .Z(new_n12582_));
  NOR2_X1    g12518(.A1(new_n12576_), .A2(new_n12581_), .ZN(new_n12583_));
  NOR2_X1    g12519(.A1(new_n12582_), .A2(new_n12583_), .ZN(new_n12584_));
  NOR2_X1    g12520(.A1(new_n12584_), .A2(new_n12574_), .ZN(new_n12585_));
  XNOR2_X1   g12521(.A1(new_n12576_), .A2(new_n12581_), .ZN(new_n12586_));
  NOR2_X1    g12522(.A1(new_n12586_), .A2(new_n12573_), .ZN(new_n12587_));
  OAI22_X1   g12523(.A1(new_n11353_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n11345_), .ZN(new_n12588_));
  NAND2_X1   g12524(.A1(new_n11370_), .A2(new_n4469_), .ZN(new_n12589_));
  AOI21_X1   g12525(.A1(new_n12589_), .A2(new_n12588_), .B(new_n4468_), .ZN(new_n12590_));
  NAND2_X1   g12526(.A1(new_n11379_), .A2(new_n12590_), .ZN(new_n12591_));
  XOR2_X1    g12527(.A1(new_n12591_), .A2(\a[17] ), .Z(new_n12592_));
  INV_X1     g12528(.I(new_n12592_), .ZN(new_n12593_));
  NOR3_X1    g12529(.A1(new_n12585_), .A2(new_n12587_), .A3(new_n12593_), .ZN(new_n12594_));
  NOR2_X1    g12530(.A1(new_n12585_), .A2(new_n12587_), .ZN(new_n12595_));
  NOR2_X1    g12531(.A1(new_n12595_), .A2(new_n12592_), .ZN(new_n12596_));
  NOR2_X1    g12532(.A1(new_n12596_), .A2(new_n12594_), .ZN(new_n12597_));
  NOR2_X1    g12533(.A1(new_n12597_), .A2(new_n12495_), .ZN(new_n12598_));
  INV_X1     g12534(.I(new_n12495_), .ZN(new_n12599_));
  XOR2_X1    g12535(.A1(new_n12595_), .A2(new_n12593_), .Z(new_n12600_));
  NOR2_X1    g12536(.A1(new_n12600_), .A2(new_n12599_), .ZN(new_n12601_));
  NOR2_X1    g12537(.A1(new_n12601_), .A2(new_n12598_), .ZN(new_n12602_));
  INV_X1     g12538(.I(new_n12602_), .ZN(new_n12603_));
  AND3_X2    g12539(.A1(new_n11463_), .A2(new_n6180_), .A3(new_n11496_), .Z(new_n12604_));
  NOR4_X1    g12540(.A1(new_n11468_), .A2(new_n6082_), .A3(new_n11461_), .A4(new_n12604_), .ZN(new_n12605_));
  XOR2_X1    g12541(.A1(new_n12605_), .A2(new_n3521_), .Z(new_n12606_));
  INV_X1     g12542(.I(new_n12606_), .ZN(new_n12607_));
  NOR2_X1    g12543(.A1(new_n12603_), .A2(new_n12607_), .ZN(new_n12608_));
  NOR2_X1    g12544(.A1(new_n12602_), .A2(new_n12606_), .ZN(new_n12609_));
  OAI21_X1   g12545(.A1(new_n12608_), .A2(new_n12609_), .B(new_n12493_), .ZN(new_n12610_));
  XOR2_X1    g12546(.A1(new_n12602_), .A2(new_n12607_), .Z(new_n12611_));
  OAI21_X1   g12547(.A1(new_n12493_), .A2(new_n12611_), .B(new_n12610_), .ZN(new_n12612_));
  INV_X1     g12548(.I(new_n12387_), .ZN(new_n12613_));
  AOI21_X1   g12549(.A1(new_n12492_), .A2(new_n12489_), .B(new_n12613_), .ZN(new_n12614_));
  XNOR2_X1   g12550(.A1(new_n12483_), .A2(new_n12488_), .ZN(new_n12615_));
  NOR2_X1    g12551(.A1(new_n12615_), .A2(new_n12387_), .ZN(new_n12616_));
  NOR2_X1    g12552(.A1(new_n12616_), .A2(new_n12614_), .ZN(new_n12617_));
  INV_X1     g12553(.I(new_n12470_), .ZN(new_n12618_));
  AOI21_X1   g12554(.A1(new_n12618_), .A2(new_n12469_), .B(new_n12392_), .ZN(new_n12619_));
  XNOR2_X1   g12555(.A1(new_n12463_), .A2(new_n12468_), .ZN(new_n12620_));
  NOR2_X1    g12556(.A1(new_n12620_), .A2(new_n12393_), .ZN(new_n12621_));
  NOR2_X1    g12557(.A1(new_n12621_), .A2(new_n12619_), .ZN(new_n12622_));
  AOI21_X1   g12558(.A1(new_n12459_), .A2(new_n12461_), .B(new_n12397_), .ZN(new_n12623_));
  INV_X1     g12559(.I(new_n12623_), .ZN(new_n12624_));
  XOR2_X1    g12560(.A1(new_n12452_), .A2(new_n12460_), .Z(new_n12625_));
  NAND2_X1   g12561(.A1(new_n12625_), .A2(new_n12397_), .ZN(new_n12626_));
  NOR2_X1    g12562(.A1(new_n11995_), .A2(new_n12006_), .ZN(new_n12627_));
  OAI21_X1   g12563(.A1(new_n12627_), .A2(new_n12431_), .B(new_n11978_), .ZN(new_n12628_));
  NOR2_X1    g12564(.A1(new_n12429_), .A2(new_n12006_), .ZN(new_n12629_));
  OAI21_X1   g12565(.A1(new_n12629_), .A2(new_n12010_), .B(new_n12427_), .ZN(new_n12630_));
  XNOR2_X1   g12566(.A1(new_n12403_), .A2(new_n12408_), .ZN(new_n12631_));
  AOI21_X1   g12567(.A1(new_n12630_), .A2(new_n12628_), .B(new_n12631_), .ZN(new_n12632_));
  INV_X1     g12568(.I(new_n12436_), .ZN(new_n12633_));
  NOR2_X1    g12569(.A1(new_n12633_), .A2(new_n12409_), .ZN(new_n12634_));
  NOR3_X1    g12570(.A1(new_n12433_), .A2(new_n12434_), .A3(new_n12634_), .ZN(new_n12635_));
  NOR2_X1    g12571(.A1(new_n12632_), .A2(new_n12635_), .ZN(new_n12636_));
  NAND3_X1   g12572(.A1(new_n11975_), .A2(new_n11973_), .A3(new_n11969_), .ZN(new_n12637_));
  OAI21_X1   g12573(.A1(new_n11958_), .A2(new_n11951_), .B(new_n11976_), .ZN(new_n12638_));
  NAND2_X1   g12574(.A1(new_n12638_), .A2(new_n12637_), .ZN(new_n12639_));
  NAND2_X1   g12575(.A1(new_n12639_), .A2(new_n12425_), .ZN(new_n12640_));
  OAI21_X1   g12576(.A1(new_n11971_), .A2(new_n12426_), .B(new_n11916_), .ZN(new_n12641_));
  OAI22_X1   g12577(.A1(new_n8751_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n10924_), .ZN(new_n12642_));
  NAND2_X1   g12578(.A1(new_n8736_), .A2(new_n3317_), .ZN(new_n12643_));
  AOI21_X1   g12579(.A1(new_n12643_), .A2(new_n12642_), .B(new_n3260_), .ZN(new_n12644_));
  NAND2_X1   g12580(.A1(new_n12118_), .A2(new_n12644_), .ZN(new_n12645_));
  XOR2_X1    g12581(.A1(new_n12645_), .A2(\a[26] ), .Z(new_n12646_));
  INV_X1     g12582(.I(new_n12646_), .ZN(new_n12647_));
  NAND3_X1   g12583(.A1(new_n12641_), .A2(new_n12640_), .A3(new_n12647_), .ZN(new_n12648_));
  OAI22_X1   g12584(.A1(new_n8710_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8718_), .ZN(new_n12649_));
  NAND2_X1   g12585(.A1(new_n8702_), .A2(new_n3312_), .ZN(new_n12650_));
  AOI21_X1   g12586(.A1(new_n12650_), .A2(new_n12649_), .B(new_n3302_), .ZN(new_n12651_));
  NAND2_X1   g12587(.A1(new_n12205_), .A2(new_n12651_), .ZN(new_n12652_));
  XOR2_X1    g12588(.A1(new_n12652_), .A2(\a[23] ), .Z(new_n12653_));
  NAND2_X1   g12589(.A1(new_n12648_), .A2(new_n12653_), .ZN(new_n12654_));
  INV_X1     g12590(.I(new_n12654_), .ZN(new_n12655_));
  AOI21_X1   g12591(.A1(new_n12637_), .A2(new_n12638_), .B(new_n11916_), .ZN(new_n12656_));
  AOI21_X1   g12592(.A1(new_n11970_), .A2(new_n11977_), .B(new_n12425_), .ZN(new_n12657_));
  NOR2_X1    g12593(.A1(new_n12656_), .A2(new_n12657_), .ZN(new_n12658_));
  INV_X1     g12594(.I(new_n12653_), .ZN(new_n12659_));
  NAND3_X1   g12595(.A1(new_n12658_), .A2(new_n12647_), .A3(new_n12659_), .ZN(new_n12660_));
  OAI21_X1   g12596(.A1(new_n12636_), .A2(new_n12655_), .B(new_n12660_), .ZN(new_n12661_));
  INV_X1     g12597(.I(new_n12661_), .ZN(new_n12662_));
  OAI22_X1   g12598(.A1(new_n3306_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n3310_), .ZN(new_n12663_));
  NAND2_X1   g12599(.A1(new_n8696_), .A2(new_n3312_), .ZN(new_n12664_));
  AOI21_X1   g12600(.A1(new_n12663_), .A2(new_n12664_), .B(new_n3302_), .ZN(new_n12665_));
  NAND2_X1   g12601(.A1(new_n11595_), .A2(new_n12665_), .ZN(new_n12666_));
  XOR2_X1    g12602(.A1(new_n12666_), .A2(\a[23] ), .Z(new_n12667_));
  NOR2_X1    g12603(.A1(new_n12662_), .A2(new_n12667_), .ZN(new_n12668_));
  XOR2_X1    g12604(.A1(new_n12450_), .A2(new_n12443_), .Z(new_n12669_));
  NAND2_X1   g12605(.A1(new_n12669_), .A2(new_n12437_), .ZN(new_n12670_));
  XOR2_X1    g12606(.A1(new_n12450_), .A2(new_n12444_), .Z(new_n12671_));
  NAND2_X1   g12607(.A1(new_n12671_), .A2(new_n12438_), .ZN(new_n12672_));
  INV_X1     g12608(.I(new_n12667_), .ZN(new_n12673_));
  NOR2_X1    g12609(.A1(new_n12661_), .A2(new_n12673_), .ZN(new_n12674_));
  INV_X1     g12610(.I(new_n12674_), .ZN(new_n12675_));
  AOI21_X1   g12611(.A1(new_n12672_), .A2(new_n12670_), .B(new_n12675_), .ZN(new_n12676_));
  OAI22_X1   g12612(.A1(new_n8673_), .A2(new_n3775_), .B1(new_n8687_), .B2(new_n3769_), .ZN(new_n12677_));
  NAND2_X1   g12613(.A1(new_n8662_), .A2(new_n4096_), .ZN(new_n12678_));
  AOI21_X1   g12614(.A1(new_n12678_), .A2(new_n12677_), .B(new_n4095_), .ZN(new_n12679_));
  NAND2_X1   g12615(.A1(new_n11624_), .A2(new_n12679_), .ZN(new_n12680_));
  XOR2_X1    g12616(.A1(new_n12680_), .A2(\a[20] ), .Z(new_n12681_));
  INV_X1     g12617(.I(new_n12681_), .ZN(new_n12682_));
  NOR3_X1    g12618(.A1(new_n12676_), .A2(new_n12668_), .A3(new_n12682_), .ZN(new_n12683_));
  AOI21_X1   g12619(.A1(new_n12624_), .A2(new_n12626_), .B(new_n12683_), .ZN(new_n12684_));
  NOR2_X1    g12620(.A1(new_n12676_), .A2(new_n12668_), .ZN(new_n12685_));
  NOR2_X1    g12621(.A1(new_n12685_), .A2(new_n12681_), .ZN(new_n12686_));
  NOR2_X1    g12622(.A1(new_n12684_), .A2(new_n12686_), .ZN(new_n12687_));
  INV_X1     g12623(.I(new_n12687_), .ZN(new_n12688_));
  AOI22_X1   g12624(.A1(new_n11311_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n11272_), .ZN(new_n12689_));
  NOR2_X1    g12625(.A1(new_n11264_), .A2(new_n4470_), .ZN(new_n12690_));
  OAI21_X1   g12626(.A1(new_n12690_), .A2(new_n12689_), .B(new_n4295_), .ZN(new_n12691_));
  NOR2_X1    g12627(.A1(new_n11310_), .A2(new_n12691_), .ZN(new_n12692_));
  XOR2_X1    g12628(.A1(new_n12692_), .A2(new_n3372_), .Z(new_n12693_));
  INV_X1     g12629(.I(new_n12693_), .ZN(new_n12694_));
  NOR2_X1    g12630(.A1(new_n12688_), .A2(new_n12694_), .ZN(new_n12695_));
  NOR2_X1    g12631(.A1(new_n12622_), .A2(new_n12695_), .ZN(new_n12696_));
  NOR2_X1    g12632(.A1(new_n12687_), .A2(new_n12693_), .ZN(new_n12697_));
  NOR2_X1    g12633(.A1(new_n12696_), .A2(new_n12697_), .ZN(new_n12698_));
  OAI22_X1   g12634(.A1(new_n11264_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n11277_), .ZN(new_n12699_));
  NAND2_X1   g12635(.A1(new_n11346_), .A2(new_n4469_), .ZN(new_n12700_));
  AOI21_X1   g12636(.A1(new_n12699_), .A2(new_n12700_), .B(new_n4468_), .ZN(new_n12701_));
  NAND2_X1   g12637(.A1(new_n11757_), .A2(new_n12701_), .ZN(new_n12702_));
  XOR2_X1    g12638(.A1(new_n12702_), .A2(\a[17] ), .Z(new_n12703_));
  NOR2_X1    g12639(.A1(new_n12698_), .A2(new_n12703_), .ZN(new_n12704_));
  INV_X1     g12640(.I(new_n12471_), .ZN(new_n12705_));
  XNOR2_X1   g12641(.A1(new_n12481_), .A2(new_n12476_), .ZN(new_n12706_));
  XOR2_X1    g12642(.A1(new_n12706_), .A2(new_n12705_), .Z(new_n12707_));
  NAND2_X1   g12643(.A1(new_n12698_), .A2(new_n12703_), .ZN(new_n12708_));
  NOR2_X1    g12644(.A1(new_n12707_), .A2(new_n12708_), .ZN(new_n12709_));
  NOR2_X1    g12645(.A1(new_n12709_), .A2(new_n12704_), .ZN(new_n12710_));
  INV_X1     g12646(.I(new_n12710_), .ZN(new_n12711_));
  NAND3_X1   g12647(.A1(new_n11359_), .A2(new_n11354_), .A3(new_n11369_), .ZN(new_n12712_));
  NAND2_X1   g12648(.A1(new_n11692_), .A2(new_n11370_), .ZN(new_n12713_));
  AOI21_X1   g12649(.A1(new_n12713_), .A2(new_n12712_), .B(new_n11461_), .ZN(new_n12714_));
  INV_X1     g12650(.I(new_n12714_), .ZN(new_n12715_));
  NOR2_X1    g12651(.A1(new_n11692_), .A2(new_n11369_), .ZN(new_n12716_));
  INV_X1     g12652(.I(new_n12716_), .ZN(new_n12717_));
  NAND3_X1   g12653(.A1(new_n12715_), .A2(new_n11463_), .A3(new_n12717_), .ZN(new_n12718_));
  OAI21_X1   g12654(.A1(new_n12714_), .A2(new_n11466_), .B(new_n12716_), .ZN(new_n12719_));
  NAND2_X1   g12655(.A1(new_n12718_), .A2(new_n12719_), .ZN(new_n12720_));
  OAI22_X1   g12656(.A1(new_n11369_), .A2(new_n6089_), .B1(new_n6091_), .B2(new_n11461_), .ZN(new_n12721_));
  NAND2_X1   g12657(.A1(new_n11694_), .A2(new_n6095_), .ZN(new_n12722_));
  AOI21_X1   g12658(.A1(new_n12721_), .A2(new_n12722_), .B(new_n6082_), .ZN(new_n12723_));
  NAND2_X1   g12659(.A1(new_n12720_), .A2(new_n12723_), .ZN(new_n12724_));
  XOR2_X1    g12660(.A1(new_n12724_), .A2(\a[14] ), .Z(new_n12725_));
  INV_X1     g12661(.I(new_n12725_), .ZN(new_n12726_));
  NOR2_X1    g12662(.A1(new_n12711_), .A2(new_n12726_), .ZN(new_n12727_));
  NOR2_X1    g12663(.A1(new_n12710_), .A2(new_n12725_), .ZN(new_n12728_));
  INV_X1     g12664(.I(new_n12728_), .ZN(new_n12729_));
  OAI21_X1   g12665(.A1(new_n12617_), .A2(new_n12727_), .B(new_n12729_), .ZN(new_n12730_));
  XNOR2_X1   g12666(.A1(new_n12730_), .A2(new_n12612_), .ZN(new_n12731_));
  INV_X1     g12667(.I(new_n12617_), .ZN(new_n12732_));
  OAI21_X1   g12668(.A1(new_n12727_), .A2(new_n12728_), .B(new_n12732_), .ZN(new_n12733_));
  NOR2_X1    g12669(.A1(new_n12710_), .A2(new_n12726_), .ZN(new_n12734_));
  NOR2_X1    g12670(.A1(new_n12711_), .A2(new_n12725_), .ZN(new_n12735_));
  OAI21_X1   g12671(.A1(new_n12735_), .A2(new_n12734_), .B(new_n12617_), .ZN(new_n12736_));
  NAND2_X1   g12672(.A1(new_n12733_), .A2(new_n12736_), .ZN(new_n12737_));
  NOR2_X1    g12673(.A1(new_n12695_), .A2(new_n12697_), .ZN(new_n12738_));
  NOR2_X1    g12674(.A1(new_n12738_), .A2(new_n12622_), .ZN(new_n12739_));
  XOR2_X1    g12675(.A1(new_n12687_), .A2(new_n12694_), .Z(new_n12740_));
  NOR3_X1    g12676(.A1(new_n12740_), .A2(new_n12619_), .A3(new_n12621_), .ZN(new_n12741_));
  OR2_X2     g12677(.A1(new_n12739_), .A2(new_n12741_), .Z(new_n12742_));
  NAND2_X1   g12678(.A1(new_n12624_), .A2(new_n12626_), .ZN(new_n12743_));
  INV_X1     g12679(.I(new_n12626_), .ZN(new_n12744_));
  OAI22_X1   g12680(.A1(new_n12686_), .A2(new_n12683_), .B1(new_n12744_), .B2(new_n12623_), .ZN(new_n12745_));
  OAI21_X1   g12681(.A1(new_n12676_), .A2(new_n12668_), .B(new_n12681_), .ZN(new_n12746_));
  NAND2_X1   g12682(.A1(new_n12685_), .A2(new_n12682_), .ZN(new_n12747_));
  AND2_X2    g12683(.A1(new_n12747_), .A2(new_n12746_), .Z(new_n12748_));
  OAI21_X1   g12684(.A1(new_n12748_), .A2(new_n12743_), .B(new_n12745_), .ZN(new_n12749_));
  INV_X1     g12685(.I(new_n12631_), .ZN(new_n12750_));
  OAI21_X1   g12686(.A1(new_n12433_), .A2(new_n12434_), .B(new_n12750_), .ZN(new_n12751_));
  INV_X1     g12687(.I(new_n12634_), .ZN(new_n12752_));
  NAND3_X1   g12688(.A1(new_n12630_), .A2(new_n12628_), .A3(new_n12752_), .ZN(new_n12753_));
  AOI22_X1   g12689(.A1(new_n12751_), .A2(new_n12753_), .B1(new_n12654_), .B2(new_n12660_), .ZN(new_n12754_));
  XOR2_X1    g12690(.A1(new_n12648_), .A2(new_n12653_), .Z(new_n12755_));
  AOI21_X1   g12691(.A1(new_n12636_), .A2(new_n12755_), .B(new_n12754_), .ZN(new_n12756_));
  XOR2_X1    g12692(.A1(new_n12658_), .A2(new_n12646_), .Z(new_n12757_));
  OAI21_X1   g12693(.A1(new_n12420_), .A2(new_n12421_), .B(new_n11913_), .ZN(new_n12758_));
  NAND3_X1   g12694(.A1(new_n11894_), .A2(new_n11898_), .A3(new_n12422_), .ZN(new_n12759_));
  AOI22_X1   g12695(.A1(new_n12758_), .A2(new_n12759_), .B1(new_n11863_), .B2(new_n11866_), .ZN(new_n12760_));
  NAND2_X1   g12696(.A1(new_n12424_), .A2(new_n11914_), .ZN(new_n12761_));
  AOI21_X1   g12697(.A1(new_n12417_), .A2(new_n12761_), .B(new_n12760_), .ZN(new_n12762_));
  NOR2_X1    g12698(.A1(new_n11865_), .A2(new_n12415_), .ZN(new_n12763_));
  AOI21_X1   g12699(.A1(new_n12413_), .A2(new_n12414_), .B(new_n12763_), .ZN(new_n12764_));
  AOI21_X1   g12700(.A1(new_n11781_), .A2(new_n11780_), .B(new_n11862_), .ZN(new_n12765_));
  NOR3_X1    g12701(.A1(new_n11785_), .A2(new_n11784_), .A3(new_n11864_), .ZN(new_n12766_));
  NOR2_X1    g12702(.A1(new_n12765_), .A2(new_n12766_), .ZN(new_n12767_));
  NOR3_X1    g12703(.A1(new_n11851_), .A2(new_n11853_), .A3(new_n12767_), .ZN(new_n12768_));
  NAND2_X1   g12704(.A1(new_n10909_), .A2(new_n10885_), .ZN(new_n12769_));
  NOR2_X1    g12705(.A1(new_n10877_), .A2(new_n10866_), .ZN(new_n12770_));
  XOR2_X1    g12706(.A1(new_n10885_), .A2(new_n10872_), .Z(new_n12771_));
  AOI21_X1   g12707(.A1(new_n12770_), .A2(new_n10886_), .B(new_n12771_), .ZN(new_n12772_));
  NAND3_X1   g12708(.A1(new_n12772_), .A2(new_n10892_), .A3(new_n12769_), .ZN(new_n12773_));
  AOI21_X1   g12709(.A1(new_n12772_), .A2(new_n12769_), .B(new_n10892_), .ZN(new_n12774_));
  INV_X1     g12710(.I(new_n12774_), .ZN(new_n12775_));
  NAND2_X1   g12711(.A1(new_n12775_), .A2(new_n12773_), .ZN(new_n12776_));
  INV_X1     g12712(.I(new_n12776_), .ZN(new_n12777_));
  NOR2_X1    g12713(.A1(new_n10892_), .A2(new_n2772_), .ZN(new_n12778_));
  NOR2_X1    g12714(.A1(new_n10885_), .A2(new_n2767_), .ZN(new_n12779_));
  AOI21_X1   g12715(.A1(new_n10872_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n12780_));
  INV_X1     g12716(.I(new_n12780_), .ZN(new_n12781_));
  NOR4_X1    g12717(.A1(new_n12777_), .A2(new_n12778_), .A3(new_n12779_), .A4(new_n12781_), .ZN(new_n12782_));
  NOR3_X1    g12718(.A1(new_n12768_), .A2(new_n12764_), .A3(new_n12782_), .ZN(new_n12783_));
  OAI21_X1   g12719(.A1(new_n12768_), .A2(new_n12764_), .B(new_n12782_), .ZN(new_n12784_));
  OAI22_X1   g12720(.A1(new_n11850_), .A2(new_n11853_), .B1(new_n12411_), .B2(new_n11828_), .ZN(new_n12785_));
  AOI21_X1   g12721(.A1(new_n11782_), .A2(new_n11826_), .B(new_n11828_), .ZN(new_n12786_));
  OAI21_X1   g12722(.A1(new_n11785_), .A2(new_n11784_), .B(new_n11852_), .ZN(new_n12787_));
  NAND3_X1   g12723(.A1(new_n11781_), .A2(new_n11780_), .A3(new_n11849_), .ZN(new_n12788_));
  NAND2_X1   g12724(.A1(new_n12787_), .A2(new_n12788_), .ZN(new_n12789_));
  NAND2_X1   g12725(.A1(new_n12789_), .A2(new_n12786_), .ZN(new_n12790_));
  NAND2_X1   g12726(.A1(new_n12790_), .A2(new_n12785_), .ZN(new_n12791_));
  AOI22_X1   g12727(.A1(new_n11781_), .A2(new_n11780_), .B1(new_n11826_), .B2(new_n11829_), .ZN(new_n12792_));
  XNOR2_X1   g12728(.A1(new_n11798_), .A2(new_n11825_), .ZN(new_n12793_));
  NOR3_X1    g12729(.A1(new_n11785_), .A2(new_n11784_), .A3(new_n12793_), .ZN(new_n12794_));
  INV_X1     g12730(.I(new_n1142_), .ZN(new_n12795_));
  INV_X1     g12731(.I(new_n2057_), .ZN(new_n12796_));
  NAND4_X1   g12732(.A1(new_n2113_), .A2(new_n2125_), .A3(new_n389_), .A4(new_n716_), .ZN(new_n12797_));
  NOR2_X1    g12733(.A1(new_n12796_), .A2(new_n12797_), .ZN(new_n12798_));
  INV_X1     g12734(.I(new_n12798_), .ZN(new_n12799_));
  NOR3_X1    g12735(.A1(new_n267_), .A2(new_n734_), .A3(new_n596_), .ZN(new_n12800_));
  NAND4_X1   g12736(.A1(new_n12800_), .A2(new_n246_), .A3(new_n272_), .A4(new_n3104_), .ZN(new_n12801_));
  NOR4_X1    g12737(.A1(new_n495_), .A2(new_n656_), .A3(new_n406_), .A4(new_n749_), .ZN(new_n12802_));
  NOR3_X1    g12738(.A1(new_n1988_), .A2(new_n366_), .A3(new_n486_), .ZN(new_n12803_));
  NAND4_X1   g12739(.A1(new_n12802_), .A2(new_n12803_), .A3(new_n4760_), .A4(new_n2970_), .ZN(new_n12804_));
  NOR4_X1    g12740(.A1(new_n12799_), .A2(new_n12091_), .A3(new_n12801_), .A4(new_n12804_), .ZN(new_n12805_));
  INV_X1     g12741(.I(new_n12805_), .ZN(new_n12806_));
  NOR3_X1    g12742(.A1(new_n12806_), .A2(new_n12795_), .A3(new_n3692_), .ZN(new_n12807_));
  INV_X1     g12743(.I(new_n12807_), .ZN(new_n12808_));
  NOR2_X1    g12744(.A1(new_n10865_), .A2(new_n8785_), .ZN(new_n12809_));
  OAI21_X1   g12745(.A1(new_n11790_), .A2(new_n12809_), .B(new_n8779_), .ZN(new_n12810_));
  NOR2_X1    g12746(.A1(new_n10875_), .A2(new_n8785_), .ZN(new_n12811_));
  NOR2_X1    g12747(.A1(new_n10865_), .A2(new_n8784_), .ZN(new_n12812_));
  OAI21_X1   g12748(.A1(new_n12811_), .A2(new_n12812_), .B(new_n8778_), .ZN(new_n12813_));
  NAND2_X1   g12749(.A1(new_n12810_), .A2(new_n12813_), .ZN(new_n12814_));
  NAND2_X1   g12750(.A1(new_n8779_), .A2(new_n3332_), .ZN(new_n12815_));
  NAND2_X1   g12751(.A1(new_n8785_), .A2(new_n3189_), .ZN(new_n12816_));
  AOI21_X1   g12752(.A1(new_n10862_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n12817_));
  NAND4_X1   g12753(.A1(new_n12814_), .A2(new_n12815_), .A3(new_n12816_), .A4(new_n12817_), .ZN(new_n12818_));
  XOR2_X1    g12754(.A1(new_n12818_), .A2(new_n12807_), .Z(new_n12819_));
  INV_X1     g12755(.I(new_n12819_), .ZN(new_n12820_));
  OAI21_X1   g12756(.A1(new_n10773_), .A2(new_n10772_), .B(new_n9530_), .ZN(new_n12821_));
  NAND3_X1   g12757(.A1(new_n10753_), .A2(new_n10770_), .A3(new_n9531_), .ZN(new_n12822_));
  NAND2_X1   g12758(.A1(new_n12821_), .A2(new_n12822_), .ZN(new_n12823_));
  NAND3_X1   g12759(.A1(new_n10792_), .A2(new_n10791_), .A3(new_n10788_), .ZN(new_n12824_));
  OAI21_X1   g12760(.A1(new_n10783_), .A2(new_n10787_), .B(new_n10789_), .ZN(new_n12825_));
  NAND2_X1   g12761(.A1(new_n12825_), .A2(new_n12824_), .ZN(new_n12826_));
  NAND3_X1   g12762(.A1(new_n12826_), .A2(new_n12823_), .A3(new_n10777_), .ZN(new_n12827_));
  AOI21_X1   g12763(.A1(new_n12826_), .A2(new_n12823_), .B(new_n10777_), .ZN(new_n12828_));
  INV_X1     g12764(.I(new_n12828_), .ZN(new_n12829_));
  NAND2_X1   g12765(.A1(new_n12829_), .A2(new_n12827_), .ZN(new_n12830_));
  OAI22_X1   g12766(.A1(new_n12826_), .A2(new_n2771_), .B1(new_n2767_), .B2(new_n10775_), .ZN(new_n12831_));
  NAND2_X1   g12767(.A1(new_n10800_), .A2(new_n3332_), .ZN(new_n12832_));
  AOI21_X1   g12768(.A1(new_n12831_), .A2(new_n12832_), .B(new_n2763_), .ZN(new_n12833_));
  NAND2_X1   g12769(.A1(new_n12830_), .A2(new_n12833_), .ZN(new_n12834_));
  NAND4_X1   g12770(.A1(new_n1404_), .A2(new_n266_), .A3(new_n1009_), .A4(new_n773_), .ZN(new_n12835_));
  NAND4_X1   g12771(.A1(new_n3877_), .A2(new_n193_), .A3(new_n806_), .A4(new_n12835_), .ZN(new_n12836_));
  NOR2_X1    g12772(.A1(new_n555_), .A2(new_n1134_), .ZN(new_n12837_));
  NOR3_X1    g12773(.A1(new_n2338_), .A2(new_n584_), .A3(new_n796_), .ZN(new_n12838_));
  NOR3_X1    g12774(.A1(new_n936_), .A2(new_n261_), .A3(new_n305_), .ZN(new_n12839_));
  NAND4_X1   g12775(.A1(new_n12837_), .A2(new_n1265_), .A3(new_n12838_), .A4(new_n12839_), .ZN(new_n12840_));
  NOR3_X1    g12776(.A1(new_n12836_), .A2(new_n12840_), .A3(new_n11814_), .ZN(new_n12841_));
  NAND3_X1   g12777(.A1(new_n12156_), .A2(new_n11729_), .A3(new_n12841_), .ZN(new_n12842_));
  NOR2_X1    g12778(.A1(new_n12834_), .A2(new_n12842_), .ZN(new_n12843_));
  OAI22_X1   g12779(.A1(new_n12826_), .A2(new_n2767_), .B1(new_n2772_), .B2(new_n10775_), .ZN(new_n12844_));
  NAND2_X1   g12780(.A1(new_n12826_), .A2(new_n10775_), .ZN(new_n12845_));
  NAND2_X1   g12781(.A1(new_n10794_), .A2(new_n12823_), .ZN(new_n12846_));
  NAND2_X1   g12782(.A1(new_n12846_), .A2(new_n12845_), .ZN(new_n12847_));
  OAI21_X1   g12783(.A1(new_n12847_), .A2(new_n2763_), .B(new_n12844_), .ZN(new_n12848_));
  NOR4_X1    g12784(.A1(new_n666_), .A2(new_n625_), .A3(new_n752_), .A4(new_n418_), .ZN(new_n12849_));
  NOR3_X1    g12785(.A1(new_n1498_), .A2(new_n1157_), .A3(new_n12849_), .ZN(new_n12850_));
  NAND3_X1   g12786(.A1(new_n3221_), .A2(new_n2632_), .A3(new_n12850_), .ZN(new_n12851_));
  INV_X1     g12787(.I(new_n2380_), .ZN(new_n12852_));
  NAND2_X1   g12788(.A1(new_n1892_), .A2(new_n872_), .ZN(new_n12853_));
  NAND3_X1   g12789(.A1(new_n2046_), .A2(new_n434_), .A3(new_n3198_), .ZN(new_n12854_));
  NOR4_X1    g12790(.A1(new_n12854_), .A2(new_n488_), .A3(new_n12852_), .A4(new_n12853_), .ZN(new_n12855_));
  NOR4_X1    g12791(.A1(new_n458_), .A2(new_n569_), .A3(new_n422_), .A4(new_n1076_), .ZN(new_n12856_));
  NOR4_X1    g12792(.A1(new_n170_), .A2(new_n955_), .A3(new_n227_), .A4(new_n310_), .ZN(new_n12857_));
  INV_X1     g12793(.I(new_n12857_), .ZN(new_n12858_));
  NAND4_X1   g12794(.A1(new_n12855_), .A2(new_n2691_), .A3(new_n12856_), .A4(new_n12858_), .ZN(new_n12859_));
  NOR2_X1    g12795(.A1(new_n12859_), .A2(new_n12851_), .ZN(new_n12860_));
  INV_X1     g12796(.I(new_n12860_), .ZN(new_n12861_));
  NAND3_X1   g12797(.A1(new_n797_), .A2(new_n250_), .A3(new_n1638_), .ZN(new_n12862_));
  NAND3_X1   g12798(.A1(new_n2341_), .A2(new_n272_), .A3(new_n707_), .ZN(new_n12863_));
  NOR4_X1    g12799(.A1(new_n12863_), .A2(new_n12862_), .A3(new_n1389_), .A4(new_n1620_), .ZN(new_n12864_));
  NOR3_X1    g12800(.A1(new_n2088_), .A2(new_n2133_), .A3(new_n2134_), .ZN(new_n12865_));
  NOR2_X1    g12801(.A1(new_n2143_), .A2(new_n2594_), .ZN(new_n12866_));
  NAND4_X1   g12802(.A1(new_n4820_), .A2(new_n12864_), .A3(new_n12865_), .A4(new_n12866_), .ZN(new_n12867_));
  NOR3_X1    g12803(.A1(new_n12861_), .A2(new_n1568_), .A3(new_n12867_), .ZN(new_n12868_));
  INV_X1     g12804(.I(new_n12868_), .ZN(new_n12869_));
  NAND2_X1   g12805(.A1(new_n12848_), .A2(new_n12869_), .ZN(new_n12870_));
  NAND2_X1   g12806(.A1(new_n12834_), .A2(new_n12842_), .ZN(new_n12871_));
  AOI21_X1   g12807(.A1(new_n12870_), .A2(new_n12871_), .B(new_n12843_), .ZN(new_n12872_));
  NAND3_X1   g12808(.A1(new_n12825_), .A2(new_n12824_), .A3(new_n10800_), .ZN(new_n12873_));
  OAI21_X1   g12809(.A1(new_n10774_), .A2(new_n10771_), .B(new_n10777_), .ZN(new_n12874_));
  NAND3_X1   g12810(.A1(new_n12821_), .A2(new_n10800_), .A3(new_n12822_), .ZN(new_n12875_));
  NAND2_X1   g12811(.A1(new_n12875_), .A2(new_n12874_), .ZN(new_n12876_));
  NAND3_X1   g12812(.A1(new_n12876_), .A2(new_n12873_), .A3(new_n10798_), .ZN(new_n12877_));
  NOR3_X1    g12813(.A1(new_n10790_), .A2(new_n10793_), .A3(new_n10777_), .ZN(new_n12878_));
  AOI21_X1   g12814(.A1(new_n12821_), .A2(new_n12822_), .B(new_n10800_), .ZN(new_n12879_));
  NOR3_X1    g12815(.A1(new_n10774_), .A2(new_n10771_), .A3(new_n10777_), .ZN(new_n12880_));
  NOR2_X1    g12816(.A1(new_n12879_), .A2(new_n12880_), .ZN(new_n12881_));
  OAI21_X1   g12817(.A1(new_n12881_), .A2(new_n12878_), .B(new_n9529_), .ZN(new_n12882_));
  NAND2_X1   g12818(.A1(new_n12882_), .A2(new_n12877_), .ZN(new_n12883_));
  NAND2_X1   g12819(.A1(new_n12823_), .A2(new_n2770_), .ZN(new_n12884_));
  NAND2_X1   g12820(.A1(new_n9529_), .A2(new_n3332_), .ZN(new_n12885_));
  AOI21_X1   g12821(.A1(new_n10800_), .A2(new_n3189_), .B(new_n2763_), .ZN(new_n12886_));
  NAND4_X1   g12822(.A1(new_n12883_), .A2(new_n12884_), .A3(new_n12885_), .A4(new_n12886_), .ZN(new_n12887_));
  INV_X1     g12823(.I(new_n11094_), .ZN(new_n12888_));
  NAND4_X1   g12824(.A1(new_n4925_), .A2(new_n2637_), .A3(new_n1173_), .A4(new_n1843_), .ZN(new_n12889_));
  NOR2_X1    g12825(.A1(new_n1487_), .A2(new_n530_), .ZN(new_n12890_));
  NAND4_X1   g12826(.A1(new_n1658_), .A2(new_n1315_), .A3(new_n351_), .A4(new_n1009_), .ZN(new_n12891_));
  NAND4_X1   g12827(.A1(new_n12890_), .A2(new_n1835_), .A3(new_n2996_), .A4(new_n12891_), .ZN(new_n12892_));
  NOR3_X1    g12828(.A1(new_n12889_), .A2(new_n3996_), .A3(new_n12892_), .ZN(new_n12893_));
  NAND4_X1   g12829(.A1(new_n2966_), .A2(new_n12893_), .A3(new_n11066_), .A4(new_n12888_), .ZN(new_n12894_));
  NAND2_X1   g12830(.A1(new_n12887_), .A2(new_n12894_), .ZN(new_n12895_));
  INV_X1     g12831(.I(new_n12895_), .ZN(new_n12896_));
  NOR2_X1    g12832(.A1(new_n12887_), .A2(new_n12894_), .ZN(new_n12897_));
  INV_X1     g12833(.I(new_n12897_), .ZN(new_n12898_));
  OAI21_X1   g12834(.A1(new_n12872_), .A2(new_n12896_), .B(new_n12898_), .ZN(new_n12899_));
  OAI21_X1   g12835(.A1(new_n10774_), .A2(new_n10771_), .B(new_n9529_), .ZN(new_n12900_));
  OAI21_X1   g12836(.A1(new_n12826_), .A2(new_n12900_), .B(new_n10777_), .ZN(new_n12901_));
  AOI21_X1   g12837(.A1(new_n12901_), .A2(new_n10799_), .B(new_n10798_), .ZN(new_n12902_));
  OAI21_X1   g12838(.A1(new_n12902_), .A2(new_n10795_), .B(new_n10839_), .ZN(new_n12903_));
  AOI21_X1   g12839(.A1(new_n12823_), .A2(new_n10800_), .B(new_n9529_), .ZN(new_n12904_));
  NOR2_X1    g12840(.A1(new_n12823_), .A2(new_n9529_), .ZN(new_n12905_));
  AOI21_X1   g12841(.A1(new_n12821_), .A2(new_n12822_), .B(new_n10798_), .ZN(new_n12906_));
  AOI21_X1   g12842(.A1(new_n10794_), .A2(new_n12906_), .B(new_n10800_), .ZN(new_n12907_));
  NOR3_X1    g12843(.A1(new_n12907_), .A2(new_n10798_), .A3(new_n12905_), .ZN(new_n12908_));
  OAI21_X1   g12844(.A1(new_n12908_), .A2(new_n12904_), .B(new_n10844_), .ZN(new_n12909_));
  NAND2_X1   g12845(.A1(new_n12909_), .A2(new_n12903_), .ZN(new_n12910_));
  NAND2_X1   g12846(.A1(new_n9529_), .A2(new_n3189_), .ZN(new_n12911_));
  NAND2_X1   g12847(.A1(new_n10839_), .A2(new_n3332_), .ZN(new_n12912_));
  AOI21_X1   g12848(.A1(new_n10800_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n12913_));
  NAND4_X1   g12849(.A1(new_n12910_), .A2(new_n12911_), .A3(new_n12912_), .A4(new_n12913_), .ZN(new_n12914_));
  INV_X1     g12850(.I(new_n11551_), .ZN(new_n12915_));
  NOR4_X1    g12851(.A1(new_n12915_), .A2(new_n490_), .A3(new_n561_), .A4(new_n744_), .ZN(new_n12916_));
  NOR4_X1    g12852(.A1(new_n135_), .A2(new_n603_), .A3(new_n487_), .A4(new_n594_), .ZN(new_n12917_));
  NAND4_X1   g12853(.A1(new_n2975_), .A2(new_n12917_), .A3(new_n358_), .A4(new_n592_), .ZN(new_n12918_));
  NOR4_X1    g12854(.A1(new_n12918_), .A2(new_n576_), .A3(new_n769_), .A4(new_n1076_), .ZN(new_n12919_));
  NOR4_X1    g12855(.A1(new_n251_), .A2(new_n147_), .A3(new_n164_), .A4(new_n330_), .ZN(new_n12920_));
  NOR4_X1    g12856(.A1(new_n573_), .A2(new_n424_), .A3(new_n70_), .A4(new_n753_), .ZN(new_n12921_));
  NOR3_X1    g12857(.A1(new_n11926_), .A2(new_n12920_), .A3(new_n12921_), .ZN(new_n12922_));
  NAND4_X1   g12858(.A1(new_n12919_), .A2(new_n12161_), .A3(new_n12922_), .A4(new_n12916_), .ZN(new_n12923_));
  INV_X1     g12859(.I(new_n12923_), .ZN(new_n12924_));
  NOR3_X1    g12860(.A1(new_n98_), .A2(new_n252_), .A3(new_n611_), .ZN(new_n12925_));
  NOR4_X1    g12861(.A1(new_n615_), .A2(new_n172_), .A3(new_n235_), .A4(new_n191_), .ZN(new_n12926_));
  NAND2_X1   g12862(.A1(new_n12926_), .A2(new_n12925_), .ZN(new_n12927_));
  NOR2_X1    g12863(.A1(new_n1245_), .A2(new_n2041_), .ZN(new_n12928_));
  NAND4_X1   g12864(.A1(new_n926_), .A2(new_n327_), .A3(new_n3662_), .A4(new_n12928_), .ZN(new_n12929_));
  NOR4_X1    g12865(.A1(new_n12929_), .A2(new_n1672_), .A3(new_n1622_), .A4(new_n12927_), .ZN(new_n12930_));
  NAND3_X1   g12866(.A1(new_n1428_), .A2(new_n12924_), .A3(new_n12930_), .ZN(new_n12931_));
  NAND2_X1   g12867(.A1(new_n12914_), .A2(new_n12931_), .ZN(new_n12932_));
  NAND2_X1   g12868(.A1(new_n12899_), .A2(new_n12932_), .ZN(new_n12933_));
  OR2_X2     g12869(.A1(new_n12914_), .A2(new_n12931_), .Z(new_n12934_));
  NAND2_X1   g12870(.A1(new_n12933_), .A2(new_n12934_), .ZN(new_n12935_));
  INV_X1     g12871(.I(new_n10846_), .ZN(new_n12936_));
  NAND4_X1   g12872(.A1(new_n12823_), .A2(new_n12825_), .A3(new_n12824_), .A4(new_n9529_), .ZN(new_n12937_));
  AOI21_X1   g12873(.A1(new_n12937_), .A2(new_n10777_), .B(new_n12905_), .ZN(new_n12938_));
  NOR3_X1    g12874(.A1(new_n12938_), .A2(new_n10798_), .A3(new_n10839_), .ZN(new_n12939_));
  INV_X1     g12875(.I(new_n10795_), .ZN(new_n12940_));
  NOR2_X1    g12876(.A1(new_n10844_), .A2(new_n12940_), .ZN(new_n12941_));
  OAI21_X1   g12877(.A1(new_n12939_), .A2(new_n12941_), .B(new_n12936_), .ZN(new_n12942_));
  OAI21_X1   g12878(.A1(new_n12938_), .A2(new_n10798_), .B(new_n10844_), .ZN(new_n12943_));
  NAND2_X1   g12879(.A1(new_n10839_), .A2(new_n12940_), .ZN(new_n12944_));
  AND2_X2    g12880(.A1(new_n12943_), .A2(new_n12944_), .Z(new_n12945_));
  OAI21_X1   g12881(.A1(new_n12945_), .A2(new_n12936_), .B(new_n12942_), .ZN(new_n12946_));
  NAND2_X1   g12882(.A1(new_n10839_), .A2(new_n3189_), .ZN(new_n12947_));
  NAND2_X1   g12883(.A1(new_n9529_), .A2(new_n2770_), .ZN(new_n12948_));
  OAI21_X1   g12884(.A1(new_n12936_), .A2(\a[31] ), .B(new_n2762_), .ZN(new_n12949_));
  NAND4_X1   g12885(.A1(new_n12946_), .A2(new_n12947_), .A3(new_n12948_), .A4(new_n12949_), .ZN(new_n12950_));
  INV_X1     g12886(.I(new_n3095_), .ZN(new_n12951_));
  NOR4_X1    g12887(.A1(new_n211_), .A2(new_n294_), .A3(new_n403_), .A4(new_n468_), .ZN(new_n12952_));
  NOR3_X1    g12888(.A1(new_n12951_), .A2(new_n3199_), .A3(new_n12952_), .ZN(new_n12953_));
  NOR4_X1    g12889(.A1(new_n1337_), .A2(new_n2234_), .A3(new_n190_), .A4(new_n604_), .ZN(new_n12954_));
  NOR4_X1    g12890(.A1(new_n3990_), .A2(new_n127_), .A3(new_n161_), .A4(new_n1185_), .ZN(new_n12955_));
  NAND4_X1   g12891(.A1(new_n1253_), .A2(new_n12953_), .A3(new_n12954_), .A4(new_n12955_), .ZN(new_n12956_));
  NOR2_X1    g12892(.A1(new_n12956_), .A2(new_n12027_), .ZN(new_n12957_));
  INV_X1     g12893(.I(new_n1575_), .ZN(new_n12958_));
  NOR4_X1    g12894(.A1(new_n12958_), .A2(new_n647_), .A3(new_n1045_), .A4(new_n4749_), .ZN(new_n12959_));
  NAND4_X1   g12895(.A1(new_n1816_), .A2(new_n429_), .A3(new_n1585_), .A4(new_n1638_), .ZN(new_n12960_));
  NOR3_X1    g12896(.A1(new_n225_), .A2(new_n1167_), .A3(new_n163_), .ZN(new_n12961_));
  NAND4_X1   g12897(.A1(new_n12959_), .A2(new_n2226_), .A3(new_n12960_), .A4(new_n12961_), .ZN(new_n12962_));
  NOR2_X1    g12898(.A1(new_n3084_), .A2(new_n12962_), .ZN(new_n12963_));
  NAND3_X1   g12899(.A1(new_n12957_), .A2(new_n11213_), .A3(new_n12963_), .ZN(new_n12964_));
  NAND2_X1   g12900(.A1(new_n12950_), .A2(new_n12964_), .ZN(new_n12965_));
  NOR2_X1    g12901(.A1(new_n12950_), .A2(new_n12964_), .ZN(new_n12966_));
  AOI21_X1   g12902(.A1(new_n12935_), .A2(new_n12965_), .B(new_n12966_), .ZN(new_n12967_));
  NAND2_X1   g12903(.A1(new_n12943_), .A2(new_n12944_), .ZN(new_n12968_));
  OAI21_X1   g12904(.A1(new_n10840_), .A2(new_n10795_), .B(new_n10846_), .ZN(new_n12969_));
  OAI21_X1   g12905(.A1(new_n12938_), .A2(new_n10798_), .B(new_n10844_), .ZN(new_n12970_));
  NAND3_X1   g12906(.A1(new_n12970_), .A2(new_n12940_), .A3(new_n12936_), .ZN(new_n12971_));
  NAND4_X1   g12907(.A1(new_n12969_), .A2(new_n12971_), .A3(new_n12968_), .A4(new_n9478_), .ZN(new_n12972_));
  NAND3_X1   g12908(.A1(new_n12969_), .A2(new_n12971_), .A3(new_n12968_), .ZN(new_n12973_));
  NAND2_X1   g12909(.A1(new_n12973_), .A2(new_n9479_), .ZN(new_n12974_));
  NAND2_X1   g12910(.A1(new_n12974_), .A2(new_n12972_), .ZN(new_n12975_));
  NAND2_X1   g12911(.A1(new_n10839_), .A2(new_n2770_), .ZN(new_n12976_));
  NAND2_X1   g12912(.A1(new_n9479_), .A2(new_n3332_), .ZN(new_n12977_));
  AOI21_X1   g12913(.A1(new_n12936_), .A2(new_n3189_), .B(new_n2764_), .ZN(new_n12978_));
  NAND4_X1   g12914(.A1(new_n12975_), .A2(new_n12976_), .A3(new_n12977_), .A4(new_n12978_), .ZN(new_n12979_));
  NOR3_X1    g12915(.A1(new_n1048_), .A2(new_n637_), .A3(new_n241_), .ZN(new_n12980_));
  NOR3_X1    g12916(.A1(new_n1984_), .A2(new_n149_), .A3(new_n264_), .ZN(new_n12981_));
  NAND4_X1   g12917(.A1(new_n360_), .A2(new_n271_), .A3(new_n1647_), .A4(new_n872_), .ZN(new_n12982_));
  NAND4_X1   g12918(.A1(new_n1366_), .A2(new_n12980_), .A3(new_n12981_), .A4(new_n12982_), .ZN(new_n12983_));
  NAND4_X1   g12919(.A1(new_n2974_), .A2(new_n1153_), .A3(new_n1416_), .A4(new_n3365_), .ZN(new_n12984_));
  NOR3_X1    g12920(.A1(new_n12984_), .A2(new_n4791_), .A3(new_n12983_), .ZN(new_n12985_));
  INV_X1     g12921(.I(new_n2679_), .ZN(new_n12986_));
  NAND4_X1   g12922(.A1(new_n233_), .A2(new_n701_), .A3(new_n435_), .A4(new_n395_), .ZN(new_n12987_));
  NAND4_X1   g12923(.A1(new_n11923_), .A2(new_n3948_), .A3(new_n4844_), .A4(new_n12987_), .ZN(new_n12988_));
  NOR3_X1    g12924(.A1(new_n2065_), .A2(new_n177_), .A3(new_n618_), .ZN(new_n12989_));
  NAND4_X1   g12925(.A1(new_n2683_), .A2(new_n12989_), .A3(new_n507_), .A4(new_n987_), .ZN(new_n12990_));
  NOR3_X1    g12926(.A1(new_n12988_), .A2(new_n12990_), .A3(new_n12986_), .ZN(new_n12991_));
  NAND2_X1   g12927(.A1(new_n1214_), .A2(new_n2835_), .ZN(new_n12992_));
  NAND4_X1   g12928(.A1(new_n1254_), .A2(new_n313_), .A3(new_n414_), .A4(new_n1156_), .ZN(new_n12993_));
  NAND2_X1   g12929(.A1(new_n6525_), .A2(new_n1781_), .ZN(new_n12994_));
  NOR4_X1    g12930(.A1(new_n12994_), .A2(new_n1914_), .A3(new_n12992_), .A4(new_n12993_), .ZN(new_n12995_));
  NAND2_X1   g12931(.A1(new_n1953_), .A2(new_n1952_), .ZN(new_n12996_));
  INV_X1     g12932(.I(new_n12521_), .ZN(new_n12997_));
  NOR4_X1    g12933(.A1(new_n437_), .A2(new_n1031_), .A3(new_n955_), .A4(new_n329_), .ZN(new_n12998_));
  NOR4_X1    g12934(.A1(new_n1084_), .A2(new_n370_), .A3(new_n374_), .A4(new_n591_), .ZN(new_n12999_));
  NOR4_X1    g12935(.A1(new_n12997_), .A2(new_n12996_), .A3(new_n12998_), .A4(new_n12999_), .ZN(new_n13000_));
  NAND4_X1   g12936(.A1(new_n13000_), .A2(new_n12985_), .A3(new_n12995_), .A4(new_n12991_), .ZN(new_n13001_));
  NAND2_X1   g12937(.A1(new_n12979_), .A2(new_n13001_), .ZN(new_n13002_));
  INV_X1     g12938(.I(new_n13002_), .ZN(new_n13003_));
  OR2_X2     g12939(.A1(new_n12979_), .A2(new_n13001_), .Z(new_n13004_));
  OAI21_X1   g12940(.A1(new_n12967_), .A2(new_n13003_), .B(new_n13004_), .ZN(new_n13005_));
  NAND2_X1   g12941(.A1(new_n12970_), .A2(new_n12940_), .ZN(new_n13006_));
  INV_X1     g12942(.I(new_n10847_), .ZN(new_n13007_));
  INV_X1     g12943(.I(new_n10848_), .ZN(new_n13008_));
  OAI21_X1   g12944(.A1(new_n13006_), .A2(new_n13007_), .B(new_n13008_), .ZN(new_n13009_));
  NAND2_X1   g12945(.A1(new_n13009_), .A2(new_n9478_), .ZN(new_n13010_));
  NAND2_X1   g12946(.A1(new_n10849_), .A2(new_n9479_), .ZN(new_n13011_));
  AOI21_X1   g12947(.A1(new_n13011_), .A2(new_n13010_), .B(new_n10853_), .ZN(new_n13012_));
  NAND2_X1   g12948(.A1(new_n10849_), .A2(new_n9478_), .ZN(new_n13013_));
  NAND2_X1   g12949(.A1(new_n13009_), .A2(new_n9479_), .ZN(new_n13014_));
  AOI21_X1   g12950(.A1(new_n13013_), .A2(new_n13014_), .B(new_n10854_), .ZN(new_n13015_));
  OR2_X2     g12951(.A1(new_n13012_), .A2(new_n13015_), .Z(new_n13016_));
  NOR2_X1    g12952(.A1(new_n10853_), .A2(new_n2772_), .ZN(new_n13017_));
  NOR2_X1    g12953(.A1(new_n9478_), .A2(new_n2767_), .ZN(new_n13018_));
  NOR2_X1    g12954(.A1(new_n10846_), .A2(new_n2771_), .ZN(new_n13019_));
  NOR4_X1    g12955(.A1(new_n13018_), .A2(new_n2763_), .A3(new_n13017_), .A4(new_n13019_), .ZN(new_n13020_));
  NAND2_X1   g12956(.A1(new_n13016_), .A2(new_n13020_), .ZN(new_n13021_));
  INV_X1     g12957(.I(new_n559_), .ZN(new_n13022_));
  NAND3_X1   g12958(.A1(new_n2175_), .A2(new_n612_), .A3(new_n1068_), .ZN(new_n13023_));
  NAND4_X1   g12959(.A1(new_n295_), .A2(new_n1601_), .A3(new_n1393_), .A4(new_n984_), .ZN(new_n13024_));
  NAND4_X1   g12960(.A1(new_n13023_), .A2(new_n13024_), .A3(new_n1430_), .A4(new_n4844_), .ZN(new_n13025_));
  NAND4_X1   g12961(.A1(new_n12850_), .A2(new_n688_), .A3(new_n720_), .A4(new_n2191_), .ZN(new_n13026_));
  NOR4_X1    g12962(.A1(new_n2993_), .A2(new_n13026_), .A3(new_n13022_), .A4(new_n13025_), .ZN(new_n13027_));
  NAND3_X1   g12963(.A1(new_n2878_), .A2(new_n13027_), .A3(new_n2890_), .ZN(new_n13028_));
  NAND2_X1   g12964(.A1(new_n13021_), .A2(new_n13028_), .ZN(new_n13029_));
  NAND2_X1   g12965(.A1(new_n13005_), .A2(new_n13029_), .ZN(new_n13030_));
  OR2_X2     g12966(.A1(new_n13021_), .A2(new_n13028_), .Z(new_n13031_));
  NAND2_X1   g12967(.A1(new_n13030_), .A2(new_n13031_), .ZN(new_n13032_));
  NOR3_X1    g12968(.A1(new_n13009_), .A2(new_n9478_), .A3(new_n10854_), .ZN(new_n13033_));
  INV_X1     g12969(.I(new_n13033_), .ZN(new_n13034_));
  NAND3_X1   g12970(.A1(new_n13009_), .A2(new_n9478_), .A3(new_n10854_), .ZN(new_n13035_));
  AOI21_X1   g12971(.A1(new_n13034_), .A2(new_n13035_), .B(new_n10861_), .ZN(new_n13036_));
  AOI21_X1   g12972(.A1(new_n13009_), .A2(new_n9478_), .B(new_n10853_), .ZN(new_n13037_));
  AOI21_X1   g12973(.A1(new_n10849_), .A2(new_n9479_), .B(new_n10854_), .ZN(new_n13038_));
  OAI21_X1   g12974(.A1(new_n13038_), .A2(new_n13037_), .B(new_n10861_), .ZN(new_n13039_));
  INV_X1     g12975(.I(new_n13039_), .ZN(new_n13040_));
  AOI21_X1   g12976(.A1(new_n9479_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n13041_));
  OAI21_X1   g12977(.A1(new_n2767_), .A2(new_n10853_), .B(new_n13041_), .ZN(new_n13042_));
  AOI21_X1   g12978(.A1(new_n3332_), .A2(new_n10862_), .B(new_n13042_), .ZN(new_n13043_));
  OAI21_X1   g12979(.A1(new_n13040_), .A2(new_n13036_), .B(new_n13043_), .ZN(new_n13044_));
  NAND2_X1   g12980(.A1(new_n1430_), .A2(new_n1828_), .ZN(new_n13045_));
  NOR3_X1    g12981(.A1(new_n2677_), .A2(new_n496_), .A3(new_n541_), .ZN(new_n13046_));
  NOR3_X1    g12982(.A1(new_n3353_), .A2(new_n615_), .A3(new_n247_), .ZN(new_n13047_));
  NOR3_X1    g12983(.A1(new_n1461_), .A2(new_n226_), .A3(new_n644_), .ZN(new_n13048_));
  NOR3_X1    g12984(.A1(new_n225_), .A2(new_n695_), .A3(new_n731_), .ZN(new_n13049_));
  NAND4_X1   g12985(.A1(new_n13046_), .A2(new_n13048_), .A3(new_n13047_), .A4(new_n13049_), .ZN(new_n13050_));
  NOR4_X1    g12986(.A1(new_n13050_), .A2(new_n1870_), .A3(new_n12266_), .A4(new_n13045_), .ZN(new_n13051_));
  NAND3_X1   g12987(.A1(new_n11811_), .A2(new_n2296_), .A3(new_n13051_), .ZN(new_n13052_));
  NAND2_X1   g12988(.A1(new_n13044_), .A2(new_n13052_), .ZN(new_n13053_));
  NAND2_X1   g12989(.A1(new_n13032_), .A2(new_n13053_), .ZN(new_n13054_));
  NOR2_X1    g12990(.A1(new_n13044_), .A2(new_n13052_), .ZN(new_n13055_));
  INV_X1     g12991(.I(new_n13055_), .ZN(new_n13056_));
  NAND2_X1   g12992(.A1(new_n13054_), .A2(new_n13056_), .ZN(new_n13057_));
  NOR2_X1    g12993(.A1(new_n13038_), .A2(new_n13037_), .ZN(new_n13058_));
  OAI21_X1   g12994(.A1(new_n13009_), .A2(new_n9478_), .B(new_n10853_), .ZN(new_n13059_));
  AOI21_X1   g12995(.A1(new_n13059_), .A2(new_n13010_), .B(new_n10862_), .ZN(new_n13060_));
  NOR3_X1    g12996(.A1(new_n10855_), .A2(new_n10850_), .A3(new_n10861_), .ZN(new_n13061_));
  NOR4_X1    g12997(.A1(new_n13061_), .A2(new_n13060_), .A3(new_n13058_), .A4(new_n8785_), .ZN(new_n13062_));
  INV_X1     g12998(.I(new_n13058_), .ZN(new_n13063_));
  NOR2_X1    g12999(.A1(new_n13061_), .A2(new_n13060_), .ZN(new_n13064_));
  AOI21_X1   g13000(.A1(new_n13064_), .A2(new_n13063_), .B(new_n8784_), .ZN(new_n13065_));
  AOI21_X1   g13001(.A1(new_n10854_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n13066_));
  OAI21_X1   g13002(.A1(new_n2767_), .A2(new_n10861_), .B(new_n13066_), .ZN(new_n13067_));
  AOI21_X1   g13003(.A1(new_n8785_), .A2(new_n3332_), .B(new_n13067_), .ZN(new_n13068_));
  OAI21_X1   g13004(.A1(new_n13065_), .A2(new_n13062_), .B(new_n13068_), .ZN(new_n13069_));
  INV_X1     g13005(.I(new_n4598_), .ZN(new_n13070_));
  NAND4_X1   g13006(.A1(new_n80_), .A2(new_n1192_), .A3(new_n1393_), .A4(new_n1009_), .ZN(new_n13071_));
  NOR3_X1    g13007(.A1(new_n1788_), .A2(new_n333_), .A3(new_n689_), .ZN(new_n13072_));
  NAND4_X1   g13008(.A1(new_n13072_), .A2(new_n765_), .A3(new_n2398_), .A4(new_n13071_), .ZN(new_n13073_));
  INV_X1     g13009(.I(new_n1559_), .ZN(new_n13074_));
  INV_X1     g13010(.I(new_n1996_), .ZN(new_n13075_));
  NAND4_X1   g13011(.A1(new_n13074_), .A2(new_n868_), .A3(new_n13075_), .A4(new_n2942_), .ZN(new_n13076_));
  NOR4_X1    g13012(.A1(new_n13076_), .A2(new_n13070_), .A3(new_n11103_), .A4(new_n13073_), .ZN(new_n13077_));
  NAND3_X1   g13013(.A1(new_n975_), .A2(new_n13077_), .A3(new_n1544_), .ZN(new_n13078_));
  NAND2_X1   g13014(.A1(new_n13069_), .A2(new_n13078_), .ZN(new_n13079_));
  INV_X1     g13015(.I(new_n13079_), .ZN(new_n13080_));
  NOR2_X1    g13016(.A1(new_n13069_), .A2(new_n13078_), .ZN(new_n13081_));
  NOR2_X1    g13017(.A1(new_n13080_), .A2(new_n13081_), .ZN(new_n13082_));
  INV_X1     g13018(.I(new_n13082_), .ZN(new_n13083_));
  NOR2_X1    g13019(.A1(new_n13057_), .A2(new_n13083_), .ZN(new_n13084_));
  INV_X1     g13020(.I(new_n13084_), .ZN(new_n13085_));
  NOR2_X1    g13021(.A1(new_n12819_), .A2(new_n13080_), .ZN(new_n13086_));
  AOI22_X1   g13022(.A1(new_n13085_), .A2(new_n13086_), .B1(new_n12820_), .B2(new_n12808_), .ZN(new_n13087_));
  INV_X1     g13023(.I(new_n13087_), .ZN(new_n13088_));
  AOI22_X1   g13024(.A1(new_n10886_), .A2(new_n2746_), .B1(new_n10889_), .B2(new_n3275_), .ZN(new_n13089_));
  NOR2_X1    g13025(.A1(new_n10899_), .A2(new_n3175_), .ZN(new_n13090_));
  OAI21_X1   g13026(.A1(new_n13090_), .A2(new_n13089_), .B(new_n2736_), .ZN(new_n13091_));
  NOR2_X1    g13027(.A1(new_n11908_), .A2(new_n13091_), .ZN(new_n13092_));
  XOR2_X1    g13028(.A1(new_n13092_), .A2(new_n74_), .Z(new_n13093_));
  INV_X1     g13029(.I(new_n13093_), .ZN(new_n13094_));
  NOR2_X1    g13030(.A1(new_n13094_), .A2(new_n13088_), .ZN(new_n13095_));
  INV_X1     g13031(.I(new_n13095_), .ZN(new_n13096_));
  OAI21_X1   g13032(.A1(new_n12792_), .A2(new_n12794_), .B(new_n13096_), .ZN(new_n13097_));
  NOR2_X1    g13033(.A1(new_n13093_), .A2(new_n13087_), .ZN(new_n13098_));
  INV_X1     g13034(.I(new_n13098_), .ZN(new_n13099_));
  INV_X1     g13035(.I(new_n12771_), .ZN(new_n13100_));
  NAND2_X1   g13036(.A1(new_n10909_), .A2(new_n13100_), .ZN(new_n13101_));
  XOR2_X1    g13037(.A1(new_n10885_), .A2(new_n10871_), .Z(new_n13102_));
  OAI21_X1   g13038(.A1(new_n10909_), .A2(new_n13102_), .B(new_n13101_), .ZN(new_n13103_));
  INV_X1     g13039(.I(new_n13103_), .ZN(new_n13104_));
  NAND2_X1   g13040(.A1(new_n10886_), .A2(new_n3332_), .ZN(new_n13105_));
  NAND2_X1   g13041(.A1(new_n10872_), .A2(new_n3189_), .ZN(new_n13106_));
  NAND2_X1   g13042(.A1(new_n8779_), .A2(new_n2770_), .ZN(new_n13107_));
  NAND4_X1   g13043(.A1(new_n13105_), .A2(new_n2764_), .A3(new_n13106_), .A4(new_n13107_), .ZN(new_n13108_));
  NOR2_X1    g13044(.A1(new_n13104_), .A2(new_n13108_), .ZN(new_n13109_));
  INV_X1     g13045(.I(new_n13109_), .ZN(new_n13110_));
  NAND3_X1   g13046(.A1(new_n13097_), .A2(new_n13099_), .A3(new_n13110_), .ZN(new_n13111_));
  AOI21_X1   g13047(.A1(new_n13097_), .A2(new_n13099_), .B(new_n13110_), .ZN(new_n13112_));
  AOI21_X1   g13048(.A1(new_n12791_), .A2(new_n13111_), .B(new_n13112_), .ZN(new_n13113_));
  AOI21_X1   g13049(.A1(new_n13113_), .A2(new_n12784_), .B(new_n12783_), .ZN(new_n13114_));
  AOI22_X1   g13050(.A1(new_n2746_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n3275_), .ZN(new_n13115_));
  NOR2_X1    g13051(.A1(new_n8758_), .A2(new_n3175_), .ZN(new_n13116_));
  OAI21_X1   g13052(.A1(new_n13115_), .A2(new_n13116_), .B(new_n2736_), .ZN(new_n13117_));
  NOR2_X1    g13053(.A1(new_n12053_), .A2(new_n13117_), .ZN(new_n13118_));
  XOR2_X1    g13054(.A1(new_n13118_), .A2(new_n74_), .Z(new_n13119_));
  INV_X1     g13055(.I(new_n13119_), .ZN(new_n13120_));
  NOR2_X1    g13056(.A1(new_n13114_), .A2(new_n13120_), .ZN(new_n13121_));
  OAI22_X1   g13057(.A1(new_n11851_), .A2(new_n11853_), .B1(new_n12415_), .B2(new_n11865_), .ZN(new_n13122_));
  OAI21_X1   g13058(.A1(new_n11785_), .A2(new_n11784_), .B(new_n11864_), .ZN(new_n13123_));
  NAND3_X1   g13059(.A1(new_n11781_), .A2(new_n11780_), .A3(new_n11862_), .ZN(new_n13124_));
  NAND2_X1   g13060(.A1(new_n13123_), .A2(new_n13124_), .ZN(new_n13125_));
  NAND3_X1   g13061(.A1(new_n12413_), .A2(new_n13125_), .A3(new_n12414_), .ZN(new_n13126_));
  INV_X1     g13062(.I(new_n12782_), .ZN(new_n13127_));
  NAND3_X1   g13063(.A1(new_n13122_), .A2(new_n13126_), .A3(new_n13127_), .ZN(new_n13128_));
  AOI21_X1   g13064(.A1(new_n13122_), .A2(new_n13126_), .B(new_n13127_), .ZN(new_n13129_));
  AOI22_X1   g13065(.A1(new_n12412_), .A2(new_n12414_), .B1(new_n11827_), .B2(new_n11829_), .ZN(new_n13130_));
  NAND2_X1   g13066(.A1(new_n11827_), .A2(new_n11829_), .ZN(new_n13131_));
  AOI21_X1   g13067(.A1(new_n11781_), .A2(new_n11780_), .B(new_n11849_), .ZN(new_n13132_));
  NOR3_X1    g13068(.A1(new_n11785_), .A2(new_n11784_), .A3(new_n11852_), .ZN(new_n13133_));
  NOR2_X1    g13069(.A1(new_n13132_), .A2(new_n13133_), .ZN(new_n13134_));
  NOR2_X1    g13070(.A1(new_n13134_), .A2(new_n13131_), .ZN(new_n13135_));
  NOR2_X1    g13071(.A1(new_n13135_), .A2(new_n13130_), .ZN(new_n13136_));
  OAI22_X1   g13072(.A1(new_n11785_), .A2(new_n11784_), .B1(new_n12410_), .B2(new_n11828_), .ZN(new_n13137_));
  INV_X1     g13073(.I(new_n12793_), .ZN(new_n13138_));
  NAND3_X1   g13074(.A1(new_n11781_), .A2(new_n11780_), .A3(new_n13138_), .ZN(new_n13139_));
  AOI21_X1   g13075(.A1(new_n13137_), .A2(new_n13139_), .B(new_n13095_), .ZN(new_n13140_));
  NOR3_X1    g13076(.A1(new_n13140_), .A2(new_n13098_), .A3(new_n13109_), .ZN(new_n13141_));
  OAI21_X1   g13077(.A1(new_n13140_), .A2(new_n13098_), .B(new_n13109_), .ZN(new_n13142_));
  OAI21_X1   g13078(.A1(new_n13136_), .A2(new_n13141_), .B(new_n13142_), .ZN(new_n13143_));
  OAI21_X1   g13079(.A1(new_n13143_), .A2(new_n13129_), .B(new_n13128_), .ZN(new_n13144_));
  NOR2_X1    g13080(.A1(new_n13144_), .A2(new_n13119_), .ZN(new_n13145_));
  OAI21_X1   g13081(.A1(new_n13145_), .A2(new_n13121_), .B(new_n12762_), .ZN(new_n13146_));
  NAND2_X1   g13082(.A1(new_n12758_), .A2(new_n12759_), .ZN(new_n13147_));
  MUX2_X1    g13083(.I0(new_n12761_), .I1(new_n13147_), .S(new_n11867_), .Z(new_n13148_));
  NAND2_X1   g13084(.A1(new_n13144_), .A2(new_n13119_), .ZN(new_n13149_));
  NAND2_X1   g13085(.A1(new_n13114_), .A2(new_n13120_), .ZN(new_n13150_));
  NAND3_X1   g13086(.A1(new_n13148_), .A2(new_n13149_), .A3(new_n13150_), .ZN(new_n13151_));
  NAND2_X1   g13087(.A1(new_n13151_), .A2(new_n13146_), .ZN(new_n13152_));
  OAI22_X1   g13088(.A1(new_n8745_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8758_), .ZN(new_n13153_));
  NAND2_X1   g13089(.A1(new_n8752_), .A2(new_n3317_), .ZN(new_n13154_));
  AOI21_X1   g13090(.A1(new_n13154_), .A2(new_n13153_), .B(new_n3260_), .ZN(new_n13155_));
  NAND2_X1   g13091(.A1(new_n12189_), .A2(new_n13155_), .ZN(new_n13156_));
  XOR2_X1    g13092(.A1(new_n13156_), .A2(\a[26] ), .Z(new_n13157_));
  OAI22_X1   g13093(.A1(new_n8774_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n10899_), .ZN(new_n13158_));
  NAND2_X1   g13094(.A1(new_n11996_), .A2(new_n2750_), .ZN(new_n13159_));
  AOI21_X1   g13095(.A1(new_n13159_), .A2(new_n13158_), .B(new_n2737_), .ZN(new_n13160_));
  NAND2_X1   g13096(.A1(new_n12001_), .A2(new_n13160_), .ZN(new_n13161_));
  XOR2_X1    g13097(.A1(new_n13161_), .A2(\a[29] ), .Z(new_n13162_));
  NOR2_X1    g13098(.A1(new_n13157_), .A2(new_n13162_), .ZN(new_n13163_));
  INV_X1     g13099(.I(new_n13163_), .ZN(new_n13164_));
  NAND3_X1   g13100(.A1(new_n13143_), .A2(new_n13128_), .A3(new_n12784_), .ZN(new_n13165_));
  OAI21_X1   g13101(.A1(new_n12783_), .A2(new_n13129_), .B(new_n13113_), .ZN(new_n13166_));
  NAND2_X1   g13102(.A1(new_n13157_), .A2(new_n13162_), .ZN(new_n13167_));
  NAND3_X1   g13103(.A1(new_n13166_), .A2(new_n13165_), .A3(new_n13167_), .ZN(new_n13168_));
  OAI22_X1   g13104(.A1(new_n8751_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8745_), .ZN(new_n13169_));
  NAND2_X1   g13105(.A1(new_n10927_), .A2(new_n3317_), .ZN(new_n13170_));
  AOI21_X1   g13106(.A1(new_n13169_), .A2(new_n13170_), .B(new_n3260_), .ZN(new_n13171_));
  NAND2_X1   g13107(.A1(new_n12072_), .A2(new_n13171_), .ZN(new_n13172_));
  XOR2_X1    g13108(.A1(new_n13172_), .A2(\a[26] ), .Z(new_n13173_));
  NAND3_X1   g13109(.A1(new_n13168_), .A2(new_n13164_), .A3(new_n13173_), .ZN(new_n13174_));
  AOI21_X1   g13110(.A1(new_n13168_), .A2(new_n13164_), .B(new_n13173_), .ZN(new_n13175_));
  AOI21_X1   g13111(.A1(new_n13152_), .A2(new_n13174_), .B(new_n13175_), .ZN(new_n13176_));
  OAI22_X1   g13112(.A1(new_n8725_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n8718_), .ZN(new_n13177_));
  NAND2_X1   g13113(.A1(new_n8711_), .A2(new_n3312_), .ZN(new_n13178_));
  AOI21_X1   g13114(.A1(new_n13178_), .A2(new_n13177_), .B(new_n3302_), .ZN(new_n13179_));
  NAND2_X1   g13115(.A1(new_n11536_), .A2(new_n13179_), .ZN(new_n13180_));
  XOR2_X1    g13116(.A1(new_n13180_), .A2(\a[23] ), .Z(new_n13181_));
  AOI21_X1   g13117(.A1(new_n13176_), .A2(new_n13181_), .B(new_n12757_), .ZN(new_n13182_));
  AOI21_X1   g13118(.A1(new_n13149_), .A2(new_n13150_), .B(new_n13148_), .ZN(new_n13183_));
  NOR3_X1    g13119(.A1(new_n13145_), .A2(new_n13121_), .A3(new_n12762_), .ZN(new_n13184_));
  OAI21_X1   g13120(.A1(new_n13183_), .A2(new_n13184_), .B(new_n13174_), .ZN(new_n13185_));
  NOR3_X1    g13121(.A1(new_n13113_), .A2(new_n13129_), .A3(new_n12783_), .ZN(new_n13186_));
  AOI21_X1   g13122(.A1(new_n13128_), .A2(new_n12784_), .B(new_n13143_), .ZN(new_n13187_));
  INV_X1     g13123(.I(new_n13167_), .ZN(new_n13188_));
  NOR3_X1    g13124(.A1(new_n13187_), .A2(new_n13186_), .A3(new_n13188_), .ZN(new_n13189_));
  INV_X1     g13125(.I(new_n13173_), .ZN(new_n13190_));
  OAI21_X1   g13126(.A1(new_n13189_), .A2(new_n13163_), .B(new_n13190_), .ZN(new_n13191_));
  AOI21_X1   g13127(.A1(new_n13185_), .A2(new_n13191_), .B(new_n13181_), .ZN(new_n13192_));
  OAI22_X1   g13128(.A1(new_n8681_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n8694_), .ZN(new_n13193_));
  NAND2_X1   g13129(.A1(new_n8688_), .A2(new_n4096_), .ZN(new_n13194_));
  AOI21_X1   g13130(.A1(new_n13194_), .A2(new_n13193_), .B(new_n4095_), .ZN(new_n13195_));
  NAND2_X1   g13131(.A1(new_n11420_), .A2(new_n13195_), .ZN(new_n13196_));
  XOR2_X1    g13132(.A1(new_n13196_), .A2(\a[20] ), .Z(new_n13197_));
  INV_X1     g13133(.I(new_n13197_), .ZN(new_n13198_));
  NOR3_X1    g13134(.A1(new_n13182_), .A2(new_n13192_), .A3(new_n13198_), .ZN(new_n13199_));
  OAI21_X1   g13135(.A1(new_n13182_), .A2(new_n13192_), .B(new_n13198_), .ZN(new_n13200_));
  OAI21_X1   g13136(.A1(new_n12756_), .A2(new_n13199_), .B(new_n13200_), .ZN(new_n13201_));
  INV_X1     g13137(.I(new_n13201_), .ZN(new_n13202_));
  OAI22_X1   g13138(.A1(new_n3769_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n3775_), .ZN(new_n13203_));
  NAND2_X1   g13139(.A1(new_n8674_), .A2(new_n4096_), .ZN(new_n13204_));
  AOI21_X1   g13140(.A1(new_n13204_), .A2(new_n13203_), .B(new_n4095_), .ZN(new_n13205_));
  NAND2_X1   g13141(.A1(new_n11431_), .A2(new_n13205_), .ZN(new_n13206_));
  XOR2_X1    g13142(.A1(new_n13206_), .A2(\a[20] ), .Z(new_n13207_));
  NOR2_X1    g13143(.A1(new_n13202_), .A2(new_n13207_), .ZN(new_n13208_));
  INV_X1     g13144(.I(new_n13208_), .ZN(new_n13209_));
  XOR2_X1    g13145(.A1(new_n12437_), .A2(new_n12667_), .Z(new_n13210_));
  NOR2_X1    g13146(.A1(new_n12671_), .A2(new_n13210_), .ZN(new_n13211_));
  XOR2_X1    g13147(.A1(new_n12437_), .A2(new_n12673_), .Z(new_n13212_));
  NOR2_X1    g13148(.A1(new_n12669_), .A2(new_n13212_), .ZN(new_n13213_));
  NOR2_X1    g13149(.A1(new_n13211_), .A2(new_n13213_), .ZN(new_n13214_));
  XOR2_X1    g13150(.A1(new_n13214_), .A2(new_n12662_), .Z(new_n13215_));
  NAND3_X1   g13151(.A1(new_n13215_), .A2(new_n13202_), .A3(new_n13207_), .ZN(new_n13216_));
  OAI22_X1   g13152(.A1(new_n11284_), .A2(new_n4291_), .B1(new_n4297_), .B2(new_n11271_), .ZN(new_n13217_));
  NAND2_X1   g13153(.A1(new_n11311_), .A2(new_n4469_), .ZN(new_n13218_));
  AOI21_X1   g13154(.A1(new_n13217_), .A2(new_n13218_), .B(new_n4468_), .ZN(new_n13219_));
  NAND2_X1   g13155(.A1(new_n11391_), .A2(new_n13219_), .ZN(new_n13220_));
  XOR2_X1    g13156(.A1(new_n13220_), .A2(\a[17] ), .Z(new_n13221_));
  NAND3_X1   g13157(.A1(new_n13216_), .A2(new_n13209_), .A3(new_n13221_), .ZN(new_n13222_));
  AOI21_X1   g13158(.A1(new_n13216_), .A2(new_n13209_), .B(new_n13221_), .ZN(new_n13223_));
  AOI21_X1   g13159(.A1(new_n12749_), .A2(new_n13222_), .B(new_n13223_), .ZN(new_n13224_));
  OAI22_X1   g13160(.A1(new_n11353_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n11345_), .ZN(new_n13225_));
  NAND2_X1   g13161(.A1(new_n11370_), .A2(new_n6090_), .ZN(new_n13226_));
  AOI21_X1   g13162(.A1(new_n13226_), .A2(new_n13225_), .B(new_n6082_), .ZN(new_n13227_));
  NAND2_X1   g13163(.A1(new_n11379_), .A2(new_n13227_), .ZN(new_n13228_));
  XOR2_X1    g13164(.A1(new_n13228_), .A2(\a[14] ), .Z(new_n13229_));
  NAND2_X1   g13165(.A1(new_n13224_), .A2(new_n13229_), .ZN(new_n13230_));
  NOR2_X1    g13166(.A1(new_n13224_), .A2(new_n13229_), .ZN(new_n13231_));
  AOI21_X1   g13167(.A1(new_n12742_), .A2(new_n13230_), .B(new_n13231_), .ZN(new_n13232_));
  INV_X1     g13168(.I(new_n12703_), .ZN(new_n13233_));
  INV_X1     g13169(.I(new_n12698_), .ZN(new_n13234_));
  NAND2_X1   g13170(.A1(new_n12706_), .A2(new_n13234_), .ZN(new_n13235_));
  NOR2_X1    g13171(.A1(new_n12706_), .A2(new_n13234_), .ZN(new_n13236_));
  INV_X1     g13172(.I(new_n13236_), .ZN(new_n13237_));
  AOI21_X1   g13173(.A1(new_n13237_), .A2(new_n13235_), .B(new_n13233_), .ZN(new_n13238_));
  INV_X1     g13174(.I(new_n13235_), .ZN(new_n13239_));
  NOR3_X1    g13175(.A1(new_n13239_), .A2(new_n13236_), .A3(new_n12703_), .ZN(new_n13240_));
  OAI21_X1   g13176(.A1(new_n13238_), .A2(new_n13240_), .B(new_n12471_), .ZN(new_n13241_));
  OAI21_X1   g13177(.A1(new_n13239_), .A2(new_n13236_), .B(new_n12703_), .ZN(new_n13242_));
  NAND3_X1   g13178(.A1(new_n13237_), .A2(new_n13233_), .A3(new_n13235_), .ZN(new_n13243_));
  NAND3_X1   g13179(.A1(new_n13242_), .A2(new_n13243_), .A3(new_n12705_), .ZN(new_n13244_));
  OAI22_X1   g13180(.A1(new_n11353_), .A2(new_n6089_), .B1(new_n6091_), .B2(new_n11697_), .ZN(new_n13245_));
  NAND2_X1   g13181(.A1(new_n11370_), .A2(new_n6095_), .ZN(new_n13246_));
  AOI21_X1   g13182(.A1(new_n13246_), .A2(new_n13245_), .B(new_n6082_), .ZN(new_n13247_));
  NAND2_X1   g13183(.A1(new_n11700_), .A2(new_n13247_), .ZN(new_n13248_));
  XOR2_X1    g13184(.A1(new_n13248_), .A2(\a[14] ), .Z(new_n13249_));
  INV_X1     g13185(.I(new_n13249_), .ZN(new_n13250_));
  AOI21_X1   g13186(.A1(new_n13241_), .A2(new_n13244_), .B(new_n13250_), .ZN(new_n13251_));
  NOR2_X1    g13187(.A1(new_n13251_), .A2(new_n13232_), .ZN(new_n13252_));
  NAND3_X1   g13188(.A1(new_n13241_), .A2(new_n13244_), .A3(new_n13250_), .ZN(new_n13253_));
  INV_X1     g13189(.I(new_n13253_), .ZN(new_n13254_));
  NOR3_X1    g13190(.A1(new_n12737_), .A2(new_n13252_), .A3(new_n13254_), .ZN(new_n13255_));
  INV_X1     g13191(.I(new_n13255_), .ZN(new_n13256_));
  INV_X1     g13192(.I(new_n13222_), .ZN(new_n13257_));
  OAI21_X1   g13193(.A1(new_n13257_), .A2(new_n13223_), .B(new_n12749_), .ZN(new_n13258_));
  INV_X1     g13194(.I(new_n12745_), .ZN(new_n13259_));
  AOI21_X1   g13195(.A1(new_n12747_), .A2(new_n12746_), .B(new_n12743_), .ZN(new_n13260_));
  NOR2_X1    g13196(.A1(new_n13259_), .A2(new_n13260_), .ZN(new_n13261_));
  INV_X1     g13197(.I(new_n13221_), .ZN(new_n13262_));
  AOI21_X1   g13198(.A1(new_n13216_), .A2(new_n13209_), .B(new_n13262_), .ZN(new_n13263_));
  NAND3_X1   g13199(.A1(new_n13216_), .A2(new_n13209_), .A3(new_n13262_), .ZN(new_n13264_));
  INV_X1     g13200(.I(new_n13264_), .ZN(new_n13265_));
  OAI21_X1   g13201(.A1(new_n13265_), .A2(new_n13263_), .B(new_n13261_), .ZN(new_n13266_));
  NAND2_X1   g13202(.A1(new_n13266_), .A2(new_n13258_), .ZN(new_n13267_));
  NAND2_X1   g13203(.A1(new_n12654_), .A2(new_n12660_), .ZN(new_n13268_));
  OAI21_X1   g13204(.A1(new_n12632_), .A2(new_n12635_), .B(new_n13268_), .ZN(new_n13269_));
  NAND3_X1   g13205(.A1(new_n12755_), .A2(new_n12751_), .A3(new_n12753_), .ZN(new_n13270_));
  NAND2_X1   g13206(.A1(new_n13270_), .A2(new_n13269_), .ZN(new_n13271_));
  XOR2_X1    g13207(.A1(new_n12658_), .A2(new_n12647_), .Z(new_n13272_));
  NOR2_X1    g13208(.A1(new_n13183_), .A2(new_n13184_), .ZN(new_n13273_));
  NOR3_X1    g13209(.A1(new_n13189_), .A2(new_n13163_), .A3(new_n13190_), .ZN(new_n13274_));
  OAI21_X1   g13210(.A1(new_n13273_), .A2(new_n13274_), .B(new_n13191_), .ZN(new_n13275_));
  INV_X1     g13211(.I(new_n13181_), .ZN(new_n13276_));
  OAI21_X1   g13212(.A1(new_n13275_), .A2(new_n13276_), .B(new_n13272_), .ZN(new_n13277_));
  NAND2_X1   g13213(.A1(new_n13275_), .A2(new_n13276_), .ZN(new_n13278_));
  AOI21_X1   g13214(.A1(new_n13277_), .A2(new_n13278_), .B(new_n13197_), .ZN(new_n13279_));
  OAI21_X1   g13215(.A1(new_n13199_), .A2(new_n13279_), .B(new_n13271_), .ZN(new_n13280_));
  AOI21_X1   g13216(.A1(new_n13277_), .A2(new_n13278_), .B(new_n13198_), .ZN(new_n13281_));
  NOR3_X1    g13217(.A1(new_n13182_), .A2(new_n13192_), .A3(new_n13197_), .ZN(new_n13282_));
  OAI21_X1   g13218(.A1(new_n13281_), .A2(new_n13282_), .B(new_n12756_), .ZN(new_n13283_));
  NAND2_X1   g13219(.A1(new_n13283_), .A2(new_n13280_), .ZN(new_n13284_));
  NAND2_X1   g13220(.A1(new_n13176_), .A2(new_n13181_), .ZN(new_n13285_));
  AOI21_X1   g13221(.A1(new_n13278_), .A2(new_n13285_), .B(new_n12757_), .ZN(new_n13286_));
  NAND2_X1   g13222(.A1(new_n13275_), .A2(new_n13181_), .ZN(new_n13287_));
  NAND3_X1   g13223(.A1(new_n13185_), .A2(new_n13191_), .A3(new_n13276_), .ZN(new_n13288_));
  AOI21_X1   g13224(.A1(new_n13287_), .A2(new_n13288_), .B(new_n13272_), .ZN(new_n13289_));
  XNOR2_X1   g13225(.A1(new_n13157_), .A2(new_n13162_), .ZN(new_n13290_));
  INV_X1     g13226(.I(new_n13290_), .ZN(new_n13291_));
  OAI21_X1   g13227(.A1(new_n13187_), .A2(new_n13186_), .B(new_n13291_), .ZN(new_n13292_));
  NOR2_X1    g13228(.A1(new_n13188_), .A2(new_n13163_), .ZN(new_n13293_));
  INV_X1     g13229(.I(new_n13293_), .ZN(new_n13294_));
  NAND3_X1   g13230(.A1(new_n13166_), .A2(new_n13165_), .A3(new_n13294_), .ZN(new_n13295_));
  OAI22_X1   g13231(.A1(new_n8758_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8766_), .ZN(new_n13296_));
  NAND2_X1   g13232(.A1(new_n8746_), .A2(new_n3317_), .ZN(new_n13297_));
  AOI21_X1   g13233(.A1(new_n13297_), .A2(new_n13296_), .B(new_n3260_), .ZN(new_n13298_));
  NAND2_X1   g13234(.A1(new_n11964_), .A2(new_n13298_), .ZN(new_n13299_));
  XOR2_X1    g13235(.A1(new_n13299_), .A2(\a[26] ), .Z(new_n13300_));
  AOI22_X1   g13236(.A1(new_n11899_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n10889_), .ZN(new_n13301_));
  NOR2_X1    g13237(.A1(new_n8774_), .A2(new_n3175_), .ZN(new_n13302_));
  OAI21_X1   g13238(.A1(new_n13302_), .A2(new_n13301_), .B(new_n2736_), .ZN(new_n13303_));
  NOR2_X1    g13239(.A1(new_n11945_), .A2(new_n13303_), .ZN(new_n13304_));
  XOR2_X1    g13240(.A1(new_n13304_), .A2(new_n74_), .Z(new_n13305_));
  NOR2_X1    g13241(.A1(new_n13300_), .A2(new_n13305_), .ZN(new_n13306_));
  NAND2_X1   g13242(.A1(new_n13097_), .A2(new_n13099_), .ZN(new_n13307_));
  NAND3_X1   g13243(.A1(new_n12790_), .A2(new_n12785_), .A3(new_n13110_), .ZN(new_n13308_));
  OAI21_X1   g13244(.A1(new_n13135_), .A2(new_n13130_), .B(new_n13109_), .ZN(new_n13309_));
  NAND3_X1   g13245(.A1(new_n13309_), .A2(new_n13308_), .A3(new_n13307_), .ZN(new_n13310_));
  INV_X1     g13246(.I(new_n13307_), .ZN(new_n13311_));
  NOR3_X1    g13247(.A1(new_n13135_), .A2(new_n13130_), .A3(new_n13109_), .ZN(new_n13312_));
  AOI21_X1   g13248(.A1(new_n12790_), .A2(new_n12785_), .B(new_n13110_), .ZN(new_n13313_));
  OAI21_X1   g13249(.A1(new_n13312_), .A2(new_n13313_), .B(new_n13311_), .ZN(new_n13314_));
  NAND2_X1   g13250(.A1(new_n13314_), .A2(new_n13310_), .ZN(new_n13315_));
  INV_X1     g13251(.I(new_n13300_), .ZN(new_n13316_));
  INV_X1     g13252(.I(new_n13305_), .ZN(new_n13317_));
  NOR2_X1    g13253(.A1(new_n13316_), .A2(new_n13317_), .ZN(new_n13318_));
  AOI21_X1   g13254(.A1(new_n13315_), .A2(new_n13318_), .B(new_n13306_), .ZN(new_n13319_));
  OAI22_X1   g13255(.A1(new_n8735_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n10924_), .ZN(new_n13320_));
  NAND2_X1   g13256(.A1(new_n8726_), .A2(new_n3312_), .ZN(new_n13321_));
  AOI21_X1   g13257(.A1(new_n13321_), .A2(new_n13320_), .B(new_n3302_), .ZN(new_n13322_));
  NAND2_X1   g13258(.A1(new_n12181_), .A2(new_n13322_), .ZN(new_n13323_));
  XOR2_X1    g13259(.A1(new_n13323_), .A2(\a[23] ), .Z(new_n13324_));
  AOI22_X1   g13260(.A1(new_n13292_), .A2(new_n13295_), .B1(new_n13319_), .B2(new_n13324_), .ZN(new_n13325_));
  NOR2_X1    g13261(.A1(new_n13319_), .A2(new_n13324_), .ZN(new_n13326_));
  NOR2_X1    g13262(.A1(new_n13325_), .A2(new_n13326_), .ZN(new_n13327_));
  INV_X1     g13263(.I(new_n13327_), .ZN(new_n13328_));
  OAI22_X1   g13264(.A1(new_n8725_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8735_), .ZN(new_n13329_));
  NAND2_X1   g13265(.A1(new_n8719_), .A2(new_n3312_), .ZN(new_n13330_));
  AOI21_X1   g13266(.A1(new_n13329_), .A2(new_n13330_), .B(new_n3302_), .ZN(new_n13331_));
  NAND2_X1   g13267(.A1(new_n12242_), .A2(new_n13331_), .ZN(new_n13332_));
  XOR2_X1    g13268(.A1(new_n13332_), .A2(\a[23] ), .Z(new_n13333_));
  INV_X1     g13269(.I(new_n13333_), .ZN(new_n13334_));
  NAND2_X1   g13270(.A1(new_n13328_), .A2(new_n13334_), .ZN(new_n13335_));
  AOI21_X1   g13271(.A1(new_n13168_), .A2(new_n13164_), .B(new_n13190_), .ZN(new_n13336_));
  NOR3_X1    g13272(.A1(new_n13189_), .A2(new_n13163_), .A3(new_n13173_), .ZN(new_n13337_));
  OAI22_X1   g13273(.A1(new_n13337_), .A2(new_n13336_), .B1(new_n13183_), .B2(new_n13184_), .ZN(new_n13338_));
  NAND2_X1   g13274(.A1(new_n13191_), .A2(new_n13174_), .ZN(new_n13339_));
  NAND2_X1   g13275(.A1(new_n13339_), .A2(new_n13273_), .ZN(new_n13340_));
  AOI21_X1   g13276(.A1(new_n13166_), .A2(new_n13165_), .B(new_n13290_), .ZN(new_n13341_));
  NOR3_X1    g13277(.A1(new_n13187_), .A2(new_n13186_), .A3(new_n13293_), .ZN(new_n13342_));
  INV_X1     g13278(.I(new_n13306_), .ZN(new_n13343_));
  NOR3_X1    g13279(.A1(new_n13312_), .A2(new_n13313_), .A3(new_n13311_), .ZN(new_n13344_));
  AOI21_X1   g13280(.A1(new_n13309_), .A2(new_n13308_), .B(new_n13307_), .ZN(new_n13345_));
  OAI21_X1   g13281(.A1(new_n13344_), .A2(new_n13345_), .B(new_n13318_), .ZN(new_n13346_));
  NAND2_X1   g13282(.A1(new_n13346_), .A2(new_n13343_), .ZN(new_n13347_));
  INV_X1     g13283(.I(new_n13324_), .ZN(new_n13348_));
  OAI22_X1   g13284(.A1(new_n13341_), .A2(new_n13342_), .B1(new_n13347_), .B2(new_n13348_), .ZN(new_n13349_));
  INV_X1     g13285(.I(new_n13326_), .ZN(new_n13350_));
  NAND3_X1   g13286(.A1(new_n13350_), .A2(new_n13349_), .A3(new_n13333_), .ZN(new_n13351_));
  NAND3_X1   g13287(.A1(new_n13340_), .A2(new_n13351_), .A3(new_n13338_), .ZN(new_n13352_));
  NAND2_X1   g13288(.A1(new_n13335_), .A2(new_n13352_), .ZN(new_n13353_));
  OAI22_X1   g13289(.A1(new_n8701_), .A2(new_n3769_), .B1(new_n8694_), .B2(new_n3775_), .ZN(new_n13354_));
  NAND2_X1   g13290(.A1(new_n8682_), .A2(new_n4096_), .ZN(new_n13355_));
  AOI21_X1   g13291(.A1(new_n13355_), .A2(new_n13354_), .B(new_n4095_), .ZN(new_n13356_));
  NAND2_X1   g13292(.A1(new_n12347_), .A2(new_n13356_), .ZN(new_n13357_));
  XOR2_X1    g13293(.A1(new_n13357_), .A2(\a[20] ), .Z(new_n13358_));
  INV_X1     g13294(.I(new_n13358_), .ZN(new_n13359_));
  OAI22_X1   g13295(.A1(new_n13286_), .A2(new_n13289_), .B1(new_n13353_), .B2(new_n13359_), .ZN(new_n13360_));
  NAND2_X1   g13296(.A1(new_n13353_), .A2(new_n13359_), .ZN(new_n13361_));
  OAI22_X1   g13297(.A1(new_n8661_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8673_), .ZN(new_n13362_));
  NAND2_X1   g13298(.A1(new_n11285_), .A2(new_n4469_), .ZN(new_n13363_));
  AOI21_X1   g13299(.A1(new_n13363_), .A2(new_n13362_), .B(new_n4468_), .ZN(new_n13364_));
  NAND2_X1   g13300(.A1(new_n11323_), .A2(new_n13364_), .ZN(new_n13365_));
  XOR2_X1    g13301(.A1(new_n13365_), .A2(\a[17] ), .Z(new_n13366_));
  NAND3_X1   g13302(.A1(new_n13360_), .A2(new_n13361_), .A3(new_n13366_), .ZN(new_n13367_));
  AOI21_X1   g13303(.A1(new_n13360_), .A2(new_n13361_), .B(new_n13366_), .ZN(new_n13368_));
  AOI21_X1   g13304(.A1(new_n13284_), .A2(new_n13367_), .B(new_n13368_), .ZN(new_n13369_));
  OAI22_X1   g13305(.A1(new_n11284_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8661_), .ZN(new_n13370_));
  NAND2_X1   g13306(.A1(new_n11272_), .A2(new_n4469_), .ZN(new_n13371_));
  AOI21_X1   g13307(.A1(new_n13370_), .A2(new_n13371_), .B(new_n4468_), .ZN(new_n13372_));
  NAND2_X1   g13308(.A1(new_n11655_), .A2(new_n13372_), .ZN(new_n13373_));
  XOR2_X1    g13309(.A1(new_n13373_), .A2(\a[17] ), .Z(new_n13374_));
  NOR2_X1    g13310(.A1(new_n13369_), .A2(new_n13374_), .ZN(new_n13375_));
  INV_X1     g13311(.I(new_n13374_), .ZN(new_n13376_));
  INV_X1     g13312(.I(new_n13207_), .ZN(new_n13377_));
  XOR2_X1    g13313(.A1(new_n12661_), .A2(new_n13377_), .Z(new_n13378_));
  XOR2_X1    g13314(.A1(new_n12661_), .A2(new_n13207_), .Z(new_n13379_));
  OR3_X2     g13315(.A1(new_n13211_), .A2(new_n13213_), .A3(new_n13379_), .Z(new_n13380_));
  OAI21_X1   g13316(.A1(new_n13214_), .A2(new_n13378_), .B(new_n13380_), .ZN(new_n13381_));
  XOR2_X1    g13317(.A1(new_n13381_), .A2(new_n13202_), .Z(new_n13382_));
  NOR2_X1    g13318(.A1(new_n13382_), .A2(new_n13376_), .ZN(new_n13383_));
  AOI21_X1   g13319(.A1(new_n13383_), .A2(new_n13369_), .B(new_n13375_), .ZN(new_n13384_));
  OAI22_X1   g13320(.A1(new_n11264_), .A2(new_n6089_), .B1(new_n6094_), .B2(new_n11345_), .ZN(new_n13385_));
  NAND2_X1   g13321(.A1(new_n11354_), .A2(new_n6090_), .ZN(new_n13386_));
  AOI21_X1   g13322(.A1(new_n13386_), .A2(new_n13385_), .B(new_n6082_), .ZN(new_n13387_));
  NAND2_X1   g13323(.A1(new_n11678_), .A2(new_n13387_), .ZN(new_n13388_));
  XOR2_X1    g13324(.A1(new_n13388_), .A2(\a[14] ), .Z(new_n13389_));
  NAND2_X1   g13325(.A1(new_n13384_), .A2(new_n13389_), .ZN(new_n13390_));
  NAND2_X1   g13326(.A1(new_n13267_), .A2(new_n13390_), .ZN(new_n13391_));
  INV_X1     g13327(.I(new_n13375_), .ZN(new_n13392_));
  XOR2_X1    g13328(.A1(new_n13381_), .A2(new_n13201_), .Z(new_n13393_));
  NAND3_X1   g13329(.A1(new_n13393_), .A2(new_n13369_), .A3(new_n13374_), .ZN(new_n13394_));
  NAND2_X1   g13330(.A1(new_n13394_), .A2(new_n13392_), .ZN(new_n13395_));
  INV_X1     g13331(.I(new_n13389_), .ZN(new_n13396_));
  NAND2_X1   g13332(.A1(new_n13395_), .A2(new_n13396_), .ZN(new_n13397_));
  NAND2_X1   g13333(.A1(new_n13391_), .A2(new_n13397_), .ZN(new_n13398_));
  INV_X1     g13334(.I(new_n13398_), .ZN(new_n13399_));
  NOR2_X1    g13335(.A1(new_n12739_), .A2(new_n12741_), .ZN(new_n13400_));
  INV_X1     g13336(.I(new_n13231_), .ZN(new_n13401_));
  AOI21_X1   g13337(.A1(new_n13230_), .A2(new_n13401_), .B(new_n13400_), .ZN(new_n13402_));
  INV_X1     g13338(.I(new_n13229_), .ZN(new_n13403_));
  NOR2_X1    g13339(.A1(new_n13224_), .A2(new_n13403_), .ZN(new_n13404_));
  INV_X1     g13340(.I(new_n13404_), .ZN(new_n13405_));
  NAND2_X1   g13341(.A1(new_n13224_), .A2(new_n13403_), .ZN(new_n13406_));
  NAND2_X1   g13342(.A1(new_n13405_), .A2(new_n13406_), .ZN(new_n13407_));
  AOI21_X1   g13343(.A1(new_n13400_), .A2(new_n13407_), .B(new_n13402_), .ZN(new_n13408_));
  AND3_X2    g13344(.A1(new_n11463_), .A2(new_n6480_), .A3(new_n12255_), .Z(new_n13409_));
  NOR4_X1    g13345(.A1(new_n11468_), .A2(new_n4707_), .A3(new_n11461_), .A4(new_n13409_), .ZN(new_n13410_));
  XOR2_X1    g13346(.A1(new_n13410_), .A2(new_n4034_), .Z(new_n13411_));
  NAND2_X1   g13347(.A1(new_n13408_), .A2(new_n13411_), .ZN(new_n13412_));
  NAND2_X1   g13348(.A1(new_n13401_), .A2(new_n13230_), .ZN(new_n13413_));
  NAND2_X1   g13349(.A1(new_n12742_), .A2(new_n13413_), .ZN(new_n13414_));
  NAND2_X1   g13350(.A1(new_n13407_), .A2(new_n13400_), .ZN(new_n13415_));
  NAND2_X1   g13351(.A1(new_n13414_), .A2(new_n13415_), .ZN(new_n13416_));
  INV_X1     g13352(.I(new_n13411_), .ZN(new_n13417_));
  NAND2_X1   g13353(.A1(new_n13416_), .A2(new_n13417_), .ZN(new_n13418_));
  AOI21_X1   g13354(.A1(new_n13412_), .A2(new_n13418_), .B(new_n13399_), .ZN(new_n13419_));
  NAND2_X1   g13355(.A1(new_n13416_), .A2(new_n13411_), .ZN(new_n13420_));
  NAND2_X1   g13356(.A1(new_n13408_), .A2(new_n13417_), .ZN(new_n13421_));
  AOI21_X1   g13357(.A1(new_n13421_), .A2(new_n13420_), .B(new_n13398_), .ZN(new_n13422_));
  NOR2_X1    g13358(.A1(new_n13395_), .A2(new_n13396_), .ZN(new_n13423_));
  NOR2_X1    g13359(.A1(new_n13384_), .A2(new_n13389_), .ZN(new_n13424_));
  OAI21_X1   g13360(.A1(new_n13423_), .A2(new_n13424_), .B(new_n13267_), .ZN(new_n13425_));
  INV_X1     g13361(.I(new_n13223_), .ZN(new_n13426_));
  AOI21_X1   g13362(.A1(new_n13426_), .A2(new_n13222_), .B(new_n13261_), .ZN(new_n13427_));
  INV_X1     g13363(.I(new_n13263_), .ZN(new_n13428_));
  AOI21_X1   g13364(.A1(new_n13428_), .A2(new_n13264_), .B(new_n12749_), .ZN(new_n13429_));
  NOR2_X1    g13365(.A1(new_n13427_), .A2(new_n13429_), .ZN(new_n13430_));
  NOR2_X1    g13366(.A1(new_n13384_), .A2(new_n13396_), .ZN(new_n13431_));
  NOR2_X1    g13367(.A1(new_n13395_), .A2(new_n13389_), .ZN(new_n13432_));
  OAI21_X1   g13368(.A1(new_n13431_), .A2(new_n13432_), .B(new_n13430_), .ZN(new_n13433_));
  NAND2_X1   g13369(.A1(new_n13433_), .A2(new_n13425_), .ZN(new_n13434_));
  NOR2_X1    g13370(.A1(new_n13275_), .A2(new_n13276_), .ZN(new_n13435_));
  OAI21_X1   g13371(.A1(new_n13435_), .A2(new_n13192_), .B(new_n13272_), .ZN(new_n13436_));
  AOI21_X1   g13372(.A1(new_n13185_), .A2(new_n13191_), .B(new_n13276_), .ZN(new_n13437_));
  AOI21_X1   g13373(.A1(new_n13146_), .A2(new_n13151_), .B(new_n13274_), .ZN(new_n13438_));
  NOR3_X1    g13374(.A1(new_n13438_), .A2(new_n13175_), .A3(new_n13181_), .ZN(new_n13439_));
  OAI21_X1   g13375(.A1(new_n13439_), .A2(new_n13437_), .B(new_n12757_), .ZN(new_n13440_));
  NOR2_X1    g13376(.A1(new_n13327_), .A2(new_n13333_), .ZN(new_n13441_));
  OAI21_X1   g13377(.A1(new_n13189_), .A2(new_n13163_), .B(new_n13173_), .ZN(new_n13442_));
  NAND3_X1   g13378(.A1(new_n13168_), .A2(new_n13164_), .A3(new_n13190_), .ZN(new_n13443_));
  AOI22_X1   g13379(.A1(new_n13442_), .A2(new_n13443_), .B1(new_n13151_), .B2(new_n13146_), .ZN(new_n13444_));
  NOR2_X1    g13380(.A1(new_n13274_), .A2(new_n13175_), .ZN(new_n13445_));
  NOR2_X1    g13381(.A1(new_n13445_), .A2(new_n13152_), .ZN(new_n13446_));
  NOR3_X1    g13382(.A1(new_n13325_), .A2(new_n13326_), .A3(new_n13334_), .ZN(new_n13447_));
  NOR3_X1    g13383(.A1(new_n13446_), .A2(new_n13444_), .A3(new_n13447_), .ZN(new_n13448_));
  NOR2_X1    g13384(.A1(new_n13448_), .A2(new_n13441_), .ZN(new_n13449_));
  AOI22_X1   g13385(.A1(new_n13449_), .A2(new_n13358_), .B1(new_n13436_), .B2(new_n13440_), .ZN(new_n13450_));
  NOR2_X1    g13386(.A1(new_n13449_), .A2(new_n13358_), .ZN(new_n13451_));
  INV_X1     g13387(.I(new_n13366_), .ZN(new_n13452_));
  NOR3_X1    g13388(.A1(new_n13450_), .A2(new_n13451_), .A3(new_n13452_), .ZN(new_n13453_));
  OAI21_X1   g13389(.A1(new_n13368_), .A2(new_n13453_), .B(new_n13284_), .ZN(new_n13454_));
  NAND3_X1   g13390(.A1(new_n13277_), .A2(new_n13278_), .A3(new_n13197_), .ZN(new_n13455_));
  AOI21_X1   g13391(.A1(new_n13455_), .A2(new_n13200_), .B(new_n12756_), .ZN(new_n13456_));
  OAI21_X1   g13392(.A1(new_n13182_), .A2(new_n13192_), .B(new_n13197_), .ZN(new_n13457_));
  NAND3_X1   g13393(.A1(new_n13277_), .A2(new_n13278_), .A3(new_n13198_), .ZN(new_n13458_));
  AOI21_X1   g13394(.A1(new_n13457_), .A2(new_n13458_), .B(new_n13271_), .ZN(new_n13459_));
  NOR2_X1    g13395(.A1(new_n13456_), .A2(new_n13459_), .ZN(new_n13460_));
  AOI21_X1   g13396(.A1(new_n13360_), .A2(new_n13361_), .B(new_n13452_), .ZN(new_n13461_));
  NOR3_X1    g13397(.A1(new_n13450_), .A2(new_n13451_), .A3(new_n13366_), .ZN(new_n13462_));
  OAI21_X1   g13398(.A1(new_n13461_), .A2(new_n13462_), .B(new_n13460_), .ZN(new_n13463_));
  NAND2_X1   g13399(.A1(new_n13463_), .A2(new_n13454_), .ZN(new_n13464_));
  NAND2_X1   g13400(.A1(new_n13436_), .A2(new_n13440_), .ZN(new_n13465_));
  NOR2_X1    g13401(.A1(new_n13353_), .A2(new_n13359_), .ZN(new_n13466_));
  OAI21_X1   g13402(.A1(new_n13466_), .A2(new_n13451_), .B(new_n13465_), .ZN(new_n13467_));
  NOR2_X1    g13403(.A1(new_n13286_), .A2(new_n13289_), .ZN(new_n13468_));
  OAI21_X1   g13404(.A1(new_n13448_), .A2(new_n13441_), .B(new_n13358_), .ZN(new_n13469_));
  NAND3_X1   g13405(.A1(new_n13335_), .A2(new_n13352_), .A3(new_n13359_), .ZN(new_n13470_));
  NAND2_X1   g13406(.A1(new_n13469_), .A2(new_n13470_), .ZN(new_n13471_));
  NAND2_X1   g13407(.A1(new_n13471_), .A2(new_n13468_), .ZN(new_n13472_));
  AOI21_X1   g13408(.A1(new_n13314_), .A2(new_n13310_), .B(new_n13317_), .ZN(new_n13473_));
  NOR3_X1    g13409(.A1(new_n13344_), .A2(new_n13345_), .A3(new_n13305_), .ZN(new_n13474_));
  OAI21_X1   g13410(.A1(new_n13474_), .A2(new_n13473_), .B(new_n13300_), .ZN(new_n13475_));
  OAI21_X1   g13411(.A1(new_n13344_), .A2(new_n13345_), .B(new_n13305_), .ZN(new_n13476_));
  NAND3_X1   g13412(.A1(new_n13314_), .A2(new_n13310_), .A3(new_n13317_), .ZN(new_n13477_));
  NAND3_X1   g13413(.A1(new_n13476_), .A2(new_n13477_), .A3(new_n13316_), .ZN(new_n13478_));
  NAND2_X1   g13414(.A1(new_n13475_), .A2(new_n13478_), .ZN(new_n13479_));
  XNOR2_X1   g13415(.A1(new_n12950_), .A2(new_n12964_), .ZN(new_n13480_));
  XNOR2_X1   g13416(.A1(new_n12950_), .A2(new_n12964_), .ZN(new_n13481_));
  NOR2_X1    g13417(.A1(new_n13481_), .A2(new_n12935_), .ZN(new_n13482_));
  AOI21_X1   g13418(.A1(new_n12935_), .A2(new_n13480_), .B(new_n13482_), .ZN(new_n13483_));
  NOR2_X1    g13419(.A1(new_n13040_), .A2(new_n13036_), .ZN(new_n13484_));
  OAI22_X1   g13420(.A1(new_n9478_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n10853_), .ZN(new_n13485_));
  NAND2_X1   g13421(.A1(new_n10862_), .A2(new_n2750_), .ZN(new_n13486_));
  AOI21_X1   g13422(.A1(new_n13485_), .A2(new_n13486_), .B(new_n2737_), .ZN(new_n13487_));
  NAND2_X1   g13423(.A1(new_n13484_), .A2(new_n13487_), .ZN(new_n13488_));
  XOR2_X1    g13424(.A1(new_n13488_), .A2(\a[29] ), .Z(new_n13489_));
  XOR2_X1    g13425(.A1(new_n13489_), .A2(new_n13483_), .Z(new_n13490_));
  OAI22_X1   g13426(.A1(new_n9478_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n10846_), .ZN(new_n13491_));
  NAND2_X1   g13427(.A1(new_n10854_), .A2(new_n2750_), .ZN(new_n13492_));
  AOI21_X1   g13428(.A1(new_n13491_), .A2(new_n13492_), .B(new_n2737_), .ZN(new_n13493_));
  NAND2_X1   g13429(.A1(new_n13016_), .A2(new_n13493_), .ZN(new_n13494_));
  XOR2_X1    g13430(.A1(new_n13494_), .A2(new_n74_), .Z(new_n13495_));
  NAND2_X1   g13431(.A1(new_n12934_), .A2(new_n12932_), .ZN(new_n13496_));
  NAND2_X1   g13432(.A1(new_n13496_), .A2(new_n12899_), .ZN(new_n13497_));
  XNOR2_X1   g13433(.A1(new_n12914_), .A2(new_n12931_), .ZN(new_n13498_));
  OAI21_X1   g13434(.A1(new_n12899_), .A2(new_n13498_), .B(new_n13497_), .ZN(new_n13499_));
  NOR2_X1    g13435(.A1(new_n13495_), .A2(new_n13499_), .ZN(new_n13500_));
  NOR2_X1    g13436(.A1(new_n12826_), .A2(new_n5021_), .ZN(new_n13501_));
  INV_X1     g13437(.I(new_n12877_), .ZN(new_n13502_));
  AOI21_X1   g13438(.A1(new_n12876_), .A2(new_n12873_), .B(new_n10798_), .ZN(new_n13503_));
  NOR2_X1    g13439(.A1(new_n13502_), .A2(new_n13503_), .ZN(new_n13504_));
  AOI22_X1   g13440(.A1(new_n12823_), .A2(new_n2746_), .B1(new_n3275_), .B2(new_n10800_), .ZN(new_n13505_));
  AOI21_X1   g13441(.A1(new_n2750_), .A2(new_n9529_), .B(new_n13505_), .ZN(new_n13506_));
  NOR3_X1    g13442(.A1(new_n13504_), .A2(new_n2737_), .A3(new_n13506_), .ZN(new_n13507_));
  NAND2_X1   g13443(.A1(new_n13507_), .A2(new_n74_), .ZN(new_n13508_));
  NOR2_X1    g13444(.A1(new_n13507_), .A2(new_n74_), .ZN(new_n13509_));
  INV_X1     g13445(.I(new_n13509_), .ZN(new_n13510_));
  AOI21_X1   g13446(.A1(new_n13510_), .A2(new_n13508_), .B(new_n13501_), .ZN(new_n13511_));
  AOI22_X1   g13447(.A1(new_n10794_), .A2(new_n2746_), .B1(new_n3275_), .B2(new_n12823_), .ZN(new_n13512_));
  AOI21_X1   g13448(.A1(new_n2750_), .A2(new_n10800_), .B(new_n13512_), .ZN(new_n13513_));
  NAND2_X1   g13449(.A1(new_n12830_), .A2(new_n2736_), .ZN(new_n13514_));
  OAI21_X1   g13450(.A1(new_n13514_), .A2(new_n13513_), .B(new_n74_), .ZN(new_n13515_));
  INV_X1     g13451(.I(new_n13515_), .ZN(new_n13516_));
  NOR3_X1    g13452(.A1(new_n13514_), .A2(new_n74_), .A3(new_n13513_), .ZN(new_n13517_));
  NOR2_X1    g13453(.A1(new_n2735_), .A2(new_n2734_), .ZN(new_n13518_));
  OAI21_X1   g13454(.A1(new_n12826_), .A2(new_n2742_), .B(new_n13518_), .ZN(new_n13519_));
  NOR2_X1    g13455(.A1(new_n12847_), .A2(new_n13519_), .ZN(new_n13520_));
  NOR2_X1    g13456(.A1(new_n12826_), .A2(new_n2734_), .ZN(new_n13521_));
  INV_X1     g13457(.I(new_n13521_), .ZN(new_n13522_));
  NAND3_X1   g13458(.A1(new_n13520_), .A2(\a[29] ), .A3(new_n13522_), .ZN(new_n13523_));
  NOR3_X1    g13459(.A1(new_n13516_), .A2(new_n13517_), .A3(new_n13523_), .ZN(new_n13524_));
  INV_X1     g13460(.I(new_n13524_), .ZN(new_n13525_));
  NAND3_X1   g13461(.A1(new_n13510_), .A2(new_n13501_), .A3(new_n13508_), .ZN(new_n13526_));
  AOI21_X1   g13462(.A1(new_n13525_), .A2(new_n13526_), .B(new_n13511_), .ZN(new_n13527_));
  INV_X1     g13463(.I(new_n13527_), .ZN(new_n13528_));
  OAI21_X1   g13464(.A1(new_n12907_), .A2(new_n12905_), .B(new_n9529_), .ZN(new_n13529_));
  AOI21_X1   g13465(.A1(new_n13529_), .A2(new_n12940_), .B(new_n10844_), .ZN(new_n13530_));
  INV_X1     g13466(.I(new_n12904_), .ZN(new_n13531_));
  NAND3_X1   g13467(.A1(new_n12901_), .A2(new_n9529_), .A3(new_n10799_), .ZN(new_n13532_));
  AOI21_X1   g13468(.A1(new_n13532_), .A2(new_n13531_), .B(new_n10839_), .ZN(new_n13533_));
  NOR2_X1    g13469(.A1(new_n13530_), .A2(new_n13533_), .ZN(new_n13534_));
  AOI22_X1   g13470(.A1(new_n9529_), .A2(new_n3275_), .B1(new_n10800_), .B2(new_n2746_), .ZN(new_n13535_));
  AOI21_X1   g13471(.A1(new_n10839_), .A2(new_n2750_), .B(new_n13535_), .ZN(new_n13536_));
  OR3_X2     g13472(.A1(new_n13534_), .A2(new_n2737_), .A3(new_n13536_), .Z(new_n13537_));
  XOR2_X1    g13473(.A1(new_n13537_), .A2(\a[29] ), .Z(new_n13538_));
  OR2_X2     g13474(.A1(new_n12848_), .A2(new_n12869_), .Z(new_n13539_));
  NAND2_X1   g13475(.A1(new_n13539_), .A2(new_n12870_), .ZN(new_n13540_));
  INV_X1     g13476(.I(new_n13540_), .ZN(new_n13541_));
  NAND2_X1   g13477(.A1(new_n13538_), .A2(new_n13541_), .ZN(new_n13542_));
  NOR2_X1    g13478(.A1(new_n13538_), .A2(new_n13541_), .ZN(new_n13543_));
  AOI21_X1   g13479(.A1(new_n13528_), .A2(new_n13542_), .B(new_n13543_), .ZN(new_n13544_));
  AOI22_X1   g13480(.A1(new_n10839_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n9529_), .ZN(new_n13545_));
  NOR2_X1    g13481(.A1(new_n10846_), .A2(new_n3175_), .ZN(new_n13546_));
  OAI21_X1   g13482(.A1(new_n13545_), .A2(new_n13546_), .B(new_n2736_), .ZN(new_n13547_));
  NOR2_X1    g13483(.A1(new_n12946_), .A2(new_n13547_), .ZN(new_n13548_));
  XOR2_X1    g13484(.A1(new_n13548_), .A2(\a[29] ), .Z(new_n13549_));
  XNOR2_X1   g13485(.A1(new_n12834_), .A2(new_n12842_), .ZN(new_n13550_));
  NOR2_X1    g13486(.A1(new_n13550_), .A2(new_n12870_), .ZN(new_n13551_));
  INV_X1     g13487(.I(new_n12843_), .ZN(new_n13552_));
  AOI22_X1   g13488(.A1(new_n13552_), .A2(new_n12871_), .B1(new_n12848_), .B2(new_n12869_), .ZN(new_n13553_));
  NOR2_X1    g13489(.A1(new_n13551_), .A2(new_n13553_), .ZN(new_n13554_));
  INV_X1     g13490(.I(new_n13554_), .ZN(new_n13555_));
  NOR2_X1    g13491(.A1(new_n13555_), .A2(new_n13549_), .ZN(new_n13556_));
  XOR2_X1    g13492(.A1(new_n13548_), .A2(new_n74_), .Z(new_n13557_));
  NOR2_X1    g13493(.A1(new_n13557_), .A2(new_n13554_), .ZN(new_n13558_));
  INV_X1     g13494(.I(new_n13558_), .ZN(new_n13559_));
  OAI21_X1   g13495(.A1(new_n13544_), .A2(new_n13556_), .B(new_n13559_), .ZN(new_n13560_));
  AOI21_X1   g13496(.A1(new_n12970_), .A2(new_n12940_), .B(new_n12936_), .ZN(new_n13561_));
  NOR3_X1    g13497(.A1(new_n10840_), .A2(new_n10795_), .A3(new_n10846_), .ZN(new_n13562_));
  NOR4_X1    g13498(.A1(new_n12945_), .A2(new_n9479_), .A3(new_n13562_), .A4(new_n13561_), .ZN(new_n13563_));
  NOR2_X1    g13499(.A1(new_n13562_), .A2(new_n13561_), .ZN(new_n13564_));
  AOI21_X1   g13500(.A1(new_n13564_), .A2(new_n12968_), .B(new_n9478_), .ZN(new_n13565_));
  NOR2_X1    g13501(.A1(new_n13565_), .A2(new_n13563_), .ZN(new_n13566_));
  OAI22_X1   g13502(.A1(new_n10844_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n10846_), .ZN(new_n13567_));
  NAND2_X1   g13503(.A1(new_n9479_), .A2(new_n2750_), .ZN(new_n13568_));
  AOI21_X1   g13504(.A1(new_n13568_), .A2(new_n13567_), .B(new_n2737_), .ZN(new_n13569_));
  NAND2_X1   g13505(.A1(new_n13566_), .A2(new_n13569_), .ZN(new_n13570_));
  XOR2_X1    g13506(.A1(new_n13570_), .A2(new_n74_), .Z(new_n13571_));
  INV_X1     g13507(.I(new_n12872_), .ZN(new_n13572_));
  OAI21_X1   g13508(.A1(new_n12896_), .A2(new_n12897_), .B(new_n13572_), .ZN(new_n13573_));
  XOR2_X1    g13509(.A1(new_n12887_), .A2(new_n12894_), .Z(new_n13574_));
  NAND2_X1   g13510(.A1(new_n13574_), .A2(new_n12872_), .ZN(new_n13575_));
  NAND2_X1   g13511(.A1(new_n13573_), .A2(new_n13575_), .ZN(new_n13576_));
  NOR2_X1    g13512(.A1(new_n13571_), .A2(new_n13576_), .ZN(new_n13577_));
  INV_X1     g13513(.I(new_n13577_), .ZN(new_n13578_));
  XOR2_X1    g13514(.A1(new_n13570_), .A2(\a[29] ), .Z(new_n13579_));
  INV_X1     g13515(.I(new_n13576_), .ZN(new_n13580_));
  NOR2_X1    g13516(.A1(new_n13579_), .A2(new_n13580_), .ZN(new_n13581_));
  AOI21_X1   g13517(.A1(new_n13560_), .A2(new_n13578_), .B(new_n13581_), .ZN(new_n13582_));
  NAND2_X1   g13518(.A1(new_n13495_), .A2(new_n13499_), .ZN(new_n13583_));
  AOI21_X1   g13519(.A1(new_n13582_), .A2(new_n13583_), .B(new_n13500_), .ZN(new_n13584_));
  OAI21_X1   g13520(.A1(new_n13483_), .A2(new_n13584_), .B(new_n13490_), .ZN(new_n13585_));
  INV_X1     g13521(.I(new_n13585_), .ZN(new_n13586_));
  AND2_X2    g13522(.A1(new_n13004_), .A2(new_n13002_), .Z(new_n13587_));
  XOR2_X1    g13523(.A1(new_n12979_), .A2(new_n13001_), .Z(new_n13588_));
  NAND2_X1   g13524(.A1(new_n13588_), .A2(new_n12967_), .ZN(new_n13589_));
  OAI21_X1   g13525(.A1(new_n12967_), .A2(new_n13587_), .B(new_n13589_), .ZN(new_n13590_));
  INV_X1     g13526(.I(new_n13590_), .ZN(new_n13591_));
  NOR2_X1    g13527(.A1(new_n13065_), .A2(new_n13062_), .ZN(new_n13592_));
  OAI22_X1   g13528(.A1(new_n10861_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n10853_), .ZN(new_n13593_));
  NAND2_X1   g13529(.A1(new_n8785_), .A2(new_n2750_), .ZN(new_n13594_));
  AOI21_X1   g13530(.A1(new_n13594_), .A2(new_n13593_), .B(new_n2737_), .ZN(new_n13595_));
  NAND2_X1   g13531(.A1(new_n13592_), .A2(new_n13595_), .ZN(new_n13596_));
  XOR2_X1    g13532(.A1(new_n13596_), .A2(\a[29] ), .Z(new_n13597_));
  NAND2_X1   g13533(.A1(new_n13591_), .A2(new_n13597_), .ZN(new_n13598_));
  NOR2_X1    g13534(.A1(new_n13591_), .A2(new_n13597_), .ZN(new_n13599_));
  AOI21_X1   g13535(.A1(new_n13586_), .A2(new_n13598_), .B(new_n13599_), .ZN(new_n13600_));
  NAND2_X1   g13536(.A1(new_n13031_), .A2(new_n13029_), .ZN(new_n13601_));
  NAND2_X1   g13537(.A1(new_n13601_), .A2(new_n13005_), .ZN(new_n13602_));
  XNOR2_X1   g13538(.A1(new_n13021_), .A2(new_n13028_), .ZN(new_n13603_));
  OAI21_X1   g13539(.A1(new_n13005_), .A2(new_n13603_), .B(new_n13602_), .ZN(new_n13604_));
  OAI22_X1   g13540(.A1(new_n8784_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n10861_), .ZN(new_n13605_));
  NAND2_X1   g13541(.A1(new_n8779_), .A2(new_n2750_), .ZN(new_n13606_));
  AOI21_X1   g13542(.A1(new_n13606_), .A2(new_n13605_), .B(new_n2737_), .ZN(new_n13607_));
  NAND2_X1   g13543(.A1(new_n12814_), .A2(new_n13607_), .ZN(new_n13608_));
  XOR2_X1    g13544(.A1(new_n13608_), .A2(new_n74_), .Z(new_n13609_));
  NOR2_X1    g13545(.A1(new_n13609_), .A2(new_n13604_), .ZN(new_n13610_));
  NAND2_X1   g13546(.A1(new_n13609_), .A2(new_n13604_), .ZN(new_n13611_));
  OAI21_X1   g13547(.A1(new_n13600_), .A2(new_n13610_), .B(new_n13611_), .ZN(new_n13612_));
  NAND2_X1   g13548(.A1(new_n13056_), .A2(new_n13053_), .ZN(new_n13613_));
  NAND2_X1   g13549(.A1(new_n13032_), .A2(new_n13613_), .ZN(new_n13614_));
  XNOR2_X1   g13550(.A1(new_n13044_), .A2(new_n13052_), .ZN(new_n13615_));
  OAI21_X1   g13551(.A1(new_n13032_), .A2(new_n13615_), .B(new_n13614_), .ZN(new_n13616_));
  AOI22_X1   g13552(.A1(new_n8779_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n8785_), .ZN(new_n13617_));
  NOR2_X1    g13553(.A1(new_n10871_), .A2(new_n3175_), .ZN(new_n13618_));
  OAI21_X1   g13554(.A1(new_n13618_), .A2(new_n13617_), .B(new_n2736_), .ZN(new_n13619_));
  NOR2_X1    g13555(.A1(new_n11794_), .A2(new_n13619_), .ZN(new_n13620_));
  XOR2_X1    g13556(.A1(new_n13620_), .A2(\a[29] ), .Z(new_n13621_));
  OR2_X2     g13557(.A1(new_n13621_), .A2(new_n13616_), .Z(new_n13622_));
  NAND2_X1   g13558(.A1(new_n13621_), .A2(new_n13616_), .ZN(new_n13623_));
  INV_X1     g13559(.I(new_n13623_), .ZN(new_n13624_));
  AOI21_X1   g13560(.A1(new_n13612_), .A2(new_n13622_), .B(new_n13624_), .ZN(new_n13625_));
  INV_X1     g13561(.I(new_n13625_), .ZN(new_n13626_));
  NAND2_X1   g13562(.A1(new_n13057_), .A2(new_n13083_), .ZN(new_n13627_));
  NAND2_X1   g13563(.A1(new_n13085_), .A2(new_n13627_), .ZN(new_n13628_));
  INV_X1     g13564(.I(new_n13628_), .ZN(new_n13629_));
  OAI22_X1   g13565(.A1(new_n10871_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8778_), .ZN(new_n13630_));
  NAND2_X1   g13566(.A1(new_n10886_), .A2(new_n2750_), .ZN(new_n13631_));
  AOI21_X1   g13567(.A1(new_n13631_), .A2(new_n13630_), .B(new_n2737_), .ZN(new_n13632_));
  NAND2_X1   g13568(.A1(new_n13103_), .A2(new_n13632_), .ZN(new_n13633_));
  XOR2_X1    g13569(.A1(new_n13633_), .A2(\a[29] ), .Z(new_n13634_));
  NAND2_X1   g13570(.A1(new_n13629_), .A2(new_n13634_), .ZN(new_n13635_));
  NAND2_X1   g13571(.A1(new_n13626_), .A2(new_n13635_), .ZN(new_n13636_));
  INV_X1     g13572(.I(new_n13634_), .ZN(new_n13637_));
  NAND2_X1   g13573(.A1(new_n13637_), .A2(new_n13628_), .ZN(new_n13638_));
  NAND2_X1   g13574(.A1(new_n13636_), .A2(new_n13638_), .ZN(new_n13639_));
  NOR2_X1    g13575(.A1(new_n13084_), .A2(new_n13080_), .ZN(new_n13640_));
  XOR2_X1    g13576(.A1(new_n13640_), .A2(new_n12807_), .Z(new_n13641_));
  XOR2_X1    g13577(.A1(new_n13641_), .A2(new_n12818_), .Z(new_n13642_));
  AOI22_X1   g13578(.A1(new_n10886_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n10872_), .ZN(new_n13643_));
  NOR2_X1    g13579(.A1(new_n10892_), .A2(new_n3175_), .ZN(new_n13644_));
  OAI21_X1   g13580(.A1(new_n13643_), .A2(new_n13644_), .B(new_n2736_), .ZN(new_n13645_));
  NOR2_X1    g13581(.A1(new_n12776_), .A2(new_n13645_), .ZN(new_n13646_));
  XOR2_X1    g13582(.A1(new_n13646_), .A2(new_n74_), .Z(new_n13647_));
  INV_X1     g13583(.I(new_n13647_), .ZN(new_n13648_));
  OR2_X2     g13584(.A1(new_n13642_), .A2(new_n13648_), .Z(new_n13649_));
  NAND2_X1   g13585(.A1(new_n13649_), .A2(new_n13639_), .ZN(new_n13650_));
  NAND2_X1   g13586(.A1(new_n13642_), .A2(new_n13648_), .ZN(new_n13651_));
  NAND2_X1   g13587(.A1(new_n13650_), .A2(new_n13651_), .ZN(new_n13652_));
  AOI22_X1   g13588(.A1(new_n3267_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n3323_), .ZN(new_n13653_));
  NOR2_X1    g13589(.A1(new_n8758_), .A2(new_n3318_), .ZN(new_n13654_));
  OAI21_X1   g13590(.A1(new_n13653_), .A2(new_n13654_), .B(new_n3259_), .ZN(new_n13655_));
  NOR2_X1    g13591(.A1(new_n12053_), .A2(new_n13655_), .ZN(new_n13656_));
  XOR2_X1    g13592(.A1(new_n13656_), .A2(new_n72_), .Z(new_n13657_));
  INV_X1     g13593(.I(new_n13657_), .ZN(new_n13658_));
  NAND2_X1   g13594(.A1(new_n13652_), .A2(new_n13658_), .ZN(new_n13659_));
  NAND2_X1   g13595(.A1(new_n13137_), .A2(new_n13139_), .ZN(new_n13660_));
  XOR2_X1    g13596(.A1(new_n13093_), .A2(new_n13087_), .Z(new_n13661_));
  NAND2_X1   g13597(.A1(new_n13660_), .A2(new_n13661_), .ZN(new_n13662_));
  NAND2_X1   g13598(.A1(new_n13096_), .A2(new_n13099_), .ZN(new_n13663_));
  NAND3_X1   g13599(.A1(new_n13137_), .A2(new_n13139_), .A3(new_n13663_), .ZN(new_n13664_));
  NOR2_X1    g13600(.A1(new_n13652_), .A2(new_n13658_), .ZN(new_n13665_));
  INV_X1     g13601(.I(new_n13665_), .ZN(new_n13666_));
  NAND3_X1   g13602(.A1(new_n13662_), .A2(new_n13664_), .A3(new_n13666_), .ZN(new_n13667_));
  NAND2_X1   g13603(.A1(new_n13667_), .A2(new_n13659_), .ZN(new_n13668_));
  OAI22_X1   g13604(.A1(new_n8751_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n10924_), .ZN(new_n13669_));
  NAND2_X1   g13605(.A1(new_n8736_), .A2(new_n3312_), .ZN(new_n13670_));
  AOI21_X1   g13606(.A1(new_n13670_), .A2(new_n13669_), .B(new_n3302_), .ZN(new_n13671_));
  NAND2_X1   g13607(.A1(new_n12118_), .A2(new_n13671_), .ZN(new_n13672_));
  XOR2_X1    g13608(.A1(new_n13672_), .A2(\a[23] ), .Z(new_n13673_));
  INV_X1     g13609(.I(new_n13673_), .ZN(new_n13674_));
  NOR2_X1    g13610(.A1(new_n13668_), .A2(new_n13674_), .ZN(new_n13675_));
  INV_X1     g13611(.I(new_n13675_), .ZN(new_n13676_));
  AOI21_X1   g13612(.A1(new_n13667_), .A2(new_n13659_), .B(new_n13673_), .ZN(new_n13677_));
  AOI21_X1   g13613(.A1(new_n13479_), .A2(new_n13676_), .B(new_n13677_), .ZN(new_n13678_));
  OAI22_X1   g13614(.A1(new_n8710_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n8718_), .ZN(new_n13679_));
  NAND2_X1   g13615(.A1(new_n8702_), .A2(new_n4096_), .ZN(new_n13680_));
  AOI21_X1   g13616(.A1(new_n13680_), .A2(new_n13679_), .B(new_n4095_), .ZN(new_n13681_));
  NAND2_X1   g13617(.A1(new_n12205_), .A2(new_n13681_), .ZN(new_n13682_));
  XOR2_X1    g13618(.A1(new_n13682_), .A2(\a[20] ), .Z(new_n13683_));
  NOR2_X1    g13619(.A1(new_n13678_), .A2(new_n13683_), .ZN(new_n13684_));
  NAND2_X1   g13620(.A1(new_n13678_), .A2(new_n13683_), .ZN(new_n13685_));
  NAND3_X1   g13621(.A1(new_n13292_), .A2(new_n13347_), .A3(new_n13295_), .ZN(new_n13686_));
  OAI21_X1   g13622(.A1(new_n13341_), .A2(new_n13342_), .B(new_n13319_), .ZN(new_n13687_));
  NAND3_X1   g13623(.A1(new_n13687_), .A2(new_n13686_), .A3(new_n13348_), .ZN(new_n13688_));
  NOR3_X1    g13624(.A1(new_n13341_), .A2(new_n13342_), .A3(new_n13319_), .ZN(new_n13689_));
  AOI21_X1   g13625(.A1(new_n13292_), .A2(new_n13295_), .B(new_n13347_), .ZN(new_n13690_));
  OAI21_X1   g13626(.A1(new_n13690_), .A2(new_n13689_), .B(new_n13324_), .ZN(new_n13691_));
  NAND2_X1   g13627(.A1(new_n13691_), .A2(new_n13688_), .ZN(new_n13692_));
  AOI21_X1   g13628(.A1(new_n13692_), .A2(new_n13685_), .B(new_n13684_), .ZN(new_n13693_));
  OAI22_X1   g13629(.A1(new_n3775_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n3769_), .ZN(new_n13694_));
  NAND2_X1   g13630(.A1(new_n8696_), .A2(new_n4096_), .ZN(new_n13695_));
  AOI21_X1   g13631(.A1(new_n13694_), .A2(new_n13695_), .B(new_n4095_), .ZN(new_n13696_));
  NAND2_X1   g13632(.A1(new_n11595_), .A2(new_n13696_), .ZN(new_n13697_));
  XOR2_X1    g13633(.A1(new_n13697_), .A2(\a[20] ), .Z(new_n13698_));
  NOR2_X1    g13634(.A1(new_n13693_), .A2(new_n13698_), .ZN(new_n13699_));
  NOR3_X1    g13635(.A1(new_n13446_), .A2(new_n13333_), .A3(new_n13444_), .ZN(new_n13700_));
  AOI21_X1   g13636(.A1(new_n13340_), .A2(new_n13338_), .B(new_n13334_), .ZN(new_n13701_));
  OAI21_X1   g13637(.A1(new_n13700_), .A2(new_n13701_), .B(new_n13327_), .ZN(new_n13702_));
  NAND3_X1   g13638(.A1(new_n13340_), .A2(new_n13334_), .A3(new_n13338_), .ZN(new_n13703_));
  OAI21_X1   g13639(.A1(new_n13446_), .A2(new_n13444_), .B(new_n13333_), .ZN(new_n13704_));
  NAND3_X1   g13640(.A1(new_n13704_), .A2(new_n13703_), .A3(new_n13328_), .ZN(new_n13705_));
  NAND2_X1   g13641(.A1(new_n13702_), .A2(new_n13705_), .ZN(new_n13706_));
  AOI22_X1   g13642(.A1(new_n13691_), .A2(new_n13688_), .B1(new_n13678_), .B2(new_n13683_), .ZN(new_n13707_));
  INV_X1     g13643(.I(new_n13698_), .ZN(new_n13708_));
  NOR3_X1    g13644(.A1(new_n13707_), .A2(new_n13684_), .A3(new_n13708_), .ZN(new_n13709_));
  AOI21_X1   g13645(.A1(new_n13706_), .A2(new_n13709_), .B(new_n13699_), .ZN(new_n13710_));
  OAI22_X1   g13646(.A1(new_n8673_), .A2(new_n4297_), .B1(new_n8687_), .B2(new_n4291_), .ZN(new_n13711_));
  NAND2_X1   g13647(.A1(new_n8662_), .A2(new_n4469_), .ZN(new_n13712_));
  AOI21_X1   g13648(.A1(new_n13712_), .A2(new_n13711_), .B(new_n4468_), .ZN(new_n13713_));
  NAND2_X1   g13649(.A1(new_n11624_), .A2(new_n13713_), .ZN(new_n13714_));
  XOR2_X1    g13650(.A1(new_n13714_), .A2(\a[17] ), .Z(new_n13715_));
  AOI22_X1   g13651(.A1(new_n13710_), .A2(new_n13715_), .B1(new_n13467_), .B2(new_n13472_), .ZN(new_n13716_));
  NOR2_X1    g13652(.A1(new_n13710_), .A2(new_n13715_), .ZN(new_n13717_));
  AOI22_X1   g13653(.A1(new_n11311_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n11272_), .ZN(new_n13718_));
  NOR2_X1    g13654(.A1(new_n11264_), .A2(new_n6091_), .ZN(new_n13719_));
  OAI21_X1   g13655(.A1(new_n13719_), .A2(new_n13718_), .B(new_n6081_), .ZN(new_n13720_));
  NOR2_X1    g13656(.A1(new_n11310_), .A2(new_n13720_), .ZN(new_n13721_));
  XOR2_X1    g13657(.A1(new_n13721_), .A2(new_n3521_), .Z(new_n13722_));
  INV_X1     g13658(.I(new_n13722_), .ZN(new_n13723_));
  NOR3_X1    g13659(.A1(new_n13716_), .A2(new_n13717_), .A3(new_n13723_), .ZN(new_n13724_));
  INV_X1     g13660(.I(new_n13724_), .ZN(new_n13725_));
  NAND2_X1   g13661(.A1(new_n13449_), .A2(new_n13358_), .ZN(new_n13726_));
  AOI21_X1   g13662(.A1(new_n13726_), .A2(new_n13361_), .B(new_n13468_), .ZN(new_n13727_));
  AOI21_X1   g13663(.A1(new_n13469_), .A2(new_n13470_), .B(new_n13465_), .ZN(new_n13728_));
  INV_X1     g13664(.I(new_n13699_), .ZN(new_n13729_));
  AOI21_X1   g13665(.A1(new_n13704_), .A2(new_n13703_), .B(new_n13328_), .ZN(new_n13730_));
  NOR3_X1    g13666(.A1(new_n13700_), .A2(new_n13701_), .A3(new_n13327_), .ZN(new_n13731_));
  OAI21_X1   g13667(.A1(new_n13731_), .A2(new_n13730_), .B(new_n13709_), .ZN(new_n13732_));
  NAND2_X1   g13668(.A1(new_n13732_), .A2(new_n13729_), .ZN(new_n13733_));
  INV_X1     g13669(.I(new_n13715_), .ZN(new_n13734_));
  OAI22_X1   g13670(.A1(new_n13733_), .A2(new_n13734_), .B1(new_n13727_), .B2(new_n13728_), .ZN(new_n13735_));
  INV_X1     g13671(.I(new_n13717_), .ZN(new_n13736_));
  AOI21_X1   g13672(.A1(new_n13736_), .A2(new_n13735_), .B(new_n13722_), .ZN(new_n13737_));
  AOI21_X1   g13673(.A1(new_n13725_), .A2(new_n13464_), .B(new_n13737_), .ZN(new_n13738_));
  OAI22_X1   g13674(.A1(new_n11264_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n11277_), .ZN(new_n13739_));
  NAND2_X1   g13675(.A1(new_n11346_), .A2(new_n6090_), .ZN(new_n13740_));
  AOI21_X1   g13676(.A1(new_n13739_), .A2(new_n13740_), .B(new_n6082_), .ZN(new_n13741_));
  NAND2_X1   g13677(.A1(new_n11757_), .A2(new_n13741_), .ZN(new_n13742_));
  XOR2_X1    g13678(.A1(new_n13742_), .A2(\a[14] ), .Z(new_n13743_));
  NOR2_X1    g13679(.A1(new_n13738_), .A2(new_n13743_), .ZN(new_n13744_));
  INV_X1     g13680(.I(new_n13738_), .ZN(new_n13745_));
  INV_X1     g13681(.I(new_n13743_), .ZN(new_n13746_));
  XOR2_X1    g13682(.A1(new_n13201_), .A2(new_n13374_), .Z(new_n13747_));
  NAND2_X1   g13683(.A1(new_n13381_), .A2(new_n13747_), .ZN(new_n13748_));
  XOR2_X1    g13684(.A1(new_n13201_), .A2(new_n13374_), .Z(new_n13749_));
  OAI21_X1   g13685(.A1(new_n13381_), .A2(new_n13749_), .B(new_n13748_), .ZN(new_n13750_));
  XOR2_X1    g13686(.A1(new_n13750_), .A2(new_n13369_), .Z(new_n13751_));
  NOR3_X1    g13687(.A1(new_n13751_), .A2(new_n13745_), .A3(new_n13746_), .ZN(new_n13752_));
  NOR2_X1    g13688(.A1(new_n13752_), .A2(new_n13744_), .ZN(new_n13753_));
  OAI22_X1   g13689(.A1(new_n11369_), .A2(new_n4716_), .B1(new_n4710_), .B2(new_n11461_), .ZN(new_n13754_));
  NAND2_X1   g13690(.A1(new_n11694_), .A2(new_n4720_), .ZN(new_n13755_));
  AOI21_X1   g13691(.A1(new_n13754_), .A2(new_n13755_), .B(new_n4707_), .ZN(new_n13756_));
  NAND2_X1   g13692(.A1(new_n12720_), .A2(new_n13756_), .ZN(new_n13757_));
  XOR2_X1    g13693(.A1(new_n13757_), .A2(\a[11] ), .Z(new_n13758_));
  NAND2_X1   g13694(.A1(new_n13753_), .A2(new_n13758_), .ZN(new_n13759_));
  INV_X1     g13695(.I(new_n13758_), .ZN(new_n13760_));
  OAI21_X1   g13696(.A1(new_n13752_), .A2(new_n13744_), .B(new_n13760_), .ZN(new_n13761_));
  INV_X1     g13697(.I(new_n13761_), .ZN(new_n13762_));
  AOI21_X1   g13698(.A1(new_n13434_), .A2(new_n13759_), .B(new_n13762_), .ZN(new_n13763_));
  NOR3_X1    g13699(.A1(new_n13419_), .A2(new_n13422_), .A3(new_n13763_), .ZN(new_n13764_));
  OAI21_X1   g13700(.A1(new_n13419_), .A2(new_n13422_), .B(new_n13763_), .ZN(new_n13765_));
  INV_X1     g13701(.I(new_n13765_), .ZN(new_n13766_));
  NOR2_X1    g13702(.A1(new_n13766_), .A2(new_n13764_), .ZN(new_n13767_));
  AOI21_X1   g13703(.A1(new_n13390_), .A2(new_n13397_), .B(new_n13430_), .ZN(new_n13768_));
  NAND2_X1   g13704(.A1(new_n13395_), .A2(new_n13389_), .ZN(new_n13769_));
  NAND2_X1   g13705(.A1(new_n13384_), .A2(new_n13396_), .ZN(new_n13770_));
  AOI21_X1   g13706(.A1(new_n13770_), .A2(new_n13769_), .B(new_n13267_), .ZN(new_n13771_));
  NOR2_X1    g13707(.A1(new_n13768_), .A2(new_n13771_), .ZN(new_n13772_));
  AOI21_X1   g13708(.A1(new_n13759_), .A2(new_n13761_), .B(new_n13772_), .ZN(new_n13773_));
  OAI21_X1   g13709(.A1(new_n13752_), .A2(new_n13744_), .B(new_n13758_), .ZN(new_n13774_));
  NAND2_X1   g13710(.A1(new_n13753_), .A2(new_n13760_), .ZN(new_n13775_));
  AOI21_X1   g13711(.A1(new_n13774_), .A2(new_n13775_), .B(new_n13434_), .ZN(new_n13776_));
  NOR2_X1    g13712(.A1(new_n13773_), .A2(new_n13776_), .ZN(new_n13777_));
  OAI21_X1   g13713(.A1(new_n13737_), .A2(new_n13724_), .B(new_n13464_), .ZN(new_n13778_));
  OAI21_X1   g13714(.A1(new_n13450_), .A2(new_n13451_), .B(new_n13452_), .ZN(new_n13779_));
  AOI21_X1   g13715(.A1(new_n13367_), .A2(new_n13779_), .B(new_n13460_), .ZN(new_n13780_));
  OAI21_X1   g13716(.A1(new_n13450_), .A2(new_n13451_), .B(new_n13366_), .ZN(new_n13781_));
  NAND3_X1   g13717(.A1(new_n13360_), .A2(new_n13361_), .A3(new_n13452_), .ZN(new_n13782_));
  AOI21_X1   g13718(.A1(new_n13782_), .A2(new_n13781_), .B(new_n13284_), .ZN(new_n13783_));
  NOR2_X1    g13719(.A1(new_n13780_), .A2(new_n13783_), .ZN(new_n13784_));
  AOI21_X1   g13720(.A1(new_n13736_), .A2(new_n13735_), .B(new_n13723_), .ZN(new_n13785_));
  NOR3_X1    g13721(.A1(new_n13716_), .A2(new_n13717_), .A3(new_n13722_), .ZN(new_n13786_));
  OAI21_X1   g13722(.A1(new_n13785_), .A2(new_n13786_), .B(new_n13784_), .ZN(new_n13787_));
  NAND2_X1   g13723(.A1(new_n13787_), .A2(new_n13778_), .ZN(new_n13788_));
  INV_X1     g13724(.I(new_n13683_), .ZN(new_n13789_));
  NAND2_X1   g13725(.A1(new_n13687_), .A2(new_n13686_), .ZN(new_n13790_));
  NOR2_X1    g13726(.A1(new_n13678_), .A2(new_n13790_), .ZN(new_n13791_));
  AOI21_X1   g13727(.A1(new_n13476_), .A2(new_n13477_), .B(new_n13316_), .ZN(new_n13792_));
  NOR3_X1    g13728(.A1(new_n13474_), .A2(new_n13473_), .A3(new_n13300_), .ZN(new_n13793_));
  OAI21_X1   g13729(.A1(new_n13793_), .A2(new_n13792_), .B(new_n13676_), .ZN(new_n13794_));
  INV_X1     g13730(.I(new_n13677_), .ZN(new_n13795_));
  NAND2_X1   g13731(.A1(new_n13794_), .A2(new_n13795_), .ZN(new_n13796_));
  NOR2_X1    g13732(.A1(new_n13690_), .A2(new_n13689_), .ZN(new_n13797_));
  NOR2_X1    g13733(.A1(new_n13797_), .A2(new_n13796_), .ZN(new_n13798_));
  OAI21_X1   g13734(.A1(new_n13798_), .A2(new_n13791_), .B(new_n13324_), .ZN(new_n13799_));
  NAND2_X1   g13735(.A1(new_n13797_), .A2(new_n13796_), .ZN(new_n13800_));
  NAND2_X1   g13736(.A1(new_n13678_), .A2(new_n13790_), .ZN(new_n13801_));
  NAND3_X1   g13737(.A1(new_n13800_), .A2(new_n13801_), .A3(new_n13348_), .ZN(new_n13802_));
  AOI21_X1   g13738(.A1(new_n13799_), .A2(new_n13802_), .B(new_n13789_), .ZN(new_n13803_));
  AOI21_X1   g13739(.A1(new_n13800_), .A2(new_n13801_), .B(new_n13348_), .ZN(new_n13804_));
  NOR3_X1    g13740(.A1(new_n13798_), .A2(new_n13791_), .A3(new_n13324_), .ZN(new_n13805_));
  NOR3_X1    g13741(.A1(new_n13804_), .A2(new_n13805_), .A3(new_n13683_), .ZN(new_n13806_));
  NOR2_X1    g13742(.A1(new_n13675_), .A2(new_n13677_), .ZN(new_n13807_));
  INV_X1     g13743(.I(new_n13807_), .ZN(new_n13808_));
  OAI21_X1   g13744(.A1(new_n13793_), .A2(new_n13792_), .B(new_n13808_), .ZN(new_n13809_));
  XOR2_X1    g13745(.A1(new_n13668_), .A2(new_n13674_), .Z(new_n13810_));
  NAND3_X1   g13746(.A1(new_n13475_), .A2(new_n13478_), .A3(new_n13810_), .ZN(new_n13811_));
  NAND2_X1   g13747(.A1(new_n13662_), .A2(new_n13664_), .ZN(new_n13812_));
  XOR2_X1    g13748(.A1(new_n13652_), .A2(new_n13657_), .Z(new_n13813_));
  INV_X1     g13749(.I(new_n13813_), .ZN(new_n13814_));
  NAND2_X1   g13750(.A1(new_n13812_), .A2(new_n13814_), .ZN(new_n13815_));
  NAND2_X1   g13751(.A1(new_n13666_), .A2(new_n13659_), .ZN(new_n13816_));
  NAND3_X1   g13752(.A1(new_n13662_), .A2(new_n13664_), .A3(new_n13816_), .ZN(new_n13817_));
  NAND2_X1   g13753(.A1(new_n13815_), .A2(new_n13817_), .ZN(new_n13818_));
  XOR2_X1    g13754(.A1(new_n13621_), .A2(new_n13616_), .Z(new_n13819_));
  AND2_X2    g13755(.A1(new_n13612_), .A2(new_n13819_), .Z(new_n13820_));
  AOI21_X1   g13756(.A1(new_n13622_), .A2(new_n13623_), .B(new_n13612_), .ZN(new_n13821_));
  NOR2_X1    g13757(.A1(new_n13820_), .A2(new_n13821_), .ZN(new_n13822_));
  INV_X1     g13758(.I(new_n13822_), .ZN(new_n13823_));
  AOI22_X1   g13759(.A1(new_n10886_), .A2(new_n3267_), .B1(new_n10889_), .B2(new_n3323_), .ZN(new_n13824_));
  NOR2_X1    g13760(.A1(new_n10899_), .A2(new_n3318_), .ZN(new_n13825_));
  OAI21_X1   g13761(.A1(new_n13825_), .A2(new_n13824_), .B(new_n3259_), .ZN(new_n13826_));
  NOR2_X1    g13762(.A1(new_n11908_), .A2(new_n13826_), .ZN(new_n13827_));
  XOR2_X1    g13763(.A1(new_n13827_), .A2(new_n72_), .Z(new_n13828_));
  NOR2_X1    g13764(.A1(new_n13823_), .A2(new_n13828_), .ZN(new_n13829_));
  XNOR2_X1   g13765(.A1(new_n13628_), .A2(new_n13634_), .ZN(new_n13830_));
  NAND2_X1   g13766(.A1(new_n13626_), .A2(new_n13830_), .ZN(new_n13831_));
  NAND2_X1   g13767(.A1(new_n13635_), .A2(new_n13638_), .ZN(new_n13832_));
  NAND2_X1   g13768(.A1(new_n13832_), .A2(new_n13625_), .ZN(new_n13833_));
  NAND2_X1   g13769(.A1(new_n13831_), .A2(new_n13833_), .ZN(new_n13834_));
  AOI22_X1   g13770(.A1(new_n11899_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n10889_), .ZN(new_n13835_));
  NOR2_X1    g13771(.A1(new_n8774_), .A2(new_n3318_), .ZN(new_n13836_));
  OAI21_X1   g13772(.A1(new_n13836_), .A2(new_n13835_), .B(new_n3259_), .ZN(new_n13837_));
  NOR2_X1    g13773(.A1(new_n11945_), .A2(new_n13837_), .ZN(new_n13838_));
  XOR2_X1    g13774(.A1(new_n13838_), .A2(new_n72_), .Z(new_n13839_));
  NAND2_X1   g13775(.A1(new_n13834_), .A2(new_n13839_), .ZN(new_n13840_));
  NOR2_X1    g13776(.A1(new_n13834_), .A2(new_n13839_), .ZN(new_n13841_));
  AOI21_X1   g13777(.A1(new_n13829_), .A2(new_n13840_), .B(new_n13841_), .ZN(new_n13842_));
  XOR2_X1    g13778(.A1(new_n13642_), .A2(new_n13647_), .Z(new_n13843_));
  AOI21_X1   g13779(.A1(new_n13636_), .A2(new_n13638_), .B(new_n13843_), .ZN(new_n13844_));
  AOI21_X1   g13780(.A1(new_n13649_), .A2(new_n13651_), .B(new_n13639_), .ZN(new_n13845_));
  NOR2_X1    g13781(.A1(new_n13844_), .A2(new_n13845_), .ZN(new_n13846_));
  OAI22_X1   g13782(.A1(new_n8774_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n10899_), .ZN(new_n13847_));
  NAND2_X1   g13783(.A1(new_n11996_), .A2(new_n3317_), .ZN(new_n13848_));
  AOI21_X1   g13784(.A1(new_n13848_), .A2(new_n13847_), .B(new_n3260_), .ZN(new_n13849_));
  NAND2_X1   g13785(.A1(new_n12001_), .A2(new_n13849_), .ZN(new_n13850_));
  XOR2_X1    g13786(.A1(new_n13850_), .A2(\a[26] ), .Z(new_n13851_));
  INV_X1     g13787(.I(new_n13851_), .ZN(new_n13852_));
  NOR2_X1    g13788(.A1(new_n13846_), .A2(new_n13852_), .ZN(new_n13853_));
  NAND2_X1   g13789(.A1(new_n13846_), .A2(new_n13852_), .ZN(new_n13854_));
  OAI21_X1   g13790(.A1(new_n13842_), .A2(new_n13853_), .B(new_n13854_), .ZN(new_n13855_));
  OAI22_X1   g13791(.A1(new_n8751_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8745_), .ZN(new_n13856_));
  NAND2_X1   g13792(.A1(new_n10927_), .A2(new_n3312_), .ZN(new_n13857_));
  AOI21_X1   g13793(.A1(new_n13856_), .A2(new_n13857_), .B(new_n3302_), .ZN(new_n13858_));
  NAND2_X1   g13794(.A1(new_n12072_), .A2(new_n13858_), .ZN(new_n13859_));
  XOR2_X1    g13795(.A1(new_n13859_), .A2(\a[23] ), .Z(new_n13860_));
  INV_X1     g13796(.I(new_n13860_), .ZN(new_n13861_));
  OR2_X2     g13797(.A1(new_n13855_), .A2(new_n13861_), .Z(new_n13862_));
  NAND2_X1   g13798(.A1(new_n13818_), .A2(new_n13862_), .ZN(new_n13863_));
  NAND2_X1   g13799(.A1(new_n13855_), .A2(new_n13861_), .ZN(new_n13864_));
  NAND2_X1   g13800(.A1(new_n13863_), .A2(new_n13864_), .ZN(new_n13865_));
  INV_X1     g13801(.I(new_n13865_), .ZN(new_n13866_));
  OAI22_X1   g13802(.A1(new_n8725_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n8718_), .ZN(new_n13867_));
  NAND2_X1   g13803(.A1(new_n8711_), .A2(new_n4096_), .ZN(new_n13868_));
  AOI21_X1   g13804(.A1(new_n13868_), .A2(new_n13867_), .B(new_n4095_), .ZN(new_n13869_));
  NAND2_X1   g13805(.A1(new_n11536_), .A2(new_n13869_), .ZN(new_n13870_));
  XOR2_X1    g13806(.A1(new_n13870_), .A2(\a[20] ), .Z(new_n13871_));
  AOI22_X1   g13807(.A1(new_n13809_), .A2(new_n13811_), .B1(new_n13866_), .B2(new_n13871_), .ZN(new_n13872_));
  NOR2_X1    g13808(.A1(new_n13866_), .A2(new_n13871_), .ZN(new_n13873_));
  OAI22_X1   g13809(.A1(new_n8681_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8694_), .ZN(new_n13874_));
  NAND2_X1   g13810(.A1(new_n8688_), .A2(new_n4469_), .ZN(new_n13875_));
  AOI21_X1   g13811(.A1(new_n13875_), .A2(new_n13874_), .B(new_n4468_), .ZN(new_n13876_));
  NAND2_X1   g13812(.A1(new_n11420_), .A2(new_n13876_), .ZN(new_n13877_));
  XOR2_X1    g13813(.A1(new_n13877_), .A2(\a[17] ), .Z(new_n13878_));
  INV_X1     g13814(.I(new_n13878_), .ZN(new_n13879_));
  NOR3_X1    g13815(.A1(new_n13872_), .A2(new_n13873_), .A3(new_n13879_), .ZN(new_n13880_));
  INV_X1     g13816(.I(new_n13880_), .ZN(new_n13881_));
  OAI21_X1   g13817(.A1(new_n13806_), .A2(new_n13803_), .B(new_n13881_), .ZN(new_n13882_));
  AOI21_X1   g13818(.A1(new_n13475_), .A2(new_n13478_), .B(new_n13807_), .ZN(new_n13883_));
  XOR2_X1    g13819(.A1(new_n13668_), .A2(new_n13673_), .Z(new_n13884_));
  NOR3_X1    g13820(.A1(new_n13793_), .A2(new_n13792_), .A3(new_n13884_), .ZN(new_n13885_));
  INV_X1     g13821(.I(new_n13871_), .ZN(new_n13886_));
  OAI22_X1   g13822(.A1(new_n13885_), .A2(new_n13883_), .B1(new_n13865_), .B2(new_n13886_), .ZN(new_n13887_));
  INV_X1     g13823(.I(new_n13873_), .ZN(new_n13888_));
  AOI21_X1   g13824(.A1(new_n13887_), .A2(new_n13888_), .B(new_n13878_), .ZN(new_n13889_));
  INV_X1     g13825(.I(new_n13889_), .ZN(new_n13890_));
  OAI22_X1   g13826(.A1(new_n4291_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n4297_), .ZN(new_n13891_));
  NAND2_X1   g13827(.A1(new_n8674_), .A2(new_n4469_), .ZN(new_n13892_));
  AOI21_X1   g13828(.A1(new_n13892_), .A2(new_n13891_), .B(new_n4468_), .ZN(new_n13893_));
  NAND2_X1   g13829(.A1(new_n11431_), .A2(new_n13893_), .ZN(new_n13894_));
  XOR2_X1    g13830(.A1(new_n13894_), .A2(\a[17] ), .Z(new_n13895_));
  AOI21_X1   g13831(.A1(new_n13882_), .A2(new_n13890_), .B(new_n13895_), .ZN(new_n13896_));
  NOR3_X1    g13832(.A1(new_n13693_), .A2(new_n13700_), .A3(new_n13701_), .ZN(new_n13897_));
  NAND2_X1   g13833(.A1(new_n13796_), .A2(new_n13789_), .ZN(new_n13898_));
  NOR2_X1    g13834(.A1(new_n13796_), .A2(new_n13789_), .ZN(new_n13899_));
  NOR3_X1    g13835(.A1(new_n13690_), .A2(new_n13689_), .A3(new_n13324_), .ZN(new_n13900_));
  AOI21_X1   g13836(.A1(new_n13687_), .A2(new_n13686_), .B(new_n13348_), .ZN(new_n13901_));
  NOR2_X1    g13837(.A1(new_n13900_), .A2(new_n13901_), .ZN(new_n13902_));
  OAI21_X1   g13838(.A1(new_n13902_), .A2(new_n13899_), .B(new_n13898_), .ZN(new_n13903_));
  AOI21_X1   g13839(.A1(new_n13703_), .A2(new_n13704_), .B(new_n13903_), .ZN(new_n13904_));
  OAI21_X1   g13840(.A1(new_n13904_), .A2(new_n13897_), .B(new_n13698_), .ZN(new_n13905_));
  NAND3_X1   g13841(.A1(new_n13903_), .A2(new_n13703_), .A3(new_n13704_), .ZN(new_n13906_));
  OAI21_X1   g13842(.A1(new_n13700_), .A2(new_n13701_), .B(new_n13693_), .ZN(new_n13907_));
  NAND3_X1   g13843(.A1(new_n13907_), .A2(new_n13906_), .A3(new_n13708_), .ZN(new_n13908_));
  AOI21_X1   g13844(.A1(new_n13905_), .A2(new_n13908_), .B(new_n13328_), .ZN(new_n13909_));
  AOI21_X1   g13845(.A1(new_n13907_), .A2(new_n13906_), .B(new_n13708_), .ZN(new_n13910_));
  NOR3_X1    g13846(.A1(new_n13904_), .A2(new_n13698_), .A3(new_n13897_), .ZN(new_n13911_));
  NOR3_X1    g13847(.A1(new_n13911_), .A2(new_n13910_), .A3(new_n13327_), .ZN(new_n13912_));
  OAI21_X1   g13848(.A1(new_n13804_), .A2(new_n13805_), .B(new_n13683_), .ZN(new_n13913_));
  NAND3_X1   g13849(.A1(new_n13799_), .A2(new_n13802_), .A3(new_n13789_), .ZN(new_n13914_));
  AOI21_X1   g13850(.A1(new_n13913_), .A2(new_n13914_), .B(new_n13880_), .ZN(new_n13915_));
  INV_X1     g13851(.I(new_n13895_), .ZN(new_n13916_));
  NOR3_X1    g13852(.A1(new_n13915_), .A2(new_n13889_), .A3(new_n13916_), .ZN(new_n13917_));
  NOR3_X1    g13853(.A1(new_n13912_), .A2(new_n13909_), .A3(new_n13917_), .ZN(new_n13918_));
  OAI22_X1   g13854(.A1(new_n11284_), .A2(new_n6089_), .B1(new_n6094_), .B2(new_n11271_), .ZN(new_n13919_));
  NAND2_X1   g13855(.A1(new_n11311_), .A2(new_n6090_), .ZN(new_n13920_));
  AOI21_X1   g13856(.A1(new_n13919_), .A2(new_n13920_), .B(new_n6082_), .ZN(new_n13921_));
  NAND2_X1   g13857(.A1(new_n11391_), .A2(new_n13921_), .ZN(new_n13922_));
  XOR2_X1    g13858(.A1(new_n13922_), .A2(\a[14] ), .Z(new_n13923_));
  INV_X1     g13859(.I(new_n13923_), .ZN(new_n13924_));
  OAI21_X1   g13860(.A1(new_n13918_), .A2(new_n13896_), .B(new_n13924_), .ZN(new_n13925_));
  NOR3_X1    g13861(.A1(new_n13918_), .A2(new_n13896_), .A3(new_n13924_), .ZN(new_n13926_));
  NOR3_X1    g13862(.A1(new_n13727_), .A2(new_n13710_), .A3(new_n13728_), .ZN(new_n13927_));
  AOI21_X1   g13863(.A1(new_n13467_), .A2(new_n13472_), .B(new_n13733_), .ZN(new_n13928_));
  NOR3_X1    g13864(.A1(new_n13928_), .A2(new_n13927_), .A3(new_n13715_), .ZN(new_n13929_));
  NAND3_X1   g13865(.A1(new_n13733_), .A2(new_n13467_), .A3(new_n13472_), .ZN(new_n13930_));
  OAI21_X1   g13866(.A1(new_n13727_), .A2(new_n13728_), .B(new_n13710_), .ZN(new_n13931_));
  AOI21_X1   g13867(.A1(new_n13931_), .A2(new_n13930_), .B(new_n13734_), .ZN(new_n13932_));
  NOR2_X1    g13868(.A1(new_n13929_), .A2(new_n13932_), .ZN(new_n13933_));
  OAI21_X1   g13869(.A1(new_n13933_), .A2(new_n13926_), .B(new_n13925_), .ZN(new_n13934_));
  OAI22_X1   g13870(.A1(new_n11353_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n11345_), .ZN(new_n13935_));
  NAND2_X1   g13871(.A1(new_n11370_), .A2(new_n4709_), .ZN(new_n13936_));
  AOI21_X1   g13872(.A1(new_n13936_), .A2(new_n13935_), .B(new_n4707_), .ZN(new_n13937_));
  NAND2_X1   g13873(.A1(new_n11379_), .A2(new_n13937_), .ZN(new_n13938_));
  XOR2_X1    g13874(.A1(new_n13938_), .A2(\a[11] ), .Z(new_n13939_));
  INV_X1     g13875(.I(new_n13939_), .ZN(new_n13940_));
  OAI21_X1   g13876(.A1(new_n13934_), .A2(new_n13940_), .B(new_n13788_), .ZN(new_n13941_));
  NAND2_X1   g13877(.A1(new_n13934_), .A2(new_n13940_), .ZN(new_n13942_));
  NAND2_X1   g13878(.A1(new_n13941_), .A2(new_n13942_), .ZN(new_n13943_));
  NOR2_X1    g13879(.A1(new_n13750_), .A2(new_n13738_), .ZN(new_n13944_));
  OR2_X2     g13880(.A1(new_n13381_), .A2(new_n13749_), .Z(new_n13945_));
  AOI21_X1   g13881(.A1(new_n13945_), .A2(new_n13748_), .B(new_n13745_), .ZN(new_n13946_));
  OAI21_X1   g13882(.A1(new_n13944_), .A2(new_n13946_), .B(new_n13743_), .ZN(new_n13947_));
  INV_X1     g13883(.I(new_n13947_), .ZN(new_n13948_));
  NOR3_X1    g13884(.A1(new_n13944_), .A2(new_n13743_), .A3(new_n13946_), .ZN(new_n13949_));
  OAI21_X1   g13885(.A1(new_n13948_), .A2(new_n13949_), .B(new_n13369_), .ZN(new_n13950_));
  INV_X1     g13886(.I(new_n13369_), .ZN(new_n13951_));
  INV_X1     g13887(.I(new_n13949_), .ZN(new_n13952_));
  NAND3_X1   g13888(.A1(new_n13952_), .A2(new_n13951_), .A3(new_n13947_), .ZN(new_n13953_));
  OAI22_X1   g13889(.A1(new_n11353_), .A2(new_n4716_), .B1(new_n4710_), .B2(new_n11697_), .ZN(new_n13954_));
  NAND2_X1   g13890(.A1(new_n11370_), .A2(new_n4720_), .ZN(new_n13955_));
  AOI21_X1   g13891(.A1(new_n13955_), .A2(new_n13954_), .B(new_n4707_), .ZN(new_n13956_));
  NAND2_X1   g13892(.A1(new_n11700_), .A2(new_n13956_), .ZN(new_n13957_));
  XOR2_X1    g13893(.A1(new_n13957_), .A2(\a[11] ), .Z(new_n13958_));
  INV_X1     g13894(.I(new_n13958_), .ZN(new_n13959_));
  AOI21_X1   g13895(.A1(new_n13950_), .A2(new_n13953_), .B(new_n13959_), .ZN(new_n13960_));
  INV_X1     g13896(.I(new_n13960_), .ZN(new_n13961_));
  NAND2_X1   g13897(.A1(new_n13961_), .A2(new_n13943_), .ZN(new_n13962_));
  NAND3_X1   g13898(.A1(new_n13950_), .A2(new_n13953_), .A3(new_n13959_), .ZN(new_n13963_));
  NAND3_X1   g13899(.A1(new_n13777_), .A2(new_n13962_), .A3(new_n13963_), .ZN(new_n13964_));
  NOR2_X1    g13900(.A1(new_n9488_), .A2(new_n9503_), .ZN(new_n13965_));
  NOR3_X1    g13901(.A1(new_n11466_), .A2(new_n9485_), .A3(new_n13965_), .ZN(new_n13966_));
  NOR3_X1    g13902(.A1(new_n13966_), .A2(new_n9482_), .A3(new_n11461_), .ZN(new_n13967_));
  INV_X1     g13903(.I(new_n13967_), .ZN(new_n13968_));
  NOR4_X1    g13904(.A1(new_n11465_), .A2(new_n11467_), .A3(\a[2] ), .A4(new_n13968_), .ZN(new_n13969_));
  NOR2_X1    g13905(.A1(new_n11465_), .A2(new_n11467_), .ZN(new_n13970_));
  AOI21_X1   g13906(.A1(new_n13970_), .A2(new_n13967_), .B(new_n4387_), .ZN(new_n13971_));
  NOR2_X1    g13907(.A1(new_n13971_), .A2(new_n13969_), .ZN(new_n13972_));
  INV_X1     g13908(.I(new_n13972_), .ZN(new_n13973_));
  AOI22_X1   g13909(.A1(new_n11354_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n11346_), .ZN(new_n13974_));
  NOR2_X1    g13910(.A1(new_n11369_), .A2(new_n6839_), .ZN(new_n13975_));
  NOR2_X1    g13911(.A1(new_n13974_), .A2(new_n13975_), .ZN(new_n13976_));
  NOR4_X1    g13912(.A1(new_n11378_), .A2(new_n6836_), .A3(new_n11375_), .A4(new_n13976_), .ZN(new_n13977_));
  XOR2_X1    g13913(.A1(new_n13977_), .A2(\a[5] ), .Z(new_n13978_));
  OAI22_X1   g13914(.A1(new_n8751_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n8745_), .ZN(new_n13979_));
  NAND2_X1   g13915(.A1(new_n10927_), .A2(new_n4096_), .ZN(new_n13980_));
  AOI21_X1   g13916(.A1(new_n13979_), .A2(new_n13980_), .B(new_n4095_), .ZN(new_n13981_));
  NAND2_X1   g13917(.A1(new_n12072_), .A2(new_n13981_), .ZN(new_n13982_));
  XOR2_X1    g13918(.A1(new_n13982_), .A2(\a[20] ), .Z(new_n13983_));
  OAI22_X1   g13919(.A1(new_n8774_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n10899_), .ZN(new_n13984_));
  NAND2_X1   g13920(.A1(new_n11996_), .A2(new_n3312_), .ZN(new_n13985_));
  AOI21_X1   g13921(.A1(new_n13985_), .A2(new_n13984_), .B(new_n3302_), .ZN(new_n13986_));
  NAND2_X1   g13922(.A1(new_n12001_), .A2(new_n13986_), .ZN(new_n13987_));
  XOR2_X1    g13923(.A1(new_n13987_), .A2(\a[23] ), .Z(new_n13988_));
  XNOR2_X1   g13924(.A1(new_n13609_), .A2(new_n13604_), .ZN(new_n13989_));
  NOR2_X1    g13925(.A1(new_n13989_), .A2(new_n13600_), .ZN(new_n13990_));
  INV_X1     g13926(.I(new_n13610_), .ZN(new_n13991_));
  NAND2_X1   g13927(.A1(new_n13991_), .A2(new_n13611_), .ZN(new_n13992_));
  AOI21_X1   g13928(.A1(new_n13600_), .A2(new_n13992_), .B(new_n13990_), .ZN(new_n13993_));
  XOR2_X1    g13929(.A1(new_n13597_), .A2(new_n13590_), .Z(new_n13994_));
  NOR2_X1    g13930(.A1(new_n13585_), .A2(new_n13994_), .ZN(new_n13995_));
  INV_X1     g13931(.I(new_n13599_), .ZN(new_n13996_));
  NAND2_X1   g13932(.A1(new_n13996_), .A2(new_n13598_), .ZN(new_n13997_));
  NAND2_X1   g13933(.A1(new_n13997_), .A2(new_n13585_), .ZN(new_n13998_));
  INV_X1     g13934(.I(new_n13998_), .ZN(new_n13999_));
  OAI22_X1   g13935(.A1(new_n10871_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8778_), .ZN(new_n14000_));
  NAND2_X1   g13936(.A1(new_n10886_), .A2(new_n3317_), .ZN(new_n14001_));
  AOI21_X1   g13937(.A1(new_n14001_), .A2(new_n14000_), .B(new_n3260_), .ZN(new_n14002_));
  NAND2_X1   g13938(.A1(new_n13103_), .A2(new_n14002_), .ZN(new_n14003_));
  XOR2_X1    g13939(.A1(new_n14003_), .A2(\a[26] ), .Z(new_n14004_));
  OAI21_X1   g13940(.A1(new_n13999_), .A2(new_n13995_), .B(new_n14004_), .ZN(new_n14005_));
  INV_X1     g13941(.I(new_n13483_), .ZN(new_n14006_));
  NOR2_X1    g13942(.A1(new_n13584_), .A2(new_n14006_), .ZN(new_n14007_));
  NAND2_X1   g13943(.A1(new_n13584_), .A2(new_n14006_), .ZN(new_n14008_));
  INV_X1     g13944(.I(new_n14008_), .ZN(new_n14009_));
  OAI21_X1   g13945(.A1(new_n14009_), .A2(new_n14007_), .B(new_n13489_), .ZN(new_n14010_));
  INV_X1     g13946(.I(new_n13489_), .ZN(new_n14011_));
  INV_X1     g13947(.I(new_n14007_), .ZN(new_n14012_));
  NAND3_X1   g13948(.A1(new_n14012_), .A2(new_n14011_), .A3(new_n14008_), .ZN(new_n14013_));
  AOI22_X1   g13949(.A1(new_n8779_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n8785_), .ZN(new_n14014_));
  NOR2_X1    g13950(.A1(new_n10871_), .A2(new_n3318_), .ZN(new_n14015_));
  OAI21_X1   g13951(.A1(new_n14015_), .A2(new_n14014_), .B(new_n3259_), .ZN(new_n14016_));
  NOR2_X1    g13952(.A1(new_n11794_), .A2(new_n14016_), .ZN(new_n14017_));
  XOR2_X1    g13953(.A1(new_n14017_), .A2(new_n72_), .Z(new_n14018_));
  INV_X1     g13954(.I(new_n14018_), .ZN(new_n14019_));
  NAND3_X1   g13955(.A1(new_n14010_), .A2(new_n14013_), .A3(new_n14019_), .ZN(new_n14020_));
  INV_X1     g13956(.I(new_n13995_), .ZN(new_n14021_));
  INV_X1     g13957(.I(new_n14004_), .ZN(new_n14022_));
  NAND3_X1   g13958(.A1(new_n14021_), .A2(new_n14022_), .A3(new_n13998_), .ZN(new_n14023_));
  NAND3_X1   g13959(.A1(new_n14005_), .A2(new_n14023_), .A3(new_n14020_), .ZN(new_n14024_));
  AOI22_X1   g13960(.A1(new_n10886_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n10872_), .ZN(new_n14025_));
  NOR2_X1    g13961(.A1(new_n10892_), .A2(new_n3318_), .ZN(new_n14026_));
  OAI21_X1   g13962(.A1(new_n14025_), .A2(new_n14026_), .B(new_n3259_), .ZN(new_n14027_));
  NOR2_X1    g13963(.A1(new_n12776_), .A2(new_n14027_), .ZN(new_n14028_));
  XOR2_X1    g13964(.A1(new_n14028_), .A2(new_n72_), .Z(new_n14029_));
  INV_X1     g13965(.I(new_n14029_), .ZN(new_n14030_));
  AOI21_X1   g13966(.A1(new_n14024_), .A2(new_n14005_), .B(new_n14030_), .ZN(new_n14031_));
  NAND3_X1   g13967(.A1(new_n14024_), .A2(new_n14005_), .A3(new_n14030_), .ZN(new_n14032_));
  INV_X1     g13968(.I(new_n14032_), .ZN(new_n14033_));
  OAI21_X1   g13969(.A1(new_n14033_), .A2(new_n14031_), .B(new_n13993_), .ZN(new_n14034_));
  INV_X1     g13970(.I(new_n13993_), .ZN(new_n14035_));
  INV_X1     g13971(.I(new_n14031_), .ZN(new_n14036_));
  NAND3_X1   g13972(.A1(new_n14036_), .A2(new_n14032_), .A3(new_n14035_), .ZN(new_n14037_));
  NAND2_X1   g13973(.A1(new_n14037_), .A2(new_n14034_), .ZN(new_n14038_));
  OAI22_X1   g13974(.A1(new_n8778_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8784_), .ZN(new_n14039_));
  OAI21_X1   g13975(.A1(new_n10871_), .A2(new_n3780_), .B(new_n14039_), .ZN(new_n14040_));
  NAND4_X1   g13976(.A1(new_n11792_), .A2(new_n3301_), .A3(new_n11793_), .A4(new_n14040_), .ZN(new_n14041_));
  XOR2_X1    g13977(.A1(new_n14041_), .A2(new_n84_), .Z(new_n14042_));
  AOI22_X1   g13978(.A1(new_n12823_), .A2(new_n3267_), .B1(new_n3323_), .B2(new_n10800_), .ZN(new_n14043_));
  NOR2_X1    g13979(.A1(new_n10798_), .A2(new_n3318_), .ZN(new_n14044_));
  OAI21_X1   g13980(.A1(new_n14043_), .A2(new_n14044_), .B(new_n3259_), .ZN(new_n14045_));
  NOR2_X1    g13981(.A1(new_n13504_), .A2(new_n14045_), .ZN(new_n14046_));
  NAND2_X1   g13982(.A1(new_n14046_), .A2(new_n72_), .ZN(new_n14047_));
  OAI21_X1   g13983(.A1(new_n13504_), .A2(new_n14045_), .B(\a[26] ), .ZN(new_n14048_));
  AOI21_X1   g13984(.A1(new_n14047_), .A2(new_n14048_), .B(new_n13521_), .ZN(new_n14049_));
  AOI22_X1   g13985(.A1(new_n10794_), .A2(new_n3267_), .B1(new_n3323_), .B2(new_n12823_), .ZN(new_n14050_));
  AOI21_X1   g13986(.A1(new_n3317_), .A2(new_n10800_), .B(new_n14050_), .ZN(new_n14051_));
  NAND2_X1   g13987(.A1(new_n12830_), .A2(new_n3259_), .ZN(new_n14052_));
  NOR2_X1    g13988(.A1(new_n14052_), .A2(new_n14051_), .ZN(new_n14053_));
  NOR2_X1    g13989(.A1(new_n3257_), .A2(new_n3258_), .ZN(new_n14054_));
  OAI21_X1   g13990(.A1(new_n12826_), .A2(new_n3322_), .B(new_n14054_), .ZN(new_n14055_));
  NOR2_X1    g13991(.A1(new_n12847_), .A2(new_n14055_), .ZN(new_n14056_));
  XOR2_X1    g13992(.A1(new_n14056_), .A2(\a[26] ), .Z(new_n14057_));
  NOR2_X1    g13993(.A1(new_n12826_), .A2(new_n3257_), .ZN(new_n14058_));
  NOR4_X1    g13994(.A1(new_n14057_), .A2(new_n72_), .A3(new_n14053_), .A4(new_n14058_), .ZN(new_n14059_));
  INV_X1     g13995(.I(new_n14059_), .ZN(new_n14060_));
  NAND3_X1   g13996(.A1(new_n14047_), .A2(new_n13521_), .A3(new_n14048_), .ZN(new_n14061_));
  AOI21_X1   g13997(.A1(new_n14060_), .A2(new_n14061_), .B(new_n14049_), .ZN(new_n14062_));
  XOR2_X1    g13998(.A1(new_n13520_), .A2(new_n74_), .Z(new_n14063_));
  NOR2_X1    g13999(.A1(new_n13521_), .A2(new_n74_), .ZN(new_n14064_));
  INV_X1     g14000(.I(new_n14064_), .ZN(new_n14065_));
  XOR2_X1    g14001(.A1(new_n14063_), .A2(new_n14065_), .Z(new_n14066_));
  AOI22_X1   g14002(.A1(new_n9529_), .A2(new_n3323_), .B1(new_n10800_), .B2(new_n3267_), .ZN(new_n14067_));
  AOI21_X1   g14003(.A1(new_n10839_), .A2(new_n3317_), .B(new_n14067_), .ZN(new_n14068_));
  NOR3_X1    g14004(.A1(new_n13534_), .A2(new_n14068_), .A3(new_n3260_), .ZN(new_n14069_));
  NAND2_X1   g14005(.A1(new_n14069_), .A2(new_n72_), .ZN(new_n14070_));
  INV_X1     g14006(.I(new_n14070_), .ZN(new_n14071_));
  NOR2_X1    g14007(.A1(new_n14069_), .A2(new_n72_), .ZN(new_n14072_));
  NOR3_X1    g14008(.A1(new_n14066_), .A2(new_n14071_), .A3(new_n14072_), .ZN(new_n14073_));
  NOR2_X1    g14009(.A1(new_n14073_), .A2(new_n14062_), .ZN(new_n14074_));
  NAND2_X1   g14010(.A1(new_n14063_), .A2(new_n14065_), .ZN(new_n14075_));
  XOR2_X1    g14011(.A1(new_n13520_), .A2(\a[29] ), .Z(new_n14076_));
  NAND2_X1   g14012(.A1(new_n14076_), .A2(new_n14064_), .ZN(new_n14077_));
  NAND2_X1   g14013(.A1(new_n14075_), .A2(new_n14077_), .ZN(new_n14078_));
  INV_X1     g14014(.I(new_n14072_), .ZN(new_n14079_));
  AOI21_X1   g14015(.A1(new_n14070_), .A2(new_n14079_), .B(new_n14078_), .ZN(new_n14080_));
  NOR2_X1    g14016(.A1(new_n14074_), .A2(new_n14080_), .ZN(new_n14081_));
  INV_X1     g14017(.I(new_n13523_), .ZN(new_n14082_));
  NOR3_X1    g14018(.A1(new_n13516_), .A2(new_n13517_), .A3(new_n14082_), .ZN(new_n14083_));
  INV_X1     g14019(.I(new_n13517_), .ZN(new_n14084_));
  AOI21_X1   g14020(.A1(new_n14084_), .A2(new_n13515_), .B(new_n13523_), .ZN(new_n14085_));
  NOR2_X1    g14021(.A1(new_n14085_), .A2(new_n14083_), .ZN(new_n14086_));
  AOI22_X1   g14022(.A1(new_n10839_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n9529_), .ZN(new_n14087_));
  NOR2_X1    g14023(.A1(new_n10846_), .A2(new_n3318_), .ZN(new_n14088_));
  OAI21_X1   g14024(.A1(new_n14087_), .A2(new_n14088_), .B(new_n3259_), .ZN(new_n14089_));
  NOR2_X1    g14025(.A1(new_n12946_), .A2(new_n14089_), .ZN(new_n14090_));
  NAND2_X1   g14026(.A1(new_n14090_), .A2(new_n72_), .ZN(new_n14091_));
  INV_X1     g14027(.I(new_n14091_), .ZN(new_n14092_));
  NOR2_X1    g14028(.A1(new_n14090_), .A2(new_n72_), .ZN(new_n14093_));
  NOR3_X1    g14029(.A1(new_n14092_), .A2(new_n14086_), .A3(new_n14093_), .ZN(new_n14094_));
  OAI21_X1   g14030(.A1(new_n14092_), .A2(new_n14093_), .B(new_n14086_), .ZN(new_n14095_));
  OAI21_X1   g14031(.A1(new_n14081_), .A2(new_n14094_), .B(new_n14095_), .ZN(new_n14096_));
  INV_X1     g14032(.I(new_n13511_), .ZN(new_n14097_));
  AOI21_X1   g14033(.A1(new_n14097_), .A2(new_n13526_), .B(new_n13525_), .ZN(new_n14098_));
  INV_X1     g14034(.I(new_n13508_), .ZN(new_n14099_));
  OR3_X2     g14035(.A1(new_n14099_), .A2(new_n13501_), .A3(new_n13509_), .Z(new_n14100_));
  OAI21_X1   g14036(.A1(new_n14099_), .A2(new_n13509_), .B(new_n13501_), .ZN(new_n14101_));
  AOI21_X1   g14037(.A1(new_n14100_), .A2(new_n14101_), .B(new_n13524_), .ZN(new_n14102_));
  NOR2_X1    g14038(.A1(new_n14098_), .A2(new_n14102_), .ZN(new_n14103_));
  INV_X1     g14039(.I(new_n14103_), .ZN(new_n14104_));
  OAI22_X1   g14040(.A1(new_n10844_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n10846_), .ZN(new_n14105_));
  NAND2_X1   g14041(.A1(new_n9479_), .A2(new_n3317_), .ZN(new_n14106_));
  AOI21_X1   g14042(.A1(new_n14106_), .A2(new_n14105_), .B(new_n3260_), .ZN(new_n14107_));
  NAND2_X1   g14043(.A1(new_n13566_), .A2(new_n14107_), .ZN(new_n14108_));
  NOR2_X1    g14044(.A1(new_n14108_), .A2(\a[26] ), .ZN(new_n14109_));
  NAND2_X1   g14045(.A1(new_n14108_), .A2(\a[26] ), .ZN(new_n14110_));
  INV_X1     g14046(.I(new_n14110_), .ZN(new_n14111_));
  NOR2_X1    g14047(.A1(new_n14111_), .A2(new_n14109_), .ZN(new_n14112_));
  NAND2_X1   g14048(.A1(new_n14104_), .A2(new_n14112_), .ZN(new_n14113_));
  NOR2_X1    g14049(.A1(new_n14104_), .A2(new_n14112_), .ZN(new_n14114_));
  AOI21_X1   g14050(.A1(new_n14096_), .A2(new_n14113_), .B(new_n14114_), .ZN(new_n14115_));
  XOR2_X1    g14051(.A1(new_n13537_), .A2(new_n74_), .Z(new_n14116_));
  NOR2_X1    g14052(.A1(new_n14116_), .A2(new_n13540_), .ZN(new_n14117_));
  OAI21_X1   g14053(.A1(new_n14117_), .A2(new_n13543_), .B(new_n13528_), .ZN(new_n14118_));
  NOR2_X1    g14054(.A1(new_n13538_), .A2(new_n13540_), .ZN(new_n14119_));
  NOR2_X1    g14055(.A1(new_n14116_), .A2(new_n13541_), .ZN(new_n14120_));
  OAI21_X1   g14056(.A1(new_n14119_), .A2(new_n14120_), .B(new_n13527_), .ZN(new_n14121_));
  NAND2_X1   g14057(.A1(new_n14118_), .A2(new_n14121_), .ZN(new_n14122_));
  OAI22_X1   g14058(.A1(new_n9478_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n10846_), .ZN(new_n14123_));
  NAND2_X1   g14059(.A1(new_n10854_), .A2(new_n3317_), .ZN(new_n14124_));
  AOI21_X1   g14060(.A1(new_n14123_), .A2(new_n14124_), .B(new_n3260_), .ZN(new_n14125_));
  NAND2_X1   g14061(.A1(new_n13016_), .A2(new_n14125_), .ZN(new_n14126_));
  XOR2_X1    g14062(.A1(new_n14126_), .A2(new_n72_), .Z(new_n14127_));
  NOR2_X1    g14063(.A1(new_n14122_), .A2(new_n14127_), .ZN(new_n14128_));
  NAND2_X1   g14064(.A1(new_n14122_), .A2(new_n14127_), .ZN(new_n14129_));
  OAI21_X1   g14065(.A1(new_n14115_), .A2(new_n14128_), .B(new_n14129_), .ZN(new_n14130_));
  OAI22_X1   g14066(.A1(new_n9478_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n10853_), .ZN(new_n14131_));
  NAND2_X1   g14067(.A1(new_n10862_), .A2(new_n3317_), .ZN(new_n14132_));
  AOI21_X1   g14068(.A1(new_n14131_), .A2(new_n14132_), .B(new_n3260_), .ZN(new_n14133_));
  NAND2_X1   g14069(.A1(new_n13484_), .A2(new_n14133_), .ZN(new_n14134_));
  XOR2_X1    g14070(.A1(new_n14134_), .A2(\a[26] ), .Z(new_n14135_));
  INV_X1     g14071(.I(new_n14135_), .ZN(new_n14136_));
  NAND2_X1   g14072(.A1(new_n13542_), .A2(new_n13528_), .ZN(new_n14137_));
  NAND2_X1   g14073(.A1(new_n14116_), .A2(new_n13540_), .ZN(new_n14138_));
  NAND2_X1   g14074(.A1(new_n13549_), .A2(new_n13554_), .ZN(new_n14139_));
  NAND2_X1   g14075(.A1(new_n13555_), .A2(new_n13557_), .ZN(new_n14140_));
  AOI22_X1   g14076(.A1(new_n14137_), .A2(new_n14138_), .B1(new_n14139_), .B2(new_n14140_), .ZN(new_n14141_));
  OAI21_X1   g14077(.A1(new_n13527_), .A2(new_n14117_), .B(new_n14138_), .ZN(new_n14142_));
  NOR2_X1    g14078(.A1(new_n13556_), .A2(new_n13558_), .ZN(new_n14143_));
  NOR2_X1    g14079(.A1(new_n14142_), .A2(new_n14143_), .ZN(new_n14144_));
  NOR2_X1    g14080(.A1(new_n14144_), .A2(new_n14141_), .ZN(new_n14145_));
  NOR2_X1    g14081(.A1(new_n14145_), .A2(new_n14136_), .ZN(new_n14146_));
  NAND2_X1   g14082(.A1(new_n14140_), .A2(new_n14139_), .ZN(new_n14147_));
  NAND2_X1   g14083(.A1(new_n14142_), .A2(new_n14147_), .ZN(new_n14148_));
  OAI21_X1   g14084(.A1(new_n14142_), .A2(new_n14143_), .B(new_n14148_), .ZN(new_n14149_));
  NOR2_X1    g14085(.A1(new_n14149_), .A2(new_n14135_), .ZN(new_n14150_));
  NOR3_X1    g14086(.A1(new_n14130_), .A2(new_n14150_), .A3(new_n14146_), .ZN(new_n14151_));
  INV_X1     g14087(.I(new_n14049_), .ZN(new_n14152_));
  INV_X1     g14088(.I(new_n14061_), .ZN(new_n14153_));
  OAI21_X1   g14089(.A1(new_n14059_), .A2(new_n14153_), .B(new_n14152_), .ZN(new_n14154_));
  NAND3_X1   g14090(.A1(new_n14078_), .A2(new_n14079_), .A3(new_n14070_), .ZN(new_n14155_));
  NAND2_X1   g14091(.A1(new_n14155_), .A2(new_n14154_), .ZN(new_n14156_));
  OAI21_X1   g14092(.A1(new_n14071_), .A2(new_n14072_), .B(new_n14066_), .ZN(new_n14157_));
  NAND2_X1   g14093(.A1(new_n14156_), .A2(new_n14157_), .ZN(new_n14158_));
  NAND3_X1   g14094(.A1(new_n14084_), .A2(new_n13515_), .A3(new_n13523_), .ZN(new_n14159_));
  OAI21_X1   g14095(.A1(new_n13516_), .A2(new_n13517_), .B(new_n14082_), .ZN(new_n14160_));
  NAND2_X1   g14096(.A1(new_n14160_), .A2(new_n14159_), .ZN(new_n14161_));
  INV_X1     g14097(.I(new_n14093_), .ZN(new_n14162_));
  NAND3_X1   g14098(.A1(new_n14162_), .A2(new_n14161_), .A3(new_n14091_), .ZN(new_n14163_));
  AOI21_X1   g14099(.A1(new_n14162_), .A2(new_n14091_), .B(new_n14161_), .ZN(new_n14164_));
  AOI21_X1   g14100(.A1(new_n14158_), .A2(new_n14163_), .B(new_n14164_), .ZN(new_n14165_));
  INV_X1     g14101(.I(new_n14109_), .ZN(new_n14166_));
  NAND2_X1   g14102(.A1(new_n14166_), .A2(new_n14110_), .ZN(new_n14167_));
  NOR2_X1    g14103(.A1(new_n14167_), .A2(new_n14103_), .ZN(new_n14168_));
  NAND2_X1   g14104(.A1(new_n14167_), .A2(new_n14103_), .ZN(new_n14169_));
  OAI21_X1   g14105(.A1(new_n14165_), .A2(new_n14168_), .B(new_n14169_), .ZN(new_n14170_));
  AOI21_X1   g14106(.A1(new_n13542_), .A2(new_n14138_), .B(new_n13527_), .ZN(new_n14171_));
  NAND2_X1   g14107(.A1(new_n14116_), .A2(new_n13541_), .ZN(new_n14172_));
  NAND2_X1   g14108(.A1(new_n13538_), .A2(new_n13540_), .ZN(new_n14173_));
  AOI21_X1   g14109(.A1(new_n14172_), .A2(new_n14173_), .B(new_n13528_), .ZN(new_n14174_));
  NOR2_X1    g14110(.A1(new_n14171_), .A2(new_n14174_), .ZN(new_n14175_));
  NOR2_X1    g14111(.A1(new_n14126_), .A2(\a[26] ), .ZN(new_n14176_));
  AOI21_X1   g14112(.A1(new_n13016_), .A2(new_n14125_), .B(new_n72_), .ZN(new_n14177_));
  NOR2_X1    g14113(.A1(new_n14176_), .A2(new_n14177_), .ZN(new_n14178_));
  NAND2_X1   g14114(.A1(new_n14175_), .A2(new_n14178_), .ZN(new_n14179_));
  NOR2_X1    g14115(.A1(new_n14175_), .A2(new_n14178_), .ZN(new_n14180_));
  AOI21_X1   g14116(.A1(new_n14170_), .A2(new_n14179_), .B(new_n14180_), .ZN(new_n14181_));
  NAND2_X1   g14117(.A1(new_n14149_), .A2(new_n14135_), .ZN(new_n14182_));
  NAND2_X1   g14118(.A1(new_n14145_), .A2(new_n14136_), .ZN(new_n14183_));
  AOI21_X1   g14119(.A1(new_n14182_), .A2(new_n14183_), .B(new_n14181_), .ZN(new_n14184_));
  NOR2_X1    g14120(.A1(new_n14184_), .A2(new_n14151_), .ZN(new_n14185_));
  NOR2_X1    g14121(.A1(new_n14185_), .A2(new_n14042_), .ZN(new_n14186_));
  AOI22_X1   g14122(.A1(new_n12823_), .A2(new_n5291_), .B1(new_n3782_), .B2(new_n10800_), .ZN(new_n14187_));
  NOR2_X1    g14123(.A1(new_n10798_), .A2(new_n3780_), .ZN(new_n14188_));
  OAI21_X1   g14124(.A1(new_n14187_), .A2(new_n14188_), .B(new_n3301_), .ZN(new_n14189_));
  NOR2_X1    g14125(.A1(new_n13504_), .A2(new_n14189_), .ZN(new_n14190_));
  NAND2_X1   g14126(.A1(new_n14190_), .A2(new_n84_), .ZN(new_n14191_));
  OAI21_X1   g14127(.A1(new_n13504_), .A2(new_n14189_), .B(\a[23] ), .ZN(new_n14192_));
  AOI21_X1   g14128(.A1(new_n14191_), .A2(new_n14192_), .B(new_n14058_), .ZN(new_n14193_));
  AOI22_X1   g14129(.A1(new_n10794_), .A2(new_n5291_), .B1(new_n3782_), .B2(new_n12823_), .ZN(new_n14194_));
  AOI21_X1   g14130(.A1(new_n3312_), .A2(new_n10800_), .B(new_n14194_), .ZN(new_n14195_));
  NAND2_X1   g14131(.A1(new_n12830_), .A2(new_n3301_), .ZN(new_n14196_));
  NOR2_X1    g14132(.A1(new_n14196_), .A2(new_n14195_), .ZN(new_n14197_));
  NOR2_X1    g14133(.A1(new_n14197_), .A2(\a[23] ), .ZN(new_n14198_));
  INV_X1     g14134(.I(new_n14198_), .ZN(new_n14199_));
  NAND2_X1   g14135(.A1(new_n14197_), .A2(\a[23] ), .ZN(new_n14200_));
  NOR2_X1    g14136(.A1(new_n3299_), .A2(new_n3300_), .ZN(new_n14201_));
  OAI21_X1   g14137(.A1(new_n12826_), .A2(new_n3306_), .B(new_n14201_), .ZN(new_n14202_));
  OR3_X2     g14138(.A1(new_n12847_), .A2(\a[23] ), .A3(new_n14202_), .Z(new_n14203_));
  OAI21_X1   g14139(.A1(new_n12847_), .A2(new_n14202_), .B(\a[23] ), .ZN(new_n14204_));
  NAND2_X1   g14140(.A1(new_n14203_), .A2(new_n14204_), .ZN(new_n14205_));
  NOR2_X1    g14141(.A1(new_n12826_), .A2(new_n3299_), .ZN(new_n14206_));
  NOR2_X1    g14142(.A1(new_n14206_), .A2(new_n84_), .ZN(new_n14207_));
  INV_X1     g14143(.I(new_n14207_), .ZN(new_n14208_));
  NOR2_X1    g14144(.A1(new_n14205_), .A2(new_n14208_), .ZN(new_n14209_));
  NAND3_X1   g14145(.A1(new_n14199_), .A2(new_n14200_), .A3(new_n14209_), .ZN(new_n14210_));
  NAND3_X1   g14146(.A1(new_n14191_), .A2(new_n14058_), .A3(new_n14192_), .ZN(new_n14211_));
  AOI21_X1   g14147(.A1(new_n14210_), .A2(new_n14211_), .B(new_n14193_), .ZN(new_n14212_));
  NOR2_X1    g14148(.A1(new_n14058_), .A2(new_n72_), .ZN(new_n14213_));
  XOR2_X1    g14149(.A1(new_n14057_), .A2(new_n14213_), .Z(new_n14214_));
  AOI22_X1   g14150(.A1(new_n9529_), .A2(new_n3782_), .B1(new_n10800_), .B2(new_n5291_), .ZN(new_n14215_));
  AOI21_X1   g14151(.A1(new_n10839_), .A2(new_n3312_), .B(new_n14215_), .ZN(new_n14216_));
  NOR2_X1    g14152(.A1(new_n14216_), .A2(new_n3302_), .ZN(new_n14217_));
  NAND2_X1   g14153(.A1(new_n12910_), .A2(new_n14217_), .ZN(new_n14218_));
  NOR2_X1    g14154(.A1(new_n14218_), .A2(\a[23] ), .ZN(new_n14219_));
  NAND2_X1   g14155(.A1(new_n14218_), .A2(\a[23] ), .ZN(new_n14220_));
  INV_X1     g14156(.I(new_n14220_), .ZN(new_n14221_));
  NOR3_X1    g14157(.A1(new_n14214_), .A2(new_n14219_), .A3(new_n14221_), .ZN(new_n14222_));
  OAI21_X1   g14158(.A1(new_n14221_), .A2(new_n14219_), .B(new_n14214_), .ZN(new_n14223_));
  OAI21_X1   g14159(.A1(new_n14212_), .A2(new_n14222_), .B(new_n14223_), .ZN(new_n14224_));
  NOR2_X1    g14160(.A1(new_n14053_), .A2(\a[26] ), .ZN(new_n14225_));
  INV_X1     g14161(.I(new_n14225_), .ZN(new_n14226_));
  NAND2_X1   g14162(.A1(new_n14053_), .A2(\a[26] ), .ZN(new_n14227_));
  NOR4_X1    g14163(.A1(new_n12847_), .A2(new_n72_), .A3(new_n14055_), .A4(new_n14058_), .ZN(new_n14228_));
  INV_X1     g14164(.I(new_n14228_), .ZN(new_n14229_));
  NAND3_X1   g14165(.A1(new_n14226_), .A2(new_n14227_), .A3(new_n14229_), .ZN(new_n14230_));
  INV_X1     g14166(.I(new_n14227_), .ZN(new_n14231_));
  OAI21_X1   g14167(.A1(new_n14231_), .A2(new_n14225_), .B(new_n14228_), .ZN(new_n14232_));
  NAND2_X1   g14168(.A1(new_n14232_), .A2(new_n14230_), .ZN(new_n14233_));
  AOI22_X1   g14169(.A1(new_n10839_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n9529_), .ZN(new_n14234_));
  NOR2_X1    g14170(.A1(new_n10846_), .A2(new_n3780_), .ZN(new_n14235_));
  OAI21_X1   g14171(.A1(new_n14234_), .A2(new_n14235_), .B(new_n3301_), .ZN(new_n14236_));
  OR3_X2     g14172(.A1(new_n12946_), .A2(\a[23] ), .A3(new_n14236_), .Z(new_n14237_));
  OAI21_X1   g14173(.A1(new_n12946_), .A2(new_n14236_), .B(\a[23] ), .ZN(new_n14238_));
  NAND2_X1   g14174(.A1(new_n14237_), .A2(new_n14238_), .ZN(new_n14239_));
  INV_X1     g14175(.I(new_n14239_), .ZN(new_n14240_));
  NAND2_X1   g14176(.A1(new_n14240_), .A2(new_n14233_), .ZN(new_n14241_));
  NOR3_X1    g14177(.A1(new_n14231_), .A2(new_n14225_), .A3(new_n14228_), .ZN(new_n14242_));
  AOI21_X1   g14178(.A1(new_n14226_), .A2(new_n14227_), .B(new_n14229_), .ZN(new_n14243_));
  NOR2_X1    g14179(.A1(new_n14243_), .A2(new_n14242_), .ZN(new_n14244_));
  NAND2_X1   g14180(.A1(new_n14244_), .A2(new_n14239_), .ZN(new_n14245_));
  INV_X1     g14181(.I(new_n14245_), .ZN(new_n14246_));
  AOI21_X1   g14182(.A1(new_n14224_), .A2(new_n14241_), .B(new_n14246_), .ZN(new_n14247_));
  NAND3_X1   g14183(.A1(new_n14047_), .A2(new_n13522_), .A3(new_n14048_), .ZN(new_n14248_));
  NAND2_X1   g14184(.A1(new_n14047_), .A2(new_n14048_), .ZN(new_n14249_));
  NAND2_X1   g14185(.A1(new_n14249_), .A2(new_n13521_), .ZN(new_n14250_));
  NAND2_X1   g14186(.A1(new_n14250_), .A2(new_n14248_), .ZN(new_n14251_));
  AOI21_X1   g14187(.A1(new_n14152_), .A2(new_n14061_), .B(new_n14059_), .ZN(new_n14252_));
  AOI21_X1   g14188(.A1(new_n14059_), .A2(new_n14251_), .B(new_n14252_), .ZN(new_n14253_));
  AOI22_X1   g14189(.A1(new_n10839_), .A2(new_n5291_), .B1(new_n12936_), .B2(new_n3782_), .ZN(new_n14254_));
  NOR2_X1    g14190(.A1(new_n9478_), .A2(new_n3780_), .ZN(new_n14255_));
  OAI21_X1   g14191(.A1(new_n14254_), .A2(new_n14255_), .B(new_n3301_), .ZN(new_n14256_));
  OR3_X2     g14192(.A1(new_n12975_), .A2(\a[23] ), .A3(new_n14256_), .Z(new_n14257_));
  OR2_X2     g14193(.A1(new_n12975_), .A2(new_n14256_), .Z(new_n14258_));
  NAND2_X1   g14194(.A1(new_n14258_), .A2(\a[23] ), .ZN(new_n14259_));
  NAND3_X1   g14195(.A1(new_n14253_), .A2(new_n14259_), .A3(new_n14257_), .ZN(new_n14260_));
  INV_X1     g14196(.I(new_n14260_), .ZN(new_n14261_));
  NAND2_X1   g14197(.A1(new_n14251_), .A2(new_n14059_), .ZN(new_n14262_));
  INV_X1     g14198(.I(new_n14252_), .ZN(new_n14263_));
  NAND2_X1   g14199(.A1(new_n14263_), .A2(new_n14262_), .ZN(new_n14264_));
  INV_X1     g14200(.I(new_n14257_), .ZN(new_n14265_));
  INV_X1     g14201(.I(new_n14259_), .ZN(new_n14266_));
  OAI21_X1   g14202(.A1(new_n14266_), .A2(new_n14265_), .B(new_n14264_), .ZN(new_n14267_));
  OAI21_X1   g14203(.A1(new_n14247_), .A2(new_n14261_), .B(new_n14267_), .ZN(new_n14268_));
  NAND3_X1   g14204(.A1(new_n14066_), .A2(new_n14079_), .A3(new_n14070_), .ZN(new_n14269_));
  OAI21_X1   g14205(.A1(new_n14071_), .A2(new_n14072_), .B(new_n14078_), .ZN(new_n14270_));
  AOI21_X1   g14206(.A1(new_n14269_), .A2(new_n14270_), .B(new_n14062_), .ZN(new_n14271_));
  INV_X1     g14207(.I(new_n14271_), .ZN(new_n14272_));
  OAI21_X1   g14208(.A1(new_n14073_), .A2(new_n14080_), .B(new_n14062_), .ZN(new_n14273_));
  NAND2_X1   g14209(.A1(new_n14272_), .A2(new_n14273_), .ZN(new_n14274_));
  OAI22_X1   g14210(.A1(new_n9478_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n10846_), .ZN(new_n14275_));
  NAND2_X1   g14211(.A1(new_n10854_), .A2(new_n3312_), .ZN(new_n14276_));
  AOI21_X1   g14212(.A1(new_n14275_), .A2(new_n14276_), .B(new_n3302_), .ZN(new_n14277_));
  NAND3_X1   g14213(.A1(new_n13016_), .A2(new_n84_), .A3(new_n14277_), .ZN(new_n14278_));
  INV_X1     g14214(.I(new_n14278_), .ZN(new_n14279_));
  AOI21_X1   g14215(.A1(new_n13016_), .A2(new_n14277_), .B(new_n84_), .ZN(new_n14280_));
  NOR2_X1    g14216(.A1(new_n14279_), .A2(new_n14280_), .ZN(new_n14281_));
  NAND2_X1   g14217(.A1(new_n14274_), .A2(new_n14281_), .ZN(new_n14282_));
  NOR2_X1    g14218(.A1(new_n14274_), .A2(new_n14281_), .ZN(new_n14283_));
  AOI21_X1   g14219(.A1(new_n14268_), .A2(new_n14282_), .B(new_n14283_), .ZN(new_n14284_));
  NAND3_X1   g14220(.A1(new_n14162_), .A2(new_n14086_), .A3(new_n14091_), .ZN(new_n14285_));
  INV_X1     g14221(.I(new_n14285_), .ZN(new_n14286_));
  AOI21_X1   g14222(.A1(new_n14162_), .A2(new_n14091_), .B(new_n14086_), .ZN(new_n14287_));
  OAI22_X1   g14223(.A1(new_n14286_), .A2(new_n14287_), .B1(new_n14074_), .B2(new_n14080_), .ZN(new_n14288_));
  NAND2_X1   g14224(.A1(new_n14095_), .A2(new_n14163_), .ZN(new_n14289_));
  NAND3_X1   g14225(.A1(new_n14289_), .A2(new_n14156_), .A3(new_n14157_), .ZN(new_n14290_));
  NAND2_X1   g14226(.A1(new_n14288_), .A2(new_n14290_), .ZN(new_n14291_));
  OAI22_X1   g14227(.A1(new_n9478_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n10853_), .ZN(new_n14292_));
  NAND2_X1   g14228(.A1(new_n10862_), .A2(new_n3312_), .ZN(new_n14293_));
  AOI21_X1   g14229(.A1(new_n14292_), .A2(new_n14293_), .B(new_n3302_), .ZN(new_n14294_));
  NAND3_X1   g14230(.A1(new_n13484_), .A2(new_n84_), .A3(new_n14294_), .ZN(new_n14295_));
  INV_X1     g14231(.I(new_n14295_), .ZN(new_n14296_));
  AOI21_X1   g14232(.A1(new_n13484_), .A2(new_n14294_), .B(new_n84_), .ZN(new_n14297_));
  NOR2_X1    g14233(.A1(new_n14296_), .A2(new_n14297_), .ZN(new_n14298_));
  NAND2_X1   g14234(.A1(new_n14291_), .A2(new_n14298_), .ZN(new_n14299_));
  INV_X1     g14235(.I(new_n14299_), .ZN(new_n14300_));
  INV_X1     g14236(.I(new_n14297_), .ZN(new_n14301_));
  NAND2_X1   g14237(.A1(new_n14301_), .A2(new_n14295_), .ZN(new_n14302_));
  NAND3_X1   g14238(.A1(new_n14302_), .A2(new_n14288_), .A3(new_n14290_), .ZN(new_n14303_));
  OAI21_X1   g14239(.A1(new_n14300_), .A2(new_n14284_), .B(new_n14303_), .ZN(new_n14304_));
  NAND2_X1   g14240(.A1(new_n14112_), .A2(new_n14103_), .ZN(new_n14305_));
  NAND2_X1   g14241(.A1(new_n14104_), .A2(new_n14167_), .ZN(new_n14306_));
  AOI21_X1   g14242(.A1(new_n14306_), .A2(new_n14305_), .B(new_n14165_), .ZN(new_n14307_));
  AOI21_X1   g14243(.A1(new_n14113_), .A2(new_n14169_), .B(new_n14096_), .ZN(new_n14308_));
  OAI22_X1   g14244(.A1(new_n10861_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n10853_), .ZN(new_n14309_));
  NAND2_X1   g14245(.A1(new_n8785_), .A2(new_n3312_), .ZN(new_n14310_));
  AOI21_X1   g14246(.A1(new_n14310_), .A2(new_n14309_), .B(new_n3302_), .ZN(new_n14311_));
  NAND2_X1   g14247(.A1(new_n13592_), .A2(new_n14311_), .ZN(new_n14312_));
  XOR2_X1    g14248(.A1(new_n14312_), .A2(\a[23] ), .Z(new_n14313_));
  OAI21_X1   g14249(.A1(new_n14307_), .A2(new_n14308_), .B(new_n14313_), .ZN(new_n14314_));
  NOR3_X1    g14250(.A1(new_n14313_), .A2(new_n14308_), .A3(new_n14307_), .ZN(new_n14315_));
  AOI21_X1   g14251(.A1(new_n14304_), .A2(new_n14314_), .B(new_n14315_), .ZN(new_n14316_));
  OAI21_X1   g14252(.A1(new_n14128_), .A2(new_n14180_), .B(new_n14170_), .ZN(new_n14317_));
  NOR2_X1    g14253(.A1(new_n14175_), .A2(new_n14127_), .ZN(new_n14318_));
  NOR2_X1    g14254(.A1(new_n14122_), .A2(new_n14178_), .ZN(new_n14319_));
  OAI21_X1   g14255(.A1(new_n14318_), .A2(new_n14319_), .B(new_n14115_), .ZN(new_n14320_));
  OAI22_X1   g14256(.A1(new_n8784_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n10861_), .ZN(new_n14321_));
  NAND2_X1   g14257(.A1(new_n8779_), .A2(new_n3312_), .ZN(new_n14322_));
  AOI21_X1   g14258(.A1(new_n14322_), .A2(new_n14321_), .B(new_n3302_), .ZN(new_n14323_));
  NAND3_X1   g14259(.A1(new_n12814_), .A2(new_n84_), .A3(new_n14323_), .ZN(new_n14324_));
  AOI21_X1   g14260(.A1(new_n12814_), .A2(new_n14323_), .B(new_n84_), .ZN(new_n14325_));
  INV_X1     g14261(.I(new_n14325_), .ZN(new_n14326_));
  NAND4_X1   g14262(.A1(new_n14320_), .A2(new_n14317_), .A3(new_n14324_), .A4(new_n14326_), .ZN(new_n14327_));
  AOI21_X1   g14263(.A1(new_n14129_), .A2(new_n14179_), .B(new_n14115_), .ZN(new_n14328_));
  NAND2_X1   g14264(.A1(new_n14122_), .A2(new_n14178_), .ZN(new_n14329_));
  NAND2_X1   g14265(.A1(new_n14175_), .A2(new_n14127_), .ZN(new_n14330_));
  AOI21_X1   g14266(.A1(new_n14330_), .A2(new_n14329_), .B(new_n14170_), .ZN(new_n14331_));
  INV_X1     g14267(.I(new_n14324_), .ZN(new_n14332_));
  OAI22_X1   g14268(.A1(new_n14328_), .A2(new_n14331_), .B1(new_n14332_), .B2(new_n14325_), .ZN(new_n14333_));
  NAND3_X1   g14269(.A1(new_n14316_), .A2(new_n14327_), .A3(new_n14333_), .ZN(new_n14334_));
  NAND3_X1   g14270(.A1(new_n14181_), .A2(new_n14182_), .A3(new_n14183_), .ZN(new_n14335_));
  OAI21_X1   g14271(.A1(new_n14146_), .A2(new_n14150_), .B(new_n14130_), .ZN(new_n14336_));
  NAND3_X1   g14272(.A1(new_n14336_), .A2(new_n14335_), .A3(new_n14042_), .ZN(new_n14337_));
  XOR2_X1    g14273(.A1(new_n14041_), .A2(\a[23] ), .Z(new_n14338_));
  OAI21_X1   g14274(.A1(new_n14184_), .A2(new_n14151_), .B(new_n14338_), .ZN(new_n14339_));
  INV_X1     g14275(.I(new_n14327_), .ZN(new_n14340_));
  AOI21_X1   g14276(.A1(new_n14337_), .A2(new_n14339_), .B(new_n14340_), .ZN(new_n14341_));
  AOI21_X1   g14277(.A1(new_n14341_), .A2(new_n14334_), .B(new_n14186_), .ZN(new_n14342_));
  OAI22_X1   g14278(.A1(new_n10871_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8778_), .ZN(new_n14343_));
  NAND2_X1   g14279(.A1(new_n10886_), .A2(new_n3312_), .ZN(new_n14344_));
  AOI21_X1   g14280(.A1(new_n14344_), .A2(new_n14343_), .B(new_n3302_), .ZN(new_n14345_));
  NAND2_X1   g14281(.A1(new_n13103_), .A2(new_n14345_), .ZN(new_n14346_));
  XOR2_X1    g14282(.A1(new_n14346_), .A2(new_n84_), .Z(new_n14347_));
  NAND2_X1   g14283(.A1(new_n13571_), .A2(new_n13580_), .ZN(new_n14348_));
  NAND2_X1   g14284(.A1(new_n13579_), .A2(new_n13576_), .ZN(new_n14349_));
  NAND2_X1   g14285(.A1(new_n14348_), .A2(new_n14349_), .ZN(new_n14350_));
  NAND2_X1   g14286(.A1(new_n14350_), .A2(new_n13560_), .ZN(new_n14351_));
  INV_X1     g14287(.I(new_n13556_), .ZN(new_n14352_));
  AOI21_X1   g14288(.A1(new_n14142_), .A2(new_n14352_), .B(new_n13558_), .ZN(new_n14353_));
  OAI21_X1   g14289(.A1(new_n13581_), .A2(new_n13577_), .B(new_n14353_), .ZN(new_n14354_));
  NAND2_X1   g14290(.A1(new_n14354_), .A2(new_n14351_), .ZN(new_n14355_));
  OAI22_X1   g14291(.A1(new_n10861_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n10853_), .ZN(new_n14356_));
  NAND2_X1   g14292(.A1(new_n8785_), .A2(new_n3317_), .ZN(new_n14357_));
  AOI21_X1   g14293(.A1(new_n14357_), .A2(new_n14356_), .B(new_n3260_), .ZN(new_n14358_));
  NAND2_X1   g14294(.A1(new_n13592_), .A2(new_n14358_), .ZN(new_n14359_));
  XOR2_X1    g14295(.A1(new_n14359_), .A2(\a[26] ), .Z(new_n14360_));
  NOR2_X1    g14296(.A1(new_n14355_), .A2(new_n14360_), .ZN(new_n14361_));
  NOR2_X1    g14297(.A1(new_n13577_), .A2(new_n13581_), .ZN(new_n14362_));
  NOR2_X1    g14298(.A1(new_n14362_), .A2(new_n13560_), .ZN(new_n14363_));
  AOI21_X1   g14299(.A1(new_n13560_), .A2(new_n14350_), .B(new_n14363_), .ZN(new_n14364_));
  INV_X1     g14300(.I(new_n14360_), .ZN(new_n14365_));
  NOR2_X1    g14301(.A1(new_n14364_), .A2(new_n14365_), .ZN(new_n14366_));
  OAI21_X1   g14302(.A1(new_n14130_), .A2(new_n14150_), .B(new_n14182_), .ZN(new_n14367_));
  NOR3_X1    g14303(.A1(new_n14366_), .A2(new_n14367_), .A3(new_n14361_), .ZN(new_n14368_));
  NAND2_X1   g14304(.A1(new_n14364_), .A2(new_n14365_), .ZN(new_n14369_));
  NAND2_X1   g14305(.A1(new_n14355_), .A2(new_n14360_), .ZN(new_n14370_));
  AOI21_X1   g14306(.A1(new_n14181_), .A2(new_n14183_), .B(new_n14146_), .ZN(new_n14371_));
  AOI21_X1   g14307(.A1(new_n14369_), .A2(new_n14370_), .B(new_n14371_), .ZN(new_n14372_));
  NOR3_X1    g14308(.A1(new_n14347_), .A2(new_n14372_), .A3(new_n14368_), .ZN(new_n14373_));
  OAI21_X1   g14309(.A1(new_n14372_), .A2(new_n14368_), .B(new_n14347_), .ZN(new_n14374_));
  OAI21_X1   g14310(.A1(new_n14342_), .A2(new_n14373_), .B(new_n14374_), .ZN(new_n14375_));
  INV_X1     g14311(.I(new_n13500_), .ZN(new_n14376_));
  NAND2_X1   g14312(.A1(new_n14376_), .A2(new_n13583_), .ZN(new_n14377_));
  XOR2_X1    g14313(.A1(new_n14377_), .A2(new_n13582_), .Z(new_n14378_));
  NAND2_X1   g14314(.A1(new_n14369_), .A2(new_n14370_), .ZN(new_n14379_));
  OAI22_X1   g14315(.A1(new_n8784_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n10861_), .ZN(new_n14380_));
  NAND2_X1   g14316(.A1(new_n8779_), .A2(new_n3317_), .ZN(new_n14381_));
  AOI21_X1   g14317(.A1(new_n14381_), .A2(new_n14380_), .B(new_n3260_), .ZN(new_n14382_));
  NAND2_X1   g14318(.A1(new_n12814_), .A2(new_n14382_), .ZN(new_n14383_));
  XOR2_X1    g14319(.A1(new_n14383_), .A2(\a[26] ), .Z(new_n14384_));
  OAI21_X1   g14320(.A1(new_n14379_), .A2(new_n14371_), .B(new_n14384_), .ZN(new_n14385_));
  INV_X1     g14321(.I(new_n14385_), .ZN(new_n14386_));
  NOR3_X1    g14322(.A1(new_n14379_), .A2(new_n14371_), .A3(new_n14384_), .ZN(new_n14387_));
  OAI21_X1   g14323(.A1(new_n14386_), .A2(new_n14387_), .B(new_n14378_), .ZN(new_n14388_));
  INV_X1     g14324(.I(new_n14378_), .ZN(new_n14389_));
  INV_X1     g14325(.I(new_n14387_), .ZN(new_n14390_));
  NAND3_X1   g14326(.A1(new_n14390_), .A2(new_n14389_), .A3(new_n14385_), .ZN(new_n14391_));
  AOI22_X1   g14327(.A1(new_n10886_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n10872_), .ZN(new_n14392_));
  NOR2_X1    g14328(.A1(new_n10892_), .A2(new_n3780_), .ZN(new_n14393_));
  OAI21_X1   g14329(.A1(new_n14392_), .A2(new_n14393_), .B(new_n3301_), .ZN(new_n14394_));
  NOR2_X1    g14330(.A1(new_n12776_), .A2(new_n14394_), .ZN(new_n14395_));
  XOR2_X1    g14331(.A1(new_n14395_), .A2(new_n84_), .Z(new_n14396_));
  NAND3_X1   g14332(.A1(new_n14388_), .A2(new_n14391_), .A3(new_n14396_), .ZN(new_n14397_));
  NAND2_X1   g14333(.A1(new_n14397_), .A2(new_n14375_), .ZN(new_n14398_));
  AOI21_X1   g14334(.A1(new_n14390_), .A2(new_n14385_), .B(new_n14389_), .ZN(new_n14399_));
  INV_X1     g14335(.I(new_n14391_), .ZN(new_n14400_));
  INV_X1     g14336(.I(new_n14396_), .ZN(new_n14401_));
  OAI21_X1   g14337(.A1(new_n14400_), .A2(new_n14399_), .B(new_n14401_), .ZN(new_n14402_));
  NAND2_X1   g14338(.A1(new_n14398_), .A2(new_n14402_), .ZN(new_n14403_));
  NAND3_X1   g14339(.A1(new_n14010_), .A2(new_n14013_), .A3(new_n14018_), .ZN(new_n14404_));
  AOI21_X1   g14340(.A1(new_n14012_), .A2(new_n14008_), .B(new_n14011_), .ZN(new_n14405_));
  INV_X1     g14341(.I(new_n14013_), .ZN(new_n14406_));
  OAI21_X1   g14342(.A1(new_n14406_), .A2(new_n14405_), .B(new_n14019_), .ZN(new_n14407_));
  AOI22_X1   g14343(.A1(new_n10886_), .A2(new_n5291_), .B1(new_n10889_), .B2(new_n3782_), .ZN(new_n14408_));
  NOR2_X1    g14344(.A1(new_n10899_), .A2(new_n3780_), .ZN(new_n14409_));
  OAI21_X1   g14345(.A1(new_n14409_), .A2(new_n14408_), .B(new_n3301_), .ZN(new_n14410_));
  NOR2_X1    g14346(.A1(new_n11908_), .A2(new_n14410_), .ZN(new_n14411_));
  XOR2_X1    g14347(.A1(new_n14411_), .A2(new_n84_), .Z(new_n14412_));
  NAND3_X1   g14348(.A1(new_n14412_), .A2(new_n14404_), .A3(new_n14407_), .ZN(new_n14413_));
  AOI21_X1   g14349(.A1(new_n14404_), .A2(new_n14407_), .B(new_n14412_), .ZN(new_n14414_));
  AOI21_X1   g14350(.A1(new_n14403_), .A2(new_n14413_), .B(new_n14414_), .ZN(new_n14415_));
  INV_X1     g14351(.I(new_n14024_), .ZN(new_n14416_));
  AOI21_X1   g14352(.A1(new_n14005_), .A2(new_n14023_), .B(new_n14020_), .ZN(new_n14417_));
  AOI22_X1   g14353(.A1(new_n11899_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n10889_), .ZN(new_n14418_));
  NOR2_X1    g14354(.A1(new_n8774_), .A2(new_n3780_), .ZN(new_n14419_));
  OAI21_X1   g14355(.A1(new_n14419_), .A2(new_n14418_), .B(new_n3301_), .ZN(new_n14420_));
  NOR2_X1    g14356(.A1(new_n11945_), .A2(new_n14420_), .ZN(new_n14421_));
  NAND2_X1   g14357(.A1(new_n14421_), .A2(new_n84_), .ZN(new_n14422_));
  INV_X1     g14358(.I(new_n14422_), .ZN(new_n14423_));
  NOR2_X1    g14359(.A1(new_n14421_), .A2(new_n84_), .ZN(new_n14424_));
  NOR4_X1    g14360(.A1(new_n14416_), .A2(new_n14417_), .A3(new_n14423_), .A4(new_n14424_), .ZN(new_n14425_));
  AOI21_X1   g14361(.A1(new_n14021_), .A2(new_n13998_), .B(new_n14022_), .ZN(new_n14426_));
  INV_X1     g14362(.I(new_n14020_), .ZN(new_n14427_));
  NOR3_X1    g14363(.A1(new_n13999_), .A2(new_n13995_), .A3(new_n14004_), .ZN(new_n14428_));
  OAI21_X1   g14364(.A1(new_n14426_), .A2(new_n14428_), .B(new_n14427_), .ZN(new_n14429_));
  INV_X1     g14365(.I(new_n14424_), .ZN(new_n14430_));
  AOI22_X1   g14366(.A1(new_n14429_), .A2(new_n14024_), .B1(new_n14430_), .B2(new_n14422_), .ZN(new_n14431_));
  NOR2_X1    g14367(.A1(new_n14425_), .A2(new_n14431_), .ZN(new_n14432_));
  NAND2_X1   g14368(.A1(new_n14415_), .A2(new_n14432_), .ZN(new_n14433_));
  INV_X1     g14369(.I(new_n13988_), .ZN(new_n14434_));
  NAND3_X1   g14370(.A1(new_n14037_), .A2(new_n14034_), .A3(new_n14434_), .ZN(new_n14435_));
  AOI21_X1   g14371(.A1(new_n14036_), .A2(new_n14032_), .B(new_n14035_), .ZN(new_n14436_));
  NOR3_X1    g14372(.A1(new_n14033_), .A2(new_n13993_), .A3(new_n14031_), .ZN(new_n14437_));
  OAI21_X1   g14373(.A1(new_n14436_), .A2(new_n14437_), .B(new_n13988_), .ZN(new_n14438_));
  AOI21_X1   g14374(.A1(new_n14438_), .A2(new_n14435_), .B(new_n14425_), .ZN(new_n14439_));
  AOI22_X1   g14375(.A1(new_n14439_), .A2(new_n14433_), .B1(new_n13988_), .B2(new_n14038_), .ZN(new_n14440_));
  INV_X1     g14376(.I(new_n13828_), .ZN(new_n14441_));
  NOR2_X1    g14377(.A1(new_n13823_), .A2(new_n14441_), .ZN(new_n14442_));
  NOR2_X1    g14378(.A1(new_n13822_), .A2(new_n13828_), .ZN(new_n14443_));
  AOI22_X1   g14379(.A1(new_n5291_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n3782_), .ZN(new_n14444_));
  NOR2_X1    g14380(.A1(new_n8758_), .A2(new_n3780_), .ZN(new_n14445_));
  OAI21_X1   g14381(.A1(new_n14444_), .A2(new_n14445_), .B(new_n3301_), .ZN(new_n14446_));
  NOR2_X1    g14382(.A1(new_n12053_), .A2(new_n14446_), .ZN(new_n14447_));
  XOR2_X1    g14383(.A1(new_n14447_), .A2(new_n84_), .Z(new_n14448_));
  INV_X1     g14384(.I(new_n14448_), .ZN(new_n14449_));
  NOR3_X1    g14385(.A1(new_n14442_), .A2(new_n14443_), .A3(new_n14449_), .ZN(new_n14450_));
  NOR2_X1    g14386(.A1(new_n14442_), .A2(new_n14443_), .ZN(new_n14451_));
  NOR2_X1    g14387(.A1(new_n14451_), .A2(new_n14448_), .ZN(new_n14452_));
  NOR2_X1    g14388(.A1(new_n14452_), .A2(new_n14450_), .ZN(new_n14453_));
  INV_X1     g14389(.I(new_n14453_), .ZN(new_n14454_));
  NAND2_X1   g14390(.A1(new_n14440_), .A2(new_n14454_), .ZN(new_n14455_));
  NAND2_X1   g14391(.A1(new_n14038_), .A2(new_n13988_), .ZN(new_n14456_));
  AOI21_X1   g14392(.A1(new_n14388_), .A2(new_n14391_), .B(new_n14396_), .ZN(new_n14457_));
  AOI21_X1   g14393(.A1(new_n14375_), .A2(new_n14397_), .B(new_n14457_), .ZN(new_n14458_));
  NAND2_X1   g14394(.A1(new_n14407_), .A2(new_n14404_), .ZN(new_n14459_));
  XOR2_X1    g14395(.A1(new_n14411_), .A2(\a[23] ), .Z(new_n14460_));
  NOR2_X1    g14396(.A1(new_n14460_), .A2(new_n14459_), .ZN(new_n14461_));
  NAND2_X1   g14397(.A1(new_n14460_), .A2(new_n14459_), .ZN(new_n14462_));
  OAI21_X1   g14398(.A1(new_n14458_), .A2(new_n14461_), .B(new_n14462_), .ZN(new_n14463_));
  NAND4_X1   g14399(.A1(new_n14429_), .A2(new_n14430_), .A3(new_n14024_), .A4(new_n14422_), .ZN(new_n14464_));
  OAI22_X1   g14400(.A1(new_n14416_), .A2(new_n14417_), .B1(new_n14423_), .B2(new_n14424_), .ZN(new_n14465_));
  NAND2_X1   g14401(.A1(new_n14465_), .A2(new_n14464_), .ZN(new_n14466_));
  NOR2_X1    g14402(.A1(new_n14463_), .A2(new_n14466_), .ZN(new_n14467_));
  NOR3_X1    g14403(.A1(new_n14436_), .A2(new_n14437_), .A3(new_n13988_), .ZN(new_n14468_));
  AOI21_X1   g14404(.A1(new_n14037_), .A2(new_n14034_), .B(new_n14434_), .ZN(new_n14469_));
  OAI21_X1   g14405(.A1(new_n14469_), .A2(new_n14468_), .B(new_n14464_), .ZN(new_n14470_));
  OAI21_X1   g14406(.A1(new_n14470_), .A2(new_n14467_), .B(new_n14456_), .ZN(new_n14471_));
  NAND2_X1   g14407(.A1(new_n14471_), .A2(new_n14453_), .ZN(new_n14472_));
  AOI21_X1   g14408(.A1(new_n14455_), .A2(new_n14472_), .B(new_n13983_), .ZN(new_n14473_));
  INV_X1     g14409(.I(new_n13983_), .ZN(new_n14474_));
  NOR2_X1    g14410(.A1(new_n14471_), .A2(new_n14453_), .ZN(new_n14475_));
  NOR2_X1    g14411(.A1(new_n14440_), .A2(new_n14454_), .ZN(new_n14476_));
  NOR3_X1    g14412(.A1(new_n14476_), .A2(new_n14475_), .A3(new_n14474_), .ZN(new_n14477_));
  OAI22_X1   g14413(.A1(new_n8725_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8735_), .ZN(new_n14478_));
  NAND2_X1   g14414(.A1(new_n8719_), .A2(new_n4469_), .ZN(new_n14479_));
  AOI21_X1   g14415(.A1(new_n14478_), .A2(new_n14479_), .B(new_n4468_), .ZN(new_n14480_));
  NAND2_X1   g14416(.A1(new_n12242_), .A2(new_n14480_), .ZN(new_n14481_));
  XOR2_X1    g14417(.A1(new_n14481_), .A2(new_n3372_), .Z(new_n14482_));
  OR3_X2     g14418(.A1(new_n14482_), .A2(new_n14477_), .A3(new_n14473_), .Z(new_n14483_));
  OAI21_X1   g14419(.A1(new_n14473_), .A2(new_n14477_), .B(new_n14482_), .ZN(new_n14484_));
  NAND2_X1   g14420(.A1(new_n14483_), .A2(new_n14484_), .ZN(new_n14485_));
  OAI22_X1   g14421(.A1(new_n8735_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n10924_), .ZN(new_n14486_));
  NAND2_X1   g14422(.A1(new_n8726_), .A2(new_n4469_), .ZN(new_n14487_));
  AOI21_X1   g14423(.A1(new_n14487_), .A2(new_n14486_), .B(new_n4468_), .ZN(new_n14488_));
  NAND2_X1   g14424(.A1(new_n12181_), .A2(new_n14488_), .ZN(new_n14489_));
  XOR2_X1    g14425(.A1(new_n14489_), .A2(new_n3372_), .Z(new_n14490_));
  INV_X1     g14426(.I(new_n14490_), .ZN(new_n14491_));
  OAI21_X1   g14427(.A1(new_n14467_), .A2(new_n14425_), .B(new_n13988_), .ZN(new_n14492_));
  NAND3_X1   g14428(.A1(new_n14433_), .A2(new_n14434_), .A3(new_n14464_), .ZN(new_n14493_));
  AOI21_X1   g14429(.A1(new_n14493_), .A2(new_n14492_), .B(new_n14038_), .ZN(new_n14494_));
  INV_X1     g14430(.I(new_n14038_), .ZN(new_n14495_));
  AOI21_X1   g14431(.A1(new_n14433_), .A2(new_n14464_), .B(new_n14434_), .ZN(new_n14496_));
  NOR3_X1    g14432(.A1(new_n14467_), .A2(new_n13988_), .A3(new_n14425_), .ZN(new_n14497_));
  NOR3_X1    g14433(.A1(new_n14496_), .A2(new_n14495_), .A3(new_n14497_), .ZN(new_n14498_));
  NOR2_X1    g14434(.A1(new_n14498_), .A2(new_n14494_), .ZN(new_n14499_));
  AOI22_X1   g14435(.A1(new_n8761_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n11996_), .ZN(new_n14500_));
  INV_X1     g14436(.I(new_n14500_), .ZN(new_n14501_));
  NAND2_X1   g14437(.A1(new_n8746_), .A2(new_n4096_), .ZN(new_n14502_));
  AOI21_X1   g14438(.A1(new_n14502_), .A2(new_n14501_), .B(new_n4095_), .ZN(new_n14503_));
  NAND3_X1   g14439(.A1(new_n11964_), .A2(new_n3035_), .A3(new_n14503_), .ZN(new_n14504_));
  NAND2_X1   g14440(.A1(new_n11964_), .A2(new_n14503_), .ZN(new_n14505_));
  NAND2_X1   g14441(.A1(new_n14505_), .A2(\a[20] ), .ZN(new_n14506_));
  NAND4_X1   g14442(.A1(new_n14465_), .A2(new_n14464_), .A3(new_n14506_), .A4(new_n14504_), .ZN(new_n14507_));
  AOI22_X1   g14443(.A1(new_n14465_), .A2(new_n14464_), .B1(new_n14506_), .B2(new_n14504_), .ZN(new_n14508_));
  INV_X1     g14444(.I(new_n14508_), .ZN(new_n14509_));
  AOI21_X1   g14445(.A1(new_n14509_), .A2(new_n14507_), .B(new_n14415_), .ZN(new_n14510_));
  XOR2_X1    g14446(.A1(new_n14505_), .A2(\a[20] ), .Z(new_n14511_));
  NAND2_X1   g14447(.A1(new_n14511_), .A2(new_n14466_), .ZN(new_n14512_));
  NAND2_X1   g14448(.A1(new_n14506_), .A2(new_n14504_), .ZN(new_n14513_));
  NAND2_X1   g14449(.A1(new_n14432_), .A2(new_n14513_), .ZN(new_n14514_));
  AOI21_X1   g14450(.A1(new_n14512_), .A2(new_n14514_), .B(new_n14463_), .ZN(new_n14515_));
  NOR2_X1    g14451(.A1(new_n14510_), .A2(new_n14515_), .ZN(new_n14516_));
  AOI22_X1   g14452(.A1(new_n3770_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n3776_), .ZN(new_n14517_));
  NOR2_X1    g14453(.A1(new_n8758_), .A2(new_n4097_), .ZN(new_n14518_));
  OAI21_X1   g14454(.A1(new_n14517_), .A2(new_n14518_), .B(new_n3773_), .ZN(new_n14519_));
  NOR2_X1    g14455(.A1(new_n12053_), .A2(new_n14519_), .ZN(new_n14520_));
  XOR2_X1    g14456(.A1(new_n14520_), .A2(new_n3035_), .Z(new_n14521_));
  XOR2_X1    g14457(.A1(new_n14412_), .A2(new_n14459_), .Z(new_n14522_));
  NAND2_X1   g14458(.A1(new_n14413_), .A2(new_n14462_), .ZN(new_n14523_));
  NAND2_X1   g14459(.A1(new_n14458_), .A2(new_n14523_), .ZN(new_n14524_));
  OAI21_X1   g14460(.A1(new_n14458_), .A2(new_n14522_), .B(new_n14524_), .ZN(new_n14525_));
  NOR2_X1    g14461(.A1(new_n14525_), .A2(new_n14521_), .ZN(new_n14526_));
  NAND2_X1   g14462(.A1(new_n14463_), .A2(new_n14432_), .ZN(new_n14527_));
  NAND2_X1   g14463(.A1(new_n14415_), .A2(new_n14466_), .ZN(new_n14528_));
  AOI21_X1   g14464(.A1(new_n14528_), .A2(new_n14527_), .B(new_n14513_), .ZN(new_n14529_));
  NOR2_X1    g14465(.A1(new_n14529_), .A2(new_n14526_), .ZN(new_n14530_));
  OAI22_X1   g14466(.A1(new_n8745_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n8758_), .ZN(new_n14531_));
  NAND2_X1   g14467(.A1(new_n8752_), .A2(new_n4096_), .ZN(new_n14532_));
  AOI21_X1   g14468(.A1(new_n14532_), .A2(new_n14531_), .B(new_n4095_), .ZN(new_n14533_));
  NAND2_X1   g14469(.A1(new_n12189_), .A2(new_n14533_), .ZN(new_n14534_));
  XOR2_X1    g14470(.A1(new_n14534_), .A2(\a[20] ), .Z(new_n14535_));
  INV_X1     g14471(.I(new_n14535_), .ZN(new_n14536_));
  AOI21_X1   g14472(.A1(new_n14530_), .A2(new_n14516_), .B(new_n14536_), .ZN(new_n14537_));
  NOR2_X1    g14473(.A1(new_n14466_), .A2(new_n14513_), .ZN(new_n14538_));
  OAI21_X1   g14474(.A1(new_n14538_), .A2(new_n14508_), .B(new_n14463_), .ZN(new_n14539_));
  NOR2_X1    g14475(.A1(new_n14432_), .A2(new_n14513_), .ZN(new_n14540_));
  NOR2_X1    g14476(.A1(new_n14511_), .A2(new_n14466_), .ZN(new_n14541_));
  OAI21_X1   g14477(.A1(new_n14541_), .A2(new_n14540_), .B(new_n14415_), .ZN(new_n14542_));
  NAND2_X1   g14478(.A1(new_n14542_), .A2(new_n14539_), .ZN(new_n14543_));
  INV_X1     g14479(.I(new_n14521_), .ZN(new_n14544_));
  NOR2_X1    g14480(.A1(new_n14522_), .A2(new_n14458_), .ZN(new_n14545_));
  NOR2_X1    g14481(.A1(new_n14414_), .A2(new_n14461_), .ZN(new_n14546_));
  NOR2_X1    g14482(.A1(new_n14403_), .A2(new_n14546_), .ZN(new_n14547_));
  NOR2_X1    g14483(.A1(new_n14547_), .A2(new_n14545_), .ZN(new_n14548_));
  NAND2_X1   g14484(.A1(new_n14548_), .A2(new_n14544_), .ZN(new_n14549_));
  NOR2_X1    g14485(.A1(new_n14415_), .A2(new_n14466_), .ZN(new_n14550_));
  NOR2_X1    g14486(.A1(new_n14463_), .A2(new_n14432_), .ZN(new_n14551_));
  OAI21_X1   g14487(.A1(new_n14550_), .A2(new_n14551_), .B(new_n14511_), .ZN(new_n14552_));
  NAND2_X1   g14488(.A1(new_n14552_), .A2(new_n14549_), .ZN(new_n14553_));
  NOR3_X1    g14489(.A1(new_n14553_), .A2(new_n14543_), .A3(new_n14535_), .ZN(new_n14554_));
  OAI21_X1   g14490(.A1(new_n14537_), .A2(new_n14554_), .B(new_n14499_), .ZN(new_n14555_));
  OAI21_X1   g14491(.A1(new_n14496_), .A2(new_n14497_), .B(new_n14495_), .ZN(new_n14556_));
  NAND3_X1   g14492(.A1(new_n14493_), .A2(new_n14038_), .A3(new_n14492_), .ZN(new_n14557_));
  NAND2_X1   g14493(.A1(new_n14556_), .A2(new_n14557_), .ZN(new_n14558_));
  OAI21_X1   g14494(.A1(new_n14553_), .A2(new_n14543_), .B(new_n14535_), .ZN(new_n14559_));
  NAND3_X1   g14495(.A1(new_n14530_), .A2(new_n14516_), .A3(new_n14536_), .ZN(new_n14560_));
  NAND3_X1   g14496(.A1(new_n14558_), .A2(new_n14559_), .A3(new_n14560_), .ZN(new_n14561_));
  NAND2_X1   g14497(.A1(new_n14555_), .A2(new_n14561_), .ZN(new_n14562_));
  NAND2_X1   g14498(.A1(new_n14562_), .A2(new_n14491_), .ZN(new_n14563_));
  NAND3_X1   g14499(.A1(new_n14555_), .A2(new_n14561_), .A3(new_n14490_), .ZN(new_n14564_));
  AOI21_X1   g14500(.A1(new_n14559_), .A2(new_n14560_), .B(new_n14558_), .ZN(new_n14565_));
  NOR3_X1    g14501(.A1(new_n14499_), .A2(new_n14537_), .A3(new_n14554_), .ZN(new_n14566_));
  OAI21_X1   g14502(.A1(new_n14565_), .A2(new_n14566_), .B(new_n14491_), .ZN(new_n14567_));
  NAND2_X1   g14503(.A1(new_n14567_), .A2(new_n14564_), .ZN(new_n14568_));
  NAND3_X1   g14504(.A1(new_n14526_), .A2(new_n14542_), .A3(new_n14539_), .ZN(new_n14569_));
  NAND2_X1   g14505(.A1(new_n14543_), .A2(new_n14549_), .ZN(new_n14570_));
  OAI22_X1   g14506(.A1(new_n8751_), .A2(new_n4291_), .B1(new_n4297_), .B2(new_n10924_), .ZN(new_n14571_));
  NAND2_X1   g14507(.A1(new_n8736_), .A2(new_n4469_), .ZN(new_n14572_));
  AOI21_X1   g14508(.A1(new_n14572_), .A2(new_n14571_), .B(new_n4468_), .ZN(new_n14573_));
  NAND2_X1   g14509(.A1(new_n12118_), .A2(new_n14573_), .ZN(new_n14574_));
  XOR2_X1    g14510(.A1(new_n14574_), .A2(\a[17] ), .Z(new_n14575_));
  NAND3_X1   g14511(.A1(new_n14570_), .A2(new_n14569_), .A3(new_n14575_), .ZN(new_n14576_));
  NOR2_X1    g14512(.A1(new_n14543_), .A2(new_n14549_), .ZN(new_n14577_));
  NOR2_X1    g14513(.A1(new_n14516_), .A2(new_n14526_), .ZN(new_n14578_));
  XOR2_X1    g14514(.A1(new_n14574_), .A2(new_n3372_), .Z(new_n14579_));
  OAI21_X1   g14515(.A1(new_n14578_), .A2(new_n14577_), .B(new_n14579_), .ZN(new_n14580_));
  NAND2_X1   g14516(.A1(new_n14580_), .A2(new_n14576_), .ZN(new_n14581_));
  NAND2_X1   g14517(.A1(new_n14525_), .A2(new_n14521_), .ZN(new_n14582_));
  INV_X1     g14518(.I(new_n14582_), .ZN(new_n14583_));
  NOR2_X1    g14519(.A1(new_n14525_), .A2(new_n14521_), .ZN(new_n14584_));
  OAI22_X1   g14520(.A1(new_n8751_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8745_), .ZN(new_n14585_));
  NAND2_X1   g14521(.A1(new_n10927_), .A2(new_n4469_), .ZN(new_n14586_));
  AOI21_X1   g14522(.A1(new_n14585_), .A2(new_n14586_), .B(new_n4468_), .ZN(new_n14587_));
  NAND2_X1   g14523(.A1(new_n12072_), .A2(new_n14587_), .ZN(new_n14588_));
  XOR2_X1    g14524(.A1(new_n14588_), .A2(\a[17] ), .Z(new_n14589_));
  OAI21_X1   g14525(.A1(new_n14583_), .A2(new_n14584_), .B(new_n14589_), .ZN(new_n14590_));
  INV_X1     g14526(.I(new_n14590_), .ZN(new_n14591_));
  NAND2_X1   g14527(.A1(new_n14548_), .A2(new_n14544_), .ZN(new_n14592_));
  XOR2_X1    g14528(.A1(new_n14588_), .A2(new_n3372_), .Z(new_n14593_));
  NAND3_X1   g14529(.A1(new_n14593_), .A2(new_n14582_), .A3(new_n14592_), .ZN(new_n14594_));
  OAI22_X1   g14530(.A1(new_n8745_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8758_), .ZN(new_n14595_));
  NAND2_X1   g14531(.A1(new_n8752_), .A2(new_n4469_), .ZN(new_n14596_));
  AOI21_X1   g14532(.A1(new_n14596_), .A2(new_n14595_), .B(new_n4468_), .ZN(new_n14597_));
  NAND2_X1   g14533(.A1(new_n12189_), .A2(new_n14597_), .ZN(new_n14598_));
  XOR2_X1    g14534(.A1(new_n14598_), .A2(\a[17] ), .Z(new_n14599_));
  INV_X1     g14535(.I(new_n14193_), .ZN(new_n14600_));
  INV_X1     g14536(.I(new_n14200_), .ZN(new_n14601_));
  INV_X1     g14537(.I(new_n14209_), .ZN(new_n14602_));
  NOR3_X1    g14538(.A1(new_n14602_), .A2(new_n14601_), .A3(new_n14198_), .ZN(new_n14603_));
  INV_X1     g14539(.I(new_n14211_), .ZN(new_n14604_));
  OAI21_X1   g14540(.A1(new_n14603_), .A2(new_n14604_), .B(new_n14600_), .ZN(new_n14605_));
  XOR2_X1    g14541(.A1(new_n14056_), .A2(new_n72_), .Z(new_n14606_));
  INV_X1     g14542(.I(new_n14213_), .ZN(new_n14607_));
  NAND2_X1   g14543(.A1(new_n14606_), .A2(new_n14607_), .ZN(new_n14608_));
  NAND2_X1   g14544(.A1(new_n14057_), .A2(new_n14213_), .ZN(new_n14609_));
  NAND2_X1   g14545(.A1(new_n14608_), .A2(new_n14609_), .ZN(new_n14610_));
  INV_X1     g14546(.I(new_n14219_), .ZN(new_n14611_));
  NAND3_X1   g14547(.A1(new_n14610_), .A2(new_n14611_), .A3(new_n14220_), .ZN(new_n14612_));
  AOI21_X1   g14548(.A1(new_n14611_), .A2(new_n14220_), .B(new_n14610_), .ZN(new_n14613_));
  AOI21_X1   g14549(.A1(new_n14605_), .A2(new_n14612_), .B(new_n14613_), .ZN(new_n14614_));
  NOR2_X1    g14550(.A1(new_n14244_), .A2(new_n14239_), .ZN(new_n14615_));
  OAI21_X1   g14551(.A1(new_n14614_), .A2(new_n14615_), .B(new_n14245_), .ZN(new_n14616_));
  AOI21_X1   g14552(.A1(new_n14257_), .A2(new_n14259_), .B(new_n14253_), .ZN(new_n14617_));
  AOI21_X1   g14553(.A1(new_n14616_), .A2(new_n14260_), .B(new_n14617_), .ZN(new_n14618_));
  AOI21_X1   g14554(.A1(new_n14157_), .A2(new_n14155_), .B(new_n14154_), .ZN(new_n14619_));
  NOR2_X1    g14555(.A1(new_n14619_), .A2(new_n14271_), .ZN(new_n14620_));
  INV_X1     g14556(.I(new_n14280_), .ZN(new_n14621_));
  NAND2_X1   g14557(.A1(new_n14621_), .A2(new_n14278_), .ZN(new_n14622_));
  NOR2_X1    g14558(.A1(new_n14622_), .A2(new_n14620_), .ZN(new_n14623_));
  NAND2_X1   g14559(.A1(new_n14622_), .A2(new_n14620_), .ZN(new_n14624_));
  OAI21_X1   g14560(.A1(new_n14618_), .A2(new_n14623_), .B(new_n14624_), .ZN(new_n14625_));
  INV_X1     g14561(.I(new_n14303_), .ZN(new_n14626_));
  AOI21_X1   g14562(.A1(new_n14625_), .A2(new_n14299_), .B(new_n14626_), .ZN(new_n14627_));
  NOR2_X1    g14563(.A1(new_n14308_), .A2(new_n14307_), .ZN(new_n14628_));
  XOR2_X1    g14564(.A1(new_n14312_), .A2(new_n84_), .Z(new_n14629_));
  NOR2_X1    g14565(.A1(new_n14628_), .A2(new_n14629_), .ZN(new_n14630_));
  NAND2_X1   g14566(.A1(new_n14628_), .A2(new_n14629_), .ZN(new_n14631_));
  OAI21_X1   g14567(.A1(new_n14627_), .A2(new_n14630_), .B(new_n14631_), .ZN(new_n14632_));
  NAND2_X1   g14568(.A1(new_n14333_), .A2(new_n14327_), .ZN(new_n14633_));
  NOR2_X1    g14569(.A1(new_n14633_), .A2(new_n14632_), .ZN(new_n14634_));
  NOR3_X1    g14570(.A1(new_n14184_), .A2(new_n14151_), .A3(new_n14338_), .ZN(new_n14635_));
  AOI21_X1   g14571(.A1(new_n14336_), .A2(new_n14335_), .B(new_n14042_), .ZN(new_n14636_));
  OAI21_X1   g14572(.A1(new_n14636_), .A2(new_n14635_), .B(new_n14327_), .ZN(new_n14637_));
  OAI22_X1   g14573(.A1(new_n14637_), .A2(new_n14634_), .B1(new_n14185_), .B2(new_n14042_), .ZN(new_n14638_));
  XOR2_X1    g14574(.A1(new_n14346_), .A2(\a[23] ), .Z(new_n14639_));
  NAND3_X1   g14575(.A1(new_n14369_), .A2(new_n14371_), .A3(new_n14370_), .ZN(new_n14640_));
  OAI21_X1   g14576(.A1(new_n14366_), .A2(new_n14361_), .B(new_n14367_), .ZN(new_n14641_));
  NAND3_X1   g14577(.A1(new_n14641_), .A2(new_n14639_), .A3(new_n14640_), .ZN(new_n14642_));
  NAND2_X1   g14578(.A1(new_n14638_), .A2(new_n14642_), .ZN(new_n14643_));
  OAI21_X1   g14579(.A1(new_n14400_), .A2(new_n14399_), .B(new_n14396_), .ZN(new_n14644_));
  NAND3_X1   g14580(.A1(new_n14401_), .A2(new_n14388_), .A3(new_n14391_), .ZN(new_n14645_));
  AOI22_X1   g14581(.A1(new_n14644_), .A2(new_n14645_), .B1(new_n14643_), .B2(new_n14374_), .ZN(new_n14646_));
  AOI21_X1   g14582(.A1(new_n14402_), .A2(new_n14397_), .B(new_n14375_), .ZN(new_n14647_));
  NOR2_X1    g14583(.A1(new_n14646_), .A2(new_n14647_), .ZN(new_n14648_));
  INV_X1     g14584(.I(new_n14648_), .ZN(new_n14649_));
  NOR3_X1    g14585(.A1(new_n14639_), .A2(new_n14372_), .A3(new_n14368_), .ZN(new_n14650_));
  AOI21_X1   g14586(.A1(new_n14640_), .A2(new_n14641_), .B(new_n14347_), .ZN(new_n14651_));
  NOR2_X1    g14587(.A1(new_n14651_), .A2(new_n14650_), .ZN(new_n14652_));
  NOR2_X1    g14588(.A1(new_n14652_), .A2(new_n14342_), .ZN(new_n14653_));
  AOI21_X1   g14589(.A1(new_n14640_), .A2(new_n14641_), .B(new_n14639_), .ZN(new_n14654_));
  NOR2_X1    g14590(.A1(new_n14654_), .A2(new_n14373_), .ZN(new_n14655_));
  NOR2_X1    g14591(.A1(new_n14638_), .A2(new_n14655_), .ZN(new_n14656_));
  INV_X1     g14592(.I(new_n11941_), .ZN(new_n14657_));
  AOI21_X1   g14593(.A1(new_n14657_), .A2(new_n11906_), .B(new_n8774_), .ZN(new_n14658_));
  AOI22_X1   g14594(.A1(new_n11899_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n10889_), .ZN(new_n14659_));
  NOR2_X1    g14595(.A1(new_n8774_), .A2(new_n4097_), .ZN(new_n14660_));
  OAI21_X1   g14596(.A1(new_n14660_), .A2(new_n14659_), .B(new_n3773_), .ZN(new_n14661_));
  NOR3_X1    g14597(.A1(new_n14658_), .A2(new_n11942_), .A3(new_n14661_), .ZN(new_n14662_));
  XOR2_X1    g14598(.A1(new_n14662_), .A2(new_n3035_), .Z(new_n14663_));
  OAI21_X1   g14599(.A1(new_n14656_), .A2(new_n14653_), .B(new_n14663_), .ZN(new_n14664_));
  AOI22_X1   g14600(.A1(new_n10886_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n10872_), .ZN(new_n14665_));
  NOR2_X1    g14601(.A1(new_n10892_), .A2(new_n4097_), .ZN(new_n14666_));
  OAI21_X1   g14602(.A1(new_n14665_), .A2(new_n14666_), .B(new_n3773_), .ZN(new_n14667_));
  NOR3_X1    g14603(.A1(new_n12776_), .A2(\a[20] ), .A3(new_n14667_), .ZN(new_n14668_));
  INV_X1     g14604(.I(new_n12773_), .ZN(new_n14669_));
  NOR3_X1    g14605(.A1(new_n14669_), .A2(new_n12774_), .A3(new_n14667_), .ZN(new_n14670_));
  NOR2_X1    g14606(.A1(new_n14670_), .A2(new_n3035_), .ZN(new_n14671_));
  NOR2_X1    g14607(.A1(new_n14668_), .A2(new_n14671_), .ZN(new_n14672_));
  INV_X1     g14608(.I(new_n14633_), .ZN(new_n14673_));
  NAND2_X1   g14609(.A1(new_n14673_), .A2(new_n14632_), .ZN(new_n14674_));
  NAND2_X1   g14610(.A1(new_n14633_), .A2(new_n14316_), .ZN(new_n14675_));
  NAND2_X1   g14611(.A1(new_n14674_), .A2(new_n14675_), .ZN(new_n14676_));
  NAND2_X1   g14612(.A1(new_n14676_), .A2(new_n14672_), .ZN(new_n14677_));
  AOI21_X1   g14613(.A1(new_n14334_), .A2(new_n14327_), .B(new_n14042_), .ZN(new_n14678_));
  AOI22_X1   g14614(.A1(new_n14320_), .A2(new_n14317_), .B1(new_n14324_), .B2(new_n14326_), .ZN(new_n14679_));
  OAI21_X1   g14615(.A1(new_n14632_), .A2(new_n14679_), .B(new_n14327_), .ZN(new_n14680_));
  NOR2_X1    g14616(.A1(new_n14680_), .A2(new_n14338_), .ZN(new_n14681_));
  OAI21_X1   g14617(.A1(new_n14678_), .A2(new_n14681_), .B(new_n14185_), .ZN(new_n14682_));
  INV_X1     g14618(.I(new_n14185_), .ZN(new_n14683_));
  NAND2_X1   g14619(.A1(new_n14680_), .A2(new_n14338_), .ZN(new_n14684_));
  NAND3_X1   g14620(.A1(new_n14334_), .A2(new_n14042_), .A3(new_n14327_), .ZN(new_n14685_));
  NAND3_X1   g14621(.A1(new_n14685_), .A2(new_n14684_), .A3(new_n14683_), .ZN(new_n14686_));
  AOI22_X1   g14622(.A1(new_n10886_), .A2(new_n3770_), .B1(new_n10889_), .B2(new_n3776_), .ZN(new_n14687_));
  NOR2_X1    g14623(.A1(new_n10899_), .A2(new_n4097_), .ZN(new_n14688_));
  OAI21_X1   g14624(.A1(new_n14688_), .A2(new_n14687_), .B(new_n3773_), .ZN(new_n14689_));
  INV_X1     g14625(.I(new_n14689_), .ZN(new_n14690_));
  NAND3_X1   g14626(.A1(new_n11903_), .A2(new_n11907_), .A3(new_n14690_), .ZN(new_n14691_));
  XOR2_X1    g14627(.A1(new_n14691_), .A2(new_n3035_), .Z(new_n14692_));
  AOI21_X1   g14628(.A1(new_n14682_), .A2(new_n14686_), .B(new_n14692_), .ZN(new_n14693_));
  NAND3_X1   g14629(.A1(new_n14682_), .A2(new_n14686_), .A3(new_n14692_), .ZN(new_n14694_));
  OAI21_X1   g14630(.A1(new_n14677_), .A2(new_n14693_), .B(new_n14694_), .ZN(new_n14695_));
  NOR2_X1    g14631(.A1(new_n14637_), .A2(new_n14634_), .ZN(new_n14696_));
  OAI22_X1   g14632(.A1(new_n14696_), .A2(new_n14186_), .B1(new_n14650_), .B2(new_n14651_), .ZN(new_n14697_));
  NAND2_X1   g14633(.A1(new_n14374_), .A2(new_n14642_), .ZN(new_n14698_));
  NAND2_X1   g14634(.A1(new_n14342_), .A2(new_n14698_), .ZN(new_n14699_));
  XOR2_X1    g14635(.A1(new_n14662_), .A2(\a[20] ), .Z(new_n14700_));
  NAND3_X1   g14636(.A1(new_n14697_), .A2(new_n14699_), .A3(new_n14700_), .ZN(new_n14701_));
  NAND2_X1   g14637(.A1(new_n14664_), .A2(new_n14701_), .ZN(new_n14702_));
  OAI21_X1   g14638(.A1(new_n14702_), .A2(new_n14695_), .B(new_n14664_), .ZN(new_n14703_));
  OAI22_X1   g14639(.A1(new_n8774_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n10899_), .ZN(new_n14704_));
  NAND2_X1   g14640(.A1(new_n11996_), .A2(new_n4096_), .ZN(new_n14705_));
  AOI21_X1   g14641(.A1(new_n14705_), .A2(new_n14704_), .B(new_n4095_), .ZN(new_n14706_));
  NAND2_X1   g14642(.A1(new_n12001_), .A2(new_n14706_), .ZN(new_n14707_));
  XOR2_X1    g14643(.A1(new_n14707_), .A2(new_n3035_), .Z(new_n14708_));
  INV_X1     g14644(.I(new_n14708_), .ZN(new_n14709_));
  NAND2_X1   g14645(.A1(new_n14703_), .A2(new_n14709_), .ZN(new_n14710_));
  INV_X1     g14646(.I(new_n14677_), .ZN(new_n14711_));
  AOI21_X1   g14647(.A1(new_n14685_), .A2(new_n14684_), .B(new_n14683_), .ZN(new_n14712_));
  NOR3_X1    g14648(.A1(new_n14678_), .A2(new_n14681_), .A3(new_n14185_), .ZN(new_n14713_));
  XOR2_X1    g14649(.A1(new_n14691_), .A2(\a[20] ), .Z(new_n14714_));
  OAI21_X1   g14650(.A1(new_n14712_), .A2(new_n14713_), .B(new_n14714_), .ZN(new_n14715_));
  NAND2_X1   g14651(.A1(new_n14715_), .A2(new_n14711_), .ZN(new_n14716_));
  NAND4_X1   g14652(.A1(new_n14716_), .A2(new_n14664_), .A3(new_n14694_), .A4(new_n14701_), .ZN(new_n14717_));
  NAND3_X1   g14653(.A1(new_n14717_), .A2(new_n14664_), .A3(new_n14708_), .ZN(new_n14718_));
  AOI21_X1   g14654(.A1(new_n14710_), .A2(new_n14718_), .B(new_n14649_), .ZN(new_n14719_));
  AOI21_X1   g14655(.A1(new_n14717_), .A2(new_n14664_), .B(new_n14708_), .ZN(new_n14720_));
  NOR2_X1    g14656(.A1(new_n14703_), .A2(new_n14709_), .ZN(new_n14721_));
  NOR3_X1    g14657(.A1(new_n14721_), .A2(new_n14720_), .A3(new_n14648_), .ZN(new_n14722_));
  NOR3_X1    g14658(.A1(new_n14722_), .A2(new_n14719_), .A3(new_n14599_), .ZN(new_n14723_));
  INV_X1     g14659(.I(new_n14599_), .ZN(new_n14724_));
  OAI21_X1   g14660(.A1(new_n14721_), .A2(new_n14720_), .B(new_n14648_), .ZN(new_n14725_));
  NAND3_X1   g14661(.A1(new_n14710_), .A2(new_n14718_), .A3(new_n14649_), .ZN(new_n14726_));
  AOI21_X1   g14662(.A1(new_n14725_), .A2(new_n14726_), .B(new_n14724_), .ZN(new_n14727_));
  NOR2_X1    g14663(.A1(new_n14702_), .A2(new_n14695_), .ZN(new_n14728_));
  AOI22_X1   g14664(.A1(new_n14716_), .A2(new_n14694_), .B1(new_n14664_), .B2(new_n14701_), .ZN(new_n14729_));
  OAI22_X1   g14665(.A1(new_n8758_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8766_), .ZN(new_n14730_));
  NAND2_X1   g14666(.A1(new_n8746_), .A2(new_n4469_), .ZN(new_n14731_));
  AOI21_X1   g14667(.A1(new_n14731_), .A2(new_n14730_), .B(new_n4468_), .ZN(new_n14732_));
  NAND2_X1   g14668(.A1(new_n11964_), .A2(new_n14732_), .ZN(new_n14733_));
  XOR2_X1    g14669(.A1(new_n14733_), .A2(new_n3372_), .Z(new_n14734_));
  NOR3_X1    g14670(.A1(new_n14728_), .A2(new_n14729_), .A3(new_n14734_), .ZN(new_n14735_));
  NAND2_X1   g14671(.A1(new_n14702_), .A2(new_n14695_), .ZN(new_n14736_));
  XOR2_X1    g14672(.A1(new_n14733_), .A2(\a[17] ), .Z(new_n14737_));
  AOI21_X1   g14673(.A1(new_n14736_), .A2(new_n14717_), .B(new_n14737_), .ZN(new_n14738_));
  AOI21_X1   g14674(.A1(new_n14715_), .A2(new_n14694_), .B(new_n14677_), .ZN(new_n14739_));
  NAND3_X1   g14675(.A1(new_n14682_), .A2(new_n14686_), .A3(new_n14714_), .ZN(new_n14740_));
  OAI21_X1   g14676(.A1(new_n14712_), .A2(new_n14713_), .B(new_n14692_), .ZN(new_n14741_));
  AOI21_X1   g14677(.A1(new_n14740_), .A2(new_n14741_), .B(new_n14711_), .ZN(new_n14742_));
  AOI22_X1   g14678(.A1(new_n4292_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n4298_), .ZN(new_n14743_));
  NOR2_X1    g14679(.A1(new_n8758_), .A2(new_n4470_), .ZN(new_n14744_));
  OAI21_X1   g14680(.A1(new_n14743_), .A2(new_n14744_), .B(new_n4295_), .ZN(new_n14745_));
  NOR2_X1    g14681(.A1(new_n12053_), .A2(new_n14745_), .ZN(new_n14746_));
  XOR2_X1    g14682(.A1(new_n14746_), .A2(\a[17] ), .Z(new_n14747_));
  NOR3_X1    g14683(.A1(new_n14742_), .A2(new_n14739_), .A3(new_n14747_), .ZN(new_n14748_));
  OAI22_X1   g14684(.A1(new_n8774_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n10899_), .ZN(new_n14749_));
  NAND2_X1   g14685(.A1(new_n11996_), .A2(new_n4469_), .ZN(new_n14750_));
  AOI21_X1   g14686(.A1(new_n14750_), .A2(new_n14749_), .B(new_n4468_), .ZN(new_n14751_));
  NAND3_X1   g14687(.A1(new_n12001_), .A2(new_n3372_), .A3(new_n14751_), .ZN(new_n14752_));
  NAND3_X1   g14688(.A1(new_n10901_), .A2(new_n10906_), .A3(new_n10903_), .ZN(new_n14753_));
  AOI21_X1   g14689(.A1(new_n12047_), .A2(new_n14753_), .B(new_n8766_), .ZN(new_n14754_));
  NAND3_X1   g14690(.A1(new_n10901_), .A2(new_n8774_), .A3(new_n10903_), .ZN(new_n14755_));
  OAI21_X1   g14691(.A1(new_n10912_), .A2(new_n10902_), .B(new_n10906_), .ZN(new_n14756_));
  AOI21_X1   g14692(.A1(new_n14756_), .A2(new_n14755_), .B(new_n11996_), .ZN(new_n14757_));
  OAI21_X1   g14693(.A1(new_n14754_), .A2(new_n14757_), .B(new_n14751_), .ZN(new_n14758_));
  NAND2_X1   g14694(.A1(new_n14758_), .A2(\a[17] ), .ZN(new_n14759_));
  NAND2_X1   g14695(.A1(new_n14759_), .A2(new_n14752_), .ZN(new_n14760_));
  NAND2_X1   g14696(.A1(new_n14670_), .A2(new_n3035_), .ZN(new_n14761_));
  OAI21_X1   g14697(.A1(new_n12776_), .A2(new_n14667_), .B(\a[20] ), .ZN(new_n14762_));
  NAND3_X1   g14698(.A1(new_n14762_), .A2(new_n14761_), .A3(new_n14632_), .ZN(new_n14763_));
  OAI21_X1   g14699(.A1(new_n14668_), .A2(new_n14671_), .B(new_n14316_), .ZN(new_n14764_));
  AOI21_X1   g14700(.A1(new_n14764_), .A2(new_n14763_), .B(new_n14633_), .ZN(new_n14765_));
  NOR3_X1    g14701(.A1(new_n14668_), .A2(new_n14671_), .A3(new_n14316_), .ZN(new_n14766_));
  AOI21_X1   g14702(.A1(new_n14762_), .A2(new_n14761_), .B(new_n14632_), .ZN(new_n14767_));
  NOR3_X1    g14703(.A1(new_n14767_), .A2(new_n14766_), .A3(new_n14673_), .ZN(new_n14768_));
  NOR2_X1    g14704(.A1(new_n14768_), .A2(new_n14765_), .ZN(new_n14769_));
  NOR2_X1    g14705(.A1(new_n14769_), .A2(new_n14760_), .ZN(new_n14770_));
  NOR2_X1    g14706(.A1(new_n12770_), .A2(new_n12771_), .ZN(new_n14771_));
  NOR2_X1    g14707(.A1(new_n10909_), .A2(new_n13102_), .ZN(new_n14772_));
  OAI22_X1   g14708(.A1(new_n10871_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8778_), .ZN(new_n14773_));
  NAND2_X1   g14709(.A1(new_n10886_), .A2(new_n4469_), .ZN(new_n14774_));
  AOI21_X1   g14710(.A1(new_n14774_), .A2(new_n14773_), .B(new_n4468_), .ZN(new_n14775_));
  OAI21_X1   g14711(.A1(new_n14771_), .A2(new_n14772_), .B(new_n14775_), .ZN(new_n14776_));
  XOR2_X1    g14712(.A1(new_n14776_), .A2(\a[17] ), .Z(new_n14777_));
  OAI22_X1   g14713(.A1(new_n10775_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n10777_), .ZN(new_n14778_));
  OAI21_X1   g14714(.A1(new_n4097_), .A2(new_n10798_), .B(new_n14778_), .ZN(new_n14779_));
  NAND3_X1   g14715(.A1(new_n12883_), .A2(new_n3773_), .A3(new_n14779_), .ZN(new_n14780_));
  NOR2_X1    g14716(.A1(new_n14780_), .A2(\a[20] ), .ZN(new_n14781_));
  INV_X1     g14717(.I(new_n14781_), .ZN(new_n14782_));
  NAND2_X1   g14718(.A1(new_n14780_), .A2(\a[20] ), .ZN(new_n14783_));
  AOI21_X1   g14719(.A1(new_n14782_), .A2(new_n14783_), .B(new_n14206_), .ZN(new_n14784_));
  INV_X1     g14720(.I(new_n14784_), .ZN(new_n14785_));
  INV_X1     g14721(.I(new_n12827_), .ZN(new_n14786_));
  NOR2_X1    g14722(.A1(new_n14786_), .A2(new_n12828_), .ZN(new_n14787_));
  AOI22_X1   g14723(.A1(new_n10794_), .A2(new_n3770_), .B1(new_n3776_), .B2(new_n12823_), .ZN(new_n14788_));
  AOI21_X1   g14724(.A1(new_n4096_), .A2(new_n10800_), .B(new_n14788_), .ZN(new_n14789_));
  NOR3_X1    g14725(.A1(new_n14789_), .A2(new_n14787_), .A3(new_n4095_), .ZN(new_n14790_));
  NOR2_X1    g14726(.A1(new_n10794_), .A2(new_n12823_), .ZN(new_n14791_));
  NOR2_X1    g14727(.A1(new_n12826_), .A2(new_n10775_), .ZN(new_n14792_));
  NOR2_X1    g14728(.A1(new_n14791_), .A2(new_n14792_), .ZN(new_n14793_));
  NAND2_X1   g14729(.A1(new_n10794_), .A2(new_n3776_), .ZN(new_n14794_));
  NOR2_X1    g14730(.A1(new_n3762_), .A2(new_n3772_), .ZN(new_n14795_));
  NAND3_X1   g14731(.A1(new_n14793_), .A2(new_n14794_), .A3(new_n14795_), .ZN(new_n14796_));
  NOR2_X1    g14732(.A1(new_n12826_), .A2(new_n3762_), .ZN(new_n14797_));
  NOR4_X1    g14733(.A1(new_n14790_), .A2(new_n3035_), .A3(new_n14796_), .A4(new_n14797_), .ZN(new_n14798_));
  INV_X1     g14734(.I(new_n14206_), .ZN(new_n14799_));
  INV_X1     g14735(.I(new_n14783_), .ZN(new_n14800_));
  NOR3_X1    g14736(.A1(new_n14800_), .A2(new_n14799_), .A3(new_n14781_), .ZN(new_n14801_));
  OAI21_X1   g14737(.A1(new_n14798_), .A2(new_n14801_), .B(new_n14785_), .ZN(new_n14802_));
  XOR2_X1    g14738(.A1(new_n14205_), .A2(new_n14208_), .Z(new_n14803_));
  AOI22_X1   g14739(.A1(new_n9529_), .A2(new_n3776_), .B1(new_n10800_), .B2(new_n3770_), .ZN(new_n14804_));
  AOI21_X1   g14740(.A1(new_n10839_), .A2(new_n4096_), .B(new_n14804_), .ZN(new_n14805_));
  OR3_X2     g14741(.A1(new_n13534_), .A2(new_n4095_), .A3(new_n14805_), .Z(new_n14806_));
  NOR2_X1    g14742(.A1(new_n14806_), .A2(\a[20] ), .ZN(new_n14807_));
  INV_X1     g14743(.I(new_n14807_), .ZN(new_n14808_));
  NAND2_X1   g14744(.A1(new_n14806_), .A2(\a[20] ), .ZN(new_n14809_));
  NAND3_X1   g14745(.A1(new_n14808_), .A2(new_n14803_), .A3(new_n14809_), .ZN(new_n14810_));
  AOI21_X1   g14746(.A1(new_n14808_), .A2(new_n14809_), .B(new_n14803_), .ZN(new_n14811_));
  AOI21_X1   g14747(.A1(new_n14802_), .A2(new_n14810_), .B(new_n14811_), .ZN(new_n14812_));
  NAND3_X1   g14748(.A1(new_n14602_), .A2(new_n14199_), .A3(new_n14200_), .ZN(new_n14813_));
  OAI21_X1   g14749(.A1(new_n14601_), .A2(new_n14198_), .B(new_n14209_), .ZN(new_n14814_));
  NAND2_X1   g14750(.A1(new_n14813_), .A2(new_n14814_), .ZN(new_n14815_));
  INV_X1     g14751(.I(new_n14815_), .ZN(new_n14816_));
  AOI22_X1   g14752(.A1(new_n10839_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n9529_), .ZN(new_n14817_));
  NOR2_X1    g14753(.A1(new_n10846_), .A2(new_n4097_), .ZN(new_n14818_));
  OAI21_X1   g14754(.A1(new_n14817_), .A2(new_n14818_), .B(new_n3773_), .ZN(new_n14819_));
  NOR2_X1    g14755(.A1(new_n12946_), .A2(new_n14819_), .ZN(new_n14820_));
  XOR2_X1    g14756(.A1(new_n14820_), .A2(\a[20] ), .Z(new_n14821_));
  NOR2_X1    g14757(.A1(new_n14816_), .A2(new_n14821_), .ZN(new_n14822_));
  NAND2_X1   g14758(.A1(new_n14816_), .A2(new_n14821_), .ZN(new_n14823_));
  OAI21_X1   g14759(.A1(new_n14812_), .A2(new_n14822_), .B(new_n14823_), .ZN(new_n14824_));
  INV_X1     g14760(.I(new_n14058_), .ZN(new_n14825_));
  NAND3_X1   g14761(.A1(new_n14191_), .A2(new_n14825_), .A3(new_n14192_), .ZN(new_n14826_));
  NAND2_X1   g14762(.A1(new_n14191_), .A2(new_n14192_), .ZN(new_n14827_));
  NAND2_X1   g14763(.A1(new_n14827_), .A2(new_n14058_), .ZN(new_n14828_));
  AOI21_X1   g14764(.A1(new_n14826_), .A2(new_n14828_), .B(new_n14210_), .ZN(new_n14829_));
  AOI21_X1   g14765(.A1(new_n14600_), .A2(new_n14211_), .B(new_n14603_), .ZN(new_n14830_));
  NOR2_X1    g14766(.A1(new_n14830_), .A2(new_n14829_), .ZN(new_n14831_));
  AOI22_X1   g14767(.A1(new_n10839_), .A2(new_n3770_), .B1(new_n12936_), .B2(new_n3776_), .ZN(new_n14832_));
  NOR2_X1    g14768(.A1(new_n9478_), .A2(new_n4097_), .ZN(new_n14833_));
  NOR2_X1    g14769(.A1(new_n14832_), .A2(new_n14833_), .ZN(new_n14834_));
  NOR2_X1    g14770(.A1(new_n14834_), .A2(new_n4095_), .ZN(new_n14835_));
  NAND2_X1   g14771(.A1(new_n13566_), .A2(new_n14835_), .ZN(new_n14836_));
  NOR2_X1    g14772(.A1(new_n14836_), .A2(\a[20] ), .ZN(new_n14837_));
  INV_X1     g14773(.I(new_n14837_), .ZN(new_n14838_));
  NAND2_X1   g14774(.A1(new_n14836_), .A2(\a[20] ), .ZN(new_n14839_));
  NAND3_X1   g14775(.A1(new_n14831_), .A2(new_n14838_), .A3(new_n14839_), .ZN(new_n14840_));
  AOI21_X1   g14776(.A1(new_n14838_), .A2(new_n14839_), .B(new_n14831_), .ZN(new_n14841_));
  AOI21_X1   g14777(.A1(new_n14824_), .A2(new_n14840_), .B(new_n14841_), .ZN(new_n14842_));
  NAND3_X1   g14778(.A1(new_n14214_), .A2(new_n14611_), .A3(new_n14220_), .ZN(new_n14843_));
  OAI21_X1   g14779(.A1(new_n14221_), .A2(new_n14219_), .B(new_n14610_), .ZN(new_n14844_));
  AOI21_X1   g14780(.A1(new_n14843_), .A2(new_n14844_), .B(new_n14212_), .ZN(new_n14845_));
  AOI21_X1   g14781(.A1(new_n14223_), .A2(new_n14612_), .B(new_n14605_), .ZN(new_n14846_));
  NOR2_X1    g14782(.A1(new_n14846_), .A2(new_n14845_), .ZN(new_n14847_));
  OAI22_X1   g14783(.A1(new_n9478_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n10846_), .ZN(new_n14848_));
  NAND2_X1   g14784(.A1(new_n10854_), .A2(new_n4096_), .ZN(new_n14849_));
  AOI21_X1   g14785(.A1(new_n14848_), .A2(new_n14849_), .B(new_n4095_), .ZN(new_n14850_));
  NAND3_X1   g14786(.A1(new_n13016_), .A2(new_n3035_), .A3(new_n14850_), .ZN(new_n14851_));
  AOI21_X1   g14787(.A1(new_n13016_), .A2(new_n14850_), .B(new_n3035_), .ZN(new_n14852_));
  INV_X1     g14788(.I(new_n14852_), .ZN(new_n14853_));
  NAND2_X1   g14789(.A1(new_n14853_), .A2(new_n14851_), .ZN(new_n14854_));
  NOR2_X1    g14790(.A1(new_n14854_), .A2(new_n14847_), .ZN(new_n14855_));
  NAND2_X1   g14791(.A1(new_n14854_), .A2(new_n14847_), .ZN(new_n14856_));
  OAI21_X1   g14792(.A1(new_n14842_), .A2(new_n14855_), .B(new_n14856_), .ZN(new_n14857_));
  NOR2_X1    g14793(.A1(new_n14222_), .A2(new_n14212_), .ZN(new_n14858_));
  NOR2_X1    g14794(.A1(new_n14233_), .A2(new_n14239_), .ZN(new_n14859_));
  NOR2_X1    g14795(.A1(new_n14240_), .A2(new_n14244_), .ZN(new_n14860_));
  OAI22_X1   g14796(.A1(new_n14859_), .A2(new_n14860_), .B1(new_n14858_), .B2(new_n14613_), .ZN(new_n14861_));
  OAI21_X1   g14797(.A1(new_n14246_), .A2(new_n14615_), .B(new_n14614_), .ZN(new_n14862_));
  NAND2_X1   g14798(.A1(new_n14862_), .A2(new_n14861_), .ZN(new_n14863_));
  OAI22_X1   g14799(.A1(new_n9478_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n10853_), .ZN(new_n14864_));
  NAND2_X1   g14800(.A1(new_n10862_), .A2(new_n4096_), .ZN(new_n14865_));
  AOI21_X1   g14801(.A1(new_n14864_), .A2(new_n14865_), .B(new_n4095_), .ZN(new_n14866_));
  NAND3_X1   g14802(.A1(new_n13484_), .A2(new_n3035_), .A3(new_n14866_), .ZN(new_n14867_));
  INV_X1     g14803(.I(new_n14867_), .ZN(new_n14868_));
  AOI21_X1   g14804(.A1(new_n13484_), .A2(new_n14866_), .B(new_n3035_), .ZN(new_n14869_));
  NOR2_X1    g14805(.A1(new_n14868_), .A2(new_n14869_), .ZN(new_n14870_));
  NAND2_X1   g14806(.A1(new_n14863_), .A2(new_n14870_), .ZN(new_n14871_));
  INV_X1     g14807(.I(new_n14869_), .ZN(new_n14872_));
  NAND2_X1   g14808(.A1(new_n14872_), .A2(new_n14867_), .ZN(new_n14873_));
  NAND3_X1   g14809(.A1(new_n14873_), .A2(new_n14862_), .A3(new_n14861_), .ZN(new_n14874_));
  INV_X1     g14810(.I(new_n14874_), .ZN(new_n14875_));
  AOI21_X1   g14811(.A1(new_n14857_), .A2(new_n14871_), .B(new_n14875_), .ZN(new_n14876_));
  NAND3_X1   g14812(.A1(new_n14264_), .A2(new_n14259_), .A3(new_n14257_), .ZN(new_n14877_));
  OAI21_X1   g14813(.A1(new_n14266_), .A2(new_n14265_), .B(new_n14253_), .ZN(new_n14878_));
  NAND2_X1   g14814(.A1(new_n14878_), .A2(new_n14877_), .ZN(new_n14879_));
  NAND2_X1   g14815(.A1(new_n14267_), .A2(new_n14260_), .ZN(new_n14880_));
  MUX2_X1    g14816(.I0(new_n14880_), .I1(new_n14879_), .S(new_n14616_), .Z(new_n14881_));
  OAI22_X1   g14817(.A1(new_n10861_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n10853_), .ZN(new_n14882_));
  NAND2_X1   g14818(.A1(new_n8785_), .A2(new_n4096_), .ZN(new_n14883_));
  AOI21_X1   g14819(.A1(new_n14883_), .A2(new_n14882_), .B(new_n4095_), .ZN(new_n14884_));
  NAND3_X1   g14820(.A1(new_n13592_), .A2(new_n3035_), .A3(new_n14884_), .ZN(new_n14885_));
  NAND2_X1   g14821(.A1(new_n13592_), .A2(new_n14884_), .ZN(new_n14886_));
  NAND2_X1   g14822(.A1(new_n14886_), .A2(\a[20] ), .ZN(new_n14887_));
  NAND2_X1   g14823(.A1(new_n14887_), .A2(new_n14885_), .ZN(new_n14888_));
  INV_X1     g14824(.I(new_n14888_), .ZN(new_n14889_));
  NAND2_X1   g14825(.A1(new_n14881_), .A2(new_n14889_), .ZN(new_n14890_));
  AOI21_X1   g14826(.A1(new_n14260_), .A2(new_n14267_), .B(new_n14616_), .ZN(new_n14891_));
  AOI21_X1   g14827(.A1(new_n14616_), .A2(new_n14879_), .B(new_n14891_), .ZN(new_n14892_));
  NAND2_X1   g14828(.A1(new_n14892_), .A2(new_n14888_), .ZN(new_n14893_));
  AOI21_X1   g14829(.A1(new_n14890_), .A2(new_n14893_), .B(new_n14876_), .ZN(new_n14894_));
  INV_X1     g14830(.I(new_n14802_), .ZN(new_n14895_));
  XOR2_X1    g14831(.A1(new_n14205_), .A2(new_n14207_), .Z(new_n14896_));
  AND2_X2    g14832(.A1(new_n14806_), .A2(\a[20] ), .Z(new_n14897_));
  NOR3_X1    g14833(.A1(new_n14897_), .A2(new_n14896_), .A3(new_n14807_), .ZN(new_n14898_));
  OAI21_X1   g14834(.A1(new_n14897_), .A2(new_n14807_), .B(new_n14896_), .ZN(new_n14899_));
  OAI21_X1   g14835(.A1(new_n14895_), .A2(new_n14898_), .B(new_n14899_), .ZN(new_n14900_));
  XOR2_X1    g14836(.A1(new_n14820_), .A2(new_n3035_), .Z(new_n14901_));
  NAND2_X1   g14837(.A1(new_n14901_), .A2(new_n14815_), .ZN(new_n14902_));
  NOR2_X1    g14838(.A1(new_n14901_), .A2(new_n14815_), .ZN(new_n14903_));
  AOI21_X1   g14839(.A1(new_n14900_), .A2(new_n14902_), .B(new_n14903_), .ZN(new_n14904_));
  NAND2_X1   g14840(.A1(new_n14828_), .A2(new_n14826_), .ZN(new_n14905_));
  NAND2_X1   g14841(.A1(new_n14905_), .A2(new_n14603_), .ZN(new_n14906_));
  OAI21_X1   g14842(.A1(new_n14193_), .A2(new_n14604_), .B(new_n14210_), .ZN(new_n14907_));
  NAND2_X1   g14843(.A1(new_n14907_), .A2(new_n14906_), .ZN(new_n14908_));
  INV_X1     g14844(.I(new_n14839_), .ZN(new_n14909_));
  NOR3_X1    g14845(.A1(new_n14908_), .A2(new_n14909_), .A3(new_n14837_), .ZN(new_n14910_));
  OAI21_X1   g14846(.A1(new_n14909_), .A2(new_n14837_), .B(new_n14908_), .ZN(new_n14911_));
  OAI21_X1   g14847(.A1(new_n14904_), .A2(new_n14910_), .B(new_n14911_), .ZN(new_n14912_));
  NOR3_X1    g14848(.A1(new_n14610_), .A2(new_n14219_), .A3(new_n14221_), .ZN(new_n14913_));
  AOI21_X1   g14849(.A1(new_n14611_), .A2(new_n14220_), .B(new_n14214_), .ZN(new_n14914_));
  OAI21_X1   g14850(.A1(new_n14914_), .A2(new_n14913_), .B(new_n14605_), .ZN(new_n14915_));
  OAI21_X1   g14851(.A1(new_n14222_), .A2(new_n14613_), .B(new_n14212_), .ZN(new_n14916_));
  NAND2_X1   g14852(.A1(new_n14915_), .A2(new_n14916_), .ZN(new_n14917_));
  INV_X1     g14853(.I(new_n14851_), .ZN(new_n14918_));
  NOR2_X1    g14854(.A1(new_n14918_), .A2(new_n14852_), .ZN(new_n14919_));
  NAND2_X1   g14855(.A1(new_n14919_), .A2(new_n14917_), .ZN(new_n14920_));
  NOR2_X1    g14856(.A1(new_n14919_), .A2(new_n14917_), .ZN(new_n14921_));
  AOI21_X1   g14857(.A1(new_n14912_), .A2(new_n14920_), .B(new_n14921_), .ZN(new_n14922_));
  AOI21_X1   g14858(.A1(new_n14861_), .A2(new_n14862_), .B(new_n14873_), .ZN(new_n14923_));
  OAI21_X1   g14859(.A1(new_n14922_), .A2(new_n14923_), .B(new_n14874_), .ZN(new_n14924_));
  NAND2_X1   g14860(.A1(new_n14892_), .A2(new_n14889_), .ZN(new_n14925_));
  NAND2_X1   g14861(.A1(new_n14881_), .A2(new_n14888_), .ZN(new_n14926_));
  AOI21_X1   g14862(.A1(new_n14926_), .A2(new_n14925_), .B(new_n14924_), .ZN(new_n14927_));
  OAI21_X1   g14863(.A1(new_n14894_), .A2(new_n14927_), .B(new_n14777_), .ZN(new_n14928_));
  INV_X1     g14864(.I(new_n14928_), .ZN(new_n14929_));
  OAI22_X1   g14865(.A1(new_n8784_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n10861_), .ZN(new_n14930_));
  NAND2_X1   g14866(.A1(new_n8779_), .A2(new_n4469_), .ZN(new_n14931_));
  AOI21_X1   g14867(.A1(new_n14931_), .A2(new_n14930_), .B(new_n4468_), .ZN(new_n14932_));
  AND3_X2    g14868(.A1(new_n12814_), .A2(new_n3372_), .A3(new_n14932_), .Z(new_n14933_));
  AOI21_X1   g14869(.A1(new_n12814_), .A2(new_n14932_), .B(new_n3372_), .ZN(new_n14934_));
  NOR2_X1    g14870(.A1(new_n14933_), .A2(new_n14934_), .ZN(new_n14935_));
  NAND2_X1   g14871(.A1(new_n14919_), .A2(new_n14847_), .ZN(new_n14936_));
  NAND2_X1   g14872(.A1(new_n14854_), .A2(new_n14917_), .ZN(new_n14937_));
  NAND2_X1   g14873(.A1(new_n14937_), .A2(new_n14936_), .ZN(new_n14938_));
  NAND2_X1   g14874(.A1(new_n14938_), .A2(new_n14912_), .ZN(new_n14939_));
  OAI21_X1   g14875(.A1(new_n14855_), .A2(new_n14921_), .B(new_n14842_), .ZN(new_n14940_));
  NAND2_X1   g14876(.A1(new_n14939_), .A2(new_n14940_), .ZN(new_n14941_));
  NAND2_X1   g14877(.A1(new_n14941_), .A2(new_n14935_), .ZN(new_n14942_));
  INV_X1     g14878(.I(new_n14797_), .ZN(new_n14943_));
  AOI22_X1   g14879(.A1(new_n12823_), .A2(new_n4292_), .B1(new_n4298_), .B2(new_n10800_), .ZN(new_n14944_));
  AOI21_X1   g14880(.A1(new_n4469_), .A2(new_n9529_), .B(new_n14944_), .ZN(new_n14945_));
  NOR3_X1    g14881(.A1(new_n13504_), .A2(new_n4468_), .A3(new_n14945_), .ZN(new_n14946_));
  NAND2_X1   g14882(.A1(new_n14946_), .A2(new_n3372_), .ZN(new_n14947_));
  NOR2_X1    g14883(.A1(new_n14946_), .A2(new_n3372_), .ZN(new_n14948_));
  INV_X1     g14884(.I(new_n14948_), .ZN(new_n14949_));
  NAND2_X1   g14885(.A1(new_n14949_), .A2(new_n14947_), .ZN(new_n14950_));
  NAND2_X1   g14886(.A1(new_n14950_), .A2(new_n14943_), .ZN(new_n14951_));
  AOI22_X1   g14887(.A1(new_n10794_), .A2(new_n4292_), .B1(new_n4298_), .B2(new_n12823_), .ZN(new_n14952_));
  AOI21_X1   g14888(.A1(new_n4469_), .A2(new_n10800_), .B(new_n14952_), .ZN(new_n14953_));
  NOR3_X1    g14889(.A1(new_n14953_), .A2(new_n14787_), .A3(new_n4468_), .ZN(new_n14954_));
  XOR2_X1    g14890(.A1(new_n14954_), .A2(\a[17] ), .Z(new_n14955_));
  NAND2_X1   g14891(.A1(new_n10794_), .A2(new_n4298_), .ZN(new_n14956_));
  NOR2_X1    g14892(.A1(new_n4284_), .A2(new_n4294_), .ZN(new_n14957_));
  NAND3_X1   g14893(.A1(new_n14793_), .A2(new_n14956_), .A3(new_n14957_), .ZN(new_n14958_));
  XOR2_X1    g14894(.A1(new_n14958_), .A2(new_n3372_), .Z(new_n14959_));
  NOR2_X1    g14895(.A1(new_n12826_), .A2(new_n4284_), .ZN(new_n14960_));
  NOR2_X1    g14896(.A1(new_n14960_), .A2(new_n3372_), .ZN(new_n14961_));
  INV_X1     g14897(.I(new_n14961_), .ZN(new_n14962_));
  NOR2_X1    g14898(.A1(new_n14959_), .A2(new_n14962_), .ZN(new_n14963_));
  NAND2_X1   g14899(.A1(new_n14963_), .A2(new_n14955_), .ZN(new_n14964_));
  INV_X1     g14900(.I(new_n14947_), .ZN(new_n14965_));
  NOR2_X1    g14901(.A1(new_n14965_), .A2(new_n14948_), .ZN(new_n14966_));
  NAND2_X1   g14902(.A1(new_n14966_), .A2(new_n14797_), .ZN(new_n14967_));
  NAND2_X1   g14903(.A1(new_n14967_), .A2(new_n14964_), .ZN(new_n14968_));
  NAND2_X1   g14904(.A1(new_n14968_), .A2(new_n14951_), .ZN(new_n14969_));
  XOR2_X1    g14905(.A1(new_n14796_), .A2(\a[20] ), .Z(new_n14970_));
  NOR2_X1    g14906(.A1(new_n14797_), .A2(new_n3035_), .ZN(new_n14971_));
  XOR2_X1    g14907(.A1(new_n14970_), .A2(new_n14971_), .Z(new_n14972_));
  AOI22_X1   g14908(.A1(new_n9529_), .A2(new_n4298_), .B1(new_n10800_), .B2(new_n4292_), .ZN(new_n14973_));
  AOI21_X1   g14909(.A1(new_n10839_), .A2(new_n4469_), .B(new_n14973_), .ZN(new_n14974_));
  OR3_X2     g14910(.A1(new_n13534_), .A2(new_n4468_), .A3(new_n14974_), .Z(new_n14975_));
  XOR2_X1    g14911(.A1(new_n14975_), .A2(\a[17] ), .Z(new_n14976_));
  NAND2_X1   g14912(.A1(new_n14976_), .A2(new_n14972_), .ZN(new_n14977_));
  NOR2_X1    g14913(.A1(new_n14976_), .A2(new_n14972_), .ZN(new_n14978_));
  AOI21_X1   g14914(.A1(new_n14969_), .A2(new_n14977_), .B(new_n14978_), .ZN(new_n14979_));
  XOR2_X1    g14915(.A1(new_n14790_), .A2(\a[20] ), .Z(new_n14980_));
  NOR3_X1    g14916(.A1(new_n14796_), .A2(new_n3035_), .A3(new_n14797_), .ZN(new_n14981_));
  INV_X1     g14917(.I(new_n14981_), .ZN(new_n14982_));
  AND2_X2    g14918(.A1(new_n14980_), .A2(new_n14982_), .Z(new_n14983_));
  NOR2_X1    g14919(.A1(new_n14980_), .A2(new_n14982_), .ZN(new_n14984_));
  NOR2_X1    g14920(.A1(new_n14983_), .A2(new_n14984_), .ZN(new_n14985_));
  AOI22_X1   g14921(.A1(new_n10839_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n9529_), .ZN(new_n14986_));
  NOR2_X1    g14922(.A1(new_n10846_), .A2(new_n4470_), .ZN(new_n14987_));
  OAI21_X1   g14923(.A1(new_n14986_), .A2(new_n14987_), .B(new_n4295_), .ZN(new_n14988_));
  NOR2_X1    g14924(.A1(new_n12946_), .A2(new_n14988_), .ZN(new_n14989_));
  XOR2_X1    g14925(.A1(new_n14989_), .A2(new_n3372_), .Z(new_n14990_));
  INV_X1     g14926(.I(new_n14990_), .ZN(new_n14991_));
  NOR2_X1    g14927(.A1(new_n14991_), .A2(new_n14985_), .ZN(new_n14992_));
  NAND2_X1   g14928(.A1(new_n14991_), .A2(new_n14985_), .ZN(new_n14993_));
  OAI21_X1   g14929(.A1(new_n14979_), .A2(new_n14992_), .B(new_n14993_), .ZN(new_n14994_));
  NAND2_X1   g14930(.A1(new_n14782_), .A2(new_n14783_), .ZN(new_n14995_));
  XOR2_X1    g14931(.A1(new_n14995_), .A2(new_n14799_), .Z(new_n14996_));
  NOR2_X1    g14932(.A1(new_n14784_), .A2(new_n14801_), .ZN(new_n14997_));
  NOR2_X1    g14933(.A1(new_n14997_), .A2(new_n14798_), .ZN(new_n14998_));
  AOI21_X1   g14934(.A1(new_n14996_), .A2(new_n14798_), .B(new_n14998_), .ZN(new_n14999_));
  AOI22_X1   g14935(.A1(new_n10839_), .A2(new_n4292_), .B1(new_n12936_), .B2(new_n4298_), .ZN(new_n15000_));
  AOI21_X1   g14936(.A1(new_n4469_), .A2(new_n9479_), .B(new_n15000_), .ZN(new_n15001_));
  OR3_X2     g14937(.A1(new_n12975_), .A2(new_n4468_), .A3(new_n15001_), .Z(new_n15002_));
  OR2_X2     g14938(.A1(new_n15002_), .A2(\a[17] ), .Z(new_n15003_));
  NAND2_X1   g14939(.A1(new_n15002_), .A2(\a[17] ), .ZN(new_n15004_));
  NAND3_X1   g14940(.A1(new_n15003_), .A2(new_n14999_), .A3(new_n15004_), .ZN(new_n15005_));
  AOI21_X1   g14941(.A1(new_n15003_), .A2(new_n15004_), .B(new_n14999_), .ZN(new_n15006_));
  AOI21_X1   g14942(.A1(new_n14994_), .A2(new_n15005_), .B(new_n15006_), .ZN(new_n15007_));
  XOR2_X1    g14943(.A1(new_n14806_), .A2(\a[20] ), .Z(new_n15008_));
  NAND2_X1   g14944(.A1(new_n15008_), .A2(new_n14896_), .ZN(new_n15009_));
  NAND2_X1   g14945(.A1(new_n14808_), .A2(new_n14809_), .ZN(new_n15010_));
  NAND2_X1   g14946(.A1(new_n15010_), .A2(new_n14803_), .ZN(new_n15011_));
  NAND2_X1   g14947(.A1(new_n15011_), .A2(new_n15009_), .ZN(new_n15012_));
  AOI21_X1   g14948(.A1(new_n14810_), .A2(new_n14899_), .B(new_n14802_), .ZN(new_n15013_));
  AOI21_X1   g14949(.A1(new_n15012_), .A2(new_n14802_), .B(new_n15013_), .ZN(new_n15014_));
  OAI22_X1   g14950(.A1(new_n9478_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n10846_), .ZN(new_n15015_));
  NAND2_X1   g14951(.A1(new_n10854_), .A2(new_n4469_), .ZN(new_n15016_));
  AOI21_X1   g14952(.A1(new_n15015_), .A2(new_n15016_), .B(new_n4468_), .ZN(new_n15017_));
  NAND2_X1   g14953(.A1(new_n13016_), .A2(new_n15017_), .ZN(new_n15018_));
  XOR2_X1    g14954(.A1(new_n15018_), .A2(new_n3372_), .Z(new_n15019_));
  NOR2_X1    g14955(.A1(new_n15019_), .A2(new_n15014_), .ZN(new_n15020_));
  NAND2_X1   g14956(.A1(new_n15019_), .A2(new_n15014_), .ZN(new_n15021_));
  OAI21_X1   g14957(.A1(new_n15007_), .A2(new_n15020_), .B(new_n15021_), .ZN(new_n15022_));
  XOR2_X1    g14958(.A1(new_n14821_), .A2(new_n14815_), .Z(new_n15023_));
  NOR2_X1    g14959(.A1(new_n15023_), .A2(new_n14812_), .ZN(new_n15024_));
  AOI21_X1   g14960(.A1(new_n14902_), .A2(new_n14823_), .B(new_n14900_), .ZN(new_n15025_));
  OAI22_X1   g14961(.A1(new_n9478_), .A2(new_n4291_), .B1(new_n4297_), .B2(new_n10853_), .ZN(new_n15026_));
  NAND2_X1   g14962(.A1(new_n10862_), .A2(new_n4469_), .ZN(new_n15027_));
  AOI21_X1   g14963(.A1(new_n15026_), .A2(new_n15027_), .B(new_n4468_), .ZN(new_n15028_));
  NAND2_X1   g14964(.A1(new_n13484_), .A2(new_n15028_), .ZN(new_n15029_));
  XOR2_X1    g14965(.A1(new_n15029_), .A2(\a[17] ), .Z(new_n15030_));
  OAI21_X1   g14966(.A1(new_n15024_), .A2(new_n15025_), .B(new_n15030_), .ZN(new_n15031_));
  NOR3_X1    g14967(.A1(new_n15030_), .A2(new_n15024_), .A3(new_n15025_), .ZN(new_n15032_));
  AOI21_X1   g14968(.A1(new_n15022_), .A2(new_n15031_), .B(new_n15032_), .ZN(new_n15033_));
  NAND2_X1   g14969(.A1(new_n14838_), .A2(new_n14839_), .ZN(new_n15034_));
  NOR2_X1    g14970(.A1(new_n15034_), .A2(new_n14831_), .ZN(new_n15035_));
  AOI21_X1   g14971(.A1(new_n14838_), .A2(new_n14839_), .B(new_n14908_), .ZN(new_n15036_));
  OAI21_X1   g14972(.A1(new_n15036_), .A2(new_n15035_), .B(new_n14824_), .ZN(new_n15037_));
  OAI21_X1   g14973(.A1(new_n14910_), .A2(new_n14841_), .B(new_n14904_), .ZN(new_n15038_));
  OAI22_X1   g14974(.A1(new_n10861_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n10853_), .ZN(new_n15039_));
  NAND2_X1   g14975(.A1(new_n8785_), .A2(new_n4469_), .ZN(new_n15040_));
  AOI21_X1   g14976(.A1(new_n15040_), .A2(new_n15039_), .B(new_n4468_), .ZN(new_n15041_));
  NAND2_X1   g14977(.A1(new_n13592_), .A2(new_n15041_), .ZN(new_n15042_));
  XOR2_X1    g14978(.A1(new_n15042_), .A2(new_n3372_), .Z(new_n15043_));
  AOI21_X1   g14979(.A1(new_n15037_), .A2(new_n15038_), .B(new_n15043_), .ZN(new_n15044_));
  NOR2_X1    g14980(.A1(new_n15033_), .A2(new_n15044_), .ZN(new_n15045_));
  NAND2_X1   g14981(.A1(new_n15037_), .A2(new_n15038_), .ZN(new_n15046_));
  XOR2_X1    g14982(.A1(new_n15042_), .A2(\a[17] ), .Z(new_n15047_));
  NOR2_X1    g14983(.A1(new_n15046_), .A2(new_n15047_), .ZN(new_n15048_));
  NOR3_X1    g14984(.A1(new_n15045_), .A2(new_n14942_), .A3(new_n15048_), .ZN(new_n15049_));
  OAI21_X1   g14985(.A1(new_n14923_), .A2(new_n14875_), .B(new_n14857_), .ZN(new_n15050_));
  NAND3_X1   g14986(.A1(new_n14870_), .A2(new_n14862_), .A3(new_n14861_), .ZN(new_n15051_));
  NOR2_X1    g14987(.A1(new_n14860_), .A2(new_n14859_), .ZN(new_n15052_));
  NOR2_X1    g14988(.A1(new_n15052_), .A2(new_n14614_), .ZN(new_n15053_));
  AOI21_X1   g14989(.A1(new_n14241_), .A2(new_n14245_), .B(new_n14224_), .ZN(new_n15054_));
  OAI21_X1   g14990(.A1(new_n15054_), .A2(new_n15053_), .B(new_n14873_), .ZN(new_n15055_));
  NAND2_X1   g14991(.A1(new_n15055_), .A2(new_n15051_), .ZN(new_n15056_));
  NAND2_X1   g14992(.A1(new_n15056_), .A2(new_n14922_), .ZN(new_n15057_));
  AOI22_X1   g14993(.A1(new_n8779_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n8785_), .ZN(new_n15058_));
  NOR2_X1    g14994(.A1(new_n10871_), .A2(new_n4470_), .ZN(new_n15059_));
  OAI21_X1   g14995(.A1(new_n15059_), .A2(new_n15058_), .B(new_n4295_), .ZN(new_n15060_));
  INV_X1     g14996(.I(new_n15060_), .ZN(new_n15061_));
  NAND3_X1   g14997(.A1(new_n11792_), .A2(new_n11793_), .A3(new_n15061_), .ZN(new_n15062_));
  XOR2_X1    g14998(.A1(new_n15062_), .A2(\a[17] ), .Z(new_n15063_));
  NAND3_X1   g14999(.A1(new_n15050_), .A2(new_n15063_), .A3(new_n15057_), .ZN(new_n15064_));
  AOI21_X1   g15000(.A1(new_n14871_), .A2(new_n14874_), .B(new_n14922_), .ZN(new_n15065_));
  AOI21_X1   g15001(.A1(new_n15051_), .A2(new_n15055_), .B(new_n14857_), .ZN(new_n15066_));
  NAND2_X1   g15002(.A1(new_n12809_), .A2(new_n8779_), .ZN(new_n15067_));
  AOI21_X1   g15003(.A1(new_n15067_), .A2(new_n11786_), .B(new_n10871_), .ZN(new_n15068_));
  INV_X1     g15004(.I(new_n11793_), .ZN(new_n15069_));
  NOR2_X1    g15005(.A1(new_n15069_), .A2(new_n15068_), .ZN(new_n15070_));
  NAND3_X1   g15006(.A1(new_n15070_), .A2(new_n3372_), .A3(new_n15061_), .ZN(new_n15071_));
  NAND2_X1   g15007(.A1(new_n15062_), .A2(\a[17] ), .ZN(new_n15072_));
  NAND2_X1   g15008(.A1(new_n15071_), .A2(new_n15072_), .ZN(new_n15073_));
  OAI21_X1   g15009(.A1(new_n15066_), .A2(new_n15065_), .B(new_n15073_), .ZN(new_n15074_));
  NAND3_X1   g15010(.A1(new_n15074_), .A2(new_n15064_), .A3(new_n14942_), .ZN(new_n15075_));
  NOR2_X1    g15011(.A1(new_n15075_), .A2(new_n15049_), .ZN(new_n15076_));
  XOR2_X1    g15012(.A1(new_n14776_), .A2(new_n3372_), .Z(new_n15077_));
  NOR2_X1    g15013(.A1(new_n14892_), .A2(new_n14888_), .ZN(new_n15078_));
  NOR2_X1    g15014(.A1(new_n14881_), .A2(new_n14889_), .ZN(new_n15079_));
  OAI21_X1   g15015(.A1(new_n15079_), .A2(new_n15078_), .B(new_n14924_), .ZN(new_n15080_));
  NOR2_X1    g15016(.A1(new_n14881_), .A2(new_n14888_), .ZN(new_n15081_));
  NOR2_X1    g15017(.A1(new_n14892_), .A2(new_n14889_), .ZN(new_n15082_));
  OAI21_X1   g15018(.A1(new_n15081_), .A2(new_n15082_), .B(new_n14876_), .ZN(new_n15083_));
  NAND3_X1   g15019(.A1(new_n15080_), .A2(new_n15083_), .A3(new_n15077_), .ZN(new_n15084_));
  OAI21_X1   g15020(.A1(new_n14894_), .A2(new_n14927_), .B(new_n14777_), .ZN(new_n15085_));
  NOR3_X1    g15021(.A1(new_n15066_), .A2(new_n15065_), .A3(new_n15073_), .ZN(new_n15086_));
  AOI21_X1   g15022(.A1(new_n15085_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n15087_));
  AOI21_X1   g15023(.A1(new_n15087_), .A2(new_n15076_), .B(new_n14929_), .ZN(new_n15088_));
  NAND2_X1   g15024(.A1(new_n14890_), .A2(new_n14924_), .ZN(new_n15089_));
  NAND2_X1   g15025(.A1(new_n15089_), .A2(new_n14893_), .ZN(new_n15090_));
  OAI22_X1   g15026(.A1(new_n8784_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n10861_), .ZN(new_n15091_));
  NAND2_X1   g15027(.A1(new_n8779_), .A2(new_n4096_), .ZN(new_n15092_));
  AOI21_X1   g15028(.A1(new_n15092_), .A2(new_n15091_), .B(new_n4095_), .ZN(new_n15093_));
  NAND3_X1   g15029(.A1(new_n12814_), .A2(new_n3035_), .A3(new_n15093_), .ZN(new_n15094_));
  AOI21_X1   g15030(.A1(new_n12814_), .A2(new_n15093_), .B(new_n3035_), .ZN(new_n15095_));
  INV_X1     g15031(.I(new_n15095_), .ZN(new_n15096_));
  NAND2_X1   g15032(.A1(new_n15096_), .A2(new_n15094_), .ZN(new_n15097_));
  NOR2_X1    g15033(.A1(new_n14274_), .A2(new_n14622_), .ZN(new_n15098_));
  NOR2_X1    g15034(.A1(new_n14281_), .A2(new_n14620_), .ZN(new_n15099_));
  OAI21_X1   g15035(.A1(new_n15098_), .A2(new_n15099_), .B(new_n14268_), .ZN(new_n15100_));
  OAI21_X1   g15036(.A1(new_n14283_), .A2(new_n14623_), .B(new_n14618_), .ZN(new_n15101_));
  NAND2_X1   g15037(.A1(new_n15100_), .A2(new_n15101_), .ZN(new_n15102_));
  NOR2_X1    g15038(.A1(new_n15102_), .A2(new_n15097_), .ZN(new_n15103_));
  INV_X1     g15039(.I(new_n15094_), .ZN(new_n15104_));
  NOR2_X1    g15040(.A1(new_n15104_), .A2(new_n15095_), .ZN(new_n15105_));
  NAND2_X1   g15041(.A1(new_n14281_), .A2(new_n14620_), .ZN(new_n15106_));
  NAND2_X1   g15042(.A1(new_n14274_), .A2(new_n14622_), .ZN(new_n15107_));
  AOI21_X1   g15043(.A1(new_n15107_), .A2(new_n15106_), .B(new_n14618_), .ZN(new_n15108_));
  AOI21_X1   g15044(.A1(new_n14282_), .A2(new_n14624_), .B(new_n14268_), .ZN(new_n15109_));
  NOR2_X1    g15045(.A1(new_n15109_), .A2(new_n15108_), .ZN(new_n15110_));
  NOR2_X1    g15046(.A1(new_n15110_), .A2(new_n15105_), .ZN(new_n15111_));
  OAI21_X1   g15047(.A1(new_n15103_), .A2(new_n15111_), .B(new_n15090_), .ZN(new_n15112_));
  NOR2_X1    g15048(.A1(new_n15078_), .A2(new_n14876_), .ZN(new_n15113_));
  NOR2_X1    g15049(.A1(new_n15113_), .A2(new_n15079_), .ZN(new_n15114_));
  NAND2_X1   g15050(.A1(new_n15102_), .A2(new_n15105_), .ZN(new_n15115_));
  NAND2_X1   g15051(.A1(new_n15110_), .A2(new_n15097_), .ZN(new_n15116_));
  NAND2_X1   g15052(.A1(new_n15116_), .A2(new_n15115_), .ZN(new_n15117_));
  NAND2_X1   g15053(.A1(new_n15117_), .A2(new_n15114_), .ZN(new_n15118_));
  AOI22_X1   g15054(.A1(new_n10886_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n10872_), .ZN(new_n15119_));
  NOR2_X1    g15055(.A1(new_n10892_), .A2(new_n4470_), .ZN(new_n15120_));
  NOR2_X1    g15056(.A1(new_n15119_), .A2(new_n15120_), .ZN(new_n15121_));
  NOR4_X1    g15057(.A1(new_n14669_), .A2(new_n12774_), .A3(new_n4468_), .A4(new_n15121_), .ZN(new_n15122_));
  XOR2_X1    g15058(.A1(new_n15122_), .A2(\a[17] ), .Z(new_n15123_));
  AOI21_X1   g15059(.A1(new_n15118_), .A2(new_n15112_), .B(new_n15123_), .ZN(new_n15124_));
  NAND3_X1   g15060(.A1(new_n15123_), .A2(new_n15112_), .A3(new_n15118_), .ZN(new_n15125_));
  OAI21_X1   g15061(.A1(new_n15088_), .A2(new_n15124_), .B(new_n15125_), .ZN(new_n15126_));
  OAI21_X1   g15062(.A1(new_n14300_), .A2(new_n14626_), .B(new_n14625_), .ZN(new_n15127_));
  NAND3_X1   g15063(.A1(new_n14298_), .A2(new_n14288_), .A3(new_n14290_), .ZN(new_n15128_));
  INV_X1     g15064(.I(new_n14287_), .ZN(new_n15129_));
  AOI22_X1   g15065(.A1(new_n15129_), .A2(new_n14285_), .B1(new_n14156_), .B2(new_n14157_), .ZN(new_n15130_));
  AOI21_X1   g15066(.A1(new_n14163_), .A2(new_n14095_), .B(new_n14158_), .ZN(new_n15131_));
  OAI21_X1   g15067(.A1(new_n15131_), .A2(new_n15130_), .B(new_n14302_), .ZN(new_n15132_));
  NAND2_X1   g15068(.A1(new_n15132_), .A2(new_n15128_), .ZN(new_n15133_));
  NAND2_X1   g15069(.A1(new_n14284_), .A2(new_n15133_), .ZN(new_n15134_));
  AOI22_X1   g15070(.A1(new_n8779_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n8785_), .ZN(new_n15135_));
  NOR2_X1    g15071(.A1(new_n10871_), .A2(new_n4097_), .ZN(new_n15136_));
  OAI21_X1   g15072(.A1(new_n15136_), .A2(new_n15135_), .B(new_n3773_), .ZN(new_n15137_));
  INV_X1     g15073(.I(new_n15137_), .ZN(new_n15138_));
  NAND4_X1   g15074(.A1(new_n11792_), .A2(new_n11793_), .A3(new_n3035_), .A4(new_n15138_), .ZN(new_n15139_));
  INV_X1     g15075(.I(new_n15139_), .ZN(new_n15140_));
  AOI21_X1   g15076(.A1(new_n15070_), .A2(new_n15138_), .B(new_n3035_), .ZN(new_n15141_));
  NOR2_X1    g15077(.A1(new_n15141_), .A2(new_n15140_), .ZN(new_n15142_));
  NAND3_X1   g15078(.A1(new_n15127_), .A2(new_n15134_), .A3(new_n15142_), .ZN(new_n15143_));
  NAND2_X1   g15079(.A1(new_n14268_), .A2(new_n14282_), .ZN(new_n15144_));
  AOI22_X1   g15080(.A1(new_n15144_), .A2(new_n14624_), .B1(new_n14299_), .B2(new_n14303_), .ZN(new_n15145_));
  NOR3_X1    g15081(.A1(new_n15131_), .A2(new_n14302_), .A3(new_n15130_), .ZN(new_n15146_));
  AOI22_X1   g15082(.A1(new_n14288_), .A2(new_n14290_), .B1(new_n14295_), .B2(new_n14301_), .ZN(new_n15147_));
  NOR2_X1    g15083(.A1(new_n15146_), .A2(new_n15147_), .ZN(new_n15148_));
  NOR2_X1    g15084(.A1(new_n15148_), .A2(new_n14625_), .ZN(new_n15149_));
  OAI21_X1   g15085(.A1(new_n11794_), .A2(new_n15137_), .B(\a[20] ), .ZN(new_n15150_));
  NAND2_X1   g15086(.A1(new_n15150_), .A2(new_n15139_), .ZN(new_n15151_));
  OAI21_X1   g15087(.A1(new_n15145_), .A2(new_n15149_), .B(new_n15151_), .ZN(new_n15152_));
  NAND2_X1   g15088(.A1(new_n15143_), .A2(new_n15152_), .ZN(new_n15153_));
  OAI21_X1   g15089(.A1(new_n15090_), .A2(new_n15110_), .B(new_n15097_), .ZN(new_n15154_));
  NOR2_X1    g15090(.A1(new_n15154_), .A2(new_n15153_), .ZN(new_n15155_));
  NAND2_X1   g15091(.A1(new_n15114_), .A2(new_n15102_), .ZN(new_n15156_));
  AOI22_X1   g15092(.A1(new_n15156_), .A2(new_n15097_), .B1(new_n15143_), .B2(new_n15152_), .ZN(new_n15157_));
  AOI22_X1   g15093(.A1(new_n10886_), .A2(new_n4292_), .B1(new_n10889_), .B2(new_n4298_), .ZN(new_n15158_));
  NOR2_X1    g15094(.A1(new_n10899_), .A2(new_n4470_), .ZN(new_n15159_));
  OR2_X2     g15095(.A1(new_n15159_), .A2(new_n15158_), .Z(new_n15160_));
  NAND4_X1   g15096(.A1(new_n11903_), .A2(new_n11907_), .A3(new_n4295_), .A4(new_n15160_), .ZN(new_n15161_));
  XOR2_X1    g15097(.A1(new_n15161_), .A2(\a[17] ), .Z(new_n15162_));
  OAI21_X1   g15098(.A1(new_n15155_), .A2(new_n15157_), .B(new_n15162_), .ZN(new_n15163_));
  NOR3_X1    g15099(.A1(new_n15162_), .A2(new_n15157_), .A3(new_n15155_), .ZN(new_n15164_));
  AOI21_X1   g15100(.A1(new_n15126_), .A2(new_n15163_), .B(new_n15164_), .ZN(new_n15165_));
  AOI22_X1   g15101(.A1(new_n11899_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n10889_), .ZN(new_n15166_));
  NOR2_X1    g15102(.A1(new_n8774_), .A2(new_n4470_), .ZN(new_n15167_));
  OAI21_X1   g15103(.A1(new_n15167_), .A2(new_n15166_), .B(new_n4295_), .ZN(new_n15168_));
  NOR4_X1    g15104(.A1(new_n14658_), .A2(\a[17] ), .A3(new_n11942_), .A4(new_n15168_), .ZN(new_n15169_));
  NOR2_X1    g15105(.A1(new_n14658_), .A2(new_n11942_), .ZN(new_n15170_));
  INV_X1     g15106(.I(new_n15168_), .ZN(new_n15171_));
  AOI21_X1   g15107(.A1(new_n15170_), .A2(new_n15171_), .B(new_n3372_), .ZN(new_n15172_));
  NOR2_X1    g15108(.A1(new_n15172_), .A2(new_n15169_), .ZN(new_n15173_));
  XOR2_X1    g15109(.A1(new_n14628_), .A2(new_n14629_), .Z(new_n15174_));
  OAI21_X1   g15110(.A1(new_n14630_), .A2(new_n14315_), .B(new_n14627_), .ZN(new_n15175_));
  INV_X1     g15111(.I(new_n15175_), .ZN(new_n15176_));
  AOI21_X1   g15112(.A1(new_n14304_), .A2(new_n15174_), .B(new_n15176_), .ZN(new_n15177_));
  NOR2_X1    g15113(.A1(new_n15110_), .A2(new_n15097_), .ZN(new_n15178_));
  NAND3_X1   g15114(.A1(new_n15178_), .A2(new_n15089_), .A3(new_n14893_), .ZN(new_n15179_));
  NOR3_X1    g15115(.A1(new_n15145_), .A2(new_n15149_), .A3(new_n15151_), .ZN(new_n15180_));
  AOI21_X1   g15116(.A1(new_n15127_), .A2(new_n15134_), .B(new_n15142_), .ZN(new_n15181_));
  NOR3_X1    g15117(.A1(new_n15181_), .A2(new_n15180_), .A3(new_n15178_), .ZN(new_n15182_));
  OAI22_X1   g15118(.A1(new_n10871_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n8778_), .ZN(new_n15183_));
  NAND2_X1   g15119(.A1(new_n10886_), .A2(new_n4096_), .ZN(new_n15184_));
  AOI21_X1   g15120(.A1(new_n15184_), .A2(new_n15183_), .B(new_n4095_), .ZN(new_n15185_));
  NAND2_X1   g15121(.A1(new_n13103_), .A2(new_n15185_), .ZN(new_n15186_));
  XOR2_X1    g15122(.A1(new_n15186_), .A2(new_n3035_), .Z(new_n15187_));
  AOI21_X1   g15123(.A1(new_n15182_), .A2(new_n15179_), .B(new_n15187_), .ZN(new_n15188_));
  NOR3_X1    g15124(.A1(new_n15113_), .A2(new_n15115_), .A3(new_n15079_), .ZN(new_n15189_));
  NAND3_X1   g15125(.A1(new_n15143_), .A2(new_n15152_), .A3(new_n15115_), .ZN(new_n15190_));
  XOR2_X1    g15126(.A1(new_n15186_), .A2(\a[20] ), .Z(new_n15191_));
  NOR3_X1    g15127(.A1(new_n15190_), .A2(new_n15189_), .A3(new_n15191_), .ZN(new_n15192_));
  OAI21_X1   g15128(.A1(new_n15188_), .A2(new_n15192_), .B(new_n15177_), .ZN(new_n15193_));
  NAND2_X1   g15129(.A1(new_n15174_), .A2(new_n14304_), .ZN(new_n15194_));
  NAND2_X1   g15130(.A1(new_n15194_), .A2(new_n15175_), .ZN(new_n15195_));
  OAI21_X1   g15131(.A1(new_n15190_), .A2(new_n15189_), .B(new_n15191_), .ZN(new_n15196_));
  NAND3_X1   g15132(.A1(new_n15182_), .A2(new_n15179_), .A3(new_n15187_), .ZN(new_n15197_));
  NAND3_X1   g15133(.A1(new_n15197_), .A2(new_n15196_), .A3(new_n15195_), .ZN(new_n15198_));
  NAND3_X1   g15134(.A1(new_n15193_), .A2(new_n15198_), .A3(new_n15173_), .ZN(new_n15199_));
  INV_X1     g15135(.I(new_n15169_), .ZN(new_n15200_));
  OAI21_X1   g15136(.A1(new_n11945_), .A2(new_n15168_), .B(\a[17] ), .ZN(new_n15201_));
  NAND2_X1   g15137(.A1(new_n15201_), .A2(new_n15200_), .ZN(new_n15202_));
  AOI21_X1   g15138(.A1(new_n15197_), .A2(new_n15196_), .B(new_n15195_), .ZN(new_n15203_));
  NOR3_X1    g15139(.A1(new_n15188_), .A2(new_n15192_), .A3(new_n15177_), .ZN(new_n15204_));
  OAI21_X1   g15140(.A1(new_n15203_), .A2(new_n15204_), .B(new_n15202_), .ZN(new_n15205_));
  NAND2_X1   g15141(.A1(new_n15205_), .A2(new_n15199_), .ZN(new_n15206_));
  NAND2_X1   g15142(.A1(new_n15165_), .A2(new_n15206_), .ZN(new_n15207_));
  NOR2_X1    g15143(.A1(new_n14758_), .A2(\a[17] ), .ZN(new_n15208_));
  AOI21_X1   g15144(.A1(new_n12001_), .A2(new_n14751_), .B(new_n3372_), .ZN(new_n15209_));
  NOR2_X1    g15145(.A1(new_n15208_), .A2(new_n15209_), .ZN(new_n15210_));
  NOR3_X1    g15146(.A1(new_n15210_), .A2(new_n14768_), .A3(new_n14765_), .ZN(new_n15211_));
  OAI21_X1   g15147(.A1(new_n14767_), .A2(new_n14766_), .B(new_n14673_), .ZN(new_n15212_));
  NAND3_X1   g15148(.A1(new_n14764_), .A2(new_n14763_), .A3(new_n14633_), .ZN(new_n15213_));
  AOI21_X1   g15149(.A1(new_n15213_), .A2(new_n15212_), .B(new_n14760_), .ZN(new_n15214_));
  NOR2_X1    g15150(.A1(new_n15214_), .A2(new_n15211_), .ZN(new_n15215_));
  OAI21_X1   g15151(.A1(new_n15203_), .A2(new_n15204_), .B(new_n15173_), .ZN(new_n15216_));
  INV_X1     g15152(.I(new_n15216_), .ZN(new_n15217_));
  NOR2_X1    g15153(.A1(new_n15215_), .A2(new_n15217_), .ZN(new_n15218_));
  AOI21_X1   g15154(.A1(new_n15207_), .A2(new_n15218_), .B(new_n14770_), .ZN(new_n15219_));
  OAI21_X1   g15155(.A1(new_n14742_), .A2(new_n14739_), .B(new_n14747_), .ZN(new_n15220_));
  AOI21_X1   g15156(.A1(new_n15219_), .A2(new_n15220_), .B(new_n14748_), .ZN(new_n15221_));
  NOR3_X1    g15157(.A1(new_n15221_), .A2(new_n14735_), .A3(new_n14738_), .ZN(new_n15222_));
  OAI22_X1   g15158(.A1(new_n14727_), .A2(new_n14723_), .B1(new_n14599_), .B2(new_n15222_), .ZN(new_n15223_));
  AOI21_X1   g15159(.A1(new_n15223_), .A2(new_n14594_), .B(new_n14591_), .ZN(new_n15224_));
  NOR2_X1    g15160(.A1(new_n15224_), .A2(new_n14581_), .ZN(new_n15225_));
  NAND3_X1   g15161(.A1(new_n14568_), .A2(new_n14576_), .A3(new_n15225_), .ZN(new_n15226_));
  AOI21_X1   g15162(.A1(new_n15226_), .A2(new_n14563_), .B(new_n14485_), .ZN(new_n15227_));
  INV_X1     g15163(.I(new_n14485_), .ZN(new_n15228_));
  INV_X1     g15164(.I(new_n15225_), .ZN(new_n15229_));
  NOR3_X1    g15165(.A1(new_n14565_), .A2(new_n14566_), .A3(new_n14491_), .ZN(new_n15230_));
  AOI21_X1   g15166(.A1(new_n14555_), .A2(new_n14561_), .B(new_n14490_), .ZN(new_n15231_));
  OAI21_X1   g15167(.A1(new_n15230_), .A2(new_n15231_), .B(new_n14576_), .ZN(new_n15232_));
  OAI21_X1   g15168(.A1(new_n15232_), .A2(new_n15229_), .B(new_n14563_), .ZN(new_n15233_));
  NOR2_X1    g15169(.A1(new_n15233_), .A2(new_n15228_), .ZN(new_n15234_));
  OAI22_X1   g15170(.A1(new_n6094_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n6089_), .ZN(new_n15235_));
  NAND2_X1   g15171(.A1(new_n8696_), .A2(new_n6090_), .ZN(new_n15236_));
  AOI21_X1   g15172(.A1(new_n15235_), .A2(new_n15236_), .B(new_n6082_), .ZN(new_n15237_));
  NAND2_X1   g15173(.A1(new_n11595_), .A2(new_n15237_), .ZN(new_n15238_));
  XOR2_X1    g15174(.A1(new_n15238_), .A2(\a[14] ), .Z(new_n15239_));
  INV_X1     g15175(.I(new_n15239_), .ZN(new_n15240_));
  NOR3_X1    g15176(.A1(new_n15234_), .A2(new_n15227_), .A3(new_n15240_), .ZN(new_n15241_));
  NAND2_X1   g15177(.A1(new_n15233_), .A2(new_n15228_), .ZN(new_n15242_));
  NAND3_X1   g15178(.A1(new_n15226_), .A2(new_n14485_), .A3(new_n14563_), .ZN(new_n15243_));
  AOI21_X1   g15179(.A1(new_n15242_), .A2(new_n15243_), .B(new_n15239_), .ZN(new_n15244_));
  OAI22_X1   g15180(.A1(new_n4716_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n4719_), .ZN(new_n15245_));
  NAND2_X1   g15181(.A1(new_n8674_), .A2(new_n4709_), .ZN(new_n15246_));
  AOI21_X1   g15182(.A1(new_n15246_), .A2(new_n15245_), .B(new_n4707_), .ZN(new_n15247_));
  NAND2_X1   g15183(.A1(new_n11431_), .A2(new_n15247_), .ZN(new_n15248_));
  XOR2_X1    g15184(.A1(new_n15248_), .A2(new_n4034_), .Z(new_n15249_));
  NOR3_X1    g15185(.A1(new_n15249_), .A2(new_n15244_), .A3(new_n15241_), .ZN(new_n15250_));
  INV_X1     g15186(.I(new_n15250_), .ZN(new_n15251_));
  OAI21_X1   g15187(.A1(new_n15241_), .A2(new_n15244_), .B(new_n15249_), .ZN(new_n15252_));
  AND2_X2    g15188(.A1(new_n15251_), .A2(new_n15252_), .Z(new_n15253_));
  OAI22_X1   g15189(.A1(new_n8681_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8694_), .ZN(new_n15254_));
  NAND2_X1   g15190(.A1(new_n8688_), .A2(new_n4709_), .ZN(new_n15255_));
  AOI21_X1   g15191(.A1(new_n15255_), .A2(new_n15254_), .B(new_n4707_), .ZN(new_n15256_));
  NAND2_X1   g15192(.A1(new_n11420_), .A2(new_n15256_), .ZN(new_n15257_));
  XOR2_X1    g15193(.A1(new_n15257_), .A2(\a[11] ), .Z(new_n15258_));
  INV_X1     g15194(.I(new_n14562_), .ZN(new_n15259_));
  AOI21_X1   g15195(.A1(new_n15225_), .A2(new_n14576_), .B(new_n14490_), .ZN(new_n15260_));
  NAND2_X1   g15196(.A1(new_n14590_), .A2(new_n14594_), .ZN(new_n15261_));
  NAND3_X1   g15197(.A1(new_n14725_), .A2(new_n14726_), .A3(new_n14724_), .ZN(new_n15262_));
  OAI21_X1   g15198(.A1(new_n14722_), .A2(new_n14719_), .B(new_n14599_), .ZN(new_n15263_));
  INV_X1     g15199(.I(new_n14735_), .ZN(new_n15264_));
  INV_X1     g15200(.I(new_n14738_), .ZN(new_n15265_));
  NOR3_X1    g15201(.A1(new_n14712_), .A2(new_n14713_), .A3(new_n14714_), .ZN(new_n15266_));
  OAI21_X1   g15202(.A1(new_n15266_), .A2(new_n14693_), .B(new_n14711_), .ZN(new_n15267_));
  NOR3_X1    g15203(.A1(new_n14712_), .A2(new_n14713_), .A3(new_n14692_), .ZN(new_n15268_));
  AOI21_X1   g15204(.A1(new_n14682_), .A2(new_n14686_), .B(new_n14714_), .ZN(new_n15269_));
  OAI21_X1   g15205(.A1(new_n15268_), .A2(new_n15269_), .B(new_n14677_), .ZN(new_n15270_));
  XOR2_X1    g15206(.A1(new_n14746_), .A2(new_n3372_), .Z(new_n15271_));
  NAND3_X1   g15207(.A1(new_n15267_), .A2(new_n15270_), .A3(new_n15271_), .ZN(new_n15272_));
  INV_X1     g15208(.I(new_n14770_), .ZN(new_n15273_));
  INV_X1     g15209(.I(new_n14935_), .ZN(new_n15274_));
  AOI21_X1   g15210(.A1(new_n14936_), .A2(new_n14937_), .B(new_n14842_), .ZN(new_n15275_));
  AOI21_X1   g15211(.A1(new_n14920_), .A2(new_n14856_), .B(new_n14912_), .ZN(new_n15276_));
  NOR2_X1    g15212(.A1(new_n15275_), .A2(new_n15276_), .ZN(new_n15277_));
  NOR2_X1    g15213(.A1(new_n15274_), .A2(new_n15277_), .ZN(new_n15278_));
  NOR2_X1    g15214(.A1(new_n14966_), .A2(new_n14797_), .ZN(new_n15279_));
  AOI21_X1   g15215(.A1(new_n14964_), .A2(new_n14967_), .B(new_n15279_), .ZN(new_n15280_));
  XNOR2_X1   g15216(.A1(new_n14970_), .A2(new_n14971_), .ZN(new_n15281_));
  XOR2_X1    g15217(.A1(new_n14975_), .A2(new_n3372_), .Z(new_n15282_));
  NOR2_X1    g15218(.A1(new_n15282_), .A2(new_n15281_), .ZN(new_n15283_));
  NAND2_X1   g15219(.A1(new_n15282_), .A2(new_n15281_), .ZN(new_n15284_));
  OAI21_X1   g15220(.A1(new_n15280_), .A2(new_n15283_), .B(new_n15284_), .ZN(new_n15285_));
  INV_X1     g15221(.I(new_n14985_), .ZN(new_n15286_));
  NAND2_X1   g15222(.A1(new_n15286_), .A2(new_n14990_), .ZN(new_n15287_));
  NOR2_X1    g15223(.A1(new_n15286_), .A2(new_n14990_), .ZN(new_n15288_));
  AOI21_X1   g15224(.A1(new_n15285_), .A2(new_n15287_), .B(new_n15288_), .ZN(new_n15289_));
  INV_X1     g15225(.I(new_n15005_), .ZN(new_n15290_));
  INV_X1     g15226(.I(new_n14999_), .ZN(new_n15291_));
  XOR2_X1    g15227(.A1(new_n15002_), .A2(new_n3372_), .Z(new_n15292_));
  NAND2_X1   g15228(.A1(new_n15292_), .A2(new_n15291_), .ZN(new_n15293_));
  OAI21_X1   g15229(.A1(new_n15290_), .A2(new_n15289_), .B(new_n15293_), .ZN(new_n15294_));
  NOR2_X1    g15230(.A1(new_n15010_), .A2(new_n14803_), .ZN(new_n15295_));
  NOR2_X1    g15231(.A1(new_n15008_), .A2(new_n14896_), .ZN(new_n15296_));
  OAI21_X1   g15232(.A1(new_n15295_), .A2(new_n15296_), .B(new_n14802_), .ZN(new_n15297_));
  OAI21_X1   g15233(.A1(new_n14898_), .A2(new_n14811_), .B(new_n14895_), .ZN(new_n15298_));
  NAND2_X1   g15234(.A1(new_n15297_), .A2(new_n15298_), .ZN(new_n15299_));
  XOR2_X1    g15235(.A1(new_n15018_), .A2(\a[17] ), .Z(new_n15300_));
  NAND2_X1   g15236(.A1(new_n15300_), .A2(new_n15299_), .ZN(new_n15301_));
  NOR2_X1    g15237(.A1(new_n15300_), .A2(new_n15299_), .ZN(new_n15302_));
  AOI21_X1   g15238(.A1(new_n15294_), .A2(new_n15301_), .B(new_n15302_), .ZN(new_n15303_));
  INV_X1     g15239(.I(new_n15031_), .ZN(new_n15304_));
  INV_X1     g15240(.I(new_n15032_), .ZN(new_n15305_));
  OAI21_X1   g15241(.A1(new_n15303_), .A2(new_n15304_), .B(new_n15305_), .ZN(new_n15306_));
  NAND2_X1   g15242(.A1(new_n15046_), .A2(new_n15047_), .ZN(new_n15307_));
  NAND2_X1   g15243(.A1(new_n15306_), .A2(new_n15307_), .ZN(new_n15308_));
  INV_X1     g15244(.I(new_n15048_), .ZN(new_n15309_));
  NAND3_X1   g15245(.A1(new_n15308_), .A2(new_n15278_), .A3(new_n15309_), .ZN(new_n15310_));
  AOI21_X1   g15246(.A1(new_n15050_), .A2(new_n15057_), .B(new_n15063_), .ZN(new_n15311_));
  NOR2_X1    g15247(.A1(new_n15311_), .A2(new_n15086_), .ZN(new_n15312_));
  NAND3_X1   g15248(.A1(new_n15310_), .A2(new_n15312_), .A3(new_n14942_), .ZN(new_n15313_));
  NOR3_X1    g15249(.A1(new_n14894_), .A2(new_n14927_), .A3(new_n14777_), .ZN(new_n15314_));
  AOI21_X1   g15250(.A1(new_n15083_), .A2(new_n15080_), .B(new_n15077_), .ZN(new_n15315_));
  OAI21_X1   g15251(.A1(new_n15314_), .A2(new_n15315_), .B(new_n15064_), .ZN(new_n15316_));
  OAI21_X1   g15252(.A1(new_n15316_), .A2(new_n15313_), .B(new_n14928_), .ZN(new_n15317_));
  NOR2_X1    g15253(.A1(new_n15111_), .A2(new_n15103_), .ZN(new_n15318_));
  NOR2_X1    g15254(.A1(new_n15318_), .A2(new_n15114_), .ZN(new_n15319_));
  AOI21_X1   g15255(.A1(new_n15115_), .A2(new_n15116_), .B(new_n15090_), .ZN(new_n15320_));
  XOR2_X1    g15256(.A1(new_n15122_), .A2(new_n3372_), .Z(new_n15321_));
  OAI21_X1   g15257(.A1(new_n15320_), .A2(new_n15319_), .B(new_n15321_), .ZN(new_n15322_));
  NOR3_X1    g15258(.A1(new_n15321_), .A2(new_n15320_), .A3(new_n15319_), .ZN(new_n15323_));
  AOI21_X1   g15259(.A1(new_n15317_), .A2(new_n15322_), .B(new_n15323_), .ZN(new_n15324_));
  INV_X1     g15260(.I(new_n15155_), .ZN(new_n15325_));
  NAND2_X1   g15261(.A1(new_n15154_), .A2(new_n15153_), .ZN(new_n15326_));
  XOR2_X1    g15262(.A1(new_n15161_), .A2(new_n3372_), .Z(new_n15327_));
  AOI21_X1   g15263(.A1(new_n15325_), .A2(new_n15326_), .B(new_n15327_), .ZN(new_n15328_));
  NAND3_X1   g15264(.A1(new_n15325_), .A2(new_n15326_), .A3(new_n15327_), .ZN(new_n15329_));
  OAI21_X1   g15265(.A1(new_n15324_), .A2(new_n15328_), .B(new_n15329_), .ZN(new_n15330_));
  NOR3_X1    g15266(.A1(new_n15203_), .A2(new_n15204_), .A3(new_n15202_), .ZN(new_n15331_));
  AOI21_X1   g15267(.A1(new_n15193_), .A2(new_n15198_), .B(new_n15173_), .ZN(new_n15332_));
  NOR2_X1    g15268(.A1(new_n15331_), .A2(new_n15332_), .ZN(new_n15333_));
  NOR2_X1    g15269(.A1(new_n15330_), .A2(new_n15333_), .ZN(new_n15334_));
  OAI21_X1   g15270(.A1(new_n15211_), .A2(new_n15214_), .B(new_n15216_), .ZN(new_n15335_));
  OAI21_X1   g15271(.A1(new_n15334_), .A2(new_n15335_), .B(new_n15273_), .ZN(new_n15336_));
  AOI21_X1   g15272(.A1(new_n15267_), .A2(new_n15270_), .B(new_n15271_), .ZN(new_n15337_));
  OAI21_X1   g15273(.A1(new_n15336_), .A2(new_n15337_), .B(new_n15272_), .ZN(new_n15338_));
  NAND3_X1   g15274(.A1(new_n15338_), .A2(new_n15264_), .A3(new_n15265_), .ZN(new_n15339_));
  AOI22_X1   g15275(.A1(new_n15263_), .A2(new_n15262_), .B1(new_n15339_), .B2(new_n14724_), .ZN(new_n15340_));
  OAI21_X1   g15276(.A1(new_n15340_), .A2(new_n15261_), .B(new_n14590_), .ZN(new_n15341_));
  NAND3_X1   g15277(.A1(new_n15341_), .A2(new_n14576_), .A3(new_n14580_), .ZN(new_n15342_));
  NOR2_X1    g15278(.A1(new_n15342_), .A2(new_n14491_), .ZN(new_n15343_));
  OAI21_X1   g15279(.A1(new_n15260_), .A2(new_n15343_), .B(new_n15259_), .ZN(new_n15344_));
  NAND2_X1   g15280(.A1(new_n15342_), .A2(new_n14491_), .ZN(new_n15345_));
  NAND3_X1   g15281(.A1(new_n15225_), .A2(new_n14490_), .A3(new_n14576_), .ZN(new_n15346_));
  NAND3_X1   g15282(.A1(new_n15346_), .A2(new_n15345_), .A3(new_n14562_), .ZN(new_n15347_));
  NAND2_X1   g15283(.A1(new_n15344_), .A2(new_n15347_), .ZN(new_n15348_));
  OAI22_X1   g15284(.A1(new_n8710_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8718_), .ZN(new_n15349_));
  NAND2_X1   g15285(.A1(new_n8702_), .A2(new_n6090_), .ZN(new_n15350_));
  AOI21_X1   g15286(.A1(new_n15350_), .A2(new_n15349_), .B(new_n6082_), .ZN(new_n15351_));
  NAND2_X1   g15287(.A1(new_n12205_), .A2(new_n15351_), .ZN(new_n15352_));
  XOR2_X1    g15288(.A1(new_n15352_), .A2(\a[14] ), .Z(new_n15353_));
  NOR2_X1    g15289(.A1(new_n15341_), .A2(new_n14581_), .ZN(new_n15354_));
  NOR3_X1    g15290(.A1(new_n14578_), .A2(new_n14577_), .A3(new_n14579_), .ZN(new_n15355_));
  AOI21_X1   g15291(.A1(new_n14570_), .A2(new_n14569_), .B(new_n14575_), .ZN(new_n15356_));
  NOR2_X1    g15292(.A1(new_n15355_), .A2(new_n15356_), .ZN(new_n15357_));
  NOR2_X1    g15293(.A1(new_n15224_), .A2(new_n15357_), .ZN(new_n15358_));
  OAI22_X1   g15294(.A1(new_n8725_), .A2(new_n6089_), .B1(new_n6094_), .B2(new_n8718_), .ZN(new_n15359_));
  NAND2_X1   g15295(.A1(new_n8711_), .A2(new_n6090_), .ZN(new_n15360_));
  AOI21_X1   g15296(.A1(new_n15360_), .A2(new_n15359_), .B(new_n6082_), .ZN(new_n15361_));
  NAND2_X1   g15297(.A1(new_n11536_), .A2(new_n15361_), .ZN(new_n15362_));
  XOR2_X1    g15298(.A1(new_n15362_), .A2(\a[14] ), .Z(new_n15363_));
  OAI21_X1   g15299(.A1(new_n15358_), .A2(new_n15354_), .B(new_n15363_), .ZN(new_n15364_));
  NAND2_X1   g15300(.A1(new_n15224_), .A2(new_n15357_), .ZN(new_n15365_));
  NAND2_X1   g15301(.A1(new_n15341_), .A2(new_n14581_), .ZN(new_n15366_));
  XOR2_X1    g15302(.A1(new_n15362_), .A2(new_n3521_), .Z(new_n15367_));
  NAND3_X1   g15303(.A1(new_n15365_), .A2(new_n15366_), .A3(new_n15367_), .ZN(new_n15368_));
  OAI22_X1   g15304(.A1(new_n8725_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8735_), .ZN(new_n15369_));
  NAND2_X1   g15305(.A1(new_n8719_), .A2(new_n6090_), .ZN(new_n15370_));
  AOI21_X1   g15306(.A1(new_n15369_), .A2(new_n15370_), .B(new_n6082_), .ZN(new_n15371_));
  NAND2_X1   g15307(.A1(new_n12242_), .A2(new_n15371_), .ZN(new_n15372_));
  XOR2_X1    g15308(.A1(new_n15372_), .A2(\a[14] ), .Z(new_n15373_));
  INV_X1     g15309(.I(new_n15373_), .ZN(new_n15374_));
  XOR2_X1    g15310(.A1(new_n15223_), .A2(new_n15261_), .Z(new_n15375_));
  NAND2_X1   g15311(.A1(new_n15375_), .A2(new_n15374_), .ZN(new_n15376_));
  NAND3_X1   g15312(.A1(new_n15364_), .A2(new_n15376_), .A3(new_n15368_), .ZN(new_n15377_));
  NAND2_X1   g15313(.A1(new_n15377_), .A2(new_n15353_), .ZN(new_n15378_));
  INV_X1     g15314(.I(new_n15353_), .ZN(new_n15379_));
  AOI21_X1   g15315(.A1(new_n15365_), .A2(new_n15366_), .B(new_n15367_), .ZN(new_n15380_));
  NOR3_X1    g15316(.A1(new_n15358_), .A2(new_n15354_), .A3(new_n15363_), .ZN(new_n15381_));
  XOR2_X1    g15317(.A1(new_n15340_), .A2(new_n15261_), .Z(new_n15382_));
  NOR2_X1    g15318(.A1(new_n15382_), .A2(new_n15373_), .ZN(new_n15383_));
  NOR3_X1    g15319(.A1(new_n15380_), .A2(new_n15381_), .A3(new_n15383_), .ZN(new_n15384_));
  NAND2_X1   g15320(.A1(new_n15384_), .A2(new_n15379_), .ZN(new_n15385_));
  AOI21_X1   g15321(.A1(new_n15385_), .A2(new_n15378_), .B(new_n15348_), .ZN(new_n15386_));
  AOI21_X1   g15322(.A1(new_n15346_), .A2(new_n15345_), .B(new_n14562_), .ZN(new_n15387_));
  NOR3_X1    g15323(.A1(new_n15260_), .A2(new_n15343_), .A3(new_n15259_), .ZN(new_n15388_));
  NOR2_X1    g15324(.A1(new_n15387_), .A2(new_n15388_), .ZN(new_n15389_));
  NOR2_X1    g15325(.A1(new_n15384_), .A2(new_n15379_), .ZN(new_n15390_));
  NOR2_X1    g15326(.A1(new_n15377_), .A2(new_n15353_), .ZN(new_n15391_));
  NOR3_X1    g15327(.A1(new_n15390_), .A2(new_n15391_), .A3(new_n15389_), .ZN(new_n15392_));
  NOR2_X1    g15328(.A1(new_n15392_), .A2(new_n15386_), .ZN(new_n15393_));
  INV_X1     g15329(.I(new_n15393_), .ZN(new_n15394_));
  NAND3_X1   g15330(.A1(new_n15364_), .A2(new_n15383_), .A3(new_n15368_), .ZN(new_n15395_));
  OAI21_X1   g15331(.A1(new_n15380_), .A2(new_n15381_), .B(new_n15376_), .ZN(new_n15396_));
  AOI22_X1   g15332(.A1(new_n8702_), .A2(new_n6480_), .B1(new_n8696_), .B2(new_n4720_), .ZN(new_n15397_));
  NOR2_X1    g15333(.A1(new_n8681_), .A2(new_n4710_), .ZN(new_n15398_));
  OAI21_X1   g15334(.A1(new_n15398_), .A2(new_n15397_), .B(new_n4706_), .ZN(new_n15399_));
  NOR3_X1    g15335(.A1(new_n11612_), .A2(\a[11] ), .A3(new_n15399_), .ZN(new_n15400_));
  NOR2_X1    g15336(.A1(new_n11612_), .A2(new_n15399_), .ZN(new_n15401_));
  NOR2_X1    g15337(.A1(new_n15401_), .A2(new_n4034_), .ZN(new_n15402_));
  NOR2_X1    g15338(.A1(new_n15402_), .A2(new_n15400_), .ZN(new_n15403_));
  NAND3_X1   g15339(.A1(new_n15396_), .A2(new_n15395_), .A3(new_n15403_), .ZN(new_n15404_));
  NOR3_X1    g15340(.A1(new_n15380_), .A2(new_n15381_), .A3(new_n15376_), .ZN(new_n15405_));
  AOI21_X1   g15341(.A1(new_n15364_), .A2(new_n15368_), .B(new_n15383_), .ZN(new_n15406_));
  INV_X1     g15342(.I(new_n15403_), .ZN(new_n15407_));
  OAI21_X1   g15343(.A1(new_n15405_), .A2(new_n15406_), .B(new_n15407_), .ZN(new_n15408_));
  NAND2_X1   g15344(.A1(new_n15408_), .A2(new_n15404_), .ZN(new_n15409_));
  NAND2_X1   g15345(.A1(new_n15382_), .A2(new_n15373_), .ZN(new_n15410_));
  NAND2_X1   g15346(.A1(new_n15375_), .A2(new_n15374_), .ZN(new_n15411_));
  OAI22_X1   g15347(.A1(new_n4719_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n4716_), .ZN(new_n15412_));
  OAI21_X1   g15348(.A1(new_n4710_), .A2(new_n8694_), .B(new_n15412_), .ZN(new_n15413_));
  NAND4_X1   g15349(.A1(new_n11592_), .A2(new_n4706_), .A3(new_n11594_), .A4(new_n15413_), .ZN(new_n15414_));
  XOR2_X1    g15350(.A1(new_n15414_), .A2(new_n4034_), .Z(new_n15415_));
  AOI21_X1   g15351(.A1(new_n15411_), .A2(new_n15410_), .B(new_n15415_), .ZN(new_n15416_));
  NOR2_X1    g15352(.A1(new_n15375_), .A2(new_n15374_), .ZN(new_n15417_));
  NOR2_X1    g15353(.A1(new_n15382_), .A2(new_n15373_), .ZN(new_n15418_));
  XOR2_X1    g15354(.A1(new_n15414_), .A2(\a[11] ), .Z(new_n15419_));
  NOR3_X1    g15355(.A1(new_n15417_), .A2(new_n15418_), .A3(new_n15419_), .ZN(new_n15420_));
  NOR2_X1    g15356(.A1(new_n15416_), .A2(new_n15420_), .ZN(new_n15421_));
  OAI22_X1   g15357(.A1(new_n8710_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8718_), .ZN(new_n15422_));
  NAND2_X1   g15358(.A1(new_n8702_), .A2(new_n4709_), .ZN(new_n15423_));
  AOI21_X1   g15359(.A1(new_n15423_), .A2(new_n15422_), .B(new_n4707_), .ZN(new_n15424_));
  NAND2_X1   g15360(.A1(new_n12205_), .A2(new_n15424_), .ZN(new_n15425_));
  XOR2_X1    g15361(.A1(new_n15425_), .A2(\a[11] ), .Z(new_n15426_));
  NAND2_X1   g15362(.A1(new_n14725_), .A2(new_n14726_), .ZN(new_n15427_));
  NAND2_X1   g15363(.A1(new_n15339_), .A2(new_n14599_), .ZN(new_n15428_));
  NAND2_X1   g15364(.A1(new_n15222_), .A2(new_n14724_), .ZN(new_n15429_));
  AOI21_X1   g15365(.A1(new_n15428_), .A2(new_n15429_), .B(new_n15427_), .ZN(new_n15430_));
  NOR2_X1    g15366(.A1(new_n14722_), .A2(new_n14719_), .ZN(new_n15431_));
  NOR2_X1    g15367(.A1(new_n15222_), .A2(new_n14724_), .ZN(new_n15432_));
  NOR2_X1    g15368(.A1(new_n15339_), .A2(new_n14599_), .ZN(new_n15433_));
  NOR3_X1    g15369(.A1(new_n15433_), .A2(new_n15432_), .A3(new_n15431_), .ZN(new_n15434_));
  NOR2_X1    g15370(.A1(new_n15434_), .A2(new_n15430_), .ZN(new_n15435_));
  NAND3_X1   g15371(.A1(new_n15221_), .A2(new_n15264_), .A3(new_n15265_), .ZN(new_n15436_));
  AOI21_X1   g15372(.A1(new_n15165_), .A2(new_n15206_), .B(new_n15335_), .ZN(new_n15437_));
  NOR4_X1    g15373(.A1(new_n15437_), .A2(new_n15337_), .A3(new_n14748_), .A4(new_n14770_), .ZN(new_n15438_));
  OAI22_X1   g15374(.A1(new_n15438_), .A2(new_n14748_), .B1(new_n14735_), .B2(new_n14738_), .ZN(new_n15439_));
  OAI22_X1   g15375(.A1(new_n8751_), .A2(new_n6089_), .B1(new_n6094_), .B2(new_n10924_), .ZN(new_n15440_));
  NAND2_X1   g15376(.A1(new_n8736_), .A2(new_n6090_), .ZN(new_n15441_));
  AOI21_X1   g15377(.A1(new_n15441_), .A2(new_n15440_), .B(new_n6082_), .ZN(new_n15442_));
  NAND3_X1   g15378(.A1(new_n12118_), .A2(new_n3521_), .A3(new_n15442_), .ZN(new_n15443_));
  AOI21_X1   g15379(.A1(new_n12118_), .A2(new_n15442_), .B(new_n3521_), .ZN(new_n15444_));
  INV_X1     g15380(.I(new_n15444_), .ZN(new_n15445_));
  NAND2_X1   g15381(.A1(new_n15445_), .A2(new_n15443_), .ZN(new_n15446_));
  AOI21_X1   g15382(.A1(new_n15436_), .A2(new_n15439_), .B(new_n15446_), .ZN(new_n15447_));
  NOR3_X1    g15383(.A1(new_n15338_), .A2(new_n14735_), .A3(new_n14738_), .ZN(new_n15448_));
  AOI21_X1   g15384(.A1(new_n15264_), .A2(new_n15265_), .B(new_n15221_), .ZN(new_n15449_));
  INV_X1     g15385(.I(new_n15443_), .ZN(new_n15450_));
  NOR2_X1    g15386(.A1(new_n15450_), .A2(new_n15444_), .ZN(new_n15451_));
  NOR3_X1    g15387(.A1(new_n15449_), .A2(new_n15448_), .A3(new_n15451_), .ZN(new_n15452_));
  OAI22_X1   g15388(.A1(new_n8751_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8745_), .ZN(new_n15453_));
  NAND2_X1   g15389(.A1(new_n10927_), .A2(new_n6090_), .ZN(new_n15454_));
  AOI21_X1   g15390(.A1(new_n15453_), .A2(new_n15454_), .B(new_n6082_), .ZN(new_n15455_));
  NAND2_X1   g15391(.A1(new_n12072_), .A2(new_n15455_), .ZN(new_n15456_));
  XOR2_X1    g15392(.A1(new_n15456_), .A2(\a[14] ), .Z(new_n15457_));
  NAND2_X1   g15393(.A1(new_n15220_), .A2(new_n15272_), .ZN(new_n15458_));
  NAND2_X1   g15394(.A1(new_n15458_), .A2(new_n15219_), .ZN(new_n15459_));
  NAND3_X1   g15395(.A1(new_n15336_), .A2(new_n15272_), .A3(new_n15220_), .ZN(new_n15460_));
  NAND2_X1   g15396(.A1(new_n15459_), .A2(new_n15460_), .ZN(new_n15461_));
  NOR2_X1    g15397(.A1(new_n15461_), .A2(new_n15457_), .ZN(new_n15462_));
  NOR3_X1    g15398(.A1(new_n15452_), .A2(new_n15447_), .A3(new_n15462_), .ZN(new_n15463_));
  OAI22_X1   g15399(.A1(new_n8735_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n10924_), .ZN(new_n15464_));
  NAND2_X1   g15400(.A1(new_n8726_), .A2(new_n6090_), .ZN(new_n15465_));
  AOI21_X1   g15401(.A1(new_n15465_), .A2(new_n15464_), .B(new_n6082_), .ZN(new_n15466_));
  AND3_X2    g15402(.A1(new_n12181_), .A2(new_n3521_), .A3(new_n15466_), .Z(new_n15467_));
  AOI21_X1   g15403(.A1(new_n12181_), .A2(new_n15466_), .B(new_n3521_), .ZN(new_n15468_));
  NOR2_X1    g15404(.A1(new_n15467_), .A2(new_n15468_), .ZN(new_n15469_));
  INV_X1     g15405(.I(new_n15469_), .ZN(new_n15470_));
  NOR2_X1    g15406(.A1(new_n15463_), .A2(new_n15470_), .ZN(new_n15471_));
  OAI21_X1   g15407(.A1(new_n15449_), .A2(new_n15448_), .B(new_n15451_), .ZN(new_n15472_));
  NAND3_X1   g15408(.A1(new_n15436_), .A2(new_n15439_), .A3(new_n15446_), .ZN(new_n15473_));
  INV_X1     g15409(.I(new_n15457_), .ZN(new_n15474_));
  AOI21_X1   g15410(.A1(new_n15272_), .A2(new_n15220_), .B(new_n15336_), .ZN(new_n15475_));
  NOR2_X1    g15411(.A1(new_n15458_), .A2(new_n15219_), .ZN(new_n15476_));
  NOR2_X1    g15412(.A1(new_n15475_), .A2(new_n15476_), .ZN(new_n15477_));
  NAND2_X1   g15413(.A1(new_n15477_), .A2(new_n15474_), .ZN(new_n15478_));
  NAND3_X1   g15414(.A1(new_n15472_), .A2(new_n15473_), .A3(new_n15478_), .ZN(new_n15479_));
  NOR2_X1    g15415(.A1(new_n15479_), .A2(new_n15469_), .ZN(new_n15480_));
  OAI21_X1   g15416(.A1(new_n15471_), .A2(new_n15480_), .B(new_n15435_), .ZN(new_n15481_));
  OAI21_X1   g15417(.A1(new_n15433_), .A2(new_n15432_), .B(new_n15431_), .ZN(new_n15482_));
  NAND3_X1   g15418(.A1(new_n15428_), .A2(new_n15429_), .A3(new_n15427_), .ZN(new_n15483_));
  NAND2_X1   g15419(.A1(new_n15482_), .A2(new_n15483_), .ZN(new_n15484_));
  NAND2_X1   g15420(.A1(new_n15479_), .A2(new_n15469_), .ZN(new_n15485_));
  NAND4_X1   g15421(.A1(new_n15470_), .A2(new_n15472_), .A3(new_n15473_), .A4(new_n15478_), .ZN(new_n15486_));
  NAND3_X1   g15422(.A1(new_n15485_), .A2(new_n15484_), .A3(new_n15486_), .ZN(new_n15487_));
  NAND2_X1   g15423(.A1(new_n15481_), .A2(new_n15487_), .ZN(new_n15488_));
  NAND3_X1   g15424(.A1(new_n15472_), .A2(new_n15473_), .A3(new_n15462_), .ZN(new_n15489_));
  OAI21_X1   g15425(.A1(new_n15452_), .A2(new_n15447_), .B(new_n15478_), .ZN(new_n15490_));
  NOR2_X1    g15426(.A1(new_n10934_), .A2(new_n11535_), .ZN(new_n15491_));
  OAI22_X1   g15427(.A1(new_n8725_), .A2(new_n4716_), .B1(new_n4719_), .B2(new_n8718_), .ZN(new_n15492_));
  NAND2_X1   g15428(.A1(new_n8711_), .A2(new_n4709_), .ZN(new_n15493_));
  AOI21_X1   g15429(.A1(new_n15493_), .A2(new_n15492_), .B(new_n4707_), .ZN(new_n15494_));
  OAI21_X1   g15430(.A1(new_n15491_), .A2(new_n11532_), .B(new_n15494_), .ZN(new_n15495_));
  XOR2_X1    g15431(.A1(new_n15495_), .A2(\a[11] ), .Z(new_n15496_));
  NAND3_X1   g15432(.A1(new_n15490_), .A2(new_n15489_), .A3(new_n15496_), .ZN(new_n15497_));
  NOR3_X1    g15433(.A1(new_n15452_), .A2(new_n15447_), .A3(new_n15478_), .ZN(new_n15498_));
  AOI21_X1   g15434(.A1(new_n15472_), .A2(new_n15473_), .B(new_n15462_), .ZN(new_n15499_));
  XOR2_X1    g15435(.A1(new_n15495_), .A2(new_n4034_), .Z(new_n15500_));
  OAI21_X1   g15436(.A1(new_n15498_), .A2(new_n15499_), .B(new_n15500_), .ZN(new_n15501_));
  NAND2_X1   g15437(.A1(new_n15501_), .A2(new_n15497_), .ZN(new_n15502_));
  NOR2_X1    g15438(.A1(new_n15477_), .A2(new_n15474_), .ZN(new_n15503_));
  NOR2_X1    g15439(.A1(new_n15461_), .A2(new_n15457_), .ZN(new_n15504_));
  OAI22_X1   g15440(.A1(new_n8725_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8735_), .ZN(new_n15505_));
  NAND2_X1   g15441(.A1(new_n8719_), .A2(new_n4709_), .ZN(new_n15506_));
  AOI21_X1   g15442(.A1(new_n15505_), .A2(new_n15506_), .B(new_n4707_), .ZN(new_n15507_));
  OAI21_X1   g15443(.A1(new_n12239_), .A2(new_n12241_), .B(new_n15507_), .ZN(new_n15508_));
  XOR2_X1    g15444(.A1(new_n15508_), .A2(\a[11] ), .Z(new_n15509_));
  OAI21_X1   g15445(.A1(new_n15503_), .A2(new_n15504_), .B(new_n15509_), .ZN(new_n15510_));
  INV_X1     g15446(.I(new_n15510_), .ZN(new_n15511_));
  NAND2_X1   g15447(.A1(new_n15461_), .A2(new_n15457_), .ZN(new_n15512_));
  NAND2_X1   g15448(.A1(new_n15477_), .A2(new_n15474_), .ZN(new_n15513_));
  XOR2_X1    g15449(.A1(new_n15508_), .A2(new_n4034_), .Z(new_n15514_));
  NAND3_X1   g15450(.A1(new_n15513_), .A2(new_n15514_), .A3(new_n15512_), .ZN(new_n15515_));
  AND2_X2    g15451(.A1(new_n15510_), .A2(new_n15515_), .Z(new_n15516_));
  OAI22_X1   g15452(.A1(new_n8735_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n10924_), .ZN(new_n15517_));
  OAI21_X1   g15453(.A1(new_n4710_), .A2(new_n8725_), .B(new_n15517_), .ZN(new_n15518_));
  NAND4_X1   g15454(.A1(new_n12178_), .A2(new_n4706_), .A3(new_n12180_), .A4(new_n15518_), .ZN(new_n15519_));
  XOR2_X1    g15455(.A1(new_n15519_), .A2(\a[11] ), .Z(new_n15520_));
  AOI21_X1   g15456(.A1(new_n15207_), .A2(new_n15216_), .B(new_n14760_), .ZN(new_n15521_));
  OAI21_X1   g15457(.A1(new_n15330_), .A2(new_n15333_), .B(new_n15216_), .ZN(new_n15522_));
  NOR2_X1    g15458(.A1(new_n15522_), .A2(new_n15210_), .ZN(new_n15523_));
  OAI21_X1   g15459(.A1(new_n15523_), .A2(new_n15521_), .B(new_n14769_), .ZN(new_n15524_));
  INV_X1     g15460(.I(new_n14769_), .ZN(new_n15525_));
  NAND2_X1   g15461(.A1(new_n15522_), .A2(new_n15210_), .ZN(new_n15526_));
  NAND3_X1   g15462(.A1(new_n15207_), .A2(new_n14760_), .A3(new_n15216_), .ZN(new_n15527_));
  NAND3_X1   g15463(.A1(new_n15526_), .A2(new_n15527_), .A3(new_n15525_), .ZN(new_n15528_));
  NAND2_X1   g15464(.A1(new_n15524_), .A2(new_n15528_), .ZN(new_n15529_));
  NOR2_X1    g15465(.A1(new_n15330_), .A2(new_n15206_), .ZN(new_n15530_));
  NOR2_X1    g15466(.A1(new_n15165_), .A2(new_n15333_), .ZN(new_n15531_));
  OAI22_X1   g15467(.A1(new_n8758_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8766_), .ZN(new_n15532_));
  NAND2_X1   g15468(.A1(new_n8746_), .A2(new_n6090_), .ZN(new_n15533_));
  AOI21_X1   g15469(.A1(new_n15533_), .A2(new_n15532_), .B(new_n6082_), .ZN(new_n15534_));
  NAND3_X1   g15470(.A1(new_n11964_), .A2(new_n3521_), .A3(new_n15534_), .ZN(new_n15535_));
  INV_X1     g15471(.I(new_n15535_), .ZN(new_n15536_));
  AOI21_X1   g15472(.A1(new_n11964_), .A2(new_n15534_), .B(new_n3521_), .ZN(new_n15537_));
  NOR2_X1    g15473(.A1(new_n15536_), .A2(new_n15537_), .ZN(new_n15538_));
  OAI21_X1   g15474(.A1(new_n15531_), .A2(new_n15530_), .B(new_n15538_), .ZN(new_n15539_));
  OAI21_X1   g15475(.A1(new_n15328_), .A2(new_n15164_), .B(new_n15126_), .ZN(new_n15540_));
  NAND3_X1   g15476(.A1(new_n15325_), .A2(new_n15326_), .A3(new_n15162_), .ZN(new_n15541_));
  OAI21_X1   g15477(.A1(new_n15155_), .A2(new_n15157_), .B(new_n15327_), .ZN(new_n15542_));
  NAND2_X1   g15478(.A1(new_n15541_), .A2(new_n15542_), .ZN(new_n15543_));
  NAND2_X1   g15479(.A1(new_n15543_), .A2(new_n15324_), .ZN(new_n15544_));
  AOI22_X1   g15480(.A1(new_n6180_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n6095_), .ZN(new_n15545_));
  NOR2_X1    g15481(.A1(new_n8758_), .A2(new_n6091_), .ZN(new_n15546_));
  OAI21_X1   g15482(.A1(new_n15545_), .A2(new_n15546_), .B(new_n6081_), .ZN(new_n15547_));
  NOR2_X1    g15483(.A1(new_n12053_), .A2(new_n15547_), .ZN(new_n15548_));
  XOR2_X1    g15484(.A1(new_n15548_), .A2(new_n3521_), .Z(new_n15549_));
  AOI21_X1   g15485(.A1(new_n15544_), .A2(new_n15540_), .B(new_n15549_), .ZN(new_n15550_));
  NOR3_X1    g15486(.A1(new_n15531_), .A2(new_n15530_), .A3(new_n15538_), .ZN(new_n15551_));
  OAI21_X1   g15487(.A1(new_n15550_), .A2(new_n15551_), .B(new_n15539_), .ZN(new_n15552_));
  OAI22_X1   g15488(.A1(new_n8745_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8758_), .ZN(new_n15553_));
  NAND2_X1   g15489(.A1(new_n8752_), .A2(new_n6090_), .ZN(new_n15554_));
  AOI21_X1   g15490(.A1(new_n15554_), .A2(new_n15553_), .B(new_n6082_), .ZN(new_n15555_));
  NAND2_X1   g15491(.A1(new_n12189_), .A2(new_n15555_), .ZN(new_n15556_));
  XOR2_X1    g15492(.A1(new_n15556_), .A2(\a[14] ), .Z(new_n15557_));
  NAND2_X1   g15493(.A1(new_n15552_), .A2(new_n15557_), .ZN(new_n15558_));
  AOI21_X1   g15494(.A1(new_n15163_), .A2(new_n15329_), .B(new_n15324_), .ZN(new_n15559_));
  AOI21_X1   g15495(.A1(new_n15541_), .A2(new_n15542_), .B(new_n15126_), .ZN(new_n15560_));
  INV_X1     g15496(.I(new_n15549_), .ZN(new_n15561_));
  OAI21_X1   g15497(.A1(new_n15559_), .A2(new_n15560_), .B(new_n15561_), .ZN(new_n15562_));
  NAND2_X1   g15498(.A1(new_n15165_), .A2(new_n15333_), .ZN(new_n15563_));
  NAND2_X1   g15499(.A1(new_n15330_), .A2(new_n15206_), .ZN(new_n15564_));
  INV_X1     g15500(.I(new_n15537_), .ZN(new_n15565_));
  NAND2_X1   g15501(.A1(new_n15565_), .A2(new_n15535_), .ZN(new_n15566_));
  NAND3_X1   g15502(.A1(new_n15563_), .A2(new_n15564_), .A3(new_n15566_), .ZN(new_n15567_));
  NAND3_X1   g15503(.A1(new_n15539_), .A2(new_n15567_), .A3(new_n15562_), .ZN(new_n15568_));
  INV_X1     g15504(.I(new_n15557_), .ZN(new_n15569_));
  NAND3_X1   g15505(.A1(new_n15568_), .A2(new_n15539_), .A3(new_n15569_), .ZN(new_n15570_));
  AOI21_X1   g15506(.A1(new_n15558_), .A2(new_n15570_), .B(new_n15529_), .ZN(new_n15571_));
  AOI21_X1   g15507(.A1(new_n15526_), .A2(new_n15527_), .B(new_n15525_), .ZN(new_n15572_));
  NOR3_X1    g15508(.A1(new_n15523_), .A2(new_n15521_), .A3(new_n14769_), .ZN(new_n15573_));
  NOR2_X1    g15509(.A1(new_n15573_), .A2(new_n15572_), .ZN(new_n15574_));
  AOI21_X1   g15510(.A1(new_n15568_), .A2(new_n15539_), .B(new_n15569_), .ZN(new_n15575_));
  NOR2_X1    g15511(.A1(new_n15552_), .A2(new_n15557_), .ZN(new_n15576_));
  NOR3_X1    g15512(.A1(new_n15576_), .A2(new_n15575_), .A3(new_n15574_), .ZN(new_n15577_));
  NOR3_X1    g15513(.A1(new_n15577_), .A2(new_n15571_), .A3(new_n15520_), .ZN(new_n15578_));
  INV_X1     g15514(.I(new_n15520_), .ZN(new_n15579_));
  OAI21_X1   g15515(.A1(new_n15576_), .A2(new_n15575_), .B(new_n15574_), .ZN(new_n15580_));
  NAND3_X1   g15516(.A1(new_n15558_), .A2(new_n15570_), .A3(new_n15529_), .ZN(new_n15581_));
  AOI21_X1   g15517(.A1(new_n15580_), .A2(new_n15581_), .B(new_n15579_), .ZN(new_n15582_));
  AOI22_X1   g15518(.A1(new_n8752_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n10927_), .ZN(new_n15583_));
  NOR2_X1    g15519(.A1(new_n8735_), .A2(new_n4710_), .ZN(new_n15584_));
  OAI21_X1   g15520(.A1(new_n15584_), .A2(new_n15583_), .B(new_n4706_), .ZN(new_n15585_));
  INV_X1     g15521(.I(new_n15585_), .ZN(new_n15586_));
  NAND3_X1   g15522(.A1(new_n12118_), .A2(new_n4034_), .A3(new_n15586_), .ZN(new_n15587_));
  OAI21_X1   g15523(.A1(new_n12322_), .A2(new_n15585_), .B(\a[11] ), .ZN(new_n15588_));
  NAND2_X1   g15524(.A1(new_n15587_), .A2(new_n15588_), .ZN(new_n15589_));
  AOI21_X1   g15525(.A1(new_n15563_), .A2(new_n15564_), .B(new_n15566_), .ZN(new_n15590_));
  OAI21_X1   g15526(.A1(new_n15590_), .A2(new_n15551_), .B(new_n15562_), .ZN(new_n15591_));
  NAND3_X1   g15527(.A1(new_n15539_), .A2(new_n15567_), .A3(new_n15550_), .ZN(new_n15592_));
  AOI21_X1   g15528(.A1(new_n15591_), .A2(new_n15592_), .B(new_n15589_), .ZN(new_n15593_));
  AOI21_X1   g15529(.A1(new_n15539_), .A2(new_n15567_), .B(new_n15550_), .ZN(new_n15594_));
  NOR3_X1    g15530(.A1(new_n15590_), .A2(new_n15551_), .A3(new_n15562_), .ZN(new_n15595_));
  NOR3_X1    g15531(.A1(new_n15595_), .A2(new_n15594_), .A3(new_n15589_), .ZN(new_n15596_));
  NOR3_X1    g15532(.A1(new_n12322_), .A2(\a[11] ), .A3(new_n15585_), .ZN(new_n15597_));
  AOI21_X1   g15533(.A1(new_n12118_), .A2(new_n15586_), .B(new_n4034_), .ZN(new_n15598_));
  NOR2_X1    g15534(.A1(new_n15598_), .A2(new_n15597_), .ZN(new_n15599_));
  AOI21_X1   g15535(.A1(new_n15591_), .A2(new_n15592_), .B(new_n15599_), .ZN(new_n15600_));
  OAI22_X1   g15536(.A1(new_n8751_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8745_), .ZN(new_n15601_));
  NAND2_X1   g15537(.A1(new_n10927_), .A2(new_n4709_), .ZN(new_n15602_));
  AOI21_X1   g15538(.A1(new_n15601_), .A2(new_n15602_), .B(new_n4707_), .ZN(new_n15603_));
  AND3_X2    g15539(.A1(new_n12072_), .A2(new_n4034_), .A3(new_n15603_), .Z(new_n15604_));
  AOI21_X1   g15540(.A1(new_n12072_), .A2(new_n15603_), .B(new_n4034_), .ZN(new_n15605_));
  NOR3_X1    g15541(.A1(new_n15559_), .A2(new_n15561_), .A3(new_n15560_), .ZN(new_n15606_));
  NOR2_X1    g15542(.A1(new_n15606_), .A2(new_n15550_), .ZN(new_n15607_));
  OAI21_X1   g15543(.A1(new_n15604_), .A2(new_n15605_), .B(new_n15607_), .ZN(new_n15608_));
  NOR3_X1    g15544(.A1(new_n15596_), .A2(new_n15600_), .A3(new_n15608_), .ZN(new_n15609_));
  NOR2_X1    g15545(.A1(new_n15609_), .A2(new_n15593_), .ZN(new_n15610_));
  OAI22_X1   g15546(.A1(new_n15578_), .A2(new_n15582_), .B1(new_n15610_), .B2(new_n15520_), .ZN(new_n15611_));
  AOI21_X1   g15547(.A1(new_n15611_), .A2(new_n15516_), .B(new_n15511_), .ZN(new_n15612_));
  NOR2_X1    g15548(.A1(new_n15612_), .A2(new_n15502_), .ZN(new_n15613_));
  XOR2_X1    g15549(.A1(new_n15425_), .A2(new_n4034_), .Z(new_n15614_));
  NAND3_X1   g15550(.A1(new_n15481_), .A2(new_n15487_), .A3(new_n15614_), .ZN(new_n15615_));
  AOI21_X1   g15551(.A1(new_n15485_), .A2(new_n15486_), .B(new_n15484_), .ZN(new_n15616_));
  NOR3_X1    g15552(.A1(new_n15471_), .A2(new_n15480_), .A3(new_n15435_), .ZN(new_n15617_));
  OAI21_X1   g15553(.A1(new_n15617_), .A2(new_n15616_), .B(new_n15426_), .ZN(new_n15618_));
  NOR3_X1    g15554(.A1(new_n15498_), .A2(new_n15499_), .A3(new_n15500_), .ZN(new_n15619_));
  AOI21_X1   g15555(.A1(new_n15618_), .A2(new_n15615_), .B(new_n15619_), .ZN(new_n15620_));
  AOI22_X1   g15556(.A1(new_n15620_), .A2(new_n15613_), .B1(new_n15426_), .B2(new_n15488_), .ZN(new_n15621_));
  AOI21_X1   g15557(.A1(new_n15621_), .A2(new_n15421_), .B(new_n15416_), .ZN(new_n15622_));
  NOR2_X1    g15558(.A1(new_n15622_), .A2(new_n15409_), .ZN(new_n15623_));
  INV_X1     g15559(.I(new_n15258_), .ZN(new_n15624_));
  OAI21_X1   g15560(.A1(new_n15390_), .A2(new_n15391_), .B(new_n15389_), .ZN(new_n15625_));
  NAND3_X1   g15561(.A1(new_n15385_), .A2(new_n15378_), .A3(new_n15348_), .ZN(new_n15626_));
  NAND3_X1   g15562(.A1(new_n15625_), .A2(new_n15626_), .A3(new_n15624_), .ZN(new_n15627_));
  OAI21_X1   g15563(.A1(new_n15392_), .A2(new_n15386_), .B(new_n15258_), .ZN(new_n15628_));
  NOR3_X1    g15564(.A1(new_n15405_), .A2(new_n15406_), .A3(new_n15407_), .ZN(new_n15629_));
  AOI21_X1   g15565(.A1(new_n15628_), .A2(new_n15627_), .B(new_n15629_), .ZN(new_n15630_));
  AOI22_X1   g15566(.A1(new_n15630_), .A2(new_n15623_), .B1(new_n15258_), .B2(new_n15394_), .ZN(new_n15631_));
  XOR2_X1    g15567(.A1(new_n15631_), .A2(new_n15253_), .Z(new_n15632_));
  OAI22_X1   g15568(.A1(new_n11284_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8661_), .ZN(new_n15633_));
  NAND2_X1   g15569(.A1(new_n11272_), .A2(new_n6784_), .ZN(new_n15634_));
  AOI21_X1   g15570(.A1(new_n15633_), .A2(new_n15634_), .B(new_n6776_), .ZN(new_n15635_));
  NAND2_X1   g15571(.A1(new_n11655_), .A2(new_n15635_), .ZN(new_n15636_));
  XOR2_X1    g15572(.A1(new_n15636_), .A2(\a[8] ), .Z(new_n15637_));
  NOR2_X1    g15573(.A1(new_n15632_), .A2(new_n15637_), .ZN(new_n15638_));
  NOR3_X1    g15574(.A1(new_n15234_), .A2(new_n15227_), .A3(new_n15239_), .ZN(new_n15639_));
  NOR3_X1    g15575(.A1(new_n14476_), .A2(new_n14475_), .A3(new_n13983_), .ZN(new_n15640_));
  INV_X1     g15576(.I(new_n15640_), .ZN(new_n15641_));
  INV_X1     g15577(.I(new_n13840_), .ZN(new_n15642_));
  OAI21_X1   g15578(.A1(new_n15642_), .A2(new_n13841_), .B(new_n13829_), .ZN(new_n15643_));
  INV_X1     g15579(.I(new_n13829_), .ZN(new_n15644_));
  INV_X1     g15580(.I(new_n13839_), .ZN(new_n15645_));
  NOR2_X1    g15581(.A1(new_n13834_), .A2(new_n15645_), .ZN(new_n15646_));
  AOI21_X1   g15582(.A1(new_n13831_), .A2(new_n13833_), .B(new_n13839_), .ZN(new_n15647_));
  OAI21_X1   g15583(.A1(new_n15646_), .A2(new_n15647_), .B(new_n15644_), .ZN(new_n15648_));
  OAI22_X1   g15584(.A1(new_n8758_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8766_), .ZN(new_n15649_));
  NAND2_X1   g15585(.A1(new_n8746_), .A2(new_n3312_), .ZN(new_n15650_));
  AOI21_X1   g15586(.A1(new_n15650_), .A2(new_n15649_), .B(new_n3302_), .ZN(new_n15651_));
  NAND2_X1   g15587(.A1(new_n11964_), .A2(new_n15651_), .ZN(new_n15652_));
  XOR2_X1    g15588(.A1(new_n15652_), .A2(\a[23] ), .Z(new_n15653_));
  NAND3_X1   g15589(.A1(new_n15643_), .A2(new_n15648_), .A3(new_n15653_), .ZN(new_n15654_));
  INV_X1     g15590(.I(new_n13841_), .ZN(new_n15655_));
  AOI21_X1   g15591(.A1(new_n15655_), .A2(new_n13840_), .B(new_n15644_), .ZN(new_n15656_));
  NOR2_X1    g15592(.A1(new_n15646_), .A2(new_n15647_), .ZN(new_n15657_));
  NOR2_X1    g15593(.A1(new_n15657_), .A2(new_n13829_), .ZN(new_n15658_));
  INV_X1     g15594(.I(new_n15653_), .ZN(new_n15659_));
  OAI21_X1   g15595(.A1(new_n15658_), .A2(new_n15656_), .B(new_n15659_), .ZN(new_n15660_));
  NAND2_X1   g15596(.A1(new_n15660_), .A2(new_n15654_), .ZN(new_n15661_));
  INV_X1     g15597(.I(new_n14450_), .ZN(new_n15662_));
  OAI21_X1   g15598(.A1(new_n14471_), .A2(new_n14452_), .B(new_n15662_), .ZN(new_n15663_));
  NOR2_X1    g15599(.A1(new_n15663_), .A2(new_n15661_), .ZN(new_n15664_));
  NOR3_X1    g15600(.A1(new_n15658_), .A2(new_n15656_), .A3(new_n15659_), .ZN(new_n15665_));
  AOI21_X1   g15601(.A1(new_n15643_), .A2(new_n15648_), .B(new_n15653_), .ZN(new_n15666_));
  NOR2_X1    g15602(.A1(new_n15665_), .A2(new_n15666_), .ZN(new_n15667_));
  AOI21_X1   g15603(.A1(new_n14440_), .A2(new_n14453_), .B(new_n14450_), .ZN(new_n15668_));
  NOR2_X1    g15604(.A1(new_n15668_), .A2(new_n15667_), .ZN(new_n15669_));
  OAI22_X1   g15605(.A1(new_n8751_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n10924_), .ZN(new_n15670_));
  NAND2_X1   g15606(.A1(new_n8736_), .A2(new_n4096_), .ZN(new_n15671_));
  AOI21_X1   g15607(.A1(new_n15671_), .A2(new_n15670_), .B(new_n4095_), .ZN(new_n15672_));
  NAND2_X1   g15608(.A1(new_n12118_), .A2(new_n15672_), .ZN(new_n15673_));
  XOR2_X1    g15609(.A1(new_n15673_), .A2(\a[20] ), .Z(new_n15674_));
  OAI21_X1   g15610(.A1(new_n15669_), .A2(new_n15664_), .B(new_n15674_), .ZN(new_n15675_));
  NAND2_X1   g15611(.A1(new_n15668_), .A2(new_n15667_), .ZN(new_n15676_));
  NAND2_X1   g15612(.A1(new_n15663_), .A2(new_n15661_), .ZN(new_n15677_));
  INV_X1     g15613(.I(new_n15674_), .ZN(new_n15678_));
  NAND3_X1   g15614(.A1(new_n15676_), .A2(new_n15677_), .A3(new_n15678_), .ZN(new_n15679_));
  AOI21_X1   g15615(.A1(new_n15675_), .A2(new_n15679_), .B(new_n15641_), .ZN(new_n15680_));
  NAND3_X1   g15616(.A1(new_n15676_), .A2(new_n15677_), .A3(new_n15674_), .ZN(new_n15681_));
  OAI21_X1   g15617(.A1(new_n15669_), .A2(new_n15664_), .B(new_n15678_), .ZN(new_n15682_));
  AOI21_X1   g15618(.A1(new_n15682_), .A2(new_n15681_), .B(new_n15640_), .ZN(new_n15683_));
  OAI22_X1   g15619(.A1(new_n8725_), .A2(new_n4291_), .B1(new_n4297_), .B2(new_n8718_), .ZN(new_n15684_));
  NAND2_X1   g15620(.A1(new_n8711_), .A2(new_n4469_), .ZN(new_n15685_));
  AOI21_X1   g15621(.A1(new_n15685_), .A2(new_n15684_), .B(new_n4468_), .ZN(new_n15686_));
  NAND2_X1   g15622(.A1(new_n11536_), .A2(new_n15686_), .ZN(new_n15687_));
  XOR2_X1    g15623(.A1(new_n15687_), .A2(\a[17] ), .Z(new_n15688_));
  INV_X1     g15624(.I(new_n15688_), .ZN(new_n15689_));
  NOR3_X1    g15625(.A1(new_n15680_), .A2(new_n15683_), .A3(new_n15689_), .ZN(new_n15690_));
  AOI21_X1   g15626(.A1(new_n15676_), .A2(new_n15677_), .B(new_n15678_), .ZN(new_n15691_));
  NOR3_X1    g15627(.A1(new_n15669_), .A2(new_n15664_), .A3(new_n15674_), .ZN(new_n15692_));
  OAI21_X1   g15628(.A1(new_n15692_), .A2(new_n15691_), .B(new_n15640_), .ZN(new_n15693_));
  NOR3_X1    g15629(.A1(new_n15669_), .A2(new_n15664_), .A3(new_n15678_), .ZN(new_n15694_));
  AOI21_X1   g15630(.A1(new_n15676_), .A2(new_n15677_), .B(new_n15674_), .ZN(new_n15695_));
  OAI21_X1   g15631(.A1(new_n15694_), .A2(new_n15695_), .B(new_n15641_), .ZN(new_n15696_));
  AOI21_X1   g15632(.A1(new_n15693_), .A2(new_n15696_), .B(new_n15688_), .ZN(new_n15697_));
  NOR2_X1    g15633(.A1(new_n15697_), .A2(new_n15690_), .ZN(new_n15698_));
  NAND3_X1   g15634(.A1(new_n15228_), .A2(new_n15226_), .A3(new_n14563_), .ZN(new_n15699_));
  NAND3_X1   g15635(.A1(new_n15699_), .A2(new_n15698_), .A3(new_n14483_), .ZN(new_n15700_));
  OR2_X2     g15636(.A1(new_n15697_), .A2(new_n15690_), .Z(new_n15701_));
  OAI21_X1   g15637(.A1(new_n15233_), .A2(new_n14485_), .B(new_n14483_), .ZN(new_n15702_));
  NAND2_X1   g15638(.A1(new_n15701_), .A2(new_n15702_), .ZN(new_n15703_));
  OAI22_X1   g15639(.A1(new_n8701_), .A2(new_n6089_), .B1(new_n8694_), .B2(new_n6094_), .ZN(new_n15704_));
  NAND2_X1   g15640(.A1(new_n8682_), .A2(new_n6090_), .ZN(new_n15705_));
  AOI21_X1   g15641(.A1(new_n15705_), .A2(new_n15704_), .B(new_n6082_), .ZN(new_n15706_));
  NAND2_X1   g15642(.A1(new_n12347_), .A2(new_n15706_), .ZN(new_n15707_));
  XOR2_X1    g15643(.A1(new_n15707_), .A2(\a[14] ), .Z(new_n15708_));
  INV_X1     g15644(.I(new_n15708_), .ZN(new_n15709_));
  AOI21_X1   g15645(.A1(new_n15703_), .A2(new_n15700_), .B(new_n15709_), .ZN(new_n15710_));
  NOR2_X1    g15646(.A1(new_n15701_), .A2(new_n15702_), .ZN(new_n15711_));
  AOI21_X1   g15647(.A1(new_n15699_), .A2(new_n14483_), .B(new_n15698_), .ZN(new_n15712_));
  NOR3_X1    g15648(.A1(new_n15711_), .A2(new_n15712_), .A3(new_n15708_), .ZN(new_n15713_));
  OAI21_X1   g15649(.A1(new_n15713_), .A2(new_n15710_), .B(new_n15639_), .ZN(new_n15714_));
  INV_X1     g15650(.I(new_n15639_), .ZN(new_n15715_));
  NOR3_X1    g15651(.A1(new_n15711_), .A2(new_n15712_), .A3(new_n15709_), .ZN(new_n15716_));
  AOI21_X1   g15652(.A1(new_n15703_), .A2(new_n15700_), .B(new_n15708_), .ZN(new_n15717_));
  OAI21_X1   g15653(.A1(new_n15716_), .A2(new_n15717_), .B(new_n15715_), .ZN(new_n15718_));
  OAI22_X1   g15654(.A1(new_n8673_), .A2(new_n4719_), .B1(new_n8687_), .B2(new_n4716_), .ZN(new_n15719_));
  NAND2_X1   g15655(.A1(new_n8662_), .A2(new_n4709_), .ZN(new_n15720_));
  AOI21_X1   g15656(.A1(new_n15720_), .A2(new_n15719_), .B(new_n4707_), .ZN(new_n15721_));
  NAND2_X1   g15657(.A1(new_n11624_), .A2(new_n15721_), .ZN(new_n15722_));
  XOR2_X1    g15658(.A1(new_n15722_), .A2(\a[11] ), .Z(new_n15723_));
  NAND3_X1   g15659(.A1(new_n15714_), .A2(new_n15718_), .A3(new_n15723_), .ZN(new_n15724_));
  OAI21_X1   g15660(.A1(new_n15711_), .A2(new_n15712_), .B(new_n15708_), .ZN(new_n15725_));
  NAND3_X1   g15661(.A1(new_n15703_), .A2(new_n15700_), .A3(new_n15709_), .ZN(new_n15726_));
  AOI21_X1   g15662(.A1(new_n15725_), .A2(new_n15726_), .B(new_n15715_), .ZN(new_n15727_));
  NAND3_X1   g15663(.A1(new_n15703_), .A2(new_n15700_), .A3(new_n15708_), .ZN(new_n15728_));
  OAI21_X1   g15664(.A1(new_n15711_), .A2(new_n15712_), .B(new_n15709_), .ZN(new_n15729_));
  AOI21_X1   g15665(.A1(new_n15729_), .A2(new_n15728_), .B(new_n15639_), .ZN(new_n15730_));
  XOR2_X1    g15666(.A1(new_n15722_), .A2(new_n4034_), .Z(new_n15731_));
  OAI21_X1   g15667(.A1(new_n15727_), .A2(new_n15730_), .B(new_n15731_), .ZN(new_n15732_));
  NAND2_X1   g15668(.A1(new_n15732_), .A2(new_n15724_), .ZN(new_n15733_));
  NAND2_X1   g15669(.A1(new_n15251_), .A2(new_n15252_), .ZN(new_n15734_));
  AOI21_X1   g15670(.A1(new_n15396_), .A2(new_n15395_), .B(new_n15403_), .ZN(new_n15735_));
  NOR2_X1    g15671(.A1(new_n15629_), .A2(new_n15735_), .ZN(new_n15736_));
  INV_X1     g15672(.I(new_n15416_), .ZN(new_n15737_));
  NAND2_X1   g15673(.A1(new_n15488_), .A2(new_n15426_), .ZN(new_n15738_));
  INV_X1     g15674(.I(new_n15613_), .ZN(new_n15739_));
  NOR3_X1    g15675(.A1(new_n15617_), .A2(new_n15616_), .A3(new_n15426_), .ZN(new_n15740_));
  AOI21_X1   g15676(.A1(new_n15481_), .A2(new_n15487_), .B(new_n15614_), .ZN(new_n15741_));
  OAI21_X1   g15677(.A1(new_n15740_), .A2(new_n15741_), .B(new_n15497_), .ZN(new_n15742_));
  OAI21_X1   g15678(.A1(new_n15742_), .A2(new_n15739_), .B(new_n15738_), .ZN(new_n15743_));
  OAI21_X1   g15679(.A1(new_n15743_), .A2(new_n15420_), .B(new_n15737_), .ZN(new_n15744_));
  NAND2_X1   g15680(.A1(new_n15744_), .A2(new_n15736_), .ZN(new_n15745_));
  NOR3_X1    g15681(.A1(new_n15392_), .A2(new_n15386_), .A3(new_n15258_), .ZN(new_n15746_));
  AOI21_X1   g15682(.A1(new_n15625_), .A2(new_n15626_), .B(new_n15624_), .ZN(new_n15747_));
  OAI21_X1   g15683(.A1(new_n15746_), .A2(new_n15747_), .B(new_n15404_), .ZN(new_n15748_));
  OAI22_X1   g15684(.A1(new_n15748_), .A2(new_n15745_), .B1(new_n15624_), .B2(new_n15393_), .ZN(new_n15749_));
  OAI21_X1   g15685(.A1(new_n15749_), .A2(new_n15734_), .B(new_n15251_), .ZN(new_n15750_));
  NOR2_X1    g15686(.A1(new_n15750_), .A2(new_n15733_), .ZN(new_n15751_));
  NOR3_X1    g15687(.A1(new_n15727_), .A2(new_n15730_), .A3(new_n15731_), .ZN(new_n15752_));
  AOI21_X1   g15688(.A1(new_n15714_), .A2(new_n15718_), .B(new_n15723_), .ZN(new_n15753_));
  NOR2_X1    g15689(.A1(new_n15753_), .A2(new_n15752_), .ZN(new_n15754_));
  AOI21_X1   g15690(.A1(new_n15631_), .A2(new_n15253_), .B(new_n15250_), .ZN(new_n15755_));
  NOR2_X1    g15691(.A1(new_n15755_), .A2(new_n15754_), .ZN(new_n15756_));
  OAI22_X1   g15692(.A1(new_n11284_), .A2(new_n6783_), .B1(new_n6788_), .B2(new_n11271_), .ZN(new_n15757_));
  NAND2_X1   g15693(.A1(new_n11311_), .A2(new_n6784_), .ZN(new_n15758_));
  AOI21_X1   g15694(.A1(new_n15757_), .A2(new_n15758_), .B(new_n6776_), .ZN(new_n15759_));
  NAND2_X1   g15695(.A1(new_n11391_), .A2(new_n15759_), .ZN(new_n15760_));
  XOR2_X1    g15696(.A1(new_n15760_), .A2(\a[8] ), .Z(new_n15761_));
  OAI21_X1   g15697(.A1(new_n15751_), .A2(new_n15756_), .B(new_n15761_), .ZN(new_n15762_));
  NOR3_X1    g15698(.A1(new_n15751_), .A2(new_n15756_), .A3(new_n15761_), .ZN(new_n15763_));
  AOI21_X1   g15699(.A1(new_n15638_), .A2(new_n15762_), .B(new_n15763_), .ZN(new_n15764_));
  AOI21_X1   g15700(.A1(new_n15639_), .A2(new_n15725_), .B(new_n15713_), .ZN(new_n15765_));
  AOI21_X1   g15701(.A1(new_n15640_), .A2(new_n15675_), .B(new_n15692_), .ZN(new_n15766_));
  NAND2_X1   g15702(.A1(new_n13846_), .A2(new_n13851_), .ZN(new_n15767_));
  OAI21_X1   g15703(.A1(new_n13844_), .A2(new_n13845_), .B(new_n13852_), .ZN(new_n15768_));
  AOI21_X1   g15704(.A1(new_n15767_), .A2(new_n15768_), .B(new_n13842_), .ZN(new_n15769_));
  INV_X1     g15705(.I(new_n13842_), .ZN(new_n15770_));
  INV_X1     g15706(.I(new_n13853_), .ZN(new_n15771_));
  AOI21_X1   g15707(.A1(new_n15771_), .A2(new_n13854_), .B(new_n15770_), .ZN(new_n15772_));
  NOR2_X1    g15708(.A1(new_n15772_), .A2(new_n15769_), .ZN(new_n15773_));
  NOR2_X1    g15709(.A1(new_n15665_), .A2(new_n15666_), .ZN(new_n15774_));
  OAI22_X1   g15710(.A1(new_n8745_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8758_), .ZN(new_n15775_));
  NAND2_X1   g15711(.A1(new_n8752_), .A2(new_n3312_), .ZN(new_n15776_));
  AOI21_X1   g15712(.A1(new_n15776_), .A2(new_n15775_), .B(new_n3302_), .ZN(new_n15777_));
  NAND2_X1   g15713(.A1(new_n12189_), .A2(new_n15777_), .ZN(new_n15778_));
  XOR2_X1    g15714(.A1(new_n15778_), .A2(\a[23] ), .Z(new_n15779_));
  INV_X1     g15715(.I(new_n15779_), .ZN(new_n15780_));
  AOI21_X1   g15716(.A1(new_n15663_), .A2(new_n15774_), .B(new_n15780_), .ZN(new_n15781_));
  NAND3_X1   g15717(.A1(new_n15663_), .A2(new_n15774_), .A3(new_n15780_), .ZN(new_n15782_));
  INV_X1     g15718(.I(new_n15782_), .ZN(new_n15783_));
  OAI21_X1   g15719(.A1(new_n15783_), .A2(new_n15781_), .B(new_n15773_), .ZN(new_n15784_));
  NOR3_X1    g15720(.A1(new_n15773_), .A2(new_n15781_), .A3(new_n15783_), .ZN(new_n15785_));
  INV_X1     g15721(.I(new_n15785_), .ZN(new_n15786_));
  OAI22_X1   g15722(.A1(new_n8735_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n10924_), .ZN(new_n15787_));
  NAND2_X1   g15723(.A1(new_n8726_), .A2(new_n4096_), .ZN(new_n15788_));
  AOI21_X1   g15724(.A1(new_n15788_), .A2(new_n15787_), .B(new_n4095_), .ZN(new_n15789_));
  NAND2_X1   g15725(.A1(new_n12181_), .A2(new_n15789_), .ZN(new_n15790_));
  XOR2_X1    g15726(.A1(new_n15790_), .A2(\a[20] ), .Z(new_n15791_));
  NAND3_X1   g15727(.A1(new_n15786_), .A2(new_n15784_), .A3(new_n15791_), .ZN(new_n15792_));
  INV_X1     g15728(.I(new_n15784_), .ZN(new_n15793_));
  INV_X1     g15729(.I(new_n15791_), .ZN(new_n15794_));
  OAI21_X1   g15730(.A1(new_n15793_), .A2(new_n15785_), .B(new_n15794_), .ZN(new_n15795_));
  AOI21_X1   g15731(.A1(new_n15795_), .A2(new_n15792_), .B(new_n15766_), .ZN(new_n15796_));
  INV_X1     g15732(.I(new_n15766_), .ZN(new_n15797_));
  OAI21_X1   g15733(.A1(new_n15793_), .A2(new_n15785_), .B(new_n15791_), .ZN(new_n15798_));
  NAND3_X1   g15734(.A1(new_n15786_), .A2(new_n15784_), .A3(new_n15794_), .ZN(new_n15799_));
  AOI21_X1   g15735(.A1(new_n15798_), .A2(new_n15799_), .B(new_n15797_), .ZN(new_n15800_));
  NOR2_X1    g15736(.A1(new_n15796_), .A2(new_n15800_), .ZN(new_n15801_));
  NOR2_X1    g15737(.A1(new_n15697_), .A2(new_n15690_), .ZN(new_n15802_));
  OAI22_X1   g15738(.A1(new_n8710_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n8718_), .ZN(new_n15803_));
  NAND2_X1   g15739(.A1(new_n8702_), .A2(new_n4469_), .ZN(new_n15804_));
  AOI21_X1   g15740(.A1(new_n15804_), .A2(new_n15803_), .B(new_n4468_), .ZN(new_n15805_));
  NAND2_X1   g15741(.A1(new_n12205_), .A2(new_n15805_), .ZN(new_n15806_));
  XOR2_X1    g15742(.A1(new_n15806_), .A2(\a[17] ), .Z(new_n15807_));
  INV_X1     g15743(.I(new_n15807_), .ZN(new_n15808_));
  AOI21_X1   g15744(.A1(new_n15702_), .A2(new_n15802_), .B(new_n15808_), .ZN(new_n15809_));
  NAND3_X1   g15745(.A1(new_n15702_), .A2(new_n15802_), .A3(new_n15808_), .ZN(new_n15810_));
  INV_X1     g15746(.I(new_n15810_), .ZN(new_n15811_));
  OAI21_X1   g15747(.A1(new_n15811_), .A2(new_n15809_), .B(new_n15801_), .ZN(new_n15812_));
  OR3_X2     g15748(.A1(new_n15811_), .A2(new_n15801_), .A3(new_n15809_), .Z(new_n15813_));
  OAI22_X1   g15749(.A1(new_n8681_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8694_), .ZN(new_n15814_));
  NAND2_X1   g15750(.A1(new_n8688_), .A2(new_n6090_), .ZN(new_n15815_));
  AOI21_X1   g15751(.A1(new_n15815_), .A2(new_n15814_), .B(new_n6082_), .ZN(new_n15816_));
  NAND2_X1   g15752(.A1(new_n11420_), .A2(new_n15816_), .ZN(new_n15817_));
  XOR2_X1    g15753(.A1(new_n15817_), .A2(\a[14] ), .Z(new_n15818_));
  NAND3_X1   g15754(.A1(new_n15813_), .A2(new_n15812_), .A3(new_n15818_), .ZN(new_n15819_));
  INV_X1     g15755(.I(new_n15812_), .ZN(new_n15820_));
  NOR3_X1    g15756(.A1(new_n15811_), .A2(new_n15801_), .A3(new_n15809_), .ZN(new_n15821_));
  INV_X1     g15757(.I(new_n15818_), .ZN(new_n15822_));
  OAI21_X1   g15758(.A1(new_n15820_), .A2(new_n15821_), .B(new_n15822_), .ZN(new_n15823_));
  AOI21_X1   g15759(.A1(new_n15823_), .A2(new_n15819_), .B(new_n15765_), .ZN(new_n15824_));
  INV_X1     g15760(.I(new_n15765_), .ZN(new_n15825_));
  OAI21_X1   g15761(.A1(new_n15820_), .A2(new_n15821_), .B(new_n15818_), .ZN(new_n15826_));
  NAND3_X1   g15762(.A1(new_n15813_), .A2(new_n15812_), .A3(new_n15822_), .ZN(new_n15827_));
  AOI21_X1   g15763(.A1(new_n15826_), .A2(new_n15827_), .B(new_n15825_), .ZN(new_n15828_));
  NOR2_X1    g15764(.A1(new_n15824_), .A2(new_n15828_), .ZN(new_n15829_));
  OAI22_X1   g15765(.A1(new_n8661_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8673_), .ZN(new_n15830_));
  NAND2_X1   g15766(.A1(new_n11285_), .A2(new_n4709_), .ZN(new_n15831_));
  AOI21_X1   g15767(.A1(new_n15831_), .A2(new_n15830_), .B(new_n4707_), .ZN(new_n15832_));
  NAND2_X1   g15768(.A1(new_n11323_), .A2(new_n15832_), .ZN(new_n15833_));
  XOR2_X1    g15769(.A1(new_n15833_), .A2(\a[11] ), .Z(new_n15834_));
  INV_X1     g15770(.I(new_n15834_), .ZN(new_n15835_));
  NOR2_X1    g15771(.A1(new_n15753_), .A2(new_n15752_), .ZN(new_n15836_));
  AOI21_X1   g15772(.A1(new_n15750_), .A2(new_n15836_), .B(new_n15835_), .ZN(new_n15837_));
  NAND2_X1   g15773(.A1(new_n15732_), .A2(new_n15724_), .ZN(new_n15838_));
  NOR3_X1    g15774(.A1(new_n15755_), .A2(new_n15834_), .A3(new_n15838_), .ZN(new_n15839_));
  OAI21_X1   g15775(.A1(new_n15837_), .A2(new_n15839_), .B(new_n15829_), .ZN(new_n15840_));
  NOR3_X1    g15776(.A1(new_n15820_), .A2(new_n15821_), .A3(new_n15822_), .ZN(new_n15841_));
  AOI21_X1   g15777(.A1(new_n15813_), .A2(new_n15812_), .B(new_n15818_), .ZN(new_n15842_));
  OAI21_X1   g15778(.A1(new_n15841_), .A2(new_n15842_), .B(new_n15825_), .ZN(new_n15843_));
  AOI21_X1   g15779(.A1(new_n15813_), .A2(new_n15812_), .B(new_n15822_), .ZN(new_n15844_));
  NOR3_X1    g15780(.A1(new_n15820_), .A2(new_n15821_), .A3(new_n15818_), .ZN(new_n15845_));
  OAI21_X1   g15781(.A1(new_n15845_), .A2(new_n15844_), .B(new_n15765_), .ZN(new_n15846_));
  NAND2_X1   g15782(.A1(new_n15843_), .A2(new_n15846_), .ZN(new_n15847_));
  OAI21_X1   g15783(.A1(new_n15755_), .A2(new_n15838_), .B(new_n15834_), .ZN(new_n15848_));
  NAND3_X1   g15784(.A1(new_n15750_), .A2(new_n15835_), .A3(new_n15836_), .ZN(new_n15849_));
  NAND3_X1   g15785(.A1(new_n15849_), .A2(new_n15848_), .A3(new_n15847_), .ZN(new_n15850_));
  AOI22_X1   g15786(.A1(new_n11311_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n11272_), .ZN(new_n15851_));
  NOR2_X1    g15787(.A1(new_n11264_), .A2(new_n6785_), .ZN(new_n15852_));
  OAI21_X1   g15788(.A1(new_n15852_), .A2(new_n15851_), .B(new_n6775_), .ZN(new_n15853_));
  NOR2_X1    g15789(.A1(new_n11310_), .A2(new_n15853_), .ZN(new_n15854_));
  XOR2_X1    g15790(.A1(new_n15854_), .A2(new_n4009_), .Z(new_n15855_));
  NAND3_X1   g15791(.A1(new_n15840_), .A2(new_n15850_), .A3(new_n15855_), .ZN(new_n15856_));
  AOI21_X1   g15792(.A1(new_n15849_), .A2(new_n15848_), .B(new_n15847_), .ZN(new_n15857_));
  NOR3_X1    g15793(.A1(new_n15837_), .A2(new_n15839_), .A3(new_n15829_), .ZN(new_n15858_));
  XOR2_X1    g15794(.A1(new_n15854_), .A2(\a[8] ), .Z(new_n15859_));
  OAI21_X1   g15795(.A1(new_n15857_), .A2(new_n15858_), .B(new_n15859_), .ZN(new_n15860_));
  AOI21_X1   g15796(.A1(new_n15856_), .A2(new_n15860_), .B(new_n15764_), .ZN(new_n15861_));
  XOR2_X1    g15797(.A1(new_n15631_), .A2(new_n15734_), .Z(new_n15862_));
  INV_X1     g15798(.I(new_n15637_), .ZN(new_n15863_));
  NAND2_X1   g15799(.A1(new_n15862_), .A2(new_n15863_), .ZN(new_n15864_));
  NAND2_X1   g15800(.A1(new_n15755_), .A2(new_n15754_), .ZN(new_n15865_));
  NAND2_X1   g15801(.A1(new_n15750_), .A2(new_n15733_), .ZN(new_n15866_));
  XOR2_X1    g15802(.A1(new_n15760_), .A2(new_n4009_), .Z(new_n15867_));
  AOI21_X1   g15803(.A1(new_n15866_), .A2(new_n15865_), .B(new_n15867_), .ZN(new_n15868_));
  NAND3_X1   g15804(.A1(new_n15866_), .A2(new_n15865_), .A3(new_n15867_), .ZN(new_n15869_));
  OAI21_X1   g15805(.A1(new_n15864_), .A2(new_n15868_), .B(new_n15869_), .ZN(new_n15870_));
  OAI21_X1   g15806(.A1(new_n15857_), .A2(new_n15858_), .B(new_n15855_), .ZN(new_n15871_));
  NAND3_X1   g15807(.A1(new_n15840_), .A2(new_n15850_), .A3(new_n15859_), .ZN(new_n15872_));
  AOI21_X1   g15808(.A1(new_n15871_), .A2(new_n15872_), .B(new_n15870_), .ZN(new_n15873_));
  NOR3_X1    g15809(.A1(new_n13978_), .A2(new_n13971_), .A3(new_n13969_), .ZN(new_n15874_));
  NOR3_X1    g15810(.A1(new_n15861_), .A2(new_n15873_), .A3(new_n15874_), .ZN(new_n15875_));
  AOI21_X1   g15811(.A1(new_n13973_), .A2(new_n13978_), .B(new_n15875_), .ZN(new_n15876_));
  NAND2_X1   g15812(.A1(new_n13973_), .A2(new_n13978_), .ZN(new_n15877_));
  NOR3_X1    g15813(.A1(new_n15857_), .A2(new_n15858_), .A3(new_n15859_), .ZN(new_n15878_));
  AOI21_X1   g15814(.A1(new_n15840_), .A2(new_n15850_), .B(new_n15855_), .ZN(new_n15879_));
  OAI21_X1   g15815(.A1(new_n15878_), .A2(new_n15879_), .B(new_n15870_), .ZN(new_n15880_));
  AOI21_X1   g15816(.A1(new_n15840_), .A2(new_n15850_), .B(new_n15859_), .ZN(new_n15881_));
  NOR3_X1    g15817(.A1(new_n15857_), .A2(new_n15858_), .A3(new_n15855_), .ZN(new_n15882_));
  OAI21_X1   g15818(.A1(new_n15882_), .A2(new_n15881_), .B(new_n15764_), .ZN(new_n15883_));
  NAND2_X1   g15819(.A1(new_n15883_), .A2(new_n15880_), .ZN(new_n15884_));
  OAI21_X1   g15820(.A1(new_n15884_), .A2(new_n15874_), .B(new_n15877_), .ZN(new_n15885_));
  OAI22_X1   g15821(.A1(new_n11264_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n11277_), .ZN(new_n15886_));
  NAND2_X1   g15822(.A1(new_n11346_), .A2(new_n6784_), .ZN(new_n15887_));
  AOI21_X1   g15823(.A1(new_n15886_), .A2(new_n15887_), .B(new_n6776_), .ZN(new_n15888_));
  NAND2_X1   g15824(.A1(new_n11757_), .A2(new_n15888_), .ZN(new_n15889_));
  XOR2_X1    g15825(.A1(new_n15889_), .A2(\a[8] ), .Z(new_n15890_));
  OAI22_X1   g15826(.A1(new_n11284_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8661_), .ZN(new_n15891_));
  NAND2_X1   g15827(.A1(new_n11272_), .A2(new_n4709_), .ZN(new_n15892_));
  AOI21_X1   g15828(.A1(new_n15891_), .A2(new_n15892_), .B(new_n4707_), .ZN(new_n15893_));
  NAND2_X1   g15829(.A1(new_n11655_), .A2(new_n15893_), .ZN(new_n15894_));
  XOR2_X1    g15830(.A1(new_n15894_), .A2(\a[11] ), .Z(new_n15895_));
  INV_X1     g15831(.I(new_n15895_), .ZN(new_n15896_));
  OAI22_X1   g15832(.A1(new_n4297_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n4291_), .ZN(new_n15897_));
  NAND2_X1   g15833(.A1(new_n8696_), .A2(new_n4469_), .ZN(new_n15898_));
  AOI21_X1   g15834(.A1(new_n15897_), .A2(new_n15898_), .B(new_n4468_), .ZN(new_n15899_));
  NAND2_X1   g15835(.A1(new_n11595_), .A2(new_n15899_), .ZN(new_n15900_));
  XOR2_X1    g15836(.A1(new_n15900_), .A2(\a[17] ), .Z(new_n15901_));
  INV_X1     g15837(.I(new_n15901_), .ZN(new_n15902_));
  OAI22_X1   g15838(.A1(new_n8725_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n8735_), .ZN(new_n15903_));
  NAND2_X1   g15839(.A1(new_n8719_), .A2(new_n4096_), .ZN(new_n15904_));
  AOI21_X1   g15840(.A1(new_n15903_), .A2(new_n15904_), .B(new_n4095_), .ZN(new_n15905_));
  NAND2_X1   g15841(.A1(new_n12242_), .A2(new_n15905_), .ZN(new_n15906_));
  XOR2_X1    g15842(.A1(new_n15906_), .A2(\a[20] ), .Z(new_n15907_));
  NAND2_X1   g15843(.A1(new_n13862_), .A2(new_n13864_), .ZN(new_n15908_));
  NAND2_X1   g15844(.A1(new_n13818_), .A2(new_n15908_), .ZN(new_n15909_));
  XOR2_X1    g15845(.A1(new_n13855_), .A2(new_n13860_), .Z(new_n15910_));
  NOR2_X1    g15846(.A1(new_n13818_), .A2(new_n15910_), .ZN(new_n15911_));
  INV_X1     g15847(.I(new_n15911_), .ZN(new_n15912_));
  NAND2_X1   g15848(.A1(new_n15798_), .A2(new_n15797_), .ZN(new_n15913_));
  NAND2_X1   g15849(.A1(new_n15913_), .A2(new_n15799_), .ZN(new_n15914_));
  NAND3_X1   g15850(.A1(new_n15912_), .A2(new_n15909_), .A3(new_n15914_), .ZN(new_n15915_));
  INV_X1     g15851(.I(new_n15915_), .ZN(new_n15916_));
  AOI21_X1   g15852(.A1(new_n15912_), .A2(new_n15909_), .B(new_n15914_), .ZN(new_n15917_));
  OAI21_X1   g15853(.A1(new_n15916_), .A2(new_n15917_), .B(new_n15907_), .ZN(new_n15918_));
  INV_X1     g15854(.I(new_n15907_), .ZN(new_n15919_));
  INV_X1     g15855(.I(new_n15909_), .ZN(new_n15920_));
  INV_X1     g15856(.I(new_n15914_), .ZN(new_n15921_));
  OAI21_X1   g15857(.A1(new_n15920_), .A2(new_n15911_), .B(new_n15921_), .ZN(new_n15922_));
  NAND3_X1   g15858(.A1(new_n15922_), .A2(new_n15915_), .A3(new_n15919_), .ZN(new_n15923_));
  AOI21_X1   g15859(.A1(new_n15918_), .A2(new_n15923_), .B(new_n15902_), .ZN(new_n15924_));
  AOI21_X1   g15860(.A1(new_n15922_), .A2(new_n15915_), .B(new_n15919_), .ZN(new_n15925_));
  INV_X1     g15861(.I(new_n15923_), .ZN(new_n15926_));
  NOR3_X1    g15862(.A1(new_n15926_), .A2(new_n15925_), .A3(new_n15901_), .ZN(new_n15927_));
  OAI22_X1   g15863(.A1(new_n6089_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n6094_), .ZN(new_n15928_));
  NAND2_X1   g15864(.A1(new_n8674_), .A2(new_n6090_), .ZN(new_n15929_));
  AOI21_X1   g15865(.A1(new_n15929_), .A2(new_n15928_), .B(new_n6082_), .ZN(new_n15930_));
  NAND2_X1   g15866(.A1(new_n11431_), .A2(new_n15930_), .ZN(new_n15931_));
  XOR2_X1    g15867(.A1(new_n15931_), .A2(\a[14] ), .Z(new_n15932_));
  OAI21_X1   g15868(.A1(new_n15927_), .A2(new_n15924_), .B(new_n15932_), .ZN(new_n15933_));
  OAI21_X1   g15869(.A1(new_n15926_), .A2(new_n15925_), .B(new_n15901_), .ZN(new_n15934_));
  NAND3_X1   g15870(.A1(new_n15918_), .A2(new_n15923_), .A3(new_n15902_), .ZN(new_n15935_));
  INV_X1     g15871(.I(new_n15932_), .ZN(new_n15936_));
  NAND3_X1   g15872(.A1(new_n15934_), .A2(new_n15935_), .A3(new_n15936_), .ZN(new_n15937_));
  AOI21_X1   g15873(.A1(new_n15825_), .A2(new_n15826_), .B(new_n15845_), .ZN(new_n15938_));
  INV_X1     g15874(.I(new_n15938_), .ZN(new_n15939_));
  NAND3_X1   g15875(.A1(new_n15933_), .A2(new_n15937_), .A3(new_n15939_), .ZN(new_n15940_));
  AOI21_X1   g15876(.A1(new_n15934_), .A2(new_n15935_), .B(new_n15936_), .ZN(new_n15941_));
  NOR3_X1    g15877(.A1(new_n15927_), .A2(new_n15924_), .A3(new_n15932_), .ZN(new_n15942_));
  OAI21_X1   g15878(.A1(new_n15942_), .A2(new_n15941_), .B(new_n15938_), .ZN(new_n15943_));
  AOI21_X1   g15879(.A1(new_n15943_), .A2(new_n15940_), .B(new_n15896_), .ZN(new_n15944_));
  NOR3_X1    g15880(.A1(new_n15942_), .A2(new_n15941_), .A3(new_n15938_), .ZN(new_n15945_));
  AOI21_X1   g15881(.A1(new_n15933_), .A2(new_n15937_), .B(new_n15939_), .ZN(new_n15946_));
  NOR3_X1    g15882(.A1(new_n15945_), .A2(new_n15946_), .A3(new_n15895_), .ZN(new_n15947_));
  OAI21_X1   g15883(.A1(new_n15947_), .A2(new_n15944_), .B(new_n15890_), .ZN(new_n15948_));
  INV_X1     g15884(.I(new_n15890_), .ZN(new_n15949_));
  OAI21_X1   g15885(.A1(new_n15945_), .A2(new_n15946_), .B(new_n15895_), .ZN(new_n15950_));
  NAND3_X1   g15886(.A1(new_n15943_), .A2(new_n15940_), .A3(new_n15896_), .ZN(new_n15951_));
  NAND3_X1   g15887(.A1(new_n15950_), .A2(new_n15951_), .A3(new_n15949_), .ZN(new_n15952_));
  NAND2_X1   g15888(.A1(new_n15948_), .A2(new_n15952_), .ZN(new_n15953_));
  NOR2_X1    g15889(.A1(new_n15881_), .A2(new_n15764_), .ZN(new_n15954_));
  OAI22_X1   g15890(.A1(new_n11353_), .A2(new_n6913_), .B1(new_n6839_), .B2(new_n11697_), .ZN(new_n15955_));
  NAND2_X1   g15891(.A1(new_n11370_), .A2(new_n8799_), .ZN(new_n15956_));
  AOI21_X1   g15892(.A1(new_n15956_), .A2(new_n15955_), .B(new_n6836_), .ZN(new_n15957_));
  OAI21_X1   g15893(.A1(new_n11696_), .A2(new_n11699_), .B(new_n15957_), .ZN(new_n15958_));
  XOR2_X1    g15894(.A1(new_n15958_), .A2(new_n65_), .Z(new_n15959_));
  NOR3_X1    g15895(.A1(new_n15954_), .A2(new_n15959_), .A3(new_n15882_), .ZN(new_n15960_));
  NAND2_X1   g15896(.A1(new_n15871_), .A2(new_n15870_), .ZN(new_n15961_));
  XOR2_X1    g15897(.A1(new_n15958_), .A2(\a[5] ), .Z(new_n15962_));
  AOI21_X1   g15898(.A1(new_n15961_), .A2(new_n15872_), .B(new_n15962_), .ZN(new_n15963_));
  OAI21_X1   g15899(.A1(new_n15963_), .A2(new_n15960_), .B(new_n15953_), .ZN(new_n15964_));
  AOI21_X1   g15900(.A1(new_n15950_), .A2(new_n15951_), .B(new_n15949_), .ZN(new_n15965_));
  NOR3_X1    g15901(.A1(new_n15947_), .A2(new_n15944_), .A3(new_n15890_), .ZN(new_n15966_));
  NOR2_X1    g15902(.A1(new_n15966_), .A2(new_n15965_), .ZN(new_n15967_));
  AOI21_X1   g15903(.A1(new_n15961_), .A2(new_n15872_), .B(new_n15959_), .ZN(new_n15968_));
  NOR3_X1    g15904(.A1(new_n15954_), .A2(new_n15962_), .A3(new_n15882_), .ZN(new_n15969_));
  OAI21_X1   g15905(.A1(new_n15968_), .A2(new_n15969_), .B(new_n15967_), .ZN(new_n15970_));
  NAND3_X1   g15906(.A1(new_n15885_), .A2(new_n15970_), .A3(new_n15964_), .ZN(new_n15971_));
  INV_X1     g15907(.I(new_n15960_), .ZN(new_n15972_));
  NAND2_X1   g15908(.A1(new_n15961_), .A2(new_n15872_), .ZN(new_n15973_));
  NAND2_X1   g15909(.A1(new_n15973_), .A2(new_n15959_), .ZN(new_n15974_));
  AOI21_X1   g15910(.A1(new_n15972_), .A2(new_n15974_), .B(new_n15967_), .ZN(new_n15975_));
  NAND2_X1   g15911(.A1(new_n15973_), .A2(new_n15962_), .ZN(new_n15976_));
  NAND3_X1   g15912(.A1(new_n15961_), .A2(new_n15959_), .A3(new_n15872_), .ZN(new_n15977_));
  AOI21_X1   g15913(.A1(new_n15976_), .A2(new_n15977_), .B(new_n15953_), .ZN(new_n15978_));
  OAI21_X1   g15914(.A1(new_n15975_), .A2(new_n15978_), .B(new_n15876_), .ZN(new_n15979_));
  NAND2_X1   g15915(.A1(new_n15979_), .A2(new_n15971_), .ZN(new_n15980_));
  NOR2_X1    g15916(.A1(new_n11308_), .A2(new_n11304_), .ZN(new_n15981_));
  AOI21_X1   g15917(.A1(new_n11302_), .A2(new_n11279_), .B(new_n11264_), .ZN(new_n15982_));
  NOR2_X1    g15918(.A1(new_n15982_), .A2(new_n15981_), .ZN(new_n15983_));
  AOI22_X1   g15919(.A1(new_n11311_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n11272_), .ZN(new_n15984_));
  NOR2_X1    g15920(.A1(new_n11264_), .A2(new_n6839_), .ZN(new_n15985_));
  OAI21_X1   g15921(.A1(new_n15985_), .A2(new_n15984_), .B(new_n6835_), .ZN(new_n15986_));
  INV_X1     g15922(.I(new_n15986_), .ZN(new_n15987_));
  NAND3_X1   g15923(.A1(new_n15983_), .A2(new_n65_), .A3(new_n15987_), .ZN(new_n15988_));
  OAI21_X1   g15924(.A1(new_n11310_), .A2(new_n15986_), .B(\a[5] ), .ZN(new_n15989_));
  NAND2_X1   g15925(.A1(new_n15988_), .A2(new_n15989_), .ZN(new_n15990_));
  OAI21_X1   g15926(.A1(new_n15745_), .A2(new_n15629_), .B(new_n15258_), .ZN(new_n15991_));
  NAND4_X1   g15927(.A1(new_n15744_), .A2(new_n15624_), .A3(new_n15404_), .A4(new_n15736_), .ZN(new_n15992_));
  AOI21_X1   g15928(.A1(new_n15991_), .A2(new_n15992_), .B(new_n15394_), .ZN(new_n15993_));
  AOI21_X1   g15929(.A1(new_n15623_), .A2(new_n15404_), .B(new_n15624_), .ZN(new_n15994_));
  INV_X1     g15930(.I(new_n15992_), .ZN(new_n15995_));
  NOR3_X1    g15931(.A1(new_n15994_), .A2(new_n15995_), .A3(new_n15393_), .ZN(new_n15996_));
  NOR2_X1    g15932(.A1(new_n15996_), .A2(new_n15993_), .ZN(new_n15997_));
  NAND2_X1   g15933(.A1(new_n15620_), .A2(new_n15613_), .ZN(new_n15998_));
  NAND3_X1   g15934(.A1(new_n15998_), .A2(new_n15421_), .A3(new_n15738_), .ZN(new_n15999_));
  NAND3_X1   g15935(.A1(new_n15999_), .A2(new_n15736_), .A3(new_n15737_), .ZN(new_n16000_));
  NAND2_X1   g15936(.A1(new_n15744_), .A2(new_n15409_), .ZN(new_n16001_));
  OAI22_X1   g15937(.A1(new_n8673_), .A2(new_n6788_), .B1(new_n8687_), .B2(new_n6783_), .ZN(new_n16002_));
  NAND2_X1   g15938(.A1(new_n8662_), .A2(new_n6784_), .ZN(new_n16003_));
  AOI21_X1   g15939(.A1(new_n16003_), .A2(new_n16002_), .B(new_n6776_), .ZN(new_n16004_));
  NAND2_X1   g15940(.A1(new_n11624_), .A2(new_n16004_), .ZN(new_n16005_));
  XOR2_X1    g15941(.A1(new_n16005_), .A2(new_n4009_), .Z(new_n16006_));
  AOI21_X1   g15942(.A1(new_n16001_), .A2(new_n16000_), .B(new_n16006_), .ZN(new_n16007_));
  NOR2_X1    g15943(.A1(new_n15744_), .A2(new_n15409_), .ZN(new_n16008_));
  NOR2_X1    g15944(.A1(new_n15622_), .A2(new_n15736_), .ZN(new_n16009_));
  XOR2_X1    g15945(.A1(new_n16005_), .A2(\a[8] ), .Z(new_n16010_));
  NOR3_X1    g15946(.A1(new_n16009_), .A2(new_n16008_), .A3(new_n16010_), .ZN(new_n16011_));
  OAI22_X1   g15947(.A1(new_n6783_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n6788_), .ZN(new_n16012_));
  NAND2_X1   g15948(.A1(new_n8674_), .A2(new_n6784_), .ZN(new_n16013_));
  AOI21_X1   g15949(.A1(new_n16013_), .A2(new_n16012_), .B(new_n6776_), .ZN(new_n16014_));
  NAND2_X1   g15950(.A1(new_n11431_), .A2(new_n16014_), .ZN(new_n16015_));
  XOR2_X1    g15951(.A1(new_n16015_), .A2(\a[8] ), .Z(new_n16016_));
  INV_X1     g15952(.I(new_n16016_), .ZN(new_n16017_));
  NAND2_X1   g15953(.A1(new_n15743_), .A2(new_n15421_), .ZN(new_n16018_));
  OR2_X2     g15954(.A1(new_n15416_), .A2(new_n15420_), .Z(new_n16019_));
  NAND2_X1   g15955(.A1(new_n15621_), .A2(new_n16019_), .ZN(new_n16020_));
  NAND3_X1   g15956(.A1(new_n16017_), .A2(new_n16020_), .A3(new_n16018_), .ZN(new_n16021_));
  INV_X1     g15957(.I(new_n16021_), .ZN(new_n16022_));
  NOR3_X1    g15958(.A1(new_n16011_), .A2(new_n16007_), .A3(new_n16022_), .ZN(new_n16023_));
  OAI22_X1   g15959(.A1(new_n8661_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8673_), .ZN(new_n16024_));
  NAND2_X1   g15960(.A1(new_n11285_), .A2(new_n6784_), .ZN(new_n16025_));
  AOI21_X1   g15961(.A1(new_n16025_), .A2(new_n16024_), .B(new_n6776_), .ZN(new_n16026_));
  NAND2_X1   g15962(.A1(new_n11323_), .A2(new_n16026_), .ZN(new_n16027_));
  XOR2_X1    g15963(.A1(new_n16027_), .A2(new_n4009_), .Z(new_n16028_));
  NOR2_X1    g15964(.A1(new_n16023_), .A2(new_n16028_), .ZN(new_n16029_));
  XOR2_X1    g15965(.A1(new_n16027_), .A2(\a[8] ), .Z(new_n16030_));
  NOR4_X1    g15966(.A1(new_n16011_), .A2(new_n16030_), .A3(new_n16007_), .A4(new_n16022_), .ZN(new_n16031_));
  OAI21_X1   g15967(.A1(new_n16029_), .A2(new_n16031_), .B(new_n15997_), .ZN(new_n16032_));
  OAI21_X1   g15968(.A1(new_n15994_), .A2(new_n15995_), .B(new_n15393_), .ZN(new_n16033_));
  NAND3_X1   g15969(.A1(new_n15991_), .A2(new_n15394_), .A3(new_n15992_), .ZN(new_n16034_));
  NAND2_X1   g15970(.A1(new_n16033_), .A2(new_n16034_), .ZN(new_n16035_));
  OAI21_X1   g15971(.A1(new_n16009_), .A2(new_n16008_), .B(new_n16010_), .ZN(new_n16036_));
  NAND3_X1   g15972(.A1(new_n16001_), .A2(new_n16006_), .A3(new_n16000_), .ZN(new_n16037_));
  NAND3_X1   g15973(.A1(new_n16036_), .A2(new_n16037_), .A3(new_n16021_), .ZN(new_n16038_));
  NAND2_X1   g15974(.A1(new_n16038_), .A2(new_n16030_), .ZN(new_n16039_));
  NAND4_X1   g15975(.A1(new_n16028_), .A2(new_n16036_), .A3(new_n16037_), .A4(new_n16021_), .ZN(new_n16040_));
  NAND3_X1   g15976(.A1(new_n16039_), .A2(new_n16035_), .A3(new_n16040_), .ZN(new_n16041_));
  NAND3_X1   g15977(.A1(new_n16032_), .A2(new_n16041_), .A3(new_n15990_), .ZN(new_n16042_));
  NOR3_X1    g15978(.A1(new_n11310_), .A2(\a[5] ), .A3(new_n15986_), .ZN(new_n16043_));
  AOI21_X1   g15979(.A1(new_n15983_), .A2(new_n15987_), .B(new_n65_), .ZN(new_n16044_));
  NOR2_X1    g15980(.A1(new_n16044_), .A2(new_n16043_), .ZN(new_n16045_));
  AOI21_X1   g15981(.A1(new_n16039_), .A2(new_n16040_), .B(new_n16035_), .ZN(new_n16046_));
  NOR3_X1    g15982(.A1(new_n16029_), .A2(new_n15997_), .A3(new_n16031_), .ZN(new_n16047_));
  OAI21_X1   g15983(.A1(new_n16046_), .A2(new_n16047_), .B(new_n16045_), .ZN(new_n16048_));
  NAND3_X1   g15984(.A1(new_n16036_), .A2(new_n16037_), .A3(new_n16022_), .ZN(new_n16049_));
  OAI21_X1   g15985(.A1(new_n16011_), .A2(new_n16007_), .B(new_n16021_), .ZN(new_n16050_));
  OAI22_X1   g15986(.A1(new_n11284_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n11271_), .ZN(new_n16051_));
  NAND2_X1   g15987(.A1(new_n11311_), .A2(new_n6838_), .ZN(new_n16052_));
  AOI21_X1   g15988(.A1(new_n16051_), .A2(new_n16052_), .B(new_n6836_), .ZN(new_n16053_));
  OAI21_X1   g15989(.A1(new_n11388_), .A2(new_n11390_), .B(new_n16053_), .ZN(new_n16054_));
  XOR2_X1    g15990(.A1(new_n16054_), .A2(\a[5] ), .Z(new_n16055_));
  NAND3_X1   g15991(.A1(new_n16050_), .A2(new_n16049_), .A3(new_n16055_), .ZN(new_n16056_));
  NOR3_X1    g15992(.A1(new_n16011_), .A2(new_n16007_), .A3(new_n16021_), .ZN(new_n16057_));
  AOI21_X1   g15993(.A1(new_n16036_), .A2(new_n16037_), .B(new_n16022_), .ZN(new_n16058_));
  XOR2_X1    g15994(.A1(new_n16054_), .A2(new_n65_), .Z(new_n16059_));
  OAI21_X1   g15995(.A1(new_n16057_), .A2(new_n16058_), .B(new_n16059_), .ZN(new_n16060_));
  AOI21_X1   g15996(.A1(new_n16020_), .A2(new_n16018_), .B(new_n16017_), .ZN(new_n16061_));
  INV_X1     g15997(.I(new_n16061_), .ZN(new_n16062_));
  NAND3_X1   g15998(.A1(new_n16017_), .A2(new_n16020_), .A3(new_n16018_), .ZN(new_n16063_));
  OAI22_X1   g15999(.A1(new_n11284_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8661_), .ZN(new_n16064_));
  NAND2_X1   g16000(.A1(new_n11272_), .A2(new_n6838_), .ZN(new_n16065_));
  AOI21_X1   g16001(.A1(new_n16064_), .A2(new_n16065_), .B(new_n6836_), .ZN(new_n16066_));
  NAND3_X1   g16002(.A1(new_n11651_), .A2(new_n11654_), .A3(new_n16066_), .ZN(new_n16067_));
  XOR2_X1    g16003(.A1(new_n16067_), .A2(new_n65_), .Z(new_n16068_));
  AOI21_X1   g16004(.A1(new_n16062_), .A2(new_n16063_), .B(new_n16068_), .ZN(new_n16069_));
  INV_X1     g16005(.I(new_n16069_), .ZN(new_n16070_));
  INV_X1     g16006(.I(new_n16063_), .ZN(new_n16071_));
  XOR2_X1    g16007(.A1(new_n16067_), .A2(\a[5] ), .Z(new_n16072_));
  NOR3_X1    g16008(.A1(new_n16072_), .A2(new_n16071_), .A3(new_n16061_), .ZN(new_n16073_));
  OAI22_X1   g16009(.A1(new_n8661_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8673_), .ZN(new_n16074_));
  NAND2_X1   g16010(.A1(new_n11285_), .A2(new_n6838_), .ZN(new_n16075_));
  AOI21_X1   g16011(.A1(new_n16075_), .A2(new_n16074_), .B(new_n6836_), .ZN(new_n16076_));
  OAI21_X1   g16012(.A1(new_n11321_), .A2(new_n11322_), .B(new_n16076_), .ZN(new_n16077_));
  XOR2_X1    g16013(.A1(new_n16077_), .A2(new_n65_), .Z(new_n16078_));
  AOI21_X1   g16014(.A1(new_n15490_), .A2(new_n15489_), .B(new_n15496_), .ZN(new_n16079_));
  NOR2_X1    g16015(.A1(new_n15619_), .A2(new_n16079_), .ZN(new_n16080_));
  NAND2_X1   g16016(.A1(new_n15510_), .A2(new_n15515_), .ZN(new_n16081_));
  NAND3_X1   g16017(.A1(new_n15580_), .A2(new_n15581_), .A3(new_n15579_), .ZN(new_n16082_));
  OAI21_X1   g16018(.A1(new_n15577_), .A2(new_n15571_), .B(new_n15520_), .ZN(new_n16083_));
  INV_X1     g16019(.I(new_n15593_), .ZN(new_n16084_));
  NAND3_X1   g16020(.A1(new_n15591_), .A2(new_n15592_), .A3(new_n15599_), .ZN(new_n16085_));
  OAI21_X1   g16021(.A1(new_n15595_), .A2(new_n15594_), .B(new_n15589_), .ZN(new_n16086_));
  NOR2_X1    g16022(.A1(new_n15604_), .A2(new_n15605_), .ZN(new_n16087_));
  NOR3_X1    g16023(.A1(new_n16087_), .A2(new_n15550_), .A3(new_n15606_), .ZN(new_n16088_));
  NAND3_X1   g16024(.A1(new_n16086_), .A2(new_n16085_), .A3(new_n16088_), .ZN(new_n16089_));
  NAND2_X1   g16025(.A1(new_n16089_), .A2(new_n16084_), .ZN(new_n16090_));
  AOI22_X1   g16026(.A1(new_n16083_), .A2(new_n16082_), .B1(new_n16090_), .B2(new_n15579_), .ZN(new_n16091_));
  OAI21_X1   g16027(.A1(new_n16091_), .A2(new_n16081_), .B(new_n15510_), .ZN(new_n16092_));
  NAND3_X1   g16028(.A1(new_n16092_), .A2(new_n15497_), .A3(new_n16080_), .ZN(new_n16093_));
  NAND2_X1   g16029(.A1(new_n16093_), .A2(new_n15426_), .ZN(new_n16094_));
  NAND4_X1   g16030(.A1(new_n16092_), .A2(new_n15614_), .A3(new_n16080_), .A4(new_n15497_), .ZN(new_n16095_));
  AOI21_X1   g16031(.A1(new_n16094_), .A2(new_n16095_), .B(new_n15488_), .ZN(new_n16096_));
  INV_X1     g16032(.I(new_n15488_), .ZN(new_n16097_));
  AOI21_X1   g16033(.A1(new_n15613_), .A2(new_n15497_), .B(new_n15614_), .ZN(new_n16098_));
  NOR4_X1    g16034(.A1(new_n15612_), .A2(new_n15426_), .A3(new_n15619_), .A4(new_n15502_), .ZN(new_n16099_));
  NOR3_X1    g16035(.A1(new_n16098_), .A2(new_n16097_), .A3(new_n16099_), .ZN(new_n16100_));
  NOR2_X1    g16036(.A1(new_n16100_), .A2(new_n16096_), .ZN(new_n16101_));
  NAND2_X1   g16037(.A1(new_n15612_), .A2(new_n16080_), .ZN(new_n16102_));
  NAND2_X1   g16038(.A1(new_n16092_), .A2(new_n15502_), .ZN(new_n16103_));
  OAI22_X1   g16039(.A1(new_n8701_), .A2(new_n6783_), .B1(new_n8694_), .B2(new_n6788_), .ZN(new_n16104_));
  NAND2_X1   g16040(.A1(new_n8682_), .A2(new_n6784_), .ZN(new_n16105_));
  AOI21_X1   g16041(.A1(new_n16105_), .A2(new_n16104_), .B(new_n6776_), .ZN(new_n16106_));
  NAND3_X1   g16042(.A1(new_n11611_), .A2(new_n11608_), .A3(new_n16106_), .ZN(new_n16107_));
  NOR2_X1    g16043(.A1(new_n16107_), .A2(\a[8] ), .ZN(new_n16108_));
  INV_X1     g16044(.I(new_n16108_), .ZN(new_n16109_));
  NAND2_X1   g16045(.A1(new_n16107_), .A2(\a[8] ), .ZN(new_n16110_));
  NAND2_X1   g16046(.A1(new_n16109_), .A2(new_n16110_), .ZN(new_n16111_));
  AOI21_X1   g16047(.A1(new_n16102_), .A2(new_n16103_), .B(new_n16111_), .ZN(new_n16112_));
  NOR2_X1    g16048(.A1(new_n16092_), .A2(new_n15502_), .ZN(new_n16113_));
  NOR2_X1    g16049(.A1(new_n15612_), .A2(new_n16080_), .ZN(new_n16114_));
  INV_X1     g16050(.I(new_n16110_), .ZN(new_n16115_));
  NOR2_X1    g16051(.A1(new_n16115_), .A2(new_n16108_), .ZN(new_n16116_));
  NOR3_X1    g16052(.A1(new_n16114_), .A2(new_n16113_), .A3(new_n16116_), .ZN(new_n16117_));
  OAI22_X1   g16053(.A1(new_n6788_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n6783_), .ZN(new_n16118_));
  OAI21_X1   g16054(.A1(new_n6785_), .A2(new_n8694_), .B(new_n16118_), .ZN(new_n16119_));
  NAND4_X1   g16055(.A1(new_n11592_), .A2(new_n6775_), .A3(new_n11594_), .A4(new_n16119_), .ZN(new_n16120_));
  XOR2_X1    g16056(.A1(new_n16120_), .A2(\a[8] ), .Z(new_n16121_));
  NAND2_X1   g16057(.A1(new_n16091_), .A2(new_n15516_), .ZN(new_n16122_));
  NAND2_X1   g16058(.A1(new_n15611_), .A2(new_n16081_), .ZN(new_n16123_));
  NAND2_X1   g16059(.A1(new_n16123_), .A2(new_n16122_), .ZN(new_n16124_));
  NOR2_X1    g16060(.A1(new_n16124_), .A2(new_n16121_), .ZN(new_n16125_));
  NOR3_X1    g16061(.A1(new_n16112_), .A2(new_n16117_), .A3(new_n16125_), .ZN(new_n16126_));
  OAI22_X1   g16062(.A1(new_n8681_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8694_), .ZN(new_n16127_));
  NAND2_X1   g16063(.A1(new_n8688_), .A2(new_n6784_), .ZN(new_n16128_));
  AOI21_X1   g16064(.A1(new_n16128_), .A2(new_n16127_), .B(new_n6776_), .ZN(new_n16129_));
  AND3_X2    g16065(.A1(new_n11420_), .A2(new_n4009_), .A3(new_n16129_), .Z(new_n16130_));
  AOI21_X1   g16066(.A1(new_n11420_), .A2(new_n16129_), .B(new_n4009_), .ZN(new_n16131_));
  NOR2_X1    g16067(.A1(new_n16130_), .A2(new_n16131_), .ZN(new_n16132_));
  INV_X1     g16068(.I(new_n16132_), .ZN(new_n16133_));
  NOR2_X1    g16069(.A1(new_n16126_), .A2(new_n16133_), .ZN(new_n16134_));
  NOR4_X1    g16070(.A1(new_n16112_), .A2(new_n16117_), .A3(new_n16125_), .A4(new_n16132_), .ZN(new_n16135_));
  OAI21_X1   g16071(.A1(new_n16134_), .A2(new_n16135_), .B(new_n16101_), .ZN(new_n16136_));
  OAI21_X1   g16072(.A1(new_n16098_), .A2(new_n16099_), .B(new_n16097_), .ZN(new_n16137_));
  NAND3_X1   g16073(.A1(new_n16094_), .A2(new_n15488_), .A3(new_n16095_), .ZN(new_n16138_));
  NAND2_X1   g16074(.A1(new_n16137_), .A2(new_n16138_), .ZN(new_n16139_));
  OAI21_X1   g16075(.A1(new_n16114_), .A2(new_n16113_), .B(new_n16116_), .ZN(new_n16140_));
  NAND3_X1   g16076(.A1(new_n16102_), .A2(new_n16103_), .A3(new_n16111_), .ZN(new_n16141_));
  INV_X1     g16077(.I(new_n16121_), .ZN(new_n16142_));
  NAND3_X1   g16078(.A1(new_n16142_), .A2(new_n16122_), .A3(new_n16123_), .ZN(new_n16143_));
  NAND3_X1   g16079(.A1(new_n16140_), .A2(new_n16141_), .A3(new_n16143_), .ZN(new_n16144_));
  NAND2_X1   g16080(.A1(new_n16144_), .A2(new_n16132_), .ZN(new_n16145_));
  NAND4_X1   g16081(.A1(new_n16133_), .A2(new_n16140_), .A3(new_n16141_), .A4(new_n16143_), .ZN(new_n16146_));
  NAND3_X1   g16082(.A1(new_n16145_), .A2(new_n16139_), .A3(new_n16146_), .ZN(new_n16147_));
  AOI21_X1   g16083(.A1(new_n16136_), .A2(new_n16147_), .B(new_n16078_), .ZN(new_n16148_));
  INV_X1     g16084(.I(new_n16148_), .ZN(new_n16149_));
  NAND3_X1   g16085(.A1(new_n16140_), .A2(new_n16141_), .A3(new_n16125_), .ZN(new_n16150_));
  INV_X1     g16086(.I(new_n16150_), .ZN(new_n16151_));
  AOI21_X1   g16087(.A1(new_n16140_), .A2(new_n16141_), .B(new_n16125_), .ZN(new_n16152_));
  OAI22_X1   g16088(.A1(new_n8673_), .A2(new_n6843_), .B1(new_n8687_), .B2(new_n6913_), .ZN(new_n16153_));
  NAND2_X1   g16089(.A1(new_n8662_), .A2(new_n6838_), .ZN(new_n16154_));
  AOI21_X1   g16090(.A1(new_n16154_), .A2(new_n16153_), .B(new_n6836_), .ZN(new_n16155_));
  NAND3_X1   g16091(.A1(new_n11624_), .A2(new_n65_), .A3(new_n16155_), .ZN(new_n16156_));
  NAND3_X1   g16092(.A1(new_n10958_), .A2(new_n10959_), .A3(new_n8661_), .ZN(new_n16157_));
  INV_X1     g16093(.I(new_n10956_), .ZN(new_n16158_));
  OAI21_X1   g16094(.A1(new_n11291_), .A2(new_n8673_), .B(new_n16158_), .ZN(new_n16159_));
  OAI21_X1   g16095(.A1(new_n16159_), .A2(new_n10947_), .B(new_n8662_), .ZN(new_n16160_));
  NAND3_X1   g16096(.A1(new_n16160_), .A2(new_n16157_), .A3(new_n16155_), .ZN(new_n16161_));
  NAND2_X1   g16097(.A1(new_n16161_), .A2(\a[5] ), .ZN(new_n16162_));
  NAND2_X1   g16098(.A1(new_n16162_), .A2(new_n16156_), .ZN(new_n16163_));
  NOR3_X1    g16099(.A1(new_n16151_), .A2(new_n16163_), .A3(new_n16152_), .ZN(new_n16164_));
  INV_X1     g16100(.I(new_n16152_), .ZN(new_n16165_));
  XOR2_X1    g16101(.A1(new_n16161_), .A2(\a[5] ), .Z(new_n16166_));
  AOI21_X1   g16102(.A1(new_n16150_), .A2(new_n16165_), .B(new_n16166_), .ZN(new_n16167_));
  NOR2_X1    g16103(.A1(new_n16167_), .A2(new_n16164_), .ZN(new_n16168_));
  NAND2_X1   g16104(.A1(new_n16124_), .A2(new_n16121_), .ZN(new_n16169_));
  NAND3_X1   g16105(.A1(new_n16142_), .A2(new_n16122_), .A3(new_n16123_), .ZN(new_n16170_));
  NAND2_X1   g16106(.A1(new_n16169_), .A2(new_n16170_), .ZN(new_n16171_));
  OAI22_X1   g16107(.A1(new_n6913_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n6843_), .ZN(new_n16172_));
  NAND2_X1   g16108(.A1(new_n8674_), .A2(new_n6838_), .ZN(new_n16173_));
  AOI21_X1   g16109(.A1(new_n16173_), .A2(new_n16172_), .B(new_n6836_), .ZN(new_n16174_));
  NAND3_X1   g16110(.A1(new_n11431_), .A2(new_n65_), .A3(new_n16174_), .ZN(new_n16175_));
  NOR2_X1    g16111(.A1(new_n10946_), .A2(new_n10956_), .ZN(new_n16176_));
  INV_X1     g16112(.I(new_n11430_), .ZN(new_n16177_));
  OAI21_X1   g16113(.A1(new_n16177_), .A2(new_n16176_), .B(new_n16174_), .ZN(new_n16178_));
  NAND2_X1   g16114(.A1(new_n16178_), .A2(\a[5] ), .ZN(new_n16179_));
  NAND3_X1   g16115(.A1(new_n16171_), .A2(new_n16175_), .A3(new_n16179_), .ZN(new_n16180_));
  NAND2_X1   g16116(.A1(new_n16179_), .A2(new_n16175_), .ZN(new_n16181_));
  NAND3_X1   g16117(.A1(new_n16181_), .A2(new_n16169_), .A3(new_n16170_), .ZN(new_n16182_));
  NAND2_X1   g16118(.A1(new_n16180_), .A2(new_n16182_), .ZN(new_n16183_));
  INV_X1     g16119(.I(new_n11418_), .ZN(new_n16184_));
  NOR2_X1    g16120(.A1(new_n10943_), .A2(new_n11419_), .ZN(new_n16185_));
  OAI22_X1   g16121(.A1(new_n8681_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8694_), .ZN(new_n16186_));
  NAND2_X1   g16122(.A1(new_n8688_), .A2(new_n6838_), .ZN(new_n16187_));
  AOI21_X1   g16123(.A1(new_n16187_), .A2(new_n16186_), .B(new_n6836_), .ZN(new_n16188_));
  OAI21_X1   g16124(.A1(new_n16184_), .A2(new_n16185_), .B(new_n16188_), .ZN(new_n16189_));
  XOR2_X1    g16125(.A1(new_n16189_), .A2(\a[5] ), .Z(new_n16190_));
  NOR2_X1    g16126(.A1(new_n15577_), .A2(new_n15571_), .ZN(new_n16191_));
  NOR2_X1    g16127(.A1(new_n15610_), .A2(new_n15579_), .ZN(new_n16192_));
  NOR2_X1    g16128(.A1(new_n16090_), .A2(new_n15520_), .ZN(new_n16193_));
  OAI21_X1   g16129(.A1(new_n16192_), .A2(new_n16193_), .B(new_n16191_), .ZN(new_n16194_));
  INV_X1     g16130(.I(new_n16191_), .ZN(new_n16195_));
  NAND2_X1   g16131(.A1(new_n16090_), .A2(new_n15520_), .ZN(new_n16196_));
  NAND2_X1   g16132(.A1(new_n15610_), .A2(new_n15579_), .ZN(new_n16197_));
  NAND3_X1   g16133(.A1(new_n16197_), .A2(new_n16196_), .A3(new_n16195_), .ZN(new_n16198_));
  NAND2_X1   g16134(.A1(new_n16194_), .A2(new_n16198_), .ZN(new_n16199_));
  AOI21_X1   g16135(.A1(new_n16086_), .A2(new_n16085_), .B(new_n16088_), .ZN(new_n16200_));
  OAI22_X1   g16136(.A1(new_n8725_), .A2(new_n6783_), .B1(new_n6788_), .B2(new_n8718_), .ZN(new_n16201_));
  NAND2_X1   g16137(.A1(new_n8711_), .A2(new_n6784_), .ZN(new_n16202_));
  AOI21_X1   g16138(.A1(new_n16202_), .A2(new_n16201_), .B(new_n6776_), .ZN(new_n16203_));
  NAND3_X1   g16139(.A1(new_n11536_), .A2(new_n4009_), .A3(new_n16203_), .ZN(new_n16204_));
  OAI21_X1   g16140(.A1(new_n15491_), .A2(new_n11532_), .B(new_n16203_), .ZN(new_n16205_));
  NAND2_X1   g16141(.A1(new_n16205_), .A2(\a[8] ), .ZN(new_n16206_));
  NAND2_X1   g16142(.A1(new_n16204_), .A2(new_n16206_), .ZN(new_n16207_));
  INV_X1     g16143(.I(new_n16207_), .ZN(new_n16208_));
  OAI21_X1   g16144(.A1(new_n15609_), .A2(new_n16200_), .B(new_n16208_), .ZN(new_n16209_));
  INV_X1     g16145(.I(new_n16200_), .ZN(new_n16210_));
  NAND3_X1   g16146(.A1(new_n16210_), .A2(new_n16089_), .A3(new_n16207_), .ZN(new_n16211_));
  XNOR2_X1   g16147(.A1(new_n16087_), .A2(new_n15607_), .ZN(new_n16212_));
  OAI22_X1   g16148(.A1(new_n8725_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8735_), .ZN(new_n16213_));
  NAND2_X1   g16149(.A1(new_n8719_), .A2(new_n6784_), .ZN(new_n16214_));
  AOI21_X1   g16150(.A1(new_n16213_), .A2(new_n16214_), .B(new_n6776_), .ZN(new_n16215_));
  NAND2_X1   g16151(.A1(new_n12242_), .A2(new_n16215_), .ZN(new_n16216_));
  XOR2_X1    g16152(.A1(new_n16216_), .A2(new_n4009_), .Z(new_n16217_));
  NAND2_X1   g16153(.A1(new_n16217_), .A2(new_n16212_), .ZN(new_n16218_));
  NAND3_X1   g16154(.A1(new_n16209_), .A2(new_n16211_), .A3(new_n16218_), .ZN(new_n16219_));
  OAI22_X1   g16155(.A1(new_n8710_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8718_), .ZN(new_n16220_));
  NAND2_X1   g16156(.A1(new_n8702_), .A2(new_n6784_), .ZN(new_n16221_));
  AOI21_X1   g16157(.A1(new_n16221_), .A2(new_n16220_), .B(new_n6776_), .ZN(new_n16222_));
  NAND2_X1   g16158(.A1(new_n12205_), .A2(new_n16222_), .ZN(new_n16223_));
  XOR2_X1    g16159(.A1(new_n16223_), .A2(\a[8] ), .Z(new_n16224_));
  NAND2_X1   g16160(.A1(new_n16219_), .A2(new_n16224_), .ZN(new_n16225_));
  AOI21_X1   g16161(.A1(new_n16210_), .A2(new_n16089_), .B(new_n16207_), .ZN(new_n16226_));
  NOR3_X1    g16162(.A1(new_n16208_), .A2(new_n15609_), .A3(new_n16200_), .ZN(new_n16227_));
  INV_X1     g16163(.I(new_n16212_), .ZN(new_n16228_));
  XOR2_X1    g16164(.A1(new_n16216_), .A2(\a[8] ), .Z(new_n16229_));
  NOR2_X1    g16165(.A1(new_n16229_), .A2(new_n16228_), .ZN(new_n16230_));
  NOR3_X1    g16166(.A1(new_n16227_), .A2(new_n16226_), .A3(new_n16230_), .ZN(new_n16231_));
  XOR2_X1    g16167(.A1(new_n16223_), .A2(new_n4009_), .Z(new_n16232_));
  NAND2_X1   g16168(.A1(new_n16231_), .A2(new_n16232_), .ZN(new_n16233_));
  AOI21_X1   g16169(.A1(new_n16225_), .A2(new_n16233_), .B(new_n16199_), .ZN(new_n16234_));
  AOI21_X1   g16170(.A1(new_n16197_), .A2(new_n16196_), .B(new_n16195_), .ZN(new_n16235_));
  NOR3_X1    g16171(.A1(new_n16192_), .A2(new_n16193_), .A3(new_n16191_), .ZN(new_n16236_));
  NOR2_X1    g16172(.A1(new_n16235_), .A2(new_n16236_), .ZN(new_n16237_));
  NOR2_X1    g16173(.A1(new_n16231_), .A2(new_n16232_), .ZN(new_n16238_));
  NOR2_X1    g16174(.A1(new_n16219_), .A2(new_n16224_), .ZN(new_n16239_));
  NOR3_X1    g16175(.A1(new_n16239_), .A2(new_n16238_), .A3(new_n16237_), .ZN(new_n16240_));
  OAI21_X1   g16176(.A1(new_n16240_), .A2(new_n16234_), .B(new_n16190_), .ZN(new_n16241_));
  OAI22_X1   g16177(.A1(new_n8701_), .A2(new_n6913_), .B1(new_n8694_), .B2(new_n6843_), .ZN(new_n16242_));
  NAND2_X1   g16178(.A1(new_n8682_), .A2(new_n6838_), .ZN(new_n16243_));
  AOI21_X1   g16179(.A1(new_n16243_), .A2(new_n16242_), .B(new_n6836_), .ZN(new_n16244_));
  NAND3_X1   g16180(.A1(new_n11611_), .A2(new_n11608_), .A3(new_n16244_), .ZN(new_n16245_));
  NOR2_X1    g16181(.A1(new_n16245_), .A2(\a[5] ), .ZN(new_n16246_));
  INV_X1     g16182(.I(new_n16246_), .ZN(new_n16247_));
  NAND2_X1   g16183(.A1(new_n16245_), .A2(\a[5] ), .ZN(new_n16248_));
  NAND2_X1   g16184(.A1(new_n16247_), .A2(new_n16248_), .ZN(new_n16249_));
  NAND3_X1   g16185(.A1(new_n16209_), .A2(new_n16211_), .A3(new_n16230_), .ZN(new_n16250_));
  INV_X1     g16186(.I(new_n16250_), .ZN(new_n16251_));
  AOI21_X1   g16187(.A1(new_n16209_), .A2(new_n16211_), .B(new_n16230_), .ZN(new_n16252_));
  NOR3_X1    g16188(.A1(new_n16251_), .A2(new_n16249_), .A3(new_n16252_), .ZN(new_n16253_));
  INV_X1     g16189(.I(new_n16248_), .ZN(new_n16254_));
  NOR2_X1    g16190(.A1(new_n16254_), .A2(new_n16246_), .ZN(new_n16255_));
  INV_X1     g16191(.I(new_n16252_), .ZN(new_n16256_));
  AOI21_X1   g16192(.A1(new_n16256_), .A2(new_n16250_), .B(new_n16255_), .ZN(new_n16257_));
  OR2_X2     g16193(.A1(new_n16257_), .A2(new_n16253_), .Z(new_n16258_));
  XOR2_X1    g16194(.A1(new_n16229_), .A2(new_n16228_), .Z(new_n16259_));
  OAI22_X1   g16195(.A1(new_n6843_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n6913_), .ZN(new_n16260_));
  NAND2_X1   g16196(.A1(new_n8696_), .A2(new_n6838_), .ZN(new_n16261_));
  AOI21_X1   g16197(.A1(new_n16260_), .A2(new_n16261_), .B(new_n6836_), .ZN(new_n16262_));
  NAND3_X1   g16198(.A1(new_n11592_), .A2(new_n11594_), .A3(new_n16262_), .ZN(new_n16263_));
  NOR2_X1    g16199(.A1(new_n16263_), .A2(\a[5] ), .ZN(new_n16264_));
  NAND2_X1   g16200(.A1(new_n16263_), .A2(\a[5] ), .ZN(new_n16265_));
  INV_X1     g16201(.I(new_n16265_), .ZN(new_n16266_));
  NOR3_X1    g16202(.A1(new_n16259_), .A2(new_n16266_), .A3(new_n16264_), .ZN(new_n16267_));
  OAI22_X1   g16203(.A1(new_n8751_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8745_), .ZN(new_n16268_));
  NAND2_X1   g16204(.A1(new_n10927_), .A2(new_n6784_), .ZN(new_n16269_));
  AOI21_X1   g16205(.A1(new_n16268_), .A2(new_n16269_), .B(new_n6776_), .ZN(new_n16270_));
  NAND2_X1   g16206(.A1(new_n12072_), .A2(new_n16270_), .ZN(new_n16271_));
  XOR2_X1    g16207(.A1(new_n16271_), .A2(\a[8] ), .Z(new_n16272_));
  INV_X1     g16208(.I(new_n16272_), .ZN(new_n16273_));
  OAI22_X1   g16209(.A1(new_n10871_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8778_), .ZN(new_n16274_));
  NAND2_X1   g16210(.A1(new_n10886_), .A2(new_n6090_), .ZN(new_n16275_));
  AOI21_X1   g16211(.A1(new_n16275_), .A2(new_n16274_), .B(new_n6082_), .ZN(new_n16276_));
  NAND2_X1   g16212(.A1(new_n13103_), .A2(new_n16276_), .ZN(new_n16277_));
  XOR2_X1    g16213(.A1(new_n16277_), .A2(new_n3521_), .Z(new_n16278_));
  AOI21_X1   g16214(.A1(new_n15309_), .A2(new_n15307_), .B(new_n15033_), .ZN(new_n16279_));
  XOR2_X1    g16215(.A1(new_n15046_), .A2(new_n15043_), .Z(new_n16280_));
  NOR2_X1    g16216(.A1(new_n16280_), .A2(new_n15306_), .ZN(new_n16281_));
  NOR2_X1    g16217(.A1(new_n16281_), .A2(new_n16279_), .ZN(new_n16282_));
  NOR2_X1    g16218(.A1(new_n16282_), .A2(new_n16278_), .ZN(new_n16283_));
  INV_X1     g16219(.I(new_n14960_), .ZN(new_n16284_));
  AOI22_X1   g16220(.A1(new_n12823_), .A2(new_n6180_), .B1(new_n6095_), .B2(new_n10800_), .ZN(new_n16285_));
  AOI21_X1   g16221(.A1(new_n6090_), .A2(new_n9529_), .B(new_n16285_), .ZN(new_n16286_));
  OR3_X2     g16222(.A1(new_n13504_), .A2(new_n6082_), .A3(new_n16286_), .Z(new_n16287_));
  XOR2_X1    g16223(.A1(new_n16287_), .A2(new_n3521_), .Z(new_n16288_));
  NAND2_X1   g16224(.A1(new_n16288_), .A2(new_n16284_), .ZN(new_n16289_));
  AOI22_X1   g16225(.A1(new_n10794_), .A2(new_n6180_), .B1(new_n6095_), .B2(new_n12823_), .ZN(new_n16290_));
  AOI21_X1   g16226(.A1(new_n6090_), .A2(new_n10800_), .B(new_n16290_), .ZN(new_n16291_));
  NOR3_X1    g16227(.A1(new_n16291_), .A2(new_n14787_), .A3(new_n6082_), .ZN(new_n16292_));
  XOR2_X1    g16228(.A1(new_n16292_), .A2(\a[14] ), .Z(new_n16293_));
  INV_X1     g16229(.I(new_n16293_), .ZN(new_n16294_));
  NAND2_X1   g16230(.A1(new_n10794_), .A2(new_n6095_), .ZN(new_n16295_));
  NOR2_X1    g16231(.A1(new_n6079_), .A2(new_n6080_), .ZN(new_n16296_));
  NAND3_X1   g16232(.A1(new_n14793_), .A2(new_n16295_), .A3(new_n16296_), .ZN(new_n16297_));
  XOR2_X1    g16233(.A1(new_n16297_), .A2(\a[14] ), .Z(new_n16298_));
  NOR2_X1    g16234(.A1(new_n12826_), .A2(new_n6079_), .ZN(new_n16299_));
  NOR2_X1    g16235(.A1(new_n16299_), .A2(new_n3521_), .ZN(new_n16300_));
  NAND2_X1   g16236(.A1(new_n16298_), .A2(new_n16300_), .ZN(new_n16301_));
  NOR2_X1    g16237(.A1(new_n16294_), .A2(new_n16301_), .ZN(new_n16302_));
  NOR2_X1    g16238(.A1(new_n16288_), .A2(new_n16284_), .ZN(new_n16303_));
  OAI21_X1   g16239(.A1(new_n16302_), .A2(new_n16303_), .B(new_n16289_), .ZN(new_n16304_));
  XOR2_X1    g16240(.A1(new_n14959_), .A2(new_n14962_), .Z(new_n16305_));
  AOI22_X1   g16241(.A1(new_n9529_), .A2(new_n6095_), .B1(new_n10800_), .B2(new_n6180_), .ZN(new_n16306_));
  AOI21_X1   g16242(.A1(new_n10839_), .A2(new_n6090_), .B(new_n16306_), .ZN(new_n16307_));
  OR3_X2     g16243(.A1(new_n13534_), .A2(new_n6082_), .A3(new_n16307_), .Z(new_n16308_));
  XOR2_X1    g16244(.A1(new_n16308_), .A2(\a[14] ), .Z(new_n16309_));
  NAND2_X1   g16245(.A1(new_n16309_), .A2(new_n16305_), .ZN(new_n16310_));
  NOR2_X1    g16246(.A1(new_n16309_), .A2(new_n16305_), .ZN(new_n16311_));
  AOI21_X1   g16247(.A1(new_n16304_), .A2(new_n16310_), .B(new_n16311_), .ZN(new_n16312_));
  AOI22_X1   g16248(.A1(new_n10839_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n9529_), .ZN(new_n16313_));
  NOR2_X1    g16249(.A1(new_n10846_), .A2(new_n6091_), .ZN(new_n16314_));
  OAI21_X1   g16250(.A1(new_n16313_), .A2(new_n16314_), .B(new_n6081_), .ZN(new_n16315_));
  NOR2_X1    g16251(.A1(new_n12946_), .A2(new_n16315_), .ZN(new_n16316_));
  XOR2_X1    g16252(.A1(new_n16316_), .A2(new_n3521_), .Z(new_n16317_));
  NOR2_X1    g16253(.A1(new_n16312_), .A2(new_n16317_), .ZN(new_n16318_));
  INV_X1     g16254(.I(new_n14955_), .ZN(new_n16319_));
  OAI21_X1   g16255(.A1(new_n14959_), .A2(new_n14962_), .B(new_n16319_), .ZN(new_n16320_));
  AOI22_X1   g16256(.A1(new_n16312_), .A2(new_n16317_), .B1(new_n14964_), .B2(new_n16320_), .ZN(new_n16321_));
  NAND2_X1   g16257(.A1(new_n14966_), .A2(new_n14943_), .ZN(new_n16322_));
  NAND2_X1   g16258(.A1(new_n14950_), .A2(new_n14797_), .ZN(new_n16323_));
  AOI21_X1   g16259(.A1(new_n16322_), .A2(new_n16323_), .B(new_n14964_), .ZN(new_n16324_));
  AOI22_X1   g16260(.A1(new_n14967_), .A2(new_n14951_), .B1(new_n14955_), .B2(new_n14963_), .ZN(new_n16325_));
  OR2_X2     g16261(.A1(new_n16325_), .A2(new_n16324_), .Z(new_n16326_));
  AOI22_X1   g16262(.A1(new_n10839_), .A2(new_n6180_), .B1(new_n12936_), .B2(new_n6095_), .ZN(new_n16327_));
  AOI21_X1   g16263(.A1(new_n6090_), .A2(new_n9479_), .B(new_n16327_), .ZN(new_n16328_));
  NOR3_X1    g16264(.A1(new_n12975_), .A2(new_n6082_), .A3(new_n16328_), .ZN(new_n16329_));
  XOR2_X1    g16265(.A1(new_n16329_), .A2(\a[14] ), .Z(new_n16330_));
  OAI22_X1   g16266(.A1(new_n16321_), .A2(new_n16318_), .B1(new_n16326_), .B2(new_n16330_), .ZN(new_n16331_));
  NAND2_X1   g16267(.A1(new_n16326_), .A2(new_n16330_), .ZN(new_n16332_));
  NAND2_X1   g16268(.A1(new_n14976_), .A2(new_n15281_), .ZN(new_n16333_));
  NAND2_X1   g16269(.A1(new_n15282_), .A2(new_n14972_), .ZN(new_n16334_));
  AOI21_X1   g16270(.A1(new_n16334_), .A2(new_n16333_), .B(new_n15280_), .ZN(new_n16335_));
  AOI21_X1   g16271(.A1(new_n15284_), .A2(new_n14977_), .B(new_n14969_), .ZN(new_n16336_));
  NOR2_X1    g16272(.A1(new_n16336_), .A2(new_n16335_), .ZN(new_n16337_));
  OAI22_X1   g16273(.A1(new_n9478_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n10846_), .ZN(new_n16338_));
  NAND2_X1   g16274(.A1(new_n10854_), .A2(new_n6090_), .ZN(new_n16339_));
  AOI21_X1   g16275(.A1(new_n16338_), .A2(new_n16339_), .B(new_n6082_), .ZN(new_n16340_));
  NAND2_X1   g16276(.A1(new_n13016_), .A2(new_n16340_), .ZN(new_n16341_));
  XOR2_X1    g16277(.A1(new_n16341_), .A2(new_n3521_), .Z(new_n16342_));
  NOR2_X1    g16278(.A1(new_n16337_), .A2(new_n16342_), .ZN(new_n16343_));
  AOI21_X1   g16279(.A1(new_n16331_), .A2(new_n16332_), .B(new_n16343_), .ZN(new_n16344_));
  AND2_X2    g16280(.A1(new_n16337_), .A2(new_n16342_), .Z(new_n16345_));
  XOR2_X1    g16281(.A1(new_n14985_), .A2(new_n14990_), .Z(new_n16346_));
  NOR2_X1    g16282(.A1(new_n16346_), .A2(new_n14979_), .ZN(new_n16347_));
  NAND2_X1   g16283(.A1(new_n15287_), .A2(new_n14993_), .ZN(new_n16348_));
  AOI21_X1   g16284(.A1(new_n14979_), .A2(new_n16348_), .B(new_n16347_), .ZN(new_n16349_));
  OAI22_X1   g16285(.A1(new_n9478_), .A2(new_n6089_), .B1(new_n6094_), .B2(new_n10853_), .ZN(new_n16350_));
  NAND2_X1   g16286(.A1(new_n10862_), .A2(new_n6090_), .ZN(new_n16351_));
  AOI21_X1   g16287(.A1(new_n16350_), .A2(new_n16351_), .B(new_n6082_), .ZN(new_n16352_));
  NAND2_X1   g16288(.A1(new_n13484_), .A2(new_n16352_), .ZN(new_n16353_));
  XOR2_X1    g16289(.A1(new_n16353_), .A2(\a[14] ), .Z(new_n16354_));
  INV_X1     g16290(.I(new_n16354_), .ZN(new_n16355_));
  NOR2_X1    g16291(.A1(new_n16349_), .A2(new_n16355_), .ZN(new_n16356_));
  INV_X1     g16292(.I(new_n16356_), .ZN(new_n16357_));
  OAI21_X1   g16293(.A1(new_n16344_), .A2(new_n16345_), .B(new_n16357_), .ZN(new_n16358_));
  NAND2_X1   g16294(.A1(new_n16349_), .A2(new_n16355_), .ZN(new_n16359_));
  XOR2_X1    g16295(.A1(new_n15292_), .A2(new_n14999_), .Z(new_n16360_));
  OAI21_X1   g16296(.A1(new_n15290_), .A2(new_n15006_), .B(new_n15289_), .ZN(new_n16361_));
  OAI21_X1   g16297(.A1(new_n15289_), .A2(new_n16360_), .B(new_n16361_), .ZN(new_n16362_));
  OAI22_X1   g16298(.A1(new_n10861_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n10853_), .ZN(new_n16363_));
  NAND2_X1   g16299(.A1(new_n8785_), .A2(new_n6090_), .ZN(new_n16364_));
  AOI21_X1   g16300(.A1(new_n16364_), .A2(new_n16363_), .B(new_n6082_), .ZN(new_n16365_));
  NAND2_X1   g16301(.A1(new_n13592_), .A2(new_n16365_), .ZN(new_n16366_));
  XOR2_X1    g16302(.A1(new_n16366_), .A2(\a[14] ), .Z(new_n16367_));
  NAND2_X1   g16303(.A1(new_n16362_), .A2(new_n16367_), .ZN(new_n16368_));
  INV_X1     g16304(.I(new_n16368_), .ZN(new_n16369_));
  AOI21_X1   g16305(.A1(new_n16358_), .A2(new_n16359_), .B(new_n16369_), .ZN(new_n16370_));
  NOR2_X1    g16306(.A1(new_n16362_), .A2(new_n16367_), .ZN(new_n16371_));
  XOR2_X1    g16307(.A1(new_n15300_), .A2(new_n15014_), .Z(new_n16372_));
  NOR2_X1    g16308(.A1(new_n16372_), .A2(new_n15007_), .ZN(new_n16373_));
  AOI21_X1   g16309(.A1(new_n15301_), .A2(new_n15021_), .B(new_n15294_), .ZN(new_n16374_));
  OAI22_X1   g16310(.A1(new_n8784_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n10861_), .ZN(new_n16375_));
  NAND2_X1   g16311(.A1(new_n8779_), .A2(new_n6090_), .ZN(new_n16376_));
  AOI21_X1   g16312(.A1(new_n16376_), .A2(new_n16375_), .B(new_n6082_), .ZN(new_n16377_));
  NAND2_X1   g16313(.A1(new_n12814_), .A2(new_n16377_), .ZN(new_n16378_));
  XOR2_X1    g16314(.A1(new_n16378_), .A2(\a[14] ), .Z(new_n16379_));
  OAI21_X1   g16315(.A1(new_n16373_), .A2(new_n16374_), .B(new_n16379_), .ZN(new_n16380_));
  OAI21_X1   g16316(.A1(new_n16370_), .A2(new_n16371_), .B(new_n16380_), .ZN(new_n16381_));
  NOR2_X1    g16317(.A1(new_n16373_), .A2(new_n16374_), .ZN(new_n16382_));
  INV_X1     g16318(.I(new_n16379_), .ZN(new_n16383_));
  NAND2_X1   g16319(.A1(new_n16382_), .A2(new_n16383_), .ZN(new_n16384_));
  OAI21_X1   g16320(.A1(new_n15304_), .A2(new_n15032_), .B(new_n15022_), .ZN(new_n16385_));
  INV_X1     g16321(.I(new_n16385_), .ZN(new_n16386_));
  NOR2_X1    g16322(.A1(new_n15024_), .A2(new_n15025_), .ZN(new_n16387_));
  XOR2_X1    g16323(.A1(new_n16387_), .A2(new_n15030_), .Z(new_n16388_));
  NOR2_X1    g16324(.A1(new_n16388_), .A2(new_n15022_), .ZN(new_n16389_));
  AOI22_X1   g16325(.A1(new_n8779_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n8785_), .ZN(new_n16390_));
  NOR2_X1    g16326(.A1(new_n10871_), .A2(new_n6091_), .ZN(new_n16391_));
  OAI21_X1   g16327(.A1(new_n16391_), .A2(new_n16390_), .B(new_n6081_), .ZN(new_n16392_));
  NOR2_X1    g16328(.A1(new_n11794_), .A2(new_n16392_), .ZN(new_n16393_));
  XOR2_X1    g16329(.A1(new_n16393_), .A2(\a[14] ), .Z(new_n16394_));
  NOR3_X1    g16330(.A1(new_n16386_), .A2(new_n16389_), .A3(new_n16394_), .ZN(new_n16395_));
  XNOR2_X1   g16331(.A1(new_n16387_), .A2(new_n15030_), .ZN(new_n16396_));
  NAND2_X1   g16332(.A1(new_n16396_), .A2(new_n15303_), .ZN(new_n16397_));
  XOR2_X1    g16333(.A1(new_n16393_), .A2(new_n3521_), .Z(new_n16398_));
  AOI21_X1   g16334(.A1(new_n16397_), .A2(new_n16385_), .B(new_n16398_), .ZN(new_n16399_));
  NOR2_X1    g16335(.A1(new_n16395_), .A2(new_n16399_), .ZN(new_n16400_));
  NAND3_X1   g16336(.A1(new_n16381_), .A2(new_n16400_), .A3(new_n16384_), .ZN(new_n16401_));
  OAI21_X1   g16337(.A1(new_n15044_), .A2(new_n15048_), .B(new_n15306_), .ZN(new_n16402_));
  XOR2_X1    g16338(.A1(new_n15046_), .A2(new_n15047_), .Z(new_n16403_));
  NAND2_X1   g16339(.A1(new_n16403_), .A2(new_n15033_), .ZN(new_n16404_));
  NAND3_X1   g16340(.A1(new_n16404_), .A2(new_n16278_), .A3(new_n16402_), .ZN(new_n16405_));
  XOR2_X1    g16341(.A1(new_n16277_), .A2(\a[14] ), .Z(new_n16406_));
  OAI21_X1   g16342(.A1(new_n16281_), .A2(new_n16279_), .B(new_n16406_), .ZN(new_n16407_));
  AOI21_X1   g16343(.A1(new_n16407_), .A2(new_n16405_), .B(new_n16395_), .ZN(new_n16408_));
  AOI21_X1   g16344(.A1(new_n16401_), .A2(new_n16408_), .B(new_n16283_), .ZN(new_n16409_));
  XOR2_X1    g16345(.A1(new_n14941_), .A2(new_n14935_), .Z(new_n16410_));
  OAI21_X1   g16346(.A1(new_n15045_), .A2(new_n15048_), .B(new_n16410_), .ZN(new_n16411_));
  NOR2_X1    g16347(.A1(new_n15045_), .A2(new_n15048_), .ZN(new_n16412_));
  NOR2_X1    g16348(.A1(new_n14941_), .A2(new_n14935_), .ZN(new_n16413_));
  OAI21_X1   g16349(.A1(new_n15278_), .A2(new_n16413_), .B(new_n16412_), .ZN(new_n16414_));
  AOI22_X1   g16350(.A1(new_n10886_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n10872_), .ZN(new_n16415_));
  NOR2_X1    g16351(.A1(new_n10892_), .A2(new_n6091_), .ZN(new_n16416_));
  OAI21_X1   g16352(.A1(new_n16415_), .A2(new_n16416_), .B(new_n6081_), .ZN(new_n16417_));
  NOR2_X1    g16353(.A1(new_n12776_), .A2(new_n16417_), .ZN(new_n16418_));
  XOR2_X1    g16354(.A1(new_n16418_), .A2(\a[14] ), .Z(new_n16419_));
  AOI21_X1   g16355(.A1(new_n16411_), .A2(new_n16414_), .B(new_n16419_), .ZN(new_n16420_));
  NAND3_X1   g16356(.A1(new_n16419_), .A2(new_n16411_), .A3(new_n16414_), .ZN(new_n16421_));
  OAI21_X1   g16357(.A1(new_n16409_), .A2(new_n16420_), .B(new_n16421_), .ZN(new_n16422_));
  NAND2_X1   g16358(.A1(new_n16412_), .A2(new_n14941_), .ZN(new_n16423_));
  NAND3_X1   g16359(.A1(new_n16423_), .A2(new_n15312_), .A3(new_n15274_), .ZN(new_n16424_));
  AOI21_X1   g16360(.A1(new_n16423_), .A2(new_n15274_), .B(new_n15312_), .ZN(new_n16425_));
  INV_X1     g16361(.I(new_n16425_), .ZN(new_n16426_));
  AOI22_X1   g16362(.A1(new_n10886_), .A2(new_n6180_), .B1(new_n10889_), .B2(new_n6095_), .ZN(new_n16427_));
  NOR2_X1    g16363(.A1(new_n10899_), .A2(new_n6091_), .ZN(new_n16428_));
  OAI21_X1   g16364(.A1(new_n16428_), .A2(new_n16427_), .B(new_n6081_), .ZN(new_n16429_));
  NOR2_X1    g16365(.A1(new_n11908_), .A2(new_n16429_), .ZN(new_n16430_));
  XOR2_X1    g16366(.A1(new_n16430_), .A2(\a[14] ), .Z(new_n16431_));
  AOI21_X1   g16367(.A1(new_n16426_), .A2(new_n16424_), .B(new_n16431_), .ZN(new_n16432_));
  INV_X1     g16368(.I(new_n16424_), .ZN(new_n16433_));
  XOR2_X1    g16369(.A1(new_n16430_), .A2(new_n3521_), .Z(new_n16434_));
  NOR3_X1    g16370(.A1(new_n16433_), .A2(new_n16434_), .A3(new_n16425_), .ZN(new_n16435_));
  OAI21_X1   g16371(.A1(new_n16432_), .A2(new_n16435_), .B(new_n16422_), .ZN(new_n16436_));
  NOR2_X1    g16372(.A1(new_n16344_), .A2(new_n16345_), .ZN(new_n16437_));
  NOR2_X1    g16373(.A1(new_n16437_), .A2(new_n16356_), .ZN(new_n16438_));
  INV_X1     g16374(.I(new_n16359_), .ZN(new_n16439_));
  OAI21_X1   g16375(.A1(new_n16438_), .A2(new_n16439_), .B(new_n16368_), .ZN(new_n16440_));
  INV_X1     g16376(.I(new_n16371_), .ZN(new_n16441_));
  INV_X1     g16377(.I(new_n16380_), .ZN(new_n16442_));
  AOI21_X1   g16378(.A1(new_n16440_), .A2(new_n16441_), .B(new_n16442_), .ZN(new_n16443_));
  INV_X1     g16379(.I(new_n16384_), .ZN(new_n16444_));
  NAND3_X1   g16380(.A1(new_n16397_), .A2(new_n16398_), .A3(new_n16385_), .ZN(new_n16445_));
  OAI21_X1   g16381(.A1(new_n16386_), .A2(new_n16389_), .B(new_n16394_), .ZN(new_n16446_));
  NAND2_X1   g16382(.A1(new_n16446_), .A2(new_n16445_), .ZN(new_n16447_));
  NOR3_X1    g16383(.A1(new_n16443_), .A2(new_n16447_), .A3(new_n16444_), .ZN(new_n16448_));
  NOR3_X1    g16384(.A1(new_n16281_), .A2(new_n16406_), .A3(new_n16279_), .ZN(new_n16449_));
  AOI21_X1   g16385(.A1(new_n16404_), .A2(new_n16402_), .B(new_n16278_), .ZN(new_n16450_));
  OAI21_X1   g16386(.A1(new_n16449_), .A2(new_n16450_), .B(new_n16445_), .ZN(new_n16451_));
  OAI22_X1   g16387(.A1(new_n16448_), .A2(new_n16451_), .B1(new_n16278_), .B2(new_n16282_), .ZN(new_n16452_));
  INV_X1     g16388(.I(new_n16420_), .ZN(new_n16453_));
  INV_X1     g16389(.I(new_n16421_), .ZN(new_n16454_));
  AOI21_X1   g16390(.A1(new_n16452_), .A2(new_n16453_), .B(new_n16454_), .ZN(new_n16455_));
  NOR3_X1    g16391(.A1(new_n16433_), .A2(new_n16431_), .A3(new_n16425_), .ZN(new_n16456_));
  AOI21_X1   g16392(.A1(new_n16426_), .A2(new_n16424_), .B(new_n16434_), .ZN(new_n16457_));
  OAI21_X1   g16393(.A1(new_n16456_), .A2(new_n16457_), .B(new_n16455_), .ZN(new_n16458_));
  AOI22_X1   g16394(.A1(new_n6480_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n4720_), .ZN(new_n16459_));
  NOR2_X1    g16395(.A1(new_n8758_), .A2(new_n4710_), .ZN(new_n16460_));
  OAI21_X1   g16396(.A1(new_n16459_), .A2(new_n16460_), .B(new_n4706_), .ZN(new_n16461_));
  NOR2_X1    g16397(.A1(new_n12053_), .A2(new_n16461_), .ZN(new_n16462_));
  XOR2_X1    g16398(.A1(new_n16462_), .A2(new_n4034_), .Z(new_n16463_));
  NAND3_X1   g16399(.A1(new_n16458_), .A2(new_n16436_), .A3(new_n16463_), .ZN(new_n16464_));
  AOI21_X1   g16400(.A1(new_n16458_), .A2(new_n16436_), .B(new_n16463_), .ZN(new_n16465_));
  INV_X1     g16401(.I(new_n16465_), .ZN(new_n16466_));
  NAND2_X1   g16402(.A1(new_n16466_), .A2(new_n16464_), .ZN(new_n16467_));
  XOR2_X1    g16403(.A1(new_n16467_), .A2(new_n16273_), .Z(new_n16468_));
  OAI22_X1   g16404(.A1(new_n8725_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8735_), .ZN(new_n16469_));
  NAND2_X1   g16405(.A1(new_n8719_), .A2(new_n6838_), .ZN(new_n16470_));
  AOI21_X1   g16406(.A1(new_n16469_), .A2(new_n16470_), .B(new_n6836_), .ZN(new_n16471_));
  NAND2_X1   g16407(.A1(new_n12242_), .A2(new_n16471_), .ZN(new_n16472_));
  XOR2_X1    g16408(.A1(new_n16472_), .A2(\a[5] ), .Z(new_n16473_));
  NOR2_X1    g16409(.A1(new_n16473_), .A2(new_n16468_), .ZN(new_n16474_));
  INV_X1     g16410(.I(new_n16435_), .ZN(new_n16475_));
  OAI21_X1   g16411(.A1(new_n16455_), .A2(new_n16432_), .B(new_n16475_), .ZN(new_n16476_));
  NOR2_X1    g16412(.A1(new_n14894_), .A2(new_n14927_), .ZN(new_n16477_));
  AOI21_X1   g16413(.A1(new_n15076_), .A2(new_n15064_), .B(new_n15077_), .ZN(new_n16478_));
  NAND3_X1   g16414(.A1(new_n15076_), .A2(new_n15077_), .A3(new_n15064_), .ZN(new_n16479_));
  INV_X1     g16415(.I(new_n16479_), .ZN(new_n16480_));
  OAI21_X1   g16416(.A1(new_n16480_), .A2(new_n16478_), .B(new_n16477_), .ZN(new_n16481_));
  INV_X1     g16417(.I(new_n16477_), .ZN(new_n16482_));
  INV_X1     g16418(.I(new_n16478_), .ZN(new_n16483_));
  NAND3_X1   g16419(.A1(new_n16483_), .A2(new_n16482_), .A3(new_n16479_), .ZN(new_n16484_));
  AOI22_X1   g16420(.A1(new_n11899_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n10889_), .ZN(new_n16485_));
  NOR2_X1    g16421(.A1(new_n8774_), .A2(new_n6091_), .ZN(new_n16486_));
  OAI21_X1   g16422(.A1(new_n16486_), .A2(new_n16485_), .B(new_n6081_), .ZN(new_n16487_));
  NOR2_X1    g16423(.A1(new_n11945_), .A2(new_n16487_), .ZN(new_n16488_));
  XOR2_X1    g16424(.A1(new_n16488_), .A2(\a[14] ), .Z(new_n16489_));
  NAND3_X1   g16425(.A1(new_n16484_), .A2(new_n16481_), .A3(new_n16489_), .ZN(new_n16490_));
  AOI21_X1   g16426(.A1(new_n16483_), .A2(new_n16479_), .B(new_n16482_), .ZN(new_n16491_));
  NOR3_X1    g16427(.A1(new_n16480_), .A2(new_n16477_), .A3(new_n16478_), .ZN(new_n16492_));
  XOR2_X1    g16428(.A1(new_n16488_), .A2(new_n3521_), .Z(new_n16493_));
  OAI21_X1   g16429(.A1(new_n16491_), .A2(new_n16492_), .B(new_n16493_), .ZN(new_n16494_));
  NAND2_X1   g16430(.A1(new_n16494_), .A2(new_n16490_), .ZN(new_n16495_));
  NOR2_X1    g16431(.A1(new_n16495_), .A2(new_n16476_), .ZN(new_n16496_));
  INV_X1     g16432(.I(new_n16432_), .ZN(new_n16497_));
  AOI21_X1   g16433(.A1(new_n16422_), .A2(new_n16497_), .B(new_n16435_), .ZN(new_n16498_));
  AOI21_X1   g16434(.A1(new_n16490_), .A2(new_n16494_), .B(new_n16498_), .ZN(new_n16499_));
  OAI22_X1   g16435(.A1(new_n8758_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8766_), .ZN(new_n16500_));
  NAND2_X1   g16436(.A1(new_n8746_), .A2(new_n4709_), .ZN(new_n16501_));
  AOI21_X1   g16437(.A1(new_n16501_), .A2(new_n16500_), .B(new_n4707_), .ZN(new_n16502_));
  NAND2_X1   g16438(.A1(new_n11964_), .A2(new_n16502_), .ZN(new_n16503_));
  XOR2_X1    g16439(.A1(new_n16503_), .A2(\a[11] ), .Z(new_n16504_));
  INV_X1     g16440(.I(new_n16504_), .ZN(new_n16505_));
  NOR3_X1    g16441(.A1(new_n16496_), .A2(new_n16499_), .A3(new_n16505_), .ZN(new_n16506_));
  NAND3_X1   g16442(.A1(new_n16498_), .A2(new_n16490_), .A3(new_n16494_), .ZN(new_n16507_));
  NAND2_X1   g16443(.A1(new_n16495_), .A2(new_n16476_), .ZN(new_n16508_));
  AOI21_X1   g16444(.A1(new_n16508_), .A2(new_n16507_), .B(new_n16504_), .ZN(new_n16509_));
  OAI21_X1   g16445(.A1(new_n16506_), .A2(new_n16509_), .B(new_n16466_), .ZN(new_n16510_));
  NAND3_X1   g16446(.A1(new_n16508_), .A2(new_n16507_), .A3(new_n16504_), .ZN(new_n16511_));
  OAI21_X1   g16447(.A1(new_n16496_), .A2(new_n16499_), .B(new_n16505_), .ZN(new_n16512_));
  NAND3_X1   g16448(.A1(new_n16512_), .A2(new_n16511_), .A3(new_n16465_), .ZN(new_n16513_));
  OAI22_X1   g16449(.A1(new_n8751_), .A2(new_n6783_), .B1(new_n6788_), .B2(new_n10924_), .ZN(new_n16514_));
  NAND2_X1   g16450(.A1(new_n8736_), .A2(new_n6784_), .ZN(new_n16515_));
  AOI21_X1   g16451(.A1(new_n16515_), .A2(new_n16514_), .B(new_n6776_), .ZN(new_n16516_));
  NAND2_X1   g16452(.A1(new_n12118_), .A2(new_n16516_), .ZN(new_n16517_));
  XOR2_X1    g16453(.A1(new_n16517_), .A2(new_n4009_), .Z(new_n16518_));
  NAND3_X1   g16454(.A1(new_n16510_), .A2(new_n16513_), .A3(new_n16518_), .ZN(new_n16519_));
  AOI21_X1   g16455(.A1(new_n16512_), .A2(new_n16511_), .B(new_n16465_), .ZN(new_n16520_));
  NOR3_X1    g16456(.A1(new_n16506_), .A2(new_n16509_), .A3(new_n16466_), .ZN(new_n16521_));
  XOR2_X1    g16457(.A1(new_n16517_), .A2(\a[8] ), .Z(new_n16522_));
  OAI21_X1   g16458(.A1(new_n16520_), .A2(new_n16521_), .B(new_n16522_), .ZN(new_n16523_));
  NOR2_X1    g16459(.A1(new_n16467_), .A2(new_n16272_), .ZN(new_n16524_));
  NAND3_X1   g16460(.A1(new_n16523_), .A2(new_n16519_), .A3(new_n16524_), .ZN(new_n16525_));
  NOR3_X1    g16461(.A1(new_n16520_), .A2(new_n16521_), .A3(new_n16522_), .ZN(new_n16526_));
  AOI21_X1   g16462(.A1(new_n16510_), .A2(new_n16513_), .B(new_n16518_), .ZN(new_n16527_));
  INV_X1     g16463(.I(new_n16524_), .ZN(new_n16528_));
  OAI21_X1   g16464(.A1(new_n16526_), .A2(new_n16527_), .B(new_n16528_), .ZN(new_n16529_));
  OAI22_X1   g16465(.A1(new_n8725_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n8718_), .ZN(new_n16530_));
  NAND2_X1   g16466(.A1(new_n8711_), .A2(new_n6838_), .ZN(new_n16531_));
  AOI21_X1   g16467(.A1(new_n16531_), .A2(new_n16530_), .B(new_n6836_), .ZN(new_n16532_));
  NAND2_X1   g16468(.A1(new_n11536_), .A2(new_n16532_), .ZN(new_n16533_));
  XOR2_X1    g16469(.A1(new_n16533_), .A2(\a[5] ), .Z(new_n16534_));
  NAND3_X1   g16470(.A1(new_n16534_), .A2(new_n16529_), .A3(new_n16525_), .ZN(new_n16535_));
  NAND2_X1   g16471(.A1(new_n16535_), .A2(new_n16474_), .ZN(new_n16536_));
  NAND2_X1   g16472(.A1(new_n16529_), .A2(new_n16525_), .ZN(new_n16537_));
  XOR2_X1    g16473(.A1(new_n16533_), .A2(new_n65_), .Z(new_n16538_));
  NAND2_X1   g16474(.A1(new_n16537_), .A2(new_n16538_), .ZN(new_n16539_));
  NAND2_X1   g16475(.A1(new_n15112_), .A2(new_n15118_), .ZN(new_n16540_));
  XOR2_X1    g16476(.A1(new_n16540_), .A2(new_n15123_), .Z(new_n16541_));
  NOR2_X1    g16477(.A1(new_n16541_), .A2(new_n15088_), .ZN(new_n16542_));
  NOR2_X1    g16478(.A1(new_n15124_), .A2(new_n15323_), .ZN(new_n16543_));
  INV_X1     g16479(.I(new_n16543_), .ZN(new_n16544_));
  AOI21_X1   g16480(.A1(new_n15088_), .A2(new_n16544_), .B(new_n16542_), .ZN(new_n16545_));
  AOI21_X1   g16481(.A1(new_n16484_), .A2(new_n16481_), .B(new_n16489_), .ZN(new_n16546_));
  AOI21_X1   g16482(.A1(new_n16498_), .A2(new_n16490_), .B(new_n16546_), .ZN(new_n16547_));
  OAI22_X1   g16483(.A1(new_n8774_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n10899_), .ZN(new_n16548_));
  NAND2_X1   g16484(.A1(new_n11996_), .A2(new_n6090_), .ZN(new_n16549_));
  AOI21_X1   g16485(.A1(new_n16549_), .A2(new_n16548_), .B(new_n6082_), .ZN(new_n16550_));
  NAND2_X1   g16486(.A1(new_n12001_), .A2(new_n16550_), .ZN(new_n16551_));
  XOR2_X1    g16487(.A1(new_n16551_), .A2(\a[14] ), .Z(new_n16552_));
  INV_X1     g16488(.I(new_n16552_), .ZN(new_n16553_));
  NOR2_X1    g16489(.A1(new_n16547_), .A2(new_n16553_), .ZN(new_n16554_));
  INV_X1     g16490(.I(new_n16490_), .ZN(new_n16555_));
  OAI21_X1   g16491(.A1(new_n16476_), .A2(new_n16555_), .B(new_n16494_), .ZN(new_n16556_));
  NOR2_X1    g16492(.A1(new_n16556_), .A2(new_n16552_), .ZN(new_n16557_));
  OAI21_X1   g16493(.A1(new_n16557_), .A2(new_n16554_), .B(new_n16545_), .ZN(new_n16558_));
  INV_X1     g16494(.I(new_n16545_), .ZN(new_n16559_));
  NAND2_X1   g16495(.A1(new_n16556_), .A2(new_n16552_), .ZN(new_n16560_));
  NAND2_X1   g16496(.A1(new_n16547_), .A2(new_n16553_), .ZN(new_n16561_));
  NAND3_X1   g16497(.A1(new_n16560_), .A2(new_n16561_), .A3(new_n16559_), .ZN(new_n16562_));
  NAND2_X1   g16498(.A1(new_n16558_), .A2(new_n16562_), .ZN(new_n16563_));
  OAI21_X1   g16499(.A1(new_n16465_), .A2(new_n16509_), .B(new_n16511_), .ZN(new_n16564_));
  OAI22_X1   g16500(.A1(new_n8745_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8758_), .ZN(new_n16565_));
  NAND2_X1   g16501(.A1(new_n8752_), .A2(new_n4709_), .ZN(new_n16566_));
  AOI21_X1   g16502(.A1(new_n16566_), .A2(new_n16565_), .B(new_n4707_), .ZN(new_n16567_));
  NAND2_X1   g16503(.A1(new_n12189_), .A2(new_n16567_), .ZN(new_n16568_));
  XOR2_X1    g16504(.A1(new_n16568_), .A2(\a[11] ), .Z(new_n16569_));
  NAND2_X1   g16505(.A1(new_n16564_), .A2(new_n16569_), .ZN(new_n16570_));
  NAND3_X1   g16506(.A1(new_n16512_), .A2(new_n16511_), .A3(new_n16466_), .ZN(new_n16571_));
  INV_X1     g16507(.I(new_n16569_), .ZN(new_n16572_));
  NAND3_X1   g16508(.A1(new_n16571_), .A2(new_n16511_), .A3(new_n16572_), .ZN(new_n16573_));
  AOI21_X1   g16509(.A1(new_n16573_), .A2(new_n16570_), .B(new_n16563_), .ZN(new_n16574_));
  AOI21_X1   g16510(.A1(new_n16560_), .A2(new_n16561_), .B(new_n16559_), .ZN(new_n16575_));
  NOR3_X1    g16511(.A1(new_n16557_), .A2(new_n16554_), .A3(new_n16545_), .ZN(new_n16576_));
  NOR2_X1    g16512(.A1(new_n16576_), .A2(new_n16575_), .ZN(new_n16577_));
  AOI21_X1   g16513(.A1(new_n16571_), .A2(new_n16511_), .B(new_n16572_), .ZN(new_n16578_));
  NOR2_X1    g16514(.A1(new_n16564_), .A2(new_n16569_), .ZN(new_n16579_));
  NOR3_X1    g16515(.A1(new_n16578_), .A2(new_n16579_), .A3(new_n16577_), .ZN(new_n16580_));
  NOR2_X1    g16516(.A1(new_n16574_), .A2(new_n16580_), .ZN(new_n16581_));
  NOR3_X1    g16517(.A1(new_n16526_), .A2(new_n16527_), .A3(new_n16524_), .ZN(new_n16582_));
  OAI22_X1   g16518(.A1(new_n8735_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n10924_), .ZN(new_n16583_));
  NAND2_X1   g16519(.A1(new_n8726_), .A2(new_n6784_), .ZN(new_n16584_));
  AOI21_X1   g16520(.A1(new_n16584_), .A2(new_n16583_), .B(new_n6776_), .ZN(new_n16585_));
  NAND2_X1   g16521(.A1(new_n12181_), .A2(new_n16585_), .ZN(new_n16586_));
  XOR2_X1    g16522(.A1(new_n16586_), .A2(\a[8] ), .Z(new_n16587_));
  INV_X1     g16523(.I(new_n16587_), .ZN(new_n16588_));
  NOR2_X1    g16524(.A1(new_n16582_), .A2(new_n16588_), .ZN(new_n16589_));
  NOR4_X1    g16525(.A1(new_n16526_), .A2(new_n16527_), .A3(new_n16587_), .A4(new_n16524_), .ZN(new_n16590_));
  OAI21_X1   g16526(.A1(new_n16589_), .A2(new_n16590_), .B(new_n16581_), .ZN(new_n16591_));
  OAI21_X1   g16527(.A1(new_n16578_), .A2(new_n16579_), .B(new_n16577_), .ZN(new_n16592_));
  NAND3_X1   g16528(.A1(new_n16573_), .A2(new_n16570_), .A3(new_n16563_), .ZN(new_n16593_));
  NAND2_X1   g16529(.A1(new_n16592_), .A2(new_n16593_), .ZN(new_n16594_));
  NAND3_X1   g16530(.A1(new_n16523_), .A2(new_n16519_), .A3(new_n16528_), .ZN(new_n16595_));
  NAND2_X1   g16531(.A1(new_n16595_), .A2(new_n16587_), .ZN(new_n16596_));
  INV_X1     g16532(.I(new_n16590_), .ZN(new_n16597_));
  NAND3_X1   g16533(.A1(new_n16597_), .A2(new_n16596_), .A3(new_n16594_), .ZN(new_n16598_));
  NAND2_X1   g16534(.A1(new_n16591_), .A2(new_n16598_), .ZN(new_n16599_));
  OAI22_X1   g16535(.A1(new_n8710_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8718_), .ZN(new_n16600_));
  NAND2_X1   g16536(.A1(new_n8702_), .A2(new_n6838_), .ZN(new_n16601_));
  AOI21_X1   g16537(.A1(new_n16601_), .A2(new_n16600_), .B(new_n6836_), .ZN(new_n16602_));
  NAND2_X1   g16538(.A1(new_n12205_), .A2(new_n16602_), .ZN(new_n16603_));
  XOR2_X1    g16539(.A1(new_n16603_), .A2(\a[5] ), .Z(new_n16604_));
  AOI22_X1   g16540(.A1(new_n16599_), .A2(new_n16604_), .B1(new_n16536_), .B2(new_n16539_), .ZN(new_n16605_));
  NOR2_X1    g16541(.A1(new_n16599_), .A2(new_n16604_), .ZN(new_n16606_));
  XOR2_X1    g16542(.A1(new_n16229_), .A2(new_n16212_), .Z(new_n16607_));
  INV_X1     g16543(.I(new_n16264_), .ZN(new_n16608_));
  NAND3_X1   g16544(.A1(new_n16607_), .A2(new_n16608_), .A3(new_n16265_), .ZN(new_n16609_));
  OAI21_X1   g16545(.A1(new_n16264_), .A2(new_n16266_), .B(new_n16259_), .ZN(new_n16610_));
  NAND2_X1   g16546(.A1(new_n16610_), .A2(new_n16609_), .ZN(new_n16611_));
  NOR3_X1    g16547(.A1(new_n16605_), .A2(new_n16606_), .A3(new_n16611_), .ZN(new_n16612_));
  NOR3_X1    g16548(.A1(new_n16612_), .A2(new_n16258_), .A3(new_n16267_), .ZN(new_n16613_));
  NOR3_X1    g16549(.A1(new_n16190_), .A2(new_n16240_), .A3(new_n16234_), .ZN(new_n16614_));
  NAND3_X1   g16550(.A1(new_n11420_), .A2(new_n65_), .A3(new_n16188_), .ZN(new_n16615_));
  NAND2_X1   g16551(.A1(new_n16189_), .A2(\a[5] ), .ZN(new_n16616_));
  NAND2_X1   g16552(.A1(new_n16616_), .A2(new_n16615_), .ZN(new_n16617_));
  OAI21_X1   g16553(.A1(new_n16239_), .A2(new_n16238_), .B(new_n16237_), .ZN(new_n16618_));
  NAND3_X1   g16554(.A1(new_n16225_), .A2(new_n16233_), .A3(new_n16199_), .ZN(new_n16619_));
  AOI21_X1   g16555(.A1(new_n16618_), .A2(new_n16619_), .B(new_n16617_), .ZN(new_n16620_));
  AOI21_X1   g16556(.A1(new_n16256_), .A2(new_n16250_), .B(new_n16249_), .ZN(new_n16621_));
  INV_X1     g16557(.I(new_n16621_), .ZN(new_n16622_));
  OAI21_X1   g16558(.A1(new_n16614_), .A2(new_n16620_), .B(new_n16622_), .ZN(new_n16623_));
  OAI21_X1   g16559(.A1(new_n16613_), .A2(new_n16623_), .B(new_n16241_), .ZN(new_n16624_));
  OAI21_X1   g16560(.A1(new_n16624_), .A2(new_n16183_), .B(new_n16180_), .ZN(new_n16625_));
  NAND2_X1   g16561(.A1(new_n16625_), .A2(new_n16168_), .ZN(new_n16626_));
  XOR2_X1    g16562(.A1(new_n16077_), .A2(\a[5] ), .Z(new_n16627_));
  AOI21_X1   g16563(.A1(new_n16145_), .A2(new_n16146_), .B(new_n16139_), .ZN(new_n16628_));
  NOR3_X1    g16564(.A1(new_n16134_), .A2(new_n16101_), .A3(new_n16135_), .ZN(new_n16629_));
  NOR3_X1    g16565(.A1(new_n16628_), .A2(new_n16629_), .A3(new_n16627_), .ZN(new_n16630_));
  AOI21_X1   g16566(.A1(new_n16136_), .A2(new_n16147_), .B(new_n16078_), .ZN(new_n16631_));
  NAND3_X1   g16567(.A1(new_n16166_), .A2(new_n16150_), .A3(new_n16165_), .ZN(new_n16632_));
  OAI21_X1   g16568(.A1(new_n16630_), .A2(new_n16631_), .B(new_n16632_), .ZN(new_n16633_));
  OAI21_X1   g16569(.A1(new_n16633_), .A2(new_n16626_), .B(new_n16149_), .ZN(new_n16634_));
  OAI21_X1   g16570(.A1(new_n16634_), .A2(new_n16073_), .B(new_n16070_), .ZN(new_n16635_));
  NAND3_X1   g16571(.A1(new_n16635_), .A2(new_n16056_), .A3(new_n16060_), .ZN(new_n16636_));
  AOI22_X1   g16572(.A1(new_n16636_), .A2(new_n15990_), .B1(new_n16048_), .B2(new_n16042_), .ZN(new_n16637_));
  NOR2_X1    g16573(.A1(new_n15632_), .A2(new_n15863_), .ZN(new_n16638_));
  NOR2_X1    g16574(.A1(new_n15862_), .A2(new_n15637_), .ZN(new_n16639_));
  OAI22_X1   g16575(.A1(new_n11264_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n11277_), .ZN(new_n16640_));
  NAND2_X1   g16576(.A1(new_n11346_), .A2(new_n6838_), .ZN(new_n16641_));
  AOI21_X1   g16577(.A1(new_n16640_), .A2(new_n16641_), .B(new_n6836_), .ZN(new_n16642_));
  AND3_X2    g16578(.A1(new_n11757_), .A2(new_n65_), .A3(new_n16642_), .Z(new_n16643_));
  AOI21_X1   g16579(.A1(new_n11757_), .A2(new_n16642_), .B(new_n65_), .ZN(new_n16644_));
  NOR2_X1    g16580(.A1(new_n16643_), .A2(new_n16644_), .ZN(new_n16645_));
  INV_X1     g16581(.I(new_n16645_), .ZN(new_n16646_));
  NOR3_X1    g16582(.A1(new_n16638_), .A2(new_n16639_), .A3(new_n16646_), .ZN(new_n16647_));
  INV_X1     g16583(.I(new_n16647_), .ZN(new_n16648_));
  INV_X1     g16584(.I(new_n16638_), .ZN(new_n16649_));
  NAND2_X1   g16585(.A1(new_n15632_), .A2(new_n15863_), .ZN(new_n16650_));
  AOI21_X1   g16586(.A1(new_n16649_), .A2(new_n16650_), .B(new_n16645_), .ZN(new_n16651_));
  AOI21_X1   g16587(.A1(new_n16637_), .A2(new_n16648_), .B(new_n16651_), .ZN(new_n16652_));
  AOI21_X1   g16588(.A1(new_n15762_), .A2(new_n15869_), .B(new_n15864_), .ZN(new_n16653_));
  NOR3_X1    g16589(.A1(new_n15751_), .A2(new_n15756_), .A3(new_n15867_), .ZN(new_n16654_));
  INV_X1     g16590(.I(new_n16654_), .ZN(new_n16655_));
  OAI21_X1   g16591(.A1(new_n15751_), .A2(new_n15756_), .B(new_n15867_), .ZN(new_n16656_));
  AOI21_X1   g16592(.A1(new_n16655_), .A2(new_n16656_), .B(new_n15638_), .ZN(new_n16657_));
  OAI22_X1   g16593(.A1(new_n11264_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n11345_), .ZN(new_n16658_));
  NAND2_X1   g16594(.A1(new_n11354_), .A2(new_n6838_), .ZN(new_n16659_));
  AOI21_X1   g16595(.A1(new_n16659_), .A2(new_n16658_), .B(new_n6836_), .ZN(new_n16660_));
  OAI21_X1   g16596(.A1(new_n11675_), .A2(new_n11677_), .B(new_n16660_), .ZN(new_n16661_));
  XOR2_X1    g16597(.A1(new_n16661_), .A2(new_n65_), .Z(new_n16662_));
  NOR3_X1    g16598(.A1(new_n16657_), .A2(new_n16662_), .A3(new_n16653_), .ZN(new_n16663_));
  OAI21_X1   g16599(.A1(new_n16657_), .A2(new_n16653_), .B(new_n16662_), .ZN(new_n16664_));
  OAI21_X1   g16600(.A1(new_n16652_), .A2(new_n16663_), .B(new_n16664_), .ZN(new_n16665_));
  NAND3_X1   g16601(.A1(new_n15883_), .A2(new_n15880_), .A3(new_n13978_), .ZN(new_n16666_));
  INV_X1     g16602(.I(new_n13978_), .ZN(new_n16667_));
  OAI21_X1   g16603(.A1(new_n15861_), .A2(new_n15873_), .B(new_n16667_), .ZN(new_n16668_));
  NAND2_X1   g16604(.A1(new_n16668_), .A2(new_n16666_), .ZN(new_n16669_));
  NAND2_X1   g16605(.A1(new_n16669_), .A2(new_n13972_), .ZN(new_n16670_));
  NOR3_X1    g16606(.A1(new_n15861_), .A2(new_n15873_), .A3(new_n16667_), .ZN(new_n16671_));
  AOI21_X1   g16607(.A1(new_n15883_), .A2(new_n15880_), .B(new_n13978_), .ZN(new_n16672_));
  NOR2_X1    g16608(.A1(new_n16672_), .A2(new_n16671_), .ZN(new_n16673_));
  NAND2_X1   g16609(.A1(new_n16673_), .A2(new_n13973_), .ZN(new_n16674_));
  AOI21_X1   g16610(.A1(new_n16674_), .A2(new_n16670_), .B(new_n16665_), .ZN(new_n16675_));
  NOR3_X1    g16611(.A1(new_n16046_), .A2(new_n16047_), .A3(new_n16045_), .ZN(new_n16676_));
  AOI21_X1   g16612(.A1(new_n16032_), .A2(new_n16041_), .B(new_n15990_), .ZN(new_n16677_));
  INV_X1     g16613(.I(new_n16056_), .ZN(new_n16678_));
  NAND2_X1   g16614(.A1(new_n16060_), .A2(new_n16056_), .ZN(new_n16679_));
  NOR2_X1    g16615(.A1(new_n16069_), .A2(new_n16073_), .ZN(new_n16680_));
  OAI21_X1   g16616(.A1(new_n16151_), .A2(new_n16152_), .B(new_n16163_), .ZN(new_n16681_));
  NAND2_X1   g16617(.A1(new_n16632_), .A2(new_n16681_), .ZN(new_n16682_));
  INV_X1     g16618(.I(new_n16180_), .ZN(new_n16683_));
  INV_X1     g16619(.I(new_n16241_), .ZN(new_n16684_));
  NOR2_X1    g16620(.A1(new_n16257_), .A2(new_n16253_), .ZN(new_n16685_));
  NAND2_X1   g16621(.A1(new_n16536_), .A2(new_n16539_), .ZN(new_n16686_));
  AOI21_X1   g16622(.A1(new_n16597_), .A2(new_n16596_), .B(new_n16594_), .ZN(new_n16687_));
  NOR3_X1    g16623(.A1(new_n16589_), .A2(new_n16581_), .A3(new_n16590_), .ZN(new_n16688_));
  OAI21_X1   g16624(.A1(new_n16687_), .A2(new_n16688_), .B(new_n16604_), .ZN(new_n16689_));
  NAND2_X1   g16625(.A1(new_n16689_), .A2(new_n16686_), .ZN(new_n16690_));
  OR3_X2     g16626(.A1(new_n16687_), .A2(new_n16688_), .A3(new_n16604_), .Z(new_n16691_));
  AOI21_X1   g16627(.A1(new_n16608_), .A2(new_n16265_), .B(new_n16607_), .ZN(new_n16692_));
  NOR2_X1    g16628(.A1(new_n16692_), .A2(new_n16267_), .ZN(new_n16693_));
  NAND3_X1   g16629(.A1(new_n16690_), .A2(new_n16691_), .A3(new_n16693_), .ZN(new_n16694_));
  NAND3_X1   g16630(.A1(new_n16694_), .A2(new_n16685_), .A3(new_n16609_), .ZN(new_n16695_));
  NAND3_X1   g16631(.A1(new_n16618_), .A2(new_n16619_), .A3(new_n16617_), .ZN(new_n16696_));
  OAI21_X1   g16632(.A1(new_n16240_), .A2(new_n16234_), .B(new_n16190_), .ZN(new_n16697_));
  AOI21_X1   g16633(.A1(new_n16697_), .A2(new_n16696_), .B(new_n16621_), .ZN(new_n16698_));
  AOI21_X1   g16634(.A1(new_n16698_), .A2(new_n16695_), .B(new_n16684_), .ZN(new_n16699_));
  AOI21_X1   g16635(.A1(new_n16699_), .A2(new_n16182_), .B(new_n16683_), .ZN(new_n16700_));
  NOR2_X1    g16636(.A1(new_n16700_), .A2(new_n16682_), .ZN(new_n16701_));
  NAND3_X1   g16637(.A1(new_n16136_), .A2(new_n16147_), .A3(new_n16078_), .ZN(new_n16702_));
  OAI21_X1   g16638(.A1(new_n16628_), .A2(new_n16629_), .B(new_n16627_), .ZN(new_n16703_));
  AOI21_X1   g16639(.A1(new_n16703_), .A2(new_n16702_), .B(new_n16164_), .ZN(new_n16704_));
  AOI21_X1   g16640(.A1(new_n16704_), .A2(new_n16701_), .B(new_n16148_), .ZN(new_n16705_));
  AOI21_X1   g16641(.A1(new_n16705_), .A2(new_n16680_), .B(new_n16069_), .ZN(new_n16706_));
  NOR3_X1    g16642(.A1(new_n16706_), .A2(new_n16678_), .A3(new_n16679_), .ZN(new_n16707_));
  OAI22_X1   g16643(.A1(new_n16707_), .A2(new_n16045_), .B1(new_n16676_), .B2(new_n16677_), .ZN(new_n16708_));
  OAI21_X1   g16644(.A1(new_n16638_), .A2(new_n16639_), .B(new_n16646_), .ZN(new_n16709_));
  OAI21_X1   g16645(.A1(new_n16708_), .A2(new_n16647_), .B(new_n16709_), .ZN(new_n16710_));
  OAI21_X1   g16646(.A1(new_n15868_), .A2(new_n15763_), .B(new_n15638_), .ZN(new_n16711_));
  AOI21_X1   g16647(.A1(new_n15866_), .A2(new_n15865_), .B(new_n15761_), .ZN(new_n16712_));
  OAI21_X1   g16648(.A1(new_n16654_), .A2(new_n16712_), .B(new_n15864_), .ZN(new_n16713_));
  AOI21_X1   g16649(.A1(new_n16711_), .A2(new_n16713_), .B(new_n16662_), .ZN(new_n16714_));
  XOR2_X1    g16650(.A1(new_n16661_), .A2(\a[5] ), .Z(new_n16715_));
  NOR3_X1    g16651(.A1(new_n16657_), .A2(new_n16653_), .A3(new_n16715_), .ZN(new_n16716_));
  OAI21_X1   g16652(.A1(new_n16714_), .A2(new_n16716_), .B(new_n16710_), .ZN(new_n16717_));
  NAND3_X1   g16653(.A1(new_n16711_), .A2(new_n16713_), .A3(new_n16715_), .ZN(new_n16718_));
  NAND2_X1   g16654(.A1(new_n16664_), .A2(new_n16718_), .ZN(new_n16719_));
  NAND2_X1   g16655(.A1(new_n16719_), .A2(new_n16652_), .ZN(new_n16720_));
  OAI22_X1   g16656(.A1(new_n11369_), .A2(new_n9485_), .B1(new_n9489_), .B2(new_n11461_), .ZN(new_n16721_));
  NAND2_X1   g16657(.A1(new_n11694_), .A2(new_n9503_), .ZN(new_n16722_));
  AOI21_X1   g16658(.A1(new_n16721_), .A2(new_n16722_), .B(new_n9482_), .ZN(new_n16723_));
  NAND2_X1   g16659(.A1(new_n12720_), .A2(new_n16723_), .ZN(new_n16724_));
  XOR2_X1    g16660(.A1(new_n16724_), .A2(new_n4387_), .Z(new_n16725_));
  NAND3_X1   g16661(.A1(new_n16725_), .A2(new_n16717_), .A3(new_n16720_), .ZN(new_n16726_));
  NAND2_X1   g16662(.A1(new_n16710_), .A2(new_n16718_), .ZN(new_n16727_));
  AOI21_X1   g16663(.A1(new_n16727_), .A2(new_n16664_), .B(new_n13973_), .ZN(new_n16728_));
  NOR2_X1    g16664(.A1(new_n16665_), .A2(new_n13972_), .ZN(new_n16729_));
  OAI21_X1   g16665(.A1(new_n16729_), .A2(new_n16728_), .B(new_n16669_), .ZN(new_n16730_));
  NOR2_X1    g16666(.A1(new_n16665_), .A2(new_n13973_), .ZN(new_n16731_));
  AOI21_X1   g16667(.A1(new_n16727_), .A2(new_n16664_), .B(new_n13972_), .ZN(new_n16732_));
  OAI21_X1   g16668(.A1(new_n16731_), .A2(new_n16732_), .B(new_n16673_), .ZN(new_n16733_));
  NAND2_X1   g16669(.A1(new_n16730_), .A2(new_n16733_), .ZN(new_n16734_));
  AOI21_X1   g16670(.A1(new_n16734_), .A2(new_n16726_), .B(new_n16675_), .ZN(new_n16735_));
  OAI21_X1   g16671(.A1(new_n16735_), .A2(new_n15876_), .B(new_n15980_), .ZN(new_n16736_));
  OAI22_X1   g16672(.A1(new_n11264_), .A2(new_n6783_), .B1(new_n6788_), .B2(new_n11345_), .ZN(new_n16737_));
  NAND2_X1   g16673(.A1(new_n11354_), .A2(new_n6784_), .ZN(new_n16738_));
  AOI21_X1   g16674(.A1(new_n16738_), .A2(new_n16737_), .B(new_n6776_), .ZN(new_n16739_));
  NAND2_X1   g16675(.A1(new_n11678_), .A2(new_n16739_), .ZN(new_n16740_));
  XOR2_X1    g16676(.A1(new_n16740_), .A2(new_n4009_), .Z(new_n16741_));
  OAI22_X1   g16677(.A1(new_n11284_), .A2(new_n4716_), .B1(new_n4719_), .B2(new_n11271_), .ZN(new_n16742_));
  NAND2_X1   g16678(.A1(new_n11311_), .A2(new_n4709_), .ZN(new_n16743_));
  AOI21_X1   g16679(.A1(new_n16742_), .A2(new_n16743_), .B(new_n4707_), .ZN(new_n16744_));
  NAND2_X1   g16680(.A1(new_n11391_), .A2(new_n16744_), .ZN(new_n16745_));
  XOR2_X1    g16681(.A1(new_n16745_), .A2(\a[11] ), .Z(new_n16746_));
  OAI22_X1   g16682(.A1(new_n8701_), .A2(new_n4291_), .B1(new_n8694_), .B2(new_n4297_), .ZN(new_n16747_));
  NAND2_X1   g16683(.A1(new_n8682_), .A2(new_n4469_), .ZN(new_n16748_));
  AOI21_X1   g16684(.A1(new_n16748_), .A2(new_n16747_), .B(new_n4468_), .ZN(new_n16749_));
  NAND2_X1   g16685(.A1(new_n12347_), .A2(new_n16749_), .ZN(new_n16750_));
  XOR2_X1    g16686(.A1(new_n16750_), .A2(\a[17] ), .Z(new_n16751_));
  NOR2_X1    g16687(.A1(new_n15920_), .A2(new_n15911_), .ZN(new_n16752_));
  NOR2_X1    g16688(.A1(new_n16752_), .A2(new_n15907_), .ZN(new_n16753_));
  NAND3_X1   g16689(.A1(new_n13809_), .A2(new_n13811_), .A3(new_n13865_), .ZN(new_n16754_));
  OAI21_X1   g16690(.A1(new_n13885_), .A2(new_n13883_), .B(new_n13866_), .ZN(new_n16755_));
  NAND3_X1   g16691(.A1(new_n16755_), .A2(new_n16754_), .A3(new_n16753_), .ZN(new_n16756_));
  INV_X1     g16692(.I(new_n16753_), .ZN(new_n16757_));
  NOR3_X1    g16693(.A1(new_n13885_), .A2(new_n13883_), .A3(new_n13866_), .ZN(new_n16758_));
  AOI21_X1   g16694(.A1(new_n13809_), .A2(new_n13811_), .B(new_n13865_), .ZN(new_n16759_));
  OAI21_X1   g16695(.A1(new_n16758_), .A2(new_n16759_), .B(new_n16757_), .ZN(new_n16760_));
  AOI21_X1   g16696(.A1(new_n16760_), .A2(new_n16756_), .B(new_n13886_), .ZN(new_n16761_));
  NOR3_X1    g16697(.A1(new_n16758_), .A2(new_n16759_), .A3(new_n16757_), .ZN(new_n16762_));
  AOI21_X1   g16698(.A1(new_n16755_), .A2(new_n16754_), .B(new_n16753_), .ZN(new_n16763_));
  NOR3_X1    g16699(.A1(new_n16762_), .A2(new_n16763_), .A3(new_n13871_), .ZN(new_n16764_));
  OAI21_X1   g16700(.A1(new_n16764_), .A2(new_n16761_), .B(new_n16751_), .ZN(new_n16765_));
  INV_X1     g16701(.I(new_n16751_), .ZN(new_n16766_));
  OAI21_X1   g16702(.A1(new_n16762_), .A2(new_n16763_), .B(new_n13871_), .ZN(new_n16767_));
  NAND3_X1   g16703(.A1(new_n16760_), .A2(new_n16756_), .A3(new_n13886_), .ZN(new_n16768_));
  NAND3_X1   g16704(.A1(new_n16767_), .A2(new_n16768_), .A3(new_n16766_), .ZN(new_n16769_));
  NOR2_X1    g16705(.A1(new_n15921_), .A2(new_n15901_), .ZN(new_n16770_));
  NAND2_X1   g16706(.A1(new_n16752_), .A2(new_n15919_), .ZN(new_n16771_));
  OAI21_X1   g16707(.A1(new_n15920_), .A2(new_n15911_), .B(new_n15907_), .ZN(new_n16772_));
  AOI22_X1   g16708(.A1(new_n16771_), .A2(new_n16772_), .B1(new_n15901_), .B2(new_n15921_), .ZN(new_n16773_));
  OAI22_X1   g16709(.A1(new_n8673_), .A2(new_n6094_), .B1(new_n8687_), .B2(new_n6089_), .ZN(new_n16774_));
  NAND2_X1   g16710(.A1(new_n8662_), .A2(new_n6090_), .ZN(new_n16775_));
  AOI21_X1   g16711(.A1(new_n16775_), .A2(new_n16774_), .B(new_n6082_), .ZN(new_n16776_));
  NAND2_X1   g16712(.A1(new_n11624_), .A2(new_n16776_), .ZN(new_n16777_));
  XOR2_X1    g16713(.A1(new_n16777_), .A2(\a[14] ), .Z(new_n16778_));
  INV_X1     g16714(.I(new_n16778_), .ZN(new_n16779_));
  NOR3_X1    g16715(.A1(new_n16773_), .A2(new_n16770_), .A3(new_n16779_), .ZN(new_n16780_));
  OAI21_X1   g16716(.A1(new_n16773_), .A2(new_n16770_), .B(new_n16779_), .ZN(new_n16781_));
  INV_X1     g16717(.I(new_n16781_), .ZN(new_n16782_));
  NOR2_X1    g16718(.A1(new_n16782_), .A2(new_n16780_), .ZN(new_n16783_));
  AOI21_X1   g16719(.A1(new_n16765_), .A2(new_n16769_), .B(new_n16783_), .ZN(new_n16784_));
  AOI21_X1   g16720(.A1(new_n16767_), .A2(new_n16768_), .B(new_n16766_), .ZN(new_n16785_));
  NOR3_X1    g16721(.A1(new_n16764_), .A2(new_n16761_), .A3(new_n16751_), .ZN(new_n16786_));
  OAI21_X1   g16722(.A1(new_n16773_), .A2(new_n16770_), .B(new_n16778_), .ZN(new_n16787_));
  INV_X1     g16723(.I(new_n16787_), .ZN(new_n16788_));
  NOR3_X1    g16724(.A1(new_n16773_), .A2(new_n16770_), .A3(new_n16778_), .ZN(new_n16789_));
  NOR2_X1    g16725(.A1(new_n16788_), .A2(new_n16789_), .ZN(new_n16790_));
  NOR3_X1    g16726(.A1(new_n16786_), .A2(new_n16785_), .A3(new_n16790_), .ZN(new_n16791_));
  AOI21_X1   g16727(.A1(new_n15934_), .A2(new_n15935_), .B(new_n15932_), .ZN(new_n16792_));
  INV_X1     g16728(.I(new_n16792_), .ZN(new_n16793_));
  NOR3_X1    g16729(.A1(new_n16791_), .A2(new_n16784_), .A3(new_n16793_), .ZN(new_n16794_));
  INV_X1     g16730(.I(new_n16780_), .ZN(new_n16795_));
  NAND2_X1   g16731(.A1(new_n16795_), .A2(new_n16781_), .ZN(new_n16796_));
  OAI21_X1   g16732(.A1(new_n16786_), .A2(new_n16785_), .B(new_n16796_), .ZN(new_n16797_));
  INV_X1     g16733(.I(new_n16789_), .ZN(new_n16798_));
  NAND2_X1   g16734(.A1(new_n16798_), .A2(new_n16787_), .ZN(new_n16799_));
  NAND3_X1   g16735(.A1(new_n16765_), .A2(new_n16769_), .A3(new_n16799_), .ZN(new_n16800_));
  AOI21_X1   g16736(.A1(new_n16797_), .A2(new_n16800_), .B(new_n16792_), .ZN(new_n16801_));
  NAND2_X1   g16737(.A1(new_n15933_), .A2(new_n15937_), .ZN(new_n16802_));
  NAND2_X1   g16738(.A1(new_n15938_), .A2(new_n15895_), .ZN(new_n16803_));
  NOR2_X1    g16739(.A1(new_n15938_), .A2(new_n15895_), .ZN(new_n16804_));
  AOI21_X1   g16740(.A1(new_n16802_), .A2(new_n16803_), .B(new_n16804_), .ZN(new_n16805_));
  NOR3_X1    g16741(.A1(new_n16794_), .A2(new_n16801_), .A3(new_n16805_), .ZN(new_n16806_));
  NAND3_X1   g16742(.A1(new_n16797_), .A2(new_n16800_), .A3(new_n16792_), .ZN(new_n16807_));
  OAI21_X1   g16743(.A1(new_n16791_), .A2(new_n16784_), .B(new_n16793_), .ZN(new_n16808_));
  INV_X1     g16744(.I(new_n16805_), .ZN(new_n16809_));
  AOI21_X1   g16745(.A1(new_n16808_), .A2(new_n16807_), .B(new_n16809_), .ZN(new_n16810_));
  OAI21_X1   g16746(.A1(new_n16806_), .A2(new_n16810_), .B(new_n16746_), .ZN(new_n16811_));
  INV_X1     g16747(.I(new_n16746_), .ZN(new_n16812_));
  NAND3_X1   g16748(.A1(new_n16808_), .A2(new_n16807_), .A3(new_n16809_), .ZN(new_n16813_));
  OAI21_X1   g16749(.A1(new_n16794_), .A2(new_n16801_), .B(new_n16805_), .ZN(new_n16814_));
  NAND3_X1   g16750(.A1(new_n16814_), .A2(new_n16813_), .A3(new_n16812_), .ZN(new_n16815_));
  AOI21_X1   g16751(.A1(new_n16811_), .A2(new_n16815_), .B(new_n16741_), .ZN(new_n16816_));
  XOR2_X1    g16752(.A1(new_n16740_), .A2(\a[8] ), .Z(new_n16817_));
  AOI21_X1   g16753(.A1(new_n16814_), .A2(new_n16813_), .B(new_n16812_), .ZN(new_n16818_));
  NOR3_X1    g16754(.A1(new_n16806_), .A2(new_n16810_), .A3(new_n16746_), .ZN(new_n16819_));
  NOR3_X1    g16755(.A1(new_n16819_), .A2(new_n16818_), .A3(new_n16817_), .ZN(new_n16820_));
  OAI21_X1   g16756(.A1(new_n15947_), .A2(new_n15944_), .B(new_n15949_), .ZN(new_n16821_));
  NOR3_X1    g16757(.A1(new_n12714_), .A2(new_n11466_), .A3(new_n12716_), .ZN(new_n16822_));
  INV_X1     g16758(.I(new_n12719_), .ZN(new_n16823_));
  OAI22_X1   g16759(.A1(new_n11369_), .A2(new_n6913_), .B1(new_n6839_), .B2(new_n11461_), .ZN(new_n16824_));
  NAND2_X1   g16760(.A1(new_n11694_), .A2(new_n8799_), .ZN(new_n16825_));
  AOI21_X1   g16761(.A1(new_n16824_), .A2(new_n16825_), .B(new_n6836_), .ZN(new_n16826_));
  OAI21_X1   g16762(.A1(new_n16823_), .A2(new_n16822_), .B(new_n16826_), .ZN(new_n16827_));
  NOR2_X1    g16763(.A1(new_n16827_), .A2(\a[5] ), .ZN(new_n16828_));
  AOI21_X1   g16764(.A1(new_n12720_), .A2(new_n16826_), .B(new_n65_), .ZN(new_n16829_));
  NOR2_X1    g16765(.A1(new_n16828_), .A2(new_n16829_), .ZN(new_n16830_));
  NAND2_X1   g16766(.A1(new_n16830_), .A2(new_n16821_), .ZN(new_n16831_));
  INV_X1     g16767(.I(new_n16831_), .ZN(new_n16832_));
  NOR2_X1    g16768(.A1(new_n16830_), .A2(new_n16821_), .ZN(new_n16833_));
  OAI22_X1   g16769(.A1(new_n16820_), .A2(new_n16816_), .B1(new_n16832_), .B2(new_n16833_), .ZN(new_n16834_));
  OAI21_X1   g16770(.A1(new_n16819_), .A2(new_n16818_), .B(new_n16817_), .ZN(new_n16835_));
  NAND3_X1   g16771(.A1(new_n16811_), .A2(new_n16815_), .A3(new_n16741_), .ZN(new_n16836_));
  XOR2_X1    g16772(.A1(new_n16830_), .A2(new_n16821_), .Z(new_n16837_));
  NAND3_X1   g16773(.A1(new_n16837_), .A2(new_n16835_), .A3(new_n16836_), .ZN(new_n16838_));
  AOI21_X1   g16774(.A1(new_n15972_), .A2(new_n15953_), .B(new_n15963_), .ZN(new_n16839_));
  NAND3_X1   g16775(.A1(new_n16834_), .A2(new_n16838_), .A3(new_n16839_), .ZN(new_n16840_));
  INV_X1     g16776(.I(new_n16840_), .ZN(new_n16841_));
  INV_X1     g16777(.I(new_n16833_), .ZN(new_n16842_));
  AOI22_X1   g16778(.A1(new_n16835_), .A2(new_n16836_), .B1(new_n16831_), .B2(new_n16842_), .ZN(new_n16843_));
  INV_X1     g16779(.I(new_n16838_), .ZN(new_n16844_));
  INV_X1     g16780(.I(new_n16839_), .ZN(new_n16845_));
  OAI21_X1   g16781(.A1(new_n16844_), .A2(new_n16843_), .B(new_n16845_), .ZN(new_n16846_));
  OAI21_X1   g16782(.A1(new_n16736_), .A2(new_n16841_), .B(new_n16846_), .ZN(new_n16847_));
  AOI22_X1   g16783(.A1(new_n11311_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n11272_), .ZN(new_n16848_));
  NOR2_X1    g16784(.A1(new_n11264_), .A2(new_n4710_), .ZN(new_n16849_));
  OAI21_X1   g16785(.A1(new_n16849_), .A2(new_n16848_), .B(new_n4706_), .ZN(new_n16850_));
  NOR2_X1    g16786(.A1(new_n11310_), .A2(new_n16850_), .ZN(new_n16851_));
  XOR2_X1    g16787(.A1(new_n16851_), .A2(new_n4034_), .Z(new_n16852_));
  OAI22_X1   g16788(.A1(new_n8661_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8673_), .ZN(new_n16853_));
  NAND2_X1   g16789(.A1(new_n11285_), .A2(new_n6090_), .ZN(new_n16854_));
  AOI21_X1   g16790(.A1(new_n16854_), .A2(new_n16853_), .B(new_n6082_), .ZN(new_n16855_));
  NAND2_X1   g16791(.A1(new_n11323_), .A2(new_n16855_), .ZN(new_n16856_));
  XOR2_X1    g16792(.A1(new_n16856_), .A2(\a[14] ), .Z(new_n16857_));
  INV_X1     g16793(.I(new_n16857_), .ZN(new_n16858_));
  OAI21_X1   g16794(.A1(new_n16786_), .A2(new_n16785_), .B(new_n16795_), .ZN(new_n16859_));
  NAND2_X1   g16795(.A1(new_n16859_), .A2(new_n16781_), .ZN(new_n16860_));
  NOR2_X1    g16796(.A1(new_n13889_), .A2(new_n13880_), .ZN(new_n16861_));
  INV_X1     g16797(.I(new_n16861_), .ZN(new_n16862_));
  OAI21_X1   g16798(.A1(new_n13806_), .A2(new_n13803_), .B(new_n16862_), .ZN(new_n16863_));
  AOI21_X1   g16799(.A1(new_n13887_), .A2(new_n13888_), .B(new_n13879_), .ZN(new_n16864_));
  NOR3_X1    g16800(.A1(new_n13872_), .A2(new_n13873_), .A3(new_n13878_), .ZN(new_n16865_));
  OR2_X2     g16801(.A1(new_n16864_), .A2(new_n16865_), .Z(new_n16866_));
  NAND3_X1   g16802(.A1(new_n13913_), .A2(new_n13914_), .A3(new_n16866_), .ZN(new_n16867_));
  NOR2_X1    g16803(.A1(new_n16757_), .A2(new_n16751_), .ZN(new_n16868_));
  NAND2_X1   g16804(.A1(new_n16757_), .A2(new_n16751_), .ZN(new_n16869_));
  NAND3_X1   g16805(.A1(new_n16755_), .A2(new_n16754_), .A3(new_n13886_), .ZN(new_n16870_));
  OAI21_X1   g16806(.A1(new_n16758_), .A2(new_n16759_), .B(new_n13871_), .ZN(new_n16871_));
  NAND2_X1   g16807(.A1(new_n16871_), .A2(new_n16870_), .ZN(new_n16872_));
  AOI21_X1   g16808(.A1(new_n16872_), .A2(new_n16869_), .B(new_n16868_), .ZN(new_n16873_));
  INV_X1     g16809(.I(new_n16873_), .ZN(new_n16874_));
  NAND3_X1   g16810(.A1(new_n16863_), .A2(new_n16867_), .A3(new_n16874_), .ZN(new_n16875_));
  AOI21_X1   g16811(.A1(new_n13913_), .A2(new_n13914_), .B(new_n16861_), .ZN(new_n16876_));
  NOR2_X1    g16812(.A1(new_n16864_), .A2(new_n16865_), .ZN(new_n16877_));
  NOR3_X1    g16813(.A1(new_n13806_), .A2(new_n13803_), .A3(new_n16877_), .ZN(new_n16878_));
  OAI21_X1   g16814(.A1(new_n16878_), .A2(new_n16876_), .B(new_n16873_), .ZN(new_n16879_));
  NAND3_X1   g16815(.A1(new_n16860_), .A2(new_n16879_), .A3(new_n16875_), .ZN(new_n16880_));
  NAND2_X1   g16816(.A1(new_n16765_), .A2(new_n16769_), .ZN(new_n16881_));
  AOI21_X1   g16817(.A1(new_n16881_), .A2(new_n16795_), .B(new_n16782_), .ZN(new_n16882_));
  NOR3_X1    g16818(.A1(new_n16878_), .A2(new_n16876_), .A3(new_n16873_), .ZN(new_n16883_));
  AOI21_X1   g16819(.A1(new_n16863_), .A2(new_n16867_), .B(new_n16874_), .ZN(new_n16884_));
  OAI21_X1   g16820(.A1(new_n16883_), .A2(new_n16884_), .B(new_n16882_), .ZN(new_n16885_));
  AOI21_X1   g16821(.A1(new_n16885_), .A2(new_n16880_), .B(new_n16858_), .ZN(new_n16886_));
  NOR3_X1    g16822(.A1(new_n16882_), .A2(new_n16883_), .A3(new_n16884_), .ZN(new_n16887_));
  AOI21_X1   g16823(.A1(new_n16875_), .A2(new_n16879_), .B(new_n16860_), .ZN(new_n16888_));
  NOR3_X1    g16824(.A1(new_n16888_), .A2(new_n16887_), .A3(new_n16857_), .ZN(new_n16889_));
  OAI21_X1   g16825(.A1(new_n16889_), .A2(new_n16886_), .B(new_n16852_), .ZN(new_n16890_));
  INV_X1     g16826(.I(new_n16852_), .ZN(new_n16891_));
  OAI21_X1   g16827(.A1(new_n16888_), .A2(new_n16887_), .B(new_n16857_), .ZN(new_n16892_));
  NAND3_X1   g16828(.A1(new_n16885_), .A2(new_n16880_), .A3(new_n16858_), .ZN(new_n16893_));
  NAND3_X1   g16829(.A1(new_n16892_), .A2(new_n16893_), .A3(new_n16891_), .ZN(new_n16894_));
  OAI22_X1   g16830(.A1(new_n16791_), .A2(new_n16784_), .B1(new_n16812_), .B2(new_n16792_), .ZN(new_n16895_));
  NOR2_X1    g16831(.A1(new_n16793_), .A2(new_n16746_), .ZN(new_n16896_));
  INV_X1     g16832(.I(new_n16896_), .ZN(new_n16897_));
  OAI22_X1   g16833(.A1(new_n11353_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n11345_), .ZN(new_n16898_));
  NAND2_X1   g16834(.A1(new_n11370_), .A2(new_n6784_), .ZN(new_n16899_));
  AOI21_X1   g16835(.A1(new_n16899_), .A2(new_n16898_), .B(new_n6776_), .ZN(new_n16900_));
  NAND2_X1   g16836(.A1(new_n11379_), .A2(new_n16900_), .ZN(new_n16901_));
  XOR2_X1    g16837(.A1(new_n16901_), .A2(\a[8] ), .Z(new_n16902_));
  NAND3_X1   g16838(.A1(new_n16895_), .A2(new_n16897_), .A3(new_n16902_), .ZN(new_n16903_));
  AOI22_X1   g16839(.A1(new_n16797_), .A2(new_n16800_), .B1(new_n16746_), .B2(new_n16793_), .ZN(new_n16904_));
  INV_X1     g16840(.I(new_n16902_), .ZN(new_n16905_));
  OAI21_X1   g16841(.A1(new_n16904_), .A2(new_n16896_), .B(new_n16905_), .ZN(new_n16906_));
  NAND2_X1   g16842(.A1(new_n16903_), .A2(new_n16906_), .ZN(new_n16907_));
  INV_X1     g16843(.I(new_n16907_), .ZN(new_n16908_));
  AOI21_X1   g16844(.A1(new_n16890_), .A2(new_n16894_), .B(new_n16908_), .ZN(new_n16909_));
  AOI21_X1   g16845(.A1(new_n16892_), .A2(new_n16893_), .B(new_n16891_), .ZN(new_n16910_));
  NOR3_X1    g16846(.A1(new_n16889_), .A2(new_n16886_), .A3(new_n16852_), .ZN(new_n16911_));
  NOR2_X1    g16847(.A1(new_n16904_), .A2(new_n16896_), .ZN(new_n16912_));
  XOR2_X1    g16848(.A1(new_n16912_), .A2(new_n16905_), .Z(new_n16913_));
  NOR3_X1    g16849(.A1(new_n16911_), .A2(new_n16913_), .A3(new_n16910_), .ZN(new_n16914_));
  NOR2_X1    g16850(.A1(new_n16914_), .A2(new_n16909_), .ZN(new_n16915_));
  NOR2_X1    g16851(.A1(new_n16817_), .A2(new_n16805_), .ZN(new_n16916_));
  NOR2_X1    g16852(.A1(new_n16741_), .A2(new_n16809_), .ZN(new_n16917_));
  NAND3_X1   g16853(.A1(new_n16808_), .A2(new_n16807_), .A3(new_n16812_), .ZN(new_n16918_));
  OAI21_X1   g16854(.A1(new_n16794_), .A2(new_n16801_), .B(new_n16746_), .ZN(new_n16919_));
  AOI21_X1   g16855(.A1(new_n16919_), .A2(new_n16918_), .B(new_n16917_), .ZN(new_n16920_));
  NOR3_X1    g16856(.A1(new_n11466_), .A2(new_n6913_), .A3(new_n11868_), .ZN(new_n16921_));
  NOR4_X1    g16857(.A1(new_n11468_), .A2(new_n6836_), .A3(new_n11461_), .A4(new_n16921_), .ZN(new_n16922_));
  XOR2_X1    g16858(.A1(new_n16922_), .A2(new_n65_), .Z(new_n16923_));
  NOR3_X1    g16859(.A1(new_n16920_), .A2(new_n16916_), .A3(new_n16923_), .ZN(new_n16924_));
  INV_X1     g16860(.I(new_n16916_), .ZN(new_n16925_));
  NAND2_X1   g16861(.A1(new_n16817_), .A2(new_n16805_), .ZN(new_n16926_));
  NOR3_X1    g16862(.A1(new_n16794_), .A2(new_n16801_), .A3(new_n16746_), .ZN(new_n16927_));
  AOI21_X1   g16863(.A1(new_n16808_), .A2(new_n16807_), .B(new_n16812_), .ZN(new_n16928_));
  OAI21_X1   g16864(.A1(new_n16927_), .A2(new_n16928_), .B(new_n16926_), .ZN(new_n16929_));
  INV_X1     g16865(.I(new_n16923_), .ZN(new_n16930_));
  AOI21_X1   g16866(.A1(new_n16929_), .A2(new_n16925_), .B(new_n16930_), .ZN(new_n16931_));
  NOR2_X1    g16867(.A1(new_n16931_), .A2(new_n16924_), .ZN(new_n16932_));
  OAI21_X1   g16868(.A1(new_n16820_), .A2(new_n16816_), .B(new_n16831_), .ZN(new_n16933_));
  NAND3_X1   g16869(.A1(new_n16933_), .A2(new_n16932_), .A3(new_n16842_), .ZN(new_n16934_));
  NAND3_X1   g16870(.A1(new_n16929_), .A2(new_n16930_), .A3(new_n16925_), .ZN(new_n16935_));
  OAI21_X1   g16871(.A1(new_n16920_), .A2(new_n16916_), .B(new_n16923_), .ZN(new_n16936_));
  NAND2_X1   g16872(.A1(new_n16935_), .A2(new_n16936_), .ZN(new_n16937_));
  AOI21_X1   g16873(.A1(new_n16835_), .A2(new_n16836_), .B(new_n16832_), .ZN(new_n16938_));
  OAI21_X1   g16874(.A1(new_n16938_), .A2(new_n16833_), .B(new_n16937_), .ZN(new_n16939_));
  AOI21_X1   g16875(.A1(new_n16934_), .A2(new_n16939_), .B(new_n16915_), .ZN(new_n16940_));
  NAND2_X1   g16876(.A1(new_n16890_), .A2(new_n16894_), .ZN(new_n16941_));
  OAI21_X1   g16877(.A1(new_n16911_), .A2(new_n16910_), .B(new_n16907_), .ZN(new_n16942_));
  OAI21_X1   g16878(.A1(new_n16941_), .A2(new_n16913_), .B(new_n16942_), .ZN(new_n16943_));
  NAND3_X1   g16879(.A1(new_n16933_), .A2(new_n16842_), .A3(new_n16937_), .ZN(new_n16944_));
  OAI21_X1   g16880(.A1(new_n16938_), .A2(new_n16833_), .B(new_n16932_), .ZN(new_n16945_));
  AOI21_X1   g16881(.A1(new_n16944_), .A2(new_n16945_), .B(new_n16943_), .ZN(new_n16946_));
  NOR2_X1    g16882(.A1(new_n16946_), .A2(new_n16940_), .ZN(new_n16947_));
  NOR2_X1    g16883(.A1(new_n16938_), .A2(new_n16833_), .ZN(new_n16948_));
  NOR3_X1    g16884(.A1(new_n16914_), .A2(new_n16909_), .A3(new_n16937_), .ZN(new_n16949_));
  OAI21_X1   g16885(.A1(new_n16914_), .A2(new_n16909_), .B(new_n16937_), .ZN(new_n16950_));
  INV_X1     g16886(.I(new_n16950_), .ZN(new_n16951_));
  OAI21_X1   g16887(.A1(new_n16951_), .A2(new_n16949_), .B(new_n16948_), .ZN(new_n16952_));
  OAI21_X1   g16888(.A1(new_n16947_), .A2(new_n16847_), .B(new_n16952_), .ZN(new_n16953_));
  NAND2_X1   g16889(.A1(new_n16941_), .A2(new_n16903_), .ZN(new_n16954_));
  NAND2_X1   g16890(.A1(new_n16954_), .A2(new_n16906_), .ZN(new_n16955_));
  AOI22_X1   g16891(.A1(new_n16863_), .A2(new_n16867_), .B1(new_n16857_), .B2(new_n16873_), .ZN(new_n16956_));
  NOR2_X1    g16892(.A1(new_n16873_), .A2(new_n16857_), .ZN(new_n16957_));
  NOR2_X1    g16893(.A1(new_n16956_), .A2(new_n16957_), .ZN(new_n16958_));
  INV_X1     g16894(.I(new_n16958_), .ZN(new_n16959_));
  OAI22_X1   g16895(.A1(new_n11264_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n11277_), .ZN(new_n16960_));
  NAND2_X1   g16896(.A1(new_n11346_), .A2(new_n4709_), .ZN(new_n16961_));
  AOI21_X1   g16897(.A1(new_n16960_), .A2(new_n16961_), .B(new_n4707_), .ZN(new_n16962_));
  NAND2_X1   g16898(.A1(new_n11757_), .A2(new_n16962_), .ZN(new_n16963_));
  XOR2_X1    g16899(.A1(new_n16963_), .A2(\a[11] ), .Z(new_n16964_));
  NOR2_X1    g16900(.A1(new_n16882_), .A2(new_n16852_), .ZN(new_n16965_));
  NAND2_X1   g16901(.A1(new_n16882_), .A2(new_n16852_), .ZN(new_n16966_));
  NAND3_X1   g16902(.A1(new_n16879_), .A2(new_n16875_), .A3(new_n16858_), .ZN(new_n16967_));
  OAI21_X1   g16903(.A1(new_n16883_), .A2(new_n16884_), .B(new_n16857_), .ZN(new_n16968_));
  NAND2_X1   g16904(.A1(new_n16968_), .A2(new_n16967_), .ZN(new_n16969_));
  AOI21_X1   g16905(.A1(new_n16969_), .A2(new_n16966_), .B(new_n16965_), .ZN(new_n16970_));
  OAI22_X1   g16906(.A1(new_n11284_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n8661_), .ZN(new_n16971_));
  NAND2_X1   g16907(.A1(new_n11272_), .A2(new_n6090_), .ZN(new_n16972_));
  AOI21_X1   g16908(.A1(new_n16971_), .A2(new_n16972_), .B(new_n6082_), .ZN(new_n16973_));
  NAND2_X1   g16909(.A1(new_n11655_), .A2(new_n16973_), .ZN(new_n16974_));
  XOR2_X1    g16910(.A1(new_n16974_), .A2(\a[14] ), .Z(new_n16975_));
  OAI21_X1   g16911(.A1(new_n13915_), .A2(new_n13889_), .B(new_n13916_), .ZN(new_n16976_));
  OAI21_X1   g16912(.A1(new_n13911_), .A2(new_n13910_), .B(new_n13327_), .ZN(new_n16977_));
  NAND3_X1   g16913(.A1(new_n13905_), .A2(new_n13908_), .A3(new_n13328_), .ZN(new_n16978_));
  NAND3_X1   g16914(.A1(new_n13882_), .A2(new_n13890_), .A3(new_n13895_), .ZN(new_n16979_));
  AOI22_X1   g16915(.A1(new_n16977_), .A2(new_n16978_), .B1(new_n16979_), .B2(new_n16976_), .ZN(new_n16980_));
  AOI21_X1   g16916(.A1(new_n13882_), .A2(new_n13890_), .B(new_n13916_), .ZN(new_n16981_));
  NOR3_X1    g16917(.A1(new_n13915_), .A2(new_n13889_), .A3(new_n13895_), .ZN(new_n16982_));
  NOR2_X1    g16918(.A1(new_n16981_), .A2(new_n16982_), .ZN(new_n16983_));
  NOR3_X1    g16919(.A1(new_n16983_), .A2(new_n13909_), .A3(new_n13912_), .ZN(new_n16984_));
  NOR3_X1    g16920(.A1(new_n16984_), .A2(new_n16975_), .A3(new_n16980_), .ZN(new_n16985_));
  INV_X1     g16921(.I(new_n16975_), .ZN(new_n16986_));
  OAI22_X1   g16922(.A1(new_n13909_), .A2(new_n13912_), .B1(new_n13896_), .B2(new_n13917_), .ZN(new_n16987_));
  OAI21_X1   g16923(.A1(new_n13915_), .A2(new_n13889_), .B(new_n13895_), .ZN(new_n16988_));
  NAND3_X1   g16924(.A1(new_n13882_), .A2(new_n13890_), .A3(new_n13916_), .ZN(new_n16989_));
  NAND2_X1   g16925(.A1(new_n16989_), .A2(new_n16988_), .ZN(new_n16990_));
  NAND3_X1   g16926(.A1(new_n16990_), .A2(new_n16977_), .A3(new_n16978_), .ZN(new_n16991_));
  AOI21_X1   g16927(.A1(new_n16991_), .A2(new_n16987_), .B(new_n16986_), .ZN(new_n16992_));
  NOR3_X1    g16928(.A1(new_n16970_), .A2(new_n16985_), .A3(new_n16992_), .ZN(new_n16993_));
  INV_X1     g16929(.I(new_n16965_), .ZN(new_n16994_));
  NOR3_X1    g16930(.A1(new_n16883_), .A2(new_n16884_), .A3(new_n16857_), .ZN(new_n16995_));
  AOI21_X1   g16931(.A1(new_n16879_), .A2(new_n16875_), .B(new_n16858_), .ZN(new_n16996_));
  OAI21_X1   g16932(.A1(new_n16995_), .A2(new_n16996_), .B(new_n16966_), .ZN(new_n16997_));
  NAND2_X1   g16933(.A1(new_n16997_), .A2(new_n16994_), .ZN(new_n16998_));
  NAND3_X1   g16934(.A1(new_n16991_), .A2(new_n16986_), .A3(new_n16987_), .ZN(new_n16999_));
  OAI21_X1   g16935(.A1(new_n16984_), .A2(new_n16980_), .B(new_n16975_), .ZN(new_n17000_));
  AOI21_X1   g16936(.A1(new_n16999_), .A2(new_n17000_), .B(new_n16998_), .ZN(new_n17001_));
  OAI21_X1   g16937(.A1(new_n17001_), .A2(new_n16993_), .B(new_n16964_), .ZN(new_n17002_));
  INV_X1     g16938(.I(new_n16964_), .ZN(new_n17003_));
  NAND3_X1   g16939(.A1(new_n16998_), .A2(new_n17000_), .A3(new_n16999_), .ZN(new_n17004_));
  OAI21_X1   g16940(.A1(new_n16985_), .A2(new_n16992_), .B(new_n16970_), .ZN(new_n17005_));
  NAND3_X1   g16941(.A1(new_n17005_), .A2(new_n17004_), .A3(new_n17003_), .ZN(new_n17006_));
  AOI21_X1   g16942(.A1(new_n17002_), .A2(new_n17006_), .B(new_n16959_), .ZN(new_n17007_));
  AOI21_X1   g16943(.A1(new_n17005_), .A2(new_n17004_), .B(new_n17003_), .ZN(new_n17008_));
  NOR3_X1    g16944(.A1(new_n17001_), .A2(new_n16993_), .A3(new_n16964_), .ZN(new_n17009_));
  NOR3_X1    g16945(.A1(new_n17009_), .A2(new_n17008_), .A3(new_n16958_), .ZN(new_n17010_));
  OAI22_X1   g16946(.A1(new_n11353_), .A2(new_n6783_), .B1(new_n6785_), .B2(new_n11697_), .ZN(new_n17011_));
  NAND2_X1   g16947(.A1(new_n11370_), .A2(new_n6789_), .ZN(new_n17012_));
  AOI21_X1   g16948(.A1(new_n17012_), .A2(new_n17011_), .B(new_n6776_), .ZN(new_n17013_));
  NAND2_X1   g16949(.A1(new_n11700_), .A2(new_n17013_), .ZN(new_n17014_));
  XOR2_X1    g16950(.A1(new_n17014_), .A2(\a[8] ), .Z(new_n17015_));
  INV_X1     g16951(.I(new_n17015_), .ZN(new_n17016_));
  NOR3_X1    g16952(.A1(new_n17010_), .A2(new_n17007_), .A3(new_n17016_), .ZN(new_n17017_));
  OAI21_X1   g16953(.A1(new_n17009_), .A2(new_n17008_), .B(new_n16958_), .ZN(new_n17018_));
  NAND3_X1   g16954(.A1(new_n17002_), .A2(new_n17006_), .A3(new_n16959_), .ZN(new_n17019_));
  AOI21_X1   g16955(.A1(new_n17018_), .A2(new_n17019_), .B(new_n17015_), .ZN(new_n17020_));
  OAI21_X1   g16956(.A1(new_n17017_), .A2(new_n17020_), .B(new_n16955_), .ZN(new_n17021_));
  INV_X1     g16957(.I(new_n16955_), .ZN(new_n17022_));
  AOI21_X1   g16958(.A1(new_n17018_), .A2(new_n17019_), .B(new_n17016_), .ZN(new_n17023_));
  NOR3_X1    g16959(.A1(new_n17010_), .A2(new_n17007_), .A3(new_n17015_), .ZN(new_n17024_));
  OAI21_X1   g16960(.A1(new_n17024_), .A2(new_n17023_), .B(new_n17022_), .ZN(new_n17025_));
  NAND3_X1   g16961(.A1(new_n16953_), .A2(new_n17021_), .A3(new_n17025_), .ZN(new_n17026_));
  NOR2_X1    g16962(.A1(new_n15975_), .A2(new_n15978_), .ZN(new_n17027_));
  INV_X1     g16963(.I(new_n17027_), .ZN(new_n17028_));
  NAND2_X1   g16964(.A1(new_n17028_), .A2(new_n15876_), .ZN(new_n17029_));
  INV_X1     g16965(.I(new_n16665_), .ZN(new_n17030_));
  NOR2_X1    g16966(.A1(new_n16673_), .A2(new_n13973_), .ZN(new_n17031_));
  NOR2_X1    g16967(.A1(new_n16669_), .A2(new_n13972_), .ZN(new_n17032_));
  OAI21_X1   g16968(.A1(new_n17031_), .A2(new_n17032_), .B(new_n17030_), .ZN(new_n17033_));
  NAND2_X1   g16969(.A1(new_n16665_), .A2(new_n13972_), .ZN(new_n17034_));
  NAND3_X1   g16970(.A1(new_n16727_), .A2(new_n13973_), .A3(new_n16664_), .ZN(new_n17035_));
  AOI21_X1   g16971(.A1(new_n17034_), .A2(new_n17035_), .B(new_n16673_), .ZN(new_n17036_));
  NAND3_X1   g16972(.A1(new_n16727_), .A2(new_n13972_), .A3(new_n16664_), .ZN(new_n17037_));
  NAND2_X1   g16973(.A1(new_n16665_), .A2(new_n13973_), .ZN(new_n17038_));
  AOI21_X1   g16974(.A1(new_n17038_), .A2(new_n17037_), .B(new_n16669_), .ZN(new_n17039_));
  OAI21_X1   g16975(.A1(new_n17036_), .A2(new_n17039_), .B(new_n16726_), .ZN(new_n17040_));
  NAND3_X1   g16976(.A1(new_n17040_), .A2(new_n15980_), .A3(new_n17033_), .ZN(new_n17041_));
  NAND2_X1   g16977(.A1(new_n17041_), .A2(new_n17029_), .ZN(new_n17042_));
  AOI21_X1   g16978(.A1(new_n16834_), .A2(new_n16838_), .B(new_n16839_), .ZN(new_n17043_));
  AOI21_X1   g16979(.A1(new_n17042_), .A2(new_n16840_), .B(new_n17043_), .ZN(new_n17044_));
  NOR3_X1    g16980(.A1(new_n16938_), .A2(new_n16937_), .A3(new_n16833_), .ZN(new_n17045_));
  AOI21_X1   g16981(.A1(new_n16933_), .A2(new_n16842_), .B(new_n16932_), .ZN(new_n17046_));
  OAI21_X1   g16982(.A1(new_n17045_), .A2(new_n17046_), .B(new_n16943_), .ZN(new_n17047_));
  NOR3_X1    g16983(.A1(new_n16938_), .A2(new_n16932_), .A3(new_n16833_), .ZN(new_n17048_));
  AOI21_X1   g16984(.A1(new_n16933_), .A2(new_n16842_), .B(new_n16937_), .ZN(new_n17049_));
  OAI21_X1   g16985(.A1(new_n17049_), .A2(new_n17048_), .B(new_n16915_), .ZN(new_n17050_));
  NAND2_X1   g16986(.A1(new_n17047_), .A2(new_n17050_), .ZN(new_n17051_));
  INV_X1     g16987(.I(new_n16948_), .ZN(new_n17052_));
  INV_X1     g16988(.I(new_n16949_), .ZN(new_n17053_));
  AOI21_X1   g16989(.A1(new_n17053_), .A2(new_n16950_), .B(new_n17052_), .ZN(new_n17054_));
  AOI21_X1   g16990(.A1(new_n17051_), .A2(new_n17044_), .B(new_n17054_), .ZN(new_n17055_));
  NAND3_X1   g16991(.A1(new_n17018_), .A2(new_n17019_), .A3(new_n17015_), .ZN(new_n17056_));
  OAI21_X1   g16992(.A1(new_n17010_), .A2(new_n17007_), .B(new_n17016_), .ZN(new_n17057_));
  AOI21_X1   g16993(.A1(new_n17057_), .A2(new_n17056_), .B(new_n17022_), .ZN(new_n17058_));
  OAI21_X1   g16994(.A1(new_n17010_), .A2(new_n17007_), .B(new_n17015_), .ZN(new_n17059_));
  NAND3_X1   g16995(.A1(new_n17018_), .A2(new_n17019_), .A3(new_n17016_), .ZN(new_n17060_));
  AOI21_X1   g16996(.A1(new_n17059_), .A2(new_n17060_), .B(new_n16955_), .ZN(new_n17061_));
  OAI21_X1   g16997(.A1(new_n17058_), .A2(new_n17061_), .B(new_n17055_), .ZN(new_n17062_));
  NAND3_X1   g16998(.A1(new_n16929_), .A2(new_n16925_), .A3(new_n16923_), .ZN(new_n17063_));
  AOI21_X1   g16999(.A1(new_n16929_), .A2(new_n16925_), .B(new_n16923_), .ZN(new_n17064_));
  AOI21_X1   g17000(.A1(new_n16943_), .A2(new_n17063_), .B(new_n17064_), .ZN(new_n17065_));
  INV_X1     g17001(.I(new_n17065_), .ZN(new_n17066_));
  AOI22_X1   g17002(.A1(new_n17062_), .A2(new_n17026_), .B1(new_n16953_), .B2(new_n17066_), .ZN(new_n17067_));
  NAND3_X1   g17003(.A1(new_n16977_), .A2(new_n16978_), .A3(new_n16979_), .ZN(new_n17068_));
  NAND2_X1   g17004(.A1(new_n13931_), .A2(new_n13930_), .ZN(new_n17069_));
  AOI21_X1   g17005(.A1(new_n16976_), .A2(new_n17068_), .B(new_n17069_), .ZN(new_n17070_));
  NOR2_X1    g17006(.A1(new_n13928_), .A2(new_n13927_), .ZN(new_n17071_));
  NOR3_X1    g17007(.A1(new_n17071_), .A2(new_n13918_), .A3(new_n13896_), .ZN(new_n17072_));
  OAI21_X1   g17008(.A1(new_n17070_), .A2(new_n17072_), .B(new_n13715_), .ZN(new_n17073_));
  OAI21_X1   g17009(.A1(new_n13896_), .A2(new_n13918_), .B(new_n17071_), .ZN(new_n17074_));
  NAND3_X1   g17010(.A1(new_n17069_), .A2(new_n17068_), .A3(new_n16976_), .ZN(new_n17075_));
  NAND3_X1   g17011(.A1(new_n17074_), .A2(new_n13734_), .A3(new_n17075_), .ZN(new_n17076_));
  AOI21_X1   g17012(.A1(new_n17076_), .A2(new_n17073_), .B(new_n13924_), .ZN(new_n17077_));
  AOI21_X1   g17013(.A1(new_n17074_), .A2(new_n17075_), .B(new_n13734_), .ZN(new_n17078_));
  NOR3_X1    g17014(.A1(new_n17070_), .A2(new_n17072_), .A3(new_n13715_), .ZN(new_n17079_));
  NOR3_X1    g17015(.A1(new_n17078_), .A2(new_n17079_), .A3(new_n13923_), .ZN(new_n17080_));
  NOR2_X1    g17016(.A1(new_n16958_), .A2(new_n16975_), .ZN(new_n17081_));
  NOR3_X1    g17017(.A1(new_n16956_), .A2(new_n16957_), .A3(new_n16986_), .ZN(new_n17082_));
  NOR3_X1    g17018(.A1(new_n16984_), .A2(new_n16980_), .A3(new_n17082_), .ZN(new_n17083_));
  OAI22_X1   g17019(.A1(new_n11264_), .A2(new_n4716_), .B1(new_n4719_), .B2(new_n11345_), .ZN(new_n17084_));
  NAND2_X1   g17020(.A1(new_n11354_), .A2(new_n4709_), .ZN(new_n17085_));
  AOI21_X1   g17021(.A1(new_n17085_), .A2(new_n17084_), .B(new_n4707_), .ZN(new_n17086_));
  NAND2_X1   g17022(.A1(new_n11678_), .A2(new_n17086_), .ZN(new_n17087_));
  XOR2_X1    g17023(.A1(new_n17087_), .A2(\a[11] ), .Z(new_n17088_));
  INV_X1     g17024(.I(new_n17088_), .ZN(new_n17089_));
  NOR3_X1    g17025(.A1(new_n17083_), .A2(new_n17081_), .A3(new_n17089_), .ZN(new_n17090_));
  INV_X1     g17026(.I(new_n17081_), .ZN(new_n17091_));
  INV_X1     g17027(.I(new_n17083_), .ZN(new_n17092_));
  AOI21_X1   g17028(.A1(new_n17092_), .A2(new_n17091_), .B(new_n17088_), .ZN(new_n17093_));
  OAI22_X1   g17029(.A1(new_n17077_), .A2(new_n17080_), .B1(new_n17093_), .B2(new_n17090_), .ZN(new_n17094_));
  OAI21_X1   g17030(.A1(new_n17078_), .A2(new_n17079_), .B(new_n13923_), .ZN(new_n17095_));
  NAND3_X1   g17031(.A1(new_n17076_), .A2(new_n17073_), .A3(new_n13924_), .ZN(new_n17096_));
  OAI21_X1   g17032(.A1(new_n17083_), .A2(new_n17081_), .B(new_n17088_), .ZN(new_n17097_));
  NAND3_X1   g17033(.A1(new_n17092_), .A2(new_n17091_), .A3(new_n17089_), .ZN(new_n17098_));
  NAND2_X1   g17034(.A1(new_n17098_), .A2(new_n17097_), .ZN(new_n17099_));
  NAND3_X1   g17035(.A1(new_n17099_), .A2(new_n17095_), .A3(new_n17096_), .ZN(new_n17100_));
  NAND2_X1   g17036(.A1(new_n17100_), .A2(new_n17094_), .ZN(new_n17101_));
  NOR2_X1    g17037(.A1(new_n16970_), .A2(new_n16964_), .ZN(new_n17102_));
  INV_X1     g17038(.I(new_n17102_), .ZN(new_n17103_));
  OAI21_X1   g17039(.A1(new_n16985_), .A2(new_n16992_), .B(new_n16958_), .ZN(new_n17104_));
  NAND3_X1   g17040(.A1(new_n17000_), .A2(new_n16999_), .A3(new_n16959_), .ZN(new_n17105_));
  NAND2_X1   g17041(.A1(new_n17104_), .A2(new_n17105_), .ZN(new_n17106_));
  NAND3_X1   g17042(.A1(new_n17106_), .A2(new_n16964_), .A3(new_n16970_), .ZN(new_n17107_));
  OAI22_X1   g17043(.A1(new_n11369_), .A2(new_n6783_), .B1(new_n6785_), .B2(new_n11461_), .ZN(new_n17108_));
  NAND2_X1   g17044(.A1(new_n11694_), .A2(new_n6789_), .ZN(new_n17109_));
  AOI21_X1   g17045(.A1(new_n17108_), .A2(new_n17109_), .B(new_n6776_), .ZN(new_n17110_));
  NAND2_X1   g17046(.A1(new_n12720_), .A2(new_n17110_), .ZN(new_n17111_));
  XOR2_X1    g17047(.A1(new_n17111_), .A2(\a[8] ), .Z(new_n17112_));
  NAND3_X1   g17048(.A1(new_n17107_), .A2(new_n17103_), .A3(new_n17112_), .ZN(new_n17113_));
  INV_X1     g17049(.I(new_n17113_), .ZN(new_n17114_));
  AOI21_X1   g17050(.A1(new_n17107_), .A2(new_n17103_), .B(new_n17112_), .ZN(new_n17115_));
  OAI21_X1   g17051(.A1(new_n17114_), .A2(new_n17115_), .B(new_n17101_), .ZN(new_n17116_));
  AND2_X2    g17052(.A1(new_n17100_), .A2(new_n17094_), .Z(new_n17117_));
  NAND2_X1   g17053(.A1(new_n17107_), .A2(new_n17103_), .ZN(new_n17118_));
  INV_X1     g17054(.I(new_n17112_), .ZN(new_n17119_));
  XOR2_X1    g17055(.A1(new_n17118_), .A2(new_n17119_), .Z(new_n17120_));
  NAND2_X1   g17056(.A1(new_n17120_), .A2(new_n17117_), .ZN(new_n17121_));
  NAND2_X1   g17057(.A1(new_n17121_), .A2(new_n17116_), .ZN(new_n17122_));
  AND3_X2    g17058(.A1(new_n11463_), .A2(new_n7530_), .A3(new_n12016_), .Z(new_n17123_));
  NOR4_X1    g17059(.A1(new_n11468_), .A2(new_n6776_), .A3(new_n11461_), .A4(new_n17123_), .ZN(new_n17124_));
  XOR2_X1    g17060(.A1(new_n17124_), .A2(new_n4009_), .Z(new_n17125_));
  OAI21_X1   g17061(.A1(new_n13716_), .A2(new_n13717_), .B(new_n13723_), .ZN(new_n17126_));
  AOI21_X1   g17062(.A1(new_n13725_), .A2(new_n17126_), .B(new_n13784_), .ZN(new_n17127_));
  OAI21_X1   g17063(.A1(new_n13716_), .A2(new_n13717_), .B(new_n13722_), .ZN(new_n17128_));
  NAND3_X1   g17064(.A1(new_n13736_), .A2(new_n13735_), .A3(new_n13723_), .ZN(new_n17129_));
  AOI21_X1   g17065(.A1(new_n17129_), .A2(new_n17128_), .B(new_n13464_), .ZN(new_n17130_));
  AOI21_X1   g17066(.A1(new_n17068_), .A2(new_n16976_), .B(new_n13923_), .ZN(new_n17131_));
  NAND3_X1   g17067(.A1(new_n17068_), .A2(new_n16976_), .A3(new_n13923_), .ZN(new_n17132_));
  NAND3_X1   g17068(.A1(new_n13931_), .A2(new_n13930_), .A3(new_n13734_), .ZN(new_n17133_));
  OAI21_X1   g17069(.A1(new_n13928_), .A2(new_n13927_), .B(new_n13715_), .ZN(new_n17134_));
  NAND2_X1   g17070(.A1(new_n17134_), .A2(new_n17133_), .ZN(new_n17135_));
  AOI21_X1   g17071(.A1(new_n17135_), .A2(new_n17132_), .B(new_n17131_), .ZN(new_n17136_));
  NOR3_X1    g17072(.A1(new_n17136_), .A2(new_n17127_), .A3(new_n17130_), .ZN(new_n17137_));
  AOI21_X1   g17073(.A1(new_n13778_), .A2(new_n13787_), .B(new_n13934_), .ZN(new_n17138_));
  NOR2_X1    g17074(.A1(new_n17138_), .A2(new_n17137_), .ZN(new_n17139_));
  AOI21_X1   g17075(.A1(new_n17095_), .A2(new_n17096_), .B(new_n17090_), .ZN(new_n17140_));
  OAI21_X1   g17076(.A1(new_n17140_), .A2(new_n17093_), .B(new_n17139_), .ZN(new_n17141_));
  INV_X1     g17077(.I(new_n17093_), .ZN(new_n17142_));
  NAND3_X1   g17078(.A1(new_n13934_), .A2(new_n13778_), .A3(new_n13787_), .ZN(new_n17143_));
  NAND2_X1   g17079(.A1(new_n13788_), .A2(new_n17136_), .ZN(new_n17144_));
  NAND2_X1   g17080(.A1(new_n17144_), .A2(new_n17143_), .ZN(new_n17145_));
  NAND3_X1   g17081(.A1(new_n17092_), .A2(new_n17091_), .A3(new_n17088_), .ZN(new_n17146_));
  OAI21_X1   g17082(.A1(new_n17077_), .A2(new_n17080_), .B(new_n17146_), .ZN(new_n17147_));
  NAND3_X1   g17083(.A1(new_n17147_), .A2(new_n17142_), .A3(new_n17145_), .ZN(new_n17148_));
  AOI21_X1   g17084(.A1(new_n17141_), .A2(new_n17148_), .B(new_n13940_), .ZN(new_n17149_));
  AOI21_X1   g17085(.A1(new_n17147_), .A2(new_n17142_), .B(new_n17145_), .ZN(new_n17150_));
  NOR3_X1    g17086(.A1(new_n17140_), .A2(new_n17093_), .A3(new_n17139_), .ZN(new_n17151_));
  NOR3_X1    g17087(.A1(new_n17150_), .A2(new_n17151_), .A3(new_n13939_), .ZN(new_n17152_));
  OAI21_X1   g17088(.A1(new_n17149_), .A2(new_n17152_), .B(new_n17125_), .ZN(new_n17153_));
  INV_X1     g17089(.I(new_n17125_), .ZN(new_n17154_));
  OAI21_X1   g17090(.A1(new_n17150_), .A2(new_n17151_), .B(new_n13939_), .ZN(new_n17155_));
  NAND3_X1   g17091(.A1(new_n17141_), .A2(new_n17148_), .A3(new_n13940_), .ZN(new_n17156_));
  NAND3_X1   g17092(.A1(new_n17155_), .A2(new_n17156_), .A3(new_n17154_), .ZN(new_n17157_));
  INV_X1     g17093(.I(new_n17115_), .ZN(new_n17158_));
  OAI21_X1   g17094(.A1(new_n17117_), .A2(new_n17114_), .B(new_n17158_), .ZN(new_n17159_));
  NAND3_X1   g17095(.A1(new_n17153_), .A2(new_n17157_), .A3(new_n17159_), .ZN(new_n17160_));
  AOI21_X1   g17096(.A1(new_n17155_), .A2(new_n17156_), .B(new_n17154_), .ZN(new_n17161_));
  NOR3_X1    g17097(.A1(new_n17149_), .A2(new_n17152_), .A3(new_n17125_), .ZN(new_n17162_));
  AOI21_X1   g17098(.A1(new_n17101_), .A2(new_n17113_), .B(new_n17115_), .ZN(new_n17163_));
  OAI21_X1   g17099(.A1(new_n17162_), .A2(new_n17161_), .B(new_n17163_), .ZN(new_n17164_));
  AOI21_X1   g17100(.A1(new_n16955_), .A2(new_n17059_), .B(new_n17024_), .ZN(new_n17165_));
  INV_X1     g17101(.I(new_n17165_), .ZN(new_n17166_));
  NAND3_X1   g17102(.A1(new_n17164_), .A2(new_n17160_), .A3(new_n17166_), .ZN(new_n17167_));
  NAND3_X1   g17103(.A1(new_n17067_), .A2(new_n17167_), .A3(new_n17122_), .ZN(new_n17168_));
  NOR3_X1    g17104(.A1(new_n17162_), .A2(new_n17161_), .A3(new_n17159_), .ZN(new_n17169_));
  INV_X1     g17105(.I(new_n17169_), .ZN(new_n17170_));
  NAND3_X1   g17106(.A1(new_n13950_), .A2(new_n13953_), .A3(new_n13958_), .ZN(new_n17171_));
  INV_X1     g17107(.I(new_n17171_), .ZN(new_n17172_));
  AOI21_X1   g17108(.A1(new_n13950_), .A2(new_n13953_), .B(new_n13958_), .ZN(new_n17173_));
  OAI21_X1   g17109(.A1(new_n17172_), .A2(new_n17173_), .B(new_n13943_), .ZN(new_n17174_));
  INV_X1     g17110(.I(new_n13943_), .ZN(new_n17175_));
  INV_X1     g17111(.I(new_n13963_), .ZN(new_n17176_));
  OAI21_X1   g17112(.A1(new_n17176_), .A2(new_n13960_), .B(new_n17175_), .ZN(new_n17177_));
  NAND2_X1   g17113(.A1(new_n17174_), .A2(new_n17177_), .ZN(new_n17178_));
  NAND3_X1   g17114(.A1(new_n17168_), .A2(new_n17170_), .A3(new_n17178_), .ZN(new_n17179_));
  AOI21_X1   g17115(.A1(new_n17168_), .A2(new_n17170_), .B(new_n17178_), .ZN(new_n17180_));
  NOR3_X1    g17116(.A1(new_n17055_), .A2(new_n17058_), .A3(new_n17061_), .ZN(new_n17181_));
  AOI21_X1   g17117(.A1(new_n17021_), .A2(new_n17025_), .B(new_n16953_), .ZN(new_n17182_));
  OAI22_X1   g17118(.A1(new_n17182_), .A2(new_n17181_), .B1(new_n17055_), .B2(new_n17065_), .ZN(new_n17183_));
  INV_X1     g17119(.I(new_n17122_), .ZN(new_n17184_));
  NOR3_X1    g17120(.A1(new_n17162_), .A2(new_n17161_), .A3(new_n17163_), .ZN(new_n17185_));
  AOI21_X1   g17121(.A1(new_n17153_), .A2(new_n17157_), .B(new_n17159_), .ZN(new_n17186_));
  NOR3_X1    g17122(.A1(new_n17185_), .A2(new_n17186_), .A3(new_n17165_), .ZN(new_n17187_));
  NOR3_X1    g17123(.A1(new_n17183_), .A2(new_n17187_), .A3(new_n17184_), .ZN(new_n17188_));
  INV_X1     g17124(.I(new_n17173_), .ZN(new_n17189_));
  AOI21_X1   g17125(.A1(new_n17189_), .A2(new_n17171_), .B(new_n17175_), .ZN(new_n17190_));
  AOI21_X1   g17126(.A1(new_n13961_), .A2(new_n13963_), .B(new_n13943_), .ZN(new_n17191_));
  NOR2_X1    g17127(.A1(new_n17190_), .A2(new_n17191_), .ZN(new_n17192_));
  NOR3_X1    g17128(.A1(new_n17188_), .A2(new_n17169_), .A3(new_n17192_), .ZN(new_n17193_));
  AOI21_X1   g17129(.A1(new_n17147_), .A2(new_n17142_), .B(new_n17125_), .ZN(new_n17194_));
  NOR3_X1    g17130(.A1(new_n17140_), .A2(new_n17093_), .A3(new_n17154_), .ZN(new_n17195_));
  XOR2_X1    g17131(.A1(new_n17145_), .A2(new_n13939_), .Z(new_n17196_));
  NOR2_X1    g17132(.A1(new_n17196_), .A2(new_n17195_), .ZN(new_n17197_));
  NOR2_X1    g17133(.A1(new_n17197_), .A2(new_n17194_), .ZN(new_n17198_));
  OAI21_X1   g17134(.A1(new_n17193_), .A2(new_n17180_), .B(new_n17198_), .ZN(new_n17199_));
  NAND2_X1   g17135(.A1(new_n13962_), .A2(new_n13963_), .ZN(new_n17200_));
  XNOR2_X1   g17136(.A1(new_n13777_), .A2(new_n17200_), .ZN(new_n17201_));
  NAND3_X1   g17137(.A1(new_n17199_), .A2(new_n17179_), .A3(new_n17201_), .ZN(new_n17202_));
  NAND3_X1   g17138(.A1(new_n17202_), .A2(new_n13767_), .A3(new_n13964_), .ZN(new_n17203_));
  INV_X1     g17139(.I(new_n13419_), .ZN(new_n17204_));
  INV_X1     g17140(.I(new_n13422_), .ZN(new_n17205_));
  NAND3_X1   g17141(.A1(new_n17204_), .A2(new_n17205_), .A3(new_n13763_), .ZN(new_n17206_));
  INV_X1     g17142(.I(new_n13232_), .ZN(new_n17207_));
  NAND2_X1   g17143(.A1(new_n13241_), .A2(new_n13244_), .ZN(new_n17208_));
  NOR2_X1    g17144(.A1(new_n17208_), .A2(new_n13250_), .ZN(new_n17209_));
  AOI21_X1   g17145(.A1(new_n13241_), .A2(new_n13244_), .B(new_n13249_), .ZN(new_n17210_));
  OAI21_X1   g17146(.A1(new_n17209_), .A2(new_n17210_), .B(new_n17207_), .ZN(new_n17211_));
  OAI21_X1   g17147(.A1(new_n13254_), .A2(new_n13251_), .B(new_n13232_), .ZN(new_n17212_));
  NAND2_X1   g17148(.A1(new_n17211_), .A2(new_n17212_), .ZN(new_n17213_));
  NAND3_X1   g17149(.A1(new_n17203_), .A2(new_n17206_), .A3(new_n17213_), .ZN(new_n17214_));
  AOI21_X1   g17150(.A1(new_n17203_), .A2(new_n17206_), .B(new_n17213_), .ZN(new_n17215_));
  INV_X1     g17151(.I(new_n13764_), .ZN(new_n17216_));
  NAND2_X1   g17152(.A1(new_n17216_), .A2(new_n13765_), .ZN(new_n17217_));
  NAND2_X1   g17153(.A1(new_n17168_), .A2(new_n17170_), .ZN(new_n17218_));
  OAI21_X1   g17154(.A1(new_n17188_), .A2(new_n17169_), .B(new_n17192_), .ZN(new_n17219_));
  NAND3_X1   g17155(.A1(new_n17168_), .A2(new_n17170_), .A3(new_n17178_), .ZN(new_n17220_));
  INV_X1     g17156(.I(new_n17198_), .ZN(new_n17221_));
  AOI22_X1   g17157(.A1(new_n17219_), .A2(new_n17220_), .B1(new_n17218_), .B2(new_n17221_), .ZN(new_n17222_));
  XOR2_X1    g17158(.A1(new_n13777_), .A2(new_n17200_), .Z(new_n17223_));
  OAI21_X1   g17159(.A1(new_n17222_), .A2(new_n17223_), .B(new_n13964_), .ZN(new_n17224_));
  OAI21_X1   g17160(.A1(new_n17224_), .A2(new_n17217_), .B(new_n17206_), .ZN(new_n17225_));
  INV_X1     g17161(.I(new_n17213_), .ZN(new_n17226_));
  NOR2_X1    g17162(.A1(new_n17225_), .A2(new_n17226_), .ZN(new_n17227_));
  NAND2_X1   g17163(.A1(new_n13412_), .A2(new_n13398_), .ZN(new_n17228_));
  AND2_X2    g17164(.A1(new_n17228_), .A2(new_n13418_), .Z(new_n17229_));
  OAI21_X1   g17165(.A1(new_n17227_), .A2(new_n17215_), .B(new_n17229_), .ZN(new_n17230_));
  NOR2_X1    g17166(.A1(new_n13252_), .A2(new_n13254_), .ZN(new_n17231_));
  AOI21_X1   g17167(.A1(new_n12733_), .A2(new_n12736_), .B(new_n17231_), .ZN(new_n17232_));
  NOR2_X1    g17168(.A1(new_n13255_), .A2(new_n17232_), .ZN(new_n17233_));
  NAND3_X1   g17169(.A1(new_n17230_), .A2(new_n17214_), .A3(new_n17233_), .ZN(new_n17234_));
  NAND3_X1   g17170(.A1(new_n17234_), .A2(new_n12731_), .A3(new_n13256_), .ZN(new_n17235_));
  NOR2_X1    g17171(.A1(new_n12730_), .A2(new_n12612_), .ZN(new_n17236_));
  INV_X1     g17172(.I(new_n17236_), .ZN(new_n17237_));
  NAND2_X1   g17173(.A1(new_n17235_), .A2(new_n17237_), .ZN(new_n17238_));
  INV_X1     g17174(.I(new_n12731_), .ZN(new_n17239_));
  NAND2_X1   g17175(.A1(new_n17225_), .A2(new_n17226_), .ZN(new_n17240_));
  NAND3_X1   g17176(.A1(new_n17203_), .A2(new_n17206_), .A3(new_n17213_), .ZN(new_n17241_));
  INV_X1     g17177(.I(new_n17229_), .ZN(new_n17242_));
  AOI22_X1   g17178(.A1(new_n17240_), .A2(new_n17241_), .B1(new_n17225_), .B2(new_n17242_), .ZN(new_n17243_));
  OAI21_X1   g17179(.A1(new_n17243_), .A2(new_n17232_), .B(new_n13256_), .ZN(new_n17244_));
  NOR2_X1    g17180(.A1(new_n17244_), .A2(new_n17239_), .ZN(new_n17245_));
  INV_X1     g17181(.I(new_n12594_), .ZN(new_n17246_));
  AOI21_X1   g17182(.A1(new_n17246_), .A2(new_n12599_), .B(new_n12596_), .ZN(new_n17247_));
  INV_X1     g17183(.I(new_n17247_), .ZN(new_n17248_));
  OAI21_X1   g17184(.A1(new_n12497_), .A2(new_n12536_), .B(new_n12538_), .ZN(new_n17249_));
  AOI21_X1   g17185(.A1(new_n11495_), .A2(new_n11504_), .B(new_n11503_), .ZN(new_n17250_));
  XNOR2_X1   g17186(.A1(new_n11483_), .A2(new_n11493_), .ZN(new_n17251_));
  NOR3_X1    g17187(.A1(new_n11502_), .A2(new_n11500_), .A3(new_n17251_), .ZN(new_n17252_));
  NOR2_X1    g17188(.A1(new_n17250_), .A2(new_n17252_), .ZN(new_n17253_));
  NAND3_X1   g17189(.A1(new_n12500_), .A2(new_n12504_), .A3(new_n12527_), .ZN(new_n17254_));
  NAND2_X1   g17190(.A1(new_n17254_), .A2(new_n12528_), .ZN(new_n17255_));
  NOR2_X1    g17191(.A1(new_n8725_), .A2(new_n2767_), .ZN(new_n17256_));
  NOR2_X1    g17192(.A1(new_n8718_), .A2(new_n2772_), .ZN(new_n17257_));
  NOR2_X1    g17193(.A1(new_n8735_), .A2(new_n2771_), .ZN(new_n17258_));
  NOR4_X1    g17194(.A1(new_n17256_), .A2(new_n2763_), .A3(new_n17257_), .A4(new_n17258_), .ZN(new_n17259_));
  NAND2_X1   g17195(.A1(new_n12242_), .A2(new_n17259_), .ZN(new_n17260_));
  XOR2_X1    g17196(.A1(new_n17255_), .A2(new_n17260_), .Z(new_n17261_));
  NOR2_X1    g17197(.A1(new_n17253_), .A2(new_n17261_), .ZN(new_n17262_));
  INV_X1     g17198(.I(new_n17253_), .ZN(new_n17263_));
  INV_X1     g17199(.I(new_n17255_), .ZN(new_n17264_));
  NOR2_X1    g17200(.A1(new_n17264_), .A2(new_n17260_), .ZN(new_n17265_));
  INV_X1     g17201(.I(new_n17265_), .ZN(new_n17266_));
  NAND2_X1   g17202(.A1(new_n17264_), .A2(new_n17260_), .ZN(new_n17267_));
  AOI21_X1   g17203(.A1(new_n17266_), .A2(new_n17267_), .B(new_n17263_), .ZN(new_n17268_));
  NOR2_X1    g17204(.A1(new_n17268_), .A2(new_n17262_), .ZN(new_n17269_));
  OAI22_X1   g17205(.A1(new_n2742_), .A2(new_n8701_), .B1(new_n8710_), .B2(new_n2747_), .ZN(new_n17270_));
  NAND2_X1   g17206(.A1(new_n8696_), .A2(new_n2750_), .ZN(new_n17271_));
  AOI21_X1   g17207(.A1(new_n17270_), .A2(new_n17271_), .B(new_n2737_), .ZN(new_n17272_));
  NAND2_X1   g17208(.A1(new_n11595_), .A2(new_n17272_), .ZN(new_n17273_));
  XOR2_X1    g17209(.A1(new_n17273_), .A2(\a[29] ), .Z(new_n17274_));
  INV_X1     g17210(.I(new_n17274_), .ZN(new_n17275_));
  XOR2_X1    g17211(.A1(new_n17269_), .A2(new_n17275_), .Z(new_n17276_));
  INV_X1     g17212(.I(new_n17276_), .ZN(new_n17277_));
  XOR2_X1    g17213(.A1(new_n17269_), .A2(new_n17274_), .Z(new_n17278_));
  NOR2_X1    g17214(.A1(new_n17249_), .A2(new_n17278_), .ZN(new_n17279_));
  AOI21_X1   g17215(.A1(new_n17249_), .A2(new_n17277_), .B(new_n17279_), .ZN(new_n17280_));
  INV_X1     g17216(.I(new_n17280_), .ZN(new_n17281_));
  AOI21_X1   g17217(.A1(new_n12540_), .A2(new_n12554_), .B(new_n12553_), .ZN(new_n17282_));
  OAI22_X1   g17218(.A1(new_n3268_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n3322_), .ZN(new_n17283_));
  NAND2_X1   g17219(.A1(new_n8674_), .A2(new_n3317_), .ZN(new_n17284_));
  AOI21_X1   g17220(.A1(new_n17284_), .A2(new_n17283_), .B(new_n3260_), .ZN(new_n17285_));
  NAND2_X1   g17221(.A1(new_n11431_), .A2(new_n17285_), .ZN(new_n17286_));
  XOR2_X1    g17222(.A1(new_n17286_), .A2(\a[26] ), .Z(new_n17287_));
  NOR2_X1    g17223(.A1(new_n17282_), .A2(new_n17287_), .ZN(new_n17288_));
  AND2_X2    g17224(.A1(new_n17282_), .A2(new_n17287_), .Z(new_n17289_));
  OAI21_X1   g17225(.A1(new_n17289_), .A2(new_n17288_), .B(new_n17281_), .ZN(new_n17290_));
  XNOR2_X1   g17226(.A1(new_n17282_), .A2(new_n17287_), .ZN(new_n17291_));
  OAI21_X1   g17227(.A1(new_n17281_), .A2(new_n17291_), .B(new_n17290_), .ZN(new_n17292_));
  NOR2_X1    g17228(.A1(new_n12568_), .A2(new_n12558_), .ZN(new_n17293_));
  NOR2_X1    g17229(.A1(new_n17293_), .A2(new_n12570_), .ZN(new_n17294_));
  OAI22_X1   g17230(.A1(new_n11284_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n8661_), .ZN(new_n17295_));
  NAND2_X1   g17231(.A1(new_n11272_), .A2(new_n3312_), .ZN(new_n17296_));
  AOI21_X1   g17232(.A1(new_n17295_), .A2(new_n17296_), .B(new_n3302_), .ZN(new_n17297_));
  NAND2_X1   g17233(.A1(new_n11655_), .A2(new_n17297_), .ZN(new_n17298_));
  XOR2_X1    g17234(.A1(new_n17298_), .A2(\a[23] ), .Z(new_n17299_));
  XOR2_X1    g17235(.A1(new_n17294_), .A2(new_n17299_), .Z(new_n17300_));
  INV_X1     g17236(.I(new_n17300_), .ZN(new_n17301_));
  XNOR2_X1   g17237(.A1(new_n17294_), .A2(new_n17299_), .ZN(new_n17302_));
  NOR2_X1    g17238(.A1(new_n17302_), .A2(new_n17292_), .ZN(new_n17303_));
  AOI21_X1   g17239(.A1(new_n17292_), .A2(new_n17301_), .B(new_n17303_), .ZN(new_n17304_));
  INV_X1     g17240(.I(new_n12582_), .ZN(new_n17305_));
  AOI21_X1   g17241(.A1(new_n17305_), .A2(new_n12573_), .B(new_n12583_), .ZN(new_n17306_));
  OAI22_X1   g17242(.A1(new_n11264_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n11277_), .ZN(new_n17307_));
  NAND2_X1   g17243(.A1(new_n11346_), .A2(new_n4096_), .ZN(new_n17308_));
  AOI21_X1   g17244(.A1(new_n17307_), .A2(new_n17308_), .B(new_n4095_), .ZN(new_n17309_));
  NAND2_X1   g17245(.A1(new_n11757_), .A2(new_n17309_), .ZN(new_n17310_));
  XOR2_X1    g17246(.A1(new_n17310_), .A2(\a[20] ), .Z(new_n17311_));
  AND2_X2    g17247(.A1(new_n17306_), .A2(new_n17311_), .Z(new_n17312_));
  NOR2_X1    g17248(.A1(new_n17306_), .A2(new_n17311_), .ZN(new_n17313_));
  NOR2_X1    g17249(.A1(new_n17312_), .A2(new_n17313_), .ZN(new_n17314_));
  NOR2_X1    g17250(.A1(new_n17314_), .A2(new_n17304_), .ZN(new_n17315_));
  XNOR2_X1   g17251(.A1(new_n17306_), .A2(new_n17311_), .ZN(new_n17316_));
  INV_X1     g17252(.I(new_n17316_), .ZN(new_n17317_));
  AOI21_X1   g17253(.A1(new_n17304_), .A2(new_n17317_), .B(new_n17315_), .ZN(new_n17318_));
  OAI22_X1   g17254(.A1(new_n11353_), .A2(new_n4291_), .B1(new_n4470_), .B2(new_n11697_), .ZN(new_n17319_));
  NAND2_X1   g17255(.A1(new_n11370_), .A2(new_n4298_), .ZN(new_n17320_));
  AOI21_X1   g17256(.A1(new_n17320_), .A2(new_n17319_), .B(new_n4468_), .ZN(new_n17321_));
  NAND2_X1   g17257(.A1(new_n11700_), .A2(new_n17321_), .ZN(new_n17322_));
  XOR2_X1    g17258(.A1(new_n17322_), .A2(\a[17] ), .Z(new_n17323_));
  XOR2_X1    g17259(.A1(new_n17318_), .A2(new_n17323_), .Z(new_n17324_));
  INV_X1     g17260(.I(new_n17324_), .ZN(new_n17325_));
  INV_X1     g17261(.I(new_n17323_), .ZN(new_n17326_));
  NOR2_X1    g17262(.A1(new_n17318_), .A2(new_n17326_), .ZN(new_n17327_));
  INV_X1     g17263(.I(new_n17327_), .ZN(new_n17328_));
  NAND2_X1   g17264(.A1(new_n17318_), .A2(new_n17326_), .ZN(new_n17329_));
  AOI21_X1   g17265(.A1(new_n17328_), .A2(new_n17329_), .B(new_n17248_), .ZN(new_n17330_));
  AOI21_X1   g17266(.A1(new_n17325_), .A2(new_n17248_), .B(new_n17330_), .ZN(new_n17331_));
  OAI21_X1   g17267(.A1(new_n17245_), .A2(new_n17236_), .B(new_n17331_), .ZN(new_n17332_));
  INV_X1     g17268(.I(new_n17331_), .ZN(new_n17333_));
  NAND3_X1   g17269(.A1(new_n17235_), .A2(new_n17237_), .A3(new_n17333_), .ZN(new_n17334_));
  INV_X1     g17270(.I(new_n12608_), .ZN(new_n17335_));
  AOI21_X1   g17271(.A1(new_n17335_), .A2(new_n12493_), .B(new_n12609_), .ZN(new_n17336_));
  INV_X1     g17272(.I(new_n17336_), .ZN(new_n17337_));
  AOI22_X1   g17273(.A1(new_n17332_), .A2(new_n17334_), .B1(new_n17238_), .B2(new_n17337_), .ZN(new_n17338_));
  OAI21_X1   g17274(.A1(new_n17247_), .A2(new_n17327_), .B(new_n17329_), .ZN(new_n17339_));
  INV_X1     g17275(.I(new_n17269_), .ZN(new_n17340_));
  OAI21_X1   g17276(.A1(new_n17340_), .A2(new_n17275_), .B(new_n17249_), .ZN(new_n17341_));
  OAI21_X1   g17277(.A1(new_n17269_), .A2(new_n17274_), .B(new_n17341_), .ZN(new_n17342_));
  AOI21_X1   g17278(.A1(new_n17253_), .A2(new_n17267_), .B(new_n17265_), .ZN(new_n17343_));
  XOR2_X1    g17279(.A1(new_n11544_), .A2(new_n11530_), .Z(new_n17344_));
  INV_X1     g17280(.I(new_n17344_), .ZN(new_n17345_));
  AOI21_X1   g17281(.A1(new_n11541_), .A2(new_n11546_), .B(new_n11506_), .ZN(new_n17346_));
  AOI21_X1   g17282(.A1(new_n11506_), .A2(new_n17345_), .B(new_n17346_), .ZN(new_n17347_));
  OAI22_X1   g17283(.A1(new_n8701_), .A2(new_n2747_), .B1(new_n8694_), .B2(new_n2742_), .ZN(new_n17348_));
  NAND2_X1   g17284(.A1(new_n8682_), .A2(new_n2750_), .ZN(new_n17349_));
  AOI21_X1   g17285(.A1(new_n17349_), .A2(new_n17348_), .B(new_n2737_), .ZN(new_n17350_));
  NAND2_X1   g17286(.A1(new_n12347_), .A2(new_n17350_), .ZN(new_n17351_));
  XOR2_X1    g17287(.A1(new_n17351_), .A2(\a[29] ), .Z(new_n17352_));
  XOR2_X1    g17288(.A1(new_n17347_), .A2(new_n17352_), .Z(new_n17353_));
  NOR2_X1    g17289(.A1(new_n17353_), .A2(new_n17343_), .ZN(new_n17354_));
  INV_X1     g17290(.I(new_n17343_), .ZN(new_n17355_));
  INV_X1     g17291(.I(new_n17352_), .ZN(new_n17356_));
  NOR2_X1    g17292(.A1(new_n17347_), .A2(new_n17356_), .ZN(new_n17357_));
  INV_X1     g17293(.I(new_n17357_), .ZN(new_n17358_));
  NAND2_X1   g17294(.A1(new_n17347_), .A2(new_n17356_), .ZN(new_n17359_));
  AOI21_X1   g17295(.A1(new_n17358_), .A2(new_n17359_), .B(new_n17355_), .ZN(new_n17360_));
  NOR2_X1    g17296(.A1(new_n17354_), .A2(new_n17360_), .ZN(new_n17361_));
  OAI22_X1   g17297(.A1(new_n8673_), .A2(new_n3322_), .B1(new_n8687_), .B2(new_n3268_), .ZN(new_n17362_));
  NAND2_X1   g17298(.A1(new_n8662_), .A2(new_n3317_), .ZN(new_n17363_));
  AOI21_X1   g17299(.A1(new_n17363_), .A2(new_n17362_), .B(new_n3260_), .ZN(new_n17364_));
  NAND2_X1   g17300(.A1(new_n11624_), .A2(new_n17364_), .ZN(new_n17365_));
  XOR2_X1    g17301(.A1(new_n17365_), .A2(\a[26] ), .Z(new_n17366_));
  INV_X1     g17302(.I(new_n17366_), .ZN(new_n17367_));
  NOR2_X1    g17303(.A1(new_n17361_), .A2(new_n17367_), .ZN(new_n17368_));
  NOR3_X1    g17304(.A1(new_n17354_), .A2(new_n17360_), .A3(new_n17366_), .ZN(new_n17369_));
  NOR2_X1    g17305(.A1(new_n17368_), .A2(new_n17369_), .ZN(new_n17370_));
  INV_X1     g17306(.I(new_n17370_), .ZN(new_n17371_));
  XOR2_X1    g17307(.A1(new_n17361_), .A2(new_n17366_), .Z(new_n17372_));
  NOR2_X1    g17308(.A1(new_n17342_), .A2(new_n17372_), .ZN(new_n17373_));
  AOI21_X1   g17309(.A1(new_n17342_), .A2(new_n17371_), .B(new_n17373_), .ZN(new_n17374_));
  NOR2_X1    g17310(.A1(new_n17289_), .A2(new_n17281_), .ZN(new_n17375_));
  NOR2_X1    g17311(.A1(new_n17375_), .A2(new_n17288_), .ZN(new_n17376_));
  OAI22_X1   g17312(.A1(new_n11284_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n11271_), .ZN(new_n17377_));
  NAND2_X1   g17313(.A1(new_n11311_), .A2(new_n3312_), .ZN(new_n17378_));
  AOI21_X1   g17314(.A1(new_n17377_), .A2(new_n17378_), .B(new_n3302_), .ZN(new_n17379_));
  NAND2_X1   g17315(.A1(new_n11391_), .A2(new_n17379_), .ZN(new_n17380_));
  XOR2_X1    g17316(.A1(new_n17380_), .A2(\a[23] ), .Z(new_n17381_));
  AND2_X2    g17317(.A1(new_n17376_), .A2(new_n17381_), .Z(new_n17382_));
  NOR2_X1    g17318(.A1(new_n17376_), .A2(new_n17381_), .ZN(new_n17383_));
  NOR2_X1    g17319(.A1(new_n17382_), .A2(new_n17383_), .ZN(new_n17384_));
  NOR2_X1    g17320(.A1(new_n17384_), .A2(new_n17374_), .ZN(new_n17385_));
  XOR2_X1    g17321(.A1(new_n17376_), .A2(new_n17381_), .Z(new_n17386_));
  AOI21_X1   g17322(.A1(new_n17374_), .A2(new_n17386_), .B(new_n17385_), .ZN(new_n17387_));
  OAI22_X1   g17323(.A1(new_n11264_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n11345_), .ZN(new_n17388_));
  NAND2_X1   g17324(.A1(new_n11354_), .A2(new_n4096_), .ZN(new_n17389_));
  AOI21_X1   g17325(.A1(new_n17389_), .A2(new_n17388_), .B(new_n4095_), .ZN(new_n17390_));
  NAND2_X1   g17326(.A1(new_n11678_), .A2(new_n17390_), .ZN(new_n17391_));
  XOR2_X1    g17327(.A1(new_n17391_), .A2(\a[20] ), .Z(new_n17392_));
  NAND2_X1   g17328(.A1(new_n17292_), .A2(new_n17299_), .ZN(new_n17393_));
  XOR2_X1    g17329(.A1(new_n17292_), .A2(new_n17299_), .Z(new_n17394_));
  NAND2_X1   g17330(.A1(new_n17394_), .A2(new_n17294_), .ZN(new_n17395_));
  NAND2_X1   g17331(.A1(new_n17395_), .A2(new_n17393_), .ZN(new_n17396_));
  XOR2_X1    g17332(.A1(new_n17396_), .A2(new_n17392_), .Z(new_n17397_));
  XNOR2_X1   g17333(.A1(new_n17397_), .A2(new_n17387_), .ZN(new_n17398_));
  INV_X1     g17334(.I(new_n17312_), .ZN(new_n17399_));
  AOI21_X1   g17335(.A1(new_n17399_), .A2(new_n17304_), .B(new_n17313_), .ZN(new_n17400_));
  OAI22_X1   g17336(.A1(new_n11369_), .A2(new_n4291_), .B1(new_n4470_), .B2(new_n11461_), .ZN(new_n17401_));
  NAND2_X1   g17337(.A1(new_n11694_), .A2(new_n4298_), .ZN(new_n17402_));
  AOI21_X1   g17338(.A1(new_n17401_), .A2(new_n17402_), .B(new_n4468_), .ZN(new_n17403_));
  NAND2_X1   g17339(.A1(new_n12720_), .A2(new_n17403_), .ZN(new_n17404_));
  XOR2_X1    g17340(.A1(new_n17404_), .A2(\a[17] ), .Z(new_n17405_));
  AND2_X2    g17341(.A1(new_n17400_), .A2(new_n17405_), .Z(new_n17406_));
  NOR2_X1    g17342(.A1(new_n17400_), .A2(new_n17405_), .ZN(new_n17407_));
  NOR2_X1    g17343(.A1(new_n17406_), .A2(new_n17407_), .ZN(new_n17408_));
  NOR2_X1    g17344(.A1(new_n17408_), .A2(new_n17398_), .ZN(new_n17409_));
  INV_X1     g17345(.I(new_n17398_), .ZN(new_n17410_));
  XNOR2_X1   g17346(.A1(new_n17400_), .A2(new_n17405_), .ZN(new_n17411_));
  NOR2_X1    g17347(.A1(new_n17411_), .A2(new_n17410_), .ZN(new_n17412_));
  NOR2_X1    g17348(.A1(new_n17409_), .A2(new_n17412_), .ZN(new_n17413_));
  INV_X1     g17349(.I(new_n17413_), .ZN(new_n17414_));
  NOR2_X1    g17350(.A1(new_n17414_), .A2(new_n17339_), .ZN(new_n17415_));
  INV_X1     g17351(.I(new_n17415_), .ZN(new_n17416_));
  INV_X1     g17352(.I(new_n17339_), .ZN(new_n17417_));
  NOR2_X1    g17353(.A1(new_n17413_), .A2(new_n17417_), .ZN(new_n17418_));
  AOI21_X1   g17354(.A1(new_n17338_), .A2(new_n17416_), .B(new_n17418_), .ZN(new_n17419_));
  INV_X1     g17355(.I(new_n17392_), .ZN(new_n17420_));
  XOR2_X1    g17356(.A1(new_n17387_), .A2(new_n17420_), .Z(new_n17421_));
  AOI21_X1   g17357(.A1(new_n17420_), .A2(new_n17396_), .B(new_n17421_), .ZN(new_n17422_));
  INV_X1     g17358(.I(new_n17422_), .ZN(new_n17423_));
  INV_X1     g17359(.I(new_n17368_), .ZN(new_n17424_));
  AOI21_X1   g17360(.A1(new_n17342_), .A2(new_n17424_), .B(new_n17369_), .ZN(new_n17425_));
  AOI22_X1   g17361(.A1(new_n11542_), .A2(new_n11546_), .B1(new_n11562_), .B2(new_n11563_), .ZN(new_n17426_));
  XOR2_X1    g17362(.A1(new_n11530_), .A2(new_n11560_), .Z(new_n17427_));
  NOR2_X1    g17363(.A1(new_n11547_), .A2(new_n17427_), .ZN(new_n17428_));
  NOR2_X1    g17364(.A1(new_n17428_), .A2(new_n17426_), .ZN(new_n17429_));
  INV_X1     g17365(.I(new_n17429_), .ZN(new_n17430_));
  OAI22_X1   g17366(.A1(new_n8681_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8694_), .ZN(new_n17431_));
  NAND2_X1   g17367(.A1(new_n8688_), .A2(new_n2750_), .ZN(new_n17432_));
  AOI21_X1   g17368(.A1(new_n17432_), .A2(new_n17431_), .B(new_n2737_), .ZN(new_n17433_));
  NAND2_X1   g17369(.A1(new_n11420_), .A2(new_n17433_), .ZN(new_n17434_));
  XOR2_X1    g17370(.A1(new_n17434_), .A2(\a[29] ), .Z(new_n17435_));
  NOR2_X1    g17371(.A1(new_n8701_), .A2(new_n2772_), .ZN(new_n17436_));
  AOI21_X1   g17372(.A1(new_n8719_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n17437_));
  OAI21_X1   g17373(.A1(new_n8710_), .A2(new_n2767_), .B(new_n17437_), .ZN(new_n17438_));
  NOR3_X1    g17374(.A1(new_n12205_), .A2(new_n17436_), .A3(new_n17438_), .ZN(new_n17439_));
  INV_X1     g17375(.I(new_n17439_), .ZN(new_n17440_));
  XOR2_X1    g17376(.A1(new_n17435_), .A2(new_n17440_), .Z(new_n17441_));
  NAND2_X1   g17377(.A1(new_n17441_), .A2(new_n17430_), .ZN(new_n17442_));
  NAND2_X1   g17378(.A1(new_n17435_), .A2(new_n17440_), .ZN(new_n17443_));
  NOR2_X1    g17379(.A1(new_n17435_), .A2(new_n17440_), .ZN(new_n17444_));
  INV_X1     g17380(.I(new_n17444_), .ZN(new_n17445_));
  NAND2_X1   g17381(.A1(new_n17445_), .A2(new_n17443_), .ZN(new_n17446_));
  NAND2_X1   g17382(.A1(new_n17446_), .A2(new_n17429_), .ZN(new_n17447_));
  NAND2_X1   g17383(.A1(new_n17447_), .A2(new_n17442_), .ZN(new_n17448_));
  OAI21_X1   g17384(.A1(new_n17343_), .A2(new_n17357_), .B(new_n17359_), .ZN(new_n17449_));
  INV_X1     g17385(.I(new_n17449_), .ZN(new_n17450_));
  OAI22_X1   g17386(.A1(new_n8661_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8673_), .ZN(new_n17451_));
  NAND2_X1   g17387(.A1(new_n11285_), .A2(new_n3317_), .ZN(new_n17452_));
  AOI21_X1   g17388(.A1(new_n17452_), .A2(new_n17451_), .B(new_n3260_), .ZN(new_n17453_));
  NAND2_X1   g17389(.A1(new_n11323_), .A2(new_n17453_), .ZN(new_n17454_));
  XOR2_X1    g17390(.A1(new_n17454_), .A2(\a[26] ), .Z(new_n17455_));
  XOR2_X1    g17391(.A1(new_n17455_), .A2(new_n17450_), .Z(new_n17456_));
  NAND2_X1   g17392(.A1(new_n17456_), .A2(new_n17448_), .ZN(new_n17457_));
  NOR2_X1    g17393(.A1(new_n17455_), .A2(new_n17450_), .ZN(new_n17458_));
  AND2_X2    g17394(.A1(new_n17455_), .A2(new_n17450_), .Z(new_n17459_));
  NOR2_X1    g17395(.A1(new_n17459_), .A2(new_n17458_), .ZN(new_n17460_));
  OAI21_X1   g17396(.A1(new_n17448_), .A2(new_n17460_), .B(new_n17457_), .ZN(new_n17461_));
  AOI22_X1   g17397(.A1(new_n11311_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n11272_), .ZN(new_n17462_));
  NOR2_X1    g17398(.A1(new_n11264_), .A2(new_n3780_), .ZN(new_n17463_));
  OAI21_X1   g17399(.A1(new_n17463_), .A2(new_n17462_), .B(new_n3301_), .ZN(new_n17464_));
  NOR2_X1    g17400(.A1(new_n11310_), .A2(new_n17464_), .ZN(new_n17465_));
  XOR2_X1    g17401(.A1(new_n17465_), .A2(new_n84_), .Z(new_n17466_));
  INV_X1     g17402(.I(new_n17466_), .ZN(new_n17467_));
  NOR2_X1    g17403(.A1(new_n17467_), .A2(new_n17461_), .ZN(new_n17468_));
  INV_X1     g17404(.I(new_n17468_), .ZN(new_n17469_));
  NAND2_X1   g17405(.A1(new_n17467_), .A2(new_n17461_), .ZN(new_n17470_));
  AOI21_X1   g17406(.A1(new_n17469_), .A2(new_n17470_), .B(new_n17425_), .ZN(new_n17471_));
  XOR2_X1    g17407(.A1(new_n17461_), .A2(new_n17466_), .Z(new_n17472_));
  INV_X1     g17408(.I(new_n17472_), .ZN(new_n17473_));
  AOI21_X1   g17409(.A1(new_n17473_), .A2(new_n17425_), .B(new_n17471_), .ZN(new_n17474_));
  NOR2_X1    g17410(.A1(new_n17382_), .A2(new_n17374_), .ZN(new_n17475_));
  NOR2_X1    g17411(.A1(new_n17475_), .A2(new_n17383_), .ZN(new_n17476_));
  INV_X1     g17412(.I(new_n17476_), .ZN(new_n17477_));
  OAI22_X1   g17413(.A1(new_n11353_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n11345_), .ZN(new_n17478_));
  NAND2_X1   g17414(.A1(new_n11370_), .A2(new_n4096_), .ZN(new_n17479_));
  AOI21_X1   g17415(.A1(new_n17479_), .A2(new_n17478_), .B(new_n4095_), .ZN(new_n17480_));
  NAND2_X1   g17416(.A1(new_n11379_), .A2(new_n17480_), .ZN(new_n17481_));
  XOR2_X1    g17417(.A1(new_n17481_), .A2(\a[20] ), .Z(new_n17482_));
  INV_X1     g17418(.I(new_n17482_), .ZN(new_n17483_));
  NOR2_X1    g17419(.A1(new_n17477_), .A2(new_n17483_), .ZN(new_n17484_));
  NOR2_X1    g17420(.A1(new_n17476_), .A2(new_n17482_), .ZN(new_n17485_));
  NOR2_X1    g17421(.A1(new_n17484_), .A2(new_n17485_), .ZN(new_n17486_));
  NOR2_X1    g17422(.A1(new_n17486_), .A2(new_n17474_), .ZN(new_n17487_));
  INV_X1     g17423(.I(new_n17474_), .ZN(new_n17488_));
  XOR2_X1    g17424(.A1(new_n17476_), .A2(new_n17483_), .Z(new_n17489_));
  NOR2_X1    g17425(.A1(new_n17489_), .A2(new_n17488_), .ZN(new_n17490_));
  NOR2_X1    g17426(.A1(new_n17487_), .A2(new_n17490_), .ZN(new_n17491_));
  AND3_X2    g17427(.A1(new_n11463_), .A2(new_n4292_), .A3(new_n11567_), .Z(new_n17492_));
  NOR4_X1    g17428(.A1(new_n11468_), .A2(new_n4468_), .A3(new_n11461_), .A4(new_n17492_), .ZN(new_n17493_));
  XOR2_X1    g17429(.A1(new_n17493_), .A2(new_n3372_), .Z(new_n17494_));
  NAND2_X1   g17430(.A1(new_n17491_), .A2(new_n17494_), .ZN(new_n17495_));
  INV_X1     g17431(.I(new_n17494_), .ZN(new_n17496_));
  OAI21_X1   g17432(.A1(new_n17487_), .A2(new_n17490_), .B(new_n17496_), .ZN(new_n17497_));
  AOI21_X1   g17433(.A1(new_n17495_), .A2(new_n17497_), .B(new_n17423_), .ZN(new_n17498_));
  XOR2_X1    g17434(.A1(new_n17491_), .A2(new_n17496_), .Z(new_n17499_));
  NOR2_X1    g17435(.A1(new_n17499_), .A2(new_n17422_), .ZN(new_n17500_));
  NOR2_X1    g17436(.A1(new_n17500_), .A2(new_n17498_), .ZN(new_n17501_));
  INV_X1     g17437(.I(new_n17501_), .ZN(new_n17502_));
  INV_X1     g17438(.I(new_n17406_), .ZN(new_n17503_));
  AOI21_X1   g17439(.A1(new_n17503_), .A2(new_n17410_), .B(new_n17407_), .ZN(new_n17504_));
  INV_X1     g17440(.I(new_n17504_), .ZN(new_n17505_));
  NOR2_X1    g17441(.A1(new_n17505_), .A2(new_n17502_), .ZN(new_n17506_));
  NOR2_X1    g17442(.A1(new_n17504_), .A2(new_n17501_), .ZN(new_n17507_));
  INV_X1     g17443(.I(new_n17507_), .ZN(new_n17508_));
  OAI21_X1   g17444(.A1(new_n17419_), .A2(new_n17506_), .B(new_n17508_), .ZN(new_n17509_));
  INV_X1     g17445(.I(new_n17485_), .ZN(new_n17510_));
  OAI21_X1   g17446(.A1(new_n17474_), .A2(new_n17484_), .B(new_n17510_), .ZN(new_n17511_));
  OAI21_X1   g17447(.A1(new_n17425_), .A2(new_n17468_), .B(new_n17470_), .ZN(new_n17512_));
  OAI22_X1   g17448(.A1(new_n11264_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n11277_), .ZN(new_n17513_));
  NAND2_X1   g17449(.A1(new_n11346_), .A2(new_n3312_), .ZN(new_n17514_));
  AOI21_X1   g17450(.A1(new_n17513_), .A2(new_n17514_), .B(new_n3302_), .ZN(new_n17515_));
  NAND2_X1   g17451(.A1(new_n11757_), .A2(new_n17515_), .ZN(new_n17516_));
  XOR2_X1    g17452(.A1(new_n17516_), .A2(\a[23] ), .Z(new_n17517_));
  INV_X1     g17453(.I(new_n17517_), .ZN(new_n17518_));
  AOI21_X1   g17454(.A1(new_n17430_), .A2(new_n17443_), .B(new_n17444_), .ZN(new_n17519_));
  AOI21_X1   g17455(.A1(new_n11601_), .A2(new_n11602_), .B(new_n11565_), .ZN(new_n17520_));
  XNOR2_X1   g17456(.A1(new_n11591_), .A2(new_n11599_), .ZN(new_n17521_));
  NOR2_X1    g17457(.A1(new_n11566_), .A2(new_n17521_), .ZN(new_n17522_));
  OAI22_X1   g17458(.A1(new_n2747_), .A2(new_n8681_), .B1(new_n8687_), .B2(new_n2742_), .ZN(new_n17523_));
  NAND2_X1   g17459(.A1(new_n8674_), .A2(new_n2750_), .ZN(new_n17524_));
  AOI21_X1   g17460(.A1(new_n17524_), .A2(new_n17523_), .B(new_n2737_), .ZN(new_n17525_));
  NAND2_X1   g17461(.A1(new_n11431_), .A2(new_n17525_), .ZN(new_n17526_));
  XOR2_X1    g17462(.A1(new_n17526_), .A2(\a[29] ), .Z(new_n17527_));
  INV_X1     g17463(.I(new_n17527_), .ZN(new_n17528_));
  NOR3_X1    g17464(.A1(new_n17528_), .A2(new_n17522_), .A3(new_n17520_), .ZN(new_n17529_));
  NOR2_X1    g17465(.A1(new_n17522_), .A2(new_n17520_), .ZN(new_n17530_));
  NOR2_X1    g17466(.A1(new_n17530_), .A2(new_n17527_), .ZN(new_n17531_));
  NOR2_X1    g17467(.A1(new_n17531_), .A2(new_n17529_), .ZN(new_n17532_));
  NOR2_X1    g17468(.A1(new_n17532_), .A2(new_n17519_), .ZN(new_n17533_));
  INV_X1     g17469(.I(new_n17519_), .ZN(new_n17534_));
  XOR2_X1    g17470(.A1(new_n17530_), .A2(new_n17528_), .Z(new_n17535_));
  NOR2_X1    g17471(.A1(new_n17535_), .A2(new_n17534_), .ZN(new_n17536_));
  NOR2_X1    g17472(.A1(new_n17536_), .A2(new_n17533_), .ZN(new_n17537_));
  NOR2_X1    g17473(.A1(new_n17459_), .A2(new_n17448_), .ZN(new_n17538_));
  NOR2_X1    g17474(.A1(new_n17538_), .A2(new_n17458_), .ZN(new_n17539_));
  OAI22_X1   g17475(.A1(new_n11284_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n8661_), .ZN(new_n17540_));
  NAND2_X1   g17476(.A1(new_n11272_), .A2(new_n3317_), .ZN(new_n17541_));
  AOI21_X1   g17477(.A1(new_n17540_), .A2(new_n17541_), .B(new_n3260_), .ZN(new_n17542_));
  NAND2_X1   g17478(.A1(new_n11655_), .A2(new_n17542_), .ZN(new_n17543_));
  XOR2_X1    g17479(.A1(new_n17543_), .A2(\a[26] ), .Z(new_n17544_));
  INV_X1     g17480(.I(new_n17544_), .ZN(new_n17545_));
  XOR2_X1    g17481(.A1(new_n17539_), .A2(new_n17545_), .Z(new_n17546_));
  NOR2_X1    g17482(.A1(new_n17546_), .A2(new_n17537_), .ZN(new_n17547_));
  INV_X1     g17483(.I(new_n17537_), .ZN(new_n17548_));
  NOR3_X1    g17484(.A1(new_n17538_), .A2(new_n17458_), .A3(new_n17545_), .ZN(new_n17549_));
  NOR2_X1    g17485(.A1(new_n17539_), .A2(new_n17544_), .ZN(new_n17550_));
  NOR2_X1    g17486(.A1(new_n17550_), .A2(new_n17549_), .ZN(new_n17551_));
  NOR2_X1    g17487(.A1(new_n17551_), .A2(new_n17548_), .ZN(new_n17552_));
  NOR2_X1    g17488(.A1(new_n17547_), .A2(new_n17552_), .ZN(new_n17553_));
  XOR2_X1    g17489(.A1(new_n17553_), .A2(new_n17518_), .Z(new_n17554_));
  XOR2_X1    g17490(.A1(new_n17554_), .A2(new_n17512_), .Z(new_n17555_));
  OAI22_X1   g17491(.A1(new_n11353_), .A2(new_n3769_), .B1(new_n4097_), .B2(new_n11697_), .ZN(new_n17556_));
  NAND2_X1   g17492(.A1(new_n11370_), .A2(new_n3776_), .ZN(new_n17557_));
  AOI21_X1   g17493(.A1(new_n17557_), .A2(new_n17556_), .B(new_n4095_), .ZN(new_n17558_));
  NAND2_X1   g17494(.A1(new_n11700_), .A2(new_n17558_), .ZN(new_n17559_));
  XOR2_X1    g17495(.A1(new_n17559_), .A2(\a[20] ), .Z(new_n17560_));
  XOR2_X1    g17496(.A1(new_n17555_), .A2(new_n17560_), .Z(new_n17561_));
  INV_X1     g17497(.I(new_n17561_), .ZN(new_n17562_));
  INV_X1     g17498(.I(new_n17560_), .ZN(new_n17563_));
  OR2_X2     g17499(.A1(new_n17555_), .A2(new_n17563_), .Z(new_n17564_));
  NAND2_X1   g17500(.A1(new_n17555_), .A2(new_n17563_), .ZN(new_n17565_));
  AOI21_X1   g17501(.A1(new_n17564_), .A2(new_n17565_), .B(new_n17511_), .ZN(new_n17566_));
  AOI21_X1   g17502(.A1(new_n17562_), .A2(new_n17511_), .B(new_n17566_), .ZN(new_n17567_));
  NAND2_X1   g17503(.A1(new_n17495_), .A2(new_n17422_), .ZN(new_n17568_));
  NAND2_X1   g17504(.A1(new_n17568_), .A2(new_n17497_), .ZN(new_n17569_));
  NOR2_X1    g17505(.A1(new_n17569_), .A2(new_n17567_), .ZN(new_n17570_));
  INV_X1     g17506(.I(new_n17570_), .ZN(new_n17571_));
  NAND2_X1   g17507(.A1(new_n17569_), .A2(new_n17567_), .ZN(new_n17572_));
  INV_X1     g17508(.I(new_n17572_), .ZN(new_n17573_));
  AOI21_X1   g17509(.A1(new_n17509_), .A2(new_n17571_), .B(new_n17573_), .ZN(new_n17574_));
  INV_X1     g17510(.I(new_n17529_), .ZN(new_n17575_));
  AOI21_X1   g17511(.A1(new_n17575_), .A2(new_n17534_), .B(new_n17531_), .ZN(new_n17576_));
  INV_X1     g17512(.I(new_n17576_), .ZN(new_n17577_));
  XOR2_X1    g17513(.A1(new_n11629_), .A2(new_n11623_), .Z(new_n17578_));
  OAI21_X1   g17514(.A1(new_n11631_), .A2(new_n11634_), .B(new_n11604_), .ZN(new_n17579_));
  OAI21_X1   g17515(.A1(new_n11604_), .A2(new_n17578_), .B(new_n17579_), .ZN(new_n17580_));
  OAI22_X1   g17516(.A1(new_n11284_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n11271_), .ZN(new_n17581_));
  NAND2_X1   g17517(.A1(new_n11311_), .A2(new_n3317_), .ZN(new_n17582_));
  AOI21_X1   g17518(.A1(new_n17581_), .A2(new_n17582_), .B(new_n3260_), .ZN(new_n17583_));
  NAND2_X1   g17519(.A1(new_n11391_), .A2(new_n17583_), .ZN(new_n17584_));
  XOR2_X1    g17520(.A1(new_n17584_), .A2(\a[26] ), .Z(new_n17585_));
  AND2_X2    g17521(.A1(new_n17580_), .A2(new_n17585_), .Z(new_n17586_));
  NOR2_X1    g17522(.A1(new_n17580_), .A2(new_n17585_), .ZN(new_n17587_));
  OAI21_X1   g17523(.A1(new_n17586_), .A2(new_n17587_), .B(new_n17577_), .ZN(new_n17588_));
  XNOR2_X1   g17524(.A1(new_n17580_), .A2(new_n17585_), .ZN(new_n17589_));
  OAI21_X1   g17525(.A1(new_n17577_), .A2(new_n17589_), .B(new_n17588_), .ZN(new_n17590_));
  INV_X1     g17526(.I(new_n17549_), .ZN(new_n17591_));
  AOI21_X1   g17527(.A1(new_n17591_), .A2(new_n17548_), .B(new_n17550_), .ZN(new_n17592_));
  INV_X1     g17528(.I(new_n17592_), .ZN(new_n17593_));
  OAI22_X1   g17529(.A1(new_n11264_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n11345_), .ZN(new_n17594_));
  NAND2_X1   g17530(.A1(new_n11354_), .A2(new_n3312_), .ZN(new_n17595_));
  AOI21_X1   g17531(.A1(new_n17595_), .A2(new_n17594_), .B(new_n3302_), .ZN(new_n17596_));
  NAND2_X1   g17532(.A1(new_n11678_), .A2(new_n17596_), .ZN(new_n17597_));
  XOR2_X1    g17533(.A1(new_n17597_), .A2(\a[23] ), .Z(new_n17598_));
  INV_X1     g17534(.I(new_n17598_), .ZN(new_n17599_));
  NOR2_X1    g17535(.A1(new_n17599_), .A2(new_n17593_), .ZN(new_n17600_));
  NOR2_X1    g17536(.A1(new_n17598_), .A2(new_n17592_), .ZN(new_n17601_));
  OAI21_X1   g17537(.A1(new_n17600_), .A2(new_n17601_), .B(new_n17590_), .ZN(new_n17602_));
  XOR2_X1    g17538(.A1(new_n17598_), .A2(new_n17593_), .Z(new_n17603_));
  OAI21_X1   g17539(.A1(new_n17590_), .A2(new_n17603_), .B(new_n17602_), .ZN(new_n17604_));
  OAI22_X1   g17540(.A1(new_n11369_), .A2(new_n3769_), .B1(new_n4097_), .B2(new_n11461_), .ZN(new_n17605_));
  NAND2_X1   g17541(.A1(new_n11694_), .A2(new_n3776_), .ZN(new_n17606_));
  AOI21_X1   g17542(.A1(new_n17605_), .A2(new_n17606_), .B(new_n4095_), .ZN(new_n17607_));
  NAND2_X1   g17543(.A1(new_n12720_), .A2(new_n17607_), .ZN(new_n17608_));
  XOR2_X1    g17544(.A1(new_n17608_), .A2(\a[20] ), .Z(new_n17609_));
  INV_X1     g17545(.I(new_n17512_), .ZN(new_n17610_));
  NOR2_X1    g17546(.A1(new_n17553_), .A2(new_n17518_), .ZN(new_n17611_));
  AOI21_X1   g17547(.A1(new_n17554_), .A2(new_n17610_), .B(new_n17611_), .ZN(new_n17612_));
  XNOR2_X1   g17548(.A1(new_n17612_), .A2(new_n17609_), .ZN(new_n17613_));
  XOR2_X1    g17549(.A1(new_n17613_), .A2(new_n17604_), .Z(new_n17614_));
  XOR2_X1    g17550(.A1(new_n17604_), .A2(new_n17609_), .Z(new_n17615_));
  INV_X1     g17551(.I(new_n17615_), .ZN(new_n17616_));
  OAI21_X1   g17552(.A1(new_n17609_), .A2(new_n17612_), .B(new_n17616_), .ZN(new_n17617_));
  XOR2_X1    g17553(.A1(new_n11644_), .A2(new_n11637_), .Z(new_n17618_));
  OAI21_X1   g17554(.A1(new_n11642_), .A2(new_n11645_), .B(new_n11635_), .ZN(new_n17619_));
  OAI21_X1   g17555(.A1(new_n11635_), .A2(new_n17618_), .B(new_n17619_), .ZN(new_n17620_));
  AOI22_X1   g17556(.A1(new_n11311_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n11272_), .ZN(new_n17621_));
  NOR2_X1    g17557(.A1(new_n11264_), .A2(new_n3318_), .ZN(new_n17622_));
  OAI21_X1   g17558(.A1(new_n17622_), .A2(new_n17621_), .B(new_n3259_), .ZN(new_n17623_));
  NOR2_X1    g17559(.A1(new_n11310_), .A2(new_n17623_), .ZN(new_n17624_));
  XOR2_X1    g17560(.A1(new_n17624_), .A2(new_n72_), .Z(new_n17625_));
  OAI22_X1   g17561(.A1(new_n8661_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n8673_), .ZN(new_n17626_));
  NAND2_X1   g17562(.A1(new_n11285_), .A2(new_n2750_), .ZN(new_n17627_));
  AOI21_X1   g17563(.A1(new_n17627_), .A2(new_n17626_), .B(new_n2737_), .ZN(new_n17628_));
  NAND2_X1   g17564(.A1(new_n11323_), .A2(new_n17628_), .ZN(new_n17629_));
  XOR2_X1    g17565(.A1(new_n17629_), .A2(\a[29] ), .Z(new_n17630_));
  XNOR2_X1   g17566(.A1(new_n17625_), .A2(new_n17630_), .ZN(new_n17631_));
  NOR2_X1    g17567(.A1(new_n17625_), .A2(new_n17630_), .ZN(new_n17632_));
  NAND2_X1   g17568(.A1(new_n17625_), .A2(new_n17630_), .ZN(new_n17633_));
  INV_X1     g17569(.I(new_n17633_), .ZN(new_n17634_));
  NOR2_X1    g17570(.A1(new_n17634_), .A2(new_n17632_), .ZN(new_n17635_));
  MUX2_X1    g17571(.I0(new_n17635_), .I1(new_n17631_), .S(new_n17620_), .Z(new_n17636_));
  NOR2_X1    g17572(.A1(new_n17586_), .A2(new_n17576_), .ZN(new_n17637_));
  NOR2_X1    g17573(.A1(new_n17637_), .A2(new_n17587_), .ZN(new_n17638_));
  OAI22_X1   g17574(.A1(new_n11353_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n11345_), .ZN(new_n17639_));
  NAND2_X1   g17575(.A1(new_n11370_), .A2(new_n3312_), .ZN(new_n17640_));
  AOI21_X1   g17576(.A1(new_n17640_), .A2(new_n17639_), .B(new_n3302_), .ZN(new_n17641_));
  NAND2_X1   g17577(.A1(new_n11379_), .A2(new_n17641_), .ZN(new_n17642_));
  XOR2_X1    g17578(.A1(new_n17642_), .A2(\a[23] ), .Z(new_n17643_));
  AND2_X2    g17579(.A1(new_n17638_), .A2(new_n17643_), .Z(new_n17644_));
  NOR2_X1    g17580(.A1(new_n17638_), .A2(new_n17643_), .ZN(new_n17645_));
  NOR2_X1    g17581(.A1(new_n17644_), .A2(new_n17645_), .ZN(new_n17646_));
  NOR2_X1    g17582(.A1(new_n17646_), .A2(new_n17636_), .ZN(new_n17647_));
  XNOR2_X1   g17583(.A1(new_n17638_), .A2(new_n17643_), .ZN(new_n17648_));
  INV_X1     g17584(.I(new_n17648_), .ZN(new_n17649_));
  AOI21_X1   g17585(.A1(new_n17636_), .A2(new_n17649_), .B(new_n17647_), .ZN(new_n17650_));
  INV_X1     g17586(.I(new_n17600_), .ZN(new_n17651_));
  AOI21_X1   g17587(.A1(new_n17651_), .A2(new_n17590_), .B(new_n17601_), .ZN(new_n17652_));
  AND3_X2    g17588(.A1(new_n11463_), .A2(new_n3770_), .A3(new_n11227_), .Z(new_n17653_));
  NOR4_X1    g17589(.A1(new_n11468_), .A2(new_n4095_), .A3(new_n11461_), .A4(new_n17653_), .ZN(new_n17654_));
  XOR2_X1    g17590(.A1(new_n17654_), .A2(new_n3035_), .Z(new_n17655_));
  AND2_X2    g17591(.A1(new_n17652_), .A2(new_n17655_), .Z(new_n17656_));
  NOR2_X1    g17592(.A1(new_n17652_), .A2(new_n17655_), .ZN(new_n17657_));
  NOR2_X1    g17593(.A1(new_n17656_), .A2(new_n17657_), .ZN(new_n17658_));
  NOR2_X1    g17594(.A1(new_n17658_), .A2(new_n17650_), .ZN(new_n17659_));
  INV_X1     g17595(.I(new_n17650_), .ZN(new_n17660_));
  XNOR2_X1   g17596(.A1(new_n17652_), .A2(new_n17655_), .ZN(new_n17661_));
  NOR2_X1    g17597(.A1(new_n17661_), .A2(new_n17660_), .ZN(new_n17662_));
  NOR2_X1    g17598(.A1(new_n17659_), .A2(new_n17662_), .ZN(new_n17663_));
  XNOR2_X1   g17599(.A1(new_n17617_), .A2(new_n17663_), .ZN(new_n17664_));
  INV_X1     g17600(.I(new_n17664_), .ZN(new_n17665_));
  NAND2_X1   g17601(.A1(new_n17564_), .A2(new_n17511_), .ZN(new_n17666_));
  NAND2_X1   g17602(.A1(new_n17666_), .A2(new_n17565_), .ZN(new_n17667_));
  INV_X1     g17603(.I(new_n17667_), .ZN(new_n17668_));
  NOR2_X1    g17604(.A1(new_n17665_), .A2(new_n17668_), .ZN(new_n17669_));
  NOR3_X1    g17605(.A1(new_n17574_), .A2(new_n17614_), .A3(new_n17669_), .ZN(new_n17670_));
  NAND2_X1   g17606(.A1(new_n17617_), .A2(new_n17663_), .ZN(new_n17671_));
  INV_X1     g17607(.I(new_n17671_), .ZN(new_n17672_));
  INV_X1     g17608(.I(new_n17645_), .ZN(new_n17673_));
  OAI21_X1   g17609(.A1(new_n17636_), .A2(new_n17644_), .B(new_n17673_), .ZN(new_n17674_));
  NOR2_X1    g17610(.A1(new_n11662_), .A2(new_n11665_), .ZN(new_n17675_));
  NOR2_X1    g17611(.A1(new_n17675_), .A2(new_n11646_), .ZN(new_n17676_));
  XOR2_X1    g17612(.A1(new_n11660_), .A2(new_n11650_), .Z(new_n17677_));
  NOR2_X1    g17613(.A1(new_n11647_), .A2(new_n17677_), .ZN(new_n17678_));
  NOR2_X1    g17614(.A1(new_n17678_), .A2(new_n17676_), .ZN(new_n17679_));
  NOR2_X1    g17615(.A1(new_n17634_), .A2(new_n17620_), .ZN(new_n17680_));
  NOR2_X1    g17616(.A1(new_n17680_), .A2(new_n17632_), .ZN(new_n17681_));
  OAI22_X1   g17617(.A1(new_n11264_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n11277_), .ZN(new_n17682_));
  NAND2_X1   g17618(.A1(new_n11346_), .A2(new_n3317_), .ZN(new_n17683_));
  AOI21_X1   g17619(.A1(new_n17682_), .A2(new_n17683_), .B(new_n3260_), .ZN(new_n17684_));
  NAND2_X1   g17620(.A1(new_n11757_), .A2(new_n17684_), .ZN(new_n17685_));
  XOR2_X1    g17621(.A1(new_n17685_), .A2(\a[26] ), .Z(new_n17686_));
  INV_X1     g17622(.I(new_n17686_), .ZN(new_n17687_));
  XOR2_X1    g17623(.A1(new_n17681_), .A2(new_n17687_), .Z(new_n17688_));
  NOR3_X1    g17624(.A1(new_n17680_), .A2(new_n17632_), .A3(new_n17687_), .ZN(new_n17689_));
  NOR2_X1    g17625(.A1(new_n17681_), .A2(new_n17686_), .ZN(new_n17690_));
  OAI21_X1   g17626(.A1(new_n17690_), .A2(new_n17689_), .B(new_n17679_), .ZN(new_n17691_));
  OAI21_X1   g17627(.A1(new_n17688_), .A2(new_n17679_), .B(new_n17691_), .ZN(new_n17692_));
  OAI22_X1   g17628(.A1(new_n11353_), .A2(new_n3310_), .B1(new_n3780_), .B2(new_n11697_), .ZN(new_n17693_));
  NAND2_X1   g17629(.A1(new_n11370_), .A2(new_n3782_), .ZN(new_n17694_));
  AOI21_X1   g17630(.A1(new_n17694_), .A2(new_n17693_), .B(new_n3302_), .ZN(new_n17695_));
  NAND2_X1   g17631(.A1(new_n11700_), .A2(new_n17695_), .ZN(new_n17696_));
  XOR2_X1    g17632(.A1(new_n17696_), .A2(\a[23] ), .Z(new_n17697_));
  XOR2_X1    g17633(.A1(new_n17692_), .A2(new_n17697_), .Z(new_n17698_));
  AND2_X2    g17634(.A1(new_n17698_), .A2(new_n17674_), .Z(new_n17699_));
  NAND2_X1   g17635(.A1(new_n17692_), .A2(new_n17697_), .ZN(new_n17700_));
  OR2_X2     g17636(.A1(new_n17692_), .A2(new_n17697_), .Z(new_n17701_));
  AOI21_X1   g17637(.A1(new_n17701_), .A2(new_n17700_), .B(new_n17674_), .ZN(new_n17702_));
  NOR2_X1    g17638(.A1(new_n17699_), .A2(new_n17702_), .ZN(new_n17703_));
  NOR3_X1    g17639(.A1(new_n17670_), .A2(new_n17672_), .A3(new_n17703_), .ZN(new_n17704_));
  INV_X1     g17640(.I(new_n17704_), .ZN(new_n17705_));
  NOR2_X1    g17641(.A1(new_n17245_), .A2(new_n17236_), .ZN(new_n17706_));
  AOI21_X1   g17642(.A1(new_n17235_), .A2(new_n17237_), .B(new_n17333_), .ZN(new_n17707_));
  NOR3_X1    g17643(.A1(new_n17245_), .A2(new_n17236_), .A3(new_n17331_), .ZN(new_n17708_));
  OAI22_X1   g17644(.A1(new_n17708_), .A2(new_n17707_), .B1(new_n17706_), .B2(new_n17336_), .ZN(new_n17709_));
  INV_X1     g17645(.I(new_n17418_), .ZN(new_n17710_));
  OAI21_X1   g17646(.A1(new_n17709_), .A2(new_n17415_), .B(new_n17710_), .ZN(new_n17711_));
  INV_X1     g17647(.I(new_n17506_), .ZN(new_n17712_));
  AOI21_X1   g17648(.A1(new_n17711_), .A2(new_n17712_), .B(new_n17507_), .ZN(new_n17713_));
  OAI21_X1   g17649(.A1(new_n17713_), .A2(new_n17570_), .B(new_n17572_), .ZN(new_n17714_));
  INV_X1     g17650(.I(new_n17614_), .ZN(new_n17715_));
  INV_X1     g17651(.I(new_n17669_), .ZN(new_n17716_));
  NAND3_X1   g17652(.A1(new_n17714_), .A2(new_n17715_), .A3(new_n17716_), .ZN(new_n17717_));
  INV_X1     g17653(.I(new_n17703_), .ZN(new_n17718_));
  AOI21_X1   g17654(.A1(new_n17717_), .A2(new_n17671_), .B(new_n17718_), .ZN(new_n17719_));
  NOR3_X1    g17655(.A1(new_n17670_), .A2(new_n17672_), .A3(new_n17703_), .ZN(new_n17720_));
  INV_X1     g17656(.I(new_n17656_), .ZN(new_n17721_));
  AOI21_X1   g17657(.A1(new_n17721_), .A2(new_n17660_), .B(new_n17657_), .ZN(new_n17722_));
  OAI21_X1   g17658(.A1(new_n17720_), .A2(new_n17719_), .B(new_n17722_), .ZN(new_n17723_));
  NAND2_X1   g17659(.A1(new_n17723_), .A2(new_n17705_), .ZN(new_n17724_));
  INV_X1     g17660(.I(new_n11685_), .ZN(new_n17725_));
  NAND2_X1   g17661(.A1(new_n17725_), .A2(new_n11684_), .ZN(new_n17726_));
  NAND2_X1   g17662(.A1(new_n17726_), .A2(new_n11667_), .ZN(new_n17727_));
  XOR2_X1    g17663(.A1(new_n11671_), .A2(new_n11683_), .Z(new_n17728_));
  NAND2_X1   g17664(.A1(new_n17728_), .A2(new_n11666_), .ZN(new_n17729_));
  NAND2_X1   g17665(.A1(new_n17727_), .A2(new_n17729_), .ZN(new_n17730_));
  INV_X1     g17666(.I(new_n17730_), .ZN(new_n17731_));
  INV_X1     g17667(.I(new_n17690_), .ZN(new_n17732_));
  OAI21_X1   g17668(.A1(new_n17679_), .A2(new_n17689_), .B(new_n17732_), .ZN(new_n17733_));
  OAI22_X1   g17669(.A1(new_n11369_), .A2(new_n3310_), .B1(new_n3780_), .B2(new_n11461_), .ZN(new_n17734_));
  NAND2_X1   g17670(.A1(new_n11694_), .A2(new_n3782_), .ZN(new_n17735_));
  AOI21_X1   g17671(.A1(new_n17734_), .A2(new_n17735_), .B(new_n3302_), .ZN(new_n17736_));
  NAND2_X1   g17672(.A1(new_n12720_), .A2(new_n17736_), .ZN(new_n17737_));
  XOR2_X1    g17673(.A1(new_n17737_), .A2(\a[23] ), .Z(new_n17738_));
  INV_X1     g17674(.I(new_n17738_), .ZN(new_n17739_));
  NOR2_X1    g17675(.A1(new_n17733_), .A2(new_n17739_), .ZN(new_n17740_));
  INV_X1     g17676(.I(new_n17740_), .ZN(new_n17741_));
  NAND2_X1   g17677(.A1(new_n17733_), .A2(new_n17739_), .ZN(new_n17742_));
  AOI21_X1   g17678(.A1(new_n17741_), .A2(new_n17742_), .B(new_n17731_), .ZN(new_n17743_));
  XOR2_X1    g17679(.A1(new_n17733_), .A2(new_n17738_), .Z(new_n17744_));
  NOR2_X1    g17680(.A1(new_n17744_), .A2(new_n17730_), .ZN(new_n17745_));
  NOR2_X1    g17681(.A1(new_n17745_), .A2(new_n17743_), .ZN(new_n17746_));
  INV_X1     g17682(.I(new_n17746_), .ZN(new_n17747_));
  INV_X1     g17683(.I(new_n11473_), .ZN(new_n17748_));
  AOI21_X1   g17684(.A1(new_n17748_), .A2(new_n11688_), .B(new_n11686_), .ZN(new_n17749_));
  XNOR2_X1   g17685(.A1(new_n11459_), .A2(new_n11472_), .ZN(new_n17750_));
  NOR2_X1    g17686(.A1(new_n17750_), .A2(new_n11687_), .ZN(new_n17751_));
  NOR2_X1    g17687(.A1(new_n17751_), .A2(new_n17749_), .ZN(new_n17752_));
  OAI21_X1   g17688(.A1(new_n17731_), .A2(new_n17740_), .B(new_n17742_), .ZN(new_n17753_));
  XOR2_X1    g17689(.A1(new_n17752_), .A2(new_n17753_), .Z(new_n17754_));
  NAND2_X1   g17690(.A1(new_n17700_), .A2(new_n17674_), .ZN(new_n17755_));
  NAND2_X1   g17691(.A1(new_n17755_), .A2(new_n17701_), .ZN(new_n17756_));
  NAND2_X1   g17692(.A1(new_n17754_), .A2(new_n17756_), .ZN(new_n17757_));
  NAND3_X1   g17693(.A1(new_n17724_), .A2(new_n17747_), .A3(new_n17757_), .ZN(new_n17758_));
  INV_X1     g17694(.I(new_n17753_), .ZN(new_n17759_));
  NAND2_X1   g17695(.A1(new_n17752_), .A2(new_n17759_), .ZN(new_n17760_));
  AOI21_X1   g17696(.A1(new_n17758_), .A2(new_n17760_), .B(new_n11777_), .ZN(new_n17761_));
  NAND3_X1   g17697(.A1(new_n17758_), .A2(new_n11777_), .A3(new_n17760_), .ZN(new_n17762_));
  INV_X1     g17698(.I(new_n17762_), .ZN(new_n17763_));
  OAI21_X1   g17699(.A1(new_n17763_), .A2(new_n17761_), .B(new_n11689_), .ZN(new_n17764_));
  INV_X1     g17700(.I(new_n11689_), .ZN(new_n17765_));
  INV_X1     g17701(.I(new_n11777_), .ZN(new_n17766_));
  NAND2_X1   g17702(.A1(new_n17758_), .A2(new_n17760_), .ZN(new_n17767_));
  NAND2_X1   g17703(.A1(new_n17767_), .A2(new_n17766_), .ZN(new_n17768_));
  NAND3_X1   g17704(.A1(new_n17768_), .A2(new_n17765_), .A3(new_n17762_), .ZN(new_n17769_));
  NAND2_X1   g17705(.A1(new_n17764_), .A2(new_n17769_), .ZN(new_n17770_));
  INV_X1     g17706(.I(new_n17756_), .ZN(new_n17771_));
  XOR2_X1    g17707(.A1(new_n17746_), .A2(new_n17771_), .Z(new_n17772_));
  XOR2_X1    g17708(.A1(new_n17746_), .A2(new_n17771_), .Z(new_n17773_));
  NOR2_X1    g17709(.A1(new_n17724_), .A2(new_n17773_), .ZN(new_n17774_));
  AOI21_X1   g17710(.A1(new_n17724_), .A2(new_n17772_), .B(new_n17774_), .ZN(new_n17775_));
  OAI21_X1   g17711(.A1(new_n17670_), .A2(new_n17672_), .B(new_n17703_), .ZN(new_n17776_));
  NAND3_X1   g17712(.A1(new_n17717_), .A2(new_n17671_), .A3(new_n17718_), .ZN(new_n17777_));
  INV_X1     g17713(.I(new_n17722_), .ZN(new_n17778_));
  NAND3_X1   g17714(.A1(new_n17776_), .A2(new_n17777_), .A3(new_n17778_), .ZN(new_n17779_));
  NAND2_X1   g17715(.A1(new_n17723_), .A2(new_n17779_), .ZN(new_n17780_));
  XNOR2_X1   g17716(.A1(new_n17569_), .A2(new_n17567_), .ZN(new_n17781_));
  NOR2_X1    g17717(.A1(new_n17713_), .A2(new_n17781_), .ZN(new_n17782_));
  AOI21_X1   g17718(.A1(new_n17571_), .A2(new_n17572_), .B(new_n17509_), .ZN(new_n17783_));
  NOR2_X1    g17719(.A1(new_n17783_), .A2(new_n17782_), .ZN(new_n17784_));
  AOI21_X1   g17720(.A1(new_n17332_), .A2(new_n17334_), .B(new_n17337_), .ZN(new_n17785_));
  NOR3_X1    g17721(.A1(new_n17708_), .A2(new_n17707_), .A3(new_n17336_), .ZN(new_n17786_));
  NOR2_X1    g17722(.A1(new_n17786_), .A2(new_n17785_), .ZN(new_n17787_));
  NAND2_X1   g17723(.A1(new_n17240_), .A2(new_n17241_), .ZN(new_n17788_));
  XOR2_X1    g17724(.A1(new_n17788_), .A2(new_n17229_), .Z(new_n17789_));
  INV_X1     g17725(.I(new_n17789_), .ZN(new_n17790_));
  INV_X1     g17726(.I(new_n17199_), .ZN(new_n17791_));
  NOR3_X1    g17727(.A1(new_n17193_), .A2(new_n17180_), .A3(new_n17198_), .ZN(new_n17792_));
  NOR2_X1    g17728(.A1(new_n17791_), .A2(new_n17792_), .ZN(new_n17793_));
  INV_X1     g17729(.I(new_n17793_), .ZN(new_n17794_));
  AOI21_X1   g17730(.A1(new_n17062_), .A2(new_n17026_), .B(new_n17066_), .ZN(new_n17795_));
  NOR3_X1    g17731(.A1(new_n17182_), .A2(new_n17181_), .A3(new_n17065_), .ZN(new_n17796_));
  NOR2_X1    g17732(.A1(new_n17796_), .A2(new_n17795_), .ZN(new_n17797_));
  INV_X1     g17733(.I(new_n17797_), .ZN(new_n17798_));
  NOR2_X1    g17734(.A1(new_n17051_), .A2(new_n16847_), .ZN(new_n17799_));
  NOR2_X1    g17735(.A1(new_n16947_), .A2(new_n17044_), .ZN(new_n17800_));
  NOR2_X1    g17736(.A1(new_n17799_), .A2(new_n17800_), .ZN(new_n17801_));
  INV_X1     g17737(.I(new_n17801_), .ZN(new_n17802_));
  INV_X1     g17738(.I(new_n16726_), .ZN(new_n17803_));
  NOR2_X1    g17739(.A1(new_n16734_), .A2(new_n17803_), .ZN(new_n17804_));
  AOI21_X1   g17740(.A1(new_n16730_), .A2(new_n16733_), .B(new_n16726_), .ZN(new_n17805_));
  NOR2_X1    g17741(.A1(new_n17804_), .A2(new_n17805_), .ZN(new_n17806_));
  INV_X1     g17742(.I(new_n17806_), .ZN(new_n17807_));
  NOR2_X1    g17743(.A1(new_n16046_), .A2(new_n16047_), .ZN(new_n17808_));
  XOR2_X1    g17744(.A1(new_n16707_), .A2(new_n16045_), .Z(new_n17809_));
  XOR2_X1    g17745(.A1(new_n17809_), .A2(new_n17808_), .Z(new_n17810_));
  OAI22_X1   g17746(.A1(new_n11353_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n11345_), .ZN(new_n17811_));
  NAND2_X1   g17747(.A1(new_n11370_), .A2(new_n9488_), .ZN(new_n17812_));
  AOI21_X1   g17748(.A1(new_n17812_), .A2(new_n17811_), .B(new_n9482_), .ZN(new_n17813_));
  NAND2_X1   g17749(.A1(new_n11379_), .A2(new_n17813_), .ZN(new_n17814_));
  XOR2_X1    g17750(.A1(new_n17814_), .A2(\a[2] ), .Z(new_n17815_));
  XOR2_X1    g17751(.A1(new_n17810_), .A2(new_n17815_), .Z(new_n17816_));
  OAI22_X1   g17752(.A1(new_n11264_), .A2(new_n9485_), .B1(new_n9483_), .B2(new_n11345_), .ZN(new_n17817_));
  NAND2_X1   g17753(.A1(new_n11354_), .A2(new_n9488_), .ZN(new_n17818_));
  AOI21_X1   g17754(.A1(new_n17818_), .A2(new_n17817_), .B(new_n9482_), .ZN(new_n17819_));
  NAND2_X1   g17755(.A1(new_n11678_), .A2(new_n17819_), .ZN(new_n17820_));
  XOR2_X1    g17756(.A1(new_n17820_), .A2(\a[2] ), .Z(new_n17821_));
  XOR2_X1    g17757(.A1(new_n16635_), .A2(new_n16679_), .Z(new_n17822_));
  INV_X1     g17758(.I(new_n17822_), .ZN(new_n17823_));
  NOR2_X1    g17759(.A1(new_n17823_), .A2(new_n17821_), .ZN(new_n17824_));
  AND2_X2    g17760(.A1(new_n17816_), .A2(new_n17824_), .Z(new_n17825_));
  NOR2_X1    g17761(.A1(new_n17816_), .A2(new_n17824_), .ZN(new_n17826_));
  OR2_X2     g17762(.A1(new_n17825_), .A2(new_n17826_), .Z(new_n17827_));
  INV_X1     g17763(.I(new_n17827_), .ZN(new_n17828_));
  NAND2_X1   g17764(.A1(new_n16136_), .A2(new_n16147_), .ZN(new_n17829_));
  NAND2_X1   g17765(.A1(new_n16701_), .A2(new_n16632_), .ZN(new_n17830_));
  XOR2_X1    g17766(.A1(new_n17830_), .A2(new_n16627_), .Z(new_n17831_));
  XOR2_X1    g17767(.A1(new_n17831_), .A2(new_n17829_), .Z(new_n17832_));
  AOI22_X1   g17768(.A1(new_n11311_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n11272_), .ZN(new_n17833_));
  NOR2_X1    g17769(.A1(new_n11264_), .A2(new_n9489_), .ZN(new_n17834_));
  OAI21_X1   g17770(.A1(new_n17834_), .A2(new_n17833_), .B(new_n6922_), .ZN(new_n17835_));
  NOR2_X1    g17771(.A1(new_n11310_), .A2(new_n17835_), .ZN(new_n17836_));
  XOR2_X1    g17772(.A1(new_n17836_), .A2(new_n4387_), .Z(new_n17837_));
  XOR2_X1    g17773(.A1(new_n17832_), .A2(new_n17837_), .Z(new_n17838_));
  OAI22_X1   g17774(.A1(new_n11284_), .A2(new_n9485_), .B1(new_n9483_), .B2(new_n11271_), .ZN(new_n17839_));
  NAND2_X1   g17775(.A1(new_n11311_), .A2(new_n9488_), .ZN(new_n17840_));
  AOI21_X1   g17776(.A1(new_n17839_), .A2(new_n17840_), .B(new_n9482_), .ZN(new_n17841_));
  NAND2_X1   g17777(.A1(new_n11391_), .A2(new_n17841_), .ZN(new_n17842_));
  XOR2_X1    g17778(.A1(new_n17842_), .A2(\a[2] ), .Z(new_n17843_));
  XOR2_X1    g17779(.A1(new_n16700_), .A2(new_n16168_), .Z(new_n17844_));
  INV_X1     g17780(.I(new_n17844_), .ZN(new_n17845_));
  NOR2_X1    g17781(.A1(new_n17845_), .A2(new_n17843_), .ZN(new_n17846_));
  AND2_X2    g17782(.A1(new_n17838_), .A2(new_n17846_), .Z(new_n17847_));
  NOR2_X1    g17783(.A1(new_n17838_), .A2(new_n17846_), .ZN(new_n17848_));
  NOR2_X1    g17784(.A1(new_n17847_), .A2(new_n17848_), .ZN(new_n17849_));
  INV_X1     g17785(.I(new_n17849_), .ZN(new_n17850_));
  XOR2_X1    g17786(.A1(new_n16699_), .A2(new_n16183_), .Z(new_n17851_));
  INV_X1     g17787(.I(new_n17851_), .ZN(new_n17852_));
  OAI22_X1   g17788(.A1(new_n8673_), .A2(new_n9483_), .B1(new_n8687_), .B2(new_n9485_), .ZN(new_n17853_));
  NAND2_X1   g17789(.A1(new_n8662_), .A2(new_n9488_), .ZN(new_n17854_));
  AOI21_X1   g17790(.A1(new_n17854_), .A2(new_n17853_), .B(new_n9482_), .ZN(new_n17855_));
  NAND2_X1   g17791(.A1(new_n11624_), .A2(new_n17855_), .ZN(new_n17856_));
  XOR2_X1    g17792(.A1(new_n17856_), .A2(\a[2] ), .Z(new_n17857_));
  INV_X1     g17793(.I(new_n17857_), .ZN(new_n17858_));
  AOI21_X1   g17794(.A1(new_n16694_), .A2(new_n16609_), .B(new_n16685_), .ZN(new_n17859_));
  NOR2_X1    g17795(.A1(new_n16613_), .A2(new_n17859_), .ZN(new_n17860_));
  NOR2_X1    g17796(.A1(new_n17858_), .A2(new_n17860_), .ZN(new_n17861_));
  INV_X1     g17797(.I(new_n17861_), .ZN(new_n17862_));
  INV_X1     g17798(.I(new_n12205_), .ZN(new_n17863_));
  NAND2_X1   g17799(.A1(new_n8702_), .A2(new_n9488_), .ZN(new_n17864_));
  NAND2_X1   g17800(.A1(new_n8711_), .A2(new_n9503_), .ZN(new_n17865_));
  AOI21_X1   g17801(.A1(new_n8719_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n17866_));
  NAND4_X1   g17802(.A1(new_n17863_), .A2(new_n17864_), .A3(new_n17865_), .A4(new_n17866_), .ZN(new_n17867_));
  XOR2_X1    g17803(.A1(new_n17867_), .A2(\a[2] ), .Z(new_n17868_));
  INV_X1     g17804(.I(new_n17868_), .ZN(new_n17869_));
  NAND2_X1   g17805(.A1(new_n8711_), .A2(new_n9488_), .ZN(new_n17870_));
  NAND2_X1   g17806(.A1(new_n8726_), .A2(new_n6925_), .ZN(new_n17871_));
  AOI21_X1   g17807(.A1(new_n8719_), .A2(new_n9503_), .B(new_n9482_), .ZN(new_n17872_));
  NAND4_X1   g17808(.A1(new_n11536_), .A2(new_n17870_), .A3(new_n17871_), .A4(new_n17872_), .ZN(new_n17873_));
  XOR2_X1    g17809(.A1(new_n17873_), .A2(\a[2] ), .Z(new_n17874_));
  INV_X1     g17810(.I(new_n17874_), .ZN(new_n17875_));
  NAND2_X1   g17811(.A1(new_n8726_), .A2(new_n9488_), .ZN(new_n17876_));
  NAND2_X1   g17812(.A1(new_n8736_), .A2(new_n9503_), .ZN(new_n17877_));
  AOI21_X1   g17813(.A1(new_n10927_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n17878_));
  NAND4_X1   g17814(.A1(new_n12500_), .A2(new_n17876_), .A3(new_n17877_), .A4(new_n17878_), .ZN(new_n17879_));
  XOR2_X1    g17815(.A1(new_n17879_), .A2(\a[2] ), .Z(new_n17880_));
  INV_X1     g17816(.I(new_n17880_), .ZN(new_n17881_));
  AOI21_X1   g17817(.A1(new_n16357_), .A2(new_n16359_), .B(new_n16437_), .ZN(new_n17882_));
  XOR2_X1    g17818(.A1(new_n16349_), .A2(new_n16355_), .Z(new_n17883_));
  AOI21_X1   g17819(.A1(new_n16437_), .A2(new_n17883_), .B(new_n17882_), .ZN(new_n17884_));
  AOI22_X1   g17820(.A1(new_n8779_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n8785_), .ZN(new_n17885_));
  NOR2_X1    g17821(.A1(new_n10871_), .A2(new_n4710_), .ZN(new_n17886_));
  OAI21_X1   g17822(.A1(new_n17886_), .A2(new_n17885_), .B(new_n4706_), .ZN(new_n17887_));
  NOR2_X1    g17823(.A1(new_n11794_), .A2(new_n17887_), .ZN(new_n17888_));
  XOR2_X1    g17824(.A1(new_n17888_), .A2(new_n4034_), .Z(new_n17889_));
  NAND2_X1   g17825(.A1(new_n17884_), .A2(new_n17889_), .ZN(new_n17890_));
  INV_X1     g17826(.I(new_n17890_), .ZN(new_n17891_));
  NOR2_X1    g17827(.A1(new_n17884_), .A2(new_n17889_), .ZN(new_n17892_));
  NOR2_X1    g17828(.A1(new_n17891_), .A2(new_n17892_), .ZN(new_n17893_));
  AOI22_X1   g17829(.A1(new_n10886_), .A2(new_n7530_), .B1(new_n10889_), .B2(new_n6789_), .ZN(new_n17894_));
  NOR2_X1    g17830(.A1(new_n10899_), .A2(new_n6785_), .ZN(new_n17895_));
  OAI21_X1   g17831(.A1(new_n17895_), .A2(new_n17894_), .B(new_n6775_), .ZN(new_n17896_));
  NOR2_X1    g17832(.A1(new_n11908_), .A2(new_n17896_), .ZN(new_n17897_));
  XOR2_X1    g17833(.A1(new_n17897_), .A2(new_n4009_), .Z(new_n17898_));
  INV_X1     g17834(.I(new_n17898_), .ZN(new_n17899_));
  INV_X1     g17835(.I(new_n16299_), .ZN(new_n17900_));
  AOI22_X1   g17836(.A1(new_n12823_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n10800_), .ZN(new_n17901_));
  AOI21_X1   g17837(.A1(new_n4709_), .A2(new_n9529_), .B(new_n17901_), .ZN(new_n17902_));
  OR3_X2     g17838(.A1(new_n13504_), .A2(new_n4707_), .A3(new_n17902_), .Z(new_n17903_));
  XOR2_X1    g17839(.A1(new_n17903_), .A2(new_n4034_), .Z(new_n17904_));
  NAND2_X1   g17840(.A1(new_n17904_), .A2(new_n17900_), .ZN(new_n17905_));
  AOI22_X1   g17841(.A1(new_n10794_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n12823_), .ZN(new_n17906_));
  AOI21_X1   g17842(.A1(new_n4709_), .A2(new_n10800_), .B(new_n17906_), .ZN(new_n17907_));
  NOR3_X1    g17843(.A1(new_n17907_), .A2(new_n14787_), .A3(new_n4707_), .ZN(new_n17908_));
  NOR2_X1    g17844(.A1(new_n4704_), .A2(new_n4705_), .ZN(new_n17909_));
  OAI21_X1   g17845(.A1(new_n12826_), .A2(new_n4719_), .B(new_n17909_), .ZN(new_n17910_));
  NOR2_X1    g17846(.A1(new_n12847_), .A2(new_n17910_), .ZN(new_n17911_));
  INV_X1     g17847(.I(new_n17911_), .ZN(new_n17912_));
  NOR2_X1    g17848(.A1(new_n12826_), .A2(new_n4704_), .ZN(new_n17913_));
  NOR4_X1    g17849(.A1(new_n17908_), .A2(new_n4034_), .A3(new_n17912_), .A4(new_n17913_), .ZN(new_n17914_));
  NOR2_X1    g17850(.A1(new_n17904_), .A2(new_n17900_), .ZN(new_n17915_));
  OAI21_X1   g17851(.A1(new_n17914_), .A2(new_n17915_), .B(new_n17905_), .ZN(new_n17916_));
  XOR2_X1    g17852(.A1(new_n16298_), .A2(new_n16300_), .Z(new_n17917_));
  AOI22_X1   g17853(.A1(new_n9529_), .A2(new_n4720_), .B1(new_n10800_), .B2(new_n6480_), .ZN(new_n17918_));
  AOI21_X1   g17854(.A1(new_n10839_), .A2(new_n4709_), .B(new_n17918_), .ZN(new_n17919_));
  OR3_X2     g17855(.A1(new_n13534_), .A2(new_n4707_), .A3(new_n17919_), .Z(new_n17920_));
  XOR2_X1    g17856(.A1(new_n17920_), .A2(\a[11] ), .Z(new_n17921_));
  NAND2_X1   g17857(.A1(new_n17921_), .A2(new_n17917_), .ZN(new_n17922_));
  NAND2_X1   g17858(.A1(new_n17922_), .A2(new_n17916_), .ZN(new_n17923_));
  INV_X1     g17859(.I(new_n17917_), .ZN(new_n17924_));
  XOR2_X1    g17860(.A1(new_n17920_), .A2(new_n4034_), .Z(new_n17925_));
  NAND2_X1   g17861(.A1(new_n17925_), .A2(new_n17924_), .ZN(new_n17926_));
  NAND2_X1   g17862(.A1(new_n17923_), .A2(new_n17926_), .ZN(new_n17927_));
  INV_X1     g17863(.I(new_n17927_), .ZN(new_n17928_));
  AOI22_X1   g17864(.A1(new_n10839_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n9529_), .ZN(new_n17929_));
  NOR2_X1    g17865(.A1(new_n10846_), .A2(new_n4710_), .ZN(new_n17930_));
  OAI21_X1   g17866(.A1(new_n17929_), .A2(new_n17930_), .B(new_n4706_), .ZN(new_n17931_));
  NOR2_X1    g17867(.A1(new_n12946_), .A2(new_n17931_), .ZN(new_n17932_));
  XOR2_X1    g17868(.A1(new_n17932_), .A2(new_n4034_), .Z(new_n17933_));
  NOR2_X1    g17869(.A1(new_n17928_), .A2(new_n17933_), .ZN(new_n17934_));
  INV_X1     g17870(.I(new_n16301_), .ZN(new_n17935_));
  NOR2_X1    g17871(.A1(new_n17935_), .A2(new_n16293_), .ZN(new_n17936_));
  NOR2_X1    g17872(.A1(new_n17936_), .A2(new_n16302_), .ZN(new_n17937_));
  AOI21_X1   g17873(.A1(new_n17928_), .A2(new_n17933_), .B(new_n17937_), .ZN(new_n17938_));
  NOR2_X1    g17874(.A1(new_n17938_), .A2(new_n17934_), .ZN(new_n17939_));
  INV_X1     g17875(.I(new_n16302_), .ZN(new_n17940_));
  XOR2_X1    g17876(.A1(new_n16288_), .A2(new_n14960_), .Z(new_n17941_));
  INV_X1     g17877(.I(new_n16289_), .ZN(new_n17942_));
  OAI21_X1   g17878(.A1(new_n17942_), .A2(new_n16303_), .B(new_n17940_), .ZN(new_n17943_));
  OAI21_X1   g17879(.A1(new_n17941_), .A2(new_n17940_), .B(new_n17943_), .ZN(new_n17944_));
  INV_X1     g17880(.I(new_n17944_), .ZN(new_n17945_));
  AOI22_X1   g17881(.A1(new_n10839_), .A2(new_n6480_), .B1(new_n12936_), .B2(new_n4720_), .ZN(new_n17946_));
  AOI21_X1   g17882(.A1(new_n4709_), .A2(new_n9479_), .B(new_n17946_), .ZN(new_n17947_));
  OR3_X2     g17883(.A1(new_n12975_), .A2(new_n4707_), .A3(new_n17947_), .Z(new_n17948_));
  XOR2_X1    g17884(.A1(new_n17948_), .A2(\a[11] ), .Z(new_n17949_));
  NAND2_X1   g17885(.A1(new_n17945_), .A2(new_n17949_), .ZN(new_n17950_));
  INV_X1     g17886(.I(new_n17950_), .ZN(new_n17951_));
  INV_X1     g17887(.I(new_n17949_), .ZN(new_n17952_));
  NAND2_X1   g17888(.A1(new_n17952_), .A2(new_n17944_), .ZN(new_n17953_));
  OAI21_X1   g17889(.A1(new_n17939_), .A2(new_n17951_), .B(new_n17953_), .ZN(new_n17954_));
  XOR2_X1    g17890(.A1(new_n16309_), .A2(new_n16305_), .Z(new_n17955_));
  INV_X1     g17891(.I(new_n16311_), .ZN(new_n17956_));
  AOI21_X1   g17892(.A1(new_n17956_), .A2(new_n16310_), .B(new_n16304_), .ZN(new_n17957_));
  AOI21_X1   g17893(.A1(new_n17955_), .A2(new_n16304_), .B(new_n17957_), .ZN(new_n17958_));
  OAI22_X1   g17894(.A1(new_n9478_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n10846_), .ZN(new_n17959_));
  NAND2_X1   g17895(.A1(new_n10854_), .A2(new_n4709_), .ZN(new_n17960_));
  AOI21_X1   g17896(.A1(new_n17959_), .A2(new_n17960_), .B(new_n4707_), .ZN(new_n17961_));
  NAND2_X1   g17897(.A1(new_n13016_), .A2(new_n17961_), .ZN(new_n17962_));
  XOR2_X1    g17898(.A1(new_n17962_), .A2(new_n4034_), .Z(new_n17963_));
  NOR2_X1    g17899(.A1(new_n17958_), .A2(new_n17963_), .ZN(new_n17964_));
  INV_X1     g17900(.I(new_n17964_), .ZN(new_n17965_));
  NAND2_X1   g17901(.A1(new_n17954_), .A2(new_n17965_), .ZN(new_n17966_));
  NAND2_X1   g17902(.A1(new_n17958_), .A2(new_n17963_), .ZN(new_n17967_));
  NAND2_X1   g17903(.A1(new_n17966_), .A2(new_n17967_), .ZN(new_n17968_));
  XNOR2_X1   g17904(.A1(new_n16312_), .A2(new_n16317_), .ZN(new_n17969_));
  XOR2_X1    g17905(.A1(new_n17969_), .A2(new_n14963_), .Z(new_n17970_));
  NOR2_X1    g17906(.A1(new_n17970_), .A2(new_n16319_), .ZN(new_n17971_));
  XNOR2_X1   g17907(.A1(new_n17969_), .A2(new_n14963_), .ZN(new_n17972_));
  NOR2_X1    g17908(.A1(new_n17972_), .A2(new_n14955_), .ZN(new_n17973_));
  OAI22_X1   g17909(.A1(new_n9478_), .A2(new_n4716_), .B1(new_n4719_), .B2(new_n10853_), .ZN(new_n17974_));
  NAND2_X1   g17910(.A1(new_n10862_), .A2(new_n4709_), .ZN(new_n17975_));
  AOI21_X1   g17911(.A1(new_n17974_), .A2(new_n17975_), .B(new_n4707_), .ZN(new_n17976_));
  NAND2_X1   g17912(.A1(new_n13484_), .A2(new_n17976_), .ZN(new_n17977_));
  XOR2_X1    g17913(.A1(new_n17977_), .A2(\a[11] ), .Z(new_n17978_));
  OAI21_X1   g17914(.A1(new_n17973_), .A2(new_n17971_), .B(new_n17978_), .ZN(new_n17979_));
  NAND2_X1   g17915(.A1(new_n17979_), .A2(new_n17968_), .ZN(new_n17980_));
  NAND2_X1   g17916(.A1(new_n17972_), .A2(new_n14955_), .ZN(new_n17981_));
  NAND2_X1   g17917(.A1(new_n17970_), .A2(new_n16319_), .ZN(new_n17982_));
  INV_X1     g17918(.I(new_n17978_), .ZN(new_n17983_));
  NAND3_X1   g17919(.A1(new_n17981_), .A2(new_n17982_), .A3(new_n17983_), .ZN(new_n17984_));
  NOR2_X1    g17920(.A1(new_n16321_), .A2(new_n16318_), .ZN(new_n17985_));
  XNOR2_X1   g17921(.A1(new_n16326_), .A2(new_n16330_), .ZN(new_n17986_));
  XNOR2_X1   g17922(.A1(new_n16326_), .A2(new_n16330_), .ZN(new_n17987_));
  NAND2_X1   g17923(.A1(new_n17987_), .A2(new_n17985_), .ZN(new_n17988_));
  OAI21_X1   g17924(.A1(new_n17985_), .A2(new_n17986_), .B(new_n17988_), .ZN(new_n17989_));
  OAI22_X1   g17925(.A1(new_n10861_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n10853_), .ZN(new_n17990_));
  NAND2_X1   g17926(.A1(new_n8785_), .A2(new_n4709_), .ZN(new_n17991_));
  AOI21_X1   g17927(.A1(new_n17991_), .A2(new_n17990_), .B(new_n4707_), .ZN(new_n17992_));
  NAND2_X1   g17928(.A1(new_n13592_), .A2(new_n17992_), .ZN(new_n17993_));
  XOR2_X1    g17929(.A1(new_n17993_), .A2(\a[11] ), .Z(new_n17994_));
  NAND2_X1   g17930(.A1(new_n17989_), .A2(new_n17994_), .ZN(new_n17995_));
  INV_X1     g17931(.I(new_n17995_), .ZN(new_n17996_));
  AOI21_X1   g17932(.A1(new_n17980_), .A2(new_n17984_), .B(new_n17996_), .ZN(new_n17997_));
  NOR2_X1    g17933(.A1(new_n17989_), .A2(new_n17994_), .ZN(new_n17998_));
  NAND2_X1   g17934(.A1(new_n16331_), .A2(new_n16332_), .ZN(new_n17999_));
  XOR2_X1    g17935(.A1(new_n16337_), .A2(new_n16342_), .Z(new_n18000_));
  NOR2_X1    g17936(.A1(new_n16345_), .A2(new_n16343_), .ZN(new_n18001_));
  NOR2_X1    g17937(.A1(new_n17999_), .A2(new_n18001_), .ZN(new_n18002_));
  AOI21_X1   g17938(.A1(new_n17999_), .A2(new_n18000_), .B(new_n18002_), .ZN(new_n18003_));
  OAI22_X1   g17939(.A1(new_n8784_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n10861_), .ZN(new_n18004_));
  NAND2_X1   g17940(.A1(new_n8779_), .A2(new_n4709_), .ZN(new_n18005_));
  AOI21_X1   g17941(.A1(new_n18005_), .A2(new_n18004_), .B(new_n4707_), .ZN(new_n18006_));
  NAND2_X1   g17942(.A1(new_n12814_), .A2(new_n18006_), .ZN(new_n18007_));
  XOR2_X1    g17943(.A1(new_n18007_), .A2(new_n4034_), .Z(new_n18008_));
  NOR2_X1    g17944(.A1(new_n18003_), .A2(new_n18008_), .ZN(new_n18009_));
  INV_X1     g17945(.I(new_n18009_), .ZN(new_n18010_));
  OAI21_X1   g17946(.A1(new_n17997_), .A2(new_n17998_), .B(new_n18010_), .ZN(new_n18011_));
  NAND2_X1   g17947(.A1(new_n18003_), .A2(new_n18008_), .ZN(new_n18012_));
  NAND2_X1   g17948(.A1(new_n18011_), .A2(new_n18012_), .ZN(new_n18013_));
  OAI22_X1   g17949(.A1(new_n10871_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8778_), .ZN(new_n18014_));
  NAND2_X1   g17950(.A1(new_n10886_), .A2(new_n6784_), .ZN(new_n18015_));
  AOI21_X1   g17951(.A1(new_n18015_), .A2(new_n18014_), .B(new_n6776_), .ZN(new_n18016_));
  NAND2_X1   g17952(.A1(new_n13103_), .A2(new_n18016_), .ZN(new_n18017_));
  XOR2_X1    g17953(.A1(new_n18017_), .A2(\a[8] ), .Z(new_n18018_));
  INV_X1     g17954(.I(new_n17998_), .ZN(new_n18019_));
  AOI22_X1   g17955(.A1(new_n17980_), .A2(new_n17984_), .B1(new_n17995_), .B2(new_n18019_), .ZN(new_n18020_));
  NAND2_X1   g17956(.A1(new_n17980_), .A2(new_n17984_), .ZN(new_n18021_));
  XNOR2_X1   g17957(.A1(new_n17989_), .A2(new_n17994_), .ZN(new_n18022_));
  NOR2_X1    g17958(.A1(new_n18021_), .A2(new_n18022_), .ZN(new_n18023_));
  NOR2_X1    g17959(.A1(new_n18023_), .A2(new_n18020_), .ZN(new_n18024_));
  INV_X1     g17960(.I(new_n18024_), .ZN(new_n18025_));
  NAND2_X1   g17961(.A1(new_n18025_), .A2(new_n18018_), .ZN(new_n18026_));
  INV_X1     g17962(.I(new_n17968_), .ZN(new_n18027_));
  AOI21_X1   g17963(.A1(new_n17979_), .A2(new_n17984_), .B(new_n18027_), .ZN(new_n18028_));
  NAND3_X1   g17964(.A1(new_n17981_), .A2(new_n17982_), .A3(new_n17978_), .ZN(new_n18029_));
  OAI21_X1   g17965(.A1(new_n17973_), .A2(new_n17971_), .B(new_n17983_), .ZN(new_n18030_));
  AOI21_X1   g17966(.A1(new_n18030_), .A2(new_n18029_), .B(new_n17968_), .ZN(new_n18031_));
  AOI22_X1   g17967(.A1(new_n8779_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n8785_), .ZN(new_n18032_));
  NOR2_X1    g17968(.A1(new_n10871_), .A2(new_n6785_), .ZN(new_n18033_));
  OAI21_X1   g17969(.A1(new_n18033_), .A2(new_n18032_), .B(new_n6775_), .ZN(new_n18034_));
  NOR2_X1    g17970(.A1(new_n11794_), .A2(new_n18034_), .ZN(new_n18035_));
  XOR2_X1    g17971(.A1(new_n18035_), .A2(new_n4009_), .Z(new_n18036_));
  INV_X1     g17972(.I(new_n18036_), .ZN(new_n18037_));
  NOR3_X1    g17973(.A1(new_n18028_), .A2(new_n18031_), .A3(new_n18037_), .ZN(new_n18038_));
  AOI21_X1   g17974(.A1(new_n17981_), .A2(new_n17982_), .B(new_n17983_), .ZN(new_n18039_));
  INV_X1     g17975(.I(new_n17984_), .ZN(new_n18040_));
  OAI21_X1   g17976(.A1(new_n18040_), .A2(new_n18039_), .B(new_n17968_), .ZN(new_n18041_));
  INV_X1     g17977(.I(new_n18031_), .ZN(new_n18042_));
  AOI21_X1   g17978(.A1(new_n18042_), .A2(new_n18041_), .B(new_n18036_), .ZN(new_n18043_));
  INV_X1     g17979(.I(new_n17939_), .ZN(new_n18044_));
  XNOR2_X1   g17980(.A1(new_n17944_), .A2(new_n17949_), .ZN(new_n18045_));
  NAND2_X1   g17981(.A1(new_n18044_), .A2(new_n18045_), .ZN(new_n18046_));
  NAND2_X1   g17982(.A1(new_n17950_), .A2(new_n17953_), .ZN(new_n18047_));
  NAND2_X1   g17983(.A1(new_n17939_), .A2(new_n18047_), .ZN(new_n18048_));
  NAND2_X1   g17984(.A1(new_n18046_), .A2(new_n18048_), .ZN(new_n18049_));
  OAI22_X1   g17985(.A1(new_n10861_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n10853_), .ZN(new_n18050_));
  NAND2_X1   g17986(.A1(new_n8785_), .A2(new_n6784_), .ZN(new_n18051_));
  AOI21_X1   g17987(.A1(new_n18051_), .A2(new_n18050_), .B(new_n6776_), .ZN(new_n18052_));
  NAND2_X1   g17988(.A1(new_n13592_), .A2(new_n18052_), .ZN(new_n18053_));
  XOR2_X1    g17989(.A1(new_n18053_), .A2(\a[8] ), .Z(new_n18054_));
  NOR2_X1    g17990(.A1(new_n18049_), .A2(new_n18054_), .ZN(new_n18055_));
  XOR2_X1    g17991(.A1(new_n17958_), .A2(new_n17963_), .Z(new_n18056_));
  NAND2_X1   g17992(.A1(new_n17954_), .A2(new_n18056_), .ZN(new_n18057_));
  INV_X1     g17993(.I(new_n17967_), .ZN(new_n18058_));
  NOR2_X1    g17994(.A1(new_n18058_), .A2(new_n17964_), .ZN(new_n18059_));
  OAI21_X1   g17995(.A1(new_n17954_), .A2(new_n18059_), .B(new_n18057_), .ZN(new_n18060_));
  OAI22_X1   g17996(.A1(new_n8784_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n10861_), .ZN(new_n18061_));
  NAND2_X1   g17997(.A1(new_n8779_), .A2(new_n6784_), .ZN(new_n18062_));
  AOI21_X1   g17998(.A1(new_n18062_), .A2(new_n18061_), .B(new_n6776_), .ZN(new_n18063_));
  NAND2_X1   g17999(.A1(new_n12814_), .A2(new_n18063_), .ZN(new_n18064_));
  XOR2_X1    g18000(.A1(new_n18064_), .A2(\a[8] ), .Z(new_n18065_));
  NAND2_X1   g18001(.A1(new_n18060_), .A2(new_n18065_), .ZN(new_n18066_));
  NOR2_X1    g18002(.A1(new_n18060_), .A2(new_n18065_), .ZN(new_n18067_));
  AOI21_X1   g18003(.A1(new_n18055_), .A2(new_n18066_), .B(new_n18067_), .ZN(new_n18068_));
  INV_X1     g18004(.I(new_n18068_), .ZN(new_n18069_));
  NOR3_X1    g18005(.A1(new_n18043_), .A2(new_n18038_), .A3(new_n18069_), .ZN(new_n18070_));
  NOR3_X1    g18006(.A1(new_n18023_), .A2(new_n18018_), .A3(new_n18020_), .ZN(new_n18071_));
  OAI21_X1   g18007(.A1(new_n18023_), .A2(new_n18020_), .B(new_n18018_), .ZN(new_n18072_));
  INV_X1     g18008(.I(new_n18072_), .ZN(new_n18073_));
  NAND3_X1   g18009(.A1(new_n18042_), .A2(new_n18041_), .A3(new_n18036_), .ZN(new_n18074_));
  OAI21_X1   g18010(.A1(new_n18073_), .A2(new_n18071_), .B(new_n18074_), .ZN(new_n18075_));
  OAI21_X1   g18011(.A1(new_n18075_), .A2(new_n18070_), .B(new_n18026_), .ZN(new_n18076_));
  XOR2_X1    g18012(.A1(new_n18003_), .A2(new_n18008_), .Z(new_n18077_));
  OAI21_X1   g18013(.A1(new_n17997_), .A2(new_n17998_), .B(new_n18077_), .ZN(new_n18078_));
  NOR2_X1    g18014(.A1(new_n17997_), .A2(new_n17998_), .ZN(new_n18079_));
  NAND2_X1   g18015(.A1(new_n18010_), .A2(new_n18012_), .ZN(new_n18080_));
  NAND2_X1   g18016(.A1(new_n18079_), .A2(new_n18080_), .ZN(new_n18081_));
  NAND2_X1   g18017(.A1(new_n18081_), .A2(new_n18078_), .ZN(new_n18082_));
  AOI22_X1   g18018(.A1(new_n10886_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n10872_), .ZN(new_n18083_));
  NOR2_X1    g18019(.A1(new_n10892_), .A2(new_n6785_), .ZN(new_n18084_));
  OAI21_X1   g18020(.A1(new_n18083_), .A2(new_n18084_), .B(new_n6775_), .ZN(new_n18085_));
  NOR2_X1    g18021(.A1(new_n12776_), .A2(new_n18085_), .ZN(new_n18086_));
  XOR2_X1    g18022(.A1(new_n18086_), .A2(new_n4009_), .Z(new_n18087_));
  NAND2_X1   g18023(.A1(new_n18082_), .A2(new_n18087_), .ZN(new_n18088_));
  NAND2_X1   g18024(.A1(new_n18076_), .A2(new_n18088_), .ZN(new_n18089_));
  NOR2_X1    g18025(.A1(new_n18082_), .A2(new_n18087_), .ZN(new_n18090_));
  INV_X1     g18026(.I(new_n18090_), .ZN(new_n18091_));
  NAND3_X1   g18027(.A1(new_n18089_), .A2(new_n18013_), .A3(new_n18091_), .ZN(new_n18092_));
  INV_X1     g18028(.I(new_n18013_), .ZN(new_n18093_));
  OAI21_X1   g18029(.A1(new_n18028_), .A2(new_n18031_), .B(new_n18037_), .ZN(new_n18094_));
  NAND3_X1   g18030(.A1(new_n18074_), .A2(new_n18094_), .A3(new_n18068_), .ZN(new_n18095_));
  INV_X1     g18031(.I(new_n18071_), .ZN(new_n18096_));
  AOI21_X1   g18032(.A1(new_n18096_), .A2(new_n18072_), .B(new_n18038_), .ZN(new_n18097_));
  NAND2_X1   g18033(.A1(new_n18097_), .A2(new_n18095_), .ZN(new_n18098_));
  INV_X1     g18034(.I(new_n18088_), .ZN(new_n18099_));
  AOI21_X1   g18035(.A1(new_n18098_), .A2(new_n18026_), .B(new_n18099_), .ZN(new_n18100_));
  OAI21_X1   g18036(.A1(new_n18100_), .A2(new_n18090_), .B(new_n18093_), .ZN(new_n18101_));
  AOI21_X1   g18037(.A1(new_n18101_), .A2(new_n18092_), .B(new_n17899_), .ZN(new_n18102_));
  NOR3_X1    g18038(.A1(new_n18100_), .A2(new_n18093_), .A3(new_n18090_), .ZN(new_n18103_));
  AOI21_X1   g18039(.A1(new_n18089_), .A2(new_n18091_), .B(new_n18013_), .ZN(new_n18104_));
  NOR3_X1    g18040(.A1(new_n18103_), .A2(new_n18104_), .A3(new_n17898_), .ZN(new_n18105_));
  OAI21_X1   g18041(.A1(new_n18105_), .A2(new_n18102_), .B(new_n17893_), .ZN(new_n18106_));
  INV_X1     g18042(.I(new_n17893_), .ZN(new_n18107_));
  OAI21_X1   g18043(.A1(new_n18103_), .A2(new_n18104_), .B(new_n17898_), .ZN(new_n18108_));
  NAND3_X1   g18044(.A1(new_n18101_), .A2(new_n18092_), .A3(new_n17899_), .ZN(new_n18109_));
  NAND3_X1   g18045(.A1(new_n18108_), .A2(new_n18109_), .A3(new_n18107_), .ZN(new_n18110_));
  AOI22_X1   g18046(.A1(new_n6846_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n8799_), .ZN(new_n18111_));
  NOR2_X1    g18047(.A1(new_n8758_), .A2(new_n6839_), .ZN(new_n18112_));
  OAI21_X1   g18048(.A1(new_n18111_), .A2(new_n18112_), .B(new_n6835_), .ZN(new_n18113_));
  NOR2_X1    g18049(.A1(new_n12053_), .A2(new_n18113_), .ZN(new_n18114_));
  XOR2_X1    g18050(.A1(new_n18114_), .A2(new_n65_), .Z(new_n18115_));
  AOI21_X1   g18051(.A1(new_n18106_), .A2(new_n18110_), .B(new_n18115_), .ZN(new_n18116_));
  AOI21_X1   g18052(.A1(new_n18089_), .A2(new_n18091_), .B(new_n17898_), .ZN(new_n18117_));
  NOR2_X1    g18053(.A1(new_n18093_), .A2(new_n18107_), .ZN(new_n18118_));
  NOR2_X1    g18054(.A1(new_n18013_), .A2(new_n17893_), .ZN(new_n18119_));
  OAI21_X1   g18055(.A1(new_n18118_), .A2(new_n18119_), .B(new_n17898_), .ZN(new_n18120_));
  NOR3_X1    g18056(.A1(new_n18100_), .A2(new_n18090_), .A3(new_n18120_), .ZN(new_n18121_));
  AOI22_X1   g18057(.A1(new_n16358_), .A2(new_n16359_), .B1(new_n16441_), .B2(new_n16368_), .ZN(new_n18122_));
  XNOR2_X1   g18058(.A1(new_n16362_), .A2(new_n16367_), .ZN(new_n18123_));
  NOR3_X1    g18059(.A1(new_n18123_), .A2(new_n16438_), .A3(new_n16439_), .ZN(new_n18124_));
  NOR2_X1    g18060(.A1(new_n18124_), .A2(new_n18122_), .ZN(new_n18125_));
  INV_X1     g18061(.I(new_n18125_), .ZN(new_n18126_));
  OAI22_X1   g18062(.A1(new_n10871_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n8778_), .ZN(new_n18127_));
  NAND2_X1   g18063(.A1(new_n10886_), .A2(new_n4709_), .ZN(new_n18128_));
  AOI21_X1   g18064(.A1(new_n18128_), .A2(new_n18127_), .B(new_n4707_), .ZN(new_n18129_));
  NAND2_X1   g18065(.A1(new_n13103_), .A2(new_n18129_), .ZN(new_n18130_));
  XOR2_X1    g18066(.A1(new_n18130_), .A2(\a[11] ), .Z(new_n18131_));
  INV_X1     g18067(.I(new_n18131_), .ZN(new_n18132_));
  NAND3_X1   g18068(.A1(new_n18011_), .A2(new_n17893_), .A3(new_n18012_), .ZN(new_n18133_));
  AOI21_X1   g18069(.A1(new_n18133_), .A2(new_n17890_), .B(new_n18132_), .ZN(new_n18134_));
  INV_X1     g18070(.I(new_n18134_), .ZN(new_n18135_));
  NAND3_X1   g18071(.A1(new_n18133_), .A2(new_n17890_), .A3(new_n18132_), .ZN(new_n18136_));
  AOI21_X1   g18072(.A1(new_n18135_), .A2(new_n18136_), .B(new_n18126_), .ZN(new_n18137_));
  INV_X1     g18073(.I(new_n18136_), .ZN(new_n18138_));
  NOR3_X1    g18074(.A1(new_n18138_), .A2(new_n18125_), .A3(new_n18134_), .ZN(new_n18139_));
  AOI22_X1   g18075(.A1(new_n11899_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n10889_), .ZN(new_n18140_));
  NOR2_X1    g18076(.A1(new_n8774_), .A2(new_n6785_), .ZN(new_n18141_));
  OAI21_X1   g18077(.A1(new_n18141_), .A2(new_n18140_), .B(new_n6775_), .ZN(new_n18142_));
  NOR2_X1    g18078(.A1(new_n11945_), .A2(new_n18142_), .ZN(new_n18143_));
  XOR2_X1    g18079(.A1(new_n18143_), .A2(new_n4009_), .Z(new_n18144_));
  NOR3_X1    g18080(.A1(new_n18137_), .A2(new_n18139_), .A3(new_n18144_), .ZN(new_n18145_));
  OAI21_X1   g18081(.A1(new_n18138_), .A2(new_n18134_), .B(new_n18125_), .ZN(new_n18146_));
  NAND3_X1   g18082(.A1(new_n18135_), .A2(new_n18126_), .A3(new_n18136_), .ZN(new_n18147_));
  INV_X1     g18083(.I(new_n18144_), .ZN(new_n18148_));
  AOI21_X1   g18084(.A1(new_n18147_), .A2(new_n18146_), .B(new_n18148_), .ZN(new_n18149_));
  NOR4_X1    g18085(.A1(new_n18121_), .A2(new_n18117_), .A3(new_n18145_), .A4(new_n18149_), .ZN(new_n18150_));
  OAI21_X1   g18086(.A1(new_n18100_), .A2(new_n18090_), .B(new_n17899_), .ZN(new_n18151_));
  INV_X1     g18087(.I(new_n18120_), .ZN(new_n18152_));
  NAND3_X1   g18088(.A1(new_n18089_), .A2(new_n18152_), .A3(new_n18091_), .ZN(new_n18153_));
  NAND3_X1   g18089(.A1(new_n18147_), .A2(new_n18146_), .A3(new_n18148_), .ZN(new_n18154_));
  OAI21_X1   g18090(.A1(new_n18137_), .A2(new_n18139_), .B(new_n18144_), .ZN(new_n18155_));
  AOI22_X1   g18091(.A1(new_n18151_), .A2(new_n18153_), .B1(new_n18154_), .B2(new_n18155_), .ZN(new_n18156_));
  OAI22_X1   g18092(.A1(new_n8758_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8766_), .ZN(new_n18157_));
  NAND2_X1   g18093(.A1(new_n8746_), .A2(new_n6838_), .ZN(new_n18158_));
  AOI21_X1   g18094(.A1(new_n18158_), .A2(new_n18157_), .B(new_n6836_), .ZN(new_n18159_));
  NAND2_X1   g18095(.A1(new_n11964_), .A2(new_n18159_), .ZN(new_n18160_));
  XOR2_X1    g18096(.A1(new_n18160_), .A2(\a[5] ), .Z(new_n18161_));
  INV_X1     g18097(.I(new_n18161_), .ZN(new_n18162_));
  NOR3_X1    g18098(.A1(new_n18156_), .A2(new_n18150_), .A3(new_n18162_), .ZN(new_n18163_));
  INV_X1     g18099(.I(new_n18163_), .ZN(new_n18164_));
  OAI21_X1   g18100(.A1(new_n18156_), .A2(new_n18150_), .B(new_n18162_), .ZN(new_n18165_));
  INV_X1     g18101(.I(new_n18165_), .ZN(new_n18166_));
  AOI21_X1   g18102(.A1(new_n18116_), .A2(new_n18164_), .B(new_n18166_), .ZN(new_n18167_));
  XOR2_X1    g18103(.A1(new_n18125_), .A2(new_n18131_), .Z(new_n18168_));
  NAND3_X1   g18104(.A1(new_n18133_), .A2(new_n17890_), .A3(new_n18168_), .ZN(new_n18169_));
  OAI21_X1   g18105(.A1(new_n18125_), .A2(new_n18132_), .B(new_n18169_), .ZN(new_n18170_));
  NAND2_X1   g18106(.A1(new_n16440_), .A2(new_n16441_), .ZN(new_n18171_));
  XOR2_X1    g18107(.A1(new_n16382_), .A2(new_n16383_), .Z(new_n18172_));
  NAND2_X1   g18108(.A1(new_n18171_), .A2(new_n18172_), .ZN(new_n18173_));
  NOR2_X1    g18109(.A1(new_n16444_), .A2(new_n16442_), .ZN(new_n18174_));
  OAI21_X1   g18110(.A1(new_n18171_), .A2(new_n18174_), .B(new_n18173_), .ZN(new_n18175_));
  AOI22_X1   g18111(.A1(new_n10886_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n10872_), .ZN(new_n18176_));
  NOR2_X1    g18112(.A1(new_n10892_), .A2(new_n4710_), .ZN(new_n18177_));
  OAI21_X1   g18113(.A1(new_n18176_), .A2(new_n18177_), .B(new_n4706_), .ZN(new_n18178_));
  NOR2_X1    g18114(.A1(new_n12776_), .A2(new_n18178_), .ZN(new_n18179_));
  XOR2_X1    g18115(.A1(new_n18179_), .A2(new_n4034_), .Z(new_n18180_));
  XNOR2_X1   g18116(.A1(new_n18175_), .A2(new_n18180_), .ZN(new_n18181_));
  INV_X1     g18117(.I(new_n18181_), .ZN(new_n18182_));
  NAND2_X1   g18118(.A1(new_n18175_), .A2(new_n18180_), .ZN(new_n18183_));
  OR2_X2     g18119(.A1(new_n18175_), .A2(new_n18180_), .Z(new_n18184_));
  NAND2_X1   g18120(.A1(new_n18184_), .A2(new_n18183_), .ZN(new_n18185_));
  INV_X1     g18121(.I(new_n18185_), .ZN(new_n18186_));
  NOR2_X1    g18122(.A1(new_n18170_), .A2(new_n18186_), .ZN(new_n18187_));
  AOI21_X1   g18123(.A1(new_n18170_), .A2(new_n18182_), .B(new_n18187_), .ZN(new_n18188_));
  NAND4_X1   g18124(.A1(new_n18151_), .A2(new_n18153_), .A3(new_n18155_), .A4(new_n18154_), .ZN(new_n18189_));
  OAI22_X1   g18125(.A1(new_n8774_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n10899_), .ZN(new_n18190_));
  NAND2_X1   g18126(.A1(new_n11996_), .A2(new_n6784_), .ZN(new_n18191_));
  AOI21_X1   g18127(.A1(new_n18191_), .A2(new_n18190_), .B(new_n6776_), .ZN(new_n18192_));
  NAND2_X1   g18128(.A1(new_n12001_), .A2(new_n18192_), .ZN(new_n18193_));
  XOR2_X1    g18129(.A1(new_n18193_), .A2(\a[8] ), .Z(new_n18194_));
  INV_X1     g18130(.I(new_n18194_), .ZN(new_n18195_));
  AOI21_X1   g18131(.A1(new_n18189_), .A2(new_n18155_), .B(new_n18195_), .ZN(new_n18196_));
  NOR3_X1    g18132(.A1(new_n18150_), .A2(new_n18149_), .A3(new_n18194_), .ZN(new_n18197_));
  OAI21_X1   g18133(.A1(new_n18197_), .A2(new_n18196_), .B(new_n18188_), .ZN(new_n18198_));
  INV_X1     g18134(.I(new_n18188_), .ZN(new_n18199_));
  OAI21_X1   g18135(.A1(new_n18150_), .A2(new_n18149_), .B(new_n18194_), .ZN(new_n18200_));
  NAND3_X1   g18136(.A1(new_n18189_), .A2(new_n18155_), .A3(new_n18195_), .ZN(new_n18201_));
  NAND3_X1   g18137(.A1(new_n18200_), .A2(new_n18201_), .A3(new_n18199_), .ZN(new_n18202_));
  OAI22_X1   g18138(.A1(new_n8745_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8758_), .ZN(new_n18203_));
  NAND2_X1   g18139(.A1(new_n8752_), .A2(new_n6838_), .ZN(new_n18204_));
  AOI21_X1   g18140(.A1(new_n18204_), .A2(new_n18203_), .B(new_n6836_), .ZN(new_n18205_));
  NAND2_X1   g18141(.A1(new_n12189_), .A2(new_n18205_), .ZN(new_n18206_));
  XOR2_X1    g18142(.A1(new_n18206_), .A2(\a[5] ), .Z(new_n18207_));
  NAND3_X1   g18143(.A1(new_n18198_), .A2(new_n18202_), .A3(new_n18207_), .ZN(new_n18208_));
  AOI21_X1   g18144(.A1(new_n18200_), .A2(new_n18201_), .B(new_n18199_), .ZN(new_n18209_));
  NOR3_X1    g18145(.A1(new_n18197_), .A2(new_n18196_), .A3(new_n18188_), .ZN(new_n18210_));
  INV_X1     g18146(.I(new_n18207_), .ZN(new_n18211_));
  OAI21_X1   g18147(.A1(new_n18210_), .A2(new_n18209_), .B(new_n18211_), .ZN(new_n18212_));
  AOI21_X1   g18148(.A1(new_n18212_), .A2(new_n18208_), .B(new_n18167_), .ZN(new_n18213_));
  AOI21_X1   g18149(.A1(new_n18108_), .A2(new_n18109_), .B(new_n18107_), .ZN(new_n18214_));
  NOR3_X1    g18150(.A1(new_n18105_), .A2(new_n18102_), .A3(new_n17893_), .ZN(new_n18215_));
  INV_X1     g18151(.I(new_n18115_), .ZN(new_n18216_));
  OAI21_X1   g18152(.A1(new_n18215_), .A2(new_n18214_), .B(new_n18216_), .ZN(new_n18217_));
  OAI21_X1   g18153(.A1(new_n18217_), .A2(new_n18163_), .B(new_n18165_), .ZN(new_n18218_));
  OAI21_X1   g18154(.A1(new_n18210_), .A2(new_n18209_), .B(new_n18207_), .ZN(new_n18219_));
  NAND3_X1   g18155(.A1(new_n18198_), .A2(new_n18202_), .A3(new_n18211_), .ZN(new_n18220_));
  AOI21_X1   g18156(.A1(new_n18219_), .A2(new_n18220_), .B(new_n18218_), .ZN(new_n18221_));
  NOR3_X1    g18157(.A1(new_n18221_), .A2(new_n18213_), .A3(new_n17880_), .ZN(new_n18222_));
  NOR3_X1    g18158(.A1(new_n18210_), .A2(new_n18209_), .A3(new_n18211_), .ZN(new_n18223_));
  AOI21_X1   g18159(.A1(new_n18198_), .A2(new_n18202_), .B(new_n18207_), .ZN(new_n18224_));
  OAI21_X1   g18160(.A1(new_n18223_), .A2(new_n18224_), .B(new_n18218_), .ZN(new_n18225_));
  AOI21_X1   g18161(.A1(new_n18198_), .A2(new_n18202_), .B(new_n18211_), .ZN(new_n18226_));
  NOR3_X1    g18162(.A1(new_n18210_), .A2(new_n18209_), .A3(new_n18207_), .ZN(new_n18227_));
  OAI21_X1   g18163(.A1(new_n18227_), .A2(new_n18226_), .B(new_n18167_), .ZN(new_n18228_));
  AOI21_X1   g18164(.A1(new_n18225_), .A2(new_n18228_), .B(new_n17881_), .ZN(new_n18229_));
  NOR2_X1    g18165(.A1(new_n18229_), .A2(new_n18222_), .ZN(new_n18230_));
  NOR2_X1    g18166(.A1(new_n18230_), .A2(new_n17881_), .ZN(new_n18231_));
  NAND2_X1   g18167(.A1(new_n8752_), .A2(new_n9488_), .ZN(new_n18232_));
  NAND2_X1   g18168(.A1(new_n8746_), .A2(new_n9503_), .ZN(new_n18233_));
  AOI21_X1   g18169(.A1(new_n8761_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n18234_));
  NAND4_X1   g18170(.A1(new_n12189_), .A2(new_n18232_), .A3(new_n18233_), .A4(new_n18234_), .ZN(new_n18235_));
  XOR2_X1    g18171(.A1(new_n18235_), .A2(\a[2] ), .Z(new_n18236_));
  NAND2_X1   g18172(.A1(new_n8746_), .A2(new_n9488_), .ZN(new_n18237_));
  NAND2_X1   g18173(.A1(new_n8761_), .A2(new_n9503_), .ZN(new_n18238_));
  AOI21_X1   g18174(.A1(new_n11996_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n18239_));
  NAND4_X1   g18175(.A1(new_n11964_), .A2(new_n18237_), .A3(new_n18238_), .A4(new_n18239_), .ZN(new_n18240_));
  XOR2_X1    g18176(.A1(new_n18240_), .A2(\a[2] ), .Z(new_n18241_));
  INV_X1     g18177(.I(new_n18241_), .ZN(new_n18242_));
  OAI22_X1   g18178(.A1(new_n8774_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n10899_), .ZN(new_n18243_));
  OAI21_X1   g18179(.A1(new_n8766_), .A2(new_n9489_), .B(new_n18243_), .ZN(new_n18244_));
  AOI21_X1   g18180(.A1(new_n12001_), .A2(new_n6922_), .B(new_n18244_), .ZN(new_n18245_));
  XOR2_X1    g18181(.A1(new_n18245_), .A2(\a[2] ), .Z(new_n18246_));
  INV_X1     g18182(.I(new_n18246_), .ZN(new_n18247_));
  XOR2_X1    g18183(.A1(new_n18049_), .A2(new_n18054_), .Z(new_n18248_));
  OAI22_X1   g18184(.A1(new_n10871_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8778_), .ZN(new_n18249_));
  NAND2_X1   g18185(.A1(new_n10886_), .A2(new_n6838_), .ZN(new_n18250_));
  AOI21_X1   g18186(.A1(new_n18250_), .A2(new_n18249_), .B(new_n6836_), .ZN(new_n18251_));
  NAND2_X1   g18187(.A1(new_n13103_), .A2(new_n18251_), .ZN(new_n18252_));
  XOR2_X1    g18188(.A1(new_n18252_), .A2(\a[5] ), .Z(new_n18253_));
  NOR2_X1    g18189(.A1(new_n18248_), .A2(new_n18253_), .ZN(new_n18254_));
  OAI22_X1   g18190(.A1(new_n10775_), .A2(new_n6783_), .B1(new_n6788_), .B2(new_n10777_), .ZN(new_n18255_));
  NAND2_X1   g18191(.A1(new_n9529_), .A2(new_n6784_), .ZN(new_n18256_));
  AOI21_X1   g18192(.A1(new_n18255_), .A2(new_n18256_), .B(new_n6776_), .ZN(new_n18257_));
  NAND3_X1   g18193(.A1(new_n12883_), .A2(new_n4009_), .A3(new_n18257_), .ZN(new_n18258_));
  OAI21_X1   g18194(.A1(new_n13502_), .A2(new_n13503_), .B(new_n18257_), .ZN(new_n18259_));
  NAND2_X1   g18195(.A1(new_n18259_), .A2(\a[8] ), .ZN(new_n18260_));
  AOI21_X1   g18196(.A1(new_n18260_), .A2(new_n18258_), .B(new_n17913_), .ZN(new_n18261_));
  NOR2_X1    g18197(.A1(new_n10775_), .A2(new_n6788_), .ZN(new_n18262_));
  NOR2_X1    g18198(.A1(new_n12826_), .A2(new_n6783_), .ZN(new_n18263_));
  OAI22_X1   g18199(.A1(new_n18263_), .A2(new_n18262_), .B1(new_n6785_), .B2(new_n10777_), .ZN(new_n18264_));
  AOI21_X1   g18200(.A1(new_n12829_), .A2(new_n12827_), .B(new_n6776_), .ZN(new_n18265_));
  NAND2_X1   g18201(.A1(new_n18265_), .A2(new_n18264_), .ZN(new_n18266_));
  NOR2_X1    g18202(.A1(new_n6773_), .A2(new_n6774_), .ZN(new_n18267_));
  OAI21_X1   g18203(.A1(new_n12826_), .A2(new_n6788_), .B(new_n18267_), .ZN(new_n18268_));
  NOR2_X1    g18204(.A1(new_n12847_), .A2(new_n18268_), .ZN(new_n18269_));
  NOR2_X1    g18205(.A1(new_n12826_), .A2(new_n6773_), .ZN(new_n18270_));
  INV_X1     g18206(.I(new_n18270_), .ZN(new_n18271_));
  NAND4_X1   g18207(.A1(new_n18266_), .A2(\a[8] ), .A3(new_n18269_), .A4(new_n18271_), .ZN(new_n18272_));
  NAND3_X1   g18208(.A1(new_n18260_), .A2(new_n18258_), .A3(new_n17913_), .ZN(new_n18273_));
  AOI21_X1   g18209(.A1(new_n18272_), .A2(new_n18273_), .B(new_n18261_), .ZN(new_n18274_));
  NAND2_X1   g18210(.A1(new_n17911_), .A2(new_n4034_), .ZN(new_n18275_));
  NOR2_X1    g18211(.A1(new_n17911_), .A2(new_n4034_), .ZN(new_n18276_));
  INV_X1     g18212(.I(new_n18276_), .ZN(new_n18277_));
  NOR2_X1    g18213(.A1(new_n17913_), .A2(new_n4034_), .ZN(new_n18278_));
  INV_X1     g18214(.I(new_n18278_), .ZN(new_n18279_));
  NAND3_X1   g18215(.A1(new_n18277_), .A2(new_n18275_), .A3(new_n18279_), .ZN(new_n18280_));
  NOR3_X1    g18216(.A1(new_n17911_), .A2(new_n4034_), .A3(new_n17913_), .ZN(new_n18281_));
  INV_X1     g18217(.I(new_n18281_), .ZN(new_n18282_));
  NAND2_X1   g18218(.A1(new_n18280_), .A2(new_n18282_), .ZN(new_n18283_));
  AOI22_X1   g18219(.A1(new_n9529_), .A2(new_n6789_), .B1(new_n10800_), .B2(new_n7530_), .ZN(new_n18284_));
  AOI21_X1   g18220(.A1(new_n10839_), .A2(new_n6784_), .B(new_n18284_), .ZN(new_n18285_));
  NOR3_X1    g18221(.A1(new_n13534_), .A2(new_n18285_), .A3(new_n6776_), .ZN(new_n18286_));
  NAND2_X1   g18222(.A1(new_n18286_), .A2(new_n4009_), .ZN(new_n18287_));
  NOR2_X1    g18223(.A1(new_n18285_), .A2(new_n6776_), .ZN(new_n18288_));
  NAND2_X1   g18224(.A1(new_n12910_), .A2(new_n18288_), .ZN(new_n18289_));
  NAND2_X1   g18225(.A1(new_n18289_), .A2(\a[8] ), .ZN(new_n18290_));
  NAND3_X1   g18226(.A1(new_n18283_), .A2(new_n18287_), .A3(new_n18290_), .ZN(new_n18291_));
  INV_X1     g18227(.I(new_n18291_), .ZN(new_n18292_));
  INV_X1     g18228(.I(new_n18275_), .ZN(new_n18293_));
  NOR3_X1    g18229(.A1(new_n18293_), .A2(new_n18276_), .A3(new_n18278_), .ZN(new_n18294_));
  NOR2_X1    g18230(.A1(new_n18294_), .A2(new_n18281_), .ZN(new_n18295_));
  NOR2_X1    g18231(.A1(new_n18289_), .A2(\a[8] ), .ZN(new_n18296_));
  NOR2_X1    g18232(.A1(new_n18286_), .A2(new_n4009_), .ZN(new_n18297_));
  OAI21_X1   g18233(.A1(new_n18296_), .A2(new_n18297_), .B(new_n18295_), .ZN(new_n18298_));
  OAI21_X1   g18234(.A1(new_n18292_), .A2(new_n18274_), .B(new_n18298_), .ZN(new_n18299_));
  XOR2_X1    g18235(.A1(new_n17908_), .A2(\a[11] ), .Z(new_n18300_));
  NOR3_X1    g18236(.A1(new_n17912_), .A2(new_n4034_), .A3(new_n17913_), .ZN(new_n18301_));
  XOR2_X1    g18237(.A1(new_n18300_), .A2(new_n18301_), .Z(new_n18302_));
  AOI22_X1   g18238(.A1(new_n10839_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n9529_), .ZN(new_n18303_));
  NOR2_X1    g18239(.A1(new_n10846_), .A2(new_n6785_), .ZN(new_n18304_));
  OAI21_X1   g18240(.A1(new_n18303_), .A2(new_n18304_), .B(new_n6775_), .ZN(new_n18305_));
  NOR2_X1    g18241(.A1(new_n12946_), .A2(new_n18305_), .ZN(new_n18306_));
  XOR2_X1    g18242(.A1(new_n18306_), .A2(new_n4009_), .Z(new_n18307_));
  NAND2_X1   g18243(.A1(new_n18302_), .A2(new_n18307_), .ZN(new_n18308_));
  NOR2_X1    g18244(.A1(new_n18302_), .A2(new_n18307_), .ZN(new_n18309_));
  AOI21_X1   g18245(.A1(new_n18299_), .A2(new_n18308_), .B(new_n18309_), .ZN(new_n18310_));
  INV_X1     g18246(.I(new_n17914_), .ZN(new_n18311_));
  XOR2_X1    g18247(.A1(new_n17904_), .A2(new_n16299_), .Z(new_n18312_));
  NOR2_X1    g18248(.A1(new_n18312_), .A2(new_n18311_), .ZN(new_n18313_));
  INV_X1     g18249(.I(new_n17915_), .ZN(new_n18314_));
  AOI21_X1   g18250(.A1(new_n18314_), .A2(new_n17905_), .B(new_n17914_), .ZN(new_n18315_));
  NOR2_X1    g18251(.A1(new_n18313_), .A2(new_n18315_), .ZN(new_n18316_));
  AOI22_X1   g18252(.A1(new_n10839_), .A2(new_n7530_), .B1(new_n12936_), .B2(new_n6789_), .ZN(new_n18317_));
  AOI21_X1   g18253(.A1(new_n6784_), .A2(new_n9479_), .B(new_n18317_), .ZN(new_n18318_));
  OR3_X2     g18254(.A1(new_n12975_), .A2(new_n6776_), .A3(new_n18318_), .Z(new_n18319_));
  XOR2_X1    g18255(.A1(new_n18319_), .A2(\a[8] ), .Z(new_n18320_));
  XNOR2_X1   g18256(.A1(new_n18316_), .A2(new_n18320_), .ZN(new_n18321_));
  OR2_X2     g18257(.A1(new_n18321_), .A2(new_n18310_), .Z(new_n18322_));
  NOR2_X1    g18258(.A1(new_n18316_), .A2(new_n18320_), .ZN(new_n18323_));
  AND2_X2    g18259(.A1(new_n18316_), .A2(new_n18320_), .Z(new_n18324_));
  OAI21_X1   g18260(.A1(new_n18324_), .A2(new_n18323_), .B(new_n18310_), .ZN(new_n18325_));
  NAND2_X1   g18261(.A1(new_n18322_), .A2(new_n18325_), .ZN(new_n18326_));
  INV_X1     g18262(.I(new_n18326_), .ZN(new_n18327_));
  OAI22_X1   g18263(.A1(new_n10861_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n10853_), .ZN(new_n18328_));
  NAND2_X1   g18264(.A1(new_n8785_), .A2(new_n6838_), .ZN(new_n18329_));
  AOI21_X1   g18265(.A1(new_n18329_), .A2(new_n18328_), .B(new_n6836_), .ZN(new_n18330_));
  NAND2_X1   g18266(.A1(new_n13592_), .A2(new_n18330_), .ZN(new_n18331_));
  XOR2_X1    g18267(.A1(new_n18331_), .A2(new_n65_), .Z(new_n18332_));
  NAND2_X1   g18268(.A1(new_n18327_), .A2(new_n18332_), .ZN(new_n18333_));
  INV_X1     g18269(.I(new_n18333_), .ZN(new_n18334_));
  XOR2_X1    g18270(.A1(new_n17921_), .A2(new_n17917_), .Z(new_n18335_));
  NAND2_X1   g18271(.A1(new_n17926_), .A2(new_n17922_), .ZN(new_n18336_));
  MUX2_X1    g18272(.I0(new_n18336_), .I1(new_n18335_), .S(new_n17916_), .Z(new_n18337_));
  OAI22_X1   g18273(.A1(new_n9478_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n10846_), .ZN(new_n18338_));
  NAND2_X1   g18274(.A1(new_n10854_), .A2(new_n6784_), .ZN(new_n18339_));
  AOI21_X1   g18275(.A1(new_n18338_), .A2(new_n18339_), .B(new_n6776_), .ZN(new_n18340_));
  NAND2_X1   g18276(.A1(new_n13016_), .A2(new_n18340_), .ZN(new_n18341_));
  XOR2_X1    g18277(.A1(new_n18341_), .A2(new_n4009_), .Z(new_n18342_));
  XOR2_X1    g18278(.A1(new_n18337_), .A2(new_n18342_), .Z(new_n18343_));
  NOR2_X1    g18279(.A1(new_n18316_), .A2(new_n18310_), .ZN(new_n18344_));
  INV_X1     g18280(.I(new_n18344_), .ZN(new_n18345_));
  NOR2_X1    g18281(.A1(new_n18343_), .A2(new_n18345_), .ZN(new_n18346_));
  XNOR2_X1   g18282(.A1(new_n18337_), .A2(new_n18342_), .ZN(new_n18347_));
  NOR2_X1    g18283(.A1(new_n18347_), .A2(new_n18344_), .ZN(new_n18348_));
  XNOR2_X1   g18284(.A1(new_n18316_), .A2(new_n18310_), .ZN(new_n18349_));
  NOR2_X1    g18285(.A1(new_n18349_), .A2(new_n18320_), .ZN(new_n18350_));
  INV_X1     g18286(.I(new_n18350_), .ZN(new_n18351_));
  NOR3_X1    g18287(.A1(new_n18348_), .A2(new_n18346_), .A3(new_n18351_), .ZN(new_n18352_));
  NAND2_X1   g18288(.A1(new_n18347_), .A2(new_n18344_), .ZN(new_n18353_));
  NAND2_X1   g18289(.A1(new_n18343_), .A2(new_n18345_), .ZN(new_n18354_));
  AOI21_X1   g18290(.A1(new_n18353_), .A2(new_n18354_), .B(new_n18350_), .ZN(new_n18355_));
  OAI22_X1   g18291(.A1(new_n8784_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n10861_), .ZN(new_n18356_));
  NAND2_X1   g18292(.A1(new_n8779_), .A2(new_n6838_), .ZN(new_n18357_));
  AOI21_X1   g18293(.A1(new_n18357_), .A2(new_n18356_), .B(new_n6836_), .ZN(new_n18358_));
  NAND2_X1   g18294(.A1(new_n12814_), .A2(new_n18358_), .ZN(new_n18359_));
  XOR2_X1    g18295(.A1(new_n18359_), .A2(\a[5] ), .Z(new_n18360_));
  OAI21_X1   g18296(.A1(new_n18352_), .A2(new_n18355_), .B(new_n18360_), .ZN(new_n18361_));
  NOR3_X1    g18297(.A1(new_n18352_), .A2(new_n18355_), .A3(new_n18360_), .ZN(new_n18362_));
  AOI21_X1   g18298(.A1(new_n18334_), .A2(new_n18361_), .B(new_n18362_), .ZN(new_n18363_));
  AOI22_X1   g18299(.A1(new_n8779_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n8785_), .ZN(new_n18364_));
  NOR2_X1    g18300(.A1(new_n10871_), .A2(new_n6839_), .ZN(new_n18365_));
  OAI21_X1   g18301(.A1(new_n18365_), .A2(new_n18364_), .B(new_n6835_), .ZN(new_n18366_));
  NOR2_X1    g18302(.A1(new_n11794_), .A2(new_n18366_), .ZN(new_n18367_));
  XOR2_X1    g18303(.A1(new_n18367_), .A2(new_n65_), .Z(new_n18368_));
  NOR2_X1    g18304(.A1(new_n17927_), .A2(new_n17933_), .ZN(new_n18369_));
  NAND2_X1   g18305(.A1(new_n17927_), .A2(new_n17933_), .ZN(new_n18370_));
  INV_X1     g18306(.I(new_n18370_), .ZN(new_n18371_));
  OAI21_X1   g18307(.A1(new_n18371_), .A2(new_n18369_), .B(new_n16301_), .ZN(new_n18372_));
  INV_X1     g18308(.I(new_n18369_), .ZN(new_n18373_));
  NAND3_X1   g18309(.A1(new_n18373_), .A2(new_n17935_), .A3(new_n18370_), .ZN(new_n18374_));
  AOI21_X1   g18310(.A1(new_n18372_), .A2(new_n18374_), .B(new_n16294_), .ZN(new_n18375_));
  AOI21_X1   g18311(.A1(new_n18373_), .A2(new_n18370_), .B(new_n17935_), .ZN(new_n18376_));
  NOR3_X1    g18312(.A1(new_n18371_), .A2(new_n16301_), .A3(new_n18369_), .ZN(new_n18377_));
  NOR3_X1    g18313(.A1(new_n18376_), .A2(new_n18377_), .A3(new_n16293_), .ZN(new_n18378_));
  NOR2_X1    g18314(.A1(new_n18375_), .A2(new_n18378_), .ZN(new_n18379_));
  NOR2_X1    g18315(.A1(new_n18324_), .A2(new_n18310_), .ZN(new_n18380_));
  INV_X1     g18316(.I(new_n18380_), .ZN(new_n18381_));
  NAND2_X1   g18317(.A1(new_n18335_), .A2(new_n17916_), .ZN(new_n18382_));
  INV_X1     g18318(.I(new_n18336_), .ZN(new_n18383_));
  OR2_X2     g18319(.A1(new_n18383_), .A2(new_n17916_), .Z(new_n18384_));
  AOI21_X1   g18320(.A1(new_n18384_), .A2(new_n18382_), .B(new_n18342_), .ZN(new_n18385_));
  NOR3_X1    g18321(.A1(new_n18343_), .A2(new_n18323_), .A3(new_n18385_), .ZN(new_n18386_));
  OAI22_X1   g18322(.A1(new_n9478_), .A2(new_n6783_), .B1(new_n6788_), .B2(new_n10853_), .ZN(new_n18387_));
  NAND2_X1   g18323(.A1(new_n10862_), .A2(new_n6784_), .ZN(new_n18388_));
  AOI21_X1   g18324(.A1(new_n18387_), .A2(new_n18388_), .B(new_n6776_), .ZN(new_n18389_));
  NAND2_X1   g18325(.A1(new_n13484_), .A2(new_n18389_), .ZN(new_n18390_));
  XOR2_X1    g18326(.A1(new_n18390_), .A2(\a[8] ), .Z(new_n18391_));
  INV_X1     g18327(.I(new_n18391_), .ZN(new_n18392_));
  AOI21_X1   g18328(.A1(new_n18386_), .A2(new_n18381_), .B(new_n18392_), .ZN(new_n18393_));
  NOR2_X1    g18329(.A1(new_n18385_), .A2(new_n18323_), .ZN(new_n18394_));
  NAND2_X1   g18330(.A1(new_n18347_), .A2(new_n18394_), .ZN(new_n18395_));
  NOR3_X1    g18331(.A1(new_n18395_), .A2(new_n18380_), .A3(new_n18391_), .ZN(new_n18396_));
  OAI21_X1   g18332(.A1(new_n18393_), .A2(new_n18396_), .B(new_n18379_), .ZN(new_n18397_));
  OR2_X2     g18333(.A1(new_n18375_), .A2(new_n18378_), .Z(new_n18398_));
  OAI21_X1   g18334(.A1(new_n18395_), .A2(new_n18380_), .B(new_n18391_), .ZN(new_n18399_));
  NAND3_X1   g18335(.A1(new_n18386_), .A2(new_n18381_), .A3(new_n18392_), .ZN(new_n18400_));
  NAND3_X1   g18336(.A1(new_n18400_), .A2(new_n18399_), .A3(new_n18398_), .ZN(new_n18401_));
  NAND3_X1   g18337(.A1(new_n18397_), .A2(new_n18401_), .A3(new_n18368_), .ZN(new_n18402_));
  INV_X1     g18338(.I(new_n18368_), .ZN(new_n18403_));
  AOI21_X1   g18339(.A1(new_n18400_), .A2(new_n18399_), .B(new_n18398_), .ZN(new_n18404_));
  NOR3_X1    g18340(.A1(new_n18393_), .A2(new_n18396_), .A3(new_n18379_), .ZN(new_n18405_));
  OAI21_X1   g18341(.A1(new_n18404_), .A2(new_n18405_), .B(new_n18403_), .ZN(new_n18406_));
  NAND3_X1   g18342(.A1(new_n18363_), .A2(new_n18406_), .A3(new_n18402_), .ZN(new_n18407_));
  NAND2_X1   g18343(.A1(new_n18248_), .A2(new_n18253_), .ZN(new_n18408_));
  INV_X1     g18344(.I(new_n18054_), .ZN(new_n18409_));
  XOR2_X1    g18345(.A1(new_n18049_), .A2(new_n18409_), .Z(new_n18410_));
  INV_X1     g18346(.I(new_n18253_), .ZN(new_n18411_));
  NAND2_X1   g18347(.A1(new_n18410_), .A2(new_n18411_), .ZN(new_n18412_));
  NOR3_X1    g18348(.A1(new_n18404_), .A2(new_n18405_), .A3(new_n18403_), .ZN(new_n18413_));
  AOI21_X1   g18349(.A1(new_n18408_), .A2(new_n18412_), .B(new_n18413_), .ZN(new_n18414_));
  AOI21_X1   g18350(.A1(new_n18414_), .A2(new_n18407_), .B(new_n18254_), .ZN(new_n18415_));
  INV_X1     g18351(.I(new_n18055_), .ZN(new_n18416_));
  NOR2_X1    g18352(.A1(new_n17954_), .A2(new_n18059_), .ZN(new_n18417_));
  AOI21_X1   g18353(.A1(new_n17954_), .A2(new_n18056_), .B(new_n18417_), .ZN(new_n18418_));
  NAND2_X1   g18354(.A1(new_n18418_), .A2(new_n18065_), .ZN(new_n18419_));
  INV_X1     g18355(.I(new_n18065_), .ZN(new_n18420_));
  NAND2_X1   g18356(.A1(new_n18060_), .A2(new_n18420_), .ZN(new_n18421_));
  AOI21_X1   g18357(.A1(new_n18419_), .A2(new_n18421_), .B(new_n18416_), .ZN(new_n18422_));
  NAND2_X1   g18358(.A1(new_n18418_), .A2(new_n18420_), .ZN(new_n18423_));
  AOI21_X1   g18359(.A1(new_n18423_), .A2(new_n18066_), .B(new_n18055_), .ZN(new_n18424_));
  AOI22_X1   g18360(.A1(new_n10886_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n10872_), .ZN(new_n18425_));
  NOR2_X1    g18361(.A1(new_n10892_), .A2(new_n6839_), .ZN(new_n18426_));
  OAI21_X1   g18362(.A1(new_n18425_), .A2(new_n18426_), .B(new_n6835_), .ZN(new_n18427_));
  NOR2_X1    g18363(.A1(new_n12776_), .A2(new_n18427_), .ZN(new_n18428_));
  XOR2_X1    g18364(.A1(new_n18428_), .A2(new_n65_), .Z(new_n18429_));
  INV_X1     g18365(.I(new_n18429_), .ZN(new_n18430_));
  NOR3_X1    g18366(.A1(new_n18422_), .A2(new_n18424_), .A3(new_n18430_), .ZN(new_n18431_));
  NOR2_X1    g18367(.A1(new_n18060_), .A2(new_n18420_), .ZN(new_n18432_));
  NOR2_X1    g18368(.A1(new_n18418_), .A2(new_n18065_), .ZN(new_n18433_));
  OAI21_X1   g18369(.A1(new_n18433_), .A2(new_n18432_), .B(new_n18055_), .ZN(new_n18434_));
  INV_X1     g18370(.I(new_n18066_), .ZN(new_n18435_));
  OAI21_X1   g18371(.A1(new_n18435_), .A2(new_n18067_), .B(new_n18416_), .ZN(new_n18436_));
  AOI21_X1   g18372(.A1(new_n18436_), .A2(new_n18434_), .B(new_n18429_), .ZN(new_n18437_));
  NOR2_X1    g18373(.A1(new_n18437_), .A2(new_n18431_), .ZN(new_n18438_));
  NOR2_X1    g18374(.A1(new_n18415_), .A2(new_n18438_), .ZN(new_n18439_));
  NAND3_X1   g18375(.A1(new_n18353_), .A2(new_n18354_), .A3(new_n18350_), .ZN(new_n18440_));
  OAI21_X1   g18376(.A1(new_n18348_), .A2(new_n18346_), .B(new_n18351_), .ZN(new_n18441_));
  INV_X1     g18377(.I(new_n18360_), .ZN(new_n18442_));
  AOI21_X1   g18378(.A1(new_n18441_), .A2(new_n18440_), .B(new_n18442_), .ZN(new_n18443_));
  NAND3_X1   g18379(.A1(new_n18441_), .A2(new_n18440_), .A3(new_n18442_), .ZN(new_n18444_));
  OAI21_X1   g18380(.A1(new_n18333_), .A2(new_n18443_), .B(new_n18444_), .ZN(new_n18445_));
  AOI21_X1   g18381(.A1(new_n18397_), .A2(new_n18401_), .B(new_n18368_), .ZN(new_n18446_));
  NOR3_X1    g18382(.A1(new_n18445_), .A2(new_n18446_), .A3(new_n18413_), .ZN(new_n18447_));
  NOR2_X1    g18383(.A1(new_n18410_), .A2(new_n18411_), .ZN(new_n18448_));
  NOR2_X1    g18384(.A1(new_n18248_), .A2(new_n18253_), .ZN(new_n18449_));
  OAI21_X1   g18385(.A1(new_n18448_), .A2(new_n18449_), .B(new_n18402_), .ZN(new_n18450_));
  OAI22_X1   g18386(.A1(new_n18450_), .A2(new_n18447_), .B1(new_n18248_), .B2(new_n18253_), .ZN(new_n18451_));
  AOI21_X1   g18387(.A1(new_n18436_), .A2(new_n18434_), .B(new_n18430_), .ZN(new_n18452_));
  NOR3_X1    g18388(.A1(new_n18422_), .A2(new_n18424_), .A3(new_n18429_), .ZN(new_n18453_));
  NOR2_X1    g18389(.A1(new_n18452_), .A2(new_n18453_), .ZN(new_n18454_));
  NOR2_X1    g18390(.A1(new_n18451_), .A2(new_n18454_), .ZN(new_n18455_));
  NOR3_X1    g18391(.A1(new_n18455_), .A2(new_n18439_), .A3(new_n18246_), .ZN(new_n18456_));
  NOR2_X1    g18392(.A1(new_n18450_), .A2(new_n18447_), .ZN(new_n18457_));
  OAI22_X1   g18393(.A1(new_n18457_), .A2(new_n18254_), .B1(new_n18431_), .B2(new_n18437_), .ZN(new_n18458_));
  OAI21_X1   g18394(.A1(new_n18422_), .A2(new_n18424_), .B(new_n18429_), .ZN(new_n18459_));
  NAND3_X1   g18395(.A1(new_n18436_), .A2(new_n18434_), .A3(new_n18430_), .ZN(new_n18460_));
  NAND2_X1   g18396(.A1(new_n18460_), .A2(new_n18459_), .ZN(new_n18461_));
  NAND2_X1   g18397(.A1(new_n18415_), .A2(new_n18461_), .ZN(new_n18462_));
  AOI21_X1   g18398(.A1(new_n18458_), .A2(new_n18462_), .B(new_n18247_), .ZN(new_n18463_));
  NOR2_X1    g18399(.A1(new_n18456_), .A2(new_n18463_), .ZN(new_n18464_));
  NOR2_X1    g18400(.A1(new_n18464_), .A2(new_n18247_), .ZN(new_n18465_));
  NAND2_X1   g18401(.A1(new_n10889_), .A2(new_n9488_), .ZN(new_n18466_));
  NAND2_X1   g18402(.A1(new_n10886_), .A2(new_n9503_), .ZN(new_n18467_));
  AOI21_X1   g18403(.A1(new_n10872_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n18468_));
  NAND4_X1   g18404(.A1(new_n12776_), .A2(new_n18466_), .A3(new_n18467_), .A4(new_n18468_), .ZN(new_n18469_));
  XOR2_X1    g18405(.A1(new_n18469_), .A2(\a[2] ), .Z(new_n18470_));
  NAND2_X1   g18406(.A1(new_n10886_), .A2(new_n9488_), .ZN(new_n18471_));
  NAND2_X1   g18407(.A1(new_n10872_), .A2(new_n9503_), .ZN(new_n18472_));
  AOI21_X1   g18408(.A1(new_n8779_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n18473_));
  NAND4_X1   g18409(.A1(new_n13103_), .A2(new_n18471_), .A3(new_n18472_), .A4(new_n18473_), .ZN(new_n18474_));
  XOR2_X1    g18410(.A1(new_n18474_), .A2(\a[2] ), .Z(new_n18475_));
  INV_X1     g18411(.I(new_n18475_), .ZN(new_n18476_));
  NAND2_X1   g18412(.A1(new_n10872_), .A2(new_n9488_), .ZN(new_n18477_));
  NAND2_X1   g18413(.A1(new_n8779_), .A2(new_n9503_), .ZN(new_n18478_));
  AOI21_X1   g18414(.A1(new_n8785_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n18479_));
  NAND4_X1   g18415(.A1(new_n11794_), .A2(new_n18477_), .A3(new_n18478_), .A4(new_n18479_), .ZN(new_n18480_));
  XOR2_X1    g18416(.A1(new_n18480_), .A2(new_n4387_), .Z(new_n18481_));
  NOR3_X1    g18417(.A1(new_n13065_), .A2(new_n9482_), .A3(new_n13062_), .ZN(new_n18482_));
  AOI22_X1   g18418(.A1(new_n10862_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n10854_), .ZN(new_n18483_));
  NOR2_X1    g18419(.A1(new_n8784_), .A2(new_n9489_), .ZN(new_n18484_));
  NOR2_X1    g18420(.A1(new_n18483_), .A2(new_n18484_), .ZN(new_n18485_));
  INV_X1     g18421(.I(new_n18485_), .ZN(new_n18486_));
  NOR3_X1    g18422(.A1(new_n18482_), .A2(new_n4387_), .A3(new_n18486_), .ZN(new_n18487_));
  OAI21_X1   g18423(.A1(new_n10855_), .A2(new_n10850_), .B(new_n10861_), .ZN(new_n18488_));
  NAND3_X1   g18424(.A1(new_n13059_), .A2(new_n13010_), .A3(new_n10862_), .ZN(new_n18489_));
  NAND4_X1   g18425(.A1(new_n13063_), .A2(new_n18488_), .A3(new_n8784_), .A4(new_n18489_), .ZN(new_n18490_));
  NAND2_X1   g18426(.A1(new_n18488_), .A2(new_n18489_), .ZN(new_n18491_));
  OAI21_X1   g18427(.A1(new_n18491_), .A2(new_n13058_), .B(new_n8785_), .ZN(new_n18492_));
  NAND3_X1   g18428(.A1(new_n18492_), .A2(new_n18490_), .A3(new_n6922_), .ZN(new_n18493_));
  AOI21_X1   g18429(.A1(new_n18493_), .A2(new_n18485_), .B(\a[2] ), .ZN(new_n18494_));
  NOR2_X1    g18430(.A1(new_n18487_), .A2(new_n18494_), .ZN(new_n18495_));
  OAI22_X1   g18431(.A1(new_n10775_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n10777_), .ZN(new_n18496_));
  NAND2_X1   g18432(.A1(new_n9529_), .A2(new_n6838_), .ZN(new_n18497_));
  AOI21_X1   g18433(.A1(new_n18496_), .A2(new_n18497_), .B(new_n6836_), .ZN(new_n18498_));
  NAND3_X1   g18434(.A1(new_n12883_), .A2(new_n65_), .A3(new_n18498_), .ZN(new_n18499_));
  INV_X1     g18435(.I(new_n18499_), .ZN(new_n18500_));
  AOI21_X1   g18436(.A1(new_n12883_), .A2(new_n18498_), .B(new_n65_), .ZN(new_n18501_));
  OAI21_X1   g18437(.A1(new_n18500_), .A2(new_n18501_), .B(new_n18271_), .ZN(new_n18502_));
  NAND2_X1   g18438(.A1(new_n12823_), .A2(new_n8799_), .ZN(new_n18503_));
  NAND2_X1   g18439(.A1(new_n10794_), .A2(new_n6846_), .ZN(new_n18504_));
  AOI22_X1   g18440(.A1(new_n18504_), .A2(new_n18503_), .B1(new_n6838_), .B2(new_n10800_), .ZN(new_n18505_));
  NOR3_X1    g18441(.A1(new_n14787_), .A2(new_n6836_), .A3(new_n18505_), .ZN(new_n18506_));
  NOR2_X1    g18442(.A1(new_n6833_), .A2(new_n6834_), .ZN(new_n18507_));
  OAI21_X1   g18443(.A1(new_n12826_), .A2(new_n6843_), .B(new_n18507_), .ZN(new_n18508_));
  NOR2_X1    g18444(.A1(new_n12847_), .A2(new_n18508_), .ZN(new_n18509_));
  INV_X1     g18445(.I(new_n18509_), .ZN(new_n18510_));
  NOR2_X1    g18446(.A1(new_n12826_), .A2(new_n6833_), .ZN(new_n18511_));
  NOR4_X1    g18447(.A1(new_n18506_), .A2(new_n18510_), .A3(new_n65_), .A4(new_n18511_), .ZN(new_n18512_));
  NOR3_X1    g18448(.A1(new_n18500_), .A2(new_n18501_), .A3(new_n18271_), .ZN(new_n18513_));
  OAI21_X1   g18449(.A1(new_n18512_), .A2(new_n18513_), .B(new_n18502_), .ZN(new_n18514_));
  INV_X1     g18450(.I(new_n18268_), .ZN(new_n18515_));
  NAND3_X1   g18451(.A1(new_n14793_), .A2(new_n18515_), .A3(new_n4009_), .ZN(new_n18516_));
  OAI21_X1   g18452(.A1(new_n12847_), .A2(new_n18268_), .B(\a[8] ), .ZN(new_n18517_));
  NOR2_X1    g18453(.A1(new_n18270_), .A2(new_n4009_), .ZN(new_n18518_));
  INV_X1     g18454(.I(new_n18518_), .ZN(new_n18519_));
  NAND3_X1   g18455(.A1(new_n18516_), .A2(new_n18517_), .A3(new_n18519_), .ZN(new_n18520_));
  NAND2_X1   g18456(.A1(new_n14793_), .A2(new_n18515_), .ZN(new_n18521_));
  NAND3_X1   g18457(.A1(new_n18521_), .A2(\a[8] ), .A3(new_n18271_), .ZN(new_n18522_));
  NAND2_X1   g18458(.A1(new_n18520_), .A2(new_n18522_), .ZN(new_n18523_));
  OAI22_X1   g18459(.A1(new_n10798_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n10777_), .ZN(new_n18524_));
  NAND2_X1   g18460(.A1(new_n10839_), .A2(new_n6838_), .ZN(new_n18525_));
  AOI21_X1   g18461(.A1(new_n18525_), .A2(new_n18524_), .B(new_n6836_), .ZN(new_n18526_));
  NAND3_X1   g18462(.A1(new_n12910_), .A2(new_n65_), .A3(new_n18526_), .ZN(new_n18527_));
  OAI21_X1   g18463(.A1(new_n13530_), .A2(new_n13533_), .B(new_n18526_), .ZN(new_n18528_));
  NAND2_X1   g18464(.A1(new_n18528_), .A2(\a[5] ), .ZN(new_n18529_));
  NAND3_X1   g18465(.A1(new_n18527_), .A2(new_n18529_), .A3(new_n18523_), .ZN(new_n18530_));
  NAND2_X1   g18466(.A1(new_n18514_), .A2(new_n18530_), .ZN(new_n18531_));
  NOR3_X1    g18467(.A1(new_n12847_), .A2(new_n18268_), .A3(\a[8] ), .ZN(new_n18532_));
  AOI21_X1   g18468(.A1(new_n14793_), .A2(new_n18515_), .B(new_n4009_), .ZN(new_n18533_));
  NOR3_X1    g18469(.A1(new_n18533_), .A2(new_n18532_), .A3(new_n18518_), .ZN(new_n18534_));
  NOR3_X1    g18470(.A1(new_n18269_), .A2(new_n4009_), .A3(new_n18270_), .ZN(new_n18535_));
  NOR2_X1    g18471(.A1(new_n18534_), .A2(new_n18535_), .ZN(new_n18536_));
  NOR2_X1    g18472(.A1(new_n18528_), .A2(\a[5] ), .ZN(new_n18537_));
  AOI21_X1   g18473(.A1(new_n12910_), .A2(new_n18526_), .B(new_n65_), .ZN(new_n18538_));
  OAI21_X1   g18474(.A1(new_n18538_), .A2(new_n18537_), .B(new_n18536_), .ZN(new_n18539_));
  AOI21_X1   g18475(.A1(new_n18265_), .A2(new_n18264_), .B(\a[8] ), .ZN(new_n18540_));
  INV_X1     g18476(.I(new_n18262_), .ZN(new_n18541_));
  NAND2_X1   g18477(.A1(new_n10794_), .A2(new_n7530_), .ZN(new_n18542_));
  AOI22_X1   g18478(.A1(new_n18542_), .A2(new_n18541_), .B1(new_n6784_), .B2(new_n10800_), .ZN(new_n18543_));
  OAI21_X1   g18479(.A1(new_n14786_), .A2(new_n12828_), .B(new_n6775_), .ZN(new_n18544_));
  NOR3_X1    g18480(.A1(new_n18544_), .A2(new_n4009_), .A3(new_n18543_), .ZN(new_n18545_));
  NOR3_X1    g18481(.A1(new_n18521_), .A2(new_n4009_), .A3(new_n18270_), .ZN(new_n18546_));
  NOR3_X1    g18482(.A1(new_n18540_), .A2(new_n18546_), .A3(new_n18545_), .ZN(new_n18547_));
  NOR4_X1    g18483(.A1(new_n18266_), .A2(new_n4009_), .A3(new_n18521_), .A4(new_n18270_), .ZN(new_n18548_));
  NOR2_X1    g18484(.A1(new_n18547_), .A2(new_n18548_), .ZN(new_n18549_));
  NAND3_X1   g18485(.A1(new_n10802_), .A2(new_n9529_), .A3(new_n10844_), .ZN(new_n18550_));
  NAND2_X1   g18486(.A1(new_n10839_), .A2(new_n10795_), .ZN(new_n18551_));
  AOI21_X1   g18487(.A1(new_n18550_), .A2(new_n18551_), .B(new_n10846_), .ZN(new_n18552_));
  AOI21_X1   g18488(.A1(new_n12943_), .A2(new_n12944_), .B(new_n12936_), .ZN(new_n18553_));
  AOI22_X1   g18489(.A1(new_n10839_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n9529_), .ZN(new_n18554_));
  NOR2_X1    g18490(.A1(new_n10846_), .A2(new_n6839_), .ZN(new_n18555_));
  OAI21_X1   g18491(.A1(new_n18554_), .A2(new_n18555_), .B(new_n6835_), .ZN(new_n18556_));
  NOR4_X1    g18492(.A1(new_n18552_), .A2(new_n18553_), .A3(new_n18556_), .A4(\a[5] ), .ZN(new_n18557_));
  NOR3_X1    g18493(.A1(new_n18552_), .A2(new_n18553_), .A3(new_n18556_), .ZN(new_n18558_));
  NOR2_X1    g18494(.A1(new_n18558_), .A2(new_n65_), .ZN(new_n18559_));
  NOR3_X1    g18495(.A1(new_n18549_), .A2(new_n18559_), .A3(new_n18557_), .ZN(new_n18560_));
  AOI21_X1   g18496(.A1(new_n18531_), .A2(new_n18539_), .B(new_n18560_), .ZN(new_n18561_));
  OAI21_X1   g18497(.A1(new_n18544_), .A2(new_n18543_), .B(new_n4009_), .ZN(new_n18562_));
  NAND3_X1   g18498(.A1(new_n18265_), .A2(\a[8] ), .A3(new_n18264_), .ZN(new_n18563_));
  NAND3_X1   g18499(.A1(new_n18269_), .A2(\a[8] ), .A3(new_n18271_), .ZN(new_n18564_));
  NAND3_X1   g18500(.A1(new_n18562_), .A2(new_n18563_), .A3(new_n18564_), .ZN(new_n18565_));
  NOR2_X1    g18501(.A1(new_n18544_), .A2(new_n18543_), .ZN(new_n18566_));
  NAND4_X1   g18502(.A1(new_n18566_), .A2(\a[8] ), .A3(new_n18269_), .A4(new_n18271_), .ZN(new_n18567_));
  NAND2_X1   g18503(.A1(new_n18565_), .A2(new_n18567_), .ZN(new_n18568_));
  INV_X1     g18504(.I(new_n18557_), .ZN(new_n18569_));
  OAI21_X1   g18505(.A1(new_n12946_), .A2(new_n18556_), .B(\a[5] ), .ZN(new_n18570_));
  AOI21_X1   g18506(.A1(new_n18570_), .A2(new_n18569_), .B(new_n18568_), .ZN(new_n18571_));
  INV_X1     g18507(.I(new_n17913_), .ZN(new_n18572_));
  NAND3_X1   g18508(.A1(new_n18260_), .A2(new_n18258_), .A3(new_n18572_), .ZN(new_n18573_));
  INV_X1     g18509(.I(new_n18258_), .ZN(new_n18574_));
  AOI21_X1   g18510(.A1(new_n12883_), .A2(new_n18257_), .B(new_n4009_), .ZN(new_n18575_));
  OAI21_X1   g18511(.A1(new_n18574_), .A2(new_n18575_), .B(new_n17913_), .ZN(new_n18576_));
  AOI21_X1   g18512(.A1(new_n18576_), .A2(new_n18573_), .B(new_n18272_), .ZN(new_n18577_));
  OAI21_X1   g18513(.A1(new_n18574_), .A2(new_n18575_), .B(new_n18572_), .ZN(new_n18578_));
  NOR3_X1    g18514(.A1(new_n18540_), .A2(new_n18545_), .A3(new_n18564_), .ZN(new_n18579_));
  AOI21_X1   g18515(.A1(new_n18578_), .A2(new_n18273_), .B(new_n18579_), .ZN(new_n18580_));
  NOR2_X1    g18516(.A1(new_n18580_), .A2(new_n18577_), .ZN(new_n18581_));
  OAI22_X1   g18517(.A1(new_n10844_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n10846_), .ZN(new_n18582_));
  NOR2_X1    g18518(.A1(new_n9478_), .A2(new_n6839_), .ZN(new_n18583_));
  INV_X1     g18519(.I(new_n18583_), .ZN(new_n18584_));
  AOI21_X1   g18520(.A1(new_n18584_), .A2(new_n18582_), .B(new_n6836_), .ZN(new_n18585_));
  INV_X1     g18521(.I(new_n18585_), .ZN(new_n18586_));
  NOR4_X1    g18522(.A1(new_n13565_), .A2(\a[5] ), .A3(new_n13563_), .A4(new_n18586_), .ZN(new_n18587_));
  AOI21_X1   g18523(.A1(new_n13566_), .A2(new_n18585_), .B(new_n65_), .ZN(new_n18588_));
  NOR3_X1    g18524(.A1(new_n18588_), .A2(new_n18581_), .A3(new_n18587_), .ZN(new_n18589_));
  NOR3_X1    g18525(.A1(new_n18574_), .A2(new_n18575_), .A3(new_n17913_), .ZN(new_n18590_));
  AOI21_X1   g18526(.A1(new_n18260_), .A2(new_n18258_), .B(new_n18572_), .ZN(new_n18591_));
  OAI21_X1   g18527(.A1(new_n18590_), .A2(new_n18591_), .B(new_n18579_), .ZN(new_n18592_));
  NOR3_X1    g18528(.A1(new_n18574_), .A2(new_n18575_), .A3(new_n18572_), .ZN(new_n18593_));
  OAI21_X1   g18529(.A1(new_n18593_), .A2(new_n18261_), .B(new_n18272_), .ZN(new_n18594_));
  NAND2_X1   g18530(.A1(new_n18592_), .A2(new_n18594_), .ZN(new_n18595_));
  NAND4_X1   g18531(.A1(new_n12974_), .A2(new_n65_), .A3(new_n12972_), .A4(new_n18585_), .ZN(new_n18596_));
  OAI21_X1   g18532(.A1(new_n12975_), .A2(new_n18586_), .B(\a[5] ), .ZN(new_n18597_));
  AOI21_X1   g18533(.A1(new_n18597_), .A2(new_n18596_), .B(new_n18595_), .ZN(new_n18598_));
  OAI22_X1   g18534(.A1(new_n18589_), .A2(new_n18598_), .B1(new_n18561_), .B2(new_n18571_), .ZN(new_n18599_));
  OAI21_X1   g18535(.A1(new_n13502_), .A2(new_n13503_), .B(new_n18498_), .ZN(new_n18600_));
  NAND2_X1   g18536(.A1(new_n18600_), .A2(\a[5] ), .ZN(new_n18601_));
  AOI21_X1   g18537(.A1(new_n18601_), .A2(new_n18499_), .B(new_n18270_), .ZN(new_n18602_));
  INV_X1     g18538(.I(new_n18505_), .ZN(new_n18603_));
  NAND3_X1   g18539(.A1(new_n18603_), .A2(new_n12830_), .A3(new_n6835_), .ZN(new_n18604_));
  INV_X1     g18540(.I(new_n18511_), .ZN(new_n18605_));
  NAND4_X1   g18541(.A1(new_n18604_), .A2(\a[5] ), .A3(new_n18509_), .A4(new_n18605_), .ZN(new_n18606_));
  NAND3_X1   g18542(.A1(new_n18601_), .A2(new_n18499_), .A3(new_n18270_), .ZN(new_n18607_));
  AOI21_X1   g18543(.A1(new_n18606_), .A2(new_n18607_), .B(new_n18602_), .ZN(new_n18608_));
  NOR3_X1    g18544(.A1(new_n18538_), .A2(new_n18537_), .A3(new_n18536_), .ZN(new_n18609_));
  OAI21_X1   g18545(.A1(new_n18608_), .A2(new_n18609_), .B(new_n18539_), .ZN(new_n18610_));
  NAND3_X1   g18546(.A1(new_n18570_), .A2(new_n18568_), .A3(new_n18569_), .ZN(new_n18611_));
  AOI21_X1   g18547(.A1(new_n18610_), .A2(new_n18611_), .B(new_n18571_), .ZN(new_n18612_));
  NOR3_X1    g18548(.A1(new_n18588_), .A2(new_n18595_), .A3(new_n18587_), .ZN(new_n18613_));
  AOI21_X1   g18549(.A1(new_n18597_), .A2(new_n18596_), .B(new_n18581_), .ZN(new_n18614_));
  OAI21_X1   g18550(.A1(new_n18613_), .A2(new_n18614_), .B(new_n18612_), .ZN(new_n18615_));
  NAND2_X1   g18551(.A1(new_n18615_), .A2(new_n18599_), .ZN(new_n18616_));
  NAND2_X1   g18552(.A1(new_n18495_), .A2(new_n18616_), .ZN(new_n18617_));
  INV_X1     g18553(.I(new_n18617_), .ZN(new_n18618_));
  NOR2_X1    g18554(.A1(new_n10853_), .A2(new_n9489_), .ZN(new_n18619_));
  NOR2_X1    g18555(.A1(new_n9478_), .A2(new_n9483_), .ZN(new_n18620_));
  NOR2_X1    g18556(.A1(new_n10846_), .A2(new_n9485_), .ZN(new_n18621_));
  NOR4_X1    g18557(.A1(new_n18620_), .A2(new_n9482_), .A3(new_n18619_), .A4(new_n18621_), .ZN(new_n18622_));
  NAND2_X1   g18558(.A1(new_n13016_), .A2(new_n18622_), .ZN(new_n18623_));
  XOR2_X1    g18559(.A1(new_n18623_), .A2(\a[2] ), .Z(new_n18624_));
  NOR2_X1    g18560(.A1(new_n10844_), .A2(new_n9483_), .ZN(new_n18625_));
  NOR2_X1    g18561(.A1(new_n10798_), .A2(new_n9485_), .ZN(new_n18626_));
  NOR2_X1    g18562(.A1(new_n10846_), .A2(new_n9489_), .ZN(new_n18627_));
  NOR4_X1    g18563(.A1(new_n18625_), .A2(new_n6922_), .A3(new_n18626_), .A4(new_n18627_), .ZN(new_n18628_));
  AOI21_X1   g18564(.A1(new_n12946_), .A2(new_n18628_), .B(new_n4387_), .ZN(new_n18629_));
  OAI21_X1   g18565(.A1(new_n18552_), .A2(new_n18553_), .B(new_n18628_), .ZN(new_n18630_));
  NOR2_X1    g18566(.A1(new_n18630_), .A2(\a[2] ), .ZN(new_n18631_));
  NOR2_X1    g18567(.A1(new_n18629_), .A2(new_n18631_), .ZN(new_n18632_));
  NOR2_X1    g18568(.A1(new_n14787_), .A2(new_n9617_), .ZN(new_n18633_));
  NAND2_X1   g18569(.A1(new_n14793_), .A2(new_n9613_), .ZN(new_n18634_));
  NAND2_X1   g18570(.A1(new_n10794_), .A2(new_n6925_), .ZN(new_n18635_));
  NAND2_X1   g18571(.A1(new_n12823_), .A2(new_n9503_), .ZN(new_n18636_));
  NOR2_X1    g18572(.A1(new_n9489_), .A2(\a[2] ), .ZN(new_n18637_));
  NAND4_X1   g18573(.A1(new_n18635_), .A2(new_n10800_), .A3(new_n18636_), .A4(new_n18637_), .ZN(new_n18638_));
  NOR2_X1    g18574(.A1(new_n10775_), .A2(new_n9623_), .ZN(new_n18639_));
  NOR2_X1    g18575(.A1(new_n6923_), .A2(\a[2] ), .ZN(new_n18640_));
  INV_X1     g18576(.I(new_n18640_), .ZN(new_n18641_));
  NOR3_X1    g18577(.A1(new_n12826_), .A2(new_n18639_), .A3(new_n18641_), .ZN(new_n18642_));
  NAND3_X1   g18578(.A1(new_n18634_), .A2(new_n18638_), .A3(new_n18642_), .ZN(new_n18643_));
  NOR3_X1    g18579(.A1(new_n18643_), .A2(new_n18605_), .A3(new_n18633_), .ZN(new_n18644_));
  AOI21_X1   g18580(.A1(new_n10800_), .A2(new_n9503_), .B(new_n9482_), .ZN(new_n18645_));
  OAI21_X1   g18581(.A1(new_n9489_), .A2(new_n10798_), .B(new_n18645_), .ZN(new_n18646_));
  AOI21_X1   g18582(.A1(new_n6925_), .A2(new_n12823_), .B(new_n18646_), .ZN(new_n18647_));
  NAND2_X1   g18583(.A1(new_n12883_), .A2(new_n18647_), .ZN(new_n18648_));
  XOR2_X1    g18584(.A1(new_n18648_), .A2(new_n4387_), .Z(new_n18649_));
  INV_X1     g18585(.I(new_n18633_), .ZN(new_n18650_));
  NAND2_X1   g18586(.A1(new_n18638_), .A2(new_n18642_), .ZN(new_n18651_));
  AOI21_X1   g18587(.A1(new_n9613_), .A2(new_n14793_), .B(new_n18651_), .ZN(new_n18652_));
  AOI21_X1   g18588(.A1(new_n18652_), .A2(new_n18650_), .B(new_n18511_), .ZN(new_n18653_));
  AOI21_X1   g18589(.A1(new_n18653_), .A2(new_n18649_), .B(new_n18644_), .ZN(new_n18654_));
  OAI22_X1   g18590(.A1(new_n10798_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n10777_), .ZN(new_n18655_));
  NAND2_X1   g18591(.A1(new_n10839_), .A2(new_n9488_), .ZN(new_n18656_));
  AOI21_X1   g18592(.A1(new_n18656_), .A2(new_n18655_), .B(new_n9482_), .ZN(new_n18657_));
  INV_X1     g18593(.I(new_n18657_), .ZN(new_n18658_));
  NOR3_X1    g18594(.A1(new_n13534_), .A2(\a[2] ), .A3(new_n18658_), .ZN(new_n18659_));
  AOI21_X1   g18595(.A1(new_n12910_), .A2(new_n18657_), .B(new_n4387_), .ZN(new_n18660_));
  NOR2_X1    g18596(.A1(new_n18660_), .A2(new_n18659_), .ZN(new_n18661_));
  NOR2_X1    g18597(.A1(new_n18654_), .A2(new_n18661_), .ZN(new_n18662_));
  NAND3_X1   g18598(.A1(new_n18509_), .A2(\a[5] ), .A3(new_n18605_), .ZN(new_n18663_));
  NOR2_X1    g18599(.A1(new_n18510_), .A2(\a[5] ), .ZN(new_n18664_));
  NOR2_X1    g18600(.A1(new_n18509_), .A2(new_n65_), .ZN(new_n18665_));
  OAI22_X1   g18601(.A1(new_n18664_), .A2(new_n18665_), .B1(new_n65_), .B2(new_n18511_), .ZN(new_n18666_));
  AOI22_X1   g18602(.A1(new_n18654_), .A2(new_n18661_), .B1(new_n18663_), .B2(new_n18666_), .ZN(new_n18667_));
  OAI21_X1   g18603(.A1(new_n18667_), .A2(new_n18662_), .B(new_n18632_), .ZN(new_n18668_));
  NOR3_X1    g18604(.A1(new_n18667_), .A2(new_n18632_), .A3(new_n18662_), .ZN(new_n18669_));
  INV_X1     g18605(.I(new_n18632_), .ZN(new_n18670_));
  NAND3_X1   g18606(.A1(new_n18652_), .A2(new_n18650_), .A3(new_n18511_), .ZN(new_n18671_));
  XOR2_X1    g18607(.A1(new_n18648_), .A2(\a[2] ), .Z(new_n18672_));
  OAI21_X1   g18608(.A1(new_n18643_), .A2(new_n18633_), .B(new_n18605_), .ZN(new_n18673_));
  OAI21_X1   g18609(.A1(new_n18672_), .A2(new_n18673_), .B(new_n18671_), .ZN(new_n18674_));
  INV_X1     g18610(.I(new_n18661_), .ZN(new_n18675_));
  NAND2_X1   g18611(.A1(new_n18675_), .A2(new_n18674_), .ZN(new_n18676_));
  NAND2_X1   g18612(.A1(new_n18666_), .A2(new_n18663_), .ZN(new_n18677_));
  OAI21_X1   g18613(.A1(new_n18675_), .A2(new_n18674_), .B(new_n18677_), .ZN(new_n18678_));
  AOI21_X1   g18614(.A1(new_n18678_), .A2(new_n18676_), .B(new_n18670_), .ZN(new_n18679_));
  XOR2_X1    g18615(.A1(new_n18506_), .A2(\a[5] ), .Z(new_n18680_));
  XOR2_X1    g18616(.A1(new_n18680_), .A2(new_n18663_), .Z(new_n18681_));
  OAI21_X1   g18617(.A1(new_n18679_), .A2(new_n18669_), .B(new_n18681_), .ZN(new_n18682_));
  AOI22_X1   g18618(.A1(new_n10839_), .A2(new_n6925_), .B1(new_n12936_), .B2(new_n9503_), .ZN(new_n18683_));
  NOR2_X1    g18619(.A1(new_n9478_), .A2(new_n9489_), .ZN(new_n18684_));
  OAI21_X1   g18620(.A1(new_n18683_), .A2(new_n18684_), .B(new_n6922_), .ZN(new_n18685_));
  NOR3_X1    g18621(.A1(new_n12975_), .A2(\a[2] ), .A3(new_n18685_), .ZN(new_n18686_));
  OAI21_X1   g18622(.A1(new_n12975_), .A2(new_n18685_), .B(\a[2] ), .ZN(new_n18687_));
  INV_X1     g18623(.I(new_n18687_), .ZN(new_n18688_));
  NOR2_X1    g18624(.A1(new_n18688_), .A2(new_n18686_), .ZN(new_n18689_));
  AOI21_X1   g18625(.A1(new_n18682_), .A2(new_n18668_), .B(new_n18689_), .ZN(new_n18690_));
  NAND3_X1   g18626(.A1(new_n18678_), .A2(new_n18676_), .A3(new_n18670_), .ZN(new_n18691_));
  OAI21_X1   g18627(.A1(new_n18667_), .A2(new_n18662_), .B(new_n18632_), .ZN(new_n18692_));
  XNOR2_X1   g18628(.A1(new_n18680_), .A2(new_n18663_), .ZN(new_n18693_));
  AOI22_X1   g18629(.A1(new_n18691_), .A2(new_n18692_), .B1(new_n18670_), .B2(new_n18693_), .ZN(new_n18694_));
  INV_X1     g18630(.I(new_n18689_), .ZN(new_n18695_));
  NOR2_X1    g18631(.A1(new_n18500_), .A2(new_n18501_), .ZN(new_n18696_));
  NOR2_X1    g18632(.A1(new_n18512_), .A2(new_n18270_), .ZN(new_n18697_));
  NOR2_X1    g18633(.A1(new_n18606_), .A2(new_n18271_), .ZN(new_n18698_));
  NOR3_X1    g18634(.A1(new_n18698_), .A2(new_n18697_), .A3(new_n18696_), .ZN(new_n18699_));
  INV_X1     g18635(.I(new_n18696_), .ZN(new_n18700_));
  NOR2_X1    g18636(.A1(new_n18698_), .A2(new_n18697_), .ZN(new_n18701_));
  NOR2_X1    g18637(.A1(new_n18701_), .A2(new_n18700_), .ZN(new_n18702_));
  NOR2_X1    g18638(.A1(new_n18702_), .A2(new_n18699_), .ZN(new_n18703_));
  NOR3_X1    g18639(.A1(new_n18694_), .A2(new_n18695_), .A3(new_n18703_), .ZN(new_n18704_));
  NOR3_X1    g18640(.A1(new_n18704_), .A2(new_n18690_), .A3(new_n18624_), .ZN(new_n18705_));
  NAND2_X1   g18641(.A1(new_n18623_), .A2(\a[2] ), .ZN(new_n18706_));
  NAND3_X1   g18642(.A1(new_n13016_), .A2(new_n4387_), .A3(new_n18622_), .ZN(new_n18707_));
  NAND2_X1   g18643(.A1(new_n18706_), .A2(new_n18707_), .ZN(new_n18708_));
  NAND2_X1   g18644(.A1(new_n18694_), .A2(new_n18695_), .ZN(new_n18709_));
  NOR3_X1    g18645(.A1(new_n18703_), .A2(new_n18686_), .A3(new_n18688_), .ZN(new_n18710_));
  NAND3_X1   g18646(.A1(new_n18682_), .A2(new_n18668_), .A3(new_n18710_), .ZN(new_n18711_));
  AOI21_X1   g18647(.A1(new_n18709_), .A2(new_n18711_), .B(new_n18708_), .ZN(new_n18712_));
  NAND2_X1   g18648(.A1(new_n18527_), .A2(new_n18529_), .ZN(new_n18713_));
  XOR2_X1    g18649(.A1(new_n18713_), .A2(new_n18523_), .Z(new_n18714_));
  NOR2_X1    g18650(.A1(new_n18714_), .A2(new_n18608_), .ZN(new_n18715_));
  AOI21_X1   g18651(.A1(new_n18527_), .A2(new_n18529_), .B(new_n18523_), .ZN(new_n18716_));
  NOR2_X1    g18652(.A1(new_n18716_), .A2(new_n18609_), .ZN(new_n18717_));
  INV_X1     g18653(.I(new_n18717_), .ZN(new_n18718_));
  AOI21_X1   g18654(.A1(new_n18608_), .A2(new_n18718_), .B(new_n18715_), .ZN(new_n18719_));
  OAI21_X1   g18655(.A1(new_n18705_), .A2(new_n18712_), .B(new_n18719_), .ZN(new_n18720_));
  NAND2_X1   g18656(.A1(new_n18709_), .A2(new_n18711_), .ZN(new_n18721_));
  INV_X1     g18657(.I(new_n13035_), .ZN(new_n18722_));
  OAI21_X1   g18658(.A1(new_n18722_), .A2(new_n13033_), .B(new_n10862_), .ZN(new_n18723_));
  NAND3_X1   g18659(.A1(new_n18723_), .A2(new_n6922_), .A3(new_n13039_), .ZN(new_n18724_));
  AOI22_X1   g18660(.A1(new_n9479_), .A2(new_n6925_), .B1(new_n10854_), .B2(new_n9503_), .ZN(new_n18725_));
  AOI21_X1   g18661(.A1(new_n9488_), .A2(new_n10862_), .B(new_n18725_), .ZN(new_n18726_));
  NAND3_X1   g18662(.A1(new_n18724_), .A2(\a[2] ), .A3(new_n18726_), .ZN(new_n18727_));
  NOR3_X1    g18663(.A1(new_n13040_), .A2(new_n13036_), .A3(new_n9482_), .ZN(new_n18728_));
  INV_X1     g18664(.I(new_n18726_), .ZN(new_n18729_));
  OAI21_X1   g18665(.A1(new_n18728_), .A2(new_n18729_), .B(new_n4387_), .ZN(new_n18730_));
  NAND2_X1   g18666(.A1(new_n18730_), .A2(new_n18727_), .ZN(new_n18731_));
  AOI21_X1   g18667(.A1(new_n18514_), .A2(new_n18530_), .B(new_n18716_), .ZN(new_n18732_));
  NAND3_X1   g18668(.A1(new_n18570_), .A2(new_n18549_), .A3(new_n18569_), .ZN(new_n18733_));
  NAND2_X1   g18669(.A1(new_n18570_), .A2(new_n18569_), .ZN(new_n18734_));
  NAND2_X1   g18670(.A1(new_n18734_), .A2(new_n18568_), .ZN(new_n18735_));
  AOI21_X1   g18671(.A1(new_n18735_), .A2(new_n18733_), .B(new_n18732_), .ZN(new_n18736_));
  OAI21_X1   g18672(.A1(new_n18557_), .A2(new_n18559_), .B(new_n18549_), .ZN(new_n18737_));
  AOI21_X1   g18673(.A1(new_n18611_), .A2(new_n18737_), .B(new_n18610_), .ZN(new_n18738_));
  NOR2_X1    g18674(.A1(new_n18736_), .A2(new_n18738_), .ZN(new_n18739_));
  NAND2_X1   g18675(.A1(new_n18731_), .A2(new_n18739_), .ZN(new_n18740_));
  NOR3_X1    g18676(.A1(new_n18728_), .A2(new_n4387_), .A3(new_n18729_), .ZN(new_n18741_));
  AOI21_X1   g18677(.A1(new_n18724_), .A2(new_n18726_), .B(\a[2] ), .ZN(new_n18742_));
  NOR2_X1    g18678(.A1(new_n18741_), .A2(new_n18742_), .ZN(new_n18743_));
  AND2_X2    g18679(.A1(new_n18735_), .A2(new_n18733_), .Z(new_n18744_));
  OAI21_X1   g18680(.A1(new_n18560_), .A2(new_n18571_), .B(new_n18732_), .ZN(new_n18745_));
  OAI21_X1   g18681(.A1(new_n18744_), .A2(new_n18732_), .B(new_n18745_), .ZN(new_n18746_));
  NAND2_X1   g18682(.A1(new_n18746_), .A2(new_n18743_), .ZN(new_n18747_));
  AOI22_X1   g18683(.A1(new_n18721_), .A2(new_n18624_), .B1(new_n18740_), .B2(new_n18747_), .ZN(new_n18748_));
  NAND3_X1   g18684(.A1(new_n18493_), .A2(\a[2] ), .A3(new_n18485_), .ZN(new_n18749_));
  OAI21_X1   g18685(.A1(new_n18482_), .A2(new_n18486_), .B(new_n4387_), .ZN(new_n18750_));
  AOI21_X1   g18686(.A1(new_n18749_), .A2(new_n18750_), .B(new_n18616_), .ZN(new_n18751_));
  NOR2_X1    g18687(.A1(new_n18609_), .A2(new_n18608_), .ZN(new_n18752_));
  OAI21_X1   g18688(.A1(new_n18752_), .A2(new_n18716_), .B(new_n18611_), .ZN(new_n18753_));
  NAND3_X1   g18689(.A1(new_n18597_), .A2(new_n18595_), .A3(new_n18596_), .ZN(new_n18754_));
  OAI21_X1   g18690(.A1(new_n18588_), .A2(new_n18587_), .B(new_n18581_), .ZN(new_n18755_));
  AOI22_X1   g18691(.A1(new_n18755_), .A2(new_n18754_), .B1(new_n18753_), .B2(new_n18737_), .ZN(new_n18756_));
  OAI21_X1   g18692(.A1(new_n18732_), .A2(new_n18560_), .B(new_n18737_), .ZN(new_n18757_));
  NAND3_X1   g18693(.A1(new_n18597_), .A2(new_n18581_), .A3(new_n18596_), .ZN(new_n18758_));
  OAI21_X1   g18694(.A1(new_n18588_), .A2(new_n18587_), .B(new_n18595_), .ZN(new_n18759_));
  AOI21_X1   g18695(.A1(new_n18758_), .A2(new_n18759_), .B(new_n18757_), .ZN(new_n18760_));
  NOR2_X1    g18696(.A1(new_n18760_), .A2(new_n18756_), .ZN(new_n18761_));
  NOR3_X1    g18697(.A1(new_n18761_), .A2(new_n18487_), .A3(new_n18494_), .ZN(new_n18762_));
  NOR2_X1    g18698(.A1(new_n18731_), .A2(new_n18739_), .ZN(new_n18763_));
  INV_X1     g18699(.I(new_n18763_), .ZN(new_n18764_));
  OAI21_X1   g18700(.A1(new_n18751_), .A2(new_n18762_), .B(new_n18764_), .ZN(new_n18765_));
  AOI21_X1   g18701(.A1(new_n18720_), .A2(new_n18748_), .B(new_n18765_), .ZN(new_n18766_));
  OAI22_X1   g18702(.A1(new_n8784_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n10861_), .ZN(new_n18767_));
  NAND2_X1   g18703(.A1(new_n8779_), .A2(new_n9488_), .ZN(new_n18768_));
  AOI21_X1   g18704(.A1(new_n18768_), .A2(new_n18767_), .B(new_n9482_), .ZN(new_n18769_));
  NAND3_X1   g18705(.A1(new_n12814_), .A2(new_n4387_), .A3(new_n18769_), .ZN(new_n18770_));
  AOI21_X1   g18706(.A1(new_n11788_), .A2(new_n11789_), .B(new_n8778_), .ZN(new_n18771_));
  NAND2_X1   g18707(.A1(new_n10865_), .A2(new_n8784_), .ZN(new_n18772_));
  NAND2_X1   g18708(.A1(new_n10875_), .A2(new_n8785_), .ZN(new_n18773_));
  AOI21_X1   g18709(.A1(new_n18773_), .A2(new_n18772_), .B(new_n8779_), .ZN(new_n18774_));
  OAI21_X1   g18710(.A1(new_n18771_), .A2(new_n18774_), .B(new_n18769_), .ZN(new_n18775_));
  NAND2_X1   g18711(.A1(new_n18775_), .A2(\a[2] ), .ZN(new_n18776_));
  NAND2_X1   g18712(.A1(new_n18770_), .A2(new_n18776_), .ZN(new_n18777_));
  OAI21_X1   g18713(.A1(new_n18766_), .A2(new_n18618_), .B(new_n18777_), .ZN(new_n18778_));
  NAND3_X1   g18714(.A1(new_n18709_), .A2(new_n18711_), .A3(new_n18708_), .ZN(new_n18779_));
  OAI21_X1   g18715(.A1(new_n18704_), .A2(new_n18690_), .B(new_n18624_), .ZN(new_n18780_));
  INV_X1     g18716(.I(new_n18719_), .ZN(new_n18781_));
  AOI21_X1   g18717(.A1(new_n18780_), .A2(new_n18779_), .B(new_n18781_), .ZN(new_n18782_));
  NAND2_X1   g18718(.A1(new_n18747_), .A2(new_n18740_), .ZN(new_n18783_));
  OAI21_X1   g18719(.A1(new_n18704_), .A2(new_n18690_), .B(new_n18624_), .ZN(new_n18784_));
  NAND2_X1   g18720(.A1(new_n18784_), .A2(new_n18783_), .ZN(new_n18785_));
  OAI21_X1   g18721(.A1(new_n18487_), .A2(new_n18494_), .B(new_n18761_), .ZN(new_n18786_));
  NAND3_X1   g18722(.A1(new_n18616_), .A2(new_n18750_), .A3(new_n18749_), .ZN(new_n18787_));
  AOI21_X1   g18723(.A1(new_n18786_), .A2(new_n18787_), .B(new_n18763_), .ZN(new_n18788_));
  OAI21_X1   g18724(.A1(new_n18782_), .A2(new_n18785_), .B(new_n18788_), .ZN(new_n18789_));
  AOI21_X1   g18725(.A1(new_n18757_), .A2(new_n18758_), .B(new_n18614_), .ZN(new_n18790_));
  INV_X1     g18726(.I(new_n18790_), .ZN(new_n18791_));
  NAND3_X1   g18727(.A1(new_n18295_), .A2(new_n18287_), .A3(new_n18290_), .ZN(new_n18792_));
  OAI21_X1   g18728(.A1(new_n18296_), .A2(new_n18297_), .B(new_n18283_), .ZN(new_n18793_));
  AOI21_X1   g18729(.A1(new_n18793_), .A2(new_n18792_), .B(new_n18274_), .ZN(new_n18794_));
  INV_X1     g18730(.I(new_n18274_), .ZN(new_n18795_));
  AOI21_X1   g18731(.A1(new_n18298_), .A2(new_n18291_), .B(new_n18795_), .ZN(new_n18796_));
  NOR2_X1    g18732(.A1(new_n18796_), .A2(new_n18794_), .ZN(new_n18797_));
  OAI22_X1   g18733(.A1(new_n9478_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n10846_), .ZN(new_n18798_));
  NAND2_X1   g18734(.A1(new_n10854_), .A2(new_n6838_), .ZN(new_n18799_));
  AOI21_X1   g18735(.A1(new_n18798_), .A2(new_n18799_), .B(new_n6836_), .ZN(new_n18800_));
  OAI21_X1   g18736(.A1(new_n13015_), .A2(new_n13012_), .B(new_n18800_), .ZN(new_n18801_));
  XOR2_X1    g18737(.A1(new_n18801_), .A2(new_n65_), .Z(new_n18802_));
  NAND2_X1   g18738(.A1(new_n18802_), .A2(new_n18797_), .ZN(new_n18803_));
  OR2_X2     g18739(.A1(new_n18796_), .A2(new_n18794_), .Z(new_n18804_));
  XOR2_X1    g18740(.A1(new_n18801_), .A2(\a[5] ), .Z(new_n18805_));
  NAND2_X1   g18741(.A1(new_n18804_), .A2(new_n18805_), .ZN(new_n18806_));
  AOI21_X1   g18742(.A1(new_n18806_), .A2(new_n18803_), .B(new_n18791_), .ZN(new_n18807_));
  NOR2_X1    g18743(.A1(new_n18804_), .A2(new_n18805_), .ZN(new_n18808_));
  NOR2_X1    g18744(.A1(new_n18802_), .A2(new_n18797_), .ZN(new_n18809_));
  NOR3_X1    g18745(.A1(new_n18808_), .A2(new_n18809_), .A3(new_n18790_), .ZN(new_n18810_));
  NOR2_X1    g18746(.A1(new_n18810_), .A2(new_n18807_), .ZN(new_n18811_));
  NOR2_X1    g18747(.A1(new_n18777_), .A2(new_n18811_), .ZN(new_n18812_));
  NAND3_X1   g18748(.A1(new_n18789_), .A2(new_n18617_), .A3(new_n18812_), .ZN(new_n18813_));
  AOI21_X1   g18749(.A1(new_n18778_), .A2(new_n18813_), .B(new_n18481_), .ZN(new_n18814_));
  INV_X1     g18750(.I(new_n18814_), .ZN(new_n18815_));
  XOR2_X1    g18751(.A1(new_n18480_), .A2(\a[2] ), .Z(new_n18816_));
  AND2_X2    g18752(.A1(new_n18770_), .A2(new_n18776_), .Z(new_n18817_));
  AOI21_X1   g18753(.A1(new_n18789_), .A2(new_n18617_), .B(new_n18817_), .ZN(new_n18818_));
  OAI21_X1   g18754(.A1(new_n18808_), .A2(new_n18809_), .B(new_n18790_), .ZN(new_n18819_));
  NAND3_X1   g18755(.A1(new_n18806_), .A2(new_n18803_), .A3(new_n18791_), .ZN(new_n18820_));
  NAND2_X1   g18756(.A1(new_n18819_), .A2(new_n18820_), .ZN(new_n18821_));
  NAND2_X1   g18757(.A1(new_n18817_), .A2(new_n18821_), .ZN(new_n18822_));
  NOR3_X1    g18758(.A1(new_n18766_), .A2(new_n18822_), .A3(new_n18618_), .ZN(new_n18823_));
  NOR3_X1    g18759(.A1(new_n18823_), .A2(new_n18818_), .A3(new_n18816_), .ZN(new_n18824_));
  AOI21_X1   g18760(.A1(new_n18778_), .A2(new_n18813_), .B(new_n18481_), .ZN(new_n18825_));
  XOR2_X1    g18761(.A1(new_n18302_), .A2(new_n18307_), .Z(new_n18826_));
  INV_X1     g18762(.I(new_n18308_), .ZN(new_n18827_));
  NOR2_X1    g18763(.A1(new_n18827_), .A2(new_n18309_), .ZN(new_n18828_));
  NOR2_X1    g18764(.A1(new_n18828_), .A2(new_n18299_), .ZN(new_n18829_));
  AOI21_X1   g18765(.A1(new_n18299_), .A2(new_n18826_), .B(new_n18829_), .ZN(new_n18830_));
  INV_X1     g18766(.I(new_n18830_), .ZN(new_n18831_));
  AOI21_X1   g18767(.A1(new_n18790_), .A2(new_n18803_), .B(new_n18809_), .ZN(new_n18832_));
  OAI22_X1   g18768(.A1(new_n9478_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n10853_), .ZN(new_n18833_));
  NAND2_X1   g18769(.A1(new_n10862_), .A2(new_n6838_), .ZN(new_n18834_));
  AOI21_X1   g18770(.A1(new_n18833_), .A2(new_n18834_), .B(new_n6836_), .ZN(new_n18835_));
  NAND2_X1   g18771(.A1(new_n13484_), .A2(new_n18835_), .ZN(new_n18836_));
  XOR2_X1    g18772(.A1(new_n18836_), .A2(\a[5] ), .Z(new_n18837_));
  INV_X1     g18773(.I(new_n18837_), .ZN(new_n18838_));
  NOR2_X1    g18774(.A1(new_n18832_), .A2(new_n18838_), .ZN(new_n18839_));
  INV_X1     g18775(.I(new_n18839_), .ZN(new_n18840_));
  NAND2_X1   g18776(.A1(new_n18832_), .A2(new_n18838_), .ZN(new_n18841_));
  AOI21_X1   g18777(.A1(new_n18840_), .A2(new_n18841_), .B(new_n18831_), .ZN(new_n18842_));
  INV_X1     g18778(.I(new_n18841_), .ZN(new_n18843_));
  NOR3_X1    g18779(.A1(new_n18843_), .A2(new_n18839_), .A3(new_n18830_), .ZN(new_n18844_));
  NOR2_X1    g18780(.A1(new_n18842_), .A2(new_n18844_), .ZN(new_n18845_));
  OAI21_X1   g18781(.A1(new_n18824_), .A2(new_n18825_), .B(new_n18845_), .ZN(new_n18846_));
  NAND3_X1   g18782(.A1(new_n18846_), .A2(new_n18476_), .A3(new_n18815_), .ZN(new_n18847_));
  NAND3_X1   g18783(.A1(new_n18778_), .A2(new_n18813_), .A3(new_n18481_), .ZN(new_n18848_));
  OAI21_X1   g18784(.A1(new_n18823_), .A2(new_n18818_), .B(new_n18816_), .ZN(new_n18849_));
  INV_X1     g18785(.I(new_n18845_), .ZN(new_n18850_));
  AOI22_X1   g18786(.A1(new_n18849_), .A2(new_n18848_), .B1(new_n18850_), .B2(new_n18481_), .ZN(new_n18851_));
  NAND2_X1   g18787(.A1(new_n18851_), .A2(new_n18475_), .ZN(new_n18852_));
  XOR2_X1    g18788(.A1(new_n18326_), .A2(new_n18332_), .Z(new_n18853_));
  AOI22_X1   g18789(.A1(new_n18847_), .A2(new_n18852_), .B1(new_n18476_), .B2(new_n18853_), .ZN(new_n18854_));
  NAND2_X1   g18790(.A1(new_n18854_), .A2(new_n18470_), .ZN(new_n18855_));
  NOR2_X1    g18791(.A1(new_n18854_), .A2(new_n18470_), .ZN(new_n18856_));
  INV_X1     g18792(.I(new_n18470_), .ZN(new_n18857_));
  NAND2_X1   g18793(.A1(new_n18851_), .A2(new_n18475_), .ZN(new_n18858_));
  AOI21_X1   g18794(.A1(new_n18849_), .A2(new_n18848_), .B(new_n18850_), .ZN(new_n18859_));
  NOR3_X1    g18795(.A1(new_n18859_), .A2(new_n18475_), .A3(new_n18814_), .ZN(new_n18860_));
  AOI21_X1   g18796(.A1(new_n18846_), .A2(new_n18815_), .B(new_n18476_), .ZN(new_n18861_));
  INV_X1     g18797(.I(new_n18853_), .ZN(new_n18862_));
  OAI21_X1   g18798(.A1(new_n18861_), .A2(new_n18860_), .B(new_n18862_), .ZN(new_n18863_));
  AOI21_X1   g18799(.A1(new_n18863_), .A2(new_n18858_), .B(new_n18857_), .ZN(new_n18864_));
  NAND3_X1   g18800(.A1(new_n18441_), .A2(new_n18440_), .A3(new_n18360_), .ZN(new_n18865_));
  OAI21_X1   g18801(.A1(new_n18352_), .A2(new_n18355_), .B(new_n18442_), .ZN(new_n18866_));
  AOI21_X1   g18802(.A1(new_n18866_), .A2(new_n18865_), .B(new_n18333_), .ZN(new_n18867_));
  AOI21_X1   g18803(.A1(new_n18361_), .A2(new_n18444_), .B(new_n18334_), .ZN(new_n18868_));
  NOR2_X1    g18804(.A1(new_n18868_), .A2(new_n18867_), .ZN(new_n18869_));
  OAI21_X1   g18805(.A1(new_n18856_), .A2(new_n18864_), .B(new_n18869_), .ZN(new_n18870_));
  AOI22_X1   g18806(.A1(new_n10886_), .A2(new_n6925_), .B1(new_n10889_), .B2(new_n9503_), .ZN(new_n18871_));
  NOR2_X1    g18807(.A1(new_n10899_), .A2(new_n9489_), .ZN(new_n18872_));
  OAI21_X1   g18808(.A1(new_n18872_), .A2(new_n18871_), .B(new_n6922_), .ZN(new_n18873_));
  NOR2_X1    g18809(.A1(new_n11908_), .A2(new_n18873_), .ZN(new_n18874_));
  XOR2_X1    g18810(.A1(new_n18874_), .A2(new_n4387_), .Z(new_n18875_));
  AOI21_X1   g18811(.A1(new_n18870_), .A2(new_n18855_), .B(new_n18875_), .ZN(new_n18876_));
  INV_X1     g18812(.I(new_n18855_), .ZN(new_n18877_));
  NAND3_X1   g18813(.A1(new_n18863_), .A2(new_n18857_), .A3(new_n18858_), .ZN(new_n18878_));
  NAND2_X1   g18814(.A1(new_n18854_), .A2(new_n18470_), .ZN(new_n18879_));
  INV_X1     g18815(.I(new_n18869_), .ZN(new_n18880_));
  AOI21_X1   g18816(.A1(new_n18879_), .A2(new_n18878_), .B(new_n18880_), .ZN(new_n18881_));
  INV_X1     g18817(.I(new_n18875_), .ZN(new_n18882_));
  OAI21_X1   g18818(.A1(new_n18413_), .A2(new_n18446_), .B(new_n18363_), .ZN(new_n18883_));
  NAND3_X1   g18819(.A1(new_n18445_), .A2(new_n18406_), .A3(new_n18402_), .ZN(new_n18884_));
  AOI21_X1   g18820(.A1(new_n18883_), .A2(new_n18884_), .B(new_n18882_), .ZN(new_n18885_));
  INV_X1     g18821(.I(new_n18885_), .ZN(new_n18886_));
  NOR3_X1    g18822(.A1(new_n18881_), .A2(new_n18877_), .A3(new_n18886_), .ZN(new_n18887_));
  AOI22_X1   g18823(.A1(new_n11899_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n10889_), .ZN(new_n18888_));
  NOR2_X1    g18824(.A1(new_n8774_), .A2(new_n9489_), .ZN(new_n18889_));
  OAI21_X1   g18825(.A1(new_n18889_), .A2(new_n18888_), .B(new_n6922_), .ZN(new_n18890_));
  NOR2_X1    g18826(.A1(new_n11945_), .A2(new_n18890_), .ZN(new_n18891_));
  XOR2_X1    g18827(.A1(new_n18891_), .A2(new_n4387_), .Z(new_n18892_));
  NOR2_X1    g18828(.A1(new_n18447_), .A2(new_n18413_), .ZN(new_n18893_));
  XOR2_X1    g18829(.A1(new_n18248_), .A2(new_n18411_), .Z(new_n18894_));
  NOR2_X1    g18830(.A1(new_n18893_), .A2(new_n18894_), .ZN(new_n18895_));
  NAND2_X1   g18831(.A1(new_n18407_), .A2(new_n18402_), .ZN(new_n18896_));
  INV_X1     g18832(.I(new_n18894_), .ZN(new_n18897_));
  NOR2_X1    g18833(.A1(new_n18897_), .A2(new_n18896_), .ZN(new_n18898_));
  OAI21_X1   g18834(.A1(new_n18898_), .A2(new_n18895_), .B(new_n18892_), .ZN(new_n18899_));
  NOR3_X1    g18835(.A1(new_n18876_), .A2(new_n18887_), .A3(new_n18899_), .ZN(new_n18900_));
  OAI21_X1   g18836(.A1(new_n18881_), .A2(new_n18877_), .B(new_n18882_), .ZN(new_n18901_));
  NAND3_X1   g18837(.A1(new_n18870_), .A2(new_n18855_), .A3(new_n18885_), .ZN(new_n18902_));
  AOI21_X1   g18838(.A1(new_n18901_), .A2(new_n18902_), .B(new_n18892_), .ZN(new_n18903_));
  NOR3_X1    g18839(.A1(new_n18903_), .A2(new_n18900_), .A3(new_n18464_), .ZN(new_n18904_));
  NAND2_X1   g18840(.A1(new_n8761_), .A2(new_n9488_), .ZN(new_n18905_));
  NAND2_X1   g18841(.A1(new_n11996_), .A2(new_n9503_), .ZN(new_n18906_));
  AOI21_X1   g18842(.A1(new_n10906_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n18907_));
  NAND4_X1   g18843(.A1(new_n12053_), .A2(new_n18905_), .A3(new_n18906_), .A4(new_n18907_), .ZN(new_n18908_));
  XOR2_X1    g18844(.A1(new_n18908_), .A2(\a[2] ), .Z(new_n18909_));
  INV_X1     g18845(.I(new_n18909_), .ZN(new_n18910_));
  OAI21_X1   g18846(.A1(new_n18904_), .A2(new_n18465_), .B(new_n18910_), .ZN(new_n18911_));
  NAND3_X1   g18847(.A1(new_n18458_), .A2(new_n18462_), .A3(new_n18247_), .ZN(new_n18912_));
  OAI21_X1   g18848(.A1(new_n18455_), .A2(new_n18439_), .B(new_n18246_), .ZN(new_n18913_));
  NAND2_X1   g18849(.A1(new_n18913_), .A2(new_n18912_), .ZN(new_n18914_));
  NAND2_X1   g18850(.A1(new_n18914_), .A2(new_n18246_), .ZN(new_n18915_));
  INV_X1     g18851(.I(new_n18892_), .ZN(new_n18916_));
  NAND2_X1   g18852(.A1(new_n18897_), .A2(new_n18896_), .ZN(new_n18917_));
  NAND2_X1   g18853(.A1(new_n18893_), .A2(new_n18894_), .ZN(new_n18918_));
  AOI21_X1   g18854(.A1(new_n18917_), .A2(new_n18918_), .B(new_n18916_), .ZN(new_n18919_));
  NAND3_X1   g18855(.A1(new_n18901_), .A2(new_n18902_), .A3(new_n18919_), .ZN(new_n18920_));
  OAI21_X1   g18856(.A1(new_n18876_), .A2(new_n18887_), .B(new_n18916_), .ZN(new_n18921_));
  NAND3_X1   g18857(.A1(new_n18921_), .A2(new_n18920_), .A3(new_n18914_), .ZN(new_n18922_));
  AOI21_X1   g18858(.A1(new_n18451_), .A2(new_n18459_), .B(new_n18453_), .ZN(new_n18923_));
  AOI22_X1   g18859(.A1(new_n10886_), .A2(new_n6846_), .B1(new_n10889_), .B2(new_n8799_), .ZN(new_n18924_));
  NOR2_X1    g18860(.A1(new_n10899_), .A2(new_n6839_), .ZN(new_n18925_));
  OAI21_X1   g18861(.A1(new_n18925_), .A2(new_n18924_), .B(new_n6835_), .ZN(new_n18926_));
  NOR2_X1    g18862(.A1(new_n11908_), .A2(new_n18926_), .ZN(new_n18927_));
  XOR2_X1    g18863(.A1(new_n18927_), .A2(new_n65_), .Z(new_n18928_));
  INV_X1     g18864(.I(new_n18928_), .ZN(new_n18929_));
  NAND3_X1   g18865(.A1(new_n18074_), .A2(new_n18069_), .A3(new_n18094_), .ZN(new_n18930_));
  OAI21_X1   g18866(.A1(new_n18043_), .A2(new_n18038_), .B(new_n18068_), .ZN(new_n18931_));
  AOI21_X1   g18867(.A1(new_n18931_), .A2(new_n18930_), .B(new_n18929_), .ZN(new_n18932_));
  NOR3_X1    g18868(.A1(new_n18043_), .A2(new_n18038_), .A3(new_n18068_), .ZN(new_n18933_));
  AOI21_X1   g18869(.A1(new_n18074_), .A2(new_n18094_), .B(new_n18069_), .ZN(new_n18934_));
  NOR3_X1    g18870(.A1(new_n18933_), .A2(new_n18934_), .A3(new_n18928_), .ZN(new_n18935_));
  OAI21_X1   g18871(.A1(new_n18932_), .A2(new_n18935_), .B(new_n18923_), .ZN(new_n18936_));
  OAI21_X1   g18872(.A1(new_n18415_), .A2(new_n18452_), .B(new_n18460_), .ZN(new_n18937_));
  OAI21_X1   g18873(.A1(new_n18933_), .A2(new_n18934_), .B(new_n18928_), .ZN(new_n18938_));
  NAND3_X1   g18874(.A1(new_n18931_), .A2(new_n18930_), .A3(new_n18929_), .ZN(new_n18939_));
  NAND3_X1   g18875(.A1(new_n18937_), .A2(new_n18938_), .A3(new_n18939_), .ZN(new_n18940_));
  AOI21_X1   g18876(.A1(new_n18936_), .A2(new_n18940_), .B(new_n18910_), .ZN(new_n18941_));
  NAND3_X1   g18877(.A1(new_n18922_), .A2(new_n18915_), .A3(new_n18941_), .ZN(new_n18942_));
  NAND3_X1   g18878(.A1(new_n18911_), .A2(new_n18942_), .A3(new_n18242_), .ZN(new_n18943_));
  AOI21_X1   g18879(.A1(new_n18922_), .A2(new_n18915_), .B(new_n18909_), .ZN(new_n18944_));
  INV_X1     g18880(.I(new_n18941_), .ZN(new_n18945_));
  NOR3_X1    g18881(.A1(new_n18904_), .A2(new_n18945_), .A3(new_n18465_), .ZN(new_n18946_));
  OAI21_X1   g18882(.A1(new_n18946_), .A2(new_n18944_), .B(new_n18241_), .ZN(new_n18947_));
  NAND2_X1   g18883(.A1(new_n18095_), .A2(new_n18074_), .ZN(new_n18948_));
  NAND2_X1   g18884(.A1(new_n18948_), .A2(new_n18018_), .ZN(new_n18949_));
  INV_X1     g18885(.I(new_n18018_), .ZN(new_n18950_));
  NOR2_X1    g18886(.A1(new_n18070_), .A2(new_n18038_), .ZN(new_n18951_));
  NAND2_X1   g18887(.A1(new_n18951_), .A2(new_n18950_), .ZN(new_n18952_));
  AOI21_X1   g18888(.A1(new_n18952_), .A2(new_n18949_), .B(new_n18025_), .ZN(new_n18953_));
  NOR2_X1    g18889(.A1(new_n18951_), .A2(new_n18950_), .ZN(new_n18954_));
  NOR2_X1    g18890(.A1(new_n18948_), .A2(new_n18018_), .ZN(new_n18955_));
  NOR3_X1    g18891(.A1(new_n18954_), .A2(new_n18955_), .A3(new_n18024_), .ZN(new_n18956_));
  AOI22_X1   g18892(.A1(new_n11899_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n10889_), .ZN(new_n18957_));
  NOR2_X1    g18893(.A1(new_n8774_), .A2(new_n6839_), .ZN(new_n18958_));
  OAI21_X1   g18894(.A1(new_n18958_), .A2(new_n18957_), .B(new_n6835_), .ZN(new_n18959_));
  NOR2_X1    g18895(.A1(new_n11945_), .A2(new_n18959_), .ZN(new_n18960_));
  XOR2_X1    g18896(.A1(new_n18960_), .A2(new_n65_), .Z(new_n18961_));
  NOR3_X1    g18897(.A1(new_n18953_), .A2(new_n18956_), .A3(new_n18961_), .ZN(new_n18962_));
  OAI21_X1   g18898(.A1(new_n18954_), .A2(new_n18955_), .B(new_n18024_), .ZN(new_n18963_));
  NAND3_X1   g18899(.A1(new_n18952_), .A2(new_n18949_), .A3(new_n18025_), .ZN(new_n18964_));
  INV_X1     g18900(.I(new_n18961_), .ZN(new_n18965_));
  AOI21_X1   g18901(.A1(new_n18963_), .A2(new_n18964_), .B(new_n18965_), .ZN(new_n18966_));
  AOI21_X1   g18902(.A1(new_n18923_), .A2(new_n18939_), .B(new_n18932_), .ZN(new_n18967_));
  INV_X1     g18903(.I(new_n18967_), .ZN(new_n18968_));
  NOR3_X1    g18904(.A1(new_n18962_), .A2(new_n18966_), .A3(new_n18968_), .ZN(new_n18969_));
  NAND3_X1   g18905(.A1(new_n18963_), .A2(new_n18964_), .A3(new_n18965_), .ZN(new_n18970_));
  OAI21_X1   g18906(.A1(new_n18953_), .A2(new_n18956_), .B(new_n18961_), .ZN(new_n18971_));
  AOI21_X1   g18907(.A1(new_n18971_), .A2(new_n18970_), .B(new_n18967_), .ZN(new_n18972_));
  NOR2_X1    g18908(.A1(new_n18969_), .A2(new_n18972_), .ZN(new_n18973_));
  INV_X1     g18909(.I(new_n18973_), .ZN(new_n18974_));
  AOI22_X1   g18910(.A1(new_n18947_), .A2(new_n18943_), .B1(new_n18242_), .B2(new_n18974_), .ZN(new_n18975_));
  NAND2_X1   g18911(.A1(new_n18975_), .A2(new_n18236_), .ZN(new_n18976_));
  AOI21_X1   g18912(.A1(new_n18911_), .A2(new_n18942_), .B(new_n18242_), .ZN(new_n18977_));
  AOI21_X1   g18913(.A1(new_n18947_), .A2(new_n18943_), .B(new_n18974_), .ZN(new_n18978_));
  NOR3_X1    g18914(.A1(new_n18978_), .A2(new_n18236_), .A3(new_n18977_), .ZN(new_n18979_));
  INV_X1     g18915(.I(new_n18236_), .ZN(new_n18980_));
  INV_X1     g18916(.I(new_n18977_), .ZN(new_n18981_));
  NOR3_X1    g18917(.A1(new_n18946_), .A2(new_n18944_), .A3(new_n18241_), .ZN(new_n18982_));
  AOI21_X1   g18918(.A1(new_n18911_), .A2(new_n18942_), .B(new_n18242_), .ZN(new_n18983_));
  OAI21_X1   g18919(.A1(new_n18982_), .A2(new_n18983_), .B(new_n18973_), .ZN(new_n18984_));
  AOI21_X1   g18920(.A1(new_n18984_), .A2(new_n18981_), .B(new_n18980_), .ZN(new_n18985_));
  INV_X1     g18921(.I(new_n18076_), .ZN(new_n18986_));
  XNOR2_X1   g18922(.A1(new_n18082_), .A2(new_n18087_), .ZN(new_n18987_));
  NOR2_X1    g18923(.A1(new_n18986_), .A2(new_n18987_), .ZN(new_n18988_));
  NAND2_X1   g18924(.A1(new_n18091_), .A2(new_n18088_), .ZN(new_n18989_));
  AOI21_X1   g18925(.A1(new_n18986_), .A2(new_n18989_), .B(new_n18988_), .ZN(new_n18990_));
  INV_X1     g18926(.I(new_n18990_), .ZN(new_n18991_));
  NOR3_X1    g18927(.A1(new_n18962_), .A2(new_n18966_), .A3(new_n18967_), .ZN(new_n18992_));
  OAI22_X1   g18928(.A1(new_n8774_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n10899_), .ZN(new_n18993_));
  NAND2_X1   g18929(.A1(new_n11996_), .A2(new_n6838_), .ZN(new_n18994_));
  AOI21_X1   g18930(.A1(new_n18994_), .A2(new_n18993_), .B(new_n6836_), .ZN(new_n18995_));
  NAND2_X1   g18931(.A1(new_n12001_), .A2(new_n18995_), .ZN(new_n18996_));
  XOR2_X1    g18932(.A1(new_n18996_), .A2(\a[5] ), .Z(new_n18997_));
  INV_X1     g18933(.I(new_n18997_), .ZN(new_n18998_));
  NOR2_X1    g18934(.A1(new_n18992_), .A2(new_n18998_), .ZN(new_n18999_));
  NOR4_X1    g18935(.A1(new_n18962_), .A2(new_n18966_), .A3(new_n18967_), .A4(new_n18997_), .ZN(new_n19000_));
  NOR2_X1    g18936(.A1(new_n18999_), .A2(new_n19000_), .ZN(new_n19001_));
  XOR2_X1    g18937(.A1(new_n19001_), .A2(new_n18991_), .Z(new_n19002_));
  OAI21_X1   g18938(.A1(new_n18985_), .A2(new_n18979_), .B(new_n19002_), .ZN(new_n19003_));
  OAI22_X1   g18939(.A1(new_n8751_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n8745_), .ZN(new_n19004_));
  NAND2_X1   g18940(.A1(new_n10927_), .A2(new_n9488_), .ZN(new_n19005_));
  AOI21_X1   g18941(.A1(new_n19004_), .A2(new_n19005_), .B(new_n9482_), .ZN(new_n19006_));
  NAND2_X1   g18942(.A1(new_n12072_), .A2(new_n19006_), .ZN(new_n19007_));
  XOR2_X1    g18943(.A1(new_n19007_), .A2(\a[2] ), .Z(new_n19008_));
  AOI21_X1   g18944(.A1(new_n19003_), .A2(new_n18976_), .B(new_n19008_), .ZN(new_n19009_));
  NAND3_X1   g18945(.A1(new_n18984_), .A2(new_n18980_), .A3(new_n18981_), .ZN(new_n19010_));
  NAND2_X1   g18946(.A1(new_n18975_), .A2(new_n18236_), .ZN(new_n19011_));
  XOR2_X1    g18947(.A1(new_n19001_), .A2(new_n18990_), .Z(new_n19012_));
  AOI22_X1   g18948(.A1(new_n19010_), .A2(new_n19011_), .B1(new_n18980_), .B2(new_n19012_), .ZN(new_n19013_));
  INV_X1     g18949(.I(new_n19008_), .ZN(new_n19014_));
  NAND3_X1   g18950(.A1(new_n18106_), .A2(new_n18110_), .A3(new_n18115_), .ZN(new_n19015_));
  AOI21_X1   g18951(.A1(new_n18217_), .A2(new_n19015_), .B(new_n19014_), .ZN(new_n19016_));
  INV_X1     g18952(.I(new_n19016_), .ZN(new_n19017_));
  NOR2_X1    g18953(.A1(new_n19013_), .A2(new_n19017_), .ZN(new_n19018_));
  OAI22_X1   g18954(.A1(new_n8751_), .A2(new_n9485_), .B1(new_n9483_), .B2(new_n10924_), .ZN(new_n19019_));
  NAND2_X1   g18955(.A1(new_n8736_), .A2(new_n9488_), .ZN(new_n19020_));
  AOI21_X1   g18956(.A1(new_n19020_), .A2(new_n19019_), .B(new_n9482_), .ZN(new_n19021_));
  NAND2_X1   g18957(.A1(new_n12118_), .A2(new_n19021_), .ZN(new_n19022_));
  XOR2_X1    g18958(.A1(new_n19022_), .A2(\a[2] ), .Z(new_n19023_));
  INV_X1     g18959(.I(new_n19023_), .ZN(new_n19024_));
  NAND3_X1   g18960(.A1(new_n18116_), .A2(new_n18164_), .A3(new_n18165_), .ZN(new_n19025_));
  OAI21_X1   g18961(.A1(new_n18163_), .A2(new_n18166_), .B(new_n18217_), .ZN(new_n19026_));
  AOI21_X1   g18962(.A1(new_n19026_), .A2(new_n19025_), .B(new_n19024_), .ZN(new_n19027_));
  INV_X1     g18963(.I(new_n19027_), .ZN(new_n19028_));
  NOR3_X1    g18964(.A1(new_n19018_), .A2(new_n19009_), .A3(new_n19028_), .ZN(new_n19029_));
  NAND2_X1   g18965(.A1(new_n19013_), .A2(new_n19014_), .ZN(new_n19030_));
  NAND3_X1   g18966(.A1(new_n19003_), .A2(new_n18976_), .A3(new_n19016_), .ZN(new_n19031_));
  AOI21_X1   g18967(.A1(new_n19030_), .A2(new_n19031_), .B(new_n19023_), .ZN(new_n19032_));
  NOR3_X1    g18968(.A1(new_n19029_), .A2(new_n19032_), .A3(new_n18230_), .ZN(new_n19033_));
  NOR2_X1    g18969(.A1(new_n8725_), .A2(new_n9483_), .ZN(new_n19034_));
  NOR2_X1    g18970(.A1(new_n8718_), .A2(new_n9489_), .ZN(new_n19035_));
  NOR2_X1    g18971(.A1(new_n8735_), .A2(new_n9485_), .ZN(new_n19036_));
  NOR4_X1    g18972(.A1(new_n19034_), .A2(new_n9482_), .A3(new_n19035_), .A4(new_n19036_), .ZN(new_n19037_));
  NAND2_X1   g18973(.A1(new_n12242_), .A2(new_n19037_), .ZN(new_n19038_));
  XOR2_X1    g18974(.A1(new_n19038_), .A2(\a[2] ), .Z(new_n19039_));
  INV_X1     g18975(.I(new_n19039_), .ZN(new_n19040_));
  OAI21_X1   g18976(.A1(new_n19033_), .A2(new_n18231_), .B(new_n19040_), .ZN(new_n19041_));
  NAND3_X1   g18977(.A1(new_n18225_), .A2(new_n18228_), .A3(new_n17881_), .ZN(new_n19042_));
  OAI21_X1   g18978(.A1(new_n18221_), .A2(new_n18213_), .B(new_n17880_), .ZN(new_n19043_));
  NAND2_X1   g18979(.A1(new_n19043_), .A2(new_n19042_), .ZN(new_n19044_));
  NAND2_X1   g18980(.A1(new_n19044_), .A2(new_n17880_), .ZN(new_n19045_));
  NAND3_X1   g18981(.A1(new_n19030_), .A2(new_n19031_), .A3(new_n19027_), .ZN(new_n19046_));
  OAI21_X1   g18982(.A1(new_n19018_), .A2(new_n19009_), .B(new_n19024_), .ZN(new_n19047_));
  NAND3_X1   g18983(.A1(new_n19047_), .A2(new_n19046_), .A3(new_n19044_), .ZN(new_n19048_));
  AOI21_X1   g18984(.A1(new_n18218_), .A2(new_n18219_), .B(new_n18227_), .ZN(new_n19049_));
  INV_X1     g18985(.I(new_n19049_), .ZN(new_n19050_));
  OAI22_X1   g18986(.A1(new_n8751_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n8745_), .ZN(new_n19051_));
  NAND2_X1   g18987(.A1(new_n10927_), .A2(new_n6838_), .ZN(new_n19052_));
  AOI21_X1   g18988(.A1(new_n19051_), .A2(new_n19052_), .B(new_n6836_), .ZN(new_n19053_));
  NAND2_X1   g18989(.A1(new_n12072_), .A2(new_n19053_), .ZN(new_n19054_));
  XOR2_X1    g18990(.A1(new_n19054_), .A2(\a[5] ), .Z(new_n19055_));
  NAND2_X1   g18991(.A1(new_n18170_), .A2(new_n18183_), .ZN(new_n19056_));
  NOR2_X1    g18992(.A1(new_n16443_), .A2(new_n16444_), .ZN(new_n19057_));
  XOR2_X1    g18993(.A1(new_n19057_), .A2(new_n16447_), .Z(new_n19058_));
  AOI22_X1   g18994(.A1(new_n10886_), .A2(new_n6480_), .B1(new_n10889_), .B2(new_n4720_), .ZN(new_n19059_));
  NOR2_X1    g18995(.A1(new_n10899_), .A2(new_n4710_), .ZN(new_n19060_));
  OAI21_X1   g18996(.A1(new_n19060_), .A2(new_n19059_), .B(new_n4706_), .ZN(new_n19061_));
  NOR2_X1    g18997(.A1(new_n11908_), .A2(new_n19061_), .ZN(new_n19062_));
  XOR2_X1    g18998(.A1(new_n19062_), .A2(new_n4034_), .Z(new_n19063_));
  INV_X1     g18999(.I(new_n19063_), .ZN(new_n19064_));
  NOR2_X1    g19000(.A1(new_n19058_), .A2(new_n19064_), .ZN(new_n19065_));
  INV_X1     g19001(.I(new_n19065_), .ZN(new_n19066_));
  NAND2_X1   g19002(.A1(new_n19058_), .A2(new_n19064_), .ZN(new_n19067_));
  AOI22_X1   g19003(.A1(new_n19056_), .A2(new_n18184_), .B1(new_n19066_), .B2(new_n19067_), .ZN(new_n19068_));
  NAND2_X1   g19004(.A1(new_n19056_), .A2(new_n18184_), .ZN(new_n19069_));
  XOR2_X1    g19005(.A1(new_n19058_), .A2(new_n19063_), .Z(new_n19070_));
  NOR2_X1    g19006(.A1(new_n19069_), .A2(new_n19070_), .ZN(new_n19071_));
  NOR2_X1    g19007(.A1(new_n19071_), .A2(new_n19068_), .ZN(new_n19072_));
  AOI22_X1   g19008(.A1(new_n7530_), .A2(new_n10906_), .B1(new_n11996_), .B2(new_n6789_), .ZN(new_n19073_));
  NOR2_X1    g19009(.A1(new_n8758_), .A2(new_n6785_), .ZN(new_n19074_));
  OAI21_X1   g19010(.A1(new_n19073_), .A2(new_n19074_), .B(new_n6775_), .ZN(new_n19075_));
  NOR2_X1    g19011(.A1(new_n12053_), .A2(new_n19075_), .ZN(new_n19076_));
  XOR2_X1    g19012(.A1(new_n19076_), .A2(new_n4009_), .Z(new_n19077_));
  NAND2_X1   g19013(.A1(new_n19072_), .A2(new_n19077_), .ZN(new_n19078_));
  OR2_X2     g19014(.A1(new_n19072_), .A2(new_n19077_), .Z(new_n19079_));
  NAND2_X1   g19015(.A1(new_n19079_), .A2(new_n19078_), .ZN(new_n19080_));
  NAND2_X1   g19016(.A1(new_n19080_), .A2(new_n19055_), .ZN(new_n19081_));
  INV_X1     g19017(.I(new_n19081_), .ZN(new_n19082_));
  NOR2_X1    g19018(.A1(new_n19080_), .A2(new_n19055_), .ZN(new_n19083_));
  NOR2_X1    g19019(.A1(new_n19082_), .A2(new_n19083_), .ZN(new_n19084_));
  NAND2_X1   g19020(.A1(new_n19050_), .A2(new_n19084_), .ZN(new_n19085_));
  OAI21_X1   g19021(.A1(new_n19082_), .A2(new_n19083_), .B(new_n19049_), .ZN(new_n19086_));
  AOI21_X1   g19022(.A1(new_n19085_), .A2(new_n19086_), .B(new_n19040_), .ZN(new_n19087_));
  NAND3_X1   g19023(.A1(new_n19048_), .A2(new_n19045_), .A3(new_n19087_), .ZN(new_n19088_));
  AOI21_X1   g19024(.A1(new_n19041_), .A2(new_n19088_), .B(new_n17875_), .ZN(new_n19089_));
  INV_X1     g19025(.I(new_n19089_), .ZN(new_n19090_));
  AOI21_X1   g19026(.A1(new_n19048_), .A2(new_n19045_), .B(new_n19039_), .ZN(new_n19091_));
  INV_X1     g19027(.I(new_n19087_), .ZN(new_n19092_));
  NOR3_X1    g19028(.A1(new_n19033_), .A2(new_n18231_), .A3(new_n19092_), .ZN(new_n19093_));
  NOR3_X1    g19029(.A1(new_n19093_), .A2(new_n19091_), .A3(new_n17874_), .ZN(new_n19094_));
  AOI21_X1   g19030(.A1(new_n19041_), .A2(new_n19088_), .B(new_n17875_), .ZN(new_n19095_));
  INV_X1     g19031(.I(new_n19067_), .ZN(new_n19096_));
  AOI21_X1   g19032(.A1(new_n19069_), .A2(new_n19066_), .B(new_n19096_), .ZN(new_n19097_));
  NOR2_X1    g19033(.A1(new_n16448_), .A2(new_n16395_), .ZN(new_n19098_));
  XOR2_X1    g19034(.A1(new_n19098_), .A2(new_n16406_), .Z(new_n19099_));
  XOR2_X1    g19035(.A1(new_n19099_), .A2(new_n16282_), .Z(new_n19100_));
  AOI22_X1   g19036(.A1(new_n11899_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n10889_), .ZN(new_n19101_));
  NOR2_X1    g19037(.A1(new_n8774_), .A2(new_n4710_), .ZN(new_n19102_));
  OAI21_X1   g19038(.A1(new_n19102_), .A2(new_n19101_), .B(new_n4706_), .ZN(new_n19103_));
  NOR2_X1    g19039(.A1(new_n11945_), .A2(new_n19103_), .ZN(new_n19104_));
  XOR2_X1    g19040(.A1(new_n19104_), .A2(new_n4034_), .Z(new_n19105_));
  INV_X1     g19041(.I(new_n19105_), .ZN(new_n19106_));
  NAND2_X1   g19042(.A1(new_n19100_), .A2(new_n19106_), .ZN(new_n19107_));
  XNOR2_X1   g19043(.A1(new_n19099_), .A2(new_n16282_), .ZN(new_n19108_));
  NAND2_X1   g19044(.A1(new_n19108_), .A2(new_n19105_), .ZN(new_n19109_));
  NAND2_X1   g19045(.A1(new_n19109_), .A2(new_n19107_), .ZN(new_n19110_));
  OAI22_X1   g19046(.A1(new_n8758_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8766_), .ZN(new_n19111_));
  NAND2_X1   g19047(.A1(new_n8746_), .A2(new_n6784_), .ZN(new_n19112_));
  AOI21_X1   g19048(.A1(new_n19112_), .A2(new_n19111_), .B(new_n6776_), .ZN(new_n19113_));
  NAND2_X1   g19049(.A1(new_n11964_), .A2(new_n19113_), .ZN(new_n19114_));
  XOR2_X1    g19050(.A1(new_n19114_), .A2(\a[8] ), .Z(new_n19115_));
  INV_X1     g19051(.I(new_n19115_), .ZN(new_n19116_));
  XOR2_X1    g19052(.A1(new_n19110_), .A2(new_n19116_), .Z(new_n19117_));
  NOR2_X1    g19053(.A1(new_n19117_), .A2(new_n19097_), .ZN(new_n19118_));
  XOR2_X1    g19054(.A1(new_n19110_), .A2(new_n19116_), .Z(new_n19119_));
  AOI21_X1   g19055(.A1(new_n19097_), .A2(new_n19119_), .B(new_n19118_), .ZN(new_n19120_));
  OAI22_X1   g19056(.A1(new_n8751_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n10924_), .ZN(new_n19121_));
  NAND2_X1   g19057(.A1(new_n8736_), .A2(new_n6838_), .ZN(new_n19122_));
  AOI21_X1   g19058(.A1(new_n19122_), .A2(new_n19121_), .B(new_n6836_), .ZN(new_n19123_));
  NAND2_X1   g19059(.A1(new_n12118_), .A2(new_n19123_), .ZN(new_n19124_));
  XOR2_X1    g19060(.A1(new_n19124_), .A2(\a[5] ), .Z(new_n19125_));
  XOR2_X1    g19061(.A1(new_n19120_), .A2(new_n19125_), .Z(new_n19126_));
  INV_X1     g19062(.I(new_n19125_), .ZN(new_n19127_));
  XOR2_X1    g19063(.A1(new_n19120_), .A2(new_n19127_), .Z(new_n19128_));
  MUX2_X1    g19064(.I0(new_n19126_), .I1(new_n19128_), .S(new_n19079_), .Z(new_n19129_));
  AOI21_X1   g19065(.A1(new_n19084_), .A2(new_n19049_), .B(new_n19082_), .ZN(new_n19130_));
  XOR2_X1    g19066(.A1(new_n19129_), .A2(new_n19130_), .Z(new_n19131_));
  OAI21_X1   g19067(.A1(new_n19094_), .A2(new_n19095_), .B(new_n19131_), .ZN(new_n19132_));
  NAND3_X1   g19068(.A1(new_n19132_), .A2(new_n17869_), .A3(new_n19090_), .ZN(new_n19133_));
  NAND3_X1   g19069(.A1(new_n19041_), .A2(new_n19088_), .A3(new_n17875_), .ZN(new_n19134_));
  OAI21_X1   g19070(.A1(new_n19093_), .A2(new_n19091_), .B(new_n17874_), .ZN(new_n19135_));
  INV_X1     g19071(.I(new_n19130_), .ZN(new_n19136_));
  XOR2_X1    g19072(.A1(new_n19129_), .A2(new_n19136_), .Z(new_n19137_));
  AOI22_X1   g19073(.A1(new_n19135_), .A2(new_n19134_), .B1(new_n17875_), .B2(new_n19137_), .ZN(new_n19138_));
  NAND2_X1   g19074(.A1(new_n19138_), .A2(new_n17868_), .ZN(new_n19139_));
  NAND2_X1   g19075(.A1(new_n16411_), .A2(new_n16414_), .ZN(new_n19140_));
  XOR2_X1    g19076(.A1(new_n19140_), .A2(new_n16419_), .Z(new_n19141_));
  NOR2_X1    g19077(.A1(new_n19141_), .A2(new_n16409_), .ZN(new_n19142_));
  NOR2_X1    g19078(.A1(new_n16454_), .A2(new_n16420_), .ZN(new_n19143_));
  NOR2_X1    g19079(.A1(new_n19143_), .A2(new_n16452_), .ZN(new_n19144_));
  NOR2_X1    g19080(.A1(new_n19142_), .A2(new_n19144_), .ZN(new_n19145_));
  NAND3_X1   g19081(.A1(new_n19097_), .A2(new_n19107_), .A3(new_n19109_), .ZN(new_n19146_));
  NAND2_X1   g19082(.A1(new_n19146_), .A2(new_n19109_), .ZN(new_n19147_));
  OAI22_X1   g19083(.A1(new_n8774_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n10899_), .ZN(new_n19148_));
  NAND2_X1   g19084(.A1(new_n11996_), .A2(new_n4709_), .ZN(new_n19149_));
  AOI21_X1   g19085(.A1(new_n19149_), .A2(new_n19148_), .B(new_n4707_), .ZN(new_n19150_));
  NAND2_X1   g19086(.A1(new_n12001_), .A2(new_n19150_), .ZN(new_n19151_));
  XOR2_X1    g19087(.A1(new_n19151_), .A2(\a[11] ), .Z(new_n19152_));
  XOR2_X1    g19088(.A1(new_n19147_), .A2(new_n19152_), .Z(new_n19153_));
  XOR2_X1    g19089(.A1(new_n19153_), .A2(new_n19145_), .Z(new_n19154_));
  XNOR2_X1   g19090(.A1(new_n19097_), .A2(new_n19110_), .ZN(new_n19155_));
  AOI22_X1   g19091(.A1(new_n19120_), .A2(new_n19079_), .B1(new_n19115_), .B2(new_n19155_), .ZN(new_n19156_));
  OAI22_X1   g19092(.A1(new_n8745_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n8758_), .ZN(new_n19157_));
  NAND2_X1   g19093(.A1(new_n8752_), .A2(new_n6784_), .ZN(new_n19158_));
  AOI21_X1   g19094(.A1(new_n19158_), .A2(new_n19157_), .B(new_n6776_), .ZN(new_n19159_));
  NAND2_X1   g19095(.A1(new_n12189_), .A2(new_n19159_), .ZN(new_n19160_));
  XOR2_X1    g19096(.A1(new_n19160_), .A2(new_n4009_), .Z(new_n19161_));
  XOR2_X1    g19097(.A1(new_n19156_), .A2(new_n19161_), .Z(new_n19162_));
  XOR2_X1    g19098(.A1(new_n19162_), .A2(new_n19154_), .Z(new_n19163_));
  XOR2_X1    g19099(.A1(new_n19120_), .A2(new_n19079_), .Z(new_n19164_));
  NAND2_X1   g19100(.A1(new_n19164_), .A2(new_n19125_), .ZN(new_n19165_));
  NAND2_X1   g19101(.A1(new_n19129_), .A2(new_n19165_), .ZN(new_n19166_));
  OAI22_X1   g19102(.A1(new_n8735_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n10924_), .ZN(new_n19167_));
  NAND2_X1   g19103(.A1(new_n8726_), .A2(new_n6838_), .ZN(new_n19168_));
  AOI21_X1   g19104(.A1(new_n19168_), .A2(new_n19167_), .B(new_n6836_), .ZN(new_n19169_));
  NAND2_X1   g19105(.A1(new_n12181_), .A2(new_n19169_), .ZN(new_n19170_));
  XOR2_X1    g19106(.A1(new_n19170_), .A2(\a[5] ), .Z(new_n19171_));
  OAI21_X1   g19107(.A1(new_n19166_), .A2(new_n19130_), .B(new_n19171_), .ZN(new_n19172_));
  INV_X1     g19108(.I(new_n19172_), .ZN(new_n19173_));
  NOR3_X1    g19109(.A1(new_n19166_), .A2(new_n19130_), .A3(new_n19171_), .ZN(new_n19174_));
  OAI21_X1   g19110(.A1(new_n19173_), .A2(new_n19174_), .B(new_n19163_), .ZN(new_n19175_));
  INV_X1     g19111(.I(new_n19163_), .ZN(new_n19176_));
  INV_X1     g19112(.I(new_n19174_), .ZN(new_n19177_));
  NAND3_X1   g19113(.A1(new_n19177_), .A2(new_n19176_), .A3(new_n19172_), .ZN(new_n19178_));
  NAND2_X1   g19114(.A1(new_n19175_), .A2(new_n19178_), .ZN(new_n19179_));
  AOI22_X1   g19115(.A1(new_n19133_), .A2(new_n19139_), .B1(new_n17869_), .B2(new_n19179_), .ZN(new_n19180_));
  OAI22_X1   g19116(.A1(new_n8701_), .A2(new_n9483_), .B1(new_n8710_), .B2(new_n9485_), .ZN(new_n19181_));
  NAND2_X1   g19117(.A1(new_n8696_), .A2(new_n9488_), .ZN(new_n19182_));
  AOI21_X1   g19118(.A1(new_n19181_), .A2(new_n19182_), .B(new_n9482_), .ZN(new_n19183_));
  NAND2_X1   g19119(.A1(new_n11595_), .A2(new_n19183_), .ZN(new_n19184_));
  XOR2_X1    g19120(.A1(new_n19184_), .A2(\a[2] ), .Z(new_n19185_));
  INV_X1     g19121(.I(new_n19185_), .ZN(new_n19186_));
  NAND2_X1   g19122(.A1(new_n19180_), .A2(new_n19186_), .ZN(new_n19187_));
  NAND2_X1   g19123(.A1(new_n19138_), .A2(new_n17868_), .ZN(new_n19188_));
  AOI21_X1   g19124(.A1(new_n19135_), .A2(new_n19134_), .B(new_n19137_), .ZN(new_n19189_));
  NOR3_X1    g19125(.A1(new_n19189_), .A2(new_n17868_), .A3(new_n19089_), .ZN(new_n19190_));
  AOI21_X1   g19126(.A1(new_n19132_), .A2(new_n19090_), .B(new_n17869_), .ZN(new_n19191_));
  AOI21_X1   g19127(.A1(new_n19177_), .A2(new_n19172_), .B(new_n19176_), .ZN(new_n19192_));
  NOR3_X1    g19128(.A1(new_n19173_), .A2(new_n19174_), .A3(new_n19163_), .ZN(new_n19193_));
  NOR2_X1    g19129(.A1(new_n19192_), .A2(new_n19193_), .ZN(new_n19194_));
  OAI21_X1   g19130(.A1(new_n19191_), .A2(new_n19190_), .B(new_n19194_), .ZN(new_n19195_));
  XOR2_X1    g19131(.A1(new_n16473_), .A2(new_n16468_), .Z(new_n19196_));
  NOR2_X1    g19132(.A1(new_n19186_), .A2(new_n19196_), .ZN(new_n19197_));
  NAND3_X1   g19133(.A1(new_n19195_), .A2(new_n19188_), .A3(new_n19197_), .ZN(new_n19198_));
  OAI22_X1   g19134(.A1(new_n8701_), .A2(new_n9485_), .B1(new_n8694_), .B2(new_n9483_), .ZN(new_n19199_));
  NAND2_X1   g19135(.A1(new_n8682_), .A2(new_n9488_), .ZN(new_n19200_));
  AOI21_X1   g19136(.A1(new_n19200_), .A2(new_n19199_), .B(new_n9482_), .ZN(new_n19201_));
  NAND2_X1   g19137(.A1(new_n12347_), .A2(new_n19201_), .ZN(new_n19202_));
  XOR2_X1    g19138(.A1(new_n19202_), .A2(\a[2] ), .Z(new_n19203_));
  AOI21_X1   g19139(.A1(new_n19187_), .A2(new_n19198_), .B(new_n19203_), .ZN(new_n19204_));
  AOI21_X1   g19140(.A1(new_n19195_), .A2(new_n19188_), .B(new_n19185_), .ZN(new_n19205_));
  NOR3_X1    g19141(.A1(new_n19180_), .A2(new_n19186_), .A3(new_n19196_), .ZN(new_n19206_));
  INV_X1     g19142(.I(new_n19203_), .ZN(new_n19207_));
  NAND2_X1   g19143(.A1(new_n16539_), .A2(new_n16535_), .ZN(new_n19208_));
  XNOR2_X1   g19144(.A1(new_n19208_), .A2(new_n16474_), .ZN(new_n19209_));
  NOR2_X1    g19145(.A1(new_n19209_), .A2(new_n19207_), .ZN(new_n19210_));
  INV_X1     g19146(.I(new_n19210_), .ZN(new_n19211_));
  NOR3_X1    g19147(.A1(new_n19206_), .A2(new_n19205_), .A3(new_n19211_), .ZN(new_n19212_));
  OAI22_X1   g19148(.A1(new_n8681_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n8694_), .ZN(new_n19213_));
  NAND2_X1   g19149(.A1(new_n8688_), .A2(new_n9488_), .ZN(new_n19214_));
  AOI21_X1   g19150(.A1(new_n19214_), .A2(new_n19213_), .B(new_n9482_), .ZN(new_n19215_));
  NAND2_X1   g19151(.A1(new_n11420_), .A2(new_n19215_), .ZN(new_n19216_));
  XOR2_X1    g19152(.A1(new_n19216_), .A2(\a[2] ), .Z(new_n19217_));
  INV_X1     g19153(.I(new_n19217_), .ZN(new_n19218_));
  OAI21_X1   g19154(.A1(new_n19212_), .A2(new_n19204_), .B(new_n19218_), .ZN(new_n19219_));
  OAI21_X1   g19155(.A1(new_n19206_), .A2(new_n19205_), .B(new_n19207_), .ZN(new_n19220_));
  NAND3_X1   g19156(.A1(new_n19187_), .A2(new_n19198_), .A3(new_n19210_), .ZN(new_n19221_));
  NAND2_X1   g19157(.A1(new_n16691_), .A2(new_n16689_), .ZN(new_n19222_));
  XNOR2_X1   g19158(.A1(new_n19222_), .A2(new_n16686_), .ZN(new_n19223_));
  NOR2_X1    g19159(.A1(new_n19223_), .A2(new_n19218_), .ZN(new_n19224_));
  NAND3_X1   g19160(.A1(new_n19220_), .A2(new_n19221_), .A3(new_n19224_), .ZN(new_n19225_));
  NAND2_X1   g19161(.A1(new_n8674_), .A2(new_n9488_), .ZN(new_n19226_));
  NAND2_X1   g19162(.A1(new_n8688_), .A2(new_n9503_), .ZN(new_n19227_));
  AOI21_X1   g19163(.A1(new_n8682_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n19228_));
  NAND4_X1   g19164(.A1(new_n11431_), .A2(new_n19226_), .A3(new_n19227_), .A4(new_n19228_), .ZN(new_n19229_));
  XOR2_X1    g19165(.A1(new_n19229_), .A2(\a[2] ), .Z(new_n19230_));
  AOI21_X1   g19166(.A1(new_n19219_), .A2(new_n19225_), .B(new_n19230_), .ZN(new_n19231_));
  AOI21_X1   g19167(.A1(new_n19220_), .A2(new_n19221_), .B(new_n19217_), .ZN(new_n19232_));
  INV_X1     g19168(.I(new_n19224_), .ZN(new_n19233_));
  NOR3_X1    g19169(.A1(new_n19212_), .A2(new_n19204_), .A3(new_n19233_), .ZN(new_n19234_));
  INV_X1     g19170(.I(new_n19230_), .ZN(new_n19235_));
  NAND2_X1   g19171(.A1(new_n16690_), .A2(new_n16691_), .ZN(new_n19236_));
  XOR2_X1    g19172(.A1(new_n19236_), .A2(new_n16693_), .Z(new_n19237_));
  NOR2_X1    g19173(.A1(new_n19237_), .A2(new_n19235_), .ZN(new_n19238_));
  INV_X1     g19174(.I(new_n19238_), .ZN(new_n19239_));
  NOR3_X1    g19175(.A1(new_n19234_), .A2(new_n19232_), .A3(new_n19239_), .ZN(new_n19240_));
  NOR3_X1    g19176(.A1(new_n19240_), .A2(new_n19231_), .A3(new_n17862_), .ZN(new_n19241_));
  NOR2_X1    g19177(.A1(new_n16240_), .A2(new_n16234_), .ZN(new_n19242_));
  NAND2_X1   g19178(.A1(new_n16695_), .A2(new_n16622_), .ZN(new_n19243_));
  XOR2_X1    g19179(.A1(new_n19243_), .A2(new_n16190_), .Z(new_n19244_));
  XNOR2_X1   g19180(.A1(new_n19244_), .A2(new_n19242_), .ZN(new_n19245_));
  INV_X1     g19181(.I(new_n19245_), .ZN(new_n19246_));
  OAI22_X1   g19182(.A1(new_n8661_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n8673_), .ZN(new_n19247_));
  NAND2_X1   g19183(.A1(new_n11285_), .A2(new_n9488_), .ZN(new_n19248_));
  AOI21_X1   g19184(.A1(new_n19248_), .A2(new_n19247_), .B(new_n9482_), .ZN(new_n19249_));
  NAND2_X1   g19185(.A1(new_n11323_), .A2(new_n19249_), .ZN(new_n19250_));
  XOR2_X1    g19186(.A1(new_n19250_), .A2(\a[2] ), .Z(new_n19251_));
  NAND2_X1   g19187(.A1(new_n19246_), .A2(new_n19251_), .ZN(new_n19252_));
  XOR2_X1    g19188(.A1(new_n19245_), .A2(new_n19251_), .Z(new_n19253_));
  INV_X1     g19189(.I(new_n19253_), .ZN(new_n19254_));
  NAND3_X1   g19190(.A1(new_n19254_), .A2(new_n17862_), .A3(new_n19252_), .ZN(new_n19255_));
  OAI22_X1   g19191(.A1(new_n11284_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n8661_), .ZN(new_n19256_));
  NAND2_X1   g19192(.A1(new_n11272_), .A2(new_n9488_), .ZN(new_n19257_));
  AOI21_X1   g19193(.A1(new_n19256_), .A2(new_n19257_), .B(new_n9482_), .ZN(new_n19258_));
  NAND2_X1   g19194(.A1(new_n11655_), .A2(new_n19258_), .ZN(new_n19259_));
  XOR2_X1    g19195(.A1(new_n19259_), .A2(\a[2] ), .Z(new_n19260_));
  OAI21_X1   g19196(.A1(new_n19241_), .A2(new_n19255_), .B(new_n19260_), .ZN(new_n19261_));
  OAI21_X1   g19197(.A1(new_n19234_), .A2(new_n19232_), .B(new_n19235_), .ZN(new_n19262_));
  NAND3_X1   g19198(.A1(new_n19219_), .A2(new_n19225_), .A3(new_n19238_), .ZN(new_n19263_));
  NAND3_X1   g19199(.A1(new_n19262_), .A2(new_n19263_), .A3(new_n17861_), .ZN(new_n19264_));
  INV_X1     g19200(.I(new_n19255_), .ZN(new_n19265_));
  INV_X1     g19201(.I(new_n19260_), .ZN(new_n19266_));
  NAND3_X1   g19202(.A1(new_n19264_), .A2(new_n19265_), .A3(new_n19266_), .ZN(new_n19267_));
  AOI21_X1   g19203(.A1(new_n19261_), .A2(new_n19267_), .B(new_n17852_), .ZN(new_n19268_));
  AOI21_X1   g19204(.A1(new_n19264_), .A2(new_n19265_), .B(new_n19266_), .ZN(new_n19269_));
  NOR3_X1    g19205(.A1(new_n19241_), .A2(new_n19255_), .A3(new_n19260_), .ZN(new_n19270_));
  NOR3_X1    g19206(.A1(new_n19270_), .A2(new_n19269_), .A3(new_n17851_), .ZN(new_n19271_));
  NOR2_X1    g19207(.A1(new_n19271_), .A2(new_n19268_), .ZN(new_n19272_));
  INV_X1     g19208(.I(new_n17843_), .ZN(new_n19273_));
  NOR2_X1    g19209(.A1(new_n19273_), .A2(new_n17844_), .ZN(new_n19274_));
  NOR2_X1    g19210(.A1(new_n17846_), .A2(new_n19274_), .ZN(new_n19275_));
  NOR3_X1    g19211(.A1(new_n19240_), .A2(new_n19231_), .A3(new_n17857_), .ZN(new_n19276_));
  AOI21_X1   g19212(.A1(new_n19262_), .A2(new_n19263_), .B(new_n17858_), .ZN(new_n19277_));
  OAI21_X1   g19213(.A1(new_n19276_), .A2(new_n19277_), .B(new_n17860_), .ZN(new_n19278_));
  NOR2_X1    g19214(.A1(new_n19278_), .A2(new_n19253_), .ZN(new_n19279_));
  NAND3_X1   g19215(.A1(new_n19262_), .A2(new_n19263_), .A3(new_n17858_), .ZN(new_n19280_));
  OAI21_X1   g19216(.A1(new_n19240_), .A2(new_n19231_), .B(new_n17857_), .ZN(new_n19281_));
  NAND2_X1   g19217(.A1(new_n19281_), .A2(new_n19280_), .ZN(new_n19282_));
  AOI21_X1   g19218(.A1(new_n19282_), .A2(new_n17860_), .B(new_n19254_), .ZN(new_n19283_));
  AOI21_X1   g19219(.A1(new_n19262_), .A2(new_n19263_), .B(new_n17857_), .ZN(new_n19284_));
  INV_X1     g19220(.I(new_n19284_), .ZN(new_n19285_));
  NOR3_X1    g19221(.A1(new_n19279_), .A2(new_n19283_), .A3(new_n19285_), .ZN(new_n19286_));
  NAND3_X1   g19222(.A1(new_n19282_), .A2(new_n17860_), .A3(new_n19254_), .ZN(new_n19287_));
  NAND2_X1   g19223(.A1(new_n19278_), .A2(new_n19253_), .ZN(new_n19288_));
  AOI21_X1   g19224(.A1(new_n19288_), .A2(new_n19287_), .B(new_n19284_), .ZN(new_n19289_));
  NOR2_X1    g19225(.A1(new_n19286_), .A2(new_n19289_), .ZN(new_n19290_));
  NOR3_X1    g19226(.A1(new_n19272_), .A2(new_n17850_), .A3(new_n19275_), .ZN(new_n19291_));
  INV_X1     g19227(.I(new_n19291_), .ZN(new_n19292_));
  XOR2_X1    g19228(.A1(new_n16634_), .A2(new_n16680_), .Z(new_n19293_));
  INV_X1     g19229(.I(new_n17837_), .ZN(new_n19294_));
  OAI22_X1   g19230(.A1(new_n17832_), .A2(new_n19294_), .B1(new_n17843_), .B2(new_n17845_), .ZN(new_n19295_));
  OAI22_X1   g19231(.A1(new_n11264_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n11277_), .ZN(new_n19296_));
  NAND2_X1   g19232(.A1(new_n11346_), .A2(new_n9488_), .ZN(new_n19297_));
  AOI21_X1   g19233(.A1(new_n19296_), .A2(new_n19297_), .B(new_n9482_), .ZN(new_n19298_));
  NAND2_X1   g19234(.A1(new_n11757_), .A2(new_n19298_), .ZN(new_n19299_));
  XOR2_X1    g19235(.A1(new_n19299_), .A2(\a[2] ), .Z(new_n19300_));
  XNOR2_X1   g19236(.A1(new_n19295_), .A2(new_n19300_), .ZN(new_n19301_));
  AND2_X2    g19237(.A1(new_n19301_), .A2(new_n19293_), .Z(new_n19302_));
  NOR2_X1    g19238(.A1(new_n19301_), .A2(new_n19293_), .ZN(new_n19303_));
  NOR2_X1    g19239(.A1(new_n19302_), .A2(new_n19303_), .ZN(new_n19304_));
  INV_X1     g19240(.I(new_n19304_), .ZN(new_n19305_));
  OAI21_X1   g19241(.A1(new_n19270_), .A2(new_n19269_), .B(new_n17851_), .ZN(new_n19306_));
  NAND3_X1   g19242(.A1(new_n19261_), .A2(new_n19267_), .A3(new_n17852_), .ZN(new_n19307_));
  NAND2_X1   g19243(.A1(new_n19306_), .A2(new_n19307_), .ZN(new_n19308_));
  NOR2_X1    g19244(.A1(new_n19308_), .A2(new_n17850_), .ZN(new_n19309_));
  INV_X1     g19245(.I(new_n19309_), .ZN(new_n19310_));
  NAND3_X1   g19246(.A1(new_n19288_), .A2(new_n19287_), .A3(new_n19284_), .ZN(new_n19311_));
  OAI21_X1   g19247(.A1(new_n19279_), .A2(new_n19283_), .B(new_n19285_), .ZN(new_n19312_));
  NAND2_X1   g19248(.A1(new_n19312_), .A2(new_n19311_), .ZN(new_n19313_));
  OAI21_X1   g19249(.A1(new_n19271_), .A2(new_n19268_), .B(new_n17850_), .ZN(new_n19314_));
  OAI21_X1   g19250(.A1(new_n19313_), .A2(new_n19314_), .B(new_n19275_), .ZN(new_n19315_));
  AOI21_X1   g19251(.A1(new_n19315_), .A2(new_n19310_), .B(new_n17849_), .ZN(new_n19316_));
  OAI21_X1   g19252(.A1(new_n19316_), .A2(new_n19305_), .B(new_n19292_), .ZN(new_n19317_));
  INV_X1     g19253(.I(new_n17821_), .ZN(new_n19318_));
  NOR2_X1    g19254(.A1(new_n19318_), .A2(new_n17822_), .ZN(new_n19319_));
  NOR2_X1    g19255(.A1(new_n19319_), .A2(new_n17824_), .ZN(new_n19320_));
  INV_X1     g19256(.I(new_n19320_), .ZN(new_n19321_));
  AOI21_X1   g19257(.A1(new_n17827_), .A2(new_n19305_), .B(new_n19321_), .ZN(new_n19322_));
  NAND2_X1   g19258(.A1(new_n17828_), .A2(new_n19304_), .ZN(new_n19323_));
  NAND2_X1   g19259(.A1(new_n19323_), .A2(new_n19321_), .ZN(new_n19324_));
  OAI21_X1   g19260(.A1(new_n19317_), .A2(new_n19322_), .B(new_n19324_), .ZN(new_n19325_));
  NAND2_X1   g19261(.A1(new_n19325_), .A2(new_n17828_), .ZN(new_n19326_));
  NOR2_X1    g19262(.A1(new_n16638_), .A2(new_n16639_), .ZN(new_n19327_));
  XOR2_X1    g19263(.A1(new_n19327_), .A2(new_n16646_), .Z(new_n19328_));
  NOR2_X1    g19264(.A1(new_n19328_), .A2(new_n16708_), .ZN(new_n19329_));
  NOR2_X1    g19265(.A1(new_n16651_), .A2(new_n16647_), .ZN(new_n19330_));
  NOR2_X1    g19266(.A1(new_n19330_), .A2(new_n16637_), .ZN(new_n19331_));
  NOR2_X1    g19267(.A1(new_n19329_), .A2(new_n19331_), .ZN(new_n19332_));
  INV_X1     g19268(.I(new_n17815_), .ZN(new_n19333_));
  OAI22_X1   g19269(.A1(new_n17810_), .A2(new_n19333_), .B1(new_n17821_), .B2(new_n17823_), .ZN(new_n19334_));
  OAI22_X1   g19270(.A1(new_n11353_), .A2(new_n9485_), .B1(new_n9489_), .B2(new_n11697_), .ZN(new_n19335_));
  NAND2_X1   g19271(.A1(new_n11370_), .A2(new_n9503_), .ZN(new_n19336_));
  AOI21_X1   g19272(.A1(new_n19336_), .A2(new_n19335_), .B(new_n9482_), .ZN(new_n19337_));
  NAND2_X1   g19273(.A1(new_n11700_), .A2(new_n19337_), .ZN(new_n19338_));
  XOR2_X1    g19274(.A1(new_n19338_), .A2(\a[2] ), .Z(new_n19339_));
  XNOR2_X1   g19275(.A1(new_n19334_), .A2(new_n19339_), .ZN(new_n19340_));
  AND2_X2    g19276(.A1(new_n19340_), .A2(new_n19332_), .Z(new_n19341_));
  NOR2_X1    g19277(.A1(new_n19340_), .A2(new_n19332_), .ZN(new_n19342_));
  NOR2_X1    g19278(.A1(new_n19341_), .A2(new_n19342_), .ZN(new_n19343_));
  OAI21_X1   g19279(.A1(new_n19325_), .A2(new_n17828_), .B(new_n19343_), .ZN(new_n19344_));
  AOI21_X1   g19280(.A1(new_n16717_), .A2(new_n16720_), .B(new_n16725_), .ZN(new_n19345_));
  NOR2_X1    g19281(.A1(new_n17803_), .A2(new_n19345_), .ZN(new_n19346_));
  OAI21_X1   g19282(.A1(new_n19343_), .A2(new_n17806_), .B(new_n19346_), .ZN(new_n19347_));
  NAND3_X1   g19283(.A1(new_n19344_), .A2(new_n19326_), .A3(new_n19347_), .ZN(new_n19348_));
  INV_X1     g19284(.I(new_n19343_), .ZN(new_n19349_));
  INV_X1     g19285(.I(new_n19346_), .ZN(new_n19350_));
  OAI21_X1   g19286(.A1(new_n19349_), .A2(new_n17807_), .B(new_n19350_), .ZN(new_n19351_));
  AOI21_X1   g19287(.A1(new_n19348_), .A2(new_n19351_), .B(new_n17807_), .ZN(new_n19352_));
  XOR2_X1    g19288(.A1(new_n16735_), .A2(new_n15885_), .Z(new_n19353_));
  NOR2_X1    g19289(.A1(new_n19353_), .A2(new_n17028_), .ZN(new_n19354_));
  AND2_X2    g19290(.A1(new_n19353_), .A2(new_n17028_), .Z(new_n19355_));
  NOR2_X1    g19291(.A1(new_n19355_), .A2(new_n19354_), .ZN(new_n19356_));
  NAND3_X1   g19292(.A1(new_n19348_), .A2(new_n17807_), .A3(new_n19351_), .ZN(new_n19357_));
  AOI21_X1   g19293(.A1(new_n19356_), .A2(new_n19357_), .B(new_n19352_), .ZN(new_n19358_));
  INV_X1     g19294(.I(new_n19356_), .ZN(new_n19359_));
  OAI21_X1   g19295(.A1(new_n16844_), .A2(new_n16843_), .B(new_n16839_), .ZN(new_n19360_));
  NAND3_X1   g19296(.A1(new_n16834_), .A2(new_n16838_), .A3(new_n16845_), .ZN(new_n19361_));
  AOI21_X1   g19297(.A1(new_n19360_), .A2(new_n19361_), .B(new_n16736_), .ZN(new_n19362_));
  AOI21_X1   g19298(.A1(new_n16840_), .A2(new_n16846_), .B(new_n17042_), .ZN(new_n19363_));
  NOR2_X1    g19299(.A1(new_n19362_), .A2(new_n19363_), .ZN(new_n19364_));
  INV_X1     g19300(.I(new_n19364_), .ZN(new_n19365_));
  AOI21_X1   g19301(.A1(new_n19359_), .A2(new_n17802_), .B(new_n19365_), .ZN(new_n19366_));
  INV_X1     g19302(.I(new_n19366_), .ZN(new_n19367_));
  AOI21_X1   g19303(.A1(new_n19356_), .A2(new_n17801_), .B(new_n19364_), .ZN(new_n19368_));
  AOI21_X1   g19304(.A1(new_n19358_), .A2(new_n19367_), .B(new_n19368_), .ZN(new_n19369_));
  AOI21_X1   g19305(.A1(new_n19369_), .A2(new_n17802_), .B(new_n17798_), .ZN(new_n19370_));
  XOR2_X1    g19306(.A1(new_n17122_), .A2(new_n17165_), .Z(new_n19371_));
  NOR2_X1    g19307(.A1(new_n19371_), .A2(new_n17183_), .ZN(new_n19372_));
  XOR2_X1    g19308(.A1(new_n17122_), .A2(new_n17166_), .Z(new_n19373_));
  NOR2_X1    g19309(.A1(new_n19373_), .A2(new_n17067_), .ZN(new_n19374_));
  NOR2_X1    g19310(.A1(new_n19372_), .A2(new_n19374_), .ZN(new_n19375_));
  OAI21_X1   g19311(.A1(new_n19369_), .A2(new_n17802_), .B(new_n17798_), .ZN(new_n19376_));
  AOI21_X1   g19312(.A1(new_n19375_), .A2(new_n19376_), .B(new_n19370_), .ZN(new_n19377_));
  NOR2_X1    g19313(.A1(new_n17185_), .A2(new_n17186_), .ZN(new_n19378_));
  NAND2_X1   g19314(.A1(new_n17067_), .A2(new_n17122_), .ZN(new_n19379_));
  XOR2_X1    g19315(.A1(new_n19379_), .A2(new_n19378_), .Z(new_n19380_));
  XOR2_X1    g19316(.A1(new_n17067_), .A2(new_n17122_), .Z(new_n19381_));
  NAND2_X1   g19317(.A1(new_n19381_), .A2(new_n17166_), .ZN(new_n19382_));
  NOR2_X1    g19318(.A1(new_n19380_), .A2(new_n19382_), .ZN(new_n19383_));
  AND2_X2    g19319(.A1(new_n19380_), .A2(new_n19382_), .Z(new_n19384_));
  NOR2_X1    g19320(.A1(new_n19384_), .A2(new_n19383_), .ZN(new_n19385_));
  INV_X1     g19321(.I(new_n19385_), .ZN(new_n19386_));
  OAI21_X1   g19322(.A1(new_n17793_), .A2(new_n19375_), .B(new_n19385_), .ZN(new_n19387_));
  NAND2_X1   g19323(.A1(new_n17793_), .A2(new_n19375_), .ZN(new_n19388_));
  AOI22_X1   g19324(.A1(new_n19377_), .A2(new_n19387_), .B1(new_n19386_), .B2(new_n19388_), .ZN(new_n19389_));
  NOR2_X1    g19325(.A1(new_n19389_), .A2(new_n17794_), .ZN(new_n19390_));
  NOR2_X1    g19326(.A1(new_n17222_), .A2(new_n17201_), .ZN(new_n19391_));
  AOI21_X1   g19327(.A1(new_n17199_), .A2(new_n17179_), .B(new_n17223_), .ZN(new_n19392_));
  NOR2_X1    g19328(.A1(new_n19391_), .A2(new_n19392_), .ZN(new_n19393_));
  INV_X1     g19329(.I(new_n19393_), .ZN(new_n19394_));
  AOI21_X1   g19330(.A1(new_n19389_), .A2(new_n17794_), .B(new_n19394_), .ZN(new_n19395_));
  NOR2_X1    g19331(.A1(new_n19395_), .A2(new_n19390_), .ZN(new_n19396_));
  NOR2_X1    g19332(.A1(new_n17224_), .A2(new_n17217_), .ZN(new_n19397_));
  AOI21_X1   g19333(.A1(new_n17202_), .A2(new_n13964_), .B(new_n13767_), .ZN(new_n19398_));
  OR2_X2     g19334(.A1(new_n19397_), .A2(new_n19398_), .Z(new_n19399_));
  INV_X1     g19335(.I(new_n19399_), .ZN(new_n19400_));
  OAI21_X1   g19336(.A1(new_n17789_), .A2(new_n19393_), .B(new_n19400_), .ZN(new_n19401_));
  AOI21_X1   g19337(.A1(new_n17789_), .A2(new_n19393_), .B(new_n19400_), .ZN(new_n19402_));
  AOI21_X1   g19338(.A1(new_n19396_), .A2(new_n19401_), .B(new_n19402_), .ZN(new_n19403_));
  NOR2_X1    g19339(.A1(new_n19403_), .A2(new_n17790_), .ZN(new_n19404_));
  OR2_X2     g19340(.A1(new_n17243_), .A2(new_n17233_), .Z(new_n19405_));
  NAND2_X1   g19341(.A1(new_n17243_), .A2(new_n17233_), .ZN(new_n19406_));
  NAND2_X1   g19342(.A1(new_n19405_), .A2(new_n19406_), .ZN(new_n19407_));
  AOI21_X1   g19343(.A1(new_n19403_), .A2(new_n17790_), .B(new_n19407_), .ZN(new_n19408_));
  NOR2_X1    g19344(.A1(new_n19408_), .A2(new_n19404_), .ZN(new_n19409_));
  INV_X1     g19345(.I(new_n19407_), .ZN(new_n19410_));
  AOI21_X1   g19346(.A1(new_n17234_), .A2(new_n13256_), .B(new_n12731_), .ZN(new_n19411_));
  NOR2_X1    g19347(.A1(new_n17245_), .A2(new_n19411_), .ZN(new_n19412_));
  OAI21_X1   g19348(.A1(new_n17787_), .A2(new_n19410_), .B(new_n19412_), .ZN(new_n19413_));
  NAND2_X1   g19349(.A1(new_n19409_), .A2(new_n19413_), .ZN(new_n19414_));
  INV_X1     g19350(.I(new_n19412_), .ZN(new_n19415_));
  NAND2_X1   g19351(.A1(new_n17787_), .A2(new_n19410_), .ZN(new_n19416_));
  NAND2_X1   g19352(.A1(new_n19416_), .A2(new_n19415_), .ZN(new_n19417_));
  NAND2_X1   g19353(.A1(new_n19414_), .A2(new_n19417_), .ZN(new_n19418_));
  NAND2_X1   g19354(.A1(new_n19418_), .A2(new_n17787_), .ZN(new_n19419_));
  XOR2_X1    g19355(.A1(new_n17413_), .A2(new_n17339_), .Z(new_n19420_));
  NOR2_X1    g19356(.A1(new_n17709_), .A2(new_n19420_), .ZN(new_n19421_));
  AOI21_X1   g19357(.A1(new_n17416_), .A2(new_n17710_), .B(new_n17338_), .ZN(new_n19422_));
  NOR2_X1    g19358(.A1(new_n19422_), .A2(new_n19421_), .ZN(new_n19423_));
  OAI21_X1   g19359(.A1(new_n19418_), .A2(new_n17787_), .B(new_n19423_), .ZN(new_n19424_));
  XNOR2_X1   g19360(.A1(new_n17504_), .A2(new_n17501_), .ZN(new_n19425_));
  NOR2_X1    g19361(.A1(new_n17419_), .A2(new_n19425_), .ZN(new_n19426_));
  AOI21_X1   g19362(.A1(new_n17712_), .A2(new_n17508_), .B(new_n17711_), .ZN(new_n19427_));
  NOR2_X1    g19363(.A1(new_n19427_), .A2(new_n19426_), .ZN(new_n19428_));
  OAI21_X1   g19364(.A1(new_n17784_), .A2(new_n19423_), .B(new_n19428_), .ZN(new_n19429_));
  AND3_X2    g19365(.A1(new_n19424_), .A2(new_n19419_), .A3(new_n19429_), .Z(new_n19430_));
  AOI21_X1   g19366(.A1(new_n17784_), .A2(new_n19423_), .B(new_n19428_), .ZN(new_n19431_));
  OAI21_X1   g19367(.A1(new_n19430_), .A2(new_n19431_), .B(new_n17784_), .ZN(new_n19432_));
  XOR2_X1    g19368(.A1(new_n17614_), .A2(new_n17667_), .Z(new_n19433_));
  NOR2_X1    g19369(.A1(new_n17574_), .A2(new_n19433_), .ZN(new_n19434_));
  XNOR2_X1   g19370(.A1(new_n17614_), .A2(new_n17667_), .ZN(new_n19435_));
  NOR2_X1    g19371(.A1(new_n17714_), .A2(new_n19435_), .ZN(new_n19436_));
  NOR2_X1    g19372(.A1(new_n19436_), .A2(new_n19434_), .ZN(new_n19437_));
  INV_X1     g19373(.I(new_n17784_), .ZN(new_n19438_));
  INV_X1     g19374(.I(new_n17787_), .ZN(new_n19439_));
  AOI22_X1   g19375(.A1(new_n19409_), .A2(new_n19413_), .B1(new_n19415_), .B2(new_n19416_), .ZN(new_n19440_));
  NOR2_X1    g19376(.A1(new_n19440_), .A2(new_n19439_), .ZN(new_n19441_));
  INV_X1     g19377(.I(new_n19423_), .ZN(new_n19442_));
  AOI21_X1   g19378(.A1(new_n19440_), .A2(new_n19439_), .B(new_n19442_), .ZN(new_n19443_));
  NOR2_X1    g19379(.A1(new_n19443_), .A2(new_n19441_), .ZN(new_n19444_));
  NAND2_X1   g19380(.A1(new_n19444_), .A2(new_n19429_), .ZN(new_n19445_));
  INV_X1     g19381(.I(new_n19431_), .ZN(new_n19446_));
  NAND3_X1   g19382(.A1(new_n19445_), .A2(new_n19438_), .A3(new_n19446_), .ZN(new_n19447_));
  NAND2_X1   g19383(.A1(new_n19447_), .A2(new_n19437_), .ZN(new_n19448_));
  NAND3_X1   g19384(.A1(new_n17714_), .A2(new_n17715_), .A3(new_n17664_), .ZN(new_n19449_));
  OAI21_X1   g19385(.A1(new_n17574_), .A2(new_n17614_), .B(new_n17665_), .ZN(new_n19450_));
  NAND2_X1   g19386(.A1(new_n19450_), .A2(new_n19449_), .ZN(new_n19451_));
  NOR2_X1    g19387(.A1(new_n17714_), .A2(new_n17614_), .ZN(new_n19452_));
  NOR2_X1    g19388(.A1(new_n17574_), .A2(new_n17715_), .ZN(new_n19453_));
  OAI21_X1   g19389(.A1(new_n19452_), .A2(new_n19453_), .B(new_n17667_), .ZN(new_n19454_));
  NOR2_X1    g19390(.A1(new_n19454_), .A2(new_n19451_), .ZN(new_n19455_));
  NOR3_X1    g19391(.A1(new_n17574_), .A2(new_n17614_), .A3(new_n17665_), .ZN(new_n19456_));
  AOI21_X1   g19392(.A1(new_n17714_), .A2(new_n17715_), .B(new_n17664_), .ZN(new_n19457_));
  NOR2_X1    g19393(.A1(new_n19457_), .A2(new_n19456_), .ZN(new_n19458_));
  NAND2_X1   g19394(.A1(new_n17574_), .A2(new_n17715_), .ZN(new_n19459_));
  NAND2_X1   g19395(.A1(new_n17714_), .A2(new_n17614_), .ZN(new_n19460_));
  AOI21_X1   g19396(.A1(new_n19460_), .A2(new_n19459_), .B(new_n17668_), .ZN(new_n19461_));
  NOR2_X1    g19397(.A1(new_n19458_), .A2(new_n19461_), .ZN(new_n19462_));
  NOR2_X1    g19398(.A1(new_n19462_), .A2(new_n19455_), .ZN(new_n19463_));
  AOI21_X1   g19399(.A1(new_n17776_), .A2(new_n17777_), .B(new_n17778_), .ZN(new_n19464_));
  NOR3_X1    g19400(.A1(new_n17720_), .A2(new_n17719_), .A3(new_n17722_), .ZN(new_n19465_));
  INV_X1     g19401(.I(new_n19437_), .ZN(new_n19466_));
  OAI21_X1   g19402(.A1(new_n19465_), .A2(new_n19464_), .B(new_n19466_), .ZN(new_n19467_));
  NAND2_X1   g19403(.A1(new_n19467_), .A2(new_n19463_), .ZN(new_n19468_));
  NAND3_X1   g19404(.A1(new_n19448_), .A2(new_n19468_), .A3(new_n19432_), .ZN(new_n19469_));
  NAND2_X1   g19405(.A1(new_n19458_), .A2(new_n19461_), .ZN(new_n19470_));
  NAND2_X1   g19406(.A1(new_n19454_), .A2(new_n19451_), .ZN(new_n19471_));
  NAND2_X1   g19407(.A1(new_n19470_), .A2(new_n19471_), .ZN(new_n19472_));
  OAI21_X1   g19408(.A1(new_n17780_), .A2(new_n19466_), .B(new_n19472_), .ZN(new_n19473_));
  AOI21_X1   g19409(.A1(new_n19469_), .A2(new_n19473_), .B(new_n17780_), .ZN(new_n19474_));
  INV_X1     g19410(.I(new_n17780_), .ZN(new_n19475_));
  AOI21_X1   g19411(.A1(new_n19444_), .A2(new_n19429_), .B(new_n19431_), .ZN(new_n19476_));
  NOR2_X1    g19412(.A1(new_n19476_), .A2(new_n19438_), .ZN(new_n19477_));
  AOI21_X1   g19413(.A1(new_n19476_), .A2(new_n19438_), .B(new_n19466_), .ZN(new_n19478_));
  AOI21_X1   g19414(.A1(new_n17780_), .A2(new_n19466_), .B(new_n19472_), .ZN(new_n19479_));
  NOR3_X1    g19415(.A1(new_n19479_), .A2(new_n19477_), .A3(new_n19478_), .ZN(new_n19480_));
  INV_X1     g19416(.I(new_n19473_), .ZN(new_n19481_));
  NOR3_X1    g19417(.A1(new_n19480_), .A2(new_n19475_), .A3(new_n19481_), .ZN(new_n19482_));
  NOR2_X1    g19418(.A1(new_n19474_), .A2(new_n17775_), .ZN(new_n19483_));
  INV_X1     g19419(.I(new_n17775_), .ZN(new_n19484_));
  OAI21_X1   g19420(.A1(new_n19480_), .A2(new_n19481_), .B(new_n19475_), .ZN(new_n19485_));
  AOI21_X1   g19421(.A1(new_n19482_), .A2(new_n19485_), .B(new_n19484_), .ZN(new_n19486_));
  NOR2_X1    g19422(.A1(new_n19486_), .A2(new_n19483_), .ZN(new_n19487_));
  NOR2_X1    g19423(.A1(new_n19464_), .A2(new_n17704_), .ZN(new_n19488_));
  INV_X1     g19424(.I(new_n17754_), .ZN(new_n19489_));
  NOR3_X1    g19425(.A1(new_n19488_), .A2(new_n17746_), .A3(new_n19489_), .ZN(new_n19490_));
  AOI21_X1   g19426(.A1(new_n17724_), .A2(new_n17747_), .B(new_n17754_), .ZN(new_n19491_));
  NOR2_X1    g19427(.A1(new_n19490_), .A2(new_n19491_), .ZN(new_n19492_));
  NAND2_X1   g19428(.A1(new_n19488_), .A2(new_n17747_), .ZN(new_n19493_));
  NAND2_X1   g19429(.A1(new_n17724_), .A2(new_n17746_), .ZN(new_n19494_));
  AOI21_X1   g19430(.A1(new_n19494_), .A2(new_n19493_), .B(new_n17771_), .ZN(new_n19495_));
  NAND2_X1   g19431(.A1(new_n19492_), .A2(new_n19495_), .ZN(new_n19496_));
  NAND3_X1   g19432(.A1(new_n17724_), .A2(new_n17747_), .A3(new_n17754_), .ZN(new_n19497_));
  OAI21_X1   g19433(.A1(new_n19488_), .A2(new_n17746_), .B(new_n19489_), .ZN(new_n19498_));
  NAND2_X1   g19434(.A1(new_n19498_), .A2(new_n19497_), .ZN(new_n19499_));
  NOR2_X1    g19435(.A1(new_n17724_), .A2(new_n17746_), .ZN(new_n19500_));
  NOR2_X1    g19436(.A1(new_n19488_), .A2(new_n17747_), .ZN(new_n19501_));
  OAI21_X1   g19437(.A1(new_n19500_), .A2(new_n19501_), .B(new_n17756_), .ZN(new_n19502_));
  NAND2_X1   g19438(.A1(new_n19502_), .A2(new_n19499_), .ZN(new_n19503_));
  AOI21_X1   g19439(.A1(new_n19496_), .A2(new_n19503_), .B(new_n19484_), .ZN(new_n19504_));
  NOR2_X1    g19440(.A1(new_n19502_), .A2(new_n19499_), .ZN(new_n19505_));
  NOR2_X1    g19441(.A1(new_n19492_), .A2(new_n19495_), .ZN(new_n19506_));
  NOR3_X1    g19442(.A1(new_n19506_), .A2(new_n19505_), .A3(new_n17775_), .ZN(new_n19507_));
  NOR2_X1    g19443(.A1(new_n19504_), .A2(new_n19507_), .ZN(new_n19508_));
  NOR3_X1    g19444(.A1(new_n19487_), .A2(new_n19508_), .A3(new_n17770_), .ZN(new_n19509_));
  AOI21_X1   g19445(.A1(new_n17768_), .A2(new_n17762_), .B(new_n17765_), .ZN(new_n19510_));
  NOR3_X1    g19446(.A1(new_n17763_), .A2(new_n11689_), .A3(new_n17761_), .ZN(new_n19511_));
  NOR2_X1    g19447(.A1(new_n19511_), .A2(new_n19510_), .ZN(new_n19512_));
  NAND2_X1   g19448(.A1(new_n19485_), .A2(new_n19484_), .ZN(new_n19513_));
  NAND2_X1   g19449(.A1(new_n19469_), .A2(new_n19473_), .ZN(new_n19514_));
  OAI21_X1   g19450(.A1(new_n19514_), .A2(new_n19475_), .B(new_n17775_), .ZN(new_n19515_));
  NAND2_X1   g19451(.A1(new_n19513_), .A2(new_n19515_), .ZN(new_n19516_));
  OAI21_X1   g19452(.A1(new_n19506_), .A2(new_n19505_), .B(new_n17775_), .ZN(new_n19517_));
  NAND3_X1   g19453(.A1(new_n19496_), .A2(new_n19503_), .A3(new_n19484_), .ZN(new_n19518_));
  NAND2_X1   g19454(.A1(new_n19517_), .A2(new_n19518_), .ZN(new_n19519_));
  AOI21_X1   g19455(.A1(new_n19516_), .A2(new_n19519_), .B(new_n19512_), .ZN(new_n19520_));
  NOR2_X1    g19456(.A1(new_n19509_), .A2(new_n19520_), .ZN(new_n19521_));
  NOR2_X1    g19457(.A1(new_n19506_), .A2(new_n19505_), .ZN(new_n19522_));
  OAI22_X1   g19458(.A1(new_n19522_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n17775_), .ZN(new_n19523_));
  NAND2_X1   g19459(.A1(new_n17770_), .A2(new_n6838_), .ZN(new_n19524_));
  AOI21_X1   g19460(.A1(new_n19524_), .A2(new_n19523_), .B(new_n6836_), .ZN(new_n19525_));
  NAND2_X1   g19461(.A1(new_n19521_), .A2(new_n19525_), .ZN(new_n19526_));
  XOR2_X1    g19462(.A1(new_n19526_), .A2(new_n65_), .Z(new_n19527_));
  NAND2_X1   g19463(.A1(new_n19348_), .A2(new_n19351_), .ZN(new_n19528_));
  OAI21_X1   g19464(.A1(new_n19528_), .A2(new_n17806_), .B(new_n19356_), .ZN(new_n19529_));
  INV_X1     g19465(.I(new_n19529_), .ZN(new_n19530_));
  NOR2_X1    g19466(.A1(new_n19352_), .A2(new_n19356_), .ZN(new_n19532_));
  OAI21_X1   g19467(.A1(new_n19530_), .A2(new_n19532_), .B(new_n19365_), .ZN(new_n19533_));
  NOR3_X1    g19468(.A1(new_n19528_), .A2(new_n17806_), .A3(new_n19359_), .ZN(new_n19534_));
  NAND2_X1   g19469(.A1(new_n19352_), .A2(new_n19359_), .ZN(new_n19535_));
  INV_X1     g19470(.I(new_n19535_), .ZN(new_n19536_));
  OAI21_X1   g19471(.A1(new_n19536_), .A2(new_n19534_), .B(new_n19364_), .ZN(new_n19537_));
  NAND2_X1   g19472(.A1(new_n19537_), .A2(new_n19533_), .ZN(new_n19538_));
  OAI22_X1   g19473(.A1(new_n19356_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n17806_), .ZN(new_n19539_));
  NAND2_X1   g19474(.A1(new_n19365_), .A2(new_n3312_), .ZN(new_n19540_));
  AOI21_X1   g19475(.A1(new_n19539_), .A2(new_n19540_), .B(new_n3302_), .ZN(new_n19541_));
  NAND2_X1   g19476(.A1(new_n19538_), .A2(new_n19541_), .ZN(new_n19542_));
  XOR2_X1    g19477(.A1(new_n19542_), .A2(new_n84_), .Z(new_n19543_));
  NOR2_X1    g19478(.A1(new_n19313_), .A2(new_n2734_), .ZN(new_n19544_));
  INV_X1     g19479(.I(new_n19275_), .ZN(new_n19545_));
  NAND3_X1   g19480(.A1(new_n19312_), .A2(new_n19311_), .A3(new_n19545_), .ZN(new_n19546_));
  OAI21_X1   g19481(.A1(new_n19271_), .A2(new_n19268_), .B(new_n19275_), .ZN(new_n19547_));
  NAND3_X1   g19482(.A1(new_n19306_), .A2(new_n19307_), .A3(new_n19545_), .ZN(new_n19548_));
  NAND2_X1   g19483(.A1(new_n19547_), .A2(new_n19548_), .ZN(new_n19549_));
  NAND3_X1   g19484(.A1(new_n19549_), .A2(new_n19546_), .A3(new_n17849_), .ZN(new_n19550_));
  AOI21_X1   g19485(.A1(new_n19549_), .A2(new_n19546_), .B(new_n17849_), .ZN(new_n19551_));
  INV_X1     g19486(.I(new_n19551_), .ZN(new_n19552_));
  NAND2_X1   g19487(.A1(new_n19552_), .A2(new_n19550_), .ZN(new_n19553_));
  OAI22_X1   g19488(.A1(new_n19272_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n19275_), .ZN(new_n19554_));
  NAND2_X1   g19489(.A1(new_n17850_), .A2(new_n3317_), .ZN(new_n19555_));
  AOI21_X1   g19490(.A1(new_n19554_), .A2(new_n19555_), .B(new_n3260_), .ZN(new_n19556_));
  NAND3_X1   g19491(.A1(new_n19553_), .A2(new_n72_), .A3(new_n19556_), .ZN(new_n19557_));
  AOI21_X1   g19492(.A1(new_n19553_), .A2(new_n19556_), .B(new_n72_), .ZN(new_n19558_));
  INV_X1     g19493(.I(new_n19558_), .ZN(new_n19559_));
  AOI21_X1   g19494(.A1(new_n19559_), .A2(new_n19557_), .B(new_n19544_), .ZN(new_n19560_));
  NAND3_X1   g19495(.A1(new_n19313_), .A2(new_n19308_), .A3(new_n19275_), .ZN(new_n19561_));
  AOI21_X1   g19496(.A1(new_n19313_), .A2(new_n19308_), .B(new_n19275_), .ZN(new_n19562_));
  INV_X1     g19497(.I(new_n19562_), .ZN(new_n19563_));
  NAND2_X1   g19498(.A1(new_n19563_), .A2(new_n19561_), .ZN(new_n19564_));
  OAI22_X1   g19499(.A1(new_n19313_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n19272_), .ZN(new_n19565_));
  NAND2_X1   g19500(.A1(new_n19545_), .A2(new_n3317_), .ZN(new_n19566_));
  NAND2_X1   g19501(.A1(new_n19565_), .A2(new_n19566_), .ZN(new_n19567_));
  NAND3_X1   g19502(.A1(new_n19564_), .A2(new_n3259_), .A3(new_n19567_), .ZN(new_n19568_));
  NAND2_X1   g19503(.A1(new_n19568_), .A2(new_n72_), .ZN(new_n19569_));
  INV_X1     g19504(.I(new_n19561_), .ZN(new_n19570_));
  NOR2_X1    g19505(.A1(new_n19570_), .A2(new_n19562_), .ZN(new_n19571_));
  NAND2_X1   g19506(.A1(new_n19567_), .A2(new_n3259_), .ZN(new_n19572_));
  NOR2_X1    g19507(.A1(new_n19572_), .A2(new_n19571_), .ZN(new_n19573_));
  NAND2_X1   g19508(.A1(new_n19573_), .A2(\a[26] ), .ZN(new_n19574_));
  NOR2_X1    g19509(.A1(new_n19290_), .A2(new_n19308_), .ZN(new_n19575_));
  NOR2_X1    g19510(.A1(new_n19313_), .A2(new_n19272_), .ZN(new_n19576_));
  NOR2_X1    g19511(.A1(new_n19575_), .A2(new_n19576_), .ZN(new_n19577_));
  NAND2_X1   g19512(.A1(new_n19290_), .A2(new_n3323_), .ZN(new_n19578_));
  NOR2_X1    g19513(.A1(new_n3257_), .A2(new_n3258_), .ZN(new_n19580_));
  NAND3_X1   g19514(.A1(new_n19577_), .A2(new_n19578_), .A3(new_n19580_), .ZN(new_n19581_));
  NOR2_X1    g19515(.A1(new_n19313_), .A2(new_n3257_), .ZN(new_n19582_));
  NOR3_X1    g19516(.A1(new_n19581_), .A2(new_n72_), .A3(new_n19582_), .ZN(new_n19583_));
  NAND3_X1   g19517(.A1(new_n19574_), .A2(new_n19569_), .A3(new_n19583_), .ZN(new_n19584_));
  NAND3_X1   g19518(.A1(new_n19559_), .A2(new_n19544_), .A3(new_n19557_), .ZN(new_n19585_));
  AOI21_X1   g19519(.A1(new_n19584_), .A2(new_n19585_), .B(new_n19560_), .ZN(new_n19586_));
  NAND2_X1   g19520(.A1(new_n19290_), .A2(new_n3275_), .ZN(new_n19587_));
  NOR2_X1    g19521(.A1(new_n2735_), .A2(new_n2734_), .ZN(new_n19588_));
  NAND3_X1   g19522(.A1(new_n19577_), .A2(new_n19587_), .A3(new_n19588_), .ZN(new_n19589_));
  NOR2_X1    g19523(.A1(new_n19589_), .A2(\a[29] ), .ZN(new_n19590_));
  NAND2_X1   g19524(.A1(new_n19313_), .A2(new_n19272_), .ZN(new_n19591_));
  NAND2_X1   g19525(.A1(new_n19290_), .A2(new_n19308_), .ZN(new_n19592_));
  NAND2_X1   g19526(.A1(new_n19592_), .A2(new_n19591_), .ZN(new_n19593_));
  NAND2_X1   g19527(.A1(new_n19587_), .A2(new_n19588_), .ZN(new_n19594_));
  NOR2_X1    g19528(.A1(new_n19593_), .A2(new_n19594_), .ZN(new_n19595_));
  NOR2_X1    g19529(.A1(new_n19595_), .A2(new_n74_), .ZN(new_n19596_));
  NOR2_X1    g19530(.A1(new_n19544_), .A2(new_n74_), .ZN(new_n19597_));
  NOR3_X1    g19531(.A1(new_n19590_), .A2(new_n19596_), .A3(new_n19597_), .ZN(new_n19598_));
  NOR3_X1    g19532(.A1(new_n19595_), .A2(new_n74_), .A3(new_n19544_), .ZN(new_n19599_));
  NOR2_X1    g19533(.A1(new_n19598_), .A2(new_n19599_), .ZN(new_n19600_));
  OAI21_X1   g19534(.A1(new_n19316_), .A2(new_n19291_), .B(new_n19305_), .ZN(new_n19601_));
  AOI21_X1   g19535(.A1(new_n19308_), .A2(new_n19545_), .B(new_n17850_), .ZN(new_n19602_));
  AOI21_X1   g19536(.A1(new_n19306_), .A2(new_n19307_), .B(new_n17849_), .ZN(new_n19603_));
  AOI21_X1   g19537(.A1(new_n19290_), .A2(new_n19603_), .B(new_n19545_), .ZN(new_n19604_));
  NOR3_X1    g19538(.A1(new_n19604_), .A2(new_n17849_), .A3(new_n19309_), .ZN(new_n19605_));
  OAI21_X1   g19539(.A1(new_n19605_), .A2(new_n19602_), .B(new_n19304_), .ZN(new_n19606_));
  NAND2_X1   g19540(.A1(new_n19606_), .A2(new_n19601_), .ZN(new_n19607_));
  AOI22_X1   g19541(.A1(new_n17850_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n19545_), .ZN(new_n19608_));
  AOI21_X1   g19542(.A1(new_n19305_), .A2(new_n3317_), .B(new_n19608_), .ZN(new_n19609_));
  NOR2_X1    g19543(.A1(new_n19609_), .A2(new_n3260_), .ZN(new_n19610_));
  NAND2_X1   g19544(.A1(new_n19607_), .A2(new_n19610_), .ZN(new_n19611_));
  NOR2_X1    g19545(.A1(new_n19611_), .A2(\a[26] ), .ZN(new_n19612_));
  OAI21_X1   g19546(.A1(new_n19604_), .A2(new_n19309_), .B(new_n17850_), .ZN(new_n19613_));
  AOI21_X1   g19547(.A1(new_n19613_), .A2(new_n19292_), .B(new_n19304_), .ZN(new_n19614_));
  INV_X1     g19548(.I(new_n19602_), .ZN(new_n19615_));
  NAND3_X1   g19549(.A1(new_n19315_), .A2(new_n17850_), .A3(new_n19310_), .ZN(new_n19616_));
  AOI21_X1   g19550(.A1(new_n19616_), .A2(new_n19615_), .B(new_n19305_), .ZN(new_n19617_));
  NOR2_X1    g19551(.A1(new_n19614_), .A2(new_n19617_), .ZN(new_n19618_));
  NOR3_X1    g19552(.A1(new_n19618_), .A2(new_n3260_), .A3(new_n19609_), .ZN(new_n19619_));
  NOR2_X1    g19553(.A1(new_n19619_), .A2(new_n72_), .ZN(new_n19620_));
  NOR3_X1    g19554(.A1(new_n19620_), .A2(new_n19612_), .A3(new_n19600_), .ZN(new_n19621_));
  OAI21_X1   g19555(.A1(new_n19620_), .A2(new_n19612_), .B(new_n19600_), .ZN(new_n19622_));
  OAI21_X1   g19556(.A1(new_n19586_), .A2(new_n19621_), .B(new_n19622_), .ZN(new_n19623_));
  OAI22_X1   g19557(.A1(new_n19313_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n19272_), .ZN(new_n19624_));
  OAI21_X1   g19558(.A1(new_n3175_), .A2(new_n19275_), .B(new_n19624_), .ZN(new_n19625_));
  NAND3_X1   g19559(.A1(new_n19564_), .A2(new_n19625_), .A3(new_n2736_), .ZN(new_n19626_));
  NAND2_X1   g19560(.A1(new_n19626_), .A2(new_n74_), .ZN(new_n19627_));
  NOR2_X1    g19561(.A1(new_n19571_), .A2(new_n2737_), .ZN(new_n19628_));
  NAND3_X1   g19562(.A1(new_n19628_), .A2(\a[29] ), .A3(new_n19625_), .ZN(new_n19629_));
  INV_X1     g19563(.I(new_n19544_), .ZN(new_n19630_));
  NAND3_X1   g19564(.A1(new_n19595_), .A2(\a[29] ), .A3(new_n19630_), .ZN(new_n19631_));
  NAND3_X1   g19565(.A1(new_n19627_), .A2(new_n19629_), .A3(new_n19631_), .ZN(new_n19632_));
  AOI21_X1   g19566(.A1(new_n19628_), .A2(new_n19625_), .B(\a[29] ), .ZN(new_n19633_));
  NOR2_X1    g19567(.A1(new_n19626_), .A2(new_n74_), .ZN(new_n19634_));
  NOR3_X1    g19568(.A1(new_n19589_), .A2(new_n74_), .A3(new_n19544_), .ZN(new_n19635_));
  OAI21_X1   g19569(.A1(new_n19634_), .A2(new_n19633_), .B(new_n19635_), .ZN(new_n19636_));
  NAND2_X1   g19570(.A1(new_n19636_), .A2(new_n19632_), .ZN(new_n19637_));
  NAND3_X1   g19571(.A1(new_n19603_), .A2(new_n19312_), .A3(new_n19311_), .ZN(new_n19638_));
  AOI21_X1   g19572(.A1(new_n19638_), .A2(new_n19275_), .B(new_n19309_), .ZN(new_n19639_));
  OAI21_X1   g19573(.A1(new_n19639_), .A2(new_n17849_), .B(new_n19304_), .ZN(new_n19640_));
  NOR2_X1    g19574(.A1(new_n19291_), .A2(new_n19304_), .ZN(new_n19641_));
  INV_X1     g19575(.I(new_n19641_), .ZN(new_n19642_));
  AND2_X2    g19576(.A1(new_n19640_), .A2(new_n19642_), .Z(new_n19643_));
  NOR3_X1    g19577(.A1(new_n19639_), .A2(new_n17849_), .A3(new_n19305_), .ZN(new_n19644_));
  NOR2_X1    g19578(.A1(new_n19292_), .A2(new_n19304_), .ZN(new_n19645_));
  OAI21_X1   g19579(.A1(new_n19644_), .A2(new_n19645_), .B(new_n19320_), .ZN(new_n19646_));
  OAI21_X1   g19580(.A1(new_n19643_), .A2(new_n19320_), .B(new_n19646_), .ZN(new_n19647_));
  OAI22_X1   g19581(.A1(new_n19304_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n17849_), .ZN(new_n19648_));
  NAND2_X1   g19582(.A1(new_n19321_), .A2(new_n3317_), .ZN(new_n19649_));
  AOI21_X1   g19583(.A1(new_n19648_), .A2(new_n19649_), .B(new_n3260_), .ZN(new_n19650_));
  NAND3_X1   g19584(.A1(new_n19647_), .A2(new_n72_), .A3(new_n19650_), .ZN(new_n19651_));
  AOI21_X1   g19585(.A1(new_n19647_), .A2(new_n19650_), .B(new_n72_), .ZN(new_n19652_));
  INV_X1     g19586(.I(new_n19652_), .ZN(new_n19653_));
  NAND3_X1   g19587(.A1(new_n19653_), .A2(new_n19637_), .A3(new_n19651_), .ZN(new_n19654_));
  AOI21_X1   g19588(.A1(new_n19653_), .A2(new_n19651_), .B(new_n19637_), .ZN(new_n19655_));
  AOI21_X1   g19589(.A1(new_n19623_), .A2(new_n19654_), .B(new_n19655_), .ZN(new_n19656_));
  NAND3_X1   g19590(.A1(new_n19627_), .A2(new_n19629_), .A3(new_n19635_), .ZN(new_n19657_));
  OAI22_X1   g19591(.A1(new_n19272_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n19275_), .ZN(new_n19658_));
  NAND2_X1   g19592(.A1(new_n17850_), .A2(new_n2750_), .ZN(new_n19659_));
  AOI21_X1   g19593(.A1(new_n19658_), .A2(new_n19659_), .B(new_n2737_), .ZN(new_n19660_));
  NAND3_X1   g19594(.A1(new_n19553_), .A2(new_n74_), .A3(new_n19660_), .ZN(new_n19661_));
  INV_X1     g19595(.I(new_n19661_), .ZN(new_n19662_));
  AOI21_X1   g19596(.A1(new_n19553_), .A2(new_n19660_), .B(new_n74_), .ZN(new_n19663_));
  NOR2_X1    g19597(.A1(new_n19313_), .A2(new_n5021_), .ZN(new_n19664_));
  INV_X1     g19598(.I(new_n19664_), .ZN(new_n19665_));
  OAI21_X1   g19599(.A1(new_n19662_), .A2(new_n19663_), .B(new_n19665_), .ZN(new_n19666_));
  INV_X1     g19600(.I(new_n19663_), .ZN(new_n19667_));
  NAND3_X1   g19601(.A1(new_n19667_), .A2(new_n19661_), .A3(new_n19664_), .ZN(new_n19668_));
  AOI21_X1   g19602(.A1(new_n19666_), .A2(new_n19668_), .B(new_n19657_), .ZN(new_n19669_));
  NOR3_X1    g19603(.A1(new_n19634_), .A2(new_n19633_), .A3(new_n19631_), .ZN(new_n19670_));
  NAND3_X1   g19604(.A1(new_n19667_), .A2(new_n19661_), .A3(new_n19665_), .ZN(new_n19671_));
  OAI21_X1   g19605(.A1(new_n19662_), .A2(new_n19663_), .B(new_n19664_), .ZN(new_n19672_));
  AOI21_X1   g19606(.A1(new_n19671_), .A2(new_n19672_), .B(new_n19670_), .ZN(new_n19673_));
  NOR2_X1    g19607(.A1(new_n19673_), .A2(new_n19669_), .ZN(new_n19674_));
  NOR2_X1    g19608(.A1(new_n19317_), .A2(new_n19320_), .ZN(new_n19675_));
  AOI21_X1   g19609(.A1(new_n19613_), .A2(new_n19304_), .B(new_n19291_), .ZN(new_n19676_));
  NOR2_X1    g19610(.A1(new_n19676_), .A2(new_n19321_), .ZN(new_n19677_));
  XOR2_X1    g19611(.A1(new_n19304_), .A2(new_n19321_), .Z(new_n19678_));
  NOR4_X1    g19612(.A1(new_n19677_), .A2(new_n19675_), .A3(new_n17827_), .A4(new_n19678_), .ZN(new_n19679_));
  NAND2_X1   g19613(.A1(new_n19676_), .A2(new_n19321_), .ZN(new_n19680_));
  AOI21_X1   g19614(.A1(new_n19317_), .A2(new_n19320_), .B(new_n19678_), .ZN(new_n19681_));
  AOI21_X1   g19615(.A1(new_n19681_), .A2(new_n19680_), .B(new_n17828_), .ZN(new_n19682_));
  OAI22_X1   g19616(.A1(new_n19304_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n19320_), .ZN(new_n19683_));
  NAND2_X1   g19617(.A1(new_n17827_), .A2(new_n3317_), .ZN(new_n19684_));
  AOI21_X1   g19618(.A1(new_n19684_), .A2(new_n19683_), .B(new_n3260_), .ZN(new_n19685_));
  OAI21_X1   g19619(.A1(new_n19679_), .A2(new_n19682_), .B(new_n19685_), .ZN(new_n19686_));
  NOR2_X1    g19620(.A1(new_n19686_), .A2(\a[26] ), .ZN(new_n19687_));
  NAND2_X1   g19621(.A1(new_n19686_), .A2(\a[26] ), .ZN(new_n19688_));
  INV_X1     g19622(.I(new_n19688_), .ZN(new_n19689_));
  NOR3_X1    g19623(.A1(new_n19689_), .A2(new_n19674_), .A3(new_n19687_), .ZN(new_n19690_));
  OAI21_X1   g19624(.A1(new_n19689_), .A2(new_n19687_), .B(new_n19674_), .ZN(new_n19691_));
  OAI21_X1   g19625(.A1(new_n19656_), .A2(new_n19690_), .B(new_n19691_), .ZN(new_n19692_));
  AOI21_X1   g19626(.A1(new_n19667_), .A2(new_n19661_), .B(new_n19664_), .ZN(new_n19693_));
  AOI21_X1   g19627(.A1(new_n19657_), .A2(new_n19668_), .B(new_n19693_), .ZN(new_n19694_));
  AOI22_X1   g19628(.A1(new_n17850_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n19545_), .ZN(new_n19695_));
  AOI21_X1   g19629(.A1(new_n19305_), .A2(new_n2750_), .B(new_n19695_), .ZN(new_n19696_));
  NOR3_X1    g19630(.A1(new_n19618_), .A2(new_n2737_), .A3(new_n19696_), .ZN(new_n19697_));
  NAND2_X1   g19631(.A1(new_n19697_), .A2(new_n74_), .ZN(new_n19698_));
  NOR2_X1    g19632(.A1(new_n19696_), .A2(new_n2737_), .ZN(new_n19699_));
  NAND2_X1   g19633(.A1(new_n19607_), .A2(new_n19699_), .ZN(new_n19700_));
  NAND2_X1   g19634(.A1(new_n19700_), .A2(\a[29] ), .ZN(new_n19701_));
  OAI22_X1   g19635(.A1(new_n19313_), .A2(new_n2767_), .B1(new_n2772_), .B2(new_n19272_), .ZN(new_n19702_));
  NAND2_X1   g19636(.A1(new_n19577_), .A2(new_n2764_), .ZN(new_n19703_));
  NOR3_X1    g19637(.A1(new_n2135_), .A2(new_n2582_), .A3(new_n1730_), .ZN(new_n19704_));
  NOR4_X1    g19638(.A1(new_n495_), .A2(new_n548_), .A3(new_n867_), .A4(new_n468_), .ZN(new_n19705_));
  INV_X1     g19639(.I(new_n19705_), .ZN(new_n19706_));
  NOR3_X1    g19640(.A1(new_n268_), .A2(new_n1236_), .A3(new_n352_), .ZN(new_n19707_));
  NOR2_X1    g19641(.A1(new_n914_), .A2(new_n1664_), .ZN(new_n19708_));
  NAND4_X1   g19642(.A1(new_n19704_), .A2(new_n19708_), .A3(new_n19706_), .A4(new_n19707_), .ZN(new_n19709_));
  NAND4_X1   g19643(.A1(new_n1371_), .A2(new_n843_), .A3(new_n502_), .A4(new_n624_), .ZN(new_n19710_));
  NAND4_X1   g19644(.A1(new_n2153_), .A2(new_n511_), .A3(new_n1327_), .A4(new_n854_), .ZN(new_n19711_));
  INV_X1     g19645(.I(new_n2433_), .ZN(new_n19712_));
  NOR4_X1    g19646(.A1(new_n1257_), .A2(new_n2083_), .A3(new_n2381_), .A4(new_n1019_), .ZN(new_n19713_));
  NAND3_X1   g19647(.A1(new_n19713_), .A2(new_n19712_), .A3(new_n12916_), .ZN(new_n19714_));
  NOR4_X1    g19648(.A1(new_n19714_), .A2(new_n19709_), .A3(new_n19711_), .A4(new_n19710_), .ZN(new_n19715_));
  INV_X1     g19649(.I(new_n3362_), .ZN(new_n19716_));
  NAND4_X1   g19650(.A1(new_n2240_), .A2(new_n207_), .A3(new_n377_), .A4(new_n1891_), .ZN(new_n19717_));
  NAND4_X1   g19651(.A1(new_n19716_), .A2(new_n19717_), .A3(new_n775_), .A4(new_n1345_), .ZN(new_n19718_));
  NOR2_X1    g19652(.A1(new_n1994_), .A2(new_n1078_), .ZN(new_n19719_));
  NAND3_X1   g19653(.A1(new_n19719_), .A2(new_n11822_), .A3(new_n2862_), .ZN(new_n19720_));
  NAND4_X1   g19654(.A1(new_n162_), .A2(new_n947_), .A3(new_n1495_), .A4(new_n3159_), .ZN(new_n19721_));
  NOR4_X1    g19655(.A1(new_n19718_), .A2(new_n12510_), .A3(new_n19721_), .A4(new_n19720_), .ZN(new_n19722_));
  NAND3_X1   g19656(.A1(new_n19715_), .A2(new_n12985_), .A3(new_n19722_), .ZN(new_n19723_));
  INV_X1     g19657(.I(new_n19723_), .ZN(new_n19724_));
  AOI21_X1   g19658(.A1(new_n19703_), .A2(new_n19702_), .B(new_n19724_), .ZN(new_n19725_));
  NAND2_X1   g19659(.A1(new_n19703_), .A2(new_n19702_), .ZN(new_n19726_));
  NOR2_X1    g19660(.A1(new_n19726_), .A2(new_n19723_), .ZN(new_n19727_));
  NOR2_X1    g19661(.A1(new_n19727_), .A2(new_n19725_), .ZN(new_n19728_));
  NAND3_X1   g19662(.A1(new_n19698_), .A2(new_n19701_), .A3(new_n19728_), .ZN(new_n19729_));
  NOR2_X1    g19663(.A1(new_n19700_), .A2(\a[29] ), .ZN(new_n19730_));
  NOR2_X1    g19664(.A1(new_n19697_), .A2(new_n74_), .ZN(new_n19731_));
  XOR2_X1    g19665(.A1(new_n19726_), .A2(new_n19724_), .Z(new_n19732_));
  OAI21_X1   g19666(.A1(new_n19731_), .A2(new_n19730_), .B(new_n19732_), .ZN(new_n19733_));
  AOI21_X1   g19667(.A1(new_n19733_), .A2(new_n19729_), .B(new_n19694_), .ZN(new_n19734_));
  NOR3_X1    g19668(.A1(new_n19662_), .A2(new_n19663_), .A3(new_n19665_), .ZN(new_n19735_));
  OAI21_X1   g19669(.A1(new_n19670_), .A2(new_n19735_), .B(new_n19666_), .ZN(new_n19736_));
  OAI21_X1   g19670(.A1(new_n19731_), .A2(new_n19730_), .B(new_n19728_), .ZN(new_n19737_));
  NAND3_X1   g19671(.A1(new_n19698_), .A2(new_n19701_), .A3(new_n19732_), .ZN(new_n19738_));
  AOI21_X1   g19672(.A1(new_n19737_), .A2(new_n19738_), .B(new_n19736_), .ZN(new_n19739_));
  NOR2_X1    g19673(.A1(new_n19739_), .A2(new_n19734_), .ZN(new_n19740_));
  INV_X1     g19674(.I(new_n19322_), .ZN(new_n19741_));
  AOI22_X1   g19675(.A1(new_n19676_), .A2(new_n19741_), .B1(new_n19321_), .B2(new_n19323_), .ZN(new_n19742_));
  NAND2_X1   g19676(.A1(new_n19742_), .A2(new_n17827_), .ZN(new_n19743_));
  AOI21_X1   g19677(.A1(new_n19743_), .A2(new_n19326_), .B(new_n19343_), .ZN(new_n19744_));
  NAND2_X1   g19678(.A1(new_n19742_), .A2(new_n17828_), .ZN(new_n19745_));
  NAND2_X1   g19679(.A1(new_n19325_), .A2(new_n17827_), .ZN(new_n19746_));
  AOI21_X1   g19680(.A1(new_n19745_), .A2(new_n19746_), .B(new_n19349_), .ZN(new_n19747_));
  OAI22_X1   g19681(.A1(new_n17828_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19320_), .ZN(new_n19748_));
  NAND2_X1   g19682(.A1(new_n19349_), .A2(new_n3317_), .ZN(new_n19749_));
  AOI21_X1   g19683(.A1(new_n19749_), .A2(new_n19748_), .B(new_n3260_), .ZN(new_n19750_));
  OAI21_X1   g19684(.A1(new_n19744_), .A2(new_n19747_), .B(new_n19750_), .ZN(new_n19751_));
  NOR2_X1    g19685(.A1(new_n19751_), .A2(\a[26] ), .ZN(new_n19752_));
  NOR2_X1    g19686(.A1(new_n19742_), .A2(new_n17827_), .ZN(new_n19753_));
  NOR2_X1    g19687(.A1(new_n19325_), .A2(new_n17828_), .ZN(new_n19754_));
  OAI21_X1   g19688(.A1(new_n19753_), .A2(new_n19754_), .B(new_n19349_), .ZN(new_n19755_));
  NOR2_X1    g19689(.A1(new_n19325_), .A2(new_n17827_), .ZN(new_n19756_));
  NAND2_X1   g19690(.A1(new_n19676_), .A2(new_n19741_), .ZN(new_n19757_));
  AOI21_X1   g19691(.A1(new_n19757_), .A2(new_n19324_), .B(new_n17828_), .ZN(new_n19758_));
  OAI21_X1   g19692(.A1(new_n19758_), .A2(new_n19756_), .B(new_n19343_), .ZN(new_n19759_));
  NAND2_X1   g19693(.A1(new_n19755_), .A2(new_n19759_), .ZN(new_n19760_));
  AOI21_X1   g19694(.A1(new_n19760_), .A2(new_n19750_), .B(new_n72_), .ZN(new_n19761_));
  NOR2_X1    g19695(.A1(new_n19752_), .A2(new_n19761_), .ZN(new_n19762_));
  NAND2_X1   g19696(.A1(new_n19762_), .A2(new_n19740_), .ZN(new_n19763_));
  NAND2_X1   g19697(.A1(new_n19692_), .A2(new_n19763_), .ZN(new_n19764_));
  NOR2_X1    g19698(.A1(new_n19762_), .A2(new_n19740_), .ZN(new_n19765_));
  INV_X1     g19699(.I(new_n19765_), .ZN(new_n19766_));
  NAND2_X1   g19700(.A1(new_n19764_), .A2(new_n19766_), .ZN(new_n19767_));
  NOR3_X1    g19701(.A1(new_n19731_), .A2(new_n19730_), .A3(new_n19732_), .ZN(new_n19768_));
  OAI21_X1   g19702(.A1(new_n19694_), .A2(new_n19768_), .B(new_n19733_), .ZN(new_n19769_));
  OAI22_X1   g19703(.A1(new_n19304_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n17849_), .ZN(new_n19770_));
  NAND2_X1   g19704(.A1(new_n19321_), .A2(new_n2750_), .ZN(new_n19771_));
  AOI21_X1   g19705(.A1(new_n19770_), .A2(new_n19771_), .B(new_n2737_), .ZN(new_n19772_));
  NAND3_X1   g19706(.A1(new_n19647_), .A2(new_n74_), .A3(new_n19772_), .ZN(new_n19773_));
  AOI21_X1   g19707(.A1(new_n19647_), .A2(new_n19772_), .B(new_n74_), .ZN(new_n19774_));
  INV_X1     g19708(.I(new_n19774_), .ZN(new_n19775_));
  OAI22_X1   g19709(.A1(new_n19313_), .A2(new_n2771_), .B1(new_n2767_), .B2(new_n19272_), .ZN(new_n19776_));
  OAI21_X1   g19710(.A1(new_n2772_), .A2(new_n19275_), .B(new_n19776_), .ZN(new_n19777_));
  NAND3_X1   g19711(.A1(new_n19564_), .A2(new_n19777_), .A3(new_n2764_), .ZN(new_n19778_));
  NAND4_X1   g19712(.A1(new_n2430_), .A2(new_n1044_), .A3(new_n1214_), .A4(new_n11507_), .ZN(new_n19779_));
  NAND2_X1   g19713(.A1(new_n8315_), .A2(new_n2849_), .ZN(new_n19780_));
  NOR2_X1    g19714(.A1(new_n19780_), .A2(new_n19779_), .ZN(new_n19781_));
  INV_X1     g19715(.I(new_n3929_), .ZN(new_n19782_));
  NAND3_X1   g19716(.A1(new_n1021_), .A2(new_n435_), .A3(new_n1059_), .ZN(new_n19783_));
  INV_X1     g19717(.I(new_n19783_), .ZN(new_n19784_));
  NOR2_X1    g19718(.A1(new_n11478_), .A2(new_n891_), .ZN(new_n19785_));
  NAND2_X1   g19719(.A1(new_n19784_), .A2(new_n19785_), .ZN(new_n19786_));
  NOR4_X1    g19720(.A1(new_n906_), .A2(new_n610_), .A3(new_n1236_), .A4(new_n1035_), .ZN(new_n19787_));
  NOR3_X1    g19721(.A1(new_n81_), .A2(new_n603_), .A3(new_n453_), .ZN(new_n19788_));
  INV_X1     g19722(.I(new_n19788_), .ZN(new_n19789_));
  NOR4_X1    g19723(.A1(new_n19786_), .A2(new_n19782_), .A3(new_n19787_), .A4(new_n19789_), .ZN(new_n19790_));
  NAND4_X1   g19724(.A1(new_n19781_), .A2(new_n19790_), .A3(new_n12985_), .A4(new_n4801_), .ZN(new_n19791_));
  INV_X1     g19725(.I(new_n19791_), .ZN(new_n19792_));
  NOR2_X1    g19726(.A1(new_n19778_), .A2(new_n19792_), .ZN(new_n19793_));
  NOR2_X1    g19727(.A1(new_n19571_), .A2(new_n2763_), .ZN(new_n19794_));
  AOI21_X1   g19728(.A1(new_n19794_), .A2(new_n19777_), .B(new_n19791_), .ZN(new_n19795_));
  OAI21_X1   g19729(.A1(new_n19793_), .A2(new_n19795_), .B(new_n19725_), .ZN(new_n19796_));
  INV_X1     g19730(.I(new_n19725_), .ZN(new_n19797_));
  AOI21_X1   g19731(.A1(new_n19794_), .A2(new_n19777_), .B(new_n19792_), .ZN(new_n19798_));
  NOR2_X1    g19732(.A1(new_n19778_), .A2(new_n19791_), .ZN(new_n19799_));
  OAI21_X1   g19733(.A1(new_n19799_), .A2(new_n19798_), .B(new_n19797_), .ZN(new_n19800_));
  NAND2_X1   g19734(.A1(new_n19800_), .A2(new_n19796_), .ZN(new_n19801_));
  AOI21_X1   g19735(.A1(new_n19773_), .A2(new_n19775_), .B(new_n19801_), .ZN(new_n19802_));
  INV_X1     g19736(.I(new_n19773_), .ZN(new_n19803_));
  NAND3_X1   g19737(.A1(new_n19794_), .A2(new_n19777_), .A3(new_n19791_), .ZN(new_n19804_));
  NAND2_X1   g19738(.A1(new_n19778_), .A2(new_n19792_), .ZN(new_n19805_));
  AOI21_X1   g19739(.A1(new_n19804_), .A2(new_n19805_), .B(new_n19797_), .ZN(new_n19806_));
  NAND2_X1   g19740(.A1(new_n19778_), .A2(new_n19791_), .ZN(new_n19807_));
  NAND3_X1   g19741(.A1(new_n19794_), .A2(new_n19777_), .A3(new_n19792_), .ZN(new_n19808_));
  AOI21_X1   g19742(.A1(new_n19807_), .A2(new_n19808_), .B(new_n19725_), .ZN(new_n19809_));
  NOR2_X1    g19743(.A1(new_n19806_), .A2(new_n19809_), .ZN(new_n19810_));
  NOR3_X1    g19744(.A1(new_n19810_), .A2(new_n19803_), .A3(new_n19774_), .ZN(new_n19811_));
  OAI21_X1   g19745(.A1(new_n19802_), .A2(new_n19811_), .B(new_n19769_), .ZN(new_n19812_));
  AOI21_X1   g19746(.A1(new_n19698_), .A2(new_n19701_), .B(new_n19728_), .ZN(new_n19813_));
  AOI21_X1   g19747(.A1(new_n19736_), .A2(new_n19729_), .B(new_n19813_), .ZN(new_n19814_));
  NOR3_X1    g19748(.A1(new_n19801_), .A2(new_n19803_), .A3(new_n19774_), .ZN(new_n19815_));
  AOI21_X1   g19749(.A1(new_n19773_), .A2(new_n19775_), .B(new_n19810_), .ZN(new_n19816_));
  OAI21_X1   g19750(.A1(new_n19815_), .A2(new_n19816_), .B(new_n19814_), .ZN(new_n19817_));
  AND2_X2    g19751(.A1(new_n19812_), .A2(new_n19817_), .Z(new_n19818_));
  OAI21_X1   g19752(.A1(new_n19325_), .A2(new_n17828_), .B(new_n19343_), .ZN(new_n19819_));
  AOI21_X1   g19753(.A1(new_n19325_), .A2(new_n17828_), .B(new_n19343_), .ZN(new_n19820_));
  INV_X1     g19754(.I(new_n19820_), .ZN(new_n19821_));
  AOI21_X1   g19755(.A1(new_n19821_), .A2(new_n19819_), .B(new_n19346_), .ZN(new_n19822_));
  NAND3_X1   g19756(.A1(new_n19742_), .A2(new_n17827_), .A3(new_n19343_), .ZN(new_n19823_));
  NAND3_X1   g19757(.A1(new_n19325_), .A2(new_n17828_), .A3(new_n19349_), .ZN(new_n19824_));
  AOI21_X1   g19758(.A1(new_n19823_), .A2(new_n19824_), .B(new_n19350_), .ZN(new_n19825_));
  OAI22_X1   g19759(.A1(new_n3322_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n3268_), .ZN(new_n19826_));
  NAND2_X1   g19760(.A1(new_n19350_), .A2(new_n3317_), .ZN(new_n19827_));
  AOI21_X1   g19761(.A1(new_n19826_), .A2(new_n19827_), .B(new_n3260_), .ZN(new_n19828_));
  OAI21_X1   g19762(.A1(new_n19822_), .A2(new_n19825_), .B(new_n19828_), .ZN(new_n19829_));
  XOR2_X1    g19763(.A1(new_n19829_), .A2(\a[26] ), .Z(new_n19830_));
  INV_X1     g19764(.I(new_n19830_), .ZN(new_n19831_));
  NOR2_X1    g19765(.A1(new_n19818_), .A2(new_n19831_), .ZN(new_n19832_));
  NAND2_X1   g19766(.A1(new_n19812_), .A2(new_n19817_), .ZN(new_n19833_));
  NOR2_X1    g19767(.A1(new_n19833_), .A2(new_n19830_), .ZN(new_n19834_));
  OAI21_X1   g19768(.A1(new_n19832_), .A2(new_n19834_), .B(new_n19767_), .ZN(new_n19835_));
  INV_X1     g19769(.I(new_n19557_), .ZN(new_n19836_));
  OAI21_X1   g19770(.A1(new_n19836_), .A2(new_n19558_), .B(new_n19630_), .ZN(new_n19837_));
  NOR2_X1    g19771(.A1(new_n19573_), .A2(\a[26] ), .ZN(new_n19838_));
  NOR2_X1    g19772(.A1(new_n19568_), .A2(new_n72_), .ZN(new_n19839_));
  NAND2_X1   g19773(.A1(new_n19578_), .A2(new_n19580_), .ZN(new_n19840_));
  NOR2_X1    g19774(.A1(new_n19593_), .A2(new_n19840_), .ZN(new_n19841_));
  INV_X1     g19775(.I(new_n19582_), .ZN(new_n19842_));
  NAND3_X1   g19776(.A1(new_n19841_), .A2(\a[26] ), .A3(new_n19842_), .ZN(new_n19843_));
  NOR3_X1    g19777(.A1(new_n19838_), .A2(new_n19839_), .A3(new_n19843_), .ZN(new_n19844_));
  NOR3_X1    g19778(.A1(new_n19836_), .A2(new_n19630_), .A3(new_n19558_), .ZN(new_n19845_));
  OAI21_X1   g19779(.A1(new_n19844_), .A2(new_n19845_), .B(new_n19837_), .ZN(new_n19846_));
  NAND2_X1   g19780(.A1(new_n19595_), .A2(new_n74_), .ZN(new_n19847_));
  NAND2_X1   g19781(.A1(new_n19589_), .A2(\a[29] ), .ZN(new_n19848_));
  INV_X1     g19782(.I(new_n19597_), .ZN(new_n19849_));
  NAND3_X1   g19783(.A1(new_n19848_), .A2(new_n19847_), .A3(new_n19849_), .ZN(new_n19850_));
  INV_X1     g19784(.I(new_n19599_), .ZN(new_n19851_));
  NAND2_X1   g19785(.A1(new_n19850_), .A2(new_n19851_), .ZN(new_n19852_));
  NAND2_X1   g19786(.A1(new_n19619_), .A2(new_n72_), .ZN(new_n19853_));
  NAND2_X1   g19787(.A1(new_n19611_), .A2(\a[26] ), .ZN(new_n19854_));
  NAND3_X1   g19788(.A1(new_n19853_), .A2(new_n19854_), .A3(new_n19852_), .ZN(new_n19855_));
  AOI21_X1   g19789(.A1(new_n19853_), .A2(new_n19854_), .B(new_n19852_), .ZN(new_n19856_));
  AOI21_X1   g19790(.A1(new_n19846_), .A2(new_n19855_), .B(new_n19856_), .ZN(new_n19857_));
  NOR3_X1    g19791(.A1(new_n19634_), .A2(new_n19633_), .A3(new_n19635_), .ZN(new_n19858_));
  AOI21_X1   g19792(.A1(new_n19627_), .A2(new_n19629_), .B(new_n19631_), .ZN(new_n19859_));
  NOR2_X1    g19793(.A1(new_n19858_), .A2(new_n19859_), .ZN(new_n19860_));
  INV_X1     g19794(.I(new_n19651_), .ZN(new_n19861_));
  NOR3_X1    g19795(.A1(new_n19860_), .A2(new_n19861_), .A3(new_n19652_), .ZN(new_n19862_));
  OAI21_X1   g19796(.A1(new_n19861_), .A2(new_n19652_), .B(new_n19860_), .ZN(new_n19863_));
  OAI21_X1   g19797(.A1(new_n19857_), .A2(new_n19862_), .B(new_n19863_), .ZN(new_n19864_));
  OAI21_X1   g19798(.A1(new_n19693_), .A2(new_n19735_), .B(new_n19670_), .ZN(new_n19865_));
  NOR3_X1    g19799(.A1(new_n19662_), .A2(new_n19663_), .A3(new_n19664_), .ZN(new_n19866_));
  AOI21_X1   g19800(.A1(new_n19667_), .A2(new_n19661_), .B(new_n19665_), .ZN(new_n19867_));
  OAI21_X1   g19801(.A1(new_n19866_), .A2(new_n19867_), .B(new_n19657_), .ZN(new_n19868_));
  NAND2_X1   g19802(.A1(new_n19865_), .A2(new_n19868_), .ZN(new_n19869_));
  INV_X1     g19803(.I(new_n19687_), .ZN(new_n19870_));
  NAND3_X1   g19804(.A1(new_n19870_), .A2(new_n19869_), .A3(new_n19688_), .ZN(new_n19871_));
  AOI21_X1   g19805(.A1(new_n19870_), .A2(new_n19688_), .B(new_n19869_), .ZN(new_n19872_));
  AOI21_X1   g19806(.A1(new_n19864_), .A2(new_n19871_), .B(new_n19872_), .ZN(new_n19873_));
  NAND3_X1   g19807(.A1(new_n19760_), .A2(new_n72_), .A3(new_n19750_), .ZN(new_n19874_));
  NAND2_X1   g19808(.A1(new_n19751_), .A2(\a[26] ), .ZN(new_n19875_));
  NAND2_X1   g19809(.A1(new_n19875_), .A2(new_n19874_), .ZN(new_n19876_));
  NOR3_X1    g19810(.A1(new_n19876_), .A2(new_n19734_), .A3(new_n19739_), .ZN(new_n19877_));
  NOR2_X1    g19811(.A1(new_n19873_), .A2(new_n19877_), .ZN(new_n19878_));
  NOR2_X1    g19812(.A1(new_n19878_), .A2(new_n19765_), .ZN(new_n19879_));
  XOR2_X1    g19813(.A1(new_n19833_), .A2(new_n19830_), .Z(new_n19880_));
  NAND2_X1   g19814(.A1(new_n19880_), .A2(new_n19879_), .ZN(new_n19881_));
  NAND3_X1   g19815(.A1(new_n19543_), .A2(new_n19881_), .A3(new_n19835_), .ZN(new_n19882_));
  XOR2_X1    g19816(.A1(new_n19542_), .A2(\a[23] ), .Z(new_n19883_));
  NAND2_X1   g19817(.A1(new_n19881_), .A2(new_n19835_), .ZN(new_n19884_));
  NAND2_X1   g19818(.A1(new_n19884_), .A2(new_n19883_), .ZN(new_n19885_));
  OAI21_X1   g19819(.A1(new_n19877_), .A2(new_n19765_), .B(new_n19692_), .ZN(new_n19886_));
  NOR2_X1    g19820(.A1(new_n19740_), .A2(new_n19876_), .ZN(new_n19887_));
  NAND2_X1   g19821(.A1(new_n19740_), .A2(new_n19876_), .ZN(new_n19888_));
  INV_X1     g19822(.I(new_n19888_), .ZN(new_n19889_));
  OAI21_X1   g19823(.A1(new_n19889_), .A2(new_n19887_), .B(new_n19873_), .ZN(new_n19890_));
  INV_X1     g19824(.I(new_n19352_), .ZN(new_n19891_));
  AOI21_X1   g19825(.A1(new_n19891_), .A2(new_n19357_), .B(new_n19356_), .ZN(new_n19892_));
  NAND3_X1   g19826(.A1(new_n19348_), .A2(new_n17806_), .A3(new_n19351_), .ZN(new_n19893_));
  NAND2_X1   g19827(.A1(new_n19528_), .A2(new_n17807_), .ZN(new_n19894_));
  AOI21_X1   g19828(.A1(new_n19894_), .A2(new_n19893_), .B(new_n19359_), .ZN(new_n19895_));
  OAI22_X1   g19829(.A1(new_n17806_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19346_), .ZN(new_n19896_));
  NAND2_X1   g19830(.A1(new_n19359_), .A2(new_n3312_), .ZN(new_n19897_));
  AOI21_X1   g19831(.A1(new_n19897_), .A2(new_n19896_), .B(new_n3302_), .ZN(new_n19898_));
  OAI21_X1   g19832(.A1(new_n19892_), .A2(new_n19895_), .B(new_n19898_), .ZN(new_n19899_));
  NOR2_X1    g19833(.A1(new_n19899_), .A2(\a[23] ), .ZN(new_n19900_));
  INV_X1     g19834(.I(new_n19900_), .ZN(new_n19901_));
  NAND2_X1   g19835(.A1(new_n19899_), .A2(\a[23] ), .ZN(new_n19902_));
  NAND4_X1   g19836(.A1(new_n19890_), .A2(new_n19886_), .A3(new_n19901_), .A4(new_n19902_), .ZN(new_n19903_));
  INV_X1     g19837(.I(new_n19819_), .ZN(new_n19904_));
  NOR2_X1    g19838(.A1(new_n19904_), .A2(new_n19820_), .ZN(new_n19905_));
  AOI21_X1   g19839(.A1(new_n19344_), .A2(new_n19326_), .B(new_n19350_), .ZN(new_n19906_));
  NAND3_X1   g19840(.A1(new_n19344_), .A2(new_n19326_), .A3(new_n19350_), .ZN(new_n19907_));
  INV_X1     g19841(.I(new_n19907_), .ZN(new_n19908_));
  NOR3_X1    g19842(.A1(new_n19908_), .A2(new_n19905_), .A3(new_n19906_), .ZN(new_n19909_));
  NAND2_X1   g19843(.A1(new_n19909_), .A2(new_n17806_), .ZN(new_n19910_));
  NAND2_X1   g19844(.A1(new_n19821_), .A2(new_n19819_), .ZN(new_n19911_));
  INV_X1     g19845(.I(new_n19906_), .ZN(new_n19912_));
  NAND3_X1   g19846(.A1(new_n19912_), .A2(new_n19911_), .A3(new_n19907_), .ZN(new_n19913_));
  NAND2_X1   g19847(.A1(new_n19913_), .A2(new_n17807_), .ZN(new_n19914_));
  NAND2_X1   g19848(.A1(new_n19910_), .A2(new_n19914_), .ZN(new_n19915_));
  AOI22_X1   g19849(.A1(new_n19349_), .A2(new_n5291_), .B1(new_n3782_), .B2(new_n19350_), .ZN(new_n19916_));
  NOR2_X1    g19850(.A1(new_n17806_), .A2(new_n3780_), .ZN(new_n19917_));
  OAI21_X1   g19851(.A1(new_n19916_), .A2(new_n19917_), .B(new_n3301_), .ZN(new_n19918_));
  NOR3_X1    g19852(.A1(new_n19915_), .A2(\a[23] ), .A3(new_n19918_), .ZN(new_n19919_));
  NOR2_X1    g19853(.A1(new_n19913_), .A2(new_n17807_), .ZN(new_n19920_));
  NOR2_X1    g19854(.A1(new_n19909_), .A2(new_n17806_), .ZN(new_n19921_));
  NOR2_X1    g19855(.A1(new_n19921_), .A2(new_n19920_), .ZN(new_n19922_));
  INV_X1     g19856(.I(new_n19918_), .ZN(new_n19923_));
  AOI21_X1   g19857(.A1(new_n19922_), .A2(new_n19923_), .B(new_n84_), .ZN(new_n19924_));
  NOR2_X1    g19858(.A1(new_n19924_), .A2(new_n19919_), .ZN(new_n19925_));
  NAND3_X1   g19859(.A1(new_n19870_), .A2(new_n19674_), .A3(new_n19688_), .ZN(new_n19926_));
  OAI21_X1   g19860(.A1(new_n19689_), .A2(new_n19687_), .B(new_n19869_), .ZN(new_n19927_));
  NAND2_X1   g19861(.A1(new_n19927_), .A2(new_n19926_), .ZN(new_n19928_));
  NAND2_X1   g19862(.A1(new_n19928_), .A2(new_n19864_), .ZN(new_n19929_));
  OAI21_X1   g19863(.A1(new_n19690_), .A2(new_n19872_), .B(new_n19656_), .ZN(new_n19930_));
  NAND2_X1   g19864(.A1(new_n19929_), .A2(new_n19930_), .ZN(new_n19931_));
  NAND2_X1   g19865(.A1(new_n19925_), .A2(new_n19931_), .ZN(new_n19932_));
  AOI21_X1   g19866(.A1(new_n19766_), .A2(new_n19763_), .B(new_n19873_), .ZN(new_n19933_));
  INV_X1     g19867(.I(new_n19740_), .ZN(new_n19934_));
  NAND2_X1   g19868(.A1(new_n19934_), .A2(new_n19762_), .ZN(new_n19935_));
  AOI21_X1   g19869(.A1(new_n19935_), .A2(new_n19888_), .B(new_n19692_), .ZN(new_n19936_));
  INV_X1     g19870(.I(new_n19902_), .ZN(new_n19937_));
  OAI22_X1   g19871(.A1(new_n19933_), .A2(new_n19936_), .B1(new_n19937_), .B2(new_n19900_), .ZN(new_n19938_));
  NAND3_X1   g19872(.A1(new_n19938_), .A2(new_n19903_), .A3(new_n19932_), .ZN(new_n19939_));
  AOI22_X1   g19873(.A1(new_n19885_), .A2(new_n19882_), .B1(new_n19543_), .B2(new_n19939_), .ZN(new_n19940_));
  NAND2_X1   g19874(.A1(new_n19358_), .A2(new_n19365_), .ZN(new_n19941_));
  NAND2_X1   g19875(.A1(new_n19357_), .A2(new_n19356_), .ZN(new_n19942_));
  NAND2_X1   g19876(.A1(new_n19942_), .A2(new_n19891_), .ZN(new_n19943_));
  NAND2_X1   g19877(.A1(new_n19943_), .A2(new_n19364_), .ZN(new_n19944_));
  XOR2_X1    g19878(.A1(new_n19356_), .A2(new_n19365_), .Z(new_n19945_));
  INV_X1     g19879(.I(new_n19945_), .ZN(new_n19946_));
  NAND4_X1   g19880(.A1(new_n19944_), .A2(new_n17801_), .A3(new_n19941_), .A4(new_n19946_), .ZN(new_n19947_));
  NOR2_X1    g19881(.A1(new_n19943_), .A2(new_n19364_), .ZN(new_n19948_));
  OAI21_X1   g19882(.A1(new_n19358_), .A2(new_n19365_), .B(new_n19946_), .ZN(new_n19949_));
  OAI21_X1   g19883(.A1(new_n19948_), .A2(new_n19949_), .B(new_n17802_), .ZN(new_n19950_));
  NAND2_X1   g19884(.A1(new_n19947_), .A2(new_n19950_), .ZN(new_n19951_));
  OAI22_X1   g19885(.A1(new_n19356_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n19364_), .ZN(new_n19952_));
  NAND2_X1   g19886(.A1(new_n17802_), .A2(new_n3312_), .ZN(new_n19953_));
  AOI21_X1   g19887(.A1(new_n19952_), .A2(new_n19953_), .B(new_n3302_), .ZN(new_n19954_));
  NAND2_X1   g19888(.A1(new_n19951_), .A2(new_n19954_), .ZN(new_n19955_));
  XOR2_X1    g19889(.A1(new_n19955_), .A2(\a[23] ), .Z(new_n19956_));
  OAI21_X1   g19890(.A1(new_n19803_), .A2(new_n19774_), .B(new_n19801_), .ZN(new_n19957_));
  OAI21_X1   g19891(.A1(new_n19814_), .A2(new_n19815_), .B(new_n19957_), .ZN(new_n19958_));
  OAI22_X1   g19892(.A1(new_n19304_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n19320_), .ZN(new_n19959_));
  NAND2_X1   g19893(.A1(new_n17827_), .A2(new_n2750_), .ZN(new_n19960_));
  AOI21_X1   g19894(.A1(new_n19960_), .A2(new_n19959_), .B(new_n2737_), .ZN(new_n19961_));
  OAI21_X1   g19895(.A1(new_n19679_), .A2(new_n19682_), .B(new_n19961_), .ZN(new_n19962_));
  NOR2_X1    g19896(.A1(new_n19962_), .A2(\a[29] ), .ZN(new_n19963_));
  INV_X1     g19897(.I(new_n19963_), .ZN(new_n19964_));
  NAND2_X1   g19898(.A1(new_n19962_), .A2(\a[29] ), .ZN(new_n19965_));
  AOI21_X1   g19899(.A1(new_n19797_), .A2(new_n19807_), .B(new_n19799_), .ZN(new_n19966_));
  AOI21_X1   g19900(.A1(new_n19545_), .A2(new_n3189_), .B(new_n2763_), .ZN(new_n19967_));
  OAI21_X1   g19901(.A1(new_n17849_), .A2(new_n2772_), .B(new_n19967_), .ZN(new_n19968_));
  AOI21_X1   g19902(.A1(new_n19308_), .A2(new_n2770_), .B(new_n19968_), .ZN(new_n19969_));
  NAND2_X1   g19903(.A1(new_n19553_), .A2(new_n19969_), .ZN(new_n19970_));
  NOR4_X1    g19904(.A1(new_n576_), .A2(new_n879_), .A3(new_n687_), .A4(new_n1620_), .ZN(new_n19971_));
  NAND4_X1   g19905(.A1(new_n469_), .A2(new_n110_), .A3(new_n182_), .A4(new_n1468_), .ZN(new_n19972_));
  NOR3_X1    g19906(.A1(new_n563_), .A2(new_n320_), .A3(new_n584_), .ZN(new_n19973_));
  AND3_X2    g19907(.A1(new_n19971_), .A2(new_n19972_), .A3(new_n19973_), .Z(new_n19974_));
  NOR4_X1    g19908(.A1(new_n2330_), .A2(new_n4752_), .A3(new_n3412_), .A4(new_n3856_), .ZN(new_n19975_));
  NAND4_X1   g19909(.A1(new_n19974_), .A2(new_n3979_), .A3(new_n4002_), .A4(new_n19975_), .ZN(new_n19976_));
  OR3_X2     g19910(.A1(new_n1455_), .A2(new_n2469_), .A3(new_n19976_), .Z(new_n19977_));
  NAND2_X1   g19911(.A1(new_n19970_), .A2(new_n19977_), .ZN(new_n19978_));
  INV_X1     g19912(.I(new_n19978_), .ZN(new_n19979_));
  NOR2_X1    g19913(.A1(new_n19970_), .A2(new_n19977_), .ZN(new_n19980_));
  NOR2_X1    g19914(.A1(new_n19979_), .A2(new_n19980_), .ZN(new_n19981_));
  XOR2_X1    g19915(.A1(new_n19970_), .A2(new_n19977_), .Z(new_n19982_));
  NAND2_X1   g19916(.A1(new_n19982_), .A2(new_n19966_), .ZN(new_n19983_));
  OAI21_X1   g19917(.A1(new_n19966_), .A2(new_n19981_), .B(new_n19983_), .ZN(new_n19984_));
  AOI21_X1   g19918(.A1(new_n19964_), .A2(new_n19965_), .B(new_n19984_), .ZN(new_n19985_));
  INV_X1     g19919(.I(new_n19965_), .ZN(new_n19986_));
  NAND2_X1   g19920(.A1(new_n19797_), .A2(new_n19807_), .ZN(new_n19987_));
  INV_X1     g19921(.I(new_n19980_), .ZN(new_n19988_));
  AOI22_X1   g19922(.A1(new_n19987_), .A2(new_n19808_), .B1(new_n19988_), .B2(new_n19978_), .ZN(new_n19989_));
  AOI21_X1   g19923(.A1(new_n19966_), .A2(new_n19982_), .B(new_n19989_), .ZN(new_n19990_));
  NOR3_X1    g19924(.A1(new_n19990_), .A2(new_n19986_), .A3(new_n19963_), .ZN(new_n19991_));
  OAI21_X1   g19925(.A1(new_n19985_), .A2(new_n19991_), .B(new_n19958_), .ZN(new_n19992_));
  NAND3_X1   g19926(.A1(new_n19810_), .A2(new_n19775_), .A3(new_n19773_), .ZN(new_n19993_));
  AOI21_X1   g19927(.A1(new_n19769_), .A2(new_n19993_), .B(new_n19816_), .ZN(new_n19994_));
  NOR3_X1    g19928(.A1(new_n19984_), .A2(new_n19986_), .A3(new_n19963_), .ZN(new_n19995_));
  AOI21_X1   g19929(.A1(new_n19964_), .A2(new_n19965_), .B(new_n19990_), .ZN(new_n19996_));
  OAI21_X1   g19930(.A1(new_n19995_), .A2(new_n19996_), .B(new_n19994_), .ZN(new_n19997_));
  NAND2_X1   g19931(.A1(new_n19997_), .A2(new_n19992_), .ZN(new_n19998_));
  AOI22_X1   g19932(.A1(new_n19349_), .A2(new_n3267_), .B1(new_n3323_), .B2(new_n19350_), .ZN(new_n19999_));
  NOR2_X1    g19933(.A1(new_n17806_), .A2(new_n3318_), .ZN(new_n20000_));
  OAI21_X1   g19934(.A1(new_n19999_), .A2(new_n20000_), .B(new_n3259_), .ZN(new_n20001_));
  NOR3_X1    g19935(.A1(new_n19915_), .A2(\a[26] ), .A3(new_n20001_), .ZN(new_n20002_));
  INV_X1     g19936(.I(new_n20001_), .ZN(new_n20003_));
  AOI21_X1   g19937(.A1(new_n19922_), .A2(new_n20003_), .B(new_n72_), .ZN(new_n20004_));
  NOR2_X1    g19938(.A1(new_n20004_), .A2(new_n20002_), .ZN(new_n20005_));
  NOR2_X1    g19939(.A1(new_n20005_), .A2(new_n19998_), .ZN(new_n20006_));
  NOR2_X1    g19940(.A1(new_n19768_), .A2(new_n19694_), .ZN(new_n20007_));
  OAI21_X1   g19941(.A1(new_n20007_), .A2(new_n19813_), .B(new_n19993_), .ZN(new_n20008_));
  OAI21_X1   g19942(.A1(new_n19963_), .A2(new_n19986_), .B(new_n19990_), .ZN(new_n20009_));
  NAND3_X1   g19943(.A1(new_n19984_), .A2(new_n19964_), .A3(new_n19965_), .ZN(new_n20010_));
  AOI22_X1   g19944(.A1(new_n20009_), .A2(new_n20010_), .B1(new_n20008_), .B2(new_n19957_), .ZN(new_n20011_));
  NAND3_X1   g19945(.A1(new_n19990_), .A2(new_n19964_), .A3(new_n19965_), .ZN(new_n20012_));
  OAI21_X1   g19946(.A1(new_n19986_), .A2(new_n19963_), .B(new_n19984_), .ZN(new_n20013_));
  AOI21_X1   g19947(.A1(new_n20012_), .A2(new_n20013_), .B(new_n19958_), .ZN(new_n20014_));
  NOR2_X1    g19948(.A1(new_n20014_), .A2(new_n20011_), .ZN(new_n20015_));
  NOR3_X1    g19949(.A1(new_n20015_), .A2(new_n20002_), .A3(new_n20004_), .ZN(new_n20016_));
  NOR2_X1    g19950(.A1(new_n20006_), .A2(new_n20016_), .ZN(new_n20017_));
  NAND3_X1   g19951(.A1(new_n19764_), .A2(new_n19766_), .A3(new_n19831_), .ZN(new_n20018_));
  OAI21_X1   g19952(.A1(new_n19878_), .A2(new_n19765_), .B(new_n19830_), .ZN(new_n20019_));
  AOI21_X1   g19953(.A1(new_n20019_), .A2(new_n20018_), .B(new_n19833_), .ZN(new_n20020_));
  NAND2_X1   g19954(.A1(new_n20017_), .A2(new_n20020_), .ZN(new_n20021_));
  OAI21_X1   g19955(.A1(new_n20002_), .A2(new_n20004_), .B(new_n20015_), .ZN(new_n20022_));
  NAND2_X1   g19956(.A1(new_n20005_), .A2(new_n19998_), .ZN(new_n20023_));
  NAND2_X1   g19957(.A1(new_n20022_), .A2(new_n20023_), .ZN(new_n20024_));
  NOR3_X1    g19958(.A1(new_n19878_), .A2(new_n19765_), .A3(new_n19830_), .ZN(new_n20025_));
  AOI21_X1   g19959(.A1(new_n19764_), .A2(new_n19766_), .B(new_n19831_), .ZN(new_n20026_));
  OAI21_X1   g19960(.A1(new_n20025_), .A2(new_n20026_), .B(new_n19818_), .ZN(new_n20027_));
  NAND2_X1   g19961(.A1(new_n20024_), .A2(new_n20027_), .ZN(new_n20028_));
  NOR2_X1    g19962(.A1(new_n19879_), .A2(new_n19830_), .ZN(new_n20029_));
  NAND3_X1   g19963(.A1(new_n20028_), .A2(new_n20021_), .A3(new_n20029_), .ZN(new_n20030_));
  NOR2_X1    g19964(.A1(new_n20024_), .A2(new_n20027_), .ZN(new_n20031_));
  NOR2_X1    g19965(.A1(new_n20017_), .A2(new_n20020_), .ZN(new_n20032_));
  INV_X1     g19966(.I(new_n20029_), .ZN(new_n20033_));
  OAI21_X1   g19967(.A1(new_n20031_), .A2(new_n20032_), .B(new_n20033_), .ZN(new_n20034_));
  NAND3_X1   g19968(.A1(new_n20034_), .A2(new_n20030_), .A3(new_n19956_), .ZN(new_n20035_));
  NAND2_X1   g19969(.A1(new_n20035_), .A2(new_n19940_), .ZN(new_n20036_));
  INV_X1     g19970(.I(new_n19956_), .ZN(new_n20037_));
  NOR3_X1    g19971(.A1(new_n20031_), .A2(new_n20032_), .A3(new_n20033_), .ZN(new_n20038_));
  AOI21_X1   g19972(.A1(new_n20028_), .A2(new_n20021_), .B(new_n20029_), .ZN(new_n20039_));
  OAI21_X1   g19973(.A1(new_n20039_), .A2(new_n20038_), .B(new_n20037_), .ZN(new_n20040_));
  NAND2_X1   g19974(.A1(new_n20036_), .A2(new_n20040_), .ZN(new_n20041_));
  NAND2_X1   g19975(.A1(new_n19369_), .A2(new_n17801_), .ZN(new_n20042_));
  NOR2_X1    g19976(.A1(new_n19369_), .A2(new_n17801_), .ZN(new_n20043_));
  INV_X1     g19977(.I(new_n20043_), .ZN(new_n20044_));
  AOI21_X1   g19978(.A1(new_n20044_), .A2(new_n20042_), .B(new_n17797_), .ZN(new_n20045_));
  INV_X1     g19979(.I(new_n19368_), .ZN(new_n20046_));
  OAI21_X1   g19980(.A1(new_n19943_), .A2(new_n19366_), .B(new_n20046_), .ZN(new_n20047_));
  NAND2_X1   g19981(.A1(new_n20047_), .A2(new_n17801_), .ZN(new_n20048_));
  NAND2_X1   g19982(.A1(new_n19369_), .A2(new_n17802_), .ZN(new_n20049_));
  AOI21_X1   g19983(.A1(new_n20048_), .A2(new_n20049_), .B(new_n17798_), .ZN(new_n20050_));
  NOR2_X1    g19984(.A1(new_n20045_), .A2(new_n20050_), .ZN(new_n20051_));
  OAI22_X1   g19985(.A1(new_n17801_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19364_), .ZN(new_n20052_));
  NAND2_X1   g19986(.A1(new_n17798_), .A2(new_n3312_), .ZN(new_n20053_));
  AOI21_X1   g19987(.A1(new_n20053_), .A2(new_n20052_), .B(new_n3302_), .ZN(new_n20054_));
  NAND2_X1   g19988(.A1(new_n20051_), .A2(new_n20054_), .ZN(new_n20055_));
  XOR2_X1    g19989(.A1(new_n20055_), .A2(new_n84_), .Z(new_n20056_));
  AOI21_X1   g19990(.A1(new_n19958_), .A2(new_n20012_), .B(new_n19996_), .ZN(new_n20057_));
  AOI22_X1   g19991(.A1(new_n17827_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n19321_), .ZN(new_n20058_));
  NOR2_X1    g19992(.A1(new_n19343_), .A2(new_n3175_), .ZN(new_n20059_));
  OAI21_X1   g19993(.A1(new_n20059_), .A2(new_n20058_), .B(new_n2736_), .ZN(new_n20060_));
  INV_X1     g19994(.I(new_n20060_), .ZN(new_n20061_));
  NAND3_X1   g19995(.A1(new_n19760_), .A2(new_n74_), .A3(new_n20061_), .ZN(new_n20062_));
  INV_X1     g19996(.I(new_n19760_), .ZN(new_n20063_));
  OAI21_X1   g19997(.A1(new_n20063_), .A2(new_n20060_), .B(\a[29] ), .ZN(new_n20064_));
  NAND2_X1   g19998(.A1(new_n20064_), .A2(new_n20062_), .ZN(new_n20065_));
  NAND2_X1   g19999(.A1(new_n19987_), .A2(new_n19808_), .ZN(new_n20066_));
  AOI21_X1   g20000(.A1(new_n20066_), .A2(new_n19978_), .B(new_n19980_), .ZN(new_n20067_));
  NAND2_X1   g20001(.A1(new_n19305_), .A2(new_n3332_), .ZN(new_n20068_));
  NAND2_X1   g20002(.A1(new_n17850_), .A2(new_n3189_), .ZN(new_n20069_));
  AOI21_X1   g20003(.A1(new_n19545_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n20070_));
  NAND4_X1   g20004(.A1(new_n19607_), .A2(new_n20068_), .A3(new_n20069_), .A4(new_n20070_), .ZN(new_n20071_));
  INV_X1     g20005(.I(new_n11243_), .ZN(new_n20072_));
  NOR3_X1    g20006(.A1(new_n98_), .A2(new_n235_), .A3(new_n307_), .ZN(new_n20073_));
  NAND3_X1   g20007(.A1(new_n2332_), .A2(new_n182_), .A3(new_n390_), .ZN(new_n20074_));
  NAND4_X1   g20008(.A1(new_n20074_), .A2(new_n4758_), .A3(new_n4397_), .A4(new_n20073_), .ZN(new_n20075_));
  NAND3_X1   g20009(.A1(new_n1150_), .A2(new_n3484_), .A3(new_n1968_), .ZN(new_n20076_));
  NOR4_X1    g20010(.A1(new_n10969_), .A2(new_n20075_), .A3(new_n10980_), .A4(new_n20076_), .ZN(new_n20077_));
  NAND3_X1   g20011(.A1(new_n12957_), .A2(new_n20072_), .A3(new_n20077_), .ZN(new_n20078_));
  NAND2_X1   g20012(.A1(new_n20071_), .A2(new_n20078_), .ZN(new_n20079_));
  INV_X1     g20013(.I(new_n20079_), .ZN(new_n20080_));
  NOR2_X1    g20014(.A1(new_n20071_), .A2(new_n20078_), .ZN(new_n20081_));
  NOR2_X1    g20015(.A1(new_n20080_), .A2(new_n20081_), .ZN(new_n20082_));
  XOR2_X1    g20016(.A1(new_n20071_), .A2(new_n20078_), .Z(new_n20083_));
  NAND2_X1   g20017(.A1(new_n20083_), .A2(new_n20067_), .ZN(new_n20084_));
  OAI21_X1   g20018(.A1(new_n20067_), .A2(new_n20082_), .B(new_n20084_), .ZN(new_n20085_));
  XNOR2_X1   g20019(.A1(new_n20065_), .A2(new_n20085_), .ZN(new_n20086_));
  NOR2_X1    g20020(.A1(new_n20086_), .A2(new_n20057_), .ZN(new_n20087_));
  OAI21_X1   g20021(.A1(new_n19994_), .A2(new_n19995_), .B(new_n20013_), .ZN(new_n20088_));
  NOR2_X1    g20022(.A1(new_n20082_), .A2(new_n20067_), .ZN(new_n20089_));
  AOI21_X1   g20023(.A1(new_n20067_), .A2(new_n20083_), .B(new_n20089_), .ZN(new_n20090_));
  NAND3_X1   g20024(.A1(new_n20090_), .A2(new_n20062_), .A3(new_n20064_), .ZN(new_n20091_));
  NAND2_X1   g20025(.A1(new_n20065_), .A2(new_n20085_), .ZN(new_n20092_));
  AOI21_X1   g20026(.A1(new_n20091_), .A2(new_n20092_), .B(new_n20088_), .ZN(new_n20093_));
  NOR2_X1    g20027(.A1(new_n20087_), .A2(new_n20093_), .ZN(new_n20094_));
  INV_X1     g20028(.I(new_n20094_), .ZN(new_n20095_));
  OR2_X2     g20029(.A1(new_n19892_), .A2(new_n19895_), .Z(new_n20096_));
  OAI22_X1   g20030(.A1(new_n17806_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19346_), .ZN(new_n20097_));
  NAND2_X1   g20031(.A1(new_n19359_), .A2(new_n3317_), .ZN(new_n20098_));
  AOI21_X1   g20032(.A1(new_n20098_), .A2(new_n20097_), .B(new_n3260_), .ZN(new_n20099_));
  NAND2_X1   g20033(.A1(new_n20096_), .A2(new_n20099_), .ZN(new_n20100_));
  XOR2_X1    g20034(.A1(new_n20100_), .A2(\a[26] ), .Z(new_n20101_));
  INV_X1     g20035(.I(new_n19832_), .ZN(new_n20102_));
  NAND2_X1   g20036(.A1(new_n19879_), .A2(new_n19832_), .ZN(new_n20103_));
  NAND4_X1   g20037(.A1(new_n20103_), .A2(new_n20102_), .A3(new_n20022_), .A4(new_n20023_), .ZN(new_n20104_));
  NAND2_X1   g20038(.A1(new_n20104_), .A2(new_n20101_), .ZN(new_n20105_));
  XOR2_X1    g20039(.A1(new_n20100_), .A2(new_n72_), .Z(new_n20106_));
  NOR3_X1    g20040(.A1(new_n20006_), .A2(new_n20016_), .A3(new_n19832_), .ZN(new_n20107_));
  NAND3_X1   g20041(.A1(new_n20107_), .A2(new_n20106_), .A3(new_n20103_), .ZN(new_n20108_));
  AOI21_X1   g20042(.A1(new_n20105_), .A2(new_n20108_), .B(new_n20095_), .ZN(new_n20109_));
  AOI21_X1   g20043(.A1(new_n20107_), .A2(new_n20103_), .B(new_n20106_), .ZN(new_n20110_));
  NOR2_X1    g20044(.A1(new_n20104_), .A2(new_n20101_), .ZN(new_n20111_));
  NOR3_X1    g20045(.A1(new_n20111_), .A2(new_n20110_), .A3(new_n20094_), .ZN(new_n20112_));
  NOR2_X1    g20046(.A1(new_n20112_), .A2(new_n20109_), .ZN(new_n20113_));
  NAND2_X1   g20047(.A1(new_n20113_), .A2(new_n20056_), .ZN(new_n20114_));
  XOR2_X1    g20048(.A1(new_n20055_), .A2(\a[23] ), .Z(new_n20115_));
  OAI21_X1   g20049(.A1(new_n20111_), .A2(new_n20110_), .B(new_n20094_), .ZN(new_n20116_));
  NAND3_X1   g20050(.A1(new_n20105_), .A2(new_n20095_), .A3(new_n20108_), .ZN(new_n20117_));
  NAND2_X1   g20051(.A1(new_n20116_), .A2(new_n20117_), .ZN(new_n20118_));
  NAND2_X1   g20052(.A1(new_n20118_), .A2(new_n20115_), .ZN(new_n20119_));
  NAND2_X1   g20053(.A1(new_n20114_), .A2(new_n20119_), .ZN(new_n20120_));
  NAND2_X1   g20054(.A1(new_n20120_), .A2(new_n20041_), .ZN(new_n20121_));
  NOR3_X1    g20055(.A1(new_n20109_), .A2(new_n20112_), .A3(new_n20056_), .ZN(new_n20122_));
  NOR2_X1    g20056(.A1(new_n20113_), .A2(new_n20115_), .ZN(new_n20123_));
  NOR2_X1    g20057(.A1(new_n20123_), .A2(new_n20122_), .ZN(new_n20124_));
  OAI21_X1   g20058(.A1(new_n20041_), .A2(new_n20124_), .B(new_n20121_), .ZN(new_n20125_));
  NOR2_X1    g20059(.A1(new_n19377_), .A2(new_n19386_), .ZN(new_n20126_));
  INV_X1     g20060(.I(new_n19375_), .ZN(new_n20127_));
  XOR2_X1    g20061(.A1(new_n19385_), .A2(new_n20127_), .Z(new_n20128_));
  AOI21_X1   g20062(.A1(new_n19377_), .A2(new_n19386_), .B(new_n20128_), .ZN(new_n20129_));
  INV_X1     g20063(.I(new_n20129_), .ZN(new_n20130_));
  NOR3_X1    g20064(.A1(new_n20130_), .A2(new_n17794_), .A3(new_n20126_), .ZN(new_n20131_));
  INV_X1     g20065(.I(new_n20126_), .ZN(new_n20132_));
  AOI21_X1   g20066(.A1(new_n20132_), .A2(new_n20129_), .B(new_n17793_), .ZN(new_n20133_));
  NOR2_X1    g20067(.A1(new_n20131_), .A2(new_n20133_), .ZN(new_n20134_));
  AOI22_X1   g20068(.A1(new_n19386_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n20127_), .ZN(new_n20135_));
  NOR2_X1    g20069(.A1(new_n17793_), .A2(new_n4097_), .ZN(new_n20136_));
  OAI21_X1   g20070(.A1(new_n20135_), .A2(new_n20136_), .B(new_n3773_), .ZN(new_n20137_));
  INV_X1     g20071(.I(new_n20137_), .ZN(new_n20138_));
  NAND2_X1   g20072(.A1(new_n20134_), .A2(new_n20138_), .ZN(new_n20139_));
  NOR2_X1    g20073(.A1(new_n20139_), .A2(\a[20] ), .ZN(new_n20140_));
  AOI21_X1   g20074(.A1(new_n20134_), .A2(new_n20138_), .B(new_n3035_), .ZN(new_n20141_));
  NOR2_X1    g20075(.A1(new_n20140_), .A2(new_n20141_), .ZN(new_n20142_));
  INV_X1     g20076(.I(new_n19882_), .ZN(new_n20143_));
  AOI21_X1   g20077(.A1(new_n19881_), .A2(new_n19835_), .B(new_n19543_), .ZN(new_n20144_));
  NOR4_X1    g20078(.A1(new_n19933_), .A2(new_n19936_), .A3(new_n19937_), .A4(new_n19900_), .ZN(new_n20145_));
  NAND3_X1   g20079(.A1(new_n19922_), .A2(new_n84_), .A3(new_n19923_), .ZN(new_n20146_));
  OAI21_X1   g20080(.A1(new_n19915_), .A2(new_n19918_), .B(\a[23] ), .ZN(new_n20147_));
  NAND2_X1   g20081(.A1(new_n20146_), .A2(new_n20147_), .ZN(new_n20148_));
  AOI21_X1   g20082(.A1(new_n19871_), .A2(new_n19691_), .B(new_n19864_), .ZN(new_n20149_));
  AOI21_X1   g20083(.A1(new_n19864_), .A2(new_n19928_), .B(new_n20149_), .ZN(new_n20150_));
  NOR2_X1    g20084(.A1(new_n20150_), .A2(new_n20148_), .ZN(new_n20151_));
  AOI22_X1   g20085(.A1(new_n19890_), .A2(new_n19886_), .B1(new_n19901_), .B2(new_n19902_), .ZN(new_n20152_));
  NOR3_X1    g20086(.A1(new_n20145_), .A2(new_n20152_), .A3(new_n20151_), .ZN(new_n20153_));
  OAI22_X1   g20087(.A1(new_n20143_), .A2(new_n20144_), .B1(new_n19883_), .B2(new_n20153_), .ZN(new_n20154_));
  NAND3_X1   g20088(.A1(new_n20034_), .A2(new_n20030_), .A3(new_n20037_), .ZN(new_n20155_));
  OAI21_X1   g20089(.A1(new_n20039_), .A2(new_n20038_), .B(new_n19956_), .ZN(new_n20156_));
  AOI21_X1   g20090(.A1(new_n20156_), .A2(new_n20155_), .B(new_n20154_), .ZN(new_n20157_));
  AOI21_X1   g20091(.A1(new_n20040_), .A2(new_n20035_), .B(new_n19940_), .ZN(new_n20158_));
  NOR2_X1    g20092(.A1(new_n19377_), .A2(new_n20128_), .ZN(new_n20159_));
  XOR2_X1    g20093(.A1(new_n19385_), .A2(new_n20127_), .Z(new_n20160_));
  AND2_X2    g20094(.A1(new_n19377_), .A2(new_n20160_), .Z(new_n20161_));
  OR2_X2     g20095(.A1(new_n20161_), .A2(new_n20159_), .Z(new_n20162_));
  OAI22_X1   g20096(.A1(new_n19375_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n17797_), .ZN(new_n20163_));
  NAND2_X1   g20097(.A1(new_n19386_), .A2(new_n4096_), .ZN(new_n20164_));
  AOI21_X1   g20098(.A1(new_n20164_), .A2(new_n20163_), .B(new_n4095_), .ZN(new_n20165_));
  NAND3_X1   g20099(.A1(new_n20162_), .A2(new_n3035_), .A3(new_n20165_), .ZN(new_n20166_));
  INV_X1     g20100(.I(new_n20166_), .ZN(new_n20167_));
  AOI21_X1   g20101(.A1(new_n20162_), .A2(new_n20165_), .B(new_n3035_), .ZN(new_n20168_));
  NOR2_X1    g20102(.A1(new_n20167_), .A2(new_n20168_), .ZN(new_n20169_));
  OAI21_X1   g20103(.A1(new_n20157_), .A2(new_n20158_), .B(new_n20169_), .ZN(new_n20170_));
  NAND2_X1   g20104(.A1(new_n20150_), .A2(new_n20148_), .ZN(new_n20171_));
  NOR3_X1    g20105(.A1(new_n20145_), .A2(new_n20152_), .A3(new_n20171_), .ZN(new_n20172_));
  NOR2_X1    g20106(.A1(new_n19925_), .A2(new_n19931_), .ZN(new_n20173_));
  AOI21_X1   g20107(.A1(new_n19938_), .A2(new_n19903_), .B(new_n20173_), .ZN(new_n20174_));
  INV_X1     g20108(.I(new_n20042_), .ZN(new_n20175_));
  OAI21_X1   g20109(.A1(new_n20175_), .A2(new_n20043_), .B(new_n17798_), .ZN(new_n20176_));
  NOR2_X1    g20110(.A1(new_n19369_), .A2(new_n17802_), .ZN(new_n20177_));
  NOR2_X1    g20111(.A1(new_n20047_), .A2(new_n17801_), .ZN(new_n20178_));
  OAI21_X1   g20112(.A1(new_n20178_), .A2(new_n20177_), .B(new_n17797_), .ZN(new_n20179_));
  AOI22_X1   g20113(.A1(new_n17802_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n19365_), .ZN(new_n20180_));
  NOR2_X1    g20114(.A1(new_n17797_), .A2(new_n4097_), .ZN(new_n20181_));
  OAI21_X1   g20115(.A1(new_n20181_), .A2(new_n20180_), .B(new_n3773_), .ZN(new_n20182_));
  INV_X1     g20116(.I(new_n20182_), .ZN(new_n20183_));
  NAND3_X1   g20117(.A1(new_n20176_), .A2(new_n20179_), .A3(new_n20183_), .ZN(new_n20184_));
  NOR2_X1    g20118(.A1(new_n20184_), .A2(\a[20] ), .ZN(new_n20185_));
  NOR3_X1    g20119(.A1(new_n20045_), .A2(new_n20050_), .A3(new_n20182_), .ZN(new_n20186_));
  NOR2_X1    g20120(.A1(new_n20186_), .A2(new_n3035_), .ZN(new_n20187_));
  NOR2_X1    g20121(.A1(new_n20187_), .A2(new_n20185_), .ZN(new_n20188_));
  NOR3_X1    g20122(.A1(new_n20188_), .A2(new_n20172_), .A3(new_n20174_), .ZN(new_n20189_));
  INV_X1     g20123(.I(new_n20189_), .ZN(new_n20190_));
  INV_X1     g20124(.I(new_n19884_), .ZN(new_n20191_));
  NOR2_X1    g20125(.A1(new_n20153_), .A2(new_n19543_), .ZN(new_n20192_));
  NOR2_X1    g20126(.A1(new_n19939_), .A2(new_n19883_), .ZN(new_n20193_));
  OAI21_X1   g20127(.A1(new_n20192_), .A2(new_n20193_), .B(new_n20191_), .ZN(new_n20194_));
  NAND2_X1   g20128(.A1(new_n19939_), .A2(new_n19883_), .ZN(new_n20195_));
  NAND2_X1   g20129(.A1(new_n20153_), .A2(new_n19543_), .ZN(new_n20196_));
  NAND3_X1   g20130(.A1(new_n20196_), .A2(new_n20195_), .A3(new_n19884_), .ZN(new_n20197_));
  NAND3_X1   g20131(.A1(new_n19369_), .A2(new_n17797_), .A3(new_n17802_), .ZN(new_n20198_));
  NAND2_X1   g20132(.A1(new_n20177_), .A2(new_n17798_), .ZN(new_n20199_));
  AOI21_X1   g20133(.A1(new_n20199_), .A2(new_n20198_), .B(new_n19375_), .ZN(new_n20200_));
  INV_X1     g20134(.I(new_n19370_), .ZN(new_n20201_));
  AOI21_X1   g20135(.A1(new_n20201_), .A2(new_n19376_), .B(new_n20127_), .ZN(new_n20202_));
  AOI22_X1   g20136(.A1(new_n17798_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n17802_), .ZN(new_n20203_));
  NOR2_X1    g20137(.A1(new_n19375_), .A2(new_n4097_), .ZN(new_n20204_));
  NOR2_X1    g20138(.A1(new_n20204_), .A2(new_n20203_), .ZN(new_n20205_));
  NOR4_X1    g20139(.A1(new_n20202_), .A2(new_n20200_), .A3(new_n4095_), .A4(new_n20205_), .ZN(new_n20206_));
  XOR2_X1    g20140(.A1(new_n20206_), .A2(\a[20] ), .Z(new_n20207_));
  AOI21_X1   g20141(.A1(new_n20194_), .A2(new_n20197_), .B(new_n20207_), .ZN(new_n20208_));
  NAND3_X1   g20142(.A1(new_n20194_), .A2(new_n20197_), .A3(new_n20207_), .ZN(new_n20209_));
  OAI21_X1   g20143(.A1(new_n20190_), .A2(new_n20208_), .B(new_n20209_), .ZN(new_n20210_));
  NOR3_X1    g20144(.A1(new_n20157_), .A2(new_n20158_), .A3(new_n20169_), .ZN(new_n20211_));
  OAI21_X1   g20145(.A1(new_n20210_), .A2(new_n20211_), .B(new_n20170_), .ZN(new_n20212_));
  NAND2_X1   g20146(.A1(new_n20212_), .A2(new_n20142_), .ZN(new_n20213_));
  INV_X1     g20147(.I(new_n20142_), .ZN(new_n20214_));
  AOI21_X1   g20148(.A1(new_n20196_), .A2(new_n20195_), .B(new_n19884_), .ZN(new_n20215_));
  NOR3_X1    g20149(.A1(new_n20192_), .A2(new_n20191_), .A3(new_n20193_), .ZN(new_n20216_));
  XOR2_X1    g20150(.A1(new_n20206_), .A2(new_n3035_), .Z(new_n20217_));
  OAI21_X1   g20151(.A1(new_n20216_), .A2(new_n20215_), .B(new_n20217_), .ZN(new_n20218_));
  NOR3_X1    g20152(.A1(new_n20216_), .A2(new_n20215_), .A3(new_n20217_), .ZN(new_n20219_));
  AOI21_X1   g20153(.A1(new_n20189_), .A2(new_n20218_), .B(new_n20219_), .ZN(new_n20220_));
  NOR3_X1    g20154(.A1(new_n20039_), .A2(new_n20038_), .A3(new_n19956_), .ZN(new_n20221_));
  AOI21_X1   g20155(.A1(new_n20034_), .A2(new_n20030_), .B(new_n20037_), .ZN(new_n20222_));
  OAI21_X1   g20156(.A1(new_n20222_), .A2(new_n20221_), .B(new_n19940_), .ZN(new_n20223_));
  NOR3_X1    g20157(.A1(new_n20038_), .A2(new_n20039_), .A3(new_n20037_), .ZN(new_n20224_));
  AOI21_X1   g20158(.A1(new_n20034_), .A2(new_n20030_), .B(new_n19956_), .ZN(new_n20225_));
  OAI21_X1   g20159(.A1(new_n20224_), .A2(new_n20225_), .B(new_n20154_), .ZN(new_n20226_));
  INV_X1     g20160(.I(new_n20168_), .ZN(new_n20227_));
  NAND2_X1   g20161(.A1(new_n20227_), .A2(new_n20166_), .ZN(new_n20228_));
  NAND3_X1   g20162(.A1(new_n20223_), .A2(new_n20226_), .A3(new_n20228_), .ZN(new_n20229_));
  NAND3_X1   g20163(.A1(new_n20229_), .A2(new_n20170_), .A3(new_n20220_), .ZN(new_n20230_));
  NAND3_X1   g20164(.A1(new_n20230_), .A2(new_n20214_), .A3(new_n20170_), .ZN(new_n20231_));
  AOI21_X1   g20165(.A1(new_n20231_), .A2(new_n20213_), .B(new_n20125_), .ZN(new_n20232_));
  NOR2_X1    g20166(.A1(new_n20124_), .A2(new_n20041_), .ZN(new_n20233_));
  AOI21_X1   g20167(.A1(new_n20041_), .A2(new_n20120_), .B(new_n20233_), .ZN(new_n20234_));
  AOI21_X1   g20168(.A1(new_n20230_), .A2(new_n20170_), .B(new_n20214_), .ZN(new_n20235_));
  NOR2_X1    g20169(.A1(new_n20212_), .A2(new_n20142_), .ZN(new_n20236_));
  NOR3_X1    g20170(.A1(new_n20235_), .A2(new_n20236_), .A3(new_n20234_), .ZN(new_n20237_));
  NOR2_X1    g20171(.A1(new_n20232_), .A2(new_n20237_), .ZN(new_n20238_));
  NOR2_X1    g20172(.A1(new_n19396_), .A2(new_n19399_), .ZN(new_n20239_));
  INV_X1     g20173(.I(new_n19389_), .ZN(new_n20240_));
  NAND2_X1   g20174(.A1(new_n20240_), .A2(new_n17793_), .ZN(new_n20241_));
  NAND2_X1   g20175(.A1(new_n19389_), .A2(new_n17794_), .ZN(new_n20242_));
  NAND2_X1   g20176(.A1(new_n20242_), .A2(new_n19393_), .ZN(new_n20243_));
  NAND2_X1   g20177(.A1(new_n20243_), .A2(new_n20241_), .ZN(new_n20244_));
  NOR2_X1    g20178(.A1(new_n20244_), .A2(new_n19400_), .ZN(new_n20245_));
  XOR2_X1    g20179(.A1(new_n19399_), .A2(new_n19393_), .Z(new_n20246_));
  NOR4_X1    g20180(.A1(new_n20245_), .A2(new_n17790_), .A3(new_n20239_), .A4(new_n20246_), .ZN(new_n20247_));
  INV_X1     g20181(.I(new_n20239_), .ZN(new_n20248_));
  NOR2_X1    g20182(.A1(new_n20245_), .A2(new_n20246_), .ZN(new_n20249_));
  AOI21_X1   g20183(.A1(new_n20249_), .A2(new_n20248_), .B(new_n17789_), .ZN(new_n20250_));
  NOR2_X1    g20184(.A1(new_n20250_), .A2(new_n20247_), .ZN(new_n20251_));
  OAI22_X1   g20185(.A1(new_n19400_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19393_), .ZN(new_n20252_));
  NAND2_X1   g20186(.A1(new_n17790_), .A2(new_n4469_), .ZN(new_n20253_));
  AOI21_X1   g20187(.A1(new_n20253_), .A2(new_n20252_), .B(new_n4468_), .ZN(new_n20254_));
  NAND3_X1   g20188(.A1(new_n20251_), .A2(new_n3372_), .A3(new_n20254_), .ZN(new_n20255_));
  NAND2_X1   g20189(.A1(new_n20251_), .A2(new_n20254_), .ZN(new_n20256_));
  NAND2_X1   g20190(.A1(new_n20256_), .A2(\a[17] ), .ZN(new_n20257_));
  NAND2_X1   g20191(.A1(new_n20257_), .A2(new_n20255_), .ZN(new_n20258_));
  AOI21_X1   g20192(.A1(new_n20223_), .A2(new_n20226_), .B(new_n20228_), .ZN(new_n20259_));
  OAI21_X1   g20193(.A1(new_n20259_), .A2(new_n20211_), .B(new_n20210_), .ZN(new_n20260_));
  INV_X1     g20194(.I(new_n20246_), .ZN(new_n20261_));
  OAI21_X1   g20195(.A1(new_n19395_), .A2(new_n19390_), .B(new_n20261_), .ZN(new_n20262_));
  XOR2_X1    g20196(.A1(new_n19399_), .A2(new_n19394_), .Z(new_n20263_));
  OAI21_X1   g20197(.A1(new_n20244_), .A2(new_n20263_), .B(new_n20262_), .ZN(new_n20264_));
  OAI22_X1   g20198(.A1(new_n19393_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n17793_), .ZN(new_n20265_));
  NAND2_X1   g20199(.A1(new_n19399_), .A2(new_n4469_), .ZN(new_n20266_));
  AOI21_X1   g20200(.A1(new_n20266_), .A2(new_n20265_), .B(new_n4468_), .ZN(new_n20267_));
  NAND2_X1   g20201(.A1(new_n20264_), .A2(new_n20267_), .ZN(new_n20268_));
  XOR2_X1    g20202(.A1(new_n20268_), .A2(\a[17] ), .Z(new_n20269_));
  NAND3_X1   g20203(.A1(new_n20260_), .A2(new_n20230_), .A3(new_n20269_), .ZN(new_n20270_));
  INV_X1     g20204(.I(new_n20270_), .ZN(new_n20271_));
  NOR3_X1    g20205(.A1(new_n20259_), .A2(new_n20211_), .A3(new_n20210_), .ZN(new_n20272_));
  AOI21_X1   g20206(.A1(new_n20229_), .A2(new_n20170_), .B(new_n20220_), .ZN(new_n20273_));
  XOR2_X1    g20207(.A1(new_n20268_), .A2(new_n3372_), .Z(new_n20274_));
  OAI21_X1   g20208(.A1(new_n20273_), .A2(new_n20272_), .B(new_n20274_), .ZN(new_n20275_));
  NAND2_X1   g20209(.A1(new_n20275_), .A2(new_n20270_), .ZN(new_n20276_));
  AOI21_X1   g20210(.A1(new_n20218_), .A2(new_n20209_), .B(new_n20190_), .ZN(new_n20277_));
  NAND3_X1   g20211(.A1(new_n20194_), .A2(new_n20197_), .A3(new_n20217_), .ZN(new_n20278_));
  OAI21_X1   g20212(.A1(new_n20216_), .A2(new_n20215_), .B(new_n20207_), .ZN(new_n20279_));
  AOI21_X1   g20213(.A1(new_n20279_), .A2(new_n20278_), .B(new_n20189_), .ZN(new_n20280_));
  NOR2_X1    g20214(.A1(new_n20240_), .A2(new_n17794_), .ZN(new_n20281_));
  NOR2_X1    g20215(.A1(new_n19389_), .A2(new_n17793_), .ZN(new_n20282_));
  OAI21_X1   g20216(.A1(new_n20281_), .A2(new_n20282_), .B(new_n19394_), .ZN(new_n20283_));
  INV_X1     g20217(.I(new_n20242_), .ZN(new_n20284_));
  OAI21_X1   g20218(.A1(new_n20284_), .A2(new_n19390_), .B(new_n19393_), .ZN(new_n20285_));
  AOI22_X1   g20219(.A1(new_n19386_), .A2(new_n4292_), .B1(new_n4298_), .B2(new_n17794_), .ZN(new_n20286_));
  NOR2_X1    g20220(.A1(new_n19393_), .A2(new_n4470_), .ZN(new_n20287_));
  OAI21_X1   g20221(.A1(new_n20286_), .A2(new_n20287_), .B(new_n4295_), .ZN(new_n20288_));
  INV_X1     g20222(.I(new_n20288_), .ZN(new_n20289_));
  NAND4_X1   g20223(.A1(new_n20283_), .A2(new_n20285_), .A3(new_n3372_), .A4(new_n20289_), .ZN(new_n20290_));
  NAND2_X1   g20224(.A1(new_n20283_), .A2(new_n20285_), .ZN(new_n20291_));
  OAI21_X1   g20225(.A1(new_n20291_), .A2(new_n20288_), .B(\a[17] ), .ZN(new_n20292_));
  NAND2_X1   g20226(.A1(new_n20292_), .A2(new_n20290_), .ZN(new_n20293_));
  NOR3_X1    g20227(.A1(new_n20277_), .A2(new_n20280_), .A3(new_n20293_), .ZN(new_n20294_));
  NAND3_X1   g20228(.A1(new_n20132_), .A2(new_n17793_), .A3(new_n20129_), .ZN(new_n20295_));
  OAI21_X1   g20229(.A1(new_n20130_), .A2(new_n20126_), .B(new_n17794_), .ZN(new_n20296_));
  OAI22_X1   g20230(.A1(new_n19385_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19375_), .ZN(new_n20297_));
  NOR2_X1    g20231(.A1(new_n17793_), .A2(new_n4470_), .ZN(new_n20298_));
  INV_X1     g20232(.I(new_n20298_), .ZN(new_n20299_));
  AOI21_X1   g20233(.A1(new_n20297_), .A2(new_n20299_), .B(new_n4468_), .ZN(new_n20300_));
  NAND3_X1   g20234(.A1(new_n20296_), .A2(new_n20295_), .A3(new_n20300_), .ZN(new_n20301_));
  NOR2_X1    g20235(.A1(new_n20301_), .A2(\a[17] ), .ZN(new_n20302_));
  INV_X1     g20236(.I(new_n20300_), .ZN(new_n20303_));
  NOR3_X1    g20237(.A1(new_n20131_), .A2(new_n20133_), .A3(new_n20303_), .ZN(new_n20304_));
  NOR2_X1    g20238(.A1(new_n20304_), .A2(new_n3372_), .ZN(new_n20305_));
  NOR2_X1    g20239(.A1(new_n20305_), .A2(new_n20302_), .ZN(new_n20306_));
  INV_X1     g20240(.I(new_n20306_), .ZN(new_n20307_));
  NOR4_X1    g20241(.A1(new_n20172_), .A2(new_n20174_), .A3(new_n20185_), .A4(new_n20187_), .ZN(new_n20308_));
  NAND3_X1   g20242(.A1(new_n19938_), .A2(new_n19903_), .A3(new_n20173_), .ZN(new_n20309_));
  OAI21_X1   g20243(.A1(new_n20145_), .A2(new_n20152_), .B(new_n20171_), .ZN(new_n20310_));
  NAND2_X1   g20244(.A1(new_n20186_), .A2(new_n3035_), .ZN(new_n20311_));
  NAND2_X1   g20245(.A1(new_n20184_), .A2(\a[20] ), .ZN(new_n20312_));
  AOI22_X1   g20246(.A1(new_n20310_), .A2(new_n20309_), .B1(new_n20311_), .B2(new_n20312_), .ZN(new_n20313_));
  NOR2_X1    g20247(.A1(new_n20308_), .A2(new_n20313_), .ZN(new_n20314_));
  NOR2_X1    g20248(.A1(new_n20307_), .A2(new_n20314_), .ZN(new_n20315_));
  OAI22_X1   g20249(.A1(new_n19356_), .A2(new_n4291_), .B1(new_n4297_), .B2(new_n19364_), .ZN(new_n20316_));
  NAND2_X1   g20250(.A1(new_n17802_), .A2(new_n4469_), .ZN(new_n20317_));
  AOI21_X1   g20251(.A1(new_n20316_), .A2(new_n20317_), .B(new_n4468_), .ZN(new_n20318_));
  NAND3_X1   g20252(.A1(new_n19951_), .A2(new_n3372_), .A3(new_n20318_), .ZN(new_n20319_));
  AOI21_X1   g20253(.A1(new_n19951_), .A2(new_n20318_), .B(new_n3372_), .ZN(new_n20320_));
  INV_X1     g20254(.I(new_n20320_), .ZN(new_n20321_));
  NAND2_X1   g20255(.A1(new_n20321_), .A2(new_n20319_), .ZN(new_n20322_));
  OAI22_X1   g20256(.A1(new_n19272_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n19275_), .ZN(new_n20323_));
  NAND2_X1   g20257(.A1(new_n17850_), .A2(new_n3312_), .ZN(new_n20324_));
  AOI21_X1   g20258(.A1(new_n20323_), .A2(new_n20324_), .B(new_n3302_), .ZN(new_n20325_));
  NAND3_X1   g20259(.A1(new_n19553_), .A2(new_n84_), .A3(new_n20325_), .ZN(new_n20326_));
  INV_X1     g20260(.I(new_n20326_), .ZN(new_n20327_));
  AOI21_X1   g20261(.A1(new_n19553_), .A2(new_n20325_), .B(new_n84_), .ZN(new_n20328_));
  OAI21_X1   g20262(.A1(new_n20327_), .A2(new_n20328_), .B(new_n19842_), .ZN(new_n20329_));
  OAI22_X1   g20263(.A1(new_n19313_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n19272_), .ZN(new_n20330_));
  OAI21_X1   g20264(.A1(new_n3780_), .A2(new_n19275_), .B(new_n20330_), .ZN(new_n20331_));
  NOR2_X1    g20265(.A1(new_n19571_), .A2(new_n3302_), .ZN(new_n20332_));
  AOI21_X1   g20266(.A1(new_n20332_), .A2(new_n20331_), .B(\a[23] ), .ZN(new_n20333_));
  NAND3_X1   g20267(.A1(new_n19564_), .A2(new_n20331_), .A3(new_n3301_), .ZN(new_n20334_));
  NOR2_X1    g20268(.A1(new_n20334_), .A2(new_n84_), .ZN(new_n20335_));
  NAND2_X1   g20269(.A1(new_n19290_), .A2(new_n3782_), .ZN(new_n20336_));
  NOR2_X1    g20270(.A1(new_n3299_), .A2(new_n3300_), .ZN(new_n20337_));
  NAND2_X1   g20271(.A1(new_n20336_), .A2(new_n20337_), .ZN(new_n20338_));
  NOR2_X1    g20272(.A1(new_n19593_), .A2(new_n20338_), .ZN(new_n20339_));
  NOR2_X1    g20273(.A1(new_n19313_), .A2(new_n3299_), .ZN(new_n20340_));
  INV_X1     g20274(.I(new_n20340_), .ZN(new_n20341_));
  NAND3_X1   g20275(.A1(new_n20339_), .A2(\a[23] ), .A3(new_n20341_), .ZN(new_n20342_));
  NOR3_X1    g20276(.A1(new_n20335_), .A2(new_n20333_), .A3(new_n20342_), .ZN(new_n20343_));
  NOR3_X1    g20277(.A1(new_n20327_), .A2(new_n19842_), .A3(new_n20328_), .ZN(new_n20344_));
  OAI21_X1   g20278(.A1(new_n20343_), .A2(new_n20344_), .B(new_n20329_), .ZN(new_n20345_));
  NAND2_X1   g20279(.A1(new_n19841_), .A2(new_n72_), .ZN(new_n20346_));
  NAND2_X1   g20280(.A1(new_n19581_), .A2(\a[26] ), .ZN(new_n20347_));
  NOR2_X1    g20281(.A1(new_n19582_), .A2(new_n72_), .ZN(new_n20348_));
  INV_X1     g20282(.I(new_n20348_), .ZN(new_n20349_));
  NAND3_X1   g20283(.A1(new_n20347_), .A2(new_n20346_), .A3(new_n20349_), .ZN(new_n20350_));
  NOR3_X1    g20284(.A1(new_n19841_), .A2(new_n72_), .A3(new_n19582_), .ZN(new_n20351_));
  INV_X1     g20285(.I(new_n20351_), .ZN(new_n20352_));
  NAND2_X1   g20286(.A1(new_n20350_), .A2(new_n20352_), .ZN(new_n20353_));
  AOI22_X1   g20287(.A1(new_n17850_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n19545_), .ZN(new_n20354_));
  AOI21_X1   g20288(.A1(new_n19305_), .A2(new_n3312_), .B(new_n20354_), .ZN(new_n20355_));
  NOR3_X1    g20289(.A1(new_n19618_), .A2(new_n3302_), .A3(new_n20355_), .ZN(new_n20356_));
  NAND2_X1   g20290(.A1(new_n20356_), .A2(new_n84_), .ZN(new_n20357_));
  NOR2_X1    g20291(.A1(new_n20355_), .A2(new_n3302_), .ZN(new_n20358_));
  NAND2_X1   g20292(.A1(new_n19607_), .A2(new_n20358_), .ZN(new_n20359_));
  NAND2_X1   g20293(.A1(new_n20359_), .A2(\a[23] ), .ZN(new_n20360_));
  NAND3_X1   g20294(.A1(new_n20357_), .A2(new_n20360_), .A3(new_n20353_), .ZN(new_n20361_));
  AOI21_X1   g20295(.A1(new_n20357_), .A2(new_n20360_), .B(new_n20353_), .ZN(new_n20362_));
  AOI21_X1   g20296(.A1(new_n20345_), .A2(new_n20361_), .B(new_n20362_), .ZN(new_n20363_));
  NOR3_X1    g20297(.A1(new_n19838_), .A2(new_n19839_), .A3(new_n19583_), .ZN(new_n20364_));
  AOI21_X1   g20298(.A1(new_n19574_), .A2(new_n19569_), .B(new_n19843_), .ZN(new_n20365_));
  NOR2_X1    g20299(.A1(new_n20364_), .A2(new_n20365_), .ZN(new_n20366_));
  OAI22_X1   g20300(.A1(new_n19304_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n17849_), .ZN(new_n20367_));
  NAND2_X1   g20301(.A1(new_n19321_), .A2(new_n3312_), .ZN(new_n20368_));
  AOI21_X1   g20302(.A1(new_n20367_), .A2(new_n20368_), .B(new_n3302_), .ZN(new_n20369_));
  NAND3_X1   g20303(.A1(new_n19647_), .A2(new_n84_), .A3(new_n20369_), .ZN(new_n20370_));
  INV_X1     g20304(.I(new_n20370_), .ZN(new_n20371_));
  AOI21_X1   g20305(.A1(new_n19647_), .A2(new_n20369_), .B(new_n84_), .ZN(new_n20372_));
  NOR3_X1    g20306(.A1(new_n20366_), .A2(new_n20371_), .A3(new_n20372_), .ZN(new_n20373_));
  OAI21_X1   g20307(.A1(new_n20371_), .A2(new_n20372_), .B(new_n20366_), .ZN(new_n20374_));
  OAI21_X1   g20308(.A1(new_n20363_), .A2(new_n20373_), .B(new_n20374_), .ZN(new_n20375_));
  NAND3_X1   g20309(.A1(new_n19559_), .A2(new_n19630_), .A3(new_n19557_), .ZN(new_n20376_));
  OAI21_X1   g20310(.A1(new_n19836_), .A2(new_n19558_), .B(new_n19544_), .ZN(new_n20377_));
  AOI21_X1   g20311(.A1(new_n20377_), .A2(new_n20376_), .B(new_n19584_), .ZN(new_n20378_));
  AOI21_X1   g20312(.A1(new_n19837_), .A2(new_n19585_), .B(new_n19844_), .ZN(new_n20379_));
  NOR2_X1    g20313(.A1(new_n20379_), .A2(new_n20378_), .ZN(new_n20380_));
  OAI22_X1   g20314(.A1(new_n19304_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n19320_), .ZN(new_n20381_));
  NAND2_X1   g20315(.A1(new_n17827_), .A2(new_n3312_), .ZN(new_n20382_));
  AOI21_X1   g20316(.A1(new_n20382_), .A2(new_n20381_), .B(new_n3302_), .ZN(new_n20383_));
  OAI21_X1   g20317(.A1(new_n19679_), .A2(new_n19682_), .B(new_n20383_), .ZN(new_n20384_));
  NOR2_X1    g20318(.A1(new_n20384_), .A2(\a[23] ), .ZN(new_n20385_));
  NAND2_X1   g20319(.A1(new_n20384_), .A2(\a[23] ), .ZN(new_n20386_));
  INV_X1     g20320(.I(new_n20386_), .ZN(new_n20387_));
  NOR3_X1    g20321(.A1(new_n20387_), .A2(new_n20380_), .A3(new_n20385_), .ZN(new_n20388_));
  NOR3_X1    g20322(.A1(new_n19836_), .A2(new_n19544_), .A3(new_n19558_), .ZN(new_n20389_));
  AOI21_X1   g20323(.A1(new_n19559_), .A2(new_n19557_), .B(new_n19630_), .ZN(new_n20390_));
  OAI21_X1   g20324(.A1(new_n20389_), .A2(new_n20390_), .B(new_n19844_), .ZN(new_n20391_));
  OAI21_X1   g20325(.A1(new_n19845_), .A2(new_n19560_), .B(new_n19584_), .ZN(new_n20392_));
  NAND2_X1   g20326(.A1(new_n20391_), .A2(new_n20392_), .ZN(new_n20393_));
  INV_X1     g20327(.I(new_n20385_), .ZN(new_n20394_));
  AOI21_X1   g20328(.A1(new_n20394_), .A2(new_n20386_), .B(new_n20393_), .ZN(new_n20395_));
  OAI21_X1   g20329(.A1(new_n20388_), .A2(new_n20395_), .B(new_n20375_), .ZN(new_n20396_));
  INV_X1     g20330(.I(new_n20328_), .ZN(new_n20397_));
  AOI21_X1   g20331(.A1(new_n20397_), .A2(new_n20326_), .B(new_n19582_), .ZN(new_n20398_));
  NAND2_X1   g20332(.A1(new_n20334_), .A2(new_n84_), .ZN(new_n20399_));
  NAND3_X1   g20333(.A1(new_n20332_), .A2(\a[23] ), .A3(new_n20331_), .ZN(new_n20400_));
  NAND3_X1   g20334(.A1(new_n19577_), .A2(new_n20336_), .A3(new_n20337_), .ZN(new_n20401_));
  NOR3_X1    g20335(.A1(new_n20401_), .A2(new_n84_), .A3(new_n20340_), .ZN(new_n20402_));
  NAND3_X1   g20336(.A1(new_n20399_), .A2(new_n20400_), .A3(new_n20402_), .ZN(new_n20403_));
  NAND3_X1   g20337(.A1(new_n20397_), .A2(new_n19582_), .A3(new_n20326_), .ZN(new_n20404_));
  AOI21_X1   g20338(.A1(new_n20403_), .A2(new_n20404_), .B(new_n20398_), .ZN(new_n20405_));
  NOR2_X1    g20339(.A1(new_n19581_), .A2(\a[26] ), .ZN(new_n20406_));
  NOR2_X1    g20340(.A1(new_n19841_), .A2(new_n72_), .ZN(new_n20407_));
  NOR3_X1    g20341(.A1(new_n20406_), .A2(new_n20407_), .A3(new_n20348_), .ZN(new_n20408_));
  NOR2_X1    g20342(.A1(new_n20408_), .A2(new_n20351_), .ZN(new_n20409_));
  NOR2_X1    g20343(.A1(new_n20359_), .A2(\a[23] ), .ZN(new_n20410_));
  NOR2_X1    g20344(.A1(new_n20356_), .A2(new_n84_), .ZN(new_n20411_));
  NOR3_X1    g20345(.A1(new_n20411_), .A2(new_n20410_), .A3(new_n20409_), .ZN(new_n20412_));
  OAI21_X1   g20346(.A1(new_n20411_), .A2(new_n20410_), .B(new_n20409_), .ZN(new_n20413_));
  OAI21_X1   g20347(.A1(new_n20405_), .A2(new_n20412_), .B(new_n20413_), .ZN(new_n20414_));
  NAND3_X1   g20348(.A1(new_n19574_), .A2(new_n19569_), .A3(new_n19843_), .ZN(new_n20415_));
  OAI21_X1   g20349(.A1(new_n19838_), .A2(new_n19839_), .B(new_n19583_), .ZN(new_n20416_));
  NAND2_X1   g20350(.A1(new_n20416_), .A2(new_n20415_), .ZN(new_n20417_));
  INV_X1     g20351(.I(new_n20372_), .ZN(new_n20418_));
  NAND3_X1   g20352(.A1(new_n20417_), .A2(new_n20418_), .A3(new_n20370_), .ZN(new_n20419_));
  AOI21_X1   g20353(.A1(new_n20370_), .A2(new_n20418_), .B(new_n20417_), .ZN(new_n20420_));
  AOI21_X1   g20354(.A1(new_n20414_), .A2(new_n20419_), .B(new_n20420_), .ZN(new_n20421_));
  NOR3_X1    g20355(.A1(new_n20387_), .A2(new_n20393_), .A3(new_n20385_), .ZN(new_n20422_));
  AOI21_X1   g20356(.A1(new_n20394_), .A2(new_n20386_), .B(new_n20380_), .ZN(new_n20423_));
  OAI21_X1   g20357(.A1(new_n20422_), .A2(new_n20423_), .B(new_n20421_), .ZN(new_n20424_));
  AOI22_X1   g20358(.A1(new_n19349_), .A2(new_n3770_), .B1(new_n3776_), .B2(new_n19350_), .ZN(new_n20425_));
  NOR2_X1    g20359(.A1(new_n17806_), .A2(new_n4097_), .ZN(new_n20426_));
  OAI21_X1   g20360(.A1(new_n20425_), .A2(new_n20426_), .B(new_n3773_), .ZN(new_n20427_));
  INV_X1     g20361(.I(new_n20427_), .ZN(new_n20428_));
  NAND3_X1   g20362(.A1(new_n19922_), .A2(new_n3035_), .A3(new_n20428_), .ZN(new_n20429_));
  OAI21_X1   g20363(.A1(new_n19915_), .A2(new_n20427_), .B(\a[20] ), .ZN(new_n20430_));
  NAND4_X1   g20364(.A1(new_n20429_), .A2(new_n20430_), .A3(new_n20424_), .A4(new_n20396_), .ZN(new_n20431_));
  INV_X1     g20365(.I(new_n20431_), .ZN(new_n20432_));
  AOI22_X1   g20366(.A1(new_n20429_), .A2(new_n20430_), .B1(new_n20424_), .B2(new_n20396_), .ZN(new_n20433_));
  NOR2_X1    g20367(.A1(new_n20432_), .A2(new_n20433_), .ZN(new_n20434_));
  NOR2_X1    g20368(.A1(new_n20322_), .A2(new_n20434_), .ZN(new_n20435_));
  OAI22_X1   g20369(.A1(new_n17806_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19346_), .ZN(new_n20436_));
  NAND2_X1   g20370(.A1(new_n19359_), .A2(new_n4469_), .ZN(new_n20437_));
  AOI21_X1   g20371(.A1(new_n20437_), .A2(new_n20436_), .B(new_n4468_), .ZN(new_n20438_));
  NAND2_X1   g20372(.A1(new_n20096_), .A2(new_n20438_), .ZN(new_n20439_));
  XOR2_X1    g20373(.A1(new_n20439_), .A2(new_n3372_), .Z(new_n20440_));
  OAI22_X1   g20374(.A1(new_n19272_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n19275_), .ZN(new_n20441_));
  NAND2_X1   g20375(.A1(new_n17850_), .A2(new_n4096_), .ZN(new_n20442_));
  AOI21_X1   g20376(.A1(new_n20441_), .A2(new_n20442_), .B(new_n4095_), .ZN(new_n20443_));
  NAND3_X1   g20377(.A1(new_n19553_), .A2(new_n3035_), .A3(new_n20443_), .ZN(new_n20444_));
  AOI21_X1   g20378(.A1(new_n19553_), .A2(new_n20443_), .B(new_n3035_), .ZN(new_n20445_));
  INV_X1     g20379(.I(new_n20445_), .ZN(new_n20446_));
  AOI21_X1   g20380(.A1(new_n20446_), .A2(new_n20444_), .B(new_n20340_), .ZN(new_n20447_));
  NAND2_X1   g20381(.A1(new_n19308_), .A2(new_n3776_), .ZN(new_n20448_));
  NAND2_X1   g20382(.A1(new_n19290_), .A2(new_n3770_), .ZN(new_n20449_));
  AOI22_X1   g20383(.A1(new_n20449_), .A2(new_n20448_), .B1(new_n4096_), .B2(new_n19545_), .ZN(new_n20450_));
  NOR3_X1    g20384(.A1(new_n19571_), .A2(new_n4095_), .A3(new_n20450_), .ZN(new_n20451_));
  NAND2_X1   g20385(.A1(new_n19290_), .A2(new_n3776_), .ZN(new_n20452_));
  NOR2_X1    g20386(.A1(new_n3762_), .A2(new_n3772_), .ZN(new_n20453_));
  NAND3_X1   g20387(.A1(new_n19577_), .A2(new_n20452_), .A3(new_n20453_), .ZN(new_n20454_));
  NOR2_X1    g20388(.A1(new_n19313_), .A2(new_n3762_), .ZN(new_n20455_));
  NOR4_X1    g20389(.A1(new_n20451_), .A2(new_n3035_), .A3(new_n20454_), .A4(new_n20455_), .ZN(new_n20456_));
  INV_X1     g20390(.I(new_n20456_), .ZN(new_n20457_));
  NAND3_X1   g20391(.A1(new_n20446_), .A2(new_n20340_), .A3(new_n20444_), .ZN(new_n20458_));
  AOI21_X1   g20392(.A1(new_n20457_), .A2(new_n20458_), .B(new_n20447_), .ZN(new_n20459_));
  NOR2_X1    g20393(.A1(new_n20401_), .A2(\a[23] ), .ZN(new_n20460_));
  NOR2_X1    g20394(.A1(new_n20339_), .A2(new_n84_), .ZN(new_n20461_));
  NOR2_X1    g20395(.A1(new_n20340_), .A2(new_n84_), .ZN(new_n20462_));
  NOR3_X1    g20396(.A1(new_n20460_), .A2(new_n20461_), .A3(new_n20462_), .ZN(new_n20463_));
  NOR3_X1    g20397(.A1(new_n20339_), .A2(new_n84_), .A3(new_n20340_), .ZN(new_n20464_));
  NOR2_X1    g20398(.A1(new_n20463_), .A2(new_n20464_), .ZN(new_n20465_));
  AOI22_X1   g20399(.A1(new_n17850_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n19545_), .ZN(new_n20466_));
  AOI21_X1   g20400(.A1(new_n19305_), .A2(new_n4096_), .B(new_n20466_), .ZN(new_n20467_));
  NOR2_X1    g20401(.A1(new_n20467_), .A2(new_n4095_), .ZN(new_n20468_));
  NAND2_X1   g20402(.A1(new_n19607_), .A2(new_n20468_), .ZN(new_n20469_));
  NOR2_X1    g20403(.A1(new_n20469_), .A2(\a[20] ), .ZN(new_n20470_));
  NOR3_X1    g20404(.A1(new_n19618_), .A2(new_n4095_), .A3(new_n20467_), .ZN(new_n20471_));
  NOR2_X1    g20405(.A1(new_n20471_), .A2(new_n3035_), .ZN(new_n20472_));
  NOR3_X1    g20406(.A1(new_n20472_), .A2(new_n20470_), .A3(new_n20465_), .ZN(new_n20473_));
  OAI21_X1   g20407(.A1(new_n20472_), .A2(new_n20470_), .B(new_n20465_), .ZN(new_n20474_));
  OAI21_X1   g20408(.A1(new_n20459_), .A2(new_n20473_), .B(new_n20474_), .ZN(new_n20475_));
  NAND3_X1   g20409(.A1(new_n20399_), .A2(new_n20400_), .A3(new_n20342_), .ZN(new_n20476_));
  OAI21_X1   g20410(.A1(new_n20335_), .A2(new_n20333_), .B(new_n20402_), .ZN(new_n20477_));
  NAND2_X1   g20411(.A1(new_n20477_), .A2(new_n20476_), .ZN(new_n20478_));
  OAI22_X1   g20412(.A1(new_n19304_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n17849_), .ZN(new_n20479_));
  NAND2_X1   g20413(.A1(new_n19321_), .A2(new_n4096_), .ZN(new_n20480_));
  AOI21_X1   g20414(.A1(new_n20479_), .A2(new_n20480_), .B(new_n4095_), .ZN(new_n20481_));
  NAND3_X1   g20415(.A1(new_n19647_), .A2(new_n3035_), .A3(new_n20481_), .ZN(new_n20482_));
  AOI21_X1   g20416(.A1(new_n19647_), .A2(new_n20481_), .B(new_n3035_), .ZN(new_n20483_));
  INV_X1     g20417(.I(new_n20483_), .ZN(new_n20484_));
  NAND3_X1   g20418(.A1(new_n20484_), .A2(new_n20478_), .A3(new_n20482_), .ZN(new_n20485_));
  AOI21_X1   g20419(.A1(new_n20484_), .A2(new_n20482_), .B(new_n20478_), .ZN(new_n20486_));
  AOI21_X1   g20420(.A1(new_n20475_), .A2(new_n20485_), .B(new_n20486_), .ZN(new_n20487_));
  NOR3_X1    g20421(.A1(new_n20327_), .A2(new_n19582_), .A3(new_n20328_), .ZN(new_n20488_));
  AOI21_X1   g20422(.A1(new_n20397_), .A2(new_n20326_), .B(new_n19842_), .ZN(new_n20489_));
  OAI21_X1   g20423(.A1(new_n20488_), .A2(new_n20489_), .B(new_n20343_), .ZN(new_n20490_));
  OAI21_X1   g20424(.A1(new_n20344_), .A2(new_n20398_), .B(new_n20403_), .ZN(new_n20491_));
  NAND2_X1   g20425(.A1(new_n20490_), .A2(new_n20491_), .ZN(new_n20492_));
  OAI22_X1   g20426(.A1(new_n19304_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n19320_), .ZN(new_n20493_));
  NAND2_X1   g20427(.A1(new_n17827_), .A2(new_n4096_), .ZN(new_n20494_));
  AOI21_X1   g20428(.A1(new_n20494_), .A2(new_n20493_), .B(new_n4095_), .ZN(new_n20495_));
  OAI21_X1   g20429(.A1(new_n19679_), .A2(new_n19682_), .B(new_n20495_), .ZN(new_n20496_));
  NOR2_X1    g20430(.A1(new_n20496_), .A2(\a[20] ), .ZN(new_n20497_));
  NAND2_X1   g20431(.A1(new_n20496_), .A2(\a[20] ), .ZN(new_n20498_));
  INV_X1     g20432(.I(new_n20498_), .ZN(new_n20499_));
  NOR3_X1    g20433(.A1(new_n20499_), .A2(new_n20492_), .A3(new_n20497_), .ZN(new_n20500_));
  OAI21_X1   g20434(.A1(new_n20499_), .A2(new_n20497_), .B(new_n20492_), .ZN(new_n20501_));
  OAI21_X1   g20435(.A1(new_n20487_), .A2(new_n20500_), .B(new_n20501_), .ZN(new_n20502_));
  NAND3_X1   g20436(.A1(new_n20357_), .A2(new_n20360_), .A3(new_n20409_), .ZN(new_n20503_));
  OAI21_X1   g20437(.A1(new_n20411_), .A2(new_n20410_), .B(new_n20353_), .ZN(new_n20504_));
  AOI21_X1   g20438(.A1(new_n20504_), .A2(new_n20503_), .B(new_n20405_), .ZN(new_n20505_));
  AOI21_X1   g20439(.A1(new_n20413_), .A2(new_n20361_), .B(new_n20345_), .ZN(new_n20506_));
  NOR2_X1    g20440(.A1(new_n20505_), .A2(new_n20506_), .ZN(new_n20507_));
  OAI22_X1   g20441(.A1(new_n17828_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19320_), .ZN(new_n20508_));
  NAND2_X1   g20442(.A1(new_n19349_), .A2(new_n4096_), .ZN(new_n20509_));
  AOI21_X1   g20443(.A1(new_n20509_), .A2(new_n20508_), .B(new_n4095_), .ZN(new_n20510_));
  NAND3_X1   g20444(.A1(new_n19760_), .A2(new_n3035_), .A3(new_n20510_), .ZN(new_n20511_));
  OAI21_X1   g20445(.A1(new_n19744_), .A2(new_n19747_), .B(new_n20510_), .ZN(new_n20512_));
  NAND2_X1   g20446(.A1(new_n20512_), .A2(\a[20] ), .ZN(new_n20513_));
  NAND2_X1   g20447(.A1(new_n20513_), .A2(new_n20511_), .ZN(new_n20514_));
  NOR2_X1    g20448(.A1(new_n20507_), .A2(new_n20514_), .ZN(new_n20515_));
  NOR3_X1    g20449(.A1(new_n20411_), .A2(new_n20410_), .A3(new_n20353_), .ZN(new_n20516_));
  AOI21_X1   g20450(.A1(new_n20357_), .A2(new_n20360_), .B(new_n20409_), .ZN(new_n20517_));
  OAI21_X1   g20451(.A1(new_n20516_), .A2(new_n20517_), .B(new_n20345_), .ZN(new_n20518_));
  OAI21_X1   g20452(.A1(new_n20412_), .A2(new_n20362_), .B(new_n20405_), .ZN(new_n20519_));
  NAND2_X1   g20453(.A1(new_n20518_), .A2(new_n20519_), .ZN(new_n20520_));
  NOR2_X1    g20454(.A1(new_n20512_), .A2(\a[20] ), .ZN(new_n20521_));
  AOI21_X1   g20455(.A1(new_n19760_), .A2(new_n20510_), .B(new_n3035_), .ZN(new_n20522_));
  NOR2_X1    g20456(.A1(new_n20521_), .A2(new_n20522_), .ZN(new_n20523_));
  NOR2_X1    g20457(.A1(new_n20523_), .A2(new_n20520_), .ZN(new_n20524_));
  NOR2_X1    g20458(.A1(new_n20524_), .A2(new_n20515_), .ZN(new_n20525_));
  XOR2_X1    g20459(.A1(new_n20525_), .A2(new_n20502_), .Z(new_n20526_));
  NOR2_X1    g20460(.A1(new_n20440_), .A2(new_n20526_), .ZN(new_n20527_));
  NOR3_X1    g20461(.A1(new_n20417_), .A2(new_n20371_), .A3(new_n20372_), .ZN(new_n20528_));
  AOI21_X1   g20462(.A1(new_n20418_), .A2(new_n20370_), .B(new_n20366_), .ZN(new_n20529_));
  OAI21_X1   g20463(.A1(new_n20528_), .A2(new_n20529_), .B(new_n20414_), .ZN(new_n20530_));
  OAI21_X1   g20464(.A1(new_n20373_), .A2(new_n20420_), .B(new_n20363_), .ZN(new_n20531_));
  NAND2_X1   g20465(.A1(new_n20530_), .A2(new_n20531_), .ZN(new_n20532_));
  NAND2_X1   g20466(.A1(new_n20523_), .A2(new_n20520_), .ZN(new_n20533_));
  OAI21_X1   g20467(.A1(new_n20502_), .A2(new_n20524_), .B(new_n20533_), .ZN(new_n20534_));
  OR2_X2     g20468(.A1(new_n19822_), .A2(new_n19825_), .Z(new_n20535_));
  OAI22_X1   g20469(.A1(new_n3775_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n3769_), .ZN(new_n20536_));
  NAND2_X1   g20470(.A1(new_n19350_), .A2(new_n4096_), .ZN(new_n20537_));
  AOI21_X1   g20471(.A1(new_n20536_), .A2(new_n20537_), .B(new_n4095_), .ZN(new_n20538_));
  NAND2_X1   g20472(.A1(new_n20535_), .A2(new_n20538_), .ZN(new_n20539_));
  NOR2_X1    g20473(.A1(new_n20539_), .A2(\a[20] ), .ZN(new_n20540_));
  AOI21_X1   g20474(.A1(new_n20535_), .A2(new_n20538_), .B(new_n3035_), .ZN(new_n20541_));
  NOR2_X1    g20475(.A1(new_n20540_), .A2(new_n20541_), .ZN(new_n20542_));
  NAND2_X1   g20476(.A1(new_n20534_), .A2(new_n20542_), .ZN(new_n20543_));
  INV_X1     g20477(.I(new_n20444_), .ZN(new_n20544_));
  OAI21_X1   g20478(.A1(new_n20544_), .A2(new_n20445_), .B(new_n20341_), .ZN(new_n20545_));
  NOR3_X1    g20479(.A1(new_n20544_), .A2(new_n20341_), .A3(new_n20445_), .ZN(new_n20546_));
  OAI21_X1   g20480(.A1(new_n20456_), .A2(new_n20546_), .B(new_n20545_), .ZN(new_n20547_));
  NAND2_X1   g20481(.A1(new_n20339_), .A2(new_n84_), .ZN(new_n20548_));
  NAND2_X1   g20482(.A1(new_n20401_), .A2(\a[23] ), .ZN(new_n20549_));
  INV_X1     g20483(.I(new_n20462_), .ZN(new_n20550_));
  NAND3_X1   g20484(.A1(new_n20549_), .A2(new_n20548_), .A3(new_n20550_), .ZN(new_n20551_));
  INV_X1     g20485(.I(new_n20464_), .ZN(new_n20552_));
  NAND2_X1   g20486(.A1(new_n20551_), .A2(new_n20552_), .ZN(new_n20553_));
  NAND2_X1   g20487(.A1(new_n20471_), .A2(new_n3035_), .ZN(new_n20554_));
  NAND2_X1   g20488(.A1(new_n20469_), .A2(\a[20] ), .ZN(new_n20555_));
  NAND3_X1   g20489(.A1(new_n20554_), .A2(new_n20555_), .A3(new_n20553_), .ZN(new_n20556_));
  AOI21_X1   g20490(.A1(new_n20554_), .A2(new_n20555_), .B(new_n20553_), .ZN(new_n20557_));
  AOI21_X1   g20491(.A1(new_n20547_), .A2(new_n20556_), .B(new_n20557_), .ZN(new_n20558_));
  INV_X1     g20492(.I(new_n20485_), .ZN(new_n20559_));
  NOR3_X1    g20493(.A1(new_n20335_), .A2(new_n20333_), .A3(new_n20402_), .ZN(new_n20560_));
  AOI21_X1   g20494(.A1(new_n20399_), .A2(new_n20400_), .B(new_n20342_), .ZN(new_n20561_));
  NOR2_X1    g20495(.A1(new_n20560_), .A2(new_n20561_), .ZN(new_n20562_));
  INV_X1     g20496(.I(new_n20482_), .ZN(new_n20563_));
  OAI21_X1   g20497(.A1(new_n20563_), .A2(new_n20483_), .B(new_n20562_), .ZN(new_n20564_));
  OAI21_X1   g20498(.A1(new_n20559_), .A2(new_n20558_), .B(new_n20564_), .ZN(new_n20565_));
  NAND3_X1   g20499(.A1(new_n20397_), .A2(new_n19842_), .A3(new_n20326_), .ZN(new_n20566_));
  OAI21_X1   g20500(.A1(new_n20327_), .A2(new_n20328_), .B(new_n19582_), .ZN(new_n20567_));
  AOI21_X1   g20501(.A1(new_n20567_), .A2(new_n20566_), .B(new_n20403_), .ZN(new_n20568_));
  AOI21_X1   g20502(.A1(new_n20329_), .A2(new_n20404_), .B(new_n20343_), .ZN(new_n20569_));
  NOR2_X1    g20503(.A1(new_n20569_), .A2(new_n20568_), .ZN(new_n20570_));
  INV_X1     g20504(.I(new_n20497_), .ZN(new_n20571_));
  NAND3_X1   g20505(.A1(new_n20571_), .A2(new_n20570_), .A3(new_n20498_), .ZN(new_n20572_));
  AOI21_X1   g20506(.A1(new_n20571_), .A2(new_n20498_), .B(new_n20570_), .ZN(new_n20573_));
  AOI21_X1   g20507(.A1(new_n20565_), .A2(new_n20572_), .B(new_n20573_), .ZN(new_n20574_));
  NAND2_X1   g20508(.A1(new_n20507_), .A2(new_n20514_), .ZN(new_n20575_));
  AOI21_X1   g20509(.A1(new_n20574_), .A2(new_n20575_), .B(new_n20515_), .ZN(new_n20576_));
  XOR2_X1    g20510(.A1(new_n20539_), .A2(new_n3035_), .Z(new_n20577_));
  NAND2_X1   g20511(.A1(new_n20576_), .A2(new_n20577_), .ZN(new_n20578_));
  AOI21_X1   g20512(.A1(new_n20578_), .A2(new_n20543_), .B(new_n20532_), .ZN(new_n20579_));
  INV_X1     g20513(.I(new_n20532_), .ZN(new_n20580_));
  NOR2_X1    g20514(.A1(new_n20576_), .A2(new_n20577_), .ZN(new_n20581_));
  NOR2_X1    g20515(.A1(new_n20534_), .A2(new_n20542_), .ZN(new_n20582_));
  NOR3_X1    g20516(.A1(new_n20581_), .A2(new_n20582_), .A3(new_n20580_), .ZN(new_n20583_));
  INV_X1     g20517(.I(new_n19532_), .ZN(new_n20584_));
  AOI21_X1   g20518(.A1(new_n20584_), .A2(new_n19529_), .B(new_n19364_), .ZN(new_n20585_));
  INV_X1     g20519(.I(new_n19534_), .ZN(new_n20586_));
  AOI21_X1   g20520(.A1(new_n20586_), .A2(new_n19535_), .B(new_n19365_), .ZN(new_n20587_));
  OAI22_X1   g20521(.A1(new_n19356_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n17806_), .ZN(new_n20588_));
  NAND2_X1   g20522(.A1(new_n19365_), .A2(new_n4469_), .ZN(new_n20589_));
  AOI21_X1   g20523(.A1(new_n20588_), .A2(new_n20589_), .B(new_n4468_), .ZN(new_n20590_));
  OAI21_X1   g20524(.A1(new_n20585_), .A2(new_n20587_), .B(new_n20590_), .ZN(new_n20591_));
  NOR2_X1    g20525(.A1(new_n20591_), .A2(\a[17] ), .ZN(new_n20592_));
  AOI21_X1   g20526(.A1(new_n19538_), .A2(new_n20590_), .B(new_n3372_), .ZN(new_n20593_));
  OR2_X2     g20527(.A1(new_n20592_), .A2(new_n20593_), .Z(new_n20594_));
  NOR3_X1    g20528(.A1(new_n20579_), .A2(new_n20583_), .A3(new_n20594_), .ZN(new_n20595_));
  OAI21_X1   g20529(.A1(new_n20581_), .A2(new_n20582_), .B(new_n20580_), .ZN(new_n20596_));
  NAND3_X1   g20530(.A1(new_n20578_), .A2(new_n20543_), .A3(new_n20532_), .ZN(new_n20597_));
  NOR2_X1    g20531(.A1(new_n20592_), .A2(new_n20593_), .ZN(new_n20598_));
  AOI21_X1   g20532(.A1(new_n20596_), .A2(new_n20597_), .B(new_n20598_), .ZN(new_n20599_));
  NOR3_X1    g20533(.A1(new_n20595_), .A2(new_n20599_), .A3(new_n20527_), .ZN(new_n20600_));
  INV_X1     g20534(.I(new_n20319_), .ZN(new_n20601_));
  OAI21_X1   g20535(.A1(new_n20601_), .A2(new_n20320_), .B(new_n20434_), .ZN(new_n20602_));
  INV_X1     g20536(.I(new_n20396_), .ZN(new_n20603_));
  NAND3_X1   g20537(.A1(new_n20394_), .A2(new_n20380_), .A3(new_n20386_), .ZN(new_n20604_));
  OAI21_X1   g20538(.A1(new_n20385_), .A2(new_n20387_), .B(new_n20393_), .ZN(new_n20605_));
  AOI21_X1   g20539(.A1(new_n20604_), .A2(new_n20605_), .B(new_n20375_), .ZN(new_n20606_));
  NOR3_X1    g20540(.A1(new_n19915_), .A2(\a[20] ), .A3(new_n20427_), .ZN(new_n20607_));
  AOI21_X1   g20541(.A1(new_n19922_), .A2(new_n20428_), .B(new_n3035_), .ZN(new_n20608_));
  OAI22_X1   g20542(.A1(new_n20603_), .A2(new_n20606_), .B1(new_n20608_), .B2(new_n20607_), .ZN(new_n20609_));
  NAND2_X1   g20543(.A1(new_n20609_), .A2(new_n20431_), .ZN(new_n20610_));
  NAND3_X1   g20544(.A1(new_n20321_), .A2(new_n20610_), .A3(new_n20319_), .ZN(new_n20611_));
  AOI21_X1   g20545(.A1(new_n20602_), .A2(new_n20611_), .B(new_n20595_), .ZN(new_n20612_));
  AOI21_X1   g20546(.A1(new_n20612_), .A2(new_n20600_), .B(new_n20435_), .ZN(new_n20613_));
  NAND2_X1   g20547(.A1(new_n20424_), .A2(new_n20396_), .ZN(new_n20614_));
  NOR2_X1    g20548(.A1(new_n20608_), .A2(new_n20607_), .ZN(new_n20615_));
  NOR2_X1    g20549(.A1(new_n20615_), .A2(new_n20614_), .ZN(new_n20616_));
  OAI22_X1   g20550(.A1(new_n17806_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19346_), .ZN(new_n20617_));
  NAND2_X1   g20551(.A1(new_n19359_), .A2(new_n4096_), .ZN(new_n20618_));
  AOI21_X1   g20552(.A1(new_n20618_), .A2(new_n20617_), .B(new_n4095_), .ZN(new_n20619_));
  OAI21_X1   g20553(.A1(new_n19892_), .A2(new_n19895_), .B(new_n20619_), .ZN(new_n20620_));
  XOR2_X1    g20554(.A1(new_n20620_), .A2(new_n3035_), .Z(new_n20621_));
  AOI21_X1   g20555(.A1(new_n20375_), .A2(new_n20604_), .B(new_n20423_), .ZN(new_n20622_));
  NAND3_X1   g20556(.A1(new_n19853_), .A2(new_n19854_), .A3(new_n19600_), .ZN(new_n20623_));
  OAI21_X1   g20557(.A1(new_n19620_), .A2(new_n19612_), .B(new_n19852_), .ZN(new_n20624_));
  AOI21_X1   g20558(.A1(new_n20624_), .A2(new_n20623_), .B(new_n19586_), .ZN(new_n20625_));
  AOI21_X1   g20559(.A1(new_n19622_), .A2(new_n19855_), .B(new_n19846_), .ZN(new_n20626_));
  NOR2_X1    g20560(.A1(new_n20625_), .A2(new_n20626_), .ZN(new_n20627_));
  OAI22_X1   g20561(.A1(new_n17828_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19320_), .ZN(new_n20628_));
  NAND2_X1   g20562(.A1(new_n19349_), .A2(new_n3312_), .ZN(new_n20629_));
  AOI21_X1   g20563(.A1(new_n20629_), .A2(new_n20628_), .B(new_n3302_), .ZN(new_n20630_));
  NAND3_X1   g20564(.A1(new_n19760_), .A2(new_n84_), .A3(new_n20630_), .ZN(new_n20631_));
  OAI21_X1   g20565(.A1(new_n19744_), .A2(new_n19747_), .B(new_n20630_), .ZN(new_n20632_));
  NAND2_X1   g20566(.A1(new_n20632_), .A2(\a[23] ), .ZN(new_n20633_));
  NAND2_X1   g20567(.A1(new_n20633_), .A2(new_n20631_), .ZN(new_n20634_));
  NOR2_X1    g20568(.A1(new_n20627_), .A2(new_n20634_), .ZN(new_n20635_));
  NOR3_X1    g20569(.A1(new_n19620_), .A2(new_n19612_), .A3(new_n19852_), .ZN(new_n20636_));
  AOI21_X1   g20570(.A1(new_n19853_), .A2(new_n19854_), .B(new_n19600_), .ZN(new_n20637_));
  OAI21_X1   g20571(.A1(new_n20636_), .A2(new_n20637_), .B(new_n19846_), .ZN(new_n20638_));
  OAI21_X1   g20572(.A1(new_n19621_), .A2(new_n19856_), .B(new_n19586_), .ZN(new_n20639_));
  NAND2_X1   g20573(.A1(new_n20638_), .A2(new_n20639_), .ZN(new_n20640_));
  NOR2_X1    g20574(.A1(new_n20632_), .A2(\a[23] ), .ZN(new_n20641_));
  AOI21_X1   g20575(.A1(new_n19760_), .A2(new_n20630_), .B(new_n84_), .ZN(new_n20642_));
  NOR2_X1    g20576(.A1(new_n20641_), .A2(new_n20642_), .ZN(new_n20643_));
  NOR2_X1    g20577(.A1(new_n20643_), .A2(new_n20640_), .ZN(new_n20644_));
  OAI21_X1   g20578(.A1(new_n20635_), .A2(new_n20644_), .B(new_n20622_), .ZN(new_n20645_));
  OAI21_X1   g20579(.A1(new_n20421_), .A2(new_n20422_), .B(new_n20605_), .ZN(new_n20646_));
  NAND2_X1   g20580(.A1(new_n20643_), .A2(new_n20640_), .ZN(new_n20647_));
  NAND2_X1   g20581(.A1(new_n20627_), .A2(new_n20634_), .ZN(new_n20648_));
  NAND3_X1   g20582(.A1(new_n20646_), .A2(new_n20647_), .A3(new_n20648_), .ZN(new_n20649_));
  NAND2_X1   g20583(.A1(new_n20645_), .A2(new_n20649_), .ZN(new_n20650_));
  NOR2_X1    g20584(.A1(new_n20650_), .A2(new_n20621_), .ZN(new_n20651_));
  XOR2_X1    g20585(.A1(new_n20620_), .A2(\a[20] ), .Z(new_n20652_));
  AOI21_X1   g20586(.A1(new_n20647_), .A2(new_n20648_), .B(new_n20646_), .ZN(new_n20653_));
  NOR3_X1    g20587(.A1(new_n20622_), .A2(new_n20644_), .A3(new_n20635_), .ZN(new_n20654_));
  NOR2_X1    g20588(.A1(new_n20653_), .A2(new_n20654_), .ZN(new_n20655_));
  NOR2_X1    g20589(.A1(new_n20655_), .A2(new_n20652_), .ZN(new_n20656_));
  OAI21_X1   g20590(.A1(new_n20651_), .A2(new_n20656_), .B(new_n20616_), .ZN(new_n20657_));
  NAND2_X1   g20591(.A1(new_n20650_), .A2(new_n20652_), .ZN(new_n20658_));
  NAND2_X1   g20592(.A1(new_n20655_), .A2(new_n20621_), .ZN(new_n20659_));
  AOI21_X1   g20593(.A1(new_n20658_), .A2(new_n20659_), .B(new_n20616_), .ZN(new_n20660_));
  INV_X1     g20594(.I(new_n20660_), .ZN(new_n20661_));
  OAI22_X1   g20595(.A1(new_n17801_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19364_), .ZN(new_n20662_));
  OAI21_X1   g20596(.A1(new_n17797_), .A2(new_n4470_), .B(new_n20662_), .ZN(new_n20663_));
  NAND4_X1   g20597(.A1(new_n20176_), .A2(new_n20179_), .A3(new_n4295_), .A4(new_n20663_), .ZN(new_n20664_));
  XOR2_X1    g20598(.A1(new_n20664_), .A2(new_n3372_), .Z(new_n20665_));
  AOI21_X1   g20599(.A1(new_n20657_), .A2(new_n20661_), .B(new_n20665_), .ZN(new_n20666_));
  NAND3_X1   g20600(.A1(new_n20665_), .A2(new_n20661_), .A3(new_n20657_), .ZN(new_n20667_));
  OAI21_X1   g20601(.A1(new_n20613_), .A2(new_n20666_), .B(new_n20667_), .ZN(new_n20668_));
  NOR3_X1    g20602(.A1(new_n19637_), .A2(new_n19861_), .A3(new_n19652_), .ZN(new_n20669_));
  AOI21_X1   g20603(.A1(new_n19651_), .A2(new_n19653_), .B(new_n19860_), .ZN(new_n20670_));
  OAI21_X1   g20604(.A1(new_n20669_), .A2(new_n20670_), .B(new_n19623_), .ZN(new_n20671_));
  OAI21_X1   g20605(.A1(new_n19862_), .A2(new_n19655_), .B(new_n19857_), .ZN(new_n20672_));
  NAND2_X1   g20606(.A1(new_n20671_), .A2(new_n20672_), .ZN(new_n20673_));
  INV_X1     g20607(.I(new_n20673_), .ZN(new_n20674_));
  AOI21_X1   g20608(.A1(new_n20622_), .A2(new_n20648_), .B(new_n20635_), .ZN(new_n20675_));
  OAI22_X1   g20609(.A1(new_n3306_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n3310_), .ZN(new_n20676_));
  NAND2_X1   g20610(.A1(new_n19350_), .A2(new_n3312_), .ZN(new_n20677_));
  AOI21_X1   g20611(.A1(new_n20676_), .A2(new_n20677_), .B(new_n3302_), .ZN(new_n20678_));
  NAND2_X1   g20612(.A1(new_n20535_), .A2(new_n20678_), .ZN(new_n20679_));
  XOR2_X1    g20613(.A1(new_n20679_), .A2(new_n84_), .Z(new_n20680_));
  NOR2_X1    g20614(.A1(new_n20675_), .A2(new_n20680_), .ZN(new_n20681_));
  OAI21_X1   g20615(.A1(new_n20646_), .A2(new_n20644_), .B(new_n20647_), .ZN(new_n20682_));
  XOR2_X1    g20616(.A1(new_n20679_), .A2(\a[23] ), .Z(new_n20683_));
  NOR2_X1    g20617(.A1(new_n20682_), .A2(new_n20683_), .ZN(new_n20684_));
  OAI21_X1   g20618(.A1(new_n20681_), .A2(new_n20684_), .B(new_n20674_), .ZN(new_n20685_));
  NAND2_X1   g20619(.A1(new_n20682_), .A2(new_n20683_), .ZN(new_n20686_));
  NAND2_X1   g20620(.A1(new_n20675_), .A2(new_n20680_), .ZN(new_n20687_));
  NAND3_X1   g20621(.A1(new_n20687_), .A2(new_n20686_), .A3(new_n20673_), .ZN(new_n20688_));
  OAI22_X1   g20622(.A1(new_n19356_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n17806_), .ZN(new_n20689_));
  NAND2_X1   g20623(.A1(new_n19365_), .A2(new_n4096_), .ZN(new_n20690_));
  AOI21_X1   g20624(.A1(new_n20689_), .A2(new_n20690_), .B(new_n4095_), .ZN(new_n20691_));
  NAND3_X1   g20625(.A1(new_n19538_), .A2(new_n3035_), .A3(new_n20691_), .ZN(new_n20692_));
  INV_X1     g20626(.I(new_n20692_), .ZN(new_n20693_));
  AOI21_X1   g20627(.A1(new_n19538_), .A2(new_n20691_), .B(new_n3035_), .ZN(new_n20694_));
  NOR2_X1    g20628(.A1(new_n20693_), .A2(new_n20694_), .ZN(new_n20695_));
  NAND3_X1   g20629(.A1(new_n20685_), .A2(new_n20688_), .A3(new_n20695_), .ZN(new_n20696_));
  AOI21_X1   g20630(.A1(new_n20687_), .A2(new_n20686_), .B(new_n20673_), .ZN(new_n20697_));
  NOR3_X1    g20631(.A1(new_n20681_), .A2(new_n20684_), .A3(new_n20674_), .ZN(new_n20698_));
  INV_X1     g20632(.I(new_n20694_), .ZN(new_n20699_));
  NAND2_X1   g20633(.A1(new_n20699_), .A2(new_n20692_), .ZN(new_n20700_));
  OAI21_X1   g20634(.A1(new_n20697_), .A2(new_n20698_), .B(new_n20700_), .ZN(new_n20701_));
  NAND2_X1   g20635(.A1(new_n20429_), .A2(new_n20430_), .ZN(new_n20702_));
  NAND3_X1   g20636(.A1(new_n20702_), .A2(new_n20396_), .A3(new_n20424_), .ZN(new_n20703_));
  AOI21_X1   g20637(.A1(new_n20703_), .A2(new_n20650_), .B(new_n20652_), .ZN(new_n20704_));
  NAND3_X1   g20638(.A1(new_n20701_), .A2(new_n20696_), .A3(new_n20704_), .ZN(new_n20705_));
  INV_X1     g20639(.I(new_n20705_), .ZN(new_n20706_));
  AOI21_X1   g20640(.A1(new_n20701_), .A2(new_n20696_), .B(new_n20704_), .ZN(new_n20707_));
  INV_X1     g20641(.I(new_n20200_), .ZN(new_n20708_));
  INV_X1     g20642(.I(new_n20202_), .ZN(new_n20709_));
  OAI22_X1   g20643(.A1(new_n17797_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n17801_), .ZN(new_n20710_));
  OAI21_X1   g20644(.A1(new_n19375_), .A2(new_n4470_), .B(new_n20710_), .ZN(new_n20711_));
  NAND4_X1   g20645(.A1(new_n20709_), .A2(new_n20708_), .A3(new_n4295_), .A4(new_n20711_), .ZN(new_n20712_));
  XOR2_X1    g20646(.A1(new_n20712_), .A2(\a[17] ), .Z(new_n20713_));
  OAI21_X1   g20647(.A1(new_n20706_), .A2(new_n20707_), .B(new_n20713_), .ZN(new_n20714_));
  NOR3_X1    g20648(.A1(new_n20706_), .A2(new_n20713_), .A3(new_n20707_), .ZN(new_n20715_));
  AOI21_X1   g20649(.A1(new_n20668_), .A2(new_n20714_), .B(new_n20715_), .ZN(new_n20716_));
  OAI22_X1   g20650(.A1(new_n19375_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n17797_), .ZN(new_n20717_));
  NAND2_X1   g20651(.A1(new_n19386_), .A2(new_n4469_), .ZN(new_n20718_));
  AOI21_X1   g20652(.A1(new_n20718_), .A2(new_n20717_), .B(new_n4468_), .ZN(new_n20719_));
  NAND3_X1   g20653(.A1(new_n20162_), .A2(new_n3372_), .A3(new_n20719_), .ZN(new_n20720_));
  AOI21_X1   g20654(.A1(new_n20162_), .A2(new_n20719_), .B(new_n3372_), .ZN(new_n20721_));
  INV_X1     g20655(.I(new_n20721_), .ZN(new_n20722_));
  NAND2_X1   g20656(.A1(new_n20722_), .A2(new_n20720_), .ZN(new_n20723_));
  NAND2_X1   g20657(.A1(new_n20150_), .A2(new_n20148_), .ZN(new_n20724_));
  NAND2_X1   g20658(.A1(new_n20724_), .A2(new_n19932_), .ZN(new_n20725_));
  NOR2_X1    g20659(.A1(new_n20655_), .A2(new_n20621_), .ZN(new_n20726_));
  NOR3_X1    g20660(.A1(new_n20616_), .A2(new_n20655_), .A3(new_n20621_), .ZN(new_n20727_));
  NOR2_X1    g20661(.A1(new_n20727_), .A2(new_n20726_), .ZN(new_n20728_));
  NAND3_X1   g20662(.A1(new_n20701_), .A2(new_n20696_), .A3(new_n20728_), .ZN(new_n20729_));
  OAI22_X1   g20663(.A1(new_n19356_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n19364_), .ZN(new_n20730_));
  NAND2_X1   g20664(.A1(new_n17802_), .A2(new_n4096_), .ZN(new_n20731_));
  AOI21_X1   g20665(.A1(new_n20730_), .A2(new_n20731_), .B(new_n4095_), .ZN(new_n20732_));
  NAND3_X1   g20666(.A1(new_n19951_), .A2(new_n3035_), .A3(new_n20732_), .ZN(new_n20733_));
  NAND2_X1   g20667(.A1(new_n19951_), .A2(new_n20732_), .ZN(new_n20734_));
  NAND2_X1   g20668(.A1(new_n20734_), .A2(\a[20] ), .ZN(new_n20735_));
  NAND2_X1   g20669(.A1(new_n20735_), .A2(new_n20733_), .ZN(new_n20736_));
  INV_X1     g20670(.I(new_n20736_), .ZN(new_n20737_));
  NAND2_X1   g20671(.A1(new_n20729_), .A2(new_n20737_), .ZN(new_n20738_));
  NAND4_X1   g20672(.A1(new_n20701_), .A2(new_n20696_), .A3(new_n20728_), .A4(new_n20736_), .ZN(new_n20739_));
  AOI21_X1   g20673(.A1(new_n20738_), .A2(new_n20739_), .B(new_n20725_), .ZN(new_n20740_));
  INV_X1     g20674(.I(new_n20725_), .ZN(new_n20741_));
  NOR3_X1    g20675(.A1(new_n20697_), .A2(new_n20698_), .A3(new_n20700_), .ZN(new_n20742_));
  AOI21_X1   g20676(.A1(new_n20685_), .A2(new_n20688_), .B(new_n20695_), .ZN(new_n20743_));
  NAND3_X1   g20677(.A1(new_n20703_), .A2(new_n20650_), .A3(new_n20652_), .ZN(new_n20744_));
  NAND2_X1   g20678(.A1(new_n20744_), .A2(new_n20658_), .ZN(new_n20745_));
  NOR3_X1    g20679(.A1(new_n20742_), .A2(new_n20743_), .A3(new_n20745_), .ZN(new_n20746_));
  NOR2_X1    g20680(.A1(new_n20746_), .A2(new_n20736_), .ZN(new_n20747_));
  INV_X1     g20681(.I(new_n20739_), .ZN(new_n20748_));
  NOR3_X1    g20682(.A1(new_n20747_), .A2(new_n20748_), .A3(new_n20741_), .ZN(new_n20749_));
  NOR3_X1    g20683(.A1(new_n20749_), .A2(new_n20740_), .A3(new_n20723_), .ZN(new_n20750_));
  INV_X1     g20684(.I(new_n20720_), .ZN(new_n20751_));
  NOR2_X1    g20685(.A1(new_n20751_), .A2(new_n20721_), .ZN(new_n20752_));
  OAI21_X1   g20686(.A1(new_n20747_), .A2(new_n20748_), .B(new_n20741_), .ZN(new_n20753_));
  NAND3_X1   g20687(.A1(new_n20738_), .A2(new_n20725_), .A3(new_n20739_), .ZN(new_n20754_));
  AOI21_X1   g20688(.A1(new_n20753_), .A2(new_n20754_), .B(new_n20752_), .ZN(new_n20755_));
  OAI21_X1   g20689(.A1(new_n20750_), .A2(new_n20755_), .B(new_n20716_), .ZN(new_n20756_));
  NAND2_X1   g20690(.A1(new_n20304_), .A2(new_n3372_), .ZN(new_n20757_));
  NAND2_X1   g20691(.A1(new_n20301_), .A2(\a[17] ), .ZN(new_n20758_));
  NAND4_X1   g20692(.A1(new_n20310_), .A2(new_n20309_), .A3(new_n20311_), .A4(new_n20312_), .ZN(new_n20759_));
  OAI22_X1   g20693(.A1(new_n20172_), .A2(new_n20174_), .B1(new_n20185_), .B2(new_n20187_), .ZN(new_n20760_));
  NAND2_X1   g20694(.A1(new_n20760_), .A2(new_n20759_), .ZN(new_n20761_));
  AOI21_X1   g20695(.A1(new_n20758_), .A2(new_n20757_), .B(new_n20761_), .ZN(new_n20762_));
  NOR3_X1    g20696(.A1(new_n20314_), .A2(new_n20305_), .A3(new_n20302_), .ZN(new_n20763_));
  NOR2_X1    g20697(.A1(new_n20762_), .A2(new_n20763_), .ZN(new_n20764_));
  AOI21_X1   g20698(.A1(new_n20753_), .A2(new_n20754_), .B(new_n20723_), .ZN(new_n20765_));
  NOR2_X1    g20699(.A1(new_n20765_), .A2(new_n20764_), .ZN(new_n20766_));
  AOI21_X1   g20700(.A1(new_n20756_), .A2(new_n20766_), .B(new_n20315_), .ZN(new_n20767_));
  OAI21_X1   g20701(.A1(new_n20219_), .A2(new_n20208_), .B(new_n20189_), .ZN(new_n20768_));
  NOR3_X1    g20702(.A1(new_n20216_), .A2(new_n20215_), .A3(new_n20207_), .ZN(new_n20769_));
  AOI21_X1   g20703(.A1(new_n20194_), .A2(new_n20197_), .B(new_n20217_), .ZN(new_n20770_));
  OAI21_X1   g20704(.A1(new_n20769_), .A2(new_n20770_), .B(new_n20190_), .ZN(new_n20771_));
  AOI22_X1   g20705(.A1(new_n20768_), .A2(new_n20771_), .B1(new_n20290_), .B2(new_n20292_), .ZN(new_n20772_));
  NOR2_X1    g20706(.A1(new_n20772_), .A2(new_n20294_), .ZN(new_n20773_));
  AOI21_X1   g20707(.A1(new_n20767_), .A2(new_n20773_), .B(new_n20294_), .ZN(new_n20774_));
  NOR3_X1    g20708(.A1(new_n20774_), .A2(new_n20276_), .A3(new_n20271_), .ZN(new_n20775_));
  NOR2_X1    g20709(.A1(new_n20775_), .A2(new_n20258_), .ZN(new_n20776_));
  NAND4_X1   g20710(.A1(new_n20768_), .A2(new_n20771_), .A3(new_n20290_), .A4(new_n20292_), .ZN(new_n20777_));
  INV_X1     g20711(.I(new_n20315_), .ZN(new_n20778_));
  NOR2_X1    g20712(.A1(new_n20601_), .A2(new_n20320_), .ZN(new_n20779_));
  NAND2_X1   g20713(.A1(new_n20779_), .A2(new_n20610_), .ZN(new_n20780_));
  XOR2_X1    g20714(.A1(new_n20439_), .A2(\a[17] ), .Z(new_n20781_));
  XOR2_X1    g20715(.A1(new_n20525_), .A2(new_n20574_), .Z(new_n20782_));
  NAND2_X1   g20716(.A1(new_n20781_), .A2(new_n20782_), .ZN(new_n20783_));
  NAND3_X1   g20717(.A1(new_n20596_), .A2(new_n20597_), .A3(new_n20598_), .ZN(new_n20784_));
  OAI21_X1   g20718(.A1(new_n20579_), .A2(new_n20583_), .B(new_n20594_), .ZN(new_n20785_));
  NAND3_X1   g20719(.A1(new_n20785_), .A2(new_n20784_), .A3(new_n20783_), .ZN(new_n20786_));
  AOI21_X1   g20720(.A1(new_n20321_), .A2(new_n20319_), .B(new_n20610_), .ZN(new_n20787_));
  NOR3_X1    g20721(.A1(new_n20434_), .A2(new_n20601_), .A3(new_n20320_), .ZN(new_n20788_));
  OAI21_X1   g20722(.A1(new_n20788_), .A2(new_n20787_), .B(new_n20784_), .ZN(new_n20789_));
  OAI21_X1   g20723(.A1(new_n20789_), .A2(new_n20786_), .B(new_n20780_), .ZN(new_n20790_));
  INV_X1     g20724(.I(new_n20657_), .ZN(new_n20791_));
  XOR2_X1    g20725(.A1(new_n20664_), .A2(\a[17] ), .Z(new_n20792_));
  OAI21_X1   g20726(.A1(new_n20791_), .A2(new_n20660_), .B(new_n20792_), .ZN(new_n20793_));
  NOR3_X1    g20727(.A1(new_n20792_), .A2(new_n20791_), .A3(new_n20660_), .ZN(new_n20794_));
  AOI21_X1   g20728(.A1(new_n20790_), .A2(new_n20793_), .B(new_n20794_), .ZN(new_n20795_));
  INV_X1     g20729(.I(new_n20704_), .ZN(new_n20796_));
  OAI21_X1   g20730(.A1(new_n20742_), .A2(new_n20743_), .B(new_n20796_), .ZN(new_n20797_));
  XOR2_X1    g20731(.A1(new_n20712_), .A2(new_n3372_), .Z(new_n20798_));
  AOI21_X1   g20732(.A1(new_n20705_), .A2(new_n20797_), .B(new_n20798_), .ZN(new_n20799_));
  NAND3_X1   g20733(.A1(new_n20798_), .A2(new_n20705_), .A3(new_n20797_), .ZN(new_n20800_));
  OAI21_X1   g20734(.A1(new_n20795_), .A2(new_n20799_), .B(new_n20800_), .ZN(new_n20801_));
  NAND3_X1   g20735(.A1(new_n20753_), .A2(new_n20754_), .A3(new_n20752_), .ZN(new_n20802_));
  OAI21_X1   g20736(.A1(new_n20749_), .A2(new_n20740_), .B(new_n20723_), .ZN(new_n20803_));
  AOI21_X1   g20737(.A1(new_n20802_), .A2(new_n20803_), .B(new_n20801_), .ZN(new_n20804_));
  NOR2_X1    g20738(.A1(new_n20749_), .A2(new_n20740_), .ZN(new_n20805_));
  OAI22_X1   g20739(.A1(new_n20805_), .A2(new_n20723_), .B1(new_n20762_), .B2(new_n20763_), .ZN(new_n20806_));
  OAI21_X1   g20740(.A1(new_n20804_), .A2(new_n20806_), .B(new_n20778_), .ZN(new_n20807_));
  OAI21_X1   g20741(.A1(new_n20277_), .A2(new_n20280_), .B(new_n20293_), .ZN(new_n20808_));
  NAND2_X1   g20742(.A1(new_n20777_), .A2(new_n20808_), .ZN(new_n20809_));
  OAI21_X1   g20743(.A1(new_n20807_), .A2(new_n20809_), .B(new_n20777_), .ZN(new_n20810_));
  NAND4_X1   g20744(.A1(new_n20810_), .A2(new_n20258_), .A3(new_n20270_), .A4(new_n20275_), .ZN(new_n20811_));
  INV_X1     g20745(.I(new_n20811_), .ZN(new_n20812_));
  OAI21_X1   g20746(.A1(new_n20776_), .A2(new_n20812_), .B(new_n20238_), .ZN(new_n20813_));
  INV_X1     g20747(.I(new_n20238_), .ZN(new_n20814_));
  XOR2_X1    g20748(.A1(new_n20256_), .A2(\a[17] ), .Z(new_n20815_));
  NAND3_X1   g20749(.A1(new_n20810_), .A2(new_n20270_), .A3(new_n20275_), .ZN(new_n20816_));
  NAND2_X1   g20750(.A1(new_n20816_), .A2(new_n20815_), .ZN(new_n20817_));
  NAND3_X1   g20751(.A1(new_n20817_), .A2(new_n20814_), .A3(new_n20811_), .ZN(new_n20818_));
  NAND2_X1   g20752(.A1(new_n20813_), .A2(new_n20818_), .ZN(new_n20819_));
  NOR2_X1    g20753(.A1(new_n19409_), .A2(new_n19415_), .ZN(new_n20820_));
  INV_X1     g20754(.I(new_n20820_), .ZN(new_n20821_));
  XOR2_X1    g20755(.A1(new_n19412_), .A2(new_n19407_), .Z(new_n20822_));
  AOI21_X1   g20756(.A1(new_n19409_), .A2(new_n19415_), .B(new_n20822_), .ZN(new_n20823_));
  NAND3_X1   g20757(.A1(new_n20821_), .A2(new_n17787_), .A3(new_n20823_), .ZN(new_n20824_));
  INV_X1     g20758(.I(new_n20824_), .ZN(new_n20825_));
  AOI21_X1   g20759(.A1(new_n20821_), .A2(new_n20823_), .B(new_n17787_), .ZN(new_n20826_));
  NOR2_X1    g20760(.A1(new_n20825_), .A2(new_n20826_), .ZN(new_n20827_));
  OAI22_X1   g20761(.A1(new_n19410_), .A2(new_n6089_), .B1(new_n19412_), .B2(new_n6094_), .ZN(new_n20828_));
  NAND2_X1   g20762(.A1(new_n19439_), .A2(new_n6090_), .ZN(new_n20829_));
  AOI21_X1   g20763(.A1(new_n20829_), .A2(new_n20828_), .B(new_n6082_), .ZN(new_n20830_));
  NAND2_X1   g20764(.A1(new_n20827_), .A2(new_n20830_), .ZN(new_n20831_));
  XOR2_X1    g20765(.A1(new_n20831_), .A2(\a[14] ), .Z(new_n20832_));
  NOR2_X1    g20766(.A1(new_n20276_), .A2(new_n20810_), .ZN(new_n20833_));
  NOR2_X1    g20767(.A1(new_n20750_), .A2(new_n20755_), .ZN(new_n20834_));
  OAI21_X1   g20768(.A1(new_n20834_), .A2(new_n20801_), .B(new_n20766_), .ZN(new_n20835_));
  NAND3_X1   g20769(.A1(new_n20835_), .A2(new_n20773_), .A3(new_n20778_), .ZN(new_n20836_));
  AOI22_X1   g20770(.A1(new_n20836_), .A2(new_n20777_), .B1(new_n20270_), .B2(new_n20275_), .ZN(new_n20837_));
  AND2_X2    g20771(.A1(new_n19396_), .A2(new_n19401_), .Z(new_n20838_));
  OAI21_X1   g20772(.A1(new_n20838_), .A2(new_n19402_), .B(new_n17789_), .ZN(new_n20839_));
  NAND2_X1   g20773(.A1(new_n19403_), .A2(new_n17790_), .ZN(new_n20840_));
  NAND2_X1   g20774(.A1(new_n20840_), .A2(new_n19410_), .ZN(new_n20841_));
  NAND2_X1   g20775(.A1(new_n20841_), .A2(new_n20839_), .ZN(new_n20842_));
  INV_X1     g20776(.I(new_n20822_), .ZN(new_n20843_));
  OAI21_X1   g20777(.A1(new_n19408_), .A2(new_n19404_), .B(new_n20843_), .ZN(new_n20844_));
  XNOR2_X1   g20778(.A1(new_n19412_), .A2(new_n19407_), .ZN(new_n20845_));
  OAI21_X1   g20779(.A1(new_n20842_), .A2(new_n20845_), .B(new_n20844_), .ZN(new_n20846_));
  OAI22_X1   g20780(.A1(new_n19410_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n17789_), .ZN(new_n20847_));
  NAND2_X1   g20781(.A1(new_n19415_), .A2(new_n6090_), .ZN(new_n20848_));
  AOI21_X1   g20782(.A1(new_n20848_), .A2(new_n20847_), .B(new_n6082_), .ZN(new_n20849_));
  NAND2_X1   g20783(.A1(new_n20846_), .A2(new_n20849_), .ZN(new_n20850_));
  XOR2_X1    g20784(.A1(new_n20850_), .A2(new_n3521_), .Z(new_n20851_));
  INV_X1     g20785(.I(new_n20851_), .ZN(new_n20852_));
  OAI21_X1   g20786(.A1(new_n20833_), .A2(new_n20837_), .B(new_n20852_), .ZN(new_n20853_));
  NAND2_X1   g20787(.A1(new_n20767_), .A2(new_n20809_), .ZN(new_n20854_));
  NAND2_X1   g20788(.A1(new_n20807_), .A2(new_n20773_), .ZN(new_n20855_));
  NAND2_X1   g20789(.A1(new_n20854_), .A2(new_n20855_), .ZN(new_n20856_));
  NAND2_X1   g20790(.A1(new_n19403_), .A2(new_n17789_), .ZN(new_n20857_));
  INV_X1     g20791(.I(new_n20857_), .ZN(new_n20858_));
  NOR2_X1    g20792(.A1(new_n19403_), .A2(new_n17789_), .ZN(new_n20859_));
  OAI21_X1   g20793(.A1(new_n20858_), .A2(new_n20859_), .B(new_n19407_), .ZN(new_n20860_));
  INV_X1     g20794(.I(new_n20840_), .ZN(new_n20861_));
  OAI21_X1   g20795(.A1(new_n20861_), .A2(new_n19404_), .B(new_n19410_), .ZN(new_n20862_));
  NAND2_X1   g20796(.A1(new_n20860_), .A2(new_n20862_), .ZN(new_n20863_));
  INV_X1     g20797(.I(new_n20863_), .ZN(new_n20864_));
  OAI22_X1   g20798(.A1(new_n17789_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n19400_), .ZN(new_n20865_));
  NOR2_X1    g20799(.A1(new_n19410_), .A2(new_n6091_), .ZN(new_n20866_));
  INV_X1     g20800(.I(new_n20866_), .ZN(new_n20867_));
  AOI21_X1   g20801(.A1(new_n20867_), .A2(new_n20865_), .B(new_n6082_), .ZN(new_n20868_));
  NAND2_X1   g20802(.A1(new_n20864_), .A2(new_n20868_), .ZN(new_n20869_));
  XOR2_X1    g20803(.A1(new_n20869_), .A2(\a[14] ), .Z(new_n20870_));
  NOR2_X1    g20804(.A1(new_n20870_), .A2(new_n20856_), .ZN(new_n20871_));
  NOR3_X1    g20805(.A1(new_n20833_), .A2(new_n20837_), .A3(new_n20852_), .ZN(new_n20872_));
  OAI21_X1   g20806(.A1(new_n20871_), .A2(new_n20872_), .B(new_n20853_), .ZN(new_n20873_));
  NAND2_X1   g20807(.A1(new_n20873_), .A2(new_n20832_), .ZN(new_n20874_));
  XOR2_X1    g20808(.A1(new_n20831_), .A2(new_n3521_), .Z(new_n20875_));
  XOR2_X1    g20809(.A1(new_n20869_), .A2(new_n3521_), .Z(new_n20876_));
  NAND3_X1   g20810(.A1(new_n20876_), .A2(new_n20854_), .A3(new_n20855_), .ZN(new_n20877_));
  NAND4_X1   g20811(.A1(new_n20836_), .A2(new_n20270_), .A3(new_n20275_), .A4(new_n20777_), .ZN(new_n20878_));
  NAND2_X1   g20812(.A1(new_n20276_), .A2(new_n20810_), .ZN(new_n20879_));
  NAND3_X1   g20813(.A1(new_n20879_), .A2(new_n20878_), .A3(new_n20851_), .ZN(new_n20880_));
  NAND3_X1   g20814(.A1(new_n20853_), .A2(new_n20880_), .A3(new_n20877_), .ZN(new_n20881_));
  NAND3_X1   g20815(.A1(new_n20881_), .A2(new_n20875_), .A3(new_n20853_), .ZN(new_n20882_));
  AOI21_X1   g20816(.A1(new_n20874_), .A2(new_n20882_), .B(new_n20819_), .ZN(new_n20883_));
  AOI21_X1   g20817(.A1(new_n20817_), .A2(new_n20811_), .B(new_n20814_), .ZN(new_n20884_));
  NOR3_X1    g20818(.A1(new_n20776_), .A2(new_n20812_), .A3(new_n20238_), .ZN(new_n20885_));
  NOR2_X1    g20819(.A1(new_n20885_), .A2(new_n20884_), .ZN(new_n20886_));
  AOI21_X1   g20820(.A1(new_n20881_), .A2(new_n20853_), .B(new_n20875_), .ZN(new_n20887_));
  NOR2_X1    g20821(.A1(new_n20873_), .A2(new_n20832_), .ZN(new_n20888_));
  NOR3_X1    g20822(.A1(new_n20888_), .A2(new_n20887_), .A3(new_n20886_), .ZN(new_n20889_));
  NOR2_X1    g20823(.A1(new_n20889_), .A2(new_n20883_), .ZN(new_n20890_));
  INV_X1     g20824(.I(new_n20890_), .ZN(new_n20891_));
  OAI21_X1   g20825(.A1(new_n19440_), .A2(new_n19439_), .B(new_n19442_), .ZN(new_n20892_));
  OAI21_X1   g20826(.A1(new_n19418_), .A2(new_n17787_), .B(new_n19423_), .ZN(new_n20893_));
  NAND2_X1   g20827(.A1(new_n20893_), .A2(new_n20892_), .ZN(new_n20894_));
  OAI21_X1   g20828(.A1(new_n19443_), .A2(new_n19441_), .B(new_n19428_), .ZN(new_n20895_));
  INV_X1     g20829(.I(new_n19428_), .ZN(new_n20896_));
  NAND3_X1   g20830(.A1(new_n19424_), .A2(new_n19419_), .A3(new_n20896_), .ZN(new_n20897_));
  NAND3_X1   g20831(.A1(new_n20897_), .A2(new_n20894_), .A3(new_n20895_), .ZN(new_n20898_));
  NOR2_X1    g20832(.A1(new_n20898_), .A2(new_n19438_), .ZN(new_n20899_));
  INV_X1     g20833(.I(new_n20892_), .ZN(new_n20900_));
  AOI21_X1   g20834(.A1(new_n19440_), .A2(new_n19439_), .B(new_n19442_), .ZN(new_n20901_));
  NOR2_X1    g20835(.A1(new_n20900_), .A2(new_n20901_), .ZN(new_n20902_));
  AOI21_X1   g20836(.A1(new_n19424_), .A2(new_n19419_), .B(new_n20896_), .ZN(new_n20903_));
  NOR3_X1    g20837(.A1(new_n19443_), .A2(new_n19441_), .A3(new_n19428_), .ZN(new_n20904_));
  NOR3_X1    g20838(.A1(new_n20902_), .A2(new_n20903_), .A3(new_n20904_), .ZN(new_n20905_));
  NOR2_X1    g20839(.A1(new_n20905_), .A2(new_n17784_), .ZN(new_n20906_));
  NOR2_X1    g20840(.A1(new_n20906_), .A2(new_n20899_), .ZN(new_n20907_));
  OAI22_X1   g20841(.A1(new_n19428_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n19423_), .ZN(new_n20908_));
  NAND2_X1   g20842(.A1(new_n19438_), .A2(new_n4709_), .ZN(new_n20909_));
  AOI21_X1   g20843(.A1(new_n20909_), .A2(new_n20908_), .B(new_n4707_), .ZN(new_n20910_));
  NAND2_X1   g20844(.A1(new_n20907_), .A2(new_n20910_), .ZN(new_n20911_));
  XOR2_X1    g20845(.A1(new_n20911_), .A2(\a[11] ), .Z(new_n20912_));
  AOI21_X1   g20846(.A1(new_n20879_), .A2(new_n20878_), .B(new_n20851_), .ZN(new_n20913_));
  OAI21_X1   g20847(.A1(new_n20872_), .A2(new_n20913_), .B(new_n20871_), .ZN(new_n20914_));
  AOI21_X1   g20848(.A1(new_n20893_), .A2(new_n20892_), .B(new_n19428_), .ZN(new_n20915_));
  NAND3_X1   g20849(.A1(new_n19440_), .A2(new_n19439_), .A3(new_n19423_), .ZN(new_n20916_));
  NAND3_X1   g20850(.A1(new_n19418_), .A2(new_n17787_), .A3(new_n19442_), .ZN(new_n20917_));
  AOI21_X1   g20851(.A1(new_n20917_), .A2(new_n20916_), .B(new_n20896_), .ZN(new_n20918_));
  OAI22_X1   g20852(.A1(new_n19423_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n17787_), .ZN(new_n20919_));
  NAND2_X1   g20853(.A1(new_n20896_), .A2(new_n4709_), .ZN(new_n20920_));
  AOI21_X1   g20854(.A1(new_n20920_), .A2(new_n20919_), .B(new_n4707_), .ZN(new_n20921_));
  OAI21_X1   g20855(.A1(new_n20915_), .A2(new_n20918_), .B(new_n20921_), .ZN(new_n20922_));
  XOR2_X1    g20856(.A1(new_n20922_), .A2(\a[11] ), .Z(new_n20923_));
  NAND3_X1   g20857(.A1(new_n20914_), .A2(new_n20881_), .A3(new_n20923_), .ZN(new_n20924_));
  NOR3_X1    g20858(.A1(new_n20872_), .A2(new_n20913_), .A3(new_n20871_), .ZN(new_n20925_));
  AOI21_X1   g20859(.A1(new_n20853_), .A2(new_n20880_), .B(new_n20877_), .ZN(new_n20926_));
  INV_X1     g20860(.I(new_n20923_), .ZN(new_n20927_));
  NOR3_X1    g20861(.A1(new_n20925_), .A2(new_n20927_), .A3(new_n20926_), .ZN(new_n20928_));
  AOI21_X1   g20862(.A1(new_n20914_), .A2(new_n20881_), .B(new_n20923_), .ZN(new_n20929_));
  NOR2_X1    g20863(.A1(new_n20928_), .A2(new_n20929_), .ZN(new_n20930_));
  INV_X1     g20864(.I(new_n20856_), .ZN(new_n20931_));
  NAND2_X1   g20865(.A1(new_n20931_), .A2(new_n20870_), .ZN(new_n20932_));
  NAND2_X1   g20866(.A1(new_n20876_), .A2(new_n20856_), .ZN(new_n20933_));
  NAND2_X1   g20867(.A1(new_n19440_), .A2(new_n17787_), .ZN(new_n20934_));
  NAND2_X1   g20868(.A1(new_n19418_), .A2(new_n19439_), .ZN(new_n20935_));
  AOI21_X1   g20869(.A1(new_n20935_), .A2(new_n20934_), .B(new_n19423_), .ZN(new_n20936_));
  NAND2_X1   g20870(.A1(new_n19440_), .A2(new_n19439_), .ZN(new_n20937_));
  AOI21_X1   g20871(.A1(new_n19419_), .A2(new_n20937_), .B(new_n19442_), .ZN(new_n20938_));
  NOR2_X1    g20872(.A1(new_n20936_), .A2(new_n20938_), .ZN(new_n20939_));
  AOI22_X1   g20873(.A1(new_n19439_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n19415_), .ZN(new_n20940_));
  NOR2_X1    g20874(.A1(new_n19423_), .A2(new_n4710_), .ZN(new_n20941_));
  OAI21_X1   g20875(.A1(new_n20941_), .A2(new_n20940_), .B(new_n4706_), .ZN(new_n20942_));
  INV_X1     g20876(.I(new_n20942_), .ZN(new_n20943_));
  NAND3_X1   g20877(.A1(new_n20939_), .A2(new_n4034_), .A3(new_n20943_), .ZN(new_n20944_));
  AOI21_X1   g20878(.A1(new_n20939_), .A2(new_n20943_), .B(new_n4034_), .ZN(new_n20945_));
  INV_X1     g20879(.I(new_n20945_), .ZN(new_n20946_));
  NAND4_X1   g20880(.A1(new_n20932_), .A2(new_n20933_), .A3(new_n20944_), .A4(new_n20946_), .ZN(new_n20947_));
  NAND2_X1   g20881(.A1(new_n20821_), .A2(new_n20823_), .ZN(new_n20948_));
  NAND2_X1   g20882(.A1(new_n20948_), .A2(new_n19439_), .ZN(new_n20949_));
  OAI22_X1   g20883(.A1(new_n19410_), .A2(new_n4716_), .B1(new_n19412_), .B2(new_n4719_), .ZN(new_n20950_));
  NAND2_X1   g20884(.A1(new_n19439_), .A2(new_n4709_), .ZN(new_n20951_));
  AOI21_X1   g20885(.A1(new_n20951_), .A2(new_n20950_), .B(new_n4707_), .ZN(new_n20952_));
  NAND3_X1   g20886(.A1(new_n20949_), .A2(new_n20824_), .A3(new_n20952_), .ZN(new_n20953_));
  XOR2_X1    g20887(.A1(new_n20953_), .A2(new_n4034_), .Z(new_n20954_));
  OAI21_X1   g20888(.A1(new_n20804_), .A2(new_n20765_), .B(new_n20306_), .ZN(new_n20955_));
  INV_X1     g20889(.I(new_n20765_), .ZN(new_n20956_));
  NAND3_X1   g20890(.A1(new_n20756_), .A2(new_n20307_), .A3(new_n20956_), .ZN(new_n20957_));
  AOI21_X1   g20891(.A1(new_n20957_), .A2(new_n20955_), .B(new_n20761_), .ZN(new_n20958_));
  AOI21_X1   g20892(.A1(new_n20756_), .A2(new_n20956_), .B(new_n20307_), .ZN(new_n20959_));
  NOR3_X1    g20893(.A1(new_n20804_), .A2(new_n20306_), .A3(new_n20765_), .ZN(new_n20960_));
  NOR3_X1    g20894(.A1(new_n20959_), .A2(new_n20960_), .A3(new_n20314_), .ZN(new_n20961_));
  NOR2_X1    g20895(.A1(new_n20958_), .A2(new_n20961_), .ZN(new_n20962_));
  AOI21_X1   g20896(.A1(new_n20714_), .A2(new_n20800_), .B(new_n20795_), .ZN(new_n20963_));
  INV_X1     g20897(.I(new_n20963_), .ZN(new_n20964_));
  NAND3_X1   g20898(.A1(new_n20713_), .A2(new_n20705_), .A3(new_n20797_), .ZN(new_n20965_));
  OAI21_X1   g20899(.A1(new_n20706_), .A2(new_n20707_), .B(new_n20798_), .ZN(new_n20966_));
  NAND2_X1   g20900(.A1(new_n20966_), .A2(new_n20965_), .ZN(new_n20967_));
  NAND2_X1   g20901(.A1(new_n20967_), .A2(new_n20795_), .ZN(new_n20968_));
  AOI22_X1   g20902(.A1(new_n19386_), .A2(new_n6180_), .B1(new_n6095_), .B2(new_n17794_), .ZN(new_n20969_));
  NOR2_X1    g20903(.A1(new_n19393_), .A2(new_n6091_), .ZN(new_n20970_));
  OAI21_X1   g20904(.A1(new_n20969_), .A2(new_n20970_), .B(new_n6081_), .ZN(new_n20971_));
  NOR2_X1    g20905(.A1(new_n20291_), .A2(new_n20971_), .ZN(new_n20972_));
  XOR2_X1    g20906(.A1(new_n20972_), .A2(new_n3521_), .Z(new_n20973_));
  AOI21_X1   g20907(.A1(new_n20964_), .A2(new_n20968_), .B(new_n20973_), .ZN(new_n20974_));
  NAND3_X1   g20908(.A1(new_n20716_), .A2(new_n20803_), .A3(new_n20802_), .ZN(new_n20975_));
  OAI21_X1   g20909(.A1(new_n20750_), .A2(new_n20755_), .B(new_n20801_), .ZN(new_n20976_));
  OAI22_X1   g20910(.A1(new_n19393_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n17793_), .ZN(new_n20977_));
  NAND2_X1   g20911(.A1(new_n19399_), .A2(new_n6090_), .ZN(new_n20978_));
  AOI21_X1   g20912(.A1(new_n20978_), .A2(new_n20977_), .B(new_n6082_), .ZN(new_n20979_));
  NAND2_X1   g20913(.A1(new_n20264_), .A2(new_n20979_), .ZN(new_n20980_));
  XOR2_X1    g20914(.A1(new_n20980_), .A2(new_n3521_), .Z(new_n20981_));
  AOI21_X1   g20915(.A1(new_n20976_), .A2(new_n20975_), .B(new_n20981_), .ZN(new_n20982_));
  NOR3_X1    g20916(.A1(new_n20801_), .A2(new_n20750_), .A3(new_n20755_), .ZN(new_n20983_));
  AOI21_X1   g20917(.A1(new_n20802_), .A2(new_n20803_), .B(new_n20716_), .ZN(new_n20984_));
  XOR2_X1    g20918(.A1(new_n20980_), .A2(\a[14] ), .Z(new_n20985_));
  NOR3_X1    g20919(.A1(new_n20984_), .A2(new_n20983_), .A3(new_n20985_), .ZN(new_n20986_));
  NOR3_X1    g20920(.A1(new_n20986_), .A2(new_n20982_), .A3(new_n20974_), .ZN(new_n20987_));
  AOI22_X1   g20921(.A1(new_n19399_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n19394_), .ZN(new_n20988_));
  NOR2_X1    g20922(.A1(new_n17789_), .A2(new_n6091_), .ZN(new_n20989_));
  OAI21_X1   g20923(.A1(new_n20989_), .A2(new_n20988_), .B(new_n6081_), .ZN(new_n20990_));
  INV_X1     g20924(.I(new_n20990_), .ZN(new_n20991_));
  NAND2_X1   g20925(.A1(new_n20251_), .A2(new_n20991_), .ZN(new_n20992_));
  XOR2_X1    g20926(.A1(new_n20992_), .A2(new_n3521_), .Z(new_n20993_));
  NOR2_X1    g20927(.A1(new_n20987_), .A2(new_n20993_), .ZN(new_n20994_));
  AOI21_X1   g20928(.A1(new_n20965_), .A2(new_n20966_), .B(new_n20668_), .ZN(new_n20995_));
  XOR2_X1    g20929(.A1(new_n20972_), .A2(\a[14] ), .Z(new_n20996_));
  OAI21_X1   g20930(.A1(new_n20995_), .A2(new_n20963_), .B(new_n20996_), .ZN(new_n20997_));
  OAI21_X1   g20931(.A1(new_n20984_), .A2(new_n20983_), .B(new_n20985_), .ZN(new_n20998_));
  NAND3_X1   g20932(.A1(new_n20976_), .A2(new_n20975_), .A3(new_n20981_), .ZN(new_n20999_));
  NAND3_X1   g20933(.A1(new_n20998_), .A2(new_n20999_), .A3(new_n20997_), .ZN(new_n21000_));
  XOR2_X1    g20934(.A1(new_n20992_), .A2(\a[14] ), .Z(new_n21001_));
  NOR2_X1    g20935(.A1(new_n21000_), .A2(new_n21001_), .ZN(new_n21002_));
  OAI21_X1   g20936(.A1(new_n20994_), .A2(new_n21002_), .B(new_n20962_), .ZN(new_n21003_));
  OAI21_X1   g20937(.A1(new_n20959_), .A2(new_n20960_), .B(new_n20314_), .ZN(new_n21004_));
  NAND3_X1   g20938(.A1(new_n20957_), .A2(new_n20955_), .A3(new_n20761_), .ZN(new_n21005_));
  NAND2_X1   g20939(.A1(new_n21004_), .A2(new_n21005_), .ZN(new_n21006_));
  NAND2_X1   g20940(.A1(new_n21000_), .A2(new_n21001_), .ZN(new_n21007_));
  NAND2_X1   g20941(.A1(new_n20987_), .A2(new_n20993_), .ZN(new_n21008_));
  NAND3_X1   g20942(.A1(new_n21006_), .A2(new_n21008_), .A3(new_n21007_), .ZN(new_n21009_));
  NAND3_X1   g20943(.A1(new_n21003_), .A2(new_n21009_), .A3(new_n20954_), .ZN(new_n21010_));
  XOR2_X1    g20944(.A1(new_n20953_), .A2(\a[11] ), .Z(new_n21011_));
  AOI21_X1   g20945(.A1(new_n21007_), .A2(new_n21008_), .B(new_n21006_), .ZN(new_n21012_));
  NOR3_X1    g20946(.A1(new_n20962_), .A2(new_n20994_), .A3(new_n21002_), .ZN(new_n21013_));
  OAI21_X1   g20947(.A1(new_n21012_), .A2(new_n21013_), .B(new_n21011_), .ZN(new_n21014_));
  OAI22_X1   g20948(.A1(new_n19410_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n17789_), .ZN(new_n21015_));
  NAND2_X1   g20949(.A1(new_n19415_), .A2(new_n4709_), .ZN(new_n21016_));
  AOI21_X1   g20950(.A1(new_n21016_), .A2(new_n21015_), .B(new_n4707_), .ZN(new_n21017_));
  NAND3_X1   g20951(.A1(new_n20846_), .A2(new_n4034_), .A3(new_n21017_), .ZN(new_n21018_));
  AOI21_X1   g20952(.A1(new_n20846_), .A2(new_n21017_), .B(new_n4034_), .ZN(new_n21019_));
  INV_X1     g20953(.I(new_n21019_), .ZN(new_n21020_));
  NAND2_X1   g20954(.A1(new_n21020_), .A2(new_n21018_), .ZN(new_n21021_));
  NAND3_X1   g20955(.A1(new_n20998_), .A2(new_n20999_), .A3(new_n20974_), .ZN(new_n21022_));
  OAI21_X1   g20956(.A1(new_n20986_), .A2(new_n20982_), .B(new_n20997_), .ZN(new_n21023_));
  AOI21_X1   g20957(.A1(new_n21023_), .A2(new_n21022_), .B(new_n21021_), .ZN(new_n21024_));
  INV_X1     g20958(.I(new_n21024_), .ZN(new_n21025_));
  INV_X1     g20959(.I(new_n21018_), .ZN(new_n21026_));
  NOR2_X1    g20960(.A1(new_n21026_), .A2(new_n21019_), .ZN(new_n21027_));
  NAND3_X1   g20961(.A1(new_n21023_), .A2(new_n21022_), .A3(new_n21027_), .ZN(new_n21028_));
  NOR3_X1    g20962(.A1(new_n20986_), .A2(new_n20982_), .A3(new_n20997_), .ZN(new_n21029_));
  AOI21_X1   g20963(.A1(new_n20998_), .A2(new_n20999_), .B(new_n20974_), .ZN(new_n21030_));
  OAI21_X1   g20964(.A1(new_n21029_), .A2(new_n21030_), .B(new_n21021_), .ZN(new_n21031_));
  NOR3_X1    g20965(.A1(new_n20996_), .A2(new_n20995_), .A3(new_n20963_), .ZN(new_n21032_));
  AOI21_X1   g20966(.A1(new_n20964_), .A2(new_n20968_), .B(new_n20973_), .ZN(new_n21033_));
  OAI22_X1   g20967(.A1(new_n17789_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n19400_), .ZN(new_n21034_));
  OAI21_X1   g20968(.A1(new_n4710_), .A2(new_n19410_), .B(new_n21034_), .ZN(new_n21035_));
  NAND4_X1   g20969(.A1(new_n20860_), .A2(new_n20862_), .A3(new_n4706_), .A4(new_n21035_), .ZN(new_n21036_));
  XOR2_X1    g20970(.A1(new_n21036_), .A2(\a[11] ), .Z(new_n21037_));
  NOR3_X1    g20971(.A1(new_n21037_), .A2(new_n21032_), .A3(new_n21033_), .ZN(new_n21038_));
  NAND3_X1   g20972(.A1(new_n21031_), .A2(new_n21028_), .A3(new_n21038_), .ZN(new_n21039_));
  NAND2_X1   g20973(.A1(new_n21039_), .A2(new_n21025_), .ZN(new_n21040_));
  AOI22_X1   g20974(.A1(new_n21014_), .A2(new_n21010_), .B1(new_n20954_), .B2(new_n21040_), .ZN(new_n21041_));
  NOR2_X1    g20975(.A1(new_n20876_), .A2(new_n20856_), .ZN(new_n21042_));
  INV_X1     g20976(.I(new_n20933_), .ZN(new_n21043_));
  INV_X1     g20977(.I(new_n20944_), .ZN(new_n21044_));
  OAI22_X1   g20978(.A1(new_n21043_), .A2(new_n21042_), .B1(new_n21044_), .B2(new_n20945_), .ZN(new_n21045_));
  NAND2_X1   g20979(.A1(new_n21045_), .A2(new_n20947_), .ZN(new_n21046_));
  OAI21_X1   g20980(.A1(new_n21041_), .A2(new_n21046_), .B(new_n20947_), .ZN(new_n21047_));
  NAND3_X1   g20981(.A1(new_n21047_), .A2(new_n20924_), .A3(new_n20930_), .ZN(new_n21048_));
  NAND2_X1   g20982(.A1(new_n21048_), .A2(new_n20912_), .ZN(new_n21049_));
  NAND3_X1   g20983(.A1(new_n20907_), .A2(new_n4034_), .A3(new_n20910_), .ZN(new_n21050_));
  NAND2_X1   g20984(.A1(new_n20911_), .A2(\a[11] ), .ZN(new_n21051_));
  NAND2_X1   g20985(.A1(new_n21051_), .A2(new_n21050_), .ZN(new_n21052_));
  NAND4_X1   g20986(.A1(new_n21047_), .A2(new_n21052_), .A3(new_n20924_), .A4(new_n20930_), .ZN(new_n21053_));
  AOI21_X1   g20987(.A1(new_n21049_), .A2(new_n21053_), .B(new_n20891_), .ZN(new_n21054_));
  OAI21_X1   g20988(.A1(new_n20925_), .A2(new_n20926_), .B(new_n20927_), .ZN(new_n21055_));
  NAND2_X1   g20989(.A1(new_n21055_), .A2(new_n20924_), .ZN(new_n21056_));
  NOR4_X1    g20990(.A1(new_n21043_), .A2(new_n21042_), .A3(new_n21044_), .A4(new_n20945_), .ZN(new_n21057_));
  NOR3_X1    g20991(.A1(new_n21012_), .A2(new_n21013_), .A3(new_n21011_), .ZN(new_n21058_));
  AOI21_X1   g20992(.A1(new_n21003_), .A2(new_n21009_), .B(new_n20954_), .ZN(new_n21059_));
  NOR3_X1    g20993(.A1(new_n21029_), .A2(new_n21030_), .A3(new_n21021_), .ZN(new_n21060_));
  AOI21_X1   g20994(.A1(new_n21023_), .A2(new_n21022_), .B(new_n21027_), .ZN(new_n21061_));
  NOR2_X1    g20995(.A1(new_n21033_), .A2(new_n21032_), .ZN(new_n21062_));
  XOR2_X1    g20996(.A1(new_n21036_), .A2(new_n4034_), .Z(new_n21063_));
  NAND2_X1   g20997(.A1(new_n21063_), .A2(new_n21062_), .ZN(new_n21064_));
  NOR3_X1    g20998(.A1(new_n21060_), .A2(new_n21061_), .A3(new_n21064_), .ZN(new_n21065_));
  NOR2_X1    g20999(.A1(new_n21065_), .A2(new_n21024_), .ZN(new_n21066_));
  OAI22_X1   g21000(.A1(new_n21059_), .A2(new_n21058_), .B1(new_n21066_), .B2(new_n21011_), .ZN(new_n21067_));
  AOI22_X1   g21001(.A1(new_n20932_), .A2(new_n20933_), .B1(new_n20944_), .B2(new_n20946_), .ZN(new_n21068_));
  NOR2_X1    g21002(.A1(new_n21057_), .A2(new_n21068_), .ZN(new_n21069_));
  AOI21_X1   g21003(.A1(new_n21067_), .A2(new_n21069_), .B(new_n21057_), .ZN(new_n21070_));
  NOR3_X1    g21004(.A1(new_n21070_), .A2(new_n20928_), .A3(new_n21056_), .ZN(new_n21071_));
  NOR2_X1    g21005(.A1(new_n21071_), .A2(new_n21052_), .ZN(new_n21072_));
  INV_X1     g21006(.I(new_n21053_), .ZN(new_n21073_));
  NOR3_X1    g21007(.A1(new_n21072_), .A2(new_n21073_), .A3(new_n20890_), .ZN(new_n21074_));
  NOR2_X1    g21008(.A1(new_n21074_), .A2(new_n21054_), .ZN(new_n21075_));
  NOR2_X1    g21009(.A1(new_n19478_), .A2(new_n19477_), .ZN(new_n21076_));
  NOR2_X1    g21010(.A1(new_n21076_), .A2(new_n19472_), .ZN(new_n21077_));
  NAND2_X1   g21011(.A1(new_n21076_), .A2(new_n19472_), .ZN(new_n21078_));
  NAND3_X1   g21012(.A1(new_n19470_), .A2(new_n19471_), .A3(new_n19466_), .ZN(new_n21079_));
  OAI21_X1   g21013(.A1(new_n19462_), .A2(new_n19455_), .B(new_n19437_), .ZN(new_n21080_));
  NAND2_X1   g21014(.A1(new_n21080_), .A2(new_n21079_), .ZN(new_n21081_));
  NAND2_X1   g21015(.A1(new_n21078_), .A2(new_n21081_), .ZN(new_n21082_));
  NOR3_X1    g21016(.A1(new_n21082_), .A2(new_n17780_), .A3(new_n21077_), .ZN(new_n21083_));
  INV_X1     g21017(.I(new_n21077_), .ZN(new_n21084_));
  INV_X1     g21018(.I(new_n21081_), .ZN(new_n21085_));
  AOI21_X1   g21019(.A1(new_n21076_), .A2(new_n19472_), .B(new_n21085_), .ZN(new_n21086_));
  AOI21_X1   g21020(.A1(new_n21084_), .A2(new_n21086_), .B(new_n19475_), .ZN(new_n21087_));
  NOR2_X1    g21021(.A1(new_n21083_), .A2(new_n21087_), .ZN(new_n21088_));
  OAI22_X1   g21022(.A1(new_n19463_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n19437_), .ZN(new_n21089_));
  NAND2_X1   g21023(.A1(new_n17780_), .A2(new_n6784_), .ZN(new_n21090_));
  AOI21_X1   g21024(.A1(new_n21089_), .A2(new_n21090_), .B(new_n6776_), .ZN(new_n21091_));
  AND3_X2    g21025(.A1(new_n21088_), .A2(new_n4009_), .A3(new_n21091_), .Z(new_n21092_));
  AOI21_X1   g21026(.A1(new_n21088_), .A2(new_n21091_), .B(new_n4009_), .ZN(new_n21093_));
  NOR2_X1    g21027(.A1(new_n21092_), .A2(new_n21093_), .ZN(new_n21094_));
  INV_X1     g21028(.I(new_n21094_), .ZN(new_n21095_));
  NAND2_X1   g21029(.A1(new_n19476_), .A2(new_n17784_), .ZN(new_n21096_));
  OAI21_X1   g21030(.A1(new_n19430_), .A2(new_n19431_), .B(new_n19438_), .ZN(new_n21097_));
  AOI21_X1   g21031(.A1(new_n21097_), .A2(new_n21096_), .B(new_n19437_), .ZN(new_n21098_));
  AOI21_X1   g21032(.A1(new_n19432_), .A2(new_n19447_), .B(new_n19466_), .ZN(new_n21099_));
  NOR2_X1    g21033(.A1(new_n21098_), .A2(new_n21099_), .ZN(new_n21100_));
  OAI22_X1   g21034(.A1(new_n17784_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n19428_), .ZN(new_n21101_));
  NAND2_X1   g21035(.A1(new_n19466_), .A2(new_n6784_), .ZN(new_n21102_));
  AOI21_X1   g21036(.A1(new_n21102_), .A2(new_n21101_), .B(new_n6776_), .ZN(new_n21103_));
  NAND2_X1   g21037(.A1(new_n21100_), .A2(new_n21103_), .ZN(new_n21104_));
  XOR2_X1    g21038(.A1(new_n21104_), .A2(\a[8] ), .Z(new_n21105_));
  NAND2_X1   g21039(.A1(new_n21067_), .A2(new_n21046_), .ZN(new_n21106_));
  NAND2_X1   g21040(.A1(new_n21041_), .A2(new_n21069_), .ZN(new_n21107_));
  NAND2_X1   g21041(.A1(new_n21107_), .A2(new_n21106_), .ZN(new_n21108_));
  NOR2_X1    g21042(.A1(new_n21108_), .A2(new_n21105_), .ZN(new_n21109_));
  NAND2_X1   g21043(.A1(new_n21070_), .A2(new_n20930_), .ZN(new_n21110_));
  NAND2_X1   g21044(.A1(new_n21047_), .A2(new_n21056_), .ZN(new_n21111_));
  OAI21_X1   g21045(.A1(new_n19478_), .A2(new_n19477_), .B(new_n21081_), .ZN(new_n21112_));
  NAND3_X1   g21046(.A1(new_n19470_), .A2(new_n19471_), .A3(new_n19437_), .ZN(new_n21113_));
  OAI21_X1   g21047(.A1(new_n19462_), .A2(new_n19455_), .B(new_n19466_), .ZN(new_n21114_));
  NAND2_X1   g21048(.A1(new_n21114_), .A2(new_n21113_), .ZN(new_n21115_));
  NAND3_X1   g21049(.A1(new_n19448_), .A2(new_n21115_), .A3(new_n19432_), .ZN(new_n21116_));
  NAND2_X1   g21050(.A1(new_n21112_), .A2(new_n21116_), .ZN(new_n21117_));
  OAI22_X1   g21051(.A1(new_n19437_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n17784_), .ZN(new_n21118_));
  NAND2_X1   g21052(.A1(new_n19472_), .A2(new_n6784_), .ZN(new_n21119_));
  AOI21_X1   g21053(.A1(new_n21119_), .A2(new_n21118_), .B(new_n6776_), .ZN(new_n21120_));
  NAND2_X1   g21054(.A1(new_n21117_), .A2(new_n21120_), .ZN(new_n21121_));
  XOR2_X1    g21055(.A1(new_n21121_), .A2(new_n4009_), .Z(new_n21122_));
  AOI21_X1   g21056(.A1(new_n21111_), .A2(new_n21110_), .B(new_n21122_), .ZN(new_n21123_));
  NOR2_X1    g21057(.A1(new_n21047_), .A2(new_n21056_), .ZN(new_n21124_));
  NOR2_X1    g21058(.A1(new_n21070_), .A2(new_n20930_), .ZN(new_n21125_));
  XOR2_X1    g21059(.A1(new_n21121_), .A2(\a[8] ), .Z(new_n21126_));
  NOR3_X1    g21060(.A1(new_n21124_), .A2(new_n21125_), .A3(new_n21126_), .ZN(new_n21127_));
  NOR3_X1    g21061(.A1(new_n21123_), .A2(new_n21127_), .A3(new_n21109_), .ZN(new_n21128_));
  NOR2_X1    g21062(.A1(new_n21128_), .A2(new_n21095_), .ZN(new_n21129_));
  XOR2_X1    g21063(.A1(new_n21104_), .A2(new_n4009_), .Z(new_n21130_));
  NAND3_X1   g21064(.A1(new_n21130_), .A2(new_n21106_), .A3(new_n21107_), .ZN(new_n21131_));
  OAI21_X1   g21065(.A1(new_n21124_), .A2(new_n21125_), .B(new_n21126_), .ZN(new_n21132_));
  NAND3_X1   g21066(.A1(new_n21111_), .A2(new_n21110_), .A3(new_n21122_), .ZN(new_n21133_));
  NAND3_X1   g21067(.A1(new_n21132_), .A2(new_n21133_), .A3(new_n21131_), .ZN(new_n21134_));
  NOR2_X1    g21068(.A1(new_n21134_), .A2(new_n21094_), .ZN(new_n21135_));
  OAI21_X1   g21069(.A1(new_n21129_), .A2(new_n21135_), .B(new_n21075_), .ZN(new_n21136_));
  OAI21_X1   g21070(.A1(new_n21072_), .A2(new_n21073_), .B(new_n20890_), .ZN(new_n21137_));
  NAND3_X1   g21071(.A1(new_n21049_), .A2(new_n20891_), .A3(new_n21053_), .ZN(new_n21138_));
  NAND2_X1   g21072(.A1(new_n21137_), .A2(new_n21138_), .ZN(new_n21139_));
  NAND2_X1   g21073(.A1(new_n21134_), .A2(new_n21094_), .ZN(new_n21140_));
  NAND2_X1   g21074(.A1(new_n21128_), .A2(new_n21095_), .ZN(new_n21141_));
  NAND3_X1   g21075(.A1(new_n21141_), .A2(new_n21140_), .A3(new_n21139_), .ZN(new_n21142_));
  NAND3_X1   g21076(.A1(new_n21136_), .A2(new_n21142_), .A3(new_n19527_), .ZN(new_n21143_));
  XOR2_X1    g21077(.A1(new_n19526_), .A2(\a[5] ), .Z(new_n21144_));
  AOI21_X1   g21078(.A1(new_n21141_), .A2(new_n21140_), .B(new_n21139_), .ZN(new_n21145_));
  NOR3_X1    g21079(.A1(new_n21129_), .A2(new_n21135_), .A3(new_n21075_), .ZN(new_n21146_));
  OAI21_X1   g21080(.A1(new_n21146_), .A2(new_n21145_), .B(new_n21144_), .ZN(new_n21147_));
  NOR3_X1    g21081(.A1(new_n21123_), .A2(new_n21127_), .A3(new_n21131_), .ZN(new_n21148_));
  AOI21_X1   g21082(.A1(new_n21132_), .A2(new_n21133_), .B(new_n21109_), .ZN(new_n21149_));
  NAND3_X1   g21083(.A1(new_n19469_), .A2(new_n17780_), .A3(new_n19473_), .ZN(new_n21150_));
  AOI21_X1   g21084(.A1(new_n17775_), .A2(new_n21150_), .B(new_n19474_), .ZN(new_n21151_));
  NOR3_X1    g21085(.A1(new_n19506_), .A2(new_n19505_), .A3(new_n19484_), .ZN(new_n21152_));
  AOI21_X1   g21086(.A1(new_n19496_), .A2(new_n19503_), .B(new_n17775_), .ZN(new_n21153_));
  OAI21_X1   g21087(.A1(new_n21152_), .A2(new_n21153_), .B(new_n21151_), .ZN(new_n21154_));
  OAI21_X1   g21088(.A1(new_n21151_), .A2(new_n19508_), .B(new_n21154_), .ZN(new_n21155_));
  OAI22_X1   g21089(.A1(new_n17775_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n19475_), .ZN(new_n21156_));
  NAND2_X1   g21090(.A1(new_n19496_), .A2(new_n19503_), .ZN(new_n21157_));
  NAND2_X1   g21091(.A1(new_n21157_), .A2(new_n6838_), .ZN(new_n21158_));
  AOI21_X1   g21092(.A1(new_n21158_), .A2(new_n21156_), .B(new_n6836_), .ZN(new_n21159_));
  AND3_X2    g21093(.A1(new_n21155_), .A2(new_n65_), .A3(new_n21159_), .Z(new_n21160_));
  AOI21_X1   g21094(.A1(new_n21155_), .A2(new_n21159_), .B(new_n65_), .ZN(new_n21161_));
  NOR4_X1    g21095(.A1(new_n21148_), .A2(new_n21149_), .A3(new_n21160_), .A4(new_n21161_), .ZN(new_n21162_));
  INV_X1     g21096(.I(new_n21162_), .ZN(new_n21163_));
  OAI22_X1   g21097(.A1(new_n21148_), .A2(new_n21149_), .B1(new_n21160_), .B2(new_n21161_), .ZN(new_n21164_));
  NAND2_X1   g21098(.A1(new_n21108_), .A2(new_n21105_), .ZN(new_n21165_));
  NAND3_X1   g21099(.A1(new_n21130_), .A2(new_n21106_), .A3(new_n21107_), .ZN(new_n21166_));
  NAND3_X1   g21100(.A1(new_n19469_), .A2(new_n19475_), .A3(new_n19473_), .ZN(new_n21167_));
  OAI21_X1   g21101(.A1(new_n19480_), .A2(new_n19481_), .B(new_n17780_), .ZN(new_n21168_));
  AOI21_X1   g21102(.A1(new_n21168_), .A2(new_n21167_), .B(new_n17775_), .ZN(new_n21169_));
  AOI21_X1   g21103(.A1(new_n19485_), .A2(new_n21150_), .B(new_n19484_), .ZN(new_n21170_));
  NOR2_X1    g21104(.A1(new_n21169_), .A2(new_n21170_), .ZN(new_n21171_));
  OAI22_X1   g21105(.A1(new_n19475_), .A2(new_n6843_), .B1(new_n19463_), .B2(new_n6913_), .ZN(new_n21172_));
  NAND2_X1   g21106(.A1(new_n19484_), .A2(new_n6838_), .ZN(new_n21173_));
  AOI21_X1   g21107(.A1(new_n21173_), .A2(new_n21172_), .B(new_n6836_), .ZN(new_n21174_));
  NAND3_X1   g21108(.A1(new_n21171_), .A2(new_n65_), .A3(new_n21174_), .ZN(new_n21175_));
  NOR3_X1    g21109(.A1(new_n19480_), .A2(new_n17780_), .A3(new_n19481_), .ZN(new_n21176_));
  AOI21_X1   g21110(.A1(new_n19469_), .A2(new_n19473_), .B(new_n19475_), .ZN(new_n21177_));
  OAI21_X1   g21111(.A1(new_n21176_), .A2(new_n21177_), .B(new_n19484_), .ZN(new_n21178_));
  OAI21_X1   g21112(.A1(new_n19482_), .A2(new_n19474_), .B(new_n17775_), .ZN(new_n21179_));
  NAND2_X1   g21113(.A1(new_n21178_), .A2(new_n21179_), .ZN(new_n21180_));
  INV_X1     g21114(.I(new_n21174_), .ZN(new_n21181_));
  OAI21_X1   g21115(.A1(new_n21180_), .A2(new_n21181_), .B(\a[5] ), .ZN(new_n21182_));
  NAND2_X1   g21116(.A1(new_n21182_), .A2(new_n21175_), .ZN(new_n21183_));
  AOI21_X1   g21117(.A1(new_n21165_), .A2(new_n21166_), .B(new_n21183_), .ZN(new_n21184_));
  INV_X1     g21118(.I(new_n21184_), .ZN(new_n21185_));
  NOR2_X1    g21119(.A1(new_n21085_), .A2(new_n21076_), .ZN(new_n21186_));
  NOR3_X1    g21120(.A1(new_n19462_), .A2(new_n19455_), .A3(new_n19466_), .ZN(new_n21187_));
  AOI21_X1   g21121(.A1(new_n19470_), .A2(new_n19471_), .B(new_n19437_), .ZN(new_n21188_));
  NOR2_X1    g21122(.A1(new_n21188_), .A2(new_n21187_), .ZN(new_n21189_));
  NOR3_X1    g21123(.A1(new_n21189_), .A2(new_n19477_), .A3(new_n19478_), .ZN(new_n21190_));
  AOI22_X1   g21124(.A1(new_n19466_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n19438_), .ZN(new_n21191_));
  AOI21_X1   g21125(.A1(new_n19472_), .A2(new_n6838_), .B(new_n21191_), .ZN(new_n21192_));
  NOR2_X1    g21126(.A1(new_n21192_), .A2(new_n6836_), .ZN(new_n21193_));
  OAI21_X1   g21127(.A1(new_n21186_), .A2(new_n21190_), .B(new_n21193_), .ZN(new_n21194_));
  NOR2_X1    g21128(.A1(new_n21194_), .A2(\a[5] ), .ZN(new_n21195_));
  AOI21_X1   g21129(.A1(new_n21117_), .A2(new_n21193_), .B(new_n65_), .ZN(new_n21196_));
  NOR2_X1    g21130(.A1(new_n21195_), .A2(new_n21196_), .ZN(new_n21197_));
  AOI21_X1   g21131(.A1(new_n21031_), .A2(new_n21028_), .B(new_n21038_), .ZN(new_n21198_));
  INV_X1     g21132(.I(new_n21198_), .ZN(new_n21199_));
  OAI22_X1   g21133(.A1(new_n19423_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n17787_), .ZN(new_n21200_));
  NAND2_X1   g21134(.A1(new_n20896_), .A2(new_n6784_), .ZN(new_n21201_));
  AOI21_X1   g21135(.A1(new_n21201_), .A2(new_n21200_), .B(new_n6776_), .ZN(new_n21202_));
  OAI21_X1   g21136(.A1(new_n20915_), .A2(new_n20918_), .B(new_n21202_), .ZN(new_n21203_));
  XOR2_X1    g21137(.A1(new_n21203_), .A2(new_n4009_), .Z(new_n21204_));
  NAND3_X1   g21138(.A1(new_n21199_), .A2(new_n21039_), .A3(new_n21204_), .ZN(new_n21205_));
  XOR2_X1    g21139(.A1(new_n21203_), .A2(\a[8] ), .Z(new_n21206_));
  OAI21_X1   g21140(.A1(new_n21065_), .A2(new_n21198_), .B(new_n21206_), .ZN(new_n21207_));
  XOR2_X1    g21141(.A1(new_n21037_), .A2(new_n21062_), .Z(new_n21208_));
  OAI22_X1   g21142(.A1(new_n17787_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n19412_), .ZN(new_n21209_));
  NAND2_X1   g21143(.A1(new_n19442_), .A2(new_n6784_), .ZN(new_n21210_));
  AOI21_X1   g21144(.A1(new_n21210_), .A2(new_n21209_), .B(new_n6776_), .ZN(new_n21211_));
  NAND3_X1   g21145(.A1(new_n20939_), .A2(new_n4009_), .A3(new_n21211_), .ZN(new_n21212_));
  AOI21_X1   g21146(.A1(new_n20939_), .A2(new_n21211_), .B(new_n4009_), .ZN(new_n21213_));
  INV_X1     g21147(.I(new_n21213_), .ZN(new_n21214_));
  AOI21_X1   g21148(.A1(new_n21214_), .A2(new_n21212_), .B(new_n21208_), .ZN(new_n21215_));
  NAND3_X1   g21149(.A1(new_n21205_), .A2(new_n21207_), .A3(new_n21215_), .ZN(new_n21216_));
  NOR3_X1    g21150(.A1(new_n21206_), .A2(new_n21065_), .A3(new_n21198_), .ZN(new_n21217_));
  AOI21_X1   g21151(.A1(new_n21199_), .A2(new_n21039_), .B(new_n21204_), .ZN(new_n21218_));
  INV_X1     g21152(.I(new_n21215_), .ZN(new_n21219_));
  OAI21_X1   g21153(.A1(new_n21218_), .A2(new_n21217_), .B(new_n21219_), .ZN(new_n21220_));
  NAND3_X1   g21154(.A1(new_n21197_), .A2(new_n21216_), .A3(new_n21220_), .ZN(new_n21221_));
  NAND3_X1   g21155(.A1(new_n21117_), .A2(new_n65_), .A3(new_n21193_), .ZN(new_n21222_));
  NAND2_X1   g21156(.A1(new_n21194_), .A2(\a[5] ), .ZN(new_n21223_));
  NAND2_X1   g21157(.A1(new_n21223_), .A2(new_n21222_), .ZN(new_n21224_));
  NOR3_X1    g21158(.A1(new_n21218_), .A2(new_n21217_), .A3(new_n21219_), .ZN(new_n21225_));
  AOI21_X1   g21159(.A1(new_n21205_), .A2(new_n21207_), .B(new_n21215_), .ZN(new_n21226_));
  OAI21_X1   g21160(.A1(new_n21225_), .A2(new_n21226_), .B(new_n21224_), .ZN(new_n21227_));
  NAND2_X1   g21161(.A1(new_n21227_), .A2(new_n21221_), .ZN(new_n21228_));
  XOR2_X1    g21162(.A1(new_n21063_), .A2(new_n21062_), .Z(new_n21229_));
  INV_X1     g21163(.I(new_n21212_), .ZN(new_n21230_));
  NOR3_X1    g21164(.A1(new_n21230_), .A2(new_n21229_), .A3(new_n21213_), .ZN(new_n21231_));
  AOI21_X1   g21165(.A1(new_n21214_), .A2(new_n21212_), .B(new_n21208_), .ZN(new_n21232_));
  NOR2_X1    g21166(.A1(new_n21232_), .A2(new_n21231_), .ZN(new_n21233_));
  AOI22_X1   g21167(.A1(new_n19438_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n20896_), .ZN(new_n21234_));
  NOR2_X1    g21168(.A1(new_n19437_), .A2(new_n6839_), .ZN(new_n21235_));
  OAI21_X1   g21169(.A1(new_n21234_), .A2(new_n21235_), .B(new_n6835_), .ZN(new_n21236_));
  NOR4_X1    g21170(.A1(new_n21098_), .A2(new_n21099_), .A3(\a[5] ), .A4(new_n21236_), .ZN(new_n21237_));
  NOR3_X1    g21171(.A1(new_n21098_), .A2(new_n21099_), .A3(new_n21236_), .ZN(new_n21238_));
  NOR2_X1    g21172(.A1(new_n21238_), .A2(new_n65_), .ZN(new_n21239_));
  NOR3_X1    g21173(.A1(new_n21239_), .A2(new_n21233_), .A3(new_n21237_), .ZN(new_n21240_));
  INV_X1     g21174(.I(new_n21240_), .ZN(new_n21241_));
  OAI21_X1   g21175(.A1(new_n21239_), .A2(new_n21237_), .B(new_n21233_), .ZN(new_n21242_));
  NAND2_X1   g21176(.A1(new_n21241_), .A2(new_n21242_), .ZN(new_n21243_));
  OAI22_X1   g21177(.A1(new_n19356_), .A2(new_n6089_), .B1(new_n6094_), .B2(new_n19364_), .ZN(new_n21244_));
  NAND2_X1   g21178(.A1(new_n17802_), .A2(new_n6090_), .ZN(new_n21245_));
  AOI21_X1   g21179(.A1(new_n21244_), .A2(new_n21245_), .B(new_n6082_), .ZN(new_n21246_));
  NAND3_X1   g21180(.A1(new_n19951_), .A2(new_n3521_), .A3(new_n21246_), .ZN(new_n21247_));
  AOI21_X1   g21181(.A1(new_n19951_), .A2(new_n21246_), .B(new_n3521_), .ZN(new_n21248_));
  INV_X1     g21182(.I(new_n21248_), .ZN(new_n21249_));
  NAND2_X1   g21183(.A1(new_n21249_), .A2(new_n21247_), .ZN(new_n21250_));
  NAND3_X1   g21184(.A1(new_n20571_), .A2(new_n20492_), .A3(new_n20498_), .ZN(new_n21251_));
  OAI21_X1   g21185(.A1(new_n20499_), .A2(new_n20497_), .B(new_n20570_), .ZN(new_n21252_));
  AOI21_X1   g21186(.A1(new_n21251_), .A2(new_n21252_), .B(new_n20487_), .ZN(new_n21253_));
  AOI21_X1   g21187(.A1(new_n20572_), .A2(new_n20501_), .B(new_n20565_), .ZN(new_n21254_));
  NOR2_X1    g21188(.A1(new_n21254_), .A2(new_n21253_), .ZN(new_n21255_));
  NOR3_X1    g21189(.A1(new_n20478_), .A2(new_n20563_), .A3(new_n20483_), .ZN(new_n21256_));
  AOI21_X1   g21190(.A1(new_n20482_), .A2(new_n20484_), .B(new_n20562_), .ZN(new_n21257_));
  OAI21_X1   g21191(.A1(new_n21256_), .A2(new_n21257_), .B(new_n20475_), .ZN(new_n21258_));
  OAI21_X1   g21192(.A1(new_n20559_), .A2(new_n20486_), .B(new_n20558_), .ZN(new_n21259_));
  NAND2_X1   g21193(.A1(new_n21258_), .A2(new_n21259_), .ZN(new_n21260_));
  OAI22_X1   g21194(.A1(new_n4297_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n4291_), .ZN(new_n21261_));
  NAND2_X1   g21195(.A1(new_n19350_), .A2(new_n4469_), .ZN(new_n21262_));
  AOI21_X1   g21196(.A1(new_n21261_), .A2(new_n21262_), .B(new_n4468_), .ZN(new_n21263_));
  OAI21_X1   g21197(.A1(new_n19822_), .A2(new_n19825_), .B(new_n21263_), .ZN(new_n21264_));
  XOR2_X1    g21198(.A1(new_n21264_), .A2(\a[17] ), .Z(new_n21265_));
  NAND2_X1   g21199(.A1(new_n21260_), .A2(new_n21265_), .ZN(new_n21266_));
  AOI22_X1   g21200(.A1(new_n19308_), .A2(new_n4292_), .B1(new_n4298_), .B2(new_n19545_), .ZN(new_n21267_));
  AOI21_X1   g21201(.A1(new_n4469_), .A2(new_n17850_), .B(new_n21267_), .ZN(new_n21268_));
  NOR2_X1    g21202(.A1(new_n21268_), .A2(new_n4468_), .ZN(new_n21269_));
  NAND2_X1   g21203(.A1(new_n19553_), .A2(new_n21269_), .ZN(new_n21270_));
  NOR2_X1    g21204(.A1(new_n21270_), .A2(\a[17] ), .ZN(new_n21271_));
  INV_X1     g21205(.I(new_n21271_), .ZN(new_n21272_));
  NAND2_X1   g21206(.A1(new_n21270_), .A2(\a[17] ), .ZN(new_n21273_));
  AOI21_X1   g21207(.A1(new_n21272_), .A2(new_n21273_), .B(new_n20455_), .ZN(new_n21274_));
  AOI22_X1   g21208(.A1(new_n19290_), .A2(new_n4292_), .B1(new_n4298_), .B2(new_n19308_), .ZN(new_n21275_));
  AOI21_X1   g21209(.A1(new_n4469_), .A2(new_n19545_), .B(new_n21275_), .ZN(new_n21276_));
  NAND2_X1   g21210(.A1(new_n19564_), .A2(new_n4295_), .ZN(new_n21277_));
  NOR2_X1    g21211(.A1(new_n21277_), .A2(new_n21276_), .ZN(new_n21278_));
  INV_X1     g21212(.I(new_n21278_), .ZN(new_n21279_));
  NOR2_X1    g21213(.A1(new_n4284_), .A2(new_n4294_), .ZN(new_n21280_));
  OAI21_X1   g21214(.A1(new_n19313_), .A2(new_n4297_), .B(new_n21280_), .ZN(new_n21281_));
  NOR2_X1    g21215(.A1(new_n19593_), .A2(new_n21281_), .ZN(new_n21282_));
  NOR2_X1    g21216(.A1(new_n19313_), .A2(new_n4284_), .ZN(new_n21283_));
  INV_X1     g21217(.I(new_n21283_), .ZN(new_n21284_));
  NAND4_X1   g21218(.A1(new_n21279_), .A2(\a[17] ), .A3(new_n21282_), .A4(new_n21284_), .ZN(new_n21285_));
  NAND3_X1   g21219(.A1(new_n21272_), .A2(new_n21273_), .A3(new_n20455_), .ZN(new_n21286_));
  AOI21_X1   g21220(.A1(new_n21285_), .A2(new_n21286_), .B(new_n21274_), .ZN(new_n21287_));
  NOR2_X1    g21221(.A1(new_n20454_), .A2(\a[20] ), .ZN(new_n21288_));
  NAND2_X1   g21222(.A1(new_n20452_), .A2(new_n20453_), .ZN(new_n21289_));
  NOR2_X1    g21223(.A1(new_n19593_), .A2(new_n21289_), .ZN(new_n21290_));
  NOR2_X1    g21224(.A1(new_n21290_), .A2(new_n3035_), .ZN(new_n21291_));
  NOR2_X1    g21225(.A1(new_n20455_), .A2(new_n3035_), .ZN(new_n21292_));
  NOR3_X1    g21226(.A1(new_n21288_), .A2(new_n21291_), .A3(new_n21292_), .ZN(new_n21293_));
  NOR3_X1    g21227(.A1(new_n21290_), .A2(new_n3035_), .A3(new_n20455_), .ZN(new_n21294_));
  NOR2_X1    g21228(.A1(new_n21293_), .A2(new_n21294_), .ZN(new_n21295_));
  AOI22_X1   g21229(.A1(new_n17850_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n19545_), .ZN(new_n21296_));
  AOI21_X1   g21230(.A1(new_n19305_), .A2(new_n4469_), .B(new_n21296_), .ZN(new_n21297_));
  NOR2_X1    g21231(.A1(new_n21297_), .A2(new_n4468_), .ZN(new_n21298_));
  NAND2_X1   g21232(.A1(new_n19607_), .A2(new_n21298_), .ZN(new_n21299_));
  NOR2_X1    g21233(.A1(new_n21299_), .A2(\a[17] ), .ZN(new_n21300_));
  NOR3_X1    g21234(.A1(new_n19618_), .A2(new_n4468_), .A3(new_n21297_), .ZN(new_n21301_));
  NOR2_X1    g21235(.A1(new_n21301_), .A2(new_n3372_), .ZN(new_n21302_));
  NOR3_X1    g21236(.A1(new_n21302_), .A2(new_n21300_), .A3(new_n21295_), .ZN(new_n21303_));
  OAI21_X1   g21237(.A1(new_n21302_), .A2(new_n21300_), .B(new_n21295_), .ZN(new_n21304_));
  OAI21_X1   g21238(.A1(new_n21287_), .A2(new_n21303_), .B(new_n21304_), .ZN(new_n21305_));
  OR3_X2     g21239(.A1(new_n19571_), .A2(new_n4095_), .A3(new_n20450_), .Z(new_n21306_));
  NAND2_X1   g21240(.A1(new_n21306_), .A2(new_n3035_), .ZN(new_n21307_));
  NAND2_X1   g21241(.A1(new_n20451_), .A2(\a[20] ), .ZN(new_n21308_));
  NOR3_X1    g21242(.A1(new_n20454_), .A2(new_n3035_), .A3(new_n20455_), .ZN(new_n21309_));
  INV_X1     g21243(.I(new_n21309_), .ZN(new_n21310_));
  NAND3_X1   g21244(.A1(new_n21307_), .A2(new_n21308_), .A3(new_n21310_), .ZN(new_n21311_));
  NOR2_X1    g21245(.A1(new_n20451_), .A2(\a[20] ), .ZN(new_n21312_));
  INV_X1     g21246(.I(new_n21308_), .ZN(new_n21313_));
  OAI21_X1   g21247(.A1(new_n21313_), .A2(new_n21312_), .B(new_n21309_), .ZN(new_n21314_));
  NAND2_X1   g21248(.A1(new_n21314_), .A2(new_n21311_), .ZN(new_n21315_));
  AOI22_X1   g21249(.A1(new_n19305_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n17850_), .ZN(new_n21316_));
  AOI21_X1   g21250(.A1(new_n4469_), .A2(new_n19321_), .B(new_n21316_), .ZN(new_n21317_));
  NOR2_X1    g21251(.A1(new_n21317_), .A2(new_n4468_), .ZN(new_n21318_));
  AND3_X2    g21252(.A1(new_n19647_), .A2(new_n3372_), .A3(new_n21318_), .Z(new_n21319_));
  AOI21_X1   g21253(.A1(new_n19647_), .A2(new_n21318_), .B(new_n3372_), .ZN(new_n21320_));
  NOR2_X1    g21254(.A1(new_n21319_), .A2(new_n21320_), .ZN(new_n21321_));
  NAND2_X1   g21255(.A1(new_n21321_), .A2(new_n21315_), .ZN(new_n21322_));
  NOR2_X1    g21256(.A1(new_n21321_), .A2(new_n21315_), .ZN(new_n21323_));
  AOI21_X1   g21257(.A1(new_n21305_), .A2(new_n21322_), .B(new_n21323_), .ZN(new_n21324_));
  NAND3_X1   g21258(.A1(new_n20446_), .A2(new_n20341_), .A3(new_n20444_), .ZN(new_n21325_));
  INV_X1     g21259(.I(new_n21325_), .ZN(new_n21326_));
  AOI21_X1   g21260(.A1(new_n20446_), .A2(new_n20444_), .B(new_n20341_), .ZN(new_n21327_));
  OAI21_X1   g21261(.A1(new_n21326_), .A2(new_n21327_), .B(new_n20456_), .ZN(new_n21328_));
  OAI21_X1   g21262(.A1(new_n20447_), .A2(new_n20546_), .B(new_n20457_), .ZN(new_n21329_));
  NAND2_X1   g21263(.A1(new_n21328_), .A2(new_n21329_), .ZN(new_n21330_));
  AOI22_X1   g21264(.A1(new_n19305_), .A2(new_n4292_), .B1(new_n4298_), .B2(new_n19321_), .ZN(new_n21331_));
  AOI21_X1   g21265(.A1(new_n4469_), .A2(new_n17827_), .B(new_n21331_), .ZN(new_n21332_));
  NOR2_X1    g21266(.A1(new_n21332_), .A2(new_n4468_), .ZN(new_n21333_));
  OAI21_X1   g21267(.A1(new_n19679_), .A2(new_n19682_), .B(new_n21333_), .ZN(new_n21334_));
  NOR2_X1    g21268(.A1(new_n21334_), .A2(\a[17] ), .ZN(new_n21335_));
  NAND2_X1   g21269(.A1(new_n21334_), .A2(\a[17] ), .ZN(new_n21336_));
  INV_X1     g21270(.I(new_n21336_), .ZN(new_n21337_));
  NOR3_X1    g21271(.A1(new_n21330_), .A2(new_n21337_), .A3(new_n21335_), .ZN(new_n21338_));
  OAI21_X1   g21272(.A1(new_n21337_), .A2(new_n21335_), .B(new_n21330_), .ZN(new_n21339_));
  OAI21_X1   g21273(.A1(new_n21324_), .A2(new_n21338_), .B(new_n21339_), .ZN(new_n21340_));
  NOR3_X1    g21274(.A1(new_n20472_), .A2(new_n20470_), .A3(new_n20553_), .ZN(new_n21341_));
  AOI21_X1   g21275(.A1(new_n20554_), .A2(new_n20555_), .B(new_n20465_), .ZN(new_n21342_));
  OAI21_X1   g21276(.A1(new_n21341_), .A2(new_n21342_), .B(new_n20547_), .ZN(new_n21343_));
  OAI21_X1   g21277(.A1(new_n20473_), .A2(new_n20557_), .B(new_n20459_), .ZN(new_n21344_));
  NAND2_X1   g21278(.A1(new_n21343_), .A2(new_n21344_), .ZN(new_n21345_));
  OAI22_X1   g21279(.A1(new_n17828_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19320_), .ZN(new_n21346_));
  NAND2_X1   g21280(.A1(new_n19349_), .A2(new_n4469_), .ZN(new_n21347_));
  AOI21_X1   g21281(.A1(new_n21347_), .A2(new_n21346_), .B(new_n4468_), .ZN(new_n21348_));
  NAND3_X1   g21282(.A1(new_n19760_), .A2(new_n3372_), .A3(new_n21348_), .ZN(new_n21349_));
  OAI21_X1   g21283(.A1(new_n19744_), .A2(new_n19747_), .B(new_n21348_), .ZN(new_n21350_));
  NAND2_X1   g21284(.A1(new_n21350_), .A2(\a[17] ), .ZN(new_n21351_));
  NAND3_X1   g21285(.A1(new_n21345_), .A2(new_n21349_), .A3(new_n21351_), .ZN(new_n21352_));
  NAND2_X1   g21286(.A1(new_n21340_), .A2(new_n21352_), .ZN(new_n21353_));
  NAND3_X1   g21287(.A1(new_n20554_), .A2(new_n20555_), .A3(new_n20465_), .ZN(new_n21354_));
  INV_X1     g21288(.I(new_n21342_), .ZN(new_n21355_));
  NAND2_X1   g21289(.A1(new_n21355_), .A2(new_n21354_), .ZN(new_n21356_));
  AOI21_X1   g21290(.A1(new_n20474_), .A2(new_n20556_), .B(new_n20547_), .ZN(new_n21357_));
  AOI21_X1   g21291(.A1(new_n21356_), .A2(new_n20547_), .B(new_n21357_), .ZN(new_n21358_));
  NAND2_X1   g21292(.A1(new_n21351_), .A2(new_n21349_), .ZN(new_n21359_));
  NAND2_X1   g21293(.A1(new_n21358_), .A2(new_n21359_), .ZN(new_n21360_));
  XOR2_X1    g21294(.A1(new_n21264_), .A2(new_n3372_), .Z(new_n21361_));
  NAND3_X1   g21295(.A1(new_n21361_), .A2(new_n21258_), .A3(new_n21259_), .ZN(new_n21362_));
  NAND4_X1   g21296(.A1(new_n21353_), .A2(new_n21266_), .A3(new_n21360_), .A4(new_n21362_), .ZN(new_n21363_));
  AOI22_X1   g21297(.A1(new_n19349_), .A2(new_n4292_), .B1(new_n4298_), .B2(new_n19350_), .ZN(new_n21364_));
  NOR2_X1    g21298(.A1(new_n17806_), .A2(new_n4470_), .ZN(new_n21365_));
  OAI21_X1   g21299(.A1(new_n21364_), .A2(new_n21365_), .B(new_n4295_), .ZN(new_n21366_));
  NOR2_X1    g21300(.A1(new_n19915_), .A2(new_n21366_), .ZN(new_n21367_));
  NAND2_X1   g21301(.A1(new_n21367_), .A2(new_n3372_), .ZN(new_n21368_));
  INV_X1     g21302(.I(new_n21366_), .ZN(new_n21369_));
  NAND2_X1   g21303(.A1(new_n19922_), .A2(new_n21369_), .ZN(new_n21370_));
  NAND2_X1   g21304(.A1(new_n21370_), .A2(\a[17] ), .ZN(new_n21371_));
  NAND2_X1   g21305(.A1(new_n21371_), .A2(new_n21368_), .ZN(new_n21372_));
  AOI21_X1   g21306(.A1(new_n21363_), .A2(new_n21266_), .B(new_n21372_), .ZN(new_n21373_));
  INV_X1     g21307(.I(new_n20455_), .ZN(new_n21374_));
  INV_X1     g21308(.I(new_n21273_), .ZN(new_n21375_));
  OAI21_X1   g21309(.A1(new_n21375_), .A2(new_n21271_), .B(new_n21374_), .ZN(new_n21376_));
  XOR2_X1    g21310(.A1(new_n21282_), .A2(\a[17] ), .Z(new_n21377_));
  NOR4_X1    g21311(.A1(new_n21377_), .A2(new_n3372_), .A3(new_n21278_), .A4(new_n21283_), .ZN(new_n21378_));
  NOR3_X1    g21312(.A1(new_n21375_), .A2(new_n21271_), .A3(new_n21374_), .ZN(new_n21379_));
  OAI21_X1   g21313(.A1(new_n21378_), .A2(new_n21379_), .B(new_n21376_), .ZN(new_n21380_));
  NAND2_X1   g21314(.A1(new_n21290_), .A2(new_n3035_), .ZN(new_n21381_));
  NAND2_X1   g21315(.A1(new_n20454_), .A2(\a[20] ), .ZN(new_n21382_));
  INV_X1     g21316(.I(new_n21292_), .ZN(new_n21383_));
  NAND3_X1   g21317(.A1(new_n21382_), .A2(new_n21381_), .A3(new_n21383_), .ZN(new_n21384_));
  INV_X1     g21318(.I(new_n21294_), .ZN(new_n21385_));
  NAND2_X1   g21319(.A1(new_n21384_), .A2(new_n21385_), .ZN(new_n21386_));
  NAND2_X1   g21320(.A1(new_n21301_), .A2(new_n3372_), .ZN(new_n21387_));
  NAND2_X1   g21321(.A1(new_n21299_), .A2(\a[17] ), .ZN(new_n21388_));
  NAND3_X1   g21322(.A1(new_n21387_), .A2(new_n21388_), .A3(new_n21386_), .ZN(new_n21389_));
  AOI21_X1   g21323(.A1(new_n21387_), .A2(new_n21388_), .B(new_n21386_), .ZN(new_n21390_));
  AOI21_X1   g21324(.A1(new_n21380_), .A2(new_n21389_), .B(new_n21390_), .ZN(new_n21391_));
  NOR3_X1    g21325(.A1(new_n21313_), .A2(new_n21312_), .A3(new_n21309_), .ZN(new_n21392_));
  AOI21_X1   g21326(.A1(new_n21307_), .A2(new_n21308_), .B(new_n21310_), .ZN(new_n21393_));
  NOR2_X1    g21327(.A1(new_n21392_), .A2(new_n21393_), .ZN(new_n21394_));
  NOR3_X1    g21328(.A1(new_n21394_), .A2(new_n21319_), .A3(new_n21320_), .ZN(new_n21395_));
  OAI21_X1   g21329(.A1(new_n21319_), .A2(new_n21320_), .B(new_n21394_), .ZN(new_n21396_));
  OAI21_X1   g21330(.A1(new_n21391_), .A2(new_n21395_), .B(new_n21396_), .ZN(new_n21397_));
  OAI21_X1   g21331(.A1(new_n20544_), .A2(new_n20445_), .B(new_n20340_), .ZN(new_n21398_));
  AOI21_X1   g21332(.A1(new_n21398_), .A2(new_n21325_), .B(new_n20457_), .ZN(new_n21399_));
  AOI21_X1   g21333(.A1(new_n20458_), .A2(new_n20545_), .B(new_n20456_), .ZN(new_n21400_));
  NOR2_X1    g21334(.A1(new_n21399_), .A2(new_n21400_), .ZN(new_n21401_));
  INV_X1     g21335(.I(new_n21335_), .ZN(new_n21402_));
  NAND3_X1   g21336(.A1(new_n21402_), .A2(new_n21401_), .A3(new_n21336_), .ZN(new_n21403_));
  AOI21_X1   g21337(.A1(new_n21402_), .A2(new_n21336_), .B(new_n21401_), .ZN(new_n21404_));
  AOI21_X1   g21338(.A1(new_n21397_), .A2(new_n21403_), .B(new_n21404_), .ZN(new_n21405_));
  NOR2_X1    g21339(.A1(new_n21358_), .A2(new_n21359_), .ZN(new_n21406_));
  OAI21_X1   g21340(.A1(new_n21405_), .A2(new_n21406_), .B(new_n21360_), .ZN(new_n21407_));
  NOR2_X1    g21341(.A1(new_n21260_), .A2(new_n21265_), .ZN(new_n21408_));
  OAI21_X1   g21342(.A1(new_n21407_), .A2(new_n21408_), .B(new_n21266_), .ZN(new_n21409_));
  NOR2_X1    g21343(.A1(new_n21370_), .A2(\a[17] ), .ZN(new_n21410_));
  NOR2_X1    g21344(.A1(new_n21367_), .A2(new_n3372_), .ZN(new_n21411_));
  NOR2_X1    g21345(.A1(new_n21410_), .A2(new_n21411_), .ZN(new_n21412_));
  NOR2_X1    g21346(.A1(new_n21409_), .A2(new_n21412_), .ZN(new_n21413_));
  OAI21_X1   g21347(.A1(new_n21373_), .A2(new_n21413_), .B(new_n21255_), .ZN(new_n21414_));
  INV_X1     g21348(.I(new_n21255_), .ZN(new_n21415_));
  NAND2_X1   g21349(.A1(new_n21409_), .A2(new_n21412_), .ZN(new_n21416_));
  NAND3_X1   g21350(.A1(new_n21363_), .A2(new_n21372_), .A3(new_n21266_), .ZN(new_n21417_));
  NAND3_X1   g21351(.A1(new_n21417_), .A2(new_n21416_), .A3(new_n21415_), .ZN(new_n21418_));
  NAND3_X1   g21352(.A1(new_n21414_), .A2(new_n21418_), .A3(new_n21250_), .ZN(new_n21419_));
  INV_X1     g21353(.I(new_n21247_), .ZN(new_n21420_));
  NOR2_X1    g21354(.A1(new_n21420_), .A2(new_n21248_), .ZN(new_n21421_));
  AOI21_X1   g21355(.A1(new_n21417_), .A2(new_n21416_), .B(new_n21415_), .ZN(new_n21422_));
  NOR3_X1    g21356(.A1(new_n21373_), .A2(new_n21413_), .A3(new_n21255_), .ZN(new_n21423_));
  OAI21_X1   g21357(.A1(new_n21422_), .A2(new_n21423_), .B(new_n21421_), .ZN(new_n21424_));
  AOI21_X1   g21358(.A1(new_n21258_), .A2(new_n21259_), .B(new_n21361_), .ZN(new_n21425_));
  NOR3_X1    g21359(.A1(new_n21407_), .A2(new_n21408_), .A3(new_n21425_), .ZN(new_n21426_));
  AOI22_X1   g21360(.A1(new_n21353_), .A2(new_n21360_), .B1(new_n21266_), .B2(new_n21362_), .ZN(new_n21427_));
  NOR2_X1    g21361(.A1(new_n21427_), .A2(new_n21426_), .ZN(new_n21428_));
  OAI22_X1   g21362(.A1(new_n19356_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n17806_), .ZN(new_n21429_));
  NAND2_X1   g21363(.A1(new_n19365_), .A2(new_n6090_), .ZN(new_n21430_));
  AOI21_X1   g21364(.A1(new_n21429_), .A2(new_n21430_), .B(new_n6082_), .ZN(new_n21431_));
  NAND3_X1   g21365(.A1(new_n19538_), .A2(new_n3521_), .A3(new_n21431_), .ZN(new_n21432_));
  INV_X1     g21366(.I(new_n21432_), .ZN(new_n21433_));
  AOI21_X1   g21367(.A1(new_n19538_), .A2(new_n21431_), .B(new_n3521_), .ZN(new_n21434_));
  NOR2_X1    g21368(.A1(new_n21433_), .A2(new_n21434_), .ZN(new_n21435_));
  NAND2_X1   g21369(.A1(new_n21428_), .A2(new_n21435_), .ZN(new_n21436_));
  OAI22_X1   g21370(.A1(new_n17806_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n19346_), .ZN(new_n21437_));
  NAND2_X1   g21371(.A1(new_n19359_), .A2(new_n6090_), .ZN(new_n21438_));
  AOI21_X1   g21372(.A1(new_n21438_), .A2(new_n21437_), .B(new_n6082_), .ZN(new_n21439_));
  NAND2_X1   g21373(.A1(new_n20096_), .A2(new_n21439_), .ZN(new_n21440_));
  XOR2_X1    g21374(.A1(new_n21440_), .A2(\a[14] ), .Z(new_n21441_));
  NOR2_X1    g21375(.A1(new_n21345_), .A2(new_n21359_), .ZN(new_n21442_));
  AOI21_X1   g21376(.A1(new_n21349_), .A2(new_n21351_), .B(new_n21358_), .ZN(new_n21443_));
  OAI21_X1   g21377(.A1(new_n21443_), .A2(new_n21442_), .B(new_n21340_), .ZN(new_n21444_));
  NAND2_X1   g21378(.A1(new_n21360_), .A2(new_n21352_), .ZN(new_n21445_));
  NAND2_X1   g21379(.A1(new_n21445_), .A2(new_n21405_), .ZN(new_n21446_));
  NAND2_X1   g21380(.A1(new_n21446_), .A2(new_n21444_), .ZN(new_n21447_));
  NAND2_X1   g21381(.A1(new_n21441_), .A2(new_n21447_), .ZN(new_n21448_));
  INV_X1     g21382(.I(new_n21434_), .ZN(new_n21449_));
  NAND2_X1   g21383(.A1(new_n21449_), .A2(new_n21432_), .ZN(new_n21450_));
  OAI21_X1   g21384(.A1(new_n21426_), .A2(new_n21427_), .B(new_n21450_), .ZN(new_n21451_));
  NAND3_X1   g21385(.A1(new_n21436_), .A2(new_n21451_), .A3(new_n21448_), .ZN(new_n21452_));
  AOI22_X1   g21386(.A1(new_n21424_), .A2(new_n21419_), .B1(new_n21452_), .B2(new_n21250_), .ZN(new_n21453_));
  INV_X1     g21387(.I(new_n20051_), .ZN(new_n21454_));
  AOI22_X1   g21388(.A1(new_n17802_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n19365_), .ZN(new_n21455_));
  NOR2_X1    g21389(.A1(new_n17797_), .A2(new_n6091_), .ZN(new_n21456_));
  OAI21_X1   g21390(.A1(new_n21456_), .A2(new_n21455_), .B(new_n6081_), .ZN(new_n21457_));
  NOR3_X1    g21391(.A1(new_n21454_), .A2(\a[14] ), .A3(new_n21457_), .ZN(new_n21458_));
  INV_X1     g21392(.I(new_n21457_), .ZN(new_n21459_));
  AOI21_X1   g21393(.A1(new_n20051_), .A2(new_n21459_), .B(new_n3521_), .ZN(new_n21460_));
  NOR2_X1    g21394(.A1(new_n21458_), .A2(new_n21460_), .ZN(new_n21461_));
  INV_X1     g21395(.I(new_n21461_), .ZN(new_n21462_));
  NAND2_X1   g21396(.A1(new_n21453_), .A2(new_n21462_), .ZN(new_n21463_));
  XOR2_X1    g21397(.A1(new_n20781_), .A2(new_n20526_), .Z(new_n21464_));
  INV_X1     g21398(.I(new_n21464_), .ZN(new_n21465_));
  OAI21_X1   g21399(.A1(new_n21453_), .A2(new_n21462_), .B(new_n21465_), .ZN(new_n21466_));
  NOR2_X1    g21400(.A1(new_n20781_), .A2(new_n20782_), .ZN(new_n21467_));
  INV_X1     g21401(.I(new_n21467_), .ZN(new_n21468_));
  NOR3_X1    g21402(.A1(new_n21468_), .A2(new_n20595_), .A3(new_n20599_), .ZN(new_n21469_));
  AOI21_X1   g21403(.A1(new_n20785_), .A2(new_n20784_), .B(new_n21467_), .ZN(new_n21470_));
  OAI22_X1   g21404(.A1(new_n17797_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n17801_), .ZN(new_n21471_));
  OAI21_X1   g21405(.A1(new_n19375_), .A2(new_n6091_), .B(new_n21471_), .ZN(new_n21472_));
  NAND4_X1   g21406(.A1(new_n20709_), .A2(new_n20708_), .A3(new_n6081_), .A4(new_n21472_), .ZN(new_n21473_));
  XOR2_X1    g21407(.A1(new_n21473_), .A2(\a[14] ), .Z(new_n21474_));
  OAI21_X1   g21408(.A1(new_n21469_), .A2(new_n21470_), .B(new_n21474_), .ZN(new_n21475_));
  NOR3_X1    g21409(.A1(new_n21474_), .A2(new_n21469_), .A3(new_n21470_), .ZN(new_n21476_));
  INV_X1     g21410(.I(new_n21476_), .ZN(new_n21477_));
  AOI22_X1   g21411(.A1(new_n21466_), .A2(new_n21463_), .B1(new_n21477_), .B2(new_n21475_), .ZN(new_n21478_));
  NOR3_X1    g21412(.A1(new_n21422_), .A2(new_n21423_), .A3(new_n21421_), .ZN(new_n21479_));
  AOI21_X1   g21413(.A1(new_n21414_), .A2(new_n21418_), .B(new_n21250_), .ZN(new_n21480_));
  NOR3_X1    g21414(.A1(new_n21450_), .A2(new_n21426_), .A3(new_n21427_), .ZN(new_n21481_));
  XOR2_X1    g21415(.A1(new_n21440_), .A2(new_n3521_), .Z(new_n21482_));
  INV_X1     g21416(.I(new_n21447_), .ZN(new_n21483_));
  NOR2_X1    g21417(.A1(new_n21483_), .A2(new_n21482_), .ZN(new_n21484_));
  NOR2_X1    g21418(.A1(new_n21428_), .A2(new_n21435_), .ZN(new_n21485_));
  NOR3_X1    g21419(.A1(new_n21485_), .A2(new_n21484_), .A3(new_n21481_), .ZN(new_n21486_));
  OAI22_X1   g21420(.A1(new_n21479_), .A2(new_n21480_), .B1(new_n21486_), .B2(new_n21421_), .ZN(new_n21487_));
  NOR2_X1    g21421(.A1(new_n21487_), .A2(new_n21461_), .ZN(new_n21488_));
  AOI21_X1   g21422(.A1(new_n21487_), .A2(new_n21461_), .B(new_n21464_), .ZN(new_n21489_));
  XOR2_X1    g21423(.A1(new_n21473_), .A2(new_n3521_), .Z(new_n21490_));
  NOR3_X1    g21424(.A1(new_n21490_), .A2(new_n21469_), .A3(new_n21470_), .ZN(new_n21491_));
  INV_X1     g21425(.I(new_n21469_), .ZN(new_n21492_));
  INV_X1     g21426(.I(new_n21470_), .ZN(new_n21493_));
  AOI21_X1   g21427(.A1(new_n21492_), .A2(new_n21493_), .B(new_n21474_), .ZN(new_n21494_));
  NOR2_X1    g21428(.A1(new_n21494_), .A2(new_n21491_), .ZN(new_n21495_));
  NOR3_X1    g21429(.A1(new_n21495_), .A2(new_n21489_), .A3(new_n21488_), .ZN(new_n21496_));
  AOI22_X1   g21430(.A1(new_n19386_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n17794_), .ZN(new_n21497_));
  NOR2_X1    g21431(.A1(new_n19393_), .A2(new_n4710_), .ZN(new_n21498_));
  OAI21_X1   g21432(.A1(new_n21497_), .A2(new_n21498_), .B(new_n4706_), .ZN(new_n21499_));
  NOR3_X1    g21433(.A1(new_n20291_), .A2(\a[11] ), .A3(new_n21499_), .ZN(new_n21500_));
  NOR2_X1    g21434(.A1(new_n20291_), .A2(new_n21499_), .ZN(new_n21501_));
  NOR2_X1    g21435(.A1(new_n21501_), .A2(new_n4034_), .ZN(new_n21502_));
  NOR2_X1    g21436(.A1(new_n21502_), .A2(new_n21500_), .ZN(new_n21503_));
  INV_X1     g21437(.I(new_n21503_), .ZN(new_n21504_));
  NOR3_X1    g21438(.A1(new_n21504_), .A2(new_n21496_), .A3(new_n21478_), .ZN(new_n21505_));
  INV_X1     g21439(.I(new_n21478_), .ZN(new_n21506_));
  INV_X1     g21440(.I(new_n21496_), .ZN(new_n21507_));
  AOI21_X1   g21441(.A1(new_n21507_), .A2(new_n21506_), .B(new_n21503_), .ZN(new_n21508_));
  OAI22_X1   g21442(.A1(new_n17789_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n19400_), .ZN(new_n21509_));
  NAND2_X1   g21443(.A1(new_n19407_), .A2(new_n6784_), .ZN(new_n21510_));
  AOI21_X1   g21444(.A1(new_n21510_), .A2(new_n21509_), .B(new_n6776_), .ZN(new_n21511_));
  NAND3_X1   g21445(.A1(new_n20860_), .A2(new_n20862_), .A3(new_n21511_), .ZN(new_n21512_));
  NOR2_X1    g21446(.A1(new_n21512_), .A2(\a[8] ), .ZN(new_n21513_));
  NAND2_X1   g21447(.A1(new_n21512_), .A2(\a[8] ), .ZN(new_n21514_));
  INV_X1     g21448(.I(new_n21514_), .ZN(new_n21515_));
  NOR2_X1    g21449(.A1(new_n21515_), .A2(new_n21513_), .ZN(new_n21516_));
  OR3_X2     g21450(.A1(new_n21516_), .A2(new_n21505_), .A3(new_n21508_), .Z(new_n21517_));
  AOI21_X1   g21451(.A1(new_n21492_), .A2(new_n21493_), .B(new_n21490_), .ZN(new_n21518_));
  AOI21_X1   g21452(.A1(new_n21466_), .A2(new_n21463_), .B(new_n21518_), .ZN(new_n21519_));
  NOR2_X1    g21453(.A1(new_n21519_), .A2(new_n21476_), .ZN(new_n21520_));
  AOI21_X1   g21454(.A1(new_n20600_), .A2(new_n20784_), .B(new_n20322_), .ZN(new_n21521_));
  NAND4_X1   g21455(.A1(new_n20785_), .A2(new_n20784_), .A3(new_n20783_), .A4(new_n20322_), .ZN(new_n21522_));
  INV_X1     g21456(.I(new_n21522_), .ZN(new_n21523_));
  OAI21_X1   g21457(.A1(new_n21521_), .A2(new_n21523_), .B(new_n20434_), .ZN(new_n21524_));
  NAND3_X1   g21458(.A1(new_n20785_), .A2(new_n20784_), .A3(new_n20783_), .ZN(new_n21525_));
  NAND2_X1   g21459(.A1(new_n21525_), .A2(new_n20779_), .ZN(new_n21526_));
  NAND3_X1   g21460(.A1(new_n21526_), .A2(new_n20610_), .A3(new_n21522_), .ZN(new_n21527_));
  OAI22_X1   g21461(.A1(new_n19375_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n17797_), .ZN(new_n21528_));
  NAND2_X1   g21462(.A1(new_n19386_), .A2(new_n6090_), .ZN(new_n21529_));
  AOI21_X1   g21463(.A1(new_n21529_), .A2(new_n21528_), .B(new_n6082_), .ZN(new_n21530_));
  NAND3_X1   g21464(.A1(new_n20162_), .A2(new_n3521_), .A3(new_n21530_), .ZN(new_n21531_));
  AOI21_X1   g21465(.A1(new_n20162_), .A2(new_n21530_), .B(new_n3521_), .ZN(new_n21532_));
  INV_X1     g21466(.I(new_n21532_), .ZN(new_n21533_));
  NAND2_X1   g21467(.A1(new_n21533_), .A2(new_n21531_), .ZN(new_n21534_));
  NAND3_X1   g21468(.A1(new_n21524_), .A2(new_n21527_), .A3(new_n21534_), .ZN(new_n21535_));
  AOI21_X1   g21469(.A1(new_n21526_), .A2(new_n21522_), .B(new_n20610_), .ZN(new_n21536_));
  NOR3_X1    g21470(.A1(new_n21521_), .A2(new_n21523_), .A3(new_n20434_), .ZN(new_n21537_));
  INV_X1     g21471(.I(new_n21531_), .ZN(new_n21538_));
  NOR2_X1    g21472(.A1(new_n21538_), .A2(new_n21532_), .ZN(new_n21539_));
  OAI21_X1   g21473(.A1(new_n21537_), .A2(new_n21536_), .B(new_n21539_), .ZN(new_n21540_));
  OAI22_X1   g21474(.A1(new_n19393_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n17793_), .ZN(new_n21541_));
  NAND2_X1   g21475(.A1(new_n19399_), .A2(new_n4709_), .ZN(new_n21542_));
  AOI21_X1   g21476(.A1(new_n21542_), .A2(new_n21541_), .B(new_n4707_), .ZN(new_n21543_));
  NAND3_X1   g21477(.A1(new_n20264_), .A2(new_n4034_), .A3(new_n21543_), .ZN(new_n21544_));
  INV_X1     g21478(.I(new_n20262_), .ZN(new_n21545_));
  NOR3_X1    g21479(.A1(new_n19395_), .A2(new_n19390_), .A3(new_n20263_), .ZN(new_n21546_));
  OAI21_X1   g21480(.A1(new_n21545_), .A2(new_n21546_), .B(new_n21543_), .ZN(new_n21547_));
  NAND2_X1   g21481(.A1(new_n21547_), .A2(\a[11] ), .ZN(new_n21548_));
  AND2_X2    g21482(.A1(new_n21548_), .A2(new_n21544_), .Z(new_n21549_));
  NAND3_X1   g21483(.A1(new_n21549_), .A2(new_n21540_), .A3(new_n21535_), .ZN(new_n21550_));
  NOR3_X1    g21484(.A1(new_n21537_), .A2(new_n21536_), .A3(new_n21539_), .ZN(new_n21551_));
  AOI21_X1   g21485(.A1(new_n21524_), .A2(new_n21527_), .B(new_n21534_), .ZN(new_n21552_));
  NAND2_X1   g21486(.A1(new_n21548_), .A2(new_n21544_), .ZN(new_n21553_));
  OAI21_X1   g21487(.A1(new_n21551_), .A2(new_n21552_), .B(new_n21553_), .ZN(new_n21554_));
  AOI21_X1   g21488(.A1(new_n21550_), .A2(new_n21554_), .B(new_n21520_), .ZN(new_n21555_));
  OAI21_X1   g21489(.A1(new_n21489_), .A2(new_n21488_), .B(new_n21475_), .ZN(new_n21556_));
  NAND2_X1   g21490(.A1(new_n21556_), .A2(new_n21477_), .ZN(new_n21557_));
  NAND3_X1   g21491(.A1(new_n21540_), .A2(new_n21535_), .A3(new_n21553_), .ZN(new_n21558_));
  OAI21_X1   g21492(.A1(new_n21551_), .A2(new_n21552_), .B(new_n21549_), .ZN(new_n21559_));
  AOI21_X1   g21493(.A1(new_n21559_), .A2(new_n21558_), .B(new_n21557_), .ZN(new_n21560_));
  OAI22_X1   g21494(.A1(new_n19410_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n17789_), .ZN(new_n21561_));
  NAND2_X1   g21495(.A1(new_n19415_), .A2(new_n6784_), .ZN(new_n21562_));
  AOI21_X1   g21496(.A1(new_n21562_), .A2(new_n21561_), .B(new_n6776_), .ZN(new_n21563_));
  NAND3_X1   g21497(.A1(new_n20846_), .A2(new_n4009_), .A3(new_n21563_), .ZN(new_n21564_));
  INV_X1     g21498(.I(new_n20844_), .ZN(new_n21565_));
  NOR3_X1    g21499(.A1(new_n19408_), .A2(new_n19404_), .A3(new_n20845_), .ZN(new_n21566_));
  OAI21_X1   g21500(.A1(new_n21565_), .A2(new_n21566_), .B(new_n21563_), .ZN(new_n21567_));
  NAND2_X1   g21501(.A1(new_n21567_), .A2(\a[8] ), .ZN(new_n21568_));
  NAND2_X1   g21502(.A1(new_n21568_), .A2(new_n21564_), .ZN(new_n21569_));
  NOR3_X1    g21503(.A1(new_n21569_), .A2(new_n21560_), .A3(new_n21555_), .ZN(new_n21570_));
  NOR3_X1    g21504(.A1(new_n21551_), .A2(new_n21552_), .A3(new_n21553_), .ZN(new_n21571_));
  AOI21_X1   g21505(.A1(new_n21535_), .A2(new_n21540_), .B(new_n21549_), .ZN(new_n21572_));
  OAI21_X1   g21506(.A1(new_n21572_), .A2(new_n21571_), .B(new_n21557_), .ZN(new_n21573_));
  NOR3_X1    g21507(.A1(new_n21549_), .A2(new_n21552_), .A3(new_n21551_), .ZN(new_n21574_));
  AOI21_X1   g21508(.A1(new_n21540_), .A2(new_n21535_), .B(new_n21553_), .ZN(new_n21575_));
  OAI21_X1   g21509(.A1(new_n21574_), .A2(new_n21575_), .B(new_n21520_), .ZN(new_n21576_));
  AOI22_X1   g21510(.A1(new_n21573_), .A2(new_n21576_), .B1(new_n21564_), .B2(new_n21568_), .ZN(new_n21577_));
  OAI21_X1   g21511(.A1(new_n21577_), .A2(new_n21570_), .B(new_n21508_), .ZN(new_n21578_));
  OAI21_X1   g21512(.A1(new_n21496_), .A2(new_n21478_), .B(new_n21504_), .ZN(new_n21579_));
  NOR2_X1    g21513(.A1(new_n21567_), .A2(\a[8] ), .ZN(new_n21580_));
  AOI21_X1   g21514(.A1(new_n20846_), .A2(new_n21563_), .B(new_n4009_), .ZN(new_n21581_));
  NOR2_X1    g21515(.A1(new_n21580_), .A2(new_n21581_), .ZN(new_n21582_));
  NOR3_X1    g21516(.A1(new_n21582_), .A2(new_n21560_), .A3(new_n21555_), .ZN(new_n21583_));
  AOI21_X1   g21517(.A1(new_n21573_), .A2(new_n21576_), .B(new_n21569_), .ZN(new_n21584_));
  OAI21_X1   g21518(.A1(new_n21584_), .A2(new_n21583_), .B(new_n21579_), .ZN(new_n21585_));
  NAND3_X1   g21519(.A1(new_n21585_), .A2(new_n21578_), .A3(new_n21517_), .ZN(new_n21586_));
  NOR3_X1    g21520(.A1(new_n21516_), .A2(new_n21505_), .A3(new_n21508_), .ZN(new_n21587_));
  NAND3_X1   g21521(.A1(new_n21582_), .A2(new_n21573_), .A3(new_n21576_), .ZN(new_n21588_));
  OAI21_X1   g21522(.A1(new_n21555_), .A2(new_n21560_), .B(new_n21569_), .ZN(new_n21589_));
  AOI21_X1   g21523(.A1(new_n21589_), .A2(new_n21588_), .B(new_n21579_), .ZN(new_n21590_));
  NAND3_X1   g21524(.A1(new_n21569_), .A2(new_n21573_), .A3(new_n21576_), .ZN(new_n21591_));
  OAI21_X1   g21525(.A1(new_n21555_), .A2(new_n21560_), .B(new_n21582_), .ZN(new_n21592_));
  AOI21_X1   g21526(.A1(new_n21592_), .A2(new_n21591_), .B(new_n21508_), .ZN(new_n21593_));
  OAI21_X1   g21527(.A1(new_n21593_), .A2(new_n21590_), .B(new_n21587_), .ZN(new_n21594_));
  NAND3_X1   g21528(.A1(new_n21507_), .A2(new_n21506_), .A3(new_n21503_), .ZN(new_n21595_));
  INV_X1     g21529(.I(new_n21513_), .ZN(new_n21596_));
  NAND4_X1   g21530(.A1(new_n21595_), .A2(new_n21579_), .A3(new_n21596_), .A4(new_n21514_), .ZN(new_n21597_));
  OAI22_X1   g21531(.A1(new_n21508_), .A2(new_n21505_), .B1(new_n21515_), .B2(new_n21513_), .ZN(new_n21598_));
  NAND2_X1   g21532(.A1(new_n21598_), .A2(new_n21597_), .ZN(new_n21599_));
  AOI22_X1   g21533(.A1(new_n19439_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n19415_), .ZN(new_n21600_));
  NOR2_X1    g21534(.A1(new_n19423_), .A2(new_n6839_), .ZN(new_n21601_));
  OAI21_X1   g21535(.A1(new_n21601_), .A2(new_n21600_), .B(new_n6835_), .ZN(new_n21602_));
  NOR4_X1    g21536(.A1(new_n20936_), .A2(new_n20938_), .A3(\a[5] ), .A4(new_n21602_), .ZN(new_n21603_));
  INV_X1     g21537(.I(new_n21602_), .ZN(new_n21604_));
  AOI21_X1   g21538(.A1(new_n20939_), .A2(new_n21604_), .B(new_n65_), .ZN(new_n21605_));
  OAI21_X1   g21539(.A1(new_n21605_), .A2(new_n21603_), .B(new_n21599_), .ZN(new_n21606_));
  OAI22_X1   g21540(.A1(new_n19423_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n17787_), .ZN(new_n21607_));
  NAND2_X1   g21541(.A1(new_n20896_), .A2(new_n6838_), .ZN(new_n21608_));
  AOI21_X1   g21542(.A1(new_n21608_), .A2(new_n21607_), .B(new_n6836_), .ZN(new_n21609_));
  OAI21_X1   g21543(.A1(new_n20915_), .A2(new_n20918_), .B(new_n21609_), .ZN(new_n21610_));
  XOR2_X1    g21544(.A1(new_n21610_), .A2(\a[5] ), .Z(new_n21611_));
  AOI22_X1   g21545(.A1(new_n21586_), .A2(new_n21594_), .B1(new_n21611_), .B2(new_n21606_), .ZN(new_n21612_));
  NOR2_X1    g21546(.A1(new_n21611_), .A2(new_n21606_), .ZN(new_n21613_));
  AOI22_X1   g21547(.A1(new_n20896_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n19442_), .ZN(new_n21614_));
  INV_X1     g21548(.I(new_n21614_), .ZN(new_n21615_));
  NAND2_X1   g21549(.A1(new_n19438_), .A2(new_n6838_), .ZN(new_n21616_));
  AOI21_X1   g21550(.A1(new_n21615_), .A2(new_n21616_), .B(new_n6836_), .ZN(new_n21617_));
  NAND3_X1   g21551(.A1(new_n20907_), .A2(new_n65_), .A3(new_n21617_), .ZN(new_n21618_));
  NAND2_X1   g21552(.A1(new_n20905_), .A2(new_n17784_), .ZN(new_n21619_));
  NAND2_X1   g21553(.A1(new_n20898_), .A2(new_n19438_), .ZN(new_n21620_));
  NAND2_X1   g21554(.A1(new_n21619_), .A2(new_n21620_), .ZN(new_n21621_));
  INV_X1     g21555(.I(new_n21617_), .ZN(new_n21622_));
  OAI21_X1   g21556(.A1(new_n21621_), .A2(new_n21622_), .B(\a[5] ), .ZN(new_n21623_));
  NAND2_X1   g21557(.A1(new_n21618_), .A2(new_n21623_), .ZN(new_n21624_));
  OAI21_X1   g21558(.A1(new_n21612_), .A2(new_n21613_), .B(new_n21624_), .ZN(new_n21625_));
  NAND2_X1   g21559(.A1(new_n20661_), .A2(new_n20657_), .ZN(new_n21626_));
  XOR2_X1    g21560(.A1(new_n21626_), .A2(new_n20665_), .Z(new_n21627_));
  NOR2_X1    g21561(.A1(new_n21627_), .A2(new_n20613_), .ZN(new_n21628_));
  NAND2_X1   g21562(.A1(new_n20793_), .A2(new_n20667_), .ZN(new_n21629_));
  AOI21_X1   g21563(.A1(new_n20613_), .A2(new_n21629_), .B(new_n21628_), .ZN(new_n21630_));
  NAND4_X1   g21564(.A1(new_n21556_), .A2(new_n21477_), .A3(new_n21535_), .A4(new_n21540_), .ZN(new_n21631_));
  INV_X1     g21565(.I(new_n20134_), .ZN(new_n21632_));
  AOI22_X1   g21566(.A1(new_n19386_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n20127_), .ZN(new_n21633_));
  NOR2_X1    g21567(.A1(new_n17793_), .A2(new_n6091_), .ZN(new_n21634_));
  OAI21_X1   g21568(.A1(new_n21633_), .A2(new_n21634_), .B(new_n6081_), .ZN(new_n21635_));
  NOR2_X1    g21569(.A1(new_n21632_), .A2(new_n21635_), .ZN(new_n21636_));
  XOR2_X1    g21570(.A1(new_n21636_), .A2(new_n3521_), .Z(new_n21637_));
  INV_X1     g21571(.I(new_n21637_), .ZN(new_n21638_));
  AOI21_X1   g21572(.A1(new_n21631_), .A2(new_n21540_), .B(new_n21638_), .ZN(new_n21639_));
  NOR4_X1    g21573(.A1(new_n21519_), .A2(new_n21551_), .A3(new_n21552_), .A4(new_n21476_), .ZN(new_n21640_));
  NOR3_X1    g21574(.A1(new_n21640_), .A2(new_n21637_), .A3(new_n21552_), .ZN(new_n21641_));
  OAI21_X1   g21575(.A1(new_n21641_), .A2(new_n21639_), .B(new_n21630_), .ZN(new_n21642_));
  INV_X1     g21576(.I(new_n21630_), .ZN(new_n21643_));
  OAI21_X1   g21577(.A1(new_n21640_), .A2(new_n21552_), .B(new_n21637_), .ZN(new_n21644_));
  NAND3_X1   g21578(.A1(new_n21631_), .A2(new_n21638_), .A3(new_n21540_), .ZN(new_n21645_));
  NAND3_X1   g21579(.A1(new_n21644_), .A2(new_n21645_), .A3(new_n21643_), .ZN(new_n21646_));
  NAND2_X1   g21580(.A1(new_n21642_), .A2(new_n21646_), .ZN(new_n21647_));
  NOR3_X1    g21581(.A1(new_n21508_), .A2(new_n21560_), .A3(new_n21555_), .ZN(new_n21648_));
  NOR2_X1    g21582(.A1(new_n21551_), .A2(new_n21552_), .ZN(new_n21649_));
  NAND2_X1   g21583(.A1(new_n21557_), .A2(new_n21649_), .ZN(new_n21650_));
  NAND2_X1   g21584(.A1(new_n21540_), .A2(new_n21535_), .ZN(new_n21651_));
  NAND2_X1   g21585(.A1(new_n21520_), .A2(new_n21651_), .ZN(new_n21652_));
  AOI21_X1   g21586(.A1(new_n21650_), .A2(new_n21652_), .B(new_n21553_), .ZN(new_n21653_));
  OAI22_X1   g21587(.A1(new_n19400_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n19393_), .ZN(new_n21654_));
  NAND2_X1   g21588(.A1(new_n17790_), .A2(new_n4709_), .ZN(new_n21655_));
  AOI21_X1   g21589(.A1(new_n21655_), .A2(new_n21654_), .B(new_n4707_), .ZN(new_n21656_));
  NAND2_X1   g21590(.A1(new_n20251_), .A2(new_n21656_), .ZN(new_n21657_));
  XOR2_X1    g21591(.A1(new_n21657_), .A2(\a[11] ), .Z(new_n21658_));
  OAI21_X1   g21592(.A1(new_n21648_), .A2(new_n21653_), .B(new_n21658_), .ZN(new_n21659_));
  NAND3_X1   g21593(.A1(new_n21573_), .A2(new_n21576_), .A3(new_n21579_), .ZN(new_n21660_));
  NOR2_X1    g21594(.A1(new_n21520_), .A2(new_n21651_), .ZN(new_n21661_));
  NOR2_X1    g21595(.A1(new_n21557_), .A2(new_n21649_), .ZN(new_n21662_));
  OAI21_X1   g21596(.A1(new_n21662_), .A2(new_n21661_), .B(new_n21549_), .ZN(new_n21663_));
  XOR2_X1    g21597(.A1(new_n21657_), .A2(new_n4034_), .Z(new_n21664_));
  NAND3_X1   g21598(.A1(new_n21660_), .A2(new_n21663_), .A3(new_n21664_), .ZN(new_n21665_));
  AOI21_X1   g21599(.A1(new_n21659_), .A2(new_n21665_), .B(new_n21647_), .ZN(new_n21666_));
  AOI21_X1   g21600(.A1(new_n21644_), .A2(new_n21645_), .B(new_n21643_), .ZN(new_n21667_));
  NOR3_X1    g21601(.A1(new_n21641_), .A2(new_n21639_), .A3(new_n21630_), .ZN(new_n21668_));
  NOR2_X1    g21602(.A1(new_n21668_), .A2(new_n21667_), .ZN(new_n21669_));
  AOI21_X1   g21603(.A1(new_n21660_), .A2(new_n21663_), .B(new_n21664_), .ZN(new_n21670_));
  NOR3_X1    g21604(.A1(new_n21648_), .A2(new_n21658_), .A3(new_n21653_), .ZN(new_n21671_));
  NOR3_X1    g21605(.A1(new_n21671_), .A2(new_n21669_), .A3(new_n21670_), .ZN(new_n21672_));
  NOR2_X1    g21606(.A1(new_n21666_), .A2(new_n21672_), .ZN(new_n21673_));
  NAND3_X1   g21607(.A1(new_n21508_), .A2(new_n21573_), .A3(new_n21576_), .ZN(new_n21674_));
  OAI21_X1   g21608(.A1(new_n21560_), .A2(new_n21555_), .B(new_n21579_), .ZN(new_n21675_));
  AOI21_X1   g21609(.A1(new_n21674_), .A2(new_n21675_), .B(new_n21569_), .ZN(new_n21676_));
  INV_X1     g21610(.I(new_n21676_), .ZN(new_n21677_));
  OAI22_X1   g21611(.A1(new_n19410_), .A2(new_n6783_), .B1(new_n19412_), .B2(new_n6788_), .ZN(new_n21678_));
  OAI21_X1   g21612(.A1(new_n17787_), .A2(new_n6785_), .B(new_n21678_), .ZN(new_n21679_));
  NAND4_X1   g21613(.A1(new_n20949_), .A2(new_n6775_), .A3(new_n20824_), .A4(new_n21679_), .ZN(new_n21680_));
  XOR2_X1    g21614(.A1(new_n21680_), .A2(new_n4009_), .Z(new_n21681_));
  AOI21_X1   g21615(.A1(new_n21586_), .A2(new_n21677_), .B(new_n21681_), .ZN(new_n21682_));
  NOR3_X1    g21616(.A1(new_n21593_), .A2(new_n21590_), .A3(new_n21587_), .ZN(new_n21683_));
  XOR2_X1    g21617(.A1(new_n21680_), .A2(\a[8] ), .Z(new_n21684_));
  NOR3_X1    g21618(.A1(new_n21683_), .A2(new_n21676_), .A3(new_n21684_), .ZN(new_n21685_));
  OAI21_X1   g21619(.A1(new_n21685_), .A2(new_n21682_), .B(new_n21673_), .ZN(new_n21686_));
  OAI21_X1   g21620(.A1(new_n21670_), .A2(new_n21671_), .B(new_n21669_), .ZN(new_n21687_));
  NAND3_X1   g21621(.A1(new_n21659_), .A2(new_n21647_), .A3(new_n21665_), .ZN(new_n21688_));
  NAND2_X1   g21622(.A1(new_n21687_), .A2(new_n21688_), .ZN(new_n21689_));
  OAI21_X1   g21623(.A1(new_n21683_), .A2(new_n21676_), .B(new_n21684_), .ZN(new_n21690_));
  NAND3_X1   g21624(.A1(new_n21586_), .A2(new_n21677_), .A3(new_n21681_), .ZN(new_n21691_));
  NAND3_X1   g21625(.A1(new_n21690_), .A2(new_n21691_), .A3(new_n21689_), .ZN(new_n21692_));
  NAND2_X1   g21626(.A1(new_n21686_), .A2(new_n21692_), .ZN(new_n21693_));
  NOR3_X1    g21627(.A1(new_n21624_), .A2(new_n21612_), .A3(new_n21613_), .ZN(new_n21694_));
  OAI21_X1   g21628(.A1(new_n21693_), .A2(new_n21694_), .B(new_n21625_), .ZN(new_n21695_));
  OAI21_X1   g21629(.A1(new_n21695_), .A2(new_n21243_), .B(new_n21241_), .ZN(new_n21696_));
  AOI21_X1   g21630(.A1(new_n21216_), .A2(new_n21220_), .B(new_n21224_), .ZN(new_n21697_));
  INV_X1     g21631(.I(new_n21697_), .ZN(new_n21698_));
  OAI21_X1   g21632(.A1(new_n21696_), .A2(new_n21228_), .B(new_n21698_), .ZN(new_n21699_));
  NOR2_X1    g21633(.A1(new_n21012_), .A2(new_n21013_), .ZN(new_n21700_));
  NOR2_X1    g21634(.A1(new_n21066_), .A2(new_n20954_), .ZN(new_n21701_));
  NOR2_X1    g21635(.A1(new_n21040_), .A2(new_n21011_), .ZN(new_n21702_));
  OAI21_X1   g21636(.A1(new_n21701_), .A2(new_n21702_), .B(new_n21700_), .ZN(new_n21703_));
  INV_X1     g21637(.I(new_n21700_), .ZN(new_n21704_));
  NAND2_X1   g21638(.A1(new_n21040_), .A2(new_n21011_), .ZN(new_n21705_));
  NAND2_X1   g21639(.A1(new_n21066_), .A2(new_n20954_), .ZN(new_n21706_));
  NAND3_X1   g21640(.A1(new_n21706_), .A2(new_n21705_), .A3(new_n21704_), .ZN(new_n21707_));
  NAND2_X1   g21641(.A1(new_n21707_), .A2(new_n21703_), .ZN(new_n21708_));
  NAND3_X1   g21642(.A1(new_n21205_), .A2(new_n21207_), .A3(new_n21219_), .ZN(new_n21709_));
  AOI22_X1   g21643(.A1(new_n20896_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n19442_), .ZN(new_n21710_));
  NOR2_X1    g21644(.A1(new_n17784_), .A2(new_n6785_), .ZN(new_n21711_));
  OAI21_X1   g21645(.A1(new_n21710_), .A2(new_n21711_), .B(new_n6775_), .ZN(new_n21712_));
  INV_X1     g21646(.I(new_n21712_), .ZN(new_n21713_));
  NAND2_X1   g21647(.A1(new_n20907_), .A2(new_n21713_), .ZN(new_n21714_));
  NOR2_X1    g21648(.A1(new_n21714_), .A2(\a[8] ), .ZN(new_n21715_));
  AOI21_X1   g21649(.A1(new_n20907_), .A2(new_n21713_), .B(new_n4009_), .ZN(new_n21716_));
  NOR2_X1    g21650(.A1(new_n21715_), .A2(new_n21716_), .ZN(new_n21717_));
  NAND2_X1   g21651(.A1(new_n21709_), .A2(new_n21717_), .ZN(new_n21718_));
  NOR3_X1    g21652(.A1(new_n21218_), .A2(new_n21217_), .A3(new_n21215_), .ZN(new_n21719_));
  INV_X1     g21653(.I(new_n21717_), .ZN(new_n21720_));
  NAND2_X1   g21654(.A1(new_n21720_), .A2(new_n21719_), .ZN(new_n21721_));
  AOI21_X1   g21655(.A1(new_n21721_), .A2(new_n21718_), .B(new_n21708_), .ZN(new_n21722_));
  AOI21_X1   g21656(.A1(new_n21706_), .A2(new_n21705_), .B(new_n21704_), .ZN(new_n21723_));
  NOR3_X1    g21657(.A1(new_n21701_), .A2(new_n21702_), .A3(new_n21700_), .ZN(new_n21724_));
  NOR2_X1    g21658(.A1(new_n21723_), .A2(new_n21724_), .ZN(new_n21725_));
  NOR2_X1    g21659(.A1(new_n21720_), .A2(new_n21719_), .ZN(new_n21726_));
  NOR2_X1    g21660(.A1(new_n21709_), .A2(new_n21717_), .ZN(new_n21727_));
  NOR3_X1    g21661(.A1(new_n21726_), .A2(new_n21725_), .A3(new_n21727_), .ZN(new_n21728_));
  NAND3_X1   g21662(.A1(new_n21084_), .A2(new_n21086_), .A3(new_n19475_), .ZN(new_n21729_));
  OAI21_X1   g21663(.A1(new_n21082_), .A2(new_n21077_), .B(new_n17780_), .ZN(new_n21730_));
  OAI22_X1   g21664(.A1(new_n19463_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n19437_), .ZN(new_n21731_));
  NAND2_X1   g21665(.A1(new_n17780_), .A2(new_n6838_), .ZN(new_n21732_));
  AOI21_X1   g21666(.A1(new_n21731_), .A2(new_n21732_), .B(new_n6836_), .ZN(new_n21733_));
  NAND3_X1   g21667(.A1(new_n21730_), .A2(new_n21729_), .A3(new_n21733_), .ZN(new_n21734_));
  XOR2_X1    g21668(.A1(new_n21734_), .A2(new_n65_), .Z(new_n21735_));
  NOR3_X1    g21669(.A1(new_n21735_), .A2(new_n21722_), .A3(new_n21728_), .ZN(new_n21736_));
  OAI21_X1   g21670(.A1(new_n21722_), .A2(new_n21728_), .B(new_n21735_), .ZN(new_n21737_));
  OAI21_X1   g21671(.A1(new_n21699_), .A2(new_n21736_), .B(new_n21737_), .ZN(new_n21738_));
  AOI21_X1   g21672(.A1(new_n21106_), .A2(new_n21107_), .B(new_n21130_), .ZN(new_n21739_));
  NOR2_X1    g21673(.A1(new_n21108_), .A2(new_n21105_), .ZN(new_n21740_));
  NOR3_X1    g21674(.A1(new_n21180_), .A2(new_n21181_), .A3(\a[5] ), .ZN(new_n21741_));
  AOI21_X1   g21675(.A1(new_n21171_), .A2(new_n21174_), .B(new_n65_), .ZN(new_n21742_));
  NOR2_X1    g21676(.A1(new_n21741_), .A2(new_n21742_), .ZN(new_n21743_));
  NOR3_X1    g21677(.A1(new_n21743_), .A2(new_n21740_), .A3(new_n21739_), .ZN(new_n21744_));
  OAI21_X1   g21678(.A1(new_n21738_), .A2(new_n21744_), .B(new_n21185_), .ZN(new_n21745_));
  NAND3_X1   g21679(.A1(new_n21745_), .A2(new_n21163_), .A3(new_n21164_), .ZN(new_n21746_));
  AOI22_X1   g21680(.A1(new_n21147_), .A2(new_n21143_), .B1(new_n21746_), .B2(new_n19527_), .ZN(new_n21747_));
  NAND2_X1   g21681(.A1(new_n20118_), .A2(new_n20056_), .ZN(new_n21748_));
  NOR2_X1    g21682(.A1(new_n20224_), .A2(new_n20154_), .ZN(new_n21749_));
  NAND3_X1   g21683(.A1(new_n20117_), .A2(new_n20116_), .A3(new_n20115_), .ZN(new_n21750_));
  OAI21_X1   g21684(.A1(new_n21749_), .A2(new_n20225_), .B(new_n21750_), .ZN(new_n21751_));
  NAND2_X1   g21685(.A1(new_n21751_), .A2(new_n21748_), .ZN(new_n21752_));
  NAND2_X1   g21686(.A1(new_n20709_), .A2(new_n20708_), .ZN(new_n21753_));
  AOI22_X1   g21687(.A1(new_n17798_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n17802_), .ZN(new_n21754_));
  NOR2_X1    g21688(.A1(new_n19375_), .A2(new_n3780_), .ZN(new_n21755_));
  OAI21_X1   g21689(.A1(new_n21755_), .A2(new_n21754_), .B(new_n3301_), .ZN(new_n21756_));
  NOR2_X1    g21690(.A1(new_n21753_), .A2(new_n21756_), .ZN(new_n21757_));
  XOR2_X1    g21691(.A1(new_n21757_), .A2(\a[23] ), .Z(new_n21758_));
  NOR2_X1    g21692(.A1(new_n20065_), .A2(new_n20085_), .ZN(new_n21759_));
  OAI21_X1   g21693(.A1(new_n20057_), .A2(new_n21759_), .B(new_n20092_), .ZN(new_n21760_));
  INV_X1     g21694(.I(new_n21760_), .ZN(new_n21761_));
  OAI22_X1   g21695(.A1(new_n2742_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n2747_), .ZN(new_n21762_));
  NAND2_X1   g21696(.A1(new_n19350_), .A2(new_n2750_), .ZN(new_n21763_));
  AOI21_X1   g21697(.A1(new_n21762_), .A2(new_n21763_), .B(new_n2737_), .ZN(new_n21764_));
  NAND3_X1   g21698(.A1(new_n20535_), .A2(new_n74_), .A3(new_n21764_), .ZN(new_n21765_));
  NAND2_X1   g21699(.A1(new_n20535_), .A2(new_n21764_), .ZN(new_n21766_));
  NAND2_X1   g21700(.A1(new_n21766_), .A2(\a[29] ), .ZN(new_n21767_));
  NAND2_X1   g21701(.A1(new_n21767_), .A2(new_n21765_), .ZN(new_n21768_));
  INV_X1     g21702(.I(new_n20081_), .ZN(new_n21769_));
  OAI21_X1   g21703(.A1(new_n20067_), .A2(new_n20080_), .B(new_n21769_), .ZN(new_n21770_));
  NOR2_X1    g21704(.A1(new_n19304_), .A2(new_n2767_), .ZN(new_n21771_));
  NOR2_X1    g21705(.A1(new_n19320_), .A2(new_n2772_), .ZN(new_n21772_));
  NOR2_X1    g21706(.A1(new_n17849_), .A2(new_n2771_), .ZN(new_n21773_));
  NOR4_X1    g21707(.A1(new_n21771_), .A2(new_n2763_), .A3(new_n21772_), .A4(new_n21773_), .ZN(new_n21774_));
  NAND2_X1   g21708(.A1(new_n19647_), .A2(new_n21774_), .ZN(new_n21775_));
  INV_X1     g21709(.I(new_n2998_), .ZN(new_n21776_));
  NAND4_X1   g21710(.A1(new_n784_), .A2(new_n2855_), .A3(new_n1329_), .A4(new_n1199_), .ZN(new_n21777_));
  NOR3_X1    g21711(.A1(new_n11550_), .A2(new_n3680_), .A3(new_n21777_), .ZN(new_n21778_));
  NAND3_X1   g21712(.A1(new_n2260_), .A2(new_n442_), .A3(new_n391_), .ZN(new_n21779_));
  NOR3_X1    g21713(.A1(new_n1508_), .A2(new_n563_), .A3(new_n422_), .ZN(new_n21780_));
  NAND4_X1   g21714(.A1(new_n21778_), .A2(new_n21776_), .A3(new_n21779_), .A4(new_n21780_), .ZN(new_n21781_));
  NOR3_X1    g21715(.A1(new_n11516_), .A2(new_n3499_), .A3(new_n21781_), .ZN(new_n21782_));
  INV_X1     g21716(.I(new_n21782_), .ZN(new_n21783_));
  NAND2_X1   g21717(.A1(new_n21775_), .A2(new_n21783_), .ZN(new_n21784_));
  NOR2_X1    g21718(.A1(new_n21775_), .A2(new_n21783_), .ZN(new_n21785_));
  INV_X1     g21719(.I(new_n21785_), .ZN(new_n21786_));
  NAND2_X1   g21720(.A1(new_n21786_), .A2(new_n21784_), .ZN(new_n21787_));
  XOR2_X1    g21721(.A1(new_n21775_), .A2(new_n21782_), .Z(new_n21788_));
  NOR2_X1    g21722(.A1(new_n21770_), .A2(new_n21788_), .ZN(new_n21789_));
  AOI21_X1   g21723(.A1(new_n21770_), .A2(new_n21787_), .B(new_n21789_), .ZN(new_n21790_));
  XOR2_X1    g21724(.A1(new_n21768_), .A2(new_n21790_), .Z(new_n21791_));
  NOR2_X1    g21725(.A1(new_n21791_), .A2(new_n21761_), .ZN(new_n21792_));
  NAND3_X1   g21726(.A1(new_n21790_), .A2(new_n21765_), .A3(new_n21767_), .ZN(new_n21793_));
  AOI21_X1   g21727(.A1(new_n21765_), .A2(new_n21767_), .B(new_n21790_), .ZN(new_n21794_));
  INV_X1     g21728(.I(new_n21794_), .ZN(new_n21795_));
  AOI21_X1   g21729(.A1(new_n21795_), .A2(new_n21793_), .B(new_n21760_), .ZN(new_n21796_));
  NOR2_X1    g21730(.A1(new_n21792_), .A2(new_n21796_), .ZN(new_n21797_));
  OAI22_X1   g21731(.A1(new_n19356_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n17806_), .ZN(new_n21798_));
  NAND2_X1   g21732(.A1(new_n19365_), .A2(new_n3317_), .ZN(new_n21799_));
  AOI21_X1   g21733(.A1(new_n21798_), .A2(new_n21799_), .B(new_n3260_), .ZN(new_n21800_));
  NAND2_X1   g21734(.A1(new_n19538_), .A2(new_n21800_), .ZN(new_n21801_));
  XOR2_X1    g21735(.A1(new_n21801_), .A2(\a[26] ), .Z(new_n21802_));
  INV_X1     g21736(.I(new_n21802_), .ZN(new_n21803_));
  XOR2_X1    g21737(.A1(new_n21797_), .A2(new_n21803_), .Z(new_n21804_));
  XOR2_X1    g21738(.A1(new_n21804_), .A2(new_n21758_), .Z(new_n21805_));
  NAND2_X1   g21739(.A1(new_n21752_), .A2(new_n21805_), .ZN(new_n21806_));
  AOI21_X1   g21740(.A1(new_n20036_), .A2(new_n20040_), .B(new_n20122_), .ZN(new_n21807_));
  NOR2_X1    g21741(.A1(new_n21807_), .A2(new_n20123_), .ZN(new_n21808_));
  NOR2_X1    g21742(.A1(new_n21804_), .A2(new_n21758_), .ZN(new_n21809_));
  XOR2_X1    g21743(.A1(new_n21757_), .A2(new_n84_), .Z(new_n21810_));
  XOR2_X1    g21744(.A1(new_n21797_), .A2(new_n21802_), .Z(new_n21811_));
  NOR2_X1    g21745(.A1(new_n21811_), .A2(new_n21810_), .ZN(new_n21812_));
  OAI21_X1   g21746(.A1(new_n21809_), .A2(new_n21812_), .B(new_n21808_), .ZN(new_n21813_));
  AOI22_X1   g21747(.A1(new_n19386_), .A2(new_n3770_), .B1(new_n3776_), .B2(new_n17794_), .ZN(new_n21814_));
  NOR2_X1    g21748(.A1(new_n19393_), .A2(new_n4097_), .ZN(new_n21815_));
  OAI21_X1   g21749(.A1(new_n21814_), .A2(new_n21815_), .B(new_n3773_), .ZN(new_n21816_));
  NOR2_X1    g21750(.A1(new_n20291_), .A2(new_n21816_), .ZN(new_n21817_));
  XOR2_X1    g21751(.A1(new_n21817_), .A2(new_n3035_), .Z(new_n21818_));
  NAND3_X1   g21752(.A1(new_n21813_), .A2(new_n21806_), .A3(new_n21818_), .ZN(new_n21819_));
  AOI21_X1   g21753(.A1(new_n21813_), .A2(new_n21806_), .B(new_n21818_), .ZN(new_n21820_));
  INV_X1     g21754(.I(new_n21820_), .ZN(new_n21821_));
  AOI22_X1   g21755(.A1(new_n17790_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n19399_), .ZN(new_n21822_));
  NOR2_X1    g21756(.A1(new_n19410_), .A2(new_n4470_), .ZN(new_n21823_));
  OAI21_X1   g21757(.A1(new_n21823_), .A2(new_n21822_), .B(new_n4295_), .ZN(new_n21824_));
  OR3_X2     g21758(.A1(new_n20863_), .A2(\a[17] ), .A3(new_n21824_), .Z(new_n21825_));
  OAI21_X1   g21759(.A1(new_n20863_), .A2(new_n21824_), .B(\a[17] ), .ZN(new_n21826_));
  NAND4_X1   g21760(.A1(new_n21821_), .A2(new_n21819_), .A3(new_n21825_), .A4(new_n21826_), .ZN(new_n21827_));
  INV_X1     g21761(.I(new_n21819_), .ZN(new_n21828_));
  NAND2_X1   g21762(.A1(new_n21825_), .A2(new_n21826_), .ZN(new_n21829_));
  OAI21_X1   g21763(.A1(new_n21828_), .A2(new_n21820_), .B(new_n21829_), .ZN(new_n21830_));
  NAND2_X1   g21764(.A1(new_n21827_), .A2(new_n21830_), .ZN(new_n21831_));
  OAI21_X1   g21765(.A1(new_n20235_), .A2(new_n20236_), .B(new_n20234_), .ZN(new_n21832_));
  NAND3_X1   g21766(.A1(new_n20231_), .A2(new_n20213_), .A3(new_n20125_), .ZN(new_n21833_));
  NAND3_X1   g21767(.A1(new_n21832_), .A2(new_n21833_), .A3(new_n20258_), .ZN(new_n21834_));
  OAI21_X1   g21768(.A1(new_n20232_), .A2(new_n20237_), .B(new_n20815_), .ZN(new_n21835_));
  AOI22_X1   g21769(.A1(new_n21835_), .A2(new_n21834_), .B1(new_n20816_), .B2(new_n20258_), .ZN(new_n21836_));
  XOR2_X1    g21770(.A1(new_n21836_), .A2(new_n21831_), .Z(new_n21837_));
  OAI22_X1   g21771(.A1(new_n17787_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n19412_), .ZN(new_n21838_));
  NAND2_X1   g21772(.A1(new_n19442_), .A2(new_n6090_), .ZN(new_n21839_));
  AOI21_X1   g21773(.A1(new_n21839_), .A2(new_n21838_), .B(new_n6082_), .ZN(new_n21840_));
  NAND2_X1   g21774(.A1(new_n20939_), .A2(new_n21840_), .ZN(new_n21841_));
  XOR2_X1    g21775(.A1(new_n21841_), .A2(\a[14] ), .Z(new_n21842_));
  INV_X1     g21776(.I(new_n21842_), .ZN(new_n21843_));
  NOR2_X1    g21777(.A1(new_n21837_), .A2(new_n21843_), .ZN(new_n21844_));
  NOR3_X1    g21778(.A1(new_n20232_), .A2(new_n20237_), .A3(new_n20815_), .ZN(new_n21845_));
  AOI21_X1   g21779(.A1(new_n21832_), .A2(new_n21833_), .B(new_n20258_), .ZN(new_n21846_));
  OAI22_X1   g21780(.A1(new_n21845_), .A2(new_n21846_), .B1(new_n20775_), .B2(new_n20815_), .ZN(new_n21847_));
  NOR2_X1    g21781(.A1(new_n21847_), .A2(new_n21831_), .ZN(new_n21848_));
  NOR3_X1    g21782(.A1(new_n21828_), .A2(new_n21820_), .A3(new_n21829_), .ZN(new_n21849_));
  AOI22_X1   g21783(.A1(new_n21821_), .A2(new_n21819_), .B1(new_n21825_), .B2(new_n21826_), .ZN(new_n21850_));
  NOR2_X1    g21784(.A1(new_n21850_), .A2(new_n21849_), .ZN(new_n21851_));
  NOR2_X1    g21785(.A1(new_n21836_), .A2(new_n21851_), .ZN(new_n21852_));
  NOR2_X1    g21786(.A1(new_n21848_), .A2(new_n21852_), .ZN(new_n21853_));
  NOR2_X1    g21787(.A1(new_n21853_), .A2(new_n21842_), .ZN(new_n21854_));
  AOI22_X1   g21788(.A1(new_n19438_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n20896_), .ZN(new_n21855_));
  AOI21_X1   g21789(.A1(new_n19466_), .A2(new_n4709_), .B(new_n21855_), .ZN(new_n21856_));
  NOR4_X1    g21790(.A1(new_n21098_), .A2(new_n21099_), .A3(new_n4707_), .A4(new_n21856_), .ZN(new_n21857_));
  XOR2_X1    g21791(.A1(new_n21857_), .A2(\a[11] ), .Z(new_n21858_));
  NOR3_X1    g21792(.A1(new_n21858_), .A2(new_n21844_), .A3(new_n21854_), .ZN(new_n21859_));
  NAND2_X1   g21793(.A1(new_n21853_), .A2(new_n21842_), .ZN(new_n21860_));
  NAND2_X1   g21794(.A1(new_n21837_), .A2(new_n21843_), .ZN(new_n21861_));
  XOR2_X1    g21795(.A1(new_n21857_), .A2(new_n4034_), .Z(new_n21862_));
  AOI21_X1   g21796(.A1(new_n21861_), .A2(new_n21860_), .B(new_n21862_), .ZN(new_n21863_));
  NOR2_X1    g21797(.A1(new_n21863_), .A2(new_n21859_), .ZN(new_n21864_));
  OAI21_X1   g21798(.A1(new_n20888_), .A2(new_n20887_), .B(new_n20886_), .ZN(new_n21865_));
  NAND3_X1   g21799(.A1(new_n20874_), .A2(new_n20882_), .A3(new_n20819_), .ZN(new_n21866_));
  NAND3_X1   g21800(.A1(new_n21865_), .A2(new_n21866_), .A3(new_n21052_), .ZN(new_n21867_));
  OAI21_X1   g21801(.A1(new_n20889_), .A2(new_n20883_), .B(new_n20912_), .ZN(new_n21868_));
  AOI22_X1   g21802(.A1(new_n21048_), .A2(new_n21052_), .B1(new_n21868_), .B2(new_n21867_), .ZN(new_n21869_));
  NAND2_X1   g21803(.A1(new_n21869_), .A2(new_n21864_), .ZN(new_n21870_));
  NAND3_X1   g21804(.A1(new_n21862_), .A2(new_n21861_), .A3(new_n21860_), .ZN(new_n21871_));
  OAI21_X1   g21805(.A1(new_n21844_), .A2(new_n21854_), .B(new_n21858_), .ZN(new_n21872_));
  NAND2_X1   g21806(.A1(new_n21872_), .A2(new_n21871_), .ZN(new_n21873_));
  NOR3_X1    g21807(.A1(new_n20889_), .A2(new_n20883_), .A3(new_n20912_), .ZN(new_n21874_));
  AOI21_X1   g21808(.A1(new_n21865_), .A2(new_n21866_), .B(new_n21052_), .ZN(new_n21875_));
  OAI22_X1   g21809(.A1(new_n21071_), .A2(new_n20912_), .B1(new_n21874_), .B2(new_n21875_), .ZN(new_n21876_));
  NAND2_X1   g21810(.A1(new_n21876_), .A2(new_n21873_), .ZN(new_n21877_));
  NAND2_X1   g21811(.A1(new_n21877_), .A2(new_n21870_), .ZN(new_n21878_));
  OAI22_X1   g21812(.A1(new_n19475_), .A2(new_n6788_), .B1(new_n19463_), .B2(new_n6783_), .ZN(new_n21879_));
  NAND2_X1   g21813(.A1(new_n19484_), .A2(new_n6784_), .ZN(new_n21880_));
  AOI21_X1   g21814(.A1(new_n21880_), .A2(new_n21879_), .B(new_n6776_), .ZN(new_n21881_));
  NAND2_X1   g21815(.A1(new_n21171_), .A2(new_n21881_), .ZN(new_n21882_));
  XOR2_X1    g21816(.A1(new_n21882_), .A2(\a[8] ), .Z(new_n21883_));
  NOR2_X1    g21817(.A1(new_n21878_), .A2(new_n21883_), .ZN(new_n21884_));
  INV_X1     g21818(.I(new_n21884_), .ZN(new_n21885_));
  NAND2_X1   g21819(.A1(new_n21878_), .A2(new_n21883_), .ZN(new_n21886_));
  OAI21_X1   g21820(.A1(new_n19512_), .A2(new_n17775_), .B(new_n19522_), .ZN(new_n21887_));
  AOI21_X1   g21821(.A1(new_n19512_), .A2(new_n17775_), .B(new_n19522_), .ZN(new_n21888_));
  AOI21_X1   g21822(.A1(new_n21151_), .A2(new_n21887_), .B(new_n21888_), .ZN(new_n21889_));
  NAND2_X1   g21823(.A1(new_n17766_), .A2(new_n17765_), .ZN(new_n21890_));
  XOR2_X1    g21824(.A1(new_n11777_), .A2(new_n17765_), .Z(new_n21891_));
  NAND3_X1   g21825(.A1(new_n17758_), .A2(new_n17760_), .A3(new_n21891_), .ZN(new_n21892_));
  OAI21_X1   g21826(.A1(new_n11752_), .A2(new_n11764_), .B(new_n11766_), .ZN(new_n21893_));
  INV_X1     g21827(.I(new_n21893_), .ZN(new_n21894_));
  AOI21_X1   g21828(.A1(new_n11749_), .A2(new_n11743_), .B(new_n11746_), .ZN(new_n21895_));
  NOR2_X1    g21829(.A1(new_n11277_), .A2(new_n2772_), .ZN(new_n21896_));
  NOR2_X1    g21830(.A1(new_n11284_), .A2(new_n2771_), .ZN(new_n21897_));
  NOR2_X1    g21831(.A1(new_n11271_), .A2(new_n2767_), .ZN(new_n21898_));
  NOR4_X1    g21832(.A1(new_n21897_), .A2(new_n2763_), .A3(new_n21896_), .A4(new_n21898_), .ZN(new_n21899_));
  NAND2_X1   g21833(.A1(new_n11391_), .A2(new_n21899_), .ZN(new_n21900_));
  AOI21_X1   g21834(.A1(new_n11713_), .A2(new_n11731_), .B(new_n11732_), .ZN(new_n21901_));
  INV_X1     g21835(.I(new_n2612_), .ZN(new_n21902_));
  INV_X1     g21836(.I(new_n4859_), .ZN(new_n21903_));
  NOR2_X1    g21837(.A1(new_n2884_), .A2(new_n2306_), .ZN(new_n21904_));
  NAND4_X1   g21838(.A1(new_n373_), .A2(new_n1805_), .A3(new_n1892_), .A4(new_n809_), .ZN(new_n21905_));
  NAND4_X1   g21839(.A1(new_n21904_), .A2(new_n2620_), .A3(new_n21903_), .A4(new_n21905_), .ZN(new_n21906_));
  NOR4_X1    g21840(.A1(new_n2582_), .A2(new_n1511_), .A3(new_n1116_), .A4(new_n1994_), .ZN(new_n21907_));
  NAND4_X1   g21841(.A1(new_n21907_), .A2(new_n1063_), .A3(new_n1753_), .A4(new_n849_), .ZN(new_n21908_));
  NOR4_X1    g21842(.A1(new_n11043_), .A2(new_n21902_), .A3(new_n21906_), .A4(new_n21908_), .ZN(new_n21909_));
  NOR2_X1    g21843(.A1(new_n581_), .A2(new_n622_), .ZN(new_n21910_));
  NAND2_X1   g21844(.A1(new_n21910_), .A2(new_n21909_), .ZN(new_n21911_));
  XOR2_X1    g21845(.A1(new_n21901_), .A2(new_n21911_), .Z(new_n21912_));
  NOR2_X1    g21846(.A1(new_n21900_), .A2(new_n21912_), .ZN(new_n21913_));
  INV_X1     g21847(.I(new_n21911_), .ZN(new_n21914_));
  NOR2_X1    g21848(.A1(new_n21901_), .A2(new_n21914_), .ZN(new_n21915_));
  NAND2_X1   g21849(.A1(new_n21901_), .A2(new_n21914_), .ZN(new_n21916_));
  INV_X1     g21850(.I(new_n21916_), .ZN(new_n21917_));
  NOR2_X1    g21851(.A1(new_n21917_), .A2(new_n21915_), .ZN(new_n21918_));
  INV_X1     g21852(.I(new_n21918_), .ZN(new_n21919_));
  AOI21_X1   g21853(.A1(new_n21900_), .A2(new_n21919_), .B(new_n21913_), .ZN(new_n21920_));
  OAI22_X1   g21854(.A1(new_n11264_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n11345_), .ZN(new_n21921_));
  NAND2_X1   g21855(.A1(new_n11354_), .A2(new_n2750_), .ZN(new_n21922_));
  AOI21_X1   g21856(.A1(new_n21922_), .A2(new_n21921_), .B(new_n2737_), .ZN(new_n21923_));
  NAND2_X1   g21857(.A1(new_n11678_), .A2(new_n21923_), .ZN(new_n21924_));
  XOR2_X1    g21858(.A1(new_n21924_), .A2(\a[29] ), .Z(new_n21925_));
  XOR2_X1    g21859(.A1(new_n21925_), .A2(new_n21920_), .Z(new_n21926_));
  NOR2_X1    g21860(.A1(new_n21926_), .A2(new_n21895_), .ZN(new_n21927_));
  INV_X1     g21861(.I(new_n21895_), .ZN(new_n21928_));
  INV_X1     g21862(.I(new_n21920_), .ZN(new_n21929_));
  NAND2_X1   g21863(.A1(new_n21925_), .A2(new_n21929_), .ZN(new_n21930_));
  OR2_X2     g21864(.A1(new_n21925_), .A2(new_n21929_), .Z(new_n21931_));
  AOI21_X1   g21865(.A1(new_n21931_), .A2(new_n21930_), .B(new_n21928_), .ZN(new_n21932_));
  NOR2_X1    g21866(.A1(new_n21927_), .A2(new_n21932_), .ZN(new_n21933_));
  OAI22_X1   g21867(.A1(new_n11369_), .A2(new_n3268_), .B1(new_n3318_), .B2(new_n11461_), .ZN(new_n21934_));
  NAND2_X1   g21868(.A1(new_n11694_), .A2(new_n3323_), .ZN(new_n21935_));
  AOI21_X1   g21869(.A1(new_n21934_), .A2(new_n21935_), .B(new_n3260_), .ZN(new_n21936_));
  NAND2_X1   g21870(.A1(new_n12720_), .A2(new_n21936_), .ZN(new_n21937_));
  XOR2_X1    g21871(.A1(new_n21937_), .A2(\a[26] ), .Z(new_n21938_));
  INV_X1     g21872(.I(new_n21938_), .ZN(new_n21939_));
  NOR2_X1    g21873(.A1(new_n21933_), .A2(new_n21939_), .ZN(new_n21940_));
  NOR3_X1    g21874(.A1(new_n21927_), .A2(new_n21938_), .A3(new_n21932_), .ZN(new_n21941_));
  NOR2_X1    g21875(.A1(new_n21940_), .A2(new_n21941_), .ZN(new_n21942_));
  NOR2_X1    g21876(.A1(new_n21942_), .A2(new_n21894_), .ZN(new_n21943_));
  XOR2_X1    g21877(.A1(new_n21933_), .A2(new_n21939_), .Z(new_n21944_));
  AOI21_X1   g21878(.A1(new_n21894_), .A2(new_n21944_), .B(new_n21943_), .ZN(new_n21945_));
  NOR2_X1    g21879(.A1(new_n11771_), .A2(new_n11774_), .ZN(new_n21946_));
  NOR2_X1    g21880(.A1(new_n21946_), .A2(new_n11772_), .ZN(new_n21947_));
  XOR2_X1    g21881(.A1(new_n21945_), .A2(new_n21947_), .Z(new_n21948_));
  INV_X1     g21882(.I(new_n21948_), .ZN(new_n21949_));
  NAND3_X1   g21883(.A1(new_n21892_), .A2(new_n21890_), .A3(new_n21949_), .ZN(new_n21950_));
  AOI21_X1   g21884(.A1(new_n21892_), .A2(new_n21890_), .B(new_n21949_), .ZN(new_n21951_));
  INV_X1     g21885(.I(new_n21951_), .ZN(new_n21952_));
  NAND2_X1   g21886(.A1(new_n21952_), .A2(new_n21950_), .ZN(new_n21953_));
  XOR2_X1    g21887(.A1(new_n17770_), .A2(new_n21953_), .Z(new_n21954_));
  NOR2_X1    g21888(.A1(new_n21889_), .A2(new_n21954_), .ZN(new_n21955_));
  INV_X1     g21889(.I(new_n21151_), .ZN(new_n21956_));
  NAND2_X1   g21890(.A1(new_n17770_), .A2(new_n19484_), .ZN(new_n21957_));
  AOI21_X1   g21891(.A1(new_n21957_), .A2(new_n19522_), .B(new_n21956_), .ZN(new_n21958_));
  INV_X1     g21892(.I(new_n21950_), .ZN(new_n21959_));
  NOR2_X1    g21893(.A1(new_n21959_), .A2(new_n21951_), .ZN(new_n21960_));
  XOR2_X1    g21894(.A1(new_n17770_), .A2(new_n21960_), .Z(new_n21961_));
  NOR3_X1    g21895(.A1(new_n21961_), .A2(new_n21958_), .A3(new_n21888_), .ZN(new_n21962_));
  NOR2_X1    g21896(.A1(new_n21955_), .A2(new_n21962_), .ZN(new_n21963_));
  OAI22_X1   g21897(.A1(new_n19512_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n19522_), .ZN(new_n21964_));
  NAND2_X1   g21898(.A1(new_n21953_), .A2(new_n6838_), .ZN(new_n21965_));
  AOI21_X1   g21899(.A1(new_n21964_), .A2(new_n21965_), .B(new_n6836_), .ZN(new_n21966_));
  NAND3_X1   g21900(.A1(new_n21963_), .A2(new_n65_), .A3(new_n21966_), .ZN(new_n21967_));
  NAND2_X1   g21901(.A1(new_n21887_), .A2(new_n21151_), .ZN(new_n21968_));
  OAI21_X1   g21902(.A1(new_n17770_), .A2(new_n19484_), .B(new_n21157_), .ZN(new_n21969_));
  NAND2_X1   g21903(.A1(new_n21968_), .A2(new_n21969_), .ZN(new_n21970_));
  XOR2_X1    g21904(.A1(new_n17770_), .A2(new_n21960_), .Z(new_n21971_));
  NAND2_X1   g21905(.A1(new_n21970_), .A2(new_n21971_), .ZN(new_n21972_));
  XOR2_X1    g21906(.A1(new_n17770_), .A2(new_n21953_), .Z(new_n21973_));
  NAND2_X1   g21907(.A1(new_n21889_), .A2(new_n21973_), .ZN(new_n21974_));
  NAND3_X1   g21908(.A1(new_n21972_), .A2(new_n21974_), .A3(new_n21966_), .ZN(new_n21975_));
  NAND2_X1   g21909(.A1(new_n21975_), .A2(\a[5] ), .ZN(new_n21976_));
  NAND2_X1   g21910(.A1(new_n21976_), .A2(new_n21967_), .ZN(new_n21977_));
  AOI21_X1   g21911(.A1(new_n21885_), .A2(new_n21886_), .B(new_n21977_), .ZN(new_n21978_));
  NOR2_X1    g21912(.A1(new_n21876_), .A2(new_n21873_), .ZN(new_n21979_));
  NOR2_X1    g21913(.A1(new_n21869_), .A2(new_n21864_), .ZN(new_n21980_));
  NOR2_X1    g21914(.A1(new_n21979_), .A2(new_n21980_), .ZN(new_n21981_));
  INV_X1     g21915(.I(new_n21883_), .ZN(new_n21982_));
  NOR2_X1    g21916(.A1(new_n21981_), .A2(new_n21982_), .ZN(new_n21983_));
  NOR2_X1    g21917(.A1(new_n21975_), .A2(\a[5] ), .ZN(new_n21984_));
  AOI21_X1   g21918(.A1(new_n21963_), .A2(new_n21966_), .B(new_n65_), .ZN(new_n21985_));
  NOR2_X1    g21919(.A1(new_n21984_), .A2(new_n21985_), .ZN(new_n21986_));
  NOR3_X1    g21920(.A1(new_n21986_), .A2(new_n21884_), .A3(new_n21983_), .ZN(new_n21987_));
  NOR2_X1    g21921(.A1(new_n21978_), .A2(new_n21987_), .ZN(new_n21988_));
  XOR2_X1    g21922(.A1(new_n21747_), .A2(new_n21988_), .Z(new_n21989_));
  INV_X1     g21923(.I(new_n21989_), .ZN(new_n21990_));
  NAND2_X1   g21924(.A1(new_n21945_), .A2(new_n21947_), .ZN(new_n21991_));
  NOR2_X1    g21925(.A1(new_n21940_), .A2(new_n21894_), .ZN(new_n21992_));
  NOR2_X1    g21926(.A1(new_n21992_), .A2(new_n21941_), .ZN(new_n21993_));
  NAND2_X1   g21927(.A1(new_n21930_), .A2(new_n21928_), .ZN(new_n21994_));
  NAND2_X1   g21928(.A1(new_n21994_), .A2(new_n21931_), .ZN(new_n21995_));
  AOI21_X1   g21929(.A1(new_n11272_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n21996_));
  OAI21_X1   g21930(.A1(new_n2767_), .A2(new_n11277_), .B(new_n21996_), .ZN(new_n21997_));
  AOI21_X1   g21931(.A1(new_n11304_), .A2(new_n3332_), .B(new_n21997_), .ZN(new_n21998_));
  NAND2_X1   g21932(.A1(new_n11310_), .A2(new_n21998_), .ZN(new_n21999_));
  INV_X1     g21933(.I(new_n2596_), .ZN(new_n22000_));
  NAND4_X1   g21934(.A1(new_n1063_), .A2(new_n272_), .A3(new_n1572_), .A4(new_n250_), .ZN(new_n22001_));
  NOR3_X1    g21935(.A1(new_n2447_), .A2(new_n447_), .A3(new_n576_), .ZN(new_n22002_));
  NOR4_X1    g21936(.A1(new_n656_), .A2(new_n1865_), .A3(new_n345_), .A4(new_n518_), .ZN(new_n22003_));
  NAND4_X1   g21937(.A1(new_n22002_), .A2(new_n2630_), .A3(new_n22001_), .A4(new_n22003_), .ZN(new_n22004_));
  NOR3_X1    g21938(.A1(new_n22004_), .A2(new_n11043_), .A3(new_n2711_), .ZN(new_n22005_));
  AOI21_X1   g21939(.A1(new_n22000_), .A2(new_n22005_), .B(new_n21911_), .ZN(new_n22006_));
  NAND2_X1   g21940(.A1(new_n22000_), .A2(new_n22005_), .ZN(new_n22007_));
  NOR2_X1    g21941(.A1(new_n22007_), .A2(new_n21914_), .ZN(new_n22008_));
  NOR2_X1    g21942(.A1(new_n22008_), .A2(new_n22006_), .ZN(new_n22009_));
  NOR2_X1    g21943(.A1(new_n21999_), .A2(new_n22009_), .ZN(new_n22010_));
  INV_X1     g21944(.I(new_n21999_), .ZN(new_n22011_));
  XOR2_X1    g21945(.A1(new_n22007_), .A2(new_n21911_), .Z(new_n22012_));
  NOR2_X1    g21946(.A1(new_n22011_), .A2(new_n22012_), .ZN(new_n22013_));
  NOR2_X1    g21947(.A1(new_n22013_), .A2(new_n22010_), .ZN(new_n22014_));
  NOR2_X1    g21948(.A1(new_n21900_), .A2(new_n21917_), .ZN(new_n22015_));
  NOR2_X1    g21949(.A1(new_n22015_), .A2(new_n21915_), .ZN(new_n22016_));
  XNOR2_X1   g21950(.A1(new_n22014_), .A2(new_n22016_), .ZN(new_n22017_));
  INV_X1     g21951(.I(new_n22017_), .ZN(new_n22018_));
  NAND2_X1   g21952(.A1(new_n22014_), .A2(new_n22016_), .ZN(new_n22019_));
  NOR2_X1    g21953(.A1(new_n22014_), .A2(new_n22016_), .ZN(new_n22020_));
  INV_X1     g21954(.I(new_n22020_), .ZN(new_n22021_));
  AOI21_X1   g21955(.A1(new_n22019_), .A2(new_n22021_), .B(new_n21995_), .ZN(new_n22022_));
  AOI21_X1   g21956(.A1(new_n21995_), .A2(new_n22018_), .B(new_n22022_), .ZN(new_n22023_));
  INV_X1     g21957(.I(new_n22023_), .ZN(new_n22024_));
  NAND2_X1   g21958(.A1(new_n3318_), .A2(new_n3322_), .ZN(new_n22025_));
  AND3_X2    g21959(.A1(new_n11463_), .A2(new_n3267_), .A3(new_n22025_), .Z(new_n22026_));
  NOR4_X1    g21960(.A1(new_n11468_), .A2(new_n3260_), .A3(new_n11461_), .A4(new_n22026_), .ZN(new_n22027_));
  XOR2_X1    g21961(.A1(new_n22027_), .A2(new_n72_), .Z(new_n22028_));
  OAI22_X1   g21962(.A1(new_n11353_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n11345_), .ZN(new_n22029_));
  NAND2_X1   g21963(.A1(new_n11370_), .A2(new_n2750_), .ZN(new_n22030_));
  AOI21_X1   g21964(.A1(new_n22030_), .A2(new_n22029_), .B(new_n2737_), .ZN(new_n22031_));
  NAND2_X1   g21965(.A1(new_n11379_), .A2(new_n22031_), .ZN(new_n22032_));
  XOR2_X1    g21966(.A1(new_n22032_), .A2(\a[29] ), .Z(new_n22033_));
  AND2_X2    g21967(.A1(new_n22028_), .A2(new_n22033_), .Z(new_n22034_));
  NOR2_X1    g21968(.A1(new_n22028_), .A2(new_n22033_), .ZN(new_n22035_));
  OAI21_X1   g21969(.A1(new_n22034_), .A2(new_n22035_), .B(new_n22024_), .ZN(new_n22036_));
  XNOR2_X1   g21970(.A1(new_n22028_), .A2(new_n22033_), .ZN(new_n22037_));
  OAI21_X1   g21971(.A1(new_n22024_), .A2(new_n22037_), .B(new_n22036_), .ZN(new_n22038_));
  XNOR2_X1   g21972(.A1(new_n22038_), .A2(new_n21993_), .ZN(new_n22039_));
  NAND3_X1   g21973(.A1(new_n21892_), .A2(new_n21890_), .A3(new_n21948_), .ZN(new_n22040_));
  NAND3_X1   g21974(.A1(new_n22040_), .A2(new_n21991_), .A3(new_n22039_), .ZN(new_n22041_));
  INV_X1     g21975(.I(new_n22039_), .ZN(new_n22042_));
  INV_X1     g21976(.I(new_n17758_), .ZN(new_n22043_));
  NAND2_X1   g21977(.A1(new_n21891_), .A2(new_n17760_), .ZN(new_n22044_));
  OAI21_X1   g21978(.A1(new_n22043_), .A2(new_n22044_), .B(new_n21890_), .ZN(new_n22045_));
  OAI21_X1   g21979(.A1(new_n22045_), .A2(new_n21949_), .B(new_n21991_), .ZN(new_n22046_));
  NAND2_X1   g21980(.A1(new_n22046_), .A2(new_n22042_), .ZN(new_n22047_));
  NAND2_X1   g21981(.A1(new_n22047_), .A2(new_n22041_), .ZN(new_n22048_));
  NOR2_X1    g21982(.A1(new_n22046_), .A2(new_n22042_), .ZN(new_n22049_));
  AOI21_X1   g21983(.A1(new_n22040_), .A2(new_n21991_), .B(new_n22039_), .ZN(new_n22050_));
  NOR2_X1    g21984(.A1(new_n22049_), .A2(new_n22050_), .ZN(new_n22051_));
  OAI21_X1   g21985(.A1(new_n22051_), .A2(new_n19512_), .B(new_n21960_), .ZN(new_n22052_));
  NAND3_X1   g21986(.A1(new_n21968_), .A2(new_n22052_), .A3(new_n21969_), .ZN(new_n22053_));
  AOI21_X1   g21987(.A1(new_n22051_), .A2(new_n19512_), .B(new_n21960_), .ZN(new_n22054_));
  INV_X1     g21988(.I(new_n22054_), .ZN(new_n22055_));
  AOI21_X1   g21989(.A1(new_n22053_), .A2(new_n22055_), .B(new_n22048_), .ZN(new_n22056_));
  NAND2_X1   g21990(.A1(new_n21995_), .A2(new_n22019_), .ZN(new_n22057_));
  NAND2_X1   g21991(.A1(new_n22057_), .A2(new_n22021_), .ZN(new_n22058_));
  INV_X1     g21992(.I(new_n22058_), .ZN(new_n22059_));
  OAI22_X1   g21993(.A1(new_n11353_), .A2(new_n2747_), .B1(new_n3175_), .B2(new_n11697_), .ZN(new_n22060_));
  NAND2_X1   g21994(.A1(new_n11370_), .A2(new_n3275_), .ZN(new_n22061_));
  AOI21_X1   g21995(.A1(new_n22061_), .A2(new_n22060_), .B(new_n2737_), .ZN(new_n22062_));
  NAND2_X1   g21996(.A1(new_n11700_), .A2(new_n22062_), .ZN(new_n22063_));
  XOR2_X1    g21997(.A1(new_n22063_), .A2(\a[29] ), .Z(new_n22064_));
  INV_X1     g21998(.I(new_n22006_), .ZN(new_n22065_));
  AOI21_X1   g21999(.A1(new_n22011_), .A2(new_n22065_), .B(new_n22008_), .ZN(new_n22066_));
  NAND2_X1   g22000(.A1(new_n11304_), .A2(new_n3189_), .ZN(new_n22067_));
  NAND2_X1   g22001(.A1(new_n11346_), .A2(new_n3332_), .ZN(new_n22068_));
  AOI21_X1   g22002(.A1(new_n11311_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n22069_));
  NAND4_X1   g22003(.A1(new_n11757_), .A2(new_n22067_), .A3(new_n22068_), .A4(new_n22069_), .ZN(new_n22070_));
  NOR3_X1    g22004(.A1(new_n22025_), .A2(new_n3259_), .A3(new_n3267_), .ZN(new_n22071_));
  NOR3_X1    g22005(.A1(new_n11461_), .A2(new_n72_), .A3(new_n22071_), .ZN(new_n22072_));
  OAI21_X1   g22006(.A1(new_n11461_), .A2(new_n22071_), .B(new_n72_), .ZN(new_n22073_));
  INV_X1     g22007(.I(new_n22073_), .ZN(new_n22074_));
  NOR2_X1    g22008(.A1(new_n22074_), .A2(new_n22072_), .ZN(new_n22075_));
  INV_X1     g22009(.I(new_n3134_), .ZN(new_n22076_));
  NOR2_X1    g22010(.A1(new_n3165_), .A2(new_n22076_), .ZN(new_n22077_));
  NOR3_X1    g22011(.A1(new_n2338_), .A2(new_n630_), .A3(new_n1168_), .ZN(new_n22078_));
  AND3_X2    g22012(.A1(new_n2706_), .A2(new_n2686_), .A3(new_n22078_), .Z(new_n22079_));
  AOI21_X1   g22013(.A1(new_n22077_), .A2(new_n22079_), .B(new_n21914_), .ZN(new_n22080_));
  NAND2_X1   g22014(.A1(new_n22079_), .A2(new_n22077_), .ZN(new_n22081_));
  NOR2_X1    g22015(.A1(new_n22081_), .A2(new_n21911_), .ZN(new_n22082_));
  NOR2_X1    g22016(.A1(new_n22082_), .A2(new_n22080_), .ZN(new_n22083_));
  NOR2_X1    g22017(.A1(new_n22075_), .A2(new_n22083_), .ZN(new_n22084_));
  XOR2_X1    g22018(.A1(new_n22081_), .A2(new_n21914_), .Z(new_n22085_));
  INV_X1     g22019(.I(new_n22085_), .ZN(new_n22086_));
  AOI21_X1   g22020(.A1(new_n22075_), .A2(new_n22086_), .B(new_n22084_), .ZN(new_n22087_));
  INV_X1     g22021(.I(new_n22087_), .ZN(new_n22088_));
  NOR2_X1    g22022(.A1(new_n22070_), .A2(new_n22088_), .ZN(new_n22089_));
  INV_X1     g22023(.I(new_n22089_), .ZN(new_n22090_));
  NAND2_X1   g22024(.A1(new_n22070_), .A2(new_n22088_), .ZN(new_n22091_));
  AOI21_X1   g22025(.A1(new_n22090_), .A2(new_n22091_), .B(new_n22066_), .ZN(new_n22092_));
  INV_X1     g22026(.I(new_n22066_), .ZN(new_n22093_));
  XOR2_X1    g22027(.A1(new_n22070_), .A2(new_n22087_), .Z(new_n22094_));
  NOR2_X1    g22028(.A1(new_n22093_), .A2(new_n22094_), .ZN(new_n22095_));
  NOR2_X1    g22029(.A1(new_n22095_), .A2(new_n22092_), .ZN(new_n22096_));
  XNOR2_X1   g22030(.A1(new_n22064_), .A2(new_n22096_), .ZN(new_n22097_));
  NOR2_X1    g22031(.A1(new_n22059_), .A2(new_n22097_), .ZN(new_n22098_));
  NAND2_X1   g22032(.A1(new_n22064_), .A2(new_n22096_), .ZN(new_n22099_));
  NOR2_X1    g22033(.A1(new_n22064_), .A2(new_n22096_), .ZN(new_n22100_));
  INV_X1     g22034(.I(new_n22100_), .ZN(new_n22101_));
  NAND2_X1   g22035(.A1(new_n22101_), .A2(new_n22099_), .ZN(new_n22102_));
  AOI21_X1   g22036(.A1(new_n22059_), .A2(new_n22102_), .B(new_n22098_), .ZN(new_n22103_));
  NAND2_X1   g22037(.A1(new_n22038_), .A2(new_n21993_), .ZN(new_n22104_));
  NOR2_X1    g22038(.A1(new_n22024_), .A2(new_n22034_), .ZN(new_n22105_));
  NOR2_X1    g22039(.A1(new_n22105_), .A2(new_n22035_), .ZN(new_n22106_));
  INV_X1     g22040(.I(new_n22106_), .ZN(new_n22107_));
  AOI21_X1   g22041(.A1(new_n22041_), .A2(new_n22104_), .B(new_n22107_), .ZN(new_n22108_));
  NAND3_X1   g22042(.A1(new_n22041_), .A2(new_n22104_), .A3(new_n22107_), .ZN(new_n22109_));
  INV_X1     g22043(.I(new_n22109_), .ZN(new_n22110_));
  OAI21_X1   g22044(.A1(new_n22110_), .A2(new_n22108_), .B(new_n22103_), .ZN(new_n22111_));
  INV_X1     g22045(.I(new_n22103_), .ZN(new_n22112_));
  INV_X1     g22046(.I(new_n22108_), .ZN(new_n22113_));
  NAND3_X1   g22047(.A1(new_n22113_), .A2(new_n22112_), .A3(new_n22109_), .ZN(new_n22114_));
  AND2_X2    g22048(.A1(new_n22114_), .A2(new_n22111_), .Z(new_n22115_));
  NAND3_X1   g22049(.A1(new_n22053_), .A2(new_n22048_), .A3(new_n22055_), .ZN(new_n22116_));
  AOI21_X1   g22050(.A1(new_n22115_), .A2(new_n22116_), .B(new_n22056_), .ZN(new_n22117_));
  NAND2_X1   g22051(.A1(new_n22114_), .A2(new_n22111_), .ZN(new_n22118_));
  AOI21_X1   g22052(.A1(new_n22058_), .A2(new_n22099_), .B(new_n22100_), .ZN(new_n22119_));
  OAI22_X1   g22053(.A1(new_n11369_), .A2(new_n2747_), .B1(new_n3175_), .B2(new_n11461_), .ZN(new_n22120_));
  NAND2_X1   g22054(.A1(new_n11694_), .A2(new_n3275_), .ZN(new_n22121_));
  AOI21_X1   g22055(.A1(new_n22120_), .A2(new_n22121_), .B(new_n2737_), .ZN(new_n22122_));
  NAND2_X1   g22056(.A1(new_n12720_), .A2(new_n22122_), .ZN(new_n22123_));
  XOR2_X1    g22057(.A1(new_n22123_), .A2(new_n74_), .Z(new_n22124_));
  AOI21_X1   g22058(.A1(new_n11346_), .A2(new_n3189_), .B(new_n2763_), .ZN(new_n22125_));
  OAI21_X1   g22059(.A1(new_n2771_), .A2(new_n11264_), .B(new_n22125_), .ZN(new_n22126_));
  AOI21_X1   g22060(.A1(new_n11354_), .A2(new_n3332_), .B(new_n22126_), .ZN(new_n22127_));
  NAND2_X1   g22061(.A1(new_n11678_), .A2(new_n22127_), .ZN(new_n22128_));
  NOR3_X1    g22062(.A1(new_n22074_), .A2(new_n22072_), .A3(new_n22080_), .ZN(new_n22129_));
  NAND4_X1   g22063(.A1(new_n22077_), .A2(new_n832_), .A3(new_n2693_), .A4(new_n3133_), .ZN(new_n22130_));
  OAI21_X1   g22064(.A1(new_n22129_), .A2(new_n22082_), .B(new_n22130_), .ZN(new_n22131_));
  NOR2_X1    g22065(.A1(new_n22129_), .A2(new_n22082_), .ZN(new_n22132_));
  INV_X1     g22066(.I(new_n22130_), .ZN(new_n22133_));
  NAND2_X1   g22067(.A1(new_n22132_), .A2(new_n22133_), .ZN(new_n22134_));
  AOI21_X1   g22068(.A1(new_n22131_), .A2(new_n22134_), .B(new_n22128_), .ZN(new_n22135_));
  INV_X1     g22069(.I(new_n22128_), .ZN(new_n22136_));
  XOR2_X1    g22070(.A1(new_n22132_), .A2(new_n22130_), .Z(new_n22137_));
  NOR2_X1    g22071(.A1(new_n22136_), .A2(new_n22137_), .ZN(new_n22138_));
  NOR2_X1    g22072(.A1(new_n22138_), .A2(new_n22135_), .ZN(new_n22139_));
  AOI21_X1   g22073(.A1(new_n22093_), .A2(new_n22091_), .B(new_n22089_), .ZN(new_n22140_));
  XOR2_X1    g22074(.A1(new_n22139_), .A2(new_n22140_), .Z(new_n22141_));
  NAND2_X1   g22075(.A1(new_n22139_), .A2(new_n22140_), .ZN(new_n22142_));
  NOR2_X1    g22076(.A1(new_n22139_), .A2(new_n22140_), .ZN(new_n22143_));
  INV_X1     g22077(.I(new_n22143_), .ZN(new_n22144_));
  NAND2_X1   g22078(.A1(new_n22144_), .A2(new_n22142_), .ZN(new_n22145_));
  MUX2_X1    g22079(.I0(new_n22145_), .I1(new_n22141_), .S(new_n22124_), .Z(new_n22146_));
  NOR2_X1    g22080(.A1(new_n22119_), .A2(new_n22146_), .ZN(new_n22147_));
  AND2_X2    g22081(.A1(new_n22119_), .A2(new_n22146_), .Z(new_n22148_));
  NOR2_X1    g22082(.A1(new_n22148_), .A2(new_n22147_), .ZN(new_n22149_));
  INV_X1     g22083(.I(new_n22149_), .ZN(new_n22150_));
  NOR2_X1    g22084(.A1(new_n22118_), .A2(new_n22150_), .ZN(new_n22151_));
  INV_X1     g22085(.I(new_n22151_), .ZN(new_n22152_));
  NAND2_X1   g22086(.A1(new_n22118_), .A2(new_n22150_), .ZN(new_n22153_));
  AOI21_X1   g22087(.A1(new_n22152_), .A2(new_n22153_), .B(new_n22117_), .ZN(new_n22154_));
  AOI21_X1   g22088(.A1(new_n22048_), .A2(new_n17770_), .B(new_n21953_), .ZN(new_n22155_));
  NOR3_X1    g22089(.A1(new_n21958_), .A2(new_n22155_), .A3(new_n21888_), .ZN(new_n22156_));
  OAI21_X1   g22090(.A1(new_n22156_), .A2(new_n22054_), .B(new_n22051_), .ZN(new_n22157_));
  NOR3_X1    g22091(.A1(new_n22156_), .A2(new_n22051_), .A3(new_n22054_), .ZN(new_n22158_));
  OAI21_X1   g22092(.A1(new_n22118_), .A2(new_n22158_), .B(new_n22157_), .ZN(new_n22159_));
  NAND2_X1   g22093(.A1(new_n22115_), .A2(new_n22150_), .ZN(new_n22160_));
  NAND2_X1   g22094(.A1(new_n22118_), .A2(new_n22149_), .ZN(new_n22161_));
  AOI21_X1   g22095(.A1(new_n22160_), .A2(new_n22161_), .B(new_n22159_), .ZN(new_n22162_));
  NOR2_X1    g22096(.A1(new_n22154_), .A2(new_n22162_), .ZN(new_n22163_));
  OAI22_X1   g22097(.A1(new_n22115_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n22051_), .ZN(new_n22164_));
  NAND2_X1   g22098(.A1(new_n22150_), .A2(new_n9488_), .ZN(new_n22165_));
  AOI21_X1   g22099(.A1(new_n22164_), .A2(new_n22165_), .B(new_n9482_), .ZN(new_n22166_));
  NAND2_X1   g22100(.A1(new_n22163_), .A2(new_n22166_), .ZN(new_n22167_));
  XOR2_X1    g22101(.A1(new_n22167_), .A2(\a[2] ), .Z(new_n22168_));
  NOR2_X1    g22102(.A1(new_n21889_), .A2(new_n21953_), .ZN(new_n22169_));
  NOR3_X1    g22103(.A1(new_n21958_), .A2(new_n21888_), .A3(new_n21960_), .ZN(new_n22170_));
  NOR4_X1    g22104(.A1(new_n22169_), .A2(new_n22170_), .A3(new_n21961_), .A4(new_n22048_), .ZN(new_n22171_));
  OAI21_X1   g22105(.A1(new_n21958_), .A2(new_n21888_), .B(new_n21960_), .ZN(new_n22172_));
  AOI21_X1   g22106(.A1(new_n21889_), .A2(new_n21953_), .B(new_n21961_), .ZN(new_n22173_));
  AOI21_X1   g22107(.A1(new_n22173_), .A2(new_n22172_), .B(new_n22051_), .ZN(new_n22174_));
  NOR2_X1    g22108(.A1(new_n22174_), .A2(new_n22171_), .ZN(new_n22175_));
  OAI22_X1   g22109(.A1(new_n19512_), .A2(new_n9485_), .B1(new_n21960_), .B2(new_n9483_), .ZN(new_n22176_));
  NAND2_X1   g22110(.A1(new_n22048_), .A2(new_n9488_), .ZN(new_n22177_));
  AOI21_X1   g22111(.A1(new_n22177_), .A2(new_n22176_), .B(new_n9482_), .ZN(new_n22178_));
  NAND2_X1   g22112(.A1(new_n22175_), .A2(new_n22178_), .ZN(new_n22179_));
  XOR2_X1    g22113(.A1(new_n22179_), .A2(\a[2] ), .Z(new_n22180_));
  INV_X1     g22114(.I(new_n22180_), .ZN(new_n22181_));
  NOR2_X1    g22115(.A1(new_n21148_), .A2(new_n21149_), .ZN(new_n22182_));
  NOR2_X1    g22116(.A1(new_n21160_), .A2(new_n21161_), .ZN(new_n22183_));
  NOR2_X1    g22117(.A1(new_n22182_), .A2(new_n22183_), .ZN(new_n22184_));
  NOR2_X1    g22118(.A1(new_n22184_), .A2(new_n21162_), .ZN(new_n22185_));
  NOR3_X1    g22119(.A1(new_n21224_), .A2(new_n21225_), .A3(new_n21226_), .ZN(new_n22186_));
  AOI21_X1   g22120(.A1(new_n21216_), .A2(new_n21220_), .B(new_n21197_), .ZN(new_n22187_));
  NOR2_X1    g22121(.A1(new_n22187_), .A2(new_n22186_), .ZN(new_n22188_));
  NAND2_X1   g22122(.A1(new_n21594_), .A2(new_n21586_), .ZN(new_n22189_));
  NAND2_X1   g22123(.A1(new_n21611_), .A2(new_n21606_), .ZN(new_n22190_));
  NAND2_X1   g22124(.A1(new_n22189_), .A2(new_n22190_), .ZN(new_n22191_));
  INV_X1     g22125(.I(new_n21613_), .ZN(new_n22192_));
  NOR3_X1    g22126(.A1(new_n21621_), .A2(\a[5] ), .A3(new_n21622_), .ZN(new_n22193_));
  AOI21_X1   g22127(.A1(new_n20907_), .A2(new_n21617_), .B(new_n65_), .ZN(new_n22194_));
  NOR2_X1    g22128(.A1(new_n22194_), .A2(new_n22193_), .ZN(new_n22195_));
  AOI21_X1   g22129(.A1(new_n22191_), .A2(new_n22192_), .B(new_n22195_), .ZN(new_n22196_));
  AOI21_X1   g22130(.A1(new_n21690_), .A2(new_n21691_), .B(new_n21689_), .ZN(new_n22197_));
  NOR3_X1    g22131(.A1(new_n21685_), .A2(new_n21682_), .A3(new_n21673_), .ZN(new_n22198_));
  NOR2_X1    g22132(.A1(new_n22198_), .A2(new_n22197_), .ZN(new_n22199_));
  NAND3_X1   g22133(.A1(new_n22191_), .A2(new_n22195_), .A3(new_n22192_), .ZN(new_n22200_));
  AOI21_X1   g22134(.A1(new_n22199_), .A2(new_n22200_), .B(new_n22196_), .ZN(new_n22201_));
  AOI21_X1   g22135(.A1(new_n22201_), .A2(new_n21242_), .B(new_n21240_), .ZN(new_n22202_));
  AOI21_X1   g22136(.A1(new_n22202_), .A2(new_n22188_), .B(new_n21697_), .ZN(new_n22203_));
  OAI21_X1   g22137(.A1(new_n21726_), .A2(new_n21727_), .B(new_n21725_), .ZN(new_n22204_));
  NAND3_X1   g22138(.A1(new_n21721_), .A2(new_n21708_), .A3(new_n21718_), .ZN(new_n22205_));
  NOR2_X1    g22139(.A1(new_n21734_), .A2(\a[5] ), .ZN(new_n22206_));
  AOI21_X1   g22140(.A1(new_n21088_), .A2(new_n21733_), .B(new_n65_), .ZN(new_n22207_));
  NOR2_X1    g22141(.A1(new_n22207_), .A2(new_n22206_), .ZN(new_n22208_));
  NAND3_X1   g22142(.A1(new_n22204_), .A2(new_n22205_), .A3(new_n22208_), .ZN(new_n22209_));
  AOI21_X1   g22143(.A1(new_n22204_), .A2(new_n22205_), .B(new_n22208_), .ZN(new_n22210_));
  AOI21_X1   g22144(.A1(new_n22203_), .A2(new_n22209_), .B(new_n22210_), .ZN(new_n22211_));
  NOR2_X1    g22145(.A1(new_n21184_), .A2(new_n21744_), .ZN(new_n22212_));
  AOI21_X1   g22146(.A1(new_n22211_), .A2(new_n22212_), .B(new_n21184_), .ZN(new_n22213_));
  XOR2_X1    g22147(.A1(new_n22185_), .A2(new_n22213_), .Z(new_n22214_));
  NAND2_X1   g22148(.A1(new_n21157_), .A2(new_n9488_), .ZN(new_n22215_));
  NAND2_X1   g22149(.A1(new_n19484_), .A2(new_n9503_), .ZN(new_n22216_));
  AOI21_X1   g22150(.A1(new_n17780_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n22217_));
  NAND4_X1   g22151(.A1(new_n21155_), .A2(new_n22215_), .A3(new_n22216_), .A4(new_n22217_), .ZN(new_n22218_));
  XOR2_X1    g22152(.A1(new_n22218_), .A2(\a[2] ), .Z(new_n22219_));
  INV_X1     g22153(.I(new_n22219_), .ZN(new_n22220_));
  NAND2_X1   g22154(.A1(new_n19438_), .A2(new_n9488_), .ZN(new_n22221_));
  NAND2_X1   g22155(.A1(new_n20896_), .A2(new_n9503_), .ZN(new_n22222_));
  AOI21_X1   g22156(.A1(new_n19442_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n22223_));
  NAND4_X1   g22157(.A1(new_n21621_), .A2(new_n22221_), .A3(new_n22222_), .A4(new_n22223_), .ZN(new_n22224_));
  XOR2_X1    g22158(.A1(new_n22224_), .A2(\a[2] ), .Z(new_n22225_));
  OR2_X2     g22159(.A1(new_n20915_), .A2(new_n20918_), .Z(new_n22226_));
  NAND2_X1   g22160(.A1(new_n20896_), .A2(new_n9488_), .ZN(new_n22227_));
  NAND2_X1   g22161(.A1(new_n19442_), .A2(new_n9503_), .ZN(new_n22228_));
  AOI21_X1   g22162(.A1(new_n19439_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n22229_));
  NAND4_X1   g22163(.A1(new_n22226_), .A2(new_n22227_), .A3(new_n22228_), .A4(new_n22229_), .ZN(new_n22230_));
  XOR2_X1    g22164(.A1(new_n22230_), .A2(\a[2] ), .Z(new_n22231_));
  INV_X1     g22165(.I(new_n22231_), .ZN(new_n22232_));
  OAI22_X1   g22166(.A1(new_n19410_), .A2(new_n9485_), .B1(new_n19412_), .B2(new_n9483_), .ZN(new_n22233_));
  OAI21_X1   g22167(.A1(new_n17787_), .A2(new_n9489_), .B(new_n22233_), .ZN(new_n22234_));
  AOI21_X1   g22168(.A1(new_n20827_), .A2(new_n6922_), .B(new_n22234_), .ZN(new_n22235_));
  XOR2_X1    g22169(.A1(new_n22235_), .A2(\a[2] ), .Z(new_n22236_));
  INV_X1     g22170(.I(new_n22236_), .ZN(new_n22237_));
  INV_X1     g22171(.I(new_n19951_), .ZN(new_n22238_));
  AOI22_X1   g22172(.A1(new_n19359_), .A2(new_n7530_), .B1(new_n6789_), .B2(new_n19365_), .ZN(new_n22239_));
  AOI21_X1   g22173(.A1(new_n6784_), .A2(new_n17802_), .B(new_n22239_), .ZN(new_n22240_));
  OR3_X2     g22174(.A1(new_n22238_), .A2(new_n6776_), .A3(new_n22240_), .Z(new_n22241_));
  XOR2_X1    g22175(.A1(new_n22241_), .A2(\a[8] ), .Z(new_n22242_));
  INV_X1     g22176(.I(new_n22242_), .ZN(new_n22243_));
  INV_X1     g22177(.I(new_n19550_), .ZN(new_n22244_));
  NOR2_X1    g22178(.A1(new_n22244_), .A2(new_n19551_), .ZN(new_n22245_));
  AOI22_X1   g22179(.A1(new_n19308_), .A2(new_n6180_), .B1(new_n6095_), .B2(new_n19545_), .ZN(new_n22246_));
  AOI21_X1   g22180(.A1(new_n6090_), .A2(new_n17850_), .B(new_n22246_), .ZN(new_n22247_));
  OR3_X2     g22181(.A1(new_n22245_), .A2(new_n6082_), .A3(new_n22247_), .Z(new_n22248_));
  XOR2_X1    g22182(.A1(new_n22248_), .A2(\a[14] ), .Z(new_n22249_));
  NOR2_X1    g22183(.A1(new_n22249_), .A2(new_n21283_), .ZN(new_n22250_));
  INV_X1     g22184(.I(new_n22250_), .ZN(new_n22251_));
  AOI22_X1   g22185(.A1(new_n19290_), .A2(new_n6180_), .B1(new_n6095_), .B2(new_n19308_), .ZN(new_n22252_));
  AOI21_X1   g22186(.A1(new_n6090_), .A2(new_n19545_), .B(new_n22252_), .ZN(new_n22253_));
  NOR3_X1    g22187(.A1(new_n22253_), .A2(new_n19571_), .A3(new_n6082_), .ZN(new_n22254_));
  XOR2_X1    g22188(.A1(new_n22254_), .A2(new_n3521_), .Z(new_n22255_));
  NOR2_X1    g22189(.A1(new_n6079_), .A2(new_n6080_), .ZN(new_n22256_));
  OAI21_X1   g22190(.A1(new_n19313_), .A2(new_n6094_), .B(new_n22256_), .ZN(new_n22257_));
  NOR2_X1    g22191(.A1(new_n19593_), .A2(new_n22257_), .ZN(new_n22258_));
  XOR2_X1    g22192(.A1(new_n22258_), .A2(new_n3521_), .Z(new_n22259_));
  NOR2_X1    g22193(.A1(new_n19313_), .A2(new_n6079_), .ZN(new_n22260_));
  NOR2_X1    g22194(.A1(new_n22260_), .A2(new_n3521_), .ZN(new_n22261_));
  NAND2_X1   g22195(.A1(new_n22259_), .A2(new_n22261_), .ZN(new_n22262_));
  NOR2_X1    g22196(.A1(new_n22255_), .A2(new_n22262_), .ZN(new_n22263_));
  AND2_X2    g22197(.A1(new_n22249_), .A2(new_n21283_), .Z(new_n22264_));
  OAI21_X1   g22198(.A1(new_n22263_), .A2(new_n22264_), .B(new_n22251_), .ZN(new_n22265_));
  NOR2_X1    g22199(.A1(new_n21283_), .A2(new_n3372_), .ZN(new_n22266_));
  XOR2_X1    g22200(.A1(new_n21377_), .A2(new_n22266_), .Z(new_n22267_));
  AOI22_X1   g22201(.A1(new_n17850_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n19545_), .ZN(new_n22268_));
  AOI21_X1   g22202(.A1(new_n19305_), .A2(new_n6090_), .B(new_n22268_), .ZN(new_n22269_));
  NOR3_X1    g22203(.A1(new_n19618_), .A2(new_n6082_), .A3(new_n22269_), .ZN(new_n22270_));
  XOR2_X1    g22204(.A1(new_n22270_), .A2(\a[14] ), .Z(new_n22271_));
  OR2_X2     g22205(.A1(new_n22271_), .A2(new_n22267_), .Z(new_n22272_));
  NAND2_X1   g22206(.A1(new_n22265_), .A2(new_n22272_), .ZN(new_n22273_));
  NAND2_X1   g22207(.A1(new_n22271_), .A2(new_n22267_), .ZN(new_n22274_));
  NAND2_X1   g22208(.A1(new_n22273_), .A2(new_n22274_), .ZN(new_n22275_));
  INV_X1     g22209(.I(new_n22275_), .ZN(new_n22276_));
  INV_X1     g22210(.I(new_n19647_), .ZN(new_n22277_));
  AOI22_X1   g22211(.A1(new_n19305_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n17850_), .ZN(new_n22278_));
  AOI21_X1   g22212(.A1(new_n6090_), .A2(new_n19321_), .B(new_n22278_), .ZN(new_n22279_));
  OR3_X2     g22213(.A1(new_n22277_), .A2(new_n6082_), .A3(new_n22279_), .Z(new_n22280_));
  XOR2_X1    g22214(.A1(new_n22280_), .A2(\a[14] ), .Z(new_n22281_));
  NOR2_X1    g22215(.A1(new_n22276_), .A2(new_n22281_), .ZN(new_n22282_));
  XOR2_X1    g22216(.A1(new_n21278_), .A2(\a[17] ), .Z(new_n22283_));
  INV_X1     g22217(.I(new_n21377_), .ZN(new_n22284_));
  NAND2_X1   g22218(.A1(new_n22284_), .A2(new_n22266_), .ZN(new_n22285_));
  INV_X1     g22219(.I(new_n22285_), .ZN(new_n22286_));
  NOR2_X1    g22220(.A1(new_n22286_), .A2(new_n22283_), .ZN(new_n22287_));
  NOR2_X1    g22221(.A1(new_n22287_), .A2(new_n21378_), .ZN(new_n22288_));
  AOI21_X1   g22222(.A1(new_n22276_), .A2(new_n22281_), .B(new_n22288_), .ZN(new_n22289_));
  NOR2_X1    g22223(.A1(new_n22289_), .A2(new_n22282_), .ZN(new_n22290_));
  NOR2_X1    g22224(.A1(new_n21375_), .A2(new_n21271_), .ZN(new_n22291_));
  XOR2_X1    g22225(.A1(new_n22291_), .A2(new_n21374_), .Z(new_n22292_));
  NOR2_X1    g22226(.A1(new_n22292_), .A2(new_n21285_), .ZN(new_n22293_));
  NOR2_X1    g22227(.A1(new_n21274_), .A2(new_n21379_), .ZN(new_n22294_));
  NOR2_X1    g22228(.A1(new_n22294_), .A2(new_n21378_), .ZN(new_n22295_));
  NOR2_X1    g22229(.A1(new_n22293_), .A2(new_n22295_), .ZN(new_n22296_));
  OR2_X2     g22230(.A1(new_n19679_), .A2(new_n19682_), .Z(new_n22297_));
  INV_X1     g22231(.I(new_n22297_), .ZN(new_n22298_));
  AOI22_X1   g22232(.A1(new_n19305_), .A2(new_n6180_), .B1(new_n6095_), .B2(new_n19321_), .ZN(new_n22299_));
  AOI21_X1   g22233(.A1(new_n6090_), .A2(new_n17827_), .B(new_n22299_), .ZN(new_n22300_));
  NOR3_X1    g22234(.A1(new_n22298_), .A2(new_n6082_), .A3(new_n22300_), .ZN(new_n22301_));
  XOR2_X1    g22235(.A1(new_n22301_), .A2(new_n3521_), .Z(new_n22302_));
  XNOR2_X1   g22236(.A1(new_n22302_), .A2(new_n22296_), .ZN(new_n22303_));
  NOR2_X1    g22237(.A1(new_n22290_), .A2(new_n22303_), .ZN(new_n22304_));
  NAND2_X1   g22238(.A1(new_n22302_), .A2(new_n22296_), .ZN(new_n22305_));
  NOR2_X1    g22239(.A1(new_n22302_), .A2(new_n22296_), .ZN(new_n22306_));
  INV_X1     g22240(.I(new_n22306_), .ZN(new_n22307_));
  NAND2_X1   g22241(.A1(new_n22307_), .A2(new_n22305_), .ZN(new_n22308_));
  AOI21_X1   g22242(.A1(new_n22290_), .A2(new_n22308_), .B(new_n22304_), .ZN(new_n22309_));
  NOR2_X1    g22243(.A1(new_n22275_), .A2(new_n22281_), .ZN(new_n22310_));
  INV_X1     g22244(.I(new_n22310_), .ZN(new_n22311_));
  NAND2_X1   g22245(.A1(new_n22275_), .A2(new_n22281_), .ZN(new_n22312_));
  AOI21_X1   g22246(.A1(new_n22311_), .A2(new_n22312_), .B(new_n22286_), .ZN(new_n22313_));
  INV_X1     g22247(.I(new_n22312_), .ZN(new_n22314_));
  NOR3_X1    g22248(.A1(new_n22314_), .A2(new_n22285_), .A3(new_n22310_), .ZN(new_n22315_));
  OAI21_X1   g22249(.A1(new_n22313_), .A2(new_n22315_), .B(new_n22283_), .ZN(new_n22316_));
  INV_X1     g22250(.I(new_n22283_), .ZN(new_n22317_));
  OAI21_X1   g22251(.A1(new_n22314_), .A2(new_n22310_), .B(new_n22285_), .ZN(new_n22318_));
  NAND3_X1   g22252(.A1(new_n22311_), .A2(new_n22286_), .A3(new_n22312_), .ZN(new_n22319_));
  NAND3_X1   g22253(.A1(new_n22318_), .A2(new_n22319_), .A3(new_n22317_), .ZN(new_n22320_));
  OAI22_X1   g22254(.A1(new_n4719_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n4716_), .ZN(new_n22321_));
  NAND2_X1   g22255(.A1(new_n19350_), .A2(new_n4709_), .ZN(new_n22322_));
  AOI21_X1   g22256(.A1(new_n22321_), .A2(new_n22322_), .B(new_n4707_), .ZN(new_n22323_));
  NAND2_X1   g22257(.A1(new_n20535_), .A2(new_n22323_), .ZN(new_n22324_));
  XOR2_X1    g22258(.A1(new_n22324_), .A2(\a[11] ), .Z(new_n22325_));
  INV_X1     g22259(.I(new_n22325_), .ZN(new_n22326_));
  AOI21_X1   g22260(.A1(new_n22316_), .A2(new_n22320_), .B(new_n22326_), .ZN(new_n22327_));
  INV_X1     g22261(.I(new_n22260_), .ZN(new_n22328_));
  AOI22_X1   g22262(.A1(new_n19308_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n19545_), .ZN(new_n22329_));
  AOI21_X1   g22263(.A1(new_n4709_), .A2(new_n17850_), .B(new_n22329_), .ZN(new_n22330_));
  OR3_X2     g22264(.A1(new_n22245_), .A2(new_n4707_), .A3(new_n22330_), .Z(new_n22331_));
  XOR2_X1    g22265(.A1(new_n22331_), .A2(new_n4034_), .Z(new_n22332_));
  NAND2_X1   g22266(.A1(new_n22332_), .A2(new_n22328_), .ZN(new_n22333_));
  AOI22_X1   g22267(.A1(new_n19290_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n19308_), .ZN(new_n22334_));
  AOI21_X1   g22268(.A1(new_n4709_), .A2(new_n19545_), .B(new_n22334_), .ZN(new_n22335_));
  NOR3_X1    g22269(.A1(new_n22335_), .A2(new_n19571_), .A3(new_n4707_), .ZN(new_n22336_));
  XOR2_X1    g22270(.A1(new_n22336_), .A2(new_n4034_), .Z(new_n22337_));
  NOR2_X1    g22271(.A1(new_n4704_), .A2(new_n4705_), .ZN(new_n22338_));
  OAI21_X1   g22272(.A1(new_n19313_), .A2(new_n4719_), .B(new_n22338_), .ZN(new_n22339_));
  NOR2_X1    g22273(.A1(new_n19593_), .A2(new_n22339_), .ZN(new_n22340_));
  XOR2_X1    g22274(.A1(new_n22340_), .A2(new_n4034_), .Z(new_n22341_));
  NOR2_X1    g22275(.A1(new_n19313_), .A2(new_n4704_), .ZN(new_n22342_));
  NOR2_X1    g22276(.A1(new_n22342_), .A2(new_n4034_), .ZN(new_n22343_));
  NAND2_X1   g22277(.A1(new_n22341_), .A2(new_n22343_), .ZN(new_n22344_));
  NOR2_X1    g22278(.A1(new_n22337_), .A2(new_n22344_), .ZN(new_n22345_));
  NOR2_X1    g22279(.A1(new_n22332_), .A2(new_n22328_), .ZN(new_n22346_));
  OAI21_X1   g22280(.A1(new_n22345_), .A2(new_n22346_), .B(new_n22333_), .ZN(new_n22347_));
  XOR2_X1    g22281(.A1(new_n22259_), .A2(new_n22261_), .Z(new_n22348_));
  AOI22_X1   g22282(.A1(new_n17850_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n19545_), .ZN(new_n22349_));
  AOI21_X1   g22283(.A1(new_n19305_), .A2(new_n4709_), .B(new_n22349_), .ZN(new_n22350_));
  NOR3_X1    g22284(.A1(new_n19618_), .A2(new_n4707_), .A3(new_n22350_), .ZN(new_n22351_));
  XOR2_X1    g22285(.A1(new_n22351_), .A2(new_n4034_), .Z(new_n22352_));
  NAND2_X1   g22286(.A1(new_n22352_), .A2(new_n22348_), .ZN(new_n22353_));
  NAND2_X1   g22287(.A1(new_n22347_), .A2(new_n22353_), .ZN(new_n22354_));
  OR2_X2     g22288(.A1(new_n22352_), .A2(new_n22348_), .Z(new_n22355_));
  NAND2_X1   g22289(.A1(new_n22354_), .A2(new_n22355_), .ZN(new_n22356_));
  INV_X1     g22290(.I(new_n22356_), .ZN(new_n22357_));
  AOI22_X1   g22291(.A1(new_n19305_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n17850_), .ZN(new_n22358_));
  AOI21_X1   g22292(.A1(new_n4709_), .A2(new_n19321_), .B(new_n22358_), .ZN(new_n22359_));
  NOR3_X1    g22293(.A1(new_n22277_), .A2(new_n4707_), .A3(new_n22359_), .ZN(new_n22360_));
  XOR2_X1    g22294(.A1(new_n22360_), .A2(new_n4034_), .Z(new_n22361_));
  NOR2_X1    g22295(.A1(new_n22357_), .A2(new_n22361_), .ZN(new_n22362_));
  INV_X1     g22296(.I(new_n22255_), .ZN(new_n22363_));
  INV_X1     g22297(.I(new_n22262_), .ZN(new_n22364_));
  NOR2_X1    g22298(.A1(new_n22363_), .A2(new_n22364_), .ZN(new_n22365_));
  NOR2_X1    g22299(.A1(new_n22365_), .A2(new_n22263_), .ZN(new_n22366_));
  AOI21_X1   g22300(.A1(new_n22357_), .A2(new_n22361_), .B(new_n22366_), .ZN(new_n22367_));
  NOR2_X1    g22301(.A1(new_n22367_), .A2(new_n22362_), .ZN(new_n22368_));
  XOR2_X1    g22302(.A1(new_n22249_), .A2(new_n21283_), .Z(new_n22369_));
  NAND2_X1   g22303(.A1(new_n22369_), .A2(new_n22263_), .ZN(new_n22370_));
  OAI22_X1   g22304(.A1(new_n22250_), .A2(new_n22264_), .B1(new_n22255_), .B2(new_n22262_), .ZN(new_n22371_));
  NAND2_X1   g22305(.A1(new_n22370_), .A2(new_n22371_), .ZN(new_n22372_));
  AOI22_X1   g22306(.A1(new_n19305_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n19321_), .ZN(new_n22373_));
  AOI21_X1   g22307(.A1(new_n4709_), .A2(new_n17827_), .B(new_n22373_), .ZN(new_n22374_));
  OR3_X2     g22308(.A1(new_n22298_), .A2(new_n4707_), .A3(new_n22374_), .Z(new_n22375_));
  XOR2_X1    g22309(.A1(new_n22375_), .A2(new_n4034_), .Z(new_n22376_));
  NOR2_X1    g22310(.A1(new_n22376_), .A2(new_n22372_), .ZN(new_n22377_));
  NAND2_X1   g22311(.A1(new_n22376_), .A2(new_n22372_), .ZN(new_n22378_));
  OAI21_X1   g22312(.A1(new_n22368_), .A2(new_n22377_), .B(new_n22378_), .ZN(new_n22379_));
  XOR2_X1    g22313(.A1(new_n22271_), .A2(new_n22267_), .Z(new_n22380_));
  AOI21_X1   g22314(.A1(new_n22272_), .A2(new_n22274_), .B(new_n22265_), .ZN(new_n22381_));
  AOI21_X1   g22315(.A1(new_n22265_), .A2(new_n22380_), .B(new_n22381_), .ZN(new_n22382_));
  AOI22_X1   g22316(.A1(new_n17827_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n19321_), .ZN(new_n22383_));
  AOI21_X1   g22317(.A1(new_n19349_), .A2(new_n4709_), .B(new_n22383_), .ZN(new_n22384_));
  NOR3_X1    g22318(.A1(new_n20063_), .A2(new_n4707_), .A3(new_n22384_), .ZN(new_n22385_));
  XOR2_X1    g22319(.A1(new_n22385_), .A2(\a[11] ), .Z(new_n22386_));
  NOR2_X1    g22320(.A1(new_n22382_), .A2(new_n22386_), .ZN(new_n22387_));
  INV_X1     g22321(.I(new_n22387_), .ZN(new_n22388_));
  NAND2_X1   g22322(.A1(new_n22379_), .A2(new_n22388_), .ZN(new_n22389_));
  NAND2_X1   g22323(.A1(new_n22382_), .A2(new_n22386_), .ZN(new_n22390_));
  NAND2_X1   g22324(.A1(new_n22389_), .A2(new_n22390_), .ZN(new_n22391_));
  INV_X1     g22325(.I(new_n22391_), .ZN(new_n22392_));
  NAND3_X1   g22326(.A1(new_n22316_), .A2(new_n22320_), .A3(new_n22326_), .ZN(new_n22393_));
  AOI21_X1   g22327(.A1(new_n22392_), .A2(new_n22393_), .B(new_n22327_), .ZN(new_n22394_));
  AOI22_X1   g22328(.A1(new_n19349_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n19350_), .ZN(new_n22395_));
  AOI21_X1   g22329(.A1(new_n4709_), .A2(new_n17807_), .B(new_n22395_), .ZN(new_n22396_));
  OR3_X2     g22330(.A1(new_n19915_), .A2(new_n4707_), .A3(new_n22396_), .Z(new_n22397_));
  XOR2_X1    g22331(.A1(new_n22397_), .A2(\a[11] ), .Z(new_n22398_));
  INV_X1     g22332(.I(new_n22398_), .ZN(new_n22399_));
  NOR2_X1    g22333(.A1(new_n22394_), .A2(new_n22399_), .ZN(new_n22400_));
  AOI21_X1   g22334(.A1(new_n22318_), .A2(new_n22319_), .B(new_n22317_), .ZN(new_n22401_));
  NOR3_X1    g22335(.A1(new_n22313_), .A2(new_n22315_), .A3(new_n22283_), .ZN(new_n22402_));
  OAI21_X1   g22336(.A1(new_n22401_), .A2(new_n22402_), .B(new_n22325_), .ZN(new_n22403_));
  NOR3_X1    g22337(.A1(new_n22401_), .A2(new_n22402_), .A3(new_n22325_), .ZN(new_n22404_));
  OAI21_X1   g22338(.A1(new_n22391_), .A2(new_n22404_), .B(new_n22403_), .ZN(new_n22405_));
  NOR2_X1    g22339(.A1(new_n22405_), .A2(new_n22398_), .ZN(new_n22406_));
  OAI21_X1   g22340(.A1(new_n22400_), .A2(new_n22406_), .B(new_n22309_), .ZN(new_n22407_));
  INV_X1     g22341(.I(new_n22309_), .ZN(new_n22408_));
  NAND2_X1   g22342(.A1(new_n22405_), .A2(new_n22398_), .ZN(new_n22409_));
  NAND2_X1   g22343(.A1(new_n22394_), .A2(new_n22399_), .ZN(new_n22410_));
  NAND3_X1   g22344(.A1(new_n22410_), .A2(new_n22409_), .A3(new_n22408_), .ZN(new_n22411_));
  NAND3_X1   g22345(.A1(new_n22407_), .A2(new_n22411_), .A3(new_n22243_), .ZN(new_n22412_));
  AOI21_X1   g22346(.A1(new_n22410_), .A2(new_n22409_), .B(new_n22408_), .ZN(new_n22413_));
  NOR3_X1    g22347(.A1(new_n22400_), .A2(new_n22406_), .A3(new_n22309_), .ZN(new_n22414_));
  OAI21_X1   g22348(.A1(new_n22414_), .A2(new_n22413_), .B(new_n22242_), .ZN(new_n22415_));
  NOR3_X1    g22349(.A1(new_n22404_), .A2(new_n22327_), .A3(new_n22391_), .ZN(new_n22416_));
  INV_X1     g22350(.I(new_n22416_), .ZN(new_n22417_));
  OAI21_X1   g22351(.A1(new_n22404_), .A2(new_n22327_), .B(new_n22391_), .ZN(new_n22418_));
  INV_X1     g22352(.I(new_n19538_), .ZN(new_n22419_));
  AOI22_X1   g22353(.A1(new_n19359_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n17807_), .ZN(new_n22420_));
  AOI21_X1   g22354(.A1(new_n6784_), .A2(new_n19365_), .B(new_n22420_), .ZN(new_n22421_));
  OR3_X2     g22355(.A1(new_n22419_), .A2(new_n6776_), .A3(new_n22421_), .Z(new_n22422_));
  XOR2_X1    g22356(.A1(new_n22422_), .A2(\a[8] ), .Z(new_n22423_));
  NAND3_X1   g22357(.A1(new_n22417_), .A2(new_n22418_), .A3(new_n22423_), .ZN(new_n22424_));
  INV_X1     g22358(.I(new_n22368_), .ZN(new_n22425_));
  AOI21_X1   g22359(.A1(new_n22370_), .A2(new_n22371_), .B(new_n22376_), .ZN(new_n22426_));
  INV_X1     g22360(.I(new_n22376_), .ZN(new_n22427_));
  NOR2_X1    g22361(.A1(new_n22427_), .A2(new_n22372_), .ZN(new_n22428_));
  OAI21_X1   g22362(.A1(new_n22426_), .A2(new_n22428_), .B(new_n22425_), .ZN(new_n22429_));
  INV_X1     g22363(.I(new_n22377_), .ZN(new_n22430_));
  NAND2_X1   g22364(.A1(new_n22430_), .A2(new_n22378_), .ZN(new_n22431_));
  NAND2_X1   g22365(.A1(new_n22431_), .A2(new_n22368_), .ZN(new_n22432_));
  NAND2_X1   g22366(.A1(new_n22429_), .A2(new_n22432_), .ZN(new_n22433_));
  AOI22_X1   g22367(.A1(new_n19349_), .A2(new_n7530_), .B1(new_n6789_), .B2(new_n19350_), .ZN(new_n22434_));
  AOI21_X1   g22368(.A1(new_n6784_), .A2(new_n17807_), .B(new_n22434_), .ZN(new_n22435_));
  OR3_X2     g22369(.A1(new_n19915_), .A2(new_n6776_), .A3(new_n22435_), .Z(new_n22436_));
  XOR2_X1    g22370(.A1(new_n22436_), .A2(\a[8] ), .Z(new_n22437_));
  NOR2_X1    g22371(.A1(new_n22433_), .A2(new_n22437_), .ZN(new_n22438_));
  INV_X1     g22372(.I(new_n22438_), .ZN(new_n22439_));
  XOR2_X1    g22373(.A1(new_n22382_), .A2(new_n22386_), .Z(new_n22440_));
  AOI21_X1   g22374(.A1(new_n22388_), .A2(new_n22390_), .B(new_n22379_), .ZN(new_n22441_));
  AOI21_X1   g22375(.A1(new_n22379_), .A2(new_n22440_), .B(new_n22441_), .ZN(new_n22442_));
  INV_X1     g22376(.I(new_n20096_), .ZN(new_n22443_));
  AOI22_X1   g22377(.A1(new_n17807_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n19350_), .ZN(new_n22444_));
  AOI21_X1   g22378(.A1(new_n19359_), .A2(new_n6784_), .B(new_n22444_), .ZN(new_n22445_));
  OR3_X2     g22379(.A1(new_n22443_), .A2(new_n6776_), .A3(new_n22445_), .Z(new_n22446_));
  XOR2_X1    g22380(.A1(new_n22446_), .A2(new_n4009_), .Z(new_n22447_));
  NOR2_X1    g22381(.A1(new_n22442_), .A2(new_n22447_), .ZN(new_n22448_));
  NAND2_X1   g22382(.A1(new_n22442_), .A2(new_n22447_), .ZN(new_n22449_));
  OAI21_X1   g22383(.A1(new_n22439_), .A2(new_n22448_), .B(new_n22449_), .ZN(new_n22450_));
  AOI21_X1   g22384(.A1(new_n22417_), .A2(new_n22418_), .B(new_n22423_), .ZN(new_n22451_));
  OAI21_X1   g22385(.A1(new_n22450_), .A2(new_n22451_), .B(new_n22424_), .ZN(new_n22452_));
  AOI22_X1   g22386(.A1(new_n22415_), .A2(new_n22412_), .B1(new_n22452_), .B2(new_n22243_), .ZN(new_n22453_));
  AOI22_X1   g22387(.A1(new_n17802_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n19365_), .ZN(new_n22454_));
  NOR2_X1    g22388(.A1(new_n17797_), .A2(new_n6785_), .ZN(new_n22455_));
  OAI21_X1   g22389(.A1(new_n22455_), .A2(new_n22454_), .B(new_n6775_), .ZN(new_n22456_));
  NOR2_X1    g22390(.A1(new_n21454_), .A2(new_n22456_), .ZN(new_n22457_));
  XOR2_X1    g22391(.A1(new_n22457_), .A2(new_n4009_), .Z(new_n22458_));
  INV_X1     g22392(.I(new_n22458_), .ZN(new_n22459_));
  NAND2_X1   g22393(.A1(new_n22453_), .A2(new_n22459_), .ZN(new_n22460_));
  AOI22_X1   g22394(.A1(new_n17807_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n19350_), .ZN(new_n22461_));
  AOI21_X1   g22395(.A1(new_n19359_), .A2(new_n4709_), .B(new_n22461_), .ZN(new_n22462_));
  OR3_X2     g22396(.A1(new_n22443_), .A2(new_n4707_), .A3(new_n22462_), .Z(new_n22463_));
  XOR2_X1    g22397(.A1(new_n22463_), .A2(\a[11] ), .Z(new_n22464_));
  OAI21_X1   g22398(.A1(new_n22289_), .A2(new_n22282_), .B(new_n22305_), .ZN(new_n22465_));
  NAND2_X1   g22399(.A1(new_n21387_), .A2(new_n21388_), .ZN(new_n22466_));
  XOR2_X1    g22400(.A1(new_n22466_), .A2(new_n21386_), .Z(new_n22467_));
  NOR2_X1    g22401(.A1(new_n22467_), .A2(new_n21287_), .ZN(new_n22468_));
  NOR2_X1    g22402(.A1(new_n21303_), .A2(new_n21390_), .ZN(new_n22469_));
  NOR2_X1    g22403(.A1(new_n22469_), .A2(new_n21380_), .ZN(new_n22470_));
  NOR2_X1    g22404(.A1(new_n22468_), .A2(new_n22470_), .ZN(new_n22471_));
  AOI22_X1   g22405(.A1(new_n17827_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n19321_), .ZN(new_n22472_));
  AOI21_X1   g22406(.A1(new_n19349_), .A2(new_n6090_), .B(new_n22472_), .ZN(new_n22473_));
  NOR3_X1    g22407(.A1(new_n20063_), .A2(new_n6082_), .A3(new_n22473_), .ZN(new_n22474_));
  XOR2_X1    g22408(.A1(new_n22474_), .A2(\a[14] ), .Z(new_n22475_));
  XNOR2_X1   g22409(.A1(new_n22475_), .A2(new_n22471_), .ZN(new_n22476_));
  AOI21_X1   g22410(.A1(new_n22465_), .A2(new_n22307_), .B(new_n22476_), .ZN(new_n22477_));
  NAND2_X1   g22411(.A1(new_n22465_), .A2(new_n22307_), .ZN(new_n22478_));
  NOR2_X1    g22412(.A1(new_n22475_), .A2(new_n22471_), .ZN(new_n22479_));
  NAND2_X1   g22413(.A1(new_n22475_), .A2(new_n22471_), .ZN(new_n22480_));
  INV_X1     g22414(.I(new_n22480_), .ZN(new_n22481_));
  NOR2_X1    g22415(.A1(new_n22481_), .A2(new_n22479_), .ZN(new_n22482_));
  NOR2_X1    g22416(.A1(new_n22478_), .A2(new_n22482_), .ZN(new_n22483_));
  NOR2_X1    g22417(.A1(new_n22483_), .A2(new_n22477_), .ZN(new_n22484_));
  XOR2_X1    g22418(.A1(new_n22484_), .A2(new_n22464_), .Z(new_n22485_));
  INV_X1     g22419(.I(new_n22485_), .ZN(new_n22486_));
  OAI21_X1   g22420(.A1(new_n22453_), .A2(new_n22459_), .B(new_n22486_), .ZN(new_n22487_));
  AOI21_X1   g22421(.A1(new_n22465_), .A2(new_n22307_), .B(new_n22479_), .ZN(new_n22488_));
  XOR2_X1    g22422(.A1(new_n21321_), .A2(new_n21394_), .Z(new_n22489_));
  NOR2_X1    g22423(.A1(new_n22489_), .A2(new_n21391_), .ZN(new_n22490_));
  NOR2_X1    g22424(.A1(new_n21323_), .A2(new_n21395_), .ZN(new_n22491_));
  INV_X1     g22425(.I(new_n22491_), .ZN(new_n22492_));
  AOI21_X1   g22426(.A1(new_n21391_), .A2(new_n22492_), .B(new_n22490_), .ZN(new_n22493_));
  INV_X1     g22427(.I(new_n22493_), .ZN(new_n22494_));
  OAI22_X1   g22428(.A1(new_n6094_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n6089_), .ZN(new_n22495_));
  NAND2_X1   g22429(.A1(new_n19350_), .A2(new_n6090_), .ZN(new_n22496_));
  AOI21_X1   g22430(.A1(new_n22495_), .A2(new_n22496_), .B(new_n6082_), .ZN(new_n22497_));
  NAND2_X1   g22431(.A1(new_n20535_), .A2(new_n22497_), .ZN(new_n22498_));
  XOR2_X1    g22432(.A1(new_n22498_), .A2(\a[14] ), .Z(new_n22499_));
  NOR2_X1    g22433(.A1(new_n22494_), .A2(new_n22499_), .ZN(new_n22500_));
  INV_X1     g22434(.I(new_n22499_), .ZN(new_n22501_));
  NOR2_X1    g22435(.A1(new_n22501_), .A2(new_n22493_), .ZN(new_n22502_));
  NOR4_X1    g22436(.A1(new_n22488_), .A2(new_n22481_), .A3(new_n22500_), .A4(new_n22502_), .ZN(new_n22503_));
  NOR2_X1    g22437(.A1(new_n22488_), .A2(new_n22481_), .ZN(new_n22504_));
  NOR2_X1    g22438(.A1(new_n22500_), .A2(new_n22502_), .ZN(new_n22505_));
  NOR2_X1    g22439(.A1(new_n22504_), .A2(new_n22505_), .ZN(new_n22506_));
  NOR2_X1    g22440(.A1(new_n22506_), .A2(new_n22503_), .ZN(new_n22507_));
  AOI22_X1   g22441(.A1(new_n19359_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n17807_), .ZN(new_n22508_));
  AOI21_X1   g22442(.A1(new_n4709_), .A2(new_n19365_), .B(new_n22508_), .ZN(new_n22509_));
  OR3_X2     g22443(.A1(new_n22419_), .A2(new_n4707_), .A3(new_n22509_), .Z(new_n22510_));
  XOR2_X1    g22444(.A1(new_n22510_), .A2(\a[11] ), .Z(new_n22511_));
  NAND2_X1   g22445(.A1(new_n22507_), .A2(new_n22511_), .ZN(new_n22512_));
  INV_X1     g22446(.I(new_n22511_), .ZN(new_n22513_));
  OAI21_X1   g22447(.A1(new_n22506_), .A2(new_n22503_), .B(new_n22513_), .ZN(new_n22514_));
  NAND2_X1   g22448(.A1(new_n22512_), .A2(new_n22514_), .ZN(new_n22515_));
  INV_X1     g22449(.I(new_n22464_), .ZN(new_n22516_));
  NAND2_X1   g22450(.A1(new_n22484_), .A2(new_n22516_), .ZN(new_n22517_));
  NOR2_X1    g22451(.A1(new_n22515_), .A2(new_n22517_), .ZN(new_n22518_));
  AOI22_X1   g22452(.A1(new_n22512_), .A2(new_n22514_), .B1(new_n22516_), .B2(new_n22484_), .ZN(new_n22519_));
  NOR2_X1    g22453(.A1(new_n22518_), .A2(new_n22519_), .ZN(new_n22520_));
  INV_X1     g22454(.I(new_n22520_), .ZN(new_n22521_));
  AOI22_X1   g22455(.A1(new_n17798_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n17802_), .ZN(new_n22522_));
  NOR2_X1    g22456(.A1(new_n19375_), .A2(new_n6785_), .ZN(new_n22523_));
  OAI21_X1   g22457(.A1(new_n22523_), .A2(new_n22522_), .B(new_n6775_), .ZN(new_n22524_));
  NOR2_X1    g22458(.A1(new_n21753_), .A2(new_n22524_), .ZN(new_n22525_));
  XOR2_X1    g22459(.A1(new_n22525_), .A2(new_n4009_), .Z(new_n22526_));
  NAND2_X1   g22460(.A1(new_n22521_), .A2(new_n22526_), .ZN(new_n22527_));
  NOR2_X1    g22461(.A1(new_n22521_), .A2(new_n22526_), .ZN(new_n22528_));
  INV_X1     g22462(.I(new_n22528_), .ZN(new_n22529_));
  AOI22_X1   g22463(.A1(new_n22529_), .A2(new_n22527_), .B1(new_n22460_), .B2(new_n22487_), .ZN(new_n22530_));
  INV_X1     g22464(.I(new_n22460_), .ZN(new_n22531_));
  INV_X1     g22465(.I(new_n22487_), .ZN(new_n22532_));
  XOR2_X1    g22466(.A1(new_n22520_), .A2(new_n22526_), .Z(new_n22533_));
  NOR3_X1    g22467(.A1(new_n22533_), .A2(new_n22531_), .A3(new_n22532_), .ZN(new_n22534_));
  AOI22_X1   g22468(.A1(new_n19386_), .A2(new_n6846_), .B1(new_n8799_), .B2(new_n17794_), .ZN(new_n22535_));
  NOR2_X1    g22469(.A1(new_n19393_), .A2(new_n6839_), .ZN(new_n22536_));
  OAI21_X1   g22470(.A1(new_n22535_), .A2(new_n22536_), .B(new_n6835_), .ZN(new_n22537_));
  NOR2_X1    g22471(.A1(new_n20291_), .A2(new_n22537_), .ZN(new_n22538_));
  XOR2_X1    g22472(.A1(new_n22538_), .A2(\a[5] ), .Z(new_n22539_));
  OAI21_X1   g22473(.A1(new_n22534_), .A2(new_n22530_), .B(new_n22539_), .ZN(new_n22540_));
  INV_X1     g22474(.I(new_n20264_), .ZN(new_n22541_));
  AOI22_X1   g22475(.A1(new_n19394_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n17794_), .ZN(new_n22542_));
  AOI21_X1   g22476(.A1(new_n6838_), .A2(new_n19399_), .B(new_n22542_), .ZN(new_n22543_));
  OR3_X2     g22477(.A1(new_n22541_), .A2(new_n6836_), .A3(new_n22543_), .Z(new_n22544_));
  XOR2_X1    g22478(.A1(new_n22544_), .A2(\a[5] ), .Z(new_n22545_));
  NOR2_X1    g22479(.A1(new_n22540_), .A2(new_n22545_), .ZN(new_n22546_));
  INV_X1     g22480(.I(new_n22546_), .ZN(new_n22547_));
  AOI22_X1   g22481(.A1(new_n22487_), .A2(new_n22460_), .B1(new_n22521_), .B2(new_n22526_), .ZN(new_n22548_));
  NOR2_X1    g22482(.A1(new_n22548_), .A2(new_n22528_), .ZN(new_n22549_));
  NOR2_X1    g22483(.A1(new_n21337_), .A2(new_n21335_), .ZN(new_n22550_));
  XOR2_X1    g22484(.A1(new_n22550_), .A2(new_n21401_), .Z(new_n22551_));
  NAND2_X1   g22485(.A1(new_n22551_), .A2(new_n21397_), .ZN(new_n22552_));
  OAI21_X1   g22486(.A1(new_n21338_), .A2(new_n21404_), .B(new_n21324_), .ZN(new_n22553_));
  NAND2_X1   g22487(.A1(new_n22552_), .A2(new_n22553_), .ZN(new_n22554_));
  AOI22_X1   g22488(.A1(new_n19349_), .A2(new_n6180_), .B1(new_n6095_), .B2(new_n19350_), .ZN(new_n22555_));
  AOI21_X1   g22489(.A1(new_n6090_), .A2(new_n17807_), .B(new_n22555_), .ZN(new_n22556_));
  OR3_X2     g22490(.A1(new_n19915_), .A2(new_n6082_), .A3(new_n22556_), .Z(new_n22557_));
  XOR2_X1    g22491(.A1(new_n22557_), .A2(\a[14] ), .Z(new_n22558_));
  OAI21_X1   g22492(.A1(new_n22503_), .A2(new_n22502_), .B(new_n22558_), .ZN(new_n22559_));
  NOR3_X1    g22493(.A1(new_n22503_), .A2(new_n22502_), .A3(new_n22558_), .ZN(new_n22560_));
  INV_X1     g22494(.I(new_n22560_), .ZN(new_n22561_));
  AOI21_X1   g22495(.A1(new_n22561_), .A2(new_n22559_), .B(new_n22554_), .ZN(new_n22562_));
  INV_X1     g22496(.I(new_n22554_), .ZN(new_n22563_));
  INV_X1     g22497(.I(new_n22559_), .ZN(new_n22564_));
  NOR3_X1    g22498(.A1(new_n22564_), .A2(new_n22560_), .A3(new_n22563_), .ZN(new_n22565_));
  NOR2_X1    g22499(.A1(new_n22562_), .A2(new_n22565_), .ZN(new_n22566_));
  AOI22_X1   g22500(.A1(new_n19359_), .A2(new_n6480_), .B1(new_n4720_), .B2(new_n19365_), .ZN(new_n22567_));
  AOI21_X1   g22501(.A1(new_n4709_), .A2(new_n17802_), .B(new_n22567_), .ZN(new_n22568_));
  OR3_X2     g22502(.A1(new_n22238_), .A2(new_n4707_), .A3(new_n22568_), .Z(new_n22569_));
  XOR2_X1    g22503(.A1(new_n22569_), .A2(\a[11] ), .Z(new_n22570_));
  OAI21_X1   g22504(.A1(new_n22483_), .A2(new_n22477_), .B(new_n22464_), .ZN(new_n22571_));
  NAND3_X1   g22505(.A1(new_n22512_), .A2(new_n22514_), .A3(new_n22571_), .ZN(new_n22572_));
  NAND2_X1   g22506(.A1(new_n22572_), .A2(new_n22570_), .ZN(new_n22573_));
  INV_X1     g22507(.I(new_n22573_), .ZN(new_n22574_));
  INV_X1     g22508(.I(new_n22570_), .ZN(new_n22575_));
  NAND4_X1   g22509(.A1(new_n22512_), .A2(new_n22514_), .A3(new_n22575_), .A4(new_n22571_), .ZN(new_n22576_));
  INV_X1     g22510(.I(new_n22576_), .ZN(new_n22577_));
  OAI21_X1   g22511(.A1(new_n22574_), .A2(new_n22577_), .B(new_n22566_), .ZN(new_n22578_));
  OR2_X2     g22512(.A1(new_n22562_), .A2(new_n22565_), .Z(new_n22579_));
  NAND3_X1   g22513(.A1(new_n22579_), .A2(new_n22573_), .A3(new_n22576_), .ZN(new_n22580_));
  OAI22_X1   g22514(.A1(new_n19375_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n17797_), .ZN(new_n22581_));
  NAND2_X1   g22515(.A1(new_n19386_), .A2(new_n6784_), .ZN(new_n22582_));
  AOI21_X1   g22516(.A1(new_n22582_), .A2(new_n22581_), .B(new_n6776_), .ZN(new_n22583_));
  NAND2_X1   g22517(.A1(new_n20162_), .A2(new_n22583_), .ZN(new_n22584_));
  XOR2_X1    g22518(.A1(new_n22584_), .A2(\a[8] ), .Z(new_n22585_));
  INV_X1     g22519(.I(new_n22585_), .ZN(new_n22586_));
  NAND3_X1   g22520(.A1(new_n22578_), .A2(new_n22580_), .A3(new_n22586_), .ZN(new_n22587_));
  AOI21_X1   g22521(.A1(new_n22573_), .A2(new_n22576_), .B(new_n22579_), .ZN(new_n22588_));
  INV_X1     g22522(.I(new_n22580_), .ZN(new_n22589_));
  OAI21_X1   g22523(.A1(new_n22589_), .A2(new_n22588_), .B(new_n22585_), .ZN(new_n22590_));
  NAND2_X1   g22524(.A1(new_n22590_), .A2(new_n22587_), .ZN(new_n22591_));
  XOR2_X1    g22525(.A1(new_n22549_), .A2(new_n22591_), .Z(new_n22592_));
  NAND2_X1   g22526(.A1(new_n22540_), .A2(new_n22545_), .ZN(new_n22593_));
  OAI21_X1   g22527(.A1(new_n22592_), .A2(new_n22593_), .B(new_n22547_), .ZN(new_n22594_));
  AOI22_X1   g22528(.A1(new_n17802_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n19365_), .ZN(new_n22595_));
  NOR2_X1    g22529(.A1(new_n17797_), .A2(new_n4710_), .ZN(new_n22596_));
  OAI21_X1   g22530(.A1(new_n22596_), .A2(new_n22595_), .B(new_n4706_), .ZN(new_n22597_));
  NOR2_X1    g22531(.A1(new_n21454_), .A2(new_n22597_), .ZN(new_n22598_));
  XOR2_X1    g22532(.A1(new_n22598_), .A2(new_n4034_), .Z(new_n22599_));
  XOR2_X1    g22533(.A1(new_n21482_), .A2(new_n21447_), .Z(new_n22600_));
  NAND2_X1   g22534(.A1(new_n22566_), .A2(new_n22575_), .ZN(new_n22601_));
  NAND2_X1   g22535(.A1(new_n22579_), .A2(new_n22570_), .ZN(new_n22602_));
  AOI22_X1   g22536(.A1(new_n22602_), .A2(new_n22601_), .B1(new_n22575_), .B2(new_n22572_), .ZN(new_n22603_));
  NAND2_X1   g22537(.A1(new_n22603_), .A2(new_n22600_), .ZN(new_n22604_));
  INV_X1     g22538(.I(new_n22604_), .ZN(new_n22605_));
  NOR2_X1    g22539(.A1(new_n22603_), .A2(new_n22600_), .ZN(new_n22606_));
  OAI21_X1   g22540(.A1(new_n22605_), .A2(new_n22606_), .B(new_n22599_), .ZN(new_n22607_));
  INV_X1     g22541(.I(new_n22599_), .ZN(new_n22608_));
  INV_X1     g22542(.I(new_n22606_), .ZN(new_n22609_));
  NAND3_X1   g22543(.A1(new_n22609_), .A2(new_n22608_), .A3(new_n22604_), .ZN(new_n22610_));
  NAND2_X1   g22544(.A1(new_n22607_), .A2(new_n22610_), .ZN(new_n22611_));
  AOI21_X1   g22545(.A1(new_n22578_), .A2(new_n22580_), .B(new_n22586_), .ZN(new_n22612_));
  NOR3_X1    g22546(.A1(new_n22548_), .A2(new_n22591_), .A3(new_n22528_), .ZN(new_n22613_));
  AOI22_X1   g22547(.A1(new_n19386_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n20127_), .ZN(new_n22614_));
  NOR2_X1    g22548(.A1(new_n17793_), .A2(new_n6785_), .ZN(new_n22615_));
  OAI21_X1   g22549(.A1(new_n22614_), .A2(new_n22615_), .B(new_n6775_), .ZN(new_n22616_));
  NOR2_X1    g22550(.A1(new_n21632_), .A2(new_n22616_), .ZN(new_n22617_));
  XOR2_X1    g22551(.A1(new_n22617_), .A2(new_n4009_), .Z(new_n22618_));
  OAI21_X1   g22552(.A1(new_n22613_), .A2(new_n22612_), .B(new_n22618_), .ZN(new_n22619_));
  OAI21_X1   g22553(.A1(new_n22532_), .A2(new_n22531_), .B(new_n22527_), .ZN(new_n22620_));
  NOR3_X1    g22554(.A1(new_n22589_), .A2(new_n22588_), .A3(new_n22585_), .ZN(new_n22621_));
  NOR2_X1    g22555(.A1(new_n22621_), .A2(new_n22612_), .ZN(new_n22622_));
  NAND3_X1   g22556(.A1(new_n22620_), .A2(new_n22529_), .A3(new_n22622_), .ZN(new_n22623_));
  INV_X1     g22557(.I(new_n22618_), .ZN(new_n22624_));
  NAND3_X1   g22558(.A1(new_n22623_), .A2(new_n22590_), .A3(new_n22624_), .ZN(new_n22625_));
  AOI21_X1   g22559(.A1(new_n22625_), .A2(new_n22619_), .B(new_n22611_), .ZN(new_n22626_));
  AOI21_X1   g22560(.A1(new_n22609_), .A2(new_n22604_), .B(new_n22608_), .ZN(new_n22627_));
  NOR3_X1    g22561(.A1(new_n22605_), .A2(new_n22599_), .A3(new_n22606_), .ZN(new_n22628_));
  NOR2_X1    g22562(.A1(new_n22627_), .A2(new_n22628_), .ZN(new_n22629_));
  AOI21_X1   g22563(.A1(new_n22623_), .A2(new_n22590_), .B(new_n22624_), .ZN(new_n22630_));
  NOR3_X1    g22564(.A1(new_n22613_), .A2(new_n22612_), .A3(new_n22618_), .ZN(new_n22631_));
  NOR3_X1    g22565(.A1(new_n22630_), .A2(new_n22631_), .A3(new_n22629_), .ZN(new_n22632_));
  OAI22_X1   g22566(.A1(new_n19400_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n19393_), .ZN(new_n22633_));
  NAND2_X1   g22567(.A1(new_n17790_), .A2(new_n6838_), .ZN(new_n22634_));
  AOI21_X1   g22568(.A1(new_n22634_), .A2(new_n22633_), .B(new_n6836_), .ZN(new_n22635_));
  NAND2_X1   g22569(.A1(new_n20251_), .A2(new_n22635_), .ZN(new_n22636_));
  XOR2_X1    g22570(.A1(new_n22636_), .A2(\a[5] ), .Z(new_n22637_));
  INV_X1     g22571(.I(new_n22637_), .ZN(new_n22638_));
  NOR3_X1    g22572(.A1(new_n22632_), .A2(new_n22626_), .A3(new_n22638_), .ZN(new_n22639_));
  OAI21_X1   g22573(.A1(new_n22630_), .A2(new_n22631_), .B(new_n22629_), .ZN(new_n22640_));
  NAND3_X1   g22574(.A1(new_n22625_), .A2(new_n22619_), .A3(new_n22611_), .ZN(new_n22641_));
  AOI21_X1   g22575(.A1(new_n22640_), .A2(new_n22641_), .B(new_n22637_), .ZN(new_n22642_));
  OAI21_X1   g22576(.A1(new_n22639_), .A2(new_n22642_), .B(new_n22594_), .ZN(new_n22643_));
  XOR2_X1    g22577(.A1(new_n22549_), .A2(new_n22622_), .Z(new_n22644_));
  INV_X1     g22578(.I(new_n22593_), .ZN(new_n22645_));
  AOI21_X1   g22579(.A1(new_n22645_), .A2(new_n22644_), .B(new_n22546_), .ZN(new_n22646_));
  AOI21_X1   g22580(.A1(new_n22640_), .A2(new_n22641_), .B(new_n22638_), .ZN(new_n22647_));
  NOR3_X1    g22581(.A1(new_n22632_), .A2(new_n22626_), .A3(new_n22637_), .ZN(new_n22648_));
  OAI21_X1   g22582(.A1(new_n22648_), .A2(new_n22647_), .B(new_n22646_), .ZN(new_n22649_));
  NAND3_X1   g22583(.A1(new_n22643_), .A2(new_n22649_), .A3(new_n22237_), .ZN(new_n22650_));
  NAND3_X1   g22584(.A1(new_n22640_), .A2(new_n22641_), .A3(new_n22637_), .ZN(new_n22651_));
  OAI21_X1   g22585(.A1(new_n22632_), .A2(new_n22626_), .B(new_n22638_), .ZN(new_n22652_));
  AOI21_X1   g22586(.A1(new_n22652_), .A2(new_n22651_), .B(new_n22646_), .ZN(new_n22653_));
  OAI21_X1   g22587(.A1(new_n22632_), .A2(new_n22626_), .B(new_n22637_), .ZN(new_n22654_));
  NAND3_X1   g22588(.A1(new_n22640_), .A2(new_n22641_), .A3(new_n22638_), .ZN(new_n22655_));
  AOI21_X1   g22589(.A1(new_n22654_), .A2(new_n22655_), .B(new_n22594_), .ZN(new_n22656_));
  OAI21_X1   g22590(.A1(new_n22656_), .A2(new_n22653_), .B(new_n22236_), .ZN(new_n22657_));
  NAND2_X1   g22591(.A1(new_n22650_), .A2(new_n22657_), .ZN(new_n22658_));
  NAND2_X1   g22592(.A1(new_n22658_), .A2(new_n22236_), .ZN(new_n22659_));
  OAI22_X1   g22593(.A1(new_n17789_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n19400_), .ZN(new_n22660_));
  OAI21_X1   g22594(.A1(new_n9489_), .A2(new_n19410_), .B(new_n22660_), .ZN(new_n22661_));
  AOI21_X1   g22595(.A1(new_n20864_), .A2(new_n6922_), .B(new_n22661_), .ZN(new_n22662_));
  XOR2_X1    g22596(.A1(new_n22662_), .A2(\a[2] ), .Z(new_n22663_));
  INV_X1     g22597(.I(new_n22663_), .ZN(new_n22664_));
  OR2_X2     g22598(.A1(new_n22534_), .A2(new_n22530_), .Z(new_n22665_));
  NOR2_X1    g22599(.A1(new_n22665_), .A2(new_n22539_), .ZN(new_n22666_));
  INV_X1     g22600(.I(new_n22666_), .ZN(new_n22667_));
  NAND3_X1   g22601(.A1(new_n22667_), .A2(new_n22540_), .A3(new_n22664_), .ZN(new_n22668_));
  INV_X1     g22602(.I(new_n22540_), .ZN(new_n22669_));
  OAI21_X1   g22603(.A1(new_n22666_), .A2(new_n22669_), .B(new_n22663_), .ZN(new_n22670_));
  NAND2_X1   g22604(.A1(new_n22668_), .A2(new_n22670_), .ZN(new_n22671_));
  NAND2_X1   g22605(.A1(new_n22671_), .A2(new_n22663_), .ZN(new_n22672_));
  INV_X1     g22606(.I(new_n20251_), .ZN(new_n22673_));
  NAND2_X1   g22607(.A1(new_n17790_), .A2(new_n9488_), .ZN(new_n22674_));
  NAND2_X1   g22608(.A1(new_n19399_), .A2(new_n9503_), .ZN(new_n22675_));
  AOI21_X1   g22609(.A1(new_n19394_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n22676_));
  NAND4_X1   g22610(.A1(new_n22673_), .A2(new_n22674_), .A3(new_n22675_), .A4(new_n22676_), .ZN(new_n22677_));
  XOR2_X1    g22611(.A1(new_n22677_), .A2(\a[2] ), .Z(new_n22678_));
  INV_X1     g22612(.I(new_n22678_), .ZN(new_n22679_));
  NAND2_X1   g22613(.A1(new_n19399_), .A2(new_n9488_), .ZN(new_n22680_));
  NAND2_X1   g22614(.A1(new_n19394_), .A2(new_n9503_), .ZN(new_n22681_));
  AOI21_X1   g22615(.A1(new_n17794_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n22682_));
  NAND4_X1   g22616(.A1(new_n20264_), .A2(new_n22680_), .A3(new_n22681_), .A4(new_n22682_), .ZN(new_n22683_));
  XOR2_X1    g22617(.A1(new_n22683_), .A2(\a[2] ), .Z(new_n22684_));
  AOI22_X1   g22618(.A1(new_n19386_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n20127_), .ZN(new_n22685_));
  AOI21_X1   g22619(.A1(new_n9488_), .A2(new_n17794_), .B(new_n22685_), .ZN(new_n22686_));
  OAI21_X1   g22620(.A1(new_n21632_), .A2(new_n9482_), .B(new_n22686_), .ZN(new_n22687_));
  XOR2_X1    g22621(.A1(new_n22687_), .A2(new_n4387_), .Z(new_n22688_));
  INV_X1     g22622(.I(new_n22688_), .ZN(new_n22689_));
  AOI22_X1   g22623(.A1(new_n19359_), .A2(new_n6846_), .B1(new_n8799_), .B2(new_n19365_), .ZN(new_n22690_));
  AOI21_X1   g22624(.A1(new_n6838_), .A2(new_n17802_), .B(new_n22690_), .ZN(new_n22691_));
  OR3_X2     g22625(.A1(new_n22238_), .A2(new_n6836_), .A3(new_n22691_), .Z(new_n22692_));
  XOR2_X1    g22626(.A1(new_n22692_), .A2(\a[5] ), .Z(new_n22693_));
  INV_X1     g22627(.I(new_n22693_), .ZN(new_n22694_));
  XNOR2_X1   g22628(.A1(new_n22433_), .A2(new_n22437_), .ZN(new_n22695_));
  NOR2_X1    g22629(.A1(new_n22695_), .A2(new_n22694_), .ZN(new_n22696_));
  AOI22_X1   g22630(.A1(new_n19290_), .A2(new_n7530_), .B1(new_n6789_), .B2(new_n19308_), .ZN(new_n22697_));
  AOI21_X1   g22631(.A1(new_n6784_), .A2(new_n19545_), .B(new_n22697_), .ZN(new_n22698_));
  NAND2_X1   g22632(.A1(new_n19564_), .A2(new_n6775_), .ZN(new_n22699_));
  NOR2_X1    g22633(.A1(new_n22699_), .A2(new_n22698_), .ZN(new_n22700_));
  NAND2_X1   g22634(.A1(new_n19290_), .A2(new_n6789_), .ZN(new_n22701_));
  NOR2_X1    g22635(.A1(new_n6773_), .A2(new_n6774_), .ZN(new_n22702_));
  NAND2_X1   g22636(.A1(new_n22701_), .A2(new_n22702_), .ZN(new_n22703_));
  NOR2_X1    g22637(.A1(new_n19593_), .A2(new_n22703_), .ZN(new_n22704_));
  INV_X1     g22638(.I(new_n22704_), .ZN(new_n22705_));
  NOR2_X1    g22639(.A1(new_n19313_), .A2(new_n6773_), .ZN(new_n22706_));
  NOR4_X1    g22640(.A1(new_n22700_), .A2(new_n4009_), .A3(new_n22705_), .A4(new_n22706_), .ZN(new_n22707_));
  NAND2_X1   g22641(.A1(new_n22707_), .A2(new_n22342_), .ZN(new_n22708_));
  NOR2_X1    g22642(.A1(new_n22707_), .A2(new_n22342_), .ZN(new_n22709_));
  OAI22_X1   g22643(.A1(new_n19272_), .A2(new_n6783_), .B1(new_n6788_), .B2(new_n19275_), .ZN(new_n22710_));
  NAND2_X1   g22644(.A1(new_n17850_), .A2(new_n6784_), .ZN(new_n22711_));
  AOI21_X1   g22645(.A1(new_n22710_), .A2(new_n22711_), .B(new_n6776_), .ZN(new_n22712_));
  NAND2_X1   g22646(.A1(new_n19553_), .A2(new_n22712_), .ZN(new_n22713_));
  XOR2_X1    g22647(.A1(new_n22713_), .A2(\a[8] ), .Z(new_n22714_));
  INV_X1     g22648(.I(new_n22714_), .ZN(new_n22715_));
  OAI21_X1   g22649(.A1(new_n22715_), .A2(new_n22709_), .B(new_n22708_), .ZN(new_n22716_));
  XNOR2_X1   g22650(.A1(new_n22341_), .A2(new_n22343_), .ZN(new_n22717_));
  NOR2_X1    g22651(.A1(new_n22716_), .A2(new_n22717_), .ZN(new_n22718_));
  INV_X1     g22652(.I(new_n22718_), .ZN(new_n22719_));
  NAND2_X1   g22653(.A1(new_n22716_), .A2(new_n22717_), .ZN(new_n22720_));
  INV_X1     g22654(.I(new_n22720_), .ZN(new_n22721_));
  NOR2_X1    g22655(.A1(new_n22716_), .A2(new_n22717_), .ZN(new_n22722_));
  AOI22_X1   g22656(.A1(new_n17850_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n19545_), .ZN(new_n22723_));
  AOI21_X1   g22657(.A1(new_n19305_), .A2(new_n6784_), .B(new_n22723_), .ZN(new_n22724_));
  OR3_X2     g22658(.A1(new_n19618_), .A2(new_n6776_), .A3(new_n22724_), .Z(new_n22725_));
  XOR2_X1    g22659(.A1(new_n22725_), .A2(\a[8] ), .Z(new_n22726_));
  OAI21_X1   g22660(.A1(new_n22721_), .A2(new_n22722_), .B(new_n22726_), .ZN(new_n22727_));
  NAND2_X1   g22661(.A1(new_n22727_), .A2(new_n22719_), .ZN(new_n22728_));
  OAI22_X1   g22662(.A1(new_n19304_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n17849_), .ZN(new_n22729_));
  NAND2_X1   g22663(.A1(new_n19321_), .A2(new_n6784_), .ZN(new_n22730_));
  AOI21_X1   g22664(.A1(new_n22729_), .A2(new_n22730_), .B(new_n6776_), .ZN(new_n22731_));
  NAND2_X1   g22665(.A1(new_n19647_), .A2(new_n22731_), .ZN(new_n22732_));
  XOR2_X1    g22666(.A1(new_n22732_), .A2(\a[8] ), .Z(new_n22733_));
  INV_X1     g22667(.I(new_n22733_), .ZN(new_n22734_));
  NAND2_X1   g22668(.A1(new_n22728_), .A2(new_n22734_), .ZN(new_n22735_));
  INV_X1     g22669(.I(new_n22345_), .ZN(new_n22736_));
  NAND2_X1   g22670(.A1(new_n22337_), .A2(new_n22344_), .ZN(new_n22737_));
  NAND2_X1   g22671(.A1(new_n22736_), .A2(new_n22737_), .ZN(new_n22738_));
  OAI21_X1   g22672(.A1(new_n22728_), .A2(new_n22734_), .B(new_n22738_), .ZN(new_n22739_));
  NAND2_X1   g22673(.A1(new_n22739_), .A2(new_n22735_), .ZN(new_n22740_));
  XOR2_X1    g22674(.A1(new_n22332_), .A2(new_n22260_), .Z(new_n22741_));
  INV_X1     g22675(.I(new_n22333_), .ZN(new_n22742_));
  OAI21_X1   g22676(.A1(new_n22742_), .A2(new_n22346_), .B(new_n22736_), .ZN(new_n22743_));
  OAI21_X1   g22677(.A1(new_n22741_), .A2(new_n22736_), .B(new_n22743_), .ZN(new_n22744_));
  AOI22_X1   g22678(.A1(new_n19305_), .A2(new_n7530_), .B1(new_n6789_), .B2(new_n19321_), .ZN(new_n22745_));
  AOI21_X1   g22679(.A1(new_n6784_), .A2(new_n17827_), .B(new_n22745_), .ZN(new_n22746_));
  NOR3_X1    g22680(.A1(new_n22298_), .A2(new_n6776_), .A3(new_n22746_), .ZN(new_n22747_));
  XOR2_X1    g22681(.A1(new_n22747_), .A2(\a[8] ), .Z(new_n22748_));
  XOR2_X1    g22682(.A1(new_n22748_), .A2(new_n22744_), .Z(new_n22749_));
  NAND2_X1   g22683(.A1(new_n22748_), .A2(new_n22744_), .ZN(new_n22750_));
  OR2_X2     g22684(.A1(new_n22748_), .A2(new_n22744_), .Z(new_n22751_));
  NAND2_X1   g22685(.A1(new_n22751_), .A2(new_n22750_), .ZN(new_n22752_));
  MUX2_X1    g22686(.I0(new_n22752_), .I1(new_n22749_), .S(new_n22740_), .Z(new_n22753_));
  AOI22_X1   g22687(.A1(new_n19349_), .A2(new_n6846_), .B1(new_n8799_), .B2(new_n19350_), .ZN(new_n22754_));
  AOI21_X1   g22688(.A1(new_n6838_), .A2(new_n17807_), .B(new_n22754_), .ZN(new_n22755_));
  NOR3_X1    g22689(.A1(new_n19915_), .A2(new_n6836_), .A3(new_n22755_), .ZN(new_n22756_));
  XOR2_X1    g22690(.A1(new_n22756_), .A2(new_n65_), .Z(new_n22757_));
  NOR2_X1    g22691(.A1(new_n22753_), .A2(new_n22757_), .ZN(new_n22758_));
  XOR2_X1    g22692(.A1(new_n22352_), .A2(new_n22348_), .Z(new_n22759_));
  AOI21_X1   g22693(.A1(new_n22353_), .A2(new_n22355_), .B(new_n22347_), .ZN(new_n22760_));
  AOI21_X1   g22694(.A1(new_n22347_), .A2(new_n22759_), .B(new_n22760_), .ZN(new_n22761_));
  AOI22_X1   g22695(.A1(new_n17827_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n19321_), .ZN(new_n22762_));
  AOI21_X1   g22696(.A1(new_n19349_), .A2(new_n6784_), .B(new_n22762_), .ZN(new_n22763_));
  NOR3_X1    g22697(.A1(new_n20063_), .A2(new_n6776_), .A3(new_n22763_), .ZN(new_n22764_));
  XOR2_X1    g22698(.A1(new_n22764_), .A2(new_n4009_), .Z(new_n22765_));
  INV_X1     g22699(.I(new_n22765_), .ZN(new_n22766_));
  NOR2_X1    g22700(.A1(new_n22766_), .A2(new_n22761_), .ZN(new_n22767_));
  NAND2_X1   g22701(.A1(new_n22766_), .A2(new_n22761_), .ZN(new_n22768_));
  INV_X1     g22702(.I(new_n22768_), .ZN(new_n22769_));
  NAND2_X1   g22703(.A1(new_n22740_), .A2(new_n22744_), .ZN(new_n22770_));
  NOR3_X1    g22704(.A1(new_n22769_), .A2(new_n22767_), .A3(new_n22770_), .ZN(new_n22771_));
  INV_X1     g22705(.I(new_n22767_), .ZN(new_n22772_));
  AOI22_X1   g22706(.A1(new_n22772_), .A2(new_n22768_), .B1(new_n22740_), .B2(new_n22744_), .ZN(new_n22773_));
  XOR2_X1    g22707(.A1(new_n22740_), .A2(new_n22744_), .Z(new_n22774_));
  NAND2_X1   g22708(.A1(new_n22774_), .A2(new_n22748_), .ZN(new_n22775_));
  NOR3_X1    g22709(.A1(new_n22775_), .A2(new_n22771_), .A3(new_n22773_), .ZN(new_n22776_));
  OAI21_X1   g22710(.A1(new_n22773_), .A2(new_n22771_), .B(new_n22775_), .ZN(new_n22777_));
  INV_X1     g22711(.I(new_n22777_), .ZN(new_n22778_));
  AOI22_X1   g22712(.A1(new_n17807_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n19350_), .ZN(new_n22779_));
  AOI21_X1   g22713(.A1(new_n19359_), .A2(new_n6838_), .B(new_n22779_), .ZN(new_n22780_));
  OR3_X2     g22714(.A1(new_n22443_), .A2(new_n6836_), .A3(new_n22780_), .Z(new_n22781_));
  XOR2_X1    g22715(.A1(new_n22781_), .A2(\a[5] ), .Z(new_n22782_));
  OAI21_X1   g22716(.A1(new_n22778_), .A2(new_n22776_), .B(new_n22782_), .ZN(new_n22783_));
  NOR3_X1    g22717(.A1(new_n22778_), .A2(new_n22776_), .A3(new_n22782_), .ZN(new_n22784_));
  AOI21_X1   g22718(.A1(new_n22758_), .A2(new_n22783_), .B(new_n22784_), .ZN(new_n22785_));
  NOR2_X1    g22719(.A1(new_n22356_), .A2(new_n22361_), .ZN(new_n22786_));
  INV_X1     g22720(.I(new_n22786_), .ZN(new_n22787_));
  NAND2_X1   g22721(.A1(new_n22356_), .A2(new_n22361_), .ZN(new_n22788_));
  AOI21_X1   g22722(.A1(new_n22787_), .A2(new_n22788_), .B(new_n22364_), .ZN(new_n22789_));
  INV_X1     g22723(.I(new_n22789_), .ZN(new_n22790_));
  NAND3_X1   g22724(.A1(new_n22787_), .A2(new_n22364_), .A3(new_n22788_), .ZN(new_n22791_));
  AOI21_X1   g22725(.A1(new_n22790_), .A2(new_n22791_), .B(new_n22255_), .ZN(new_n22792_));
  INV_X1     g22726(.I(new_n22788_), .ZN(new_n22793_));
  NOR3_X1    g22727(.A1(new_n22793_), .A2(new_n22262_), .A3(new_n22786_), .ZN(new_n22794_));
  NOR3_X1    g22728(.A1(new_n22789_), .A2(new_n22794_), .A3(new_n22363_), .ZN(new_n22795_));
  NOR2_X1    g22729(.A1(new_n22792_), .A2(new_n22795_), .ZN(new_n22796_));
  INV_X1     g22730(.I(new_n22796_), .ZN(new_n22797_));
  NAND2_X1   g22731(.A1(new_n22740_), .A2(new_n22751_), .ZN(new_n22798_));
  INV_X1     g22732(.I(new_n22798_), .ZN(new_n22799_));
  NAND3_X1   g22733(.A1(new_n22772_), .A2(new_n22750_), .A3(new_n22768_), .ZN(new_n22800_));
  OAI22_X1   g22734(.A1(new_n6788_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n6783_), .ZN(new_n22801_));
  NAND2_X1   g22735(.A1(new_n19350_), .A2(new_n6784_), .ZN(new_n22802_));
  AOI21_X1   g22736(.A1(new_n22801_), .A2(new_n22802_), .B(new_n6776_), .ZN(new_n22803_));
  NAND2_X1   g22737(.A1(new_n20535_), .A2(new_n22803_), .ZN(new_n22804_));
  XOR2_X1    g22738(.A1(new_n22804_), .A2(\a[8] ), .Z(new_n22805_));
  OAI21_X1   g22739(.A1(new_n22799_), .A2(new_n22800_), .B(new_n22805_), .ZN(new_n22806_));
  NOR3_X1    g22740(.A1(new_n22799_), .A2(new_n22800_), .A3(new_n22805_), .ZN(new_n22807_));
  INV_X1     g22741(.I(new_n22807_), .ZN(new_n22808_));
  AOI21_X1   g22742(.A1(new_n22806_), .A2(new_n22808_), .B(new_n22797_), .ZN(new_n22809_));
  INV_X1     g22743(.I(new_n22806_), .ZN(new_n22810_));
  NOR3_X1    g22744(.A1(new_n22810_), .A2(new_n22807_), .A3(new_n22796_), .ZN(new_n22811_));
  AOI22_X1   g22745(.A1(new_n19359_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n17807_), .ZN(new_n22812_));
  AOI21_X1   g22746(.A1(new_n6838_), .A2(new_n19365_), .B(new_n22812_), .ZN(new_n22813_));
  OR3_X2     g22747(.A1(new_n22419_), .A2(new_n6836_), .A3(new_n22813_), .Z(new_n22814_));
  XOR2_X1    g22748(.A1(new_n22814_), .A2(\a[5] ), .Z(new_n22815_));
  INV_X1     g22749(.I(new_n22815_), .ZN(new_n22816_));
  NOR3_X1    g22750(.A1(new_n22809_), .A2(new_n22811_), .A3(new_n22816_), .ZN(new_n22817_));
  OAI21_X1   g22751(.A1(new_n22810_), .A2(new_n22807_), .B(new_n22796_), .ZN(new_n22818_));
  NAND3_X1   g22752(.A1(new_n22797_), .A2(new_n22808_), .A3(new_n22806_), .ZN(new_n22819_));
  AOI21_X1   g22753(.A1(new_n22819_), .A2(new_n22818_), .B(new_n22815_), .ZN(new_n22820_));
  NOR2_X1    g22754(.A1(new_n22817_), .A2(new_n22820_), .ZN(new_n22821_));
  XOR2_X1    g22755(.A1(new_n22433_), .A2(new_n22437_), .Z(new_n22822_));
  NOR2_X1    g22756(.A1(new_n22822_), .A2(new_n22693_), .ZN(new_n22823_));
  NOR2_X1    g22757(.A1(new_n22695_), .A2(new_n22694_), .ZN(new_n22824_));
  NAND3_X1   g22758(.A1(new_n22819_), .A2(new_n22818_), .A3(new_n22815_), .ZN(new_n22825_));
  OAI21_X1   g22759(.A1(new_n22824_), .A2(new_n22823_), .B(new_n22825_), .ZN(new_n22826_));
  AOI21_X1   g22760(.A1(new_n22785_), .A2(new_n22821_), .B(new_n22826_), .ZN(new_n22827_));
  NAND2_X1   g22761(.A1(new_n22440_), .A2(new_n22379_), .ZN(new_n22828_));
  INV_X1     g22762(.I(new_n22390_), .ZN(new_n22829_));
  NOR2_X1    g22763(.A1(new_n22829_), .A2(new_n22387_), .ZN(new_n22830_));
  OAI21_X1   g22764(.A1(new_n22379_), .A2(new_n22830_), .B(new_n22828_), .ZN(new_n22831_));
  NOR2_X1    g22765(.A1(new_n22831_), .A2(new_n22447_), .ZN(new_n22832_));
  INV_X1     g22766(.I(new_n22447_), .ZN(new_n22833_));
  NOR2_X1    g22767(.A1(new_n22442_), .A2(new_n22833_), .ZN(new_n22834_));
  OAI21_X1   g22768(.A1(new_n22834_), .A2(new_n22832_), .B(new_n22438_), .ZN(new_n22835_));
  NOR2_X1    g22769(.A1(new_n22831_), .A2(new_n22833_), .ZN(new_n22836_));
  OAI21_X1   g22770(.A1(new_n22448_), .A2(new_n22836_), .B(new_n22439_), .ZN(new_n22837_));
  AOI22_X1   g22771(.A1(new_n17802_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n19365_), .ZN(new_n22838_));
  NOR2_X1    g22772(.A1(new_n17797_), .A2(new_n6839_), .ZN(new_n22839_));
  OAI21_X1   g22773(.A1(new_n22839_), .A2(new_n22838_), .B(new_n6835_), .ZN(new_n22840_));
  NOR2_X1    g22774(.A1(new_n21454_), .A2(new_n22840_), .ZN(new_n22841_));
  XOR2_X1    g22775(.A1(new_n22841_), .A2(new_n65_), .Z(new_n22842_));
  NAND3_X1   g22776(.A1(new_n22837_), .A2(new_n22835_), .A3(new_n22842_), .ZN(new_n22843_));
  NAND2_X1   g22777(.A1(new_n22442_), .A2(new_n22833_), .ZN(new_n22844_));
  NAND2_X1   g22778(.A1(new_n22831_), .A2(new_n22447_), .ZN(new_n22845_));
  AOI21_X1   g22779(.A1(new_n22844_), .A2(new_n22845_), .B(new_n22439_), .ZN(new_n22846_));
  NAND2_X1   g22780(.A1(new_n22831_), .A2(new_n22833_), .ZN(new_n22847_));
  AOI21_X1   g22781(.A1(new_n22449_), .A2(new_n22847_), .B(new_n22438_), .ZN(new_n22848_));
  INV_X1     g22782(.I(new_n22842_), .ZN(new_n22849_));
  OAI21_X1   g22783(.A1(new_n22846_), .A2(new_n22848_), .B(new_n22849_), .ZN(new_n22850_));
  NAND2_X1   g22784(.A1(new_n22850_), .A2(new_n22843_), .ZN(new_n22851_));
  OAI21_X1   g22785(.A1(new_n22827_), .A2(new_n22696_), .B(new_n22851_), .ZN(new_n22852_));
  INV_X1     g22786(.I(new_n22696_), .ZN(new_n22853_));
  INV_X1     g22787(.I(new_n22758_), .ZN(new_n22854_));
  INV_X1     g22788(.I(new_n22776_), .ZN(new_n22855_));
  INV_X1     g22789(.I(new_n22782_), .ZN(new_n22856_));
  AOI21_X1   g22790(.A1(new_n22855_), .A2(new_n22777_), .B(new_n22856_), .ZN(new_n22857_));
  NAND3_X1   g22791(.A1(new_n22855_), .A2(new_n22777_), .A3(new_n22856_), .ZN(new_n22858_));
  OAI21_X1   g22792(.A1(new_n22854_), .A2(new_n22857_), .B(new_n22858_), .ZN(new_n22859_));
  INV_X1     g22793(.I(new_n22821_), .ZN(new_n22860_));
  NAND2_X1   g22794(.A1(new_n22695_), .A2(new_n22694_), .ZN(new_n22861_));
  NAND2_X1   g22795(.A1(new_n22822_), .A2(new_n22693_), .ZN(new_n22862_));
  AOI21_X1   g22796(.A1(new_n22861_), .A2(new_n22862_), .B(new_n22817_), .ZN(new_n22863_));
  OAI21_X1   g22797(.A1(new_n22860_), .A2(new_n22859_), .B(new_n22863_), .ZN(new_n22864_));
  OAI21_X1   g22798(.A1(new_n22846_), .A2(new_n22848_), .B(new_n22842_), .ZN(new_n22865_));
  NAND3_X1   g22799(.A1(new_n22837_), .A2(new_n22835_), .A3(new_n22849_), .ZN(new_n22866_));
  NAND2_X1   g22800(.A1(new_n22865_), .A2(new_n22866_), .ZN(new_n22867_));
  NAND3_X1   g22801(.A1(new_n22864_), .A2(new_n22853_), .A3(new_n22867_), .ZN(new_n22868_));
  NAND3_X1   g22802(.A1(new_n22852_), .A2(new_n22868_), .A3(new_n22689_), .ZN(new_n22869_));
  AOI22_X1   g22803(.A1(new_n22864_), .A2(new_n22853_), .B1(new_n22843_), .B2(new_n22850_), .ZN(new_n22870_));
  AOI21_X1   g22804(.A1(new_n22837_), .A2(new_n22835_), .B(new_n22849_), .ZN(new_n22871_));
  NOR3_X1    g22805(.A1(new_n22846_), .A2(new_n22848_), .A3(new_n22842_), .ZN(new_n22872_));
  NOR2_X1    g22806(.A1(new_n22871_), .A2(new_n22872_), .ZN(new_n22873_));
  NOR3_X1    g22807(.A1(new_n22827_), .A2(new_n22696_), .A3(new_n22873_), .ZN(new_n22874_));
  OAI21_X1   g22808(.A1(new_n22870_), .A2(new_n22874_), .B(new_n22688_), .ZN(new_n22875_));
  NAND2_X1   g22809(.A1(new_n22875_), .A2(new_n22869_), .ZN(new_n22876_));
  NAND2_X1   g22810(.A1(new_n22876_), .A2(new_n22688_), .ZN(new_n22877_));
  NAND2_X1   g22811(.A1(new_n17798_), .A2(new_n9488_), .ZN(new_n22878_));
  NAND2_X1   g22812(.A1(new_n17802_), .A2(new_n9503_), .ZN(new_n22879_));
  AOI21_X1   g22813(.A1(new_n19365_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n22880_));
  NAND4_X1   g22814(.A1(new_n21454_), .A2(new_n22878_), .A3(new_n22879_), .A4(new_n22880_), .ZN(new_n22881_));
  XOR2_X1    g22815(.A1(new_n22881_), .A2(\a[2] ), .Z(new_n22882_));
  NAND2_X1   g22816(.A1(new_n17802_), .A2(new_n9488_), .ZN(new_n22883_));
  NAND2_X1   g22817(.A1(new_n19365_), .A2(new_n9503_), .ZN(new_n22884_));
  AOI21_X1   g22818(.A1(new_n19359_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n22885_));
  NAND4_X1   g22819(.A1(new_n19951_), .A2(new_n22883_), .A3(new_n22884_), .A4(new_n22885_), .ZN(new_n22886_));
  XOR2_X1    g22820(.A1(new_n22886_), .A2(\a[2] ), .Z(new_n22887_));
  INV_X1     g22821(.I(new_n22887_), .ZN(new_n22888_));
  NAND2_X1   g22822(.A1(new_n19365_), .A2(new_n9488_), .ZN(new_n22889_));
  NAND2_X1   g22823(.A1(new_n19359_), .A2(new_n9503_), .ZN(new_n22890_));
  AOI21_X1   g22824(.A1(new_n17807_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n22891_));
  NAND4_X1   g22825(.A1(new_n19538_), .A2(new_n22889_), .A3(new_n22890_), .A4(new_n22891_), .ZN(new_n22892_));
  XOR2_X1    g22826(.A1(new_n22892_), .A2(\a[2] ), .Z(new_n22893_));
  INV_X1     g22827(.I(new_n22893_), .ZN(new_n22894_));
  AOI21_X1   g22828(.A1(new_n19321_), .A2(new_n6925_), .B(new_n9482_), .ZN(new_n22895_));
  OAI21_X1   g22829(.A1(new_n17828_), .A2(new_n9483_), .B(new_n22895_), .ZN(new_n22896_));
  AOI21_X1   g22830(.A1(new_n9488_), .A2(new_n19349_), .B(new_n22896_), .ZN(new_n22897_));
  NAND2_X1   g22831(.A1(new_n19760_), .A2(new_n22897_), .ZN(new_n22898_));
  XOR2_X1    g22832(.A1(new_n22898_), .A2(new_n4387_), .Z(new_n22899_));
  AOI21_X1   g22833(.A1(new_n19640_), .A2(new_n19642_), .B(new_n19320_), .ZN(new_n22900_));
  INV_X1     g22834(.I(new_n19646_), .ZN(new_n22901_));
  NOR2_X1    g22835(.A1(new_n19304_), .A2(new_n9483_), .ZN(new_n22902_));
  NOR2_X1    g22836(.A1(new_n19320_), .A2(new_n9489_), .ZN(new_n22903_));
  NOR2_X1    g22837(.A1(new_n17849_), .A2(new_n9485_), .ZN(new_n22904_));
  NOR4_X1    g22838(.A1(new_n22902_), .A2(new_n9482_), .A3(new_n22903_), .A4(new_n22904_), .ZN(new_n22905_));
  OAI21_X1   g22839(.A1(new_n22901_), .A2(new_n22900_), .B(new_n22905_), .ZN(new_n22906_));
  NAND2_X1   g22840(.A1(new_n22906_), .A2(\a[2] ), .ZN(new_n22907_));
  NAND3_X1   g22841(.A1(new_n19647_), .A2(new_n4387_), .A3(new_n22905_), .ZN(new_n22908_));
  NAND2_X1   g22842(.A1(new_n22907_), .A2(new_n22908_), .ZN(new_n22909_));
  NOR2_X1    g22843(.A1(new_n19313_), .A2(new_n6833_), .ZN(new_n22910_));
  INV_X1     g22844(.I(new_n22910_), .ZN(new_n22911_));
  AOI21_X1   g22845(.A1(new_n19563_), .A2(new_n19561_), .B(new_n9617_), .ZN(new_n22912_));
  NAND3_X1   g22846(.A1(new_n19592_), .A2(new_n19591_), .A3(new_n9613_), .ZN(new_n22913_));
  NAND2_X1   g22847(.A1(new_n19545_), .A2(new_n18637_), .ZN(new_n22914_));
  AOI21_X1   g22848(.A1(new_n19308_), .A2(new_n9503_), .B(new_n22914_), .ZN(new_n22915_));
  OAI21_X1   g22849(.A1(new_n9485_), .A2(new_n19313_), .B(new_n22915_), .ZN(new_n22916_));
  NOR2_X1    g22850(.A1(new_n19272_), .A2(new_n9623_), .ZN(new_n22917_));
  NOR3_X1    g22851(.A1(new_n19313_), .A2(new_n22917_), .A3(new_n18641_), .ZN(new_n22918_));
  NAND3_X1   g22852(.A1(new_n22913_), .A2(new_n22916_), .A3(new_n22918_), .ZN(new_n22919_));
  NOR3_X1    g22853(.A1(new_n22919_), .A2(new_n22912_), .A3(new_n22911_), .ZN(new_n22920_));
  AOI21_X1   g22854(.A1(new_n19545_), .A2(new_n9503_), .B(new_n9482_), .ZN(new_n22921_));
  OAI21_X1   g22855(.A1(new_n17849_), .A2(new_n9489_), .B(new_n22921_), .ZN(new_n22922_));
  AOI21_X1   g22856(.A1(new_n19308_), .A2(new_n6925_), .B(new_n22922_), .ZN(new_n22923_));
  OAI21_X1   g22857(.A1(new_n22244_), .A2(new_n19551_), .B(new_n22923_), .ZN(new_n22924_));
  NAND2_X1   g22858(.A1(new_n22924_), .A2(\a[2] ), .ZN(new_n22925_));
  NAND3_X1   g22859(.A1(new_n19553_), .A2(new_n4387_), .A3(new_n22923_), .ZN(new_n22926_));
  OAI21_X1   g22860(.A1(new_n22919_), .A2(new_n22912_), .B(new_n22911_), .ZN(new_n22927_));
  AOI21_X1   g22861(.A1(new_n22925_), .A2(new_n22926_), .B(new_n22927_), .ZN(new_n22928_));
  AOI22_X1   g22862(.A1(new_n17850_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n19545_), .ZN(new_n22929_));
  INV_X1     g22863(.I(new_n22929_), .ZN(new_n22930_));
  NAND2_X1   g22864(.A1(new_n19305_), .A2(new_n9488_), .ZN(new_n22931_));
  AOI21_X1   g22865(.A1(new_n22931_), .A2(new_n22930_), .B(new_n9482_), .ZN(new_n22932_));
  OAI21_X1   g22866(.A1(new_n19614_), .A2(new_n19617_), .B(new_n22932_), .ZN(new_n22933_));
  NOR2_X1    g22867(.A1(new_n22933_), .A2(\a[2] ), .ZN(new_n22934_));
  AOI21_X1   g22868(.A1(new_n19607_), .A2(new_n22932_), .B(new_n4387_), .ZN(new_n22935_));
  OAI22_X1   g22869(.A1(new_n22920_), .A2(new_n22928_), .B1(new_n22935_), .B2(new_n22934_), .ZN(new_n22936_));
  NAND2_X1   g22870(.A1(new_n19564_), .A2(new_n9613_), .ZN(new_n22937_));
  INV_X1     g22871(.I(new_n22919_), .ZN(new_n22938_));
  NAND3_X1   g22872(.A1(new_n22938_), .A2(new_n22937_), .A3(new_n22910_), .ZN(new_n22939_));
  AOI21_X1   g22873(.A1(new_n19553_), .A2(new_n22923_), .B(new_n4387_), .ZN(new_n22940_));
  NOR2_X1    g22874(.A1(new_n22924_), .A2(\a[2] ), .ZN(new_n22941_));
  NOR2_X1    g22875(.A1(new_n22940_), .A2(new_n22941_), .ZN(new_n22942_));
  OAI21_X1   g22876(.A1(new_n22942_), .A2(new_n22927_), .B(new_n22939_), .ZN(new_n22943_));
  NAND3_X1   g22877(.A1(new_n19607_), .A2(new_n4387_), .A3(new_n22932_), .ZN(new_n22944_));
  NAND2_X1   g22878(.A1(new_n22933_), .A2(\a[2] ), .ZN(new_n22945_));
  NAND2_X1   g22879(.A1(new_n22944_), .A2(new_n22945_), .ZN(new_n22946_));
  NAND2_X1   g22880(.A1(new_n19290_), .A2(new_n8799_), .ZN(new_n22947_));
  NOR2_X1    g22881(.A1(new_n6833_), .A2(new_n6834_), .ZN(new_n22948_));
  NAND3_X1   g22882(.A1(new_n19577_), .A2(new_n22947_), .A3(new_n22948_), .ZN(new_n22949_));
  NOR3_X1    g22883(.A1(new_n22949_), .A2(new_n65_), .A3(new_n22910_), .ZN(new_n22950_));
  INV_X1     g22884(.I(new_n22950_), .ZN(new_n22951_));
  NOR2_X1    g22885(.A1(new_n22949_), .A2(\a[5] ), .ZN(new_n22952_));
  NAND2_X1   g22886(.A1(new_n22947_), .A2(new_n22948_), .ZN(new_n22953_));
  NOR2_X1    g22887(.A1(new_n19593_), .A2(new_n22953_), .ZN(new_n22954_));
  NOR2_X1    g22888(.A1(new_n22954_), .A2(new_n65_), .ZN(new_n22955_));
  NAND2_X1   g22889(.A1(new_n22911_), .A2(\a[5] ), .ZN(new_n22956_));
  OAI21_X1   g22890(.A1(new_n22952_), .A2(new_n22955_), .B(new_n22956_), .ZN(new_n22957_));
  NAND2_X1   g22891(.A1(new_n22957_), .A2(new_n22951_), .ZN(new_n22958_));
  OAI21_X1   g22892(.A1(new_n22946_), .A2(new_n22943_), .B(new_n22958_), .ZN(new_n22959_));
  NAND3_X1   g22893(.A1(new_n22959_), .A2(new_n22909_), .A3(new_n22936_), .ZN(new_n22960_));
  AOI21_X1   g22894(.A1(new_n19647_), .A2(new_n22905_), .B(new_n4387_), .ZN(new_n22961_));
  NOR2_X1    g22895(.A1(new_n22906_), .A2(\a[2] ), .ZN(new_n22962_));
  NOR2_X1    g22896(.A1(new_n22962_), .A2(new_n22961_), .ZN(new_n22963_));
  NAND2_X1   g22897(.A1(new_n22926_), .A2(new_n22925_), .ZN(new_n22964_));
  INV_X1     g22898(.I(new_n22927_), .ZN(new_n22965_));
  AOI21_X1   g22899(.A1(new_n22964_), .A2(new_n22965_), .B(new_n22920_), .ZN(new_n22966_));
  NOR2_X1    g22900(.A1(new_n22935_), .A2(new_n22934_), .ZN(new_n22967_));
  NOR2_X1    g22901(.A1(new_n22967_), .A2(new_n22966_), .ZN(new_n22968_));
  NAND2_X1   g22902(.A1(new_n22954_), .A2(new_n65_), .ZN(new_n22969_));
  NAND2_X1   g22903(.A1(new_n22949_), .A2(\a[5] ), .ZN(new_n22970_));
  AOI22_X1   g22904(.A1(new_n22970_), .A2(new_n22969_), .B1(\a[5] ), .B2(new_n22911_), .ZN(new_n22971_));
  NOR2_X1    g22905(.A1(new_n22971_), .A2(new_n22950_), .ZN(new_n22972_));
  AOI21_X1   g22906(.A1(new_n22967_), .A2(new_n22966_), .B(new_n22972_), .ZN(new_n22973_));
  OAI21_X1   g22907(.A1(new_n22973_), .A2(new_n22968_), .B(new_n22963_), .ZN(new_n22974_));
  NOR2_X1    g22908(.A1(new_n19272_), .A2(new_n6843_), .ZN(new_n22975_));
  NOR2_X1    g22909(.A1(new_n19313_), .A2(new_n6913_), .ZN(new_n22976_));
  OAI22_X1   g22910(.A1(new_n22976_), .A2(new_n22975_), .B1(new_n6839_), .B2(new_n19275_), .ZN(new_n22977_));
  NAND3_X1   g22911(.A1(new_n19564_), .A2(new_n6835_), .A3(new_n22977_), .ZN(new_n22978_));
  XOR2_X1    g22912(.A1(new_n22978_), .A2(\a[5] ), .Z(new_n22979_));
  XOR2_X1    g22913(.A1(new_n22979_), .A2(new_n22951_), .Z(new_n22980_));
  AOI22_X1   g22914(.A1(new_n22974_), .A2(new_n22960_), .B1(new_n22909_), .B2(new_n22980_), .ZN(new_n22981_));
  OAI22_X1   g22915(.A1(new_n19304_), .A2(new_n9485_), .B1(new_n9483_), .B2(new_n19320_), .ZN(new_n22982_));
  NAND2_X1   g22916(.A1(new_n17827_), .A2(new_n9488_), .ZN(new_n22983_));
  AOI21_X1   g22917(.A1(new_n22983_), .A2(new_n22982_), .B(new_n9482_), .ZN(new_n22984_));
  OAI21_X1   g22918(.A1(new_n19679_), .A2(new_n19682_), .B(new_n22984_), .ZN(new_n22985_));
  NOR2_X1    g22919(.A1(new_n22985_), .A2(\a[2] ), .ZN(new_n22986_));
  INV_X1     g22920(.I(new_n22986_), .ZN(new_n22987_));
  NAND2_X1   g22921(.A1(new_n22985_), .A2(\a[2] ), .ZN(new_n22988_));
  NAND2_X1   g22922(.A1(new_n22987_), .A2(new_n22988_), .ZN(new_n22989_));
  NAND2_X1   g22923(.A1(new_n22981_), .A2(new_n22989_), .ZN(new_n22990_));
  OAI21_X1   g22924(.A1(new_n22973_), .A2(new_n22968_), .B(new_n22963_), .ZN(new_n22991_));
  NOR3_X1    g22925(.A1(new_n22973_), .A2(new_n22968_), .A3(new_n22963_), .ZN(new_n22992_));
  AOI21_X1   g22926(.A1(new_n22959_), .A2(new_n22936_), .B(new_n22909_), .ZN(new_n22993_));
  XOR2_X1    g22927(.A1(new_n22979_), .A2(new_n22950_), .Z(new_n22994_));
  OAI21_X1   g22928(.A1(new_n22992_), .A2(new_n22993_), .B(new_n22994_), .ZN(new_n22995_));
  AOI21_X1   g22929(.A1(new_n22297_), .A2(new_n22984_), .B(new_n4387_), .ZN(new_n22996_));
  OAI22_X1   g22930(.A1(new_n19272_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n19275_), .ZN(new_n22997_));
  NAND2_X1   g22931(.A1(new_n17850_), .A2(new_n6838_), .ZN(new_n22998_));
  AOI21_X1   g22932(.A1(new_n22997_), .A2(new_n22998_), .B(new_n6836_), .ZN(new_n22999_));
  NAND3_X1   g22933(.A1(new_n19553_), .A2(new_n65_), .A3(new_n22999_), .ZN(new_n23000_));
  NAND2_X1   g22934(.A1(new_n19553_), .A2(new_n22999_), .ZN(new_n23001_));
  NAND2_X1   g22935(.A1(new_n23001_), .A2(\a[5] ), .ZN(new_n23002_));
  NAND2_X1   g22936(.A1(new_n23002_), .A2(new_n23000_), .ZN(new_n23003_));
  INV_X1     g22937(.I(new_n23003_), .ZN(new_n23004_));
  INV_X1     g22938(.I(new_n22977_), .ZN(new_n23005_));
  NOR3_X1    g22939(.A1(new_n23005_), .A2(new_n19571_), .A3(new_n6836_), .ZN(new_n23006_));
  NOR4_X1    g22940(.A1(new_n23006_), .A2(new_n65_), .A3(new_n22910_), .A4(new_n22949_), .ZN(new_n23007_));
  NOR2_X1    g22941(.A1(new_n23007_), .A2(new_n22706_), .ZN(new_n23008_));
  INV_X1     g22942(.I(new_n22706_), .ZN(new_n23009_));
  NAND4_X1   g22943(.A1(new_n22978_), .A2(\a[5] ), .A3(new_n22911_), .A4(new_n22954_), .ZN(new_n23010_));
  NOR2_X1    g22944(.A1(new_n23010_), .A2(new_n23009_), .ZN(new_n23011_));
  NOR3_X1    g22945(.A1(new_n23004_), .A2(new_n23008_), .A3(new_n23011_), .ZN(new_n23012_));
  NAND2_X1   g22946(.A1(new_n23010_), .A2(new_n23009_), .ZN(new_n23013_));
  NAND2_X1   g22947(.A1(new_n23007_), .A2(new_n22706_), .ZN(new_n23014_));
  AOI21_X1   g22948(.A1(new_n23014_), .A2(new_n23013_), .B(new_n23003_), .ZN(new_n23015_));
  NOR2_X1    g22949(.A1(new_n23012_), .A2(new_n23015_), .ZN(new_n23016_));
  NOR3_X1    g22950(.A1(new_n23016_), .A2(new_n22996_), .A3(new_n22986_), .ZN(new_n23017_));
  NAND3_X1   g22951(.A1(new_n22995_), .A2(new_n22991_), .A3(new_n23017_), .ZN(new_n23018_));
  NAND3_X1   g22952(.A1(new_n22990_), .A2(new_n23018_), .A3(new_n22899_), .ZN(new_n23019_));
  XOR2_X1    g22953(.A1(new_n22898_), .A2(\a[2] ), .Z(new_n23020_));
  AOI22_X1   g22954(.A1(new_n22995_), .A2(new_n22991_), .B1(new_n22987_), .B2(new_n22988_), .ZN(new_n23021_));
  NAND3_X1   g22955(.A1(new_n23014_), .A2(new_n23003_), .A3(new_n23013_), .ZN(new_n23022_));
  OAI21_X1   g22956(.A1(new_n23008_), .A2(new_n23011_), .B(new_n23004_), .ZN(new_n23023_));
  NAND2_X1   g22957(.A1(new_n23023_), .A2(new_n23022_), .ZN(new_n23024_));
  NAND3_X1   g22958(.A1(new_n23024_), .A2(new_n22987_), .A3(new_n22988_), .ZN(new_n23025_));
  NOR2_X1    g22959(.A1(new_n22981_), .A2(new_n23025_), .ZN(new_n23026_));
  OAI21_X1   g22960(.A1(new_n23021_), .A2(new_n23026_), .B(new_n23020_), .ZN(new_n23027_));
  NAND2_X1   g22961(.A1(new_n23003_), .A2(new_n23009_), .ZN(new_n23028_));
  NOR2_X1    g22962(.A1(new_n23003_), .A2(new_n23009_), .ZN(new_n23029_));
  OAI21_X1   g22963(.A1(new_n23007_), .A2(new_n23029_), .B(new_n23028_), .ZN(new_n23030_));
  INV_X1     g22964(.I(new_n23030_), .ZN(new_n23031_));
  XOR2_X1    g22965(.A1(new_n22704_), .A2(\a[8] ), .Z(new_n23032_));
  NOR2_X1    g22966(.A1(new_n22706_), .A2(new_n4009_), .ZN(new_n23033_));
  NOR2_X1    g22967(.A1(new_n23032_), .A2(new_n23033_), .ZN(new_n23034_));
  XOR2_X1    g22968(.A1(new_n22704_), .A2(new_n4009_), .Z(new_n23035_));
  INV_X1     g22969(.I(new_n23033_), .ZN(new_n23036_));
  NOR2_X1    g22970(.A1(new_n23035_), .A2(new_n23036_), .ZN(new_n23037_));
  NOR2_X1    g22971(.A1(new_n23034_), .A2(new_n23037_), .ZN(new_n23038_));
  AOI22_X1   g22972(.A1(new_n17850_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n19545_), .ZN(new_n23039_));
  AOI21_X1   g22973(.A1(new_n19305_), .A2(new_n6838_), .B(new_n23039_), .ZN(new_n23040_));
  NOR3_X1    g22974(.A1(new_n19618_), .A2(new_n6836_), .A3(new_n23040_), .ZN(new_n23041_));
  NAND2_X1   g22975(.A1(new_n23041_), .A2(new_n65_), .ZN(new_n23042_));
  NOR2_X1    g22976(.A1(new_n23041_), .A2(new_n65_), .ZN(new_n23043_));
  INV_X1     g22977(.I(new_n23043_), .ZN(new_n23044_));
  NAND3_X1   g22978(.A1(new_n23038_), .A2(new_n23042_), .A3(new_n23044_), .ZN(new_n23045_));
  NAND2_X1   g22979(.A1(new_n23035_), .A2(new_n23036_), .ZN(new_n23046_));
  NAND2_X1   g22980(.A1(new_n23032_), .A2(new_n23033_), .ZN(new_n23047_));
  NAND2_X1   g22981(.A1(new_n23046_), .A2(new_n23047_), .ZN(new_n23048_));
  INV_X1     g22982(.I(new_n23042_), .ZN(new_n23049_));
  OAI21_X1   g22983(.A1(new_n23049_), .A2(new_n23043_), .B(new_n23048_), .ZN(new_n23050_));
  AOI21_X1   g22984(.A1(new_n23045_), .A2(new_n23050_), .B(new_n23031_), .ZN(new_n23051_));
  NAND3_X1   g22985(.A1(new_n23048_), .A2(new_n23044_), .A3(new_n23042_), .ZN(new_n23052_));
  OAI21_X1   g22986(.A1(new_n23049_), .A2(new_n23043_), .B(new_n23038_), .ZN(new_n23053_));
  AOI21_X1   g22987(.A1(new_n23053_), .A2(new_n23052_), .B(new_n23030_), .ZN(new_n23054_));
  NOR2_X1    g22988(.A1(new_n23051_), .A2(new_n23054_), .ZN(new_n23055_));
  INV_X1     g22989(.I(new_n23055_), .ZN(new_n23056_));
  AOI22_X1   g22990(.A1(new_n23027_), .A2(new_n23019_), .B1(new_n22899_), .B2(new_n23056_), .ZN(new_n23057_));
  NAND2_X1   g22991(.A1(new_n23052_), .A2(new_n23030_), .ZN(new_n23058_));
  NAND2_X1   g22992(.A1(new_n23058_), .A2(new_n23053_), .ZN(new_n23059_));
  OAI21_X1   g22993(.A1(new_n22699_), .A2(new_n22698_), .B(new_n4009_), .ZN(new_n23060_));
  NAND2_X1   g22994(.A1(new_n22700_), .A2(\a[8] ), .ZN(new_n23061_));
  NAND3_X1   g22995(.A1(new_n22704_), .A2(\a[8] ), .A3(new_n23009_), .ZN(new_n23062_));
  NAND3_X1   g22996(.A1(new_n23061_), .A2(new_n23060_), .A3(new_n23062_), .ZN(new_n23063_));
  NAND4_X1   g22997(.A1(new_n22700_), .A2(\a[8] ), .A3(new_n22704_), .A4(new_n23009_), .ZN(new_n23064_));
  NAND2_X1   g22998(.A1(new_n23063_), .A2(new_n23064_), .ZN(new_n23065_));
  INV_X1     g22999(.I(new_n23065_), .ZN(new_n23066_));
  OAI22_X1   g23000(.A1(new_n19304_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n17849_), .ZN(new_n23067_));
  NAND2_X1   g23001(.A1(new_n19321_), .A2(new_n6838_), .ZN(new_n23068_));
  AOI21_X1   g23002(.A1(new_n23067_), .A2(new_n23068_), .B(new_n6836_), .ZN(new_n23069_));
  NAND2_X1   g23003(.A1(new_n19647_), .A2(new_n23069_), .ZN(new_n23070_));
  NOR2_X1    g23004(.A1(new_n23070_), .A2(\a[5] ), .ZN(new_n23071_));
  INV_X1     g23005(.I(new_n23071_), .ZN(new_n23072_));
  NAND2_X1   g23006(.A1(new_n23070_), .A2(\a[5] ), .ZN(new_n23073_));
  NAND3_X1   g23007(.A1(new_n23066_), .A2(new_n23072_), .A3(new_n23073_), .ZN(new_n23074_));
  INV_X1     g23008(.I(new_n23073_), .ZN(new_n23075_));
  OAI21_X1   g23009(.A1(new_n23075_), .A2(new_n23071_), .B(new_n23065_), .ZN(new_n23076_));
  NAND2_X1   g23010(.A1(new_n23074_), .A2(new_n23076_), .ZN(new_n23077_));
  NAND2_X1   g23011(.A1(new_n23059_), .A2(new_n23077_), .ZN(new_n23078_));
  AOI21_X1   g23012(.A1(new_n23042_), .A2(new_n23044_), .B(new_n23048_), .ZN(new_n23079_));
  AOI21_X1   g23013(.A1(new_n23030_), .A2(new_n23052_), .B(new_n23079_), .ZN(new_n23080_));
  NOR3_X1    g23014(.A1(new_n23066_), .A2(new_n23071_), .A3(new_n23075_), .ZN(new_n23081_));
  AOI21_X1   g23015(.A1(new_n23072_), .A2(new_n23073_), .B(new_n23065_), .ZN(new_n23082_));
  OAI21_X1   g23016(.A1(new_n23081_), .A2(new_n23082_), .B(new_n23080_), .ZN(new_n23083_));
  NAND2_X1   g23017(.A1(new_n23083_), .A2(new_n23078_), .ZN(new_n23084_));
  OAI22_X1   g23018(.A1(new_n9483_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n9485_), .ZN(new_n23085_));
  NAND2_X1   g23019(.A1(new_n19350_), .A2(new_n9488_), .ZN(new_n23086_));
  AOI21_X1   g23020(.A1(new_n23085_), .A2(new_n23086_), .B(new_n9482_), .ZN(new_n23087_));
  NAND2_X1   g23021(.A1(new_n20535_), .A2(new_n23087_), .ZN(new_n23088_));
  XOR2_X1    g23022(.A1(new_n23088_), .A2(\a[2] ), .Z(new_n23089_));
  NAND2_X1   g23023(.A1(new_n23084_), .A2(new_n23089_), .ZN(new_n23090_));
  NOR2_X1    g23024(.A1(new_n23084_), .A2(new_n23089_), .ZN(new_n23091_));
  AOI21_X1   g23025(.A1(new_n23057_), .A2(new_n23090_), .B(new_n23091_), .ZN(new_n23092_));
  INV_X1     g23026(.I(new_n23081_), .ZN(new_n23093_));
  AOI21_X1   g23027(.A1(new_n23059_), .A2(new_n23093_), .B(new_n23082_), .ZN(new_n23094_));
  INV_X1     g23028(.I(new_n22342_), .ZN(new_n23095_));
  INV_X1     g23029(.I(new_n23062_), .ZN(new_n23096_));
  NAND3_X1   g23030(.A1(new_n23061_), .A2(new_n23060_), .A3(new_n23096_), .ZN(new_n23097_));
  NAND2_X1   g23031(.A1(new_n23097_), .A2(new_n23095_), .ZN(new_n23098_));
  NAND3_X1   g23032(.A1(new_n23098_), .A2(new_n22708_), .A3(new_n22714_), .ZN(new_n23099_));
  INV_X1     g23033(.I(new_n22708_), .ZN(new_n23100_));
  OAI21_X1   g23034(.A1(new_n23100_), .A2(new_n22709_), .B(new_n22715_), .ZN(new_n23101_));
  NAND2_X1   g23035(.A1(new_n23101_), .A2(new_n23099_), .ZN(new_n23102_));
  OAI22_X1   g23036(.A1(new_n19304_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n19320_), .ZN(new_n23103_));
  NAND2_X1   g23037(.A1(new_n17827_), .A2(new_n6838_), .ZN(new_n23104_));
  AOI21_X1   g23038(.A1(new_n23104_), .A2(new_n23103_), .B(new_n6836_), .ZN(new_n23105_));
  NAND3_X1   g23039(.A1(new_n22297_), .A2(new_n65_), .A3(new_n23105_), .ZN(new_n23106_));
  AOI21_X1   g23040(.A1(new_n22297_), .A2(new_n23105_), .B(new_n65_), .ZN(new_n23107_));
  INV_X1     g23041(.I(new_n23107_), .ZN(new_n23108_));
  NAND3_X1   g23042(.A1(new_n23102_), .A2(new_n23106_), .A3(new_n23108_), .ZN(new_n23109_));
  NOR3_X1    g23043(.A1(new_n23100_), .A2(new_n22709_), .A3(new_n22715_), .ZN(new_n23110_));
  AOI21_X1   g23044(.A1(new_n23098_), .A2(new_n22708_), .B(new_n22714_), .ZN(new_n23111_));
  NOR2_X1    g23045(.A1(new_n23110_), .A2(new_n23111_), .ZN(new_n23112_));
  INV_X1     g23046(.I(new_n23106_), .ZN(new_n23113_));
  OAI21_X1   g23047(.A1(new_n23113_), .A2(new_n23107_), .B(new_n23112_), .ZN(new_n23114_));
  AOI21_X1   g23048(.A1(new_n23109_), .A2(new_n23114_), .B(new_n23094_), .ZN(new_n23115_));
  INV_X1     g23049(.I(new_n23082_), .ZN(new_n23116_));
  OAI21_X1   g23050(.A1(new_n23080_), .A2(new_n23081_), .B(new_n23116_), .ZN(new_n23117_));
  NAND3_X1   g23051(.A1(new_n23112_), .A2(new_n23106_), .A3(new_n23108_), .ZN(new_n23118_));
  OAI21_X1   g23052(.A1(new_n23107_), .A2(new_n23113_), .B(new_n23102_), .ZN(new_n23119_));
  AOI21_X1   g23053(.A1(new_n23118_), .A2(new_n23119_), .B(new_n23117_), .ZN(new_n23120_));
  NOR2_X1    g23054(.A1(new_n23115_), .A2(new_n23120_), .ZN(new_n23121_));
  AOI22_X1   g23055(.A1(new_n19349_), .A2(new_n6925_), .B1(new_n9503_), .B2(new_n19350_), .ZN(new_n23122_));
  NOR2_X1    g23056(.A1(new_n17806_), .A2(new_n9489_), .ZN(new_n23123_));
  OAI21_X1   g23057(.A1(new_n23122_), .A2(new_n23123_), .B(new_n6922_), .ZN(new_n23124_));
  NOR2_X1    g23058(.A1(new_n19915_), .A2(new_n23124_), .ZN(new_n23125_));
  NAND2_X1   g23059(.A1(new_n23125_), .A2(new_n4387_), .ZN(new_n23126_));
  OAI21_X1   g23060(.A1(new_n19915_), .A2(new_n23124_), .B(\a[2] ), .ZN(new_n23127_));
  NAND2_X1   g23061(.A1(new_n23126_), .A2(new_n23127_), .ZN(new_n23128_));
  NOR2_X1    g23062(.A1(new_n23121_), .A2(new_n23128_), .ZN(new_n23129_));
  NAND2_X1   g23063(.A1(new_n23121_), .A2(new_n23128_), .ZN(new_n23130_));
  OAI21_X1   g23064(.A1(new_n23092_), .A2(new_n23129_), .B(new_n23130_), .ZN(new_n23131_));
  OAI22_X1   g23065(.A1(new_n17806_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n19346_), .ZN(new_n23132_));
  NAND2_X1   g23066(.A1(new_n19359_), .A2(new_n9488_), .ZN(new_n23133_));
  AOI21_X1   g23067(.A1(new_n23133_), .A2(new_n23132_), .B(new_n9482_), .ZN(new_n23134_));
  NAND3_X1   g23068(.A1(new_n20096_), .A2(new_n4387_), .A3(new_n23134_), .ZN(new_n23135_));
  NAND2_X1   g23069(.A1(new_n20096_), .A2(new_n23134_), .ZN(new_n23136_));
  NAND2_X1   g23070(.A1(new_n23136_), .A2(\a[2] ), .ZN(new_n23137_));
  NAND2_X1   g23071(.A1(new_n23137_), .A2(new_n23135_), .ZN(new_n23138_));
  NAND2_X1   g23072(.A1(new_n23131_), .A2(new_n23138_), .ZN(new_n23139_));
  NOR3_X1    g23073(.A1(new_n23021_), .A2(new_n23026_), .A3(new_n23020_), .ZN(new_n23140_));
  AOI21_X1   g23074(.A1(new_n22990_), .A2(new_n23018_), .B(new_n22899_), .ZN(new_n23141_));
  OAI22_X1   g23075(.A1(new_n23140_), .A2(new_n23141_), .B1(new_n23020_), .B2(new_n23055_), .ZN(new_n23142_));
  AOI21_X1   g23076(.A1(new_n23074_), .A2(new_n23076_), .B(new_n23080_), .ZN(new_n23143_));
  AOI21_X1   g23077(.A1(new_n23093_), .A2(new_n23116_), .B(new_n23059_), .ZN(new_n23144_));
  NOR2_X1    g23078(.A1(new_n23144_), .A2(new_n23143_), .ZN(new_n23145_));
  XOR2_X1    g23079(.A1(new_n23088_), .A2(new_n4387_), .Z(new_n23146_));
  NOR2_X1    g23080(.A1(new_n23145_), .A2(new_n23146_), .ZN(new_n23147_));
  NAND2_X1   g23081(.A1(new_n23145_), .A2(new_n23146_), .ZN(new_n23148_));
  OAI21_X1   g23082(.A1(new_n23142_), .A2(new_n23147_), .B(new_n23148_), .ZN(new_n23149_));
  NAND2_X1   g23083(.A1(new_n23114_), .A2(new_n23109_), .ZN(new_n23150_));
  NAND2_X1   g23084(.A1(new_n23119_), .A2(new_n23118_), .ZN(new_n23151_));
  MUX2_X1    g23085(.I0(new_n23151_), .I1(new_n23150_), .S(new_n23117_), .Z(new_n23152_));
  NAND3_X1   g23086(.A1(new_n23152_), .A2(new_n23126_), .A3(new_n23127_), .ZN(new_n23153_));
  NAND2_X1   g23087(.A1(new_n23149_), .A2(new_n23153_), .ZN(new_n23154_));
  INV_X1     g23088(.I(new_n22722_), .ZN(new_n23155_));
  INV_X1     g23089(.I(new_n22726_), .ZN(new_n23156_));
  NAND3_X1   g23090(.A1(new_n23155_), .A2(new_n22720_), .A3(new_n23156_), .ZN(new_n23157_));
  OAI22_X1   g23091(.A1(new_n17828_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n19320_), .ZN(new_n23158_));
  NAND2_X1   g23092(.A1(new_n19349_), .A2(new_n6838_), .ZN(new_n23159_));
  AOI21_X1   g23093(.A1(new_n23159_), .A2(new_n23158_), .B(new_n6836_), .ZN(new_n23160_));
  NAND2_X1   g23094(.A1(new_n19760_), .A2(new_n23160_), .ZN(new_n23161_));
  XOR2_X1    g23095(.A1(new_n23161_), .A2(new_n65_), .Z(new_n23162_));
  NAND3_X1   g23096(.A1(new_n23162_), .A2(new_n22727_), .A3(new_n23157_), .ZN(new_n23163_));
  AOI21_X1   g23097(.A1(new_n23155_), .A2(new_n22720_), .B(new_n23156_), .ZN(new_n23164_));
  NOR3_X1    g23098(.A1(new_n22721_), .A2(new_n22722_), .A3(new_n22726_), .ZN(new_n23165_));
  XOR2_X1    g23099(.A1(new_n23161_), .A2(\a[5] ), .Z(new_n23166_));
  OAI21_X1   g23100(.A1(new_n23164_), .A2(new_n23165_), .B(new_n23166_), .ZN(new_n23167_));
  NAND2_X1   g23101(.A1(new_n23167_), .A2(new_n23163_), .ZN(new_n23168_));
  NAND2_X1   g23102(.A1(new_n23117_), .A2(new_n23118_), .ZN(new_n23169_));
  NAND3_X1   g23103(.A1(new_n23168_), .A2(new_n23119_), .A3(new_n23169_), .ZN(new_n23170_));
  NAND2_X1   g23104(.A1(new_n23169_), .A2(new_n23119_), .ZN(new_n23171_));
  NAND3_X1   g23105(.A1(new_n23171_), .A2(new_n23167_), .A3(new_n23163_), .ZN(new_n23172_));
  AOI21_X1   g23106(.A1(new_n23170_), .A2(new_n23172_), .B(new_n23138_), .ZN(new_n23173_));
  NAND3_X1   g23107(.A1(new_n23154_), .A2(new_n23130_), .A3(new_n23173_), .ZN(new_n23174_));
  AOI21_X1   g23108(.A1(new_n23174_), .A2(new_n23139_), .B(new_n22894_), .ZN(new_n23175_));
  INV_X1     g23109(.I(new_n23175_), .ZN(new_n23176_));
  XOR2_X1    g23110(.A1(new_n23136_), .A2(\a[2] ), .Z(new_n23177_));
  AOI21_X1   g23111(.A1(new_n23154_), .A2(new_n23130_), .B(new_n23177_), .ZN(new_n23178_));
  AOI21_X1   g23112(.A1(new_n23163_), .A2(new_n23167_), .B(new_n23171_), .ZN(new_n23179_));
  INV_X1     g23113(.I(new_n23172_), .ZN(new_n23180_));
  OAI21_X1   g23114(.A1(new_n23180_), .A2(new_n23179_), .B(new_n23177_), .ZN(new_n23181_));
  NOR2_X1    g23115(.A1(new_n23131_), .A2(new_n23181_), .ZN(new_n23182_));
  NOR3_X1    g23116(.A1(new_n23178_), .A2(new_n23182_), .A3(new_n22893_), .ZN(new_n23183_));
  AOI21_X1   g23117(.A1(new_n23174_), .A2(new_n23139_), .B(new_n22894_), .ZN(new_n23184_));
  INV_X1     g23118(.I(new_n22337_), .ZN(new_n23185_));
  INV_X1     g23119(.I(new_n22344_), .ZN(new_n23186_));
  NAND3_X1   g23120(.A1(new_n22727_), .A2(new_n22719_), .A3(new_n22734_), .ZN(new_n23187_));
  OAI21_X1   g23121(.A1(new_n23164_), .A2(new_n22718_), .B(new_n22733_), .ZN(new_n23188_));
  AOI21_X1   g23122(.A1(new_n23188_), .A2(new_n23187_), .B(new_n23186_), .ZN(new_n23189_));
  NOR3_X1    g23123(.A1(new_n23164_), .A2(new_n22718_), .A3(new_n22733_), .ZN(new_n23190_));
  AOI21_X1   g23124(.A1(new_n22727_), .A2(new_n22719_), .B(new_n22734_), .ZN(new_n23191_));
  NOR3_X1    g23125(.A1(new_n23190_), .A2(new_n23191_), .A3(new_n22344_), .ZN(new_n23192_));
  OAI21_X1   g23126(.A1(new_n23192_), .A2(new_n23189_), .B(new_n23185_), .ZN(new_n23193_));
  OAI21_X1   g23127(.A1(new_n23190_), .A2(new_n23191_), .B(new_n22344_), .ZN(new_n23194_));
  NAND3_X1   g23128(.A1(new_n23188_), .A2(new_n23187_), .A3(new_n23186_), .ZN(new_n23195_));
  NAND3_X1   g23129(.A1(new_n23194_), .A2(new_n23195_), .A3(new_n22337_), .ZN(new_n23196_));
  NAND2_X1   g23130(.A1(new_n23193_), .A2(new_n23196_), .ZN(new_n23197_));
  NAND4_X1   g23131(.A1(new_n23167_), .A2(new_n23163_), .A3(new_n23169_), .A4(new_n23119_), .ZN(new_n23198_));
  OAI22_X1   g23132(.A1(new_n6843_), .A2(new_n19343_), .B1(new_n17828_), .B2(new_n6913_), .ZN(new_n23199_));
  NAND2_X1   g23133(.A1(new_n19350_), .A2(new_n6838_), .ZN(new_n23200_));
  AOI21_X1   g23134(.A1(new_n23199_), .A2(new_n23200_), .B(new_n6836_), .ZN(new_n23201_));
  NAND2_X1   g23135(.A1(new_n20535_), .A2(new_n23201_), .ZN(new_n23202_));
  XOR2_X1    g23136(.A1(new_n23202_), .A2(\a[5] ), .Z(new_n23203_));
  INV_X1     g23137(.I(new_n23203_), .ZN(new_n23204_));
  AOI21_X1   g23138(.A1(new_n23198_), .A2(new_n23167_), .B(new_n23204_), .ZN(new_n23205_));
  INV_X1     g23139(.I(new_n23205_), .ZN(new_n23206_));
  NAND3_X1   g23140(.A1(new_n23198_), .A2(new_n23167_), .A3(new_n23204_), .ZN(new_n23207_));
  AOI21_X1   g23141(.A1(new_n23206_), .A2(new_n23207_), .B(new_n23197_), .ZN(new_n23208_));
  AOI21_X1   g23142(.A1(new_n23194_), .A2(new_n23195_), .B(new_n22337_), .ZN(new_n23209_));
  NOR3_X1    g23143(.A1(new_n23192_), .A2(new_n23189_), .A3(new_n23185_), .ZN(new_n23210_));
  NOR2_X1    g23144(.A1(new_n23210_), .A2(new_n23209_), .ZN(new_n23211_));
  INV_X1     g23145(.I(new_n23207_), .ZN(new_n23212_));
  NOR3_X1    g23146(.A1(new_n23211_), .A2(new_n23212_), .A3(new_n23205_), .ZN(new_n23213_));
  NOR2_X1    g23147(.A1(new_n23208_), .A2(new_n23213_), .ZN(new_n23214_));
  OAI21_X1   g23148(.A1(new_n23183_), .A2(new_n23184_), .B(new_n23214_), .ZN(new_n23215_));
  NAND3_X1   g23149(.A1(new_n23215_), .A2(new_n23176_), .A3(new_n22888_), .ZN(new_n23216_));
  NAND3_X1   g23150(.A1(new_n23174_), .A2(new_n23139_), .A3(new_n22894_), .ZN(new_n23217_));
  OAI21_X1   g23151(.A1(new_n23178_), .A2(new_n23182_), .B(new_n22893_), .ZN(new_n23218_));
  OAI21_X1   g23152(.A1(new_n23205_), .A2(new_n23212_), .B(new_n23211_), .ZN(new_n23219_));
  NAND3_X1   g23153(.A1(new_n23197_), .A2(new_n23206_), .A3(new_n23207_), .ZN(new_n23220_));
  NAND2_X1   g23154(.A1(new_n23219_), .A2(new_n23220_), .ZN(new_n23221_));
  AOI22_X1   g23155(.A1(new_n23218_), .A2(new_n23217_), .B1(new_n22894_), .B2(new_n23221_), .ZN(new_n23222_));
  NAND2_X1   g23156(.A1(new_n23222_), .A2(new_n22887_), .ZN(new_n23223_));
  NAND2_X1   g23157(.A1(new_n22753_), .A2(new_n22757_), .ZN(new_n23224_));
  NAND2_X1   g23158(.A1(new_n22854_), .A2(new_n23224_), .ZN(new_n23225_));
  AOI22_X1   g23159(.A1(new_n23216_), .A2(new_n23223_), .B1(new_n23225_), .B2(new_n22888_), .ZN(new_n23226_));
  NAND2_X1   g23160(.A1(new_n23226_), .A2(new_n22882_), .ZN(new_n23227_));
  INV_X1     g23161(.I(new_n23227_), .ZN(new_n23228_));
  INV_X1     g23162(.I(new_n22882_), .ZN(new_n23229_));
  NAND2_X1   g23163(.A1(new_n23222_), .A2(new_n22887_), .ZN(new_n23230_));
  AOI21_X1   g23164(.A1(new_n23218_), .A2(new_n23217_), .B(new_n23221_), .ZN(new_n23231_));
  NOR3_X1    g23165(.A1(new_n23231_), .A2(new_n22887_), .A3(new_n23175_), .ZN(new_n23232_));
  AOI21_X1   g23166(.A1(new_n23215_), .A2(new_n23176_), .B(new_n22888_), .ZN(new_n23233_));
  INV_X1     g23167(.I(new_n23225_), .ZN(new_n23234_));
  OAI21_X1   g23168(.A1(new_n23233_), .A2(new_n23232_), .B(new_n23234_), .ZN(new_n23235_));
  NAND3_X1   g23169(.A1(new_n23235_), .A2(new_n23229_), .A3(new_n23230_), .ZN(new_n23236_));
  NAND2_X1   g23170(.A1(new_n23226_), .A2(new_n22882_), .ZN(new_n23237_));
  NAND3_X1   g23171(.A1(new_n22855_), .A2(new_n22777_), .A3(new_n22782_), .ZN(new_n23238_));
  INV_X1     g23172(.I(new_n23238_), .ZN(new_n23239_));
  AOI21_X1   g23173(.A1(new_n22855_), .A2(new_n22777_), .B(new_n22782_), .ZN(new_n23240_));
  OAI21_X1   g23174(.A1(new_n23239_), .A2(new_n23240_), .B(new_n22758_), .ZN(new_n23241_));
  OAI21_X1   g23175(.A1(new_n22784_), .A2(new_n22857_), .B(new_n22854_), .ZN(new_n23242_));
  NAND2_X1   g23176(.A1(new_n23241_), .A2(new_n23242_), .ZN(new_n23243_));
  AOI21_X1   g23177(.A1(new_n23237_), .A2(new_n23236_), .B(new_n23243_), .ZN(new_n23244_));
  AOI22_X1   g23178(.A1(new_n17798_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n17802_), .ZN(new_n23245_));
  NOR2_X1    g23179(.A1(new_n19375_), .A2(new_n9489_), .ZN(new_n23246_));
  OAI21_X1   g23180(.A1(new_n23246_), .A2(new_n23245_), .B(new_n6922_), .ZN(new_n23247_));
  NOR2_X1    g23181(.A1(new_n21753_), .A2(new_n23247_), .ZN(new_n23248_));
  XOR2_X1    g23182(.A1(new_n23248_), .A2(new_n4387_), .Z(new_n23249_));
  INV_X1     g23183(.I(new_n23249_), .ZN(new_n23250_));
  OAI21_X1   g23184(.A1(new_n23244_), .A2(new_n23228_), .B(new_n23250_), .ZN(new_n23251_));
  NOR2_X1    g23185(.A1(new_n23226_), .A2(new_n22882_), .ZN(new_n23252_));
  AOI21_X1   g23186(.A1(new_n23235_), .A2(new_n23230_), .B(new_n23229_), .ZN(new_n23253_));
  INV_X1     g23187(.I(new_n23240_), .ZN(new_n23254_));
  NAND2_X1   g23188(.A1(new_n23254_), .A2(new_n23238_), .ZN(new_n23255_));
  AOI21_X1   g23189(.A1(new_n22783_), .A2(new_n22858_), .B(new_n22758_), .ZN(new_n23256_));
  AOI21_X1   g23190(.A1(new_n23255_), .A2(new_n22758_), .B(new_n23256_), .ZN(new_n23257_));
  OAI21_X1   g23191(.A1(new_n23252_), .A2(new_n23253_), .B(new_n23257_), .ZN(new_n23258_));
  NAND2_X1   g23192(.A1(new_n22785_), .A2(new_n22860_), .ZN(new_n23259_));
  NAND2_X1   g23193(.A1(new_n22859_), .A2(new_n22821_), .ZN(new_n23260_));
  AOI21_X1   g23194(.A1(new_n23259_), .A2(new_n23260_), .B(new_n23250_), .ZN(new_n23261_));
  NAND3_X1   g23195(.A1(new_n23258_), .A2(new_n23227_), .A3(new_n23261_), .ZN(new_n23262_));
  OAI22_X1   g23196(.A1(new_n19375_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n17797_), .ZN(new_n23263_));
  NAND2_X1   g23197(.A1(new_n19386_), .A2(new_n9488_), .ZN(new_n23264_));
  AOI21_X1   g23198(.A1(new_n23264_), .A2(new_n23263_), .B(new_n9482_), .ZN(new_n23265_));
  NAND2_X1   g23199(.A1(new_n20162_), .A2(new_n23265_), .ZN(new_n23266_));
  XOR2_X1    g23200(.A1(new_n23266_), .A2(\a[2] ), .Z(new_n23267_));
  INV_X1     g23201(.I(new_n23267_), .ZN(new_n23268_));
  NOR2_X1    g23202(.A1(new_n22860_), .A2(new_n22859_), .ZN(new_n23269_));
  XOR2_X1    g23203(.A1(new_n22822_), .A2(new_n22694_), .Z(new_n23270_));
  INV_X1     g23204(.I(new_n23270_), .ZN(new_n23271_));
  OAI21_X1   g23205(.A1(new_n23269_), .A2(new_n22817_), .B(new_n23271_), .ZN(new_n23272_));
  NAND2_X1   g23206(.A1(new_n22785_), .A2(new_n22821_), .ZN(new_n23273_));
  NAND3_X1   g23207(.A1(new_n23273_), .A2(new_n22825_), .A3(new_n23270_), .ZN(new_n23274_));
  AOI21_X1   g23208(.A1(new_n23272_), .A2(new_n23274_), .B(new_n23268_), .ZN(new_n23275_));
  NAND3_X1   g23209(.A1(new_n23251_), .A2(new_n23262_), .A3(new_n23275_), .ZN(new_n23276_));
  AOI21_X1   g23210(.A1(new_n23258_), .A2(new_n23227_), .B(new_n23249_), .ZN(new_n23277_));
  NOR2_X1    g23211(.A1(new_n22859_), .A2(new_n22821_), .ZN(new_n23278_));
  NOR2_X1    g23212(.A1(new_n22785_), .A2(new_n22860_), .ZN(new_n23279_));
  OAI21_X1   g23213(.A1(new_n23279_), .A2(new_n23278_), .B(new_n23249_), .ZN(new_n23280_));
  NOR3_X1    g23214(.A1(new_n23244_), .A2(new_n23228_), .A3(new_n23280_), .ZN(new_n23281_));
  OAI21_X1   g23215(.A1(new_n23277_), .A2(new_n23281_), .B(new_n23268_), .ZN(new_n23282_));
  NAND3_X1   g23216(.A1(new_n23282_), .A2(new_n23276_), .A3(new_n22876_), .ZN(new_n23283_));
  NAND2_X1   g23217(.A1(new_n19394_), .A2(new_n9488_), .ZN(new_n23284_));
  NAND2_X1   g23218(.A1(new_n17794_), .A2(new_n9503_), .ZN(new_n23285_));
  AOI21_X1   g23219(.A1(new_n19386_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n23286_));
  NAND4_X1   g23220(.A1(new_n20291_), .A2(new_n23284_), .A3(new_n23285_), .A4(new_n23286_), .ZN(new_n23287_));
  XOR2_X1    g23221(.A1(new_n23287_), .A2(\a[2] ), .Z(new_n23288_));
  AOI21_X1   g23222(.A1(new_n23283_), .A2(new_n22877_), .B(new_n23288_), .ZN(new_n23289_));
  NOR3_X1    g23223(.A1(new_n22870_), .A2(new_n22874_), .A3(new_n22688_), .ZN(new_n23290_));
  AOI21_X1   g23224(.A1(new_n22852_), .A2(new_n22868_), .B(new_n22689_), .ZN(new_n23291_));
  NOR2_X1    g23225(.A1(new_n23290_), .A2(new_n23291_), .ZN(new_n23292_));
  NOR2_X1    g23226(.A1(new_n23292_), .A2(new_n22689_), .ZN(new_n23293_));
  AOI21_X1   g23227(.A1(new_n23273_), .A2(new_n22825_), .B(new_n23270_), .ZN(new_n23294_));
  NOR3_X1    g23228(.A1(new_n23269_), .A2(new_n23271_), .A3(new_n22817_), .ZN(new_n23295_));
  OAI21_X1   g23229(.A1(new_n23295_), .A2(new_n23294_), .B(new_n23267_), .ZN(new_n23296_));
  NOR3_X1    g23230(.A1(new_n23277_), .A2(new_n23281_), .A3(new_n23296_), .ZN(new_n23297_));
  AOI21_X1   g23231(.A1(new_n23251_), .A2(new_n23262_), .B(new_n23267_), .ZN(new_n23298_));
  NOR3_X1    g23232(.A1(new_n23298_), .A2(new_n23297_), .A3(new_n23292_), .ZN(new_n23299_));
  NAND2_X1   g23233(.A1(new_n22864_), .A2(new_n22853_), .ZN(new_n23300_));
  AOI21_X1   g23234(.A1(new_n23300_), .A2(new_n22865_), .B(new_n22872_), .ZN(new_n23301_));
  AOI22_X1   g23235(.A1(new_n17798_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n17802_), .ZN(new_n23302_));
  NOR2_X1    g23236(.A1(new_n19375_), .A2(new_n6839_), .ZN(new_n23303_));
  OAI21_X1   g23237(.A1(new_n23303_), .A2(new_n23302_), .B(new_n6835_), .ZN(new_n23304_));
  NOR2_X1    g23238(.A1(new_n21753_), .A2(new_n23304_), .ZN(new_n23305_));
  XOR2_X1    g23239(.A1(new_n23305_), .A2(new_n65_), .Z(new_n23306_));
  INV_X1     g23240(.I(new_n23306_), .ZN(new_n23307_));
  INV_X1     g23241(.I(new_n22418_), .ZN(new_n23308_));
  INV_X1     g23242(.I(new_n22423_), .ZN(new_n23309_));
  NOR3_X1    g23243(.A1(new_n23308_), .A2(new_n22416_), .A3(new_n23309_), .ZN(new_n23310_));
  AOI21_X1   g23244(.A1(new_n22438_), .A2(new_n22847_), .B(new_n22836_), .ZN(new_n23311_));
  OAI21_X1   g23245(.A1(new_n23310_), .A2(new_n22451_), .B(new_n23311_), .ZN(new_n23312_));
  OAI21_X1   g23246(.A1(new_n23308_), .A2(new_n22416_), .B(new_n23309_), .ZN(new_n23313_));
  NAND3_X1   g23247(.A1(new_n23313_), .A2(new_n22424_), .A3(new_n22450_), .ZN(new_n23314_));
  AOI21_X1   g23248(.A1(new_n23312_), .A2(new_n23314_), .B(new_n23307_), .ZN(new_n23315_));
  AOI21_X1   g23249(.A1(new_n23313_), .A2(new_n22424_), .B(new_n22450_), .ZN(new_n23316_));
  NOR3_X1    g23250(.A1(new_n23310_), .A2(new_n22451_), .A3(new_n23311_), .ZN(new_n23317_));
  NOR3_X1    g23251(.A1(new_n23317_), .A2(new_n23316_), .A3(new_n23306_), .ZN(new_n23318_));
  NOR2_X1    g23252(.A1(new_n23318_), .A2(new_n23315_), .ZN(new_n23319_));
  INV_X1     g23253(.I(new_n23319_), .ZN(new_n23320_));
  NAND2_X1   g23254(.A1(new_n23301_), .A2(new_n23320_), .ZN(new_n23321_));
  INV_X1     g23255(.I(new_n23321_), .ZN(new_n23322_));
  NOR2_X1    g23256(.A1(new_n23301_), .A2(new_n23320_), .ZN(new_n23323_));
  OAI21_X1   g23257(.A1(new_n23322_), .A2(new_n23323_), .B(new_n23288_), .ZN(new_n23324_));
  NOR3_X1    g23258(.A1(new_n23299_), .A2(new_n23324_), .A3(new_n23293_), .ZN(new_n23325_));
  NOR3_X1    g23259(.A1(new_n23325_), .A2(new_n23289_), .A3(new_n22684_), .ZN(new_n23326_));
  INV_X1     g23260(.I(new_n22684_), .ZN(new_n23327_));
  INV_X1     g23261(.I(new_n23288_), .ZN(new_n23328_));
  OAI21_X1   g23262(.A1(new_n23299_), .A2(new_n23293_), .B(new_n23328_), .ZN(new_n23329_));
  OAI21_X1   g23263(.A1(new_n22827_), .A2(new_n22696_), .B(new_n22865_), .ZN(new_n23330_));
  NAND2_X1   g23264(.A1(new_n23330_), .A2(new_n22866_), .ZN(new_n23331_));
  NAND2_X1   g23265(.A1(new_n23331_), .A2(new_n23319_), .ZN(new_n23332_));
  AOI21_X1   g23266(.A1(new_n23332_), .A2(new_n23321_), .B(new_n23328_), .ZN(new_n23333_));
  NAND3_X1   g23267(.A1(new_n23283_), .A2(new_n22877_), .A3(new_n23333_), .ZN(new_n23334_));
  AOI21_X1   g23268(.A1(new_n23329_), .A2(new_n23334_), .B(new_n23327_), .ZN(new_n23335_));
  NOR2_X1    g23269(.A1(new_n22414_), .A2(new_n22413_), .ZN(new_n23336_));
  INV_X1     g23270(.I(new_n23336_), .ZN(new_n23337_));
  XOR2_X1    g23271(.A1(new_n22452_), .A2(new_n22242_), .Z(new_n23338_));
  NOR2_X1    g23272(.A1(new_n23338_), .A2(new_n23337_), .ZN(new_n23339_));
  XOR2_X1    g23273(.A1(new_n22452_), .A2(new_n22243_), .Z(new_n23340_));
  NOR2_X1    g23274(.A1(new_n23340_), .A2(new_n23336_), .ZN(new_n23341_));
  OAI22_X1   g23275(.A1(new_n19375_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n17797_), .ZN(new_n23342_));
  NAND2_X1   g23276(.A1(new_n19386_), .A2(new_n6838_), .ZN(new_n23343_));
  AOI21_X1   g23277(.A1(new_n23343_), .A2(new_n23342_), .B(new_n6836_), .ZN(new_n23344_));
  NAND2_X1   g23278(.A1(new_n20162_), .A2(new_n23344_), .ZN(new_n23345_));
  XOR2_X1    g23279(.A1(new_n23345_), .A2(\a[5] ), .Z(new_n23346_));
  NOR3_X1    g23280(.A1(new_n23339_), .A2(new_n23341_), .A3(new_n23346_), .ZN(new_n23347_));
  NAND2_X1   g23281(.A1(new_n23340_), .A2(new_n23336_), .ZN(new_n23348_));
  NAND2_X1   g23282(.A1(new_n23338_), .A2(new_n23337_), .ZN(new_n23349_));
  INV_X1     g23283(.I(new_n23346_), .ZN(new_n23350_));
  AOI21_X1   g23284(.A1(new_n23348_), .A2(new_n23349_), .B(new_n23350_), .ZN(new_n23351_));
  AOI21_X1   g23285(.A1(new_n23301_), .A2(new_n23319_), .B(new_n23315_), .ZN(new_n23352_));
  INV_X1     g23286(.I(new_n23352_), .ZN(new_n23353_));
  NOR3_X1    g23287(.A1(new_n23353_), .A2(new_n23347_), .A3(new_n23351_), .ZN(new_n23354_));
  INV_X1     g23288(.I(new_n23347_), .ZN(new_n23355_));
  OAI21_X1   g23289(.A1(new_n23339_), .A2(new_n23341_), .B(new_n23346_), .ZN(new_n23356_));
  AOI21_X1   g23290(.A1(new_n23355_), .A2(new_n23356_), .B(new_n23352_), .ZN(new_n23357_));
  NOR2_X1    g23291(.A1(new_n23357_), .A2(new_n23354_), .ZN(new_n23358_));
  OAI22_X1   g23292(.A1(new_n23326_), .A2(new_n23335_), .B1(new_n23358_), .B2(new_n22684_), .ZN(new_n23359_));
  NAND2_X1   g23293(.A1(new_n23359_), .A2(new_n22679_), .ZN(new_n23360_));
  NAND3_X1   g23294(.A1(new_n23329_), .A2(new_n23334_), .A3(new_n23327_), .ZN(new_n23361_));
  OAI21_X1   g23295(.A1(new_n23325_), .A2(new_n23289_), .B(new_n22684_), .ZN(new_n23362_));
  INV_X1     g23296(.I(new_n23358_), .ZN(new_n23363_));
  AOI22_X1   g23297(.A1(new_n23362_), .A2(new_n23361_), .B1(new_n23327_), .B2(new_n23363_), .ZN(new_n23364_));
  NAND2_X1   g23298(.A1(new_n23364_), .A2(new_n22678_), .ZN(new_n23365_));
  XOR2_X1    g23299(.A1(new_n22453_), .A2(new_n22485_), .Z(new_n23366_));
  XOR2_X1    g23300(.A1(new_n23366_), .A2(new_n22459_), .Z(new_n23367_));
  INV_X1     g23301(.I(new_n23367_), .ZN(new_n23368_));
  NOR2_X1    g23302(.A1(new_n23351_), .A2(new_n23347_), .ZN(new_n23369_));
  AOI22_X1   g23303(.A1(new_n19386_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n20127_), .ZN(new_n23370_));
  NOR2_X1    g23304(.A1(new_n17793_), .A2(new_n6839_), .ZN(new_n23371_));
  OAI21_X1   g23305(.A1(new_n23370_), .A2(new_n23371_), .B(new_n6835_), .ZN(new_n23372_));
  NOR2_X1    g23306(.A1(new_n21632_), .A2(new_n23372_), .ZN(new_n23373_));
  XOR2_X1    g23307(.A1(new_n23373_), .A2(new_n65_), .Z(new_n23374_));
  INV_X1     g23308(.I(new_n23374_), .ZN(new_n23375_));
  AOI21_X1   g23309(.A1(new_n23369_), .A2(new_n23353_), .B(new_n23375_), .ZN(new_n23376_));
  INV_X1     g23310(.I(new_n23376_), .ZN(new_n23377_));
  NAND3_X1   g23311(.A1(new_n23369_), .A2(new_n23353_), .A3(new_n23375_), .ZN(new_n23378_));
  AOI21_X1   g23312(.A1(new_n23377_), .A2(new_n23378_), .B(new_n23368_), .ZN(new_n23379_));
  INV_X1     g23313(.I(new_n23378_), .ZN(new_n23380_));
  NOR3_X1    g23314(.A1(new_n23380_), .A2(new_n23367_), .A3(new_n23376_), .ZN(new_n23381_));
  NOR2_X1    g23315(.A1(new_n23379_), .A2(new_n23381_), .ZN(new_n23382_));
  INV_X1     g23316(.I(new_n23382_), .ZN(new_n23383_));
  AOI21_X1   g23317(.A1(new_n23360_), .A2(new_n23365_), .B(new_n23383_), .ZN(new_n23384_));
  OAI21_X1   g23318(.A1(new_n22679_), .A2(new_n23359_), .B(new_n22671_), .ZN(new_n23385_));
  OAI21_X1   g23319(.A1(new_n23384_), .A2(new_n23385_), .B(new_n22672_), .ZN(new_n23386_));
  OAI22_X1   g23320(.A1(new_n19410_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n17789_), .ZN(new_n23387_));
  NAND2_X1   g23321(.A1(new_n19415_), .A2(new_n9488_), .ZN(new_n23388_));
  AOI21_X1   g23322(.A1(new_n23388_), .A2(new_n23387_), .B(new_n9482_), .ZN(new_n23389_));
  NAND2_X1   g23323(.A1(new_n20846_), .A2(new_n23389_), .ZN(new_n23390_));
  XOR2_X1    g23324(.A1(new_n23390_), .A2(\a[2] ), .Z(new_n23391_));
  INV_X1     g23325(.I(new_n23391_), .ZN(new_n23392_));
  INV_X1     g23326(.I(new_n22545_), .ZN(new_n23393_));
  XOR2_X1    g23327(.A1(new_n22591_), .A2(new_n23393_), .Z(new_n23394_));
  XOR2_X1    g23328(.A1(new_n22591_), .A2(new_n23393_), .Z(new_n23395_));
  NAND2_X1   g23329(.A1(new_n23395_), .A2(new_n22549_), .ZN(new_n23396_));
  OAI21_X1   g23330(.A1(new_n22549_), .A2(new_n23394_), .B(new_n23396_), .ZN(new_n23397_));
  XOR2_X1    g23331(.A1(new_n23397_), .A2(new_n22540_), .Z(new_n23398_));
  NOR2_X1    g23332(.A1(new_n23398_), .A2(new_n23392_), .ZN(new_n23399_));
  INV_X1     g23333(.I(new_n23399_), .ZN(new_n23400_));
  NOR2_X1    g23334(.A1(new_n23386_), .A2(new_n23400_), .ZN(new_n23401_));
  NOR3_X1    g23335(.A1(new_n22666_), .A2(new_n22669_), .A3(new_n22663_), .ZN(new_n23402_));
  INV_X1     g23336(.I(new_n22670_), .ZN(new_n23403_));
  NOR2_X1    g23337(.A1(new_n23403_), .A2(new_n23402_), .ZN(new_n23404_));
  NOR2_X1    g23338(.A1(new_n23404_), .A2(new_n22664_), .ZN(new_n23405_));
  NOR2_X1    g23339(.A1(new_n23364_), .A2(new_n22678_), .ZN(new_n23406_));
  NOR2_X1    g23340(.A1(new_n23359_), .A2(new_n22679_), .ZN(new_n23407_));
  OAI21_X1   g23341(.A1(new_n23407_), .A2(new_n23406_), .B(new_n23382_), .ZN(new_n23408_));
  AOI21_X1   g23342(.A1(new_n22678_), .A2(new_n23364_), .B(new_n23404_), .ZN(new_n23409_));
  AOI21_X1   g23343(.A1(new_n23408_), .A2(new_n23409_), .B(new_n23405_), .ZN(new_n23410_));
  OAI21_X1   g23344(.A1(new_n23410_), .A2(new_n23391_), .B(new_n22658_), .ZN(new_n23411_));
  OAI21_X1   g23345(.A1(new_n23411_), .A2(new_n23401_), .B(new_n22659_), .ZN(new_n23412_));
  INV_X1     g23346(.I(new_n20939_), .ZN(new_n23413_));
  NAND2_X1   g23347(.A1(new_n19442_), .A2(new_n9488_), .ZN(new_n23414_));
  NAND2_X1   g23348(.A1(new_n19439_), .A2(new_n9503_), .ZN(new_n23415_));
  AOI21_X1   g23349(.A1(new_n19415_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n23416_));
  NAND4_X1   g23350(.A1(new_n23413_), .A2(new_n23414_), .A3(new_n23415_), .A4(new_n23416_), .ZN(new_n23417_));
  XOR2_X1    g23351(.A1(new_n23417_), .A2(\a[2] ), .Z(new_n23418_));
  INV_X1     g23352(.I(new_n23418_), .ZN(new_n23419_));
  NAND2_X1   g23353(.A1(new_n23412_), .A2(new_n23419_), .ZN(new_n23420_));
  NAND2_X1   g23354(.A1(new_n23410_), .A2(new_n23399_), .ZN(new_n23421_));
  NOR3_X1    g23355(.A1(new_n22656_), .A2(new_n22653_), .A3(new_n22236_), .ZN(new_n23422_));
  AOI21_X1   g23356(.A1(new_n22643_), .A2(new_n22649_), .B(new_n22237_), .ZN(new_n23423_));
  NOR2_X1    g23357(.A1(new_n23423_), .A2(new_n23422_), .ZN(new_n23424_));
  AOI21_X1   g23358(.A1(new_n23386_), .A2(new_n23392_), .B(new_n23424_), .ZN(new_n23425_));
  NAND2_X1   g23359(.A1(new_n23425_), .A2(new_n23421_), .ZN(new_n23426_));
  OAI21_X1   g23360(.A1(new_n22646_), .A2(new_n22647_), .B(new_n22655_), .ZN(new_n23427_));
  OAI22_X1   g23361(.A1(new_n17789_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n19400_), .ZN(new_n23428_));
  NAND2_X1   g23362(.A1(new_n19407_), .A2(new_n6838_), .ZN(new_n23429_));
  AOI21_X1   g23363(.A1(new_n23429_), .A2(new_n23428_), .B(new_n6836_), .ZN(new_n23430_));
  NAND2_X1   g23364(.A1(new_n20864_), .A2(new_n23430_), .ZN(new_n23431_));
  XOR2_X1    g23365(.A1(new_n23431_), .A2(\a[5] ), .Z(new_n23432_));
  INV_X1     g23366(.I(new_n23432_), .ZN(new_n23433_));
  NAND2_X1   g23367(.A1(new_n22603_), .A2(new_n22608_), .ZN(new_n23434_));
  NOR2_X1    g23368(.A1(new_n22603_), .A2(new_n22608_), .ZN(new_n23435_));
  OAI21_X1   g23369(.A1(new_n22600_), .A2(new_n23435_), .B(new_n23434_), .ZN(new_n23436_));
  NOR2_X1    g23370(.A1(new_n21485_), .A2(new_n21481_), .ZN(new_n23437_));
  NOR2_X1    g23371(.A1(new_n21441_), .A2(new_n21447_), .ZN(new_n23438_));
  XOR2_X1    g23372(.A1(new_n23437_), .A2(new_n23438_), .Z(new_n23439_));
  AOI22_X1   g23373(.A1(new_n17798_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n17802_), .ZN(new_n23440_));
  NOR2_X1    g23374(.A1(new_n19375_), .A2(new_n4710_), .ZN(new_n23441_));
  OAI21_X1   g23375(.A1(new_n23441_), .A2(new_n23440_), .B(new_n4706_), .ZN(new_n23442_));
  NOR2_X1    g23376(.A1(new_n21753_), .A2(new_n23442_), .ZN(new_n23443_));
  XOR2_X1    g23377(.A1(new_n23443_), .A2(\a[11] ), .Z(new_n23444_));
  OR2_X2     g23378(.A1(new_n23439_), .A2(new_n23444_), .Z(new_n23445_));
  NAND2_X1   g23379(.A1(new_n23439_), .A2(new_n23444_), .ZN(new_n23446_));
  NAND2_X1   g23380(.A1(new_n23445_), .A2(new_n23446_), .ZN(new_n23447_));
  NAND2_X1   g23381(.A1(new_n23436_), .A2(new_n23447_), .ZN(new_n23448_));
  XNOR2_X1   g23382(.A1(new_n23439_), .A2(new_n23444_), .ZN(new_n23449_));
  OR2_X2     g23383(.A1(new_n23436_), .A2(new_n23449_), .Z(new_n23450_));
  AOI22_X1   g23384(.A1(new_n19386_), .A2(new_n7530_), .B1(new_n6789_), .B2(new_n17794_), .ZN(new_n23451_));
  NOR2_X1    g23385(.A1(new_n19393_), .A2(new_n6785_), .ZN(new_n23452_));
  OAI21_X1   g23386(.A1(new_n23451_), .A2(new_n23452_), .B(new_n6775_), .ZN(new_n23453_));
  NOR2_X1    g23387(.A1(new_n20291_), .A2(new_n23453_), .ZN(new_n23454_));
  XOR2_X1    g23388(.A1(new_n23454_), .A2(new_n4009_), .Z(new_n23455_));
  NAND3_X1   g23389(.A1(new_n23450_), .A2(new_n23448_), .A3(new_n23455_), .ZN(new_n23456_));
  AOI21_X1   g23390(.A1(new_n23450_), .A2(new_n23448_), .B(new_n23455_), .ZN(new_n23457_));
  INV_X1     g23391(.I(new_n23457_), .ZN(new_n23458_));
  AOI21_X1   g23392(.A1(new_n23458_), .A2(new_n23456_), .B(new_n23433_), .ZN(new_n23459_));
  INV_X1     g23393(.I(new_n23456_), .ZN(new_n23460_));
  NOR3_X1    g23394(.A1(new_n23460_), .A2(new_n23432_), .A3(new_n23457_), .ZN(new_n23461_));
  NOR2_X1    g23395(.A1(new_n23459_), .A2(new_n23461_), .ZN(new_n23462_));
  XOR2_X1    g23396(.A1(new_n23462_), .A2(new_n23427_), .Z(new_n23463_));
  NOR2_X1    g23397(.A1(new_n23463_), .A2(new_n23419_), .ZN(new_n23464_));
  NAND3_X1   g23398(.A1(new_n23426_), .A2(new_n22659_), .A3(new_n23464_), .ZN(new_n23465_));
  NAND3_X1   g23399(.A1(new_n23420_), .A2(new_n23465_), .A3(new_n22232_), .ZN(new_n23466_));
  AOI21_X1   g23400(.A1(new_n23426_), .A2(new_n22659_), .B(new_n23418_), .ZN(new_n23467_));
  NOR3_X1    g23401(.A1(new_n23412_), .A2(new_n23463_), .A3(new_n23419_), .ZN(new_n23468_));
  OAI21_X1   g23402(.A1(new_n23468_), .A2(new_n23467_), .B(new_n22231_), .ZN(new_n23469_));
  NAND2_X1   g23403(.A1(new_n23436_), .A2(new_n23445_), .ZN(new_n23470_));
  NAND2_X1   g23404(.A1(new_n23470_), .A2(new_n23446_), .ZN(new_n23471_));
  INV_X1     g23405(.I(new_n23471_), .ZN(new_n23472_));
  NOR2_X1    g23406(.A1(new_n21422_), .A2(new_n21423_), .ZN(new_n23473_));
  XOR2_X1    g23407(.A1(new_n21486_), .A2(new_n21421_), .Z(new_n23474_));
  XOR2_X1    g23408(.A1(new_n23474_), .A2(new_n23473_), .Z(new_n23475_));
  OAI22_X1   g23409(.A1(new_n19375_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n17797_), .ZN(new_n23476_));
  NAND2_X1   g23410(.A1(new_n19386_), .A2(new_n4709_), .ZN(new_n23477_));
  AOI21_X1   g23411(.A1(new_n23477_), .A2(new_n23476_), .B(new_n4707_), .ZN(new_n23478_));
  NAND2_X1   g23412(.A1(new_n20162_), .A2(new_n23478_), .ZN(new_n23479_));
  XOR2_X1    g23413(.A1(new_n23479_), .A2(\a[11] ), .Z(new_n23480_));
  INV_X1     g23414(.I(new_n23480_), .ZN(new_n23481_));
  NAND2_X1   g23415(.A1(new_n23475_), .A2(new_n23481_), .ZN(new_n23482_));
  OR2_X2     g23416(.A1(new_n23475_), .A2(new_n23481_), .Z(new_n23483_));
  NAND2_X1   g23417(.A1(new_n23483_), .A2(new_n23482_), .ZN(new_n23484_));
  AOI22_X1   g23418(.A1(new_n19394_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n17794_), .ZN(new_n23485_));
  AOI21_X1   g23419(.A1(new_n6784_), .A2(new_n19399_), .B(new_n23485_), .ZN(new_n23486_));
  OR3_X2     g23420(.A1(new_n22541_), .A2(new_n6776_), .A3(new_n23486_), .Z(new_n23487_));
  XOR2_X1    g23421(.A1(new_n23487_), .A2(\a[8] ), .Z(new_n23488_));
  INV_X1     g23422(.I(new_n23488_), .ZN(new_n23489_));
  XOR2_X1    g23423(.A1(new_n23484_), .A2(new_n23489_), .Z(new_n23490_));
  NOR2_X1    g23424(.A1(new_n23472_), .A2(new_n23490_), .ZN(new_n23491_));
  XOR2_X1    g23425(.A1(new_n23484_), .A2(new_n23488_), .Z(new_n23492_));
  NOR2_X1    g23426(.A1(new_n23471_), .A2(new_n23492_), .ZN(new_n23493_));
  NOR2_X1    g23427(.A1(new_n23491_), .A2(new_n23493_), .ZN(new_n23494_));
  OAI22_X1   g23428(.A1(new_n19410_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n17789_), .ZN(new_n23495_));
  NAND2_X1   g23429(.A1(new_n19415_), .A2(new_n6838_), .ZN(new_n23496_));
  AOI21_X1   g23430(.A1(new_n23496_), .A2(new_n23495_), .B(new_n6836_), .ZN(new_n23497_));
  NAND2_X1   g23431(.A1(new_n20846_), .A2(new_n23497_), .ZN(new_n23498_));
  XOR2_X1    g23432(.A1(new_n23498_), .A2(\a[5] ), .Z(new_n23499_));
  XOR2_X1    g23433(.A1(new_n23494_), .A2(new_n23499_), .Z(new_n23500_));
  XOR2_X1    g23434(.A1(new_n23494_), .A2(new_n23499_), .Z(new_n23501_));
  NAND2_X1   g23435(.A1(new_n23501_), .A2(new_n23458_), .ZN(new_n23502_));
  OAI21_X1   g23436(.A1(new_n23500_), .A2(new_n23458_), .B(new_n23502_), .ZN(new_n23503_));
  NAND2_X1   g23437(.A1(new_n22654_), .A2(new_n22594_), .ZN(new_n23504_));
  NAND3_X1   g23438(.A1(new_n23462_), .A2(new_n22655_), .A3(new_n23504_), .ZN(new_n23505_));
  INV_X1     g23439(.I(new_n23505_), .ZN(new_n23506_));
  NOR2_X1    g23440(.A1(new_n23506_), .A2(new_n23459_), .ZN(new_n23507_));
  XNOR2_X1   g23441(.A1(new_n23503_), .A2(new_n23507_), .ZN(new_n23508_));
  INV_X1     g23442(.I(new_n23508_), .ZN(new_n23509_));
  AOI22_X1   g23443(.A1(new_n23469_), .A2(new_n23466_), .B1(new_n22232_), .B2(new_n23509_), .ZN(new_n23510_));
  NAND2_X1   g23444(.A1(new_n23510_), .A2(new_n22225_), .ZN(new_n23511_));
  AOI21_X1   g23445(.A1(new_n23420_), .A2(new_n23465_), .B(new_n22232_), .ZN(new_n23512_));
  AOI21_X1   g23446(.A1(new_n23469_), .A2(new_n23466_), .B(new_n23509_), .ZN(new_n23513_));
  NOR3_X1    g23447(.A1(new_n23513_), .A2(new_n22225_), .A3(new_n23512_), .ZN(new_n23514_));
  INV_X1     g23448(.I(new_n22225_), .ZN(new_n23515_));
  INV_X1     g23449(.I(new_n23512_), .ZN(new_n23516_));
  NOR3_X1    g23450(.A1(new_n23468_), .A2(new_n23467_), .A3(new_n22231_), .ZN(new_n23517_));
  AOI21_X1   g23451(.A1(new_n23420_), .A2(new_n23465_), .B(new_n22232_), .ZN(new_n23518_));
  OAI21_X1   g23452(.A1(new_n23517_), .A2(new_n23518_), .B(new_n23508_), .ZN(new_n23519_));
  AOI21_X1   g23453(.A1(new_n23519_), .A2(new_n23516_), .B(new_n23515_), .ZN(new_n23520_));
  XOR2_X1    g23454(.A1(new_n21453_), .A2(new_n21464_), .Z(new_n23521_));
  XOR2_X1    g23455(.A1(new_n23521_), .A2(new_n21462_), .Z(new_n23522_));
  INV_X1     g23456(.I(new_n23522_), .ZN(new_n23523_));
  NAND3_X1   g23457(.A1(new_n23472_), .A2(new_n23482_), .A3(new_n23483_), .ZN(new_n23524_));
  NAND2_X1   g23458(.A1(new_n23524_), .A2(new_n23483_), .ZN(new_n23525_));
  AOI22_X1   g23459(.A1(new_n19386_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n20127_), .ZN(new_n23526_));
  NOR2_X1    g23460(.A1(new_n17793_), .A2(new_n4710_), .ZN(new_n23527_));
  OAI21_X1   g23461(.A1(new_n23526_), .A2(new_n23527_), .B(new_n4706_), .ZN(new_n23528_));
  NOR2_X1    g23462(.A1(new_n21632_), .A2(new_n23528_), .ZN(new_n23529_));
  XOR2_X1    g23463(.A1(new_n23529_), .A2(new_n4034_), .Z(new_n23530_));
  NAND2_X1   g23464(.A1(new_n23525_), .A2(new_n23530_), .ZN(new_n23531_));
  NOR2_X1    g23465(.A1(new_n23525_), .A2(new_n23530_), .ZN(new_n23532_));
  INV_X1     g23466(.I(new_n23532_), .ZN(new_n23533_));
  NAND2_X1   g23467(.A1(new_n23533_), .A2(new_n23531_), .ZN(new_n23534_));
  XOR2_X1    g23468(.A1(new_n23534_), .A2(new_n23523_), .Z(new_n23535_));
  INV_X1     g23469(.I(new_n23494_), .ZN(new_n23536_));
  XNOR2_X1   g23470(.A1(new_n23471_), .A2(new_n23484_), .ZN(new_n23537_));
  OAI22_X1   g23471(.A1(new_n23536_), .A2(new_n23457_), .B1(new_n23489_), .B2(new_n23537_), .ZN(new_n23538_));
  OAI22_X1   g23472(.A1(new_n19400_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n19393_), .ZN(new_n23539_));
  NAND2_X1   g23473(.A1(new_n17790_), .A2(new_n6784_), .ZN(new_n23540_));
  AOI21_X1   g23474(.A1(new_n23540_), .A2(new_n23539_), .B(new_n6776_), .ZN(new_n23541_));
  NAND2_X1   g23475(.A1(new_n20251_), .A2(new_n23541_), .ZN(new_n23542_));
  XOR2_X1    g23476(.A1(new_n23542_), .A2(\a[8] ), .Z(new_n23543_));
  XOR2_X1    g23477(.A1(new_n23538_), .A2(new_n23543_), .Z(new_n23544_));
  XNOR2_X1   g23478(.A1(new_n23535_), .A2(new_n23544_), .ZN(new_n23545_));
  INV_X1     g23479(.I(new_n23499_), .ZN(new_n23546_));
  XOR2_X1    g23480(.A1(new_n23494_), .A2(new_n23457_), .Z(new_n23547_));
  OAI22_X1   g23481(.A1(new_n23506_), .A2(new_n23459_), .B1(new_n23546_), .B2(new_n23547_), .ZN(new_n23548_));
  NOR2_X1    g23482(.A1(new_n23503_), .A2(new_n23548_), .ZN(new_n23549_));
  OAI22_X1   g23483(.A1(new_n19410_), .A2(new_n6913_), .B1(new_n19412_), .B2(new_n6843_), .ZN(new_n23550_));
  NAND2_X1   g23484(.A1(new_n19439_), .A2(new_n6838_), .ZN(new_n23551_));
  AOI21_X1   g23485(.A1(new_n23551_), .A2(new_n23550_), .B(new_n6836_), .ZN(new_n23552_));
  NAND2_X1   g23486(.A1(new_n20827_), .A2(new_n23552_), .ZN(new_n23553_));
  XOR2_X1    g23487(.A1(new_n23553_), .A2(\a[5] ), .Z(new_n23554_));
  INV_X1     g23488(.I(new_n23554_), .ZN(new_n23555_));
  NOR2_X1    g23489(.A1(new_n23549_), .A2(new_n23555_), .ZN(new_n23556_));
  INV_X1     g23490(.I(new_n23556_), .ZN(new_n23557_));
  NAND2_X1   g23491(.A1(new_n23549_), .A2(new_n23555_), .ZN(new_n23558_));
  AOI21_X1   g23492(.A1(new_n23558_), .A2(new_n23557_), .B(new_n23545_), .ZN(new_n23559_));
  XOR2_X1    g23493(.A1(new_n23535_), .A2(new_n23544_), .Z(new_n23560_));
  INV_X1     g23494(.I(new_n23558_), .ZN(new_n23561_));
  NOR3_X1    g23495(.A1(new_n23560_), .A2(new_n23561_), .A3(new_n23556_), .ZN(new_n23562_));
  NOR2_X1    g23496(.A1(new_n23559_), .A2(new_n23562_), .ZN(new_n23563_));
  OAI21_X1   g23497(.A1(new_n23520_), .A2(new_n23514_), .B(new_n23563_), .ZN(new_n23564_));
  INV_X1     g23498(.I(new_n21100_), .ZN(new_n23565_));
  AOI22_X1   g23499(.A1(new_n19438_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n20896_), .ZN(new_n23566_));
  NOR2_X1    g23500(.A1(new_n19437_), .A2(new_n9489_), .ZN(new_n23567_));
  OAI21_X1   g23501(.A1(new_n23566_), .A2(new_n23567_), .B(new_n6922_), .ZN(new_n23568_));
  NOR3_X1    g23502(.A1(new_n23565_), .A2(\a[2] ), .A3(new_n23568_), .ZN(new_n23569_));
  NOR2_X1    g23503(.A1(new_n23565_), .A2(new_n23568_), .ZN(new_n23570_));
  NOR2_X1    g23504(.A1(new_n23570_), .A2(new_n4387_), .ZN(new_n23571_));
  NOR2_X1    g23505(.A1(new_n23571_), .A2(new_n23569_), .ZN(new_n23572_));
  AOI21_X1   g23506(.A1(new_n23564_), .A2(new_n23511_), .B(new_n23572_), .ZN(new_n23573_));
  NAND3_X1   g23507(.A1(new_n23519_), .A2(new_n23516_), .A3(new_n23515_), .ZN(new_n23574_));
  NAND2_X1   g23508(.A1(new_n23510_), .A2(new_n22225_), .ZN(new_n23575_));
  INV_X1     g23509(.I(new_n23563_), .ZN(new_n23576_));
  AOI22_X1   g23510(.A1(new_n23574_), .A2(new_n23575_), .B1(new_n23576_), .B2(new_n23515_), .ZN(new_n23577_));
  INV_X1     g23511(.I(new_n23572_), .ZN(new_n23578_));
  OR3_X2     g23512(.A1(new_n21605_), .A2(new_n21599_), .A3(new_n21603_), .Z(new_n23579_));
  AND2_X2    g23513(.A1(new_n23579_), .A2(new_n21606_), .Z(new_n23580_));
  NOR2_X1    g23514(.A1(new_n23578_), .A2(new_n23580_), .ZN(new_n23581_));
  INV_X1     g23515(.I(new_n23581_), .ZN(new_n23582_));
  NOR2_X1    g23516(.A1(new_n23577_), .A2(new_n23582_), .ZN(new_n23583_));
  OAI22_X1   g23517(.A1(new_n19437_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n17784_), .ZN(new_n23584_));
  NAND2_X1   g23518(.A1(new_n19472_), .A2(new_n9488_), .ZN(new_n23585_));
  AOI21_X1   g23519(.A1(new_n23585_), .A2(new_n23584_), .B(new_n9482_), .ZN(new_n23586_));
  NAND2_X1   g23520(.A1(new_n21117_), .A2(new_n23586_), .ZN(new_n23587_));
  XOR2_X1    g23521(.A1(new_n23587_), .A2(\a[2] ), .Z(new_n23588_));
  INV_X1     g23522(.I(new_n23588_), .ZN(new_n23589_));
  OAI21_X1   g23523(.A1(new_n23583_), .A2(new_n23573_), .B(new_n23589_), .ZN(new_n23590_));
  NAND2_X1   g23524(.A1(new_n23577_), .A2(new_n23578_), .ZN(new_n23591_));
  NAND3_X1   g23525(.A1(new_n23564_), .A2(new_n23511_), .A3(new_n23581_), .ZN(new_n23592_));
  XNOR2_X1   g23526(.A1(new_n22189_), .A2(new_n21611_), .ZN(new_n23593_));
  XNOR2_X1   g23527(.A1(new_n23593_), .A2(new_n21606_), .ZN(new_n23594_));
  NOR2_X1    g23528(.A1(new_n23594_), .A2(new_n23589_), .ZN(new_n23595_));
  NAND3_X1   g23529(.A1(new_n23591_), .A2(new_n23592_), .A3(new_n23595_), .ZN(new_n23596_));
  OAI22_X1   g23530(.A1(new_n19463_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n19437_), .ZN(new_n23597_));
  NAND2_X1   g23531(.A1(new_n17780_), .A2(new_n9488_), .ZN(new_n23598_));
  AOI21_X1   g23532(.A1(new_n23597_), .A2(new_n23598_), .B(new_n9482_), .ZN(new_n23599_));
  NAND2_X1   g23533(.A1(new_n21088_), .A2(new_n23599_), .ZN(new_n23600_));
  XOR2_X1    g23534(.A1(new_n23600_), .A2(\a[2] ), .Z(new_n23601_));
  AOI21_X1   g23535(.A1(new_n23590_), .A2(new_n23596_), .B(new_n23601_), .ZN(new_n23602_));
  AOI21_X1   g23536(.A1(new_n23591_), .A2(new_n23592_), .B(new_n23588_), .ZN(new_n23603_));
  INV_X1     g23537(.I(new_n23595_), .ZN(new_n23604_));
  NOR3_X1    g23538(.A1(new_n23583_), .A2(new_n23573_), .A3(new_n23604_), .ZN(new_n23605_));
  INV_X1     g23539(.I(new_n23601_), .ZN(new_n23606_));
  NAND2_X1   g23540(.A1(new_n22191_), .A2(new_n22192_), .ZN(new_n23607_));
  XOR2_X1    g23541(.A1(new_n21693_), .A2(new_n22195_), .Z(new_n23608_));
  XOR2_X1    g23542(.A1(new_n23608_), .A2(new_n23607_), .Z(new_n23609_));
  NOR2_X1    g23543(.A1(new_n23609_), .A2(new_n23606_), .ZN(new_n23610_));
  INV_X1     g23544(.I(new_n23610_), .ZN(new_n23611_));
  NOR3_X1    g23545(.A1(new_n23605_), .A2(new_n23603_), .A3(new_n23611_), .ZN(new_n23612_));
  NAND2_X1   g23546(.A1(new_n19484_), .A2(new_n9488_), .ZN(new_n23613_));
  NAND2_X1   g23547(.A1(new_n17780_), .A2(new_n9503_), .ZN(new_n23614_));
  AOI21_X1   g23548(.A1(new_n19472_), .A2(new_n6925_), .B(new_n6922_), .ZN(new_n23615_));
  NAND4_X1   g23549(.A1(new_n21180_), .A2(new_n23613_), .A3(new_n23614_), .A4(new_n23615_), .ZN(new_n23616_));
  XOR2_X1    g23550(.A1(new_n23616_), .A2(\a[2] ), .Z(new_n23617_));
  INV_X1     g23551(.I(new_n23617_), .ZN(new_n23618_));
  OAI21_X1   g23552(.A1(new_n23612_), .A2(new_n23602_), .B(new_n23618_), .ZN(new_n23619_));
  OAI21_X1   g23553(.A1(new_n23605_), .A2(new_n23603_), .B(new_n23606_), .ZN(new_n23620_));
  NAND3_X1   g23554(.A1(new_n23590_), .A2(new_n23596_), .A3(new_n23610_), .ZN(new_n23621_));
  XOR2_X1    g23555(.A1(new_n22201_), .A2(new_n21243_), .Z(new_n23622_));
  NOR2_X1    g23556(.A1(new_n23618_), .A2(new_n23622_), .ZN(new_n23623_));
  NAND3_X1   g23557(.A1(new_n23620_), .A2(new_n23621_), .A3(new_n23623_), .ZN(new_n23624_));
  NAND3_X1   g23558(.A1(new_n23619_), .A2(new_n23624_), .A3(new_n22220_), .ZN(new_n23625_));
  AOI21_X1   g23559(.A1(new_n23620_), .A2(new_n23621_), .B(new_n23617_), .ZN(new_n23626_));
  INV_X1     g23560(.I(new_n23623_), .ZN(new_n23627_));
  NOR3_X1    g23561(.A1(new_n23612_), .A2(new_n23602_), .A3(new_n23627_), .ZN(new_n23628_));
  OAI21_X1   g23562(.A1(new_n23628_), .A2(new_n23626_), .B(new_n22219_), .ZN(new_n23629_));
  XOR2_X1    g23563(.A1(new_n21696_), .A2(new_n21228_), .Z(new_n23630_));
  INV_X1     g23564(.I(new_n23630_), .ZN(new_n23631_));
  AOI22_X1   g23565(.A1(new_n23629_), .A2(new_n23625_), .B1(new_n22220_), .B2(new_n23631_), .ZN(new_n23632_));
  OAI22_X1   g23566(.A1(new_n19522_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n17775_), .ZN(new_n23633_));
  NAND2_X1   g23567(.A1(new_n17770_), .A2(new_n9488_), .ZN(new_n23634_));
  AOI21_X1   g23568(.A1(new_n23634_), .A2(new_n23633_), .B(new_n9482_), .ZN(new_n23635_));
  NAND2_X1   g23569(.A1(new_n19521_), .A2(new_n23635_), .ZN(new_n23636_));
  XOR2_X1    g23570(.A1(new_n23636_), .A2(\a[2] ), .Z(new_n23637_));
  INV_X1     g23571(.I(new_n23637_), .ZN(new_n23638_));
  NAND2_X1   g23572(.A1(new_n23632_), .A2(new_n23638_), .ZN(new_n23639_));
  OAI21_X1   g23573(.A1(new_n23628_), .A2(new_n23626_), .B(new_n22219_), .ZN(new_n23640_));
  NOR3_X1    g23574(.A1(new_n23628_), .A2(new_n23626_), .A3(new_n22219_), .ZN(new_n23641_));
  AOI21_X1   g23575(.A1(new_n23619_), .A2(new_n23624_), .B(new_n22220_), .ZN(new_n23642_));
  OAI21_X1   g23576(.A1(new_n23641_), .A2(new_n23642_), .B(new_n23630_), .ZN(new_n23643_));
  NOR2_X1    g23577(.A1(new_n21736_), .A2(new_n22210_), .ZN(new_n23644_));
  XOR2_X1    g23578(.A1(new_n23644_), .A2(new_n22203_), .Z(new_n23645_));
  NOR2_X1    g23579(.A1(new_n23645_), .A2(new_n23638_), .ZN(new_n23646_));
  NAND3_X1   g23580(.A1(new_n23643_), .A2(new_n23640_), .A3(new_n23646_), .ZN(new_n23647_));
  OAI22_X1   g23581(.A1(new_n19512_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n19522_), .ZN(new_n23648_));
  NAND2_X1   g23582(.A1(new_n21953_), .A2(new_n9488_), .ZN(new_n23649_));
  AOI21_X1   g23583(.A1(new_n23648_), .A2(new_n23649_), .B(new_n9482_), .ZN(new_n23650_));
  NAND2_X1   g23584(.A1(new_n21963_), .A2(new_n23650_), .ZN(new_n23651_));
  XOR2_X1    g23585(.A1(new_n23651_), .A2(\a[2] ), .Z(new_n23652_));
  AOI21_X1   g23586(.A1(new_n23647_), .A2(new_n23639_), .B(new_n23652_), .ZN(new_n23653_));
  AOI21_X1   g23587(.A1(new_n23643_), .A2(new_n23640_), .B(new_n23637_), .ZN(new_n23654_));
  INV_X1     g23588(.I(new_n23646_), .ZN(new_n23655_));
  NOR2_X1    g23589(.A1(new_n23632_), .A2(new_n23655_), .ZN(new_n23656_));
  INV_X1     g23590(.I(new_n23652_), .ZN(new_n23657_));
  XOR2_X1    g23591(.A1(new_n21738_), .A2(new_n22212_), .Z(new_n23658_));
  NOR2_X1    g23592(.A1(new_n23657_), .A2(new_n23658_), .ZN(new_n23659_));
  INV_X1     g23593(.I(new_n23659_), .ZN(new_n23660_));
  NOR3_X1    g23594(.A1(new_n23654_), .A2(new_n23656_), .A3(new_n23660_), .ZN(new_n23661_));
  NOR4_X1    g23595(.A1(new_n23653_), .A2(new_n23661_), .A3(new_n22181_), .A4(new_n22214_), .ZN(new_n23662_));
  NOR2_X1    g23596(.A1(new_n22181_), .A2(new_n22214_), .ZN(new_n23663_));
  NOR2_X1    g23597(.A1(new_n21146_), .A2(new_n21145_), .ZN(new_n23664_));
  XOR2_X1    g23598(.A1(new_n21746_), .A2(new_n19527_), .Z(new_n23665_));
  XOR2_X1    g23599(.A1(new_n23665_), .A2(new_n23664_), .Z(new_n23666_));
  INV_X1     g23600(.I(new_n23666_), .ZN(new_n23667_));
  AOI21_X1   g23601(.A1(new_n21889_), .A2(new_n22052_), .B(new_n22054_), .ZN(new_n23668_));
  NAND2_X1   g23602(.A1(new_n23668_), .A2(new_n22051_), .ZN(new_n23669_));
  NAND2_X1   g23603(.A1(new_n22053_), .A2(new_n22055_), .ZN(new_n23670_));
  NAND2_X1   g23604(.A1(new_n23670_), .A2(new_n22048_), .ZN(new_n23671_));
  AOI21_X1   g23605(.A1(new_n23671_), .A2(new_n23669_), .B(new_n22115_), .ZN(new_n23672_));
  AOI21_X1   g23606(.A1(new_n22157_), .A2(new_n22116_), .B(new_n22118_), .ZN(new_n23673_));
  NOR2_X1    g23607(.A1(new_n23672_), .A2(new_n23673_), .ZN(new_n23674_));
  INV_X1     g23608(.I(new_n23674_), .ZN(new_n23675_));
  AOI22_X1   g23609(.A1(new_n22048_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n21953_), .ZN(new_n23676_));
  NOR2_X1    g23610(.A1(new_n22115_), .A2(new_n9489_), .ZN(new_n23677_));
  OAI21_X1   g23611(.A1(new_n23677_), .A2(new_n23676_), .B(new_n6922_), .ZN(new_n23678_));
  NOR2_X1    g23612(.A1(new_n23675_), .A2(new_n23678_), .ZN(new_n23679_));
  XOR2_X1    g23613(.A1(new_n23679_), .A2(new_n4387_), .Z(new_n23680_));
  NAND2_X1   g23614(.A1(new_n23667_), .A2(new_n23680_), .ZN(new_n23681_));
  INV_X1     g23615(.I(new_n23681_), .ZN(new_n23682_));
  NOR2_X1    g23616(.A1(new_n23667_), .A2(new_n23680_), .ZN(new_n23683_));
  NOR3_X1    g23617(.A1(new_n23682_), .A2(new_n23663_), .A3(new_n23683_), .ZN(new_n23684_));
  INV_X1     g23618(.I(new_n23684_), .ZN(new_n23685_));
  OAI21_X1   g23619(.A1(new_n23662_), .A2(new_n23685_), .B(new_n22168_), .ZN(new_n23686_));
  INV_X1     g23620(.I(new_n22168_), .ZN(new_n23687_));
  OAI21_X1   g23621(.A1(new_n23654_), .A2(new_n23656_), .B(new_n23657_), .ZN(new_n23688_));
  NAND3_X1   g23622(.A1(new_n23647_), .A2(new_n23639_), .A3(new_n23659_), .ZN(new_n23689_));
  NAND3_X1   g23623(.A1(new_n23688_), .A2(new_n23689_), .A3(new_n23663_), .ZN(new_n23690_));
  NAND3_X1   g23624(.A1(new_n23690_), .A2(new_n23687_), .A3(new_n23684_), .ZN(new_n23691_));
  AOI21_X1   g23625(.A1(new_n23686_), .A2(new_n23691_), .B(new_n21990_), .ZN(new_n23692_));
  AOI21_X1   g23626(.A1(new_n23690_), .A2(new_n23684_), .B(new_n23687_), .ZN(new_n23693_));
  NOR3_X1    g23627(.A1(new_n23662_), .A2(new_n22168_), .A3(new_n23685_), .ZN(new_n23694_));
  NOR3_X1    g23628(.A1(new_n23694_), .A2(new_n23693_), .A3(new_n21989_), .ZN(new_n23695_));
  NOR2_X1    g23629(.A1(new_n23695_), .A2(new_n23692_), .ZN(new_n23696_));
  NOR2_X1    g23630(.A1(new_n23682_), .A2(new_n23683_), .ZN(new_n23697_));
  NAND3_X1   g23631(.A1(new_n23688_), .A2(new_n23689_), .A3(new_n22181_), .ZN(new_n23698_));
  OAI21_X1   g23632(.A1(new_n23653_), .A2(new_n23661_), .B(new_n22180_), .ZN(new_n23699_));
  NAND2_X1   g23633(.A1(new_n23699_), .A2(new_n23698_), .ZN(new_n23700_));
  NAND3_X1   g23634(.A1(new_n23700_), .A2(new_n22214_), .A3(new_n23697_), .ZN(new_n23701_));
  INV_X1     g23635(.I(new_n23697_), .ZN(new_n23702_));
  NOR3_X1    g23636(.A1(new_n23653_), .A2(new_n23661_), .A3(new_n22180_), .ZN(new_n23703_));
  AOI21_X1   g23637(.A1(new_n23688_), .A2(new_n23689_), .B(new_n22181_), .ZN(new_n23704_));
  OAI21_X1   g23638(.A1(new_n23703_), .A2(new_n23704_), .B(new_n22214_), .ZN(new_n23705_));
  NAND2_X1   g23639(.A1(new_n23705_), .A2(new_n23702_), .ZN(new_n23706_));
  AOI21_X1   g23640(.A1(new_n23688_), .A2(new_n23689_), .B(new_n22180_), .ZN(new_n23707_));
  NAND3_X1   g23641(.A1(new_n23706_), .A2(new_n23701_), .A3(new_n23707_), .ZN(new_n23708_));
  NOR2_X1    g23642(.A1(new_n23705_), .A2(new_n23702_), .ZN(new_n23709_));
  AOI21_X1   g23643(.A1(new_n23700_), .A2(new_n22214_), .B(new_n23697_), .ZN(new_n23710_));
  INV_X1     g23644(.I(new_n23707_), .ZN(new_n23711_));
  OAI21_X1   g23645(.A1(new_n23709_), .A2(new_n23710_), .B(new_n23711_), .ZN(new_n23712_));
  NAND2_X1   g23646(.A1(new_n23712_), .A2(new_n23708_), .ZN(new_n23713_));
  XOR2_X1    g23647(.A1(new_n23713_), .A2(new_n23696_), .Z(\result[0] ));
  NOR2_X1    g23648(.A1(new_n21837_), .A2(new_n21842_), .ZN(new_n23715_));
  INV_X1     g23649(.I(new_n21818_), .ZN(new_n23716_));
  NAND3_X1   g23650(.A1(new_n21813_), .A2(new_n21806_), .A3(new_n23716_), .ZN(new_n23717_));
  INV_X1     g23651(.I(new_n21812_), .ZN(new_n23718_));
  NAND2_X1   g23652(.A1(new_n21811_), .A2(new_n21810_), .ZN(new_n23719_));
  OAI21_X1   g23653(.A1(new_n21807_), .A2(new_n20123_), .B(new_n23719_), .ZN(new_n23720_));
  OAI22_X1   g23654(.A1(new_n19375_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n17797_), .ZN(new_n23721_));
  NAND2_X1   g23655(.A1(new_n19386_), .A2(new_n3312_), .ZN(new_n23722_));
  AOI21_X1   g23656(.A1(new_n23722_), .A2(new_n23721_), .B(new_n3302_), .ZN(new_n23723_));
  OAI21_X1   g23657(.A1(new_n20161_), .A2(new_n20159_), .B(new_n23723_), .ZN(new_n23724_));
  XOR2_X1    g23658(.A1(new_n23724_), .A2(\a[23] ), .Z(new_n23725_));
  NAND2_X1   g23659(.A1(new_n20091_), .A2(new_n20088_), .ZN(new_n23726_));
  NAND2_X1   g23660(.A1(new_n21770_), .A2(new_n21787_), .ZN(new_n23727_));
  OAI21_X1   g23661(.A1(new_n21770_), .A2(new_n21788_), .B(new_n23727_), .ZN(new_n23728_));
  NOR2_X1    g23662(.A1(new_n21768_), .A2(new_n23728_), .ZN(new_n23729_));
  AOI21_X1   g23663(.A1(new_n20092_), .A2(new_n23726_), .B(new_n23729_), .ZN(new_n23730_));
  OAI21_X1   g23664(.A1(new_n19966_), .A2(new_n19979_), .B(new_n19988_), .ZN(new_n23731_));
  AOI21_X1   g23665(.A1(new_n23731_), .A2(new_n20079_), .B(new_n20081_), .ZN(new_n23732_));
  INV_X1     g23666(.I(new_n21784_), .ZN(new_n23733_));
  OAI21_X1   g23667(.A1(new_n23732_), .A2(new_n23733_), .B(new_n21786_), .ZN(new_n23734_));
  AOI21_X1   g23668(.A1(new_n19321_), .A2(new_n3189_), .B(new_n2763_), .ZN(new_n23735_));
  OAI21_X1   g23669(.A1(new_n19304_), .A2(new_n2771_), .B(new_n23735_), .ZN(new_n23736_));
  AOI21_X1   g23670(.A1(new_n17827_), .A2(new_n3332_), .B(new_n23736_), .ZN(new_n23737_));
  NAND2_X1   g23671(.A1(new_n22297_), .A2(new_n23737_), .ZN(new_n23738_));
  INV_X1     g23672(.I(new_n1594_), .ZN(new_n23739_));
  NAND3_X1   g23673(.A1(new_n2339_), .A2(new_n1767_), .A3(new_n1416_), .ZN(new_n23740_));
  NAND4_X1   g23674(.A1(new_n1816_), .A2(new_n842_), .A3(new_n409_), .A4(new_n508_), .ZN(new_n23741_));
  NOR4_X1    g23675(.A1(new_n23740_), .A2(new_n3203_), .A3(new_n1328_), .A4(new_n23741_), .ZN(new_n23742_));
  INV_X1     g23676(.I(new_n1569_), .ZN(new_n23743_));
  NOR4_X1    g23677(.A1(new_n202_), .A2(new_n172_), .A3(new_n731_), .A4(new_n594_), .ZN(new_n23744_));
  NOR3_X1    g23678(.A1(new_n2524_), .A2(new_n23743_), .A3(new_n23744_), .ZN(new_n23745_));
  NAND4_X1   g23679(.A1(new_n23742_), .A2(new_n4885_), .A3(new_n23745_), .A4(new_n4784_), .ZN(new_n23746_));
  NOR4_X1    g23680(.A1(new_n11933_), .A2(new_n728_), .A3(new_n23739_), .A4(new_n23746_), .ZN(new_n23747_));
  INV_X1     g23681(.I(new_n23747_), .ZN(new_n23748_));
  NAND2_X1   g23682(.A1(new_n23738_), .A2(new_n23748_), .ZN(new_n23749_));
  NOR2_X1    g23683(.A1(new_n23738_), .A2(new_n23748_), .ZN(new_n23750_));
  INV_X1     g23684(.I(new_n23750_), .ZN(new_n23751_));
  NAND2_X1   g23685(.A1(new_n23751_), .A2(new_n23749_), .ZN(new_n23752_));
  NAND3_X1   g23686(.A1(new_n22297_), .A2(new_n23737_), .A3(new_n23748_), .ZN(new_n23753_));
  NAND2_X1   g23687(.A1(new_n23738_), .A2(new_n23747_), .ZN(new_n23754_));
  AOI21_X1   g23688(.A1(new_n23753_), .A2(new_n23754_), .B(new_n23734_), .ZN(new_n23755_));
  AOI21_X1   g23689(.A1(new_n23734_), .A2(new_n23752_), .B(new_n23755_), .ZN(new_n23756_));
  AOI22_X1   g23690(.A1(new_n19349_), .A2(new_n2746_), .B1(new_n3275_), .B2(new_n19350_), .ZN(new_n23757_));
  NOR2_X1    g23691(.A1(new_n17806_), .A2(new_n3175_), .ZN(new_n23758_));
  OAI21_X1   g23692(.A1(new_n23757_), .A2(new_n23758_), .B(new_n2736_), .ZN(new_n23759_));
  INV_X1     g23693(.I(new_n23759_), .ZN(new_n23760_));
  NAND3_X1   g23694(.A1(new_n19922_), .A2(new_n74_), .A3(new_n23760_), .ZN(new_n23761_));
  INV_X1     g23695(.I(new_n23761_), .ZN(new_n23762_));
  AOI21_X1   g23696(.A1(new_n19922_), .A2(new_n23760_), .B(new_n74_), .ZN(new_n23763_));
  NOR3_X1    g23697(.A1(new_n23762_), .A2(new_n23756_), .A3(new_n23763_), .ZN(new_n23764_));
  INV_X1     g23698(.I(new_n23749_), .ZN(new_n23765_));
  OAI21_X1   g23699(.A1(new_n23765_), .A2(new_n23750_), .B(new_n23734_), .ZN(new_n23766_));
  INV_X1     g23700(.I(new_n23734_), .ZN(new_n23767_));
  NAND2_X1   g23701(.A1(new_n23754_), .A2(new_n23753_), .ZN(new_n23768_));
  NAND2_X1   g23702(.A1(new_n23767_), .A2(new_n23768_), .ZN(new_n23769_));
  NAND2_X1   g23703(.A1(new_n23769_), .A2(new_n23766_), .ZN(new_n23770_));
  INV_X1     g23704(.I(new_n23763_), .ZN(new_n23771_));
  AOI21_X1   g23705(.A1(new_n23771_), .A2(new_n23761_), .B(new_n23770_), .ZN(new_n23772_));
  OAI22_X1   g23706(.A1(new_n23730_), .A2(new_n21794_), .B1(new_n23772_), .B2(new_n23764_), .ZN(new_n23773_));
  AOI21_X1   g23707(.A1(new_n21760_), .A2(new_n21793_), .B(new_n21794_), .ZN(new_n23774_));
  NOR3_X1    g23708(.A1(new_n23762_), .A2(new_n23770_), .A3(new_n23763_), .ZN(new_n23775_));
  OAI21_X1   g23709(.A1(new_n23762_), .A2(new_n23763_), .B(new_n23770_), .ZN(new_n23776_));
  INV_X1     g23710(.I(new_n23776_), .ZN(new_n23777_));
  OAI21_X1   g23711(.A1(new_n23777_), .A2(new_n23775_), .B(new_n23774_), .ZN(new_n23778_));
  OAI22_X1   g23712(.A1(new_n19356_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n19364_), .ZN(new_n23779_));
  NAND2_X1   g23713(.A1(new_n17802_), .A2(new_n3317_), .ZN(new_n23780_));
  AOI21_X1   g23714(.A1(new_n23779_), .A2(new_n23780_), .B(new_n3260_), .ZN(new_n23781_));
  NAND2_X1   g23715(.A1(new_n19951_), .A2(new_n23781_), .ZN(new_n23782_));
  XOR2_X1    g23716(.A1(new_n23782_), .A2(new_n72_), .Z(new_n23783_));
  NAND3_X1   g23717(.A1(new_n23783_), .A2(new_n23773_), .A3(new_n23778_), .ZN(new_n23784_));
  NAND2_X1   g23718(.A1(new_n23778_), .A2(new_n23773_), .ZN(new_n23785_));
  XOR2_X1    g23719(.A1(new_n23782_), .A2(\a[26] ), .Z(new_n23786_));
  NAND2_X1   g23720(.A1(new_n23785_), .A2(new_n23786_), .ZN(new_n23787_));
  NAND4_X1   g23721(.A1(new_n23787_), .A2(new_n21797_), .A3(new_n23784_), .A4(new_n21803_), .ZN(new_n23788_));
  NAND2_X1   g23722(.A1(new_n21797_), .A2(new_n21803_), .ZN(new_n23789_));
  NOR2_X1    g23723(.A1(new_n23785_), .A2(new_n23786_), .ZN(new_n23790_));
  AOI21_X1   g23724(.A1(new_n23773_), .A2(new_n23778_), .B(new_n23783_), .ZN(new_n23791_));
  OAI21_X1   g23725(.A1(new_n23790_), .A2(new_n23791_), .B(new_n23789_), .ZN(new_n23792_));
  NAND3_X1   g23726(.A1(new_n23788_), .A2(new_n23792_), .A3(new_n23725_), .ZN(new_n23793_));
  INV_X1     g23727(.I(new_n23725_), .ZN(new_n23794_));
  NOR3_X1    g23728(.A1(new_n23790_), .A2(new_n23791_), .A3(new_n23789_), .ZN(new_n23795_));
  AOI22_X1   g23729(.A1(new_n23787_), .A2(new_n23784_), .B1(new_n21797_), .B2(new_n21803_), .ZN(new_n23796_));
  OAI21_X1   g23730(.A1(new_n23796_), .A2(new_n23795_), .B(new_n23794_), .ZN(new_n23797_));
  NAND2_X1   g23731(.A1(new_n23797_), .A2(new_n23793_), .ZN(new_n23798_));
  NAND3_X1   g23732(.A1(new_n23720_), .A2(new_n23798_), .A3(new_n23718_), .ZN(new_n23799_));
  AOI21_X1   g23733(.A1(new_n21751_), .A2(new_n21748_), .B(new_n21809_), .ZN(new_n23800_));
  NOR3_X1    g23734(.A1(new_n23796_), .A2(new_n23795_), .A3(new_n23794_), .ZN(new_n23801_));
  AOI21_X1   g23735(.A1(new_n23788_), .A2(new_n23792_), .B(new_n23725_), .ZN(new_n23802_));
  NOR2_X1    g23736(.A1(new_n23801_), .A2(new_n23802_), .ZN(new_n23803_));
  OAI21_X1   g23737(.A1(new_n23800_), .A2(new_n21812_), .B(new_n23803_), .ZN(new_n23804_));
  OAI22_X1   g23738(.A1(new_n19393_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n17793_), .ZN(new_n23805_));
  NAND2_X1   g23739(.A1(new_n19399_), .A2(new_n4096_), .ZN(new_n23806_));
  AOI21_X1   g23740(.A1(new_n23806_), .A2(new_n23805_), .B(new_n4095_), .ZN(new_n23807_));
  NAND2_X1   g23741(.A1(new_n20264_), .A2(new_n23807_), .ZN(new_n23808_));
  XOR2_X1    g23742(.A1(new_n23808_), .A2(\a[20] ), .Z(new_n23809_));
  INV_X1     g23743(.I(new_n23809_), .ZN(new_n23810_));
  NAND3_X1   g23744(.A1(new_n23804_), .A2(new_n23799_), .A3(new_n23810_), .ZN(new_n23811_));
  NOR3_X1    g23745(.A1(new_n23800_), .A2(new_n21812_), .A3(new_n23803_), .ZN(new_n23812_));
  AOI21_X1   g23746(.A1(new_n23720_), .A2(new_n23718_), .B(new_n23798_), .ZN(new_n23813_));
  OAI21_X1   g23747(.A1(new_n23812_), .A2(new_n23813_), .B(new_n23809_), .ZN(new_n23814_));
  NAND3_X1   g23748(.A1(new_n23814_), .A2(new_n23811_), .A3(new_n23717_), .ZN(new_n23815_));
  XOR2_X1    g23749(.A1(new_n21804_), .A2(new_n21810_), .Z(new_n23816_));
  NOR2_X1    g23750(.A1(new_n21808_), .A2(new_n23816_), .ZN(new_n23817_));
  AOI21_X1   g23751(.A1(new_n23719_), .A2(new_n23718_), .B(new_n21752_), .ZN(new_n23818_));
  NOR3_X1    g23752(.A1(new_n23818_), .A2(new_n23817_), .A3(new_n21818_), .ZN(new_n23819_));
  NOR3_X1    g23753(.A1(new_n23812_), .A2(new_n23813_), .A3(new_n23809_), .ZN(new_n23820_));
  AOI21_X1   g23754(.A1(new_n23804_), .A2(new_n23799_), .B(new_n23810_), .ZN(new_n23821_));
  OAI21_X1   g23755(.A1(new_n23820_), .A2(new_n23821_), .B(new_n23819_), .ZN(new_n23822_));
  OAI22_X1   g23756(.A1(new_n19410_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n17789_), .ZN(new_n23823_));
  NAND2_X1   g23757(.A1(new_n19415_), .A2(new_n4469_), .ZN(new_n23824_));
  AOI21_X1   g23758(.A1(new_n23824_), .A2(new_n23823_), .B(new_n4468_), .ZN(new_n23825_));
  NAND2_X1   g23759(.A1(new_n20846_), .A2(new_n23825_), .ZN(new_n23826_));
  XOR2_X1    g23760(.A1(new_n23826_), .A2(new_n3372_), .Z(new_n23827_));
  INV_X1     g23761(.I(new_n23827_), .ZN(new_n23828_));
  NAND3_X1   g23762(.A1(new_n23828_), .A2(new_n23822_), .A3(new_n23815_), .ZN(new_n23829_));
  NOR3_X1    g23763(.A1(new_n23819_), .A2(new_n23820_), .A3(new_n23821_), .ZN(new_n23830_));
  AOI21_X1   g23764(.A1(new_n23814_), .A2(new_n23811_), .B(new_n23717_), .ZN(new_n23831_));
  OAI21_X1   g23765(.A1(new_n23830_), .A2(new_n23831_), .B(new_n23827_), .ZN(new_n23832_));
  NAND2_X1   g23766(.A1(new_n23829_), .A2(new_n23832_), .ZN(new_n23833_));
  OAI21_X1   g23767(.A1(new_n21836_), .A2(new_n21831_), .B(new_n21827_), .ZN(new_n23834_));
  NOR2_X1    g23768(.A1(new_n23834_), .A2(new_n23833_), .ZN(new_n23835_));
  NOR3_X1    g23769(.A1(new_n23830_), .A2(new_n23831_), .A3(new_n23827_), .ZN(new_n23836_));
  AOI21_X1   g23770(.A1(new_n23822_), .A2(new_n23815_), .B(new_n23828_), .ZN(new_n23837_));
  NOR2_X1    g23771(.A1(new_n23837_), .A2(new_n23836_), .ZN(new_n23838_));
  AOI21_X1   g23772(.A1(new_n21847_), .A2(new_n21851_), .B(new_n21849_), .ZN(new_n23839_));
  NOR2_X1    g23773(.A1(new_n23839_), .A2(new_n23838_), .ZN(new_n23840_));
  OAI22_X1   g23774(.A1(new_n19423_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n17787_), .ZN(new_n23841_));
  NAND2_X1   g23775(.A1(new_n20896_), .A2(new_n6090_), .ZN(new_n23842_));
  AOI21_X1   g23776(.A1(new_n23842_), .A2(new_n23841_), .B(new_n6082_), .ZN(new_n23843_));
  NAND2_X1   g23777(.A1(new_n22226_), .A2(new_n23843_), .ZN(new_n23844_));
  XOR2_X1    g23778(.A1(new_n23844_), .A2(\a[14] ), .Z(new_n23845_));
  NOR3_X1    g23779(.A1(new_n23840_), .A2(new_n23835_), .A3(new_n23845_), .ZN(new_n23846_));
  NAND2_X1   g23780(.A1(new_n21847_), .A2(new_n21851_), .ZN(new_n23847_));
  NAND3_X1   g23781(.A1(new_n23847_), .A2(new_n21827_), .A3(new_n23838_), .ZN(new_n23848_));
  NAND2_X1   g23782(.A1(new_n23834_), .A2(new_n23833_), .ZN(new_n23849_));
  XOR2_X1    g23783(.A1(new_n23844_), .A2(new_n3521_), .Z(new_n23850_));
  AOI21_X1   g23784(.A1(new_n23848_), .A2(new_n23849_), .B(new_n23850_), .ZN(new_n23851_));
  NOR3_X1    g23785(.A1(new_n23846_), .A2(new_n23851_), .A3(new_n23715_), .ZN(new_n23852_));
  NAND2_X1   g23786(.A1(new_n21853_), .A2(new_n21843_), .ZN(new_n23853_));
  NAND3_X1   g23787(.A1(new_n23848_), .A2(new_n23849_), .A3(new_n23850_), .ZN(new_n23854_));
  OAI21_X1   g23788(.A1(new_n23840_), .A2(new_n23835_), .B(new_n23845_), .ZN(new_n23855_));
  AOI21_X1   g23789(.A1(new_n23855_), .A2(new_n23854_), .B(new_n23853_), .ZN(new_n23856_));
  OAI22_X1   g23790(.A1(new_n19437_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n17784_), .ZN(new_n23857_));
  NAND2_X1   g23791(.A1(new_n19472_), .A2(new_n4709_), .ZN(new_n23858_));
  AOI21_X1   g23792(.A1(new_n23858_), .A2(new_n23857_), .B(new_n4707_), .ZN(new_n23859_));
  NAND2_X1   g23793(.A1(new_n21117_), .A2(new_n23859_), .ZN(new_n23860_));
  XOR2_X1    g23794(.A1(new_n23860_), .A2(new_n4034_), .Z(new_n23861_));
  NOR3_X1    g23795(.A1(new_n23852_), .A2(new_n23856_), .A3(new_n23861_), .ZN(new_n23862_));
  NAND3_X1   g23796(.A1(new_n23855_), .A2(new_n23854_), .A3(new_n23853_), .ZN(new_n23863_));
  OAI21_X1   g23797(.A1(new_n23846_), .A2(new_n23851_), .B(new_n23715_), .ZN(new_n23864_));
  XOR2_X1    g23798(.A1(new_n23860_), .A2(\a[11] ), .Z(new_n23865_));
  AOI21_X1   g23799(.A1(new_n23864_), .A2(new_n23863_), .B(new_n23865_), .ZN(new_n23866_));
  NOR2_X1    g23800(.A1(new_n23862_), .A2(new_n23866_), .ZN(new_n23867_));
  AOI21_X1   g23801(.A1(new_n21876_), .A2(new_n21864_), .B(new_n21859_), .ZN(new_n23868_));
  NAND2_X1   g23802(.A1(new_n23868_), .A2(new_n23867_), .ZN(new_n23869_));
  NAND3_X1   g23803(.A1(new_n23864_), .A2(new_n23863_), .A3(new_n23865_), .ZN(new_n23870_));
  OAI21_X1   g23804(.A1(new_n23852_), .A2(new_n23856_), .B(new_n23861_), .ZN(new_n23871_));
  NAND2_X1   g23805(.A1(new_n23871_), .A2(new_n23870_), .ZN(new_n23872_));
  OAI21_X1   g23806(.A1(new_n21869_), .A2(new_n21873_), .B(new_n21871_), .ZN(new_n23873_));
  NAND2_X1   g23807(.A1(new_n23873_), .A2(new_n23872_), .ZN(new_n23874_));
  OAI22_X1   g23808(.A1(new_n17775_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n19475_), .ZN(new_n23875_));
  NAND2_X1   g23809(.A1(new_n21157_), .A2(new_n6784_), .ZN(new_n23876_));
  AOI21_X1   g23810(.A1(new_n23876_), .A2(new_n23875_), .B(new_n6776_), .ZN(new_n23877_));
  NAND3_X1   g23811(.A1(new_n21155_), .A2(new_n4009_), .A3(new_n23877_), .ZN(new_n23878_));
  AOI21_X1   g23812(.A1(new_n21155_), .A2(new_n23877_), .B(new_n4009_), .ZN(new_n23879_));
  INV_X1     g23813(.I(new_n23879_), .ZN(new_n23880_));
  NAND2_X1   g23814(.A1(new_n23880_), .A2(new_n23878_), .ZN(new_n23881_));
  NAND3_X1   g23815(.A1(new_n23869_), .A2(new_n23874_), .A3(new_n23881_), .ZN(new_n23882_));
  NOR2_X1    g23816(.A1(new_n23873_), .A2(new_n23872_), .ZN(new_n23883_));
  NOR2_X1    g23817(.A1(new_n23868_), .A2(new_n23867_), .ZN(new_n23884_));
  INV_X1     g23818(.I(new_n23878_), .ZN(new_n23885_));
  NOR2_X1    g23819(.A1(new_n23885_), .A2(new_n23879_), .ZN(new_n23886_));
  OAI21_X1   g23820(.A1(new_n23884_), .A2(new_n23883_), .B(new_n23886_), .ZN(new_n23887_));
  NOR2_X1    g23821(.A1(new_n21878_), .A2(new_n21883_), .ZN(new_n23888_));
  NAND3_X1   g23822(.A1(new_n23887_), .A2(new_n23882_), .A3(new_n23888_), .ZN(new_n23889_));
  NOR3_X1    g23823(.A1(new_n23884_), .A2(new_n23883_), .A3(new_n23886_), .ZN(new_n23890_));
  AOI21_X1   g23824(.A1(new_n23869_), .A2(new_n23874_), .B(new_n23881_), .ZN(new_n23891_));
  NAND2_X1   g23825(.A1(new_n21981_), .A2(new_n21982_), .ZN(new_n23892_));
  OAI21_X1   g23826(.A1(new_n23891_), .A2(new_n23890_), .B(new_n23892_), .ZN(new_n23893_));
  OAI22_X1   g23827(.A1(new_n19512_), .A2(new_n6913_), .B1(new_n21960_), .B2(new_n6843_), .ZN(new_n23894_));
  NAND2_X1   g23828(.A1(new_n22048_), .A2(new_n6838_), .ZN(new_n23895_));
  AOI21_X1   g23829(.A1(new_n23895_), .A2(new_n23894_), .B(new_n6836_), .ZN(new_n23896_));
  INV_X1     g23830(.I(new_n23896_), .ZN(new_n23897_));
  NOR4_X1    g23831(.A1(new_n22174_), .A2(new_n22171_), .A3(\a[5] ), .A4(new_n23897_), .ZN(new_n23898_));
  INV_X1     g23832(.I(new_n23898_), .ZN(new_n23899_));
  NAND3_X1   g23833(.A1(new_n22173_), .A2(new_n22051_), .A3(new_n22172_), .ZN(new_n23900_));
  OAI21_X1   g23834(.A1(new_n21970_), .A2(new_n21960_), .B(new_n21973_), .ZN(new_n23901_));
  OAI21_X1   g23835(.A1(new_n23901_), .A2(new_n22169_), .B(new_n22048_), .ZN(new_n23902_));
  NAND3_X1   g23836(.A1(new_n23902_), .A2(new_n23900_), .A3(new_n23896_), .ZN(new_n23903_));
  NAND2_X1   g23837(.A1(new_n23903_), .A2(\a[5] ), .ZN(new_n23904_));
  NAND4_X1   g23838(.A1(new_n23893_), .A2(new_n23889_), .A3(new_n23899_), .A4(new_n23904_), .ZN(new_n23905_));
  NOR3_X1    g23839(.A1(new_n23891_), .A2(new_n23890_), .A3(new_n23892_), .ZN(new_n23906_));
  AOI21_X1   g23840(.A1(new_n23887_), .A2(new_n23882_), .B(new_n23888_), .ZN(new_n23907_));
  NAND2_X1   g23841(.A1(new_n23904_), .A2(new_n23899_), .ZN(new_n23908_));
  OAI21_X1   g23842(.A1(new_n23906_), .A2(new_n23907_), .B(new_n23908_), .ZN(new_n23909_));
  NAND2_X1   g23843(.A1(new_n23909_), .A2(new_n23905_), .ZN(new_n23910_));
  NOR3_X1    g23844(.A1(new_n21146_), .A2(new_n21145_), .A3(new_n21144_), .ZN(new_n23911_));
  AOI21_X1   g23845(.A1(new_n21136_), .A2(new_n21142_), .B(new_n19527_), .ZN(new_n23912_));
  NOR3_X1    g23846(.A1(new_n22213_), .A2(new_n22184_), .A3(new_n21162_), .ZN(new_n23913_));
  OAI22_X1   g23847(.A1(new_n23911_), .A2(new_n23912_), .B1(new_n23913_), .B2(new_n21144_), .ZN(new_n23914_));
  AOI21_X1   g23848(.A1(new_n23914_), .A2(new_n21988_), .B(new_n21978_), .ZN(new_n23915_));
  XOR2_X1    g23849(.A1(new_n23915_), .A2(new_n23910_), .Z(new_n23916_));
  NAND2_X1   g23850(.A1(new_n22159_), .A2(new_n22153_), .ZN(new_n23917_));
  AOI21_X1   g23851(.A1(new_n22124_), .A2(new_n22142_), .B(new_n22143_), .ZN(new_n23918_));
  NAND2_X1   g23852(.A1(new_n22136_), .A2(new_n22134_), .ZN(new_n23919_));
  NOR2_X1    g23853(.A1(new_n3155_), .A2(new_n3135_), .ZN(new_n23920_));
  NOR2_X1    g23854(.A1(new_n22130_), .A2(new_n23920_), .ZN(new_n23921_));
  INV_X1     g23855(.I(new_n23921_), .ZN(new_n23922_));
  INV_X1     g23856(.I(new_n23920_), .ZN(new_n23923_));
  NOR2_X1    g23857(.A1(new_n22133_), .A2(new_n23923_), .ZN(new_n23924_));
  INV_X1     g23858(.I(new_n23924_), .ZN(new_n23925_));
  AOI22_X1   g23859(.A1(new_n23919_), .A2(new_n22131_), .B1(new_n23922_), .B2(new_n23925_), .ZN(new_n23926_));
  NAND2_X1   g23860(.A1(new_n23919_), .A2(new_n22131_), .ZN(new_n23927_));
  XNOR2_X1   g23861(.A1(new_n22130_), .A2(new_n23920_), .ZN(new_n23928_));
  NOR2_X1    g23862(.A1(new_n23927_), .A2(new_n23928_), .ZN(new_n23929_));
  OAI21_X1   g23863(.A1(new_n3275_), .A2(new_n2750_), .B(new_n2746_), .ZN(new_n23930_));
  NOR2_X1    g23864(.A1(new_n11466_), .A2(new_n23930_), .ZN(new_n23931_));
  NOR4_X1    g23865(.A1(new_n11468_), .A2(new_n2737_), .A3(new_n11461_), .A4(new_n23931_), .ZN(new_n23932_));
  XOR2_X1    g23866(.A1(new_n23932_), .A2(\a[29] ), .Z(new_n23933_));
  NOR2_X1    g23867(.A1(new_n11369_), .A2(new_n2772_), .ZN(new_n23934_));
  AOI21_X1   g23868(.A1(new_n11346_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n23935_));
  OAI21_X1   g23869(.A1(new_n11353_), .A2(new_n2767_), .B(new_n23935_), .ZN(new_n23936_));
  NOR3_X1    g23870(.A1(new_n11379_), .A2(new_n23934_), .A3(new_n23936_), .ZN(new_n23937_));
  NOR2_X1    g23871(.A1(new_n23933_), .A2(new_n23937_), .ZN(new_n23938_));
  AND2_X2    g23872(.A1(new_n23933_), .A2(new_n23937_), .Z(new_n23939_));
  OAI22_X1   g23873(.A1(new_n23939_), .A2(new_n23938_), .B1(new_n23926_), .B2(new_n23929_), .ZN(new_n23940_));
  NOR2_X1    g23874(.A1(new_n23929_), .A2(new_n23926_), .ZN(new_n23941_));
  XOR2_X1    g23875(.A1(new_n23933_), .A2(new_n23937_), .Z(new_n23942_));
  NAND2_X1   g23876(.A1(new_n23942_), .A2(new_n23941_), .ZN(new_n23943_));
  NAND2_X1   g23877(.A1(new_n23943_), .A2(new_n23940_), .ZN(new_n23944_));
  XOR2_X1    g23878(.A1(new_n23944_), .A2(new_n23918_), .Z(new_n23945_));
  AND2_X2    g23879(.A1(new_n23945_), .A2(new_n22147_), .Z(new_n23946_));
  NOR2_X1    g23880(.A1(new_n23945_), .A2(new_n22147_), .ZN(new_n23947_));
  NOR2_X1    g23881(.A1(new_n23946_), .A2(new_n23947_), .ZN(new_n23948_));
  XOR2_X1    g23882(.A1(new_n23948_), .A2(new_n22150_), .Z(new_n23949_));
  AOI21_X1   g23883(.A1(new_n23917_), .A2(new_n22152_), .B(new_n23949_), .ZN(new_n23950_));
  INV_X1     g23884(.I(new_n22153_), .ZN(new_n23951_));
  NOR2_X1    g23885(.A1(new_n22117_), .A2(new_n23951_), .ZN(new_n23952_));
  XOR2_X1    g23886(.A1(new_n23948_), .A2(new_n22149_), .Z(new_n23953_));
  NOR3_X1    g23887(.A1(new_n23952_), .A2(new_n22151_), .A3(new_n23953_), .ZN(new_n23954_));
  OR2_X2     g23888(.A1(new_n23954_), .A2(new_n23950_), .Z(new_n23955_));
  OAI22_X1   g23889(.A1(new_n22115_), .A2(new_n9485_), .B1(new_n9483_), .B2(new_n22149_), .ZN(new_n23956_));
  INV_X1     g23890(.I(new_n23948_), .ZN(new_n23957_));
  NAND2_X1   g23891(.A1(new_n23957_), .A2(new_n9488_), .ZN(new_n23958_));
  AOI21_X1   g23892(.A1(new_n23956_), .A2(new_n23958_), .B(new_n9482_), .ZN(new_n23959_));
  NAND2_X1   g23893(.A1(new_n23955_), .A2(new_n23959_), .ZN(new_n23960_));
  XOR2_X1    g23894(.A1(new_n23960_), .A2(\a[2] ), .Z(new_n23961_));
  XNOR2_X1   g23895(.A1(new_n23916_), .A2(new_n23961_), .ZN(new_n23962_));
  INV_X1     g23896(.I(new_n23962_), .ZN(new_n23963_));
  OAI21_X1   g23897(.A1(new_n23713_), .A2(new_n23696_), .B(new_n23963_), .ZN(new_n23964_));
  NOR3_X1    g23898(.A1(new_n23709_), .A2(new_n23710_), .A3(new_n23711_), .ZN(new_n23965_));
  AOI21_X1   g23899(.A1(new_n23706_), .A2(new_n23701_), .B(new_n23707_), .ZN(new_n23966_));
  NOR3_X1    g23900(.A1(new_n23696_), .A2(new_n23965_), .A3(new_n23966_), .ZN(new_n23967_));
  NAND2_X1   g23901(.A1(new_n23967_), .A2(new_n23962_), .ZN(new_n23968_));
  NAND2_X1   g23902(.A1(new_n23968_), .A2(new_n23964_), .ZN(\result[1] ));
  OAI21_X1   g23903(.A1(new_n21761_), .A2(new_n23729_), .B(new_n21795_), .ZN(new_n23970_));
  INV_X1     g23904(.I(new_n23775_), .ZN(new_n23971_));
  AOI21_X1   g23905(.A1(new_n23970_), .A2(new_n23971_), .B(new_n23777_), .ZN(new_n23972_));
  AOI21_X1   g23906(.A1(new_n23734_), .A2(new_n23749_), .B(new_n23750_), .ZN(new_n23973_));
  INV_X1     g23907(.I(new_n23973_), .ZN(new_n23974_));
  AOI21_X1   g23908(.A1(new_n19321_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n23975_));
  OAI21_X1   g23909(.A1(new_n17828_), .A2(new_n2767_), .B(new_n23975_), .ZN(new_n23976_));
  AOI21_X1   g23910(.A1(new_n3332_), .A2(new_n19349_), .B(new_n23976_), .ZN(new_n23977_));
  NAND2_X1   g23911(.A1(new_n19760_), .A2(new_n23977_), .ZN(new_n23978_));
  INV_X1     g23912(.I(new_n1551_), .ZN(new_n23979_));
  NOR4_X1    g23913(.A1(new_n1257_), .A2(new_n254_), .A3(new_n23979_), .A4(new_n2284_), .ZN(new_n23980_));
  NOR4_X1    g23914(.A1(new_n1969_), .A2(new_n11816_), .A3(new_n214_), .A4(new_n376_), .ZN(new_n23981_));
  NAND3_X1   g23915(.A1(new_n23980_), .A2(new_n2218_), .A3(new_n23981_), .ZN(new_n23982_));
  INV_X1     g23916(.I(new_n23982_), .ZN(new_n23983_));
  NAND2_X1   g23917(.A1(new_n11489_), .A2(new_n1173_), .ZN(new_n23984_));
  NOR4_X1    g23918(.A1(new_n2963_), .A2(new_n23984_), .A3(new_n4861_), .A4(new_n12032_), .ZN(new_n23985_));
  NAND4_X1   g23919(.A1(new_n2196_), .A2(new_n23983_), .A3(new_n23985_), .A4(new_n2980_), .ZN(new_n23986_));
  NAND2_X1   g23920(.A1(new_n23978_), .A2(new_n23986_), .ZN(new_n23987_));
  NOR2_X1    g23921(.A1(new_n23978_), .A2(new_n23986_), .ZN(new_n23988_));
  INV_X1     g23922(.I(new_n23988_), .ZN(new_n23989_));
  NAND2_X1   g23923(.A1(new_n23989_), .A2(new_n23987_), .ZN(new_n23990_));
  XNOR2_X1   g23924(.A1(new_n23978_), .A2(new_n23986_), .ZN(new_n23991_));
  NOR2_X1    g23925(.A1(new_n23974_), .A2(new_n23991_), .ZN(new_n23992_));
  AOI21_X1   g23926(.A1(new_n23974_), .A2(new_n23990_), .B(new_n23992_), .ZN(new_n23993_));
  OAI22_X1   g23927(.A1(new_n17806_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19346_), .ZN(new_n23994_));
  NAND2_X1   g23928(.A1(new_n19359_), .A2(new_n2750_), .ZN(new_n23995_));
  AOI21_X1   g23929(.A1(new_n23995_), .A2(new_n23994_), .B(new_n2737_), .ZN(new_n23996_));
  NAND2_X1   g23930(.A1(new_n20096_), .A2(new_n23996_), .ZN(new_n23997_));
  NOR2_X1    g23931(.A1(new_n23997_), .A2(\a[29] ), .ZN(new_n23998_));
  NAND2_X1   g23932(.A1(new_n23997_), .A2(\a[29] ), .ZN(new_n23999_));
  INV_X1     g23933(.I(new_n23999_), .ZN(new_n24000_));
  NOR3_X1    g23934(.A1(new_n24000_), .A2(new_n23993_), .A3(new_n23998_), .ZN(new_n24001_));
  NAND2_X1   g23935(.A1(new_n23974_), .A2(new_n23990_), .ZN(new_n24002_));
  OAI21_X1   g23936(.A1(new_n23974_), .A2(new_n23991_), .B(new_n24002_), .ZN(new_n24003_));
  INV_X1     g23937(.I(new_n23998_), .ZN(new_n24004_));
  AOI21_X1   g23938(.A1(new_n24004_), .A2(new_n23999_), .B(new_n24003_), .ZN(new_n24005_));
  NOR2_X1    g23939(.A1(new_n24005_), .A2(new_n24001_), .ZN(new_n24006_));
  NOR2_X1    g23940(.A1(new_n24006_), .A2(new_n23972_), .ZN(new_n24007_));
  NAND3_X1   g23941(.A1(new_n24004_), .A2(new_n23993_), .A3(new_n23999_), .ZN(new_n24008_));
  OAI21_X1   g23942(.A1(new_n24000_), .A2(new_n23998_), .B(new_n24003_), .ZN(new_n24009_));
  NAND2_X1   g23943(.A1(new_n24009_), .A2(new_n24008_), .ZN(new_n24010_));
  AOI21_X1   g23944(.A1(new_n23972_), .A2(new_n24010_), .B(new_n24007_), .ZN(new_n24011_));
  INV_X1     g23945(.I(new_n24011_), .ZN(new_n24012_));
  AOI22_X1   g23946(.A1(new_n17802_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n19365_), .ZN(new_n24013_));
  NOR2_X1    g23947(.A1(new_n17797_), .A2(new_n3318_), .ZN(new_n24014_));
  OAI21_X1   g23948(.A1(new_n24014_), .A2(new_n24013_), .B(new_n3259_), .ZN(new_n24015_));
  NOR3_X1    g23949(.A1(new_n21454_), .A2(\a[26] ), .A3(new_n24015_), .ZN(new_n24016_));
  INV_X1     g23950(.I(new_n24015_), .ZN(new_n24017_));
  AOI21_X1   g23951(.A1(new_n20051_), .A2(new_n24017_), .B(new_n72_), .ZN(new_n24018_));
  NOR2_X1    g23952(.A1(new_n24016_), .A2(new_n24018_), .ZN(new_n24019_));
  OAI21_X1   g23953(.A1(new_n21792_), .A2(new_n21796_), .B(new_n21802_), .ZN(new_n24020_));
  NAND3_X1   g23954(.A1(new_n23787_), .A2(new_n23784_), .A3(new_n24020_), .ZN(new_n24021_));
  NAND2_X1   g23955(.A1(new_n24021_), .A2(new_n24019_), .ZN(new_n24022_));
  INV_X1     g23956(.I(new_n24019_), .ZN(new_n24023_));
  NAND4_X1   g23957(.A1(new_n24023_), .A2(new_n23787_), .A3(new_n23784_), .A4(new_n24020_), .ZN(new_n24024_));
  AOI21_X1   g23958(.A1(new_n24022_), .A2(new_n24024_), .B(new_n24012_), .ZN(new_n24025_));
  INV_X1     g23959(.I(new_n24020_), .ZN(new_n24026_));
  NOR3_X1    g23960(.A1(new_n23790_), .A2(new_n23791_), .A3(new_n24026_), .ZN(new_n24027_));
  NOR2_X1    g23961(.A1(new_n24027_), .A2(new_n24023_), .ZN(new_n24028_));
  NOR2_X1    g23962(.A1(new_n24021_), .A2(new_n24019_), .ZN(new_n24029_));
  NOR3_X1    g23963(.A1(new_n24028_), .A2(new_n24029_), .A3(new_n24011_), .ZN(new_n24030_));
  NOR2_X1    g23964(.A1(new_n24030_), .A2(new_n24025_), .ZN(new_n24031_));
  OAI22_X1   g23965(.A1(new_n19385_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19375_), .ZN(new_n24032_));
  NAND2_X1   g23966(.A1(new_n17794_), .A2(new_n3312_), .ZN(new_n24033_));
  AOI21_X1   g23967(.A1(new_n24032_), .A2(new_n24033_), .B(new_n3302_), .ZN(new_n24034_));
  NAND2_X1   g23968(.A1(new_n20134_), .A2(new_n24034_), .ZN(new_n24035_));
  XOR2_X1    g23969(.A1(new_n24035_), .A2(new_n84_), .Z(new_n24036_));
  NAND3_X1   g23970(.A1(new_n23720_), .A2(new_n23803_), .A3(new_n23718_), .ZN(new_n24037_));
  AOI21_X1   g23971(.A1(new_n24037_), .A2(new_n23793_), .B(new_n24036_), .ZN(new_n24038_));
  XOR2_X1    g23972(.A1(new_n24035_), .A2(\a[23] ), .Z(new_n24039_));
  NOR3_X1    g23973(.A1(new_n23800_), .A2(new_n21812_), .A3(new_n23798_), .ZN(new_n24040_));
  NOR3_X1    g23974(.A1(new_n24040_), .A2(new_n23801_), .A3(new_n24039_), .ZN(new_n24041_));
  OAI21_X1   g23975(.A1(new_n24041_), .A2(new_n24038_), .B(new_n24031_), .ZN(new_n24042_));
  INV_X1     g23976(.I(new_n24031_), .ZN(new_n24043_));
  OAI21_X1   g23977(.A1(new_n24040_), .A2(new_n23801_), .B(new_n24039_), .ZN(new_n24044_));
  NAND3_X1   g23978(.A1(new_n24037_), .A2(new_n23793_), .A3(new_n24036_), .ZN(new_n24045_));
  NAND3_X1   g23979(.A1(new_n24044_), .A2(new_n24045_), .A3(new_n24043_), .ZN(new_n24046_));
  NAND2_X1   g23980(.A1(new_n24042_), .A2(new_n24046_), .ZN(new_n24047_));
  OAI22_X1   g23981(.A1(new_n19400_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19393_), .ZN(new_n24048_));
  NAND2_X1   g23982(.A1(new_n17790_), .A2(new_n4096_), .ZN(new_n24049_));
  AOI21_X1   g23983(.A1(new_n24049_), .A2(new_n24048_), .B(new_n4095_), .ZN(new_n24050_));
  NAND2_X1   g23984(.A1(new_n20251_), .A2(new_n24050_), .ZN(new_n24051_));
  XOR2_X1    g23985(.A1(new_n24051_), .A2(new_n3035_), .Z(new_n24052_));
  INV_X1     g23986(.I(new_n24052_), .ZN(new_n24053_));
  OAI21_X1   g23987(.A1(new_n23819_), .A2(new_n23820_), .B(new_n23814_), .ZN(new_n24054_));
  NAND2_X1   g23988(.A1(new_n24054_), .A2(new_n24053_), .ZN(new_n24055_));
  NAND3_X1   g23989(.A1(new_n23815_), .A2(new_n23814_), .A3(new_n24052_), .ZN(new_n24056_));
  AOI21_X1   g23990(.A1(new_n24055_), .A2(new_n24056_), .B(new_n24047_), .ZN(new_n24057_));
  AOI21_X1   g23991(.A1(new_n24044_), .A2(new_n24045_), .B(new_n24043_), .ZN(new_n24058_));
  NOR3_X1    g23992(.A1(new_n24041_), .A2(new_n24038_), .A3(new_n24031_), .ZN(new_n24059_));
  NOR2_X1    g23993(.A1(new_n24059_), .A2(new_n24058_), .ZN(new_n24060_));
  AOI21_X1   g23994(.A1(new_n23815_), .A2(new_n23814_), .B(new_n24052_), .ZN(new_n24061_));
  NOR2_X1    g23995(.A1(new_n24054_), .A2(new_n24053_), .ZN(new_n24062_));
  NOR3_X1    g23996(.A1(new_n24061_), .A2(new_n24062_), .A3(new_n24060_), .ZN(new_n24063_));
  NOR2_X1    g23997(.A1(new_n24063_), .A2(new_n24057_), .ZN(new_n24064_));
  OAI22_X1   g23998(.A1(new_n19410_), .A2(new_n4291_), .B1(new_n19412_), .B2(new_n4297_), .ZN(new_n24065_));
  NAND2_X1   g23999(.A1(new_n19439_), .A2(new_n4469_), .ZN(new_n24066_));
  AOI21_X1   g24000(.A1(new_n24066_), .A2(new_n24065_), .B(new_n4468_), .ZN(new_n24067_));
  NAND2_X1   g24001(.A1(new_n20827_), .A2(new_n24067_), .ZN(new_n24068_));
  XOR2_X1    g24002(.A1(new_n24068_), .A2(new_n3372_), .Z(new_n24069_));
  NOR3_X1    g24003(.A1(new_n23839_), .A2(new_n23836_), .A3(new_n23833_), .ZN(new_n24070_));
  NOR2_X1    g24004(.A1(new_n24070_), .A2(new_n24069_), .ZN(new_n24071_));
  NAND4_X1   g24005(.A1(new_n23834_), .A2(new_n23829_), .A3(new_n23838_), .A4(new_n24069_), .ZN(new_n24072_));
  INV_X1     g24006(.I(new_n24072_), .ZN(new_n24073_));
  OAI21_X1   g24007(.A1(new_n24071_), .A2(new_n24073_), .B(new_n24064_), .ZN(new_n24074_));
  INV_X1     g24008(.I(new_n24064_), .ZN(new_n24075_));
  XOR2_X1    g24009(.A1(new_n24068_), .A2(\a[17] ), .Z(new_n24076_));
  NAND3_X1   g24010(.A1(new_n23834_), .A2(new_n23829_), .A3(new_n23838_), .ZN(new_n24077_));
  NAND2_X1   g24011(.A1(new_n24077_), .A2(new_n24076_), .ZN(new_n24078_));
  NAND3_X1   g24012(.A1(new_n24078_), .A2(new_n24075_), .A3(new_n24072_), .ZN(new_n24079_));
  NAND2_X1   g24013(.A1(new_n24074_), .A2(new_n24079_), .ZN(new_n24080_));
  OAI22_X1   g24014(.A1(new_n19428_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n19423_), .ZN(new_n24081_));
  NAND2_X1   g24015(.A1(new_n19438_), .A2(new_n6090_), .ZN(new_n24082_));
  AOI21_X1   g24016(.A1(new_n24082_), .A2(new_n24081_), .B(new_n6082_), .ZN(new_n24083_));
  NAND2_X1   g24017(.A1(new_n20907_), .A2(new_n24083_), .ZN(new_n24084_));
  XOR2_X1    g24018(.A1(new_n24084_), .A2(\a[14] ), .Z(new_n24085_));
  OAI21_X1   g24019(.A1(new_n23715_), .A2(new_n23846_), .B(new_n23855_), .ZN(new_n24086_));
  NAND2_X1   g24020(.A1(new_n24086_), .A2(new_n24085_), .ZN(new_n24087_));
  INV_X1     g24021(.I(new_n24085_), .ZN(new_n24088_));
  NAND3_X1   g24022(.A1(new_n23863_), .A2(new_n23855_), .A3(new_n24088_), .ZN(new_n24089_));
  AOI21_X1   g24023(.A1(new_n24087_), .A2(new_n24089_), .B(new_n24080_), .ZN(new_n24090_));
  AOI21_X1   g24024(.A1(new_n24078_), .A2(new_n24072_), .B(new_n24075_), .ZN(new_n24091_));
  NOR3_X1    g24025(.A1(new_n24071_), .A2(new_n24073_), .A3(new_n24064_), .ZN(new_n24092_));
  NOR2_X1    g24026(.A1(new_n24092_), .A2(new_n24091_), .ZN(new_n24093_));
  AOI21_X1   g24027(.A1(new_n23863_), .A2(new_n23855_), .B(new_n24088_), .ZN(new_n24094_));
  NOR2_X1    g24028(.A1(new_n24086_), .A2(new_n24085_), .ZN(new_n24095_));
  NOR3_X1    g24029(.A1(new_n24095_), .A2(new_n24094_), .A3(new_n24093_), .ZN(new_n24096_));
  NOR2_X1    g24030(.A1(new_n24096_), .A2(new_n24090_), .ZN(new_n24097_));
  OAI22_X1   g24031(.A1(new_n19463_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n19437_), .ZN(new_n24098_));
  NAND2_X1   g24032(.A1(new_n17780_), .A2(new_n4709_), .ZN(new_n24099_));
  AOI21_X1   g24033(.A1(new_n24098_), .A2(new_n24099_), .B(new_n4707_), .ZN(new_n24100_));
  NAND2_X1   g24034(.A1(new_n21088_), .A2(new_n24100_), .ZN(new_n24101_));
  XOR2_X1    g24035(.A1(new_n24101_), .A2(new_n4034_), .Z(new_n24102_));
  NOR3_X1    g24036(.A1(new_n23868_), .A2(new_n23862_), .A3(new_n23872_), .ZN(new_n24103_));
  NOR2_X1    g24037(.A1(new_n24103_), .A2(new_n24102_), .ZN(new_n24104_));
  XOR2_X1    g24038(.A1(new_n24101_), .A2(\a[11] ), .Z(new_n24105_));
  NOR4_X1    g24039(.A1(new_n23868_), .A2(new_n23862_), .A3(new_n23872_), .A4(new_n24105_), .ZN(new_n24106_));
  OAI21_X1   g24040(.A1(new_n24104_), .A2(new_n24106_), .B(new_n24097_), .ZN(new_n24107_));
  INV_X1     g24041(.I(new_n24097_), .ZN(new_n24108_));
  NAND3_X1   g24042(.A1(new_n23873_), .A2(new_n23870_), .A3(new_n23871_), .ZN(new_n24109_));
  NAND2_X1   g24043(.A1(new_n24109_), .A2(new_n24105_), .ZN(new_n24110_));
  NAND4_X1   g24044(.A1(new_n23873_), .A2(new_n23870_), .A3(new_n23867_), .A4(new_n24102_), .ZN(new_n24111_));
  NAND3_X1   g24045(.A1(new_n24110_), .A2(new_n24108_), .A3(new_n24111_), .ZN(new_n24112_));
  NAND2_X1   g24046(.A1(new_n24107_), .A2(new_n24112_), .ZN(new_n24113_));
  OAI22_X1   g24047(.A1(new_n19522_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n17775_), .ZN(new_n24114_));
  NAND2_X1   g24048(.A1(new_n17770_), .A2(new_n6784_), .ZN(new_n24115_));
  AOI21_X1   g24049(.A1(new_n24115_), .A2(new_n24114_), .B(new_n6776_), .ZN(new_n24116_));
  NAND2_X1   g24050(.A1(new_n19521_), .A2(new_n24116_), .ZN(new_n24117_));
  XOR2_X1    g24051(.A1(new_n24117_), .A2(\a[8] ), .Z(new_n24118_));
  NAND3_X1   g24052(.A1(new_n23887_), .A2(new_n23882_), .A3(new_n23892_), .ZN(new_n24119_));
  NAND2_X1   g24053(.A1(new_n24119_), .A2(new_n24118_), .ZN(new_n24120_));
  INV_X1     g24054(.I(new_n24118_), .ZN(new_n24121_));
  NAND4_X1   g24055(.A1(new_n24121_), .A2(new_n23887_), .A3(new_n23882_), .A4(new_n23892_), .ZN(new_n24122_));
  AOI21_X1   g24056(.A1(new_n24120_), .A2(new_n24122_), .B(new_n24113_), .ZN(new_n24123_));
  AOI21_X1   g24057(.A1(new_n24110_), .A2(new_n24111_), .B(new_n24108_), .ZN(new_n24124_));
  NOR3_X1    g24058(.A1(new_n24104_), .A2(new_n24097_), .A3(new_n24106_), .ZN(new_n24125_));
  NOR2_X1    g24059(.A1(new_n24125_), .A2(new_n24124_), .ZN(new_n24126_));
  NOR3_X1    g24060(.A1(new_n23891_), .A2(new_n23890_), .A3(new_n23888_), .ZN(new_n24127_));
  NOR2_X1    g24061(.A1(new_n24127_), .A2(new_n24121_), .ZN(new_n24128_));
  NOR4_X1    g24062(.A1(new_n23891_), .A2(new_n23890_), .A3(new_n23888_), .A4(new_n24118_), .ZN(new_n24129_));
  NOR3_X1    g24063(.A1(new_n24128_), .A2(new_n24126_), .A3(new_n24129_), .ZN(new_n24130_));
  NOR2_X1    g24064(.A1(new_n24123_), .A2(new_n24130_), .ZN(new_n24131_));
  AOI22_X1   g24065(.A1(new_n22048_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n21953_), .ZN(new_n24132_));
  AOI21_X1   g24066(.A1(new_n22118_), .A2(new_n6838_), .B(new_n24132_), .ZN(new_n24133_));
  NOR4_X1    g24067(.A1(new_n23672_), .A2(new_n6836_), .A3(new_n23673_), .A4(new_n24133_), .ZN(new_n24134_));
  XOR2_X1    g24068(.A1(new_n24134_), .A2(new_n65_), .Z(new_n24135_));
  INV_X1     g24069(.I(new_n21978_), .ZN(new_n24136_));
  OAI21_X1   g24070(.A1(new_n21747_), .A2(new_n21987_), .B(new_n24136_), .ZN(new_n24137_));
  NAND3_X1   g24071(.A1(new_n24137_), .A2(new_n23905_), .A3(new_n23909_), .ZN(new_n24138_));
  XOR2_X1    g24072(.A1(new_n24138_), .A2(new_n24135_), .Z(new_n24139_));
  XNOR2_X1   g24073(.A1(new_n24139_), .A2(new_n24131_), .ZN(new_n24140_));
  NOR2_X1    g24074(.A1(new_n23938_), .A2(new_n23941_), .ZN(new_n24141_));
  NOR2_X1    g24075(.A1(new_n24141_), .A2(new_n23939_), .ZN(new_n24142_));
  NAND2_X1   g24076(.A1(new_n23927_), .A2(new_n23925_), .ZN(new_n24143_));
  NAND2_X1   g24077(.A1(new_n24143_), .A2(new_n23922_), .ZN(new_n24144_));
  NOR2_X1    g24078(.A1(new_n11369_), .A2(new_n2767_), .ZN(new_n24145_));
  NOR2_X1    g24079(.A1(new_n11697_), .A2(new_n2772_), .ZN(new_n24146_));
  NOR2_X1    g24080(.A1(new_n11353_), .A2(new_n2771_), .ZN(new_n24147_));
  NOR4_X1    g24081(.A1(new_n24145_), .A2(new_n2763_), .A3(new_n24146_), .A4(new_n24147_), .ZN(new_n24148_));
  NAND2_X1   g24082(.A1(new_n11700_), .A2(new_n24148_), .ZN(new_n24149_));
  NOR2_X1    g24083(.A1(new_n2738_), .A2(new_n2740_), .ZN(new_n24150_));
  NAND4_X1   g24084(.A1(new_n11226_), .A2(new_n2734_), .A3(new_n2735_), .A4(new_n24150_), .ZN(new_n24151_));
  XOR2_X1    g24085(.A1(new_n24151_), .A2(new_n11222_), .Z(new_n24152_));
  XOR2_X1    g24086(.A1(new_n24152_), .A2(\a[29] ), .Z(new_n24153_));
  XOR2_X1    g24087(.A1(new_n24153_), .A2(new_n23920_), .Z(new_n24154_));
  INV_X1     g24088(.I(new_n24154_), .ZN(new_n24155_));
  XOR2_X1    g24089(.A1(new_n24149_), .A2(new_n24155_), .Z(new_n24156_));
  NAND2_X1   g24090(.A1(new_n24144_), .A2(new_n24156_), .ZN(new_n24157_));
  XOR2_X1    g24091(.A1(new_n24149_), .A2(new_n24155_), .Z(new_n24158_));
  OAI21_X1   g24092(.A1(new_n24144_), .A2(new_n24158_), .B(new_n24157_), .ZN(new_n24159_));
  INV_X1     g24093(.I(new_n23918_), .ZN(new_n24160_));
  NOR2_X1    g24094(.A1(new_n23944_), .A2(new_n24160_), .ZN(new_n24161_));
  NOR2_X1    g24095(.A1(new_n24161_), .A2(new_n22147_), .ZN(new_n24162_));
  XNOR2_X1   g24096(.A1(new_n24162_), .A2(new_n24159_), .ZN(new_n24163_));
  NAND2_X1   g24097(.A1(new_n24163_), .A2(new_n24142_), .ZN(new_n24164_));
  INV_X1     g24098(.I(new_n24164_), .ZN(new_n24165_));
  NOR2_X1    g24099(.A1(new_n24163_), .A2(new_n24142_), .ZN(new_n24166_));
  NOR2_X1    g24100(.A1(new_n24165_), .A2(new_n24166_), .ZN(new_n24167_));
  INV_X1     g24101(.I(new_n23949_), .ZN(new_n24168_));
  AOI21_X1   g24102(.A1(new_n22159_), .A2(new_n22115_), .B(new_n22149_), .ZN(new_n24169_));
  AOI21_X1   g24103(.A1(new_n22117_), .A2(new_n22118_), .B(new_n22150_), .ZN(new_n24170_));
  OAI21_X1   g24104(.A1(new_n24170_), .A2(new_n24169_), .B(new_n24168_), .ZN(new_n24171_));
  XOR2_X1    g24105(.A1(new_n24171_), .A2(new_n24167_), .Z(new_n24172_));
  OAI22_X1   g24106(.A1(new_n23948_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n22149_), .ZN(new_n24173_));
  INV_X1     g24107(.I(new_n24167_), .ZN(new_n24174_));
  NAND2_X1   g24108(.A1(new_n24174_), .A2(new_n9488_), .ZN(new_n24175_));
  AOI21_X1   g24109(.A1(new_n24175_), .A2(new_n24173_), .B(new_n9482_), .ZN(new_n24176_));
  NAND2_X1   g24110(.A1(new_n24172_), .A2(new_n24176_), .ZN(new_n24177_));
  XOR2_X1    g24111(.A1(new_n24177_), .A2(\a[2] ), .Z(new_n24178_));
  XOR2_X1    g24112(.A1(new_n24140_), .A2(new_n24178_), .Z(new_n24179_));
  NOR2_X1    g24113(.A1(new_n23916_), .A2(new_n23961_), .ZN(new_n24180_));
  XOR2_X1    g24114(.A1(new_n24179_), .A2(new_n24180_), .Z(new_n24181_));
  XOR2_X1    g24115(.A1(new_n23964_), .A2(new_n24181_), .Z(\result[2] ));
  NOR2_X1    g24116(.A1(new_n23964_), .A2(new_n24181_), .ZN(new_n24183_));
  XOR2_X1    g24117(.A1(new_n24134_), .A2(\a[5] ), .Z(new_n24184_));
  OAI21_X1   g24118(.A1(new_n24128_), .A2(new_n24129_), .B(new_n24126_), .ZN(new_n24185_));
  NAND3_X1   g24119(.A1(new_n24120_), .A2(new_n24113_), .A3(new_n24122_), .ZN(new_n24186_));
  NAND3_X1   g24120(.A1(new_n24185_), .A2(new_n24186_), .A3(new_n24184_), .ZN(new_n24187_));
  OAI21_X1   g24121(.A1(new_n24123_), .A2(new_n24130_), .B(new_n24135_), .ZN(new_n24188_));
  AOI22_X1   g24122(.A1(new_n24138_), .A2(new_n24184_), .B1(new_n24188_), .B2(new_n24187_), .ZN(new_n24189_));
  NOR2_X1    g24123(.A1(new_n24031_), .A2(new_n24036_), .ZN(new_n24190_));
  OAI21_X1   g24124(.A1(new_n24028_), .A2(new_n24029_), .B(new_n24011_), .ZN(new_n24191_));
  NAND3_X1   g24125(.A1(new_n24022_), .A2(new_n24012_), .A3(new_n24024_), .ZN(new_n24192_));
  NAND3_X1   g24126(.A1(new_n24191_), .A2(new_n24192_), .A3(new_n24036_), .ZN(new_n24193_));
  OAI21_X1   g24127(.A1(new_n24030_), .A2(new_n24025_), .B(new_n24039_), .ZN(new_n24194_));
  AOI21_X1   g24128(.A1(new_n24194_), .A2(new_n24193_), .B(new_n23801_), .ZN(new_n24195_));
  AOI21_X1   g24129(.A1(new_n24195_), .A2(new_n24037_), .B(new_n24190_), .ZN(new_n24196_));
  OAI21_X1   g24130(.A1(new_n23774_), .A2(new_n23775_), .B(new_n23776_), .ZN(new_n24197_));
  AOI21_X1   g24131(.A1(new_n24004_), .A2(new_n23999_), .B(new_n23993_), .ZN(new_n24198_));
  AOI21_X1   g24132(.A1(new_n24197_), .A2(new_n24008_), .B(new_n24198_), .ZN(new_n24199_));
  INV_X1     g24133(.I(new_n23987_), .ZN(new_n24200_));
  OAI21_X1   g24134(.A1(new_n23973_), .A2(new_n24200_), .B(new_n23989_), .ZN(new_n24201_));
  NAND2_X1   g24135(.A1(new_n19349_), .A2(new_n3189_), .ZN(new_n24202_));
  NAND2_X1   g24136(.A1(new_n2762_), .A2(\a[31] ), .ZN(new_n24203_));
  AOI21_X1   g24137(.A1(new_n17827_), .A2(new_n2770_), .B(new_n24203_), .ZN(new_n24204_));
  NAND3_X1   g24138(.A1(new_n20535_), .A2(new_n24202_), .A3(new_n24204_), .ZN(new_n24205_));
  NOR4_X1    g24139(.A1(new_n837_), .A2(new_n170_), .A3(new_n306_), .A4(new_n506_), .ZN(new_n24206_));
  NAND4_X1   g24140(.A1(new_n2286_), .A2(new_n3678_), .A3(new_n24206_), .A4(new_n2297_), .ZN(new_n24207_));
  NOR4_X1    g24141(.A1(new_n4886_), .A2(new_n525_), .A3(new_n491_), .A4(new_n561_), .ZN(new_n24208_));
  NAND4_X1   g24142(.A1(new_n24208_), .A2(new_n537_), .A3(new_n957_), .A4(new_n1551_), .ZN(new_n24209_));
  NOR3_X1    g24143(.A1(new_n24209_), .A2(new_n24207_), .A3(new_n12801_), .ZN(new_n24210_));
  NAND4_X1   g24144(.A1(new_n4868_), .A2(new_n24210_), .A3(new_n2015_), .A4(new_n2890_), .ZN(new_n24211_));
  NAND2_X1   g24145(.A1(new_n24205_), .A2(new_n24211_), .ZN(new_n24212_));
  NOR2_X1    g24146(.A1(new_n24205_), .A2(new_n24211_), .ZN(new_n24213_));
  INV_X1     g24147(.I(new_n24213_), .ZN(new_n24214_));
  NAND2_X1   g24148(.A1(new_n24214_), .A2(new_n24212_), .ZN(new_n24215_));
  XNOR2_X1   g24149(.A1(new_n24205_), .A2(new_n24211_), .ZN(new_n24216_));
  NOR2_X1    g24150(.A1(new_n24216_), .A2(new_n24201_), .ZN(new_n24217_));
  AOI21_X1   g24151(.A1(new_n24201_), .A2(new_n24215_), .B(new_n24217_), .ZN(new_n24218_));
  AOI22_X1   g24152(.A1(new_n19359_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n17807_), .ZN(new_n24219_));
  NOR2_X1    g24153(.A1(new_n19364_), .A2(new_n3175_), .ZN(new_n24220_));
  OAI21_X1   g24154(.A1(new_n24219_), .A2(new_n24220_), .B(new_n2736_), .ZN(new_n24221_));
  INV_X1     g24155(.I(new_n24221_), .ZN(new_n24222_));
  NAND3_X1   g24156(.A1(new_n19538_), .A2(new_n74_), .A3(new_n24222_), .ZN(new_n24223_));
  INV_X1     g24157(.I(new_n24223_), .ZN(new_n24224_));
  AOI21_X1   g24158(.A1(new_n19538_), .A2(new_n24222_), .B(new_n74_), .ZN(new_n24225_));
  NOR2_X1    g24159(.A1(new_n24224_), .A2(new_n24225_), .ZN(new_n24226_));
  INV_X1     g24160(.I(new_n24226_), .ZN(new_n24227_));
  XOR2_X1    g24161(.A1(new_n24218_), .A2(new_n24227_), .Z(new_n24228_));
  NAND2_X1   g24162(.A1(new_n24215_), .A2(new_n24201_), .ZN(new_n24229_));
  OAI21_X1   g24163(.A1(new_n24201_), .A2(new_n24216_), .B(new_n24229_), .ZN(new_n24230_));
  NOR2_X1    g24164(.A1(new_n24227_), .A2(new_n24230_), .ZN(new_n24231_));
  NOR2_X1    g24165(.A1(new_n24218_), .A2(new_n24226_), .ZN(new_n24232_));
  OAI21_X1   g24166(.A1(new_n24231_), .A2(new_n24232_), .B(new_n24199_), .ZN(new_n24233_));
  OAI21_X1   g24167(.A1(new_n24199_), .A2(new_n24228_), .B(new_n24233_), .ZN(new_n24234_));
  AOI22_X1   g24168(.A1(new_n17798_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n17802_), .ZN(new_n24235_));
  NOR2_X1    g24169(.A1(new_n19375_), .A2(new_n3318_), .ZN(new_n24236_));
  OAI21_X1   g24170(.A1(new_n24236_), .A2(new_n24235_), .B(new_n3259_), .ZN(new_n24237_));
  NOR2_X1    g24171(.A1(new_n21753_), .A2(new_n24237_), .ZN(new_n24238_));
  XOR2_X1    g24172(.A1(new_n24238_), .A2(new_n72_), .Z(new_n24239_));
  XOR2_X1    g24173(.A1(new_n24234_), .A2(new_n24239_), .Z(new_n24240_));
  AOI22_X1   g24174(.A1(new_n19386_), .A2(new_n5291_), .B1(new_n3782_), .B2(new_n17794_), .ZN(new_n24241_));
  NOR2_X1    g24175(.A1(new_n19393_), .A2(new_n3780_), .ZN(new_n24242_));
  OAI21_X1   g24176(.A1(new_n24241_), .A2(new_n24242_), .B(new_n3301_), .ZN(new_n24243_));
  NOR2_X1    g24177(.A1(new_n20291_), .A2(new_n24243_), .ZN(new_n24244_));
  XOR2_X1    g24178(.A1(new_n24244_), .A2(\a[23] ), .Z(new_n24245_));
  NOR2_X1    g24179(.A1(new_n24240_), .A2(new_n24245_), .ZN(new_n24246_));
  INV_X1     g24180(.I(new_n24246_), .ZN(new_n24247_));
  NAND2_X1   g24181(.A1(new_n24240_), .A2(new_n24245_), .ZN(new_n24248_));
  NAND2_X1   g24182(.A1(new_n24247_), .A2(new_n24248_), .ZN(new_n24249_));
  NAND2_X1   g24183(.A1(new_n24196_), .A2(new_n24249_), .ZN(new_n24250_));
  NOR3_X1    g24184(.A1(new_n24030_), .A2(new_n24025_), .A3(new_n24039_), .ZN(new_n24251_));
  AOI21_X1   g24185(.A1(new_n24191_), .A2(new_n24192_), .B(new_n24036_), .ZN(new_n24252_));
  OAI21_X1   g24186(.A1(new_n24252_), .A2(new_n24251_), .B(new_n23793_), .ZN(new_n24253_));
  OAI22_X1   g24187(.A1(new_n24253_), .A2(new_n24040_), .B1(new_n24031_), .B2(new_n24036_), .ZN(new_n24254_));
  XOR2_X1    g24188(.A1(new_n24240_), .A2(new_n24245_), .Z(new_n24255_));
  NAND2_X1   g24189(.A1(new_n24254_), .A2(new_n24255_), .ZN(new_n24256_));
  NAND2_X1   g24190(.A1(new_n24256_), .A2(new_n24250_), .ZN(new_n24257_));
  OAI22_X1   g24191(.A1(new_n17789_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19400_), .ZN(new_n24258_));
  NAND2_X1   g24192(.A1(new_n19407_), .A2(new_n4096_), .ZN(new_n24259_));
  AOI21_X1   g24193(.A1(new_n24259_), .A2(new_n24258_), .B(new_n4095_), .ZN(new_n24260_));
  NAND2_X1   g24194(.A1(new_n20864_), .A2(new_n24260_), .ZN(new_n24261_));
  XOR2_X1    g24195(.A1(new_n24261_), .A2(\a[20] ), .Z(new_n24262_));
  NOR2_X1    g24196(.A1(new_n24257_), .A2(new_n24262_), .ZN(new_n24263_));
  XOR2_X1    g24197(.A1(new_n24196_), .A2(new_n24249_), .Z(new_n24264_));
  INV_X1     g24198(.I(new_n24262_), .ZN(new_n24265_));
  NOR2_X1    g24199(.A1(new_n24264_), .A2(new_n24265_), .ZN(new_n24266_));
  OAI22_X1   g24200(.A1(new_n17787_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19412_), .ZN(new_n24267_));
  NAND2_X1   g24201(.A1(new_n19442_), .A2(new_n4469_), .ZN(new_n24268_));
  AOI21_X1   g24202(.A1(new_n24268_), .A2(new_n24267_), .B(new_n4468_), .ZN(new_n24269_));
  NAND2_X1   g24203(.A1(new_n20939_), .A2(new_n24269_), .ZN(new_n24270_));
  XOR2_X1    g24204(.A1(new_n24270_), .A2(\a[17] ), .Z(new_n24271_));
  OAI21_X1   g24205(.A1(new_n24263_), .A2(new_n24266_), .B(new_n24271_), .ZN(new_n24272_));
  NAND2_X1   g24206(.A1(new_n24264_), .A2(new_n24265_), .ZN(new_n24273_));
  NAND2_X1   g24207(.A1(new_n24257_), .A2(new_n24262_), .ZN(new_n24274_));
  XOR2_X1    g24208(.A1(new_n24270_), .A2(new_n3372_), .Z(new_n24275_));
  NAND3_X1   g24209(.A1(new_n24273_), .A2(new_n24275_), .A3(new_n24274_), .ZN(new_n24276_));
  NAND2_X1   g24210(.A1(new_n24272_), .A2(new_n24276_), .ZN(new_n24277_));
  OAI21_X1   g24211(.A1(new_n24062_), .A2(new_n24061_), .B(new_n24060_), .ZN(new_n24278_));
  NAND3_X1   g24212(.A1(new_n24056_), .A2(new_n24055_), .A3(new_n24047_), .ZN(new_n24279_));
  NAND3_X1   g24213(.A1(new_n24278_), .A2(new_n24279_), .A3(new_n24069_), .ZN(new_n24280_));
  OAI21_X1   g24214(.A1(new_n24063_), .A2(new_n24057_), .B(new_n24076_), .ZN(new_n24281_));
  NAND2_X1   g24215(.A1(new_n24281_), .A2(new_n24280_), .ZN(new_n24282_));
  NOR2_X1    g24216(.A1(new_n24064_), .A2(new_n24069_), .ZN(new_n24283_));
  AOI21_X1   g24217(.A1(new_n24282_), .A2(new_n24070_), .B(new_n24283_), .ZN(new_n24284_));
  NOR2_X1    g24218(.A1(new_n24284_), .A2(new_n24277_), .ZN(new_n24285_));
  AOI21_X1   g24219(.A1(new_n24273_), .A2(new_n24274_), .B(new_n24275_), .ZN(new_n24286_));
  NOR3_X1    g24220(.A1(new_n24266_), .A2(new_n24271_), .A3(new_n24263_), .ZN(new_n24287_));
  NOR2_X1    g24221(.A1(new_n24286_), .A2(new_n24287_), .ZN(new_n24288_));
  AOI22_X1   g24222(.A1(new_n24077_), .A2(new_n24069_), .B1(new_n24280_), .B2(new_n24281_), .ZN(new_n24289_));
  NOR2_X1    g24223(.A1(new_n24289_), .A2(new_n24288_), .ZN(new_n24290_));
  OAI22_X1   g24224(.A1(new_n17784_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n19428_), .ZN(new_n24291_));
  NAND2_X1   g24225(.A1(new_n19466_), .A2(new_n6090_), .ZN(new_n24292_));
  AOI21_X1   g24226(.A1(new_n24292_), .A2(new_n24291_), .B(new_n6082_), .ZN(new_n24293_));
  NAND2_X1   g24227(.A1(new_n21100_), .A2(new_n24293_), .ZN(new_n24294_));
  XOR2_X1    g24228(.A1(new_n24294_), .A2(\a[14] ), .Z(new_n24295_));
  NOR3_X1    g24229(.A1(new_n24285_), .A2(new_n24290_), .A3(new_n24295_), .ZN(new_n24296_));
  INV_X1     g24230(.I(new_n24296_), .ZN(new_n24297_));
  OAI21_X1   g24231(.A1(new_n24285_), .A2(new_n24290_), .B(new_n24295_), .ZN(new_n24298_));
  OAI22_X1   g24232(.A1(new_n19475_), .A2(new_n4719_), .B1(new_n19463_), .B2(new_n4716_), .ZN(new_n24299_));
  NAND2_X1   g24233(.A1(new_n19484_), .A2(new_n4709_), .ZN(new_n24300_));
  AOI21_X1   g24234(.A1(new_n24300_), .A2(new_n24299_), .B(new_n4707_), .ZN(new_n24301_));
  NAND2_X1   g24235(.A1(new_n21171_), .A2(new_n24301_), .ZN(new_n24302_));
  XOR2_X1    g24236(.A1(new_n24302_), .A2(new_n4034_), .Z(new_n24303_));
  AOI21_X1   g24237(.A1(new_n24297_), .A2(new_n24298_), .B(new_n24303_), .ZN(new_n24304_));
  INV_X1     g24238(.I(new_n24298_), .ZN(new_n24305_));
  XOR2_X1    g24239(.A1(new_n24302_), .A2(\a[11] ), .Z(new_n24306_));
  NOR3_X1    g24240(.A1(new_n24306_), .A2(new_n24305_), .A3(new_n24296_), .ZN(new_n24307_));
  NOR2_X1    g24241(.A1(new_n24304_), .A2(new_n24307_), .ZN(new_n24308_));
  OAI21_X1   g24242(.A1(new_n24095_), .A2(new_n24094_), .B(new_n24093_), .ZN(new_n24309_));
  NAND3_X1   g24243(.A1(new_n24087_), .A2(new_n24089_), .A3(new_n24080_), .ZN(new_n24310_));
  NAND3_X1   g24244(.A1(new_n24309_), .A2(new_n24310_), .A3(new_n24102_), .ZN(new_n24311_));
  OAI21_X1   g24245(.A1(new_n24096_), .A2(new_n24090_), .B(new_n24105_), .ZN(new_n24312_));
  AOI22_X1   g24246(.A1(new_n24109_), .A2(new_n24102_), .B1(new_n24312_), .B2(new_n24311_), .ZN(new_n24313_));
  XOR2_X1    g24247(.A1(new_n24313_), .A2(new_n24308_), .Z(new_n24314_));
  OAI22_X1   g24248(.A1(new_n19512_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n19522_), .ZN(new_n24315_));
  NAND2_X1   g24249(.A1(new_n21953_), .A2(new_n6784_), .ZN(new_n24316_));
  AOI21_X1   g24250(.A1(new_n24315_), .A2(new_n24316_), .B(new_n6776_), .ZN(new_n24317_));
  NAND2_X1   g24251(.A1(new_n21963_), .A2(new_n24317_), .ZN(new_n24318_));
  XOR2_X1    g24252(.A1(new_n24318_), .A2(\a[8] ), .Z(new_n24319_));
  INV_X1     g24253(.I(new_n24319_), .ZN(new_n24320_));
  NAND2_X1   g24254(.A1(new_n24314_), .A2(new_n24320_), .ZN(new_n24321_));
  NAND2_X1   g24255(.A1(new_n24313_), .A2(new_n24308_), .ZN(new_n24322_));
  OAI21_X1   g24256(.A1(new_n24296_), .A2(new_n24305_), .B(new_n24306_), .ZN(new_n24323_));
  NAND3_X1   g24257(.A1(new_n24303_), .A2(new_n24297_), .A3(new_n24298_), .ZN(new_n24324_));
  NAND2_X1   g24258(.A1(new_n24323_), .A2(new_n24324_), .ZN(new_n24325_));
  NOR3_X1    g24259(.A1(new_n24096_), .A2(new_n24090_), .A3(new_n24105_), .ZN(new_n24326_));
  AOI21_X1   g24260(.A1(new_n24309_), .A2(new_n24310_), .B(new_n24102_), .ZN(new_n24327_));
  OAI22_X1   g24261(.A1(new_n24103_), .A2(new_n24105_), .B1(new_n24326_), .B2(new_n24327_), .ZN(new_n24328_));
  NAND2_X1   g24262(.A1(new_n24328_), .A2(new_n24325_), .ZN(new_n24329_));
  NAND2_X1   g24263(.A1(new_n24329_), .A2(new_n24322_), .ZN(new_n24330_));
  NAND2_X1   g24264(.A1(new_n24330_), .A2(new_n24319_), .ZN(new_n24331_));
  OAI22_X1   g24265(.A1(new_n22115_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n22051_), .ZN(new_n24332_));
  OAI21_X1   g24266(.A1(new_n6839_), .A2(new_n22149_), .B(new_n24332_), .ZN(new_n24333_));
  NAND4_X1   g24267(.A1(new_n22163_), .A2(new_n65_), .A3(new_n6835_), .A4(new_n24333_), .ZN(new_n24334_));
  OAI21_X1   g24268(.A1(new_n22151_), .A2(new_n23951_), .B(new_n22159_), .ZN(new_n24335_));
  NAND2_X1   g24269(.A1(new_n22160_), .A2(new_n22161_), .ZN(new_n24336_));
  NAND2_X1   g24270(.A1(new_n22117_), .A2(new_n24336_), .ZN(new_n24337_));
  NAND4_X1   g24271(.A1(new_n24335_), .A2(new_n6835_), .A3(new_n24337_), .A4(new_n24333_), .ZN(new_n24338_));
  NAND2_X1   g24272(.A1(new_n24338_), .A2(\a[5] ), .ZN(new_n24339_));
  NAND2_X1   g24273(.A1(new_n24334_), .A2(new_n24339_), .ZN(new_n24340_));
  AOI21_X1   g24274(.A1(new_n24331_), .A2(new_n24321_), .B(new_n24340_), .ZN(new_n24341_));
  NOR2_X1    g24275(.A1(new_n24330_), .A2(new_n24319_), .ZN(new_n24342_));
  NOR2_X1    g24276(.A1(new_n24314_), .A2(new_n24320_), .ZN(new_n24343_));
  XOR2_X1    g24277(.A1(new_n24338_), .A2(\a[5] ), .Z(new_n24344_));
  NOR3_X1    g24278(.A1(new_n24344_), .A2(new_n24343_), .A3(new_n24342_), .ZN(new_n24345_));
  NOR2_X1    g24279(.A1(new_n24345_), .A2(new_n24341_), .ZN(new_n24346_));
  XOR2_X1    g24280(.A1(new_n24189_), .A2(new_n24346_), .Z(new_n24347_));
  NAND2_X1   g24281(.A1(new_n24162_), .A2(new_n24159_), .ZN(new_n24348_));
  AOI21_X1   g24282(.A1(new_n2760_), .A2(new_n2761_), .B(new_n2769_), .ZN(new_n24349_));
  OAI21_X1   g24283(.A1(new_n11697_), .A2(new_n2767_), .B(new_n24349_), .ZN(new_n24350_));
  AOI21_X1   g24284(.A1(new_n11370_), .A2(new_n2770_), .B(new_n24350_), .ZN(new_n24351_));
  NAND2_X1   g24285(.A1(new_n12720_), .A2(new_n24351_), .ZN(new_n24352_));
  NOR2_X1    g24286(.A1(new_n23923_), .A2(new_n11221_), .ZN(new_n24353_));
  XOR2_X1    g24287(.A1(new_n24151_), .A2(\a[29] ), .Z(new_n24354_));
  AOI21_X1   g24288(.A1(new_n11221_), .A2(new_n23923_), .B(new_n24354_), .ZN(new_n24355_));
  NOR2_X1    g24289(.A1(new_n24355_), .A2(new_n24353_), .ZN(new_n24356_));
  INV_X1     g24290(.I(new_n24356_), .ZN(new_n24357_));
  NAND2_X1   g24291(.A1(new_n24357_), .A2(new_n3141_), .ZN(new_n24358_));
  NOR2_X1    g24292(.A1(new_n24357_), .A2(new_n3141_), .ZN(new_n24359_));
  INV_X1     g24293(.I(new_n24359_), .ZN(new_n24360_));
  AOI21_X1   g24294(.A1(new_n24358_), .A2(new_n24360_), .B(new_n24352_), .ZN(new_n24361_));
  XOR2_X1    g24295(.A1(new_n24356_), .A2(new_n3141_), .Z(new_n24362_));
  AOI21_X1   g24296(.A1(new_n12720_), .A2(new_n24351_), .B(new_n24362_), .ZN(new_n24363_));
  NOR2_X1    g24297(.A1(new_n24361_), .A2(new_n24363_), .ZN(new_n24364_));
  NOR2_X1    g24298(.A1(new_n24149_), .A2(new_n24155_), .ZN(new_n24365_));
  NAND2_X1   g24299(.A1(new_n24149_), .A2(new_n24155_), .ZN(new_n24366_));
  AOI21_X1   g24300(.A1(new_n24144_), .A2(new_n24366_), .B(new_n24365_), .ZN(new_n24367_));
  XNOR2_X1   g24301(.A1(new_n24367_), .A2(new_n24364_), .ZN(new_n24368_));
  AOI21_X1   g24302(.A1(new_n24164_), .A2(new_n24348_), .B(new_n24368_), .ZN(new_n24369_));
  NAND2_X1   g24303(.A1(new_n24164_), .A2(new_n24348_), .ZN(new_n24370_));
  NAND2_X1   g24304(.A1(new_n24367_), .A2(new_n24364_), .ZN(new_n24371_));
  INV_X1     g24305(.I(new_n24364_), .ZN(new_n24372_));
  INV_X1     g24306(.I(new_n24367_), .ZN(new_n24373_));
  NAND2_X1   g24307(.A1(new_n24373_), .A2(new_n24372_), .ZN(new_n24374_));
  AOI21_X1   g24308(.A1(new_n24371_), .A2(new_n24374_), .B(new_n24370_), .ZN(new_n24375_));
  NOR2_X1    g24309(.A1(new_n24375_), .A2(new_n24369_), .ZN(new_n24376_));
  AOI21_X1   g24310(.A1(new_n24174_), .A2(new_n22150_), .B(new_n23957_), .ZN(new_n24377_));
  INV_X1     g24311(.I(new_n24377_), .ZN(new_n24378_));
  NAND3_X1   g24312(.A1(new_n23917_), .A2(new_n22152_), .A3(new_n24378_), .ZN(new_n24379_));
  AOI21_X1   g24313(.A1(new_n24167_), .A2(new_n22149_), .B(new_n23948_), .ZN(new_n24380_));
  INV_X1     g24314(.I(new_n24380_), .ZN(new_n24381_));
  NAND3_X1   g24315(.A1(new_n24379_), .A2(new_n24167_), .A3(new_n24381_), .ZN(new_n24382_));
  NOR3_X1    g24316(.A1(new_n23952_), .A2(new_n22151_), .A3(new_n24377_), .ZN(new_n24383_));
  OAI21_X1   g24317(.A1(new_n24383_), .A2(new_n24380_), .B(new_n24174_), .ZN(new_n24384_));
  AOI21_X1   g24318(.A1(new_n24384_), .A2(new_n24382_), .B(new_n24376_), .ZN(new_n24385_));
  INV_X1     g24319(.I(new_n24376_), .ZN(new_n24386_));
  OAI21_X1   g24320(.A1(new_n24383_), .A2(new_n24380_), .B(new_n24167_), .ZN(new_n24387_));
  NAND3_X1   g24321(.A1(new_n24379_), .A2(new_n24174_), .A3(new_n24381_), .ZN(new_n24388_));
  AOI21_X1   g24322(.A1(new_n24387_), .A2(new_n24388_), .B(new_n24386_), .ZN(new_n24389_));
  NOR2_X1    g24323(.A1(new_n24385_), .A2(new_n24389_), .ZN(new_n24390_));
  INV_X1     g24324(.I(new_n24390_), .ZN(new_n24391_));
  AOI22_X1   g24325(.A1(new_n24174_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n23957_), .ZN(new_n24392_));
  NOR2_X1    g24326(.A1(new_n24376_), .A2(new_n9489_), .ZN(new_n24393_));
  OAI21_X1   g24327(.A1(new_n24393_), .A2(new_n24392_), .B(new_n6922_), .ZN(new_n24394_));
  NOR2_X1    g24328(.A1(new_n24391_), .A2(new_n24394_), .ZN(new_n24395_));
  XOR2_X1    g24329(.A1(new_n24395_), .A2(\a[2] ), .Z(new_n24396_));
  INV_X1     g24330(.I(new_n24140_), .ZN(new_n24397_));
  AOI21_X1   g24331(.A1(new_n24397_), .A2(new_n24178_), .B(new_n24180_), .ZN(new_n24398_));
  XOR2_X1    g24332(.A1(new_n24398_), .A2(new_n24396_), .Z(new_n24399_));
  XNOR2_X1   g24333(.A1(new_n24399_), .A2(new_n24347_), .ZN(new_n24400_));
  INV_X1     g24334(.I(new_n24400_), .ZN(new_n24401_));
  XOR2_X1    g24335(.A1(new_n24183_), .A2(new_n24401_), .Z(\result[3] ));
  NOR2_X1    g24336(.A1(new_n24234_), .A2(new_n24239_), .ZN(new_n24403_));
  AOI21_X1   g24337(.A1(new_n24201_), .A2(new_n24212_), .B(new_n24213_), .ZN(new_n24404_));
  AOI21_X1   g24338(.A1(new_n19350_), .A2(new_n3189_), .B(new_n2764_), .ZN(new_n24405_));
  OAI21_X1   g24339(.A1(new_n19343_), .A2(new_n2771_), .B(new_n24405_), .ZN(new_n24406_));
  AOI21_X1   g24340(.A1(new_n3332_), .A2(new_n17807_), .B(new_n24406_), .ZN(new_n24407_));
  NOR2_X1    g24341(.A1(new_n2598_), .A2(new_n1995_), .ZN(new_n24408_));
  NAND2_X1   g24342(.A1(new_n599_), .A2(new_n271_), .ZN(new_n24409_));
  NOR4_X1    g24343(.A1(new_n988_), .A2(new_n369_), .A3(new_n656_), .A4(new_n24409_), .ZN(new_n24410_));
  NAND4_X1   g24344(.A1(new_n24410_), .A2(new_n646_), .A3(new_n24408_), .A4(new_n852_), .ZN(new_n24411_));
  NAND4_X1   g24345(.A1(new_n2339_), .A2(new_n454_), .A3(new_n725_), .A4(new_n2012_), .ZN(new_n24412_));
  NOR4_X1    g24346(.A1(new_n398_), .A2(new_n388_), .A3(new_n376_), .A4(new_n468_), .ZN(new_n24413_));
  NOR4_X1    g24347(.A1(new_n482_), .A2(new_n475_), .A3(new_n560_), .A4(new_n163_), .ZN(new_n24414_));
  OR3_X2     g24348(.A1(new_n24412_), .A2(new_n24413_), .A3(new_n24414_), .Z(new_n24415_));
  NAND4_X1   g24349(.A1(new_n385_), .A2(new_n690_), .A3(new_n842_), .A4(new_n1647_), .ZN(new_n24416_));
  NAND4_X1   g24350(.A1(new_n1207_), .A2(new_n416_), .A3(new_n1310_), .A4(new_n24416_), .ZN(new_n24417_));
  NOR4_X1    g24351(.A1(new_n24415_), .A2(new_n2182_), .A3(new_n24411_), .A4(new_n24417_), .ZN(new_n24418_));
  NAND3_X1   g24352(.A1(new_n3446_), .A2(new_n3017_), .A3(new_n24418_), .ZN(new_n24419_));
  INV_X1     g24353(.I(new_n24419_), .ZN(new_n24420_));
  AOI21_X1   g24354(.A1(new_n19915_), .A2(new_n24407_), .B(new_n24420_), .ZN(new_n24421_));
  NAND3_X1   g24355(.A1(new_n19915_), .A2(new_n24407_), .A3(new_n24420_), .ZN(new_n24422_));
  INV_X1     g24356(.I(new_n24422_), .ZN(new_n24423_));
  NOR2_X1    g24357(.A1(new_n24423_), .A2(new_n24421_), .ZN(new_n24424_));
  NAND2_X1   g24358(.A1(new_n24424_), .A2(new_n24404_), .ZN(new_n24425_));
  INV_X1     g24359(.I(new_n24404_), .ZN(new_n24426_));
  INV_X1     g24360(.I(new_n24421_), .ZN(new_n24427_));
  NAND2_X1   g24361(.A1(new_n24427_), .A2(new_n24422_), .ZN(new_n24428_));
  NAND2_X1   g24362(.A1(new_n24426_), .A2(new_n24428_), .ZN(new_n24429_));
  NAND2_X1   g24363(.A1(new_n24429_), .A2(new_n24425_), .ZN(new_n24430_));
  OAI22_X1   g24364(.A1(new_n19356_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n19364_), .ZN(new_n24431_));
  NAND2_X1   g24365(.A1(new_n17802_), .A2(new_n2750_), .ZN(new_n24432_));
  AOI21_X1   g24366(.A1(new_n24431_), .A2(new_n24432_), .B(new_n2737_), .ZN(new_n24433_));
  NAND2_X1   g24367(.A1(new_n19951_), .A2(new_n24433_), .ZN(new_n24434_));
  NOR2_X1    g24368(.A1(new_n24434_), .A2(\a[29] ), .ZN(new_n24435_));
  INV_X1     g24369(.I(new_n24435_), .ZN(new_n24436_));
  NAND2_X1   g24370(.A1(new_n24434_), .A2(\a[29] ), .ZN(new_n24437_));
  AOI21_X1   g24371(.A1(new_n24436_), .A2(new_n24437_), .B(new_n24430_), .ZN(new_n24438_));
  XOR2_X1    g24372(.A1(new_n24424_), .A2(new_n24404_), .Z(new_n24439_));
  INV_X1     g24373(.I(new_n24437_), .ZN(new_n24440_));
  NOR3_X1    g24374(.A1(new_n24439_), .A2(new_n24440_), .A3(new_n24435_), .ZN(new_n24441_));
  NOR4_X1    g24375(.A1(new_n24438_), .A2(new_n24441_), .A3(new_n24199_), .A4(new_n24218_), .ZN(new_n24442_));
  OAI22_X1   g24376(.A1(new_n24438_), .A2(new_n24441_), .B1(new_n24199_), .B2(new_n24218_), .ZN(new_n24443_));
  INV_X1     g24377(.I(new_n24443_), .ZN(new_n24444_));
  NAND2_X1   g24378(.A1(new_n24197_), .A2(new_n24008_), .ZN(new_n24445_));
  NAND2_X1   g24379(.A1(new_n24445_), .A2(new_n24009_), .ZN(new_n24446_));
  NOR2_X1    g24380(.A1(new_n24446_), .A2(new_n24218_), .ZN(new_n24447_));
  NOR2_X1    g24381(.A1(new_n24199_), .A2(new_n24230_), .ZN(new_n24448_));
  OAI21_X1   g24382(.A1(new_n24447_), .A2(new_n24448_), .B(new_n24227_), .ZN(new_n24449_));
  NOR3_X1    g24383(.A1(new_n24449_), .A2(new_n24444_), .A3(new_n24442_), .ZN(new_n24450_));
  OAI21_X1   g24384(.A1(new_n24435_), .A2(new_n24440_), .B(new_n24439_), .ZN(new_n24451_));
  NAND3_X1   g24385(.A1(new_n24430_), .A2(new_n24436_), .A3(new_n24437_), .ZN(new_n24452_));
  NOR2_X1    g24386(.A1(new_n24199_), .A2(new_n24218_), .ZN(new_n24453_));
  NAND3_X1   g24387(.A1(new_n24453_), .A2(new_n24451_), .A3(new_n24452_), .ZN(new_n24454_));
  XOR2_X1    g24388(.A1(new_n24199_), .A2(new_n24218_), .Z(new_n24455_));
  AOI22_X1   g24389(.A1(new_n24455_), .A2(new_n24227_), .B1(new_n24454_), .B2(new_n24443_), .ZN(new_n24456_));
  OAI22_X1   g24390(.A1(new_n19375_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n17797_), .ZN(new_n24457_));
  NAND2_X1   g24391(.A1(new_n19386_), .A2(new_n3317_), .ZN(new_n24458_));
  AOI21_X1   g24392(.A1(new_n24458_), .A2(new_n24457_), .B(new_n3260_), .ZN(new_n24459_));
  NAND2_X1   g24393(.A1(new_n20162_), .A2(new_n24459_), .ZN(new_n24460_));
  XOR2_X1    g24394(.A1(new_n24460_), .A2(\a[26] ), .Z(new_n24461_));
  NOR3_X1    g24395(.A1(new_n24450_), .A2(new_n24456_), .A3(new_n24461_), .ZN(new_n24462_));
  NAND4_X1   g24396(.A1(new_n24455_), .A2(new_n24443_), .A3(new_n24454_), .A4(new_n24227_), .ZN(new_n24463_));
  OAI21_X1   g24397(.A1(new_n24442_), .A2(new_n24444_), .B(new_n24449_), .ZN(new_n24464_));
  INV_X1     g24398(.I(new_n24461_), .ZN(new_n24465_));
  AOI21_X1   g24399(.A1(new_n24464_), .A2(new_n24463_), .B(new_n24465_), .ZN(new_n24466_));
  NOR3_X1    g24400(.A1(new_n24466_), .A2(new_n24462_), .A3(new_n24403_), .ZN(new_n24467_));
  INV_X1     g24401(.I(new_n24403_), .ZN(new_n24468_));
  NAND3_X1   g24402(.A1(new_n24464_), .A2(new_n24463_), .A3(new_n24465_), .ZN(new_n24469_));
  OAI21_X1   g24403(.A1(new_n24450_), .A2(new_n24456_), .B(new_n24461_), .ZN(new_n24470_));
  AOI21_X1   g24404(.A1(new_n24469_), .A2(new_n24470_), .B(new_n24468_), .ZN(new_n24471_));
  OAI22_X1   g24405(.A1(new_n19393_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n17793_), .ZN(new_n24472_));
  NAND2_X1   g24406(.A1(new_n19399_), .A2(new_n3312_), .ZN(new_n24473_));
  AOI21_X1   g24407(.A1(new_n24473_), .A2(new_n24472_), .B(new_n3302_), .ZN(new_n24474_));
  NAND2_X1   g24408(.A1(new_n20264_), .A2(new_n24474_), .ZN(new_n24475_));
  XOR2_X1    g24409(.A1(new_n24475_), .A2(\a[23] ), .Z(new_n24476_));
  INV_X1     g24410(.I(new_n24476_), .ZN(new_n24477_));
  NOR3_X1    g24411(.A1(new_n24471_), .A2(new_n24467_), .A3(new_n24477_), .ZN(new_n24478_));
  NAND3_X1   g24412(.A1(new_n24469_), .A2(new_n24470_), .A3(new_n24468_), .ZN(new_n24479_));
  OAI21_X1   g24413(.A1(new_n24466_), .A2(new_n24462_), .B(new_n24403_), .ZN(new_n24480_));
  AOI21_X1   g24414(.A1(new_n24480_), .A2(new_n24479_), .B(new_n24476_), .ZN(new_n24481_));
  NOR2_X1    g24415(.A1(new_n24478_), .A2(new_n24481_), .ZN(new_n24482_));
  AOI21_X1   g24416(.A1(new_n24196_), .A2(new_n24255_), .B(new_n24246_), .ZN(new_n24483_));
  NAND2_X1   g24417(.A1(new_n24483_), .A2(new_n24482_), .ZN(new_n24484_));
  NAND3_X1   g24418(.A1(new_n24480_), .A2(new_n24479_), .A3(new_n24476_), .ZN(new_n24485_));
  OAI21_X1   g24419(.A1(new_n24471_), .A2(new_n24467_), .B(new_n24477_), .ZN(new_n24486_));
  NAND2_X1   g24420(.A1(new_n24486_), .A2(new_n24485_), .ZN(new_n24487_));
  OAI21_X1   g24421(.A1(new_n24254_), .A2(new_n24249_), .B(new_n24247_), .ZN(new_n24488_));
  NAND2_X1   g24422(.A1(new_n24488_), .A2(new_n24487_), .ZN(new_n24489_));
  OAI22_X1   g24423(.A1(new_n19410_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n17789_), .ZN(new_n24490_));
  NAND2_X1   g24424(.A1(new_n19415_), .A2(new_n4096_), .ZN(new_n24491_));
  AOI21_X1   g24425(.A1(new_n24491_), .A2(new_n24490_), .B(new_n4095_), .ZN(new_n24492_));
  NAND2_X1   g24426(.A1(new_n20846_), .A2(new_n24492_), .ZN(new_n24493_));
  XOR2_X1    g24427(.A1(new_n24493_), .A2(\a[20] ), .Z(new_n24494_));
  INV_X1     g24428(.I(new_n24494_), .ZN(new_n24495_));
  NAND3_X1   g24429(.A1(new_n24489_), .A2(new_n24484_), .A3(new_n24495_), .ZN(new_n24496_));
  NOR2_X1    g24430(.A1(new_n24488_), .A2(new_n24487_), .ZN(new_n24497_));
  NOR2_X1    g24431(.A1(new_n24483_), .A2(new_n24482_), .ZN(new_n24498_));
  OAI21_X1   g24432(.A1(new_n24497_), .A2(new_n24498_), .B(new_n24494_), .ZN(new_n24499_));
  NOR2_X1    g24433(.A1(new_n24257_), .A2(new_n24262_), .ZN(new_n24500_));
  NAND3_X1   g24434(.A1(new_n24499_), .A2(new_n24496_), .A3(new_n24500_), .ZN(new_n24501_));
  NOR3_X1    g24435(.A1(new_n24497_), .A2(new_n24498_), .A3(new_n24494_), .ZN(new_n24502_));
  AOI21_X1   g24436(.A1(new_n24489_), .A2(new_n24484_), .B(new_n24495_), .ZN(new_n24503_));
  NAND2_X1   g24437(.A1(new_n24264_), .A2(new_n24265_), .ZN(new_n24504_));
  OAI21_X1   g24438(.A1(new_n24502_), .A2(new_n24503_), .B(new_n24504_), .ZN(new_n24505_));
  OAI22_X1   g24439(.A1(new_n19423_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n17787_), .ZN(new_n24506_));
  NAND2_X1   g24440(.A1(new_n20896_), .A2(new_n4469_), .ZN(new_n24507_));
  AOI21_X1   g24441(.A1(new_n24507_), .A2(new_n24506_), .B(new_n4468_), .ZN(new_n24508_));
  NAND2_X1   g24442(.A1(new_n22226_), .A2(new_n24508_), .ZN(new_n24509_));
  XOR2_X1    g24443(.A1(new_n24509_), .A2(\a[17] ), .Z(new_n24510_));
  NAND3_X1   g24444(.A1(new_n24505_), .A2(new_n24501_), .A3(new_n24510_), .ZN(new_n24511_));
  NOR3_X1    g24445(.A1(new_n24502_), .A2(new_n24503_), .A3(new_n24504_), .ZN(new_n24512_));
  AOI21_X1   g24446(.A1(new_n24499_), .A2(new_n24496_), .B(new_n24500_), .ZN(new_n24513_));
  XOR2_X1    g24447(.A1(new_n24509_), .A2(new_n3372_), .Z(new_n24514_));
  OAI21_X1   g24448(.A1(new_n24512_), .A2(new_n24513_), .B(new_n24514_), .ZN(new_n24515_));
  NAND2_X1   g24449(.A1(new_n24515_), .A2(new_n24511_), .ZN(new_n24516_));
  OAI21_X1   g24450(.A1(new_n24289_), .A2(new_n24277_), .B(new_n24272_), .ZN(new_n24517_));
  NOR2_X1    g24451(.A1(new_n24517_), .A2(new_n24516_), .ZN(new_n24518_));
  NOR3_X1    g24452(.A1(new_n24512_), .A2(new_n24513_), .A3(new_n24514_), .ZN(new_n24519_));
  AOI21_X1   g24453(.A1(new_n24505_), .A2(new_n24501_), .B(new_n24510_), .ZN(new_n24520_));
  NOR2_X1    g24454(.A1(new_n24519_), .A2(new_n24520_), .ZN(new_n24521_));
  AOI21_X1   g24455(.A1(new_n24284_), .A2(new_n24288_), .B(new_n24286_), .ZN(new_n24522_));
  NOR2_X1    g24456(.A1(new_n24522_), .A2(new_n24521_), .ZN(new_n24523_));
  OAI22_X1   g24457(.A1(new_n19437_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n17784_), .ZN(new_n24524_));
  NAND2_X1   g24458(.A1(new_n19472_), .A2(new_n6090_), .ZN(new_n24525_));
  AOI21_X1   g24459(.A1(new_n24525_), .A2(new_n24524_), .B(new_n6082_), .ZN(new_n24526_));
  NAND2_X1   g24460(.A1(new_n21117_), .A2(new_n24526_), .ZN(new_n24527_));
  XOR2_X1    g24461(.A1(new_n24527_), .A2(\a[14] ), .Z(new_n24528_));
  NOR3_X1    g24462(.A1(new_n24523_), .A2(new_n24518_), .A3(new_n24528_), .ZN(new_n24529_));
  INV_X1     g24463(.I(new_n24283_), .ZN(new_n24530_));
  NAND2_X1   g24464(.A1(new_n24282_), .A2(new_n24070_), .ZN(new_n24531_));
  NAND3_X1   g24465(.A1(new_n24531_), .A2(new_n24288_), .A3(new_n24530_), .ZN(new_n24532_));
  NAND3_X1   g24466(.A1(new_n24532_), .A2(new_n24272_), .A3(new_n24521_), .ZN(new_n24533_));
  NAND2_X1   g24467(.A1(new_n24517_), .A2(new_n24516_), .ZN(new_n24534_));
  INV_X1     g24468(.I(new_n24528_), .ZN(new_n24535_));
  AOI21_X1   g24469(.A1(new_n24533_), .A2(new_n24534_), .B(new_n24535_), .ZN(new_n24536_));
  NOR3_X1    g24470(.A1(new_n24285_), .A2(new_n24290_), .A3(new_n24295_), .ZN(new_n24537_));
  INV_X1     g24471(.I(new_n24537_), .ZN(new_n24538_));
  NOR3_X1    g24472(.A1(new_n24529_), .A2(new_n24536_), .A3(new_n24538_), .ZN(new_n24539_));
  NAND3_X1   g24473(.A1(new_n24533_), .A2(new_n24534_), .A3(new_n24535_), .ZN(new_n24540_));
  OAI21_X1   g24474(.A1(new_n24523_), .A2(new_n24518_), .B(new_n24528_), .ZN(new_n24541_));
  AOI21_X1   g24475(.A1(new_n24541_), .A2(new_n24540_), .B(new_n24537_), .ZN(new_n24542_));
  NOR2_X1    g24476(.A1(new_n19508_), .A2(new_n21151_), .ZN(new_n24543_));
  NOR2_X1    g24477(.A1(new_n21153_), .A2(new_n21152_), .ZN(new_n24544_));
  NOR2_X1    g24478(.A1(new_n21956_), .A2(new_n24544_), .ZN(new_n24545_));
  OAI22_X1   g24479(.A1(new_n17775_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n19475_), .ZN(new_n24546_));
  NAND2_X1   g24480(.A1(new_n21157_), .A2(new_n4709_), .ZN(new_n24547_));
  AOI21_X1   g24481(.A1(new_n24547_), .A2(new_n24546_), .B(new_n4707_), .ZN(new_n24548_));
  OAI21_X1   g24482(.A1(new_n24545_), .A2(new_n24543_), .B(new_n24548_), .ZN(new_n24549_));
  XOR2_X1    g24483(.A1(new_n24549_), .A2(new_n4034_), .Z(new_n24550_));
  NOR3_X1    g24484(.A1(new_n24539_), .A2(new_n24542_), .A3(new_n24550_), .ZN(new_n24551_));
  NAND3_X1   g24485(.A1(new_n24541_), .A2(new_n24540_), .A3(new_n24537_), .ZN(new_n24552_));
  OAI21_X1   g24486(.A1(new_n24529_), .A2(new_n24536_), .B(new_n24538_), .ZN(new_n24553_));
  XOR2_X1    g24487(.A1(new_n24549_), .A2(\a[11] ), .Z(new_n24554_));
  AOI21_X1   g24488(.A1(new_n24553_), .A2(new_n24552_), .B(new_n24554_), .ZN(new_n24555_));
  NOR2_X1    g24489(.A1(new_n24551_), .A2(new_n24555_), .ZN(new_n24556_));
  AOI21_X1   g24490(.A1(new_n24328_), .A2(new_n24308_), .B(new_n24304_), .ZN(new_n24557_));
  NAND2_X1   g24491(.A1(new_n24557_), .A2(new_n24556_), .ZN(new_n24558_));
  NAND3_X1   g24492(.A1(new_n24553_), .A2(new_n24552_), .A3(new_n24554_), .ZN(new_n24559_));
  OAI21_X1   g24493(.A1(new_n24539_), .A2(new_n24542_), .B(new_n24550_), .ZN(new_n24560_));
  NAND2_X1   g24494(.A1(new_n24560_), .A2(new_n24559_), .ZN(new_n24561_));
  OAI21_X1   g24495(.A1(new_n24313_), .A2(new_n24325_), .B(new_n24323_), .ZN(new_n24562_));
  NAND2_X1   g24496(.A1(new_n24562_), .A2(new_n24561_), .ZN(new_n24563_));
  OAI22_X1   g24497(.A1(new_n19512_), .A2(new_n6783_), .B1(new_n21960_), .B2(new_n6788_), .ZN(new_n24564_));
  NAND2_X1   g24498(.A1(new_n22048_), .A2(new_n6784_), .ZN(new_n24565_));
  AOI21_X1   g24499(.A1(new_n24565_), .A2(new_n24564_), .B(new_n6776_), .ZN(new_n24566_));
  NAND2_X1   g24500(.A1(new_n22175_), .A2(new_n24566_), .ZN(new_n24567_));
  XOR2_X1    g24501(.A1(new_n24567_), .A2(new_n4009_), .Z(new_n24568_));
  NAND3_X1   g24502(.A1(new_n24558_), .A2(new_n24568_), .A3(new_n24563_), .ZN(new_n24569_));
  NOR2_X1    g24503(.A1(new_n24562_), .A2(new_n24561_), .ZN(new_n24570_));
  NOR2_X1    g24504(.A1(new_n24557_), .A2(new_n24556_), .ZN(new_n24571_));
  XOR2_X1    g24505(.A1(new_n24567_), .A2(\a[8] ), .Z(new_n24572_));
  OAI21_X1   g24506(.A1(new_n24571_), .A2(new_n24570_), .B(new_n24572_), .ZN(new_n24573_));
  NOR2_X1    g24507(.A1(new_n24330_), .A2(new_n24319_), .ZN(new_n24574_));
  NAND3_X1   g24508(.A1(new_n24573_), .A2(new_n24569_), .A3(new_n24574_), .ZN(new_n24575_));
  NOR3_X1    g24509(.A1(new_n24571_), .A2(new_n24570_), .A3(new_n24572_), .ZN(new_n24576_));
  AOI21_X1   g24510(.A1(new_n24558_), .A2(new_n24563_), .B(new_n24568_), .ZN(new_n24577_));
  NAND2_X1   g24511(.A1(new_n24314_), .A2(new_n24320_), .ZN(new_n24578_));
  OAI21_X1   g24512(.A1(new_n24576_), .A2(new_n24577_), .B(new_n24578_), .ZN(new_n24579_));
  OAI22_X1   g24513(.A1(new_n22115_), .A2(new_n6913_), .B1(new_n6843_), .B2(new_n22149_), .ZN(new_n24580_));
  NAND2_X1   g24514(.A1(new_n23957_), .A2(new_n6838_), .ZN(new_n24581_));
  AOI21_X1   g24515(.A1(new_n24580_), .A2(new_n24581_), .B(new_n6836_), .ZN(new_n24582_));
  OAI21_X1   g24516(.A1(new_n23954_), .A2(new_n23950_), .B(new_n24582_), .ZN(new_n24583_));
  XOR2_X1    g24517(.A1(new_n24583_), .A2(\a[5] ), .Z(new_n24584_));
  NAND3_X1   g24518(.A1(new_n24579_), .A2(new_n24575_), .A3(new_n24584_), .ZN(new_n24585_));
  NOR3_X1    g24519(.A1(new_n24576_), .A2(new_n24577_), .A3(new_n24578_), .ZN(new_n24586_));
  AOI21_X1   g24520(.A1(new_n24573_), .A2(new_n24569_), .B(new_n24574_), .ZN(new_n24587_));
  XOR2_X1    g24521(.A1(new_n24583_), .A2(new_n65_), .Z(new_n24588_));
  OAI21_X1   g24522(.A1(new_n24586_), .A2(new_n24587_), .B(new_n24588_), .ZN(new_n24589_));
  NAND2_X1   g24523(.A1(new_n24589_), .A2(new_n24585_), .ZN(new_n24590_));
  INV_X1     g24524(.I(new_n23905_), .ZN(new_n24591_));
  NOR3_X1    g24525(.A1(new_n23915_), .A2(new_n23910_), .A3(new_n24591_), .ZN(new_n24592_));
  NOR3_X1    g24526(.A1(new_n24123_), .A2(new_n24130_), .A3(new_n24135_), .ZN(new_n24593_));
  AOI21_X1   g24527(.A1(new_n24185_), .A2(new_n24186_), .B(new_n24184_), .ZN(new_n24594_));
  OAI22_X1   g24528(.A1(new_n24592_), .A2(new_n24135_), .B1(new_n24593_), .B2(new_n24594_), .ZN(new_n24595_));
  AOI21_X1   g24529(.A1(new_n24595_), .A2(new_n24346_), .B(new_n24341_), .ZN(new_n24596_));
  XOR2_X1    g24530(.A1(new_n24596_), .A2(new_n24590_), .Z(new_n24597_));
  NOR3_X1    g24531(.A1(new_n24383_), .A2(new_n24167_), .A3(new_n24380_), .ZN(new_n24598_));
  OAI21_X1   g24532(.A1(new_n24386_), .A2(new_n24598_), .B(new_n24387_), .ZN(new_n24599_));
  INV_X1     g24533(.I(new_n3141_), .ZN(new_n24600_));
  NAND2_X1   g24534(.A1(new_n2772_), .A2(new_n2767_), .ZN(new_n24601_));
  AOI22_X1   g24535(.A1(new_n11694_), .A2(new_n2770_), .B1(new_n11226_), .B2(new_n24601_), .ZN(new_n24602_));
  OAI21_X1   g24536(.A1(new_n13970_), .A2(new_n2764_), .B(new_n24602_), .ZN(new_n24603_));
  XOR2_X1    g24537(.A1(new_n24603_), .A2(new_n24600_), .Z(new_n24604_));
  OAI21_X1   g24538(.A1(new_n24352_), .A2(new_n24359_), .B(new_n24358_), .ZN(new_n24605_));
  XNOR2_X1   g24539(.A1(new_n24605_), .A2(new_n24604_), .ZN(new_n24606_));
  NAND2_X1   g24540(.A1(new_n24370_), .A2(new_n24372_), .ZN(new_n24607_));
  XOR2_X1    g24541(.A1(new_n24607_), .A2(new_n24606_), .Z(new_n24608_));
  XOR2_X1    g24542(.A1(new_n24370_), .A2(new_n24372_), .Z(new_n24609_));
  NAND2_X1   g24543(.A1(new_n24609_), .A2(new_n24373_), .ZN(new_n24610_));
  NOR2_X1    g24544(.A1(new_n24610_), .A2(new_n24608_), .ZN(new_n24611_));
  AND2_X2    g24545(.A1(new_n24610_), .A2(new_n24608_), .Z(new_n24612_));
  NOR2_X1    g24546(.A1(new_n24612_), .A2(new_n24611_), .ZN(new_n24613_));
  XOR2_X1    g24547(.A1(new_n24613_), .A2(new_n24386_), .Z(new_n24614_));
  INV_X1     g24548(.I(new_n24614_), .ZN(new_n24615_));
  NAND2_X1   g24549(.A1(new_n24599_), .A2(new_n24615_), .ZN(new_n24616_));
  XOR2_X1    g24550(.A1(new_n24613_), .A2(new_n24376_), .Z(new_n24617_));
  OAI21_X1   g24551(.A1(new_n24599_), .A2(new_n24617_), .B(new_n24616_), .ZN(new_n24618_));
  OAI22_X1   g24552(.A1(new_n24376_), .A2(new_n9483_), .B1(new_n9485_), .B2(new_n24167_), .ZN(new_n24619_));
  INV_X1     g24553(.I(new_n24613_), .ZN(new_n24620_));
  NAND2_X1   g24554(.A1(new_n24620_), .A2(new_n9488_), .ZN(new_n24621_));
  AOI21_X1   g24555(.A1(new_n24621_), .A2(new_n24619_), .B(new_n9482_), .ZN(new_n24622_));
  NAND2_X1   g24556(.A1(new_n24618_), .A2(new_n24622_), .ZN(new_n24623_));
  XOR2_X1    g24557(.A1(new_n24623_), .A2(\a[2] ), .Z(new_n24624_));
  INV_X1     g24558(.I(new_n24624_), .ZN(new_n24625_));
  XOR2_X1    g24559(.A1(new_n24597_), .A2(new_n24625_), .Z(new_n24626_));
  INV_X1     g24560(.I(new_n24626_), .ZN(new_n24627_));
  NOR4_X1    g24561(.A1(new_n23964_), .A2(new_n24181_), .A3(new_n24400_), .A4(new_n24627_), .ZN(new_n24628_));
  INV_X1     g24562(.I(new_n24628_), .ZN(new_n24629_));
  OAI21_X1   g24563(.A1(new_n23694_), .A2(new_n23693_), .B(new_n21989_), .ZN(new_n24630_));
  NAND3_X1   g24564(.A1(new_n23686_), .A2(new_n23691_), .A3(new_n21990_), .ZN(new_n24631_));
  NAND2_X1   g24565(.A1(new_n24630_), .A2(new_n24631_), .ZN(new_n24632_));
  NAND3_X1   g24566(.A1(new_n24632_), .A2(new_n23712_), .A3(new_n23708_), .ZN(new_n24633_));
  INV_X1     g24567(.I(new_n24181_), .ZN(new_n24634_));
  NAND4_X1   g24568(.A1(new_n24633_), .A2(new_n23963_), .A3(new_n24634_), .A4(new_n24401_), .ZN(new_n24635_));
  NAND2_X1   g24569(.A1(new_n24635_), .A2(new_n24627_), .ZN(new_n24636_));
  NAND2_X1   g24570(.A1(new_n24629_), .A2(new_n24636_), .ZN(\result[4] ));
  NAND3_X1   g24571(.A1(new_n24451_), .A2(new_n24452_), .A3(new_n24227_), .ZN(new_n24638_));
  NAND3_X1   g24572(.A1(new_n24638_), .A2(new_n24446_), .A3(new_n24230_), .ZN(new_n24639_));
  NAND3_X1   g24573(.A1(new_n24439_), .A2(new_n24436_), .A3(new_n24437_), .ZN(new_n24640_));
  AOI21_X1   g24574(.A1(new_n19350_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n24641_));
  OAI21_X1   g24575(.A1(new_n2767_), .A2(new_n17806_), .B(new_n24641_), .ZN(new_n24642_));
  AOI21_X1   g24576(.A1(new_n19359_), .A2(new_n3332_), .B(new_n24642_), .ZN(new_n24643_));
  NOR4_X1    g24577(.A1(new_n402_), .A2(new_n523_), .A3(new_n1154_), .A4(new_n2323_), .ZN(new_n24644_));
  NOR4_X1    g24578(.A1(new_n217_), .A2(new_n591_), .A3(new_n119_), .A4(new_n782_), .ZN(new_n24645_));
  NOR3_X1    g24579(.A1(new_n774_), .A2(new_n752_), .A3(new_n488_), .ZN(new_n24646_));
  INV_X1     g24580(.I(new_n24646_), .ZN(new_n24647_));
  NAND2_X1   g24581(.A1(new_n1212_), .A2(new_n221_), .ZN(new_n24648_));
  NOR4_X1    g24582(.A1(new_n24647_), .A2(new_n2445_), .A3(new_n24645_), .A4(new_n24648_), .ZN(new_n24649_));
  NAND4_X1   g24583(.A1(new_n24644_), .A2(new_n2827_), .A3(new_n2872_), .A4(new_n24649_), .ZN(new_n24650_));
  NOR3_X1    g24584(.A1(new_n24650_), .A2(new_n3974_), .A3(new_n12923_), .ZN(new_n24651_));
  AOI21_X1   g24585(.A1(new_n20096_), .A2(new_n24643_), .B(new_n24651_), .ZN(new_n24652_));
  NAND3_X1   g24586(.A1(new_n20096_), .A2(new_n24643_), .A3(new_n24651_), .ZN(new_n24653_));
  INV_X1     g24587(.I(new_n24653_), .ZN(new_n24654_));
  NOR2_X1    g24588(.A1(new_n24654_), .A2(new_n24652_), .ZN(new_n24655_));
  INV_X1     g24589(.I(new_n24652_), .ZN(new_n24656_));
  AOI21_X1   g24590(.A1(new_n24656_), .A2(new_n24653_), .B(new_n24421_), .ZN(new_n24657_));
  AOI21_X1   g24591(.A1(new_n24404_), .A2(new_n24422_), .B(new_n24421_), .ZN(new_n24658_));
  INV_X1     g24592(.I(new_n24658_), .ZN(new_n24659_));
  AOI22_X1   g24593(.A1(new_n24659_), .A2(new_n24655_), .B1(new_n24425_), .B2(new_n24657_), .ZN(new_n24660_));
  OAI22_X1   g24594(.A1(new_n17801_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19364_), .ZN(new_n24661_));
  OAI21_X1   g24595(.A1(new_n17797_), .A2(new_n3175_), .B(new_n24661_), .ZN(new_n24662_));
  NAND4_X1   g24596(.A1(new_n20176_), .A2(new_n20179_), .A3(new_n2736_), .A4(new_n24662_), .ZN(new_n24663_));
  XOR2_X1    g24597(.A1(new_n24663_), .A2(\a[29] ), .Z(new_n24664_));
  XOR2_X1    g24598(.A1(new_n24664_), .A2(new_n24660_), .Z(new_n24665_));
  NAND3_X1   g24599(.A1(new_n24639_), .A2(new_n24665_), .A3(new_n24640_), .ZN(new_n24666_));
  NOR3_X1    g24600(.A1(new_n24438_), .A2(new_n24441_), .A3(new_n24226_), .ZN(new_n24667_));
  NOR3_X1    g24601(.A1(new_n24667_), .A2(new_n24199_), .A3(new_n24218_), .ZN(new_n24668_));
  INV_X1     g24602(.I(new_n24640_), .ZN(new_n24669_));
  XOR2_X1    g24603(.A1(new_n24663_), .A2(new_n74_), .Z(new_n24670_));
  XOR2_X1    g24604(.A1(new_n24670_), .A2(new_n24660_), .Z(new_n24671_));
  OAI21_X1   g24605(.A1(new_n24668_), .A2(new_n24669_), .B(new_n24671_), .ZN(new_n24672_));
  OAI22_X1   g24606(.A1(new_n19385_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19375_), .ZN(new_n24673_));
  NAND2_X1   g24607(.A1(new_n17794_), .A2(new_n3317_), .ZN(new_n24674_));
  AOI21_X1   g24608(.A1(new_n24673_), .A2(new_n24674_), .B(new_n3260_), .ZN(new_n24675_));
  NAND2_X1   g24609(.A1(new_n20134_), .A2(new_n24675_), .ZN(new_n24676_));
  XOR2_X1    g24610(.A1(new_n24676_), .A2(new_n72_), .Z(new_n24677_));
  NAND3_X1   g24611(.A1(new_n24672_), .A2(new_n24666_), .A3(new_n24677_), .ZN(new_n24678_));
  NOR3_X1    g24612(.A1(new_n24668_), .A2(new_n24671_), .A3(new_n24669_), .ZN(new_n24679_));
  AOI21_X1   g24613(.A1(new_n24639_), .A2(new_n24640_), .B(new_n24665_), .ZN(new_n24680_));
  XOR2_X1    g24614(.A1(new_n24676_), .A2(\a[26] ), .Z(new_n24681_));
  OAI21_X1   g24615(.A1(new_n24680_), .A2(new_n24679_), .B(new_n24681_), .ZN(new_n24682_));
  NAND2_X1   g24616(.A1(new_n24682_), .A2(new_n24678_), .ZN(new_n24683_));
  AOI21_X1   g24617(.A1(new_n24468_), .A2(new_n24469_), .B(new_n24466_), .ZN(new_n24684_));
  NAND2_X1   g24618(.A1(new_n24684_), .A2(new_n24683_), .ZN(new_n24685_));
  NOR3_X1    g24619(.A1(new_n24680_), .A2(new_n24679_), .A3(new_n24681_), .ZN(new_n24686_));
  AOI21_X1   g24620(.A1(new_n24672_), .A2(new_n24666_), .B(new_n24677_), .ZN(new_n24687_));
  NOR2_X1    g24621(.A1(new_n24686_), .A2(new_n24687_), .ZN(new_n24688_));
  OAI21_X1   g24622(.A1(new_n24403_), .A2(new_n24462_), .B(new_n24470_), .ZN(new_n24689_));
  NAND2_X1   g24623(.A1(new_n24689_), .A2(new_n24688_), .ZN(new_n24690_));
  OAI22_X1   g24624(.A1(new_n19400_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19393_), .ZN(new_n24691_));
  NAND2_X1   g24625(.A1(new_n17790_), .A2(new_n3312_), .ZN(new_n24692_));
  AOI21_X1   g24626(.A1(new_n24692_), .A2(new_n24691_), .B(new_n3302_), .ZN(new_n24693_));
  NAND3_X1   g24627(.A1(new_n20251_), .A2(new_n84_), .A3(new_n24693_), .ZN(new_n24694_));
  INV_X1     g24628(.I(new_n24694_), .ZN(new_n24695_));
  AOI21_X1   g24629(.A1(new_n20251_), .A2(new_n24693_), .B(new_n84_), .ZN(new_n24696_));
  NOR2_X1    g24630(.A1(new_n24695_), .A2(new_n24696_), .ZN(new_n24697_));
  NAND3_X1   g24631(.A1(new_n24685_), .A2(new_n24690_), .A3(new_n24697_), .ZN(new_n24698_));
  NOR2_X1    g24632(.A1(new_n24689_), .A2(new_n24688_), .ZN(new_n24699_));
  NOR2_X1    g24633(.A1(new_n24684_), .A2(new_n24683_), .ZN(new_n24700_));
  INV_X1     g24634(.I(new_n24696_), .ZN(new_n24701_));
  NAND2_X1   g24635(.A1(new_n24701_), .A2(new_n24694_), .ZN(new_n24702_));
  OAI21_X1   g24636(.A1(new_n24700_), .A2(new_n24699_), .B(new_n24702_), .ZN(new_n24703_));
  NAND2_X1   g24637(.A1(new_n24703_), .A2(new_n24698_), .ZN(new_n24704_));
  NAND3_X1   g24638(.A1(new_n24488_), .A2(new_n24485_), .A3(new_n24482_), .ZN(new_n24705_));
  NAND2_X1   g24639(.A1(new_n24705_), .A2(new_n24704_), .ZN(new_n24706_));
  NOR3_X1    g24640(.A1(new_n24700_), .A2(new_n24699_), .A3(new_n24702_), .ZN(new_n24707_));
  AOI21_X1   g24641(.A1(new_n24685_), .A2(new_n24690_), .B(new_n24697_), .ZN(new_n24708_));
  NOR2_X1    g24642(.A1(new_n24707_), .A2(new_n24708_), .ZN(new_n24709_));
  NOR2_X1    g24643(.A1(new_n24483_), .A2(new_n24487_), .ZN(new_n24710_));
  NAND3_X1   g24644(.A1(new_n24710_), .A2(new_n24709_), .A3(new_n24485_), .ZN(new_n24711_));
  OAI22_X1   g24645(.A1(new_n19410_), .A2(new_n3769_), .B1(new_n19412_), .B2(new_n3775_), .ZN(new_n24712_));
  NAND2_X1   g24646(.A1(new_n19439_), .A2(new_n4096_), .ZN(new_n24713_));
  AOI21_X1   g24647(.A1(new_n24713_), .A2(new_n24712_), .B(new_n4095_), .ZN(new_n24714_));
  NAND2_X1   g24648(.A1(new_n20827_), .A2(new_n24714_), .ZN(new_n24715_));
  XOR2_X1    g24649(.A1(new_n24715_), .A2(new_n3035_), .Z(new_n24716_));
  NAND3_X1   g24650(.A1(new_n24706_), .A2(new_n24711_), .A3(new_n24716_), .ZN(new_n24717_));
  AOI21_X1   g24651(.A1(new_n24710_), .A2(new_n24485_), .B(new_n24709_), .ZN(new_n24718_));
  NOR4_X1    g24652(.A1(new_n24704_), .A2(new_n24478_), .A3(new_n24487_), .A4(new_n24483_), .ZN(new_n24719_));
  XOR2_X1    g24653(.A1(new_n24715_), .A2(\a[20] ), .Z(new_n24720_));
  OAI21_X1   g24654(.A1(new_n24718_), .A2(new_n24719_), .B(new_n24720_), .ZN(new_n24721_));
  NAND3_X1   g24655(.A1(new_n24499_), .A2(new_n24504_), .A3(new_n24496_), .ZN(new_n24722_));
  AOI21_X1   g24656(.A1(new_n24717_), .A2(new_n24721_), .B(new_n24722_), .ZN(new_n24723_));
  NOR3_X1    g24657(.A1(new_n24718_), .A2(new_n24719_), .A3(new_n24720_), .ZN(new_n24724_));
  AOI21_X1   g24658(.A1(new_n24706_), .A2(new_n24711_), .B(new_n24716_), .ZN(new_n24725_));
  NOR3_X1    g24659(.A1(new_n24502_), .A2(new_n24503_), .A3(new_n24500_), .ZN(new_n24726_));
  NOR3_X1    g24660(.A1(new_n24726_), .A2(new_n24725_), .A3(new_n24724_), .ZN(new_n24727_));
  NOR2_X1    g24661(.A1(new_n24723_), .A2(new_n24727_), .ZN(new_n24728_));
  INV_X1     g24662(.I(new_n24728_), .ZN(new_n24729_));
  OAI22_X1   g24663(.A1(new_n19428_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19423_), .ZN(new_n24730_));
  NAND2_X1   g24664(.A1(new_n19438_), .A2(new_n4469_), .ZN(new_n24731_));
  AOI21_X1   g24665(.A1(new_n24731_), .A2(new_n24730_), .B(new_n4468_), .ZN(new_n24732_));
  AND3_X2    g24666(.A1(new_n20907_), .A2(new_n3372_), .A3(new_n24732_), .Z(new_n24733_));
  AOI21_X1   g24667(.A1(new_n20907_), .A2(new_n24732_), .B(new_n3372_), .ZN(new_n24734_));
  NOR2_X1    g24668(.A1(new_n24733_), .A2(new_n24734_), .ZN(new_n24735_));
  NAND3_X1   g24669(.A1(new_n24517_), .A2(new_n24511_), .A3(new_n24515_), .ZN(new_n24736_));
  NAND2_X1   g24670(.A1(new_n24736_), .A2(new_n24735_), .ZN(new_n24737_));
  INV_X1     g24671(.I(new_n24735_), .ZN(new_n24738_));
  NOR2_X1    g24672(.A1(new_n24522_), .A2(new_n24516_), .ZN(new_n24739_));
  NAND3_X1   g24673(.A1(new_n24739_), .A2(new_n24511_), .A3(new_n24738_), .ZN(new_n24740_));
  AOI21_X1   g24674(.A1(new_n24740_), .A2(new_n24737_), .B(new_n24729_), .ZN(new_n24741_));
  AOI21_X1   g24675(.A1(new_n24739_), .A2(new_n24511_), .B(new_n24738_), .ZN(new_n24742_));
  NOR2_X1    g24676(.A1(new_n24736_), .A2(new_n24735_), .ZN(new_n24743_));
  NOR3_X1    g24677(.A1(new_n24742_), .A2(new_n24728_), .A3(new_n24743_), .ZN(new_n24744_));
  OAI22_X1   g24678(.A1(new_n19463_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n19437_), .ZN(new_n24745_));
  NAND2_X1   g24679(.A1(new_n17780_), .A2(new_n6090_), .ZN(new_n24746_));
  AOI21_X1   g24680(.A1(new_n24745_), .A2(new_n24746_), .B(new_n6082_), .ZN(new_n24747_));
  NAND2_X1   g24681(.A1(new_n21088_), .A2(new_n24747_), .ZN(new_n24748_));
  XOR2_X1    g24682(.A1(new_n24748_), .A2(\a[14] ), .Z(new_n24749_));
  NOR3_X1    g24683(.A1(new_n24744_), .A2(new_n24741_), .A3(new_n24749_), .ZN(new_n24750_));
  OAI21_X1   g24684(.A1(new_n24742_), .A2(new_n24743_), .B(new_n24728_), .ZN(new_n24751_));
  NAND3_X1   g24685(.A1(new_n24740_), .A2(new_n24729_), .A3(new_n24737_), .ZN(new_n24752_));
  INV_X1     g24686(.I(new_n24749_), .ZN(new_n24753_));
  AOI21_X1   g24687(.A1(new_n24751_), .A2(new_n24752_), .B(new_n24753_), .ZN(new_n24754_));
  NOR3_X1    g24688(.A1(new_n24529_), .A2(new_n24536_), .A3(new_n24537_), .ZN(new_n24755_));
  OAI21_X1   g24689(.A1(new_n24750_), .A2(new_n24754_), .B(new_n24755_), .ZN(new_n24756_));
  NAND3_X1   g24690(.A1(new_n24751_), .A2(new_n24752_), .A3(new_n24753_), .ZN(new_n24757_));
  OAI21_X1   g24691(.A1(new_n24744_), .A2(new_n24741_), .B(new_n24749_), .ZN(new_n24758_));
  INV_X1     g24692(.I(new_n24755_), .ZN(new_n24759_));
  NAND3_X1   g24693(.A1(new_n24758_), .A2(new_n24757_), .A3(new_n24759_), .ZN(new_n24760_));
  NAND2_X1   g24694(.A1(new_n24756_), .A2(new_n24760_), .ZN(new_n24761_));
  INV_X1     g24695(.I(new_n24761_), .ZN(new_n24762_));
  OAI22_X1   g24696(.A1(new_n19522_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n17775_), .ZN(new_n24763_));
  NAND2_X1   g24697(.A1(new_n17770_), .A2(new_n4709_), .ZN(new_n24764_));
  AOI21_X1   g24698(.A1(new_n24764_), .A2(new_n24763_), .B(new_n4707_), .ZN(new_n24765_));
  NAND2_X1   g24699(.A1(new_n19521_), .A2(new_n24765_), .ZN(new_n24766_));
  XOR2_X1    g24700(.A1(new_n24766_), .A2(\a[11] ), .Z(new_n24767_));
  INV_X1     g24701(.I(new_n24767_), .ZN(new_n24768_));
  NOR2_X1    g24702(.A1(new_n24557_), .A2(new_n24561_), .ZN(new_n24769_));
  AOI21_X1   g24703(.A1(new_n24769_), .A2(new_n24559_), .B(new_n24768_), .ZN(new_n24770_));
  NOR4_X1    g24704(.A1(new_n24557_), .A2(new_n24551_), .A3(new_n24561_), .A4(new_n24767_), .ZN(new_n24771_));
  OAI21_X1   g24705(.A1(new_n24770_), .A2(new_n24771_), .B(new_n24762_), .ZN(new_n24772_));
  NAND3_X1   g24706(.A1(new_n24562_), .A2(new_n24559_), .A3(new_n24556_), .ZN(new_n24773_));
  NAND2_X1   g24707(.A1(new_n24773_), .A2(new_n24767_), .ZN(new_n24774_));
  NAND4_X1   g24708(.A1(new_n24562_), .A2(new_n24559_), .A3(new_n24556_), .A4(new_n24768_), .ZN(new_n24775_));
  NAND3_X1   g24709(.A1(new_n24774_), .A2(new_n24761_), .A3(new_n24775_), .ZN(new_n24776_));
  AOI22_X1   g24710(.A1(new_n22048_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n21953_), .ZN(new_n24777_));
  NOR2_X1    g24711(.A1(new_n22115_), .A2(new_n6785_), .ZN(new_n24778_));
  OAI21_X1   g24712(.A1(new_n24778_), .A2(new_n24777_), .B(new_n6775_), .ZN(new_n24779_));
  NOR2_X1    g24713(.A1(new_n23675_), .A2(new_n24779_), .ZN(new_n24780_));
  XOR2_X1    g24714(.A1(new_n24780_), .A2(\a[8] ), .Z(new_n24781_));
  NAND3_X1   g24715(.A1(new_n24772_), .A2(new_n24776_), .A3(new_n24781_), .ZN(new_n24782_));
  AOI21_X1   g24716(.A1(new_n24774_), .A2(new_n24775_), .B(new_n24761_), .ZN(new_n24783_));
  NOR3_X1    g24717(.A1(new_n24770_), .A2(new_n24762_), .A3(new_n24771_), .ZN(new_n24784_));
  XOR2_X1    g24718(.A1(new_n24780_), .A2(new_n4009_), .Z(new_n24785_));
  OAI21_X1   g24719(.A1(new_n24784_), .A2(new_n24783_), .B(new_n24785_), .ZN(new_n24786_));
  NAND3_X1   g24720(.A1(new_n24573_), .A2(new_n24569_), .A3(new_n24578_), .ZN(new_n24787_));
  AOI21_X1   g24721(.A1(new_n24786_), .A2(new_n24782_), .B(new_n24787_), .ZN(new_n24788_));
  NOR3_X1    g24722(.A1(new_n24784_), .A2(new_n24783_), .A3(new_n24785_), .ZN(new_n24789_));
  AOI21_X1   g24723(.A1(new_n24772_), .A2(new_n24776_), .B(new_n24781_), .ZN(new_n24790_));
  INV_X1     g24724(.I(new_n24787_), .ZN(new_n24791_));
  NOR3_X1    g24725(.A1(new_n24789_), .A2(new_n24790_), .A3(new_n24791_), .ZN(new_n24792_));
  NOR2_X1    g24726(.A1(new_n24792_), .A2(new_n24788_), .ZN(new_n24793_));
  OAI22_X1   g24727(.A1(new_n23948_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n22149_), .ZN(new_n24794_));
  NAND2_X1   g24728(.A1(new_n24174_), .A2(new_n6838_), .ZN(new_n24795_));
  AOI21_X1   g24729(.A1(new_n24795_), .A2(new_n24794_), .B(new_n6836_), .ZN(new_n24796_));
  NAND2_X1   g24730(.A1(new_n24172_), .A2(new_n24796_), .ZN(new_n24797_));
  XOR2_X1    g24731(.A1(new_n24797_), .A2(new_n65_), .Z(new_n24798_));
  INV_X1     g24732(.I(new_n24585_), .ZN(new_n24799_));
  NOR3_X1    g24733(.A1(new_n24596_), .A2(new_n24590_), .A3(new_n24799_), .ZN(new_n24800_));
  NOR2_X1    g24734(.A1(new_n24800_), .A2(new_n24798_), .ZN(new_n24801_));
  XOR2_X1    g24735(.A1(new_n24797_), .A2(\a[5] ), .Z(new_n24802_));
  NOR4_X1    g24736(.A1(new_n24596_), .A2(new_n24590_), .A3(new_n24799_), .A4(new_n24802_), .ZN(new_n24803_));
  OAI21_X1   g24737(.A1(new_n24801_), .A2(new_n24803_), .B(new_n24793_), .ZN(new_n24804_));
  INV_X1     g24738(.I(new_n24793_), .ZN(new_n24805_));
  INV_X1     g24739(.I(new_n24341_), .ZN(new_n24806_));
  OAI21_X1   g24740(.A1(new_n24189_), .A2(new_n24345_), .B(new_n24806_), .ZN(new_n24807_));
  NAND3_X1   g24741(.A1(new_n24807_), .A2(new_n24585_), .A3(new_n24589_), .ZN(new_n24808_));
  NAND2_X1   g24742(.A1(new_n24808_), .A2(new_n24802_), .ZN(new_n24809_));
  NAND4_X1   g24743(.A1(new_n24807_), .A2(new_n24585_), .A3(new_n24589_), .A4(new_n24798_), .ZN(new_n24810_));
  NAND3_X1   g24744(.A1(new_n24809_), .A2(new_n24805_), .A3(new_n24810_), .ZN(new_n24811_));
  NAND2_X1   g24745(.A1(new_n24804_), .A2(new_n24811_), .ZN(new_n24812_));
  NAND2_X1   g24746(.A1(new_n354_), .A2(new_n2769_), .ZN(new_n24813_));
  NAND2_X1   g24747(.A1(new_n11226_), .A2(new_n24813_), .ZN(new_n24814_));
  NAND2_X1   g24748(.A1(new_n24603_), .A2(new_n24600_), .ZN(new_n24815_));
  NOR2_X1    g24749(.A1(new_n24814_), .A2(new_n3141_), .ZN(new_n24816_));
  AOI22_X1   g24750(.A1(new_n24815_), .A2(new_n24814_), .B1(new_n24603_), .B2(new_n24816_), .ZN(new_n24817_));
  NAND2_X1   g24751(.A1(new_n24370_), .A2(new_n24371_), .ZN(new_n24818_));
  NAND2_X1   g24752(.A1(new_n24818_), .A2(new_n24374_), .ZN(new_n24819_));
  NAND2_X1   g24753(.A1(new_n24819_), .A2(new_n24604_), .ZN(new_n24820_));
  XOR2_X1    g24754(.A1(new_n24820_), .A2(new_n24817_), .Z(new_n24821_));
  XOR2_X1    g24755(.A1(new_n24819_), .A2(new_n24604_), .Z(new_n24822_));
  NAND2_X1   g24756(.A1(new_n24822_), .A2(new_n24605_), .ZN(new_n24823_));
  NOR2_X1    g24757(.A1(new_n24821_), .A2(new_n24823_), .ZN(new_n24824_));
  AND2_X2    g24758(.A1(new_n24821_), .A2(new_n24823_), .Z(new_n24825_));
  NOR2_X1    g24759(.A1(new_n24825_), .A2(new_n24824_), .ZN(new_n24826_));
  NAND2_X1   g24760(.A1(new_n24387_), .A2(new_n24386_), .ZN(new_n24827_));
  AOI21_X1   g24761(.A1(new_n24379_), .A2(new_n24381_), .B(new_n24174_), .ZN(new_n24828_));
  OAI21_X1   g24762(.A1(new_n24828_), .A2(new_n24388_), .B(new_n24376_), .ZN(new_n24829_));
  NAND2_X1   g24763(.A1(new_n24829_), .A2(new_n24827_), .ZN(new_n24830_));
  AND3_X2    g24764(.A1(new_n24830_), .A2(new_n24615_), .A3(new_n24826_), .Z(new_n24831_));
  AOI21_X1   g24765(.A1(new_n24830_), .A2(new_n24615_), .B(new_n24826_), .ZN(new_n24832_));
  NOR2_X1    g24766(.A1(new_n24831_), .A2(new_n24832_), .ZN(new_n24833_));
  AOI22_X1   g24767(.A1(new_n24620_), .A2(new_n9503_), .B1(new_n6925_), .B2(new_n24386_), .ZN(new_n24834_));
  OR2_X2     g24768(.A1(new_n24825_), .A2(new_n24824_), .Z(new_n24835_));
  NOR2_X1    g24769(.A1(new_n24835_), .A2(new_n9489_), .ZN(new_n24836_));
  OAI21_X1   g24770(.A1(new_n24836_), .A2(new_n24834_), .B(new_n6922_), .ZN(new_n24837_));
  INV_X1     g24771(.I(new_n24837_), .ZN(new_n24838_));
  NAND2_X1   g24772(.A1(new_n24833_), .A2(new_n24838_), .ZN(new_n24839_));
  XOR2_X1    g24773(.A1(new_n24839_), .A2(\a[2] ), .Z(new_n24840_));
  XNOR2_X1   g24774(.A1(new_n24812_), .A2(new_n24840_), .ZN(new_n24841_));
  NOR2_X1    g24775(.A1(new_n24597_), .A2(new_n24624_), .ZN(new_n24842_));
  XOR2_X1    g24776(.A1(new_n24841_), .A2(new_n24842_), .Z(new_n24843_));
  INV_X1     g24777(.I(new_n24843_), .ZN(new_n24844_));
  XOR2_X1    g24778(.A1(new_n24628_), .A2(new_n24844_), .Z(\result[5] ));
  NAND2_X1   g24779(.A1(new_n24628_), .A2(new_n24844_), .ZN(new_n24846_));
  OAI21_X1   g24780(.A1(new_n24789_), .A2(new_n24790_), .B(new_n24791_), .ZN(new_n24847_));
  NAND3_X1   g24781(.A1(new_n24786_), .A2(new_n24782_), .A3(new_n24787_), .ZN(new_n24848_));
  NAND3_X1   g24782(.A1(new_n24847_), .A2(new_n24848_), .A3(new_n24798_), .ZN(new_n24849_));
  OAI21_X1   g24783(.A1(new_n24792_), .A2(new_n24788_), .B(new_n24802_), .ZN(new_n24850_));
  AOI22_X1   g24784(.A1(new_n24798_), .A2(new_n24808_), .B1(new_n24850_), .B2(new_n24849_), .ZN(new_n24851_));
  NAND3_X1   g24785(.A1(new_n24756_), .A2(new_n24760_), .A3(new_n24768_), .ZN(new_n24852_));
  AOI21_X1   g24786(.A1(new_n24756_), .A2(new_n24760_), .B(new_n24768_), .ZN(new_n24853_));
  INV_X1     g24787(.I(new_n24853_), .ZN(new_n24854_));
  AOI22_X1   g24788(.A1(new_n24854_), .A2(new_n24852_), .B1(new_n24768_), .B2(new_n24773_), .ZN(new_n24855_));
  OAI21_X1   g24789(.A1(new_n24724_), .A2(new_n24725_), .B(new_n24726_), .ZN(new_n24856_));
  NAND3_X1   g24790(.A1(new_n24722_), .A2(new_n24721_), .A3(new_n24717_), .ZN(new_n24857_));
  NAND3_X1   g24791(.A1(new_n24856_), .A2(new_n24857_), .A3(new_n24738_), .ZN(new_n24858_));
  OAI21_X1   g24792(.A1(new_n24723_), .A2(new_n24727_), .B(new_n24735_), .ZN(new_n24859_));
  AOI22_X1   g24793(.A1(new_n24736_), .A2(new_n24738_), .B1(new_n24858_), .B2(new_n24859_), .ZN(new_n24860_));
  NAND2_X1   g24794(.A1(new_n19365_), .A2(new_n3332_), .ZN(new_n24861_));
  NAND2_X1   g24795(.A1(new_n19359_), .A2(new_n3189_), .ZN(new_n24862_));
  NAND2_X1   g24796(.A1(new_n17807_), .A2(new_n2770_), .ZN(new_n24863_));
  NAND4_X1   g24797(.A1(new_n24862_), .A2(new_n2764_), .A3(new_n24861_), .A4(new_n24863_), .ZN(new_n24864_));
  INV_X1     g24798(.I(new_n24864_), .ZN(new_n24865_));
  NAND2_X1   g24799(.A1(new_n19538_), .A2(new_n24865_), .ZN(new_n24866_));
  INV_X1     g24800(.I(new_n24866_), .ZN(new_n24867_));
  NOR2_X1    g24801(.A1(new_n914_), .A2(new_n956_), .ZN(new_n24868_));
  NAND4_X1   g24802(.A1(new_n24208_), .A2(new_n2597_), .A3(new_n12034_), .A4(new_n24868_), .ZN(new_n24869_));
  NAND4_X1   g24803(.A1(new_n1305_), .A2(new_n739_), .A3(new_n665_), .A4(new_n221_), .ZN(new_n24870_));
  NOR2_X1    g24804(.A1(new_n867_), .A2(new_n485_), .ZN(new_n24871_));
  NAND4_X1   g24805(.A1(new_n327_), .A2(new_n24870_), .A3(new_n1441_), .A4(new_n24871_), .ZN(new_n24872_));
  NOR4_X1    g24806(.A1(new_n3687_), .A2(new_n563_), .A3(new_n1043_), .A4(new_n647_), .ZN(new_n24873_));
  NAND4_X1   g24807(.A1(new_n248_), .A2(new_n1628_), .A3(new_n342_), .A4(new_n761_), .ZN(new_n24874_));
  NAND4_X1   g24808(.A1(new_n1018_), .A2(new_n188_), .A3(new_n1106_), .A4(new_n1322_), .ZN(new_n24875_));
  NAND3_X1   g24809(.A1(new_n24873_), .A2(new_n24874_), .A3(new_n24875_), .ZN(new_n24876_));
  NAND3_X1   g24810(.A1(new_n3860_), .A2(new_n1594_), .A3(new_n11833_), .ZN(new_n24877_));
  NOR4_X1    g24811(.A1(new_n24877_), .A2(new_n24869_), .A3(new_n24872_), .A4(new_n24876_), .ZN(new_n24878_));
  INV_X1     g24812(.I(new_n24878_), .ZN(new_n24879_));
  OAI21_X1   g24813(.A1(new_n24658_), .A2(new_n24654_), .B(new_n24656_), .ZN(new_n24880_));
  NAND2_X1   g24814(.A1(new_n24880_), .A2(new_n24879_), .ZN(new_n24881_));
  NOR2_X1    g24815(.A1(new_n24880_), .A2(new_n24879_), .ZN(new_n24882_));
  INV_X1     g24816(.I(new_n24882_), .ZN(new_n24883_));
  AOI21_X1   g24817(.A1(new_n24883_), .A2(new_n24881_), .B(new_n24867_), .ZN(new_n24884_));
  INV_X1     g24818(.I(new_n24881_), .ZN(new_n24885_));
  NOR3_X1    g24819(.A1(new_n24885_), .A2(new_n24866_), .A3(new_n24882_), .ZN(new_n24886_));
  NOR2_X1    g24820(.A1(new_n24884_), .A2(new_n24886_), .ZN(new_n24887_));
  AOI22_X1   g24821(.A1(new_n17798_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n17802_), .ZN(new_n24888_));
  NOR2_X1    g24822(.A1(new_n19375_), .A2(new_n3175_), .ZN(new_n24889_));
  OAI21_X1   g24823(.A1(new_n24889_), .A2(new_n24888_), .B(new_n2736_), .ZN(new_n24890_));
  NOR2_X1    g24824(.A1(new_n21753_), .A2(new_n24890_), .ZN(new_n24891_));
  XOR2_X1    g24825(.A1(new_n24891_), .A2(new_n74_), .Z(new_n24892_));
  OAI21_X1   g24826(.A1(new_n24668_), .A2(new_n24669_), .B(new_n24665_), .ZN(new_n24893_));
  NAND2_X1   g24827(.A1(new_n24664_), .A2(new_n24660_), .ZN(new_n24894_));
  NAND2_X1   g24828(.A1(new_n24893_), .A2(new_n24894_), .ZN(new_n24895_));
  XOR2_X1    g24829(.A1(new_n24895_), .A2(new_n24892_), .Z(new_n24896_));
  XOR2_X1    g24830(.A1(new_n24896_), .A2(new_n24887_), .Z(new_n24897_));
  AOI22_X1   g24831(.A1(new_n19386_), .A2(new_n3267_), .B1(new_n3323_), .B2(new_n17794_), .ZN(new_n24898_));
  NOR2_X1    g24832(.A1(new_n19393_), .A2(new_n3318_), .ZN(new_n24899_));
  OAI21_X1   g24833(.A1(new_n24898_), .A2(new_n24899_), .B(new_n3259_), .ZN(new_n24900_));
  NOR2_X1    g24834(.A1(new_n20291_), .A2(new_n24900_), .ZN(new_n24901_));
  XOR2_X1    g24835(.A1(new_n24901_), .A2(new_n72_), .Z(new_n24902_));
  NAND2_X1   g24836(.A1(new_n24690_), .A2(new_n24682_), .ZN(new_n24903_));
  NAND2_X1   g24837(.A1(new_n24903_), .A2(new_n24902_), .ZN(new_n24904_));
  INV_X1     g24838(.I(new_n24902_), .ZN(new_n24905_));
  NOR2_X1    g24839(.A1(new_n24700_), .A2(new_n24687_), .ZN(new_n24906_));
  NAND2_X1   g24840(.A1(new_n24906_), .A2(new_n24905_), .ZN(new_n24907_));
  AOI21_X1   g24841(.A1(new_n24904_), .A2(new_n24907_), .B(new_n24897_), .ZN(new_n24908_));
  XNOR2_X1   g24842(.A1(new_n24896_), .A2(new_n24887_), .ZN(new_n24909_));
  NOR2_X1    g24843(.A1(new_n24906_), .A2(new_n24905_), .ZN(new_n24910_));
  NOR2_X1    g24844(.A1(new_n24903_), .A2(new_n24902_), .ZN(new_n24911_));
  NOR3_X1    g24845(.A1(new_n24909_), .A2(new_n24911_), .A3(new_n24910_), .ZN(new_n24912_));
  NOR2_X1    g24846(.A1(new_n24908_), .A2(new_n24912_), .ZN(new_n24913_));
  OAI22_X1   g24847(.A1(new_n17789_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19400_), .ZN(new_n24914_));
  NAND2_X1   g24848(.A1(new_n19407_), .A2(new_n3312_), .ZN(new_n24915_));
  AOI21_X1   g24849(.A1(new_n24915_), .A2(new_n24914_), .B(new_n3302_), .ZN(new_n24916_));
  NAND2_X1   g24850(.A1(new_n20864_), .A2(new_n24916_), .ZN(new_n24917_));
  XOR2_X1    g24851(.A1(new_n24917_), .A2(\a[23] ), .Z(new_n24918_));
  INV_X1     g24852(.I(new_n24918_), .ZN(new_n24919_));
  NAND2_X1   g24853(.A1(new_n24705_), .A2(new_n24709_), .ZN(new_n24920_));
  AOI21_X1   g24854(.A1(new_n24920_), .A2(new_n24698_), .B(new_n24919_), .ZN(new_n24921_));
  AOI21_X1   g24855(.A1(new_n24710_), .A2(new_n24485_), .B(new_n24704_), .ZN(new_n24922_));
  NOR3_X1    g24856(.A1(new_n24922_), .A2(new_n24707_), .A3(new_n24918_), .ZN(new_n24923_));
  OAI21_X1   g24857(.A1(new_n24921_), .A2(new_n24923_), .B(new_n24913_), .ZN(new_n24924_));
  OAI21_X1   g24858(.A1(new_n24910_), .A2(new_n24911_), .B(new_n24909_), .ZN(new_n24925_));
  NAND3_X1   g24859(.A1(new_n24897_), .A2(new_n24907_), .A3(new_n24904_), .ZN(new_n24926_));
  NAND2_X1   g24860(.A1(new_n24925_), .A2(new_n24926_), .ZN(new_n24927_));
  OAI21_X1   g24861(.A1(new_n24922_), .A2(new_n24707_), .B(new_n24918_), .ZN(new_n24928_));
  NAND3_X1   g24862(.A1(new_n24920_), .A2(new_n24698_), .A3(new_n24919_), .ZN(new_n24929_));
  NAND3_X1   g24863(.A1(new_n24929_), .A2(new_n24928_), .A3(new_n24927_), .ZN(new_n24930_));
  NAND2_X1   g24864(.A1(new_n24924_), .A2(new_n24930_), .ZN(new_n24931_));
  OAI22_X1   g24865(.A1(new_n17787_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19412_), .ZN(new_n24932_));
  NAND2_X1   g24866(.A1(new_n19442_), .A2(new_n4096_), .ZN(new_n24933_));
  AOI21_X1   g24867(.A1(new_n24933_), .A2(new_n24932_), .B(new_n4095_), .ZN(new_n24934_));
  NAND2_X1   g24868(.A1(new_n20939_), .A2(new_n24934_), .ZN(new_n24935_));
  XOR2_X1    g24869(.A1(new_n24935_), .A2(\a[20] ), .Z(new_n24936_));
  OAI21_X1   g24870(.A1(new_n24726_), .A2(new_n24724_), .B(new_n24721_), .ZN(new_n24937_));
  NAND2_X1   g24871(.A1(new_n24937_), .A2(new_n24936_), .ZN(new_n24938_));
  INV_X1     g24872(.I(new_n24936_), .ZN(new_n24939_));
  AOI21_X1   g24873(.A1(new_n24722_), .A2(new_n24717_), .B(new_n24725_), .ZN(new_n24940_));
  NAND2_X1   g24874(.A1(new_n24940_), .A2(new_n24939_), .ZN(new_n24941_));
  AOI21_X1   g24875(.A1(new_n24941_), .A2(new_n24938_), .B(new_n24931_), .ZN(new_n24942_));
  AOI21_X1   g24876(.A1(new_n24929_), .A2(new_n24928_), .B(new_n24927_), .ZN(new_n24943_));
  NOR3_X1    g24877(.A1(new_n24921_), .A2(new_n24923_), .A3(new_n24913_), .ZN(new_n24944_));
  NOR2_X1    g24878(.A1(new_n24943_), .A2(new_n24944_), .ZN(new_n24945_));
  NOR2_X1    g24879(.A1(new_n24940_), .A2(new_n24939_), .ZN(new_n24946_));
  NOR2_X1    g24880(.A1(new_n24937_), .A2(new_n24936_), .ZN(new_n24947_));
  NOR3_X1    g24881(.A1(new_n24946_), .A2(new_n24947_), .A3(new_n24945_), .ZN(new_n24948_));
  NOR2_X1    g24882(.A1(new_n24948_), .A2(new_n24942_), .ZN(new_n24949_));
  INV_X1     g24883(.I(new_n24949_), .ZN(new_n24950_));
  OAI22_X1   g24884(.A1(new_n17784_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19428_), .ZN(new_n24951_));
  NAND2_X1   g24885(.A1(new_n19466_), .A2(new_n4469_), .ZN(new_n24952_));
  AOI21_X1   g24886(.A1(new_n24952_), .A2(new_n24951_), .B(new_n4468_), .ZN(new_n24953_));
  NAND2_X1   g24887(.A1(new_n21100_), .A2(new_n24953_), .ZN(new_n24954_));
  XOR2_X1    g24888(.A1(new_n24954_), .A2(\a[17] ), .Z(new_n24955_));
  INV_X1     g24889(.I(new_n24955_), .ZN(new_n24956_));
  NOR2_X1    g24890(.A1(new_n24950_), .A2(new_n24956_), .ZN(new_n24957_));
  NOR2_X1    g24891(.A1(new_n24949_), .A2(new_n24955_), .ZN(new_n24958_));
  OAI21_X1   g24892(.A1(new_n24957_), .A2(new_n24958_), .B(new_n24860_), .ZN(new_n24959_));
  OAI21_X1   g24893(.A1(new_n24946_), .A2(new_n24947_), .B(new_n24945_), .ZN(new_n24960_));
  NAND3_X1   g24894(.A1(new_n24938_), .A2(new_n24941_), .A3(new_n24931_), .ZN(new_n24961_));
  AOI21_X1   g24895(.A1(new_n24960_), .A2(new_n24961_), .B(new_n24956_), .ZN(new_n24962_));
  NOR3_X1    g24896(.A1(new_n24948_), .A2(new_n24942_), .A3(new_n24955_), .ZN(new_n24963_));
  NOR2_X1    g24897(.A1(new_n24962_), .A2(new_n24963_), .ZN(new_n24964_));
  OR2_X2     g24898(.A1(new_n24964_), .A2(new_n24860_), .Z(new_n24965_));
  NAND2_X1   g24899(.A1(new_n24965_), .A2(new_n24959_), .ZN(new_n24966_));
  INV_X1     g24900(.I(new_n24966_), .ZN(new_n24967_));
  OAI22_X1   g24901(.A1(new_n19475_), .A2(new_n6094_), .B1(new_n19463_), .B2(new_n6089_), .ZN(new_n24968_));
  NAND2_X1   g24902(.A1(new_n19484_), .A2(new_n6090_), .ZN(new_n24969_));
  AOI21_X1   g24903(.A1(new_n24969_), .A2(new_n24968_), .B(new_n6082_), .ZN(new_n24970_));
  NAND2_X1   g24904(.A1(new_n21171_), .A2(new_n24970_), .ZN(new_n24971_));
  XOR2_X1    g24905(.A1(new_n24971_), .A2(\a[14] ), .Z(new_n24972_));
  INV_X1     g24906(.I(new_n24972_), .ZN(new_n24973_));
  AOI21_X1   g24907(.A1(new_n24760_), .A2(new_n24758_), .B(new_n24973_), .ZN(new_n24974_));
  OAI21_X1   g24908(.A1(new_n24750_), .A2(new_n24755_), .B(new_n24758_), .ZN(new_n24975_));
  NOR2_X1    g24909(.A1(new_n24975_), .A2(new_n24972_), .ZN(new_n24976_));
  OAI21_X1   g24910(.A1(new_n24976_), .A2(new_n24974_), .B(new_n24967_), .ZN(new_n24977_));
  NAND2_X1   g24911(.A1(new_n24975_), .A2(new_n24972_), .ZN(new_n24978_));
  NAND3_X1   g24912(.A1(new_n24760_), .A2(new_n24758_), .A3(new_n24973_), .ZN(new_n24979_));
  NAND3_X1   g24913(.A1(new_n24978_), .A2(new_n24979_), .A3(new_n24966_), .ZN(new_n24980_));
  OAI22_X1   g24914(.A1(new_n19512_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n19522_), .ZN(new_n24981_));
  NAND2_X1   g24915(.A1(new_n21953_), .A2(new_n4709_), .ZN(new_n24982_));
  AOI21_X1   g24916(.A1(new_n24981_), .A2(new_n24982_), .B(new_n4707_), .ZN(new_n24983_));
  NAND2_X1   g24917(.A1(new_n21963_), .A2(new_n24983_), .ZN(new_n24984_));
  XOR2_X1    g24918(.A1(new_n24984_), .A2(\a[11] ), .Z(new_n24985_));
  NAND3_X1   g24919(.A1(new_n24977_), .A2(new_n24980_), .A3(new_n24985_), .ZN(new_n24986_));
  INV_X1     g24920(.I(new_n24986_), .ZN(new_n24987_));
  AOI21_X1   g24921(.A1(new_n24977_), .A2(new_n24980_), .B(new_n24985_), .ZN(new_n24988_));
  OAI21_X1   g24922(.A1(new_n24987_), .A2(new_n24988_), .B(new_n24855_), .ZN(new_n24989_));
  INV_X1     g24923(.I(new_n24855_), .ZN(new_n24990_));
  AOI21_X1   g24924(.A1(new_n24978_), .A2(new_n24979_), .B(new_n24966_), .ZN(new_n24991_));
  NOR3_X1    g24925(.A1(new_n24976_), .A2(new_n24974_), .A3(new_n24967_), .ZN(new_n24992_));
  OAI21_X1   g24926(.A1(new_n24992_), .A2(new_n24991_), .B(new_n24985_), .ZN(new_n24993_));
  INV_X1     g24927(.I(new_n24985_), .ZN(new_n24994_));
  NAND3_X1   g24928(.A1(new_n24977_), .A2(new_n24980_), .A3(new_n24994_), .ZN(new_n24995_));
  NAND2_X1   g24929(.A1(new_n24993_), .A2(new_n24995_), .ZN(new_n24996_));
  NAND2_X1   g24930(.A1(new_n24996_), .A2(new_n24990_), .ZN(new_n24997_));
  NAND2_X1   g24931(.A1(new_n24997_), .A2(new_n24989_), .ZN(new_n24998_));
  OAI22_X1   g24932(.A1(new_n22115_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n22051_), .ZN(new_n24999_));
  NAND2_X1   g24933(.A1(new_n22150_), .A2(new_n6784_), .ZN(new_n25000_));
  AOI21_X1   g24934(.A1(new_n24999_), .A2(new_n25000_), .B(new_n6776_), .ZN(new_n25001_));
  NAND2_X1   g24935(.A1(new_n22163_), .A2(new_n25001_), .ZN(new_n25002_));
  XOR2_X1    g24936(.A1(new_n25002_), .A2(\a[8] ), .Z(new_n25003_));
  OAI21_X1   g24937(.A1(new_n24789_), .A2(new_n24791_), .B(new_n24786_), .ZN(new_n25004_));
  NAND2_X1   g24938(.A1(new_n25004_), .A2(new_n25003_), .ZN(new_n25005_));
  INV_X1     g24939(.I(new_n25003_), .ZN(new_n25006_));
  NAND3_X1   g24940(.A1(new_n24848_), .A2(new_n24786_), .A3(new_n25006_), .ZN(new_n25007_));
  AOI21_X1   g24941(.A1(new_n25005_), .A2(new_n25007_), .B(new_n24998_), .ZN(new_n25008_));
  INV_X1     g24942(.I(new_n24988_), .ZN(new_n25009_));
  AOI21_X1   g24943(.A1(new_n25009_), .A2(new_n24986_), .B(new_n24990_), .ZN(new_n25010_));
  AOI21_X1   g24944(.A1(new_n24990_), .A2(new_n24996_), .B(new_n25010_), .ZN(new_n25011_));
  AOI21_X1   g24945(.A1(new_n24848_), .A2(new_n24786_), .B(new_n25006_), .ZN(new_n25012_));
  NOR2_X1    g24946(.A1(new_n25004_), .A2(new_n25003_), .ZN(new_n25013_));
  NOR3_X1    g24947(.A1(new_n25013_), .A2(new_n25012_), .A3(new_n25011_), .ZN(new_n25014_));
  AOI21_X1   g24948(.A1(new_n24376_), .A2(new_n24388_), .B(new_n24828_), .ZN(new_n25015_));
  AOI21_X1   g24949(.A1(new_n25015_), .A2(new_n24826_), .B(new_n24386_), .ZN(new_n25017_));
  OAI22_X1   g24950(.A1(new_n24835_), .A2(new_n13965_), .B1(new_n9485_), .B2(new_n24613_), .ZN(new_n25018_));
  NAND2_X1   g24951(.A1(new_n25018_), .A2(new_n6922_), .ZN(new_n25019_));
  NOR2_X1    g24952(.A1(new_n25017_), .A2(new_n25019_), .ZN(new_n25020_));
  NAND2_X1   g24953(.A1(new_n25020_), .A2(new_n4387_), .ZN(new_n25021_));
  OAI21_X1   g24954(.A1(new_n25017_), .A2(new_n25019_), .B(\a[2] ), .ZN(new_n25022_));
  NAND2_X1   g24955(.A1(new_n25021_), .A2(new_n25022_), .ZN(new_n25023_));
  AOI22_X1   g24956(.A1(new_n24174_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n23957_), .ZN(new_n25024_));
  NOR2_X1    g24957(.A1(new_n24376_), .A2(new_n6839_), .ZN(new_n25025_));
  OAI21_X1   g24958(.A1(new_n25025_), .A2(new_n25024_), .B(new_n6835_), .ZN(new_n25026_));
  NOR3_X1    g24959(.A1(new_n24385_), .A2(new_n24389_), .A3(new_n25026_), .ZN(new_n25027_));
  XOR2_X1    g24960(.A1(new_n25027_), .A2(new_n65_), .Z(new_n25028_));
  NAND2_X1   g24961(.A1(new_n25023_), .A2(new_n25028_), .ZN(new_n25029_));
  NOR3_X1    g24962(.A1(new_n25017_), .A2(\a[2] ), .A3(new_n25019_), .ZN(new_n25030_));
  INV_X1     g24963(.I(new_n25022_), .ZN(new_n25031_));
  NOR2_X1    g24964(.A1(new_n25031_), .A2(new_n25030_), .ZN(new_n25032_));
  XOR2_X1    g24965(.A1(new_n25027_), .A2(\a[5] ), .Z(new_n25033_));
  NAND2_X1   g24966(.A1(new_n25032_), .A2(new_n25033_), .ZN(new_n25034_));
  NAND2_X1   g24967(.A1(new_n25034_), .A2(new_n25029_), .ZN(new_n25035_));
  OAI21_X1   g24968(.A1(new_n25014_), .A2(new_n25008_), .B(new_n25035_), .ZN(new_n25036_));
  OAI21_X1   g24969(.A1(new_n25013_), .A2(new_n25012_), .B(new_n25011_), .ZN(new_n25037_));
  NAND3_X1   g24970(.A1(new_n25005_), .A2(new_n25007_), .A3(new_n24998_), .ZN(new_n25038_));
  NAND3_X1   g24971(.A1(new_n25028_), .A2(new_n25021_), .A3(new_n25022_), .ZN(new_n25039_));
  NAND2_X1   g24972(.A1(new_n25023_), .A2(new_n25033_), .ZN(new_n25040_));
  NAND2_X1   g24973(.A1(new_n25040_), .A2(new_n25039_), .ZN(new_n25041_));
  NAND3_X1   g24974(.A1(new_n25037_), .A2(new_n25038_), .A3(new_n25041_), .ZN(new_n25042_));
  NAND2_X1   g24975(.A1(new_n25036_), .A2(new_n25042_), .ZN(new_n25043_));
  AOI21_X1   g24976(.A1(new_n24812_), .A2(new_n24840_), .B(new_n24842_), .ZN(new_n25044_));
  XOR2_X1    g24977(.A1(new_n25044_), .A2(new_n25043_), .Z(new_n25045_));
  XOR2_X1    g24978(.A1(new_n25045_), .A2(new_n24851_), .Z(new_n25046_));
  XOR2_X1    g24979(.A1(new_n24846_), .A2(new_n25046_), .Z(\result[6] ));
  OAI22_X1   g24980(.A1(new_n24376_), .A2(new_n6843_), .B1(new_n6913_), .B2(new_n24167_), .ZN(new_n25048_));
  NAND2_X1   g24981(.A1(new_n24620_), .A2(new_n6838_), .ZN(new_n25049_));
  AOI21_X1   g24982(.A1(new_n25049_), .A2(new_n25048_), .B(new_n6836_), .ZN(new_n25050_));
  NAND2_X1   g24983(.A1(new_n24618_), .A2(new_n25050_), .ZN(new_n25051_));
  XOR2_X1    g24984(.A1(new_n25051_), .A2(new_n65_), .Z(new_n25052_));
  OAI22_X1   g24985(.A1(new_n22115_), .A2(new_n6783_), .B1(new_n6788_), .B2(new_n22149_), .ZN(new_n25053_));
  NAND2_X1   g24986(.A1(new_n23957_), .A2(new_n6784_), .ZN(new_n25054_));
  AOI21_X1   g24987(.A1(new_n25053_), .A2(new_n25054_), .B(new_n6776_), .ZN(new_n25055_));
  NAND2_X1   g24988(.A1(new_n23955_), .A2(new_n25055_), .ZN(new_n25056_));
  XOR2_X1    g24989(.A1(new_n25056_), .A2(\a[8] ), .Z(new_n25057_));
  OAI22_X1   g24990(.A1(new_n19512_), .A2(new_n4716_), .B1(new_n21960_), .B2(new_n4719_), .ZN(new_n25058_));
  NAND2_X1   g24991(.A1(new_n22048_), .A2(new_n4709_), .ZN(new_n25059_));
  AOI21_X1   g24992(.A1(new_n25059_), .A2(new_n25058_), .B(new_n4707_), .ZN(new_n25060_));
  NAND2_X1   g24993(.A1(new_n22175_), .A2(new_n25060_), .ZN(new_n25061_));
  XOR2_X1    g24994(.A1(new_n25061_), .A2(\a[11] ), .Z(new_n25062_));
  INV_X1     g24995(.I(new_n25062_), .ZN(new_n25063_));
  OAI22_X1   g24996(.A1(new_n17775_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n19475_), .ZN(new_n25064_));
  NAND2_X1   g24997(.A1(new_n21157_), .A2(new_n6090_), .ZN(new_n25065_));
  AOI21_X1   g24998(.A1(new_n25065_), .A2(new_n25064_), .B(new_n6082_), .ZN(new_n25066_));
  AND3_X2    g24999(.A1(new_n21155_), .A2(new_n3521_), .A3(new_n25066_), .Z(new_n25067_));
  AOI21_X1   g25000(.A1(new_n21155_), .A2(new_n25066_), .B(new_n3521_), .ZN(new_n25068_));
  NOR2_X1    g25001(.A1(new_n25067_), .A2(new_n25068_), .ZN(new_n25069_));
  INV_X1     g25002(.I(new_n25069_), .ZN(new_n25070_));
  OAI22_X1   g25003(.A1(new_n19437_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n17784_), .ZN(new_n25071_));
  NAND2_X1   g25004(.A1(new_n19472_), .A2(new_n4469_), .ZN(new_n25072_));
  AOI21_X1   g25005(.A1(new_n25072_), .A2(new_n25071_), .B(new_n4468_), .ZN(new_n25073_));
  NAND2_X1   g25006(.A1(new_n21117_), .A2(new_n25073_), .ZN(new_n25074_));
  XOR2_X1    g25007(.A1(new_n25074_), .A2(\a[17] ), .Z(new_n25075_));
  OAI22_X1   g25008(.A1(new_n19423_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n17787_), .ZN(new_n25076_));
  NAND2_X1   g25009(.A1(new_n20896_), .A2(new_n4096_), .ZN(new_n25077_));
  AOI21_X1   g25010(.A1(new_n25077_), .A2(new_n25076_), .B(new_n4095_), .ZN(new_n25078_));
  NAND3_X1   g25011(.A1(new_n22226_), .A2(new_n3035_), .A3(new_n25078_), .ZN(new_n25079_));
  NAND2_X1   g25012(.A1(new_n22226_), .A2(new_n25078_), .ZN(new_n25080_));
  NAND2_X1   g25013(.A1(new_n25080_), .A2(\a[20] ), .ZN(new_n25081_));
  NAND2_X1   g25014(.A1(new_n25081_), .A2(new_n25079_), .ZN(new_n25082_));
  OAI22_X1   g25015(.A1(new_n19410_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n17789_), .ZN(new_n25083_));
  NAND2_X1   g25016(.A1(new_n19415_), .A2(new_n3312_), .ZN(new_n25084_));
  AOI21_X1   g25017(.A1(new_n25084_), .A2(new_n25083_), .B(new_n3302_), .ZN(new_n25085_));
  NAND2_X1   g25018(.A1(new_n20846_), .A2(new_n25085_), .ZN(new_n25086_));
  XOR2_X1    g25019(.A1(new_n25086_), .A2(\a[23] ), .Z(new_n25087_));
  OAI22_X1   g25020(.A1(new_n19393_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n17793_), .ZN(new_n25088_));
  NAND2_X1   g25021(.A1(new_n19399_), .A2(new_n3317_), .ZN(new_n25089_));
  AOI21_X1   g25022(.A1(new_n25089_), .A2(new_n25088_), .B(new_n3260_), .ZN(new_n25090_));
  NAND2_X1   g25023(.A1(new_n20264_), .A2(new_n25090_), .ZN(new_n25091_));
  XOR2_X1    g25024(.A1(new_n25091_), .A2(\a[26] ), .Z(new_n25092_));
  NOR2_X1    g25025(.A1(new_n24835_), .A2(new_n11783_), .ZN(new_n25093_));
  AOI21_X1   g25026(.A1(new_n24826_), .A2(new_n6924_), .B(\a[2] ), .ZN(new_n25094_));
  NOR2_X1    g25027(.A1(new_n25093_), .A2(new_n25094_), .ZN(new_n25095_));
  NAND2_X1   g25028(.A1(new_n17802_), .A2(new_n3332_), .ZN(new_n25096_));
  NAND2_X1   g25029(.A1(new_n19365_), .A2(new_n3189_), .ZN(new_n25097_));
  AOI21_X1   g25030(.A1(new_n19359_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n25098_));
  NAND3_X1   g25031(.A1(new_n25098_), .A2(new_n25096_), .A3(new_n25097_), .ZN(new_n25099_));
  INV_X1     g25032(.I(new_n25099_), .ZN(new_n25100_));
  NAND2_X1   g25033(.A1(new_n19951_), .A2(new_n25100_), .ZN(new_n25101_));
  INV_X1     g25034(.I(new_n25101_), .ZN(new_n25102_));
  NAND4_X1   g25035(.A1(new_n373_), .A2(new_n934_), .A3(new_n1572_), .A4(new_n1325_), .ZN(new_n25103_));
  NAND4_X1   g25036(.A1(new_n2130_), .A2(new_n4843_), .A3(new_n11576_), .A4(new_n25103_), .ZN(new_n25104_));
  NOR3_X1    g25037(.A1(new_n12958_), .A2(new_n1486_), .A3(new_n1561_), .ZN(new_n25105_));
  NOR3_X1    g25038(.A1(new_n549_), .A2(new_n456_), .A3(new_n397_), .ZN(new_n25106_));
  NAND4_X1   g25039(.A1(new_n25105_), .A2(new_n777_), .A3(new_n2606_), .A4(new_n25106_), .ZN(new_n25107_));
  OR2_X2     g25040(.A1(new_n1517_), .A2(new_n2696_), .Z(new_n25108_));
  NOR4_X1    g25041(.A1(new_n25108_), .A2(new_n10988_), .A3(new_n25104_), .A4(new_n25107_), .ZN(new_n25109_));
  NAND3_X1   g25042(.A1(new_n25109_), .A2(new_n1762_), .A3(new_n2585_), .ZN(new_n25110_));
  INV_X1     g25043(.I(new_n25110_), .ZN(new_n25111_));
  NOR2_X1    g25044(.A1(new_n25102_), .A2(new_n25111_), .ZN(new_n25112_));
  NOR2_X1    g25045(.A1(new_n25101_), .A2(new_n25110_), .ZN(new_n25113_));
  NOR2_X1    g25046(.A1(new_n25112_), .A2(new_n25113_), .ZN(new_n25114_));
  XOR2_X1    g25047(.A1(new_n25101_), .A2(new_n25110_), .Z(new_n25115_));
  NAND2_X1   g25048(.A1(new_n25115_), .A2(new_n25095_), .ZN(new_n25116_));
  OAI21_X1   g25049(.A1(new_n25095_), .A2(new_n25114_), .B(new_n25116_), .ZN(new_n25117_));
  OAI22_X1   g25050(.A1(new_n19375_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n17797_), .ZN(new_n25118_));
  NAND2_X1   g25051(.A1(new_n19386_), .A2(new_n2750_), .ZN(new_n25119_));
  AOI21_X1   g25052(.A1(new_n25119_), .A2(new_n25118_), .B(new_n2737_), .ZN(new_n25120_));
  NAND3_X1   g25053(.A1(new_n20162_), .A2(new_n74_), .A3(new_n25120_), .ZN(new_n25121_));
  INV_X1     g25054(.I(new_n25121_), .ZN(new_n25122_));
  AOI21_X1   g25055(.A1(new_n20162_), .A2(new_n25120_), .B(new_n74_), .ZN(new_n25123_));
  INV_X1     g25056(.I(new_n24880_), .ZN(new_n25124_));
  XOR2_X1    g25057(.A1(new_n24866_), .A2(new_n24879_), .Z(new_n25125_));
  OAI21_X1   g25058(.A1(new_n25124_), .A2(new_n24879_), .B(new_n25125_), .ZN(new_n25126_));
  OAI21_X1   g25059(.A1(new_n25122_), .A2(new_n25123_), .B(new_n25126_), .ZN(new_n25127_));
  INV_X1     g25060(.I(new_n25127_), .ZN(new_n25128_));
  NOR3_X1    g25061(.A1(new_n25122_), .A2(new_n25123_), .A3(new_n25126_), .ZN(new_n25129_));
  OAI21_X1   g25062(.A1(new_n25128_), .A2(new_n25129_), .B(new_n25117_), .ZN(new_n25130_));
  INV_X1     g25063(.I(new_n25117_), .ZN(new_n25131_));
  INV_X1     g25064(.I(new_n25126_), .ZN(new_n25132_));
  NOR3_X1    g25065(.A1(new_n25122_), .A2(new_n25132_), .A3(new_n25123_), .ZN(new_n25133_));
  INV_X1     g25066(.I(new_n25123_), .ZN(new_n25134_));
  AOI21_X1   g25067(.A1(new_n25134_), .A2(new_n25121_), .B(new_n25126_), .ZN(new_n25135_));
  OAI21_X1   g25068(.A1(new_n25133_), .A2(new_n25135_), .B(new_n25131_), .ZN(new_n25136_));
  NAND2_X1   g25069(.A1(new_n25130_), .A2(new_n25136_), .ZN(new_n25137_));
  XOR2_X1    g25070(.A1(new_n24891_), .A2(\a[29] ), .Z(new_n25138_));
  AOI21_X1   g25071(.A1(new_n24639_), .A2(new_n24640_), .B(new_n24671_), .ZN(new_n25139_));
  NOR3_X1    g25072(.A1(new_n24892_), .A2(new_n24884_), .A3(new_n24886_), .ZN(new_n25140_));
  OAI21_X1   g25073(.A1(new_n24885_), .A2(new_n24882_), .B(new_n24866_), .ZN(new_n25141_));
  NAND3_X1   g25074(.A1(new_n24883_), .A2(new_n24867_), .A3(new_n24881_), .ZN(new_n25142_));
  AOI21_X1   g25075(.A1(new_n25141_), .A2(new_n25142_), .B(new_n25138_), .ZN(new_n25143_));
  OAI21_X1   g25076(.A1(new_n25143_), .A2(new_n25140_), .B(new_n24894_), .ZN(new_n25144_));
  OAI22_X1   g25077(.A1(new_n25144_), .A2(new_n25139_), .B1(new_n24887_), .B2(new_n25138_), .ZN(new_n25145_));
  NOR2_X1    g25078(.A1(new_n25145_), .A2(new_n25137_), .ZN(new_n25146_));
  INV_X1     g25079(.I(new_n25129_), .ZN(new_n25147_));
  AOI21_X1   g25080(.A1(new_n25147_), .A2(new_n25127_), .B(new_n25131_), .ZN(new_n25148_));
  INV_X1     g25081(.I(new_n25136_), .ZN(new_n25149_));
  NOR2_X1    g25082(.A1(new_n25149_), .A2(new_n25148_), .ZN(new_n25150_));
  NOR2_X1    g25083(.A1(new_n24887_), .A2(new_n25138_), .ZN(new_n25151_));
  NAND3_X1   g25084(.A1(new_n25138_), .A2(new_n25141_), .A3(new_n25142_), .ZN(new_n25152_));
  OAI21_X1   g25085(.A1(new_n24886_), .A2(new_n24884_), .B(new_n24892_), .ZN(new_n25153_));
  AOI22_X1   g25086(.A1(new_n25153_), .A2(new_n25152_), .B1(new_n24660_), .B2(new_n24664_), .ZN(new_n25154_));
  AOI21_X1   g25087(.A1(new_n25154_), .A2(new_n24893_), .B(new_n25151_), .ZN(new_n25155_));
  NOR2_X1    g25088(.A1(new_n25155_), .A2(new_n25150_), .ZN(new_n25156_));
  OAI21_X1   g25089(.A1(new_n25156_), .A2(new_n25146_), .B(new_n25092_), .ZN(new_n25157_));
  INV_X1     g25090(.I(new_n25092_), .ZN(new_n25158_));
  NAND2_X1   g25091(.A1(new_n25155_), .A2(new_n25150_), .ZN(new_n25159_));
  NAND2_X1   g25092(.A1(new_n25145_), .A2(new_n25137_), .ZN(new_n25160_));
  NAND3_X1   g25093(.A1(new_n25159_), .A2(new_n25160_), .A3(new_n25158_), .ZN(new_n25161_));
  NAND2_X1   g25094(.A1(new_n25157_), .A2(new_n25161_), .ZN(new_n25162_));
  NAND2_X1   g25095(.A1(new_n25162_), .A2(new_n25087_), .ZN(new_n25163_));
  INV_X1     g25096(.I(new_n25087_), .ZN(new_n25164_));
  AOI21_X1   g25097(.A1(new_n25159_), .A2(new_n25160_), .B(new_n25158_), .ZN(new_n25165_));
  NOR3_X1    g25098(.A1(new_n25156_), .A2(new_n25146_), .A3(new_n25092_), .ZN(new_n25166_));
  NOR2_X1    g25099(.A1(new_n25165_), .A2(new_n25166_), .ZN(new_n25167_));
  NAND2_X1   g25100(.A1(new_n25167_), .A2(new_n25164_), .ZN(new_n25168_));
  NAND2_X1   g25101(.A1(new_n25168_), .A2(new_n25163_), .ZN(new_n25169_));
  XNOR2_X1   g25102(.A1(new_n25082_), .A2(new_n25169_), .ZN(new_n25170_));
  INV_X1     g25103(.I(new_n25170_), .ZN(new_n25171_));
  OAI21_X1   g25104(.A1(new_n24948_), .A2(new_n24942_), .B(new_n24955_), .ZN(new_n25172_));
  AOI21_X1   g25105(.A1(new_n24860_), .A2(new_n25172_), .B(new_n24963_), .ZN(new_n25173_));
  NOR2_X1    g25106(.A1(new_n25173_), .A2(new_n25171_), .ZN(new_n25174_));
  NAND2_X1   g25107(.A1(new_n24729_), .A2(new_n24735_), .ZN(new_n25175_));
  NAND2_X1   g25108(.A1(new_n24859_), .A2(new_n24858_), .ZN(new_n25176_));
  NAND3_X1   g25109(.A1(new_n24739_), .A2(new_n25176_), .A3(new_n24511_), .ZN(new_n25177_));
  AOI21_X1   g25110(.A1(new_n25177_), .A2(new_n25175_), .B(new_n24962_), .ZN(new_n25178_));
  NOR3_X1    g25111(.A1(new_n25178_), .A2(new_n24963_), .A3(new_n25170_), .ZN(new_n25179_));
  OAI21_X1   g25112(.A1(new_n25179_), .A2(new_n25174_), .B(new_n25075_), .ZN(new_n25180_));
  INV_X1     g25113(.I(new_n25075_), .ZN(new_n25181_));
  OAI21_X1   g25114(.A1(new_n25178_), .A2(new_n24963_), .B(new_n25170_), .ZN(new_n25182_));
  NAND2_X1   g25115(.A1(new_n25173_), .A2(new_n25171_), .ZN(new_n25183_));
  NAND3_X1   g25116(.A1(new_n25182_), .A2(new_n25183_), .A3(new_n25181_), .ZN(new_n25184_));
  AOI21_X1   g25117(.A1(new_n25180_), .A2(new_n25184_), .B(new_n25070_), .ZN(new_n25185_));
  AOI21_X1   g25118(.A1(new_n25182_), .A2(new_n25183_), .B(new_n25181_), .ZN(new_n25186_));
  NOR3_X1    g25119(.A1(new_n25179_), .A2(new_n25174_), .A3(new_n25075_), .ZN(new_n25187_));
  NOR3_X1    g25120(.A1(new_n25187_), .A2(new_n25186_), .A3(new_n25069_), .ZN(new_n25188_));
  NOR2_X1    g25121(.A1(new_n25188_), .A2(new_n25185_), .ZN(new_n25189_));
  NAND2_X1   g25122(.A1(new_n24993_), .A2(new_n24855_), .ZN(new_n25190_));
  NAND2_X1   g25123(.A1(new_n25190_), .A2(new_n24995_), .ZN(new_n25191_));
  NAND2_X1   g25124(.A1(new_n25191_), .A2(new_n25189_), .ZN(new_n25192_));
  OAI21_X1   g25125(.A1(new_n25187_), .A2(new_n25186_), .B(new_n25069_), .ZN(new_n25193_));
  NAND3_X1   g25126(.A1(new_n25180_), .A2(new_n25184_), .A3(new_n25070_), .ZN(new_n25194_));
  NAND2_X1   g25127(.A1(new_n25193_), .A2(new_n25194_), .ZN(new_n25195_));
  NOR3_X1    g25128(.A1(new_n24992_), .A2(new_n24991_), .A3(new_n24985_), .ZN(new_n25196_));
  AOI21_X1   g25129(.A1(new_n24855_), .A2(new_n24993_), .B(new_n25196_), .ZN(new_n25197_));
  NAND2_X1   g25130(.A1(new_n25197_), .A2(new_n25195_), .ZN(new_n25198_));
  AOI21_X1   g25131(.A1(new_n25192_), .A2(new_n25198_), .B(new_n25063_), .ZN(new_n25199_));
  NOR2_X1    g25132(.A1(new_n25197_), .A2(new_n25195_), .ZN(new_n25200_));
  NOR2_X1    g25133(.A1(new_n25191_), .A2(new_n25189_), .ZN(new_n25201_));
  NOR3_X1    g25134(.A1(new_n25201_), .A2(new_n25062_), .A3(new_n25200_), .ZN(new_n25202_));
  OAI21_X1   g25135(.A1(new_n25202_), .A2(new_n25199_), .B(new_n25057_), .ZN(new_n25203_));
  INV_X1     g25136(.I(new_n25057_), .ZN(new_n25204_));
  OAI21_X1   g25137(.A1(new_n25201_), .A2(new_n25200_), .B(new_n25062_), .ZN(new_n25205_));
  NAND3_X1   g25138(.A1(new_n25192_), .A2(new_n25063_), .A3(new_n25198_), .ZN(new_n25206_));
  NAND3_X1   g25139(.A1(new_n25205_), .A2(new_n25206_), .A3(new_n25204_), .ZN(new_n25207_));
  NAND2_X1   g25140(.A1(new_n25203_), .A2(new_n25207_), .ZN(new_n25208_));
  XOR2_X1    g25141(.A1(new_n25208_), .A2(new_n25052_), .Z(new_n25209_));
  NAND3_X1   g25142(.A1(new_n25037_), .A2(new_n25038_), .A3(new_n25039_), .ZN(new_n25210_));
  NAND2_X1   g25143(.A1(new_n25210_), .A2(new_n25040_), .ZN(new_n25211_));
  INV_X1     g25144(.I(new_n25211_), .ZN(new_n25212_));
  XOR2_X1    g25145(.A1(new_n25209_), .A2(new_n25212_), .Z(new_n25213_));
  NAND2_X1   g25146(.A1(new_n24850_), .A2(new_n24849_), .ZN(new_n25214_));
  NOR2_X1    g25147(.A1(new_n24793_), .A2(new_n24798_), .ZN(new_n25215_));
  AOI21_X1   g25148(.A1(new_n25214_), .A2(new_n24800_), .B(new_n25215_), .ZN(new_n25216_));
  NOR2_X1    g25149(.A1(new_n25032_), .A2(new_n25033_), .ZN(new_n25217_));
  NOR3_X1    g25150(.A1(new_n25028_), .A2(new_n25030_), .A3(new_n25031_), .ZN(new_n25218_));
  NOR2_X1    g25151(.A1(new_n25217_), .A2(new_n25218_), .ZN(new_n25219_));
  AOI21_X1   g25152(.A1(new_n25037_), .A2(new_n25038_), .B(new_n25219_), .ZN(new_n25220_));
  NOR2_X1    g25153(.A1(new_n25023_), .A2(new_n25033_), .ZN(new_n25221_));
  NOR2_X1    g25154(.A1(new_n25032_), .A2(new_n25028_), .ZN(new_n25222_));
  NOR2_X1    g25155(.A1(new_n25222_), .A2(new_n25221_), .ZN(new_n25223_));
  NOR3_X1    g25156(.A1(new_n25008_), .A2(new_n25014_), .A3(new_n25223_), .ZN(new_n25224_));
  OAI21_X1   g25157(.A1(new_n25224_), .A2(new_n25220_), .B(new_n25216_), .ZN(new_n25225_));
  NAND3_X1   g25158(.A1(new_n25036_), .A2(new_n25042_), .A3(new_n24851_), .ZN(new_n25226_));
  NAND2_X1   g25159(.A1(new_n25225_), .A2(new_n25226_), .ZN(new_n25227_));
  NOR2_X1    g25160(.A1(new_n25043_), .A2(new_n25216_), .ZN(new_n25228_));
  AOI21_X1   g25161(.A1(new_n25227_), .A2(new_n25044_), .B(new_n25228_), .ZN(new_n25229_));
  NOR4_X1    g25162(.A1(new_n24635_), .A2(new_n24627_), .A3(new_n24843_), .A4(new_n25046_), .ZN(new_n25230_));
  XOR2_X1    g25163(.A1(new_n25230_), .A2(new_n25229_), .Z(new_n25231_));
  XOR2_X1    g25164(.A1(new_n25231_), .A2(new_n25213_), .Z(\result[7] ));
  INV_X1     g25165(.I(new_n25046_), .ZN(new_n25233_));
  INV_X1     g25166(.I(new_n24842_), .ZN(new_n25234_));
  AOI21_X1   g25167(.A1(new_n24809_), .A2(new_n24810_), .B(new_n24805_), .ZN(new_n25235_));
  NOR3_X1    g25168(.A1(new_n24801_), .A2(new_n24793_), .A3(new_n24803_), .ZN(new_n25236_));
  OAI21_X1   g25169(.A1(new_n25236_), .A2(new_n25235_), .B(new_n24840_), .ZN(new_n25237_));
  NAND2_X1   g25170(.A1(new_n25237_), .A2(new_n25234_), .ZN(new_n25238_));
  AOI22_X1   g25171(.A1(new_n25238_), .A2(new_n25043_), .B1(new_n25225_), .B2(new_n25226_), .ZN(new_n25239_));
  XOR2_X1    g25172(.A1(new_n25213_), .A2(new_n25239_), .Z(new_n25240_));
  NAND4_X1   g25173(.A1(new_n24628_), .A2(new_n24844_), .A3(new_n25233_), .A4(new_n25240_), .ZN(new_n25241_));
  AOI21_X1   g25174(.A1(new_n25205_), .A2(new_n25206_), .B(new_n25204_), .ZN(new_n25242_));
  NOR3_X1    g25175(.A1(new_n25202_), .A2(new_n25199_), .A3(new_n25057_), .ZN(new_n25243_));
  OAI21_X1   g25176(.A1(new_n25243_), .A2(new_n25242_), .B(new_n25052_), .ZN(new_n25244_));
  AOI22_X1   g25177(.A1(new_n24620_), .A2(new_n8799_), .B1(new_n6846_), .B2(new_n24386_), .ZN(new_n25245_));
  NOR2_X1    g25178(.A1(new_n24835_), .A2(new_n6839_), .ZN(new_n25246_));
  OAI21_X1   g25179(.A1(new_n25246_), .A2(new_n25245_), .B(new_n6835_), .ZN(new_n25247_));
  NOR3_X1    g25180(.A1(new_n24831_), .A2(new_n24832_), .A3(new_n25247_), .ZN(new_n25248_));
  XOR2_X1    g25181(.A1(new_n25248_), .A2(\a[5] ), .Z(new_n25249_));
  NOR2_X1    g25182(.A1(new_n24171_), .A2(new_n24174_), .ZN(new_n25250_));
  OAI21_X1   g25183(.A1(new_n22117_), .A2(new_n22118_), .B(new_n22150_), .ZN(new_n25251_));
  OAI21_X1   g25184(.A1(new_n22159_), .A2(new_n22115_), .B(new_n22149_), .ZN(new_n25252_));
  NAND2_X1   g25185(.A1(new_n25251_), .A2(new_n25252_), .ZN(new_n25253_));
  AOI21_X1   g25186(.A1(new_n25253_), .A2(new_n24168_), .B(new_n24167_), .ZN(new_n25254_));
  OAI22_X1   g25187(.A1(new_n23948_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n22149_), .ZN(new_n25255_));
  NAND2_X1   g25188(.A1(new_n24174_), .A2(new_n6784_), .ZN(new_n25256_));
  AOI21_X1   g25189(.A1(new_n25256_), .A2(new_n25255_), .B(new_n6776_), .ZN(new_n25257_));
  OAI21_X1   g25190(.A1(new_n25250_), .A2(new_n25254_), .B(new_n25257_), .ZN(new_n25258_));
  XOR2_X1    g25191(.A1(new_n25258_), .A2(new_n4009_), .Z(new_n25259_));
  AOI22_X1   g25192(.A1(new_n22048_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n21953_), .ZN(new_n25260_));
  AOI21_X1   g25193(.A1(new_n22118_), .A2(new_n4709_), .B(new_n25260_), .ZN(new_n25261_));
  NOR4_X1    g25194(.A1(new_n23672_), .A2(new_n4707_), .A3(new_n23673_), .A4(new_n25261_), .ZN(new_n25262_));
  XOR2_X1    g25195(.A1(new_n25262_), .A2(new_n4034_), .Z(new_n25263_));
  NOR2_X1    g25196(.A1(new_n25173_), .A2(new_n25069_), .ZN(new_n25264_));
  XOR2_X1    g25197(.A1(new_n25075_), .A2(new_n25171_), .Z(new_n25265_));
  AOI21_X1   g25198(.A1(new_n25173_), .A2(new_n25069_), .B(new_n25265_), .ZN(new_n25266_));
  NOR2_X1    g25199(.A1(new_n25266_), .A2(new_n25264_), .ZN(new_n25267_));
  NAND3_X1   g25200(.A1(new_n19516_), .A2(new_n19519_), .A3(new_n19512_), .ZN(new_n25268_));
  OAI21_X1   g25201(.A1(new_n19487_), .A2(new_n19508_), .B(new_n17770_), .ZN(new_n25269_));
  OAI22_X1   g25202(.A1(new_n19522_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n17775_), .ZN(new_n25270_));
  OAI21_X1   g25203(.A1(new_n19511_), .A2(new_n19510_), .B(new_n6090_), .ZN(new_n25271_));
  AOI21_X1   g25204(.A1(new_n25270_), .A2(new_n25271_), .B(new_n6082_), .ZN(new_n25272_));
  NAND3_X1   g25205(.A1(new_n25269_), .A2(new_n25272_), .A3(new_n25268_), .ZN(new_n25273_));
  XOR2_X1    g25206(.A1(new_n25273_), .A2(new_n3521_), .Z(new_n25274_));
  OAI22_X1   g25207(.A1(new_n19463_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19437_), .ZN(new_n25275_));
  NAND2_X1   g25208(.A1(new_n17780_), .A2(new_n4469_), .ZN(new_n25276_));
  AOI21_X1   g25209(.A1(new_n25275_), .A2(new_n25276_), .B(new_n4468_), .ZN(new_n25277_));
  NAND3_X1   g25210(.A1(new_n21730_), .A2(new_n21729_), .A3(new_n25277_), .ZN(new_n25278_));
  XOR2_X1    g25211(.A1(new_n25278_), .A2(\a[17] ), .Z(new_n25279_));
  OAI22_X1   g25212(.A1(new_n19428_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19423_), .ZN(new_n25280_));
  NAND2_X1   g25213(.A1(new_n19438_), .A2(new_n4096_), .ZN(new_n25281_));
  AOI21_X1   g25214(.A1(new_n25281_), .A2(new_n25280_), .B(new_n4095_), .ZN(new_n25282_));
  NAND2_X1   g25215(.A1(new_n20907_), .A2(new_n25282_), .ZN(new_n25283_));
  XOR2_X1    g25216(.A1(new_n25283_), .A2(\a[20] ), .Z(new_n25284_));
  NOR2_X1    g25217(.A1(new_n25155_), .A2(new_n25092_), .ZN(new_n25285_));
  AOI21_X1   g25218(.A1(new_n25155_), .A2(new_n25092_), .B(new_n25137_), .ZN(new_n25286_));
  NOR2_X1    g25219(.A1(new_n25286_), .A2(new_n25285_), .ZN(new_n25287_));
  INV_X1     g25220(.I(new_n25287_), .ZN(new_n25288_));
  AOI22_X1   g25221(.A1(new_n19415_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n19407_), .ZN(new_n25289_));
  NOR2_X1    g25222(.A1(new_n17787_), .A2(new_n3780_), .ZN(new_n25290_));
  OAI21_X1   g25223(.A1(new_n25290_), .A2(new_n25289_), .B(new_n3301_), .ZN(new_n25291_));
  INV_X1     g25224(.I(new_n25291_), .ZN(new_n25292_));
  NAND3_X1   g25225(.A1(new_n20827_), .A2(new_n84_), .A3(new_n25292_), .ZN(new_n25293_));
  NAND2_X1   g25226(.A1(new_n20949_), .A2(new_n20824_), .ZN(new_n25294_));
  OAI21_X1   g25227(.A1(new_n25294_), .A2(new_n25291_), .B(\a[23] ), .ZN(new_n25295_));
  NAND2_X1   g25228(.A1(new_n25295_), .A2(new_n25293_), .ZN(new_n25296_));
  INV_X1     g25229(.I(new_n25296_), .ZN(new_n25297_));
  OAI22_X1   g25230(.A1(new_n19400_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19393_), .ZN(new_n25298_));
  NAND2_X1   g25231(.A1(new_n17790_), .A2(new_n3317_), .ZN(new_n25299_));
  AOI21_X1   g25232(.A1(new_n25299_), .A2(new_n25298_), .B(new_n3260_), .ZN(new_n25300_));
  NAND3_X1   g25233(.A1(new_n20251_), .A2(new_n72_), .A3(new_n25300_), .ZN(new_n25301_));
  NAND2_X1   g25234(.A1(new_n20251_), .A2(new_n25300_), .ZN(new_n25302_));
  NAND2_X1   g25235(.A1(new_n25302_), .A2(\a[26] ), .ZN(new_n25303_));
  NAND2_X1   g25236(.A1(new_n25303_), .A2(new_n25301_), .ZN(new_n25304_));
  AOI22_X1   g25237(.A1(new_n19386_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n20127_), .ZN(new_n25305_));
  NOR2_X1    g25238(.A1(new_n17793_), .A2(new_n3175_), .ZN(new_n25306_));
  OAI21_X1   g25239(.A1(new_n25305_), .A2(new_n25306_), .B(new_n2736_), .ZN(new_n25307_));
  NOR3_X1    g25240(.A1(new_n21632_), .A2(\a[29] ), .A3(new_n25307_), .ZN(new_n25308_));
  OAI21_X1   g25241(.A1(new_n21632_), .A2(new_n25307_), .B(\a[29] ), .ZN(new_n25309_));
  INV_X1     g25242(.I(new_n25309_), .ZN(new_n25310_));
  NOR2_X1    g25243(.A1(new_n25310_), .A2(new_n25308_), .ZN(new_n25311_));
  INV_X1     g25244(.I(new_n25311_), .ZN(new_n25312_));
  INV_X1     g25245(.I(new_n25113_), .ZN(new_n25313_));
  OR2_X2     g25246(.A1(new_n25093_), .A2(new_n25094_), .Z(new_n25314_));
  OAI21_X1   g25247(.A1(new_n25102_), .A2(new_n25111_), .B(new_n25314_), .ZN(new_n25315_));
  NOR4_X1    g25248(.A1(new_n573_), .A2(new_n791_), .A3(new_n703_), .A4(new_n561_), .ZN(new_n25316_));
  NOR2_X1    g25249(.A1(new_n286_), .A2(new_n163_), .ZN(new_n25317_));
  INV_X1     g25250(.I(new_n25317_), .ZN(new_n25318_));
  NOR4_X1    g25251(.A1(new_n19789_), .A2(new_n1784_), .A3(new_n25316_), .A4(new_n25318_), .ZN(new_n25319_));
  NOR4_X1    g25252(.A1(new_n23979_), .A2(new_n2480_), .A3(new_n3938_), .A4(new_n1914_), .ZN(new_n25320_));
  NOR4_X1    g25253(.A1(new_n3213_), .A2(new_n1339_), .A3(new_n2232_), .A4(new_n1858_), .ZN(new_n25321_));
  NOR2_X1    g25254(.A1(new_n304_), .A2(new_n398_), .ZN(new_n25322_));
  NAND4_X1   g25255(.A1(new_n11727_), .A2(new_n25322_), .A3(new_n545_), .A4(new_n628_), .ZN(new_n25323_));
  NOR2_X1    g25256(.A1(new_n1293_), .A2(new_n25323_), .ZN(new_n25324_));
  NAND4_X1   g25257(.A1(new_n25324_), .A2(new_n25319_), .A3(new_n25320_), .A4(new_n25321_), .ZN(new_n25325_));
  NOR3_X1    g25258(.A1(new_n12506_), .A2(new_n12861_), .A3(new_n25325_), .ZN(new_n25326_));
  NOR2_X1    g25259(.A1(new_n25314_), .A2(new_n25326_), .ZN(new_n25327_));
  INV_X1     g25260(.I(new_n25326_), .ZN(new_n25328_));
  NOR2_X1    g25261(.A1(new_n25095_), .A2(new_n25328_), .ZN(new_n25329_));
  NOR2_X1    g25262(.A1(new_n25327_), .A2(new_n25329_), .ZN(new_n25330_));
  AOI21_X1   g25263(.A1(new_n25313_), .A2(new_n25315_), .B(new_n25330_), .ZN(new_n25331_));
  NAND2_X1   g25264(.A1(new_n25315_), .A2(new_n25313_), .ZN(new_n25332_));
  XOR2_X1    g25265(.A1(new_n25095_), .A2(new_n25326_), .Z(new_n25333_));
  NOR2_X1    g25266(.A1(new_n25332_), .A2(new_n25333_), .ZN(new_n25334_));
  NAND2_X1   g25267(.A1(new_n17798_), .A2(new_n3332_), .ZN(new_n25335_));
  OAI21_X1   g25268(.A1(new_n19364_), .A2(new_n2771_), .B(new_n2763_), .ZN(new_n25336_));
  AOI21_X1   g25269(.A1(new_n17802_), .A2(new_n3189_), .B(new_n25336_), .ZN(new_n25337_));
  NAND3_X1   g25270(.A1(new_n21454_), .A2(new_n25335_), .A3(new_n25337_), .ZN(new_n25338_));
  INV_X1     g25271(.I(new_n25338_), .ZN(new_n25339_));
  NOR3_X1    g25272(.A1(new_n25331_), .A2(new_n25334_), .A3(new_n25339_), .ZN(new_n25340_));
  OAI21_X1   g25273(.A1(new_n25331_), .A2(new_n25334_), .B(new_n25339_), .ZN(new_n25341_));
  INV_X1     g25274(.I(new_n25341_), .ZN(new_n25342_));
  NOR2_X1    g25275(.A1(new_n25342_), .A2(new_n25340_), .ZN(new_n25343_));
  NOR2_X1    g25276(.A1(new_n25131_), .A2(new_n25133_), .ZN(new_n25344_));
  OAI21_X1   g25277(.A1(new_n25344_), .A2(new_n25135_), .B(new_n25343_), .ZN(new_n25345_));
  INV_X1     g25278(.I(new_n25331_), .ZN(new_n25346_));
  INV_X1     g25279(.I(new_n25334_), .ZN(new_n25347_));
  NAND3_X1   g25280(.A1(new_n25346_), .A2(new_n25347_), .A3(new_n25338_), .ZN(new_n25348_));
  NAND2_X1   g25281(.A1(new_n25348_), .A2(new_n25341_), .ZN(new_n25349_));
  NOR2_X1    g25282(.A1(new_n25344_), .A2(new_n25135_), .ZN(new_n25350_));
  NAND2_X1   g25283(.A1(new_n25350_), .A2(new_n25349_), .ZN(new_n25351_));
  AOI21_X1   g25284(.A1(new_n25345_), .A2(new_n25351_), .B(new_n25312_), .ZN(new_n25352_));
  NOR2_X1    g25285(.A1(new_n25350_), .A2(new_n25349_), .ZN(new_n25353_));
  NOR3_X1    g25286(.A1(new_n25343_), .A2(new_n25344_), .A3(new_n25135_), .ZN(new_n25354_));
  NOR3_X1    g25287(.A1(new_n25353_), .A2(new_n25354_), .A3(new_n25311_), .ZN(new_n25355_));
  NOR2_X1    g25288(.A1(new_n25352_), .A2(new_n25355_), .ZN(new_n25356_));
  NOR2_X1    g25289(.A1(new_n25356_), .A2(new_n25304_), .ZN(new_n25357_));
  INV_X1     g25290(.I(new_n25304_), .ZN(new_n25358_));
  OAI21_X1   g25291(.A1(new_n25353_), .A2(new_n25354_), .B(new_n25311_), .ZN(new_n25359_));
  NAND3_X1   g25292(.A1(new_n25345_), .A2(new_n25351_), .A3(new_n25312_), .ZN(new_n25360_));
  NAND2_X1   g25293(.A1(new_n25360_), .A2(new_n25359_), .ZN(new_n25361_));
  NOR2_X1    g25294(.A1(new_n25358_), .A2(new_n25361_), .ZN(new_n25362_));
  NOR4_X1    g25295(.A1(new_n25167_), .A2(new_n25362_), .A3(new_n25357_), .A4(new_n25087_), .ZN(new_n25363_));
  NAND2_X1   g25296(.A1(new_n25358_), .A2(new_n25361_), .ZN(new_n25364_));
  NAND2_X1   g25297(.A1(new_n25356_), .A2(new_n25304_), .ZN(new_n25365_));
  AOI22_X1   g25298(.A1(new_n25162_), .A2(new_n25164_), .B1(new_n25364_), .B2(new_n25365_), .ZN(new_n25366_));
  OAI21_X1   g25299(.A1(new_n25366_), .A2(new_n25363_), .B(new_n25297_), .ZN(new_n25367_));
  NAND4_X1   g25300(.A1(new_n25162_), .A2(new_n25364_), .A3(new_n25365_), .A4(new_n25164_), .ZN(new_n25368_));
  OAI22_X1   g25301(.A1(new_n25167_), .A2(new_n25087_), .B1(new_n25362_), .B2(new_n25357_), .ZN(new_n25369_));
  NAND3_X1   g25302(.A1(new_n25369_), .A2(new_n25368_), .A3(new_n25296_), .ZN(new_n25370_));
  AOI21_X1   g25303(.A1(new_n25367_), .A2(new_n25370_), .B(new_n25288_), .ZN(new_n25371_));
  AOI21_X1   g25304(.A1(new_n25369_), .A2(new_n25368_), .B(new_n25296_), .ZN(new_n25372_));
  NOR3_X1    g25305(.A1(new_n25366_), .A2(new_n25363_), .A3(new_n25297_), .ZN(new_n25373_));
  NOR3_X1    g25306(.A1(new_n25373_), .A2(new_n25372_), .A3(new_n25287_), .ZN(new_n25374_));
  AOI22_X1   g25307(.A1(new_n25081_), .A2(new_n25079_), .B1(new_n25163_), .B2(new_n25168_), .ZN(new_n25375_));
  INV_X1     g25308(.I(new_n25375_), .ZN(new_n25376_));
  NOR3_X1    g25309(.A1(new_n25374_), .A2(new_n25371_), .A3(new_n25376_), .ZN(new_n25377_));
  OAI21_X1   g25310(.A1(new_n25373_), .A2(new_n25372_), .B(new_n25287_), .ZN(new_n25378_));
  NAND3_X1   g25311(.A1(new_n25367_), .A2(new_n25370_), .A3(new_n25288_), .ZN(new_n25379_));
  AOI21_X1   g25312(.A1(new_n25378_), .A2(new_n25379_), .B(new_n25375_), .ZN(new_n25380_));
  OAI21_X1   g25313(.A1(new_n25377_), .A2(new_n25380_), .B(new_n25284_), .ZN(new_n25381_));
  XOR2_X1    g25314(.A1(new_n25283_), .A2(new_n3035_), .Z(new_n25382_));
  NAND3_X1   g25315(.A1(new_n25378_), .A2(new_n25379_), .A3(new_n25375_), .ZN(new_n25383_));
  OAI21_X1   g25316(.A1(new_n25374_), .A2(new_n25371_), .B(new_n25376_), .ZN(new_n25384_));
  NAND3_X1   g25317(.A1(new_n25384_), .A2(new_n25383_), .A3(new_n25382_), .ZN(new_n25385_));
  NAND2_X1   g25318(.A1(new_n25381_), .A2(new_n25385_), .ZN(new_n25386_));
  NAND2_X1   g25319(.A1(new_n25386_), .A2(new_n25279_), .ZN(new_n25387_));
  XOR2_X1    g25320(.A1(new_n25278_), .A2(new_n3372_), .Z(new_n25388_));
  NAND3_X1   g25321(.A1(new_n25388_), .A2(new_n25381_), .A3(new_n25385_), .ZN(new_n25389_));
  NOR2_X1    g25322(.A1(new_n25075_), .A2(new_n25170_), .ZN(new_n25390_));
  NAND3_X1   g25323(.A1(new_n25387_), .A2(new_n25389_), .A3(new_n25390_), .ZN(new_n25391_));
  AOI21_X1   g25324(.A1(new_n25381_), .A2(new_n25385_), .B(new_n25388_), .ZN(new_n25392_));
  NOR2_X1    g25325(.A1(new_n25386_), .A2(new_n25279_), .ZN(new_n25393_));
  INV_X1     g25326(.I(new_n25390_), .ZN(new_n25394_));
  OAI21_X1   g25327(.A1(new_n25392_), .A2(new_n25393_), .B(new_n25394_), .ZN(new_n25395_));
  AOI21_X1   g25328(.A1(new_n25395_), .A2(new_n25391_), .B(new_n25274_), .ZN(new_n25396_));
  XOR2_X1    g25329(.A1(new_n25273_), .A2(\a[14] ), .Z(new_n25397_));
  NOR3_X1    g25330(.A1(new_n25392_), .A2(new_n25393_), .A3(new_n25394_), .ZN(new_n25398_));
  AOI21_X1   g25331(.A1(new_n25387_), .A2(new_n25389_), .B(new_n25390_), .ZN(new_n25399_));
  NOR3_X1    g25332(.A1(new_n25398_), .A2(new_n25399_), .A3(new_n25397_), .ZN(new_n25400_));
  NOR2_X1    g25333(.A1(new_n25400_), .A2(new_n25396_), .ZN(new_n25401_));
  XOR2_X1    g25334(.A1(new_n25401_), .A2(new_n25267_), .Z(new_n25402_));
  NOR3_X1    g25335(.A1(new_n25402_), .A2(new_n25189_), .A3(new_n25062_), .ZN(new_n25403_));
  NOR3_X1    g25336(.A1(new_n25401_), .A2(new_n25264_), .A3(new_n25266_), .ZN(new_n25404_));
  NOR3_X1    g25337(.A1(new_n25267_), .A2(new_n25396_), .A3(new_n25400_), .ZN(new_n25405_));
  NOR2_X1    g25338(.A1(new_n25404_), .A2(new_n25405_), .ZN(new_n25406_));
  AOI21_X1   g25339(.A1(new_n25195_), .A2(new_n25063_), .B(new_n25406_), .ZN(new_n25407_));
  OAI21_X1   g25340(.A1(new_n25403_), .A2(new_n25407_), .B(new_n25263_), .ZN(new_n25408_));
  XOR2_X1    g25341(.A1(new_n25262_), .A2(\a[11] ), .Z(new_n25409_));
  NAND3_X1   g25342(.A1(new_n25195_), .A2(new_n25406_), .A3(new_n25063_), .ZN(new_n25410_));
  OAI21_X1   g25343(.A1(new_n25189_), .A2(new_n25062_), .B(new_n25402_), .ZN(new_n25411_));
  NAND3_X1   g25344(.A1(new_n25411_), .A2(new_n25410_), .A3(new_n25409_), .ZN(new_n25412_));
  AOI21_X1   g25345(.A1(new_n25408_), .A2(new_n25412_), .B(new_n25259_), .ZN(new_n25413_));
  XOR2_X1    g25346(.A1(new_n25258_), .A2(\a[8] ), .Z(new_n25414_));
  AOI21_X1   g25347(.A1(new_n25411_), .A2(new_n25410_), .B(new_n25409_), .ZN(new_n25415_));
  NOR3_X1    g25348(.A1(new_n25403_), .A2(new_n25407_), .A3(new_n25263_), .ZN(new_n25416_));
  NOR3_X1    g25349(.A1(new_n25416_), .A2(new_n25415_), .A3(new_n25414_), .ZN(new_n25417_));
  NOR2_X1    g25350(.A1(new_n25417_), .A2(new_n25413_), .ZN(new_n25418_));
  XOR2_X1    g25351(.A1(new_n25195_), .A2(new_n25062_), .Z(new_n25419_));
  AOI21_X1   g25352(.A1(new_n25197_), .A2(new_n25057_), .B(new_n25419_), .ZN(new_n25420_));
  NOR2_X1    g25353(.A1(new_n25197_), .A2(new_n25057_), .ZN(new_n25421_));
  OAI21_X1   g25354(.A1(new_n25420_), .A2(new_n25421_), .B(new_n25418_), .ZN(new_n25422_));
  OAI21_X1   g25355(.A1(new_n25415_), .A2(new_n25416_), .B(new_n25414_), .ZN(new_n25423_));
  NAND3_X1   g25356(.A1(new_n25408_), .A2(new_n25412_), .A3(new_n25259_), .ZN(new_n25424_));
  NAND2_X1   g25357(.A1(new_n25423_), .A2(new_n25424_), .ZN(new_n25425_));
  NOR2_X1    g25358(.A1(new_n25420_), .A2(new_n25421_), .ZN(new_n25426_));
  NAND2_X1   g25359(.A1(new_n25425_), .A2(new_n25426_), .ZN(new_n25427_));
  AOI21_X1   g25360(.A1(new_n25422_), .A2(new_n25427_), .B(new_n25249_), .ZN(new_n25428_));
  NOR4_X1    g25361(.A1(new_n24831_), .A2(new_n24832_), .A3(\a[5] ), .A4(new_n25247_), .ZN(new_n25429_));
  NOR2_X1    g25362(.A1(new_n25248_), .A2(new_n65_), .ZN(new_n25430_));
  NOR2_X1    g25363(.A1(new_n25430_), .A2(new_n25429_), .ZN(new_n25431_));
  NOR2_X1    g25364(.A1(new_n25425_), .A2(new_n25426_), .ZN(new_n25432_));
  NOR3_X1    g25365(.A1(new_n25418_), .A2(new_n25420_), .A3(new_n25421_), .ZN(new_n25433_));
  NOR3_X1    g25366(.A1(new_n25433_), .A2(new_n25432_), .A3(new_n25431_), .ZN(new_n25434_));
  OAI21_X1   g25367(.A1(new_n25428_), .A2(new_n25434_), .B(new_n25244_), .ZN(new_n25435_));
  OAI21_X1   g25368(.A1(new_n25433_), .A2(new_n25432_), .B(new_n25431_), .ZN(new_n25436_));
  NAND3_X1   g25369(.A1(new_n25422_), .A2(new_n25249_), .A3(new_n25427_), .ZN(new_n25437_));
  NAND4_X1   g25370(.A1(new_n25208_), .A2(new_n25437_), .A3(new_n25436_), .A4(new_n25052_), .ZN(new_n25438_));
  NAND2_X1   g25371(.A1(new_n25435_), .A2(new_n25438_), .ZN(new_n25439_));
  XNOR2_X1   g25372(.A1(new_n25208_), .A2(new_n25052_), .ZN(new_n25440_));
  NOR2_X1    g25373(.A1(new_n25229_), .A2(new_n25440_), .ZN(new_n25441_));
  XOR2_X1    g25374(.A1(new_n25441_), .A2(new_n25439_), .Z(new_n25442_));
  XOR2_X1    g25375(.A1(new_n25229_), .A2(new_n25440_), .Z(new_n25443_));
  NAND2_X1   g25376(.A1(new_n25443_), .A2(new_n25211_), .ZN(new_n25444_));
  XOR2_X1    g25377(.A1(new_n25442_), .A2(new_n25444_), .Z(new_n25445_));
  XOR2_X1    g25378(.A1(new_n25241_), .A2(new_n25445_), .Z(\result[8] ));
  NOR2_X1    g25379(.A1(new_n25241_), .A2(new_n25445_), .ZN(new_n25447_));
  NAND3_X1   g25380(.A1(new_n25435_), .A2(new_n25211_), .A3(new_n25438_), .ZN(new_n25448_));
  NAND3_X1   g25381(.A1(new_n25239_), .A2(new_n25209_), .A3(new_n25448_), .ZN(new_n25449_));
  NAND2_X1   g25382(.A1(new_n25249_), .A2(new_n25426_), .ZN(new_n25450_));
  OAI21_X1   g25383(.A1(new_n25420_), .A2(new_n25421_), .B(new_n25431_), .ZN(new_n25451_));
  NAND3_X1   g25384(.A1(new_n25450_), .A2(new_n25451_), .A3(new_n25425_), .ZN(new_n25452_));
  NOR3_X1    g25385(.A1(new_n25431_), .A2(new_n25420_), .A3(new_n25421_), .ZN(new_n25453_));
  NOR2_X1    g25386(.A1(new_n25249_), .A2(new_n25426_), .ZN(new_n25454_));
  OAI21_X1   g25387(.A1(new_n25454_), .A2(new_n25453_), .B(new_n25418_), .ZN(new_n25455_));
  NAND3_X1   g25388(.A1(new_n25452_), .A2(new_n25455_), .A3(new_n25244_), .ZN(new_n25456_));
  INV_X1     g25389(.I(new_n25456_), .ZN(new_n25457_));
  OAI22_X1   g25390(.A1(new_n24167_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n23948_), .ZN(new_n25458_));
  NAND2_X1   g25391(.A1(new_n24386_), .A2(new_n6784_), .ZN(new_n25459_));
  AOI21_X1   g25392(.A1(new_n25459_), .A2(new_n25458_), .B(new_n6776_), .ZN(new_n25460_));
  NAND2_X1   g25393(.A1(new_n24390_), .A2(new_n25460_), .ZN(new_n25461_));
  XOR2_X1    g25394(.A1(new_n25461_), .A2(new_n4009_), .Z(new_n25462_));
  OAI22_X1   g25395(.A1(new_n22115_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n22051_), .ZN(new_n25463_));
  NAND2_X1   g25396(.A1(new_n22150_), .A2(new_n4709_), .ZN(new_n25464_));
  AOI21_X1   g25397(.A1(new_n25463_), .A2(new_n25464_), .B(new_n4707_), .ZN(new_n25465_));
  NAND2_X1   g25398(.A1(new_n22163_), .A2(new_n25465_), .ZN(new_n25466_));
  XOR2_X1    g25399(.A1(new_n25466_), .A2(\a[11] ), .Z(new_n25467_));
  NAND2_X1   g25400(.A1(new_n25388_), .A2(new_n25375_), .ZN(new_n25468_));
  NAND2_X1   g25401(.A1(new_n25378_), .A2(new_n25379_), .ZN(new_n25469_));
  XOR2_X1    g25402(.A1(new_n25469_), .A2(new_n25382_), .Z(new_n25470_));
  OAI21_X1   g25403(.A1(new_n25388_), .A2(new_n25375_), .B(new_n25470_), .ZN(new_n25471_));
  NAND2_X1   g25404(.A1(new_n25471_), .A2(new_n25468_), .ZN(new_n25472_));
  INV_X1     g25405(.I(new_n25472_), .ZN(new_n25473_));
  OAI22_X1   g25406(.A1(new_n19512_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n19522_), .ZN(new_n25474_));
  OAI21_X1   g25407(.A1(new_n6091_), .A2(new_n21960_), .B(new_n25474_), .ZN(new_n25475_));
  NAND3_X1   g25408(.A1(new_n21963_), .A2(new_n6081_), .A3(new_n25475_), .ZN(new_n25476_));
  XOR2_X1    g25409(.A1(new_n25476_), .A2(new_n3521_), .Z(new_n25477_));
  OAI22_X1   g25410(.A1(new_n19475_), .A2(new_n4297_), .B1(new_n19463_), .B2(new_n4291_), .ZN(new_n25478_));
  NAND2_X1   g25411(.A1(new_n19484_), .A2(new_n4469_), .ZN(new_n25479_));
  AOI21_X1   g25412(.A1(new_n25479_), .A2(new_n25478_), .B(new_n4468_), .ZN(new_n25480_));
  NAND2_X1   g25413(.A1(new_n21171_), .A2(new_n25480_), .ZN(new_n25481_));
  XOR2_X1    g25414(.A1(new_n25481_), .A2(\a[17] ), .Z(new_n25482_));
  INV_X1     g25415(.I(new_n25482_), .ZN(new_n25483_));
  OAI22_X1   g25416(.A1(new_n17784_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19428_), .ZN(new_n25484_));
  NAND2_X1   g25417(.A1(new_n19466_), .A2(new_n4096_), .ZN(new_n25485_));
  AOI21_X1   g25418(.A1(new_n25485_), .A2(new_n25484_), .B(new_n4095_), .ZN(new_n25486_));
  NAND2_X1   g25419(.A1(new_n21100_), .A2(new_n25486_), .ZN(new_n25487_));
  XOR2_X1    g25420(.A1(new_n25487_), .A2(\a[20] ), .Z(new_n25488_));
  OAI22_X1   g25421(.A1(new_n17789_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19400_), .ZN(new_n25489_));
  NAND2_X1   g25422(.A1(new_n19407_), .A2(new_n3317_), .ZN(new_n25490_));
  AOI21_X1   g25423(.A1(new_n25490_), .A2(new_n25489_), .B(new_n3260_), .ZN(new_n25491_));
  NAND2_X1   g25424(.A1(new_n20864_), .A2(new_n25491_), .ZN(new_n25492_));
  XOR2_X1    g25425(.A1(new_n25492_), .A2(\a[26] ), .Z(new_n25493_));
  AOI22_X1   g25426(.A1(new_n19386_), .A2(new_n2746_), .B1(new_n3275_), .B2(new_n17794_), .ZN(new_n25494_));
  NOR2_X1    g25427(.A1(new_n19393_), .A2(new_n3175_), .ZN(new_n25495_));
  OAI21_X1   g25428(.A1(new_n25494_), .A2(new_n25495_), .B(new_n2736_), .ZN(new_n25496_));
  NOR2_X1    g25429(.A1(new_n20291_), .A2(new_n25496_), .ZN(new_n25497_));
  XOR2_X1    g25430(.A1(new_n25497_), .A2(new_n74_), .Z(new_n25498_));
  INV_X1     g25431(.I(new_n25498_), .ZN(new_n25499_));
  NAND2_X1   g25432(.A1(new_n20127_), .A2(new_n3332_), .ZN(new_n25500_));
  NAND2_X1   g25433(.A1(new_n17798_), .A2(new_n3189_), .ZN(new_n25501_));
  AOI21_X1   g25434(.A1(new_n17802_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n25502_));
  NAND4_X1   g25435(.A1(new_n21753_), .A2(new_n25500_), .A3(new_n25501_), .A4(new_n25502_), .ZN(new_n25503_));
  INV_X1     g25436(.I(new_n25503_), .ZN(new_n25504_));
  INV_X1     g25437(.I(new_n2840_), .ZN(new_n25505_));
  NAND4_X1   g25438(.A1(new_n1565_), .A2(new_n1263_), .A3(new_n537_), .A4(new_n1321_), .ZN(new_n25506_));
  NOR3_X1    g25439(.A1(new_n25505_), .A2(new_n11840_), .A3(new_n25506_), .ZN(new_n25507_));
  NAND3_X1   g25440(.A1(new_n1658_), .A2(new_n1796_), .A3(new_n187_), .ZN(new_n25508_));
  NAND2_X1   g25441(.A1(new_n358_), .A2(new_n231_), .ZN(new_n25509_));
  NOR4_X1    g25442(.A1(new_n11926_), .A2(new_n1788_), .A3(new_n25508_), .A4(new_n25509_), .ZN(new_n25510_));
  NAND4_X1   g25443(.A1(new_n25507_), .A2(new_n1006_), .A3(new_n3931_), .A4(new_n25510_), .ZN(new_n25511_));
  NOR3_X1    g25444(.A1(new_n1052_), .A2(new_n25511_), .A3(new_n2085_), .ZN(new_n25512_));
  INV_X1     g25445(.I(new_n25329_), .ZN(new_n25513_));
  OAI21_X1   g25446(.A1(new_n25314_), .A2(new_n25326_), .B(new_n25332_), .ZN(new_n25514_));
  NAND3_X1   g25447(.A1(new_n25514_), .A2(new_n25314_), .A3(new_n25513_), .ZN(new_n25515_));
  NAND3_X1   g25448(.A1(new_n25332_), .A2(new_n25095_), .A3(new_n25326_), .ZN(new_n25516_));
  AOI21_X1   g25449(.A1(new_n25515_), .A2(new_n25516_), .B(new_n25512_), .ZN(new_n25517_));
  INV_X1     g25450(.I(new_n25517_), .ZN(new_n25518_));
  NAND3_X1   g25451(.A1(new_n25515_), .A2(new_n25512_), .A3(new_n25516_), .ZN(new_n25519_));
  AOI21_X1   g25452(.A1(new_n25518_), .A2(new_n25519_), .B(new_n25504_), .ZN(new_n25520_));
  INV_X1     g25453(.I(new_n25519_), .ZN(new_n25521_));
  NOR3_X1    g25454(.A1(new_n25521_), .A2(new_n25517_), .A3(new_n25503_), .ZN(new_n25522_));
  NOR2_X1    g25455(.A1(new_n25520_), .A2(new_n25522_), .ZN(new_n25523_));
  AOI22_X1   g25456(.A1(new_n25350_), .A2(new_n25338_), .B1(new_n25346_), .B2(new_n25347_), .ZN(new_n25524_));
  NOR2_X1    g25457(.A1(new_n25350_), .A2(new_n25338_), .ZN(new_n25525_));
  OAI21_X1   g25458(.A1(new_n25524_), .A2(new_n25525_), .B(new_n25523_), .ZN(new_n25526_));
  NOR2_X1    g25459(.A1(new_n25524_), .A2(new_n25525_), .ZN(new_n25527_));
  OAI21_X1   g25460(.A1(new_n25520_), .A2(new_n25522_), .B(new_n25527_), .ZN(new_n25528_));
  AOI21_X1   g25461(.A1(new_n25528_), .A2(new_n25526_), .B(new_n25499_), .ZN(new_n25529_));
  NAND3_X1   g25462(.A1(new_n25528_), .A2(new_n25526_), .A3(new_n25499_), .ZN(new_n25530_));
  INV_X1     g25463(.I(new_n25530_), .ZN(new_n25531_));
  OAI21_X1   g25464(.A1(new_n25531_), .A2(new_n25529_), .B(new_n25493_), .ZN(new_n25532_));
  INV_X1     g25465(.I(new_n25493_), .ZN(new_n25533_));
  INV_X1     g25466(.I(new_n25529_), .ZN(new_n25534_));
  NAND3_X1   g25467(.A1(new_n25534_), .A2(new_n25533_), .A3(new_n25530_), .ZN(new_n25535_));
  NAND2_X1   g25468(.A1(new_n25535_), .A2(new_n25532_), .ZN(new_n25536_));
  NOR2_X1    g25469(.A1(new_n25358_), .A2(new_n25311_), .ZN(new_n25537_));
  NOR2_X1    g25470(.A1(new_n25304_), .A2(new_n25359_), .ZN(new_n25538_));
  NOR2_X1    g25471(.A1(new_n25537_), .A2(new_n25538_), .ZN(new_n25539_));
  INV_X1     g25472(.I(new_n25539_), .ZN(new_n25540_));
  AOI22_X1   g25473(.A1(new_n19439_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n19415_), .ZN(new_n25541_));
  NOR2_X1    g25474(.A1(new_n19423_), .A2(new_n3780_), .ZN(new_n25542_));
  OAI21_X1   g25475(.A1(new_n25542_), .A2(new_n25541_), .B(new_n3301_), .ZN(new_n25543_));
  INV_X1     g25476(.I(new_n25543_), .ZN(new_n25544_));
  NAND2_X1   g25477(.A1(new_n20939_), .A2(new_n25544_), .ZN(new_n25545_));
  NOR2_X1    g25478(.A1(new_n25545_), .A2(\a[23] ), .ZN(new_n25546_));
  INV_X1     g25479(.I(new_n25546_), .ZN(new_n25547_));
  NAND2_X1   g25480(.A1(new_n25545_), .A2(\a[23] ), .ZN(new_n25548_));
  NAND2_X1   g25481(.A1(new_n25547_), .A2(new_n25548_), .ZN(new_n25549_));
  NOR2_X1    g25482(.A1(new_n25549_), .A2(new_n25540_), .ZN(new_n25550_));
  INV_X1     g25483(.I(new_n25548_), .ZN(new_n25551_));
  NOR2_X1    g25484(.A1(new_n25551_), .A2(new_n25546_), .ZN(new_n25552_));
  NOR2_X1    g25485(.A1(new_n25552_), .A2(new_n25539_), .ZN(new_n25553_));
  OAI21_X1   g25486(.A1(new_n25553_), .A2(new_n25550_), .B(new_n25536_), .ZN(new_n25554_));
  AOI21_X1   g25487(.A1(new_n25534_), .A2(new_n25530_), .B(new_n25533_), .ZN(new_n25555_));
  NOR3_X1    g25488(.A1(new_n25531_), .A2(new_n25493_), .A3(new_n25529_), .ZN(new_n25556_));
  NOR2_X1    g25489(.A1(new_n25555_), .A2(new_n25556_), .ZN(new_n25557_));
  NOR2_X1    g25490(.A1(new_n25549_), .A2(new_n25539_), .ZN(new_n25558_));
  NOR2_X1    g25491(.A1(new_n25552_), .A2(new_n25540_), .ZN(new_n25559_));
  OAI21_X1   g25492(.A1(new_n25559_), .A2(new_n25558_), .B(new_n25557_), .ZN(new_n25560_));
  NAND2_X1   g25493(.A1(new_n25364_), .A2(new_n25365_), .ZN(new_n25561_));
  NOR2_X1    g25494(.A1(new_n25296_), .A2(new_n25288_), .ZN(new_n25562_));
  INV_X1     g25495(.I(new_n25562_), .ZN(new_n25563_));
  NOR2_X1    g25496(.A1(new_n25297_), .A2(new_n25287_), .ZN(new_n25564_));
  AOI21_X1   g25497(.A1(new_n25561_), .A2(new_n25563_), .B(new_n25564_), .ZN(new_n25565_));
  INV_X1     g25498(.I(new_n25565_), .ZN(new_n25566_));
  NAND3_X1   g25499(.A1(new_n25560_), .A2(new_n25554_), .A3(new_n25566_), .ZN(new_n25567_));
  INV_X1     g25500(.I(new_n25550_), .ZN(new_n25568_));
  NAND2_X1   g25501(.A1(new_n25549_), .A2(new_n25540_), .ZN(new_n25569_));
  AOI21_X1   g25502(.A1(new_n25568_), .A2(new_n25569_), .B(new_n25557_), .ZN(new_n25570_));
  NAND2_X1   g25503(.A1(new_n25552_), .A2(new_n25540_), .ZN(new_n25571_));
  NAND2_X1   g25504(.A1(new_n25549_), .A2(new_n25539_), .ZN(new_n25572_));
  AOI21_X1   g25505(.A1(new_n25571_), .A2(new_n25572_), .B(new_n25536_), .ZN(new_n25573_));
  OAI21_X1   g25506(.A1(new_n25570_), .A2(new_n25573_), .B(new_n25565_), .ZN(new_n25574_));
  NAND2_X1   g25507(.A1(new_n25574_), .A2(new_n25567_), .ZN(new_n25575_));
  OAI21_X1   g25508(.A1(new_n25564_), .A2(new_n25562_), .B(new_n25561_), .ZN(new_n25576_));
  XOR2_X1    g25509(.A1(new_n25296_), .A2(new_n25287_), .Z(new_n25577_));
  OAI21_X1   g25510(.A1(new_n25577_), .A2(new_n25561_), .B(new_n25576_), .ZN(new_n25578_));
  NAND2_X1   g25511(.A1(new_n25162_), .A2(new_n25164_), .ZN(new_n25579_));
  NAND2_X1   g25512(.A1(new_n25284_), .A2(new_n25579_), .ZN(new_n25580_));
  NOR2_X1    g25513(.A1(new_n25284_), .A2(new_n25579_), .ZN(new_n25581_));
  AOI21_X1   g25514(.A1(new_n25578_), .A2(new_n25580_), .B(new_n25581_), .ZN(new_n25582_));
  NOR2_X1    g25515(.A1(new_n25575_), .A2(new_n25582_), .ZN(new_n25583_));
  NOR3_X1    g25516(.A1(new_n25570_), .A2(new_n25573_), .A3(new_n25565_), .ZN(new_n25584_));
  AOI21_X1   g25517(.A1(new_n25560_), .A2(new_n25554_), .B(new_n25566_), .ZN(new_n25585_));
  NOR2_X1    g25518(.A1(new_n25584_), .A2(new_n25585_), .ZN(new_n25586_));
  NAND2_X1   g25519(.A1(new_n25580_), .A2(new_n25578_), .ZN(new_n25587_));
  INV_X1     g25520(.I(new_n25581_), .ZN(new_n25588_));
  NAND2_X1   g25521(.A1(new_n25587_), .A2(new_n25588_), .ZN(new_n25589_));
  NOR2_X1    g25522(.A1(new_n25586_), .A2(new_n25589_), .ZN(new_n25590_));
  OAI21_X1   g25523(.A1(new_n25590_), .A2(new_n25583_), .B(new_n25488_), .ZN(new_n25591_));
  INV_X1     g25524(.I(new_n25488_), .ZN(new_n25592_));
  NAND2_X1   g25525(.A1(new_n25586_), .A2(new_n25589_), .ZN(new_n25593_));
  NAND2_X1   g25526(.A1(new_n25575_), .A2(new_n25582_), .ZN(new_n25594_));
  NAND3_X1   g25527(.A1(new_n25593_), .A2(new_n25594_), .A3(new_n25592_), .ZN(new_n25595_));
  AOI21_X1   g25528(.A1(new_n25591_), .A2(new_n25595_), .B(new_n25483_), .ZN(new_n25596_));
  AOI21_X1   g25529(.A1(new_n25593_), .A2(new_n25594_), .B(new_n25592_), .ZN(new_n25597_));
  NOR3_X1    g25530(.A1(new_n25590_), .A2(new_n25583_), .A3(new_n25488_), .ZN(new_n25598_));
  NOR3_X1    g25531(.A1(new_n25597_), .A2(new_n25598_), .A3(new_n25482_), .ZN(new_n25599_));
  NOR2_X1    g25532(.A1(new_n25599_), .A2(new_n25596_), .ZN(new_n25600_));
  NOR2_X1    g25533(.A1(new_n25392_), .A2(new_n25393_), .ZN(new_n25601_));
  NOR2_X1    g25534(.A1(new_n25274_), .A2(new_n25390_), .ZN(new_n25602_));
  NAND2_X1   g25535(.A1(new_n25274_), .A2(new_n25390_), .ZN(new_n25603_));
  OAI21_X1   g25536(.A1(new_n25601_), .A2(new_n25602_), .B(new_n25603_), .ZN(new_n25604_));
  NAND2_X1   g25537(.A1(new_n25600_), .A2(new_n25604_), .ZN(new_n25605_));
  OAI21_X1   g25538(.A1(new_n25597_), .A2(new_n25598_), .B(new_n25482_), .ZN(new_n25606_));
  NAND3_X1   g25539(.A1(new_n25591_), .A2(new_n25595_), .A3(new_n25483_), .ZN(new_n25607_));
  NAND2_X1   g25540(.A1(new_n25606_), .A2(new_n25607_), .ZN(new_n25608_));
  INV_X1     g25541(.I(new_n25601_), .ZN(new_n25609_));
  NAND2_X1   g25542(.A1(new_n25397_), .A2(new_n25394_), .ZN(new_n25610_));
  NOR2_X1    g25543(.A1(new_n25397_), .A2(new_n25394_), .ZN(new_n25611_));
  AOI21_X1   g25544(.A1(new_n25609_), .A2(new_n25610_), .B(new_n25611_), .ZN(new_n25612_));
  NAND2_X1   g25545(.A1(new_n25608_), .A2(new_n25612_), .ZN(new_n25613_));
  AOI21_X1   g25546(.A1(new_n25613_), .A2(new_n25605_), .B(new_n25477_), .ZN(new_n25614_));
  XOR2_X1    g25547(.A1(new_n25476_), .A2(\a[14] ), .Z(new_n25615_));
  NOR2_X1    g25548(.A1(new_n25608_), .A2(new_n25612_), .ZN(new_n25616_));
  NOR2_X1    g25549(.A1(new_n25600_), .A2(new_n25604_), .ZN(new_n25617_));
  NOR3_X1    g25550(.A1(new_n25616_), .A2(new_n25617_), .A3(new_n25615_), .ZN(new_n25618_));
  OAI21_X1   g25551(.A1(new_n25614_), .A2(new_n25618_), .B(new_n25473_), .ZN(new_n25619_));
  OAI21_X1   g25552(.A1(new_n25616_), .A2(new_n25617_), .B(new_n25615_), .ZN(new_n25620_));
  NAND3_X1   g25553(.A1(new_n25613_), .A2(new_n25605_), .A3(new_n25477_), .ZN(new_n25621_));
  NAND3_X1   g25554(.A1(new_n25620_), .A2(new_n25621_), .A3(new_n25472_), .ZN(new_n25622_));
  INV_X1     g25555(.I(new_n25267_), .ZN(new_n25623_));
  OAI21_X1   g25556(.A1(new_n25611_), .A2(new_n25602_), .B(new_n25609_), .ZN(new_n25624_));
  XOR2_X1    g25557(.A1(new_n25397_), .A2(new_n25390_), .Z(new_n25625_));
  OAI21_X1   g25558(.A1(new_n25625_), .A2(new_n25609_), .B(new_n25624_), .ZN(new_n25626_));
  OAI21_X1   g25559(.A1(new_n25409_), .A2(new_n25623_), .B(new_n25626_), .ZN(new_n25627_));
  NAND2_X1   g25560(.A1(new_n25409_), .A2(new_n25623_), .ZN(new_n25628_));
  NAND2_X1   g25561(.A1(new_n25627_), .A2(new_n25628_), .ZN(new_n25629_));
  NAND3_X1   g25562(.A1(new_n25629_), .A2(new_n25619_), .A3(new_n25622_), .ZN(new_n25630_));
  INV_X1     g25563(.I(new_n25630_), .ZN(new_n25631_));
  AOI21_X1   g25564(.A1(new_n25619_), .A2(new_n25622_), .B(new_n25629_), .ZN(new_n25632_));
  OAI21_X1   g25565(.A1(new_n25631_), .A2(new_n25632_), .B(new_n25467_), .ZN(new_n25633_));
  INV_X1     g25566(.I(new_n25467_), .ZN(new_n25634_));
  NAND2_X1   g25567(.A1(new_n25619_), .A2(new_n25622_), .ZN(new_n25635_));
  NAND3_X1   g25568(.A1(new_n25635_), .A2(new_n25627_), .A3(new_n25628_), .ZN(new_n25636_));
  NAND3_X1   g25569(.A1(new_n25636_), .A2(new_n25634_), .A3(new_n25630_), .ZN(new_n25637_));
  AOI21_X1   g25570(.A1(new_n25633_), .A2(new_n25637_), .B(new_n25462_), .ZN(new_n25638_));
  XOR2_X1    g25571(.A1(new_n25461_), .A2(\a[8] ), .Z(new_n25639_));
  AOI21_X1   g25572(.A1(new_n25636_), .A2(new_n25630_), .B(new_n25634_), .ZN(new_n25640_));
  NOR3_X1    g25573(.A1(new_n25631_), .A2(new_n25632_), .A3(new_n25467_), .ZN(new_n25641_));
  NOR3_X1    g25574(.A1(new_n25641_), .A2(new_n25640_), .A3(new_n25639_), .ZN(new_n25642_));
  NOR2_X1    g25575(.A1(new_n25189_), .A2(new_n25062_), .ZN(new_n25643_));
  NAND2_X1   g25576(.A1(new_n25259_), .A2(new_n25643_), .ZN(new_n25644_));
  XOR2_X1    g25577(.A1(new_n25406_), .A2(new_n25263_), .Z(new_n25645_));
  OAI21_X1   g25578(.A1(new_n25259_), .A2(new_n25643_), .B(new_n25645_), .ZN(new_n25646_));
  OAI21_X1   g25579(.A1(new_n24599_), .A2(new_n24835_), .B(new_n24376_), .ZN(new_n25647_));
  NOR2_X1    g25580(.A1(new_n24613_), .A2(new_n6913_), .ZN(new_n25648_));
  NOR2_X1    g25581(.A1(new_n24835_), .A2(new_n11868_), .ZN(new_n25649_));
  OAI21_X1   g25582(.A1(new_n25649_), .A2(new_n25648_), .B(new_n6835_), .ZN(new_n25650_));
  INV_X1     g25583(.I(new_n25650_), .ZN(new_n25651_));
  NAND3_X1   g25584(.A1(new_n25647_), .A2(new_n65_), .A3(new_n25651_), .ZN(new_n25652_));
  OAI21_X1   g25585(.A1(new_n25017_), .A2(new_n25650_), .B(\a[5] ), .ZN(new_n25653_));
  NAND2_X1   g25586(.A1(new_n25652_), .A2(new_n25653_), .ZN(new_n25654_));
  NAND3_X1   g25587(.A1(new_n25646_), .A2(new_n25644_), .A3(new_n25654_), .ZN(new_n25655_));
  INV_X1     g25588(.I(new_n25643_), .ZN(new_n25656_));
  NOR2_X1    g25589(.A1(new_n25414_), .A2(new_n25656_), .ZN(new_n25657_));
  XOR2_X1    g25590(.A1(new_n25406_), .A2(new_n25409_), .Z(new_n25658_));
  AOI21_X1   g25591(.A1(new_n25414_), .A2(new_n25656_), .B(new_n25658_), .ZN(new_n25659_));
  NOR3_X1    g25592(.A1(new_n25017_), .A2(\a[5] ), .A3(new_n25650_), .ZN(new_n25660_));
  AOI21_X1   g25593(.A1(new_n25647_), .A2(new_n25651_), .B(new_n65_), .ZN(new_n25661_));
  NOR2_X1    g25594(.A1(new_n25661_), .A2(new_n25660_), .ZN(new_n25662_));
  OAI21_X1   g25595(.A1(new_n25659_), .A2(new_n25657_), .B(new_n25662_), .ZN(new_n25663_));
  NAND2_X1   g25596(.A1(new_n25663_), .A2(new_n25655_), .ZN(new_n25664_));
  AOI21_X1   g25597(.A1(new_n25431_), .A2(new_n25426_), .B(new_n25418_), .ZN(new_n25665_));
  NOR2_X1    g25598(.A1(new_n25431_), .A2(new_n25426_), .ZN(new_n25666_));
  NOR2_X1    g25599(.A1(new_n25665_), .A2(new_n25666_), .ZN(new_n25667_));
  XOR2_X1    g25600(.A1(new_n25667_), .A2(new_n25664_), .Z(new_n25668_));
  OAI21_X1   g25601(.A1(new_n25638_), .A2(new_n25642_), .B(new_n25668_), .ZN(new_n25669_));
  OAI21_X1   g25602(.A1(new_n25641_), .A2(new_n25640_), .B(new_n25639_), .ZN(new_n25670_));
  NAND3_X1   g25603(.A1(new_n25633_), .A2(new_n25637_), .A3(new_n25462_), .ZN(new_n25671_));
  NOR3_X1    g25604(.A1(new_n25659_), .A2(new_n25657_), .A3(new_n25662_), .ZN(new_n25672_));
  AOI21_X1   g25605(.A1(new_n25646_), .A2(new_n25644_), .B(new_n25654_), .ZN(new_n25673_));
  NOR2_X1    g25606(.A1(new_n25672_), .A2(new_n25673_), .ZN(new_n25674_));
  XOR2_X1    g25607(.A1(new_n25667_), .A2(new_n25674_), .Z(new_n25675_));
  NAND3_X1   g25608(.A1(new_n25675_), .A2(new_n25670_), .A3(new_n25671_), .ZN(new_n25676_));
  NAND2_X1   g25609(.A1(new_n25669_), .A2(new_n25676_), .ZN(new_n25677_));
  AND3_X2    g25610(.A1(new_n25677_), .A2(new_n25449_), .A3(new_n25457_), .Z(new_n25678_));
  AOI21_X1   g25611(.A1(new_n25449_), .A2(new_n25457_), .B(new_n25677_), .ZN(new_n25679_));
  NOR2_X1    g25612(.A1(new_n25678_), .A2(new_n25679_), .ZN(new_n25680_));
  INV_X1     g25613(.I(new_n25680_), .ZN(new_n25681_));
  XOR2_X1    g25614(.A1(new_n25447_), .A2(new_n25681_), .Z(\result[9] ));
  AOI22_X1   g25615(.A1(new_n25208_), .A2(new_n25052_), .B1(new_n25437_), .B2(new_n25436_), .ZN(new_n25683_));
  NOR3_X1    g25616(.A1(new_n25244_), .A2(new_n25428_), .A3(new_n25434_), .ZN(new_n25684_));
  NOR3_X1    g25617(.A1(new_n25683_), .A2(new_n25684_), .A3(new_n25212_), .ZN(new_n25685_));
  NOR3_X1    g25618(.A1(new_n25229_), .A2(new_n25440_), .A3(new_n25685_), .ZN(new_n25686_));
  INV_X1     g25619(.I(new_n25667_), .ZN(new_n25687_));
  NAND3_X1   g25620(.A1(new_n25664_), .A2(new_n25670_), .A3(new_n25671_), .ZN(new_n25688_));
  OAI21_X1   g25621(.A1(new_n25638_), .A2(new_n25642_), .B(new_n25674_), .ZN(new_n25689_));
  NAND2_X1   g25622(.A1(new_n25689_), .A2(new_n25688_), .ZN(new_n25690_));
  INV_X1     g25623(.I(new_n25690_), .ZN(new_n25691_));
  NOR2_X1    g25624(.A1(new_n25691_), .A2(new_n25687_), .ZN(new_n25692_));
  INV_X1     g25625(.I(new_n25692_), .ZN(new_n25693_));
  NOR2_X1    g25626(.A1(new_n25690_), .A2(new_n25667_), .ZN(new_n25694_));
  NOR2_X1    g25627(.A1(new_n25691_), .A2(new_n25687_), .ZN(new_n25695_));
  OAI21_X1   g25628(.A1(new_n25694_), .A2(new_n25695_), .B(new_n25457_), .ZN(new_n25696_));
  OAI21_X1   g25629(.A1(new_n25686_), .A2(new_n25696_), .B(new_n25693_), .ZN(new_n25697_));
  NAND2_X1   g25630(.A1(new_n25646_), .A2(new_n25644_), .ZN(new_n25698_));
  OAI22_X1   g25631(.A1(new_n25642_), .A2(new_n25638_), .B1(new_n25698_), .B2(new_n25654_), .ZN(new_n25699_));
  NAND2_X1   g25632(.A1(new_n25698_), .A2(new_n25654_), .ZN(new_n25700_));
  NAND2_X1   g25633(.A1(new_n25699_), .A2(new_n25700_), .ZN(new_n25701_));
  NAND2_X1   g25634(.A1(new_n25462_), .A2(new_n25629_), .ZN(new_n25702_));
  NOR2_X1    g25635(.A1(new_n25462_), .A2(new_n25629_), .ZN(new_n25703_));
  XOR2_X1    g25636(.A1(new_n25635_), .A2(new_n25467_), .Z(new_n25704_));
  OAI21_X1   g25637(.A1(new_n25703_), .A2(new_n25704_), .B(new_n25702_), .ZN(new_n25705_));
  OAI22_X1   g25638(.A1(new_n24376_), .A2(new_n6788_), .B1(new_n6783_), .B2(new_n24167_), .ZN(new_n25706_));
  NAND2_X1   g25639(.A1(new_n24620_), .A2(new_n6784_), .ZN(new_n25707_));
  AOI21_X1   g25640(.A1(new_n25707_), .A2(new_n25706_), .B(new_n6776_), .ZN(new_n25708_));
  NAND2_X1   g25641(.A1(new_n24618_), .A2(new_n25708_), .ZN(new_n25709_));
  XOR2_X1    g25642(.A1(new_n25709_), .A2(new_n4009_), .Z(new_n25710_));
  INV_X1     g25643(.I(new_n25710_), .ZN(new_n25711_));
  AOI22_X1   g25644(.A1(new_n25488_), .A2(new_n25565_), .B1(new_n25554_), .B2(new_n25560_), .ZN(new_n25712_));
  NOR2_X1    g25645(.A1(new_n25488_), .A2(new_n25565_), .ZN(new_n25713_));
  NOR2_X1    g25646(.A1(new_n25712_), .A2(new_n25713_), .ZN(new_n25714_));
  INV_X1     g25647(.I(new_n25714_), .ZN(new_n25715_));
  OAI22_X1   g25648(.A1(new_n17775_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19475_), .ZN(new_n25716_));
  NAND2_X1   g25649(.A1(new_n21157_), .A2(new_n4469_), .ZN(new_n25717_));
  AOI21_X1   g25650(.A1(new_n25717_), .A2(new_n25716_), .B(new_n4468_), .ZN(new_n25718_));
  NAND2_X1   g25651(.A1(new_n21155_), .A2(new_n25718_), .ZN(new_n25719_));
  XOR2_X1    g25652(.A1(new_n25719_), .A2(\a[17] ), .Z(new_n25720_));
  OAI22_X1   g25653(.A1(new_n19437_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n17784_), .ZN(new_n25721_));
  NAND2_X1   g25654(.A1(new_n19472_), .A2(new_n4096_), .ZN(new_n25722_));
  AOI21_X1   g25655(.A1(new_n25722_), .A2(new_n25721_), .B(new_n4095_), .ZN(new_n25723_));
  NAND2_X1   g25656(.A1(new_n21117_), .A2(new_n25723_), .ZN(new_n25724_));
  XOR2_X1    g25657(.A1(new_n25724_), .A2(\a[20] ), .Z(new_n25725_));
  OAI22_X1   g25658(.A1(new_n19423_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n17787_), .ZN(new_n25726_));
  NAND2_X1   g25659(.A1(new_n20896_), .A2(new_n3312_), .ZN(new_n25727_));
  AOI21_X1   g25660(.A1(new_n25727_), .A2(new_n25726_), .B(new_n3302_), .ZN(new_n25728_));
  NAND2_X1   g25661(.A1(new_n22226_), .A2(new_n25728_), .ZN(new_n25729_));
  XOR2_X1    g25662(.A1(new_n25729_), .A2(\a[23] ), .Z(new_n25730_));
  INV_X1     g25663(.I(new_n25730_), .ZN(new_n25731_));
  OAI22_X1   g25664(.A1(new_n19410_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n17789_), .ZN(new_n25732_));
  NAND2_X1   g25665(.A1(new_n19415_), .A2(new_n3317_), .ZN(new_n25733_));
  AOI21_X1   g25666(.A1(new_n25733_), .A2(new_n25732_), .B(new_n3260_), .ZN(new_n25734_));
  NAND2_X1   g25667(.A1(new_n20846_), .A2(new_n25734_), .ZN(new_n25735_));
  XOR2_X1    g25668(.A1(new_n25735_), .A2(\a[26] ), .Z(new_n25736_));
  AOI22_X1   g25669(.A1(new_n19394_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n17794_), .ZN(new_n25737_));
  AOI21_X1   g25670(.A1(new_n2750_), .A2(new_n19399_), .B(new_n25737_), .ZN(new_n25738_));
  OR3_X2     g25671(.A1(new_n22541_), .A2(new_n2737_), .A3(new_n25738_), .Z(new_n25739_));
  XOR2_X1    g25672(.A1(new_n25739_), .A2(\a[29] ), .Z(new_n25740_));
  INV_X1     g25673(.I(new_n25740_), .ZN(new_n25741_));
  NAND2_X1   g25674(.A1(new_n25514_), .A2(new_n25513_), .ZN(new_n25742_));
  XOR2_X1    g25675(.A1(new_n25095_), .A2(new_n25512_), .Z(new_n25743_));
  NAND2_X1   g25676(.A1(new_n25742_), .A2(new_n25743_), .ZN(new_n25744_));
  NOR2_X1    g25677(.A1(new_n25742_), .A2(new_n25743_), .ZN(new_n25745_));
  NOR2_X1    g25678(.A1(new_n25745_), .A2(new_n25504_), .ZN(new_n25746_));
  NAND2_X1   g25679(.A1(new_n25746_), .A2(new_n25744_), .ZN(new_n25747_));
  AOI21_X1   g25680(.A1(new_n25523_), .A2(new_n25527_), .B(new_n25747_), .ZN(new_n25748_));
  INV_X1     g25681(.I(new_n25512_), .ZN(new_n25749_));
  AOI22_X1   g25682(.A1(new_n25514_), .A2(new_n25513_), .B1(new_n25095_), .B2(new_n25749_), .ZN(new_n25750_));
  AOI21_X1   g25683(.A1(new_n25314_), .A2(new_n25512_), .B(new_n25750_), .ZN(new_n25751_));
  NOR2_X1    g25684(.A1(new_n24835_), .A2(new_n11870_), .ZN(new_n25752_));
  OAI22_X1   g25685(.A1(new_n25752_), .A2(\a[5] ), .B1(new_n11887_), .B2(new_n24835_), .ZN(new_n25753_));
  INV_X1     g25686(.I(new_n19709_), .ZN(new_n25754_));
  NOR4_X1    g25687(.A1(new_n446_), .A2(new_n251_), .A3(new_n944_), .A4(new_n906_), .ZN(new_n25755_));
  NAND2_X1   g25688(.A1(new_n2398_), .A2(new_n3459_), .ZN(new_n25756_));
  NOR4_X1    g25689(.A1(new_n25756_), .A2(new_n25755_), .A3(new_n369_), .A4(new_n1589_), .ZN(new_n25757_));
  NAND2_X1   g25690(.A1(new_n1751_), .A2(new_n2428_), .ZN(new_n25758_));
  NOR3_X1    g25691(.A1(new_n3512_), .A2(new_n25758_), .A3(new_n3855_), .ZN(new_n25759_));
  NAND4_X1   g25692(.A1(new_n25754_), .A2(new_n11485_), .A3(new_n25757_), .A4(new_n25759_), .ZN(new_n25760_));
  NOR3_X1    g25693(.A1(new_n2222_), .A2(new_n2948_), .A3(new_n25760_), .ZN(new_n25761_));
  XOR2_X1    g25694(.A1(new_n25753_), .A2(new_n25761_), .Z(new_n25762_));
  NOR2_X1    g25695(.A1(new_n25762_), .A2(new_n25095_), .ZN(new_n25763_));
  INV_X1     g25696(.I(new_n25761_), .ZN(new_n25764_));
  NAND2_X1   g25697(.A1(new_n25753_), .A2(new_n25764_), .ZN(new_n25765_));
  OR2_X2     g25698(.A1(new_n25753_), .A2(new_n25764_), .Z(new_n25766_));
  AOI21_X1   g25699(.A1(new_n25766_), .A2(new_n25765_), .B(new_n25314_), .ZN(new_n25767_));
  NOR2_X1    g25700(.A1(new_n25763_), .A2(new_n25767_), .ZN(new_n25768_));
  NAND2_X1   g25701(.A1(new_n19386_), .A2(new_n3332_), .ZN(new_n25769_));
  NAND2_X1   g25702(.A1(new_n20127_), .A2(new_n3189_), .ZN(new_n25770_));
  AOI21_X1   g25703(.A1(new_n17798_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n25771_));
  NAND4_X1   g25704(.A1(new_n20162_), .A2(new_n25769_), .A3(new_n25770_), .A4(new_n25771_), .ZN(new_n25772_));
  XNOR2_X1   g25705(.A1(new_n25768_), .A2(new_n25772_), .ZN(new_n25773_));
  NAND2_X1   g25706(.A1(new_n25768_), .A2(new_n25772_), .ZN(new_n25774_));
  OR2_X2     g25707(.A1(new_n25768_), .A2(new_n25772_), .Z(new_n25775_));
  NAND2_X1   g25708(.A1(new_n25775_), .A2(new_n25774_), .ZN(new_n25776_));
  NAND2_X1   g25709(.A1(new_n25776_), .A2(new_n25751_), .ZN(new_n25777_));
  OAI21_X1   g25710(.A1(new_n25751_), .A2(new_n25773_), .B(new_n25777_), .ZN(new_n25778_));
  XOR2_X1    g25711(.A1(new_n25748_), .A2(new_n25778_), .Z(new_n25779_));
  NOR2_X1    g25712(.A1(new_n25493_), .A2(new_n25498_), .ZN(new_n25780_));
  NOR2_X1    g25713(.A1(new_n25534_), .A2(new_n25533_), .ZN(new_n25781_));
  NOR2_X1    g25714(.A1(new_n25781_), .A2(new_n25780_), .ZN(new_n25782_));
  INV_X1     g25715(.I(new_n25782_), .ZN(new_n25783_));
  NAND2_X1   g25716(.A1(new_n25783_), .A2(new_n25779_), .ZN(new_n25784_));
  INV_X1     g25717(.I(new_n25779_), .ZN(new_n25785_));
  NAND2_X1   g25718(.A1(new_n25782_), .A2(new_n25785_), .ZN(new_n25786_));
  AOI21_X1   g25719(.A1(new_n25784_), .A2(new_n25786_), .B(new_n25741_), .ZN(new_n25787_));
  NAND3_X1   g25720(.A1(new_n25784_), .A2(new_n25741_), .A3(new_n25786_), .ZN(new_n25788_));
  INV_X1     g25721(.I(new_n25788_), .ZN(new_n25789_));
  OAI21_X1   g25722(.A1(new_n25789_), .A2(new_n25787_), .B(new_n25736_), .ZN(new_n25790_));
  INV_X1     g25723(.I(new_n25736_), .ZN(new_n25791_));
  NAND2_X1   g25724(.A1(new_n25784_), .A2(new_n25786_), .ZN(new_n25792_));
  NAND2_X1   g25725(.A1(new_n25792_), .A2(new_n25740_), .ZN(new_n25793_));
  NAND3_X1   g25726(.A1(new_n25793_), .A2(new_n25791_), .A3(new_n25788_), .ZN(new_n25794_));
  AOI21_X1   g25727(.A1(new_n25568_), .A2(new_n25536_), .B(new_n25553_), .ZN(new_n25795_));
  INV_X1     g25728(.I(new_n25795_), .ZN(new_n25796_));
  NAND3_X1   g25729(.A1(new_n25790_), .A2(new_n25794_), .A3(new_n25796_), .ZN(new_n25797_));
  AOI21_X1   g25730(.A1(new_n25793_), .A2(new_n25788_), .B(new_n25791_), .ZN(new_n25798_));
  NOR3_X1    g25731(.A1(new_n25789_), .A2(new_n25736_), .A3(new_n25787_), .ZN(new_n25799_));
  OAI21_X1   g25732(.A1(new_n25799_), .A2(new_n25798_), .B(new_n25795_), .ZN(new_n25800_));
  AOI21_X1   g25733(.A1(new_n25800_), .A2(new_n25797_), .B(new_n25731_), .ZN(new_n25801_));
  NOR3_X1    g25734(.A1(new_n25799_), .A2(new_n25798_), .A3(new_n25795_), .ZN(new_n25802_));
  AOI21_X1   g25735(.A1(new_n25790_), .A2(new_n25794_), .B(new_n25796_), .ZN(new_n25803_));
  NOR3_X1    g25736(.A1(new_n25802_), .A2(new_n25803_), .A3(new_n25730_), .ZN(new_n25804_));
  OAI21_X1   g25737(.A1(new_n25804_), .A2(new_n25801_), .B(new_n25725_), .ZN(new_n25805_));
  INV_X1     g25738(.I(new_n25725_), .ZN(new_n25806_));
  OAI21_X1   g25739(.A1(new_n25802_), .A2(new_n25803_), .B(new_n25730_), .ZN(new_n25807_));
  NAND3_X1   g25740(.A1(new_n25800_), .A2(new_n25797_), .A3(new_n25731_), .ZN(new_n25808_));
  NAND3_X1   g25741(.A1(new_n25807_), .A2(new_n25808_), .A3(new_n25806_), .ZN(new_n25809_));
  NAND2_X1   g25742(.A1(new_n25805_), .A2(new_n25809_), .ZN(new_n25810_));
  NOR2_X1    g25743(.A1(new_n25482_), .A2(new_n25582_), .ZN(new_n25811_));
  NAND2_X1   g25744(.A1(new_n25482_), .A2(new_n25582_), .ZN(new_n25812_));
  XOR2_X1    g25745(.A1(new_n25575_), .A2(new_n25592_), .Z(new_n25813_));
  AOI21_X1   g25746(.A1(new_n25813_), .A2(new_n25812_), .B(new_n25811_), .ZN(new_n25814_));
  NOR2_X1    g25747(.A1(new_n25810_), .A2(new_n25814_), .ZN(new_n25815_));
  AOI21_X1   g25748(.A1(new_n25807_), .A2(new_n25808_), .B(new_n25806_), .ZN(new_n25816_));
  NOR3_X1    g25749(.A1(new_n25804_), .A2(new_n25801_), .A3(new_n25725_), .ZN(new_n25817_));
  NOR2_X1    g25750(.A1(new_n25817_), .A2(new_n25816_), .ZN(new_n25818_));
  INV_X1     g25751(.I(new_n25814_), .ZN(new_n25819_));
  NOR2_X1    g25752(.A1(new_n25818_), .A2(new_n25819_), .ZN(new_n25820_));
  OAI21_X1   g25753(.A1(new_n25820_), .A2(new_n25815_), .B(new_n25720_), .ZN(new_n25821_));
  INV_X1     g25754(.I(new_n25720_), .ZN(new_n25822_));
  NAND2_X1   g25755(.A1(new_n25818_), .A2(new_n25819_), .ZN(new_n25823_));
  NAND2_X1   g25756(.A1(new_n25810_), .A2(new_n25814_), .ZN(new_n25824_));
  NAND3_X1   g25757(.A1(new_n25823_), .A2(new_n25824_), .A3(new_n25822_), .ZN(new_n25825_));
  AOI21_X1   g25758(.A1(new_n25821_), .A2(new_n25825_), .B(new_n25715_), .ZN(new_n25826_));
  AOI21_X1   g25759(.A1(new_n25823_), .A2(new_n25824_), .B(new_n25822_), .ZN(new_n25827_));
  NOR3_X1    g25760(.A1(new_n25820_), .A2(new_n25815_), .A3(new_n25720_), .ZN(new_n25828_));
  NOR3_X1    g25761(.A1(new_n25827_), .A2(new_n25828_), .A3(new_n25714_), .ZN(new_n25829_));
  NOR2_X1    g25762(.A1(new_n25829_), .A2(new_n25826_), .ZN(new_n25830_));
  OAI22_X1   g25763(.A1(new_n19512_), .A2(new_n6089_), .B1(new_n21960_), .B2(new_n6094_), .ZN(new_n25831_));
  NAND2_X1   g25764(.A1(new_n22048_), .A2(new_n6090_), .ZN(new_n25832_));
  AOI21_X1   g25765(.A1(new_n25832_), .A2(new_n25831_), .B(new_n6082_), .ZN(new_n25833_));
  NAND2_X1   g25766(.A1(new_n22175_), .A2(new_n25833_), .ZN(new_n25834_));
  XOR2_X1    g25767(.A1(new_n25834_), .A2(\a[14] ), .Z(new_n25835_));
  INV_X1     g25768(.I(new_n25835_), .ZN(new_n25836_));
  NOR2_X1    g25769(.A1(new_n25600_), .A2(new_n25473_), .ZN(new_n25837_));
  INV_X1     g25770(.I(new_n25837_), .ZN(new_n25838_));
  NOR2_X1    g25771(.A1(new_n25836_), .A2(new_n25838_), .ZN(new_n25839_));
  NOR2_X1    g25772(.A1(new_n25835_), .A2(new_n25837_), .ZN(new_n25840_));
  XOR2_X1    g25773(.A1(new_n25608_), .A2(new_n25473_), .Z(new_n25841_));
  NOR2_X1    g25774(.A1(new_n25841_), .A2(new_n25615_), .ZN(new_n25842_));
  INV_X1     g25775(.I(new_n25842_), .ZN(new_n25843_));
  NOR3_X1    g25776(.A1(new_n25843_), .A2(new_n25839_), .A3(new_n25840_), .ZN(new_n25844_));
  INV_X1     g25777(.I(new_n25839_), .ZN(new_n25845_));
  INV_X1     g25778(.I(new_n25840_), .ZN(new_n25846_));
  AOI21_X1   g25779(.A1(new_n25845_), .A2(new_n25846_), .B(new_n25842_), .ZN(new_n25847_));
  OAI22_X1   g25780(.A1(new_n22115_), .A2(new_n4716_), .B1(new_n4719_), .B2(new_n22149_), .ZN(new_n25848_));
  NAND2_X1   g25781(.A1(new_n23957_), .A2(new_n4709_), .ZN(new_n25849_));
  AOI21_X1   g25782(.A1(new_n25848_), .A2(new_n25849_), .B(new_n4707_), .ZN(new_n25850_));
  NAND2_X1   g25783(.A1(new_n23955_), .A2(new_n25850_), .ZN(new_n25851_));
  XOR2_X1    g25784(.A1(new_n25851_), .A2(\a[11] ), .Z(new_n25852_));
  OAI21_X1   g25785(.A1(new_n25844_), .A2(new_n25847_), .B(new_n25852_), .ZN(new_n25853_));
  NAND3_X1   g25786(.A1(new_n25845_), .A2(new_n25846_), .A3(new_n25842_), .ZN(new_n25854_));
  OAI21_X1   g25787(.A1(new_n25839_), .A2(new_n25840_), .B(new_n25843_), .ZN(new_n25855_));
  XOR2_X1    g25788(.A1(new_n25851_), .A2(new_n4034_), .Z(new_n25856_));
  NAND3_X1   g25789(.A1(new_n25855_), .A2(new_n25854_), .A3(new_n25856_), .ZN(new_n25857_));
  AOI21_X1   g25790(.A1(new_n25857_), .A2(new_n25853_), .B(new_n25830_), .ZN(new_n25858_));
  OAI21_X1   g25791(.A1(new_n25827_), .A2(new_n25828_), .B(new_n25714_), .ZN(new_n25859_));
  NAND3_X1   g25792(.A1(new_n25821_), .A2(new_n25825_), .A3(new_n25715_), .ZN(new_n25860_));
  NAND2_X1   g25793(.A1(new_n25859_), .A2(new_n25860_), .ZN(new_n25861_));
  NAND3_X1   g25794(.A1(new_n25855_), .A2(new_n25854_), .A3(new_n25852_), .ZN(new_n25862_));
  OAI21_X1   g25795(.A1(new_n25844_), .A2(new_n25847_), .B(new_n25856_), .ZN(new_n25863_));
  AOI21_X1   g25796(.A1(new_n25862_), .A2(new_n25863_), .B(new_n25861_), .ZN(new_n25864_));
  NOR2_X1    g25797(.A1(new_n25477_), .A2(new_n25472_), .ZN(new_n25865_));
  NOR2_X1    g25798(.A1(new_n25615_), .A2(new_n25473_), .ZN(new_n25866_));
  OAI21_X1   g25799(.A1(new_n25865_), .A2(new_n25866_), .B(new_n25608_), .ZN(new_n25867_));
  XOR2_X1    g25800(.A1(new_n25615_), .A2(new_n25472_), .Z(new_n25868_));
  OAI21_X1   g25801(.A1(new_n25608_), .A2(new_n25868_), .B(new_n25867_), .ZN(new_n25869_));
  NAND2_X1   g25802(.A1(new_n25467_), .A2(new_n25612_), .ZN(new_n25870_));
  NOR2_X1    g25803(.A1(new_n25467_), .A2(new_n25612_), .ZN(new_n25871_));
  AOI21_X1   g25804(.A1(new_n25869_), .A2(new_n25870_), .B(new_n25871_), .ZN(new_n25872_));
  NOR3_X1    g25805(.A1(new_n25858_), .A2(new_n25864_), .A3(new_n25872_), .ZN(new_n25873_));
  AOI21_X1   g25806(.A1(new_n25855_), .A2(new_n25854_), .B(new_n25856_), .ZN(new_n25874_));
  NOR3_X1    g25807(.A1(new_n25844_), .A2(new_n25847_), .A3(new_n25852_), .ZN(new_n25875_));
  OAI21_X1   g25808(.A1(new_n25874_), .A2(new_n25875_), .B(new_n25861_), .ZN(new_n25876_));
  NOR3_X1    g25809(.A1(new_n25844_), .A2(new_n25847_), .A3(new_n25856_), .ZN(new_n25877_));
  AOI21_X1   g25810(.A1(new_n25855_), .A2(new_n25854_), .B(new_n25852_), .ZN(new_n25878_));
  OAI21_X1   g25811(.A1(new_n25878_), .A2(new_n25877_), .B(new_n25830_), .ZN(new_n25879_));
  INV_X1     g25812(.I(new_n25872_), .ZN(new_n25880_));
  AOI21_X1   g25813(.A1(new_n25876_), .A2(new_n25879_), .B(new_n25880_), .ZN(new_n25881_));
  OAI21_X1   g25814(.A1(new_n25881_), .A2(new_n25873_), .B(new_n25711_), .ZN(new_n25882_));
  NAND3_X1   g25815(.A1(new_n25876_), .A2(new_n25879_), .A3(new_n25880_), .ZN(new_n25883_));
  OAI21_X1   g25816(.A1(new_n25858_), .A2(new_n25864_), .B(new_n25872_), .ZN(new_n25884_));
  NAND3_X1   g25817(.A1(new_n25884_), .A2(new_n25883_), .A3(new_n25710_), .ZN(new_n25885_));
  AOI21_X1   g25818(.A1(new_n25882_), .A2(new_n25885_), .B(new_n25705_), .ZN(new_n25886_));
  INV_X1     g25819(.I(new_n25705_), .ZN(new_n25887_));
  AOI21_X1   g25820(.A1(new_n25884_), .A2(new_n25883_), .B(new_n25710_), .ZN(new_n25888_));
  NOR3_X1    g25821(.A1(new_n25881_), .A2(new_n25873_), .A3(new_n25711_), .ZN(new_n25889_));
  NOR3_X1    g25822(.A1(new_n25889_), .A2(new_n25888_), .A3(new_n25887_), .ZN(new_n25890_));
  NOR2_X1    g25823(.A1(new_n25890_), .A2(new_n25886_), .ZN(new_n25891_));
  XNOR2_X1   g25824(.A1(new_n25891_), .A2(new_n25701_), .ZN(new_n25892_));
  INV_X1     g25825(.I(new_n25445_), .ZN(new_n25893_));
  NAND4_X1   g25826(.A1(new_n25230_), .A2(new_n25240_), .A3(new_n25893_), .A4(new_n25681_), .ZN(new_n25894_));
  XOR2_X1    g25827(.A1(new_n25894_), .A2(new_n25892_), .Z(new_n25895_));
  XOR2_X1    g25828(.A1(new_n25895_), .A2(new_n25697_), .Z(\result[10] ));
  XOR2_X1    g25829(.A1(new_n25697_), .A2(new_n25892_), .Z(new_n25897_));
  INV_X1     g25830(.I(new_n25897_), .ZN(new_n25898_));
  NOR4_X1    g25831(.A1(new_n25241_), .A2(new_n25445_), .A3(new_n25680_), .A4(new_n25898_), .ZN(new_n25899_));
  NAND2_X1   g25832(.A1(new_n25705_), .A2(new_n25710_), .ZN(new_n25900_));
  OAI21_X1   g25833(.A1(new_n25882_), .A2(new_n25705_), .B(new_n25900_), .ZN(new_n25901_));
  AOI22_X1   g25834(.A1(new_n24620_), .A2(new_n6789_), .B1(new_n7530_), .B2(new_n24386_), .ZN(new_n25902_));
  NOR2_X1    g25835(.A1(new_n24835_), .A2(new_n6785_), .ZN(new_n25903_));
  OAI21_X1   g25836(.A1(new_n25903_), .A2(new_n25902_), .B(new_n6775_), .ZN(new_n25904_));
  INV_X1     g25837(.I(new_n25904_), .ZN(new_n25905_));
  NAND2_X1   g25838(.A1(new_n24833_), .A2(new_n25905_), .ZN(new_n25906_));
  NOR2_X1    g25839(.A1(new_n25906_), .A2(\a[8] ), .ZN(new_n25907_));
  AOI21_X1   g25840(.A1(new_n24833_), .A2(new_n25905_), .B(new_n4009_), .ZN(new_n25908_));
  NOR2_X1    g25841(.A1(new_n25907_), .A2(new_n25908_), .ZN(new_n25909_));
  OAI22_X1   g25842(.A1(new_n23948_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n22149_), .ZN(new_n25910_));
  NAND2_X1   g25843(.A1(new_n24174_), .A2(new_n4709_), .ZN(new_n25911_));
  AOI21_X1   g25844(.A1(new_n25911_), .A2(new_n25910_), .B(new_n4707_), .ZN(new_n25912_));
  NAND2_X1   g25845(.A1(new_n24172_), .A2(new_n25912_), .ZN(new_n25913_));
  XOR2_X1    g25846(.A1(new_n25913_), .A2(\a[11] ), .Z(new_n25914_));
  INV_X1     g25847(.I(new_n25914_), .ZN(new_n25915_));
  AOI22_X1   g25848(.A1(new_n22048_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n21953_), .ZN(new_n25916_));
  NOR2_X1    g25849(.A1(new_n22115_), .A2(new_n6091_), .ZN(new_n25917_));
  OAI21_X1   g25850(.A1(new_n25917_), .A2(new_n25916_), .B(new_n6081_), .ZN(new_n25918_));
  NOR2_X1    g25851(.A1(new_n23675_), .A2(new_n25918_), .ZN(new_n25919_));
  XOR2_X1    g25852(.A1(new_n25919_), .A2(new_n3521_), .Z(new_n25920_));
  NOR2_X1    g25853(.A1(new_n25814_), .A2(new_n25720_), .ZN(new_n25921_));
  OAI21_X1   g25854(.A1(new_n25817_), .A2(new_n25816_), .B(new_n25714_), .ZN(new_n25922_));
  NAND3_X1   g25855(.A1(new_n25805_), .A2(new_n25809_), .A3(new_n25715_), .ZN(new_n25923_));
  AOI21_X1   g25856(.A1(new_n25922_), .A2(new_n25923_), .B(new_n25822_), .ZN(new_n25924_));
  AOI21_X1   g25857(.A1(new_n25924_), .A2(new_n25814_), .B(new_n25921_), .ZN(new_n25925_));
  INV_X1     g25858(.I(new_n19521_), .ZN(new_n25926_));
  AOI22_X1   g25859(.A1(new_n21157_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n19484_), .ZN(new_n25927_));
  NOR2_X1    g25860(.A1(new_n19512_), .A2(new_n4470_), .ZN(new_n25928_));
  OAI21_X1   g25861(.A1(new_n25928_), .A2(new_n25927_), .B(new_n4295_), .ZN(new_n25929_));
  NOR2_X1    g25862(.A1(new_n25926_), .A2(new_n25929_), .ZN(new_n25930_));
  NAND2_X1   g25863(.A1(new_n25930_), .A2(new_n3372_), .ZN(new_n25931_));
  NOR2_X1    g25864(.A1(new_n25930_), .A2(new_n3372_), .ZN(new_n25932_));
  INV_X1     g25865(.I(new_n25932_), .ZN(new_n25933_));
  NAND2_X1   g25866(.A1(new_n25933_), .A2(new_n25931_), .ZN(new_n25934_));
  OAI22_X1   g25867(.A1(new_n19428_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19423_), .ZN(new_n25935_));
  NAND2_X1   g25868(.A1(new_n19438_), .A2(new_n3312_), .ZN(new_n25936_));
  AOI21_X1   g25869(.A1(new_n25936_), .A2(new_n25935_), .B(new_n3302_), .ZN(new_n25937_));
  NAND2_X1   g25870(.A1(new_n20907_), .A2(new_n25937_), .ZN(new_n25938_));
  XOR2_X1    g25871(.A1(new_n25938_), .A2(\a[23] ), .Z(new_n25939_));
  OAI22_X1   g25872(.A1(new_n19410_), .A2(new_n3268_), .B1(new_n19412_), .B2(new_n3322_), .ZN(new_n25940_));
  NAND2_X1   g25873(.A1(new_n19439_), .A2(new_n3317_), .ZN(new_n25941_));
  AOI21_X1   g25874(.A1(new_n25941_), .A2(new_n25940_), .B(new_n3260_), .ZN(new_n25942_));
  NAND2_X1   g25875(.A1(new_n20827_), .A2(new_n25942_), .ZN(new_n25943_));
  XOR2_X1    g25876(.A1(new_n25943_), .A2(\a[26] ), .Z(new_n25944_));
  INV_X1     g25877(.I(new_n25944_), .ZN(new_n25945_));
  NAND2_X1   g25878(.A1(new_n25778_), .A2(new_n25740_), .ZN(new_n25946_));
  NOR2_X1    g25879(.A1(new_n25778_), .A2(new_n25740_), .ZN(new_n25947_));
  AOI21_X1   g25880(.A1(new_n25748_), .A2(new_n25946_), .B(new_n25947_), .ZN(new_n25948_));
  INV_X1     g25881(.I(new_n25774_), .ZN(new_n25949_));
  OAI21_X1   g25882(.A1(new_n25751_), .A2(new_n25949_), .B(new_n25775_), .ZN(new_n25950_));
  NAND2_X1   g25883(.A1(new_n25765_), .A2(new_n25095_), .ZN(new_n25951_));
  NAND2_X1   g25884(.A1(new_n25951_), .A2(new_n25766_), .ZN(new_n25952_));
  INV_X1     g25885(.I(new_n25952_), .ZN(new_n25953_));
  NAND2_X1   g25886(.A1(new_n17794_), .A2(new_n3332_), .ZN(new_n25954_));
  NAND2_X1   g25887(.A1(new_n19386_), .A2(new_n3189_), .ZN(new_n25955_));
  AOI21_X1   g25888(.A1(new_n20127_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n25956_));
  NAND4_X1   g25889(.A1(new_n21632_), .A2(new_n25954_), .A3(new_n25955_), .A4(new_n25956_), .ZN(new_n25957_));
  NAND4_X1   g25890(.A1(new_n4576_), .A2(new_n1097_), .A3(new_n1549_), .A4(new_n2479_), .ZN(new_n25958_));
  INV_X1     g25891(.I(new_n1235_), .ZN(new_n25959_));
  NOR4_X1    g25892(.A1(new_n866_), .A2(new_n560_), .A3(new_n561_), .A4(new_n92_), .ZN(new_n25960_));
  NOR4_X1    g25893(.A1(new_n25960_), .A2(new_n25959_), .A3(new_n3470_), .A4(new_n642_), .ZN(new_n25961_));
  INV_X1     g25894(.I(new_n25961_), .ZN(new_n25962_));
  NOR4_X1    g25895(.A1(new_n4851_), .A2(new_n25958_), .A3(new_n25962_), .A4(new_n2536_), .ZN(new_n25963_));
  INV_X1     g25896(.I(new_n25963_), .ZN(new_n25964_));
  NOR4_X1    g25897(.A1(new_n2976_), .A2(new_n2291_), .A3(new_n769_), .A4(new_n1417_), .ZN(new_n25965_));
  NAND3_X1   g25898(.A1(new_n25965_), .A2(new_n1148_), .A3(new_n4892_), .ZN(new_n25966_));
  NAND2_X1   g25899(.A1(new_n2213_), .A2(new_n706_), .ZN(new_n25967_));
  NOR4_X1    g25900(.A1(new_n25967_), .A2(new_n752_), .A3(new_n801_), .A4(new_n607_), .ZN(new_n25968_));
  NAND4_X1   g25901(.A1(new_n358_), .A2(new_n2178_), .A3(new_n1816_), .A4(new_n1706_), .ZN(new_n25969_));
  NAND3_X1   g25902(.A1(new_n25968_), .A2(new_n3008_), .A3(new_n25969_), .ZN(new_n25970_));
  NOR4_X1    g25903(.A1(new_n25964_), .A2(new_n1406_), .A3(new_n25970_), .A4(new_n25966_), .ZN(new_n25971_));
  NAND2_X1   g25904(.A1(new_n25971_), .A2(new_n942_), .ZN(new_n25972_));
  INV_X1     g25905(.I(new_n25972_), .ZN(new_n25973_));
  XOR2_X1    g25906(.A1(new_n25957_), .A2(new_n25973_), .Z(new_n25974_));
  NOR2_X1    g25907(.A1(new_n25974_), .A2(new_n25953_), .ZN(new_n25975_));
  XOR2_X1    g25908(.A1(new_n25957_), .A2(new_n25973_), .Z(new_n25976_));
  AOI21_X1   g25909(.A1(new_n25953_), .A2(new_n25976_), .B(new_n25975_), .ZN(new_n25977_));
  OAI22_X1   g25910(.A1(new_n19400_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19393_), .ZN(new_n25978_));
  NAND2_X1   g25911(.A1(new_n17790_), .A2(new_n2750_), .ZN(new_n25979_));
  AOI21_X1   g25912(.A1(new_n25979_), .A2(new_n25978_), .B(new_n2737_), .ZN(new_n25980_));
  NAND2_X1   g25913(.A1(new_n20251_), .A2(new_n25980_), .ZN(new_n25981_));
  XOR2_X1    g25914(.A1(new_n25981_), .A2(\a[29] ), .Z(new_n25982_));
  XOR2_X1    g25915(.A1(new_n25982_), .A2(new_n25977_), .Z(new_n25983_));
  AND2_X2    g25916(.A1(new_n25983_), .A2(new_n25950_), .Z(new_n25984_));
  NAND2_X1   g25917(.A1(new_n25982_), .A2(new_n25977_), .ZN(new_n25985_));
  OR2_X2     g25918(.A1(new_n25982_), .A2(new_n25977_), .Z(new_n25986_));
  AOI21_X1   g25919(.A1(new_n25986_), .A2(new_n25985_), .B(new_n25950_), .ZN(new_n25987_));
  NOR2_X1    g25920(.A1(new_n25984_), .A2(new_n25987_), .ZN(new_n25988_));
  XOR2_X1    g25921(.A1(new_n25988_), .A2(new_n25948_), .Z(new_n25989_));
  NOR2_X1    g25922(.A1(new_n25782_), .A2(new_n25736_), .ZN(new_n25990_));
  INV_X1     g25923(.I(new_n25990_), .ZN(new_n25991_));
  NOR2_X1    g25924(.A1(new_n25783_), .A2(new_n25791_), .ZN(new_n25992_));
  XOR2_X1    g25925(.A1(new_n25779_), .A2(new_n25741_), .Z(new_n25993_));
  OAI21_X1   g25926(.A1(new_n25993_), .A2(new_n25992_), .B(new_n25991_), .ZN(new_n25994_));
  NAND2_X1   g25927(.A1(new_n25994_), .A2(new_n25989_), .ZN(new_n25995_));
  NOR2_X1    g25928(.A1(new_n25994_), .A2(new_n25989_), .ZN(new_n25996_));
  INV_X1     g25929(.I(new_n25996_), .ZN(new_n25997_));
  AOI21_X1   g25930(.A1(new_n25997_), .A2(new_n25995_), .B(new_n25945_), .ZN(new_n25998_));
  INV_X1     g25931(.I(new_n25995_), .ZN(new_n25999_));
  NOR3_X1    g25932(.A1(new_n25999_), .A2(new_n25996_), .A3(new_n25944_), .ZN(new_n26000_));
  OAI21_X1   g25933(.A1(new_n25998_), .A2(new_n26000_), .B(new_n25939_), .ZN(new_n26001_));
  INV_X1     g25934(.I(new_n25939_), .ZN(new_n26002_));
  OAI21_X1   g25935(.A1(new_n25999_), .A2(new_n25996_), .B(new_n25944_), .ZN(new_n26003_));
  NAND3_X1   g25936(.A1(new_n25997_), .A2(new_n25995_), .A3(new_n25945_), .ZN(new_n26004_));
  NAND3_X1   g25937(.A1(new_n26003_), .A2(new_n26004_), .A3(new_n26002_), .ZN(new_n26005_));
  NAND2_X1   g25938(.A1(new_n26001_), .A2(new_n26005_), .ZN(new_n26006_));
  NOR2_X1    g25939(.A1(new_n25799_), .A2(new_n25798_), .ZN(new_n26007_));
  NAND2_X1   g25940(.A1(new_n25796_), .A2(new_n25731_), .ZN(new_n26008_));
  INV_X1     g25941(.I(new_n26008_), .ZN(new_n26009_));
  NAND2_X1   g25942(.A1(new_n25795_), .A2(new_n25730_), .ZN(new_n26010_));
  AOI21_X1   g25943(.A1(new_n26007_), .A2(new_n26010_), .B(new_n26009_), .ZN(new_n26011_));
  OAI22_X1   g25944(.A1(new_n19463_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19437_), .ZN(new_n26012_));
  NAND2_X1   g25945(.A1(new_n17780_), .A2(new_n4096_), .ZN(new_n26013_));
  AOI21_X1   g25946(.A1(new_n26012_), .A2(new_n26013_), .B(new_n4095_), .ZN(new_n26014_));
  NAND2_X1   g25947(.A1(new_n21088_), .A2(new_n26014_), .ZN(new_n26015_));
  XOR2_X1    g25948(.A1(new_n26015_), .A2(\a[20] ), .Z(new_n26016_));
  NAND2_X1   g25949(.A1(new_n26011_), .A2(new_n26016_), .ZN(new_n26017_));
  INV_X1     g25950(.I(new_n26017_), .ZN(new_n26018_));
  NOR2_X1    g25951(.A1(new_n26011_), .A2(new_n26016_), .ZN(new_n26019_));
  OAI21_X1   g25952(.A1(new_n26018_), .A2(new_n26019_), .B(new_n26006_), .ZN(new_n26020_));
  AOI21_X1   g25953(.A1(new_n26003_), .A2(new_n26004_), .B(new_n26002_), .ZN(new_n26021_));
  NOR3_X1    g25954(.A1(new_n25998_), .A2(new_n26000_), .A3(new_n25939_), .ZN(new_n26022_));
  NOR2_X1    g25955(.A1(new_n26021_), .A2(new_n26022_), .ZN(new_n26023_));
  INV_X1     g25956(.I(new_n26016_), .ZN(new_n26024_));
  NOR2_X1    g25957(.A1(new_n26011_), .A2(new_n26024_), .ZN(new_n26025_));
  NAND2_X1   g25958(.A1(new_n26011_), .A2(new_n26024_), .ZN(new_n26026_));
  INV_X1     g25959(.I(new_n26026_), .ZN(new_n26027_));
  OAI21_X1   g25960(.A1(new_n26027_), .A2(new_n26025_), .B(new_n26023_), .ZN(new_n26028_));
  NOR2_X1    g25961(.A1(new_n25714_), .A2(new_n25725_), .ZN(new_n26029_));
  INV_X1     g25962(.I(new_n26029_), .ZN(new_n26030_));
  NOR2_X1    g25963(.A1(new_n25715_), .A2(new_n25806_), .ZN(new_n26031_));
  INV_X1     g25964(.I(new_n26010_), .ZN(new_n26032_));
  OAI22_X1   g25965(.A1(new_n25799_), .A2(new_n25798_), .B1(new_n26009_), .B2(new_n26032_), .ZN(new_n26033_));
  XOR2_X1    g25966(.A1(new_n25795_), .A2(new_n25730_), .Z(new_n26034_));
  NAND2_X1   g25967(.A1(new_n26007_), .A2(new_n26034_), .ZN(new_n26035_));
  NAND2_X1   g25968(.A1(new_n26035_), .A2(new_n26033_), .ZN(new_n26036_));
  OAI21_X1   g25969(.A1(new_n26036_), .A2(new_n26031_), .B(new_n26030_), .ZN(new_n26037_));
  NAND3_X1   g25970(.A1(new_n26028_), .A2(new_n26020_), .A3(new_n26037_), .ZN(new_n26038_));
  INV_X1     g25971(.I(new_n26019_), .ZN(new_n26039_));
  AOI21_X1   g25972(.A1(new_n26039_), .A2(new_n26017_), .B(new_n26023_), .ZN(new_n26040_));
  INV_X1     g25973(.I(new_n26025_), .ZN(new_n26041_));
  AOI21_X1   g25974(.A1(new_n26041_), .A2(new_n26026_), .B(new_n26006_), .ZN(new_n26042_));
  INV_X1     g25975(.I(new_n26037_), .ZN(new_n26043_));
  OAI21_X1   g25976(.A1(new_n26040_), .A2(new_n26042_), .B(new_n26043_), .ZN(new_n26044_));
  AOI21_X1   g25977(.A1(new_n26044_), .A2(new_n26038_), .B(new_n25934_), .ZN(new_n26045_));
  INV_X1     g25978(.I(new_n25934_), .ZN(new_n26046_));
  NOR3_X1    g25979(.A1(new_n26040_), .A2(new_n26042_), .A3(new_n26043_), .ZN(new_n26047_));
  AOI21_X1   g25980(.A1(new_n26028_), .A2(new_n26020_), .B(new_n26037_), .ZN(new_n26048_));
  NOR3_X1    g25981(.A1(new_n26048_), .A2(new_n26047_), .A3(new_n26046_), .ZN(new_n26049_));
  OAI21_X1   g25982(.A1(new_n26049_), .A2(new_n26045_), .B(new_n25925_), .ZN(new_n26050_));
  INV_X1     g25983(.I(new_n25925_), .ZN(new_n26051_));
  OAI21_X1   g25984(.A1(new_n26048_), .A2(new_n26047_), .B(new_n26046_), .ZN(new_n26052_));
  NAND3_X1   g25985(.A1(new_n26044_), .A2(new_n26038_), .A3(new_n25934_), .ZN(new_n26053_));
  NAND3_X1   g25986(.A1(new_n26051_), .A2(new_n26052_), .A3(new_n26053_), .ZN(new_n26054_));
  NAND2_X1   g25987(.A1(new_n26054_), .A2(new_n26050_), .ZN(new_n26055_));
  NOR2_X1    g25988(.A1(new_n25865_), .A2(new_n25600_), .ZN(new_n26056_));
  NOR2_X1    g25989(.A1(new_n26056_), .A2(new_n25866_), .ZN(new_n26057_));
  NOR2_X1    g25990(.A1(new_n26057_), .A2(new_n25835_), .ZN(new_n26058_));
  NAND2_X1   g25991(.A1(new_n26057_), .A2(new_n25835_), .ZN(new_n26059_));
  AOI21_X1   g25992(.A1(new_n25830_), .A2(new_n26059_), .B(new_n26058_), .ZN(new_n26060_));
  NOR2_X1    g25993(.A1(new_n26060_), .A2(new_n26055_), .ZN(new_n26061_));
  AOI21_X1   g25994(.A1(new_n26052_), .A2(new_n26053_), .B(new_n26051_), .ZN(new_n26062_));
  NOR3_X1    g25995(.A1(new_n26049_), .A2(new_n26045_), .A3(new_n25925_), .ZN(new_n26063_));
  NOR2_X1    g25996(.A1(new_n26062_), .A2(new_n26063_), .ZN(new_n26064_));
  INV_X1     g25997(.I(new_n26058_), .ZN(new_n26065_));
  NAND3_X1   g25998(.A1(new_n25859_), .A2(new_n25860_), .A3(new_n26059_), .ZN(new_n26066_));
  NAND2_X1   g25999(.A1(new_n26066_), .A2(new_n26065_), .ZN(new_n26067_));
  NOR2_X1    g26000(.A1(new_n26064_), .A2(new_n26067_), .ZN(new_n26068_));
  OAI21_X1   g26001(.A1(new_n26061_), .A2(new_n26068_), .B(new_n25920_), .ZN(new_n26069_));
  INV_X1     g26002(.I(new_n25920_), .ZN(new_n26070_));
  NAND2_X1   g26003(.A1(new_n26064_), .A2(new_n26067_), .ZN(new_n26071_));
  NAND3_X1   g26004(.A1(new_n26055_), .A2(new_n26065_), .A3(new_n26066_), .ZN(new_n26072_));
  NAND3_X1   g26005(.A1(new_n26071_), .A2(new_n26072_), .A3(new_n26070_), .ZN(new_n26073_));
  AOI21_X1   g26006(.A1(new_n26069_), .A2(new_n26073_), .B(new_n25915_), .ZN(new_n26074_));
  AOI21_X1   g26007(.A1(new_n26071_), .A2(new_n26072_), .B(new_n26070_), .ZN(new_n26075_));
  NOR3_X1    g26008(.A1(new_n26061_), .A2(new_n26068_), .A3(new_n25920_), .ZN(new_n26076_));
  NOR3_X1    g26009(.A1(new_n26076_), .A2(new_n26075_), .A3(new_n25914_), .ZN(new_n26077_));
  NOR2_X1    g26010(.A1(new_n25872_), .A2(new_n25852_), .ZN(new_n26078_));
  NAND2_X1   g26011(.A1(new_n25872_), .A2(new_n25852_), .ZN(new_n26079_));
  OAI21_X1   g26012(.A1(new_n25844_), .A2(new_n25847_), .B(new_n25830_), .ZN(new_n26080_));
  NAND3_X1   g26013(.A1(new_n25855_), .A2(new_n25861_), .A3(new_n25854_), .ZN(new_n26081_));
  NAND2_X1   g26014(.A1(new_n26080_), .A2(new_n26081_), .ZN(new_n26082_));
  AOI21_X1   g26015(.A1(new_n26082_), .A2(new_n26079_), .B(new_n26078_), .ZN(new_n26083_));
  NOR3_X1    g26016(.A1(new_n26074_), .A2(new_n26077_), .A3(new_n26083_), .ZN(new_n26084_));
  OAI21_X1   g26017(.A1(new_n26076_), .A2(new_n26075_), .B(new_n25914_), .ZN(new_n26085_));
  NAND3_X1   g26018(.A1(new_n26069_), .A2(new_n26073_), .A3(new_n25915_), .ZN(new_n26086_));
  INV_X1     g26019(.I(new_n26083_), .ZN(new_n26087_));
  AOI21_X1   g26020(.A1(new_n26085_), .A2(new_n26086_), .B(new_n26087_), .ZN(new_n26088_));
  OAI21_X1   g26021(.A1(new_n26084_), .A2(new_n26088_), .B(new_n25909_), .ZN(new_n26089_));
  INV_X1     g26022(.I(new_n25909_), .ZN(new_n26090_));
  NAND3_X1   g26023(.A1(new_n26085_), .A2(new_n26086_), .A3(new_n26087_), .ZN(new_n26091_));
  OAI21_X1   g26024(.A1(new_n26074_), .A2(new_n26077_), .B(new_n26083_), .ZN(new_n26092_));
  NAND3_X1   g26025(.A1(new_n26092_), .A2(new_n26091_), .A3(new_n26090_), .ZN(new_n26093_));
  AOI21_X1   g26026(.A1(new_n26089_), .A2(new_n26093_), .B(new_n25901_), .ZN(new_n26094_));
  INV_X1     g26027(.I(new_n25901_), .ZN(new_n26095_));
  AOI21_X1   g26028(.A1(new_n26092_), .A2(new_n26091_), .B(new_n26090_), .ZN(new_n26096_));
  NOR3_X1    g26029(.A1(new_n26084_), .A2(new_n26088_), .A3(new_n25909_), .ZN(new_n26097_));
  NOR3_X1    g26030(.A1(new_n26097_), .A2(new_n26096_), .A3(new_n26095_), .ZN(new_n26098_));
  NOR2_X1    g26031(.A1(new_n26098_), .A2(new_n26094_), .ZN(new_n26099_));
  OAI21_X1   g26032(.A1(new_n25697_), .A2(new_n25891_), .B(new_n25701_), .ZN(new_n26100_));
  XNOR2_X1   g26033(.A1(new_n26100_), .A2(new_n26099_), .ZN(new_n26101_));
  INV_X1     g26034(.I(new_n26101_), .ZN(new_n26102_));
  XOR2_X1    g26035(.A1(new_n25899_), .A2(new_n26102_), .Z(\result[11] ));
  NAND2_X1   g26036(.A1(new_n25899_), .A2(new_n26102_), .ZN(new_n26104_));
  NOR2_X1    g26037(.A1(new_n25891_), .A2(new_n25701_), .ZN(new_n26105_));
  INV_X1     g26038(.I(new_n26105_), .ZN(new_n26106_));
  NOR3_X1    g26039(.A1(new_n26098_), .A2(new_n26094_), .A3(new_n26105_), .ZN(new_n26107_));
  OAI21_X1   g26040(.A1(new_n25697_), .A2(new_n26106_), .B(new_n26107_), .ZN(new_n26108_));
  NOR2_X1    g26041(.A1(new_n26074_), .A2(new_n26077_), .ZN(new_n26109_));
  XOR2_X1    g26042(.A1(new_n26083_), .A2(new_n25909_), .Z(new_n26110_));
  OR2_X2     g26043(.A1(new_n26110_), .A2(new_n26109_), .Z(new_n26111_));
  NAND2_X1   g26044(.A1(new_n26110_), .A2(new_n26109_), .ZN(new_n26112_));
  NAND3_X1   g26045(.A1(new_n26111_), .A2(new_n26112_), .A3(new_n26095_), .ZN(new_n26113_));
  OAI22_X1   g26046(.A1(new_n19475_), .A2(new_n3775_), .B1(new_n19463_), .B2(new_n3769_), .ZN(new_n26114_));
  NAND2_X1   g26047(.A1(new_n19484_), .A2(new_n4096_), .ZN(new_n26115_));
  AOI21_X1   g26048(.A1(new_n26115_), .A2(new_n26114_), .B(new_n4095_), .ZN(new_n26116_));
  NAND2_X1   g26049(.A1(new_n21171_), .A2(new_n26116_), .ZN(new_n26117_));
  XOR2_X1    g26050(.A1(new_n26117_), .A2(\a[20] ), .Z(new_n26118_));
  OAI22_X1   g26051(.A1(new_n17784_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19428_), .ZN(new_n26119_));
  NAND2_X1   g26052(.A1(new_n19466_), .A2(new_n3312_), .ZN(new_n26120_));
  AOI21_X1   g26053(.A1(new_n26120_), .A2(new_n26119_), .B(new_n3302_), .ZN(new_n26121_));
  NAND2_X1   g26054(.A1(new_n21100_), .A2(new_n26121_), .ZN(new_n26122_));
  XOR2_X1    g26055(.A1(new_n26122_), .A2(\a[23] ), .Z(new_n26123_));
  INV_X1     g26056(.I(new_n26123_), .ZN(new_n26124_));
  OAI22_X1   g26057(.A1(new_n17787_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19412_), .ZN(new_n26125_));
  NAND2_X1   g26058(.A1(new_n19442_), .A2(new_n3317_), .ZN(new_n26126_));
  AOI21_X1   g26059(.A1(new_n26126_), .A2(new_n26125_), .B(new_n3260_), .ZN(new_n26127_));
  NAND2_X1   g26060(.A1(new_n20939_), .A2(new_n26127_), .ZN(new_n26128_));
  XOR2_X1    g26061(.A1(new_n26128_), .A2(\a[26] ), .Z(new_n26129_));
  INV_X1     g26062(.I(new_n26129_), .ZN(new_n26130_));
  OAI22_X1   g26063(.A1(new_n17789_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19400_), .ZN(new_n26131_));
  NAND2_X1   g26064(.A1(new_n19407_), .A2(new_n2750_), .ZN(new_n26132_));
  AOI21_X1   g26065(.A1(new_n26132_), .A2(new_n26131_), .B(new_n2737_), .ZN(new_n26133_));
  NAND2_X1   g26066(.A1(new_n20864_), .A2(new_n26133_), .ZN(new_n26134_));
  XOR2_X1    g26067(.A1(new_n26134_), .A2(\a[29] ), .Z(new_n26135_));
  NAND2_X1   g26068(.A1(new_n25985_), .A2(new_n25950_), .ZN(new_n26136_));
  NAND2_X1   g26069(.A1(new_n26136_), .A2(new_n25986_), .ZN(new_n26137_));
  NOR2_X1    g26070(.A1(new_n437_), .A2(new_n506_), .ZN(new_n26138_));
  NOR4_X1    g26071(.A1(new_n90_), .A2(new_n255_), .A3(new_n1031_), .A4(new_n902_), .ZN(new_n26139_));
  NAND4_X1   g26072(.A1(new_n26139_), .A2(new_n922_), .A3(new_n655_), .A4(new_n26138_), .ZN(new_n26140_));
  NOR2_X1    g26073(.A1(new_n3220_), .A2(new_n1730_), .ZN(new_n26141_));
  NAND4_X1   g26074(.A1(new_n26141_), .A2(new_n1606_), .A3(new_n2478_), .A4(new_n2444_), .ZN(new_n26142_));
  NOR4_X1    g26075(.A1(new_n26142_), .A2(new_n1552_), .A3(new_n12266_), .A4(new_n26140_), .ZN(new_n26143_));
  NOR4_X1    g26076(.A1(new_n482_), .A2(new_n698_), .A3(new_n721_), .A4(new_n640_), .ZN(new_n26144_));
  NOR2_X1    g26077(.A1(new_n124_), .A2(new_n682_), .ZN(new_n26145_));
  NAND4_X1   g26078(.A1(new_n26145_), .A2(new_n992_), .A3(new_n408_), .A4(new_n325_), .ZN(new_n26146_));
  NOR2_X1    g26079(.A1(new_n26146_), .A2(new_n26144_), .ZN(new_n26147_));
  INV_X1     g26080(.I(new_n10984_), .ZN(new_n26148_));
  NOR4_X1    g26081(.A1(new_n238_), .A2(new_n603_), .A3(new_n553_), .A4(new_n456_), .ZN(new_n26149_));
  NOR4_X1    g26082(.A1(new_n740_), .A2(new_n670_), .A3(new_n783_), .A4(new_n330_), .ZN(new_n26150_));
  NOR4_X1    g26083(.A1(new_n26148_), .A2(new_n4937_), .A3(new_n26149_), .A4(new_n26150_), .ZN(new_n26151_));
  NAND3_X1   g26084(.A1(new_n26151_), .A2(new_n26147_), .A3(new_n2926_), .ZN(new_n26152_));
  NOR2_X1    g26085(.A1(new_n26152_), .A2(new_n2853_), .ZN(new_n26153_));
  NAND3_X1   g26086(.A1(new_n26153_), .A2(new_n11474_), .A3(new_n26143_), .ZN(new_n26154_));
  XOR2_X1    g26087(.A1(new_n25952_), .A2(new_n25972_), .Z(new_n26155_));
  OAI21_X1   g26088(.A1(new_n25957_), .A2(new_n25952_), .B(new_n26155_), .ZN(new_n26156_));
  AOI21_X1   g26089(.A1(new_n25952_), .A2(new_n25957_), .B(new_n26156_), .ZN(new_n26157_));
  XOR2_X1    g26090(.A1(new_n26157_), .A2(new_n26154_), .Z(new_n26158_));
  NAND2_X1   g26091(.A1(new_n19394_), .A2(new_n3332_), .ZN(new_n26159_));
  NAND2_X1   g26092(.A1(new_n17794_), .A2(new_n3189_), .ZN(new_n26160_));
  AOI21_X1   g26093(.A1(new_n19386_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n26161_));
  NAND4_X1   g26094(.A1(new_n20291_), .A2(new_n26159_), .A3(new_n26160_), .A4(new_n26161_), .ZN(new_n26162_));
  XOR2_X1    g26095(.A1(new_n26158_), .A2(new_n26162_), .Z(new_n26163_));
  XOR2_X1    g26096(.A1(new_n26137_), .A2(new_n26163_), .Z(new_n26164_));
  XOR2_X1    g26097(.A1(new_n26164_), .A2(new_n26135_), .Z(new_n26165_));
  XOR2_X1    g26098(.A1(new_n26165_), .A2(new_n26130_), .Z(new_n26166_));
  INV_X1     g26099(.I(new_n25988_), .ZN(new_n26167_));
  AOI21_X1   g26100(.A1(new_n26167_), .A2(new_n25944_), .B(new_n25948_), .ZN(new_n26168_));
  NOR2_X1    g26101(.A1(new_n26167_), .A2(new_n25944_), .ZN(new_n26169_));
  NOR2_X1    g26102(.A1(new_n26168_), .A2(new_n26169_), .ZN(new_n26170_));
  XOR2_X1    g26103(.A1(new_n26166_), .A2(new_n26170_), .Z(new_n26171_));
  INV_X1     g26104(.I(new_n25994_), .ZN(new_n26172_));
  NOR2_X1    g26105(.A1(new_n26172_), .A2(new_n25939_), .ZN(new_n26173_));
  NAND2_X1   g26106(.A1(new_n26172_), .A2(new_n25939_), .ZN(new_n26174_));
  XOR2_X1    g26107(.A1(new_n25989_), .A2(new_n25944_), .Z(new_n26175_));
  AOI21_X1   g26108(.A1(new_n26175_), .A2(new_n26174_), .B(new_n26173_), .ZN(new_n26176_));
  XOR2_X1    g26109(.A1(new_n26171_), .A2(new_n26176_), .Z(new_n26177_));
  NOR2_X1    g26110(.A1(new_n26177_), .A2(new_n26124_), .ZN(new_n26178_));
  INV_X1     g26111(.I(new_n26170_), .ZN(new_n26179_));
  XOR2_X1    g26112(.A1(new_n26166_), .A2(new_n26179_), .Z(new_n26180_));
  XOR2_X1    g26113(.A1(new_n26180_), .A2(new_n26176_), .Z(new_n26181_));
  NOR2_X1    g26114(.A1(new_n26181_), .A2(new_n26123_), .ZN(new_n26182_));
  OAI21_X1   g26115(.A1(new_n26178_), .A2(new_n26182_), .B(new_n26118_), .ZN(new_n26183_));
  INV_X1     g26116(.I(new_n26118_), .ZN(new_n26184_));
  NAND2_X1   g26117(.A1(new_n26181_), .A2(new_n26123_), .ZN(new_n26185_));
  NAND2_X1   g26118(.A1(new_n26177_), .A2(new_n26124_), .ZN(new_n26186_));
  NAND3_X1   g26119(.A1(new_n26185_), .A2(new_n26186_), .A3(new_n26184_), .ZN(new_n26187_));
  OAI21_X1   g26120(.A1(new_n26023_), .A2(new_n26018_), .B(new_n26039_), .ZN(new_n26188_));
  OAI22_X1   g26121(.A1(new_n19512_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n19522_), .ZN(new_n26189_));
  NAND2_X1   g26122(.A1(new_n21953_), .A2(new_n4469_), .ZN(new_n26190_));
  AOI21_X1   g26123(.A1(new_n26189_), .A2(new_n26190_), .B(new_n4468_), .ZN(new_n26191_));
  NAND2_X1   g26124(.A1(new_n21963_), .A2(new_n26191_), .ZN(new_n26192_));
  NOR2_X1    g26125(.A1(new_n26192_), .A2(\a[17] ), .ZN(new_n26193_));
  AOI21_X1   g26126(.A1(new_n21963_), .A2(new_n26191_), .B(new_n3372_), .ZN(new_n26194_));
  NOR2_X1    g26127(.A1(new_n26193_), .A2(new_n26194_), .ZN(new_n26195_));
  INV_X1     g26128(.I(new_n26195_), .ZN(new_n26196_));
  OR2_X2     g26129(.A1(new_n26188_), .A2(new_n26196_), .Z(new_n26197_));
  NAND2_X1   g26130(.A1(new_n26188_), .A2(new_n26196_), .ZN(new_n26198_));
  AOI22_X1   g26131(.A1(new_n26183_), .A2(new_n26187_), .B1(new_n26197_), .B2(new_n26198_), .ZN(new_n26199_));
  NAND2_X1   g26132(.A1(new_n26183_), .A2(new_n26187_), .ZN(new_n26200_));
  XOR2_X1    g26133(.A1(new_n26188_), .A2(new_n26195_), .Z(new_n26201_));
  NOR2_X1    g26134(.A1(new_n26200_), .A2(new_n26201_), .ZN(new_n26202_));
  NOR2_X1    g26135(.A1(new_n26040_), .A2(new_n26042_), .ZN(new_n26203_));
  NOR2_X1    g26136(.A1(new_n26037_), .A2(new_n25934_), .ZN(new_n26204_));
  NAND2_X1   g26137(.A1(new_n26037_), .A2(new_n25934_), .ZN(new_n26205_));
  OAI21_X1   g26138(.A1(new_n26203_), .A2(new_n26204_), .B(new_n26205_), .ZN(new_n26206_));
  OAI22_X1   g26139(.A1(new_n22115_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n22051_), .ZN(new_n26207_));
  NAND2_X1   g26140(.A1(new_n22150_), .A2(new_n6090_), .ZN(new_n26208_));
  AOI21_X1   g26141(.A1(new_n26207_), .A2(new_n26208_), .B(new_n6082_), .ZN(new_n26209_));
  NAND2_X1   g26142(.A1(new_n22163_), .A2(new_n26209_), .ZN(new_n26210_));
  XOR2_X1    g26143(.A1(new_n26210_), .A2(new_n3521_), .Z(new_n26211_));
  NOR2_X1    g26144(.A1(new_n26211_), .A2(new_n26206_), .ZN(new_n26212_));
  NAND2_X1   g26145(.A1(new_n26211_), .A2(new_n26206_), .ZN(new_n26213_));
  INV_X1     g26146(.I(new_n26213_), .ZN(new_n26214_));
  OAI22_X1   g26147(.A1(new_n26202_), .A2(new_n26199_), .B1(new_n26214_), .B2(new_n26212_), .ZN(new_n26215_));
  NOR2_X1    g26148(.A1(new_n26202_), .A2(new_n26199_), .ZN(new_n26216_));
  XOR2_X1    g26149(.A1(new_n26211_), .A2(new_n26206_), .Z(new_n26217_));
  NAND2_X1   g26150(.A1(new_n26216_), .A2(new_n26217_), .ZN(new_n26218_));
  NAND2_X1   g26151(.A1(new_n26218_), .A2(new_n26215_), .ZN(new_n26219_));
  INV_X1     g26152(.I(new_n26203_), .ZN(new_n26220_));
  NOR2_X1    g26153(.A1(new_n26043_), .A2(new_n26046_), .ZN(new_n26221_));
  OAI21_X1   g26154(.A1(new_n26204_), .A2(new_n26221_), .B(new_n26220_), .ZN(new_n26222_));
  XNOR2_X1   g26155(.A1(new_n26037_), .A2(new_n25934_), .ZN(new_n26223_));
  OAI21_X1   g26156(.A1(new_n26220_), .A2(new_n26223_), .B(new_n26222_), .ZN(new_n26224_));
  NAND2_X1   g26157(.A1(new_n25920_), .A2(new_n25925_), .ZN(new_n26225_));
  NOR2_X1    g26158(.A1(new_n25920_), .A2(new_n25925_), .ZN(new_n26226_));
  AOI21_X1   g26159(.A1(new_n26224_), .A2(new_n26225_), .B(new_n26226_), .ZN(new_n26227_));
  AOI22_X1   g26160(.A1(new_n24174_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n23957_), .ZN(new_n26228_));
  NOR2_X1    g26161(.A1(new_n24376_), .A2(new_n4710_), .ZN(new_n26229_));
  OAI21_X1   g26162(.A1(new_n26229_), .A2(new_n26228_), .B(new_n4706_), .ZN(new_n26230_));
  NOR3_X1    g26163(.A1(new_n24391_), .A2(\a[11] ), .A3(new_n26230_), .ZN(new_n26231_));
  INV_X1     g26164(.I(new_n26230_), .ZN(new_n26232_));
  AOI21_X1   g26165(.A1(new_n24390_), .A2(new_n26232_), .B(new_n4034_), .ZN(new_n26233_));
  NOR2_X1    g26166(.A1(new_n26231_), .A2(new_n26233_), .ZN(new_n26234_));
  XNOR2_X1   g26167(.A1(new_n26234_), .A2(new_n26227_), .ZN(new_n26235_));
  NAND2_X1   g26168(.A1(new_n26235_), .A2(new_n26219_), .ZN(new_n26236_));
  XNOR2_X1   g26169(.A1(new_n26227_), .A2(new_n26234_), .ZN(new_n26237_));
  OAI21_X1   g26170(.A1(new_n26219_), .A2(new_n26237_), .B(new_n26236_), .ZN(new_n26238_));
  INV_X1     g26171(.I(new_n26238_), .ZN(new_n26239_));
  NOR2_X1    g26172(.A1(new_n26060_), .A2(new_n25914_), .ZN(new_n26240_));
  NAND2_X1   g26173(.A1(new_n26064_), .A2(new_n26070_), .ZN(new_n26241_));
  NAND2_X1   g26174(.A1(new_n26055_), .A2(new_n25920_), .ZN(new_n26242_));
  AOI22_X1   g26175(.A1(new_n26241_), .A2(new_n26242_), .B1(new_n25914_), .B2(new_n26060_), .ZN(new_n26243_));
  AOI22_X1   g26176(.A1(new_n24826_), .A2(new_n12016_), .B1(new_n7530_), .B2(new_n24620_), .ZN(new_n26244_));
  OR3_X2     g26177(.A1(new_n25017_), .A2(new_n6776_), .A3(new_n26244_), .Z(new_n26245_));
  XOR2_X1    g26178(.A1(new_n26245_), .A2(\a[8] ), .Z(new_n26246_));
  NOR3_X1    g26179(.A1(new_n26243_), .A2(new_n26240_), .A3(new_n26246_), .ZN(new_n26247_));
  NOR2_X1    g26180(.A1(new_n26243_), .A2(new_n26240_), .ZN(new_n26248_));
  INV_X1     g26181(.I(new_n26246_), .ZN(new_n26249_));
  NOR2_X1    g26182(.A1(new_n26248_), .A2(new_n26249_), .ZN(new_n26250_));
  NOR2_X1    g26183(.A1(new_n26250_), .A2(new_n26247_), .ZN(new_n26251_));
  NOR2_X1    g26184(.A1(new_n26087_), .A2(new_n26090_), .ZN(new_n26252_));
  NOR2_X1    g26185(.A1(new_n26109_), .A2(new_n26252_), .ZN(new_n26253_));
  NOR2_X1    g26186(.A1(new_n26083_), .A2(new_n25909_), .ZN(new_n26254_));
  NOR2_X1    g26187(.A1(new_n26253_), .A2(new_n26254_), .ZN(new_n26255_));
  XOR2_X1    g26188(.A1(new_n26255_), .A2(new_n26251_), .Z(new_n26256_));
  NOR2_X1    g26189(.A1(new_n26256_), .A2(new_n26239_), .ZN(new_n26257_));
  XOR2_X1    g26190(.A1(new_n26255_), .A2(new_n26251_), .Z(new_n26258_));
  AOI21_X1   g26191(.A1(new_n26239_), .A2(new_n26258_), .B(new_n26257_), .ZN(new_n26259_));
  OR3_X2     g26192(.A1(new_n26259_), .A2(new_n26108_), .A3(new_n26113_), .Z(new_n26260_));
  OAI21_X1   g26193(.A1(new_n26108_), .A2(new_n26113_), .B(new_n26259_), .ZN(new_n26261_));
  NAND2_X1   g26194(.A1(new_n26260_), .A2(new_n26261_), .ZN(new_n26262_));
  INV_X1     g26195(.I(new_n26262_), .ZN(new_n26263_));
  XOR2_X1    g26196(.A1(new_n26104_), .A2(new_n26263_), .Z(\result[12] ));
  XOR2_X1    g26197(.A1(new_n25690_), .A2(new_n25667_), .Z(new_n26265_));
  NOR2_X1    g26198(.A1(new_n26265_), .A2(new_n25456_), .ZN(new_n26266_));
  AOI21_X1   g26199(.A1(new_n25449_), .A2(new_n26266_), .B(new_n25692_), .ZN(new_n26267_));
  OR3_X2     g26200(.A1(new_n26098_), .A2(new_n26094_), .A3(new_n26105_), .Z(new_n26268_));
  AOI21_X1   g26201(.A1(new_n26267_), .A2(new_n26105_), .B(new_n26268_), .ZN(new_n26269_));
  INV_X1     g26202(.I(new_n26255_), .ZN(new_n26270_));
  NOR2_X1    g26203(.A1(new_n26238_), .A2(new_n26251_), .ZN(new_n26271_));
  INV_X1     g26204(.I(new_n26271_), .ZN(new_n26272_));
  NAND2_X1   g26205(.A1(new_n26238_), .A2(new_n26251_), .ZN(new_n26273_));
  AOI21_X1   g26206(.A1(new_n26272_), .A2(new_n26273_), .B(new_n26270_), .ZN(new_n26274_));
  NAND3_X1   g26207(.A1(new_n26270_), .A2(new_n26272_), .A3(new_n26273_), .ZN(new_n26275_));
  INV_X1     g26208(.I(new_n26273_), .ZN(new_n26276_));
  OAI21_X1   g26209(.A1(new_n26276_), .A2(new_n26271_), .B(new_n26255_), .ZN(new_n26277_));
  AOI21_X1   g26210(.A1(new_n26275_), .A2(new_n26277_), .B(new_n26113_), .ZN(new_n26278_));
  AOI21_X1   g26211(.A1(new_n26269_), .A2(new_n26278_), .B(new_n26274_), .ZN(new_n26279_));
  NAND2_X1   g26212(.A1(new_n26248_), .A2(new_n26246_), .ZN(new_n26280_));
  NOR2_X1    g26213(.A1(new_n26248_), .A2(new_n26246_), .ZN(new_n26281_));
  AOI21_X1   g26214(.A1(new_n26238_), .A2(new_n26280_), .B(new_n26281_), .ZN(new_n26282_));
  OAI22_X1   g26215(.A1(new_n19437_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n17784_), .ZN(new_n26283_));
  NAND2_X1   g26216(.A1(new_n19472_), .A2(new_n3312_), .ZN(new_n26284_));
  AOI21_X1   g26217(.A1(new_n26284_), .A2(new_n26283_), .B(new_n3302_), .ZN(new_n26285_));
  NAND2_X1   g26218(.A1(new_n21117_), .A2(new_n26285_), .ZN(new_n26286_));
  XOR2_X1    g26219(.A1(new_n26286_), .A2(\a[23] ), .Z(new_n26287_));
  INV_X1     g26220(.I(new_n26287_), .ZN(new_n26288_));
  OAI22_X1   g26221(.A1(new_n19423_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n17787_), .ZN(new_n26289_));
  NAND2_X1   g26222(.A1(new_n20896_), .A2(new_n3317_), .ZN(new_n26290_));
  AOI21_X1   g26223(.A1(new_n26290_), .A2(new_n26289_), .B(new_n3260_), .ZN(new_n26291_));
  NAND2_X1   g26224(.A1(new_n22226_), .A2(new_n26291_), .ZN(new_n26292_));
  XOR2_X1    g26225(.A1(new_n26292_), .A2(\a[26] ), .Z(new_n26293_));
  INV_X1     g26226(.I(new_n26293_), .ZN(new_n26294_));
  OAI22_X1   g26227(.A1(new_n19410_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n17789_), .ZN(new_n26295_));
  NAND2_X1   g26228(.A1(new_n19415_), .A2(new_n2750_), .ZN(new_n26296_));
  AOI21_X1   g26229(.A1(new_n26296_), .A2(new_n26295_), .B(new_n2737_), .ZN(new_n26297_));
  NAND2_X1   g26230(.A1(new_n20846_), .A2(new_n26297_), .ZN(new_n26298_));
  XOR2_X1    g26231(.A1(new_n26298_), .A2(new_n74_), .Z(new_n26299_));
  NAND2_X1   g26232(.A1(new_n19399_), .A2(new_n3332_), .ZN(new_n26300_));
  NAND2_X1   g26233(.A1(new_n19394_), .A2(new_n3189_), .ZN(new_n26301_));
  AOI21_X1   g26234(.A1(new_n17794_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n26302_));
  NAND4_X1   g26235(.A1(new_n20264_), .A2(new_n26300_), .A3(new_n26301_), .A4(new_n26302_), .ZN(new_n26303_));
  NOR4_X1    g26236(.A1(new_n25957_), .A2(new_n25953_), .A3(new_n25973_), .A4(new_n26154_), .ZN(new_n26304_));
  AND3_X2    g26237(.A1(new_n25957_), .A2(new_n25953_), .A3(new_n26154_), .Z(new_n26305_));
  NOR2_X1    g26238(.A1(new_n26305_), .A2(new_n26304_), .ZN(new_n26306_));
  NOR2_X1    g26239(.A1(new_n24835_), .A2(new_n12019_), .ZN(new_n26307_));
  AOI21_X1   g26240(.A1(new_n24826_), .A2(new_n12021_), .B(\a[8] ), .ZN(new_n26308_));
  NOR2_X1    g26241(.A1(new_n26307_), .A2(new_n26308_), .ZN(new_n26309_));
  NOR2_X1    g26242(.A1(new_n2429_), .A2(new_n552_), .ZN(new_n26310_));
  NOR4_X1    g26243(.A1(new_n26310_), .A2(new_n1384_), .A3(new_n4022_), .A4(new_n11523_), .ZN(new_n26311_));
  NOR4_X1    g26244(.A1(new_n525_), .A2(new_n465_), .A3(new_n946_), .A4(new_n1865_), .ZN(new_n26312_));
  AND3_X2    g26245(.A1(new_n26312_), .A2(new_n859_), .A3(new_n2540_), .Z(new_n26313_));
  NAND4_X1   g26246(.A1(new_n26313_), .A2(new_n26311_), .A3(new_n2170_), .A4(new_n11513_), .ZN(new_n26314_));
  NOR3_X1    g26247(.A1(new_n760_), .A2(new_n4744_), .A3(new_n26314_), .ZN(new_n26315_));
  NOR2_X1    g26248(.A1(new_n25973_), .A2(new_n26315_), .ZN(new_n26316_));
  INV_X1     g26249(.I(new_n26315_), .ZN(new_n26317_));
  NOR2_X1    g26250(.A1(new_n25972_), .A2(new_n26317_), .ZN(new_n26318_));
  NOR2_X1    g26251(.A1(new_n26316_), .A2(new_n26318_), .ZN(new_n26319_));
  NOR2_X1    g26252(.A1(new_n26309_), .A2(new_n26319_), .ZN(new_n26320_));
  XOR2_X1    g26253(.A1(new_n25972_), .A2(new_n26315_), .Z(new_n26321_));
  INV_X1     g26254(.I(new_n26321_), .ZN(new_n26322_));
  AOI21_X1   g26255(.A1(new_n26309_), .A2(new_n26322_), .B(new_n26320_), .ZN(new_n26323_));
  NOR2_X1    g26256(.A1(new_n26306_), .A2(new_n26323_), .ZN(new_n26324_));
  INV_X1     g26257(.I(new_n26324_), .ZN(new_n26325_));
  NAND2_X1   g26258(.A1(new_n26306_), .A2(new_n26323_), .ZN(new_n26326_));
  NAND2_X1   g26259(.A1(new_n26325_), .A2(new_n26326_), .ZN(new_n26327_));
  XOR2_X1    g26260(.A1(new_n26327_), .A2(new_n26303_), .Z(new_n26328_));
  XOR2_X1    g26261(.A1(new_n26328_), .A2(new_n26299_), .Z(new_n26329_));
  INV_X1     g26262(.I(new_n26158_), .ZN(new_n26330_));
  NAND2_X1   g26263(.A1(new_n26330_), .A2(new_n26162_), .ZN(new_n26331_));
  OAI21_X1   g26264(.A1(new_n26137_), .A2(new_n26163_), .B(new_n26331_), .ZN(new_n26332_));
  XOR2_X1    g26265(.A1(new_n26329_), .A2(new_n26332_), .Z(new_n26333_));
  NOR2_X1    g26266(.A1(new_n26129_), .A2(new_n26135_), .ZN(new_n26334_));
  AND3_X2    g26267(.A1(new_n26164_), .A2(new_n26129_), .A3(new_n26135_), .Z(new_n26335_));
  NOR2_X1    g26268(.A1(new_n26335_), .A2(new_n26334_), .ZN(new_n26336_));
  XOR2_X1    g26269(.A1(new_n26336_), .A2(new_n26333_), .Z(new_n26337_));
  XOR2_X1    g26270(.A1(new_n26337_), .A2(new_n26294_), .Z(new_n26338_));
  XOR2_X1    g26271(.A1(new_n26338_), .A2(new_n26288_), .Z(new_n26339_));
  NOR2_X1    g26272(.A1(new_n26166_), .A2(new_n26170_), .ZN(new_n26340_));
  NAND2_X1   g26273(.A1(new_n26339_), .A2(new_n26340_), .ZN(new_n26341_));
  XOR2_X1    g26274(.A1(new_n26338_), .A2(new_n26287_), .Z(new_n26342_));
  INV_X1     g26275(.I(new_n26340_), .ZN(new_n26343_));
  NAND2_X1   g26276(.A1(new_n26342_), .A2(new_n26343_), .ZN(new_n26344_));
  NOR2_X1    g26277(.A1(new_n26180_), .A2(new_n26123_), .ZN(new_n26345_));
  NAND3_X1   g26278(.A1(new_n26341_), .A2(new_n26344_), .A3(new_n26345_), .ZN(new_n26346_));
  NOR2_X1    g26279(.A1(new_n26342_), .A2(new_n26343_), .ZN(new_n26347_));
  NOR2_X1    g26280(.A1(new_n26339_), .A2(new_n26340_), .ZN(new_n26348_));
  INV_X1     g26281(.I(new_n26345_), .ZN(new_n26349_));
  OAI21_X1   g26282(.A1(new_n26347_), .A2(new_n26348_), .B(new_n26349_), .ZN(new_n26350_));
  NAND2_X1   g26283(.A1(new_n26350_), .A2(new_n26346_), .ZN(new_n26351_));
  NOR2_X1    g26284(.A1(new_n26176_), .A2(new_n26118_), .ZN(new_n26352_));
  NAND2_X1   g26285(.A1(new_n26180_), .A2(new_n26124_), .ZN(new_n26353_));
  NAND2_X1   g26286(.A1(new_n26171_), .A2(new_n26123_), .ZN(new_n26354_));
  AOI22_X1   g26287(.A1(new_n26353_), .A2(new_n26354_), .B1(new_n26118_), .B2(new_n26176_), .ZN(new_n26355_));
  NOR2_X1    g26288(.A1(new_n26355_), .A2(new_n26352_), .ZN(new_n26356_));
  OAI22_X1   g26289(.A1(new_n17775_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19475_), .ZN(new_n26357_));
  NAND2_X1   g26290(.A1(new_n21157_), .A2(new_n4096_), .ZN(new_n26358_));
  AOI21_X1   g26291(.A1(new_n26358_), .A2(new_n26357_), .B(new_n4095_), .ZN(new_n26359_));
  NAND2_X1   g26292(.A1(new_n21155_), .A2(new_n26359_), .ZN(new_n26360_));
  XOR2_X1    g26293(.A1(new_n26360_), .A2(\a[20] ), .Z(new_n26361_));
  NAND2_X1   g26294(.A1(new_n26356_), .A2(new_n26361_), .ZN(new_n26362_));
  NOR2_X1    g26295(.A1(new_n26356_), .A2(new_n26361_), .ZN(new_n26363_));
  INV_X1     g26296(.I(new_n26363_), .ZN(new_n26364_));
  NAND2_X1   g26297(.A1(new_n26364_), .A2(new_n26362_), .ZN(new_n26365_));
  NAND2_X1   g26298(.A1(new_n26365_), .A2(new_n26351_), .ZN(new_n26366_));
  NOR3_X1    g26299(.A1(new_n26347_), .A2(new_n26348_), .A3(new_n26349_), .ZN(new_n26367_));
  AOI21_X1   g26300(.A1(new_n26341_), .A2(new_n26344_), .B(new_n26345_), .ZN(new_n26368_));
  NOR2_X1    g26301(.A1(new_n26368_), .A2(new_n26367_), .ZN(new_n26369_));
  OAI21_X1   g26302(.A1(new_n26355_), .A2(new_n26352_), .B(new_n26361_), .ZN(new_n26370_));
  INV_X1     g26303(.I(new_n26361_), .ZN(new_n26371_));
  NAND2_X1   g26304(.A1(new_n26356_), .A2(new_n26371_), .ZN(new_n26372_));
  NAND2_X1   g26305(.A1(new_n26372_), .A2(new_n26370_), .ZN(new_n26373_));
  NAND2_X1   g26306(.A1(new_n26369_), .A2(new_n26373_), .ZN(new_n26374_));
  NAND2_X1   g26307(.A1(new_n26366_), .A2(new_n26374_), .ZN(new_n26375_));
  INV_X1     g26308(.I(new_n26375_), .ZN(new_n26376_));
  OAI22_X1   g26309(.A1(new_n22115_), .A2(new_n6089_), .B1(new_n6094_), .B2(new_n22149_), .ZN(new_n26377_));
  NAND2_X1   g26310(.A1(new_n23957_), .A2(new_n6090_), .ZN(new_n26378_));
  AOI21_X1   g26311(.A1(new_n26377_), .A2(new_n26378_), .B(new_n6082_), .ZN(new_n26379_));
  NAND2_X1   g26312(.A1(new_n23955_), .A2(new_n26379_), .ZN(new_n26380_));
  XOR2_X1    g26313(.A1(new_n26380_), .A2(\a[14] ), .Z(new_n26381_));
  INV_X1     g26314(.I(new_n26381_), .ZN(new_n26382_));
  NAND2_X1   g26315(.A1(new_n26200_), .A2(new_n26197_), .ZN(new_n26383_));
  OAI22_X1   g26316(.A1(new_n19512_), .A2(new_n4291_), .B1(new_n21960_), .B2(new_n4297_), .ZN(new_n26384_));
  NAND2_X1   g26317(.A1(new_n22048_), .A2(new_n4469_), .ZN(new_n26385_));
  AOI21_X1   g26318(.A1(new_n26385_), .A2(new_n26384_), .B(new_n4468_), .ZN(new_n26386_));
  NAND2_X1   g26319(.A1(new_n22175_), .A2(new_n26386_), .ZN(new_n26387_));
  XOR2_X1    g26320(.A1(new_n26387_), .A2(\a[17] ), .Z(new_n26388_));
  NAND3_X1   g26321(.A1(new_n26383_), .A2(new_n26198_), .A3(new_n26388_), .ZN(new_n26389_));
  INV_X1     g26322(.I(new_n26389_), .ZN(new_n26390_));
  AOI21_X1   g26323(.A1(new_n26383_), .A2(new_n26198_), .B(new_n26388_), .ZN(new_n26391_));
  NOR2_X1    g26324(.A1(new_n26390_), .A2(new_n26391_), .ZN(new_n26392_));
  OAI21_X1   g26325(.A1(new_n26216_), .A2(new_n26212_), .B(new_n26213_), .ZN(new_n26393_));
  NAND2_X1   g26326(.A1(new_n26392_), .A2(new_n26393_), .ZN(new_n26394_));
  INV_X1     g26327(.I(new_n26391_), .ZN(new_n26395_));
  NAND2_X1   g26328(.A1(new_n26395_), .A2(new_n26389_), .ZN(new_n26396_));
  INV_X1     g26329(.I(new_n26393_), .ZN(new_n26397_));
  NAND2_X1   g26330(.A1(new_n26397_), .A2(new_n26396_), .ZN(new_n26398_));
  AOI21_X1   g26331(.A1(new_n26398_), .A2(new_n26394_), .B(new_n26382_), .ZN(new_n26399_));
  NOR2_X1    g26332(.A1(new_n26397_), .A2(new_n26396_), .ZN(new_n26400_));
  NOR2_X1    g26333(.A1(new_n26392_), .A2(new_n26393_), .ZN(new_n26401_));
  NOR3_X1    g26334(.A1(new_n26400_), .A2(new_n26401_), .A3(new_n26381_), .ZN(new_n26402_));
  OAI21_X1   g26335(.A1(new_n26402_), .A2(new_n26399_), .B(new_n26376_), .ZN(new_n26403_));
  OAI21_X1   g26336(.A1(new_n26400_), .A2(new_n26401_), .B(new_n26381_), .ZN(new_n26404_));
  NAND3_X1   g26337(.A1(new_n26398_), .A2(new_n26394_), .A3(new_n26382_), .ZN(new_n26405_));
  NAND3_X1   g26338(.A1(new_n26404_), .A2(new_n26405_), .A3(new_n26375_), .ZN(new_n26406_));
  NAND2_X1   g26339(.A1(new_n26403_), .A2(new_n26406_), .ZN(new_n26407_));
  INV_X1     g26340(.I(new_n26407_), .ZN(new_n26408_));
  INV_X1     g26341(.I(new_n26227_), .ZN(new_n26409_));
  OAI22_X1   g26342(.A1(new_n24376_), .A2(new_n4719_), .B1(new_n4716_), .B2(new_n24167_), .ZN(new_n26410_));
  NAND2_X1   g26343(.A1(new_n24620_), .A2(new_n4709_), .ZN(new_n26411_));
  AOI21_X1   g26344(.A1(new_n26411_), .A2(new_n26410_), .B(new_n4707_), .ZN(new_n26412_));
  NAND2_X1   g26345(.A1(new_n24618_), .A2(new_n26412_), .ZN(new_n26413_));
  XOR2_X1    g26346(.A1(new_n26413_), .A2(\a[11] ), .Z(new_n26414_));
  NAND3_X1   g26347(.A1(new_n26219_), .A2(new_n26409_), .A3(new_n26414_), .ZN(new_n26415_));
  INV_X1     g26348(.I(new_n26415_), .ZN(new_n26416_));
  AOI21_X1   g26349(.A1(new_n26219_), .A2(new_n26409_), .B(new_n26414_), .ZN(new_n26417_));
  NAND3_X1   g26350(.A1(new_n26409_), .A2(new_n26218_), .A3(new_n26215_), .ZN(new_n26418_));
  NAND2_X1   g26351(.A1(new_n26219_), .A2(new_n26227_), .ZN(new_n26419_));
  AOI21_X1   g26352(.A1(new_n26419_), .A2(new_n26418_), .B(new_n26234_), .ZN(new_n26420_));
  INV_X1     g26353(.I(new_n26420_), .ZN(new_n26421_));
  NOR3_X1    g26354(.A1(new_n26421_), .A2(new_n26416_), .A3(new_n26417_), .ZN(new_n26422_));
  NOR2_X1    g26355(.A1(new_n26416_), .A2(new_n26417_), .ZN(new_n26423_));
  NOR2_X1    g26356(.A1(new_n26423_), .A2(new_n26420_), .ZN(new_n26424_));
  NOR2_X1    g26357(.A1(new_n26422_), .A2(new_n26424_), .ZN(new_n26425_));
  NAND2_X1   g26358(.A1(new_n26408_), .A2(new_n26425_), .ZN(new_n26426_));
  INV_X1     g26359(.I(new_n26426_), .ZN(new_n26427_));
  OAI21_X1   g26360(.A1(new_n26422_), .A2(new_n26424_), .B(new_n26407_), .ZN(new_n26428_));
  INV_X1     g26361(.I(new_n26428_), .ZN(new_n26429_));
  NOR2_X1    g26362(.A1(new_n26427_), .A2(new_n26429_), .ZN(new_n26430_));
  XOR2_X1    g26363(.A1(new_n26430_), .A2(new_n26282_), .Z(new_n26431_));
  NOR4_X1    g26364(.A1(new_n25894_), .A2(new_n25898_), .A3(new_n26101_), .A4(new_n26263_), .ZN(new_n26432_));
  XOR2_X1    g26365(.A1(new_n26432_), .A2(new_n26431_), .Z(new_n26433_));
  XOR2_X1    g26366(.A1(new_n26433_), .A2(new_n26279_), .Z(\result[13] ));
  INV_X1     g26367(.I(new_n26274_), .ZN(new_n26435_));
  INV_X1     g26368(.I(new_n26113_), .ZN(new_n26436_));
  NOR3_X1    g26369(.A1(new_n26276_), .A2(new_n26255_), .A3(new_n26271_), .ZN(new_n26437_));
  AOI21_X1   g26370(.A1(new_n26272_), .A2(new_n26273_), .B(new_n26270_), .ZN(new_n26438_));
  OAI21_X1   g26371(.A1(new_n26438_), .A2(new_n26437_), .B(new_n26436_), .ZN(new_n26439_));
  OAI21_X1   g26372(.A1(new_n26108_), .A2(new_n26439_), .B(new_n26435_), .ZN(new_n26440_));
  XOR2_X1    g26373(.A1(new_n26431_), .A2(new_n26440_), .Z(new_n26441_));
  NAND4_X1   g26374(.A1(new_n25899_), .A2(new_n26102_), .A3(new_n26262_), .A4(new_n26441_), .ZN(new_n26442_));
  NOR3_X1    g26375(.A1(new_n26307_), .A2(new_n26308_), .A3(new_n26316_), .ZN(new_n26443_));
  NOR2_X1    g26376(.A1(new_n26443_), .A2(new_n26318_), .ZN(new_n26444_));
  INV_X1     g26377(.I(new_n26444_), .ZN(new_n26445_));
  NAND2_X1   g26378(.A1(new_n17790_), .A2(new_n3332_), .ZN(new_n26446_));
  NAND2_X1   g26379(.A1(new_n19399_), .A2(new_n3189_), .ZN(new_n26447_));
  AOI21_X1   g26380(.A1(new_n19394_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n26448_));
  NAND4_X1   g26381(.A1(new_n22673_), .A2(new_n26446_), .A3(new_n26447_), .A4(new_n26448_), .ZN(new_n26449_));
  INV_X1     g26382(.I(new_n12981_), .ZN(new_n26450_));
  NOR4_X1    g26383(.A1(new_n782_), .A2(new_n213_), .A3(new_n1236_), .A4(new_n640_), .ZN(new_n26451_));
  NOR4_X1    g26384(.A1(new_n229_), .A2(new_n26450_), .A3(new_n3419_), .A4(new_n26451_), .ZN(new_n26452_));
  NAND3_X1   g26385(.A1(new_n3676_), .A2(new_n1658_), .A3(new_n378_), .ZN(new_n26453_));
  NOR4_X1    g26386(.A1(new_n3670_), .A2(new_n558_), .A3(new_n3685_), .A4(new_n26453_), .ZN(new_n26454_));
  AND4_X2    g26387(.A1(new_n478_), .A2(new_n12265_), .A3(new_n26452_), .A4(new_n26454_), .Z(new_n26455_));
  NAND2_X1   g26388(.A1(new_n2281_), .A2(new_n26455_), .ZN(new_n26456_));
  INV_X1     g26389(.I(new_n26456_), .ZN(new_n26457_));
  XOR2_X1    g26390(.A1(new_n26449_), .A2(new_n26457_), .Z(new_n26458_));
  INV_X1     g26391(.I(new_n26458_), .ZN(new_n26459_));
  XOR2_X1    g26392(.A1(new_n26449_), .A2(new_n26456_), .Z(new_n26460_));
  NOR2_X1    g26393(.A1(new_n26460_), .A2(new_n26445_), .ZN(new_n26461_));
  AOI21_X1   g26394(.A1(new_n26445_), .A2(new_n26459_), .B(new_n26461_), .ZN(new_n26462_));
  OAI22_X1   g26395(.A1(new_n19410_), .A2(new_n2747_), .B1(new_n19412_), .B2(new_n2742_), .ZN(new_n26463_));
  NAND2_X1   g26396(.A1(new_n19439_), .A2(new_n2750_), .ZN(new_n26464_));
  AOI21_X1   g26397(.A1(new_n26464_), .A2(new_n26463_), .B(new_n2737_), .ZN(new_n26465_));
  NAND2_X1   g26398(.A1(new_n20827_), .A2(new_n26465_), .ZN(new_n26466_));
  XOR2_X1    g26399(.A1(new_n26466_), .A2(new_n74_), .Z(new_n26467_));
  XOR2_X1    g26400(.A1(new_n26306_), .A2(new_n26323_), .Z(new_n26468_));
  AOI21_X1   g26401(.A1(new_n26468_), .A2(new_n26303_), .B(new_n26324_), .ZN(new_n26469_));
  INV_X1     g26402(.I(new_n26469_), .ZN(new_n26470_));
  XOR2_X1    g26403(.A1(new_n26467_), .A2(new_n26470_), .Z(new_n26471_));
  XOR2_X1    g26404(.A1(new_n26471_), .A2(new_n26462_), .Z(new_n26472_));
  OAI22_X1   g26405(.A1(new_n19428_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19423_), .ZN(new_n26473_));
  NAND2_X1   g26406(.A1(new_n19438_), .A2(new_n3317_), .ZN(new_n26474_));
  AOI21_X1   g26407(.A1(new_n26474_), .A2(new_n26473_), .B(new_n3260_), .ZN(new_n26475_));
  NAND2_X1   g26408(.A1(new_n20907_), .A2(new_n26475_), .ZN(new_n26476_));
  XOR2_X1    g26409(.A1(new_n26476_), .A2(\a[26] ), .Z(new_n26477_));
  XOR2_X1    g26410(.A1(new_n26303_), .A2(new_n26323_), .Z(new_n26478_));
  XNOR2_X1   g26411(.A1(new_n26478_), .A2(new_n26306_), .ZN(new_n26479_));
  OR2_X2     g26412(.A1(new_n26299_), .A2(new_n26479_), .Z(new_n26480_));
  NAND3_X1   g26413(.A1(new_n26329_), .A2(new_n26332_), .A3(new_n26480_), .ZN(new_n26481_));
  XOR2_X1    g26414(.A1(new_n26477_), .A2(new_n26481_), .Z(new_n26482_));
  XOR2_X1    g26415(.A1(new_n26482_), .A2(new_n26472_), .Z(new_n26483_));
  NOR2_X1    g26416(.A1(new_n26336_), .A2(new_n26293_), .ZN(new_n26484_));
  AOI21_X1   g26417(.A1(new_n26336_), .A2(new_n26293_), .B(new_n26333_), .ZN(new_n26485_));
  NOR2_X1    g26418(.A1(new_n26485_), .A2(new_n26484_), .ZN(new_n26486_));
  OAI22_X1   g26419(.A1(new_n19463_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19437_), .ZN(new_n26487_));
  NAND2_X1   g26420(.A1(new_n17780_), .A2(new_n3312_), .ZN(new_n26488_));
  AOI21_X1   g26421(.A1(new_n26487_), .A2(new_n26488_), .B(new_n3302_), .ZN(new_n26489_));
  NAND2_X1   g26422(.A1(new_n21088_), .A2(new_n26489_), .ZN(new_n26490_));
  XOR2_X1    g26423(.A1(new_n26490_), .A2(\a[23] ), .Z(new_n26491_));
  NAND2_X1   g26424(.A1(new_n26486_), .A2(new_n26491_), .ZN(new_n26492_));
  OR2_X2     g26425(.A1(new_n26486_), .A2(new_n26491_), .Z(new_n26493_));
  NAND2_X1   g26426(.A1(new_n26493_), .A2(new_n26492_), .ZN(new_n26494_));
  XOR2_X1    g26427(.A1(new_n26486_), .A2(new_n26491_), .Z(new_n26495_));
  MUX2_X1    g26428(.I0(new_n26495_), .I1(new_n26494_), .S(new_n26483_), .Z(new_n26496_));
  OAI22_X1   g26429(.A1(new_n19522_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n17775_), .ZN(new_n26497_));
  NAND2_X1   g26430(.A1(new_n17770_), .A2(new_n4096_), .ZN(new_n26498_));
  AOI21_X1   g26431(.A1(new_n26498_), .A2(new_n26497_), .B(new_n4095_), .ZN(new_n26499_));
  NAND2_X1   g26432(.A1(new_n19521_), .A2(new_n26499_), .ZN(new_n26500_));
  XOR2_X1    g26433(.A1(new_n26500_), .A2(\a[20] ), .Z(new_n26501_));
  INV_X1     g26434(.I(new_n26501_), .ZN(new_n26502_));
  NOR2_X1    g26435(.A1(new_n26170_), .A2(new_n26123_), .ZN(new_n26503_));
  AOI21_X1   g26436(.A1(new_n26123_), .A2(new_n26170_), .B(new_n26166_), .ZN(new_n26504_));
  XOR2_X1    g26437(.A1(new_n26336_), .A2(new_n26294_), .Z(new_n26505_));
  XOR2_X1    g26438(.A1(new_n26505_), .A2(new_n26333_), .Z(new_n26506_));
  NOR2_X1    g26439(.A1(new_n26506_), .A2(new_n26288_), .ZN(new_n26507_));
  NOR4_X1    g26440(.A1(new_n26342_), .A2(new_n26503_), .A3(new_n26504_), .A4(new_n26507_), .ZN(new_n26508_));
  XOR2_X1    g26441(.A1(new_n26508_), .A2(new_n26502_), .Z(new_n26509_));
  XOR2_X1    g26442(.A1(new_n26509_), .A2(new_n26496_), .Z(new_n26510_));
  AOI21_X1   g26443(.A1(new_n26369_), .A2(new_n26362_), .B(new_n26363_), .ZN(new_n26511_));
  AOI22_X1   g26444(.A1(new_n22048_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n21953_), .ZN(new_n26512_));
  NOR2_X1    g26445(.A1(new_n22115_), .A2(new_n4470_), .ZN(new_n26513_));
  OAI21_X1   g26446(.A1(new_n26513_), .A2(new_n26512_), .B(new_n4295_), .ZN(new_n26514_));
  NOR2_X1    g26447(.A1(new_n23675_), .A2(new_n26514_), .ZN(new_n26515_));
  XOR2_X1    g26448(.A1(new_n26515_), .A2(new_n3372_), .Z(new_n26516_));
  NAND2_X1   g26449(.A1(new_n26511_), .A2(new_n26516_), .ZN(new_n26517_));
  NOR2_X1    g26450(.A1(new_n26511_), .A2(new_n26516_), .ZN(new_n26518_));
  INV_X1     g26451(.I(new_n26518_), .ZN(new_n26519_));
  AOI21_X1   g26452(.A1(new_n26519_), .A2(new_n26517_), .B(new_n26510_), .ZN(new_n26520_));
  XOR2_X1    g26453(.A1(new_n26511_), .A2(new_n26516_), .Z(new_n26521_));
  AOI21_X1   g26454(.A1(new_n26521_), .A2(new_n26510_), .B(new_n26520_), .ZN(new_n26522_));
  OAI21_X1   g26455(.A1(new_n26375_), .A2(new_n26390_), .B(new_n26395_), .ZN(new_n26523_));
  OAI22_X1   g26456(.A1(new_n23948_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n22149_), .ZN(new_n26524_));
  NAND2_X1   g26457(.A1(new_n24174_), .A2(new_n6090_), .ZN(new_n26525_));
  AOI21_X1   g26458(.A1(new_n26525_), .A2(new_n26524_), .B(new_n6082_), .ZN(new_n26526_));
  NAND2_X1   g26459(.A1(new_n24172_), .A2(new_n26526_), .ZN(new_n26527_));
  XOR2_X1    g26460(.A1(new_n26527_), .A2(\a[14] ), .Z(new_n26528_));
  INV_X1     g26461(.I(new_n26528_), .ZN(new_n26529_));
  NOR2_X1    g26462(.A1(new_n26523_), .A2(new_n26529_), .ZN(new_n26530_));
  INV_X1     g26463(.I(new_n26530_), .ZN(new_n26531_));
  NAND2_X1   g26464(.A1(new_n26523_), .A2(new_n26529_), .ZN(new_n26532_));
  AOI21_X1   g26465(.A1(new_n26531_), .A2(new_n26532_), .B(new_n26522_), .ZN(new_n26533_));
  XNOR2_X1   g26466(.A1(new_n26509_), .A2(new_n26496_), .ZN(new_n26534_));
  INV_X1     g26467(.I(new_n26517_), .ZN(new_n26535_));
  OAI21_X1   g26468(.A1(new_n26535_), .A2(new_n26518_), .B(new_n26534_), .ZN(new_n26536_));
  INV_X1     g26469(.I(new_n26516_), .ZN(new_n26537_));
  NOR2_X1    g26470(.A1(new_n26511_), .A2(new_n26537_), .ZN(new_n26538_));
  AND2_X2    g26471(.A1(new_n26511_), .A2(new_n26537_), .Z(new_n26539_));
  OAI21_X1   g26472(.A1(new_n26539_), .A2(new_n26538_), .B(new_n26510_), .ZN(new_n26540_));
  NAND2_X1   g26473(.A1(new_n26536_), .A2(new_n26540_), .ZN(new_n26541_));
  NAND2_X1   g26474(.A1(new_n26523_), .A2(new_n26528_), .ZN(new_n26542_));
  NOR2_X1    g26475(.A1(new_n26523_), .A2(new_n26528_), .ZN(new_n26543_));
  INV_X1     g26476(.I(new_n26543_), .ZN(new_n26544_));
  AOI21_X1   g26477(.A1(new_n26544_), .A2(new_n26542_), .B(new_n26541_), .ZN(new_n26545_));
  NOR2_X1    g26478(.A1(new_n26533_), .A2(new_n26545_), .ZN(new_n26546_));
  NOR2_X1    g26479(.A1(new_n26397_), .A2(new_n26381_), .ZN(new_n26547_));
  INV_X1     g26480(.I(new_n26547_), .ZN(new_n26548_));
  NOR2_X1    g26481(.A1(new_n26393_), .A2(new_n26382_), .ZN(new_n26549_));
  NOR2_X1    g26482(.A1(new_n26396_), .A2(new_n26376_), .ZN(new_n26550_));
  NOR2_X1    g26483(.A1(new_n26392_), .A2(new_n26375_), .ZN(new_n26551_));
  NOR2_X1    g26484(.A1(new_n26550_), .A2(new_n26551_), .ZN(new_n26552_));
  OAI21_X1   g26485(.A1(new_n26552_), .A2(new_n26549_), .B(new_n26548_), .ZN(new_n26553_));
  INV_X1     g26486(.I(new_n24833_), .ZN(new_n26554_));
  AOI22_X1   g26487(.A1(new_n24620_), .A2(new_n4720_), .B1(new_n6480_), .B2(new_n24386_), .ZN(new_n26555_));
  NOR2_X1    g26488(.A1(new_n24835_), .A2(new_n4710_), .ZN(new_n26556_));
  OAI21_X1   g26489(.A1(new_n26556_), .A2(new_n26555_), .B(new_n4706_), .ZN(new_n26557_));
  NOR2_X1    g26490(.A1(new_n26554_), .A2(new_n26557_), .ZN(new_n26558_));
  XOR2_X1    g26491(.A1(new_n26558_), .A2(new_n4034_), .Z(new_n26559_));
  INV_X1     g26492(.I(new_n26559_), .ZN(new_n26560_));
  NOR2_X1    g26493(.A1(new_n26553_), .A2(new_n26560_), .ZN(new_n26561_));
  INV_X1     g26494(.I(new_n26561_), .ZN(new_n26562_));
  NAND2_X1   g26495(.A1(new_n26553_), .A2(new_n26560_), .ZN(new_n26563_));
  AOI21_X1   g26496(.A1(new_n26562_), .A2(new_n26563_), .B(new_n26546_), .ZN(new_n26564_));
  INV_X1     g26497(.I(new_n26532_), .ZN(new_n26565_));
  OAI21_X1   g26498(.A1(new_n26565_), .A2(new_n26530_), .B(new_n26541_), .ZN(new_n26566_));
  INV_X1     g26499(.I(new_n26542_), .ZN(new_n26567_));
  OAI21_X1   g26500(.A1(new_n26567_), .A2(new_n26543_), .B(new_n26522_), .ZN(new_n26568_));
  NAND2_X1   g26501(.A1(new_n26568_), .A2(new_n26566_), .ZN(new_n26569_));
  NAND2_X1   g26502(.A1(new_n26553_), .A2(new_n26559_), .ZN(new_n26570_));
  NOR2_X1    g26503(.A1(new_n26553_), .A2(new_n26559_), .ZN(new_n26571_));
  INV_X1     g26504(.I(new_n26571_), .ZN(new_n26572_));
  AOI21_X1   g26505(.A1(new_n26572_), .A2(new_n26570_), .B(new_n26569_), .ZN(new_n26573_));
  NOR2_X1    g26506(.A1(new_n26227_), .A2(new_n26234_), .ZN(new_n26574_));
  AOI22_X1   g26507(.A1(new_n26218_), .A2(new_n26215_), .B1(new_n26227_), .B2(new_n26234_), .ZN(new_n26575_));
  NOR2_X1    g26508(.A1(new_n26575_), .A2(new_n26574_), .ZN(new_n26576_));
  OR2_X2     g26509(.A1(new_n26576_), .A2(new_n26414_), .Z(new_n26577_));
  NAND2_X1   g26510(.A1(new_n26576_), .A2(new_n26414_), .ZN(new_n26578_));
  NAND3_X1   g26511(.A1(new_n26403_), .A2(new_n26406_), .A3(new_n26578_), .ZN(new_n26579_));
  NAND2_X1   g26512(.A1(new_n26579_), .A2(new_n26577_), .ZN(new_n26580_));
  NOR3_X1    g26513(.A1(new_n26564_), .A2(new_n26573_), .A3(new_n26580_), .ZN(new_n26581_));
  INV_X1     g26514(.I(new_n26549_), .ZN(new_n26582_));
  XOR2_X1    g26515(.A1(new_n26392_), .A2(new_n26376_), .Z(new_n26583_));
  AOI21_X1   g26516(.A1(new_n26583_), .A2(new_n26582_), .B(new_n26547_), .ZN(new_n26584_));
  NOR2_X1    g26517(.A1(new_n26584_), .A2(new_n26559_), .ZN(new_n26585_));
  OAI22_X1   g26518(.A1(new_n26585_), .A2(new_n26561_), .B1(new_n26533_), .B2(new_n26545_), .ZN(new_n26586_));
  INV_X1     g26519(.I(new_n26570_), .ZN(new_n26587_));
  OAI21_X1   g26520(.A1(new_n26587_), .A2(new_n26571_), .B(new_n26546_), .ZN(new_n26588_));
  AOI22_X1   g26521(.A1(new_n26588_), .A2(new_n26586_), .B1(new_n26577_), .B2(new_n26579_), .ZN(new_n26589_));
  NOR2_X1    g26522(.A1(new_n26589_), .A2(new_n26581_), .ZN(new_n26590_));
  INV_X1     g26523(.I(new_n26282_), .ZN(new_n26591_));
  OAI21_X1   g26524(.A1(new_n26440_), .A2(new_n26430_), .B(new_n26591_), .ZN(new_n26592_));
  XNOR2_X1   g26525(.A1(new_n26592_), .A2(new_n26590_), .ZN(new_n26593_));
  XOR2_X1    g26526(.A1(new_n26442_), .A2(new_n26593_), .Z(\result[14] ));
  XOR2_X1    g26527(.A1(new_n26462_), .A2(new_n26467_), .Z(new_n26595_));
  AOI21_X1   g26528(.A1(new_n26467_), .A2(new_n26470_), .B(new_n26595_), .ZN(new_n26596_));
  NOR3_X1    g26529(.A1(new_n770_), .A2(new_n937_), .A3(new_n796_), .ZN(new_n26597_));
  NOR3_X1    g26530(.A1(new_n1787_), .A2(new_n788_), .A3(new_n288_), .ZN(new_n26598_));
  NAND2_X1   g26531(.A1(new_n26598_), .A2(new_n26597_), .ZN(new_n26599_));
  NOR3_X1    g26532(.A1(new_n26599_), .A2(new_n530_), .A3(new_n1987_), .ZN(new_n26600_));
  NOR4_X1    g26533(.A1(new_n1498_), .A2(new_n1045_), .A3(new_n1266_), .A4(new_n1944_), .ZN(new_n26601_));
  NOR4_X1    g26534(.A1(new_n458_), .A2(new_n879_), .A3(new_n400_), .A4(new_n1527_), .ZN(new_n26602_));
  NOR2_X1    g26535(.A1(new_n11522_), .A2(new_n11806_), .ZN(new_n26603_));
  NAND4_X1   g26536(.A1(new_n26603_), .A2(new_n26600_), .A3(new_n26601_), .A4(new_n26602_), .ZN(new_n26604_));
  NOR3_X1    g26537(.A1(new_n26604_), .A2(new_n25964_), .A3(new_n3974_), .ZN(new_n26605_));
  INV_X1     g26538(.I(new_n26605_), .ZN(new_n26606_));
  XOR2_X1    g26539(.A1(new_n26444_), .A2(new_n26457_), .Z(new_n26607_));
  OAI21_X1   g26540(.A1(new_n26449_), .A2(new_n26445_), .B(new_n26607_), .ZN(new_n26608_));
  AOI21_X1   g26541(.A1(new_n26445_), .A2(new_n26449_), .B(new_n26608_), .ZN(new_n26609_));
  XOR2_X1    g26542(.A1(new_n26609_), .A2(new_n26606_), .Z(new_n26610_));
  INV_X1     g26543(.I(new_n26610_), .ZN(new_n26611_));
  AOI22_X1   g26544(.A1(new_n19439_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n19415_), .ZN(new_n26612_));
  NOR2_X1    g26545(.A1(new_n19423_), .A2(new_n3175_), .ZN(new_n26613_));
  OAI21_X1   g26546(.A1(new_n26613_), .A2(new_n26612_), .B(new_n2736_), .ZN(new_n26614_));
  INV_X1     g26547(.I(new_n26614_), .ZN(new_n26615_));
  NAND2_X1   g26548(.A1(new_n20939_), .A2(new_n26615_), .ZN(new_n26616_));
  XOR2_X1    g26549(.A1(new_n26616_), .A2(\a[29] ), .Z(new_n26617_));
  NAND2_X1   g26550(.A1(new_n19407_), .A2(new_n3332_), .ZN(new_n26618_));
  NAND2_X1   g26551(.A1(new_n17790_), .A2(new_n3189_), .ZN(new_n26619_));
  AOI21_X1   g26552(.A1(new_n19399_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n26620_));
  NAND4_X1   g26553(.A1(new_n20863_), .A2(new_n26618_), .A3(new_n26619_), .A4(new_n26620_), .ZN(new_n26621_));
  XNOR2_X1   g26554(.A1(new_n26617_), .A2(new_n26621_), .ZN(new_n26622_));
  NOR2_X1    g26555(.A1(new_n26622_), .A2(new_n26611_), .ZN(new_n26623_));
  NAND2_X1   g26556(.A1(new_n26617_), .A2(new_n26621_), .ZN(new_n26624_));
  OR2_X2     g26557(.A1(new_n26617_), .A2(new_n26621_), .Z(new_n26625_));
  AOI21_X1   g26558(.A1(new_n26625_), .A2(new_n26624_), .B(new_n26610_), .ZN(new_n26626_));
  NOR2_X1    g26559(.A1(new_n26623_), .A2(new_n26626_), .ZN(new_n26627_));
  OAI22_X1   g26560(.A1(new_n17784_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19428_), .ZN(new_n26628_));
  NAND2_X1   g26561(.A1(new_n19466_), .A2(new_n3317_), .ZN(new_n26629_));
  AOI21_X1   g26562(.A1(new_n26629_), .A2(new_n26628_), .B(new_n3260_), .ZN(new_n26630_));
  NAND2_X1   g26563(.A1(new_n21100_), .A2(new_n26630_), .ZN(new_n26631_));
  XOR2_X1    g26564(.A1(new_n26631_), .A2(\a[26] ), .Z(new_n26632_));
  INV_X1     g26565(.I(new_n26632_), .ZN(new_n26633_));
  NOR2_X1    g26566(.A1(new_n26627_), .A2(new_n26633_), .ZN(new_n26634_));
  NOR3_X1    g26567(.A1(new_n26623_), .A2(new_n26626_), .A3(new_n26632_), .ZN(new_n26635_));
  OAI21_X1   g26568(.A1(new_n26634_), .A2(new_n26635_), .B(new_n26596_), .ZN(new_n26636_));
  XOR2_X1    g26569(.A1(new_n26627_), .A2(new_n26632_), .Z(new_n26637_));
  OAI21_X1   g26570(.A1(new_n26637_), .A2(new_n26596_), .B(new_n26636_), .ZN(new_n26638_));
  OAI22_X1   g26571(.A1(new_n19475_), .A2(new_n3306_), .B1(new_n19463_), .B2(new_n3310_), .ZN(new_n26639_));
  NAND2_X1   g26572(.A1(new_n19484_), .A2(new_n3312_), .ZN(new_n26640_));
  AOI21_X1   g26573(.A1(new_n26640_), .A2(new_n26639_), .B(new_n3302_), .ZN(new_n26641_));
  NAND2_X1   g26574(.A1(new_n21171_), .A2(new_n26641_), .ZN(new_n26642_));
  XOR2_X1    g26575(.A1(new_n26642_), .A2(\a[23] ), .Z(new_n26643_));
  XOR2_X1    g26576(.A1(new_n26638_), .A2(new_n26643_), .Z(new_n26644_));
  NAND2_X1   g26577(.A1(new_n26492_), .A2(new_n26483_), .ZN(new_n26645_));
  NAND2_X1   g26578(.A1(new_n26645_), .A2(new_n26493_), .ZN(new_n26646_));
  OAI22_X1   g26579(.A1(new_n19512_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n19522_), .ZN(new_n26647_));
  NAND2_X1   g26580(.A1(new_n21953_), .A2(new_n4096_), .ZN(new_n26648_));
  AOI21_X1   g26581(.A1(new_n26647_), .A2(new_n26648_), .B(new_n4095_), .ZN(new_n26649_));
  NAND2_X1   g26582(.A1(new_n21963_), .A2(new_n26649_), .ZN(new_n26650_));
  XOR2_X1    g26583(.A1(new_n26650_), .A2(new_n3035_), .Z(new_n26651_));
  NOR2_X1    g26584(.A1(new_n26651_), .A2(new_n26646_), .ZN(new_n26652_));
  INV_X1     g26585(.I(new_n26652_), .ZN(new_n26653_));
  NAND2_X1   g26586(.A1(new_n26651_), .A2(new_n26646_), .ZN(new_n26654_));
  AOI21_X1   g26587(.A1(new_n26653_), .A2(new_n26654_), .B(new_n26644_), .ZN(new_n26655_));
  XOR2_X1    g26588(.A1(new_n26651_), .A2(new_n26646_), .Z(new_n26656_));
  AOI21_X1   g26589(.A1(new_n26644_), .A2(new_n26656_), .B(new_n26655_), .ZN(new_n26657_));
  NAND2_X1   g26590(.A1(new_n26496_), .A2(new_n26501_), .ZN(new_n26658_));
  XOR2_X1    g26591(.A1(new_n26496_), .A2(new_n26502_), .Z(new_n26659_));
  NAND2_X1   g26592(.A1(new_n26659_), .A2(new_n26508_), .ZN(new_n26660_));
  NAND2_X1   g26593(.A1(new_n26660_), .A2(new_n26658_), .ZN(new_n26661_));
  OAI22_X1   g26594(.A1(new_n22115_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n22051_), .ZN(new_n26662_));
  NAND2_X1   g26595(.A1(new_n22150_), .A2(new_n4469_), .ZN(new_n26663_));
  AOI21_X1   g26596(.A1(new_n26662_), .A2(new_n26663_), .B(new_n4468_), .ZN(new_n26664_));
  NAND2_X1   g26597(.A1(new_n22163_), .A2(new_n26664_), .ZN(new_n26665_));
  XOR2_X1    g26598(.A1(new_n26665_), .A2(new_n3372_), .Z(new_n26666_));
  NOR2_X1    g26599(.A1(new_n26661_), .A2(new_n26666_), .ZN(new_n26667_));
  AND2_X2    g26600(.A1(new_n26661_), .A2(new_n26666_), .Z(new_n26668_));
  NOR2_X1    g26601(.A1(new_n26668_), .A2(new_n26667_), .ZN(new_n26669_));
  NOR2_X1    g26602(.A1(new_n26669_), .A2(new_n26657_), .ZN(new_n26670_));
  XOR2_X1    g26603(.A1(new_n26661_), .A2(new_n26666_), .Z(new_n26671_));
  AOI21_X1   g26604(.A1(new_n26657_), .A2(new_n26671_), .B(new_n26670_), .ZN(new_n26672_));
  INV_X1     g26605(.I(new_n26672_), .ZN(new_n26673_));
  AOI21_X1   g26606(.A1(new_n26534_), .A2(new_n26517_), .B(new_n26518_), .ZN(new_n26674_));
  AOI22_X1   g26607(.A1(new_n24174_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n23957_), .ZN(new_n26675_));
  NOR2_X1    g26608(.A1(new_n24376_), .A2(new_n6091_), .ZN(new_n26676_));
  NOR2_X1    g26609(.A1(new_n26676_), .A2(new_n26675_), .ZN(new_n26677_));
  OR3_X2     g26610(.A1(new_n24391_), .A2(new_n6082_), .A3(new_n26677_), .Z(new_n26678_));
  XOR2_X1    g26611(.A1(new_n26678_), .A2(\a[14] ), .Z(new_n26679_));
  NAND2_X1   g26612(.A1(new_n26674_), .A2(new_n26679_), .ZN(new_n26680_));
  OR2_X2     g26613(.A1(new_n26674_), .A2(new_n26679_), .Z(new_n26681_));
  NAND2_X1   g26614(.A1(new_n26681_), .A2(new_n26680_), .ZN(new_n26682_));
  NAND2_X1   g26615(.A1(new_n26682_), .A2(new_n26673_), .ZN(new_n26683_));
  XOR2_X1    g26616(.A1(new_n26674_), .A2(new_n26679_), .Z(new_n26684_));
  NAND2_X1   g26617(.A1(new_n26684_), .A2(new_n26672_), .ZN(new_n26685_));
  NAND2_X1   g26618(.A1(new_n26683_), .A2(new_n26685_), .ZN(new_n26686_));
  OAI21_X1   g26619(.A1(new_n26522_), .A2(new_n26530_), .B(new_n26532_), .ZN(new_n26687_));
  AOI22_X1   g26620(.A1(new_n24826_), .A2(new_n12255_), .B1(new_n6480_), .B2(new_n24620_), .ZN(new_n26688_));
  OR3_X2     g26621(.A1(new_n25017_), .A2(new_n4707_), .A3(new_n26688_), .Z(new_n26689_));
  XOR2_X1    g26622(.A1(new_n26689_), .A2(\a[11] ), .Z(new_n26690_));
  INV_X1     g26623(.I(new_n26690_), .ZN(new_n26691_));
  NOR2_X1    g26624(.A1(new_n26687_), .A2(new_n26691_), .ZN(new_n26692_));
  NAND2_X1   g26625(.A1(new_n26687_), .A2(new_n26691_), .ZN(new_n26693_));
  INV_X1     g26626(.I(new_n26693_), .ZN(new_n26694_));
  OAI21_X1   g26627(.A1(new_n26692_), .A2(new_n26694_), .B(new_n26686_), .ZN(new_n26695_));
  INV_X1     g26628(.I(new_n26686_), .ZN(new_n26696_));
  XOR2_X1    g26629(.A1(new_n26687_), .A2(new_n26691_), .Z(new_n26697_));
  NAND2_X1   g26630(.A1(new_n26696_), .A2(new_n26697_), .ZN(new_n26698_));
  NAND2_X1   g26631(.A1(new_n26698_), .A2(new_n26695_), .ZN(new_n26699_));
  AOI21_X1   g26632(.A1(new_n26562_), .A2(new_n26569_), .B(new_n26585_), .ZN(new_n26700_));
  INV_X1     g26633(.I(new_n26700_), .ZN(new_n26701_));
  AOI21_X1   g26634(.A1(new_n26426_), .A2(new_n26428_), .B(new_n26591_), .ZN(new_n26702_));
  INV_X1     g26635(.I(new_n26702_), .ZN(new_n26703_));
  NOR3_X1    g26636(.A1(new_n26589_), .A2(new_n26702_), .A3(new_n26581_), .ZN(new_n26704_));
  OAI21_X1   g26637(.A1(new_n26440_), .A2(new_n26703_), .B(new_n26704_), .ZN(new_n26705_));
  NOR2_X1    g26638(.A1(new_n26705_), .A2(new_n26581_), .ZN(new_n26706_));
  XOR2_X1    g26639(.A1(new_n26706_), .A2(new_n26701_), .Z(new_n26707_));
  XOR2_X1    g26640(.A1(new_n26707_), .A2(new_n26699_), .Z(new_n26708_));
  INV_X1     g26641(.I(new_n26708_), .ZN(new_n26709_));
  NOR2_X1    g26642(.A1(new_n26442_), .A2(new_n26593_), .ZN(new_n26710_));
  XOR2_X1    g26643(.A1(new_n26710_), .A2(new_n26709_), .Z(\result[15] ));
  NAND2_X1   g26644(.A1(new_n26699_), .A2(new_n26700_), .ZN(new_n26712_));
  INV_X1     g26645(.I(new_n26581_), .ZN(new_n26713_));
  NAND3_X1   g26646(.A1(new_n26698_), .A2(new_n26701_), .A3(new_n26695_), .ZN(new_n26714_));
  INV_X1     g26647(.I(new_n26714_), .ZN(new_n26715_));
  AOI21_X1   g26648(.A1(new_n26698_), .A2(new_n26695_), .B(new_n26701_), .ZN(new_n26716_));
  OAI21_X1   g26649(.A1(new_n26715_), .A2(new_n26716_), .B(new_n26713_), .ZN(new_n26717_));
  OAI21_X1   g26650(.A1(new_n26705_), .A2(new_n26717_), .B(new_n26712_), .ZN(new_n26718_));
  OAI21_X1   g26651(.A1(new_n26696_), .A2(new_n26692_), .B(new_n26693_), .ZN(new_n26719_));
  INV_X1     g26652(.I(new_n26719_), .ZN(new_n26720_));
  INV_X1     g26653(.I(new_n26643_), .ZN(new_n26721_));
  NAND2_X1   g26654(.A1(new_n26638_), .A2(new_n26721_), .ZN(new_n26722_));
  OAI22_X1   g26655(.A1(new_n19437_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n17784_), .ZN(new_n26723_));
  NAND2_X1   g26656(.A1(new_n19472_), .A2(new_n3317_), .ZN(new_n26724_));
  AOI21_X1   g26657(.A1(new_n26724_), .A2(new_n26723_), .B(new_n3260_), .ZN(new_n26725_));
  NAND2_X1   g26658(.A1(new_n21117_), .A2(new_n26725_), .ZN(new_n26726_));
  XOR2_X1    g26659(.A1(new_n26726_), .A2(\a[26] ), .Z(new_n26727_));
  OAI22_X1   g26660(.A1(new_n19423_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n17787_), .ZN(new_n26728_));
  NAND2_X1   g26661(.A1(new_n20896_), .A2(new_n2750_), .ZN(new_n26729_));
  AOI21_X1   g26662(.A1(new_n26729_), .A2(new_n26728_), .B(new_n2737_), .ZN(new_n26730_));
  NAND2_X1   g26663(.A1(new_n22226_), .A2(new_n26730_), .ZN(new_n26731_));
  XOR2_X1    g26664(.A1(new_n26731_), .A2(\a[29] ), .Z(new_n26732_));
  NAND2_X1   g26665(.A1(new_n26624_), .A2(new_n26610_), .ZN(new_n26733_));
  NAND2_X1   g26666(.A1(new_n26733_), .A2(new_n26625_), .ZN(new_n26734_));
  NOR4_X1    g26667(.A1(new_n26449_), .A2(new_n26444_), .A3(new_n26457_), .A4(new_n26606_), .ZN(new_n26735_));
  NOR2_X1    g26668(.A1(new_n26445_), .A2(new_n26605_), .ZN(new_n26736_));
  AOI21_X1   g26669(.A1(new_n26449_), .A2(new_n26736_), .B(new_n26735_), .ZN(new_n26737_));
  NOR2_X1    g26670(.A1(new_n24835_), .A2(new_n12256_), .ZN(new_n26738_));
  OAI22_X1   g26671(.A1(new_n26738_), .A2(\a[11] ), .B1(new_n12258_), .B2(new_n24835_), .ZN(new_n26739_));
  INV_X1     g26672(.I(new_n2520_), .ZN(new_n26740_));
  INV_X1     g26673(.I(new_n1348_), .ZN(new_n26741_));
  INV_X1     g26674(.I(new_n3837_), .ZN(new_n26742_));
  NAND4_X1   g26675(.A1(new_n874_), .A2(new_n775_), .A3(new_n1701_), .A4(new_n2192_), .ZN(new_n26743_));
  NOR4_X1    g26676(.A1(new_n573_), .A2(new_n86_), .A3(new_n782_), .A4(new_n238_), .ZN(new_n26744_));
  NOR3_X1    g26677(.A1(new_n26743_), .A2(new_n26742_), .A3(new_n26744_), .ZN(new_n26745_));
  NOR4_X1    g26678(.A1(new_n2090_), .A2(new_n1247_), .A3(new_n1996_), .A4(new_n3855_), .ZN(new_n26746_));
  NAND4_X1   g26679(.A1(new_n26746_), .A2(new_n26741_), .A3(new_n3850_), .A4(new_n26745_), .ZN(new_n26747_));
  NOR3_X1    g26680(.A1(new_n26740_), .A2(new_n26747_), .A3(new_n1378_), .ZN(new_n26748_));
  NOR2_X1    g26681(.A1(new_n26457_), .A2(new_n26748_), .ZN(new_n26749_));
  INV_X1     g26682(.I(new_n26748_), .ZN(new_n26750_));
  NOR2_X1    g26683(.A1(new_n26456_), .A2(new_n26750_), .ZN(new_n26751_));
  NOR2_X1    g26684(.A1(new_n26749_), .A2(new_n26751_), .ZN(new_n26752_));
  INV_X1     g26685(.I(new_n26752_), .ZN(new_n26753_));
  XOR2_X1    g26686(.A1(new_n26456_), .A2(new_n26748_), .Z(new_n26754_));
  NOR2_X1    g26687(.A1(new_n26739_), .A2(new_n26754_), .ZN(new_n26755_));
  AOI21_X1   g26688(.A1(new_n26739_), .A2(new_n26753_), .B(new_n26755_), .ZN(new_n26756_));
  INV_X1     g26689(.I(new_n26756_), .ZN(new_n26757_));
  NAND2_X1   g26690(.A1(new_n19415_), .A2(new_n3332_), .ZN(new_n26758_));
  NAND2_X1   g26691(.A1(new_n19407_), .A2(new_n3189_), .ZN(new_n26759_));
  AOI21_X1   g26692(.A1(new_n17790_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n26760_));
  NAND4_X1   g26693(.A1(new_n20846_), .A2(new_n26758_), .A3(new_n26759_), .A4(new_n26760_), .ZN(new_n26761_));
  NAND2_X1   g26694(.A1(new_n26761_), .A2(new_n26757_), .ZN(new_n26762_));
  INV_X1     g26695(.I(new_n26762_), .ZN(new_n26763_));
  NOR2_X1    g26696(.A1(new_n26761_), .A2(new_n26757_), .ZN(new_n26764_));
  NOR2_X1    g26697(.A1(new_n26763_), .A2(new_n26764_), .ZN(new_n26765_));
  INV_X1     g26698(.I(new_n26765_), .ZN(new_n26766_));
  XOR2_X1    g26699(.A1(new_n26761_), .A2(new_n26756_), .Z(new_n26767_));
  NOR2_X1    g26700(.A1(new_n26737_), .A2(new_n26767_), .ZN(new_n26768_));
  AOI21_X1   g26701(.A1(new_n26737_), .A2(new_n26766_), .B(new_n26768_), .ZN(new_n26769_));
  INV_X1     g26702(.I(new_n26769_), .ZN(new_n26770_));
  XOR2_X1    g26703(.A1(new_n26734_), .A2(new_n26770_), .Z(new_n26771_));
  XOR2_X1    g26704(.A1(new_n26771_), .A2(new_n26732_), .Z(new_n26772_));
  XNOR2_X1   g26705(.A1(new_n26772_), .A2(new_n26727_), .ZN(new_n26773_));
  NOR2_X1    g26706(.A1(new_n26627_), .A2(new_n26596_), .ZN(new_n26774_));
  NOR2_X1    g26707(.A1(new_n26774_), .A2(new_n26632_), .ZN(new_n26775_));
  XOR2_X1    g26708(.A1(new_n26773_), .A2(new_n26775_), .Z(new_n26776_));
  OAI22_X1   g26709(.A1(new_n17775_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19475_), .ZN(new_n26777_));
  NAND2_X1   g26710(.A1(new_n21157_), .A2(new_n3312_), .ZN(new_n26778_));
  AOI21_X1   g26711(.A1(new_n26778_), .A2(new_n26777_), .B(new_n3302_), .ZN(new_n26779_));
  NAND2_X1   g26712(.A1(new_n21155_), .A2(new_n26779_), .ZN(new_n26780_));
  XOR2_X1    g26713(.A1(new_n26780_), .A2(\a[23] ), .Z(new_n26781_));
  XOR2_X1    g26714(.A1(new_n26776_), .A2(new_n26781_), .Z(new_n26782_));
  INV_X1     g26715(.I(new_n26781_), .ZN(new_n26783_));
  OR2_X2     g26716(.A1(new_n26776_), .A2(new_n26783_), .Z(new_n26784_));
  NAND2_X1   g26717(.A1(new_n26776_), .A2(new_n26783_), .ZN(new_n26785_));
  NAND2_X1   g26718(.A1(new_n26784_), .A2(new_n26785_), .ZN(new_n26786_));
  NAND2_X1   g26719(.A1(new_n26786_), .A2(new_n26722_), .ZN(new_n26787_));
  OAI21_X1   g26720(.A1(new_n26722_), .A2(new_n26782_), .B(new_n26787_), .ZN(new_n26788_));
  OAI22_X1   g26721(.A1(new_n22115_), .A2(new_n4291_), .B1(new_n4297_), .B2(new_n22149_), .ZN(new_n26789_));
  NAND2_X1   g26722(.A1(new_n23957_), .A2(new_n4469_), .ZN(new_n26790_));
  AOI21_X1   g26723(.A1(new_n26789_), .A2(new_n26790_), .B(new_n4468_), .ZN(new_n26791_));
  NAND2_X1   g26724(.A1(new_n23955_), .A2(new_n26791_), .ZN(new_n26792_));
  XOR2_X1    g26725(.A1(new_n26792_), .A2(\a[17] ), .Z(new_n26793_));
  OAI21_X1   g26726(.A1(new_n26644_), .A2(new_n26652_), .B(new_n26654_), .ZN(new_n26794_));
  OAI22_X1   g26727(.A1(new_n19512_), .A2(new_n3769_), .B1(new_n21960_), .B2(new_n3775_), .ZN(new_n26795_));
  NAND2_X1   g26728(.A1(new_n22048_), .A2(new_n4096_), .ZN(new_n26796_));
  AOI21_X1   g26729(.A1(new_n26796_), .A2(new_n26795_), .B(new_n4095_), .ZN(new_n26797_));
  NAND2_X1   g26730(.A1(new_n22175_), .A2(new_n26797_), .ZN(new_n26798_));
  XOR2_X1    g26731(.A1(new_n26798_), .A2(\a[20] ), .Z(new_n26799_));
  INV_X1     g26732(.I(new_n26799_), .ZN(new_n26800_));
  NOR2_X1    g26733(.A1(new_n26794_), .A2(new_n26800_), .ZN(new_n26801_));
  NAND2_X1   g26734(.A1(new_n26794_), .A2(new_n26800_), .ZN(new_n26802_));
  INV_X1     g26735(.I(new_n26802_), .ZN(new_n26803_));
  NOR2_X1    g26736(.A1(new_n26803_), .A2(new_n26801_), .ZN(new_n26804_));
  NOR2_X1    g26737(.A1(new_n26667_), .A2(new_n26657_), .ZN(new_n26805_));
  NOR2_X1    g26738(.A1(new_n26805_), .A2(new_n26668_), .ZN(new_n26806_));
  XNOR2_X1   g26739(.A1(new_n26806_), .A2(new_n26804_), .ZN(new_n26807_));
  XOR2_X1    g26740(.A1(new_n26807_), .A2(new_n26793_), .Z(new_n26808_));
  XOR2_X1    g26741(.A1(new_n26808_), .A2(new_n26788_), .Z(new_n26809_));
  NAND2_X1   g26742(.A1(new_n26673_), .A2(new_n26680_), .ZN(new_n26810_));
  NAND2_X1   g26743(.A1(new_n26810_), .A2(new_n26681_), .ZN(new_n26811_));
  OAI22_X1   g26744(.A1(new_n24376_), .A2(new_n6094_), .B1(new_n6089_), .B2(new_n24167_), .ZN(new_n26812_));
  NAND2_X1   g26745(.A1(new_n24620_), .A2(new_n6090_), .ZN(new_n26813_));
  AOI21_X1   g26746(.A1(new_n26813_), .A2(new_n26812_), .B(new_n6082_), .ZN(new_n26814_));
  NAND2_X1   g26747(.A1(new_n24618_), .A2(new_n26814_), .ZN(new_n26815_));
  XOR2_X1    g26748(.A1(new_n26815_), .A2(\a[14] ), .Z(new_n26816_));
  INV_X1     g26749(.I(new_n26816_), .ZN(new_n26817_));
  NOR2_X1    g26750(.A1(new_n26811_), .A2(new_n26817_), .ZN(new_n26818_));
  INV_X1     g26751(.I(new_n26818_), .ZN(new_n26819_));
  NAND2_X1   g26752(.A1(new_n26811_), .A2(new_n26817_), .ZN(new_n26820_));
  NAND2_X1   g26753(.A1(new_n26819_), .A2(new_n26820_), .ZN(new_n26821_));
  NAND2_X1   g26754(.A1(new_n26809_), .A2(new_n26821_), .ZN(new_n26822_));
  INV_X1     g26755(.I(new_n26822_), .ZN(new_n26823_));
  XOR2_X1    g26756(.A1(new_n26811_), .A2(new_n26816_), .Z(new_n26824_));
  NOR2_X1    g26757(.A1(new_n26809_), .A2(new_n26824_), .ZN(new_n26825_));
  NOR2_X1    g26758(.A1(new_n26823_), .A2(new_n26825_), .ZN(new_n26826_));
  XOR2_X1    g26759(.A1(new_n26826_), .A2(new_n26720_), .Z(new_n26827_));
  INV_X1     g26760(.I(new_n26593_), .ZN(new_n26828_));
  NAND4_X1   g26761(.A1(new_n26432_), .A2(new_n26441_), .A3(new_n26828_), .A4(new_n26709_), .ZN(new_n26829_));
  XOR2_X1    g26762(.A1(new_n26829_), .A2(new_n26827_), .Z(new_n26830_));
  XOR2_X1    g26763(.A1(new_n26830_), .A2(new_n26718_), .Z(\result[16] ));
  XOR2_X1    g26764(.A1(new_n26827_), .A2(new_n26718_), .Z(new_n26832_));
  INV_X1     g26765(.I(new_n26832_), .ZN(new_n26833_));
  NOR4_X1    g26766(.A1(new_n26442_), .A2(new_n26593_), .A3(new_n26708_), .A4(new_n26833_), .ZN(new_n26834_));
  NOR2_X1    g26767(.A1(new_n26776_), .A2(new_n26783_), .ZN(new_n26835_));
  OAI21_X1   g26768(.A1(new_n26722_), .A2(new_n26835_), .B(new_n26785_), .ZN(new_n26836_));
  AOI21_X1   g26769(.A1(new_n26737_), .A2(new_n26762_), .B(new_n26764_), .ZN(new_n26837_));
  NOR2_X1    g26770(.A1(new_n26739_), .A2(new_n26749_), .ZN(new_n26838_));
  NOR2_X1    g26771(.A1(new_n26838_), .A2(new_n26751_), .ZN(new_n26839_));
  NAND2_X1   g26772(.A1(new_n19439_), .A2(new_n3332_), .ZN(new_n26840_));
  NAND2_X1   g26773(.A1(new_n19415_), .A2(new_n3189_), .ZN(new_n26841_));
  AOI21_X1   g26774(.A1(new_n19407_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n26842_));
  NAND4_X1   g26775(.A1(new_n25294_), .A2(new_n26840_), .A3(new_n26841_), .A4(new_n26842_), .ZN(new_n26843_));
  INV_X1     g26776(.I(new_n11808_), .ZN(new_n26844_));
  NAND3_X1   g26777(.A1(new_n624_), .A2(new_n250_), .A3(new_n1212_), .ZN(new_n26845_));
  NOR4_X1    g26778(.A1(new_n26845_), .A2(new_n214_), .A3(new_n406_), .A4(new_n1262_), .ZN(new_n26846_));
  INV_X1     g26779(.I(new_n1690_), .ZN(new_n26847_));
  INV_X1     g26780(.I(new_n11403_), .ZN(new_n26848_));
  NOR4_X1    g26781(.A1(new_n26848_), .A2(new_n200_), .A3(new_n26847_), .A4(new_n1595_), .ZN(new_n26849_));
  NAND4_X1   g26782(.A1(new_n26849_), .A2(new_n263_), .A3(new_n2691_), .A4(new_n26846_), .ZN(new_n26850_));
  NOR4_X1    g26783(.A1(new_n10997_), .A2(new_n26850_), .A3(new_n24415_), .A4(new_n24872_), .ZN(new_n26851_));
  NAND2_X1   g26784(.A1(new_n26851_), .A2(new_n26844_), .ZN(new_n26852_));
  INV_X1     g26785(.I(new_n26852_), .ZN(new_n26853_));
  NOR2_X1    g26786(.A1(new_n26843_), .A2(new_n26853_), .ZN(new_n26854_));
  NAND2_X1   g26787(.A1(new_n26843_), .A2(new_n26853_), .ZN(new_n26855_));
  INV_X1     g26788(.I(new_n26855_), .ZN(new_n26856_));
  NOR2_X1    g26789(.A1(new_n26856_), .A2(new_n26854_), .ZN(new_n26857_));
  XOR2_X1    g26790(.A1(new_n26843_), .A2(new_n26852_), .Z(new_n26858_));
  MUX2_X1    g26791(.I0(new_n26857_), .I1(new_n26858_), .S(new_n26839_), .Z(new_n26859_));
  OAI22_X1   g26792(.A1(new_n19428_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19423_), .ZN(new_n26860_));
  NAND2_X1   g26793(.A1(new_n19438_), .A2(new_n2750_), .ZN(new_n26861_));
  AOI21_X1   g26794(.A1(new_n26861_), .A2(new_n26860_), .B(new_n2737_), .ZN(new_n26862_));
  NAND2_X1   g26795(.A1(new_n20907_), .A2(new_n26862_), .ZN(new_n26863_));
  XOR2_X1    g26796(.A1(new_n26863_), .A2(\a[29] ), .Z(new_n26864_));
  XNOR2_X1   g26797(.A1(new_n26864_), .A2(new_n26859_), .ZN(new_n26865_));
  NAND2_X1   g26798(.A1(new_n26864_), .A2(new_n26859_), .ZN(new_n26866_));
  OR2_X2     g26799(.A1(new_n26864_), .A2(new_n26859_), .Z(new_n26867_));
  NAND2_X1   g26800(.A1(new_n26867_), .A2(new_n26866_), .ZN(new_n26868_));
  NAND2_X1   g26801(.A1(new_n26868_), .A2(new_n26837_), .ZN(new_n26869_));
  OAI21_X1   g26802(.A1(new_n26837_), .A2(new_n26865_), .B(new_n26869_), .ZN(new_n26870_));
  OAI22_X1   g26803(.A1(new_n19463_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19437_), .ZN(new_n26871_));
  NAND2_X1   g26804(.A1(new_n17780_), .A2(new_n3317_), .ZN(new_n26872_));
  AOI21_X1   g26805(.A1(new_n26871_), .A2(new_n26872_), .B(new_n3260_), .ZN(new_n26873_));
  NAND2_X1   g26806(.A1(new_n21088_), .A2(new_n26873_), .ZN(new_n26874_));
  XOR2_X1    g26807(.A1(new_n26874_), .A2(\a[26] ), .Z(new_n26875_));
  NOR2_X1    g26808(.A1(new_n26734_), .A2(new_n26770_), .ZN(new_n26876_));
  AOI21_X1   g26809(.A1(new_n26771_), .A2(new_n26732_), .B(new_n26876_), .ZN(new_n26877_));
  XNOR2_X1   g26810(.A1(new_n26877_), .A2(new_n26875_), .ZN(new_n26878_));
  XOR2_X1    g26811(.A1(new_n26878_), .A2(new_n26870_), .Z(new_n26879_));
  OAI22_X1   g26812(.A1(new_n19522_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n17775_), .ZN(new_n26880_));
  NAND2_X1   g26813(.A1(new_n17770_), .A2(new_n3312_), .ZN(new_n26881_));
  AOI21_X1   g26814(.A1(new_n26881_), .A2(new_n26880_), .B(new_n3302_), .ZN(new_n26882_));
  NAND2_X1   g26815(.A1(new_n19521_), .A2(new_n26882_), .ZN(new_n26883_));
  XOR2_X1    g26816(.A1(new_n26883_), .A2(\a[23] ), .Z(new_n26884_));
  NOR3_X1    g26817(.A1(new_n26627_), .A2(new_n26596_), .A3(new_n26633_), .ZN(new_n26885_));
  NOR2_X1    g26818(.A1(new_n26885_), .A2(new_n26634_), .ZN(new_n26886_));
  XNOR2_X1   g26819(.A1(new_n26732_), .A2(new_n26769_), .ZN(new_n26887_));
  XOR2_X1    g26820(.A1(new_n26887_), .A2(new_n26734_), .Z(new_n26888_));
  NAND4_X1   g26821(.A1(new_n26772_), .A2(new_n26727_), .A3(new_n26886_), .A4(new_n26888_), .ZN(new_n26889_));
  XOR2_X1    g26822(.A1(new_n26889_), .A2(new_n26884_), .Z(new_n26890_));
  XOR2_X1    g26823(.A1(new_n26879_), .A2(new_n26890_), .Z(new_n26891_));
  AOI22_X1   g26824(.A1(new_n22048_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n21953_), .ZN(new_n26892_));
  NOR2_X1    g26825(.A1(new_n22115_), .A2(new_n4097_), .ZN(new_n26893_));
  OAI21_X1   g26826(.A1(new_n26893_), .A2(new_n26892_), .B(new_n3773_), .ZN(new_n26894_));
  NOR2_X1    g26827(.A1(new_n23675_), .A2(new_n26894_), .ZN(new_n26895_));
  XOR2_X1    g26828(.A1(new_n26895_), .A2(new_n3035_), .Z(new_n26896_));
  INV_X1     g26829(.I(new_n26896_), .ZN(new_n26897_));
  NOR2_X1    g26830(.A1(new_n26897_), .A2(new_n26891_), .ZN(new_n26898_));
  NAND2_X1   g26831(.A1(new_n26897_), .A2(new_n26891_), .ZN(new_n26899_));
  INV_X1     g26832(.I(new_n26899_), .ZN(new_n26900_));
  OAI21_X1   g26833(.A1(new_n26900_), .A2(new_n26898_), .B(new_n26836_), .ZN(new_n26901_));
  XOR2_X1    g26834(.A1(new_n26891_), .A2(new_n26896_), .Z(new_n26902_));
  OAI21_X1   g26835(.A1(new_n26902_), .A2(new_n26836_), .B(new_n26901_), .ZN(new_n26903_));
  OAI21_X1   g26836(.A1(new_n26788_), .A2(new_n26801_), .B(new_n26802_), .ZN(new_n26904_));
  INV_X1     g26837(.I(new_n26904_), .ZN(new_n26905_));
  OAI22_X1   g26838(.A1(new_n23948_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n22149_), .ZN(new_n26906_));
  NAND2_X1   g26839(.A1(new_n24174_), .A2(new_n4469_), .ZN(new_n26907_));
  AOI21_X1   g26840(.A1(new_n26907_), .A2(new_n26906_), .B(new_n4468_), .ZN(new_n26908_));
  NAND2_X1   g26841(.A1(new_n24172_), .A2(new_n26908_), .ZN(new_n26909_));
  XOR2_X1    g26842(.A1(new_n26909_), .A2(\a[17] ), .Z(new_n26910_));
  NAND2_X1   g26843(.A1(new_n26905_), .A2(new_n26910_), .ZN(new_n26911_));
  INV_X1     g26844(.I(new_n26910_), .ZN(new_n26912_));
  NAND2_X1   g26845(.A1(new_n26904_), .A2(new_n26912_), .ZN(new_n26913_));
  NAND2_X1   g26846(.A1(new_n26911_), .A2(new_n26913_), .ZN(new_n26914_));
  NAND2_X1   g26847(.A1(new_n26914_), .A2(new_n26903_), .ZN(new_n26915_));
  XOR2_X1    g26848(.A1(new_n26904_), .A2(new_n26910_), .Z(new_n26916_));
  OR2_X2     g26849(.A1(new_n26916_), .A2(new_n26903_), .Z(new_n26917_));
  NOR2_X1    g26850(.A1(new_n26806_), .A2(new_n26793_), .ZN(new_n26918_));
  NAND2_X1   g26851(.A1(new_n26806_), .A2(new_n26793_), .ZN(new_n26919_));
  XNOR2_X1   g26852(.A1(new_n26788_), .A2(new_n26804_), .ZN(new_n26920_));
  AOI21_X1   g26853(.A1(new_n26920_), .A2(new_n26919_), .B(new_n26918_), .ZN(new_n26921_));
  AOI22_X1   g26854(.A1(new_n24620_), .A2(new_n6095_), .B1(new_n6180_), .B2(new_n24386_), .ZN(new_n26922_));
  NOR2_X1    g26855(.A1(new_n24835_), .A2(new_n6091_), .ZN(new_n26923_));
  OAI21_X1   g26856(.A1(new_n26923_), .A2(new_n26922_), .B(new_n6081_), .ZN(new_n26924_));
  NOR2_X1    g26857(.A1(new_n26554_), .A2(new_n26924_), .ZN(new_n26925_));
  XOR2_X1    g26858(.A1(new_n26925_), .A2(new_n3521_), .Z(new_n26926_));
  NAND2_X1   g26859(.A1(new_n26921_), .A2(new_n26926_), .ZN(new_n26927_));
  OR2_X2     g26860(.A1(new_n26921_), .A2(new_n26926_), .Z(new_n26928_));
  AOI22_X1   g26861(.A1(new_n26928_), .A2(new_n26927_), .B1(new_n26917_), .B2(new_n26915_), .ZN(new_n26929_));
  OAI21_X1   g26862(.A1(new_n26903_), .A2(new_n26916_), .B(new_n26915_), .ZN(new_n26930_));
  XNOR2_X1   g26863(.A1(new_n26921_), .A2(new_n26926_), .ZN(new_n26931_));
  NOR2_X1    g26864(.A1(new_n26931_), .A2(new_n26930_), .ZN(new_n26932_));
  NOR2_X1    g26865(.A1(new_n26932_), .A2(new_n26929_), .ZN(new_n26933_));
  INV_X1     g26866(.I(new_n26933_), .ZN(new_n26934_));
  OAI21_X1   g26867(.A1(new_n26809_), .A2(new_n26818_), .B(new_n26820_), .ZN(new_n26935_));
  NOR2_X1    g26868(.A1(new_n26935_), .A2(new_n26934_), .ZN(new_n26936_));
  XNOR2_X1   g26869(.A1(new_n26808_), .A2(new_n26788_), .ZN(new_n26937_));
  NAND2_X1   g26870(.A1(new_n26937_), .A2(new_n26819_), .ZN(new_n26938_));
  AOI21_X1   g26871(.A1(new_n26938_), .A2(new_n26820_), .B(new_n26933_), .ZN(new_n26939_));
  NOR2_X1    g26872(.A1(new_n26939_), .A2(new_n26936_), .ZN(new_n26940_));
  OAI21_X1   g26873(.A1(new_n26718_), .A2(new_n26826_), .B(new_n26719_), .ZN(new_n26941_));
  XNOR2_X1   g26874(.A1(new_n26941_), .A2(new_n26940_), .ZN(new_n26942_));
  INV_X1     g26875(.I(new_n26942_), .ZN(new_n26943_));
  XOR2_X1    g26876(.A1(new_n26834_), .A2(new_n26943_), .Z(\result[17] ));
  NAND2_X1   g26877(.A1(new_n26834_), .A2(new_n26943_), .ZN(new_n26945_));
  INV_X1     g26878(.I(new_n26898_), .ZN(new_n26946_));
  AOI21_X1   g26879(.A1(new_n26836_), .A2(new_n26946_), .B(new_n26900_), .ZN(new_n26947_));
  INV_X1     g26880(.I(new_n26947_), .ZN(new_n26948_));
  INV_X1     g26881(.I(new_n26837_), .ZN(new_n26949_));
  NAND2_X1   g26882(.A1(new_n26866_), .A2(new_n26949_), .ZN(new_n26950_));
  NAND2_X1   g26883(.A1(new_n26950_), .A2(new_n26867_), .ZN(new_n26951_));
  NOR2_X1    g26884(.A1(new_n26856_), .A2(new_n26839_), .ZN(new_n26952_));
  NOR2_X1    g26885(.A1(new_n26952_), .A2(new_n26854_), .ZN(new_n26953_));
  AOI21_X1   g26886(.A1(new_n19415_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n26954_));
  OAI21_X1   g26887(.A1(new_n17787_), .A2(new_n2767_), .B(new_n26954_), .ZN(new_n26955_));
  AOI21_X1   g26888(.A1(new_n19442_), .A2(new_n3332_), .B(new_n26955_), .ZN(new_n26956_));
  NAND2_X1   g26889(.A1(new_n23413_), .A2(new_n26956_), .ZN(new_n26957_));
  INV_X1     g26890(.I(new_n589_), .ZN(new_n26958_));
  NAND3_X1   g26891(.A1(new_n3101_), .A2(new_n1955_), .A3(new_n10999_), .ZN(new_n26959_));
  NAND4_X1   g26892(.A1(new_n2119_), .A2(new_n436_), .A3(new_n521_), .A4(new_n856_), .ZN(new_n26960_));
  NAND4_X1   g26893(.A1(new_n675_), .A2(new_n707_), .A3(new_n985_), .A4(new_n378_), .ZN(new_n26961_));
  NAND2_X1   g26894(.A1(new_n26960_), .A2(new_n26961_), .ZN(new_n26962_));
  NOR4_X1    g26895(.A1(new_n2094_), .A2(new_n2794_), .A3(new_n26959_), .A4(new_n26962_), .ZN(new_n26963_));
  NAND3_X1   g26896(.A1(new_n26963_), .A2(new_n1731_), .A3(new_n1736_), .ZN(new_n26964_));
  NOR4_X1    g26897(.A1(new_n26964_), .A2(new_n26958_), .A3(new_n19782_), .A4(new_n11057_), .ZN(new_n26965_));
  NAND2_X1   g26898(.A1(new_n26965_), .A2(new_n3029_), .ZN(new_n26966_));
  NAND2_X1   g26899(.A1(new_n26853_), .A2(new_n26966_), .ZN(new_n26967_));
  NAND3_X1   g26900(.A1(new_n26852_), .A2(new_n3029_), .A3(new_n26965_), .ZN(new_n26968_));
  AOI21_X1   g26901(.A1(new_n26967_), .A2(new_n26968_), .B(new_n26957_), .ZN(new_n26969_));
  XNOR2_X1   g26902(.A1(new_n26852_), .A2(new_n26966_), .ZN(new_n26970_));
  AOI21_X1   g26903(.A1(new_n26957_), .A2(new_n26970_), .B(new_n26969_), .ZN(new_n26971_));
  XNOR2_X1   g26904(.A1(new_n26971_), .A2(new_n26953_), .ZN(new_n26972_));
  INV_X1     g26905(.I(new_n26972_), .ZN(new_n26973_));
  INV_X1     g26906(.I(new_n26953_), .ZN(new_n26974_));
  INV_X1     g26907(.I(new_n26971_), .ZN(new_n26975_));
  NOR2_X1    g26908(.A1(new_n26975_), .A2(new_n26974_), .ZN(new_n26976_));
  NOR2_X1    g26909(.A1(new_n26971_), .A2(new_n26953_), .ZN(new_n26977_));
  NOR2_X1    g26910(.A1(new_n26976_), .A2(new_n26977_), .ZN(new_n26978_));
  NOR2_X1    g26911(.A1(new_n26951_), .A2(new_n26978_), .ZN(new_n26979_));
  AOI21_X1   g26912(.A1(new_n26951_), .A2(new_n26973_), .B(new_n26979_), .ZN(new_n26980_));
  OAI22_X1   g26913(.A1(new_n19475_), .A2(new_n3322_), .B1(new_n19463_), .B2(new_n3268_), .ZN(new_n26981_));
  NAND2_X1   g26914(.A1(new_n19484_), .A2(new_n3317_), .ZN(new_n26982_));
  AOI21_X1   g26915(.A1(new_n26982_), .A2(new_n26981_), .B(new_n3260_), .ZN(new_n26983_));
  NAND2_X1   g26916(.A1(new_n21171_), .A2(new_n26983_), .ZN(new_n26984_));
  XOR2_X1    g26917(.A1(new_n26984_), .A2(new_n72_), .Z(new_n26985_));
  OAI22_X1   g26918(.A1(new_n17784_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19428_), .ZN(new_n26986_));
  NAND2_X1   g26919(.A1(new_n19466_), .A2(new_n2750_), .ZN(new_n26987_));
  AOI21_X1   g26920(.A1(new_n26987_), .A2(new_n26986_), .B(new_n2737_), .ZN(new_n26988_));
  NAND2_X1   g26921(.A1(new_n21100_), .A2(new_n26988_), .ZN(new_n26989_));
  XOR2_X1    g26922(.A1(new_n26989_), .A2(\a[29] ), .Z(new_n26990_));
  XOR2_X1    g26923(.A1(new_n26985_), .A2(new_n26990_), .Z(new_n26991_));
  NOR2_X1    g26924(.A1(new_n26991_), .A2(new_n26980_), .ZN(new_n26992_));
  INV_X1     g26925(.I(new_n26990_), .ZN(new_n26993_));
  NOR2_X1    g26926(.A1(new_n26985_), .A2(new_n26993_), .ZN(new_n26994_));
  INV_X1     g26927(.I(new_n26994_), .ZN(new_n26995_));
  NAND2_X1   g26928(.A1(new_n26985_), .A2(new_n26993_), .ZN(new_n26996_));
  NAND2_X1   g26929(.A1(new_n26995_), .A2(new_n26996_), .ZN(new_n26997_));
  AOI21_X1   g26930(.A1(new_n26980_), .A2(new_n26997_), .B(new_n26992_), .ZN(new_n26998_));
  OAI22_X1   g26931(.A1(new_n19512_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n19522_), .ZN(new_n26999_));
  NAND2_X1   g26932(.A1(new_n21953_), .A2(new_n3312_), .ZN(new_n27000_));
  AOI21_X1   g26933(.A1(new_n26999_), .A2(new_n27000_), .B(new_n3302_), .ZN(new_n27001_));
  NAND2_X1   g26934(.A1(new_n21963_), .A2(new_n27001_), .ZN(new_n27002_));
  XOR2_X1    g26935(.A1(new_n27002_), .A2(\a[23] ), .Z(new_n27003_));
  XNOR2_X1   g26936(.A1(new_n26998_), .A2(new_n27003_), .ZN(new_n27004_));
  INV_X1     g26937(.I(new_n26889_), .ZN(new_n27005_));
  XOR2_X1    g26938(.A1(new_n26879_), .A2(new_n26884_), .Z(new_n27006_));
  OAI21_X1   g26939(.A1(new_n26884_), .A2(new_n27005_), .B(new_n27006_), .ZN(new_n27007_));
  OAI22_X1   g26940(.A1(new_n22115_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n22051_), .ZN(new_n27008_));
  NAND2_X1   g26941(.A1(new_n22150_), .A2(new_n4096_), .ZN(new_n27009_));
  AOI21_X1   g26942(.A1(new_n27008_), .A2(new_n27009_), .B(new_n4095_), .ZN(new_n27010_));
  NAND2_X1   g26943(.A1(new_n22163_), .A2(new_n27010_), .ZN(new_n27011_));
  XOR2_X1    g26944(.A1(new_n27011_), .A2(\a[20] ), .Z(new_n27012_));
  NAND2_X1   g26945(.A1(new_n27007_), .A2(new_n27012_), .ZN(new_n27013_));
  INV_X1     g26946(.I(new_n27007_), .ZN(new_n27014_));
  INV_X1     g26947(.I(new_n27012_), .ZN(new_n27015_));
  NAND2_X1   g26948(.A1(new_n27014_), .A2(new_n27015_), .ZN(new_n27016_));
  AOI21_X1   g26949(.A1(new_n27016_), .A2(new_n27013_), .B(new_n27004_), .ZN(new_n27017_));
  INV_X1     g26950(.I(new_n27004_), .ZN(new_n27018_));
  XOR2_X1    g26951(.A1(new_n27007_), .A2(new_n27015_), .Z(new_n27019_));
  NOR2_X1    g26952(.A1(new_n27019_), .A2(new_n27018_), .ZN(new_n27020_));
  NOR2_X1    g26953(.A1(new_n27020_), .A2(new_n27017_), .ZN(new_n27021_));
  AOI22_X1   g26954(.A1(new_n24174_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n23957_), .ZN(new_n27022_));
  NOR2_X1    g26955(.A1(new_n24376_), .A2(new_n4470_), .ZN(new_n27023_));
  OAI21_X1   g26956(.A1(new_n27023_), .A2(new_n27022_), .B(new_n4295_), .ZN(new_n27024_));
  NOR2_X1    g26957(.A1(new_n24391_), .A2(new_n27024_), .ZN(new_n27025_));
  XOR2_X1    g26958(.A1(new_n27025_), .A2(new_n3372_), .Z(new_n27026_));
  NAND2_X1   g26959(.A1(new_n27021_), .A2(new_n27026_), .ZN(new_n27027_));
  NOR2_X1    g26960(.A1(new_n27021_), .A2(new_n27026_), .ZN(new_n27028_));
  INV_X1     g26961(.I(new_n27028_), .ZN(new_n27029_));
  NAND2_X1   g26962(.A1(new_n27029_), .A2(new_n27027_), .ZN(new_n27030_));
  NAND2_X1   g26963(.A1(new_n27030_), .A2(new_n26948_), .ZN(new_n27031_));
  XNOR2_X1   g26964(.A1(new_n27021_), .A2(new_n27026_), .ZN(new_n27032_));
  OAI21_X1   g26965(.A1(new_n26948_), .A2(new_n27032_), .B(new_n27031_), .ZN(new_n27033_));
  INV_X1     g26966(.I(new_n26913_), .ZN(new_n27034_));
  AND2_X2    g26967(.A1(new_n26911_), .A2(new_n26903_), .Z(new_n27035_));
  NOR2_X1    g26968(.A1(new_n27035_), .A2(new_n27034_), .ZN(new_n27036_));
  INV_X1     g26969(.I(new_n27036_), .ZN(new_n27037_));
  AOI22_X1   g26970(.A1(new_n24826_), .A2(new_n11496_), .B1(new_n6180_), .B2(new_n24620_), .ZN(new_n27038_));
  OR3_X2     g26971(.A1(new_n25017_), .A2(new_n6082_), .A3(new_n27038_), .Z(new_n27039_));
  XOR2_X1    g26972(.A1(new_n27039_), .A2(\a[14] ), .Z(new_n27040_));
  INV_X1     g26973(.I(new_n27040_), .ZN(new_n27041_));
  NOR2_X1    g26974(.A1(new_n27037_), .A2(new_n27041_), .ZN(new_n27042_));
  NOR2_X1    g26975(.A1(new_n27036_), .A2(new_n27040_), .ZN(new_n27043_));
  OAI21_X1   g26976(.A1(new_n27042_), .A2(new_n27043_), .B(new_n27033_), .ZN(new_n27044_));
  XOR2_X1    g26977(.A1(new_n27036_), .A2(new_n27041_), .Z(new_n27045_));
  OR2_X2     g26978(.A1(new_n27045_), .A2(new_n27033_), .Z(new_n27046_));
  NAND2_X1   g26979(.A1(new_n27046_), .A2(new_n27044_), .ZN(new_n27047_));
  NAND2_X1   g26980(.A1(new_n26930_), .A2(new_n26927_), .ZN(new_n27048_));
  NAND2_X1   g26981(.A1(new_n27048_), .A2(new_n26928_), .ZN(new_n27049_));
  OAI21_X1   g26982(.A1(new_n26823_), .A2(new_n26825_), .B(new_n26720_), .ZN(new_n27050_));
  OR2_X2     g26983(.A1(new_n26809_), .A2(new_n26824_), .Z(new_n27051_));
  AOI21_X1   g26984(.A1(new_n27051_), .A2(new_n26822_), .B(new_n26719_), .ZN(new_n27052_));
  NOR3_X1    g26985(.A1(new_n27052_), .A2(new_n26936_), .A3(new_n26939_), .ZN(new_n27053_));
  OAI21_X1   g26986(.A1(new_n26718_), .A2(new_n27050_), .B(new_n27053_), .ZN(new_n27054_));
  NOR2_X1    g26987(.A1(new_n27054_), .A2(new_n26936_), .ZN(new_n27055_));
  XOR2_X1    g26988(.A1(new_n27055_), .A2(new_n27049_), .Z(new_n27056_));
  XOR2_X1    g26989(.A1(new_n27056_), .A2(new_n27047_), .Z(new_n27057_));
  XOR2_X1    g26990(.A1(new_n26945_), .A2(new_n27057_), .Z(\result[18] ));
  OR3_X2     g26991(.A1(new_n26589_), .A2(new_n26702_), .A3(new_n26581_), .Z(new_n27059_));
  AOI21_X1   g26992(.A1(new_n26279_), .A2(new_n26702_), .B(new_n27059_), .ZN(new_n27060_));
  INV_X1     g26993(.I(new_n26712_), .ZN(new_n27061_));
  INV_X1     g26994(.I(new_n26695_), .ZN(new_n27062_));
  XOR2_X1    g26995(.A1(new_n26687_), .A2(new_n26690_), .Z(new_n27063_));
  NOR2_X1    g26996(.A1(new_n27063_), .A2(new_n26686_), .ZN(new_n27064_));
  OAI21_X1   g26997(.A1(new_n27062_), .A2(new_n27064_), .B(new_n26700_), .ZN(new_n27065_));
  AOI21_X1   g26998(.A1(new_n27065_), .A2(new_n26714_), .B(new_n26581_), .ZN(new_n27066_));
  AOI21_X1   g26999(.A1(new_n27060_), .A2(new_n27066_), .B(new_n27061_), .ZN(new_n27067_));
  NAND2_X1   g27000(.A1(new_n26940_), .A2(new_n27050_), .ZN(new_n27068_));
  AOI21_X1   g27001(.A1(new_n27067_), .A2(new_n27052_), .B(new_n27068_), .ZN(new_n27069_));
  AOI21_X1   g27002(.A1(new_n27046_), .A2(new_n27044_), .B(new_n27049_), .ZN(new_n27070_));
  NAND3_X1   g27003(.A1(new_n27046_), .A2(new_n27044_), .A3(new_n27049_), .ZN(new_n27071_));
  AOI21_X1   g27004(.A1(new_n27046_), .A2(new_n27044_), .B(new_n27049_), .ZN(new_n27072_));
  INV_X1     g27005(.I(new_n27072_), .ZN(new_n27073_));
  AOI21_X1   g27006(.A1(new_n27073_), .A2(new_n27071_), .B(new_n26936_), .ZN(new_n27074_));
  AOI21_X1   g27007(.A1(new_n27069_), .A2(new_n27074_), .B(new_n27070_), .ZN(new_n27075_));
  OAI21_X1   g27008(.A1(new_n27037_), .A2(new_n27041_), .B(new_n27033_), .ZN(new_n27076_));
  OAI21_X1   g27009(.A1(new_n27036_), .A2(new_n27040_), .B(new_n27076_), .ZN(new_n27077_));
  AOI21_X1   g27010(.A1(new_n27021_), .A2(new_n27026_), .B(new_n26947_), .ZN(new_n27078_));
  NOR2_X1    g27011(.A1(new_n27078_), .A2(new_n27028_), .ZN(new_n27079_));
  INV_X1     g27012(.I(new_n27079_), .ZN(new_n27080_));
  NOR2_X1    g27013(.A1(new_n26998_), .A2(new_n27003_), .ZN(new_n27081_));
  OAI22_X1   g27014(.A1(new_n19512_), .A2(new_n3310_), .B1(new_n21960_), .B2(new_n3306_), .ZN(new_n27082_));
  NAND2_X1   g27015(.A1(new_n22048_), .A2(new_n3312_), .ZN(new_n27083_));
  AOI21_X1   g27016(.A1(new_n27083_), .A2(new_n27082_), .B(new_n3302_), .ZN(new_n27084_));
  NAND2_X1   g27017(.A1(new_n22175_), .A2(new_n27084_), .ZN(new_n27085_));
  XOR2_X1    g27018(.A1(new_n27085_), .A2(\a[23] ), .Z(new_n27086_));
  INV_X1     g27019(.I(new_n27086_), .ZN(new_n27087_));
  NOR2_X1    g27020(.A1(new_n27087_), .A2(new_n27081_), .ZN(new_n27088_));
  NAND2_X1   g27021(.A1(new_n27087_), .A2(new_n27081_), .ZN(new_n27089_));
  INV_X1     g27022(.I(new_n27089_), .ZN(new_n27090_));
  NOR2_X1    g27023(.A1(new_n27090_), .A2(new_n27088_), .ZN(new_n27091_));
  OAI21_X1   g27024(.A1(new_n26974_), .A2(new_n26975_), .B(new_n26951_), .ZN(new_n27092_));
  OAI21_X1   g27025(.A1(new_n26953_), .A2(new_n26971_), .B(new_n27092_), .ZN(new_n27093_));
  NOR2_X1    g27026(.A1(new_n24835_), .A2(new_n11497_), .ZN(new_n27094_));
  OAI22_X1   g27027(.A1(new_n27094_), .A2(\a[14] ), .B1(new_n11499_), .B2(new_n24835_), .ZN(new_n27095_));
  INV_X1     g27028(.I(new_n1280_), .ZN(new_n27096_));
  NAND3_X1   g27029(.A1(new_n2946_), .A2(new_n1871_), .A3(new_n745_), .ZN(new_n27097_));
  NOR3_X1    g27030(.A1(new_n801_), .A2(new_n764_), .A3(new_n310_), .ZN(new_n27098_));
  NAND4_X1   g27031(.A1(new_n12152_), .A2(new_n1205_), .A3(new_n11856_), .A4(new_n27098_), .ZN(new_n27099_));
  NAND2_X1   g27032(.A1(new_n4858_), .A2(new_n2443_), .ZN(new_n27100_));
  NOR4_X1    g27033(.A1(new_n27100_), .A2(new_n12514_), .A3(new_n27097_), .A4(new_n27099_), .ZN(new_n27101_));
  AOI21_X1   g27034(.A1(new_n27096_), .A2(new_n27101_), .B(new_n26853_), .ZN(new_n27102_));
  NAND2_X1   g27035(.A1(new_n27096_), .A2(new_n27101_), .ZN(new_n27103_));
  NOR2_X1    g27036(.A1(new_n26852_), .A2(new_n27103_), .ZN(new_n27104_));
  NOR2_X1    g27037(.A1(new_n27102_), .A2(new_n27104_), .ZN(new_n27105_));
  INV_X1     g27038(.I(new_n27105_), .ZN(new_n27106_));
  XNOR2_X1   g27039(.A1(new_n26852_), .A2(new_n27103_), .ZN(new_n27107_));
  NOR2_X1    g27040(.A1(new_n27095_), .A2(new_n27107_), .ZN(new_n27108_));
  AOI21_X1   g27041(.A1(new_n27095_), .A2(new_n27106_), .B(new_n27108_), .ZN(new_n27109_));
  NAND3_X1   g27042(.A1(new_n23413_), .A2(new_n26956_), .A3(new_n26967_), .ZN(new_n27110_));
  NAND2_X1   g27043(.A1(new_n27110_), .A2(new_n26968_), .ZN(new_n27111_));
  INV_X1     g27044(.I(new_n22226_), .ZN(new_n27112_));
  NOR2_X1    g27045(.A1(new_n19428_), .A2(new_n2772_), .ZN(new_n27113_));
  NOR2_X1    g27046(.A1(new_n19423_), .A2(new_n2767_), .ZN(new_n27114_));
  OAI21_X1   g27047(.A1(new_n17787_), .A2(new_n2771_), .B(new_n2764_), .ZN(new_n27115_));
  NOR4_X1    g27048(.A1(new_n27112_), .A2(new_n27113_), .A3(new_n27114_), .A4(new_n27115_), .ZN(new_n27116_));
  XNOR2_X1   g27049(.A1(new_n27116_), .A2(new_n27111_), .ZN(new_n27117_));
  NOR2_X1    g27050(.A1(new_n27117_), .A2(new_n27109_), .ZN(new_n27118_));
  INV_X1     g27051(.I(new_n27109_), .ZN(new_n27119_));
  NOR2_X1    g27052(.A1(new_n27116_), .A2(new_n27111_), .ZN(new_n27120_));
  INV_X1     g27053(.I(new_n27120_), .ZN(new_n27121_));
  NAND2_X1   g27054(.A1(new_n27116_), .A2(new_n27111_), .ZN(new_n27122_));
  AOI21_X1   g27055(.A1(new_n27121_), .A2(new_n27122_), .B(new_n27119_), .ZN(new_n27123_));
  NOR2_X1    g27056(.A1(new_n27118_), .A2(new_n27123_), .ZN(new_n27124_));
  OAI22_X1   g27057(.A1(new_n19437_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n17784_), .ZN(new_n27125_));
  NAND2_X1   g27058(.A1(new_n19472_), .A2(new_n2750_), .ZN(new_n27126_));
  AOI21_X1   g27059(.A1(new_n27126_), .A2(new_n27125_), .B(new_n2737_), .ZN(new_n27127_));
  NAND2_X1   g27060(.A1(new_n21117_), .A2(new_n27127_), .ZN(new_n27128_));
  XOR2_X1    g27061(.A1(new_n27128_), .A2(\a[29] ), .Z(new_n27129_));
  XNOR2_X1   g27062(.A1(new_n27124_), .A2(new_n27129_), .ZN(new_n27130_));
  INV_X1     g27063(.I(new_n27130_), .ZN(new_n27131_));
  INV_X1     g27064(.I(new_n27124_), .ZN(new_n27132_));
  INV_X1     g27065(.I(new_n27129_), .ZN(new_n27133_));
  NOR2_X1    g27066(.A1(new_n27132_), .A2(new_n27133_), .ZN(new_n27134_));
  NOR2_X1    g27067(.A1(new_n27124_), .A2(new_n27129_), .ZN(new_n27135_));
  NOR2_X1    g27068(.A1(new_n27134_), .A2(new_n27135_), .ZN(new_n27136_));
  NOR2_X1    g27069(.A1(new_n27093_), .A2(new_n27136_), .ZN(new_n27137_));
  AOI21_X1   g27070(.A1(new_n27093_), .A2(new_n27131_), .B(new_n27137_), .ZN(new_n27138_));
  INV_X1     g27071(.I(new_n26996_), .ZN(new_n27139_));
  AOI21_X1   g27072(.A1(new_n26980_), .A2(new_n26995_), .B(new_n27139_), .ZN(new_n27140_));
  OAI22_X1   g27073(.A1(new_n17775_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19475_), .ZN(new_n27141_));
  NAND2_X1   g27074(.A1(new_n21157_), .A2(new_n3317_), .ZN(new_n27142_));
  AOI21_X1   g27075(.A1(new_n27142_), .A2(new_n27141_), .B(new_n3260_), .ZN(new_n27143_));
  NAND2_X1   g27076(.A1(new_n21155_), .A2(new_n27143_), .ZN(new_n27144_));
  XOR2_X1    g27077(.A1(new_n27144_), .A2(\a[26] ), .Z(new_n27145_));
  NAND2_X1   g27078(.A1(new_n27140_), .A2(new_n27145_), .ZN(new_n27146_));
  NOR2_X1    g27079(.A1(new_n27140_), .A2(new_n27145_), .ZN(new_n27147_));
  INV_X1     g27080(.I(new_n27147_), .ZN(new_n27148_));
  AOI21_X1   g27081(.A1(new_n27148_), .A2(new_n27146_), .B(new_n27138_), .ZN(new_n27149_));
  INV_X1     g27082(.I(new_n27138_), .ZN(new_n27150_));
  XNOR2_X1   g27083(.A1(new_n27140_), .A2(new_n27145_), .ZN(new_n27151_));
  NOR2_X1    g27084(.A1(new_n27151_), .A2(new_n27150_), .ZN(new_n27152_));
  NOR2_X1    g27085(.A1(new_n27152_), .A2(new_n27149_), .ZN(new_n27153_));
  INV_X1     g27086(.I(new_n27153_), .ZN(new_n27154_));
  OAI22_X1   g27087(.A1(new_n22115_), .A2(new_n3769_), .B1(new_n3775_), .B2(new_n22149_), .ZN(new_n27155_));
  NAND2_X1   g27088(.A1(new_n23957_), .A2(new_n4096_), .ZN(new_n27156_));
  AOI21_X1   g27089(.A1(new_n27155_), .A2(new_n27156_), .B(new_n4095_), .ZN(new_n27157_));
  NAND2_X1   g27090(.A1(new_n23955_), .A2(new_n27157_), .ZN(new_n27158_));
  XOR2_X1    g27091(.A1(new_n27158_), .A2(\a[20] ), .Z(new_n27159_));
  XOR2_X1    g27092(.A1(new_n27159_), .A2(new_n27154_), .Z(new_n27160_));
  NOR2_X1    g27093(.A1(new_n27160_), .A2(new_n27091_), .ZN(new_n27161_));
  XOR2_X1    g27094(.A1(new_n27159_), .A2(new_n27153_), .Z(new_n27162_));
  NOR3_X1    g27095(.A1(new_n27162_), .A2(new_n27088_), .A3(new_n27090_), .ZN(new_n27163_));
  NOR2_X1    g27096(.A1(new_n27163_), .A2(new_n27161_), .ZN(new_n27164_));
  NAND2_X1   g27097(.A1(new_n27014_), .A2(new_n27018_), .ZN(new_n27165_));
  XNOR2_X1   g27098(.A1(new_n27164_), .A2(new_n27165_), .ZN(new_n27166_));
  XOR2_X1    g27099(.A1(new_n27007_), .A2(new_n27018_), .Z(new_n27167_));
  NOR2_X1    g27100(.A1(new_n27167_), .A2(new_n27012_), .ZN(new_n27168_));
  AND2_X2    g27101(.A1(new_n27166_), .A2(new_n27168_), .Z(new_n27169_));
  NOR2_X1    g27102(.A1(new_n27166_), .A2(new_n27168_), .ZN(new_n27170_));
  NOR2_X1    g27103(.A1(new_n27169_), .A2(new_n27170_), .ZN(new_n27171_));
  OAI22_X1   g27104(.A1(new_n24376_), .A2(new_n4297_), .B1(new_n4291_), .B2(new_n24167_), .ZN(new_n27172_));
  NAND2_X1   g27105(.A1(new_n24620_), .A2(new_n4469_), .ZN(new_n27173_));
  AOI21_X1   g27106(.A1(new_n27173_), .A2(new_n27172_), .B(new_n4468_), .ZN(new_n27174_));
  NAND2_X1   g27107(.A1(new_n24618_), .A2(new_n27174_), .ZN(new_n27175_));
  XOR2_X1    g27108(.A1(new_n27175_), .A2(\a[17] ), .Z(new_n27176_));
  INV_X1     g27109(.I(new_n27176_), .ZN(new_n27177_));
  XOR2_X1    g27110(.A1(new_n27171_), .A2(new_n27177_), .Z(new_n27178_));
  INV_X1     g27111(.I(new_n27171_), .ZN(new_n27179_));
  NAND2_X1   g27112(.A1(new_n27179_), .A2(new_n27176_), .ZN(new_n27180_));
  NAND2_X1   g27113(.A1(new_n27171_), .A2(new_n27177_), .ZN(new_n27181_));
  AOI21_X1   g27114(.A1(new_n27180_), .A2(new_n27181_), .B(new_n27080_), .ZN(new_n27182_));
  AOI21_X1   g27115(.A1(new_n27080_), .A2(new_n27178_), .B(new_n27182_), .ZN(new_n27183_));
  XNOR2_X1   g27116(.A1(new_n27183_), .A2(new_n27077_), .ZN(new_n27184_));
  NOR4_X1    g27117(.A1(new_n26829_), .A2(new_n26833_), .A3(new_n26942_), .A4(new_n27057_), .ZN(new_n27185_));
  XOR2_X1    g27118(.A1(new_n27185_), .A2(new_n27184_), .Z(new_n27186_));
  XOR2_X1    g27119(.A1(new_n27186_), .A2(new_n27075_), .Z(\result[19] ));
  INV_X1     g27120(.I(new_n27057_), .ZN(new_n27188_));
  INV_X1     g27121(.I(new_n27070_), .ZN(new_n27189_));
  INV_X1     g27122(.I(new_n27071_), .ZN(new_n27190_));
  OAI22_X1   g27123(.A1(new_n27190_), .A2(new_n27072_), .B1(new_n26934_), .B2(new_n26935_), .ZN(new_n27191_));
  OAI21_X1   g27124(.A1(new_n27054_), .A2(new_n27191_), .B(new_n27189_), .ZN(new_n27192_));
  XOR2_X1    g27125(.A1(new_n27192_), .A2(new_n27184_), .Z(new_n27193_));
  NAND4_X1   g27126(.A1(new_n26834_), .A2(new_n26943_), .A3(new_n27188_), .A4(new_n27193_), .ZN(new_n27194_));
  INV_X1     g27127(.I(new_n27134_), .ZN(new_n27195_));
  AOI21_X1   g27128(.A1(new_n27093_), .A2(new_n27195_), .B(new_n27135_), .ZN(new_n27196_));
  INV_X1     g27129(.I(new_n27196_), .ZN(new_n27197_));
  NOR2_X1    g27130(.A1(new_n27095_), .A2(new_n27102_), .ZN(new_n27198_));
  NOR2_X1    g27131(.A1(new_n27198_), .A2(new_n27104_), .ZN(new_n27199_));
  NOR2_X1    g27132(.A1(new_n17784_), .A2(new_n2772_), .ZN(new_n27200_));
  NOR2_X1    g27133(.A1(new_n19428_), .A2(new_n2767_), .ZN(new_n27201_));
  NOR2_X1    g27134(.A1(new_n19423_), .A2(new_n2771_), .ZN(new_n27202_));
  NOR4_X1    g27135(.A1(new_n27200_), .A2(new_n2764_), .A3(new_n27201_), .A4(new_n27202_), .ZN(new_n27203_));
  NOR4_X1    g27136(.A1(new_n576_), .A2(new_n663_), .A3(new_n1620_), .A4(new_n1784_), .ZN(new_n27204_));
  NAND4_X1   g27137(.A1(new_n3198_), .A2(new_n1189_), .A3(new_n395_), .A4(new_n1436_), .ZN(new_n27205_));
  INV_X1     g27138(.I(new_n619_), .ZN(new_n27206_));
  NOR4_X1    g27139(.A1(new_n27206_), .A2(new_n650_), .A3(new_n1185_), .A4(new_n1902_), .ZN(new_n27207_));
  NAND4_X1   g27140(.A1(new_n27207_), .A2(new_n1402_), .A3(new_n27204_), .A4(new_n27205_), .ZN(new_n27208_));
  NAND2_X1   g27141(.A1(new_n11925_), .A2(new_n4380_), .ZN(new_n27209_));
  NOR4_X1    g27142(.A1(new_n27209_), .A2(new_n27208_), .A3(new_n4744_), .A4(new_n3854_), .ZN(new_n27210_));
  INV_X1     g27143(.I(new_n27210_), .ZN(new_n27211_));
  NAND3_X1   g27144(.A1(new_n21621_), .A2(new_n27203_), .A3(new_n27211_), .ZN(new_n27212_));
  NAND2_X1   g27145(.A1(new_n21621_), .A2(new_n27203_), .ZN(new_n27213_));
  NAND2_X1   g27146(.A1(new_n27213_), .A2(new_n27210_), .ZN(new_n27214_));
  AOI21_X1   g27147(.A1(new_n27214_), .A2(new_n27212_), .B(new_n27199_), .ZN(new_n27215_));
  XOR2_X1    g27148(.A1(new_n27213_), .A2(new_n27211_), .Z(new_n27216_));
  NOR3_X1    g27149(.A1(new_n27216_), .A2(new_n27104_), .A3(new_n27198_), .ZN(new_n27217_));
  NOR2_X1    g27150(.A1(new_n27217_), .A2(new_n27215_), .ZN(new_n27218_));
  OAI21_X1   g27151(.A1(new_n27119_), .A2(new_n27120_), .B(new_n27122_), .ZN(new_n27219_));
  OAI22_X1   g27152(.A1(new_n19463_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19437_), .ZN(new_n27220_));
  NAND2_X1   g27153(.A1(new_n17780_), .A2(new_n2750_), .ZN(new_n27221_));
  AOI21_X1   g27154(.A1(new_n27220_), .A2(new_n27221_), .B(new_n2737_), .ZN(new_n27222_));
  NAND2_X1   g27155(.A1(new_n21088_), .A2(new_n27222_), .ZN(new_n27223_));
  XOR2_X1    g27156(.A1(new_n27223_), .A2(\a[29] ), .Z(new_n27224_));
  XOR2_X1    g27157(.A1(new_n27224_), .A2(new_n27219_), .Z(new_n27225_));
  NOR2_X1    g27158(.A1(new_n27225_), .A2(new_n27218_), .ZN(new_n27226_));
  INV_X1     g27159(.I(new_n27218_), .ZN(new_n27227_));
  INV_X1     g27160(.I(new_n27224_), .ZN(new_n27228_));
  NOR2_X1    g27161(.A1(new_n27228_), .A2(new_n27219_), .ZN(new_n27229_));
  INV_X1     g27162(.I(new_n27229_), .ZN(new_n27230_));
  NAND2_X1   g27163(.A1(new_n27228_), .A2(new_n27219_), .ZN(new_n27231_));
  AOI21_X1   g27164(.A1(new_n27230_), .A2(new_n27231_), .B(new_n27227_), .ZN(new_n27232_));
  NOR2_X1    g27165(.A1(new_n27232_), .A2(new_n27226_), .ZN(new_n27233_));
  INV_X1     g27166(.I(new_n27233_), .ZN(new_n27234_));
  OAI22_X1   g27167(.A1(new_n19522_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n17775_), .ZN(new_n27235_));
  NAND2_X1   g27168(.A1(new_n17770_), .A2(new_n3317_), .ZN(new_n27236_));
  AOI21_X1   g27169(.A1(new_n27236_), .A2(new_n27235_), .B(new_n3260_), .ZN(new_n27237_));
  NAND2_X1   g27170(.A1(new_n19521_), .A2(new_n27237_), .ZN(new_n27238_));
  XOR2_X1    g27171(.A1(new_n27238_), .A2(\a[26] ), .Z(new_n27239_));
  NAND2_X1   g27172(.A1(new_n27234_), .A2(new_n27239_), .ZN(new_n27240_));
  NOR2_X1    g27173(.A1(new_n27234_), .A2(new_n27239_), .ZN(new_n27241_));
  INV_X1     g27174(.I(new_n27241_), .ZN(new_n27242_));
  NAND2_X1   g27175(.A1(new_n27242_), .A2(new_n27240_), .ZN(new_n27243_));
  NAND2_X1   g27176(.A1(new_n27243_), .A2(new_n27197_), .ZN(new_n27244_));
  XOR2_X1    g27177(.A1(new_n27233_), .A2(new_n27239_), .Z(new_n27245_));
  OAI21_X1   g27178(.A1(new_n27197_), .A2(new_n27245_), .B(new_n27244_), .ZN(new_n27246_));
  INV_X1     g27179(.I(new_n27246_), .ZN(new_n27247_));
  NAND2_X1   g27180(.A1(new_n27138_), .A2(new_n27146_), .ZN(new_n27248_));
  NAND2_X1   g27181(.A1(new_n27248_), .A2(new_n27148_), .ZN(new_n27249_));
  AOI22_X1   g27182(.A1(new_n22048_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n21953_), .ZN(new_n27250_));
  NOR2_X1    g27183(.A1(new_n22115_), .A2(new_n3780_), .ZN(new_n27251_));
  OAI21_X1   g27184(.A1(new_n27251_), .A2(new_n27250_), .B(new_n3301_), .ZN(new_n27252_));
  NOR2_X1    g27185(.A1(new_n23675_), .A2(new_n27252_), .ZN(new_n27253_));
  XOR2_X1    g27186(.A1(new_n27253_), .A2(new_n84_), .Z(new_n27254_));
  INV_X1     g27187(.I(new_n27254_), .ZN(new_n27255_));
  NOR2_X1    g27188(.A1(new_n27255_), .A2(new_n27249_), .ZN(new_n27256_));
  INV_X1     g27189(.I(new_n27256_), .ZN(new_n27257_));
  NAND2_X1   g27190(.A1(new_n27255_), .A2(new_n27249_), .ZN(new_n27258_));
  AOI21_X1   g27191(.A1(new_n27257_), .A2(new_n27258_), .B(new_n27247_), .ZN(new_n27259_));
  XOR2_X1    g27192(.A1(new_n27254_), .A2(new_n27249_), .Z(new_n27260_));
  INV_X1     g27193(.I(new_n27260_), .ZN(new_n27261_));
  AOI21_X1   g27194(.A1(new_n27247_), .A2(new_n27261_), .B(new_n27259_), .ZN(new_n27262_));
  INV_X1     g27195(.I(new_n27262_), .ZN(new_n27263_));
  OAI21_X1   g27196(.A1(new_n27154_), .A2(new_n27088_), .B(new_n27089_), .ZN(new_n27264_));
  OAI22_X1   g27197(.A1(new_n23948_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n22149_), .ZN(new_n27265_));
  NAND2_X1   g27198(.A1(new_n24174_), .A2(new_n4096_), .ZN(new_n27266_));
  AOI21_X1   g27199(.A1(new_n27266_), .A2(new_n27265_), .B(new_n4095_), .ZN(new_n27267_));
  NAND2_X1   g27200(.A1(new_n24172_), .A2(new_n27267_), .ZN(new_n27268_));
  XOR2_X1    g27201(.A1(new_n27268_), .A2(\a[20] ), .Z(new_n27269_));
  INV_X1     g27202(.I(new_n27269_), .ZN(new_n27270_));
  NOR2_X1    g27203(.A1(new_n27270_), .A2(new_n27264_), .ZN(new_n27271_));
  NAND2_X1   g27204(.A1(new_n27270_), .A2(new_n27264_), .ZN(new_n27272_));
  INV_X1     g27205(.I(new_n27272_), .ZN(new_n27273_));
  OAI21_X1   g27206(.A1(new_n27271_), .A2(new_n27273_), .B(new_n27263_), .ZN(new_n27274_));
  XOR2_X1    g27207(.A1(new_n27269_), .A2(new_n27264_), .Z(new_n27275_));
  OAI21_X1   g27208(.A1(new_n27263_), .A2(new_n27275_), .B(new_n27274_), .ZN(new_n27276_));
  AOI22_X1   g27209(.A1(new_n24620_), .A2(new_n4298_), .B1(new_n4292_), .B2(new_n24386_), .ZN(new_n27277_));
  NOR2_X1    g27210(.A1(new_n24835_), .A2(new_n4470_), .ZN(new_n27278_));
  OAI21_X1   g27211(.A1(new_n27278_), .A2(new_n27277_), .B(new_n4295_), .ZN(new_n27279_));
  NOR2_X1    g27212(.A1(new_n26554_), .A2(new_n27279_), .ZN(new_n27280_));
  XOR2_X1    g27213(.A1(new_n27280_), .A2(new_n3372_), .Z(new_n27281_));
  NAND2_X1   g27214(.A1(new_n27013_), .A2(new_n27018_), .ZN(new_n27282_));
  INV_X1     g27215(.I(new_n27159_), .ZN(new_n27283_));
  XOR2_X1    g27216(.A1(new_n27091_), .A2(new_n27153_), .Z(new_n27284_));
  NOR2_X1    g27217(.A1(new_n27284_), .A2(new_n27283_), .ZN(new_n27285_));
  INV_X1     g27218(.I(new_n27285_), .ZN(new_n27286_));
  NAND4_X1   g27219(.A1(new_n27164_), .A2(new_n27016_), .A3(new_n27282_), .A4(new_n27286_), .ZN(new_n27287_));
  XOR2_X1    g27220(.A1(new_n27287_), .A2(new_n27281_), .Z(new_n27288_));
  XOR2_X1    g27221(.A1(new_n27276_), .A2(new_n27288_), .Z(new_n27289_));
  XOR2_X1    g27222(.A1(new_n27079_), .A2(new_n27177_), .Z(new_n27290_));
  NOR2_X1    g27223(.A1(new_n27179_), .A2(new_n27290_), .ZN(new_n27291_));
  NAND2_X1   g27224(.A1(new_n27291_), .A2(new_n27289_), .ZN(new_n27292_));
  INV_X1     g27225(.I(new_n27292_), .ZN(new_n27293_));
  NOR2_X1    g27226(.A1(new_n27291_), .A2(new_n27289_), .ZN(new_n27294_));
  NOR4_X1    g27227(.A1(new_n27293_), .A2(new_n27079_), .A3(new_n27294_), .A4(new_n27176_), .ZN(new_n27295_));
  INV_X1     g27228(.I(new_n27294_), .ZN(new_n27296_));
  AOI22_X1   g27229(.A1(new_n27296_), .A2(new_n27292_), .B1(new_n27080_), .B2(new_n27177_), .ZN(new_n27297_));
  NOR2_X1    g27230(.A1(new_n27297_), .A2(new_n27295_), .ZN(new_n27298_));
  XOR2_X1    g27231(.A1(new_n27192_), .A2(new_n27077_), .Z(new_n27299_));
  NAND3_X1   g27232(.A1(new_n27299_), .A2(new_n27183_), .A3(new_n27298_), .ZN(new_n27300_));
  AOI21_X1   g27233(.A1(new_n27299_), .A2(new_n27183_), .B(new_n27298_), .ZN(new_n27301_));
  INV_X1     g27234(.I(new_n27301_), .ZN(new_n27302_));
  NAND2_X1   g27235(.A1(new_n27192_), .A2(new_n27077_), .ZN(new_n27303_));
  INV_X1     g27236(.I(new_n27303_), .ZN(new_n27304_));
  NAND3_X1   g27237(.A1(new_n27302_), .A2(new_n27300_), .A3(new_n27304_), .ZN(new_n27305_));
  INV_X1     g27238(.I(new_n27300_), .ZN(new_n27306_));
  OAI21_X1   g27239(.A1(new_n27306_), .A2(new_n27301_), .B(new_n27303_), .ZN(new_n27307_));
  NAND2_X1   g27240(.A1(new_n27305_), .A2(new_n27307_), .ZN(new_n27308_));
  INV_X1     g27241(.I(new_n27308_), .ZN(new_n27309_));
  XOR2_X1    g27242(.A1(new_n27194_), .A2(new_n27309_), .Z(\result[20] ));
  XOR2_X1    g27243(.A1(new_n27276_), .A2(new_n27281_), .Z(new_n27311_));
  NAND2_X1   g27244(.A1(new_n27276_), .A2(new_n27281_), .ZN(new_n27312_));
  OAI21_X1   g27245(.A1(new_n27311_), .A2(new_n27287_), .B(new_n27312_), .ZN(new_n27313_));
  INV_X1     g27246(.I(new_n27313_), .ZN(new_n27314_));
  AOI21_X1   g27247(.A1(new_n27197_), .A2(new_n27240_), .B(new_n27241_), .ZN(new_n27315_));
  INV_X1     g27248(.I(new_n27315_), .ZN(new_n27316_));
  OAI21_X1   g27249(.A1(new_n27104_), .A2(new_n27198_), .B(new_n27214_), .ZN(new_n27317_));
  NAND2_X1   g27250(.A1(new_n27317_), .A2(new_n27212_), .ZN(new_n27318_));
  INV_X1     g27251(.I(new_n2581_), .ZN(new_n27319_));
  NAND4_X1   g27252(.A1(new_n382_), .A2(new_n1759_), .A3(new_n432_), .A4(new_n871_), .ZN(new_n27320_));
  NOR3_X1    g27253(.A1(new_n1245_), .A2(new_n98_), .A3(new_n782_), .ZN(new_n27321_));
  NAND4_X1   g27254(.A1(new_n27321_), .A2(new_n706_), .A3(new_n924_), .A4(new_n27320_), .ZN(new_n27322_));
  NOR2_X1    g27255(.A1(new_n200_), .A2(new_n1172_), .ZN(new_n27323_));
  NAND4_X1   g27256(.A1(new_n1742_), .A2(new_n27323_), .A3(new_n1576_), .A4(new_n2233_), .ZN(new_n27324_));
  NOR4_X1    g27257(.A1(new_n27322_), .A2(new_n27324_), .A3(new_n3212_), .A4(new_n27319_), .ZN(new_n27325_));
  NOR2_X1    g27258(.A1(new_n12024_), .A2(new_n3941_), .ZN(new_n27326_));
  NAND2_X1   g27259(.A1(new_n27326_), .A2(new_n27325_), .ZN(new_n27327_));
  INV_X1     g27260(.I(new_n27327_), .ZN(new_n27328_));
  NOR2_X1    g27261(.A1(new_n27328_), .A2(new_n27211_), .ZN(new_n27329_));
  NOR2_X1    g27262(.A1(new_n27327_), .A2(new_n27210_), .ZN(new_n27330_));
  NOR2_X1    g27263(.A1(new_n27329_), .A2(new_n27330_), .ZN(new_n27331_));
  INV_X1     g27264(.I(new_n27331_), .ZN(new_n27332_));
  XNOR2_X1   g27265(.A1(new_n27327_), .A2(new_n27210_), .ZN(new_n27333_));
  NOR2_X1    g27266(.A1(new_n27318_), .A2(new_n27333_), .ZN(new_n27334_));
  AOI21_X1   g27267(.A1(new_n27318_), .A2(new_n27332_), .B(new_n27334_), .ZN(new_n27335_));
  AOI22_X1   g27268(.A1(new_n17780_), .A2(new_n3275_), .B1(new_n19472_), .B2(new_n2746_), .ZN(new_n27336_));
  NOR2_X1    g27269(.A1(new_n17775_), .A2(new_n3175_), .ZN(new_n27337_));
  OAI21_X1   g27270(.A1(new_n27337_), .A2(new_n27336_), .B(new_n2736_), .ZN(new_n27338_));
  NOR2_X1    g27271(.A1(new_n21180_), .A2(new_n27338_), .ZN(new_n27339_));
  XOR2_X1    g27272(.A1(new_n27339_), .A2(new_n74_), .Z(new_n27340_));
  NOR2_X1    g27273(.A1(new_n19437_), .A2(new_n2772_), .ZN(new_n27341_));
  NOR2_X1    g27274(.A1(new_n17784_), .A2(new_n2767_), .ZN(new_n27342_));
  AOI21_X1   g27275(.A1(new_n20896_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n27343_));
  INV_X1     g27276(.I(new_n27343_), .ZN(new_n27344_));
  NOR4_X1    g27277(.A1(new_n21100_), .A2(new_n27341_), .A3(new_n27342_), .A4(new_n27344_), .ZN(new_n27345_));
  XOR2_X1    g27278(.A1(new_n27340_), .A2(new_n27345_), .Z(new_n27346_));
  NOR2_X1    g27279(.A1(new_n27346_), .A2(new_n27335_), .ZN(new_n27347_));
  INV_X1     g27280(.I(new_n27335_), .ZN(new_n27348_));
  INV_X1     g27281(.I(new_n27345_), .ZN(new_n27349_));
  NAND2_X1   g27282(.A1(new_n27340_), .A2(new_n27349_), .ZN(new_n27350_));
  NOR2_X1    g27283(.A1(new_n27340_), .A2(new_n27349_), .ZN(new_n27351_));
  INV_X1     g27284(.I(new_n27351_), .ZN(new_n27352_));
  AOI21_X1   g27285(.A1(new_n27352_), .A2(new_n27350_), .B(new_n27348_), .ZN(new_n27353_));
  NOR2_X1    g27286(.A1(new_n27347_), .A2(new_n27353_), .ZN(new_n27354_));
  OAI21_X1   g27287(.A1(new_n27218_), .A2(new_n27229_), .B(new_n27231_), .ZN(new_n27355_));
  OAI22_X1   g27288(.A1(new_n19512_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n19522_), .ZN(new_n27356_));
  NAND2_X1   g27289(.A1(new_n21953_), .A2(new_n3317_), .ZN(new_n27357_));
  AOI21_X1   g27290(.A1(new_n27356_), .A2(new_n27357_), .B(new_n3260_), .ZN(new_n27358_));
  NAND2_X1   g27291(.A1(new_n21963_), .A2(new_n27358_), .ZN(new_n27359_));
  XOR2_X1    g27292(.A1(new_n27359_), .A2(\a[26] ), .Z(new_n27360_));
  XOR2_X1    g27293(.A1(new_n27360_), .A2(new_n27355_), .Z(new_n27361_));
  NOR2_X1    g27294(.A1(new_n27361_), .A2(new_n27354_), .ZN(new_n27362_));
  INV_X1     g27295(.I(new_n27354_), .ZN(new_n27363_));
  INV_X1     g27296(.I(new_n27360_), .ZN(new_n27364_));
  NOR2_X1    g27297(.A1(new_n27364_), .A2(new_n27355_), .ZN(new_n27365_));
  INV_X1     g27298(.I(new_n27365_), .ZN(new_n27366_));
  NAND2_X1   g27299(.A1(new_n27364_), .A2(new_n27355_), .ZN(new_n27367_));
  AOI21_X1   g27300(.A1(new_n27366_), .A2(new_n27367_), .B(new_n27363_), .ZN(new_n27368_));
  NOR2_X1    g27301(.A1(new_n27368_), .A2(new_n27362_), .ZN(new_n27369_));
  OAI22_X1   g27302(.A1(new_n22115_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n22051_), .ZN(new_n27370_));
  NAND2_X1   g27303(.A1(new_n22150_), .A2(new_n3312_), .ZN(new_n27371_));
  AOI21_X1   g27304(.A1(new_n27370_), .A2(new_n27371_), .B(new_n3302_), .ZN(new_n27372_));
  NAND2_X1   g27305(.A1(new_n22163_), .A2(new_n27372_), .ZN(new_n27373_));
  XOR2_X1    g27306(.A1(new_n27373_), .A2(\a[23] ), .Z(new_n27374_));
  XOR2_X1    g27307(.A1(new_n27369_), .A2(new_n27374_), .Z(new_n27375_));
  INV_X1     g27308(.I(new_n27375_), .ZN(new_n27376_));
  XNOR2_X1   g27309(.A1(new_n27369_), .A2(new_n27374_), .ZN(new_n27377_));
  NOR2_X1    g27310(.A1(new_n27377_), .A2(new_n27316_), .ZN(new_n27378_));
  AOI21_X1   g27311(.A1(new_n27316_), .A2(new_n27376_), .B(new_n27378_), .ZN(new_n27379_));
  OAI21_X1   g27312(.A1(new_n27247_), .A2(new_n27256_), .B(new_n27258_), .ZN(new_n27380_));
  AOI22_X1   g27313(.A1(new_n24174_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n23957_), .ZN(new_n27381_));
  NOR2_X1    g27314(.A1(new_n24376_), .A2(new_n4097_), .ZN(new_n27382_));
  OAI21_X1   g27315(.A1(new_n27382_), .A2(new_n27381_), .B(new_n3773_), .ZN(new_n27383_));
  NOR3_X1    g27316(.A1(new_n24391_), .A2(\a[20] ), .A3(new_n27383_), .ZN(new_n27384_));
  NOR2_X1    g27317(.A1(new_n24391_), .A2(new_n27383_), .ZN(new_n27385_));
  NOR2_X1    g27318(.A1(new_n27385_), .A2(new_n3035_), .ZN(new_n27386_));
  NOR3_X1    g27319(.A1(new_n27380_), .A2(new_n27384_), .A3(new_n27386_), .ZN(new_n27387_));
  INV_X1     g27320(.I(new_n27380_), .ZN(new_n27388_));
  NOR2_X1    g27321(.A1(new_n27386_), .A2(new_n27384_), .ZN(new_n27389_));
  NOR2_X1    g27322(.A1(new_n27388_), .A2(new_n27389_), .ZN(new_n27390_));
  NOR2_X1    g27323(.A1(new_n27390_), .A2(new_n27387_), .ZN(new_n27391_));
  NOR2_X1    g27324(.A1(new_n27391_), .A2(new_n27379_), .ZN(new_n27392_));
  INV_X1     g27325(.I(new_n27379_), .ZN(new_n27393_));
  XOR2_X1    g27326(.A1(new_n27380_), .A2(new_n27389_), .Z(new_n27394_));
  NOR2_X1    g27327(.A1(new_n27394_), .A2(new_n27393_), .ZN(new_n27395_));
  NOR2_X1    g27328(.A1(new_n27392_), .A2(new_n27395_), .ZN(new_n27396_));
  OAI21_X1   g27329(.A1(new_n27262_), .A2(new_n27271_), .B(new_n27272_), .ZN(new_n27397_));
  AOI22_X1   g27330(.A1(new_n24826_), .A2(new_n11567_), .B1(new_n4292_), .B2(new_n24620_), .ZN(new_n27398_));
  OR3_X2     g27331(.A1(new_n25017_), .A2(new_n4468_), .A3(new_n27398_), .Z(new_n27399_));
  XOR2_X1    g27332(.A1(new_n27399_), .A2(\a[17] ), .Z(new_n27400_));
  INV_X1     g27333(.I(new_n27400_), .ZN(new_n27401_));
  NOR2_X1    g27334(.A1(new_n27397_), .A2(new_n27401_), .ZN(new_n27402_));
  INV_X1     g27335(.I(new_n27402_), .ZN(new_n27403_));
  NAND2_X1   g27336(.A1(new_n27397_), .A2(new_n27401_), .ZN(new_n27404_));
  AOI21_X1   g27337(.A1(new_n27403_), .A2(new_n27404_), .B(new_n27396_), .ZN(new_n27405_));
  XOR2_X1    g27338(.A1(new_n27397_), .A2(new_n27400_), .Z(new_n27406_));
  NOR3_X1    g27339(.A1(new_n27406_), .A2(new_n27392_), .A3(new_n27395_), .ZN(new_n27407_));
  NOR2_X1    g27340(.A1(new_n27407_), .A2(new_n27405_), .ZN(new_n27408_));
  INV_X1     g27341(.I(new_n27408_), .ZN(new_n27409_));
  NOR2_X1    g27342(.A1(new_n27183_), .A2(new_n27077_), .ZN(new_n27410_));
  INV_X1     g27343(.I(new_n27410_), .ZN(new_n27411_));
  NOR3_X1    g27344(.A1(new_n27410_), .A2(new_n27295_), .A3(new_n27297_), .ZN(new_n27412_));
  OAI21_X1   g27345(.A1(new_n27192_), .A2(new_n27411_), .B(new_n27412_), .ZN(new_n27413_));
  NOR2_X1    g27346(.A1(new_n27180_), .A2(new_n27080_), .ZN(new_n27414_));
  INV_X1     g27347(.I(new_n27414_), .ZN(new_n27415_));
  AND3_X2    g27348(.A1(new_n27415_), .A2(new_n27180_), .A3(new_n27289_), .Z(new_n27416_));
  INV_X1     g27349(.I(new_n27416_), .ZN(new_n27417_));
  NOR2_X1    g27350(.A1(new_n27413_), .A2(new_n27417_), .ZN(new_n27418_));
  XOR2_X1    g27351(.A1(new_n27418_), .A2(new_n27409_), .Z(new_n27419_));
  XOR2_X1    g27352(.A1(new_n27419_), .A2(new_n27314_), .Z(new_n27420_));
  NOR2_X1    g27353(.A1(new_n27194_), .A2(new_n27309_), .ZN(new_n27421_));
  XOR2_X1    g27354(.A1(new_n27421_), .A2(new_n27420_), .Z(\result[21] ));
  NOR2_X1    g27355(.A1(new_n27314_), .A2(new_n27409_), .ZN(new_n27423_));
  INV_X1     g27356(.I(new_n27423_), .ZN(new_n27424_));
  XOR2_X1    g27357(.A1(new_n27313_), .A2(new_n27408_), .Z(new_n27425_));
  NOR2_X1    g27358(.A1(new_n27417_), .A2(new_n27425_), .ZN(new_n27426_));
  INV_X1     g27359(.I(new_n27426_), .ZN(new_n27427_));
  OAI21_X1   g27360(.A1(new_n27413_), .A2(new_n27427_), .B(new_n27424_), .ZN(new_n27428_));
  OAI21_X1   g27361(.A1(new_n27396_), .A2(new_n27402_), .B(new_n27404_), .ZN(new_n27429_));
  INV_X1     g27362(.I(new_n27429_), .ZN(new_n27430_));
  INV_X1     g27363(.I(new_n27387_), .ZN(new_n27431_));
  AOI21_X1   g27364(.A1(new_n27393_), .A2(new_n27431_), .B(new_n27390_), .ZN(new_n27432_));
  INV_X1     g27365(.I(new_n27432_), .ZN(new_n27433_));
  OAI21_X1   g27366(.A1(new_n27363_), .A2(new_n27365_), .B(new_n27367_), .ZN(new_n27434_));
  OAI22_X1   g27367(.A1(new_n19512_), .A2(new_n3268_), .B1(new_n21960_), .B2(new_n3322_), .ZN(new_n27435_));
  NAND2_X1   g27368(.A1(new_n22048_), .A2(new_n3317_), .ZN(new_n27436_));
  AOI21_X1   g27369(.A1(new_n27436_), .A2(new_n27435_), .B(new_n3260_), .ZN(new_n27437_));
  NAND2_X1   g27370(.A1(new_n22175_), .A2(new_n27437_), .ZN(new_n27438_));
  XOR2_X1    g27371(.A1(new_n27438_), .A2(\a[26] ), .Z(new_n27439_));
  INV_X1     g27372(.I(new_n27439_), .ZN(new_n27440_));
  NOR2_X1    g27373(.A1(new_n27434_), .A2(new_n27440_), .ZN(new_n27441_));
  NAND2_X1   g27374(.A1(new_n27434_), .A2(new_n27440_), .ZN(new_n27442_));
  INV_X1     g27375(.I(new_n27442_), .ZN(new_n27443_));
  NOR2_X1    g27376(.A1(new_n27443_), .A2(new_n27441_), .ZN(new_n27444_));
  NAND2_X1   g27377(.A1(new_n27350_), .A2(new_n27348_), .ZN(new_n27445_));
  NAND2_X1   g27378(.A1(new_n27445_), .A2(new_n27352_), .ZN(new_n27446_));
  INV_X1     g27379(.I(new_n27329_), .ZN(new_n27447_));
  OAI21_X1   g27380(.A1(new_n27210_), .A2(new_n27327_), .B(new_n27318_), .ZN(new_n27448_));
  NAND2_X1   g27381(.A1(new_n27448_), .A2(new_n27447_), .ZN(new_n27449_));
  INV_X1     g27382(.I(new_n27449_), .ZN(new_n27450_));
  NOR2_X1    g27383(.A1(new_n24835_), .A2(new_n11568_), .ZN(new_n27451_));
  OAI22_X1   g27384(.A1(new_n27451_), .A2(\a[17] ), .B1(new_n11570_), .B2(new_n24835_), .ZN(new_n27452_));
  NOR3_X1    g27385(.A1(new_n866_), .A2(new_n326_), .A3(new_n731_), .ZN(new_n27453_));
  NOR3_X1    g27386(.A1(new_n3213_), .A2(new_n76_), .A3(new_n125_), .ZN(new_n27454_));
  NAND4_X1   g27387(.A1(new_n1208_), .A2(new_n19973_), .A3(new_n27454_), .A4(new_n27453_), .ZN(new_n27455_));
  NAND2_X1   g27388(.A1(new_n2477_), .A2(new_n1785_), .ZN(new_n27456_));
  NOR4_X1    g27389(.A1(new_n916_), .A2(new_n10974_), .A3(new_n27456_), .A4(new_n27455_), .ZN(new_n27457_));
  NOR2_X1    g27390(.A1(new_n8323_), .A2(new_n3683_), .ZN(new_n27458_));
  NAND2_X1   g27391(.A1(new_n27458_), .A2(new_n27457_), .ZN(new_n27459_));
  NAND2_X1   g27392(.A1(new_n27459_), .A2(new_n27327_), .ZN(new_n27460_));
  INV_X1     g27393(.I(new_n27460_), .ZN(new_n27461_));
  NOR2_X1    g27394(.A1(new_n27459_), .A2(new_n27327_), .ZN(new_n27462_));
  OAI21_X1   g27395(.A1(new_n27461_), .A2(new_n27462_), .B(new_n27452_), .ZN(new_n27463_));
  XOR2_X1    g27396(.A1(new_n27459_), .A2(new_n27328_), .Z(new_n27464_));
  OAI21_X1   g27397(.A1(new_n27452_), .A2(new_n27464_), .B(new_n27463_), .ZN(new_n27465_));
  NAND2_X1   g27398(.A1(new_n19472_), .A2(new_n3332_), .ZN(new_n27466_));
  NAND2_X1   g27399(.A1(new_n19466_), .A2(new_n3189_), .ZN(new_n27467_));
  AOI21_X1   g27400(.A1(new_n19438_), .A2(new_n2770_), .B(new_n2763_), .ZN(new_n27468_));
  NAND4_X1   g27401(.A1(new_n21117_), .A2(new_n27466_), .A3(new_n27467_), .A4(new_n27468_), .ZN(new_n27469_));
  NAND2_X1   g27402(.A1(new_n27469_), .A2(new_n27465_), .ZN(new_n27470_));
  NOR2_X1    g27403(.A1(new_n27469_), .A2(new_n27465_), .ZN(new_n27471_));
  INV_X1     g27404(.I(new_n27471_), .ZN(new_n27472_));
  AOI21_X1   g27405(.A1(new_n27470_), .A2(new_n27472_), .B(new_n27450_), .ZN(new_n27473_));
  XOR2_X1    g27406(.A1(new_n27469_), .A2(new_n27465_), .Z(new_n27474_));
  AOI21_X1   g27407(.A1(new_n27450_), .A2(new_n27474_), .B(new_n27473_), .ZN(new_n27475_));
  XOR2_X1    g27408(.A1(new_n27475_), .A2(new_n27446_), .Z(new_n27476_));
  OAI22_X1   g27409(.A1(new_n17775_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19475_), .ZN(new_n27477_));
  NAND2_X1   g27410(.A1(new_n21157_), .A2(new_n2750_), .ZN(new_n27478_));
  AOI21_X1   g27411(.A1(new_n27478_), .A2(new_n27477_), .B(new_n2737_), .ZN(new_n27479_));
  NAND2_X1   g27412(.A1(new_n21155_), .A2(new_n27479_), .ZN(new_n27480_));
  XOR2_X1    g27413(.A1(new_n27480_), .A2(\a[29] ), .Z(new_n27481_));
  INV_X1     g27414(.I(new_n27481_), .ZN(new_n27482_));
  XOR2_X1    g27415(.A1(new_n27476_), .A2(new_n27482_), .Z(new_n27483_));
  OAI22_X1   g27416(.A1(new_n22115_), .A2(new_n3310_), .B1(new_n3306_), .B2(new_n22149_), .ZN(new_n27484_));
  NAND2_X1   g27417(.A1(new_n23957_), .A2(new_n3312_), .ZN(new_n27485_));
  AOI21_X1   g27418(.A1(new_n27484_), .A2(new_n27485_), .B(new_n3302_), .ZN(new_n27486_));
  NAND2_X1   g27419(.A1(new_n23955_), .A2(new_n27486_), .ZN(new_n27487_));
  XOR2_X1    g27420(.A1(new_n27487_), .A2(\a[23] ), .Z(new_n27488_));
  XOR2_X1    g27421(.A1(new_n27488_), .A2(new_n27483_), .Z(new_n27489_));
  INV_X1     g27422(.I(new_n27489_), .ZN(new_n27490_));
  INV_X1     g27423(.I(new_n27483_), .ZN(new_n27491_));
  XOR2_X1    g27424(.A1(new_n27488_), .A2(new_n27491_), .Z(new_n27492_));
  NAND2_X1   g27425(.A1(new_n27492_), .A2(new_n27444_), .ZN(new_n27493_));
  OAI21_X1   g27426(.A1(new_n27444_), .A2(new_n27490_), .B(new_n27493_), .ZN(new_n27494_));
  NOR2_X1    g27427(.A1(new_n27369_), .A2(new_n27315_), .ZN(new_n27495_));
  INV_X1     g27428(.I(new_n27495_), .ZN(new_n27496_));
  XOR2_X1    g27429(.A1(new_n27494_), .A2(new_n27496_), .Z(new_n27497_));
  XOR2_X1    g27430(.A1(new_n27369_), .A2(new_n27316_), .Z(new_n27498_));
  NOR2_X1    g27431(.A1(new_n27498_), .A2(new_n27374_), .ZN(new_n27499_));
  XOR2_X1    g27432(.A1(new_n27497_), .A2(new_n27499_), .Z(new_n27500_));
  OAI22_X1   g27433(.A1(new_n24376_), .A2(new_n3775_), .B1(new_n3769_), .B2(new_n24167_), .ZN(new_n27501_));
  NAND2_X1   g27434(.A1(new_n24620_), .A2(new_n4096_), .ZN(new_n27502_));
  AOI21_X1   g27435(.A1(new_n27502_), .A2(new_n27501_), .B(new_n4095_), .ZN(new_n27503_));
  NAND2_X1   g27436(.A1(new_n24618_), .A2(new_n27503_), .ZN(new_n27504_));
  XOR2_X1    g27437(.A1(new_n27504_), .A2(\a[20] ), .Z(new_n27505_));
  INV_X1     g27438(.I(new_n27505_), .ZN(new_n27506_));
  XOR2_X1    g27439(.A1(new_n27500_), .A2(new_n27506_), .Z(new_n27507_));
  NOR2_X1    g27440(.A1(new_n27500_), .A2(new_n27506_), .ZN(new_n27508_));
  INV_X1     g27441(.I(new_n27508_), .ZN(new_n27509_));
  NAND2_X1   g27442(.A1(new_n27500_), .A2(new_n27506_), .ZN(new_n27510_));
  AOI21_X1   g27443(.A1(new_n27509_), .A2(new_n27510_), .B(new_n27433_), .ZN(new_n27511_));
  AOI21_X1   g27444(.A1(new_n27433_), .A2(new_n27507_), .B(new_n27511_), .ZN(new_n27512_));
  XOR2_X1    g27445(.A1(new_n27512_), .A2(new_n27430_), .Z(new_n27513_));
  NAND4_X1   g27446(.A1(new_n27185_), .A2(new_n27193_), .A3(new_n27420_), .A4(new_n27308_), .ZN(new_n27514_));
  XOR2_X1    g27447(.A1(new_n27514_), .A2(new_n27513_), .Z(new_n27515_));
  XOR2_X1    g27448(.A1(new_n27515_), .A2(new_n27428_), .Z(\result[22] ));
  XOR2_X1    g27449(.A1(new_n27419_), .A2(new_n27313_), .Z(new_n27517_));
  XOR2_X1    g27450(.A1(new_n27428_), .A2(new_n27513_), .Z(new_n27518_));
  INV_X1     g27451(.I(new_n27518_), .ZN(new_n27519_));
  NOR4_X1    g27452(.A1(new_n27194_), .A2(new_n27309_), .A3(new_n27517_), .A4(new_n27519_), .ZN(new_n27520_));
  AOI21_X1   g27453(.A1(new_n27449_), .A2(new_n27470_), .B(new_n27471_), .ZN(new_n27521_));
  INV_X1     g27454(.I(new_n27452_), .ZN(new_n27522_));
  AOI21_X1   g27455(.A1(new_n27522_), .A2(new_n27460_), .B(new_n27462_), .ZN(new_n27523_));
  INV_X1     g27456(.I(new_n27523_), .ZN(new_n27524_));
  NOR2_X1    g27457(.A1(new_n19475_), .A2(new_n2772_), .ZN(new_n27525_));
  NOR2_X1    g27458(.A1(new_n19463_), .A2(new_n2767_), .ZN(new_n27526_));
  OAI21_X1   g27459(.A1(new_n19437_), .A2(new_n2771_), .B(new_n2763_), .ZN(new_n27527_));
  OR4_X2     g27460(.A1(new_n21088_), .A2(new_n27525_), .A3(new_n27526_), .A4(new_n27527_), .Z(new_n27528_));
  INV_X1     g27461(.I(new_n6539_), .ZN(new_n27529_));
  NOR2_X1    g27462(.A1(new_n939_), .A2(new_n114_), .ZN(new_n27530_));
  NAND3_X1   g27463(.A1(new_n1495_), .A2(new_n356_), .A3(new_n842_), .ZN(new_n27531_));
  NOR4_X1    g27464(.A1(new_n906_), .A2(new_n198_), .A3(new_n136_), .A4(new_n776_), .ZN(new_n27532_));
  NOR4_X1    g27465(.A1(new_n27531_), .A2(new_n314_), .A3(new_n1932_), .A4(new_n27532_), .ZN(new_n27533_));
  NAND3_X1   g27466(.A1(new_n27533_), .A2(new_n3365_), .A3(new_n27530_), .ZN(new_n27534_));
  NOR4_X1    g27467(.A1(new_n27529_), .A2(new_n1874_), .A3(new_n2519_), .A4(new_n27534_), .ZN(new_n27535_));
  NAND2_X1   g27468(.A1(new_n27535_), .A2(new_n26143_), .ZN(new_n27536_));
  INV_X1     g27469(.I(new_n27536_), .ZN(new_n27537_));
  NOR2_X1    g27470(.A1(new_n27528_), .A2(new_n27537_), .ZN(new_n27538_));
  NAND2_X1   g27471(.A1(new_n27528_), .A2(new_n27537_), .ZN(new_n27539_));
  INV_X1     g27472(.I(new_n27539_), .ZN(new_n27540_));
  OAI21_X1   g27473(.A1(new_n27540_), .A2(new_n27538_), .B(new_n27524_), .ZN(new_n27541_));
  XOR2_X1    g27474(.A1(new_n27528_), .A2(new_n27536_), .Z(new_n27542_));
  OAI21_X1   g27475(.A1(new_n27524_), .A2(new_n27542_), .B(new_n27541_), .ZN(new_n27543_));
  AOI22_X1   g27476(.A1(new_n21157_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n19484_), .ZN(new_n27544_));
  NOR2_X1    g27477(.A1(new_n19512_), .A2(new_n3175_), .ZN(new_n27545_));
  OAI21_X1   g27478(.A1(new_n27545_), .A2(new_n27544_), .B(new_n2736_), .ZN(new_n27546_));
  NOR3_X1    g27479(.A1(new_n25926_), .A2(\a[29] ), .A3(new_n27546_), .ZN(new_n27547_));
  NOR2_X1    g27480(.A1(new_n25926_), .A2(new_n27546_), .ZN(new_n27548_));
  NOR2_X1    g27481(.A1(new_n27548_), .A2(new_n74_), .ZN(new_n27549_));
  NOR2_X1    g27482(.A1(new_n27549_), .A2(new_n27547_), .ZN(new_n27550_));
  XOR2_X1    g27483(.A1(new_n27543_), .A2(new_n27550_), .Z(new_n27551_));
  NOR2_X1    g27484(.A1(new_n27551_), .A2(new_n27521_), .ZN(new_n27552_));
  INV_X1     g27485(.I(new_n27550_), .ZN(new_n27553_));
  NOR2_X1    g27486(.A1(new_n27553_), .A2(new_n27543_), .ZN(new_n27554_));
  INV_X1     g27487(.I(new_n27554_), .ZN(new_n27555_));
  NAND2_X1   g27488(.A1(new_n27553_), .A2(new_n27543_), .ZN(new_n27556_));
  NAND2_X1   g27489(.A1(new_n27555_), .A2(new_n27556_), .ZN(new_n27557_));
  AOI21_X1   g27490(.A1(new_n27521_), .A2(new_n27557_), .B(new_n27552_), .ZN(new_n27558_));
  AOI22_X1   g27491(.A1(new_n22048_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n21953_), .ZN(new_n27559_));
  NOR2_X1    g27492(.A1(new_n22115_), .A2(new_n3318_), .ZN(new_n27560_));
  OAI21_X1   g27493(.A1(new_n27560_), .A2(new_n27559_), .B(new_n3259_), .ZN(new_n27561_));
  NOR2_X1    g27494(.A1(new_n23675_), .A2(new_n27561_), .ZN(new_n27562_));
  XOR2_X1    g27495(.A1(new_n27562_), .A2(\a[26] ), .Z(new_n27563_));
  INV_X1     g27496(.I(new_n27475_), .ZN(new_n27564_));
  NOR2_X1    g27497(.A1(new_n27564_), .A2(new_n27446_), .ZN(new_n27565_));
  NOR2_X1    g27498(.A1(new_n27476_), .A2(new_n27482_), .ZN(new_n27566_));
  NOR2_X1    g27499(.A1(new_n27566_), .A2(new_n27565_), .ZN(new_n27567_));
  XOR2_X1    g27500(.A1(new_n27567_), .A2(new_n27563_), .Z(new_n27568_));
  XNOR2_X1   g27501(.A1(new_n27568_), .A2(new_n27558_), .ZN(new_n27569_));
  INV_X1     g27502(.I(new_n27569_), .ZN(new_n27570_));
  OAI21_X1   g27503(.A1(new_n27483_), .A2(new_n27441_), .B(new_n27442_), .ZN(new_n27571_));
  OAI22_X1   g27504(.A1(new_n23948_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n22149_), .ZN(new_n27572_));
  NAND2_X1   g27505(.A1(new_n24174_), .A2(new_n3312_), .ZN(new_n27573_));
  AOI21_X1   g27506(.A1(new_n27573_), .A2(new_n27572_), .B(new_n3302_), .ZN(new_n27574_));
  NAND2_X1   g27507(.A1(new_n24172_), .A2(new_n27574_), .ZN(new_n27575_));
  XOR2_X1    g27508(.A1(new_n27575_), .A2(\a[23] ), .Z(new_n27576_));
  INV_X1     g27509(.I(new_n27576_), .ZN(new_n27577_));
  NOR2_X1    g27510(.A1(new_n27577_), .A2(new_n27571_), .ZN(new_n27578_));
  NAND2_X1   g27511(.A1(new_n27577_), .A2(new_n27571_), .ZN(new_n27579_));
  INV_X1     g27512(.I(new_n27579_), .ZN(new_n27580_));
  OAI21_X1   g27513(.A1(new_n27578_), .A2(new_n27580_), .B(new_n27570_), .ZN(new_n27581_));
  XOR2_X1    g27514(.A1(new_n27576_), .A2(new_n27571_), .Z(new_n27582_));
  OAI21_X1   g27515(.A1(new_n27570_), .A2(new_n27582_), .B(new_n27581_), .ZN(new_n27583_));
  AOI22_X1   g27516(.A1(new_n24620_), .A2(new_n3776_), .B1(new_n3770_), .B2(new_n24386_), .ZN(new_n27584_));
  NOR2_X1    g27517(.A1(new_n24835_), .A2(new_n4097_), .ZN(new_n27585_));
  OAI21_X1   g27518(.A1(new_n27585_), .A2(new_n27584_), .B(new_n3773_), .ZN(new_n27586_));
  NOR2_X1    g27519(.A1(new_n26554_), .A2(new_n27586_), .ZN(new_n27587_));
  XOR2_X1    g27520(.A1(new_n27587_), .A2(new_n3035_), .Z(new_n27588_));
  INV_X1     g27521(.I(new_n27588_), .ZN(new_n27589_));
  INV_X1     g27522(.I(new_n27488_), .ZN(new_n27590_));
  NOR3_X1    g27523(.A1(new_n27316_), .A2(new_n27362_), .A3(new_n27368_), .ZN(new_n27591_));
  NOR3_X1    g27524(.A1(new_n27494_), .A2(new_n27374_), .A3(new_n27591_), .ZN(new_n27592_));
  XOR2_X1    g27525(.A1(new_n27444_), .A2(new_n27491_), .Z(new_n27593_));
  OAI22_X1   g27526(.A1(new_n27592_), .A2(new_n27496_), .B1(new_n27590_), .B2(new_n27593_), .ZN(new_n27594_));
  XOR2_X1    g27527(.A1(new_n27594_), .A2(new_n27589_), .Z(new_n27595_));
  XOR2_X1    g27528(.A1(new_n27595_), .A2(new_n27583_), .Z(new_n27596_));
  XOR2_X1    g27529(.A1(new_n27432_), .A2(new_n27505_), .Z(new_n27597_));
  NAND2_X1   g27530(.A1(new_n27500_), .A2(new_n27597_), .ZN(new_n27598_));
  XOR2_X1    g27531(.A1(new_n27596_), .A2(new_n27598_), .Z(new_n27599_));
  NAND2_X1   g27532(.A1(new_n27433_), .A2(new_n27506_), .ZN(new_n27600_));
  XOR2_X1    g27533(.A1(new_n27599_), .A2(new_n27600_), .Z(new_n27601_));
  INV_X1     g27534(.I(new_n27601_), .ZN(new_n27602_));
  XOR2_X1    g27535(.A1(new_n27428_), .A2(new_n27429_), .Z(new_n27603_));
  NAND3_X1   g27536(.A1(new_n27603_), .A2(new_n27512_), .A3(new_n27602_), .ZN(new_n27604_));
  NOR2_X1    g27537(.A1(new_n27428_), .A2(new_n27430_), .ZN(new_n27605_));
  INV_X1     g27538(.I(new_n27412_), .ZN(new_n27606_));
  AOI21_X1   g27539(.A1(new_n27075_), .A2(new_n27410_), .B(new_n27606_), .ZN(new_n27607_));
  AOI21_X1   g27540(.A1(new_n27607_), .A2(new_n27426_), .B(new_n27423_), .ZN(new_n27608_));
  NOR2_X1    g27541(.A1(new_n27608_), .A2(new_n27429_), .ZN(new_n27609_));
  OAI21_X1   g27542(.A1(new_n27609_), .A2(new_n27605_), .B(new_n27512_), .ZN(new_n27610_));
  NAND2_X1   g27543(.A1(new_n27610_), .A2(new_n27601_), .ZN(new_n27611_));
  NOR2_X1    g27544(.A1(new_n27608_), .A2(new_n27430_), .ZN(new_n27612_));
  NAND3_X1   g27545(.A1(new_n27604_), .A2(new_n27611_), .A3(new_n27612_), .ZN(new_n27613_));
  NOR2_X1    g27546(.A1(new_n27610_), .A2(new_n27601_), .ZN(new_n27614_));
  AOI21_X1   g27547(.A1(new_n27603_), .A2(new_n27512_), .B(new_n27602_), .ZN(new_n27615_));
  INV_X1     g27548(.I(new_n27612_), .ZN(new_n27616_));
  OAI21_X1   g27549(.A1(new_n27615_), .A2(new_n27614_), .B(new_n27616_), .ZN(new_n27617_));
  NAND2_X1   g27550(.A1(new_n27617_), .A2(new_n27613_), .ZN(new_n27618_));
  XOR2_X1    g27551(.A1(new_n27520_), .A2(new_n27618_), .Z(\result[23] ));
  NAND2_X1   g27552(.A1(new_n27520_), .A2(new_n27618_), .ZN(new_n27620_));
  OAI21_X1   g27553(.A1(new_n27521_), .A2(new_n27554_), .B(new_n27556_), .ZN(new_n27621_));
  NOR2_X1    g27554(.A1(new_n27540_), .A2(new_n27523_), .ZN(new_n27622_));
  NOR2_X1    g27555(.A1(new_n27622_), .A2(new_n27538_), .ZN(new_n27623_));
  NOR2_X1    g27556(.A1(new_n17775_), .A2(new_n2772_), .ZN(new_n27624_));
  NOR2_X1    g27557(.A1(new_n19475_), .A2(new_n2767_), .ZN(new_n27625_));
  NOR2_X1    g27558(.A1(new_n19463_), .A2(new_n2771_), .ZN(new_n27626_));
  NOR4_X1    g27559(.A1(new_n27624_), .A2(new_n2764_), .A3(new_n27625_), .A4(new_n27626_), .ZN(new_n27627_));
  NAND2_X1   g27560(.A1(new_n21180_), .A2(new_n27627_), .ZN(new_n27628_));
  NAND4_X1   g27561(.A1(new_n868_), .A2(new_n1662_), .A3(new_n773_), .A4(new_n1856_), .ZN(new_n27629_));
  NOR4_X1    g27562(.A1(new_n1138_), .A2(new_n333_), .A3(new_n1167_), .A4(new_n518_), .ZN(new_n27630_));
  NAND2_X1   g27563(.A1(new_n27321_), .A2(new_n10987_), .ZN(new_n27631_));
  INV_X1     g27564(.I(new_n25323_), .ZN(new_n27632_));
  NAND2_X1   g27565(.A1(new_n27632_), .A2(new_n8320_), .ZN(new_n27633_));
  NOR4_X1    g27566(.A1(new_n27633_), .A2(new_n27629_), .A3(new_n27631_), .A4(new_n27630_), .ZN(new_n27634_));
  NAND4_X1   g27567(.A1(new_n4943_), .A2(new_n942_), .A3(new_n3464_), .A4(new_n27634_), .ZN(new_n27635_));
  NAND2_X1   g27568(.A1(new_n27537_), .A2(new_n27635_), .ZN(new_n27636_));
  OR2_X2     g27569(.A1(new_n27537_), .A2(new_n27635_), .Z(new_n27637_));
  AOI21_X1   g27570(.A1(new_n27636_), .A2(new_n27637_), .B(new_n27628_), .ZN(new_n27638_));
  INV_X1     g27571(.I(new_n27628_), .ZN(new_n27639_));
  XOR2_X1    g27572(.A1(new_n27536_), .A2(new_n27635_), .Z(new_n27640_));
  NOR2_X1    g27573(.A1(new_n27639_), .A2(new_n27640_), .ZN(new_n27641_));
  NOR2_X1    g27574(.A1(new_n27641_), .A2(new_n27638_), .ZN(new_n27642_));
  XOR2_X1    g27575(.A1(new_n27623_), .A2(new_n27642_), .Z(new_n27643_));
  NAND2_X1   g27576(.A1(new_n27621_), .A2(new_n27643_), .ZN(new_n27644_));
  NOR4_X1    g27577(.A1(new_n27622_), .A2(new_n27538_), .A3(new_n27638_), .A4(new_n27641_), .ZN(new_n27645_));
  NOR2_X1    g27578(.A1(new_n27623_), .A2(new_n27642_), .ZN(new_n27646_));
  NOR2_X1    g27579(.A1(new_n27646_), .A2(new_n27645_), .ZN(new_n27647_));
  OAI21_X1   g27580(.A1(new_n27621_), .A2(new_n27647_), .B(new_n27644_), .ZN(new_n27648_));
  OAI22_X1   g27581(.A1(new_n22115_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n22051_), .ZN(new_n27649_));
  NAND2_X1   g27582(.A1(new_n22150_), .A2(new_n3317_), .ZN(new_n27650_));
  AOI21_X1   g27583(.A1(new_n27649_), .A2(new_n27650_), .B(new_n3260_), .ZN(new_n27651_));
  NAND2_X1   g27584(.A1(new_n22163_), .A2(new_n27651_), .ZN(new_n27652_));
  XOR2_X1    g27585(.A1(new_n27652_), .A2(\a[26] ), .Z(new_n27653_));
  OAI22_X1   g27586(.A1(new_n19512_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n19522_), .ZN(new_n27654_));
  NAND2_X1   g27587(.A1(new_n21953_), .A2(new_n2750_), .ZN(new_n27655_));
  AOI21_X1   g27588(.A1(new_n27654_), .A2(new_n27655_), .B(new_n2737_), .ZN(new_n27656_));
  NAND2_X1   g27589(.A1(new_n21963_), .A2(new_n27656_), .ZN(new_n27657_));
  XOR2_X1    g27590(.A1(new_n27657_), .A2(\a[29] ), .Z(new_n27658_));
  XOR2_X1    g27591(.A1(new_n27653_), .A2(new_n27658_), .Z(new_n27659_));
  NAND2_X1   g27592(.A1(new_n27659_), .A2(new_n27648_), .ZN(new_n27660_));
  AND2_X2    g27593(.A1(new_n27653_), .A2(new_n27658_), .Z(new_n27661_));
  NOR2_X1    g27594(.A1(new_n27653_), .A2(new_n27658_), .ZN(new_n27662_));
  NOR2_X1    g27595(.A1(new_n27661_), .A2(new_n27662_), .ZN(new_n27663_));
  OAI21_X1   g27596(.A1(new_n27648_), .A2(new_n27663_), .B(new_n27660_), .ZN(new_n27664_));
  AOI22_X1   g27597(.A1(new_n24174_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n23957_), .ZN(new_n27665_));
  NOR2_X1    g27598(.A1(new_n24376_), .A2(new_n3780_), .ZN(new_n27666_));
  OAI21_X1   g27599(.A1(new_n27666_), .A2(new_n27665_), .B(new_n3301_), .ZN(new_n27667_));
  NOR2_X1    g27600(.A1(new_n24391_), .A2(new_n27667_), .ZN(new_n27668_));
  XOR2_X1    g27601(.A1(new_n27668_), .A2(new_n84_), .Z(new_n27669_));
  XOR2_X1    g27602(.A1(new_n27664_), .A2(new_n27669_), .Z(new_n27670_));
  OAI21_X1   g27603(.A1(new_n27569_), .A2(new_n27578_), .B(new_n27579_), .ZN(new_n27671_));
  AOI22_X1   g27604(.A1(new_n24826_), .A2(new_n11227_), .B1(new_n3770_), .B2(new_n24620_), .ZN(new_n27672_));
  OR3_X2     g27605(.A1(new_n25017_), .A2(new_n4095_), .A3(new_n27672_), .Z(new_n27673_));
  XOR2_X1    g27606(.A1(new_n27673_), .A2(\a[20] ), .Z(new_n27674_));
  INV_X1     g27607(.I(new_n27674_), .ZN(new_n27675_));
  NOR2_X1    g27608(.A1(new_n27671_), .A2(new_n27675_), .ZN(new_n27676_));
  INV_X1     g27609(.I(new_n27676_), .ZN(new_n27677_));
  NAND2_X1   g27610(.A1(new_n27671_), .A2(new_n27675_), .ZN(new_n27678_));
  AOI21_X1   g27611(.A1(new_n27677_), .A2(new_n27678_), .B(new_n27670_), .ZN(new_n27679_));
  XOR2_X1    g27612(.A1(new_n27671_), .A2(new_n27674_), .Z(new_n27680_));
  INV_X1     g27613(.I(new_n27680_), .ZN(new_n27681_));
  AOI21_X1   g27614(.A1(new_n27681_), .A2(new_n27670_), .B(new_n27679_), .ZN(new_n27682_));
  INV_X1     g27615(.I(new_n27682_), .ZN(new_n27683_));
  XOR2_X1    g27616(.A1(new_n27583_), .A2(new_n27588_), .Z(new_n27684_));
  AOI21_X1   g27617(.A1(new_n27589_), .A2(new_n27594_), .B(new_n27684_), .ZN(new_n27685_));
  INV_X1     g27618(.I(new_n27685_), .ZN(new_n27686_));
  NOR2_X1    g27619(.A1(new_n27512_), .A2(new_n27429_), .ZN(new_n27687_));
  INV_X1     g27620(.I(new_n27687_), .ZN(new_n27688_));
  NOR2_X1    g27621(.A1(new_n27601_), .A2(new_n27687_), .ZN(new_n27689_));
  OAI21_X1   g27622(.A1(new_n27428_), .A2(new_n27688_), .B(new_n27689_), .ZN(new_n27690_));
  NOR2_X1    g27623(.A1(new_n27509_), .A2(new_n27433_), .ZN(new_n27691_));
  NOR3_X1    g27624(.A1(new_n27691_), .A2(new_n27596_), .A3(new_n27508_), .ZN(new_n27692_));
  INV_X1     g27625(.I(new_n27692_), .ZN(new_n27693_));
  NOR2_X1    g27626(.A1(new_n27690_), .A2(new_n27693_), .ZN(new_n27694_));
  INV_X1     g27627(.I(new_n27694_), .ZN(new_n27695_));
  NAND2_X1   g27628(.A1(new_n27695_), .A2(new_n27686_), .ZN(new_n27696_));
  NAND2_X1   g27629(.A1(new_n27694_), .A2(new_n27685_), .ZN(new_n27697_));
  AOI21_X1   g27630(.A1(new_n27696_), .A2(new_n27697_), .B(new_n27683_), .ZN(new_n27698_));
  NOR2_X1    g27631(.A1(new_n27694_), .A2(new_n27685_), .ZN(new_n27699_));
  INV_X1     g27632(.I(new_n27697_), .ZN(new_n27700_));
  NOR3_X1    g27633(.A1(new_n27700_), .A2(new_n27682_), .A3(new_n27699_), .ZN(new_n27701_));
  NOR2_X1    g27634(.A1(new_n27701_), .A2(new_n27698_), .ZN(new_n27702_));
  XOR2_X1    g27635(.A1(new_n27620_), .A2(new_n27702_), .Z(\result[24] ));
  NOR2_X1    g27636(.A1(new_n27685_), .A2(new_n27682_), .ZN(new_n27704_));
  INV_X1     g27637(.I(new_n27704_), .ZN(new_n27705_));
  XOR2_X1    g27638(.A1(new_n27685_), .A2(new_n27682_), .Z(new_n27706_));
  NOR2_X1    g27639(.A1(new_n27693_), .A2(new_n27706_), .ZN(new_n27707_));
  INV_X1     g27640(.I(new_n27707_), .ZN(new_n27708_));
  OAI21_X1   g27641(.A1(new_n27690_), .A2(new_n27708_), .B(new_n27705_), .ZN(new_n27709_));
  OAI21_X1   g27642(.A1(new_n27670_), .A2(new_n27676_), .B(new_n27678_), .ZN(new_n27710_));
  INV_X1     g27643(.I(new_n27710_), .ZN(new_n27711_));
  INV_X1     g27644(.I(new_n27621_), .ZN(new_n27712_));
  NOR2_X1    g27645(.A1(new_n27712_), .A2(new_n27645_), .ZN(new_n27713_));
  NOR2_X1    g27646(.A1(new_n27713_), .A2(new_n27646_), .ZN(new_n27714_));
  INV_X1     g27647(.I(new_n11229_), .ZN(new_n27715_));
  NOR2_X1    g27648(.A1(new_n24835_), .A2(new_n11228_), .ZN(new_n27716_));
  OAI22_X1   g27649(.A1(new_n27716_), .A2(\a[20] ), .B1(new_n27715_), .B2(new_n24835_), .ZN(new_n27717_));
  INV_X1     g27650(.I(new_n12918_), .ZN(new_n27718_));
  NAND3_X1   g27651(.A1(new_n27718_), .A2(new_n1742_), .A3(new_n11834_), .ZN(new_n27719_));
  NAND4_X1   g27652(.A1(new_n2375_), .A2(new_n451_), .A3(new_n1892_), .A4(new_n985_), .ZN(new_n27720_));
  NAND3_X1   g27653(.A1(new_n11578_), .A2(new_n27720_), .A3(new_n661_), .ZN(new_n27721_));
  INV_X1     g27654(.I(new_n1079_), .ZN(new_n27722_));
  NOR4_X1    g27655(.A1(new_n950_), .A2(new_n510_), .A3(new_n634_), .A4(new_n1160_), .ZN(new_n27723_));
  NAND4_X1   g27656(.A1(new_n27723_), .A2(new_n473_), .A3(new_n959_), .A4(new_n27722_), .ZN(new_n27724_));
  NOR4_X1    g27657(.A1(new_n27724_), .A2(new_n2426_), .A3(new_n27719_), .A4(new_n27721_), .ZN(new_n27725_));
  NAND2_X1   g27658(.A1(new_n27725_), .A2(new_n3491_), .ZN(new_n27726_));
  NAND2_X1   g27659(.A1(new_n27536_), .A2(new_n27726_), .ZN(new_n27727_));
  INV_X1     g27660(.I(new_n27727_), .ZN(new_n27728_));
  NOR2_X1    g27661(.A1(new_n27536_), .A2(new_n27726_), .ZN(new_n27729_));
  NOR2_X1    g27662(.A1(new_n27728_), .A2(new_n27729_), .ZN(new_n27730_));
  INV_X1     g27663(.I(new_n27730_), .ZN(new_n27731_));
  XNOR2_X1   g27664(.A1(new_n27536_), .A2(new_n27726_), .ZN(new_n27732_));
  NOR2_X1    g27665(.A1(new_n27717_), .A2(new_n27732_), .ZN(new_n27733_));
  AOI21_X1   g27666(.A1(new_n27717_), .A2(new_n27731_), .B(new_n27733_), .ZN(new_n27734_));
  NAND2_X1   g27667(.A1(new_n27639_), .A2(new_n27636_), .ZN(new_n27735_));
  NAND2_X1   g27668(.A1(new_n27735_), .A2(new_n27637_), .ZN(new_n27736_));
  NAND2_X1   g27669(.A1(new_n21157_), .A2(new_n3332_), .ZN(new_n27737_));
  OAI21_X1   g27670(.A1(new_n19475_), .A2(new_n2771_), .B(new_n2764_), .ZN(new_n27738_));
  AOI21_X1   g27671(.A1(new_n19484_), .A2(new_n3189_), .B(new_n27738_), .ZN(new_n27739_));
  AND3_X2    g27672(.A1(new_n21155_), .A2(new_n27737_), .A3(new_n27739_), .Z(new_n27740_));
  XNOR2_X1   g27673(.A1(new_n27740_), .A2(new_n27736_), .ZN(new_n27741_));
  NOR2_X1    g27674(.A1(new_n27741_), .A2(new_n27734_), .ZN(new_n27742_));
  INV_X1     g27675(.I(new_n27734_), .ZN(new_n27743_));
  NOR2_X1    g27676(.A1(new_n27740_), .A2(new_n27736_), .ZN(new_n27744_));
  INV_X1     g27677(.I(new_n27744_), .ZN(new_n27745_));
  NAND2_X1   g27678(.A1(new_n27740_), .A2(new_n27736_), .ZN(new_n27746_));
  AOI21_X1   g27679(.A1(new_n27745_), .A2(new_n27746_), .B(new_n27743_), .ZN(new_n27747_));
  NOR2_X1    g27680(.A1(new_n27742_), .A2(new_n27747_), .ZN(new_n27748_));
  OAI22_X1   g27681(.A1(new_n19512_), .A2(new_n2747_), .B1(new_n21960_), .B2(new_n2742_), .ZN(new_n27749_));
  NAND2_X1   g27682(.A1(new_n22048_), .A2(new_n2750_), .ZN(new_n27750_));
  AOI21_X1   g27683(.A1(new_n27750_), .A2(new_n27749_), .B(new_n2737_), .ZN(new_n27751_));
  NAND2_X1   g27684(.A1(new_n22175_), .A2(new_n27751_), .ZN(new_n27752_));
  XOR2_X1    g27685(.A1(new_n27752_), .A2(\a[29] ), .Z(new_n27753_));
  AND2_X2    g27686(.A1(new_n27753_), .A2(new_n27748_), .Z(new_n27754_));
  NOR2_X1    g27687(.A1(new_n27753_), .A2(new_n27748_), .ZN(new_n27755_));
  NOR2_X1    g27688(.A1(new_n27754_), .A2(new_n27755_), .ZN(new_n27756_));
  NOR2_X1    g27689(.A1(new_n27714_), .A2(new_n27756_), .ZN(new_n27757_));
  INV_X1     g27690(.I(new_n27714_), .ZN(new_n27758_));
  XNOR2_X1   g27691(.A1(new_n27753_), .A2(new_n27748_), .ZN(new_n27759_));
  NOR2_X1    g27692(.A1(new_n27758_), .A2(new_n27759_), .ZN(new_n27760_));
  NOR2_X1    g27693(.A1(new_n27760_), .A2(new_n27757_), .ZN(new_n27761_));
  INV_X1     g27694(.I(new_n27761_), .ZN(new_n27762_));
  NOR2_X1    g27695(.A1(new_n27661_), .A2(new_n27648_), .ZN(new_n27763_));
  NOR2_X1    g27696(.A1(new_n27763_), .A2(new_n27662_), .ZN(new_n27764_));
  OAI22_X1   g27697(.A1(new_n22115_), .A2(new_n3268_), .B1(new_n3322_), .B2(new_n22149_), .ZN(new_n27765_));
  NAND2_X1   g27698(.A1(new_n23957_), .A2(new_n3317_), .ZN(new_n27766_));
  AOI21_X1   g27699(.A1(new_n27765_), .A2(new_n27766_), .B(new_n3260_), .ZN(new_n27767_));
  NAND2_X1   g27700(.A1(new_n23955_), .A2(new_n27767_), .ZN(new_n27768_));
  XOR2_X1    g27701(.A1(new_n27768_), .A2(\a[26] ), .Z(new_n27769_));
  INV_X1     g27702(.I(new_n27769_), .ZN(new_n27770_));
  XOR2_X1    g27703(.A1(new_n27764_), .A2(new_n27770_), .Z(new_n27771_));
  INV_X1     g27704(.I(new_n27771_), .ZN(new_n27772_));
  NOR3_X1    g27705(.A1(new_n27763_), .A2(new_n27662_), .A3(new_n27770_), .ZN(new_n27773_));
  NOR2_X1    g27706(.A1(new_n27764_), .A2(new_n27769_), .ZN(new_n27774_));
  NOR2_X1    g27707(.A1(new_n27774_), .A2(new_n27773_), .ZN(new_n27775_));
  NOR2_X1    g27708(.A1(new_n27775_), .A2(new_n27762_), .ZN(new_n27776_));
  AOI21_X1   g27709(.A1(new_n27772_), .A2(new_n27762_), .B(new_n27776_), .ZN(new_n27777_));
  INV_X1     g27710(.I(new_n27664_), .ZN(new_n27778_));
  NOR2_X1    g27711(.A1(new_n27778_), .A2(new_n27669_), .ZN(new_n27779_));
  OAI22_X1   g27712(.A1(new_n24376_), .A2(new_n3306_), .B1(new_n3310_), .B2(new_n24167_), .ZN(new_n27780_));
  NAND2_X1   g27713(.A1(new_n24620_), .A2(new_n3312_), .ZN(new_n27781_));
  AOI21_X1   g27714(.A1(new_n27781_), .A2(new_n27780_), .B(new_n3302_), .ZN(new_n27782_));
  NAND2_X1   g27715(.A1(new_n24618_), .A2(new_n27782_), .ZN(new_n27783_));
  XOR2_X1    g27716(.A1(new_n27783_), .A2(\a[23] ), .Z(new_n27784_));
  INV_X1     g27717(.I(new_n27784_), .ZN(new_n27785_));
  NOR2_X1    g27718(.A1(new_n27779_), .A2(new_n27785_), .ZN(new_n27786_));
  INV_X1     g27719(.I(new_n27786_), .ZN(new_n27787_));
  NAND2_X1   g27720(.A1(new_n27779_), .A2(new_n27785_), .ZN(new_n27788_));
  AOI21_X1   g27721(.A1(new_n27787_), .A2(new_n27788_), .B(new_n27777_), .ZN(new_n27789_));
  INV_X1     g27722(.I(new_n27777_), .ZN(new_n27790_));
  XOR2_X1    g27723(.A1(new_n27779_), .A2(new_n27784_), .Z(new_n27791_));
  NOR2_X1    g27724(.A1(new_n27791_), .A2(new_n27790_), .ZN(new_n27792_));
  NOR2_X1    g27725(.A1(new_n27792_), .A2(new_n27789_), .ZN(new_n27793_));
  XOR2_X1    g27726(.A1(new_n27793_), .A2(new_n27711_), .Z(new_n27794_));
  NOR3_X1    g27727(.A1(new_n27615_), .A2(new_n27614_), .A3(new_n27616_), .ZN(new_n27795_));
  AOI21_X1   g27728(.A1(new_n27604_), .A2(new_n27611_), .B(new_n27612_), .ZN(new_n27796_));
  NOR2_X1    g27729(.A1(new_n27796_), .A2(new_n27795_), .ZN(new_n27797_));
  NOR4_X1    g27730(.A1(new_n27514_), .A2(new_n27519_), .A3(new_n27702_), .A4(new_n27797_), .ZN(new_n27798_));
  NAND2_X1   g27731(.A1(new_n27798_), .A2(new_n27794_), .ZN(new_n27799_));
  INV_X1     g27732(.I(new_n27794_), .ZN(new_n27800_));
  NOR4_X1    g27733(.A1(new_n23967_), .A2(new_n23962_), .A3(new_n24181_), .A4(new_n24400_), .ZN(new_n27801_));
  NAND4_X1   g27734(.A1(new_n27801_), .A2(new_n24626_), .A3(new_n24844_), .A4(new_n25233_), .ZN(new_n27802_));
  INV_X1     g27735(.I(new_n25240_), .ZN(new_n27803_));
  NOR4_X1    g27736(.A1(new_n27802_), .A2(new_n27803_), .A3(new_n25445_), .A4(new_n25680_), .ZN(new_n27804_));
  NAND4_X1   g27737(.A1(new_n27804_), .A2(new_n25897_), .A3(new_n26102_), .A4(new_n26262_), .ZN(new_n27805_));
  INV_X1     g27738(.I(new_n26441_), .ZN(new_n27806_));
  NOR4_X1    g27739(.A1(new_n27805_), .A2(new_n27806_), .A3(new_n26593_), .A4(new_n26708_), .ZN(new_n27807_));
  NAND4_X1   g27740(.A1(new_n27807_), .A2(new_n26832_), .A3(new_n26943_), .A4(new_n27188_), .ZN(new_n27808_));
  INV_X1     g27741(.I(new_n27193_), .ZN(new_n27809_));
  NOR4_X1    g27742(.A1(new_n27808_), .A2(new_n27809_), .A3(new_n27309_), .A4(new_n27517_), .ZN(new_n27810_));
  OAI21_X1   g27743(.A1(new_n27700_), .A2(new_n27699_), .B(new_n27682_), .ZN(new_n27811_));
  NAND3_X1   g27744(.A1(new_n27696_), .A2(new_n27683_), .A3(new_n27697_), .ZN(new_n27812_));
  NAND2_X1   g27745(.A1(new_n27811_), .A2(new_n27812_), .ZN(new_n27813_));
  NAND4_X1   g27746(.A1(new_n27810_), .A2(new_n27518_), .A3(new_n27618_), .A4(new_n27813_), .ZN(new_n27814_));
  NAND2_X1   g27747(.A1(new_n27814_), .A2(new_n27800_), .ZN(new_n27815_));
  NAND2_X1   g27748(.A1(new_n27815_), .A2(new_n27799_), .ZN(new_n27816_));
  XOR2_X1    g27749(.A1(new_n27816_), .A2(new_n27709_), .Z(\result[25] ));
  XOR2_X1    g27750(.A1(new_n27709_), .A2(new_n27794_), .Z(new_n27818_));
  NAND4_X1   g27751(.A1(new_n27520_), .A2(new_n27618_), .A3(new_n27813_), .A4(new_n27818_), .ZN(new_n27819_));
  INV_X1     g27752(.I(new_n27754_), .ZN(new_n27820_));
  AOI21_X1   g27753(.A1(new_n27758_), .A2(new_n27820_), .B(new_n27755_), .ZN(new_n27821_));
  NOR2_X1    g27754(.A1(new_n27717_), .A2(new_n27728_), .ZN(new_n27822_));
  NOR2_X1    g27755(.A1(new_n27822_), .A2(new_n27729_), .ZN(new_n27823_));
  NOR2_X1    g27756(.A1(new_n19512_), .A2(new_n2772_), .ZN(new_n27824_));
  NOR2_X1    g27757(.A1(new_n19522_), .A2(new_n2767_), .ZN(new_n27825_));
  NOR2_X1    g27758(.A1(new_n17775_), .A2(new_n2771_), .ZN(new_n27826_));
  NOR4_X1    g27759(.A1(new_n27824_), .A2(new_n2764_), .A3(new_n27825_), .A4(new_n27826_), .ZN(new_n27827_));
  INV_X1     g27760(.I(new_n8323_), .ZN(new_n27828_));
  INV_X1     g27761(.I(new_n12855_), .ZN(new_n27829_));
  NAND3_X1   g27762(.A1(new_n773_), .A2(new_n551_), .A3(new_n669_), .ZN(new_n27830_));
  NOR4_X1    g27763(.A1(new_n27830_), .A2(new_n1247_), .A3(new_n1167_), .A4(new_n298_), .ZN(new_n27831_));
  INV_X1     g27764(.I(new_n3671_), .ZN(new_n27832_));
  NOR4_X1    g27765(.A1(new_n11045_), .A2(new_n27832_), .A3(new_n226_), .A4(new_n644_), .ZN(new_n27833_));
  NAND4_X1   g27766(.A1(new_n27833_), .A2(new_n1534_), .A3(new_n2337_), .A4(new_n27831_), .ZN(new_n27834_));
  NAND2_X1   g27767(.A1(new_n2264_), .A2(new_n11723_), .ZN(new_n27835_));
  NOR4_X1    g27768(.A1(new_n27835_), .A2(new_n2941_), .A3(new_n27829_), .A4(new_n27834_), .ZN(new_n27836_));
  NAND2_X1   g27769(.A1(new_n27828_), .A2(new_n27836_), .ZN(new_n27837_));
  NAND3_X1   g27770(.A1(new_n25926_), .A2(new_n27827_), .A3(new_n27837_), .ZN(new_n27838_));
  NAND2_X1   g27771(.A1(new_n25926_), .A2(new_n27827_), .ZN(new_n27839_));
  INV_X1     g27772(.I(new_n27837_), .ZN(new_n27840_));
  NAND2_X1   g27773(.A1(new_n27839_), .A2(new_n27840_), .ZN(new_n27841_));
  AOI21_X1   g27774(.A1(new_n27841_), .A2(new_n27838_), .B(new_n27823_), .ZN(new_n27842_));
  XOR2_X1    g27775(.A1(new_n27839_), .A2(new_n27837_), .Z(new_n27843_));
  NOR3_X1    g27776(.A1(new_n27843_), .A2(new_n27729_), .A3(new_n27822_), .ZN(new_n27844_));
  NOR2_X1    g27777(.A1(new_n27844_), .A2(new_n27842_), .ZN(new_n27845_));
  INV_X1     g27778(.I(new_n27845_), .ZN(new_n27846_));
  OAI21_X1   g27779(.A1(new_n27743_), .A2(new_n27744_), .B(new_n27746_), .ZN(new_n27847_));
  AOI22_X1   g27780(.A1(new_n22048_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n21953_), .ZN(new_n27848_));
  NOR2_X1    g27781(.A1(new_n22115_), .A2(new_n3175_), .ZN(new_n27849_));
  OAI21_X1   g27782(.A1(new_n27849_), .A2(new_n27848_), .B(new_n2736_), .ZN(new_n27850_));
  NOR3_X1    g27783(.A1(new_n23675_), .A2(\a[29] ), .A3(new_n27850_), .ZN(new_n27851_));
  NOR2_X1    g27784(.A1(new_n23675_), .A2(new_n27850_), .ZN(new_n27852_));
  NOR2_X1    g27785(.A1(new_n27852_), .A2(new_n74_), .ZN(new_n27853_));
  NOR2_X1    g27786(.A1(new_n27853_), .A2(new_n27851_), .ZN(new_n27854_));
  XOR2_X1    g27787(.A1(new_n27854_), .A2(new_n27847_), .Z(new_n27855_));
  INV_X1     g27788(.I(new_n27855_), .ZN(new_n27856_));
  INV_X1     g27789(.I(new_n27854_), .ZN(new_n27857_));
  NOR2_X1    g27790(.A1(new_n27857_), .A2(new_n27847_), .ZN(new_n27858_));
  INV_X1     g27791(.I(new_n27858_), .ZN(new_n27859_));
  NAND2_X1   g27792(.A1(new_n27857_), .A2(new_n27847_), .ZN(new_n27860_));
  AOI21_X1   g27793(.A1(new_n27859_), .A2(new_n27860_), .B(new_n27846_), .ZN(new_n27861_));
  AOI21_X1   g27794(.A1(new_n27846_), .A2(new_n27856_), .B(new_n27861_), .ZN(new_n27862_));
  OAI22_X1   g27795(.A1(new_n23948_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n22149_), .ZN(new_n27863_));
  NAND2_X1   g27796(.A1(new_n24174_), .A2(new_n3317_), .ZN(new_n27864_));
  AOI21_X1   g27797(.A1(new_n27864_), .A2(new_n27863_), .B(new_n3260_), .ZN(new_n27865_));
  NAND2_X1   g27798(.A1(new_n24172_), .A2(new_n27865_), .ZN(new_n27866_));
  XOR2_X1    g27799(.A1(new_n27866_), .A2(\a[26] ), .Z(new_n27867_));
  INV_X1     g27800(.I(new_n27867_), .ZN(new_n27868_));
  NOR2_X1    g27801(.A1(new_n27862_), .A2(new_n27868_), .ZN(new_n27869_));
  INV_X1     g27802(.I(new_n27862_), .ZN(new_n27870_));
  NOR2_X1    g27803(.A1(new_n27870_), .A2(new_n27867_), .ZN(new_n27871_));
  NOR2_X1    g27804(.A1(new_n27871_), .A2(new_n27869_), .ZN(new_n27872_));
  NOR2_X1    g27805(.A1(new_n27872_), .A2(new_n27821_), .ZN(new_n27873_));
  INV_X1     g27806(.I(new_n27821_), .ZN(new_n27874_));
  XOR2_X1    g27807(.A1(new_n27862_), .A2(new_n27867_), .Z(new_n27875_));
  NOR2_X1    g27808(.A1(new_n27875_), .A2(new_n27874_), .ZN(new_n27876_));
  NOR2_X1    g27809(.A1(new_n27873_), .A2(new_n27876_), .ZN(new_n27877_));
  NOR2_X1    g27810(.A1(new_n27773_), .A2(new_n27761_), .ZN(new_n27878_));
  AOI22_X1   g27811(.A1(new_n24620_), .A2(new_n3782_), .B1(new_n5291_), .B2(new_n24386_), .ZN(new_n27879_));
  NOR2_X1    g27812(.A1(new_n24835_), .A2(new_n3780_), .ZN(new_n27880_));
  OAI21_X1   g27813(.A1(new_n27880_), .A2(new_n27879_), .B(new_n3301_), .ZN(new_n27881_));
  NOR2_X1    g27814(.A1(new_n26554_), .A2(new_n27881_), .ZN(new_n27882_));
  XOR2_X1    g27815(.A1(new_n27882_), .A2(new_n84_), .Z(new_n27883_));
  INV_X1     g27816(.I(new_n27883_), .ZN(new_n27884_));
  NOR3_X1    g27817(.A1(new_n27884_), .A2(new_n27774_), .A3(new_n27878_), .ZN(new_n27885_));
  NOR2_X1    g27818(.A1(new_n27878_), .A2(new_n27774_), .ZN(new_n27886_));
  NOR2_X1    g27819(.A1(new_n27883_), .A2(new_n27886_), .ZN(new_n27887_));
  NOR2_X1    g27820(.A1(new_n27885_), .A2(new_n27887_), .ZN(new_n27888_));
  NOR2_X1    g27821(.A1(new_n27888_), .A2(new_n27877_), .ZN(new_n27889_));
  INV_X1     g27822(.I(new_n27877_), .ZN(new_n27890_));
  XNOR2_X1   g27823(.A1(new_n27883_), .A2(new_n27886_), .ZN(new_n27891_));
  NOR2_X1    g27824(.A1(new_n27890_), .A2(new_n27891_), .ZN(new_n27892_));
  NOR2_X1    g27825(.A1(new_n27892_), .A2(new_n27889_), .ZN(new_n27893_));
  INV_X1     g27826(.I(new_n27893_), .ZN(new_n27894_));
  OAI21_X1   g27827(.A1(new_n27790_), .A2(new_n27786_), .B(new_n27788_), .ZN(new_n27895_));
  NOR2_X1    g27828(.A1(new_n27894_), .A2(new_n27895_), .ZN(new_n27896_));
  INV_X1     g27829(.I(new_n27896_), .ZN(new_n27897_));
  NAND2_X1   g27830(.A1(new_n27894_), .A2(new_n27895_), .ZN(new_n27898_));
  AND2_X2    g27831(.A1(new_n27897_), .A2(new_n27898_), .Z(new_n27899_));
  INV_X1     g27832(.I(new_n27899_), .ZN(new_n27900_));
  OAI21_X1   g27833(.A1(new_n27709_), .A2(new_n27793_), .B(new_n27710_), .ZN(new_n27901_));
  XOR2_X1    g27834(.A1(new_n27901_), .A2(new_n27900_), .Z(new_n27902_));
  XOR2_X1    g27835(.A1(new_n27819_), .A2(new_n27902_), .Z(\result[26] ));
  INV_X1     g27836(.I(new_n27869_), .ZN(new_n27904_));
  AOI21_X1   g27837(.A1(new_n27874_), .A2(new_n27904_), .B(new_n27871_), .ZN(new_n27905_));
  OAI21_X1   g27838(.A1(new_n27729_), .A2(new_n27822_), .B(new_n27841_), .ZN(new_n27906_));
  NAND2_X1   g27839(.A1(new_n27906_), .A2(new_n27838_), .ZN(new_n27907_));
  INV_X1     g27840(.I(new_n19722_), .ZN(new_n27908_));
  INV_X1     g27841(.I(new_n26147_), .ZN(new_n27909_));
  INV_X1     g27842(.I(new_n12998_), .ZN(new_n27910_));
  NOR4_X1    g27843(.A1(new_n1264_), .A2(new_n1247_), .A3(new_n1944_), .A4(new_n2551_), .ZN(new_n27911_));
  NAND2_X1   g27844(.A1(new_n295_), .A2(new_n302_), .ZN(new_n27912_));
  NOR4_X1    g27845(.A1(new_n2396_), .A2(new_n27912_), .A3(new_n804_), .A4(new_n544_), .ZN(new_n27913_));
  NAND4_X1   g27846(.A1(new_n1921_), .A2(new_n276_), .A3(new_n1066_), .A4(new_n423_), .ZN(new_n27914_));
  NAND4_X1   g27847(.A1(new_n27911_), .A2(new_n27913_), .A3(new_n27910_), .A4(new_n27914_), .ZN(new_n27915_));
  NOR4_X1    g27848(.A1(new_n27908_), .A2(new_n21906_), .A3(new_n27915_), .A4(new_n27909_), .ZN(new_n27916_));
  NAND2_X1   g27849(.A1(new_n27916_), .A2(new_n3415_), .ZN(new_n27917_));
  INV_X1     g27850(.I(new_n27917_), .ZN(new_n27918_));
  NOR2_X1    g27851(.A1(new_n27837_), .A2(new_n27918_), .ZN(new_n27919_));
  NOR2_X1    g27852(.A1(new_n27840_), .A2(new_n27917_), .ZN(new_n27920_));
  NOR2_X1    g27853(.A1(new_n27920_), .A2(new_n27919_), .ZN(new_n27921_));
  INV_X1     g27854(.I(new_n27921_), .ZN(new_n27922_));
  XOR2_X1    g27855(.A1(new_n27837_), .A2(new_n27917_), .Z(new_n27923_));
  NOR2_X1    g27856(.A1(new_n27907_), .A2(new_n27923_), .ZN(new_n27924_));
  AOI21_X1   g27857(.A1(new_n27907_), .A2(new_n27922_), .B(new_n27924_), .ZN(new_n27925_));
  OAI21_X1   g27858(.A1(new_n27845_), .A2(new_n27858_), .B(new_n27860_), .ZN(new_n27926_));
  NOR2_X1    g27859(.A1(new_n19512_), .A2(new_n2767_), .ZN(new_n27927_));
  NOR2_X1    g27860(.A1(new_n21960_), .A2(new_n2772_), .ZN(new_n27928_));
  OAI21_X1   g27861(.A1(new_n19522_), .A2(new_n2771_), .B(new_n2763_), .ZN(new_n27929_));
  NOR4_X1    g27862(.A1(new_n21963_), .A2(new_n27927_), .A3(new_n27928_), .A4(new_n27929_), .ZN(new_n27930_));
  XNOR2_X1   g27863(.A1(new_n27926_), .A2(new_n27930_), .ZN(new_n27931_));
  NOR2_X1    g27864(.A1(new_n27931_), .A2(new_n27925_), .ZN(new_n27932_));
  INV_X1     g27865(.I(new_n27925_), .ZN(new_n27933_));
  NOR2_X1    g27866(.A1(new_n27926_), .A2(new_n27930_), .ZN(new_n27934_));
  INV_X1     g27867(.I(new_n27934_), .ZN(new_n27935_));
  NAND2_X1   g27868(.A1(new_n27926_), .A2(new_n27930_), .ZN(new_n27936_));
  AOI21_X1   g27869(.A1(new_n27935_), .A2(new_n27936_), .B(new_n27933_), .ZN(new_n27937_));
  NOR2_X1    g27870(.A1(new_n27932_), .A2(new_n27937_), .ZN(new_n27938_));
  INV_X1     g27871(.I(new_n27938_), .ZN(new_n27939_));
  AOI22_X1   g27872(.A1(new_n24174_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n23957_), .ZN(new_n27940_));
  NOR2_X1    g27873(.A1(new_n24376_), .A2(new_n3318_), .ZN(new_n27941_));
  OAI21_X1   g27874(.A1(new_n27941_), .A2(new_n27940_), .B(new_n3259_), .ZN(new_n27942_));
  NOR2_X1    g27875(.A1(new_n24391_), .A2(new_n27942_), .ZN(new_n27943_));
  XOR2_X1    g27876(.A1(new_n27943_), .A2(new_n72_), .Z(new_n27944_));
  OAI22_X1   g27877(.A1(new_n22115_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n22051_), .ZN(new_n27945_));
  NAND2_X1   g27878(.A1(new_n22150_), .A2(new_n2750_), .ZN(new_n27946_));
  AOI21_X1   g27879(.A1(new_n27945_), .A2(new_n27946_), .B(new_n2737_), .ZN(new_n27947_));
  NAND2_X1   g27880(.A1(new_n22163_), .A2(new_n27947_), .ZN(new_n27948_));
  XOR2_X1    g27881(.A1(new_n27948_), .A2(\a[29] ), .Z(new_n27949_));
  XOR2_X1    g27882(.A1(new_n27944_), .A2(new_n27949_), .Z(new_n27950_));
  AND2_X2    g27883(.A1(new_n27944_), .A2(new_n27949_), .Z(new_n27951_));
  NOR2_X1    g27884(.A1(new_n27944_), .A2(new_n27949_), .ZN(new_n27952_));
  NOR2_X1    g27885(.A1(new_n27951_), .A2(new_n27952_), .ZN(new_n27953_));
  NOR2_X1    g27886(.A1(new_n27939_), .A2(new_n27953_), .ZN(new_n27954_));
  AOI21_X1   g27887(.A1(new_n27939_), .A2(new_n27950_), .B(new_n27954_), .ZN(new_n27955_));
  AOI22_X1   g27888(.A1(new_n24826_), .A2(new_n11469_), .B1(new_n5291_), .B2(new_n24620_), .ZN(new_n27956_));
  NOR3_X1    g27889(.A1(new_n25017_), .A2(new_n3302_), .A3(new_n27956_), .ZN(new_n27957_));
  XOR2_X1    g27890(.A1(new_n27957_), .A2(new_n84_), .Z(new_n27958_));
  NAND2_X1   g27891(.A1(new_n27955_), .A2(new_n27958_), .ZN(new_n27959_));
  NOR2_X1    g27892(.A1(new_n27955_), .A2(new_n27958_), .ZN(new_n27960_));
  INV_X1     g27893(.I(new_n27960_), .ZN(new_n27961_));
  AOI21_X1   g27894(.A1(new_n27961_), .A2(new_n27959_), .B(new_n27905_), .ZN(new_n27962_));
  INV_X1     g27895(.I(new_n27905_), .ZN(new_n27963_));
  XNOR2_X1   g27896(.A1(new_n27955_), .A2(new_n27958_), .ZN(new_n27964_));
  NOR2_X1    g27897(.A1(new_n27964_), .A2(new_n27963_), .ZN(new_n27965_));
  NOR2_X1    g27898(.A1(new_n27965_), .A2(new_n27962_), .ZN(new_n27966_));
  INV_X1     g27899(.I(new_n27885_), .ZN(new_n27967_));
  AOI21_X1   g27900(.A1(new_n27890_), .A2(new_n27967_), .B(new_n27887_), .ZN(new_n27968_));
  NOR2_X1    g27901(.A1(new_n27793_), .A2(new_n27710_), .ZN(new_n27969_));
  INV_X1     g27902(.I(new_n27969_), .ZN(new_n27970_));
  NOR2_X1    g27903(.A1(new_n27900_), .A2(new_n27969_), .ZN(new_n27971_));
  OAI21_X1   g27904(.A1(new_n27709_), .A2(new_n27970_), .B(new_n27971_), .ZN(new_n27972_));
  OAI21_X1   g27905(.A1(new_n27972_), .A2(new_n27896_), .B(new_n27968_), .ZN(new_n27973_));
  INV_X1     g27906(.I(new_n27973_), .ZN(new_n27974_));
  INV_X1     g27907(.I(new_n27968_), .ZN(new_n27975_));
  NAND2_X1   g27908(.A1(new_n26267_), .A2(new_n26105_), .ZN(new_n27976_));
  NAND3_X1   g27909(.A1(new_n27976_), .A2(new_n26278_), .A3(new_n26107_), .ZN(new_n27977_));
  NAND3_X1   g27910(.A1(new_n27977_), .A2(new_n26435_), .A3(new_n26702_), .ZN(new_n27978_));
  NAND3_X1   g27911(.A1(new_n27978_), .A2(new_n26704_), .A3(new_n27066_), .ZN(new_n27979_));
  NAND3_X1   g27912(.A1(new_n27979_), .A2(new_n26712_), .A3(new_n27052_), .ZN(new_n27980_));
  NAND3_X1   g27913(.A1(new_n27980_), .A2(new_n27074_), .A3(new_n27053_), .ZN(new_n27981_));
  NAND3_X1   g27914(.A1(new_n27981_), .A2(new_n27189_), .A3(new_n27410_), .ZN(new_n27982_));
  NAND3_X1   g27915(.A1(new_n27982_), .A2(new_n27412_), .A3(new_n27426_), .ZN(new_n27983_));
  NAND3_X1   g27916(.A1(new_n27983_), .A2(new_n27424_), .A3(new_n27687_), .ZN(new_n27984_));
  NAND3_X1   g27917(.A1(new_n27984_), .A2(new_n27689_), .A3(new_n27707_), .ZN(new_n27985_));
  NAND3_X1   g27918(.A1(new_n27985_), .A2(new_n27705_), .A3(new_n27969_), .ZN(new_n27986_));
  NAND4_X1   g27919(.A1(new_n27986_), .A2(new_n27897_), .A3(new_n27975_), .A4(new_n27971_), .ZN(new_n27987_));
  INV_X1     g27920(.I(new_n27987_), .ZN(new_n27988_));
  OAI21_X1   g27921(.A1(new_n27974_), .A2(new_n27988_), .B(new_n27966_), .ZN(new_n27989_));
  INV_X1     g27922(.I(new_n27966_), .ZN(new_n27990_));
  NAND3_X1   g27923(.A1(new_n27973_), .A2(new_n27990_), .A3(new_n27987_), .ZN(new_n27991_));
  NAND2_X1   g27924(.A1(new_n27989_), .A2(new_n27991_), .ZN(new_n27992_));
  NOR2_X1    g27925(.A1(new_n27819_), .A2(new_n27902_), .ZN(new_n27993_));
  XOR2_X1    g27926(.A1(new_n27993_), .A2(new_n27992_), .Z(\result[27] ));
  INV_X1     g27927(.I(new_n27689_), .ZN(new_n27995_));
  AOI21_X1   g27928(.A1(new_n27608_), .A2(new_n27687_), .B(new_n27995_), .ZN(new_n27996_));
  AOI21_X1   g27929(.A1(new_n27996_), .A2(new_n27707_), .B(new_n27704_), .ZN(new_n27997_));
  INV_X1     g27930(.I(new_n27971_), .ZN(new_n27998_));
  AOI21_X1   g27931(.A1(new_n27997_), .A2(new_n27969_), .B(new_n27998_), .ZN(new_n27999_));
  NOR2_X1    g27932(.A1(new_n27966_), .A2(new_n27975_), .ZN(new_n28000_));
  XOR2_X1    g27933(.A1(new_n27966_), .A2(new_n27975_), .Z(new_n28001_));
  NOR2_X1    g27934(.A1(new_n28001_), .A2(new_n27896_), .ZN(new_n28002_));
  AOI21_X1   g27935(.A1(new_n27999_), .A2(new_n28002_), .B(new_n28000_), .ZN(new_n28003_));
  NAND2_X1   g27936(.A1(new_n27959_), .A2(new_n27963_), .ZN(new_n28004_));
  NAND2_X1   g27937(.A1(new_n28004_), .A2(new_n27961_), .ZN(new_n28005_));
  INV_X1     g27938(.I(new_n27951_), .ZN(new_n28006_));
  AOI21_X1   g27939(.A1(new_n27938_), .A2(new_n28006_), .B(new_n27952_), .ZN(new_n28007_));
  INV_X1     g27940(.I(new_n28007_), .ZN(new_n28008_));
  INV_X1     g27941(.I(new_n27919_), .ZN(new_n28009_));
  OAI21_X1   g27942(.A1(new_n27840_), .A2(new_n27917_), .B(new_n27907_), .ZN(new_n28010_));
  INV_X1     g27943(.I(new_n22175_), .ZN(new_n28011_));
  INV_X1     g27944(.I(new_n11710_), .ZN(new_n28012_));
  NOR2_X1    g27945(.A1(new_n24835_), .A2(new_n11709_), .ZN(new_n28013_));
  OAI22_X1   g27946(.A1(new_n28013_), .A2(\a[23] ), .B1(new_n28012_), .B2(new_n24835_), .ZN(new_n28014_));
  INV_X1     g27947(.I(new_n2681_), .ZN(new_n28015_));
  NOR4_X1    g27948(.A1(new_n633_), .A2(new_n638_), .A3(new_n226_), .A4(new_n744_), .ZN(new_n28016_));
  NAND4_X1   g27949(.A1(new_n269_), .A2(new_n507_), .A3(new_n1068_), .A4(new_n1059_), .ZN(new_n28017_));
  NAND4_X1   g27950(.A1(new_n3684_), .A2(new_n1321_), .A3(new_n716_), .A4(new_n1699_), .ZN(new_n28018_));
  NOR3_X1    g27951(.A1(new_n28018_), .A2(new_n28016_), .A3(new_n28017_), .ZN(new_n28019_));
  NAND4_X1   g27952(.A1(new_n11042_), .A2(new_n28015_), .A3(new_n3161_), .A4(new_n28019_), .ZN(new_n28020_));
  NAND2_X1   g27953(.A1(new_n28020_), .A2(new_n27917_), .ZN(new_n28021_));
  INV_X1     g27954(.I(new_n28021_), .ZN(new_n28022_));
  NOR2_X1    g27955(.A1(new_n28020_), .A2(new_n27917_), .ZN(new_n28023_));
  NOR2_X1    g27956(.A1(new_n28022_), .A2(new_n28023_), .ZN(new_n28024_));
  INV_X1     g27957(.I(new_n28024_), .ZN(new_n28025_));
  XOR2_X1    g27958(.A1(new_n28020_), .A2(new_n27918_), .Z(new_n28026_));
  NOR2_X1    g27959(.A1(new_n28014_), .A2(new_n28026_), .ZN(new_n28027_));
  AOI21_X1   g27960(.A1(new_n28014_), .A2(new_n28025_), .B(new_n28027_), .ZN(new_n28028_));
  NOR2_X1    g27961(.A1(new_n22051_), .A2(new_n2772_), .ZN(new_n28029_));
  NOR2_X1    g27962(.A1(new_n19512_), .A2(new_n2771_), .ZN(new_n28030_));
  NOR2_X1    g27963(.A1(new_n21960_), .A2(new_n2767_), .ZN(new_n28031_));
  NOR4_X1    g27964(.A1(new_n28029_), .A2(new_n2764_), .A3(new_n28030_), .A4(new_n28031_), .ZN(new_n28032_));
  AOI21_X1   g27965(.A1(new_n28011_), .A2(new_n28032_), .B(new_n28028_), .ZN(new_n28033_));
  INV_X1     g27966(.I(new_n28033_), .ZN(new_n28034_));
  INV_X1     g27967(.I(new_n28028_), .ZN(new_n28035_));
  NAND2_X1   g27968(.A1(new_n28011_), .A2(new_n28032_), .ZN(new_n28036_));
  NOR2_X1    g27969(.A1(new_n28036_), .A2(new_n28035_), .ZN(new_n28037_));
  INV_X1     g27970(.I(new_n28037_), .ZN(new_n28038_));
  AOI22_X1   g27971(.A1(new_n28034_), .A2(new_n28038_), .B1(new_n28009_), .B2(new_n28010_), .ZN(new_n28039_));
  NAND2_X1   g27972(.A1(new_n28010_), .A2(new_n28009_), .ZN(new_n28040_));
  XOR2_X1    g27973(.A1(new_n28036_), .A2(new_n28028_), .Z(new_n28041_));
  NOR2_X1    g27974(.A1(new_n28040_), .A2(new_n28041_), .ZN(new_n28042_));
  NOR2_X1    g27975(.A1(new_n28042_), .A2(new_n28039_), .ZN(new_n28043_));
  OAI21_X1   g27976(.A1(new_n27925_), .A2(new_n27934_), .B(new_n27936_), .ZN(new_n28044_));
  OAI22_X1   g27977(.A1(new_n22115_), .A2(new_n2747_), .B1(new_n2742_), .B2(new_n22149_), .ZN(new_n28045_));
  NAND2_X1   g27978(.A1(new_n23957_), .A2(new_n2750_), .ZN(new_n28046_));
  AOI21_X1   g27979(.A1(new_n28045_), .A2(new_n28046_), .B(new_n2737_), .ZN(new_n28047_));
  NAND2_X1   g27980(.A1(new_n23955_), .A2(new_n28047_), .ZN(new_n28048_));
  XOR2_X1    g27981(.A1(new_n28048_), .A2(\a[29] ), .Z(new_n28049_));
  INV_X1     g27982(.I(new_n28049_), .ZN(new_n28050_));
  NOR2_X1    g27983(.A1(new_n28044_), .A2(new_n28050_), .ZN(new_n28051_));
  INV_X1     g27984(.I(new_n28051_), .ZN(new_n28052_));
  NAND2_X1   g27985(.A1(new_n28044_), .A2(new_n28050_), .ZN(new_n28053_));
  AOI21_X1   g27986(.A1(new_n28052_), .A2(new_n28053_), .B(new_n28043_), .ZN(new_n28054_));
  XOR2_X1    g27987(.A1(new_n28044_), .A2(new_n28049_), .Z(new_n28055_));
  NOR3_X1    g27988(.A1(new_n28055_), .A2(new_n28039_), .A3(new_n28042_), .ZN(new_n28056_));
  OAI22_X1   g27989(.A1(new_n24376_), .A2(new_n3322_), .B1(new_n3268_), .B2(new_n24167_), .ZN(new_n28057_));
  NAND2_X1   g27990(.A1(new_n24620_), .A2(new_n3317_), .ZN(new_n28058_));
  AOI21_X1   g27991(.A1(new_n28058_), .A2(new_n28057_), .B(new_n3260_), .ZN(new_n28059_));
  NAND2_X1   g27992(.A1(new_n24618_), .A2(new_n28059_), .ZN(new_n28060_));
  XOR2_X1    g27993(.A1(new_n28060_), .A2(\a[26] ), .Z(new_n28061_));
  INV_X1     g27994(.I(new_n28061_), .ZN(new_n28062_));
  NOR3_X1    g27995(.A1(new_n28056_), .A2(new_n28054_), .A3(new_n28062_), .ZN(new_n28063_));
  NOR2_X1    g27996(.A1(new_n28056_), .A2(new_n28054_), .ZN(new_n28064_));
  NOR2_X1    g27997(.A1(new_n28064_), .A2(new_n28061_), .ZN(new_n28065_));
  OAI21_X1   g27998(.A1(new_n28065_), .A2(new_n28063_), .B(new_n28008_), .ZN(new_n28066_));
  XOR2_X1    g27999(.A1(new_n28064_), .A2(new_n28062_), .Z(new_n28067_));
  OAI21_X1   g28000(.A1(new_n28067_), .A2(new_n28008_), .B(new_n28066_), .ZN(new_n28068_));
  XNOR2_X1   g28001(.A1(new_n28005_), .A2(new_n28068_), .ZN(new_n28069_));
  INV_X1     g28002(.I(new_n28069_), .ZN(new_n28070_));
  INV_X1     g28003(.I(new_n27902_), .ZN(new_n28071_));
  NAND4_X1   g28004(.A1(new_n27798_), .A2(new_n27818_), .A3(new_n27992_), .A4(new_n28071_), .ZN(new_n28072_));
  NOR2_X1    g28005(.A1(new_n28072_), .A2(new_n28070_), .ZN(new_n28073_));
  INV_X1     g28006(.I(new_n27818_), .ZN(new_n28074_));
  AOI21_X1   g28007(.A1(new_n27973_), .A2(new_n27987_), .B(new_n27990_), .ZN(new_n28075_));
  INV_X1     g28008(.I(new_n27991_), .ZN(new_n28076_));
  NOR2_X1    g28009(.A1(new_n28076_), .A2(new_n28075_), .ZN(new_n28077_));
  NOR4_X1    g28010(.A1(new_n27814_), .A2(new_n28074_), .A3(new_n27902_), .A4(new_n28077_), .ZN(new_n28078_));
  NOR2_X1    g28011(.A1(new_n28078_), .A2(new_n28069_), .ZN(new_n28079_));
  OAI21_X1   g28012(.A1(new_n28079_), .A2(new_n28073_), .B(new_n28003_), .ZN(new_n28080_));
  INV_X1     g28013(.I(new_n28000_), .ZN(new_n28081_));
  INV_X1     g28014(.I(new_n28002_), .ZN(new_n28082_));
  OAI21_X1   g28015(.A1(new_n27972_), .A2(new_n28082_), .B(new_n28081_), .ZN(new_n28083_));
  NOR2_X1    g28016(.A1(new_n27814_), .A2(new_n28074_), .ZN(new_n28084_));
  NAND4_X1   g28017(.A1(new_n28084_), .A2(new_n28071_), .A3(new_n27992_), .A4(new_n28069_), .ZN(new_n28085_));
  NAND2_X1   g28018(.A1(new_n28072_), .A2(new_n28070_), .ZN(new_n28086_));
  NAND3_X1   g28019(.A1(new_n28085_), .A2(new_n28086_), .A3(new_n28083_), .ZN(new_n28087_));
  NAND2_X1   g28020(.A1(new_n28080_), .A2(new_n28087_), .ZN(\result[28] ));
  XOR2_X1    g28021(.A1(new_n28083_), .A2(new_n28069_), .Z(new_n28089_));
  INV_X1     g28022(.I(new_n28089_), .ZN(new_n28090_));
  NOR4_X1    g28023(.A1(new_n27819_), .A2(new_n27902_), .A3(new_n28077_), .A4(new_n28090_), .ZN(new_n28091_));
  OAI21_X1   g28024(.A1(new_n28043_), .A2(new_n28051_), .B(new_n28053_), .ZN(new_n28092_));
  INV_X1     g28025(.I(new_n28092_), .ZN(new_n28093_));
  AOI21_X1   g28026(.A1(new_n28040_), .A2(new_n28034_), .B(new_n28037_), .ZN(new_n28094_));
  NOR2_X1    g28027(.A1(new_n28014_), .A2(new_n28022_), .ZN(new_n28095_));
  NOR2_X1    g28028(.A1(new_n28095_), .A2(new_n28023_), .ZN(new_n28096_));
  NAND2_X1   g28029(.A1(new_n22118_), .A2(new_n3332_), .ZN(new_n28097_));
  NAND2_X1   g28030(.A1(new_n22048_), .A2(new_n3189_), .ZN(new_n28098_));
  AOI21_X1   g28031(.A1(new_n21953_), .A2(new_n2770_), .B(new_n2764_), .ZN(new_n28099_));
  NAND4_X1   g28032(.A1(new_n23675_), .A2(new_n28097_), .A3(new_n28098_), .A4(new_n28099_), .ZN(new_n28100_));
  NAND2_X1   g28033(.A1(new_n2148_), .A2(new_n1380_), .ZN(new_n28101_));
  NAND2_X1   g28034(.A1(new_n688_), .A2(new_n653_), .ZN(new_n28102_));
  NOR4_X1    g28035(.A1(new_n945_), .A2(new_n217_), .A3(new_n330_), .A4(new_n610_), .ZN(new_n28103_));
  INV_X1     g28036(.I(new_n28103_), .ZN(new_n28104_));
  NAND2_X1   g28037(.A1(new_n11982_), .A2(new_n28104_), .ZN(new_n28105_));
  NAND4_X1   g28038(.A1(new_n4798_), .A2(new_n827_), .A3(new_n1700_), .A4(new_n1810_), .ZN(new_n28106_));
  NOR4_X1    g28039(.A1(new_n28106_), .A2(new_n28101_), .A3(new_n28102_), .A4(new_n28105_), .ZN(new_n28107_));
  NAND4_X1   g28040(.A1(new_n28107_), .A2(new_n12991_), .A3(new_n2662_), .A4(new_n2675_), .ZN(new_n28108_));
  NOR3_X1    g28041(.A1(new_n3165_), .A2(new_n28108_), .A3(new_n22076_), .ZN(new_n28109_));
  NOR2_X1    g28042(.A1(new_n28100_), .A2(new_n28109_), .ZN(new_n28110_));
  NAND2_X1   g28043(.A1(new_n28100_), .A2(new_n28109_), .ZN(new_n28111_));
  INV_X1     g28044(.I(new_n28111_), .ZN(new_n28112_));
  NOR2_X1    g28045(.A1(new_n28112_), .A2(new_n28110_), .ZN(new_n28113_));
  NOR2_X1    g28046(.A1(new_n28113_), .A2(new_n28096_), .ZN(new_n28114_));
  INV_X1     g28047(.I(new_n28109_), .ZN(new_n28115_));
  XOR2_X1    g28048(.A1(new_n28100_), .A2(new_n28115_), .Z(new_n28116_));
  INV_X1     g28049(.I(new_n28116_), .ZN(new_n28117_));
  AOI21_X1   g28050(.A1(new_n28096_), .A2(new_n28117_), .B(new_n28114_), .ZN(new_n28118_));
  OAI22_X1   g28051(.A1(new_n23948_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n22149_), .ZN(new_n28119_));
  NAND2_X1   g28052(.A1(new_n24174_), .A2(new_n2750_), .ZN(new_n28120_));
  AOI21_X1   g28053(.A1(new_n28120_), .A2(new_n28119_), .B(new_n2737_), .ZN(new_n28121_));
  NAND2_X1   g28054(.A1(new_n24172_), .A2(new_n28121_), .ZN(new_n28122_));
  XOR2_X1    g28055(.A1(new_n28122_), .A2(\a[29] ), .Z(new_n28123_));
  XNOR2_X1   g28056(.A1(new_n28118_), .A2(new_n28123_), .ZN(new_n28124_));
  AND2_X2    g28057(.A1(new_n28118_), .A2(new_n28123_), .Z(new_n28125_));
  NOR2_X1    g28058(.A1(new_n28118_), .A2(new_n28123_), .ZN(new_n28126_));
  OAI21_X1   g28059(.A1(new_n28125_), .A2(new_n28126_), .B(new_n28094_), .ZN(new_n28127_));
  OAI21_X1   g28060(.A1(new_n28094_), .A2(new_n28124_), .B(new_n28127_), .ZN(new_n28128_));
  AOI22_X1   g28061(.A1(new_n24620_), .A2(new_n3323_), .B1(new_n3267_), .B2(new_n24386_), .ZN(new_n28129_));
  NOR2_X1    g28062(.A1(new_n24835_), .A2(new_n3318_), .ZN(new_n28130_));
  OAI21_X1   g28063(.A1(new_n28130_), .A2(new_n28129_), .B(new_n3259_), .ZN(new_n28131_));
  NOR2_X1    g28064(.A1(new_n26554_), .A2(new_n28131_), .ZN(new_n28132_));
  XOR2_X1    g28065(.A1(new_n28132_), .A2(new_n72_), .Z(new_n28133_));
  NAND2_X1   g28066(.A1(new_n28128_), .A2(new_n28133_), .ZN(new_n28134_));
  NOR2_X1    g28067(.A1(new_n28128_), .A2(new_n28133_), .ZN(new_n28135_));
  INV_X1     g28068(.I(new_n28135_), .ZN(new_n28136_));
  AOI21_X1   g28069(.A1(new_n28136_), .A2(new_n28134_), .B(new_n28093_), .ZN(new_n28137_));
  XOR2_X1    g28070(.A1(new_n28128_), .A2(new_n28133_), .Z(new_n28138_));
  AOI21_X1   g28071(.A1(new_n28093_), .A2(new_n28138_), .B(new_n28137_), .ZN(new_n28139_));
  NOR2_X1    g28072(.A1(new_n28063_), .A2(new_n28007_), .ZN(new_n28140_));
  NOR2_X1    g28073(.A1(new_n28140_), .A2(new_n28065_), .ZN(new_n28141_));
  NAND2_X1   g28074(.A1(new_n28141_), .A2(new_n28139_), .ZN(new_n28142_));
  OR2_X2     g28075(.A1(new_n28141_), .A2(new_n28139_), .Z(new_n28143_));
  AND2_X2    g28076(.A1(new_n28143_), .A2(new_n28142_), .Z(new_n28144_));
  NAND3_X1   g28077(.A1(new_n28083_), .A2(new_n28005_), .A3(new_n28144_), .ZN(new_n28145_));
  INV_X1     g28078(.I(new_n28005_), .ZN(new_n28146_));
  INV_X1     g28079(.I(new_n28144_), .ZN(new_n28147_));
  OAI21_X1   g28080(.A1(new_n28003_), .A2(new_n28146_), .B(new_n28147_), .ZN(new_n28148_));
  NAND3_X1   g28081(.A1(new_n27986_), .A2(new_n27971_), .A3(new_n28002_), .ZN(new_n28149_));
  NAND3_X1   g28082(.A1(new_n28149_), .A2(new_n28081_), .A3(new_n28005_), .ZN(new_n28150_));
  NAND2_X1   g28083(.A1(new_n28083_), .A2(new_n28146_), .ZN(new_n28151_));
  NAND2_X1   g28084(.A1(new_n28151_), .A2(new_n28150_), .ZN(new_n28152_));
  NAND4_X1   g28085(.A1(new_n28152_), .A2(new_n28068_), .A3(new_n28148_), .A4(new_n28145_), .ZN(new_n28153_));
  NAND2_X1   g28086(.A1(new_n28148_), .A2(new_n28145_), .ZN(new_n28154_));
  NOR2_X1    g28087(.A1(new_n28083_), .A2(new_n28146_), .ZN(new_n28155_));
  AOI21_X1   g28088(.A1(new_n28149_), .A2(new_n28081_), .B(new_n28005_), .ZN(new_n28156_));
  OAI21_X1   g28089(.A1(new_n28155_), .A2(new_n28156_), .B(new_n28068_), .ZN(new_n28157_));
  NAND2_X1   g28090(.A1(new_n28154_), .A2(new_n28157_), .ZN(new_n28158_));
  NAND2_X1   g28091(.A1(new_n28158_), .A2(new_n28153_), .ZN(new_n28159_));
  XOR2_X1    g28092(.A1(new_n28091_), .A2(new_n28159_), .Z(\result[29] ));
  NAND2_X1   g28093(.A1(new_n28078_), .A2(new_n28089_), .ZN(new_n28161_));
  INV_X1     g28094(.I(new_n28159_), .ZN(new_n28162_));
  NOR2_X1    g28095(.A1(new_n28125_), .A2(new_n28094_), .ZN(new_n28163_));
  NOR2_X1    g28096(.A1(new_n28163_), .A2(new_n28126_), .ZN(new_n28164_));
  NOR2_X1    g28097(.A1(new_n28112_), .A2(new_n28096_), .ZN(new_n28165_));
  NOR2_X1    g28098(.A1(new_n28165_), .A2(new_n28110_), .ZN(new_n28166_));
  NAND4_X1   g28099(.A1(new_n3152_), .A2(new_n1444_), .A3(new_n2697_), .A4(new_n11030_), .ZN(new_n28167_));
  NOR4_X1    g28100(.A1(new_n28167_), .A2(new_n3141_), .A3(new_n2036_), .A4(new_n2672_), .ZN(new_n28168_));
  NAND2_X1   g28101(.A1(new_n22077_), .A2(new_n28168_), .ZN(new_n28169_));
  XOR2_X1    g28102(.A1(new_n28169_), .A2(new_n28109_), .Z(new_n28170_));
  NOR2_X1    g28103(.A1(new_n28166_), .A2(new_n28170_), .ZN(new_n28171_));
  XNOR2_X1   g28104(.A1(new_n28169_), .A2(new_n28109_), .ZN(new_n28172_));
  INV_X1     g28105(.I(new_n28172_), .ZN(new_n28173_));
  AOI21_X1   g28106(.A1(new_n28166_), .A2(new_n28173_), .B(new_n28171_), .ZN(new_n28174_));
  NOR2_X1    g28107(.A1(new_n22115_), .A2(new_n2767_), .ZN(new_n28175_));
  NOR2_X1    g28108(.A1(new_n22051_), .A2(new_n2771_), .ZN(new_n28176_));
  OAI21_X1   g28109(.A1(new_n22149_), .A2(new_n2772_), .B(new_n2763_), .ZN(new_n28177_));
  NOR4_X1    g28110(.A1(new_n22163_), .A2(new_n28175_), .A3(new_n28176_), .A4(new_n28177_), .ZN(new_n28178_));
  XOR2_X1    g28111(.A1(new_n28174_), .A2(new_n28178_), .Z(new_n28179_));
  NOR2_X1    g28112(.A1(new_n28164_), .A2(new_n28179_), .ZN(new_n28180_));
  XNOR2_X1   g28113(.A1(new_n28174_), .A2(new_n28178_), .ZN(new_n28181_));
  NOR3_X1    g28114(.A1(new_n28181_), .A2(new_n28126_), .A3(new_n28163_), .ZN(new_n28182_));
  NOR2_X1    g28115(.A1(new_n28182_), .A2(new_n28180_), .ZN(new_n28183_));
  AOI22_X1   g28116(.A1(new_n24826_), .A2(new_n22025_), .B1(new_n3267_), .B2(new_n24620_), .ZN(new_n28184_));
  OR3_X2     g28117(.A1(new_n25017_), .A2(new_n3260_), .A3(new_n28184_), .Z(new_n28185_));
  XOR2_X1    g28118(.A1(new_n28185_), .A2(\a[26] ), .Z(new_n28186_));
  AOI22_X1   g28119(.A1(new_n24174_), .A2(new_n3275_), .B1(new_n2746_), .B2(new_n23957_), .ZN(new_n28187_));
  NOR2_X1    g28120(.A1(new_n24376_), .A2(new_n3175_), .ZN(new_n28188_));
  OAI21_X1   g28121(.A1(new_n28188_), .A2(new_n28187_), .B(new_n2736_), .ZN(new_n28189_));
  NOR2_X1    g28122(.A1(new_n24391_), .A2(new_n28189_), .ZN(new_n28190_));
  XOR2_X1    g28123(.A1(new_n28190_), .A2(new_n74_), .Z(new_n28191_));
  XOR2_X1    g28124(.A1(new_n28186_), .A2(new_n28191_), .Z(new_n28192_));
  NOR2_X1    g28125(.A1(new_n28183_), .A2(new_n28192_), .ZN(new_n28193_));
  XNOR2_X1   g28126(.A1(new_n28186_), .A2(new_n28191_), .ZN(new_n28194_));
  INV_X1     g28127(.I(new_n28194_), .ZN(new_n28195_));
  AOI21_X1   g28128(.A1(new_n28183_), .A2(new_n28195_), .B(new_n28193_), .ZN(new_n28196_));
  AOI21_X1   g28129(.A1(new_n28092_), .A2(new_n28134_), .B(new_n28135_), .ZN(new_n28197_));
  INV_X1     g28130(.I(new_n28197_), .ZN(new_n28198_));
  NOR2_X1    g28131(.A1(new_n28005_), .A2(new_n28068_), .ZN(new_n28199_));
  INV_X1     g28132(.I(new_n28199_), .ZN(new_n28200_));
  NAND2_X1   g28133(.A1(new_n28083_), .A2(new_n28200_), .ZN(new_n28201_));
  NAND2_X1   g28134(.A1(new_n28005_), .A2(new_n28068_), .ZN(new_n28202_));
  NAND3_X1   g28135(.A1(new_n28202_), .A2(new_n28142_), .A3(new_n28143_), .ZN(new_n28203_));
  INV_X1     g28136(.I(new_n28203_), .ZN(new_n28204_));
  AOI21_X1   g28137(.A1(new_n28201_), .A2(new_n28204_), .B(new_n28198_), .ZN(new_n28205_));
  AOI21_X1   g28138(.A1(new_n28149_), .A2(new_n28081_), .B(new_n28199_), .ZN(new_n28206_));
  NOR3_X1    g28139(.A1(new_n28206_), .A2(new_n28197_), .A3(new_n28203_), .ZN(new_n28207_));
  OAI21_X1   g28140(.A1(new_n28205_), .A2(new_n28207_), .B(new_n28196_), .ZN(new_n28208_));
  INV_X1     g28141(.I(new_n28196_), .ZN(new_n28209_));
  OAI21_X1   g28142(.A1(new_n28206_), .A2(new_n28203_), .B(new_n28197_), .ZN(new_n28210_));
  NAND3_X1   g28143(.A1(new_n28201_), .A2(new_n28198_), .A3(new_n28204_), .ZN(new_n28211_));
  NAND3_X1   g28144(.A1(new_n28211_), .A2(new_n28209_), .A3(new_n28210_), .ZN(new_n28212_));
  NAND2_X1   g28145(.A1(new_n28208_), .A2(new_n28212_), .ZN(new_n28213_));
  OAI21_X1   g28146(.A1(new_n28161_), .A2(new_n28162_), .B(new_n28213_), .ZN(new_n28214_));
  NAND4_X1   g28147(.A1(new_n28091_), .A2(new_n28159_), .A3(new_n28208_), .A4(new_n28212_), .ZN(new_n28215_));
  NAND2_X1   g28148(.A1(new_n28214_), .A2(new_n28215_), .ZN(\result[30] ));
  NOR2_X1    g28149(.A1(new_n28164_), .A2(new_n28174_), .ZN(new_n28217_));
  XOR2_X1    g28150(.A1(new_n28217_), .A2(\a[29] ), .Z(new_n28218_));
  XOR2_X1    g28151(.A1(new_n28164_), .A2(new_n28174_), .Z(new_n28219_));
  NAND2_X1   g28152(.A1(new_n28219_), .A2(new_n28178_), .ZN(new_n28220_));
  XOR2_X1    g28153(.A1(new_n28218_), .A2(new_n28220_), .Z(new_n28221_));
  OAI22_X1   g28154(.A1(new_n24376_), .A2(new_n2742_), .B1(new_n2747_), .B2(new_n24167_), .ZN(new_n28222_));
  NAND2_X1   g28155(.A1(new_n24620_), .A2(new_n2750_), .ZN(new_n28223_));
  AOI21_X1   g28156(.A1(new_n28223_), .A2(new_n28222_), .B(new_n2737_), .ZN(new_n28224_));
  NAND2_X1   g28157(.A1(new_n24618_), .A2(new_n28224_), .ZN(new_n28225_));
  XOR2_X1    g28158(.A1(new_n28221_), .A2(new_n28225_), .Z(new_n28226_));
  NAND3_X1   g28159(.A1(new_n3166_), .A2(new_n1572_), .A3(new_n3133_), .ZN(new_n28227_));
  XOR2_X1    g28160(.A1(new_n28227_), .A2(\a[26] ), .Z(new_n28228_));
  NOR2_X1    g28161(.A1(new_n24835_), .A2(new_n22071_), .ZN(new_n28229_));
  XOR2_X1    g28162(.A1(new_n28229_), .A2(new_n28115_), .Z(new_n28230_));
  XOR2_X1    g28163(.A1(new_n28230_), .A2(new_n28228_), .Z(new_n28231_));
  NOR3_X1    g28164(.A1(new_n28182_), .A2(new_n28180_), .A3(new_n28186_), .ZN(new_n28232_));
  XOR2_X1    g28165(.A1(new_n28232_), .A2(new_n28231_), .Z(new_n28233_));
  INV_X1     g28166(.I(new_n28191_), .ZN(new_n28234_));
  INV_X1     g28167(.I(new_n28186_), .ZN(new_n28235_));
  NOR2_X1    g28168(.A1(new_n28183_), .A2(new_n28235_), .ZN(new_n28236_));
  NOR3_X1    g28169(.A1(new_n28236_), .A2(new_n28232_), .A3(new_n28234_), .ZN(new_n28237_));
  XNOR2_X1   g28170(.A1(new_n28233_), .A2(new_n28237_), .ZN(new_n28238_));
  NAND2_X1   g28171(.A1(new_n22118_), .A2(new_n2770_), .ZN(new_n28239_));
  NAND2_X1   g28172(.A1(new_n23957_), .A2(new_n3332_), .ZN(new_n28240_));
  AOI21_X1   g28173(.A1(new_n22150_), .A2(new_n3189_), .B(new_n2763_), .ZN(new_n28241_));
  NAND4_X1   g28174(.A1(new_n23955_), .A2(new_n28239_), .A3(new_n28240_), .A4(new_n28241_), .ZN(new_n28242_));
  XOR2_X1    g28175(.A1(new_n28166_), .A2(new_n28169_), .Z(new_n28243_));
  NAND2_X1   g28176(.A1(new_n28243_), .A2(new_n28115_), .ZN(new_n28244_));
  XNOR2_X1   g28177(.A1(new_n28244_), .A2(new_n28242_), .ZN(new_n28245_));
  NOR2_X1    g28178(.A1(new_n28166_), .A2(new_n28169_), .ZN(new_n28246_));
  XOR2_X1    g28179(.A1(new_n28245_), .A2(new_n28246_), .Z(new_n28247_));
  XNOR2_X1   g28180(.A1(new_n28238_), .A2(new_n28247_), .ZN(new_n28248_));
  INV_X1     g28181(.I(new_n28248_), .ZN(new_n28249_));
  XOR2_X1    g28182(.A1(new_n28238_), .A2(new_n28247_), .Z(new_n28250_));
  NOR2_X1    g28183(.A1(new_n28250_), .A2(new_n28226_), .ZN(new_n28251_));
  AOI21_X1   g28184(.A1(new_n28226_), .A2(new_n28249_), .B(new_n28251_), .ZN(new_n28252_));
  NAND4_X1   g28185(.A1(new_n28091_), .A2(new_n28159_), .A3(new_n28213_), .A4(new_n28252_), .ZN(new_n28253_));
  INV_X1     g28186(.I(new_n28252_), .ZN(new_n28254_));
  NAND4_X1   g28187(.A1(new_n28078_), .A2(new_n28089_), .A3(new_n28159_), .A4(new_n28213_), .ZN(new_n28255_));
  NAND2_X1   g28188(.A1(new_n28255_), .A2(new_n28254_), .ZN(new_n28256_));
  NAND2_X1   g28189(.A1(new_n28256_), .A2(new_n28253_), .ZN(\result[31] ));
endmodule


